-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
qtuLg3+71X/iuE1c2x6pSQ8k6OCp1l+HPkx82vjluHYvarCznUoWWjrqywiZA/fF8bwedZxFN6Xs
kYa5Z/CPohKyFyfNJDfcbmXI3I/I6ECZX5YnM83yf/MGM0y1yThFEY4iCa8JJ3x5BCgICGywWhyn
UJ79VJ+mq1aAnoFbSNb5yk9V/VuGXyzw84W6A/dj5twptqWqr1Y1az1h+hyzFB7GzFKCcDOwlst2
eo00FQYcag3504qRw5bAKJ3tAefhahUpgUm+fE1RGB/2OjFrEjDsowKS6pBDIBJJpDR7V3Cs3wO+
pLuCtkmuIlFBKYV4xmm3TbqOiVzq5cjJ+iJHRQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 10256)
`protect data_block
Nlyf6SxAYsYZNo90JniEl5laXayoh4S9TkjwYH1oBlOxSq6z2nOkKq3QQ0vn4/k7ImP4VfqPA2fm
WZS3p9PxW0Nv6/Xc3kuQ15XtO/pjBhmdS7/x5/y1ePj/NyKTsjiYauMnHNI9AD9fqBeMWAR4s+rw
rx1cW1iA6VO4DhIwp5fxRcT55LHqTc9yCe/bIHOs1QVL+Ypt52lhn7jk3+RUTClWJn5nYMuELkhI
jSwWcadER6/TRKeUn4iCfwuTSNdRmvd1uwan8OF4E/5KoQSwuqH9dcE2a4TUgsexEHPGzL4eQgW8
I2y4yntYaHsPDAjrYjWAsy48hhDekO7lWZ4jjiAwuDjid7yOiZ/eiNb6/ZurqxSXbBx8cEw+G8QE
MxfmQmjS6pWpvUGea/Kc0Ie1+VHDf733GgDqBPrKYov02kMGC+cD+rSdLhvPf4X3bfVNygGMC9uG
aFaQWtCdNcvB5cG9UWnYMhg/34YaRI9YvO9LCvgLNttCvNYt5D7Qy8RyVqljK6lEhrtk+5VY5ayo
nOo6/bx4jBffoRYbUboIlzm8kLgcH1ENg09yxPgUws39rbEP+fRQSHb95vgw1E6GzfPDreJvV3PP
YVDbKdzwoo25qagG9O2TNxBD3OJa1rEJ7uUnecTU2d1ltCrO2A1nH08z6kyqFDzXTXurL3SFeR1x
LQyK8TE3DDUXkpzsHJ/pTU3CrqUkWAGaWrucTzfUFqBRVHYx2YNJltXZNmtHCVwhSHRa/mzyoGxc
+EEhNwmepApc9QYdVohDJs74yT2v/rcULrUQuyI2RoWp4hKUyNqVwuKYfOS63uTy3xTVAq90AgGk
h1lhdImyjJaHXHVDYEjwPShMRqq27Jy/LNad063y+jE0IzrGOgMCpq7TIlo8uFPuDRm5+tQp5nJ4
cvVRgP5cGSm4cber6j7NhRi+eH9mhMJk6ewWQz4WL3dR0mWCfMlebCT8W6jmss2AE4vzVpSta894
A5X2F0zI5UqR50M16zzufeyUDL5BS/FWYZiyjK4MysBPgeXYB2MVlL5mvMbbDn0ctvM6KPWpeSdV
2wphDavxU7NdrhHVlyIG6r1yhxu2FsHRLhNMMDj8R9+tuQbXQYhA0DRcTbO+ukFBpHDm6JUPpEo9
HiFGjFRiS5gzbejB7e6yzFDQySs3kipK2MZ3Sym14js1Td2aoNuNIeH+0jW70acfL/umr2FynfGw
rwLcUkPfm0GSvHl+s7a0TOh6NGepUYnx1Q6ymdnyyrEO5KKbVd/VQe2D+9kZfN/cSaDd7R//LSx/
hVKieN9x+3mon6uACcjhEjz68soiTtXi3BO3Ekxj3S+YeVe8bKbSw49Iat6YhhbKCWBnu3OPx3hP
QmPCdOxfdW+0IbjeLOKrn691Xji3XjMYCJ0I2T+XPCtMQ3JObaZzWi4EH9uo5ROZ5eALb0QnpEyh
19eW07BCC5oS8GHsbFxp8V7g2s8+MOiEr5C3WHSMBSINq8gKXvalu7qsfMrqwj76Kw7eAteO5TkX
GGRXjn85RVj5WEiV2Xe/J4tZf2Papi1hY2cOsVk52UgSl3Rp/YgZVGBQc1eowBQi4mYI48R+wiNN
cq0TcELtEXokdOKfFwVozuSfSR7s6jisFML7Q93AJoWZN6SOGYs9fdDElKAlFXfs1vCFpyrO//5F
mkJkumq3AAIs5Zu+0UTC2tr0K7J4vuzWU2aLOPoclc+FKIMQVnLLMX7qbFo687V0f9sFHiAFaRLG
NBxgMhQFx0L7CPpvKfDcUnImYVDUoqF1DVTnYbnogNqWzx7Upurq6hjvmQeUNbrwU0fZ27ojqfyo
iaGupn5qaaBRfX145M1B2eXalgHvh5nsuik1he/xZkb+KOLLUTFzlX/CECphUzV6Q9IkN4/KiIky
Nxw/SiDFIspXmUYTMl8utPElqGg83etNw+WY5uGt75MsOcxBdu6GZYuOx1rBzjn9GNUl8oS6x3iV
Tp9QsT7Fpi3fvl/7wZxpGaAfjpNgbkoe/hZvgB72X/9qwgVUyZMDxXULzxYtMUiYIxZbDnMSivip
TwdrS0XEQ4AfLVpI+sL1DRZ+ZzLhyoSvt8wvpXVgE4ac3N4BUo8yFD2WeS1KIQcurJAWkSzC1g2M
1yLuKdzwaOHsNvr6191pQIpOUfa8fSmmoVOO52HiuAlwar6tRWxYiy+POlR0+Kv557CJzcmNp8pD
autuiQTiTvwwKPDHZp7GcoUx8GbiDqXnq6b+u3LZHGOas7dwd2KxTbrVe+Zl8KZhwgRLjL28Hfd+
3M04Vd3gRC1eeJEjNqA0gXLri4BngaBoDYYR2Thxr5UU26VxiqPYveJLw7DgO7KXUG5r+xOI3Hjf
CUC8wW6A9AAHCW6T1yz1Pf7w7BGAbV3oU1v/vTc3wRp+x8Byq1/WI2pA/96YZOe/I7fuG1+aSk3M
OXLcyV1v7UdrIhiVGKD5KjhGh3kPRG3iIPDj12aSaVmX2oOJ35Ztw240yyBzDj2sEObAG3d25taf
TDdmRLC2/fFPmvDxadOzUamqEW83vCIrZxdjsKDjOS6Aj7Sy3fazRoftxWny/QSzgkK5vgBXafFU
jaxGBsLvOx7eaDdeyRwPyOLO1+wcniC/58/8pWGVPjc+GOA9Sp4JAneC9k2DN6F65HAGK9i327nG
qXhyjVUjaRMtroUd3sYnYDhk0+5pyHgIO3epLW/MVqF8yWf8saENXwYxLH3JJiF+CycNA2cNi/6n
TeD/o8XxLpECdAQaHtOcXxJaXUQLej5g79cZv+FYn7hLyRFWyOp0nyFxgBLOsuevx5h/rJijX8/J
XOEuRZ3RsU8XKpA3JNd9fE55xF9VzIEqRnIKHzJ+BwZSG3/tlokn1WHWp2Fq/QsnYJaD+GpIyj1r
s5tKE1qReBt2lAvh3lWNRBcAG/Wd1gJ30325S1JoRMt9TP5rI7XT4zQEFCrXpRWpOdxCUFjx8+jm
IJbHamCqXpo+Q8EmyIr3cu3Goxy2wdnOK80tRCiPi/4cA8Um69gFL5SRoM2m5BQGlWP/URlbd/WK
2INyOLSyx8dBJIwtLHb/1KFKG1GZ5iZybYxSeebmjEt0OD17hdIbx1JNI2t3uwXbSJfEs+GanoPj
rRTfiqhrDHYNBsT2JjGLEvfSwvhwzZQpC9OHLzHiPUQ9GtqWn+sUKqp+r/a4prEbBEZQ44IkiQI6
x2p+Gy2sQQ+hxzrQw175Y2poSGz6iRu0UBazHcRO5VXHmV8/SYRg2BBmxbkBnpnvhyPQGIt5E5r1
eFemHP00tAQQIXqUHFP94J9CUJikTwbB/AsyUFtt9lEb2w7lWd553becTeHmLx7qQnh55cQVnRzI
il6riNR+nuGVZVrHbWHPQXm5M1wtXYekFj8bt+GN/RlnZNSttpoDQ0wlLOuNmTCk4Wqo1VKe4M/p
CfNUYonOPsHH0XgcnQ9/3SLAOYCaTBdpl63qi4Q9Xsn7Woec6+DxY0r+mgqdbA2e0TlxrMmBM7QH
uRYhmdlFjeyKMQVny6z8txCeMLGE4CCXUwVGYAX4CGdEoXdSty7FkLVmkkK1s7CRGCnafyeHie/n
YLwxeLRA5vGTi3Wf6iLfmFxUmediIi653oho2HtwRXwNrwvOrVuHSOXYGQRSj4e8VyPA5rqX50Cs
NYCXYq8atYssqtKXpqawzjTZTjDWVVgQydLcPQfnG2C0YEViCOyGcxTsucwI0K9J7U6Xll5suKXw
wYzI4HVapt8nHwiJ7+LGsM8R2BdcbxlplP/l2NCmEXYcGjFa92JLKXyw+aeaD+M4DD7XQNXWQ3yr
xj4eG4ihqFyWgILUjrp9wmpVpqGv3PIfeo37jom9SDTGYYDjPQXSR3WYvFxuim6DrB57Kt+P8c1K
X9JZ5YwBBkkNEtdfd06asSBjHqK4FKIjK+BsLOLuDJ4eDAOM9ii+2fCo58Nxe+rKyxYOoBNxITcJ
KwwTeqbIXXRBiXjr0FYC5FveLv6BhgKKfFrQVDaCMY1LCzKyov3connFJYDLNhjQ9i+C5T5+drHi
cFVpm0mrbz5a9V7wshPNXvR218/q9g2FERIPGwjA4ed7snDMeQFKkbzIFJTeunOgRO84Np06WpBg
eAWi5MzCtyojOEx/h7mFvyUrX3lHT1C/i6qRxfQpGhJTRJFiexFomIfPmRMS5mmk16lJ5uVHaSo5
Z8LVMXEbSUCJHVElcL3JhSSlaa1S3ywoBtDim0ZpHhCD0DcQe5JBqiUNn88esygcfeVCGxqlIxv5
O1kxnes6u4aG1vgTV/hpfn7Sd/5cV3iyMBMwSNp1uAWLBuKMw5gGaNAeVisFQ1MBJQVH6YgisZM7
UxEr04bZTFtqie8ITBLW6sIq5c34L1Dp846m5Lp9NcAC6ix8D5FdQasT/1sHrotD4VbjLRQDUbQv
fiKafEj58wgHgSDTCgyGNWb2/CArrDUNXoQiXVxWoiR6KFCUbkXKDOdkHEe6KmrSG1OOV45PbQfS
psBTExumFg7BSVb0VO/M6zWYm87HWG/C4Y5vfaxI89yUO/bKArjlPDDE85XMgFhwP33RTDLMs5fm
gDt6d4/V/FFieNyEs668gckNb/jktn8pjwdrci0B6jo+X8xak5Sgv8PMi304cz6mdQkU7LLJKOba
9oS9eHsdaagFGjQ3Qr/gD3V7ocHq3y+7V2FjAfecf+pUOzev7YfBoxwbnVtPpDvhNfCnTw0/on1e
6WCaEzCbuTOpFYez6F+3MGOpdPWCJK3GpAxoGa8A1TiUrSQbmiZT7AHoSD04Asxwpm2eeGSbeUeh
ReINYqZZskdcgOWQCwhlWqazHWjC+qpxnljRJhTNFVdLy6b4ugvs1UiAZawmqGULbmtyOEvwe5kR
v2dBm8KdIyCXPOiHebRArZQ3g4cWPzjbItdDQKJG948IULG8/lEguP9Kes99uMiqiOZ8MnoDTiHp
SDyja9B0X8vYejZMnBFNxT6h1Pts3dFiLBbSDO901zjEJn4SPXtQht+klciqAkKjEhXLc+lvt1wN
O1HY5xlow9IEqzGyhrGCXO1IveGEwuxWp/9r7faH/+52dUry5XNQbLqw39wqhoFkDqdpKYkS+q3p
6DJTVxj9shdXEecwSQl3HjXPePCgEnhJ48b60a5wA7ZO2HwxGS6KIbTnmkAVZoNYLP9oI5khxmo1
GyRJ5dHgIeO4z5UGC/E/TcuoyNo6bW7Xy7tGUX7eIjQsq2KxLwBnW5KVTO670iZt2o1w26DUeVTR
ULneklnqKQx0nQerTG/9rrNf907Le4Y27/HCtw9TkFBbBP/ybcxtIwyRE4IqEWxeuNycCwi3tYbW
B2NgtdjtneUw/g8BU71uQ45fwWhP4HnfMDxiE8Xzci9bH0uCEYS+eFcPOpxi95pRhgAn47B8wHxb
fUQH+37sa/vs3coIBez4VMCeK/5hOEBcAzqg+xN6p5aR6+tSGlQ81YOP5ndxy87UDB0sIpPIyfVK
VGYOqltfXMzWOXgDYc91ZWXV91WyuX0zS7nkgrsFjv+Am+ejPwWdRmz+bl+bWm/uevNxfnMLXnOO
YlOs9ofU0mdRdY/f6rrNaGjHUwYHAXArr7STvIDBUIZXPbFLLoNemPbFxZol+35TDhHxUqFqd6D8
mcrOoY3uHYuhs1Sp8VqaYytMUrB+6RG6apxApWbXQPo41Z2/zplsLFcfUeBwhpO5CHKitMGZbZUx
djkUpfJD1LTjB/+Vfd3/jplhXJq7Lbi+o+nCiFey6b7Q4E+WAe/TQTM8S065rmVwqIhsYrrx50zL
AJwCVx1Qq9K9xQUztDmNu263g6BhdntLRHR6UijVeOAEBXJGqIPeP9ejEAPVm0eqWTH7mGJEGn5c
W73IviSZH6Y/7K8iDIgErVJhfQCBBPhjG8o/i0PbSSWWqu1P4qbOrrm/tzymBOGGZxEQS1qk8+Vy
zmpn1FIl80P8eetx6AS8iTIcZQ1xTN8Jb52Xl2AMe9buH1FeLwIsGjyOouAdCnX3WpuTu1e5cNcG
AVsa4rbiZVwynp90k7SnMRb2+MfpxCuzHdgUiAIBXtAHUISaeJvBH6Si5p5bt5OUq2F/jqc1B9tv
Yo/jbpePuYlveiu6TRe4qCwiCzEtV08syHt8iAqnEnt0tKL6vrnm7TQDxDBTrugGgSHIRzFCscwK
9aooRxZCdpOHYhGNhtVpeGnL9CWKbqmO4sgA2UB0R/0UwuWUtFfxbetX8pundJnFCVvNu/YFyTxX
1tJm9B2WbarbwK22NZIHqO/5EahWjc2w25LMw8vsm15kTigSW/oCh4Z3rbNHFL6ko3U6R9snkUCk
9zPjxk/uXQtJ/sSXKdVXoXZOMdTftnaC4txFZXMnzKDzlklkr/ezYuLk1hJFleMEZ4Q/2eQSZeg8
YMRNOTyx88oohvNLPYaqhEcIBb5+WCcUmRjbKPFYmktqXtD6COAZH9kzih2LK+7pGuwLt6KCfJQj
Zbea/edtFCmcaaPVg6ZC5CCyRAf1pY+488NIDMWV0QW8bOl2dAMJaY4GgHUk7oQdBH7Dp4Td3tsW
g/zv4RKz0qiLHcqzsLwjVSk1/XKXd3tTsF275dWKACQaxjCJEgwi1VG1TxEVP+86H3jsGAI1O/xQ
hj2Jz9h1l7AlZnpWWY353Xo9S+ZHA5a69GZgUj4Rz8eqQ6ZF5tHxDCoRfxn8aIaoqZ6QJ2wg9ahY
YfKfr8LbTqRrPuUX/IBIBCCVh9DlKyonG5S5SUg/QgUVGE3tvkYX8jRpOUsH6vsrV2O+EGhoBjtv
h/eYE+14j6f5ceLqEzO+M2IHCZdkCq02bCjszX5GJRDn11sGikWi6U+VxoG6Dtjyl/fH4tbxsqBp
owqM7gN5j4E+lJKWoubFEWf1XgGpuffQs8VHYxOoBahcYbE7k6/l6+MMBSgsMVpLbjk3xtsJ7TkA
OcbayZ/S9RYanWNFZYfvycoeEJDowbgY5xYQnPehqvz81lcQdAOPuxfM4eGWVGZkEflRUr/CgrwX
/kKs3hDf8CCPupP4S83g2ULNbnOcUBeUPZ05T0QiFTBj03ymZXAv8zVw8VQ+cmvywwEcs4iTaMtU
lqbPURHjaf+qwcZDrJvwiUAtHBJ8/NlJ7MeMEQc9t+DbVpb2O+o5hiZ0hKOFULZKVPmeBH7AhTKq
91mgUo+G+SMZ822hOv5AvVSPUFM0LcyttTWTyb4+j7txpW81hxNW2bIwdaC4eKCjjZw+dphDYlAy
KxmxKT0y19oPACNk2tlOaVb5cU4/eNjTDRgSZVI0+pmhynLyIWMonAqueSm5UIK0XTCne+0CbOTp
q+ys8HX6q/y97/Kz4lHlWK9OtFwN5VdYP3CGITm0M7hizvvmokTXjPv9btnrbcssJmnC4QrYUxL7
i48AmHStjWNgISo8oG/5zBszwPLKCySNiu9ZOy3TCw94l/vuzIUzqrqu+7JxAbnPygkPgPFpxHQv
ugmEZDpM2ZPu7/udvzrU3xcHzjyDJR7kFzsRQxDklP1PNc1xyu1a7Ezu0ouqwcADHPRFtDka8vSw
K2VVGQaq9wev/A4RsxGpytG/jP7XoW0MTPVB1uEP6UCe7nGqiC2dZSQcLUxkdds6bY0Kp/+HKHbu
KAXPGfu9muSdFxdENKosgBz/zHG8A6Fv1iocU16dsfuZ9rfuo2RKuuhi7OP7A918IpKJcxpSnziP
S0N4dtZfXINwFb68Ut+ScevCHkm3y1oXm9J/50OWbXC8jbyFjsJ7vrUTXxTGWDrhKjEh/jQz2biQ
m/kDX8GexubPnTt2ol0mNWZigH95k4Dcw57JThke3N+ZCSOAM/mPRvSsSiljGFH228z/uKALxI8I
z3xHqg99t/C7BWntBBY36Og4v+1/RGQosglXm6Yh5dinkF58U1+9Wu3jAJsmbKBCBMqAkfAV4jhR
L0Ygpn6oftDEbThcQvtjJYwLXJTibY0VDkqjLGY1IyfbntUj6P7JobLOK4TmLoqZdgLg8gm2BlKD
qwogRG6p73njGxdOzR31UiJ9Sp+YOXc8WwRgww4tHpe1e7t/mCJKmebi6G8YJpVSRg7hO627DMU7
DdgfEEeytRkTsuTHw/2//4DwcT5nGl+irwGnmOI/wzADx6oBeILXOiPiG1CeM6fH/wJMDXnTsvJ8
uBgE2HueZHR0qUB5UZnu6jNEUhrn+Nu36t9+GyNxWfDmE2/oXAoTyLd7GVUoHgham+bqYiB/MkMS
qSckw7R6PMA3r3QyPXNRcIPA1lk/C12+brk0uKu7qJxvyvlXG2bEArqUx/IjCqcCS+Tcdnoxbuwk
3nGyctx4Brje++ArfofP5ANZ6WMaPtyj9jQVCYv34mAMwaheMCVik/wfcHSZIrDkVmfi7GT0V+Bq
25VjYLkDG9guali0Lx+dKbyed0jOimm+v5IuWt5FcHMX56i4hqa0zm624fnRNzJxCJXq6e2sOARK
k25pdaq+4G3JdqPdtl9XNALdcZ4GpvXlEYV0+jC8Sf6mVK83dK18RGIzZQL2cM9KVFaAYsIt/rr/
j3QlazUHQknAvv0Wrh/BjJgPgw7d0pUoC/yzLRLIxPNDtuF4b/ZlQvg/bLxbbxe4C+ap8xicOdg7
tDosYAPXkIq0nedGKu/mznUJgDlP5i87iy2X4FJGhZudIii1p27O+FPBe7e9MskmQgdfrlBMHbIA
aOuHJuJtGJmPT4WzYlvLP63dP08G2p0HAgYEWarwGvHkUzjYpfFYn44W2hGpyRVBLcyuBj/Ymwgf
Zkb1P32a10EkIABVd17rsA5yu0mPcMKfKlSZG+EkgyK/rVQuu0QK6kJoOPvEgJBlPB/jsfeaQXWq
c+1iPwNwf++hhFIuYG/1apn9FDRE69UUccI5dPBKNaplb6cy2vn98YDqXLhAeNtxUXy3utb5MAQk
1iXxzpB38uvrrTf+lNThfKu/QtfXttMZ/M7M0Ep5OIAjFNGCJcgo493P3sY7zknBR8zoqTzJztIq
lvPhch++xlvVSPXmqndvCvIhg7G/QXwohDXVOtFUOfEpU2mfRUStjbbKzq3NqrjR6mbD8fHReWC9
YP0H27HltOQNBBJ4myXnkBG8ToZz/PITyjmmHAHWAi03FzmY6FghGjWbWOIxHRs3PchKCipGRPxo
jgy3pDv9idc2Sv2PNpz46seCh3Zs0wJ0PjnC8sBeD723afEo9jd0zTrRRDkaviDYSfEnALQqUrkp
rc965Wg6qFfvmpUOz7L3UmjBMBMKI/vB+zM924UepUQM4GF0ijsqwOQGDgf4jLsxTFrIbBOOc7/p
y5wp3EF8XN2ZxH4Hw4GGlnmqZOshWrM6YhWzkv/WrGxt6CFvfnPsXxCeSL79AK8mnDj2ptNMrxDx
LpE0DHi/tUqcr5RuyAmnXG6RxgsmgUBdn+iS+qZsqMNBqZSZERjJ0v+FeVA8sig7/YQKuPt73X8D
GH1RpvfJBUCA7nhItgYZX+eux/EhT44eJv2q9helc2N2vC/iiKg+JTJ6w42yk0Yn8m51i2n40rzT
TgQWGiottKdH3h3tkFP+/Z3kBsQQxM/yvXhqagcgkbIeKCzfkz/XBoDtSQ9VWWaDIBeLXgo/ZTT1
QSHbNZ1wNUEfk4bQt1cE/rDfkA9e2ES8uaDWb4eKrxMrapaOkF2+x0lb59cOTJXblqKWJyadbV2u
pNrxFRoLayY6+z9eYz0SOCOmZfT1mtWNM/Sa/cd3zTTlGzgCC4jVhQZAt553CQOU6dMdzVpNejL9
F4a8BIq1DZ/zFfi6EbY/17mUKR7ky+Hw0eAdJ/wLymdn/KgSNNmmzkohowcZ71JhpjXhne4cB96R
AdVkKcWbXlWxbYryg9zcEjxay5yryPW25Um/5n+krftPDvPngaC0A9WQqJJp7y9BcFbAl+x+IDnl
mZli4WaWiLEHbdVIjj3LMC3YCH8BYTXJjNhDl7R+7JhgpFD9iGrevTdHu+Tj0UKsvpCJj+Fuiq+B
XM3P9NibKzB07BdlLtNgwbmrCEBksnEooyaSSoQRLVMwG0YVo7fMDW5d0MFuPYb1bhemKJYuT9f5
j3uHOZv1qaeGXDLxmhpgP6RASSMQSUNMHXxM7Zy0+7rv3G6m54YjYWKA6PlQ31m/QV8IxuJC4omt
5iVy9utb72KvsJFxhYHMkIM/IfcrsHJ7nmyy4BZ0K1sHS3uqvj6uiRaY9SWotyRFdE7PLKUqh2tE
TR2e+MDED3pjyCxxV4ktOcplL9KC8e5HgMTQo3v9GSAA51frpFo0kiTS3y7EBt7qMw9Vl0VvNwyG
eeW1L2MRxXAJWdNA2hXcuXTbMFlTl7DSxkHG9t4rmnPtUS/xMPC+tmCiroYTCWFM1K2McypTHk3R
LI2YnalASX0xuRgJ2VEx5zy1U7wktCLneIP4Hn+CmIlQsuEZ9Uzn1LkprBnJxze7lzVM0Vk7DRSZ
9FIbsEAJiax270uw9Q6C7sUxSkGGLQAyEReRsrTTOakEKWfBVR/UE2705Hr9raAMIYrDeLw5n3m3
lCTmv5faYmLrM7jihD4x+YywaEdLSa9v9dn5AXS8T5q+lM/tjj8WANDoLnVgGPoMBnUhF2KyH6AP
ibNektQ7TY0Yc4Ja6vURYV3CFJeMuskI4Qfcr+ZUx4uKxDAoXYUSNi3yXFavf0wP387YewfvbX+R
cIni9UYa+HKOM8if//C6O+vTw54thZkl49lKj54wE1z2ck7owtH5IzBO6b/40GDPAlfQR+KMyG8W
5vcwHF5wIPxt8KeCCEwdBFcCE54u1JqS5fTlK5Sli38ajEJn1WGr2D5tZaatQYXslqZ2ItEO+zCd
EXuYqdS23N9mIPzxuSYpyzYoGqjcazcvFfJ2u51JbKbAuPXvALImJGKUs38NEU+w87IzELGGDaCG
e8u5QrTGzs9PeQThYKl2STtXdbjdk5QVkIzhQZHN71sd2aGO1VuXLUXxWxlXZZnbo6bYaF9+VqHp
yZGIkBfGeaZS+Wq8RQyy9bDGrO0dteL5QH2ACT14y4nA3hu4anAXxjHYvQ4JMoGKNfazgvPIGAii
15V7Mdgd0gAB4BaUtTSYRd3lL/cf2Zydu/+Zjjw1Qs1oX/fIBB3+irIQB5Cpqy+7IRBYg0OzJmSt
k69UWcBBkSeloPsTZn3zp7UrAXzOo5cBEH4Ac5US3V1jog7L1BkBqP6TF80oMQ0nIzZeqXNjHkVb
RaNEgkIlUVW2Vwghwv1Il/2paTg7vAG/AmG32MNZZL5ucIgM4v3xVg9T1YVlm41ZNUaYT9MMet3A
vqy0m2Zjjc+aIg8/omqs1xoT5WPc/Kw1pGYx/AdqAKCPFdnU60EJpsE/SJgkWVT+tCN5E7wo6EdX
XSYVtgl9YYEFr3ahJACunqbbMlQKjJl4fvDUUizDxx4fjDbCOI7k0qJOaKj0Yk9dla0lIiigo74e
Gn4ksVZse5GK0tpOlxSaQXXg2mrJ2jE0xNGnM9JlTjUTgIql9umCir4eoX7oKjE8XE5ayRYLiUtq
PIKHVVuXz9ma+tOT80hv2BiLjimWQkJwMkeEUfyN4WL2uljHNgUqSf1DKfHAzC+iTLNkGXBt3Oc5
/TQa7cIk8iGk94mwMyGrU20RABDls64Ds32zxQzC4pHcvK8oczI49zv4INUTFhWtYc4tfuWsvr3c
p+U7IBMwjWOHzpt6iKVHchzWIw0EDE84E2N/ysMiJNdtf004k5iCX12othAAjo/JRrJH7i4NIiCx
rnB63EPA7cbAbamXg14aA3uOvybk4W4eX7RDrpjfThOsZbRsCgCiyhA0s/sMoJDp2MfX8RCl1Doj
UC9QEKbBT40ZrIa0OmcBC0nfp3K2Xkuoy1ILZ0DhGWwoSBOpY74mtAHKNUUIALti2zO4i+DY1nAh
lAmzuxUx1fESbEFlhglc2Foy2YFcZ0OtFo/uWW9wkbDlIlTUIH75gs6Bz1EdsThCtQzJLN11KMPQ
004Pp99n7FRwK6WHxFCq5h9mvRtsUvqoZvPB69GUHl6c75wPr6WFjYfISVrInLP1KTgjsB8VfmEw
vEMf/ShDmCc3dGsHLik5NLBIjPQ6dFYRzVPvXDyY0T0cTPff7xZHfjqJCxdbaR5T72KeITPiCAgn
b1ToAArddmnrflo7IE27DL5LiSDoB0ph3qh4WJDFkZqIhk5Y+Oejm67YFy7XXwvZnu4Ypnvw+8Bd
p8KS8Y+qgAlNfHsuS6VZxaGGT3kGFRSb8VfiDPEmD9x+SDyOOmEwrHutpL5g5BX9A94EoQAtjtMR
NxsURU4gKDU6P4OSu5t8hqHXdzw9MWSahmwAqiHnGVwpO6SdYcdQZbJWT4lnfAcWmA0S2pMGX/KT
Vvsajcq9ztPLK7QLBJQXNdegBS9h7nu1JpV3at5+t1Js35NI8h6RaeWiAQThGJTBSlrPiBPgKctU
3A0o5t74Jd6Hy+BLyVt9izbJ8C/JQGjmdrgoy1zb5ty4Du0NEjGJHwePjHF73JDyX3sYLyvqZF7I
PScDDychut/fsze6fYnh5VzjsyM0EzM8lXAS24P1QrUpucVFnnhpSux4TNmrVjl9T4PJq8/wugVa
BIOu9kZwCtWenjuWXRqmQTCkADb7seLX0RWPt5CsmZmERaBJ3Ol38Sm2UYnY81sKFKRNS87SMnQz
rmSGRtRY+UlLw6DVtWPh3SXBxseSWBmGWRCoSxjex8eLYP048oqs1BwwlHIyisDg1FQCg+/zaPtj
bSW7qKcawXXV+8xFdxgQ2lh/nVdvcI+mhFQ5bhkOE54UWnjYlVYsRcfjOKuvzA5TG6WIHFfuVCGv
ASD1zzcHOKZf6NtroNYTNNTQL91d7mz3fzPeId8lq5XR4/xfdCP4Ukx/lcikVEpuF25Cx+rkkXAc
pzY1Dl9ErtL9TOvd//D2+CKFKxZqsvlUtDJHV/XZ8iRyBSv5VrCsfLehuiVVCIJzJo2SF5RhZrnz
MzIHhQurxFixww7IBuOvxgbpAjxJ9Ckwn2QH1EYn2E2lvjjgdfhrpd/C5K6g4Y1Wm1cvtSGyjhdh
mOZEK5CatKpc0QFbx0vC48ln1uHJuoZGDX/pS4RcOGk1X86lMXcRPOumJda7xS2H0gG9o1knsS8u
VrNIMVukP5JHZ5r4oO0D+NlI8YFe5EPuQiG3ymJYcqCKVowYldjR9TuYl51iispPGkLtyqb+T6Sx
ZtaC0lo/rzROCF+G0w0IcdNwCYolxVkfo1T1QNVTL6fvYjKCy4kIDdBxPW5biI0hDMG9/DLOUmvy
/pTjKuX3nE/hlpOozaCWCIsxTmtXOlSOSbabAngoasdWzZTtsMa8OoK4LIgWUXO1HDOF0UY1PXMA
4NYz2mQlDEmatDFY0f79gA/U7iTU5i6q3CKBby9oJU2ogPl/2xcgfotv6PPekRfJ40HKN9wI6h2S
mYQv48p6dmEUVD+sEOOi0i4rpQmg/dMq5fMCSeodW7wxDBTYqMKZyFkgwys+BgrKxYYqi7EcZbn8
ZetdvZovUr+RSB4kPTtC4F3IqyPnB/9POvoVUYPFIWtPBtSLa9yR+WbK+ddabhAeOptHFY0Ka8NR
VFfZ4A3HgLxH8tSPThyyOCQsbyupZskkPmse+aYd/3wdDauZSkhaj9rVKLVFI+N9CF7ZjlU6pWGQ
PL049wr7NZ2DOgaAbUAjB+xwosTHd4p3YD6+cCecVogsBJXDSZoDEj3WkbO8z2jF9Q53x5I=
`protect end_protected
