-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
0N1YSJtnh3iYtJ0hu8LC1CcRMm/XGkX6mxKA8H5QhtPpx82ilgNxVzLdEY72bc3Q1UlfTEQPdZhZ
aQjEymepPNvXm/TI3EAMOAnyEtwofqWbATXtN+2//JAts2KpXSfxye76QxRXRBqS61Voipo9Fi9H
iMkSxmt/PFO9Vx1vQef0oJL0Zk2cCQIUfycqsPEOVg4xszaWrEUdc9JFrI6od47gBQiyGEIYQK5m
/ZXrkkkSqYtP6BfT9Wqdv6TJTQb3Y42QaP0CVqWkLNuo6VKgrM3FSEPA75S+HMUYs9lveUoT+GMC
dsI0k5N7aoysS19oc8INGSBv3tB/2I2JZpw6uQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5280)
`protect data_block
End9IzNLrgj9I16Hv1a8rPigCO27Wr7mp3z4kl7OlWpl9L15pa6KUJpXv6rWjfNmGwj13SsGKwbc
IquCk2pEp6UUpZecFQFyozOP/EfzbWSGg6BVpwZymCM7Qu+hJvkk7D+YkWwQWJjHUY/tVWzbVLPf
TiXQ9KU2UGYQDhuoK5Bmp33yqXVl6LXnavpuxKopaw9tqE7bgFM8ohPgr5YX2QRmQqtmUvudydlQ
1T98iot9DK+Er6P6Ic0zcEjBZL8TOquvfon/I/aKhkDJ1sz1dua49qF09524CpJnBQXosh+iQVeD
Rv7tf1Of+g1QINTQh0XFRRC+itfXyydy5JvdTRNLwXCe+1MXMehqkqPWknggLlC+ievgVI9Hk1oV
oFL5EczLMac3fVtSVLKrjWwEJqzfMAIv2v7Sea2KfKMUkbg1igUFwDhw19J+8IfMxw5ANFIMnXj7
Jpxb0DDCwkp7GWAYmt0A30r7zEhASdtp3XdbQZ7mJ0rBXU1KnDqvQ+QydpjGZqJ/WDpmT+OKSZ9v
VdbxcPqf/x886+6brOY6bAIHHfUHDAdf93yYs+bbtGWoO/J81mm0uXPiJmF00solQauALrZCSBGU
nsnx2zsA0zjiBZqQ79E8GE+1Ukwbgpp0pITzWbf39+BmTpdCTCixvDHAIQV+lMGSWmWPfoqklGCr
hezh2CblnozbVARnOtgiiiZX9PRcqz7lgIVxqSMcQL/frBKybdlkTSmStAHNHCaq+q5G5rT5GJIe
198DTDNfBEFLF7zBxYj44u6o/3GnkQpkBP+mdbsrWML4nqVJh/QVkmFIonE0D5Wf5lsPoNnWq4RZ
nrgSMaW8jnBe4njXtO54TR2X6F+odzuHWBeX+tuhPRePHVK0yEvBWzuIvhJsPY3I5X3yncIX/3Ah
n/Q8IXM7be3FCB+Q7aoBJ2d1BxUgGGzWk49zI7J3UXHqPxsYuNfjwTVxG3BFuzerZW+J0zFv1XRS
h38ZHm1eLzIF+r1T2QTbdGeeR6jSFRae1a24+EdY6pPBg5N7Jf5RO/CpV5LPA/Bc0/UZSBQtOREf
zVzhg+cZyfP0TI8VJSYBK1rqDu2SeDiJuiFBTfsP+Gk7D4zyvG6rqtlhbD3Ocl0wJIE0RWSsK+Xf
CLWyIj/iOJ498VdBfkmmMx+jdx0qcct52RgG57lwHJBOAK4p6GDU+j8tEV32DxCybRjo/MtJ2m1h
Qsr+/Z/qqOcfa7U7DG8Mqf4kYi6Bj0oiCW8P72rVk/XzKKUs7znXd2GgV1L8GT7+Dq4+d73PG2hb
Er1y7aStqplwaqN/f4XXYOSyJRKa2DMteEqEPfvn+PoxvzSXLx0Du3QfH7bhOp8LjIGl8RYy96aN
fHx674NrMhAqqVo1MQGNOA+v/Dfx8hHJLsoRNF86V80tnnUtEhO/kxiAbqZbSJ/VwQ/m4axGHCp1
PJ5xq7aeWEncjpEb11lQl8giaq2RE+yMVfEfto2eUmBpbba80q0aqkorMO0wr0viqbsh+p3ZzcAv
AUwZDKEbr0shC2HwHqWV9CJCbMZIsE8Cx93oSaZ3t/jVeroqFHMKzTi5kZewoJZglem8Hlj9LhaV
Faqk22oV9DBaV6z5Kxps8BVqNnid9g35OkHn4kXjlDzSkggA8ipkc9cdCEmKC1agISTFxqGqc6Ga
jNZi1xk5TFQPDZo1jri/Ao+rs9ZThQJ1u1+YUIgIE8yfG+Xhgh3F4yhzidCbEf7ZHuUZVh8BDXzs
7TrrtTwCqy8LUS6VBNTyTgjC9rjZ2QB4XUFdiCYd00mktS73b2SkW40z/n2mLYinJ4IsD48+pOZ9
JAJE2n0JdmXmeRZc4P8xBPXafTpK5Nqr5t5OdNe8aAgo9XTY77ZlEEZaHttSnyXT70Bubar/o96O
oWuLRmZuz7fl9sbakCflnq0iVQLqtSsMH1DUzfB2fmwvZCtLsPaF5mQL68csaO21muQwXufoXzwI
X3VJxZx8fnrYI2P5JYagMwrweAS6vms+khMZXUbdaGn43stG8d7E6v+xZcw4a9wz9vR3QjJtrmP3
NPjUsX4s6bl5NZGdWNX1c8/UigSVi3EZ1TMO/+yBoRHLKtW5UP8UT+ndqCpOIFd+dU/DaQpGIdWx
hAFyDrn71q5/nL5FACXV+QvsUYbzHqTc+jxsx7wgJiHgaQSpmPGhlfR1HR3IyhV3DWlXfX0asctd
VTYyr7fyYHuvMgGwtSVYTu6cZ4Y73vwVHQONQrsmxqHmTjwsJSx/V+rk5mj1lGDNoxMyugAOVZ5G
eukkq7JDvUGJYwsX4TNJZNgNc5B/5HsnAIaZzK4KNlhPdbV/R3lfwrl3cBcxRmNEmXaAzwLrGf3Z
TC4cF7dRaO6k5rSMhpMOi1lhVywfVbyQz2geKwWMIzbECxfPuWEhej0GHBFJN4+654BYRTsxeay+
qTSmg2F0Hlhx2zuRSEraHcOgs7d44Vs9ECaUuQ0/W2z5BxWOlnqdf9Mu3LDGof1usZ1+d8/OlD7n
1R/P2qKGgp9Cj46K0F7yogSG/b/DP8OF5e8uppZifCXGWM/v2OTb7w0Jg8aRZiJj1RteXpKtW5JV
T3jZrPCn75V4HBD5lvQt4rfSwV4MG+Qa6/l6tXAiS0y1neB1ysEiP2mPHDnUKvTVzTKXVMx8BW0C
g63zn4ukeOcZwks11WSi0mLWJY8Cr7TRE5lz8QPU6Z/ARiMnuTIRnCDQMC98VsJlvVxHpKiHcLwi
AyL/sDdjko41Co4l4IJgvGiXH7F5w0faULCo2k/au2VmgJCuv8NfIc0dPSR2pITY5oboi+RaIrcc
+BFHIQYu2bA92IhqtF1i/qQN3ryjIgq7ejVlwndKRJMeJN011c2hLCcK5DdNrRXxsQfZiaZ1NIJK
g0stOFkDTZ9qk9qvfDqtUxKpGJhEpTK5EVsA3whAT2Ma2mzo5+wtbYVyBGoL4pyQuJT6FUgM24BM
66wkmj09Flx/EBJc5uKJ+BLBaNLYlvHTIK4YEAkXp6JNaHDc3GQ/E+d7rJxMEq4bmIzupumjMTRr
GaYIqBZFEu8ufMKYENP8lGt49Ox/PZiRvxI3o2mZvpRCbC7AyFBNW64THn7yihtTaH7sXcLPcrY3
qCFE3lsvKhv+rKA2d0ME1hm7JHEoX5prp5EUQ4eYbqQuOwCpKeNP/B5NFiCK0W9P7wxXPdUgFCJF
o30+gmCdWTiuS2IA/UbFm/Kw3MX5m8Iy9pTyU6LEJL8L4a8tcRANMlQejBdxau6cOrJ/zuxqkyuo
kV7FrrfbmM/wSjGaNBxUXcaInoOqi3IcDzYgr6FPoOhA4U2a3CJibXKTxOSxVIJDQITW2vGT+Eo+
pBeq5lYlMdOKpne1F3pKLUQdrmzePNgGZMnHRh8LdE8v+W0/SOVOPD1zZlmuPSFh0RbN2ffIiNRo
6cK2i/q1FoWXay6M8hDnASRRWvH2UeIdGLMIW8tTSjuBFGyEGW9ddh4ma3NCuPrRrEoO5P1EQXhl
pDzqQNrhSn1aQ1wO0vRcpTqN5/vc07gzEnpRPGKhBPMiV9lINFeDctEJ8k2tsn+BGkIt75tYRcFH
MUlJVWtdQTsd212vx+GmBw8fCPTtI+Sh2pbHXZRBOdzprZ9zUGRfgR9NEEmCOLhLLbwDKSPFLEkJ
4Tud3rPm5gMFoAY2vKxdli6HvyOYQYcOK985stFhUGdMlPHOkA7pXigndwWme1ZLc4/uXZE6GFWl
rdJvQ7rQguYDG1IRIs383bBKX+n7dCu17EIMe9xMkTXcv1j9Y7oV+lxlSzoz11hQBWX7zUef4GuP
bHY9eq2Hb+rOiCOtMMlfeuneKP8jXgfDNIwGtu7vkLAKofqNcB7RMJ8kI5FlazhjNHSU6ScPELim
kX3D9slTTBL55RH8/odOejJ7zOubGiceBU+4ygVtX1thzyC5JHQ5tl0bVEjmw0MAQIfqukMl5NaB
6g1qz1kcy/V1BTocVzVZiNIMMpQtQYUcaFKMQNy3V8gJ2KDg49z4J+G0EEd5h/eyQLHVTyLseHtk
5uZ1E/QpJTMNUMlfGjy0UZFCzKOG1CmYe1YdeWOKYTC2+Fysft//FNYnQZGtSR5D99QS8d2iubcg
VMK7Mmv+CRZSAgcePQMCltpQRafNHdEpmzJHMFDAnr3FwNYaT4cQVazwsfhzRdTWaPPw4fq4H4jN
kwOOXGrNXYGeQmAzzAWxiFe2zHs0hHTPfAm7OfeZ4E9yAAa5tWiHv3ApvAGv/O2jdDvQRnO8hmAR
xyPhKehD5qORRnrkaYONQER4vAgfr25Xuf2uedzv5e8M/Ki4PZaDro2MunlEVTgiPV7Azl2+vHmN
jnK85tpLmUHhA6WEL0FnoKl9JeHlbdJhV0eN0Q8dZz3XmdWQCZ/qjUxMvSbZXojP3mkZzTo9greT
HqO14VPW/hYuLdcDj//TtmyKdL+ZenxX0wdni0apnXmVhxK6wbXEv4TchzqAZj+a0OtN4XTAZxuH
U0VW55v1wkGyTZvzEHmYorPQJeeap2IlQnuDIAiocdig+fjtzqsU+05/cDYTshV359ufDqoJRopX
ZKyWpXyKYWNdGpTVFgF5uUgH7yPwjDQeiFRsRJ4eoMzqiPfjoAdl5lkPSkEEJTPzizm01SzgcIiX
kBaFV1k7VRFrcCRCCwBReMKaMOa35GUke1F+6vcWCcl2yz1SrWC/f0/1S9D8y+fxqLOPEKEkLG0N
6k95Oqexcc2IhaPK3uBEE3tN7H2JP/QpKGdXtTTaFPvb06fe7waW/tqtAV4sMifgDl3nsE+RxHmw
SaRnhcY3E/bkEK6XoJdaa8P/IQY1lu+AdOaUuZl1t8r1ucBirpDpK5WBw9kLQEGXKGZYMTs9rdyB
WAo6fArHFxYIYVH2cFrRKt11Cn2h8+eZOsIK0tVOytXTyB3DzO6BMXN1OMAjRX5lCY8YLR0NFC0o
5MZPhmDAKJqLrCuzU+VO544LcJbJVfa0uVlZgdgaSMxQnLoPBlMge94pRHyoGNrIXgS8WURTGqLQ
yLhaBty0CkOq4NgGXhlciUadFXWfYr/sqrIlC10wQZ3+1Y3NWx2dbdL7Ad7sHCZhQ8k/H1+rpPIr
DQdKU8FiAoDyYNWxXsqp6tbXMsiUrr3/nfSxJDNSpEB2sZOh4hp0kNxjOp3PCUbxJRMKi/20p8dE
AhVRXg8PY3ltL9uL2O8QFAFUl2q8bZKJMr8na2EuUldepgVVIfTXSCP2xzr4J3CuyCV+xtS5ODKT
AHLCO/xqQgujM44nnw8JSCKy4LsAo/z2Hq6kdlNYn7FH4rG9Mc0dKceWGrfgVraXjZGMwx5/6JR2
C4EUEza0iSTenBYbhSkAQumWcQPmOuLJ/kcDn3nPRiZepzHTjx7Rv09cs9DKbnduvyWU9qK3ILkR
CyPfqKEo4m1uZXE7ZpyUizaFIZFhgeCdkHUDimMAqsYODW5626ShGje1mEqEPYTCBQtW10Uk8taB
1+/NU61eQT0JL7HmoqORFQ5JCp2MkgkgRhzEWIidehhm7y8z+Nuzb69bXccZPKZivpnhjYCdFWQp
/K2K/FKZLlx15G/I1bEoISfA9HHxCnJk0DMhFvKKnNkiuxAvl+WtWPODgX0JIpkzFozWfb/sKG1s
QbcrSQyUJMjzGUf9rTbgqPlYcfb+tZ8f9Hs72gEEROJY5gx2sj1AxWByZi3gEKwWq8hSx+RsNqBY
FbIicLD5/dIO8Eu37wnAuwM+xI39tqWthkeQVcW5tGDGJ0ddYNAs617f15q2ORZYhtuheVG/od9j
UiaaOu6gsZXpZ21Vl2o2HDQMVlIuZZ3VVzD025poefkOonD9d5eZy57ChV3YCMJwhxCD5AYgkgjt
iKnV5vt/NNH2F0FnDzcHG4oA+TTE6NAs+9/Fc8CFrghQdwbWWRlEX5SUjM4nRj1USIGZLkWVp2J8
Rp8dAEPAQc6703bhBIhUr1sfNKq2Yy8wJQdoxbV3/BPAqICQJO+zs3KJHhRPqfHxOpUwEQ7P5ZKg
iGVrHt6C+3iNpqSZvudZPJwABBX17tGnijr2xCIW1rY+JcoficAOM0j0E0jYCdkUjg5iSWZ7hEBg
PrhDaI9u60H9lKrpl4QonnZ9erWz6iqsI8pL08YBoWaHsWZLKuXbYzf7d9VDBX+xH1KxcaX46U26
4bxY3OfSSHK/nH7GsYs7gHR14srXhRKUe7M4XoFULfl9Q2pDpfaaLCsswzgohAtoujX+VJEtKgg2
QPJi0GPXrw4iAsADnIxZ568+l+rIzZzzo8NDlE+3ySC7kdJrlEZP9JKWv8wdEsRk8ZrpbDE6i6OQ
JqxUHew2qz+S45aqY173yrsQsDR1ZTxYYghute20u7ZgQ7FPgOtbdGKvCGNfZFuuqYUPoCL+t5bo
y3fndJOOG4TD6tr9cISnV5RbEJtsNgV1alQKh61Jj+LuLFbGJJcwwRtb0I7CIx4mcyzaNPmkx2rB
QtMpupIMyb1ziytY5IFpoNVvnEsqXoRqUkz7Ow4rGvkrAYyN7oZs/ihQJaKCTlZ1xo++X6Gxa45m
EsWTjzEfh08uAJLZG40faERjUpNKoBEvdghhlM9xlWLBo9YOHybTAf9+ZHB1kLK+Ls8zDhwHgDhL
Pa/JOhc0ZK2wclh2RBByAEHw8P57hpRoWVNpoyA0qXC4ZEoFB4/CuySyxHIyxaFyWWz8LRGLega8
ih4Xs2Nv/rpDQa22OOU0Hpb3ws6hJajQ9wzXcuYjMf+qhPGEmyliss9PPExI0fcSUJWcYHFshbIX
wbevwn04TVzaBI065F95371BYcXFxI1GFA1HY5vg4AoDpQ3BXFmXwrq9rBVXcpaacMN7RFBMJ1it
OLtVz/F92H2yVx1RwO8D1LRiM6e76m7UJnE0lV0cJY1Q+cAWjbO84fNwVJjdYXy01kimIVozQ8E2
ZIwFy6cz9R8Z5oYeUBiLxqAPC3vS1NgIRXD94MhJRXjVgfrmHcXzGjU9LoUo18ifUPxSD0ucujU0
j+FuhNx6r7LiAIHVvSP5Y2Z77ykVuzWYX9SMJLqYcoJpm5HK
`protect end_protected
