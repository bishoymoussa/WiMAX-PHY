-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
gyTCIkJ1yj+bPCuGYslh+nsR0Ru08EoabZyoZ9MeRD9A9fkuJaxsb9u+Pejx/pmWg4J2V1ucjuYM
IqKQapT3jHJ6Y7ca0cp8yuo++9lBf5xEICxHSsW3D6+4gynLFd273zSmWmoiSZKMfdDIKFNH0jJp
VqEYkSk1q9DEIaCfBZImbxWWjYKyEH2fD3MjlrhFft6cJPrMF9V4p76W1G3OGZJ+pGBZEBksMMgw
wa6nfAAMO3TynTBsYiQnlnKVwWa2xJ5xx3VJqz+21DGfkW0+C393MVQMh6iCSVW8IzBewLcj2v2R
qgjqmjt6ySLMqxqNw83BEbOfnbOZdQZpu/F/kg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 23808)
`protect data_block
rCD6Ytld4JkY0ANMyr4Lu6AdzrJZjmTOBDnTrL8ox0KJPMnWT9D3tm+CN0bm0wmF+djfMYYdmkuN
IvU77l22TSKLsUhb4xUUgEPUvN1/4pjF/RirnfDRQFFdFJh1uhW89aC4NE+jXvvD9TFPQWBwV5Mk
kx9KCFHpzhz3Syms45tkIUk/hj+TkmfhvqhrFLiopXpGJZ6I0Lt6JiiC8HN6MJ/t3WZcaI+k6/zY
ASN3KrugU/8JD0SGhq5qg3V8kfiOnSzfrO0qU0caRQNhIlSRLNLS03Vzeaz2kkH7dK+oGN+zMjtT
7PeuaJxy6YaANYpQYN4hrMj0ZMpz5AmTzgcYCbAB1hLDWnjzfyM385wMzZYtk035IIurnhwnXHoE
m215UlgfqebrPt9zAhHwvXDCLZsSW8m1VINbNHWiZVT3LnvvbZr1vdc3i9K9HO+vhmPovFldCCFn
DEDZ3t57qHsnARWox5E+wLret1CW9hCsbKbTNPLVw3ddZyE5e6L48LYKez86XyYlpilxXhy8S8F0
DHmcCgVzh3N8nZewjXt6d8vxoU0VDPD4V7ZhTdSB84Gnmi+raVpGvtU356Q7NAeRi+K2OrY3o3hk
Ew66GmsiT3TNSxE+zo0XHZhEr4Vi4atqBIhw3bB+DSkASeV3td2+oeUyMDmdNemZHWBFV1ZQL84m
E/2w45569wx9NdpCiESAYJTLYEldUIRsnM5KjzyBSfsv8YkoLNn7PmVfMBF3D8KibBJIv+ZCt+wU
qL4QU8V9PhFGftdGpGNgeXxuIRTePHyzYUH2HPHk70pvbsPcUax+NqBQB5/88yPzgLZ82og+oVEk
KTdHNoiqbt76Fcq0nQboma0WV9dhIX4pNdJnXpxL+3TUtHuYnWRG0nSef2/2+XSmR021QkwKyEET
pqIZCfCTK2NTRkEDKiJ9cO2Zpgg1LyzgpGile4QhAcnUlsQOtHuyh/VbSweM9era9NAGsRs/ySQ2
PanawFA42lpyC0WxqPe8HPi/UiERrn5oU6M+Y+MsTBHgmsoyq7yZJ04BK1bMl9Z4ck34PktBUNBu
Zpof/hHoaR+R6emLidd8clYP5EzdLwkT5PuTJJhZErZ19cwZ/WDv4gJVgEfNbBttIJh1RJjiPTA3
Vm21RLntFyeVmroCwF7hQfsZIaRDAo/UZpcswwvtTS1tsB4lD2kVheVhSK5xUXtUkgFvg/c6Dhjh
ssV3fMIWsNRCO0dUcQp1rKk5McMoUlJz2mVbjlQEfG+HrlIczbBqGqxYXxIMy0pAAQYPQIpuHG+z
SueENONnGFq3AKI+HbiG9zPgAO8XXtYm7Z6hg7GdEbwbqeAhPEeumbnOHu89s3LBXcjv/vOOhIAZ
MSzdZeY3H6FQHBO8QShNSS2bqJdG32VUgqP3K9aho93AZH/zO9YurO42HImKZHq9uOaNMU0+Buqn
NjNHHPrl0ztQi/E4quc2oN2wWQ2TuGOHwo1T2dnQMy1emMLtvFCnjG78eErwrmGPDbK1SxW+e6Hh
uHVdvHy3zkcLqJ3Gr5pw83RGcHx7TD/W840VyesEq9hWCVKRcI4aSCN1cJnM+ltKAdZhN5XXoDb0
Gi705y9GBuG1VU3LNNkj/BPzYj4C/5eEbxbpRKNZahFt7DMFlLPIakZsg/hQOxHIg50fNtz7goA5
11mFV9qlHqhXFhDMH9bFjdKWuaNJx+10igkhfFAFx5rv1ydQZOE8iO0eRGhuBpgXk5XF0vNKDnex
CejZVNdwRl/wWUHWkgcG4Hh85g1g4x3RroDMISzWuRUlqE/P4/Jj44iAwtfvwl4H8wF7S+nwXddi
f/kMbU182y281YcOKU8EAig+JfAJMRMQf6929kJt/MPNsXRsFpZ+muqE0Tb+8nZtQAH/j7VUEe9j
WmkER+pF1ut6gPPOCLFQJYoKXb/o+5AJIgPPd0wznf8OoyGou7k7iiVO7Fs8QZPpmUZ64Uzx9I7q
SjRLZO/5gRJK8ZSa9MXChK6M9sBh23Y5GsizGg3VxTy7rGMqmeZiy9dAWhv2NsEtyz0SvG0KOx5d
osCPuWLZdNDT41decP3bodqAX5A0reN5L49l9qyp2lRhSqurU26PSx1tacvbJoSu3BJ1TO1Bx9hK
+5BYgGnvAUFvcrISUFPV/qb043J77rVzBjRCnA2Z4t1uHuA9LmqCtUfDcsq2XUYWmqiiQu21HsT0
73UroBzMZNlcKNCaUmwIsS/rwd9SU+eLj8BeYcxjgQz9vXpaLrEP6IS/YIT0yji2PnkkK5keAJ2k
jIW1yZJ7IGYJ9G5pU+/tfUg84VrL98rCS/3utruF/USD6jQQQAYdgxk9p8N42jEyQCWE7Kbw2NPW
0VPnDKTWoL5zcXzfXhRL12H6jllJXC7W+wge0lWp84L3Cffu9XlKliuBdAYfHIjrArAL9SmkxeSS
tzIRag93bQ2aJzdKT8pnMB7UuOVof7wJtRyLkc2/gKO2PNIed13B1+gI/pTNoCE0xqFQhVFc3lXU
rdAgD4P/ojJaobIuYygNHKtlcokRvP96PVeSuaC2ej6LIueC+cw71dKYGCaXfhD2LrLnpT6nE0G8
TRK6V1/dlJlZSgIp3m1Aw+y/6FH45GZEyIuEMf8rMEfNSjJ1cViII/ipmNeq+HDJtaXxI8Uww2Uf
t0UT49P0M/usigEYIkwl+JE4SnrClZqJ96nxfIh2z/whFwtYLTv0Uv3YouIrk1H7NFZI/L4qc4O1
/WFcEyT93oimOM973qnEDbXcGPiBlobDrtM0VQKGlq1Neyyyl/QvjILpz4i4c6KOsLuI/+HEooDE
o/KXbgqaTcG4hSGX3oHlqZ0EvIah/R1MX4wf3qAUFqO0R5dUt293PUK2A0i+TYLzQZ3Y9MVk/Lsg
/JeAzE/x1Qmo1EvPRKTWo1UUuR+ARmyTm4XhwMzJLDpCW3SNqQEJC04kjbTjs+431d0LOeHQLYVG
+drl3ffXF25FZma3V3vgoCV72dGtbDWZI79GKPIhUHQwJY9kHUI6Xpqw8gCsIeu0RXuNC/WY6xYK
xtjLSZ95VDGKTmoHySfuApAuVC5yXrSOHDe6WVBJ/usAUHefV8vN1JjLE1MUpYKqdVOgI2zApjFm
joIvsLXkK4mPuVRABx2dCIOsyzrbPhkW7Ll3k5r9FowWMLH+m+pPLKmdpZMUeIdpprBSS0lSECz5
5xunidkgyTjvLNmcwSTz7h1ONxIxXSXMk06794FTXXc1EfrwPiXne/nuA5Bb3MP7EE9b0iilxq4D
YCqn5cPeh0UQwtKRVPrpdKq76WjExWV106dvuRmlmKF9pMQHL/ZwwjsJx2BdIIQRBy7GYcg/Bv5u
Tsd5N8QPo/rcNkTKOYGJ7+tH0J0nx0ftpltpycGGiFXSaRrI/D8qagMkTq0gcbJTF6McYIDIeYzD
b5l8iqHUtdas2xeMQLSRfZ0zdjsvVsAPQIoc1WXJ0osN0F/nvw2LzhCOLRSxsraef5BgrafM6g6u
80hK3h/JY1wkN09/ffHt+icQDSBHY690nM+R6nY9FkGcCIljtaDBrlBCeBYoY+qSpKRvG9NCkZjU
Gh8gV58tU1AjpU7hNSuyBWWRnTq/brdVmrRRyA9zLNZcvv83Qe32AyOGdif9SB02i4zFKDtDbyRl
bQ07Iv2JjgPTfRHGSfKIC0Pm2HSPdO86lwsq5oCiY16VmH/GW83GAzdHvIL7CathdT+EEHDEHMp4
G4Ae1lD5aitjblTYguJSPS0rauQjFnU396vqpA/YjJGNlZeZvH4vjzf7ioMhvEG0O0jIqLMsySHI
GsCMEv9plh0mPCUGMbWRuQ8Rttb1nRA64qbGWdCsP47ZX6lG1G+/hyXSS1sOut8rX5n8w8xdgios
8hXAC3o2hSmt3KgXBrK3bQhUUv88WHqZPvUhgGyDCbSEYcH14gMj8zo3+HjksCkH1f9Zz++yLpDV
q/scsknihY5rBad2PUVp4LlCbuvDr/ES17mredeVJ4c/7VWZwpOvUoKrCPl+0PZE0sMuURGyWGXL
/vYW4No+in8Fs1c9Wc9B8VhhM5YVKGMnmg0KvhLAchDrhBOMdkK9le97Q+IFoMoqNe+e+AXWP71P
9FFL97kylyl1oNtgIQnpONhj0y3F7/Sfijh4kgfcH5lwmqqrZv4SLt5fcq75RcDMdgBOzNsAu62e
h56jp6lWeK/FEHHnIMaPPi/aPmivut1yRaNKG0zAn6HxMkzxZlBCqOlXkYSZG7w36z+tTas5hfk0
YQQPPV8VZQY7Rwc3lw7dOy5MV3rk6b7OmWgdA0g9YoQxMAkNM+8PTxjzPuZT8WKb1cif9JG7H9nM
VBDNZRsrijR/+sz39iUOBnyoNfMFtVOmMp0FcR6IIs4YQ30Uuo3OPXvT1Qldb+ZtK9llNVcGhXyK
q51G1O8Jh1FThRmHYgu1n/9UIl9NbT/Een3VbaQS+B7KUvOfAVct8qUn2+Jr28dGSVRbXVM+s8y0
m7+YA0okE7Jt5xr47H189khL+F4W3g1sf/DgDg8cKixdUp/dCEwHRLMMBborWsnvrqvZU1GtiV5S
7dEm2o4nhGZTDF/BtilrHw9eabLJnPSEDANhv4rwNiiy7qmaFe4wEEWMc2zt/nMDE7oWC3ijZtWL
kf6TZBBFMYhqs833WYQsKy9oII9ZYCFYGNkU6rwOaropNPVHxY4orAuErBCmm0AkLyKyxItDUIUt
j227YzPlHBsXgsWId3cwnMOO2MxtZVZQEHv3ZsFbQVSxhMotenoj5Jj3aJi7NPyIZbpEZW+GktEg
2VPuG76D2gxFT/qgD8kxJ4Gkzz+oYlCjw4n/2RnXcZVhA6b0GoB19Aqn+nm8N93r6LW4/d8Tb8y4
ovV40+GvyGlmA+pmPIlhSY0yADkKQ43RlyXt108KXVfya+KJAFT5lAt8EHYkZ5QcmzCdd6P2OTQA
F1i5qJjBeEJTuQhHmooVNnNcsVfxFof9Hc5r0RbbnDIEyTyy9jgVNfAnat+mm2M8P9QkctJgmFNq
kezTED6Dq4nKshklC1fRRFroXEW17X0QJXYnOF71kFyRnzeIpMyAUlB6TqgP9OY0QsE90X6hoOeY
vkfw8s23pOK76EBmKYEGMA2PzwiXM2mBONmmenjTTh8tR03iR9rcjakpYSBv8r827N8lOH2RGKLF
7cViTkPfbzZCf3NVQdByX+t5Keu4ZcvUyD5Q0BP/Wa46Q/ATOy5Qdt0PYaYI4tjvImg0bELSTrSD
/oDBOH0vwQRTq4sCIgIGOhm3ozuGz9rE2HLgaB8xTGgp6G+nsR909POhlrB6qpXoK6JGQ5jAqFYO
kCNFup+QB2md/s/w7oYXxcubsW6TLwF/47QJwyTWHUDUYDzrv5TpXy/o1QXPaYYyj8Xbi2QP/rtS
Roew0+KwfcxZkUa720ZLT91xP9zD/MPwSsEJcy8y6kI5m/1SS3oCguRhCd9vK7LwgB7E26j6pWvd
i8TZaCa5P4/KOEYTjkXtrBQHDxZEPDjAteK+mwNiXUES09a8PfAuGTgTmZCkwMMxt97TKbSPGHgO
5Z24/XiGjMbz5Jj2D863W6ViXGJZUj1rq9LZVEJgmiCHb1iC78uxjbR3XF6hOxn5wVZR7Ynb6/i8
Tge25G125hUzBb1q682MErsGCptvzF7UHGsLxNUOW+UbK4B3bk89kGoQHG6B//rZIiouLoc4pUqA
Gwvzraip66PL/MiVGJwVlkxuYwY8IBt0mZd/O5gd9BywFrhvwYZmpEz9aySjh1Gj0PwUWZfWWzUY
OXvc83AU9KdJpFqVnWdVDkesp0m+CJHfovm0/Kv446js6Gzo2T4zfpftm8DVRo0ePF+bb6+ZgxMY
zBQnlF6i9qvxdzSUPhRzkVlBjNExFXtP5NMqsgYBbDLXVnowxDgg5HXxVtFM8bndJvYuCAHRGqra
86mT/IR39JJcNY6bCX5QFsWj2CcnMebMQbz2g4kg23hfhzCOo9a/P7RyEWZx7TuGMi+jnVmZjrRr
w+EaTtVsQus/c/7haUagvCYgE2avMOLQnyod8vLdZndoEB8dtyZHna15ZdhYVerb3yULoPMtzHSJ
pRUi5jEEgkQ8lSSp03ov9qSjuJ9acvrqBCdmpHxO2J4oyqn/lCwS+IHuOrSWyV9qselsQ8zMnvvW
KdJYQffw/tfgAXMBQ7fKeptJvvGsn8leb2PCvXj7NWyqMasMuvJ1ssmjP+fBrOf0TlX5DlkqkYNu
mRnJhnMLlKCTSOQpmOktckJKu+8AqaXY64EoT6SnbuSXWgi3fnEguARcxb5hOVbW0ywUtrGSbn5K
FDkGR0V8c52713HjgUZbZT90zpkpLDqOz8Rz4jUEN9/9IPBUiTAiZGcZwDWFOT1SwhUwKZmuJ46Z
i5ITaq2Jza3qxJTXoBbJM0xRWoHnIZr4koNCbY+i76kqu3gXHI1tsf8VS6aC46/hD7ZxuEWgrP8x
kQVzcbCB0WFjhf619luyrNZs3zlbTCfsq8T1XP9PfQsH0j6YYa4xfgez5kYi0VHUJ70wZzgt7cK6
3SrVYkSBXR24u5NBKem52LPXPUt75A61KPZ9rizT1YCPrWeilsUm1morkFY3en0uOL3M6DdOZBRn
6AlUxiNYzHX549enHBAMP/A4ajmfLC5y8/3a3GmI8UJqBmVIi46w61+yUUqel6ZcNS7WSBmocaho
3IvN2psjfonymX7kyODwhAHS3SaKwafDS7Cm9J5Vh2Pr0wg4DxNto2fsQe0SVocIsBiqnAoxVZ+Y
pzh9EE8Y7aYQRqDVGaLp6ZQUgXd82c5MtKnXIbqussnSpuJvZ4d0qgu3eickGrBqX2oaHFuOuwvx
LAl+MQOBWcXmu/8ZqGPcdUR7KkvdWoscT3V1jSyy1wfYySSOzaV6UX/XgrqG7vq9miNaDtfA2sp/
GVd5qtHETmFo2Wt63hCGM8SLSDM7EzMXQ/zOjg1CvdWs3AqjH2nml61na0aMADwA4JFU4NwEqEqo
Ge4bE+wF+nPTdCQCmDPYexGbFs4Ip1kkcn4Uigb2uQlBd+Wn+77RPSq4mTUckw3HJgebRmMOXlqE
EgcgjwK+U3dus2UIcOuKE6kuSg39cf74vJULgupTPiX9b9GceyY0wTzsQWztJmMQjm5Gm+/QtKJr
NAGoIVFDhd+D0U52Fpzp9jAzgt2CZCb3w6I/Wvkm7GKlacI+V33iDPLjmW8fVcrLRIxJzKR+chlg
3mjGSfNMIaT05/9qehPggVopzryTfz5gLqIarv+CS495baMW2PXfM0ZslPV+EDPPexhxB4E/mNEq
V4bR2NLPCZ0hbRUjRGUflE4HXet/fuYmm142KQCsD8PyzDnrKnu4DyKeKRKhrbIiHhzdQ1RCFOc7
HUYAnmbZLbwDixTygAj3glqc7N1msSMOUw6cJA/AqllZAGeIaSSMeUsuOwdhhr7lra7M8PZ38vJl
WjPDi/BtYFOmDvzh2/b0ffZuj5ByIZpRY3H5peA/xf5YNQ/Tir47FTxGADMbOu6R/8tX2n3OGRZN
ktjrD8OxHf2hYZ3Bkb1u6J5Ii5MNy4CMjkwL0bgKSRd3iAR2uMRjQVyk10V0ZMUDHW0CuBtUGrIj
k7Uww1bL7gvM6raCJXyoxC++SXtb9vVgR4miGwOz6TwFhp34OI1sMxbJCFZa7Jeu0a96bT+cz42S
WmBNRQONP+Av4q0hQDION8V8V0TFKJuoR4NxaZ/snyohPg471FB82dquhq5Vv2xJfBbtmps6nZKS
xlV7BHBRaD7sZg7uxU7Co+1Tg6sz9a2QohGeEjjLol4PdakC3EMPr00yuOT7QJ+mYDpo5bs6VC1T
3UcTmt+eaxYmUJ/nH4mErX5a6D41APfM6F0aiioQKWOmd/ap7oI5gNIETFpskHkVavXC83lmXT+f
iGUfBZ0X5dEO+aYJMZm3xJn9cOswDqQz0exbGZzSeWstkm4dvvk5xiTqyjc3zrULp6yWVEoWoBVB
5/aENfKt3NN+mLEp/58VQaKdAKSqVWWHN+IbrOCgyVZeqO7w7US9uEPX+K+ZM2AB7gvBbw+OC1/6
E5fBrJD+UineFp5vynx6Hh65Dv9sOcAkPTUodg8O/Fx1IK0xWh/ncDxCETi5BZRBOWguq7G/gHg+
Dh4sZi3MmnXiWXXwY7SIzdsiqVDny/zSqj1+XlTe5fklWxIaknlokJOu4WWSYTQUgGev+/Y/CWiO
zXwm2qaso4x57MHb3GITltFYuGQQNA9oPMc6a3ESi7tfS70sqwaBtUqdyc3k3IQZrkY58/xrPg7r
UmkG4YWTo9dz5KCWWDfM0Nmg1fwsz0Dc2+1QPVHY+jVUz5xxHkAwrqGCHgxeBJ/F7XJSNSzuU4BP
I1Msc4X/QahGb214N5oFyE0ch5i9xxYnKYxSDHMWSVvBzYqIqX+ilXzxLgzJc4YB1krXQXgXhbD9
cjNBk+tVgisw6SldbGS4qVnpUFtWLPTgwdlyur5WvGF7rAMSdNb+5TxNBrSV1KiCPjKSN8r+9Q8s
FZrqAs5QO9N7+8GTCZgj61jBGabJ+vJpQJNOVD9fGxP71e/LdDsPfZgNddur7T8/gkdOPOHMx7tY
Ln0on3xdx26M+hidyscvbLKx6T9J5qOup05rYS21v4D/kPucyC1qU+gpbyG95J0dxQP7xACBn8pt
Mt7eR93S5RHacX/WozMoTBp06T227R9RCVj8BTYUpJi2RMUv21kFVXwcwo70N9EpKuevQHYD2V1e
gZyf0CayCeIxuM/1ruZCN9pxv977PYwaFKj+ga9s+xNmZrXVnvnZr3zrFFn68pxA30qdiHFuacKD
1gy+jroHn5pYXCjWVQn4r5EYQ96mEfphfOosJryKktjwfa5RqMqLCATMfPU3EMTR6q4aETV5BuDD
jW0+2trQdQdYro4WcjyBsYPy0TuszJH6FADpoCd2AwME1QVjI0237V5yILpJrKEtcR06zCxYP30n
sWZFMmTBoVXlJnMkkM8GxQ42oYhro4HrB492e6Edob85ISBXpH5GXMCGcnC8ADVOPDfBAsrfakhr
ixd7XW0CUB2+kSrLFROVDFx7ugsM83PF8pN3FoEE1uKnhvSX3yKkPXplC14Ljb1byTIKyt3cBQ7j
9ny0jesb11ki6sg1qoryUl64ilQQrEkpXq4D6ApSjjWympJ6HJ53s8YrZPKCGVNde9kVz64gGsxG
eq1/5KZeBVA8/N4qV/9iL3X/LqJNWICKtTXA8foWY3iY6aFwUfFrEJx4++hoy1MGvEpmP8bY+XAq
DxvFi23IMvq2B9ZLtxzYTKhtFz+u+dRX/nKbDNNydzknQr4PldFkW5T46J0fwIvmAS/wvzHs+KVF
6rIY+ubFCP2uS6l9k4L++DDljcT5BMr6MPO6QeBthrOZI0l857ONMmZDBk847v+VwFBHrjgaqVyp
lGEq4XFsueR/EXdWz+QjipAVtnGbCsPco6yyP5cLyyihYfVKjWzLr7ZszAYCDKNaAv8tLaqx9bRK
kLB6aGPpbOrWwXap7p0d9qFIeCbn1I6rtFt3ENjmSCIXSPqkkFwTNrOK5IvSWNI5jDVcX6gG5gcK
2wUTpLGpfLeWBVzqdOvdHPynb87csybTJMb/T9nxCyVZA9o4yYOMOWGFtKl1meCfQFgMUbyJgcL1
M8bRFVXDO0WUqYF8rBilidaU570SUDkoVPDugFvFyYBD4YyZxZtBC+47Tg+qWjW46wKapBB0DP4b
YZr+5t/34ydoEEewdxXtTWXJLQoi+98sUE3/ElcDCwnCeh9hbMNn2NTXxtAbfVAv02xWiTqysqYc
k74dtY449QW7VsPlFgxZkaqaP/IAtvC0J/kGW72L0m8pi3uzcsPqZv3MZjnpd0ODqjQlFk8ThAme
iUz+X23ZxNeRVKPA0e2+74BeGbqEy3AkTG2MtRZ1IL76Fw2zQ7DdWNytv8YGyQj7B7z7OYTTRSH3
IJBWaW74WimLqoN9gAX1F+6vgRzYwwt3DwtPaheBMX9YV3X21VbIZhHkxbDqdg2pkAML7IEuNv0B
wzTmcPRcT8sBz5n4kmbbkeBctNo7sXM11cHeaxBjRiImtSlHgnW5CMX0PofrR6brPNx+uhfjKsPd
4aOYqLiUWq/XRaVxP+ZTZpWAAq/JSqh806G5x7Vw78cToeWanESqd4p+Kav44UCLWagN58dbI5xN
oqQrT6nI5htxyg2GoMsfrTpONtF+JAQX+tPHbLBqTd4YXEf5vY8jAfakUuwBr8NPGpv0mrSzoLgP
MM0KROSly5M+SXkIDaOwrbOvqSBxxXPrE2l3mPdQE2Q1OkHrP3Gx3ZcrIg35DvdzUIYwzw5iq0AK
ufxi7477mLhgiabouWRjhsIVimJ0jV8mR6zIuW0LBc5/apZ2Vfqag0ZXIZA1/AJFzWZvpozjRJYY
/IQhcVmV6AhJOOwLETuwLZj1mAEGK00CrmQV45B+2GpzKRbSnDC3sl1xuKjLltJB++G7CAUO6duA
wMb/gK2nszE+7n42+M6WD7ZHxjIgtv/kYCkltJvV0Yme2/Ak8ck7HFWFdOB2O1OnBHsulY09rYjm
gk1uW1mXpKReBQRCJ8zv5tnw0he0GxSV5IlG5pHCm0+dm9cLKUVKShMOFmcTIfLnPQYXayN9/n3O
Q6KvshB3LT7bH27yQV0y9aBMp0qAyR7ulDHCvdRoKhFH/3Q0xUpNAUXr0iXQY1WB59+RCdjCjOgF
DpUhdp655d4ocpTXBtLCKJBevSDdTzTV05tFD9M64DJsd+CwvbqWiZ8ueGPVq8nOIad3o0iGwxGz
W4U6OXu8NuWBDY7JgV+f0huxu5soggVD3r4oX047EyHJFf/a+r4/8Uk5seJMVRC5dsZGsxeOOaKb
z5RARwEhui2wgKlYTf0NSzw9ZHHANNU+zKS4T2SInVOHn++qcz+m2pjpOa1lftDdZ6yTZi3h8d43
9j+xlv+iyBp3QX5ozXhf3HZVW9Ytt4xzhfT3zgynnC9zNZP6/WM8VFSSs5w2fSnuwYbTSI1vWIkU
dX/Kze1SSxH+5+Kq6nOVnBqbQ2I9XKI3H3M1ZFsqWscSp0qyKCqo0y2t3HWJX45wxmsLzF3UteGc
cDAfb7mkT8clWXx6Y01JsORlCNaVBCguWLD/6Xglkk4C7u/y33sklHA5MN+XxEh3P/guFWDnykeI
r7edbyPEATIhDZJejDgGzlstxHAo9IvuHAVFj+8UcyVaw18LBqQTi0NjALVfWxn66/l671ZnIxQM
GIXmEUmc+9gOceaYI1oMU2IB/tRZLkbqv2mGwJr75TMPaY43Vud6WI8tK4Ss5m3yH6sj6s5+otES
j2jXfuuE4f66RrgjjmSKfZ30+bmmzmzNuFvYrRp24VT4hDmnTKgsWRA7QHO7ieU7cDfY6hkOQsvu
O5phVq3dWX6cY0lGvh1JI991CMMuN37YznvUIcBYeGOF+sptkS3CdnKrxeabuZuB1xjjvpnspxbX
RACoYnoTwMeTHZwR+Vs3RZ7K3POwspdsUjWyWt3CNX3ObDHqqlCK2QgQ6zr9O5ATSLKo0QR5+lk7
Oo8U5QQ8l/ddhWgp9lgjM2dHBOeFwc8HEoQJHG0aBR2OX787lohsyrjaDClgZkZz5JEDsfSdrMQz
t7nAHm3Q9IZ+35JhmC2GG0MPw7A3g4Qee7BWACQzcJ4ov8pWH4PmMWx1D/L55ZZD1q7R3u9ssdUH
TsuFOuyPUFtF/b+Ej9psppW/4ORui4nUNzMFZ4AQ8gN+xEdJ87nSHxuQVh18X1F1uD6HESWx30mq
EKm9tbevmxKBKfNC1QU7gAiSwQalYD1xx6Ksy6nSXCs10AEggVMZLSTHxKt/oLZYasANOT8keuiz
7BHJ7sseDxc8T87/FTW+xw2kSbUnSqtKHLRavEDYioop7tL04xzVps0dQbIWoGhTPO1JdGMwPteS
UZ6Pmf0IKTP8XRPH65PRdH5mgqYawIE9PYEeab2lK0NsNzllJ6DYIivpgl4mtPbLW3+k4bJWubTS
fwpNT5eMfk319AoWUTffUjUNPfJA1o/h8fPye8A7vkyMzcHJezlNaJgDzLVVl3Cxy8yHCjSaae++
4T0AQspekm5wyzz7P7bGO/cp07HctMGpV8+8RK+Yg5tBRRZSyVQLsUuO6DIChif3MjT/cpxWe3Eh
CoL98rRozyG7P52+ycbNFh19cxWxy2yWi/DWf/AobT1rVTKs3L/J5L9kSow/8JZgzn9zvb56jvZw
ozTLueab0cSlKAw2e356v6ysV2L1ey2rMZTHGw7fqMA6zaT/9IqFwHBu9Ef3y9vxeQyoqMRadwrE
LEJW/3HmIKAPmjtu9idVhpDNyH/pvBHNnvzlD2jFM7i39FklItmfpfQmlWxGQ2dbqeHnkjktKv5i
RG6AlBf7JV0r+aECVjaPA2xj/p2FSMxiTHMC3jB4QY8CmDcK8hHDM14kvEY8uq+K1RWhQ5sp1aNy
gqJ4rwBrHqvB7hF3lEIaX/SqUdrCTTfN9wvoY3MVdIgIgWAu+qfluAu3u4jBmqdWjwPct/7/MtUo
tyNsBW90ku7/FOgmDQdgK1/VF+ZajWVtz0HnySZYaUSkWy/rPAnKd6B6UFi0mOrmDLH2nR8InOVG
CSz7j78i8zAB6sXDo1osJjaLi+hHL+ydLBOu/Ow9l6pKao4MydEk106hClUaYpF9ZKBZZ9enJZ2D
XtWklPHRckXvBSmNXMpd9q9ABaSp45IrPlu4LTJx017YApppSd3TORnETZEXw82htHibHc2xpZSN
LDpM15cLxLSePZNq6xiR+lLvTHvzZgpe55qJ27j0jRrVcitz93IpDDC1sot0mSkj1ecQiCDJzsLw
+zfvKtfDWLBVqC39d/uN2cnqHMvKAe4it3qnFNxIQtbB80VtYP8G0XZ3MedroNI19HhQiHxnisBN
zMJpMiuGzYovqsQVnzUQIlJRPdOlSo3mSywDTlBkoMf4McbgFh/FjEgZ7bUaWil6YXq3NKCClwzN
GqKbh7HYLwqktjeQ0EIGAFmJ+Qdc4xjdUqISURdGxAsVmcEiiaILvNCqjvaGz+mpmdYldIcKRSy1
mWr9CHk/cPRpVMhdBBkVB6Crg4PwKAmTrClfI/vVMSQE2cch8RL7O2+kXLVruSepYi+Ij7fmmphJ
4Z84zOY85dOz5UYOGojhmA101VU6egJtoNBIjF7zfYtFGokqc4ZZJbeJZxLSrpSKvUU2un+BPMPD
oT1rVDH0aU0frU/2u4aO8albWiTR1tuBZktuvD+nX2uI1z+fnsesB2R/hPAgngrV8LJ8w4BVfnPL
jmRhcmWZFzl1QL8pfT7BVPBt5hPgB0pVeJt9ssrH674rGqpWV9N4PIlhnfSiYXUIcu/SPGuuhUWU
jlZ0itMzF1xfmm6jdPzxQF1dPwe7lmdJ/YFieECuOgVaigh+NNVRUZMfmoB/wgvow0c/y3zO2ov6
eAXBrUVUxdr1lk4Bn+t6U+vONtvhB6mpH0YU8KAcBcB8wlqb27gobF0A7gh/FtpLhN4gJuyEJGTw
M/WPnRe54NqkuCwdcdQa3T4W3Br3HbbwooEktGJxWp/liKLn4R/5wKv3iSPVdQ0Qou9UzxsTIUGx
zJ2AAESzUsCiq9Ffuyy4FdgxvlqZtBsW+uiW9Jb637LWWLZJPSvDDq5Z6DJEz3jsrGWXIfT68C+c
DeI24VX1Q9F0Y5CoxniW8uYZqBlXAMx2ZbpPEb+mnIaUFkqY60xu7P4rQNM2nz6fpUGnY09jw6i5
sWzkVEYjYUqd5M2Uk/jiBQTErKy3Tc8I8mX6lHVPf578ODEf0vrEkH9w5I/yuFUNPP0cdkiBb42X
hwtYQpYsjiyhysqKkvICgu73DkvKlknqr8Xj3Ikg4Anni6XnrUEQdHliBR1L5WnB6uN60bxLQv3Z
qxgSayWMi3i2E3zV/CEQH+V4IGsw+LlOdaBLWijrnpGAJCOYN33UTEO/osp7tRVnm7nBWQwv9h1p
Hlr+BTBl6Lq0CbieAp/cBlQMBJO5EqAXMRfhanqlXAp8/YIe3n/1/xi03gWNPA4dNw14YWWFurC3
U/OpCbHWzbHI6ImuWy6PZg8rsiDoFJR6JHogiae6zCe+afqZQkO7RS+NvjaJlPiTEJOCYplP/k3/
0hhnbmWB4KmT7R5XAoxWO+JXMgEIOMPh+Bf6yDYjulYT5TTX6HfOCE9z3xXpkcg6zV8sntcpa7Mw
eNnESWplnhA6lDGn5kbK/Y5fGcRcrm0WTd7Tn5H6x9UB1mKPUf18GUg2xIqX7UKgOum5T6PtdE/5
0H/N3+/epYAj8Q+bSE8RNK6dj+7kJ0+lUOXOamQs9/Lmn/YxQ1gnNZB7qsLRW/FTO8DcpgbdATNh
dt22S3CXH1K1lRP5vWA/G0NZWV/fpLCU/KC2XLB1rhcG3l0Udh9wHmNdFdlNen4AtCT4YJN6/O+E
nFk+WX7f1OUtZi1w/B9Kc4WgALBt5YnnQIZ12WEAScsruMcbbIyM08ChRS37s1f7+8tqDiD87/MA
wrUO406OIjJjTccpImmfcijsveVwuG2kHXhJ0r8CicmyG41V8eM0zcEYEB2aBcwiFG1/kFzb3P28
Ssw3WrsLOyK0XWmt61gOt3E9/vsb9ULVpJBYZ7Jrjvv6SjcSfJ7d1xlK0ywoZkEuWqstXA1UOEqv
oJVliLEHaVs9yNrIPmGwvSCFAveT7SHs0Q6Fh+xHCkzNDEKl1DHbM8Zke00vKptG9WrwBMlBz0Gf
CkIVCzbtPnIz+3vJmDhZsSfwK1gOSmK8E2FmdSb2nxr5YKb/gcsuXkwwwKfilB0eT2sPiCiR+dYD
qt3gBIOP4l208b6ERAPyJd0cTldaxpmXkPkD+h0lpAjsBSCyrzdHkXMWAMWbANWzBvWTthf6TGhL
NB7+tIYPhU4dDfzRIUIAECI3sW30D1mTjlOEedh8Rrpr4DnYRcXfPQgnN79eIjM5aDfSgUS9/fx4
xe4Tja3LqiT03sTdajwG0rGRtBGJwM5740eAQqMUjk3L9im9VBH28c0YOJay8jT57vnRY7hhzEq5
mFtgSDCvkKQXiSB184kJh8xugtwij+NFFHGgovGP04yNLxc7SbLLnOCDVDzTpCRv/hlo/IzqffT7
jwfFnn/8Sd9rm2cfFoxvChFKTow9QsmHyocXLWKo23dIhPb+ZFuoTKyinYrpF3mras5QHW8+9NDB
fZNy2JNvIZ9rnfbDSGNqkjM/XgVIhkJnRvYEqUbUjfyaXBa2Z+FnQ43DWBEXUTjJhYRKeQZV8tIr
Um4vaFvgyjRtGHlBA4GJh+V0WIGaRnuzn2m05Pa/zqjIl/uOXrafeBEVT66sNGQXPwkVOdb07lQS
z9CX+4OFdkle0GpFX8qSoZw4w//jMtW+pTdD/Bz+MZG/2vlvHmtrB6vtkI0dEqjDebGfEa0mhY9W
tTknRvpcXR2/RSO7GDM8RsaMVd1cU1gQQthW2ypIWDiph6lq5wrvdOLkJnHAScrmLq4pWXvuZO01
lYVghmF6QtoOlZkxz80Vwyt89HYHNV6v/6UbcVxb+C/QLmAk1D2umVwx849t4VCnBDv37IlBFkRw
3aL0pL/l+05qNdLWGWNSEFsq6pB13uEMEpQKxz2269iod3Ic1R5KPoN8cC2lthCy1Eo8HpDi4JYB
IbTmaePabINTuQDqVbboU6h9Cu+9EuVVWdcERkZ5s3vzUk5OsjmWqyYtzn+ZyjpBCxTVHZO4axzI
kF7Rp/bSVF6eBzfoG6+5CU6etktYEQWEC9Ch9XM+ir0ATv2hmoj2ItVZzITeGP2pJaAXRPAHtFlH
VAoYx+3ahM1YMt/7RQTkIhZAdTh28M8ORYZ+RBWYvxl7JrTTfBFSm3fzc5iTraMQdgkHHrbA8qTr
HLyb4fZ7zPFDV57Qm6l/HfI2LCgECxvIu/46NyVf8ZxxRjAUrACJe6E6gtGNIQuy39i9FZE75SxI
/+cOTjrGsmdeSW8Ljqv2fog0/cgE2qzOhoyHaVdE7TqXXVSJ/6I0/5GPfnwdZG6DEdTtvtseCL2I
MwBdi0/Ea0IQKk97WddC6mCphTUieh4uB6paM+QSAMpG3iZZpLVSQx4CzQCGXECG0x7y92EimWTN
KJ3WZRq9TzN/5/+qsaH/fZRttEEzy5F8fkhX/moDHrJh6Jg0IS0jRrnIaTFBOZEEJH+2INOBHvSs
GN+PD0MDRCqmDG0Ha/+BtuwClP9/VGE3YEqeR4ZOMNsQ3CEwdQtbS6tGw063nUJfJDHH4JoWtDU4
hrh0KePla3aJv7G0oz2tvB73U+NU847pNknDUEuS8dO9FG6bXTv9FHYup/yh3V9u3lbDbRFJaLEm
+FcsPHc5/taHJYt/DV5qt+s1cRzUAoJSu4NbEV7w000NOe8N9kXtcrjgXGENiG+aY5ulNXH75kzd
/xcqvAKQEgsLTaT1bpz3Sy7+6rZnjkwp3v8GyeXOwG9Lrfy2kM63QKo5QxQESCPT5FjC9JhL1Viz
n2PZM7ocT+aqgikNt5q8320jslg6sYliXeh/Z6gs7DcyA0EaADGeO9hd14LUotzCS1Y4+lWwFQ/t
GyTDm9evz0Ys5fI2c0OBlTSDVmFR7kkum6+TngilvO/KZm8kQqfRcA9wTUgFkycscam9/XMGCTsU
BBkM3tEbOMBLcngFZfDwjk2SYM6MMv3bLtZKq/GC7MWNbogAPDcSkOnM523Q6tRG+d0iwa0buT+E
v5YpkDnaA4Hi0YENTCq2lBnVkETfqph3q2MXuna6yOU8SSrXAbDOwXmNXc/fkRYshqwuPoFdl7N/
8EodEQKqqpfZox+3ZsXsjHAYa8nCfdaT5e3FNJGWJXL7phV+m4g9kBPuXf7OJd5zgmyPe4+qp27E
mrNYzbIgJPbi1oySEWXuS3BEKABmiOc7cASXaMDE8e2deF3XStTVA41irtqOQdftgGUDuH3qCtu/
MUgLRbl5OLVTubh68Eh2voRv6x10IimVFs66K/flu7O1YoUtYnPs8Mk9GWKB3vjFwTPietnmnAJP
u1Hjxf02sHuZTBxYUNnJKeS9OJ3s+qUxWjjWdmCBxXN5HvMsatgFil1/aI6fFjhqLXuN4Nsyg3l/
Y+mo5t5Cf/9cyE6mqqes++9LDfVR+aURlkoOOn5nYjynbNFtzA0zhNeeSrbhory0lnTbGjzpscu9
TgCzc3HM56o6T4gtFoQ5cLFf7VEthzqBzEsz6035V6TMJqMYaqP0oxnSnJNsUPZoMGboeDJSWvG9
3piveOVI9Hxbdf81Rb4iksXMzv2wNSfiBu3MN97BojqQMsVsDadEDhCPgcW+W/5lCRUUYyk5zDUa
W71qXD6PDnigwy3UKpUnONSEw/buYEAl+TevKI+IbPapUMOnrGVVgNXvlWT0NbFw9wX/ThJO1oVy
0Tuv9WPZNSV5f/h+3RdMwgI8KL/mS7c5dsRMWZ5MZouZi+2UYWmXfBD1LROLyERb0ApJe36gydbz
qiZZt4O3nASAWPCvhTnQhesbEhdRTbAELpv2h9LZnxlfgPPrToMT5lfqoJKuYAfieS+EXZGNHJVg
9N1Vpx60AR3dkmcWrE8S1o4NDmeG05CtMZkjqbmVoBRKQI5xH3O/wqAkdHDtipt2YNMhaAtILk9s
80ccM8hpcVRLMm3AwNrPcYngdlnt1d6dx+KCeX2DqNZ6J7sFcUtg/eaXEXMifBS7Sd2QDgRmk4Qa
+79z76l+QHJ5t8kPoY4oOgUn0zFNECSXq2H7UBevksJiQxXCq/PFCnluSwtYAw5wtZnzJwyuHrim
jGj/2r5biIDE5XhfQ7yGtWiWpmxpk5QkvHoOiIGudnhB1JK0DpKU74JsDqW40XclnGB1oKZG0jlu
ZQYNECDxOLi2VcZ63mQ+bhh8kp9UaRUp8hqUEjyUFjNA+ghnuiGL00D+QAspMlvZf1mhQfFD3GIF
LbQmFTqTaiABMPeln0ZiCLtWAB/55vHY0kYLgPey238dR+eEPWHdbLzh6DzAdQ40lEU/Up8L5Ayi
ZA+eDjqDQIsLTzWW/k+DRpx7d2gadcU76xGKKx0091a5SZEinnawaVDGYVXsDvd48lcCiacYFjzc
GXp9LPRljIggBgvDcu0gUKCzKAFK8OGXesuQJzaf58ZEiB60ceaWcnNEqM5dtt/agqkrs2BmMpfU
+nl55CUuPB2PXeCGYQl6rI9rf7JzgKl7g1DIXo/Z5MnCT8OkoQGxQI3+rtCRghqjDAtrdZY+a9oo
06rM+1Gx/BhTQy9U7pb7lwMR3GYsrSPk3HuaXQTH4ZCxE4u/gliQ9mH5KDVuPGiRz2GkSkTWR2Ek
zwVpSSMlJV4LBSSiQdJ3GrZaP6t8WZ34DUP1fwsom5ninB2EFo9mVBZAZRs1wb72YMQsibKFThTM
PCSdFUSgtvBFRGrojvQqQS70q9AbFbrIuIXtUfUgzCFbGr9fLaVMkSEwQ6cPKyb7HnAjBpLfvZql
RuuQKi85doE8W7VGrUBtPqr3eSEaQ2t36xPpx4olEkxeUKLje912+45rk9200pqp7nL0oQDFJV3z
YW9tXQ96jQ7K0g+IUJhX9jC+55K40MmSS0X5y+OJO942Dx34mhT27b4RebnAY4JPcDZ1P/sFRfRp
RB+eDa81JvFKuQM1zoZ96xWU/7Qb+F220jp5LL9QNp9pq42EWzospRsQtbmu+1z6UWeBbyGBGowW
Dgyi6J7wqM6lwgDSADivPygUc+QEwYCO3JpOjUrzmBo/Xay351ENq4neL5qn4+phUCWcmt2yqLiV
NgXmWwXAddweEm9O+XGDUnLLD54yqJdnqQ06H5GBPW3wqLL7Ltg3pVQYEHprHkvlEgIJ405sUJpE
pR+c8QAcWvtkUcjydExE9ru+BJaExYpDHKx6uy8TaVS0RVZ05/Ve+OHqYN8kiunGNCKwBdKYa40B
uZaam+eVUeCTaBVoRZWLi3hbzIN1+TNWbcjrz0ReB13KDwQImuZxlfGyp94bQUquoz26GrMj4BHV
tTnUxTiKXzjLXNqjD5shI427xDh7vVjT6Df9RPPavUCW4MeC0iStGZIge0Dsb+BLnav9dX3q2JGf
cKK2s2479OSSAM5s8a25SsaVvjXzqhqvmt0EpPsb4HplLpS57U28EJ9zUrUi6LA6rZdoOS0EY8ts
5fq27sF41llr4JU8gjZf593aZF98Ij/U/B0Kh4ZBQF8ieGwOUV5+wLHFw+zWXTdMbPFLcS4g/CSn
k5qXyp7vkNvF9OU/5qhZj90lO27kWfACkq63cFYFYyN/Wsn6sY1MgG2+i3CbxYQyrLvz8uFqaiS8
dQ3nhpgEQ6UKP7RFeq6eA8kRNcjdDmscsyHahgfA4XVVHNvkpJkbq01dOasfDg2lB72r1RRekfZQ
eUpXdj2OFR3PsXqj+Uog8DWw+W3ZVniB2ETUPv/pCMMufcdEEJGpUYEQh9/SyZ5A0haZKj5CEVoG
/Lg/M1RzXvuXXjswq6ykidXY/SFCoUddtzH+rlRwdTEuK3DoY2GkhhVGEYpGoiu6ONNH3PRRbtv0
JDkWQrGq4JQ3qVFmVFyKKvI2TKxN/VYbAXyBxE25fHaE0QrQQWtjDPxE049w1/ho5F2TEIYk9flV
MRBplfu4ZSvKGWHO6mrPpb42cCDS+ia6HkO1cvgqseOKK377H/KO12dm7rzVve758+MTDCgqcWac
QL7R9kU5wDhuNwtuhZEc+fA22Kq0YAIxbixHhsyAIlCCkaBp6vpdWIjIAGqJm7pigGnwpI/Rpke1
EJuve6kFHMZn03F1TxfQ5N5DsFKKAr/Vyg7GZ5bTVT8GMz4Fe4dhn/L9ckEZ7uKC4uzfHN9t8lWZ
rjYME80kVizZmwh8IVZSDZB/OZhGLixEl4jO7yWQyTO3JdlsctEonBpjkkzq9OyjogzrZ53y+M4A
GsrGVu+GxEvIVXbwCkyeF2vkVDoXBRRE7yr0Y8XDFVN4beICJE2VtmSFnTVR2hZg84ahek7iFO3g
bM0FPYIibvce0LHFlg2jgAOb78fujlhRa22EzvWc81insApyIV03/AF28Vobq+S+/Q0bKIcNXWRL
cXlkcgrEW1/hJ5Z6C1ZY/tViNi5B9TWvkNP6mP1/D3yumHli4exXvp3VDi+0iPSLS4UvkXmTa860
PFSTdXgWmF0oXxCKLh8CP7ACZ7q2WW+bqGPIBNmXlJXIe6w0RcDau/KPLyR5CircKd6C3AnbJwtc
l0TFFnI2kD+J0VLhl0+iF1exguAtZZ/LgJbPLGMsDQeTVrEalEtGUxmJlOuTmFkbLa3X/fUWA5No
MAAVlUL5nUqOOquBxPgKzgCKp41z0GCioLA/PVqi2EoxS/RCDMLd3o6hgxRTNn3sHJZLrgNyMAIy
4ZKwOhB1gYMFuYrjj9pV0muNmVCLMj/9DNKVbq3bGI/VIDwtaGCJz80q3xB9dRdQnnTh5OBY4bUg
8M27NviBiY86N6e2+eOpqRv2+2FXb9hzA3+KdawkMZT6KRrBiQLtPFRy7Z4wa2cW3I6kI8oFu43R
W/98U8iBE1yftF434unuCwAP9S7RpcMPsX4vVIwDOi+y7xTwQTwZw+AAHAuHdoP7cZMOTEcnY5x3
3Nx0D+6BU9qEkjSTMGKncUXCgLqGjrPEzcz8/j8qUdffGSQL1SFY3D2ntDhBgnEBsm/gF8VcDebM
UJiTzSNztbjKrRi0eiMxrCH+Ek7wfDENrDfQ217RvKs82K8zIqPWZSC0ctzOHxP3g/DalGmM+i0t
MKYq3J5koYORnzKoo9lACIh+lZJ3Q1r3MuZHQV8hhGmzFJaPPvgwdcpwBJ7Lu92gQHsnkRXlKlv/
dMSOvo9NuxXcCCLLocZBGaqyzpyWRsjMDWef/44VSKpqfe+Jg9YgSNYbD03Ae4JlHPBmRyIdFiXy
YcqmL4+HTJixxMlvAWxN9kwFLOX8u6hLP+x5J05LFhoBFf61+g3J2UW33ax08IeekLcKnV59/1on
3Hd9ndFX0AKe9d+kHLKGjN05NrWxi1xE+l0buP2lTS9QZ0fSNSiBRpthlrvAvXF6oFYBapmch602
GnllLRgX36MxAv7Ww89oYKy3Xl0pORSvCVQ7YEGDbVpz0BFnbB8tPoA7zfdsyzvWrPDu+mNrDs/o
mSKM2UG+1+zgS70bet3syKCKXMpknIZCDL82EysUIQTXC6Dr5RbcTUKjuHH18e2eSxNABTql3rH9
QzXrWf9DtduaJq9HWUkin8yLOJMhffLZ18AZfeqKcbL+Mylto7sGa5frynGRnAzE73Nw/oR/PT/i
8K49JOgAiijOUMzYrkYTJ0C7wKBnQSOQse0WJiElUJS6s8I0GeuK0rmw3i7iJs7AQMOUJNX9q0KG
ME+thYERMBf/h6RX10NNmcNMeuNfDbpzCW/0zPCxrMJFk4uBgj0v+s37cBeHzq5guy7L51Fc61r0
uF7wv3K36XH0pyBI9K1KWHaXhZVdVK6FNDcmibE0MV7NIF+2Odh9zryoXyDZ+RScrzzZygKT0DnP
EwjZw4E09wl+lMnETJroNWTrS1LQ8aj4IjfPt0dmqvWyZKO0OnDF828HwE04kXPsUBQJzPyoNmUk
3MoJ8ZmLhK/ZsN7sGWCvnl39NHCBlUGdDU7MEoRPEAY3s9vDPoMr4wWen8h2rhReusaXG7dpiDR5
BmOA9hVfQNLkoYhHalvHfTEk8xWzHkI5NLQiaxBY2MXuk1qnMft/UGm9bCV8BATPo6hvaKOfLiQ9
+t+rh+BqMIUYINXvormgUDWtcB3ksGLc9i7zeLgSuAW2z4LBzshz0IOJ8rgsHLgS8/FERP9Eb6Pg
VdKDdFTYXOYie9zNhiPLn/6Q0Q04/uYijTpdi/+UwFrle6DSHZnmCWAhywL5e+zDQv0aCGCRQYDz
3LLDEEtz+KnBJM1XoDd+6uRW8zUhjSLUkiPslLhN1L1wcmohjFVDY/Lsjbpc7lwiMtFuknSa1TVu
dEuaevLqiqc2sHl1CykCaWzWXnq38nJPYpgnQRHPxdTcgNzILZFjlAdE0DKDhOr/Vww79Kp7UBlt
cfuQqy1duMkU7PbGsSOJ9RGn9E/uRsIezZ7g2A9PPSMcsBv4PafdrlYT+8fGMPZzxdHuvYR1nFBc
UZHbdtb05sLAP1wrrAbuLkT95GjGOD75UiDbN2HbbXICzFfuCUpT/VEIEJyP0UJTRVtmFev0xHBO
2TfOBQ+ZOcYlmgTzyL503s9/b3wuk5itl43vS4Rp+zDM75vmokzeM1oybPl91MA+/xkyqbC6ww58
lyy/DoUfzCRlaRehaJkSvy0jjf59nxj1u7k9s6MkBNwPB5Zq7vPq+OR/C8Aeyjhs4t0n+vrShZuB
06aRGE+MNYGGk8ToBao/bH7gfX7CeQfSB0V5YzegZHOHxISpUPL9Os5tf0yH4Gdvqzgt9dkF8aTo
jaSiIjb+m1Bj4TVjFNZGzohRgDwZw9yKC3NrP5GT7nbG0Y3A+GoC7M1l8kaiHNQj0tuDz1E9A2jj
Upzj5rjpV/19qWcphDTv1K/QUZOG3/nGe7wUHEV4Syyqrnik/3QRy2LqbzCBQZrf8Y8jbxBl6ild
4yoKL1O/c1DTnDy04D3qq9BwN/qqE8lDluOlh52I/6EjEQw9O7f08WbnrUgH5hmNXKlQn+e1HgTs
FY8r/wFQIwvUzzh1OeZ3yrq7QSk3WJQUUyyM7g+r2btLxr8w0owRBe4TmzIOtZ2FbqN/yjQfs1NE
3gWHcWXue/bWKMJo4AIVFp7s0NFVvSLpFfOD4uyebbRE+oARuYY2FFu4B4HYDYgdWDDFV8xV9X4l
ANLbrhvSL8eVw0DdgTxeUe4QyGg08pKvzPxGzK17T6vpYLkymqux3QxQIU77IWRfgfiX9GzusY7t
T+rYZrlkJECQ6cKy2QBZCvi8fUkVgsv/ppvVwa8dldmBquXZzbDbBZV1mtzQvazIQemc3IeXcENp
l6R4dNTR4n1q3AMMH30G3OCddpcMenmvMk0dk+2Wx4IPUy1Dy6KoUev/feTnR4sWyC53ycRbVC06
VC+9hegM51G1a7vegEfZq+V+WdujrJKI3NJ/24+5AwCHwvvc5l9MtVsWlJ+pvPx42CSjBjeLv+lT
fH3KKr5MVV6lsVhbJwrxH5Ef/eKDN/s7lcHEcgcpeZrx0ZR7B4PnaNBRGrt25jDsbpLdcgbwlmRw
OhyWrkDLV72WfHiU5ABUscwGpYQtvBgePNtEK5DMkejVo+ZjVr0fd9LrT5Kw+w8zNK0QQqNo2Bac
ESodDQPraEREXewDHSin9B+dANpJRBNUWmulXaRVResXmb4JQX97p73OPT6e7AylDV56Yc0dqpyt
5LShkGCxD+IpSUA/2J3Kemcwv/7alACgJQpHQlFLGP2FjD717lFepEJcX7GA/trC6PdCu12yKWdF
ZJiTrevebrXT74LbGj2BlSL+ZeVyfe61s6ZC63BZgObeJeVc/tfAID5EYGT0nSfGHGQ71JQF2W/J
wU4AJ8eM/c51X6Qjn97nuyuw7e1H0HkJIhIy8o2/o1iL2I9l/m+0rB+QPM1sbx1BgcnEayO6nMf6
n4Xa9QQawYldS5a6Wp+7Cp4VqzOTeMevtl/tGZX0Qeie9rCQBB7DZeqJQYRa4jLtQtrzPCYziWPN
AK6xRvvEIkQKragqOPRtuggYfpyUJ/K23VdVuz5S523KdL3ETwBn8RYpqGcMaHI5Bzu90WKIjh2G
buu8xsBxXprn3j77GVFDyrI+qjd+DfXOk6NTqFr+Bm8qAAdUW3LgJYCxNmyTA++ieQwOhDyOxYTX
xAQmfP5BElajJ1SqQKga8lxlE0XVTOcA9ZsGlfiP9kEbQQhmeZhwufaXa5eW7cUhqVDe9nP15ZhT
cVTiHgn4AsYJ7Esb0I/Bkfc2tPjD4F9ld3Tpdxj3xKHcS8IzyQOZ2nOjMKnzJZZHYL4Bw42ligBa
TlFVewXM1kP8dKVIxT0CTZCOVDRUI5rddpVWqwKSLkL0zzu4lWGFjscAxROe3Pjp51dY7S1LNE8L
a+ks/rpunufCGHJYKtvxemUTTCs+1VLpuNvXuHc8xM+vjktvl3w/WEA0tQhABPuWwgLGZK+g6Nbi
2cO49z+JGS6BJkRI5oqSHnzFiLxML2KJFR8XwVp5I/JGkDqXFssvS1gqV1Pnhlng2vCsqcUb715q
SXqpKtUoqGrOpWliWpH3hY0UY/qcSS/O1M1VNzwgaRIUagTTdaFY0PP/eA3OjTVayFhuQafJGY6l
lhFrnIYrxA55AR1bF78WT+FMd9iycvxI9B4fcauqEEyuiErchCU/8mZ9dDQCkTW1k+KGlF5Zzc7i
cZVFJcddienAKnfM21q/qAx+LWQ64DSK4sehAgStpVQQIqHlPvzixl1xG93aH+XWaPobHtgBgiil
mSHqt5q2pi9Ufu+BEiaYFp9PrDrjZELizYb+abq9cxt9dVCRvwkN4pLwwcjqDIFJtF5hBjSLBnPz
zPl+NrSCnyMN9c5qcI+vYLAs8oobQSQhDeZQvgsoAKtzJFuiqBV9jf07Hq0icom7LhgbiF9AxYGX
m28xlasyDi2vhm2NVGxcfWX+hVT4O/SvXKy3nywmUmNu2GPPciFjUt9Nhcv1OXCJVzibFu7i5e89
ifktBPLB4BpmuaSVmwsGO+uUUvmWHZ5mOaZYeBrW6ZoU01p290I3GESgxjxXuL4CK7EXEObF0Z1S
GVAZSyZ772EpWr8XqWwdXSYomyH1Y4+ZfXmtBm6Aikt2GC/2jrm02qzapnZS9blO7PYYmne6HEdq
uSbWYaLA1WWBJNyAqBthHr0k817yQSXvmN64i/zEVobzClwpKrx7Py6Qgbz4C9axkaGhdymhQhel
XGDJ5LnoCC/sq6WkwC3XIdbDI+B/GFKepsMPf7NQNlhv0bvQ2ZjX1sUx9aqjxOtaAHxzP1a/yfAe
s9Gm27oJULj9moCXAlubpxS4WJ7m+/2prXCEN5DKLOWk8aSNjf1Hz7hjwC3/5DvfxhIpyILeudS/
MAmRkq3AagZVDiyM5OgCI9Kto9lmxeMSc+Ots+uAMHKyTZP6pQ9NqVNrjF5zlJHzK1b79iRiceku
wBS0PBPmXLcSRs7/hi7CzxX0tFO1HOgCWGG7dSil+nKJT0zU1Oq6slOWWoc5yjwqikdy85wuzT3b
Ql7gmGV4+wOvJ6ZLej4JUpOaiu4Yd6LO6zFnygOs2Ca6TxvZ0doT4S0jNafoAMp5+obB27+4MIRA
qNKzr6JSeMrcGa7AeZp5zfbn/pD8Cu8gokuixGvxi3KK4LDm3pwaZqexqwzeGVKkgioeEdV8w0oS
RWIeWZO6ExZhlIGLBswE6m91OOSxJuhI1Fw99OL/uW+UzCS/gDlJCKY0JOUyYBmHGn53WpL8OInu
pCK8l3eObgSRv7EoQYPK+vzPXoTDds5d8Lt+cm1GsUe4pGihBVLgYoDlcK97nEsu2KunZFinpWW7
4tbB4ydss/vPvf09KWfUtiF/7EkaoFF9oZTP++X46Ot0FxnWOtSpe2gu96kYg3Wo7VnrG4i57jrk
pQuZyk0xKKhjsXzll3xKKyEUp+jvSXgE/uQr7hPFWj602uk0t1fYsCwv6q9m24WdQ44GWxraeWOq
j7tPCHKOnnG6Ftz/aYIbg/ZkMoMdZ5fR/rqr0c1TlkcyCpU56E+hoAEZKEqrvIlOwT/Cee+x+8vD
eLkIpSdbHQku7m5l056UdSUHsyuXkfNAABO94uuwvDEWRY4+HNZ+gz+YV4hRcLd+qFIYU5xKgnJI
2KMg/Ck9MrAS4twiPzexOgia+UnPYIBl12WuA1Ba2w/Mbu/CyL3sqe1/3VomYjRCTD6VhaBmMsbo
HEyxFk/ktWcoaJYhH2i9SrfgZqpUKDZUfKp0eR9wfkt4xX70kb74WArXri0U0BTpCvMLaZuuG5/T
LV5ybPMWFwGULKyPMrXGD2yRmjCAF6fStj+QcKrVMIUeUq2FJmCPgCs1WKc6wFEzuHUt6KJ8a75z
3HK744vBSOBhNBxj/RZOh/QhY4cSjGPVzv0AExIRZujOKn5d5O2WQBmqkm0BP7Y5dXNcyLu242t+
GpYr4LlgU7Qy3d8FSXfFRf/lM/dFcOmiMuTaAeZoJjPHuPFlv08F0cXgmZKEqRR4LMsPEp8KzQi1
OFvWkOhi4nih9sEB1C8HarRbHzRYfA1CZ9w0L5sXIRrK3mbv88pvANiEUju0xUlQrWqkZSMgSF7s
Y5CjrGXru129Zpez/dmVNFijXsujafplYaRjABJ82CNYxJUPhhUx70klqm8/FTmkCJ0olojVNLrG
QCFn8LdTIIDvV6WWOCOlSHW+j3W+gR0hNCHcjuqugfS4xYV27/HDQBTDWmdQLp9ang9a3vkEjyp7
9KDtSE8kCJYw4suWssBu7f1eda1lAQRNkdQjyDHKyermKp+Yi9NTLVSAEVuBpUKpOJTotfWA/rOe
03k1AsthZvxaYGh+AmYGMxvztXuDNhixmvVhg8PrwfXLeaYy3HtmOZYXEsPqMJHKGRbP3TbF0Djc
kbKX8pAgbb3JMTIKa2JjSlGAN15DZ0Rv3LcMzM4ey9kKai0KeiQekVFdsSuhmdUQVVkOODgC7sR4
nltxa7e3eYvM+Lx0Dh2pp9MsnpLlJgTYBqoE/53HpbTZEc/0nLGBbWOZ8aYinWO8omEcZbV8XFJB
MZ8TxC3uKAhEWNDRFZTzsuwRiEhK4sCBebwWx+KO480SS+0v8XpLOFA0d/N/1H4lS3uL95gSMB6c
5x2YWk+IQPZe8Zjep7vrwb+KzLgtiVr7khQraf2LrdS716l3pgc5LB3AXOu+xmIlQc4dF9aqduxa
nqOTVXG3Yk0701fJj9yFLKpNyqWL3ql000AKmfmRkHSDC+QYtmdB/ujWy62WIhptY7z/aLXdxCE6
UtS0xsxXcTEMnpE15R1MGxsh7oH2wpQznIcAlT/jIct3JeHT5NPX0pjqrgZGGO1whYxAk045Di2I
DgCcMqdEwjA6TgXGogdmiQt7yyQ4+cvIvRDdRrGUPg8idT23fBmcLVZ4QWba0TuxCg4ktk1Qkx9W
cCzuOCQhLOyQjl3eKHiUpPShCtwtYpXlp2r4J9YI1zi9qjhZfwZ+Q2svW7BzAEELqL2Dtxm7e4YB
Ul1ThLt2vup88k75QIzNIp0WhUEIAQlmuR1xp67lIiXfdmC5+9LgAVtUMzVGU3tn3e0niG4HSOFD
ZUxRDgyfRuUBL8NDz49TsEtlIwttVdkwlCdiJN9XtIx1JUfuuCiO3fCSBr1tWfi/egWgqPNsipKr
C/LAD9Z1xBEu0KxD5+208AmBHdlu4jSHZqN1ZctqZ3kl60egmxbWColYx7M6RWhKglj0OAL0ARyc
3glMK8JR2IsSznujzGt1LGrc4d0fxk4j/bQWJ5VPkyALOkiFr/lAMJshtQy6DAzfdQKnvKYjb7Q+
v6/PwjrSyDCqXJra3NoAop9ITjGjzkbRZM0DRFix6LYncSbqGerLaPulRJwP58FSUvd/EtZ3mjSX
F4vsmOZexJThpVyqEgoZND4tDl+jBeC1raI6FitHXos96TRj5m1XAGCuVIe62JgrsKsb+lsOeyyr
r+GkIGuWbpDobkjnh1pDDGA8v+F1CU0fI9DLkSp39aJ8eg1LGdUd81Jdf07Qi8ec1bqmiKklFXjj
VVFItOcY/Y4q/yAvOhtbmynKkKkPORdO8uU+eeS5rYzEcQEAeY9Xb+AoF8wzyJZ5yll10F5u8Mc0
WW+PVys80FCvIqzaE8o0wrnuwwbGxq2rd/kgQU3jET1MURF8CNAuoMrRigt+aVQB1du+yQ1nYg0v
aaF9b7v+HWh/eY23B97A7TWsmcpC2JErUlYper8TJ+QIeWoO12NELQi/gokO26/qeBDB+vvSDgjl
lUQTThRcBl34SPaj08BmsD7UKsGDlzK6Dd1MWTuA0jDSN0/HOu1AddknrqznDa9gbGStHaIYpOT0
TrNSr8/6teV4XRceJJXWP5GRXH/QOux4/x/WIprnur6ZeuLIchMeDaicFxrH7brWrtRvPjKLlOgu
D7yu69fJKsZsQcxS2vQ/ic7uRFfDDEieG3QXD4j3dFVbPpOBwyVWZZQ/gdp6zSSPTfYiXFY4P/xy
5xnziJy0wd1f0WC+avdMNkQ0DuZxPyhw3C45Mg2YxFbQw7pen+QzSXpMbTX+rKt2UTEMKQYF2WdE
F3FVS8swqXpNUYFH+0XBWbwS3YzjJs4P9hCoiozDs6ZlUrIOPEKhI1KdvwSnhjweqkABPtWF75V8
VIX8FsouU9QozggjmmiXJyEYcol79lKM3Bcj1SE7G1IUog0GFFEqDaHj/SnQ1lao69LVbbDF9K3O
X+Gz+1Qhh7dXnV249CoNEoEsWWyHgPv6SnoJlwcozNQpkVjwT3ltqw9NvY3Gbdu1wNMpE4qrA5o0
7YFXzfqM+AFGvhrcqCzQuO+iz1ANRts2A40ZGerBLv669S3yd6y9gFU0TJ1XfTKAqsRveijTpHQx
l7K5cXO1drT2Z301ebyGYZwBngcXPnLmIwHYVRWpfJKBWo65n7gzdCvdEymsZUboHiKGKi2Fkxnk
wEES1g8IYXBnBqPr0yVHP0KypS1TEKOId1t1pmUjpO1EetV056b+h4o/6z+b/h5lo6kofVZAzm7y
U0mXXdigRXckuYFvjJpTi1ybYhn/29PVNc3tzUH/N8YTYUD2CYMO+DizHfSn6noDLdPI4EIBFFfW
e3xatgDvyy17BdEvr/jZ5o8CEYLk1kO/f0drDWU5/jweAxfPSImmU1hKZkgphjmI5LM/KwCqsNAR
fo4CwIpk5j+GR00YGvxsTc0LQIvRwKLFPLYpcbf/G1TUW45v1yvijXzDU/Qz39nlhu5EjdvyH9Us
FqvKtgmZKcl1o7c3wuf+tpuwnM6DuNa9N/EjBTznmQm5251enrMaGUwG1UioRGsbDWixdF/vFloC
4g9QaBVzPTDJiKzyMdd88Rwv8TZTR1cU91dHVsCfjPyWmej0J5ZYBPq02GucUfn3CeuV1uwR3NII
DXMAzdFVTjAdm3Gxppb9Ix2xeLqK23Y7ZomO9zffm3R+La4EGMTlsDL63vCd5ZzXJKbrBLOh4dhv
RJBab7tw/r9OUsN+CIUd32QBqr4cINK0T60aGkK82jaaVWlEMlyz0DaJ4Ad96cdAnZq9udg5UYqx
S5ARKwzhIGDeQXL9PE0Zy+pOI1Zi82b8HnIRlJnEdYVI1eblsolW2Df4sSdCidvkqxo71zr40e/D
ezA8Nx3eqSUXJ2zUmKZeL0Efi/nb8gEknlFbM/cKiBGNOQdvmLWfWworhWQIc4K3jMh96VutsrYs
hOimfipNWD8jR9u4tzdicsitc3+WSgzQmG8DsDDm6uO2xCFp8J2I5Iz9kt5lMF+l4XsTZklVOGS3
CRtE+uQSp4kCDaucJI4eKHaoEiXcr+pl+z0PmwWfhmIZClWw/sBvKDM1tMQ5yHHFViOYPMzCn7K/
HU1Hk85RY+pn3OHBB1rs5xMks0Bk0DR+xu/pN0hCmBjo5o+tCP2X32zfccyCTCzsQEyAiVL5RpPL
vZyK8xPwEe3V9UM2bijVs2rjsJEKACX/7xfznOE15SiEffTCWKBNw07K2uwXWgeJg1r04LrqLPq1
i3fi8LjyAjMvE3ChoDHv/GMZQCCVP0r4Jjjfyy6QyC4iKB+C4Yc3B21uKLYTH2tOMHwBpjMYsQxa
zZ2ntV16Bz6T4+f9Ow0pL4pYB3z/RCUb2b1izT+z6RpSdGy/UFc4jW6sA4yi/4qOUcS2pSBxQnJq
2R6BjKqvgjbmx5CwUXOG0SZj8BXBXgE2fUd4TecDCYphe0MqLtLB3JcLj99fWH0a4peFHa0QWspb
+YZPU5ycWZAgW63cCpigP75oR5+06tIyVJtS7JGdqWGgUh/0oUY8ol9RGFlMhXNpkkjTtf+7bhO5
0LfWHfMHYvis24cISxe36eI+ZoAGS87tSHCCaO8bmbAYKjLNmeGx3JAogY9SEeeTKR+GBspTo0oJ
5TS7+nu1yNURnoOe08sk8UhQU60FUNNVPBg1ER8vo1r553VKjivjSzQqTPW2Lxp7cfNdhEEpTOP9
a4/Q7dySuv3cOC4kq8Eti7T4P5ZGtEsqY2bwx99kDFwn8yHHvPYXWLTxcRchyO/GvqS1aDgYtwte
I3gmMrbd7PSDje29Jr0uCdRakwSl7GjTA02TJ/3brOj4n7JS61pRsD76aFYX68UWz09PW+O0IkoK
cR5eVCW98dEoP3SAVUW3ba/9bD7hba2C76bwyN8LqhN4M0QLGUnOrcq9pBJChI2XrINQRI6sdfLV
vRH0ZgH5XgmlE1a0N6WWcuCZ13j1ZL8lwyduwq2xpV+pkGwuvjeiXsGBUc5vil2d1LebE2hGeJHE
XLVIVmYFoqR1ZTp08iDG4LcMTJ3muoA/IvMDOGgNf7KfD1yhRzzre+GbmKv0GaR0NVvtGjoh/f8W
g9cfzPsR6yXO9i7pv4/SxBHwFKsBz5/TW7O67dUbZBS50qfjvevyegyzsWQL8JGKcCLODj7qaTSN
+s2nnTUcUdtl4RO7ktZFZqaunhsQ21G6qpxRjMEkQavlYXtDrisYPsabO3I8rapbVkD/vXgZg0nT
OtBFF49Y1Tsmk4Qd/S+1ld7fqF8cVTYyeU1Lb8Ghv/Y9hS3OdyTsixlq4ElyXNvaRXUM9QIxEIXP
xz0yRmT/PzqT5qPTZwKR3Qr4XpbLRdkJDVfUu9+ISlW8PkSnW3dUhXdy3euGWIy9D8s8LyN0hswP
aMSYGS/3UVbNEy6yCWdLo1H4KCJ/LgcFI0JDuGyy7dpbk1nDXgXv5lmlI4Wtn7qLNcbQIC25XT9U
peRNej5CPhiq0S3KyzLkMMvjwaWx5akbH03VhisUMjMZA2QgVMv52/CDChNKZZginxMYn2JSRRFC
7na6JxssJX645sNrs5V8u7qYxz0o1FkaoFH709VLiXxi/yxN5nPlZh2prnA9MxmgibGTJ6Vi5lH/
KZuMrSsnmHM7PGathxNb01CZqGOVNddWlHVPzFU7ueyqlATyA51IfOudd8FmgGfVWhYXDjPwZCMW
esVxrRGbJUmL5hFuta4rm4j1S1xYfGhmSGNzv2UlZI4sFFi6jgYaqJg8+k+TYMak9kaLHsRyQdQH
o7+Tk88+ZCyGulLKscv+V6o8dzfLaQEU7kwFPTc13i3M3yfc3JbrtDYP0lttcUcfLaLSDp5DgexO
UwgSmCvN3ksB07Wrl/uvaQ1lGdRXjJiQdZSbvZAIIhn2dc1f3GqirYOkl3BsrrDnYYV/UgfIH+K/
QIaYCXI4DbiBJXGybvwmxGLYH2cJ/+hEtYwQDwjjpj+lkbqPxhqnml6yHPCEPyDTVqbI6P5BSR5k
LybwCyBCGBhAkVzBUHGQObANo4f52nFwNYlqeD3Rkri1A3wqGdvdRG+jW04H+e07gvE84s+Y/mau
jiKkDWB1tubJFqjguXkp0IhzHk3CGL0xMQ3CTxnWVR9ddtNMO0Ih0eGvcriWXm+HzS8eJQSN72ay
HOqthNDMsEtJI+HgLo0Kfxe2vjXeoiDYqDLjLZemVHAbO+aMQWcYU1rzUCsBPN4bPLSs1xuU1J57
v2exM9DCf5pPhzCIARFC22nLGhoersAKuDTKPLI7SOrWwWGlqI55M7G85t3O2TnRYy2O7QEm/b60
ACTvh+Wm5Vkj6d7r78GB8t3thYwhYKfS7gd8T8ogQenWttJOXqHi
`protect end_protected
