��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$Rx�y�<��wA�*;�x���@�̦�W�X�fa�M-$u����n~�%���P�$��W��kYَ���P7�?UMfT��q�6�U��k�>����~�\N�(�����X�e���/6U|)�X2pF�]$h���d.���9E��WG��L�X"]�Ad����ľS���8od����e�GT?y	7�������ݵ�^��R�q^]�鍦�����s�ae���h��L��P_���ާ��YЭF���'\��68�b�[����w8�[X��V�F�0͘3����q諵�uW� �h�u\V�?@��_6G�_�*�G���B�絉�f������[�G��U&�����~�F��AׯK1�`c��[<��FY���4I� �#�G��x[X�=�Q1��`��R>(�w����R�O�?����7�,(�H\�#h(W�EH=�������yq��Ѿ��aF����:�U~m<|��.��0=�P/���4ǆ���T(���'V��KWق�����<�1q;�����I��:�y@�HSK.�ݿ�Iu��g�o �=��Tg;������"���N���PRݖ�)Ú�gQ�x���*�ʠ�3�rkY1�B~�t_����GD �޶���6���ޯ2{ڸ��~��Z讋7/�_'��� ��?�!=7� �ܗZ�t�Kj���<ɼF3�W��չر�[�c�8)�&��7sW5=29��-jsڈе�߂&.�.��c��a8QA��1�Tk\Ǐ�Jq���ѥb#�[<�s�hpg==
�$�法���L⽱��#��3|�a}�D��V"�l��Y,݀�R��4���O)M���h�5��_�֠��-�������1�>_�l��lH�����n��a[�1{��l���F�KQe~��g'P��2AH|���s��A�,�N��N�Dcw#��X+�)���S�RnY�]��ᆧML;0�J�=��]ԫt�?�?��*�]cV����@ʞh�ut�me>|x�D{�Mmg��I��	�_Y�_�ڳ���ц"�gw��[���^�����is���`�6SÐ0���Yɣʝ��5���=�>��5w=�G����6�0o��3�Ƌ��`�ӹ����ȳ(@fYHd�m���0�
�����=�<:j��%�v}��}ܒq��߿CsC�6d�� ��!i��e
/�A��tYv�1��
]p�$]�34�U��u^HH�|+~_�Ī���Y����)Q���QD}� �k�+,X���D���s�
�v�/�֘�'
W��	׾�qJ��� �B�o�X^�r$4�=��e����`2ٲ~"8��k�:Z���$P;L^�1PBDg �R'�>��=�,;���B�J�;�	�h����?�4A���D��@!�J��݁��{�En�c�W}�8��PQ}Ӏ��_�� pt��.�H^uBSr<�������M꾐?��~˳�VSx�=1��������;��)*zp��|�9A� �a��U��	�9
R�i*>�	���ExXdxwGJ @�x8��>�:(6�����:��nXկF�a+5��'?
���ʱ���EP����h(���rŲ���\0EV�-����"^��|���g�[��9�R9q�s�'Ӻ��/�5�|�tMt�������r���(�
UFl�s�v�W,�H���%�y��g�i���®�xA�Ѫ���wPU</��/�*ʠ�l�4�s@��YP�}��_�B��d�pc�0M�9x����6p�E, �\����T��'/7��q�B&S���N�B�N��fl�5zqu]� �*j�Uߦ��F�n�C��/����5}PF���鎧у�t[��-�D��9LC9m(�_䦫�	Ýi^h�.���F+���+[꣓/�|x���ʵ>���[�_��ݯ��)�b\�?��	a�Q����6n�+g�u�a��B��֑���ÌR�V��p:#�)5���T�=N��L�3�����5�;�)\6�V=}ct�����̺�e8ț��*��+Z)ޜQVU���� #�0��+v>��ߏ�?��D'L1���d�լ(����ek�2|��/0�0����5�@�+�ݚM�G�{�10�trapr��/V�Tg�p�ߜ�bV�BiO-�+l�!O/*D5Y\�/�`v/N̫�x>��wI� ��3�-g	����A�3�'�DB�0ٮ�r��U�ߺ(�'�@G�WI����:���z�T�WN�����*P��*3����_�i��h5}�Y���̊t!�Q�D$i-�A#��5��#������)^:!׉�g%�m�~#�{��01�ZQD��.��pw�bK��Q�0l;F�H-���L�4�ꣿ��4����6�T�m���Ξ|1�dӠ�$��bo����n+dq�暋� x[>���
`u���<@�xJ��);9�>a=�&�鸼E�7/H3� ������"�X/y*G�jv}`1I��c��4�S��v(�f���jp�S`뾡D�H�I�J8B1���*c�J{wB� �u��s����(pg{;�r��1��`i3Ɉ�+y/�fv���%'v2�{�c��U�G9�+�{-d!�:k�,�3�^�n%�џ�#��F���;gT�Q���ֱ�)���?����	<gV���E����S��ri�68�Y��P��?M��PT��;��}p�8i^.��MF�/)Z�->���dDy�Z�~�iܫc�xN����0$�DI�@�ݜ�b&�s\���P"�H3��`#�-˯ ��l��� ��bӄM}��H?�����쭴qϝ��>��"2�P��,o6�����8T)*�����-4B��b�C���Ģ�E�ᗤ� c�&<O9P ����8�|::C]�J�l��v(D��j������,�BRB�u�%{�_�V��t�6�,���F� Q/�neU;����М�N��1�T��Z�ZfTO���ε�Y[��Fp�r.Q��Ӟ5$��L �G�ӗ���O����[�U<'�Hϱ( ����P���*��T���\�Ŵ�n%��e"[����R�)ԓaUM����7l��'�+�>3B�!��ܞ������d�0�YS��{c����\��C-2�y���~a��x;pfK�`����D�V+v���d0�H�JE��)�y����4j�0#�x��諆�$잱jY4Ǜ��U]N��t�ݭ�N��fD蝥i���p"��Ң�7�xB�^� ��h]O����E��`S�ݼD3�����	�aE;�Dc?!�j����D��%���ь�����"�$>�ܶ����w��+�_֤�������T�������a&���l�>{3���g��$�-��|v����{�\���`���������xw������<�w 7\���[��C��p'J����:�k���B��}�����T�Ī�n���a� Ԯ8�r{s7mO�F��@lKb!=����"̅iC2�6\���K�&�<��w`�#��W<�@k;���z2rn���W�	l�C�(f!�H��f���
�� ~� |`s^��y��R�);���z5;��*<Ԥ�..�|��Ȝ��R�<P�F������;��ڕ�����u� �̻^�L�ݜ[���J$�����o��8�s$!�&��B���4�O��?�6�>p_f�V�U�Dd��WlV�F]rQ�w�ԃ_ޯ�C�R��ՍI%c��v��Q5Oߎ���wu��?H</V��=)M�J�D�D��h9��Z�aw:I��w|�m�������w��\�AY�A���+!�C��U��ʋk:tE%�V,1fȔ��ձ{Z��a�_ó�C&#�Wy��J�]���6P�kus����O�TcQU3��q��R{���4%���䄊n��	�mrbp���^��4��Q���q��.��<ׅ��#�r=I������T�k�*`S��+,��1�]��ƶ�Z��%���v�֦&s	����s!�0t����������.e�N� �r�xTa:!�l}}h��ŗ�kXk����+��&�[i�	�o�� ��\�=(��M�ӃPB_Z����	&dy&u�A�lce�4f�x�{�pp gԹ;���v���p����w�ǒ��1U�Hv	
!T���Zb��[E��o�_9�ƃ������l�AX�&i����u7��|U�H"'���Պi�R$a ���I�\B�^vK��Ɠ�9P��� ��Ѐ]c316�k��+e����8��[���얚����$�G�p�4�*�5()p��p+���zƋ�!LS�}�|w�.
���Zt��!���>�k�ƚ�Ʀ*0"�Y�xY5�y����2Q��2@���t_�5���Eo�<;1V��^t�uLn,d��{����>��2�4fb��j��.�n�{��l;����蘞��7���'uS\��=��NV�1_�q%"���K�����j�t��l�ѢI4�"�y��bꬓ�)�������|~�
D�;�(o� ��W.k!ҿ�[f��r�]��HI�Ҍc|�k��8�0g>��2�&��S(	c�R5z�����IQ���f<�g^2��+�;n蛔�t����,��@����������G�7�oSO��[��hb�jp��w��<B�����Z�nqα��K�-��+�toކ�~v4�+���	3�0SK�Yw�N�°Z�:hw"S(�$�S�)n����to�s�_L���R���i �����O"7@Z�枅A�W.��Q�͊��e��1x�����	����:s��i���J&���9ט�\܄1^�y����~H���K.5S�8��ޫ��Mo؋�(R/�%�i�o�3�\_���<�s8k�����n�Ҁf�����)XNQ�y�cڗ���zyӒ� ��Q�*�
�d�౑4�|��~�O��i�5F����~�Ps����Kf�K�^�	�;E��|�Pr�	� O�*�C��tX�������q�ũT!1���C�i�Կ�F`��Ii���O韠��s�'��^���m\#��I($���x�v8�~+mF�:�\q#�d��wR��	f�P�w����Ѷ���y~F���w�|yO�C�O$R8�I�"�D��D�Ev#K^ֻ�;E0Ru�RR;|WD�l�>�������ô�	��s~,C�>��3ur�1��)��O���˒���j��j3�]��o7*���)W�q* ���R��X���>!�)Y��y��p��Z����Խ��3[�C�����%,�I(�����P�WWȦ&}�}��Ǚ��ִ� Ū�)�Ā���y�\"򪂸?�9�)J�K��'��mi��$�F��*��)j��LM���(4J���!��$������/ ��~o�L�"�~]VhY����$���&n�.�/ҩ>��[6E�(7�{��r�Ԫxܝ4u��
���>(�<S	�P���g/�4L=�殿+�&�S�󘱎��_*��a)�#�{��kD�]�� �����/�6:.�@��D��e�o��	 A�K@%yr;�)����z%�YM/{q8XAJ��rQ`�RCo,7���n}ܿ?U�\Zޣ��w�ĥ���s�]�u�9`�������z$q����$�a��b���<�Pn���`���c2HO(Q謆�`�H:���aE�~�gR�ywR��^�a�iL5����"L+)�J�f9r���e�qU�9�I�#b�9)�M�Z-^��וf�2%��b����u���H$.l�$!~\ҶQ�*���� ���ˮ� ĩ������H��QƐ���m�z�̚ko�o�Etԟ%4<a�7����s�&i��rlbQ��Vr��BM�~����V�����uz��U��kwذ�<%�)X7k��2���	�!�>L����M[��Q'�����#)&m�a���3R>,%?g̤,�X�AVԨ+w���i�]�*��4��ڿ.��qq��VCN�+̑���4;�r�
�g�۟���~1U&���3^|,���)���\�4����ϑz$Zl�72=[�p��5�feA���CHWz�Bxr��ˌo$�+�}����q�n2��%銘.���՚�&��Bi���gí� �E���6 T�明D�%�-N��?�̤Ie�U�	���0��s�h�����nY
o�Cg�y|�D�-m����AIW�b6~����ox��d)��68&e.�ȯ B�&��6t��(��'?��_˗��������I�[У] �P�"���_ZQ+g�~�Q������Q*�'���m
���K�P̯aQ}�t�m1� �>��
"k�LCUu�70��m�uh�I(�V�_���5��>�Y������u�~{[� ���@ 
l�M
���6.�h��v�g~uu�ϙmj[BEh��ޙk4����#M��m�T�I���L�����[dDSy�F�'�m�y G��;��SWMf��ߊ��l�'������8�b���<��� @9�6��BP&i��B�.�+V�݇�W�$h?���+��������y�������v�hΤ#��h�H�Z��"M�_n` (X��	�(-�o��l+��[˟2�ɝ����H%܋1䲈�@U?K��=�E�~+��k��L�P;�`��Y�%�_$R�骏2�͙мy��(��,d9��:�k/G�7���U�4�E���3.3,��E�k�����dؚ�vd�+R0��>Z�/�)�Z� �>��@K�ˎjI̘��`����z'���	��C��4�¾q3����W�g˺�4�>|�B�<�ה���Ѓ���Ze`��9O�\e����H�%HV�DP��SB���U)�Q�"��v��B���u��w�y܏1Y�HpΔ��S����OT��g<[/FH$�E��K?�|g/�y��fB�I�Q��	X`��K4�b��(��S>ANsB�zp5��P|��φT�#��ˣZ����@۰�D�o^�Uy�~d�`�ϊQ���:bB�u��i �W�Y�Ma�Qx�y|���%����/�DD����m��3�~|�����Ųp���s0��?�����}mL�"���P)Mݯ4羍�?��=�;�Jb�q���\�?��	�˾�t��d/�Jg��xmV:� а�?���CQp����e�PA� �2aD��aP�."����,�b����F�R�� �xR(��}U��^�����o�m�!�,g�h�z�Q�bj��IK��K2	<	��^r�1�J���Rv�?�klxn��r��`�+a=8��Oe%4��=pV�����"/)�#�gLf@"��t�@�4ώzh$O��_i�U�#�Æ���ޕ6��Ue���{o��Gv�|@����踇De�����9s�*�?���,r��`b����Ð��*�D����"I%
͌Y�(ZH�a!����-���^�Y�"��fQ=!]T]��*Z2�����P��Z���gZ�������g��x�с��ګQ��`y��n�=Ւ�E�(�+�VW���jvPp���)�m��c� �rN��Kex�~Z/��p�*tq�'A/�E@�N�ZYM�L1g��琉uν=ߴqG�r�9͑f�N#����o�*��>�浱�D���:��0��Z/���OT�[��I�s�#�_ݽ�YO��Zɺ��V�ڻ��f�d�ň��p'!V�]s��g \t��餞�s���Bc#�<mSk���l�"�ϟ��\�03��B����@C���ӯ��&���A���'0�f�6�]�&��{d���gmG�e�kF#w<P��M�U�8X/���}C�V�4�t�q$L߻���ZkyE�*q��\����j���%R�~3�t+�Dƈ�F*	r��m@�k�6�Y�&�9U%( �<���]��- H�}�-��+��mEH��?h2
��p�i�8SWA{&f_@p?f9��!���S���c�o�Gnp����ZiGU��}�ɾ,�u��C���A�O��4~e��q��$-�`x�u�w�/���|��	�J���:��V#��U'������5��5����cA���v��eQM�?_Y��M_6cA�������]k���1���UN4���c齿;���J!��R�1^����ݪ�ˬ�b0���+ĂU�����]ģ�yh����6��d�-Ǳf�h}��Y?I����d��aR -WE�r|~�i�_��5�NA&Cm���(�츿]i�|4�����ĥ�W�N�n�S��NX��{O�>�����.}��� �Z�Ӯ$)
珲H�8\���,p'W�50se� ,�\����Kz��r���Fa���Իb7pҨ��Z�o_Y��˳���s@�O-[Tw�G@<�!<fRi��8`��Bo~�*S�[�.gX�@7�q�0ܑ�&�Z�Ɛ,ª>c�r߳-��JS����p!���D0Q"&(�z�ʿ��Fx�f	m6��:��
��ؔO Q+��G�?CCx���˼����)x��)p�_PD�8O��YP����ޖ��ʔ�-�֪�@���Rg�2�\!��j�b:�Hg��[�-x���������`Ξr�#o�g�m�8��B����n{���Y��&K��,Q}�X�����((�6�5�ur*zD��G�g�y�-'�d4p�?wP�����`�j�"�b�di�V��B����%U�S��%��#GIo6�6oE�J}:Q����82M: �.MU*,��(.��\�I�����&�������73�vX{�q!��8I�DG�;��g�ۘ>a�)4x����|K]�Z�il�/�ɳu�gO ���j8ݘQ�w�E�H�"�R̋V	�����!<#0ܬz��c=��L�|�$����|?�N�C�m�E�}��G^[�Q a����z�2��ֵ봋d���N!y�YA�^�x��ީN�G��;�!A�������l��QPR�����tҕk����m
�Z��V$9ǚ�B�H�4@����=oY{���l@��KCk2��4ht���6���4K���&�}v ��b��jt�C.�)��u�H����ZO�5�qDzX�<��qΞyF�ѽ@�]��[���;����'7�H�=-%UY|X�.9! �Zu�g�mYw�4:T(oK�<�y�6���C�_Ƶ��b���Kz�[�t>8;$�W��0�Z����V"K9g�=�M���8��OU�_aG�"�"6����TP��o�!���jk!��͎*'���� �BQ:i�w�0^�p�.�aMI,�~�h4��\�9�|ơP��:T>�s�*w� 3MT���]�/�������ܱ5|F�R@$���y쿍�F^"i�͒I
�x��}�qD��\�1`G�IENS,�~qiEM�[Ū�����Wa°�`ښ��+��'��^�1O������ؘ=�.�Q�f�����9]xh׿"��غ�"[٬���e,]ʫ
��P^��D��g���6�`^�!Y�%',%yӚ�>}hb�L�J�nH�H���ce~W�<0Ri���Z�"-��}s���)Q*ǌϋ�6�u^�<w����?g@�w��Xnt1�pÓ׊C�N4T�X["I���Kϝ���Q�J�4[���QxS��Fh,�M�ns%UG��o�w���J\�Ǻ�>Y�
u����}�Klz<�ƴwX"�F�,����l
�W�wۥ �Kn���Y
�wh%֎�,�f8B��VU�!y���a..&�����r���)4�L��G��1V�<ʞ߇cHQ��r5�!�oJ�y.�s��� ��g���c�h�y�d��7	G� $0�~�+�N�M� �̍�8�1znr��n�N
�xg�)��<�
c���������&K��`g��l�X�u0g�hr�^k���3���2���\J��̹�7?c�<�8�Y�Ic��U���Q����)������خ�
;�/�6�O[_�[G�#�X�{��K�ܶC�A�[̿E���d��8ݸ"�]U��$8��C���/���φ;�bFn�>$~���\o;�)�ϙ��1S(��Q��E<��ՙü|6�߆X��d,�jp���m��E�+�)i�ʊk��I2?���z��<����-�mƁT���r������A�\�p�+�����I��1�O]�uY����yҏΓdC�PA<��g�T�	�p塟}E6��$���р����tr�+�<a%�}�S��q��#B�e-+\����^���D�Y���9�bXנ�l�.{�����h�F5l�_�8��W���G�n��Ē:�/S��.g0��Q� ���V;����Fs�P4�>{�%X	[��q���u���lv��WZ�xB�f7�np���{rؾLGat!ԩ�|������S��",���]|��9H��C�<Ί�Pkxmh��1A�)dKD$�R�UBS!�fnL<w~�[�b%3r쨎�v;h�3�(e~�h���Y�漽4�jXi��ד�٬)���I%S$/&�������В˜8��*rԄ	)�H3Q�s�y5i�S_�ך��Y~c�춏S���r�r}v6�Y�a�iO�v+8Np��wI����ص4*�+�[oq�t
���w�����`����W�|^�pQɳ�K����͆a�Qm�%�kVH�:�(��`�׵+�'+�W(�{��	^�P
�z�J���=�C��<7�N�Y {g���>�>W?�M�?����������d+���S*�j��\�Y�f�����
�dj}���Ϯ�����,M�M�x!�p���#��.Vg���T(T��^y�9�I�)8c֥���+��z��k�19��bB2��s؟��4/�z�:ײ+��R���x���v2mzӟVx4m	�F]i�Jp�'��1�M�ŀ���N��oD3i����@��i.!�1w�r���y�Nz*��SɝKa��c��G?ԙ�� �"������;FkdON(ŉf�7�Ei��� ���䑕7��DE #��|�Cx�*�3ޜ�?!�[��,�>�,�8��`B>i���g���(C�%!mق!?��R�Z��l荤�򣓬 _o�)U�%��Ch������F�����[�Ӣ�[ѷ��:�A�[��ɿC�|p�9��dD��~��l�g�<��"�߶X��raBk̓!@�CdQ^
���.��^��g'�,�q|��z^��`Q@/ڃQI�Iyڄ�s�!��+a(�7��94�B��"L�D��&{ȴ�,qu�a؆���j�݁�zG������;2츃��{�G��P�¶���w�^�L�������"	���bYj�»)�	� �o@�%���*$Ο�=�Etz����N�����5�7A�i�1οs*z2d�'8,:�@!�f������1���$�3
SHIsy� k��x��|!<+�⑀�����?(��F� (8�]�^�����9㨘yb1�7�ȁ�T���F��#뱭`�m(,8;�텧_���>�/�i5y�),�t���
������~�P��������Z�I���}Cѵ۷��!��M������: ���()}��@p1�۝�ӡ�L����kT&�n���ۈ���g�ع��'\/9sr���X|����+Ӛ`�y�5/���F��U̾����!6���n�d
�h}f�o'�d��U�]�	�M����1J�o��k��?�
���,,^��;��(�d��ܬe[?�i�Y5��/�q�s�����ν�P���1�:N~�J�b*"e!i�����n��k.�PYk�����nN���06t+����ڦ�E�tҦ�W��}s�Y;�;l[Dڊ��zY}Ә�H1�K��'>�4���j����9y�hH-�<�,}�śы�Jh=A��'�B�})�8Z�H�4������tu̷��g�%Ϙ0��C�N�E�TQ,�U���X��4��T�oA�����4k�vbFͿ��,{��9�|�3�/�侇���
����Y��mv�k�oo���oOz��"x�K2���ۇ��3$ؿ���I�V��`��#�r�/nܯ���@)UNl�@L��E�ծ�WO��ȡ�I�r��ю�&'�)����s�]n#��L�[=c��<>��$�4�H����y� `]�2�0AU�}�@��Av=Q>D��+0����=�L��rS����9�-}��D���t��$��,*�Y�^��~Yf��m�Ù�ӻ�p-�4�-���x&�V	�l$@5`d(q꒎n�\S:��M�~˘(�rO��C��>5U��̪�����n��N���t��)�n�똯t1�m���N�s�$�z�i�,�I����\ʖu��;Ń7��φ��lM)#@��8l��,p�T�Pͭk�b[���z�i>�V�K����£����p��!Zn�=�ߜ� 5�sW�:)��f�}m��k�I9Oz�魦�i�}6����$/�a�k���|u(�%ר����kc��H,k@˫+/%�J,~1��S�<�A��(�]��o�����PR����Н� �5���QQ.����R���o��)|��6�>'eE�ɳq��S��
u��Nh�@3���oo���p��d��>�_޶˿W�ߘw,��*��W���v�7clregUAsY��|#pt%���.���-��)cm�QX�C�.tWy+�ū��Γ�z�K�<���y�/�/�YhwD��r�
��l⛽t��;١
,Gy_�'��"��Ӭ=Ԯ'L8r$788��Lm��r"�I��<]�U��
�f�V����j�	+$!S[�U������*�9c/��rI7�*����3��e�9c��T�k��EE]@/���f�)G��7=]L�mIf�R�v��$E���i�~�g�0���p���a����f�s�e7d 6�kI7�ѿ������,������y)���� �=���I8ɠ�::�:\EH;ņL�,����X�	�(�ǪQ�U�8�4*��2���j�w�
 )U�y*&�G�N+�E����^Sj����/!��eY��*u���1�bS���8]���r�O���x��o�4�Y�{��A�J��(V.M9 ��Y���'��0�Q�4sz���<-��G�}G�	����il��j�?�[�<I	�J7�O�+�ɶ�*��Z`ǆ�#!��#��h��y�߼�.̠�^����[Y~���e؁�H����}/?���!W�
6��a���� _ꓑ�o��4�c�K;�s�3'��gm�D�~~og�_��b�JIʌ;�ݕ����HC�Z����TI��>:K�dV��W�$A汵�ച-	~(S�@'!�����*Iv��Ŕ�7�kILY�b���&��=���Z:��7~�\����n���D�9(�C4�c[-���+�.q�ُl�Q;�f��M��ǳ����Gę�3�w�#��jm�;�����h���LpA�����F���)�X
�,������͸�:J��y-�y:�G@�/�!�x�=gO��oXy�(]��%xȏCmC#����8��#)h�u��b���ޟŕE/G����cvl3�e�}��kQJ]���N�/��z+zK&���%<q��K`mĭ��.�y݁*�&᫔��k�ߞ�����@O�e�JQ��}W�YdtZf06y_��Kf��+u�x��$H�kk��`�@�џ��]�=`A�����tZ���)=[��݇�}w���MY�u˘�q�]`�oE[8X��`c���_�{M�G]^�t1|��)Ehv@��z}���_��A_�~w�5N�>ֻh1II��w��P�R�.���B�Tߓ���v�Z�7k"�L��?m��r�����?
����:��X<"�tKW\�3����,��%-��SGB
�^T?�葿�G����Pz�÷��ҾηF�/9[i�P�G�z)�l�[�c❼���&`��{���O����c��;u���c��n���� � ?5w����J
Ծ��dïzջh��6�.u�*�<�'#��K�����m�e�Bߋ�65$e�m�����0F��������"�ם��ޡ�8�.c�����6�q���c�xZ�K�����O���a��\d��:1z`i�"�_~���w޳�����E�!7��K�����Q��.���\�t������r��?���-`ɏ��j�
F�h{�`�+_�Th�PE�yp�]�VlGCfme�=�˼w��i�Qұn��3�3ã��'�:�R	@5�eL�oVT�~�'�t�dgR��O�����Q��+?�)nsHWBPz��_B��m��v*T�e���(a��$����&[y������U�1�c$aKm��p*����Ż #�/�l1�]z0|8-f����W��ŏ����*��[�;w�0m��:�o�o��O�� ,T�˒��3x��!�/��Ui;��ǁ�s�);�6�)H���2.:@���y'��Q��кȸ���w��oߴb�ơ��܅�����#3��k&}�¡I]�5�2c(�ޘ��z�uub�)��ie@%G?�"G�2;�$�іPUɃk���&��lJ\��g9��`b��	~
���ϋ}[�H!x����jnpx�5�yZ� F�G?���8��D׋����Z�s�S.9����7��1j���-�ۮQ�4��۸2��
�}�ݭѨZ���[�gM4a�$�e�l�T�(��tq۳�I���/�n�YP��N�+�$��*&�46��#:x0�*Tߏ|�8M,���田H�gSE+��P��3��8� S {V@I>����Yn�	�4zv�p�j&���T��&�U�=��EPBT�F��ox��\��6� Э��բ�![���-y�\��TD�<ߴ�Dq<���3��ز}��[j�)��l��!|���Q��Kp}I�C�d6��t�KFx�f�i)Tf��b�R�H��Vf��8�
�:����������9�I���l�M�܀��a��mс����(�G{t,JD�[�ȏ��pX������.̭:�.�-�$]{7}ì�B���;���-|49�S~
�"P�b�� �QJ𢷸݁����/����L������x\�C�~���[�9+,�_.Y���\�r��߳�P�s��%���V�Q��0�b�Nt5�"�$�|uMsc�}ӏqmv��(?W`鮁��S]P=����Aܐ�[�y�V����Dt=sǩ��K$���+"��xl]�֩�"J�z�� �4b�����7Y��'g���jv?����yĖ�xΞ�g~}K�2w�\��5B>eU��J#@6g��v�:�!_	80�q|��o��h��L��vm�h�y]����bU��G�x�ٶOF�0�k�H[�:�T#�L^c<��R����7қn"&1O�wr�$M��Ch��Q�KK��"Dۨ�5��1�|^����-�ͭ4yz!�L�%����h�R��. �]?��+�sY�`�jJ>��QLU���ִ�)�#5�^/)x��UD�;��^<4O�#/��5��ȿt��'��E���(�F������ogÂ��U�Mq�Bŗm7�v�!�����_Q��y����G,Fċ��v��T���@�gc6/�E<���01G�rQ�r?`WN�JnSۻ�L����7��gӠ~^��Ĵ]pf:�"��D�k�i�Pg����֌7�����{�mrO ��/��b�C�'�`оR(��c�+�k��h��n����el�4�7�O�#l����J���d��a5�{yKX<p���`J���	2 sZ�|��+��0����v���dХ��0��f����i���ێ7}7�"�& N�Ib�j�ǉx��� ���~�a.�hcm��<��Q<�)��'g#��DZN@Xh*'.-�/J(�{Q�2���w�7ܲ5s �ӌ)+f$�ey���x�
�
�^��:�X,�Z�Ї�7����$������atס�?���|ؽG�l�ۧo��[����!����d�}*���	8pA>�u^5#�'%!�V>e'M�!ڬ�~o���M�F0���I�����}FY�st�V]�?k�1�G:e<���Yy\%��Y��D��|a0=���>
��m5Y�x�!y*3B�e�y��f5�Fp��)Z.Vӳx2~*qAߥ~Lz�
i�\vi�L�}���6�0�3��f��_vxn��[Tʹ��G�BǾ��N�#M��Xa��7nO,��7_~	�M�glQ�Ъ�A�.��Z�����ΧK��;�PC���n���
��E5��������S���>����*x������C�^*���I���-2����W���+�ٰ
x�z�@mi������75;���Ĭt�k$��KL��iQ��bߺ���`�)��[�[RYIlg�ߙ�rO�Y��(I���B4D��E��5�xM��_.K G�`϶��Af�I�N��C�lL�o���F8�x����)���R�ݯ�� ��ȥ����)̇[�a�A(�b����1�O��-�4���3B:�C��]S��xx.b��˻��p��O�
��7o�N:oU�v�CZ^��x/ia_*�=�!P�'�bv0^�Y����) �4�"��c���8�	b�X_)�8��#�mU��[l�2&��AS/�?�`1��E�MG��#�M��*�@�W�������f��y���{��}�?Ց6��q�&
2�,?��
�C�m�g��P �� ��s������qH�Ň��:3��g���p�������
q >�O�덀\P�m��ӱ���L
�!�_�4*��?��sW��8�I2]�8&j�8IÆf��fB��c�YZ���J�ٗ�+89��}<�"|LR)�?7zg���J�M�?������=HmĿ�Vz�FB�^ ���pR-L�ΫL�x�~*u޺�o�]�9�i��qї9S��F�S�L�� (��Xcb�E^���'��'���M��]�BmK���̽SW��6�a0�|���������&��/nm���Z��Ւ!���_#�7݇_����d���o�ǧ��B��w"��+���t�?u�aΠxdK�����6Z%+گ��Gv�y���?��r�~]��%�0�a]U�:n��w�$�g��
��>��a�a~�% �*G��y��;2_�b9���o�u��~׭�X��3_��FMRpς^i�ODM��G�� N�ۑ2~�8�������o2���3��K����*��Ls� 2�>'%���ٞ|�� P%�'��En�#���������>��7�.ケ/�l?�H�.�f��Bn\�L��W���
4X�9�0��CNe:V��:��@	�ɗ$_xdG�����ka˯>`�Ә�i����b�i�u���J4�w6�>�ט0�-/��+H�S[��Z9b�(��FAf���c����E^�����P�i.w��F���9��k�e�4:��t!� >˗�E^�r> �f��BX��#�&3�Y�	�m􅉊̰�uby��v��=��w�8+߹��1��l��JFE1}�~�΢�ǨT���}���E����|�Mv<�y?"}9f��'Egd
:3�ҨW���2{>W�}At{��;���M�=Fބ Qa,~ �yͫ25."H3�޶�Ȉ����mf���{)]<����5P���!�oN�th)0V��*���"���#��r���;�RˍcL�_��C�� ϶BLH�%�_�ٴ\����#�2Mg�����T��w����/P�RY4m��н���˰%�T/�D�D�0��I�r�-�cU\�5�șD�erV�����T3�H{��2��:��� ��gxM	��
5[�ݢ4)��N�F������z��e���y�$�&sN�h�FY���d�Q.Og��w��0� ^�� ΄!��B�׊��s �Ed��Hu�똏��:�tj���u�C�-�U��������$�g�W!Y�����@oR�ǫ�{_p��vסϽwIU�\�>�/��O"�Z�}�7�1��j����=�|�yӂ�] Bhd��L/`�J�<$�U�7����6.���u��7�fѤ�{rxI�b��2W�uv�T[�1����-R��K6Q���ӈJ��7*�1��x
	���5z:�Y��N�0�>���<�Vg�w�yVL '��X�gkGl5���X/�4U�=��~��~x~,|f�7��f5EJ9��Rã��Go!�/�;#픹U�M����h�=j�~ۼ�!�`�`x$l�3����Mw�r/`�����J�U>��
�&�p�40��koi����Ӹ�X!��j��ȿzY>P^ޘa􄣶#1���x%)~a��3��An+b,��	<�B=��G�8�4���\��˱�ޒs1!E��_���AU
`?֗�n]��#� (�*���K<I��  +�iqr��n���*ܪ�|
A�m[)5p�J����g�4�����gE�	H�����S�9w��e�bW{V��A1��0_b������G&���ѻ:����1B�N�����(`���E!��t�n)� ���E�����VO+��2��J���:)h^U���ix��5,-��]��	l�̓��Bg�s�V]G�85��ݓ�׶HoA�<}���8^�i&���[�1r�����)��%�(�8����:P U���%iۤ4���
��n�r6y�$�Cm�b�P=<�Z�w�NYu8�ap�QxЊx˧�L+\�.6]��t�N��b�*�3vW�$�����|I"���~l�\k'�`���`���i��#�^BGLH.!)8�kV��a�0K��1��H�,(x)�p�=�'���;�4�p��&o�C�jVZ�#mC�~��X7��'�/|%��V$����S���E�SY��$,vşSޤF��Y[/��h��y�7��Q'����m����Kpk;7ȧ<�ʣV���Z$!Q������!��nƐ蒛Ë�
S�0��u(��:�B@tt���JT,l���k�[������G�zT���X^#��S�%/B�_�σ��Ja8i�9�ҧ�uʰ6#W�j�yl�9�%�`i��hr�x����,X���ckE���oІ�/�۟p`#��Q�E�h6���f�R�SL4\`X��U tXf tw*�,��~��4<~v�i �M:��3�M"��LY�J��:�mWlz]��������n|�E���[��W[%�"D�A9j�����H��W1�;C���D;�d�_��(ẫv�9��\�Aա�Bւ����@�ˀC�Us�b�����`��<��ü{�(���8��F���js������A�<_�-�)��Cئ�r�&%'�l����(h?͏\�KDe�@4Ob�I4��	�#Qմ5���C�ʂ�vg��phV��6o����j	"_�#SJ�L{g1�jP�,J��R���q,����k@�͋|�j�D��r�s���-���+*�b�E{��G�l���0I�_֙]�jAw� ��=�I�HY-�l>L�⋧;��\�%�U�?Y���օ��x~@ax�U��ĊR�;Mxݯ-���E�xE���?�\�b�zۧ
�<�V��-%v{u�j�8`����,�o��w��KA9t%���Y�QD������N#���D��8��z��#��-a��ë0>�;G�AE"C��|�B�٬Vҏ����v�V#�ãuȱ(�N.��a�1�G�}�r����c��x;�m�x��w�p��g�.��VS��I��|�7��G���}����zk�����؆d���ef��&o #c$���jT�1q��7n�Q�Pt�;d؏u�hU�V�Ijb�R����<��~,QM��r�;�~����8Dob�볍�S��5��x �� �>���v�ۜ.Y�J:�I�����3�f ]u�� ���"��p�� y�ta�#�Q�*��=��F~1?�Fَ��Rd�R1�������RV�
)�S;�iq��1)Q�"�� f�$�v,�p�l�G�p�9���(���D��� �����{x75`�(FG�FM$��3{���^�|gWʕ���|�ߟq�	]Z�妛m�$G;���#��jÐ{2��)3t��}*?���ff�{k񛭆SxL���ԏK�b����e{�DHo�!G=I��w L j�F�d#�|��aZ����b����M�����q(�o������
���M�x����^�'	C��ҷ��Fn��~�6ڳ��E�M�x�l��[��%>�b�VN�}����z�Q���ۋ���eg�L'���Dk.R|���88�~��	D;EVIu2�E>>�l��F'_��R^�\{��� "g�'=�����gf��bJ���G81-�����Yw?
-���$�3�S"��h`��ꂀ���K���A$�}H��,��.W�����N��'��h�Wx:�?�c�{��YGD�g���������o߸��6�&k*�=��"��?׏}Os~|��(��>�I�An߆�[�d���!P=�C��|&o�ڈ�7ёO3H���(�[L3o?�K���h½Z���7v�Yd�C5�M=�z#����}�yy��y�U����;�}�>,��|�*��Q��O��"?/C�w�M�<f�����?���!��O�IMݑ�ij�:�i���e�u���L���I�jBu����/V��?~�t�.@�|:�Dɒ���Cq>�rl&AC����"x���k�W�v�b�g�������.�Hi��б6���u��
"U��hNe�U����n����ļ���hÝDΓ}x5�)���$�f�$��?��0y���iX�~3JGfH^�`�X�\�V����������$>{��w�t��/%���b`�ɷX�S�b�B�����e�����*���O�M��MݾR;���^�o3�?��{��y*���W~�/|w��[ഛ_=u\B#�f�T�J�+��A�M��z��xA��S��Fsf��ݟ�[�:�Lb�`n]�R�ۀ��w����qC�L�E� ��X o���m�G����d�������+ {�O�J�en��l`��p�R�/�6�s�\e��=�ץ�"\�0����*���2A�����w�j=�w�����\�n�s� �����*�oB ��d�g��<��B�{�s��OʭM_fwe^�nԶ���S�d��=�E8`+&6z�o��.:N�4)JV�He�'m��#�+��a�٠�9�3�)ycp&:I�ve�P����kiO��_���AJ
{K�A/���Gj�|z�r1}a����B�4��n����=%T��/cK��q	X��u�
Xk�dֈ�������%�\�q�>~�1T�YY>	���^���㊰�w�����np��*~:{Je_Pi]I+;�-mC�9���wf '�ͰM!���U��*\"�ZΛ�v{x��>�f�3>Ae�U��1�{�BU�����"�m�jԡ��F��7���pD��A{38��yHW���)eÛI��5�+��(4��['���#آ.�x��~6)u^��v}�U�?���~�^��q*��!pu�q<s���t��6n��0�2ed&��=�?�8�L�@��,ĦV�+L8�J{œ�r�J�H�ΐ]������e� '}w֕9�\��0��MkW�}B&H��V��V����.(M^��j~Y����x��9`�Ig��ג����ަ�f�7��R���6�M��1|e�Ҫ}'?!Opt�+������4��/t�G�r�as��X���f���U�Xh6 ����z�T�H�M n��c�>P�Ն��K�e��0����<hnu�w��8�; ��9�э��3�=��~�3�}�$I���+�k ��U�j�����v�]�AHz���o7ŧ�;�\�#����¨WPF��A��l�>d�u*<��ލ[C�J��.CrׯL�0��P!XS9&`2�H�D+7�;�2$�M��c�9t��h��"P@�8�5���-!������vS��'W�SRyq�#���s{�y��l5�Xd�����=Օс�wC��0�����	�R(���
'O�6&�>�g[y�ݐq9H���^QۀeL��@�Љ"��Q�+�!�Jw�\�R*�5�<w�/�'�L"�}:D2I|�\�������T���W�Q	" +�x��.d��cO��HԌ���T����;
wQ5,�}�l�
��!"űbe'���)�9p>
t�"�ƽ�>%��Ѕ�\r8+�7-�3EJk}���Ds�YJe��~�D1����(����F��L��.����Ph���2<��j>��Vuʳ��$�	�y��9��[�ï�>�$�t����%S �9W�W�7������ɚ���@�UR�v7s�=��*2�)A�U_$O�Q�� Z�H9�K�p��{�uD��v�7�m.�)�����X���x.�{�_��(MF��Y��"�YRJ�<��x��<BF��|��'�wPN��q��ǒf��ȶ\�� �3N���n4��g4˺?B���ܦ�"W��MFxvD������c`q)��kׇ'\�1fc������O����|���\��򰜲�f��i��3�{m2������/�5K=���i���`�I阎��R�Ը=ԏ@�/�+v!��΂  _Ne�?�4#�PճO���ؕ~��8ch��hᚈ��,? Y��c_�M�J�hL�
d2a}��t�ih��Y��"OM*�"�1Q��a8F��ba�b�֭��M���tF�t>Ɋ��/j�P<��(d����q���(X�ʾ���&�#�;�}PP��1�0�i���3�!�����O�:��Tsg�����o��8��\BTeK��1�s�����<kK����+�X��[��h�X���l7�z����FK��~�`�#djLy�h̃#��;3��s��~2��S7u;P��W�m�T@��N���5bf�M<��w��IJ/F��g�Koь�1`|re�X��s�����뎜���� �r���""���+�[Coq+�j6����l E����a���5K��N1�h�&n�&���<�0-�6NRx�1k��#@����0�Hh@�w��6*��g�E.28�L���F�Pͮ�K-��~��^H�"0@`F!��$���^\�����5 ��(l�y�3"���W�۔M5�֗o��S4�>�CYGu��:���y/fOX�7�(��c�c)������;��)�,�7l*��÷���
�,���F���������u��H.�hM�d��/��EB��?3����\��=}�6�Ρ���d>/�������L�po=a@��JSM{D��q��@���&�#RD"@QΝ F��F���DP���.I�~�'$�*��N�tnމE�N�)+���5g�Ɛg`��%l�<����״� ��}�+Gr=&�>`ȁȢ���)m5ʨ'�h��Dl�2q?����m��MT8I�\"�KrTN�1�Έ�e>�kf������ʮ$�?Wq�����%S��묙f�s��Yok3��Y��_x/RS�1�53Yݯ�H�Qf@5X5�k�*{�
���4X�<��� ��@��.���ͷD�����0M+�Rj��Y
2�|�,�R:[ͻWJDhog3EJt3�jj5��]/H����]���nRܳ� ��v���?u�}~N"��.V�Q����\(	��D��x!�e�u�mn�l�/��I��d?@��>m�w��%��O��>�	y����+�ց9Ό��L
2����~�\D�Ԑ�r���(��L�n�����0ۺ0x��_�0�p\��t+xaT��|�h>�O��EZpշ�#�,���n���u�b08�w�ic��cJ���t���l��N�ȳI!'�Y�7��wn2 kEcx ��f��eo����̿Z:z��7'�������j���e#��BA����t���@������&����r��=Ύu}�u��أ�z�U9<c��F�ԐL+�u3>w���8���E��]{&���LXQ7�oD���� �H�A��.�<l% �� n6�;	���	���u�W�h�i8Y����vN{,���H�0��u%���:�q�EW��V����^n��Ǒi��2%?�CC���'��a^�N+( �,lޱG%�*܎�̜�Po�T*R.�����~���~`er�Q�Oh<G�����uc���b4\鐇4H﨨jn�����$^��X���3:���ΛZt��(6��h������P�k
��;�H�j��N�0V�--�pE7u���Bt��U������w.0� �E5�����~��� s5�f�{=|�����X�5Qٕ�x�ŀ���M��UYr��ӤO�z̹���b\���:�P�%S.b�ff���2��]b��TV�+ ��Ə�]�;�J�8����o���d�z>�U��X�KRB�7����' �Mȡ-R��W�R���m��o_+�§{7zA���Qr`T�{����B�alQ�29"J�?�d����z0�a��s��飈[��KцX�۷n���M��#�)�{�N�I��^xm��C���_:y�hJ��J����=��/���4�����^P>7�/�%�AD�p�v��&&����d� -�|���o�(\o�x5�^�C�����G���~(���7��"�-��A�;,�6��a���K.+n�s�ۜ��1����>'uH��Wŕ�@3���l���!v�HE��ҙ�n�;�H�����n�&Ujb䴴Y,��ʄ�g���G��g68�l9ssi9_O�Qm��0y��}���f���Zؤ'�v��Nb<�����
�� ����`�E(����$-���鶍� T*%ggd��X���LOY[9�U�@������;p��C>��o��	��D��1�P>�K�����0�H�@9��?�)�N.����@a��6�*" �r�Ty�S*��@
a���]P�����g�����l��4 �l���>;Fp-U(*�?�u�¢�;���}��`�z�6�V	@����B�l���o7��],���R,� �ĎL��s�#� ���A��y�8�@Ϙ�A�[��nNzS��[�d��|�4��ϲ�HJ�Ę_.&՜e6��:h]� ��R�$ N�+���471�:�����7U����$򜕌;Y24��P��e�|FV0�(l�\�3@��?&]�7d9�v��ct?`��][Վ�zzʥw��`���������i<�2��b�(�n����u���A!���W�VƏ}�Z�#�T�W�BKn �*�<)F..�7C��!����V	�� �4�yx�Ef�[���N���1d��t,�X�1< �n�y�2 C�顔�L߇����Fd-xM����^�I�E�K���f��c��i��6���i�CP�x�����2�3�>1-���@t�:ך����� ��t�r��y���S�$G�7��]A�*�'(���؊�+-�/+r�� 5I�#�#��'P���g��b���*�w\���k�H3q/�pX�q(���~71�ƋB��U����^�]����k����C�i��ІG��`wł�?}�I{`�`!P吲)&�6Bǂ/�?����VYЭ���4��@3��xL�)9z<�	�/�2�V���<��I"FuDJ����L��������H�ϖ]RPK1Y�"?����CiA�����OcY�QȰ'�t\���"b*����c�A����޴c;kPm,p�>�!��˟��E�'?��;D����)���Ӹ�Ϫ0W��W�O|�Á���%ˇ�ԉY��ꔟ�Lc�}Y�&�2�l�u��5v�T}������$��8T[�C~A���ŪL��t'q�(<=���XZu�V�e��0�$5kZ�+��`��rm�����kLu�k�[h�6�ԧ��l����?��6�0�L���� �}��+�!1mv�ۑ�׾��v'91�y�ڥ:�aܖkF�.���`�#��2O#j꣏�^�2y�����'��y�5�zB [�q����t�]���U��%�.�@��t�9o L9�f��Ci�C�T��l;-�ݺ��Y&oJT�qL�	�����cTE�����g$%�9A4��nkp����,�4�~ �=p7��Z��mu�Lą(+���|��Ԣ����������.*�b�e��`ڋ�$V L��@p��9�[��C�X�o3���Z ����-�� �^�ǹ�)�22J�v�rVa���K�&	�ts6�lwX�L)g�f域IP6��P�>�W�gfn���6��:tݾ�S��z\A;���4G2������v��:"(�]��g���儊��2��e;5å����δ#��_��ip,���:�U<����0L����4c*����A�E�!�;NБ�U��5�*�Э\6 6�=g��)�*�d�N�6�ȏ��i�..ҫޖ�X"�r�p��_�d2 y!QOL��W�7N�?:Q���Jտ�wW���>�~��f
�Hۑ�n�q�Н�;�3��e�2���8M� �D,�e���!�5/rz���͕�1D7�{�8{�\��SM���̗^#{!q-�zׁ$����,��3�/,�`K��=�X�rJ�B�J�k��|�$��OK����	AV�jp�G��='�	��w;����Û�t�|H���o���Gvi�?����N�9�.Z��#n<v�rŖW(�X�LN��ڍ��m{���`	�*/Mc�ۛp���R��89R�sE����uI��� ���`.�/�7>pCDj�;��e���;�6��7����
���W�����{�'���k�R�Q��ʑ����U~E�S���!�'\I���tF��0���b��F�K�P���p��\o�bT��B�{� *Wl�(�}z86���o�ݏ�?�jIm���W��Ԓmn�Kﯫ����1C��>��q���6�C ��$6J�ِp��cmzM�w���@�t19UT�C�~@EM��66��a]]��Tvh�bZ�F9�Z�i����uU܄5��()�+Y¼t��ˉ`y�U���7�^O��;R;~S�?]0���Ww�w?tj)��ܱ	�>`��pMMC)���2���K%���s���xx
�	��ܾ5�K������;���+i<��@��Z��X�,T� w�5�Д�PW�n��|[���q˶����|B�R�$8��IY�Z�w˲����Rc�&�SF�͉dL��y\.�r�K��Q�X6D)��`9�`�����R���P�*�f�U �]r>k�Y�̠X�m��AwZ:� v�O��]�:UA?��k"�Q-��"��<�+� ���g$i��z�������įzl�T]��S�7M�r8aU�I�ß�8�qD����$0�x�on"��[&��,�=��=��"���t �@�^��Ä��9���$���2J�M��r�ۋ���zG
����oy���Ե_����U ��S��ݹ����ݧ�+�����?y{�Q���G"��A�>	�1b�a7��j�Is��J��*��ߌJ�~^'	��)tD����%�����5�4�����q��q�} �8>��5%�o�"�.�W�?`��d��~ ����o۞w.Xkߧ����k]*'�FbB�\քf������*�ʺ	���@�^�d^����$�����r!�����kN�Pw�Q��-�7>�;v��U��Ⱊ�m����zwCe�2bHSŊe�O0��B��׫d �^ �d8����,{�鴃����9b����򎼐�J�_3.��Hc���<��'�[�g�1�	&�Ђ]��[اv&�abmK5O��!��X�Z���YM���T����y�����!�T�s�rڌ�.�i�!��~=-td%��4�L-��P`�1ql�����t�C��Bc�����
��[����H���)]$�y\(�ÔYh��w"�JN{_���>4Z��y��={�;iE-$�T���^�����Dq������q�Us�r,I:�W��E=��i��/�ixp���МR�ۈ�����x�i�kƸ���J��t�WY��3�B�rJ�v&�v�Zf���{��^]١�"� ���ܠ�},H&�d
�m"vM�����l��vM|�`�L�
z:a5�}7�FQD$�+�u(G��q�v6\&�����^�]9��{@�x�9�b�v�����oӎ�������GSe��&䯝�ŋ����x��k��]�מ����O�M�,~\|X�:��7�&\9���^n}�*�o1u�)Q�2��YvQ%!�3����Y����B�?f�;0A8y����)��n���9�q�#Ln[&���r��	��ݴ��E(h�ܙ��k	��A�yv�V�8L%5b�B��(�@kEq����Q�F�G�p
'.x��kŕ�����/'��)���}죝Ռ������U[�+�$Tz��4�ߗ���x2�dh�V�7� !�?e�{��5ȕ�҆?�ոb+V3(׻ɪK0�#��x��Q�}R9߭��J2uPY��:a���FU XI~L�>��h�o��J�
��z<`Q}_�(po�g����|�x{�;Be�W��tu�t�D4�@V��	� �Y�E|�q�P���$�{0���j��D"˄teg��7��ɸ�8�f�������uɛ�B�1�+w�·s8X���-��3�ߣwA� �.�p�U��1�|7����j@\�p%��9~��FS����� fi���Z��w����d����Z�'e����PU[�%�e�X����y�6sY�������ː�x�D�|�y18�9�`�Q#���o����� �k�C"|����5���C��z�V�0j2��>�z랋�ڂ,;ql��Q��.�%0�5��A�-��p2?���Σ�w�T�=2(f >�K��5�LS-lV����4:D�vZ�����~D��p�D|��fL(uwQ5և�)Mܘ��~���i@��s�{љ݂��-y�\~B�6�O�p0cX����@��D'�etU�O&�P:S�~ �=�0���i#�IZŢ��B]����ٳՅ�S���@Fݐ����$>�S"�����Tց2�]`υ���Ue��W�t�9���b�RA�f�����}�q+�j-2Q�XZ�W���>��­�+ͽ����4����bSm�ػ�Yy[�����h`��ZCm�g/���l�/���������\q����h�f:��~bK�f�	����2�L,�jb���!���Uݢ�U_ j:��&��6�=dT"j3\j�gs͑�T��9�֬�Qp�Ʃ�9���a�sKϡf,zS�:2�P�ݲ��q�ġ���Y�&�6��1���<��;�zw0F�L��q�4�+K8LK!�f�z�	�x��k�e3�L���:}��ʖCИmMu����NMs�ȇ2 �A��.퓛���-U��q���ZWݤ��v�W�ӿ<j��NB:�:!i�fmmF]K��(Ǟv�\WW����'�h�Vul��.gg��>=o"dz���rT��GN��_�8M���sK��B�ЂD�&�	�O�@ܮid3V�tf�ڂ#i���a�l �#�+�S�[��΅?������Dh��)��&T1��5��N%7�o<��܎�'�i�T׿��@�m4W}��+��a�F��u�y8b�&i�$�����d��0��{�6`���B�r������p����T6ڼ�����<4��]������ >�!a�L7�y(�3�Rzz���r=��x�$&d�j��U�1<֙���8JNi����d�&��C��S.����h4=�~��,&�Z�2oҩ8)�cdpց}?b�|��7���r�[��_�Sb��&O��	U�D��4o�F�QR3��dD�X����4O������i&M��8�m�88�������F(�6��Q&" Z�<��P[���X����tLp:P�B����b�O����>��;9�1���YqW����kGU]$��d]~���;?�����[���&�r���j(�v2�A��H�o�d�*��F���S�Ҍ��
%*�o����ދ�m�F��	��� �Sl9D�\����+�P�=}� .��,Z�"�s5��J��7�!�Hm�T)u�%m�p��Od�q���!��%�]Pڭf�<�&�b�o�/��	}�\�_b�G��U�hS��v��oP_�#��r�s�w�	_�f,�I�bFHG}j����-QV�ڴ��MF���_�������uw���E�e@���ϩ��xG2��^���-Z��!�3��ޕ�LW4f�B4nU:���Y��襧�"�W��H��0o$D(s���b���n�&9�r�B���Q;$6�x�#Ō�=�E\���<�6_�<���4�u³��]��R4��Z�و-k�	ũ�r�y7"v��x�
 aW�Sf���nsa�SbMH4<k)��p]?k������L��i�<u���Y�Cb��+G����ږ���)�y��{Nc؞�8:���.��D��	��	�d(nz�F7�q�4�?+!���>*>U��$ Z�믓�lj/�K_�O�p�x��cT[�T��ݨ�e]Oȣ����pK�q�F����-l�y�lh��ri�<���!�Z�~��%�,,��ZKHy�s �5zM௠"a�{^J�������v�s:r
�M1��j~�?'Q��ܪ�k���ӈee�s������ ���M�dS��L�F1}O��d�ftgZ��MG*G&��/cKTKenct?�)�\[�����"�|���X�d��z��$����v�Mwg'�p�T��+���� 2���"OvpF X�y���w���V
E57|��0�����ʹIP4�I��߱�C���FQf��N鐐��c�Ƶ�U�)��@p�S�Màzà�q��P?2�:��"��I����6�tʥL���	�l�W���
>%m�a���M�^?d�t�]L�����->���ʡ�����<����̑�S5J��?��v��`��m}�w�Z�9Ċ�'�3�))[��PكQ�7Jj6�(vR��7�a�T�!u���&L�&�b��T�Aq�E�^V��J��p/_5y��&`0И�5�	�j�<z��=�qQL�Ab�S��v�B��8Us>*�jz˕-�|`����VKI
���=�K����_Ws/�e���l\*��͇f���2���+&��u��r_C��܇�l���E��08�&n��e������I��$o�w"fm_��)�R��^�Nc�P���hd��zĈ�5�>��X��">��%������C|�V�PYP3	��ک��h�S�H�
O`tt����ߝ�o�SA��!���J���W6痱v���^�s�!�m��������[���6�%pxE!��<��T2pٸO�Q*�����i/�{c���K�c7���A�J����ʯm�T���q,,0�r"��U?��U�Hϊ;�ޅ�z�~�vK��3�N��s�a��Nz�+���o�H�oV����]��`$fH�px$-���J*�ym��rb3��=\vTu�&GH��`{q��\f�ll�:P����M=�Tχ�e�1�=Fx�na�0
ܵ��
A�z:��i~����w(C�\���G��З\H8;�>��?`�vV'������J|�K�]��J�Ys�V�|���Rd�Թ��&��+��p�Y
�'o�ofW~&biJ�B��B�<�J�[�+�kǠ�W@�g	:lab�C��s+�i�[�'���Ų�+dd��v��!�Q�K#�fuA�m�P��=)p��^���y��C�3��Fܶؗ+�Ě�����f���{,�Qi�}BFD�0ۉVZ:FQ��c����h�=ռ�3��'�*��@XМ��fc];`H�F���^��+�-��TZ,�����I��Gf;dx�nG��x�i�;���x������+��-�t����4�&���wݙ�k�_�D�+[�����N�k��]@�!���}����e�kl%�yN]�.s��:�n�)Qɱ��EJ�d^���4`2\�J0�U^����eS�����H���� �,�"	�VJ$��`*��Zo�^�U����%Q�QӴ�u�T��n@JW��if����*{������ꭶ�aZ���@�x�j��=O��؅�;/�`p_��1�?��%x���}�)9G�Dٳ`��㙆i� ��x[֙��S3O��?����+F.90T��j����Y�(j9�&^��W�����0����yc{�0l�;U�?Q���/�n� �&s��l��2���&�V�u%;��u�����d��_�Xww���Y�C�1-�f��Qm��{_����*�uB�� ���^)FX4u�
>&���%���%U�k�h�=xKWY�Ҙv���\��T�4�vh?E_���p�}4��a�����J/��2�Kߓ�
����}f�&�Gg�C�<)�
��B$��`�k0����*�dj|iE*SV��6�|��ke��A� ��QQߥ��L�F�@c40r�C	=�~֎�).m�m��u|6��5�[o"l��}��/�mP��Ҁ��ō�t;~uB[�48�N�s���a*S�F�q�:o�Άx��8�G�^�=�F���Y���πE�ʶ�/�ψ_�o֓3m��c��'V�تelX��nC��u>�o��8��,L���*�,چӫ���P,����#ᪧ�����o��%�3�U1���L���;@��o�SѤG랰��wcVY��z�Oq��ǂ��2*��}&>:ꂕԑp�}�u��㴓fZO��Q��c�4Af��Ç{��ȟ���`*�2�"w%7ڐ�Q���Xh��l3}opm?��#1l�.n����b�Ͷ)r����������E�k��{���꭮4����$�r�Z~��p��jVQ�����l��0�}�5�{7�$؁Z�[8���� ��+G\�6�ӊצ
l����j�E�1g���X�_���\���h;�J�+�^��t۟�E�0] ����e��c()	dT�`-�����T[�*z�@�}��u�E�Q0���֦��}0�9������@��l�l4�v|ˑS����x���`8���Q*�ۿjl��a;u8H���Ϭ��+�gI��� "E3����&�3�\�.G�I�Z������Լ*��|i���^th!�n�/�EcS�8���I��d:d���@*a���9�!���Pf�&u b��p���.�{*`���e:Bݹ�L�C���"sR��w,ތ����Đ�G܂x�r���?��1ˇ��j�Vu��4����i勘Cn�`�L��� �Ӓ�G��"=$��tD`/�y:΅k	+�&?�sI��r�Ʉ�g���&�d�?�dx�TO��\��F /~E���wO"�����m���{p�Iz�glU.޲�:�5�1��/�Ϟ��"z4+H���N7�7�Ӷ�o��Z{Y�X6e{:�9E����B=J`���{�%_f�r���	�����s�BTL@�eC�.���ݥ� !���@�Q����ڰS$ԂߣI-<y�c�޸��d��ox�^�4�g��V~�E��AMu� �VB�H@i�M˿�c�a��u��
�l" \[{s��J�9x�����i>c���	,|�,�Iÿ6Hۧ��ç\}�<�����Qk���r�Ԍ�"��6M�sM&X�p�dj���Ǳ]Ǳ
���:A'P'���KM�U����U���3"�/_�,���1_��S��tǞ �j��o����̬�O�$w��@����j
�k>�@(%]�bWf�S+��dq{pYP��*E�?�Yo�y�"J�üy���+�S�JKQ��VM�������#���{{�f�Q2_NWW�z*�y�kIϵ��M1:�hR�ۺܧau@}��;����.#�H1��!��2fգ���{*[#xýƯ|�d�8T����6�+n�QJ�΄ɽ½�v�aO�sz���oX/$�����<�t�H�"����� zU!s�0�z�:�C,���#���A�؃��eb�u��a�q̣n���4y�x��̧��(�P��@O`-乵5�;��P�{
�֮���p$A���{�,��*d�M	=y�J�آ��i�j�pɦ쬯�x���i%��{���|jчN��|	:�]|P6�	�۴,HKB��g���!�H�L�C�4gO'7�G0LF������Ol
�����'j���,�2m|��mY��Q�~��*��C�A,]r�,/�<��wd,�0�)e	�$K�Aւ6X$0mR�\-,��+h�x�X�#�Ţ�!	w������ �k�&ݻ��z|](��Z-�Ub�-��Rv<3w��<��[d0�;󖳣��$M���[����L����R|!������dYpV��<��&�<K��'�+1���#�i%�Do��g\Z�|F헇^�]ዶ����#^'�8��tSvBL��|3������N�(�Лǐ-T��v���P4^ԅ=�)�=�r!�k�JF�j	j�4Q`�A��8�J���(W�g�ˊd���w=*��E��̿�ew"n.nb�y��a��к���..�$r���mlx��(��s���u��j�A8�D����Dn1�oפ�߇�ˌn]���3D޼Ҋ8��hP���w�T<�q8�el��5���}b�G�"!��q-��c�{%�)j�e�f�G�io��Q �i�� ~#9�/_UN��E��/E{�����6�ǂ�~#�Z6K�G��[��~�_��k��?�]էk��Y�T�0$�Vf���@=p�׾b�S>�<xn��?�HH.Ń�p q�Tj�u���3�.IF����JA3F�op*A����`�;�.��/<�;����#��X�c��&ȸ<d�i�4�*M�Dn��3�
nYЕ���j&xcF��Q��瞹�3G{}T�����a	D2�**�%��Z�1B��Y�Q)�҆�/�	��ۺ�R�6 �Tb��ɈB�!�봸��%(����#��J���N)��wz�җ�-A��a��}�����e����7�9��^���0�Wu���_Ԝ�A�y���6n��TGG�t�W�p|��op�9��,穼�ɔ\�r�ݤ$��Ƒu��0Mu�,K�&�Nu�P���7��|I�ʙDL{yeb.�����p����+�p�����T����Qq�Ί�mv�"8�j�N��ɘ���0J�&~|��7嫿U7��=�-�n�A ��J0o{���>6 �:�F�۟3 s��E�$��S"�3Ԓ�P ���H���A�����֨j�M�fr���ymI�>�B){��@ħKu.�ì�{1�X[[�ư#yeL4*:p�x�݅�,�R�w��"���a�RgN�y�r�r��K+	�KJ���,{9�v�^S��'ݫ9�eʖE��\����9�
������7|�wu�)��VJ�'zDgMZ�(���=�Ŀ�,���0}���ː癠:��1n���C�6�O���d:~�n��C���ԮZ��3Q��q!*��&���D�l�����M�$;6����t���e3��8��Y���pI8�84q�:���� 5��: ���S�GK%�4`4�|�=���**��a+m���7d�F>f��-�c��^�
2~���Kq���8��ٹS�m}���������S2s��Ʌ�V/89�X�,��-�Yæ�\#���0n���Y�č���j�23��R�/�~��5f/�
��,�:��si��N�p[z1b~d�� h���C����=b7�>���!���e]rcF��}֚�Ƒ�����a�iU+G0���*	4�e��fPT;ٙ��`���:��:�S���{�# ���$�S��n�C�*��A���r��	�^&��}�e����t���NX����d���= >���v.�g�E]�¯�V�L>��9�m�K�z�5c['������B������0|�[h[��g& �L5n��o�Q1y��~�c)2\�?�Q6OR�k�nnV����^�Î<keєRǰ�`���j��I��g�,@�����1��NA�]x��;��h ��D�x�gu�A%亵#���!��SB������Hg���WzP#��U�����i�ؙ������q:��ȴ��3���`hU�Z{op]���
)R�ձy��fٕ�l&_�q[[����DjC�"h��+􍘸+��;��H�TҼT:�V5�Y��LT�(;�n,��xG�>��5Sc���īWC�50��"���L� ��}��}~ �|�`�w��|���=�K�P�g���/ՙ=t?C������#�[���O:�u�M�ؗ�>)�`m������{��!Th	d,	��1(D�p�
�n!�^Gũ�/{��su�X]�f�r�=c�	[�N�úK�Y�0���;+��efU�s}�Y],����Q-�����r�*;vw-m)ޱ'�>�U�B.M�.y����F-g�$���[��u?Yf�V��{���q��SfȔV��/��T31�K�ZAw:^Jܵ/��E��t:"UO���rT23���K��	e�e�!r)M�2o/�Ǝ���$_bTr�2�T7�q^T!*�������to7����Pa�]�ܷ�p?�Ih;@�r*��w�ʭe
�Hw*��N������ �����ZS���ln7g5�u�)ɗ����l52��+r��P��x��	9J�oT>'���mp�cK�KV��� c�y�!93Ӻ`&��/?LA�~�ne�S6�|pM���vud����o�*��σ~Z�)���쭁X;�M����e	�//T�dw|�g�?`�N	��xK^���ǅ�W����m�di�К�p�E7Aߗ��g�I�CZ����.a��:2ݾ�I�f�Ak3}Y��O��c;Pk��(NS�t�j��H�����l=���I�~�ƚH�;X��X�l�N|7w��Rpb�_�G���r��,�a��"T'~�H[�Lz�D~%��,Oi־��\����W���$�O�}q��'���hF�R��q��?��
�s�՞2�?�u�d�Ϫ�R����q�M��^s�-�Jcڠ�ю�2~�vT	����W�i�o�� ���c؀�&�C�$-�^��X}�+����ز��O,�u"7FF�되?v��eKS�js�kC�T������FV8��Fj�����&��<��Q��gߍ��s�xo�v��0�UlV��g�A
yA6�[e�G������=�|�0>����m�f�>��_��S�s 1d�M�o���R-���Ou 29��>F:��z�V)�sU��2 %"7�l
�y[��c1�bDª����c�b�i)4VN<��.2;���s�lSn~2G��؜��}�����a�	��2I�������^Ee����e���_�=Д�< H~϶���(����&�_C��8�Nb� q�n�'/MI�㬄Q">�x�7����y��AWwq�r7��h��������G#	
!�ZY�i�;���|-D3��g^0K�l��j���֟{����șU��6~!k�M�u0>"�s$*�ǽX ���:&�M$�������k�\.�gV����3&(����%I���S
��g,P�z:�}���)ϊ����k��&�F�����~g'�L��5h��|Y;�7s#%�ml��K��"<�)٤���v�{{f���K�����Ի�t��ka	�1�W(b�c�����17�9۷ƣo!��N8H&GQM&,%�!������{��½�t^����A���������C�����?��=4��yb�	e�O�~��(�Ss]�r�J�j��C�jq�>�;s�-!L�I����� �����,�u�F�rg1]�`�_P��ہҺ��^�r�/��6�]\���Yu5]�&��-VS{����>�i��1]���C��K�;>�)���dlyo�i[a	���m`�_����6&
�˳F+IEm�q�����جm[��������0��h/n��6�|5UK�BGe��6=���:BFN�:c)턘�^2[2ҝ�+oZ&um';/��#��w�5�O Թq�����~;;^	�/=@{s�~���Α��[�2ޛ[EH� ���3���T6������n
P!����E��i����o��Hu�/���;��LA^M[:U��6z�.�l�.�tI�}����H-�������HN����4��B����%��d�����l�2q��
O���� {������K��(��i߲��N�VC��ܧǠ��)���۠�b؉m�E��bF��mJpV�����+�2 �HwE��|>�F�RM�Fϝ ��˄��}=�n�j8��E�`��3����Nɥ/���@��Ӂ�E<,�1�t���'������˃Ê�od�����I62��-	 P"��a�lʗ�pL��>��<�����P:~��B�Hhm>�%�-������-7��ʪ��ko�՘��"C�6��S�7�y����å�<v������rd1Bh�c��f�h"A���b5����3�I�z��aS^�R[d�����Ϙ2���u�VS~�Nw0<z������mIut�3R��!_��Ưh��u|_m���1���.���L��M��>�j<�H<��\t��~��P��հ��!���<=�۳P��
��A}��U���A���X-�gɞ@��,�Y���9�>T!r>�+޴����)u,������z�5��xM[�KnY��h3_N�^K�-�@4���zL���� W�5����TD�j�����I
=��u��2$�����~�ti���
�Tɶ�tUT�x�pST͒;z���;��>�A�Ht��*~^��Ѽ	;Qb�����LG!|;g�c�b|9�w:��,����k\��o@�g��3�����t��+1p����?��%@�xt�	K �@˧�(M|�����N/�쉶�x"ԟ��GPƝ�VW`2�+��E���0�� °׌���*� ��~��L����4���x��P� ����"y
�S�?1�SSi�� ��z�Լ����<�!Ǜ_���� ��~U]J��*�"k�u���3M	��m���޳*�ׇCPgiU��������{����)�q�M��:}_��6����^�1�t�0W3b�#�ڂf�ի¨u6��z��#xsi�w%�Nt���������v)�b_�*5�J�v��hY1 -�O��A�{�b�0��<]p�M9.�A����P���h׻Eg0�xxо�2�J�.����$FB8�؟�ӄ	"[.g���n��.	������VQ�M��(����,�NLWߓ�	"%ՙ[��W���h�l���_p�H��2��^���K	�d�@��a2���	դ��}Yk�*1Y�	�'��Q��QT]���C�%.g��8*\�T7�����2��Bzu��&�pǐ ��U���h߫�7@i5Ɇ?��p��n���7%:�.�dz�?v%bP��7��\J#LTi�t�|���-�^�f�]NySve���
�Cgآ���K�re��\�����=0�P��C&:}����#�BR7�1zv��Sк9�߅#ލ/��Qrq�
���rg�	W+�x��Gq���)�����m��P�5S�!$>��'�(ς` ���s,����) o���A�9���_�ϟ$o�Z���}w���-�Cc;Q�;�9�_v�>�ѫ��C�oW���7�R��ʖ�p�_���^*Lϋ<rn��%�{C��r�GI�*~{f�w�r.Y�9�a�?�ԵI�����=Y�o��$��S��Nr�+p�dW$-�-������lb�89gתf��ww�I�4�4`��ɐ�f.v �K���G����� i�SH�4�VN(�l6��i�"�%��ECɗ>gL$��΁u����<�[����f��ܦ8�Q�#ʵAS��]'r��|ʪ��������������^�n^HT<��v���h�ﾯ6?��l�s����"�Qh,@��⯯J�_���H��K>���z����O�m�h��g��&�T��e�U�C�j_S_ˁ��ͼ��e-��C�*%��EG�1\;<qX������-��y%��r��G[��K�M���G��P�s�TfA)��4��-" ͍�;��Z� t�XE��v��Z�q��7�z���0,���{���r�6^��a�s�~t��K�Ay�<�V��|���ö�h�3)��q5����޾�����B57Ć�_��1X��]���j�b�_�l���� �&[¹^s K��C_��T����L0���1�*��� Vo��9Pk�����M{��ۂ�h/'=҃��f��Yȭe8��O�U>����wZ'�Y�5��욂��+�d�Q���4�����������dF�7&�d\��EF�݇r4r��ª�+�	�r�x��ױm�z� �\#o��]�&\>\��x1��K�8�ӫ���'6U�3q��x�.E��35>D�qZn2��A�<m�",����9+9Ox�� 6�HUY�a��Llv�1�Z��lq��퀍�rk]�U����-I�S���)�_�dP�[�1��M��b=	]�(��X�㍆��)�!c�c�:TkY�����<�����_E��*��!e�ju��K������G"��}�*'"A�蠶h=;}��es a�Xƻ�q�t~�� ��d�n�=��`}�Ʊ� �����}y#)hU9�?������<@��*m`M[O��6d�������۴x|�[�I�iwՃ�;�X���Qd�͜���aVA^Y�OEdy8&���]�LDR_���`?em%�w�y
\�`�{�{�����mp������)�e�p�=�LB��3AUh����:Iӵn�.&�$K�J	�,�"l�P�<���F�rU�H�mnx�E��
����U��*�m��N���շ��}�V��LE�!�{ok�,���؈6��g1��w����8g�J.�H|�κ�����W���T�(�nh����Cl�L�b�'���.����q�G��J��RǓ֔H/A�1Z�~�f���xN��v[���W�ZF���to�{M��ϩq)}Fy�؏#w�F���6�x=͍���cq���d�4u�N)Lr�XN?@�>�T0�����C�t�E*Q	��n"�B��Ec�^V慈 �C�
�w�g AԿ���=a�	}�ǯ��i�N�$�vB��YA�W�ZY�p3����n*�*G(��D�FGk) j>"�De;6-��8��7��\r�h����	�z8����ODT��_��2A>Z0��{F���7�b�ɱ�a�\�]� *�!U,Ǧv�*.�\a��x@c���1�;¬�v��t�� e���!���~����A؉q�p�9�?�&Q�$�Ăæ8J=e�$(����]��[��4`�@cb��vbY�}��p`2��L��!���YO0��ÎBx�oo؀ô(!��M�,5���/����X����U`b5u�Վq���?�m��^v���"�@R�ք����G�]��
Y��=��X�������4:!�(氝4���Xy�+7|�v�����A"�{�����'��r+V�Ǔ6��v�������qd4�t��L��Y��.TA`4�ϐ1?x)���!�2H��2>�Q�o�i�;��\� �L�0��D�� �ܨ�aBg��"SR��t�d���0����M"���lf
Ҹ��ްǟL	��S�����1h1��F�a��6%| �������ޯ�p�[�)�0}aƨ�/�Q&8wJ�����V	��S!���1�:��J�엄6�X4:��x��f�|�f ?t"�I���ކ�4Ͽ���XV����8��Y�?�2Y�_��?��%��SnU��ٙrC��*�V{x����.�Y�K$|��Ԃ|O[K7 ��8�-% ��W�h�^ҭ�G�X�?�uN�o�\��a`'2�1�P�����%+��F2��w��+h�ԫ6��zv2�h���_�y���=J\!�]��5���� �%���;�?�]��?8p������.��
i2�ZÏ�m;1��s-:��^u�n��V�K%t�g\�e6Ʌ�hp���k�&d'Lds=B#j����^�ǽ$%��ڢ 	�gi�)�h�/ȸ7D��c�k|rf¯;� c��y5l�a.�v"�{r�n����:����s�|Y�T��m�e,A[ZR5˔[���x��8��(�#��Dp=�� ������(��(���2ӹ%A�p�Xycr�(L��J�ƶMThEG)��9�j(����6�/|S���{q�I|b	R��+��J�qE�ݶ��؝D�9�cyE���r�Ќ�׬�e�U;t���Xp�Pɱ7Z)c-hU�R���J�w�.����4���dP&_@�oF���U_g��w��7�2W��cp�Q�_,�+}��p��}��"�yek|���ʔ�|D[�;�ō�;���y��z�(ը��F�q�[p}j�b�-v��h�v��ײ��+�;,T�*��c噜��Cv�[��hǳ��ꫥ� ��t���)tH{?��%��+i#{����`�w�->�}������Z���F���ubNc/���x�򟟻uOs��ny���P��[�!� �y0�w���79���+�g�
�Iډs1��\���"��m��˶�3J��B�B�3w_��<��3>,���`��ű��Ng�ם\����3����=�e�ŧ��K���M�JfO^]]�{ʭ�޲����Y���� *v�b��Xw���!��=c"�7��5_�/{�Ô�3��Cr�K��
z#�D��3{�!n��M�2�ϛ���6��7��B������C�ڞ]��U� ��R� ������Ν���m��3q��y0�ª5���N!�a�U��쬤�s�O��l�`�@��r���l!i	�*�p���k��g��P�}t��u>�i���li )7��H�ю�WZ�'/���l��jD�����[�5_E��k��b��c����$Ү�mĸ������'��3	z�gK�p�'K�!���X54����uޘH-cd���`�#~Jb��˦]�� L���󨰚)��Vei�gf�$qԙ�P4�y���P��4�.�%�ULE~٤ Sy� �Y�_����hڪ}�@F4��B�Ֆ8���jЮ	��' �u���a���|�{��y���Ĥ9�\[s%��������}"�#B�I�ぴ���Y��_�������j��5�C˫>n%-ӽ\V���8�8 ��4Z;�����fz���e��d�g��9|q��y��xt�wH����i��<<;
�I�s�m��P����ȉ�f�D-u�����g	ܟ%$�sILTH�}����uv���bO�AXG�r5��˲���O�6�_#q�NB`~�ڄ�AZBNb녯���p�`�e���x��'z��-=WrBy�nfFf�IsN�}��z� hX��]�5�%ו����O��$���I�PMu(V.��.���z���6\գ���ͼ(6"8�"��:^����m�&9a��Z�M���5��<pS3�JgX����Gďh�>�3�Yq�/�0��0.i�Q���0���}Yv[�2����nB4|��{��a���_����W�֣Y��������4G5��rL�����$�/�N"rx�OT���[�.��F�P��s����!d�	�WFo*x)1/��MF_�$n��1�	��E�|#�s"��A{e2��nE��}�#F��Ϣo��bs� �U��kg(9�>JW$\��`��"i;��GɘeQ����I�$ڶ���.� e`�9����N��sE���Ð@�@&�fg�G2V�&�W�U��Zֶwt!�*��w��di�h�"�#�Ƅ��Ǭ��J}�����	��C�<�sza����z"Yz�pRO�V����a�G�}8�+��ϲ�
cjV��E��;8QI�����P���rMǷ6�e7��1�%~ұV�߼��6e�Ta��|�@I��r�[�LzS_M�i��er��X� ��f~�v���G�A�-�ۃ���qO�Y(�iX^�b!��M��ܟ�������f��'��r�:q P�PY�3�j-S�X��3�mU���$�]�}'=�vTkK�>���h	ZzI�ɉb�/��YN�pa�����?b����^z!��V�=|�Lb��Eڄ���,�d̎@N�A޿�8g�04��^��@lJt\v�Vo/4�Z��m�'�[�Ƅ*8X���y���{�v��>Q��P����E�ml��
a�/ѻQ�����L�%[߼$����&0���#V�/�q�8�i���V��53�LYU�0*��qR�Ǭ
l���(kEc�>Rz�THҩ�7`��½6n�)��"s�Rg�oy��h���H��o�_�L/1��ބ/cw���Q0MK�((z��/c橀�����T�x-�:Dj%�?f���%"O}M� �A����V��f2i�gl�L�|����ʎ�!�n�^�9��M�;|�zn�s%�۰GÊ���Q������y�J��+?Ƶjk���a��]u	���4:/�U�2��4zX�c�jFՠ�|I]*��@pdr��R1T��`j������^��'�jpj�L?z���ᤠZӲ�U��u�����+"h��e�pk�����I�J�C=�t��5���>�����=;�АoR�U�d����v���5����܆8I���9��Z�)�!��ٱ�ͳ
���dB]T/8���e��x /�7dOo��������<�!���#�.#���
�n��4vL�%A�'���߱�'�GG��l#�h�>�sp���R����{��:�P����9Z:�N;���R�]һ�/��>�s�/��<�6��$��<��$f�Y0���ߢ��4���&V/'����%øL�$�m\{�8p��s�k��=Aα�����u]_F ����jI���[�v�������-��	��DL�A����61��yg�`��&�rQ=߁;ApRـ�Y��)ƈ�AG_���G��j�
�r1^l}��[k9p�e�g�Tb���${�3�gGLf@:�j��s%j���T�c1>�A�c+�9/��>�93����2ؕ��%kT�W�}��y$	'�U�*�>�O�$b�NA�+�_@��D�	�_˹��%����K��%�cu�V��%����1�\�N���N���C/a�)�Ҳ���s�(��h��*���pyl�5P�Q�_� ʰ�P;z���Q��f�����j�����/M�جS���1��,�I�g��f������K]�<�?�9P.�_��8��$�fsw��uq�Z��&7����{Yh� ᙔ��j��u�J���21��ґ̼d���`:����o�i�GE�Z�M��H`<H7#�h�n���>�,�Q"��0�3�D	U��W6 l~ ���<%wMFt�R��}E�<�e�M�0\�v�!'>��gH	��"l9�CMw*% �syNX*������~6n�}�#��Yӳ֟M1���ڽHoc�/�Ng���9ģ�[���&�*%�A������|��2x��W1���o怤c4h$Q�c��3�14gϖ >;������L�T�n����T�E�$��&��'�H*n��6Wqh΂&g?f�h$�G��U��_��
�]��VxV��5yTȦ#�o�ʣ��J�F�n�R�R;Qbj��9�dg�'A�IO$�/��DS��̃����*&s�c��c��sq��B2���^k�M�5%PA�L��:�o�[ssU^���o�Q��8��Gy�x�;K4�y�	Bd��J�����F�	�p���ܛo���`���/�P2����h$�p�;��_&�6!�y:�M��7�.r�&�uL���FA\����d)�ձ��>�����%R�D�A=�\P�l��K�Xd�#:#�_���c�T����zU)�;�����5W{w��9�����*��-bSd`��ݖ[��CF�3�`�zhu��NQ[6��+N���s�'����E��q k&;s�a��rTꜩ�ݢ�Oˡ�t!*��k�պ�Zn1B��
���O��R��]��C�u�i��V�����n� ���P���1�i;o�6=<���R:�Vߩe�4�u�>U%��ɽ�6��¤��*J*�O�,�l7�h3˯��%<	-J�Q�z����d�k�Uە�L��,���i�x��^#j/��rBҘ]8�/��?,QYտ��vd �2&�Lr�8� �RZ����Ym�(�/[#�|�Z�h�/��+<>k.�e����~ijc_�g��Yw)���vüAf_�(�⽔���O�rl㜁��>G���}�Efhj�»�LG8��JMt���oӇ�[J�����{�f�/��i�jw�&G������A)�XG淥U|��Dzh0ͥFGK~e2Aj+���`]C"%���|�g�u�^��͠���tW�A�4�z���x��;�(�0)�5�������� �2#�!���-r��$�9V#�����������9�(|��m��bF���?X}}Z�lz�@C��7��ټ2a:jj����ρ������z^b�\m�<�o�� �	�o�3��p����!�î�E��<b���}����!��f�tK�"� ޜ�1u}:��LxG�>&M�=Ů����� ���!Ck�(�
l�L���}i�C�§J�GX�oj HSl�o'��I��7�e�[a3i��a�Ȇ[Th�'}#�k��rY3�(�|�f�+��wV�Z�
:��S�WͱOU;��39���������\�\��|�(��Б)%Yx[0bP�dJ��HkX�ƀ��3�J��Z�=y4�.�!q_s�#}F2�ҁ�И����VH�T�n�3�@q��,��z�Z�Ȁ/c�'NH����l�S50�g�BH}W`�n����܀�4�t��$h��n8� g3m�� ���xMdyB�c����7���۔�$�|�D�'V��~'��D��x<����1eZ�.�)s�&.j�pB��emV����;����.V-(����~�dJ����b^��y&�VW������w�)Z�y��|���Ot�Ug��xKT�����=��"6/ͯF� �3���\�|����hy�8�֣%�؁�|�N6�����!���oE��R4غ:�� �Y4~��KǄ�\ZM�m}~�r���F�r�p�T���������2��=�!%\��grڬ����TJb�z�v��z��u2�n��U�aO�Cz��-w�� sYku6��L�]\�=��c�$
�q��!&�v��OXs�6�W,nd$;�g��#;�a�a�<�X��2�n3c;�px-[��C��߶|hu�?LB+S�/#g�?����g3�,B���r��F��g�H�����l�[�ǩ�*����$�
�]�K�0�$�[���v�J�yM�	}�Tϼ�<�2�����e�$�BY�_6��עf#Ƶ�i�]���b��(�_HQ�P���G{�4=�|��B~����TY��N��n@G��W����$��%�ߙ+��8Y�N��v�vZ��������������K��	>Ƶ�l���$RQ��9v�W���-Z��2�xWOn	_�e����m�Rc��ʹ;�:0�h+M9�`S3���Ǔз� ��qe�fC��ƿ�8���w�Y\��>�����U��(>
��yg�%��p�=q�M�R,E�x�čw=��ޥ�
z�)�\�Ik��!�=j9tCN�:y��*�������]�2�9D��cz���&�\����=�p�C�����./ǲ�l�����@�-��u��-���k��fcK���b�.rdO�����'�]��+mL^7W���B����WhT��@�X�b��Ը}��-���7yG|^����ܣ��!Q��+ȏٸ�U-$W�OQp���0w��ҽ�ö��(B��=r(���W#�SyX%Iq�ٟ~�O>�=�Ab�z;��0ָu�e�(l~�ƺ1$��:I��U�}��[�P&-餳�"�h3M�t�=�-F!x�8��x��[�1Z�)#�8t�j��뛅$��-;�-�.በGj�!��_$s�&�]���M(Z@	 �.єl}�e� �sG���a�|�-��$`On�fʴ�'-s2g�{�O@h��x	�/�\K`,����_Qe�x�`Σ��E��Ò�mƟ��D�eWte%+y��
N㷖@W�?C+?�4�̆���V�8�F\�D|���	�iԑn�~���.mN�I�����0�`�c��p���kV�s�vg�'���}Hy��p���Y�oG󋩱�6y&Js	�j����7Q����q���f���㩣�m"���'Ϲ�R����c���Bg��"�)"���G���'�D�6��(��ꥠ�H�r�M2glG�b`��BQE;s�f�6�,>V�0��RŘ!`�m��u~�$���u7�v�(�nX�3���¨���$U)�<�&<n�ЩINvPֵtj]H����+5��۪9�4 �b?!� Q�3�z�>4P���>��	�m���Hqj�j���졊�zګ(�8�>�/���21Fl�a�>�}B���V`�2����3l�#�ńw�=͝�_�|,��["i���a�Y[K��@�^%��!͗2��+5m� ݮnս�ޠ�o8��_r���e1��W|;!K����7���g�ȊB���j��ҳoyy���5饙��d�S�LX��N���y�򒠦������>�L�G�����*�W#:I�D8���\�͢y��;�� �bO����e%�U!�I�z6�(�_�t�(nah[��Rqg�lO���{ОZE/�$�Ӗ�k� ?|��R#��"X��V���Ϝ}g�(��%ny�4�lOi�XbQm�l�֬5f�����ɸZތ}��a�h��]��S�&�.b9�&�▽Y}��}�E�n>g`*�$Vd���K���6Ư�"���A�`hb���S3����SG�z>�a�����Ӛ]�w�6�l����-PRg`I�;9M����Q4�L���-@��\z�Ci�>*f����jQ����b@�����& �8�~w�����n������W�b��Ú�p������t0�V�T�/x@�#��QM�e�n�-ݥ��v�Z��Ƒ�� ,&��B3��>)���� #�:\�	�:z��v��	e!���ۦ��У����Ʃ;U]�3�&B`K��X/�bQ��bQ�ͫb+:sf���D��w��|5 ��^	�c�v=�w(}<�,.Y�[N��\��~�R�A5�B�x�/�d���.��0��*K �"+X�>�d��	���Y��C}�X!ｈ����%�p�Y�x�goxN�^��lk�|�s�wyw�o���婟���$.5G<��g��8��e���{�k�a-M��1Q�V4D���*e�;��7��[����"���.X5$pS�	�C�+v�r���+16��C�cL�(������02\�%-��"@B�Dx������eTq@��s��k�qDa\,T`�A�វ�")�j���Fy��=a��di�KHSDrM�b�ޜ>T����-1���sc���e�k��T&G��܋	�t��<H�>?��B���g������	���a-��$�r���|�4?|3(-눿�/{0�2p�����K���a��iPq�:��1���|���mͺ쾟S��,�x�7M�F��icy)+�baS�8Lh_0K�d��Ʉ�Q����uW�_��8��̞��x�£���6,�Lix7�Ի�ɧ��A����'�d �ͨ<j��O���*p�� F��;��-��[�&�4�Öw0))�p�<�"&<�+�M@#�� ��'r�bgW�Ɲ�(����%K�0(�bY�?>R��󹦀���ɡw(ϛ�=;���a�mǸ�-)�Ϡqx�c�ͯ�$o�S�����Ȋ_�f8�9��7�Pl{dڲ�|֕����b��l��$A{���y:ء�RB�t�`�d��|�O҉�Ft���R=�����!V<Ǌ������Ȭ��<�pi�u�[%U��(3��N��d0������b���?(O�|�dg/A��bM�I�quna�5����/x��WtS'�ևJ�n8A�N�E��弡y
ފ�D�W�e��f�[�dԽI���BH?f�W�@XM*���'F�O��#5�PRܦ&�G�kτ88p��lh�v����9�?�)�PB�:G����ƭ���z�=�$��:�h������xwhz�Fſb�X�i���l�;X��'�w�Χ1L�+%��N�h6a��C��d% m&�m���,�H�L��~`�V�Qw����(���{�!��ƝϨs3�f�S �������F�{��=L9t���������c <�C-Ĩ���?S�M���Y�؅/Ţ� ���P�����(ıAؑ�@{¤2��`!�"B7���t�H�٦*�d{#��,/��.N�C/Y�Ʒ������`�z��d�	}�b�������Z6��3�n��"R Λҧ�Q���g�.��ვ�3Ԉ����~��-"��3�)͞�f�����Z���ɸqyM{�j^`3�ٷ�n��+�;�2"|:��s%�0N�'S�om�J��;�p�V$r6���	1%p
�G5)����l���*������T�4�ZD'���1��]0��*ȵ*Џ�(p��=4��n#Ct<�����s5鸲8�O��)����[~�T]�vud.��w��s�^,�k&��G����e2g�l��Q+mU/C�le�i=��\sk���p{sW��2�P�G�@i⿻�^��?۝�7��ZaY@��6�\�jV�i|N
e�w���;Z+h�X<����n�����I����	����:��j�J��頠SN+Y8�����ē5"է�v6S�T׍��6�o�e�C'��]C=�Ҋ:��1>� >iXR{n��N�(��.���iK�X��P�P��e8�X1��A^5��'��@;wH/4ZN���C��աt�M��ۍ�	�h�>�I����Uֲ%&"-�F�,���4�����y\�s �����^�B��k��B�+G�ԙ����fM��&���1|�� Ȭ���\�[�;��D0��:0Z|�u
L �K�� �y�0��ٶs �:�b�#�z�#�g�'HHGMv�!���f�A��{�_-$��j���i;޻E�>>n��1���{9��7�$�3�Rݹm��|W۞��KnL�L�gE/����n�˶{Fgq�m�.����4�)���%���2T���|*�cl]��2O�O�Z���Ĳ�{�r��;g�4�Koް-�\(������Lyw�s��Ǘ�=2\T��N`�@�$��Q�_Ȏ�&�K�@��rHv�ה1���P��StS���oٔ�ȧu*�sp>�-�U?B}S��Y��ŃU)f`k�~�P�n�
?A���J"MC��;G�� �P�m��p�z]H�Ŗ~��k Ɋ����\�����Bh<�c�S5A��5�(M�*���cL��Yy�&�|����\�xC���_ynm�յΉ۰�UөN��xhTA�(z�-�'8`�a-意�9�:F5f�q׹��`�2�ϡj2����X3�E��7[�#������an&g}4�� �ڙ�L���m�'e�A�2�Z���8d�|j�)�#�-i��m��C��>f~��r	/!!S�5z3�"��Gq���O��ǯ�-�q�i1�ҁw@�h$񩩮y\�}��P3���';j�G߁u,��ȸCɥiz��0�S��h�Ǿ�1_7�;:�������/.�c���x��;�`��݄�=Q���`����1���srEjϙ��Yd�$�
�v�� -���xC'yG�g-�B9���xq�$P�?d�-�U�@ �����6���e����ɅG�S��p	w�kb�nɋ�[)����t�~N'~�������eE�-�
aWY��*����s��N��I�3~w��k�P�_�J!J^vgV9��N���������<�F���L�R����i��%/Ե�βuw��
ap��8�#bA��/��Z��x�)�_�<!f�4h���Z�&�PZ�߱��Y�2Ș�Ro9���$�)#~3�kX貨�
�:dD�!@�|��s���Jb�D���#��rڴ��k��j���iw�@Z�P�/Z+����N�V��jmx'r�;cպB6��@�{�>S���!�@=$6��'�_;�W/ֽ�v�S�A��2�,57c�i����)]Pw2J�3��o�� e�	�s2��
Y�\��T��#�ߤ:O������f�b9��U+���J,���g�s�	c�X�����vLHެ��}��X�"������ �=���#k0���X@�r���_�?���~�^��RL�
�}����uk��P�8]�'�n�ߙ�z���ᑦL��f+%9�t�p3[?0q��x>.`b�Tat)���I5����Xd�9�����,z��d\%Z)�AC�`�/v�f뻟:���ro4���5���~��(�����ivH�T��(��辇Nq�a�RF�r�'����J������'�M���eTגJC��^	}-e���\ʱ]n¿�G����A�{[�P,�Ov���hd��i=������k:��ܖ9V�<�$B5�R$���Z�tn�`���`׼�C��G��SA���]�O�@Z�nQ}�����ŉ^�lm�>�=��95^������㞚�|�rNζ�w��{*�!�ɜCv�=2�'��~���D)}V��XB"�0�J�Y�<��_�9�,4b��������ǹc,��m.7&~��p1xY�9���y�i4��ڏO`���v���t�V:���H�ߊcxe#��7�i
�9��}O��e�qx{�!��\X����/�	_P�|\"�A?bX��b#X�ÔJ�0�,zL�����rVt�����
��C�c�̱}���c��&lQ�Z_�U�&�~�������i�n9�"F������\F�\_���3�x�o����O[2Å��eg!,e��o̭�w,ڝ뮝����x���f��J��$��W���Տ�u�
ő��#�8�}�������I�v��2}VF�C\O��m*���F"I���tBj���O�LBB2�+%l	�(����j�>3�+Pp�[խq(���A�����R`~��lP�T��sۃ�ԳD���Ov%��I����R�9���"[�,;A N�N�>@�m�I�08�aa�Ξ��g����|��b�<+�=h�KT{�U�ZZ���G�s�-�"h�S��zY� �vP��w�I)z�M�r�9@E���_����WN�X�GH	�1eb�G9���I�<��4�#�䐉o�L�P������n3�z0���$s�P�ax�����XhMf�X@�]��S�3:��p rS�|�e�lg4���tը@��㠢����e�<<C�LX@�@~�B<�ݢ�84%�.��u�蟗k�FO��U�R��N�XH3�� ��~
eЕʫ"բŷZ�i��EE�œFx������in�@UQ��B��,~�ؘmo�.�.W��W�J��
�P�6LF�.�b�"O�����+�.�T�1�j���(��@Fo3�̛c��Q�����:�'0��*�T�٪�Y�h�r
�7*M<�[3M�y���/X�_��AK��3-d����/#�M6-�+[
+ irؗ7D.V�`s�h��:��9��'�f���?3�Od
h}?��KD�i�\�(����	^�	�R�X�mk�_�R���?Ke#��1�;G�ŭ�u+��"������Ji'r4a{(�^�\�e[���Ƅ��R!R�`#.�j/@�-s2~rB��x8�2$ݽ���(/��z�œ�Xv.��x=h������9k�!
�z'�S�/�6��j�Z�L�����ǜ9pf��[GU��^��qy��#��p��};&�3S���$�(6n�'��SX�J���I�*þ�)��"6�^�H.�޶��?1��[�6ޤX��!k��1&,��&B&a�_�I�,窕|��SCgG���]�Ԉ?��ԧ��$N$#�Ej��a�;��&[���ۆ��L�cL�uq��<�S#¼�8&����RHv�+���<%c�i��'S�w�F��XO �ZL����B�OY�60+�v0����"@�����+hm�݃��Y����Wj�4BOu�ҋ��z�q֨���d�ՠ�˘�Zۚ��/z�T?�-u'��kr<ȳ"��CՀ+�ˠ���0蹲����K܃�_@���G�<����mu�hL���[C.h#n�UІ�(<ÃZ�gq �������[�q0��u�~��3{�L��/�	U��aO����Y�z�Qw�o|��f��ρA�iJ{�����j1�������F	�߷��`�ml.lY
�y����+Z*g���Ƿ�Pi�S>���vo_�n�^ܳ#�4݉�E�C55��7�G�6�Y�Â
ޤv`��[��^D�q�xn�j�nTӀ��b���_�kXL�ೇ���,�l�:���x���`�P���QMz|��g�!��cOq�����lu,h����OV���P��)Qk�9@�6-�ט4͐&��q�_��ń�����+�Sb�J��~��jl��-���_�]ֈ��+,��jC/�t�F�8�i8G{����II�;~Se�8�f����^pu#�r[�t�`Pt�����ި��>t��G�:J��vCHK@� �w0�}���K����L�*�LS�:[Ӄ
4}��G����"3�$̧mI�r����H2�^ࣅ$fL1j�����v�'�3�AQHg�j�m�`��Y��UJ�
q6e��`}�ջPg*pM��c]�ގ��	Ű�M�Z(���,a�j��k�a2�n(�ֳt����� u���(�?��B$:)�#���9�o
�yjg�C����~'=�,���o�{B'}�Q��kl*p{�{�OV
8�y(�
��/W��� N�N�FR�εh�O�~��aLF�U�Q��Ba�R�MA��g�s�'zg�*ۆrρ:��O@����0K.��Vr��|�%,I�WtL� ȓ�'��ו�å&tJ����+�/�RKq42���S�۷�.�0���{$���a���v�7JJg� �ˬV*o��6���Ȥ70�?�92veh���R��*{�����[~HBa���xz�j����Drه���#\��p��4���ŘG��7M\�MD�	ָ^��R�^���.S��` R[���DH�%,��;��]|���,��}H)�������z
�<��u��X��	"�s�5�.��,���Gc�6.F��4V̕u�Ĩ������yY��Q�s�}6H�;Lx`eƋ��+\w��Q�=�=��w`#�c�0G��K���_h��9IH9'�o*A�D��0���M`�1�m����`��jk�eό�_�����L1VbNF��FQ��U����~8�J�(�Fkמ^�|�a�m�'k Nt���Is�̓� ��x�x&d�E~�p�wԭ	\������n〗u�s�9HG��/����]2���̏�_�T��dHG#E�%׃Cak��C��0e����(C��'�v(oQ%1Ȳ���u'	ӿKk \u�{�m��V�(��0��ن8�_�e���Қу.+���g�=
��r�ƔAF;�a�UxC-�6��V���x{Z�(�&FGu^|O&���^�ȯ��S��3�=y�O��?QY�q��(�!��5�#���#�����V(zi;T�$_Vfd�	�ӹb���+��'kN�����_uF*��E���Ke�Jt4��0�oz��??۲��[	1��'ZOe��EI��_��s�X@[����$��Au�Ӟ���P��.c�;M�@]<���=���OcjwA�l�)
�����.㲏�S���vh�}�28��M8��Y����
ͿV,-�U�b֌���b�B�dX;p)xƑFQ�a+�[�ʗ{9o�W��e1[��4],C44~#�nNow)9@����$\�ۡ&�Ds=�}��(����A4�`�[�O7��Sez�� ��I�V�?�݇��=qVj���m��T�k�ܣ��v�a�ή����!L��%X��w�o)^b�$C|���Y�(E���vb���q�r�{;���
󾹿���բ��ur���ӎd������M"7Ƶ��v���l7עM��-��c�#D�V��_Ӈ��:�O��LW����u����tzr]&�I'�r,����7��Xf/�tX���Ցb�`4.��(�\vi	�^f�T�	���}���x��b����<4.�}�~��C�������_]t�.K�>ǥ����7M�%F�fn?�Q�5�A|�� <���{���������>����]8'���:�[3_��-`�꡶�d7� ���/2��z��2z3��Tw#;�܎Ň�Ăi��LUx�����P��� )=��&2�%���V�@٭��{;��sI��kv����l���e(c�B�je�b¬ ��֭6H<j��b�G�+,{�݈�I����I���Ć��?j�b�S�Ɍ~vj�#?��T��U�'��?�]9�\%�OY|�U��������Ck1f����B|�ޛ���L��d�[;��I����������&���C�f��V�ŰVp$ 58w�w�|�ʱU\5��r�*M��I�v��$>���j\a�А��_6<��(9U�p�2��R�uHf����4�.�=�,~4���z��Sz�e;/$\��ROL>*8���; 궈Y����-È�~��O��[�����c�Pt����߹{��XjX^�P���|1�K���F���$M�맓�N�	5�1Qрxa�/
�E܂h�@5D�Y'�}���ޟWI�ы���^��`��M��<�
��Lp��d�b��z'�w�sٵ��'���w�Wjq��!n��H���!��r��e�{��v�*�:.D?l*-�V3#!���pqB���g�����eQrc"�)��C�*�\�Y��}\�F�~�hr#y��o]�X��b��O�O�\��Z���d��Z3�W�Ld8,�1����{|��=N9��S�E��y���#�e��W���M��y�R��S:�9g���5���'~�5ur���b���ϔ��c��U4�{s��|�J��.9�6�Ԝ���ގ�%��X��K;���Q=������6�N�MH�]s�0%����O
�*����-�\�;��/����Z�V�$v��}�D`�+0|w^�&a�"�1�
R�D��	�#� �� ]�����ϐ�������s�a*��5�ғ��$r4l��Q6ɚ`���Ζ� Ю���tap1���:�?W�O�� j���cQrS��3ؔ���mQ�|��4>����v]�9f����E���d?0�S�a���)�������|�4�QGg�>�U�_�^w�eW��T]qqFv���s�u�b�-��Ǐ�	&����ű?ב ��LP���V�	�H|~}�*n����l�� �YIt�-����+�|�L'�&�~Fͨ��$R1�u��d<��ԗӾ��y'⪉��7n �Y��e����g��.�a`#��g�Q�A_	E�S��p5T7C�ae��̇�����K�S.�9@ o	�FVt�ǚ,��2����QxTzӔD���j����t���c��*�MWEێ��;���俏詚\F3
fl�N5�e�)�ޯ���*l�A��mi�omdX�O�˾���)�6u9��Vl�Jݮ��VĢ��J8_��?c���X`}R��aQ�xb��Zn:)=�N�.�͊�@�@2S㖮�o�\�Ƚ�/�=����P�RI{��QJ��t�{�w��àRއ�3cK�oAX<�7��Ztx��1�}f�� n��w�a^���9,�����V��^J=U�!�
�Z���z�+�:e|���С�%�LKП��٦��^t%*>7R.>x�'����
{s�}�#��{y���vJ�^������~�1 �q���
rqE��~�>˺)1��h5�Zw;L=s�j�"G�=�6,�Gty۴��]�*�������j�p�!����A�Fl
�l`��⢯�g\�>?�t�P	|�d- _NS��,�E�[�{�Zn�]��P<rR_�>'d,b�9T�MRf2;�n�j�V-���G�N{2��!u��}P�>,��t�����}�\B��x�#�u��o��� ��n@H�6)�I�jA�F�]�X`���+��_x��3�5����.(Ƙ@�As!H͡��N�C�ð��8+�Gog|���턱�3ЛO������Ex�ǣ�~�)��	����l �, ��W� �.�D�G��pFV��y���ag�S���ex��$��y9���-EO�ݹ-�j�a0������c�c�Y5ǩA=�U,�=ҩ;r��2e���O�8�O޼���	�C鱐A`/pa�߷W���K���"���3��ry�X��rz��hQR��gwfj7��+1߬lkLM��]2G�g皃��XA���z�sh�#e��z/5!L!�����=!ТG�R�cicE���M���e��ȸ}���w=����>��)�;(�o/������z�l���� g���(����X �-"��a���t�g�`�d
��!�Vp8v� �z<q��j-{��c�flm�%K�r��V=B~�ř��E��n�Zbݣq��KJL㬏Y��Hx��@j0� �M0�n�k�ͯ���S�2#}�H�)\�<ڥz�(��$̗��y��aA^�,<�^�1�4	T�����z��ahߙ��n����O�j�e �Mqx%���\�����9a2����Q��Q1�#94}Q�}��T"m	�Uw��%[ց���4��,�'�W���c�|��mE�E�l��:<�Z�_k�����Q��0�4M�|�V'�D�/H 17{	39GԔ�n����uPw"��&uh I�&�ٍ����@a�"�f�=%E
�b	D��]b�.0g�޽��!�g��5��n���qB
�iJ�����[�;���=���A}�#r��ȱ
����Po֪�ޔF-ȜwΫ��J��gmBQ�4&1�ogxp�6ت���c!�O�Ƈ�1��`���;V֦�$I��2�E��:��߫� �G�|@�ݺ�^K��&}A�������_P�!S�@p	=M���ǑCG���H"��'V�jN�n2�����M�a�s|�8�~�}�(�1�4���-��;���?������\,�=����I�c�-����E�߽>����Լ6��-�4�pQeȗ龥M�K��t���6T�v�ڵ�
B+i�9J���Ǆ�ᖫ�A�Mo[S�cH���%�ȳq�o� �c�蟎������>e?x%@�G>V8���NN܃�PR���2G�n��d����:ޤ����#��_�,5)�I'H-?y���zH��XT-x�f	�w�{G�ݻZs�adF�?�mJxf�o��JM��Vj�Ș��S|��G8�Nܳ��c�wE�+T<����\�K�ӣ��� 1�� ����S�v��Uy�+ۨ������V�<�,��V��:jW��ܿ��j��O��¸sg�~��l՟��Z��ԅG�>~����Ի��� ���#�X|�t��ng#u6e����QDc�����H������^ߺ9����/�����?]�摀r>��4*ұ6�\��q�>�s�fSn�4��4^7��>��f�E�ERT-�'T��_@�Kmv#Y��w�q���Uʛ4[�k��R��$ �QI�eM�{1G\x?��T�2��}�o,u? �-�vD���V��r!��a�4	Ç�Z�]ȔǱ7z^���s���PX7f��!L ��ƨ��֍�KH\魟�+r��Yop/�O�Ȯִ��[�z*jx����3�ǧ����CR�dp�u^�/��Df�5'6�h��wo2�F�U�U�	�,��I����z5���'C�FY��JH�.e�;m*����t�ڸ�#
Q��[��13�*a~�c�ٞ�1��'0M�s0_�ǽ���0� �q���_*�c����ƚ������-a�r�"p��rTs��=8$�h��c�Z�\y���cb�KU���8]B��l�[gz��1ϳ�-�~wmd��! lTW�f�1NKCr��h
B��M�<�`��W�̹"��K��Q��	�q7|&W��-�KMw�!e�y��@L>�����Z�Q��@�d&�[����&�ev�;bJ��b���k��9���Hd_j91�.�C�_uY�0_ZA�^7��g�@P�vu�f�E0�m�B|o̞=i��S��p&��뿾3fz���۳�G�( ���%�O��Q��q�:Dz�Koe���D\�x��:jĴ.mg���E ������%�on �g����e�\���n�I�tLw�Y�s����#Oٟ�wʝZ4��[Zd^�?0��z��Ac0�\Ծ��_��ƛ�)��y�[���T;mɤ�ڳ˿0޸��)G�Ӄ���ef�@o��0��7)*,��c�.Ȼ����
��;C���32��J4�L�+̑%�l��RI����#�/�V3�-��~�%��{"�M?��5<���[�"�gX֪����=�͞bm.N��4(M|RV�Օ�2~�׍�!<LO�a~�׹���"4�qQ����J"�j����d�9P*s�5��Դv�b��Z:g�F���9k��P�6?�\�]��.�f=�>.:@R	��U�7*S~£��k�yT
s����G�{Ş�����Y��epk�
X��fBtIXB�9��Q���"���1��LQ6�p�����%$<��{�c|y�Э?6dؔ`.J����,�-tqrG�)\�F� l�����}7����w'&��8i`5�n<�	�^���6�彉YST�����5y[�>GXF��6�l��!�,��39���	���Z��+�O�li��gF�ׄ<�	?KV��T=��Q��C^`͢e�
��p�d���,��rJB��\ֻ��mI�	'�le��b���y�.>G�\�,V�T���$�2�=u_ �r��'�_��(W��k(�!ؕh��P�f"�'.�S��A�v���
y����Y�q��/����F�LA�:;IR�
Sz~a�	l4W'_H�0go_�Z4�E���{��CYV�H=�'{9f� �j*��Lʶb�9�E�h�O�S�eN��,�Ͽ��McP����8o2D��?\\i���?X��F�i��+��.T��r:�k 9e�רp=4|�H����+N�t�/�ʕ����tU�'�UxB�+׃��&���K��#_��d��^�:�e�7Q��#�_g-x	�+����.��z�6��ӫ�'G����c(��V�4k��W�X�)޸�?��d��H�*Ύ�zG�Wz�[ϟ�kL�r4���n��rAo;p��j�X��9��F�7b�E����e&٨�1LT}���ʷ�.���+6M�"�⣣�΋ѺgU� ��<Ud���܀��"�4�nR�a��a�Hq��C@�W;rF�<�CN"_����jo�N���u�s��ǎn(���<���ۼL)��V�\�Mt���Q{�����n��80�i������-y�rI&�lz���E�SDw���!<Mi)��K��Xf.����nQC��N2���f]��Cȟh��=d��� !|p�?7N�w���	5G6�U�U��b��=r��^�m���`#����3�QO�J�j�����s��#.z�:h��ζ�\����$0����Y���R�f�Y%��7���}
����l2���h�U��)��nM:#Ο��S4����JE�<�ۺm��]�9�.�`�wΥu�S���0�����}�̻��!T�$>o	75�DT�x�����Ѥf�@P�w*}���;�(딷��oŬ��]r�P�����Y�WoK�m�86H(��N���2�����ܻ��hG[ږ�sn����d�$eW5��g��.���h�A;:�w�t��\;�OC�)�:/)����ϧ"�1� 2��h���T1�vZ��9����l���@��e]@I�H�6�[�eS\��Շ���M�R_�g�V��]s�s�2?�������5�(v۷6N8h?e�X��#j��x/	�v���Q�L�X��[���1��xd��ɘ(�jy87��]���h�qG?��L+�{����78�Ȍ���-b��t�%m �9�\{� �c��?�Ts��@�i8.�pb,��t�����ʶEe��W����䍷���ro�+o��Zť��9?��a�2�W���"��x�Q����^
��j�O�O�u	�_���My��9�cיL���.`�%`�8?v�Z7NYa]�������g�(4���$	ٳn��d��NR��=��O�Kʗ���z��G�h��*!�q�9�X��>��V8X��U+ǭ�[����1O��e���x�D�O�'q�� ��W�� 7M�a���(
��1�����;ѷ�� ?-ؗɓ�yyk1��yu�|g!zi����֋�P_̉*~�7w�Y#�P����k�>����%�lݱ�$�����P�#>�b�2��> �A&�(�g���M���W?�� �]�AĶX�
�`�����K�'�M+aT��o��6�)�J�9�1� {�k?s-,*K*�]�}-g�i��4�ת�-�� ���*���2��0��䥒��'����m���B��������7�����j�^3���W�I�'/^��nϋh�w� m�p�y��Jw�!�P��׋v���E��Ժ�]�0���G*��K�v�f̋$CV�9Cn�[��K��D�l�cd���ހa��+"�M-	���S�G'N����˗fO�_���.�t�#$�lE�����^���R(>�;@����4ԅ�XoEl��.�.�O	��>ut_J��b%����|�������+��8x����¿H�T�V��4�9�lJw҅�DT�,�O�ˁ�iE�R��S-��#����v�-�S4��؁Y��c����Lw���O<J�IF�5�I`��<���'� �`
eI��`$�Gn� ���r!���_��@q����|�ɞ�v0�9e]���%ט�Tne�?�B�+��yx$�5������]�Q!+ʦ�K�R��������YE�g�?�o7�$u�8`�<���wt�:�����lzKF8$�zF�E�N���?�,���}���?>�R2�Ֆ՞��������-�����q�C����8��y�C��BI�,g�,\)�tҙCAlb��$�y�#]@�'�bZ�z���[�>+�b�`g.�<�ol���t[�+�$sj�]w�=1WWx�Xy���,p;uD�j� �s����]�Sp�pMcA�]<�V���"O�i�B]:۔��E.���� �RL�mq���mi��!?��� �)aT�axE�&�pW����!a�����=V ���R����;�TWZH�Ep�+@ʶ�9�g���M~�%}d}���i��5��q&����E+]P`F�KS��r~��oٶy
e*7�7x�z�^!x��s����z܈�	/ׁ{�{��G�����\q�W�����Vd$�N4ߞVH#�p<�ԟ[?/�;A`�A9����[r�X�8��`s�#պ��8b���s;o*[^����@�Ր�W?>,����-�&g.
�SGl��1��J��Ճ'\��S�]+� �*�%����z������-y3.���
Rm��Đ��ܡ��w��a��!��^�Bo��t�p�[{,���a��՚�C�c��=<�W&xZ��,05l��u.����y``2�ʢ���B��o+�}��E/��d�{�^kE^���r��o��t��Q+�
�F��[���-2�܎�n���>i�¥��/Z���?�C��
���D(y��nwҫqA��i%%2i�NM�Xz�Y��4`�-|Z��o�A��6|�+�>��iA�U�"Ҫ^�X��7k���j��Y���������O���c��rB�8��lL����(��&Cl��ɐ���V��
��ZZ}�`���f�I2��V0gґ����R�̵�[���Ǖ��>�D\�>w���i�dcbbldz��.�=>Ee��p����z>C�V�_ )�P��4����:r�x�:���Ժ�GWo�$��XAH3z���#��}0uM���[dDpI�a1�������7[h�GE�B-46��4�V	ZO�:�)]o���`���1�;� fY&�K�����4CU]S��!��1DC1�x�����y��(����)� ��^QOm"�2����C�)�:�_1Gy1Y�����Ө�M�`�曎8��?z�2�:g�䶡?"�)��T�9�w�r��KϽ̛v1����V4P�Və�|7��ius�}�Z���S���+:�t-�l���h�;A����Jh|d�gh�ߊ��}dp~b�F����?��ӆ`8\�iC�l�������~�y����?�	�IT@���B��#���+��+�Z��_t6pC������GB�q%��m�Q�$���@Uv{��#>���pA\�.�Ƚ��1������=[�]�c���-�,E�Z�L��PC�>A�0w�V�S�~wl�tH��œ���0����e�v3FJ�-��|?X��������E�v�t�q���`�p���@��U��T�n��>ƾ�}R3�=�-����腡�����'ae��>��Ҟ7$�]� xÜ�yM�v�c^����6���\���?e�Ȣ����y��zD�-.���A�g�jo�Q��|̞�!��h���ߛ���R���կ������t�BP�N�D�}DV/U�47F���|�&�C�P�ڑ�Q�"˶J�YIB��w��o��uD��g�X��A[k0M�ǆ֝I�3�?���<
|/����>�a����0����@�Ƽ���ܦE0�����*f�#b��.C�ϰfA��!�'�j�m@�ڽ���E/��#Ϸ��(!0PxI�B!���.�О�����k�S��纕acI|y+�_ӻJk
'���`����>|֋��g �|<(�)�����|#����eĵ�i��X2�%�u�YYXvj��gN+�
����Sv������cx!\�`�@Ĭ5k=կ;�p��џ�O\�S왞7��[�)q��w�� Դ���i��d��S�T#+���{���@]�
�>�G��z����[��LX���O6f.��{^�p����O�/�s�I%���2�އ�|Zn����A�蚟��x7~G���\iG��*ֺ�w?1?Qw~���ʴz�O�iqi4���K�j3~��_c�̄+dտTT�`�%�@�j��nL;�0�65>�"J��x�y0�Jf�VW�1�,=���y�(B<Y�Nc	����!�/���1����̗��h����O\�+HO�z�`L=��qCYC{x��i�	n�փ�5�jN FM-M��ل
��σ�_\���Ԛgd`Y����oD��F���	�D"N�-tѯ�H����I! ˨���U3�j��ygS�|��\A�V��K�	&S�V	�2��s�MH]{�C��Bi�0&�>�q.ϊ���w�%  &X�2#k'��'�p �I�$j2 �K>��#�5��_ȟ-Ļ���!ؕ��������S�=�N�z'8�6j޽*{�NJ��'��]��>��m���X����,�+��������RU���==�0�,)�PI��=�Y5���,h���ug�A���px�>���k�Wt��Q���� ���Dj[B�-�A`8\���߮:
�:ZT_�7�$�U�R�>�����F��>���[�;��Z^�;Е����_e���C(��w��|���������EN'n`�Wt��OQ�=b������1U�'�7�b�}dYk)WC�oI�n|9�ұj�z�|�~�rۯ�>\��7��$3���[w�H�Xd��HJ�˕=1��ZtE�Q ����~��7����Wf�Xs\�OfW�X��&��¦�I��&�N�O�O3S��F�}��\�_m��N��-�&��`]sM�I�m�j��e��!0���}��JERkx�mL����cAʦ'�T4u��6?M�?"0l��Jѩ��[yE�u�.M!6Wd����A�ɗ&i/q&�y>'h l��d3��i��[�'�KkF �X��m��ǎ���	\���D��
)��_��hc���c�|z�+�^a�&��{/�@:�*��i��Wg���$ĸxQ��P�IÙ��m�������Sİ5w�Ҵ��/؆!��?�м3l�m����Gk��vf-��w�C������O��I�q�rI��b�i)�CU V�������=�,%����-7�h��*�NON����a�˔37:v_ �=<�4������r��W_ֹ��ϓX55��f����J��h�;1|X��#�2Z��oع�Ӡn~Y%M�pp .x*�X���3�U�RAxo cǡ2���<���ѽ��!�S���5��w۰�`8�M�p�S �������X�G��|�J]��@?��3��~������lI�?j1~G���r���E^���60���F��}
ͅ
��:�ҧ��U��6 �%7$&X���J2�R�{%��%�8P�Qtx���Me��[�Ș�qD��j^�6�*�KF��/��!zIԥQ5����Rf9x\?C�^���>��6��*��<p#$��Rv[��a��G˿�-��*���p��Lc����H�������!���e�|� ���Sأ�����෰l�u���9�����'6�"�1�����df��֦dcȵ�]��v�l~f�������v��H��c- uS�9j��\��9lZ���wi��q]��x�T�K�����&��t�k���Zk�;���Ok���J��J�KY(B"�"A�����P��l"�&Xbk ��.b���T'.y�M7~,�Tj�Qݹʻ��#Z�R��x�7DF1�SO-ռ�1�WȆAJ0mS���g���<�|"�R.��e�aC�
����c��	]l)�#���+'�*������>	�`�����m�2����a���SSu�d��C��S�B8ӂEز�vo�)߇��qw�櫡��s{,[�Ab�>������Q��V�
�4R�)�e�5Ы-�(j�����=�^�ݙzX��E^��?�4����d�%��0��c12e�vɛl��3��3���ٕԳ��BwJ'j�м����{�=>x���?f"G��Yٓv���b�ԙ/Ukn>1@^�!��l�v6�����u��6����n���+p!󹦗���X�|ݙ��}�(׾2»���H�|I[j��i��������q,��,Q�Rp�ݍ��|��7D�N�}v���|/	�	ٵ�lo9�1�kn5�Z� �+��o�7A����v0}(e�Ǩe[��I(�Z�T.`��+��~�Mwx%�,����r��.D��n����l�}I����;�u�!�!6�;�s�ӎ���v%r�{�6�+M������Ʌv�Tb�2��9*�N����z���Mu��W+��iA�y��W>��@l�^-�.�D����6n���yP�W"��!�r�6��T]a";�����aEqK�㚥xՂ�e+4�$� f�4�ꄇ�`'�i��T؞������r:�Vjl��-�|�9A)l�h����X���-w���	[���uT�������GO���&�
��tX1��z�81���� )<*L �]��&\p8A��7c�>�\�����&�@(�{数�1wvr	���*�%�aP���G.3��FT���D��a�4�uv`��5����|A*��iG��%@��z��fk�m��2������B�����)py����x�_�!_��_e@N.�[����ʃ2�puئ���z��NՑ�?g�f�}7� 5T	b6 v 9�^��!��G9�vi�0�M�	�V~}��K�m����i�~����U"��!�"p|��1Ǆ��;.:Ӳ��+͹ݥ�՜#B�9p���VqO���+:	��V��З��R���O��;,4��^�O	ZGzQ�����f
�44�8'!��֬�i8m3�8�au��w�B�g= nT�b�
��R:Dꔯޣ4���^��q(h�x�1�Č���si�q�������7pAa�0k���[�a���#�o�� �-���_�:-�~|���f)i{NiJAeߓ�ö�R�h�uę�>Q7�>��ۛ��J0�Lq��:�f��	'���g�Ps���������?:~��kR\���P�!�\��LlF7NJ�6���f2��E+Ntb�R�p�Ij��/�ual�6䅢�!��ѷ�k�e� ���*U��ٯ��v����[u�7G�g��n���,\Uf��͠7e!IE;�6C%"A��"��Iވ02��<�U�M�U��M`/�|T��9�{���]+^k��^��;�:��a�3r�p����m�W��3�=#<�_�*�r�{D�9�IᑈWb9��R��2�'Rm��{a��O��$�f�wfmF�2B�\����@���m�a\qD�n�Xy�~u�xE"������P$��!���6v��Tb�&��=�?��2^<%����O��/7��Ǖ c^��ɚEU.-�G"T,��'q*,}�-xp��v��T�c�p�U��	�_�U;>/�����`��Qs^ԸO�
��shI��b�v��C]j��\�1�+W��Vs)���P ��p.!���('ct:@@�pHY�3�0Dȁ�(��8g�������R0e^�~�/=��pT�4�5��Z^�*rV�����Z)!؅�N p��MK<ڽ6L-� bG�d�lMxw�6&�k���%n-�V�碵�c�Z3
fWt�V��{kA�u�s��f�5��a�� d-��$MI�`�@O�>�΢ڃ�:�R'�����`����F��B!x?�U��D��H�(ep+�����4�1�&�(D'MȠB�궕�f�d�kL�*��g�&d����᛭�vt�!^ʪ��?�.��M��˝?\P��:�\M��='�2�R�EnZ^������.E��GGf(���`�F��"��;�[��9��X��U��p���q�
ˣ[���qL>\�YE9U�=&��ˬ���g<�a������%`����p��Ig�{Is��?H�덿�:ºn�yc�J��#�B"�$�V�x�2@W{�q]Ӹj�m�R�喇r<`�JY�MNUr���ۓ���i��S�~E�@��M���q����jY1���Qȥّ�wc��f3�VåI��������g��ի!������?}�`1�d�U�KG,+v��������f*��ZP|���ұ0r�ă,�l���:&�x���Z�P������\ ��P�Ŕj,HƇ���Q��'�s~5��ܰ�TI;g�~���r�Q�V��X��څ	�\eښ#��H�(�s5����z��Oz����B[�TV��鍰�6�����HO��*��Ha�V��w�0�w�������cX�Or��U��58U��%}# ��	�/������ۀ���K;>׵����:�C%�ث#����	�]��ׇ�ihj��tv@5��@���I�U�D�!��-;~�P��c}<���V`���@�s1�5�ōJ��?�K��|�@L�No�d
���XN�i���g�,8@�_G�<"�#�4��\���S��C���L޴�� \3���������!1�x���( *늜�RƎ)�4��v/6es!aq�d"����-{?�N��N� 
(����鏹&؋AV2�n�g����X1\w	��X�塥!3\ކԹ��vZ!�k3���n3�HЋ�;���m211˽Q�[-��T���-�˯�]���!����(����~�(������@-�$5
[5(�d�q�7���O���C�'��
㼰6?�(��M�6o���a�Ԕ������J'S�t;^�u�Z�/��=�֓��4%lu�MZ����(�u�ڮ�.����+S�YK𓦗�6#����5�h��a�51�(�1�XMx�P���L����z��Ƶ��T�Q
���Yϸ���B��������� �j�U�oP���\b�}���n���qޓ;n�x_�5,J�h>w�[H��+�u�����ߡ�(��<��B=��.�[Kr�_�W]�vDdu���	���-�Bt�V�qQ��T�۟(H�`�Xm��������hn���btE��!��rs'l��3��5��dl����Ԇ�x��zq̇�?m��H���2����t���|����P�������j�����^R��djw�,ur)�'�h�~��8�[��i= ���f�Ve)��̥�e��L���!���*�/�`���#�vG����(L5U�3$�ƅM�on)M��U�3��_�dJ=9]����%C�R}+��_#��qp5j�q :�R��f(2�V����;��D��w�k�ン	q0A���U�����90�[$�2�����J�y��S�&�3u.����'dx�-o�E4�s��6=�נpA�������ii� էϱ����$iL�E![>���
�ܪ�	����~��F�X�-���񂯿p�����ҡ�/�{05��E��A�{��lE�c$�y��g�+h�lz��*���G��:��d6r��l?|���qM�vř����M
�&����>-(��!y֞��^�E�*<��t��m�b U�������w��6V����4�� �f�zPI�ߊ���r���ï��g(�>�	�N+ì]�}Ҏg��kz��A��N�J*��uUФ
Aur���q����LV�qX��vj/�{/+f4{�l�Y?��4���[�U���~�����f��ȭ��9ĴB�s W�����+��������ߙjX����*��P2�ɍf,��C��������ݶQ=�M���- %yd��G�0ر$�-BZ��2벦
,�\L��bE@繷�z��"oTI����z�}��x�}0�������b��g"7����5]����C�M;m[Y>�Y햃"�bU	��q��T O�������M�7.n�7��������D�HLG�BX@��?�E8N���3r�]���s�r�.����N�K*�,+m�ٚ0`v������C�1f��W&�6E�p��-����3�>=v�bg�����5�@�w%�)Z�_8�de��чm�'dX���{�&N��4�F�#o}�?�>\�8֯E_B=�9F����x�#�ֽ���D��S��Ŧ�O�����QE�s��6�-xm�,)�Y�|K����<R��,�g
��{���sY?x	{|�i�y;{�>"}��ir�K������Z�]�����v���$,y���<�9T�~N2��<�!.�&���a��Ɏ�����VT�	5�,�_ �7�k-��$\��߾FI7���g'�
��|�����Ku@���P1�����_�ǭ&h�I�DD�_ڄ��!ʝ����翭���t ��u���t��FVΥ8��ܯ>/]Ci�1�8��FƊ'ed�;k��:���/=�c�E����g+_����W!cf֙'����9*���� I,^ݞ��Q�f#!_�Q̙�+��fۯ>o�$��I,*A��W`��T�M3���/��c	�ڧe�g���Y=2.l��7K�v��g��9���
L�եj����Ãou���EA)-�aA�^�D&�i#kj����3�Y����!��æ�3>�6Ĉ>���2���ڛ+�����v��t#w�v�1kk����n��K�J����L�2�V�`�g�V���{޺m;ׅ�7TkJ�<(u��?�k���O�z�F��s:)o�bu"�Ҏ���U��A��uf��Y3��oA9������\h�E]���o����՛�PZ}�SZC8J*?���a�Y1��Y�u�$���S�#OPp�a��cА+�k�.NDǤق_���-����*Y����5M��⧫��T��.r��n*J�ʹ��Wd��5��g���-_�W����V�I�C�/�9J*�w�.����Ee���R���B� j.n�ڂ�]����H�e�W�f�4=���a�(��̭�IE��55D��@;X:���NݷmR�m*����˒��|-Ҷ�JԻ<��ʦ��z�8��v���K�$�B`��a�{�|�=(���0���.�hq7�~��C{N*5�����Y2��2�F��m�l-y�������2?��`�����Y:�i�g�5�y�+��o1�p��%juz�Q�Ҹ��$:��_8v�� [���H�N��M�̣LG	P��N*:�5Y�M;.Ù�,9�� I"���
�8�6y�؎��h�|.fW�Se�\�.��^![<�>U�Q�_n~x��i�1,�,�VK�cL�码�r
�"=/3���3���U�<���'[��ŬNGH�9=<#t����.e�7$@�֠�mm�3ˤU"a+��<-G�rڛ8 �Ӆ4V�d���ᏸ�?g�\�EjO�
�YT@s4uf���en5��)3i������p�4#��$�Ю�e�N1b�N@�N�����Șz ��>W�_�.S��}�ٕ��%�W	h��zpI�r�<{2r[�f����{jh�A����G@E�bÃz{�;���y���h����f���E�q�������q�t�8x$�N%��.O���18g��M��
8�S�i9#(�|��Z��䎝�]Hf�g���f�M���>�K��Ty�w���Nd�2=�Y)�"�i���:3��f�+w70��Dv���_P\�E�7J"�Vm�R{���%�%���E{@k����=�m? ������&`�-�G��g^\.����o�/&��c-ly�7N]%6E0��g��uuq��U Az��90��$����ݭ�oܧ � B`#+�ޠ$�u���77{�`a@Ғ�Hj��[��e)��aR�ִG����%��X�q������E� ���;�;�&�*vD����X,|.�CX́ʊ#���"]�_�3u>����Pj 3��Ή@E��c:s���8<MM�D,�ܺjYm�,�K���,/���б-9B0%��d���t��{[����N�����t�T.^��3��dS��h/��~��Y�l���ηfЭW������~�nu�!��,}�����32��.��V/)�����g�+؇(�y��B�9�S�W����"t=Q�ُ�{��A�+nOJ��ͫmBV<��~���хl��5�U�
Ld�R�_���'���8�p��d8���ׇӰ�II��ך+�1�e.3�+����̏��)�,��˜�e�Ԕ&��V s��;5]��_�VK;�,��f��p)-�yLQ�*"ǯ`����B��K���:/�	x�1~�����?au]���\�s�$m����a�³]ӟ.3��%�8���D��N��G���}Wc����L��P�w��X&y��d��m$FZ�3��/%��g0�@�n����2ܫ-�Wh�E�����r��T�M;zL����{�`,���8�	NF��`������ys(�i��+k��L	(��t7�QӜ��U��� �(��.W���P��G����Y_<���B����P�U��j����x�d���(.c��q�tD�I�<�4�e�HN�����5z��C8b}�+V�O+��T-��Y�+�����������#~4(y��\&��e���@7#���tC�5��Y=<olϚ�;?ֳ%�Hu_�߿n���w��ɂr�C�D$���OMN�f��0�]a�6^��)�!gU�&��,^|A�{��j
X\�Ѝ&ӱ��Tƻ��_
��g�=fE�t��)��@>.��a�h~9G=T�A�l�)����3�.���6^�N�q���k��?�l�ܨv\�A�R�D�_�h�M��H̎�R��q��Ov/��/��9*�w�d��Ħ�ٗ�͹t�w�m���IB*5@�*��{��̶U�ӓ�F��_�z5����G蕮^P���!T��,;r��8��bmP��k,���1�n1�(nƖ.z/j,1įOw��N�$�I��ST�$L(|�RHc����
>���Q�7�^��W��{���$�'�=�y�X�Q^���S���n���0������8.��ɧ3/,�ُ��c�c������]EY�Y%��.���wP�ԭ�H��V[��"�V>���S�#�| ��1��<�~���)�M��,�T�9,tr�T���Y������H��m�� D��0i�#����j��=�~ʩ�t�_Q$���c��9�sp�F�W�7�� b�Z)�n�={�`�Hv�;��|&�a��i����;K @�kR��& �"��u�J�i��=�;�4D��x�v�ρ�-��/���A^�M�QNs<�����hx�'���V�)��@*BJ�������y(�k���}"I��?*��h��߽�R��*�^�Sϻ����tb�l���2Qهc��<�}�G�s�֊
�X��b���ot�#�9�3�] k*o��E������*q^�<I��Q��+���$>��SPe��c�N��J�D�%���ң�HH�.�/Է@3ŉU�p�`,s���Q�����允���N:T��r	������S�C:��u����X6}��K�Ǭ�;[ȶ`ǘ��=�DFM��ųd�!Ar���J�TA�a�G��Iˮ�q�\ml��J3n]�Miɟh����df�Ky\A�NL�If�w'VvG��h4���.��B��aB�ŕ��^.ƚ����a����dЯC����"���"4g
�QZb~:��:�=N7��	B��Kz����}�^���X%O=B0�*�V��b��sYA��3�E���0���4�E0r|���?y��_��
0 �z_�k�� f�^����9:�
>u�$`��)�
9b�0������[����6Wwмa:T��~1Zm�Dw� ��I��'��� ])�n@����,~H�UCQbyK5b^�h����I�:�J���sK;�}�?���R��������\��x�"��7t��ظ��Z���\^aFiA�-��C��g��_��WWCģ<�,5:=��Zd�le.�X����mo`a�e��.5�(�ه��B���{���\�t���@�[���|�#`r�%�׷������^b�w� �涶l5g'_'�EF�h����"]��Y�r}s����]'E�½1m�Y�ߚ��w٩T�0o-�C�mL�YNE��}��PBXL��^i��<bJ������pDr��n!}�����zn�Ujй�@)�Ӷ��U��+��7���=�K�c����1q�kY�k4ߜ1��K���NĘ/�&Ia#�v��*�+Q��M��d�t���LX���%P���n<ڠ���Y���.2u �K��wB��-�qq�8�s�ӯ�H���ش,\̢�=�м�F)8r+ׁa�v�����
���F�3A�]C�L�:�@C�����}˗ �ݓ���^lYf�p�/C����՗T��i�#B!a�Qȼ�Oz���J�_eRS&��������h~E)+l�2�C5�ΰ�Tj���)�!5�$�[�*�1�I��L%�����[���hNm��v���3�!����sE��FI,�Q
h��DMu{J��b^�*7�nB��`�$�l*K���=�{�ھYj*��wr¬z�9��M����r!��_} m�M,aiaۮ����g�t������fgm9��bz9T���Kڂ.����
�bC=��<Z�� D�E�s��	.��"	,m˜����*	=��o�s_g���� ����ye/�z���[]�o�X�:a�W��X� V���;��ʇe�>R���a���qSd��y>�N�~E`m"BU�KzZ���E!?+Xu��E�2����Τ��)K�~u Ҥ Q[��,�{ �Z|}kpKM�h@Zw�~���}�
�����y1��WW���.���(rq�f����ER�/�>X7U���*�
���ꈵ4F�cq��Db��]��. #�J�^!i�3"�a�V��߼�yk�r�S-#����P����O�E��i[�)u�M��ij>!]ӼH���G��W�����T�
!J��s�x�.xf�"��O�1t��57Y�����Ώ̭���᯶���͑�R��y[ m�Ӭ��2�ҷ�@�;��Ua�q�	���\�a��Vi�Z� b�*<,�>���ݶG��['����vj�=R�����Mq�x�u��=!=6��o�e���PJ�)_��f��V"�9�Cv�i��6{��C�/ <�v���Kl�[t3��<��/`Z��xtS�D���B�k��2��?���H���R�P����u�)#2�5*h��@�w���.J�qoЍ�����$�*s�^�S%��j��&3��O�^}����c���%�z؝=����_�y2M+U��hn���:�]��3���r�t��(��$��N��9�V���*��Q�L#�RA�6.��wxG;������C �Y���-��������qax�����Z��n���J��ʖ�`S��qcH�)U2�+����ǥ�~����<oLl*o��%���)CTM�S��Cȸ���W��Y�m�֫��:�"��ٰ�£g��}�}�qiq�U҆��-��.��-�@8����ܥ�H��0�ϩ��޹�����|�+r\A�.|��yĂl�Wl'�?N��k��48�Cc���J�
h���W����Ce7�Hǋ��	��,�#�5����*#��U��
c��t2�-�-Ϩ���&~�O�k�P�����@��$W�S`3/��P��י�֥L[�?ا~n\"e��"K�	-R���%��!���O��F���V��U�S���ٺZ�����M
$�0~����=c�Ԭ؊��o�.u��Z�p�oj�,lg���-�h�1����n;�u5����Xtt��t*Z:�2��¿�H�p2��-�J	�-�{��G�����̽V�dc:�x,���˪�<z����cu���VY 
7�5��x!���]����݈�	�E��N*ͧl1�2}Oz�	H�:`�J��(S��A�/�1�d��*�7f���ɀ%���@x� �Yf��ð�	'�JM��D�&b�%��_�R���B�Dt<xGŉj&[�țs��3�