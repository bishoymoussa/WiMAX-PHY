��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$Rx�y�<��wA�*;�x���@�̦?N����~�ɌZ�08/���\�K�}���a��p��?�����>4*�ǚ{�����BHU{L���G�bY^/�Ԗ��5$
�4Q�?�4�u_����6��|{f�ɸ0��I��8q ���p�=�k�Ws�lAVP(��������ܸV����{�[&sz�{�+���#��-ҙu�v��s6ؖ���<H�sAU���\�*�R�]�x���MM�*��b�{��6J��\��ĵ�[+Aҳ�-v!�]���}>�~�k|+�T�������u=p�3�QKi�Sc�t�~[��_��ן/+D�i7n �D��+�د����&`lX'uL�F������LӶ�vT
���m_�\{T8�c\���z���	/�|��m�(��_�iv��Q,����C�s�1�"�]6\E�#�!�� ��21��@��[(���Q�����9��t9���v"Q㔘����4o�yT(I�Y%���ad���Ҵ�swlC�ɡ��ĕ���r�i�im��}�Q�m�D2l1Y&Z�?��"����-�?��ZQ�9蒣B� �.d��V�sڎ��֘�T�PN)}���#��{s􎔓�U�I�E����ZM��GcT�4%@�SU��42�(���_�=��P1O3$yڷ|_���2���ꆟUL{��x;&����q��L�@�G�sA6-XZiV��XEn�{� �E�z��o~@SphMk,H�D'*�6M��bC/���Q��R͔�yWe�+ ���-�=���]�saެ�T���I:_ܑ'D,����G���d�h���a��k<��9�\Р���p5m}#�#F�/�r2��'�h'�,$�U�='�����+P&���n#�uߡ�-��qv�X��j�J-*���fĻ�5n���$�"�p�O��"�z?S�T��h*ē�l�	e��-C��_�br:����� "��:Ǥ@Cy+5�s��"�ܚ3ui� 8(��iC?���O>!6�!0�y%O�~��W?#��9D�y1!=���5��E��&�Ev��A�a{,�}_K�x�����BPֲ�{�8�8��N=���:�)/=8����6k9\��B���Q_~�o	�Q�{DfmK��â:�j����w\F@>0��~�J4��d�}�ǌ���[��^���P���P�&>�`:�Q��+l
@W	�Ӽ�%H,r�'�q;�e��AW�=E�A0�d�q��� �N�B���w#.K���Zr|�����Dyy�Q�'v"�u�~@U�7X!Z��j����w�_���E��w=��h�y�yɩII� H�CW���dwႉ�mbuz@<��Ni���,�=G�<jmgl:��Ę���a0Cb��z3�s!�FԒ�h&Е�q/��8���a�Q��<����Hr]�_L�~7f���P-ܿ�RyhĆ��P�Q�����Yay�K��%��+̒ak�}H����P�V���Ӳ��ɿf�AH �3���=%h4�J�Į\�3�>�W�7��m`W�Xf�4������g 2�1�YhKz�ٜ1��`�y�)� P	k]��.	MČ�uXa��M������D*x\�N-u�$�I�³��+;pJV	����d���D8"D�L�^�}�n3�'���\�S�X��)�����̻�ȧ>@�a�AK~`��2u����:sOx�a{�I�Q�W�ׁ�_����D[�'Fa��o���'��5_��#U��|�����!ō�F�u�c5�Eu�}*�k\�a�Pw���P��j�8��_�kKe�gR��!��k�?�$�<��0L�=Zg��]�+xC@��֏�,u.[tF���c�z�w�1h�(�Dҫ(�I��x�ιA���Ch�wQ7U6�[��cPΒw���Ӏ���@���!J��&�]JՓg@��"�3����No����SXE����Lx9s	�}�+�A�e3w��>�����k�pB!c<�L��G��0�
o
����@O��	3Lž]�f�PD0foB��qNF/��i�[����dV.�z��{|.I�
A~�m��ު(���ƸgQ�JG�B�bUr�vq2c�:�p�3�[�cl�8K�*ŲQ����v�b���![��Ac�����ؿ��c�*z��#���e���d�-��	�}$֡�]������A��^��J/�[���k�
��0�>�@����ʀ�ݪ�r��Ϭɭ��x�٨Ww3r�����kԀ�}�m��Cjd�횭��^�����<���I�i<��_fR�EE$��107>�H�^/QM3���crwyQ�ٻ�?~�/|{� ߧ�0��{ǽ���fڇ��x�f��;�wum=��i�+��s�
����|���e�9�u5�S˄&*PB!k�x&�M*	!D�[�;y/���������sQ�z��eM4�	�W|���\Mz���A�g��#e�����+ٯBz�~ta�*ɧv��������V#���+O�#�9m]��vq�Ws���9��m�c90������Y�Y~&Ȫ
[k�P
�Q){��Xf�����]���v��&�-�|32��a�;4���Y_��H	��n��\��!a��e���ձ�@`�7*.x�ȭ�Զʵ�yS�u�w���F5W#�^,�������u�x�Ro~!��h1K�4�=����l��l�(��3��Q�j��Н���8o*�h<���x�:��QQ���@[��=�����SփG�|��L@��w@��W�����YT�V��Za�|`��Z��<M��v�h[�2�k��ٌ�k�T��n&G��
x�JՁ%�_<�Hq~�m��{�S���u��{O�e�Ów~��آ�7`��ߗ6:���:6'�zD�H����@`]&识��dޜKy2���V&{�'Myș���ZFv�n8rUl�'Q�^�v�1;�[��ЂF̮�֑������?j>�T��  ��	+89�g�d��*��Mr�;pÂ
x�;�~a��c�hq�.��w_��ZX�1�P��~��%�8
�/GΧ��J�j�(j+�b�	z��h�S����V���T�����Ϸ|+��������~nn��t�7�t &g�>a��&�7�HA��<�_����ϓ|&!&r�5:9;�k�����,�u�忮�S��`P��X3�K8�9�Yv����\W�޿ow%���ܜ�/��O7#/vE=3�����RM֣�HFw�����-� �/F}#o�͊����-A�M�V[�_�gfo�iɓg����
t�{�zq
C$^��]~�V#?X��K��dkv,�e�o2�����3�������HG[���E3�t���r��%rA�@���⒛"�+��:�2m\������"eT�;U4D�V�&�S�dJ�oY.�0~�����NG0�k2���ҟ)j���U��W���I|2�㨇}��?���%7W>N��"�C��5x�:�9&l�z�Ӈ\��ř�ĢROǶ��L����)J_�tN*�d3E�c\�q����te��օퟙ�ڬh8����H�=3��`�'��]^�D�/K:g
'^�_?l�*֪�@ �A7smA��&U6{�B�Ѐm�U'�t�z�m<��?I<tJ�cV&���39M����QYa�s��W�dXC��;�ϔ��BUvD�b�wm!v����ԕ�J�X�b߁��"E��+�*1��tX8JB��%�y����b�K�oe	�����X�	�x�H�K?��咆�O����e�|�y�h"8;p.7	�r�+��)0��6��^��n�_�������gJP̆�ə�������yː��G�s;澳^�˹/�z��U�,�`�7��+=����V�+o$�q���2U4��f��B�?�U��@U�ERTX��T^LU0L�z伫ed�V���w�Ʊ%���o�A�F@p�s��Y'�7f-��SF�$dr|%$S/;#���Y\lID�;�{Ǭ��Ɯs�t1";M��R5I��df�p�������Ċ"f}6g�-��_�����+�y��/�ȓPG�6��=$6os�v���*:�&�HC�8W��J��2��X�Dݗ�4��v�����O=��VPr�k<𞗯��M�� ���U��P��9�٧Kg�B�"������ڳ�DS�ݬm�ԯ�-�x�V<�	�Ɩ�.��s����������2x� uY���w�+�erV��$ 1ȟ$�946L�]���,e.�F�"�d��J�R�0W����8l�����d�ճےO��m��C$)�>Y�����QZn��E�MZ�\lA�Ek�t͜�����dp�N�͠[�]$F�?���m�C����ն�&*�`����Y/�i_Zv�����e}��;�ȫe��8i����`��u�5)���Y���3'�:����%���0����	��}�G�����U���(�)��=M����{����'���#��i��=���޸cW\=��ڎ3����ZL%�k�gh���M$eӱ���u��_�jE)Ycz�T��R��Jy�h���h����҉����I��|fIO����s�����ڻ��̀�J'MaZD��z��aM)6l��JR7��.�!
�͙X��nA}�i`���3w�IsN!GyL�m��i�����Q��|�t�y�w"���_vA���Jt��K�Z�~d��֩�
g�fU�f��cܸ��c�[�"Kѩ?������f�<�Q�<���E��7g�"��Xrn�{�E���me�u:�ܦ�$��T[o�s�:6��Ps��j�\D�Ұ�6O��i9�
t{��V�F�v��o��Qo�g6����F1�j�¸"w��ٱ��F��s�>dj5j�ݧ� "��x�8o��sN5�[W�W}+\��
@�e6��?�ֲ(���cN�Nw���]�4ͬn�Hm���)����oۺ��L��IM�v�nDX�ݿ��ߨ�.9��wc*�DXSsC[o�$���S��^Q6��^!R�6{*=fP���Cq(d��.(��B��0dq�k^0�hm�t8�O�nI��n�����~Pö�!|q���y]:x��3��+k�,f?����k8�`?��8!	DB)܉�S$���)f��dj�
i�sKF4���DX� ��n�m ���$ly�$�ǥO�>�1�3�����A�M��9n��f�!��T�r!>7�sp\���L,�o�*h�iӮ&���<��aI[��B}�4��E5O�XN�e	���� �K<�2���v�u�x� �O��gmY�ii>���"���-h�7�ap2��wT.W���p���8�3���؏��x�/!���Z�s �R�
% ��F���K��m�$j9/�\��fT|�_�d=��i�x�@��T߭���j}�)�VP��P�q�A��V�;�cH���g���]��T�j�_Q>�Ԑ�~�&���I�7�z�4��R�M�y�W�"{�)e�b����h�ֱ��b�U�]l���袅}��SCOb8 F_JF�B��P��U�vzL�'d���%���b�4\I
Գ�s��ړ�7��hɻO
G8w(�-w����ԡ>�Ey��}RCD��;'q(.�V�{�jپ��mՇs�o��I���{��1ρԒ9�M���2��(�2�)�G,�❜�\T��>M� ��H�z��F���O�B�E]���2��'��m�४n�&�_��z��S��$g�DP��G�b�o��a�]G�9n�� ��9�q{U���+ G�i)�ӏ�XO�@�5*L�C���^S%�����Q�x�oD�l�v2�2�6��<y:)�,sM/���_�;5�"�����;��]�,��l�r�~ ���F���a������;:c���^��
$?l�M�*$�t�S������(4|m�N8KC�3T��vB�^����mB��1���}.�},��?U��BtqǓUS�%
ldGE/:91�}���+��c���2ta^^��Lij��˲/.0�#R�-^�K&t� �b>��Hʼ�B��yR�}�Q�����Xdhlf=Jk���#�	�/^�#6�W�����Z5����#�*�좍J�1T�4�����7�h���N9z�y�՘.�����;�r��S�E���#s�)��-���E�R\g�������,�Ң��A��r��>9���A
=n�"~�������#�rT��^����!z@|�Wn�'�������c�@1��uӄU�^t��M���z���I��*,.��S^�<��aT��g�-�d0hJ�Ь4�6�cn=#̚"P����0������V�䵈7���٘l��^��l-w#��K�m��o�ڈ��:Qʇ%�,hX!��a8�.�j(s��3�[x�F1���	F疽XHa^�	}>p�$�b�р�p0GՑp�����Q4{�OQE�y�խ|��AK�Ar�t^T��'S����kO�%�<Z�<_ö���S߈��*ܒ��?ѫ�^_���3���h�����
�,���Y�Jc1Q}�B�_�^/�+@��0n�eK���Es��9���,�u�a��������c��?H)/+A'.d$�=�S�T�,�V�w���~x�����H�(4m:מ���q�kmaa%�\�����-a(s�"TMp���Ӊ)��n����H���7��e-��V�Z�ު>�[[��Q.kkuT��@��S��trOk/U���co��$��բ�4���y�u%�I��]w5ýc�t5X�[9(hHf:�/C%gi�EF]��� ���S���7K��:,n�!7<%��d*��j�肯�~h�7���[;426'��5I3
(s�d��"~1�y��V�Ԧ'���RX��F�x�E�d1j3��6���+���^�C��}��P��)�T���s�
5X�ɱۑ���N?��x戃3������	>wɔ��X�vI7�.DM%t�}���e�)���8���C�H��zQf�f�e/�HaL>�(y�pen��"E�dy���xj,T� �\�1{^b�Ʉ8����,ȍ�<-$`�Y�`�EOCH�6�o�|=�X�$O�F�h���P���n9%uC� ���5W�v��b��e9�Z	���cWֵ��w���GF�)�]���t��"�*�&�r;T���nT��ߒ����ύC���Ԟ���;lﱇ���K{R����j��NM�!��W�<;)�(0G'��1�Rɿ�L��)���j2�IR��� &�B��EŦ_pK��K�a3�z�����x]�Fs���3�c@t2j!!Z�B����%U��.0��O���FRZUE*{�ދԭ����/�p_�f0#��x���m>,#E���F$^����+4�[@P ��27^��$?�O�kk?�'�����	/?�t���� �3��4߯so4�E��Ɋ*P�ǁF4��Y��Y�.�D��	��m��	Ey"{J��v���X���� �^������
ݷ�c���J��`]�_�W�kۺ����{��҆��7;L��Y�	V�-͸�� �����A�せ_��(T�Ė��$� �զ�