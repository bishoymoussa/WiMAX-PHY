-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
ZfFRVnvl1zO1vFKKTZ8zTba7QpsNf/CJH1m5CZsilqub44aSc5eWCCfvG5qUI1caqmLPV6ux4TkD
2Fb7YIQ1PlReW98a1cmv6JkbooTmRgGo3quTW5itk4qHHiqkAMxpC82hMzJG1JrPbZ4zSD1H4oxw
IugHpLP27A/WdOiBcFvpaWvwMircMxRxI3pTDwVP7K/mlrtIotAgH4GU0663R4ut216OvnIQs4tw
c7x10by+DnwAGr0jQd58pk9hNlLmwYQhjtY/beINbRXPqj4pwiqMWXdje2d0VN46inhDUzuXBbvC
ARFKfXV3Fv4NI3fEoEtMUlKikFqN3bJw8TbdNw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4672)
`protect data_block
+lX4phCrrcUnFRFfMFqE8vLYAWVr8HA+pcAvRWDWaEl5QVFQRvTfvM43Xc07byqu0sBlVdm2sNHk
aAj8E84X6ETMaqucHCo/2tExtFlqODSy/hteKGBM6JX4yLdWRnXzVAcKo96mktzF7/Byo0Pb2HVs
Q178SWWWm90sZIAF19IUgAV/HXKXErYIKnKNwmx3sD72C0Q5G/ysmgCEbHlfKQspgwmKBvVfAriF
bsP91eRRqO9hC53z0FQPCumTVL92EEt+Qh0gtQInX8vDBqQMNxOKqqsC6/BOjU846Cqyz6Kk1lkg
LtPl9tNo2UFiB9KlHPtzHTEmvmy5D4HMKnxNJ/rFvPDPYSW8+E97NGJd1EmYHNsxKPe2fPZzRqnw
nY1RopeWlZH9aafCF1U636Rh0ZAwnhZ5gks15a+FMQX4ic/YuGQESDRq9VM0DKmHaphZICfFV5P9
bB4R/7bWTs1tN1sjFxdwDE034huF99R8Di7pXEAJnZ76Cgy7k09Zy5svMjtEN3Y3RsbHpxJi9vhT
G4ADV4D2f5Hv/u31tUbFMBFERqG83GrCST6XEVbeKLRVO16vxwPwOJdy6cnDyRruPmz7NPI75sXJ
qboJwFce8kqaMB4QNPWe66YK5Df0866c7PvllNcr466a0xSNchyjR1D1+eR6fmNU3OWM6p99aeme
3ExaG/A8vUS6c1r9ar5SGnPE8lfpKYKZCWuDzqNMM/XdINjoYtS80tsHHvtTx/HkW2/2zdZWfHiN
rASj5wKoRCfxy4YbRygCxYJK7rz4xnAzRFv7688o2hCkYPPU12sBEdaVOgZ5DiCBxjmaclZTqnYD
eAXc0A8JHmkyGFdFKDcupe0sQX/75zjWAVSL26/pW/UCJQCYy9J21yxmGFVI4zz2jAbqUWNXhz9g
i5W0nVKibW2gz5QopWgDJO00sU+9OpiH9a21C5HGwmZost1f9UpbXBHydcvbxm8xhnOCC4O1fm+7
ilw380LMlqP0fUSFnVkXjc7vL/pr8jxsBUS1QxIrDu43tV0RclrNUZaThV06wXvdjveFXA6d+UOT
6xboiRrgAGdGOB3YIhL10Zwhx/MywaJlOq8++QB9GQo0OLPM1E3FQZvruPRdeBOOdxyEVC5MX7Pb
GLJ1ds+HgXU2Fr5xh9u+zD6+nlHvok77EJyOqS5qenwIkt90eD4wrsruyB45ULvcwVFNPu3Ka+Oi
YW0UWjv7l2Q94jDPvhu+5X/pfEUXq6Qre09URsuLPJ0f5i8Vze57H2+nVui0dGZxSvTR5xcL3SCy
hehjiQTWZh2bRQ//smECMwwivGE7yTR5CPNl1A2HQcAf445zEzxc3BO0xmwTi0AJli7UbZcEoA9O
GGd4zUWRxpALqy/8lQTYKXfUswpxFrrNZXyDPxVoxvwHuhwAzZDDb2IOwdDcJ3amy+lN3XHpok3L
PhRm/JWYfD4TJPbT325553I/GAmQkwd/mKanRC2tsOE5pwTM7Fvlf2FaGDbDBU1RoWWwgt+vDp8V
cpVSWetKnirmQ9gGPH9Kzh6F8cjZEaRET9NzZlGqAyK0VGA0OgGMrzzfMavuxwzmHOsnnnbG7+eO
76Q0gdhRCtyS5uO+hIHt5eMFA7FZJGpW8djZEbCsLejJUdjDbbmkEXngN2MLC1kqfKOXNCIxe81r
PLG8Wf0nBb/epQ43+yAAU6jmv9o50oGKVHX0e6RErpAStFhsM1nrAs5pV8roeQQHMMmUHbVcwPMy
OXemt+uK1brCOjw4ft1EAQK3yP9DiJA/sf6dzktcXjDbPIw5rrLTSRkD4uzOS9dzYN/8YOJ72YCe
hyfkG5SzP/HOnCMfFMSXIUkXGWZownr31NL+I4aHj3sDbIhUrE38MMbVb6oXeo1oUiR/HN5S3vHk
VMOjy/WJIjomlgzhXJ+wjvdTlcg0idv9nnERl9NMegSFJAhT9ym6GtSqotRX8/sLlrwPUulQKWVT
ZmlZ4o3lRDTBBs7jUHqC1WugOkmSLACPVr53jnC0+upcKv4QVeDPMijM7qBOPdrbzFW+Q2l4fi7r
dDasFhaJjy8Zc2+0nzgZeKwwoqJSaVgHxa3kWbIKHHuTIvuSiueA4qgZQDaOBlyHGGJMFx2mPC4g
7eZe7rAwoWI+0aOBZjT8e3piBMj8FUqv8hE+M/s9mXF7Sj0iu1dtq3DlD2M6oaLLWyAaPP//iSqQ
ScWFNrtGA/EftUEquISzDCGkpFILiyc584VYSTZPxWr3cQddB/imusmeRdXPKGX0LqGgie6NFNLM
IMt4jwreUijkzXTUa7UNqFr11LB7vPuKsJ95UE7C0npU6RpViwC+4xL17e6H8ciUhjOZjwBu57qC
bVTCBbUFkJlcSBLTTwuQgbyKDe7pCTvCltkYk2xI0I41+sUqMdulZPLeh0B+m3gsRa7BfAozSEdg
Mwqtl8VFNyGNMaqH5g6g1tq5TyFdROv7btob7w65bQjrcbDZWK6gKsKVzhb/cd3sL+0YcbEWSBvc
OPaabwPB5M+eXywxH3BmPT/xbskmd0AIq0kwYz+M5XEFVW+NRTIQY0YIOojc6DmDWLi2ajkQYANN
r0f2/lYzNQFkGt2B0IE7Po6xEouJfxk0VpL6rpSP1hAKO1PPt5Gmp1WP899orwFsaQPEFa3nBmG+
0Zu3tG9zAnU9vO3PloTqkhPritUqm+K4si4N7jCCV5KHGFP9UAz1YMd98IJUDMZWpFbWfoAKJOCg
0G9P598YZzmvmH1fvN8oMcXiaUdrP1jg/Qk/JkwzReqOqXJWBSRgIzxN83EF94e4DyDJShrW+iua
EaqqQBg2lgo+c+8aM/0f2YP71ZDlGbAHq3UROG5Y1s88MlrYfo2YShRlZDwVZalnPCYzoDfzmLmE
ZQody0VTn6BUXuypVwPf22E1OqMe0CufK4dhraz3+uixBFn7+6IcOh1IQZBitM8YC7bokweJfQ4v
wU38OzTb4sSWThgIrQaI2fhRoQh4pevUj6g6B7fZn6Rse4LY1QuksVTSVnghgmcYUdcnBtnC2Ym+
jchqdiH2sbk//WSyDGBOuj8sxIz+BSD/w7JU5gVwu2sWVTjUPn0Rb7AotqKu5BmQa7Yo3cJ2nZjX
DbmNB1p4X7JBR8i1ag5Qjij/VG41eexp9MOdWc4W/FR6HSimd8QXOssRwqGJLvE7nh8nNWjlEj+U
bWa0lGOV86LzZjYCj0BZ2+nFRPlbjuTU/Xi9XDtS3r5jeWJJtYD+xfaEU8NZO9gawm4iuAowQK6/
tXLzV/OTnL812EMnM/gO62CD5TCpbkK4kq4YeQpp0NH1AfofsMlmBqONHVdYxsBN/UW2EQWVYjk+
p19aRwO/lF8rEnMVRgTt11+JwId8y1pt7p0mexGG0LueTx0cF6rkCBuU4OPV0bM9onkT0jYTDwHR
4b3TqwFD3x+zQhqrffjFxll0bRVBiC5lldhVZsFsUUXv/PEhRGKv9iG7kIIxpV/d1qF8GhSmtNXL
lHEKfZgay8ZPG1m2uPm6eo0SbGrPRH9Ts2u8gu5c6RGgwdN91HqEh6O/O28Rpyt03tLaQsz6fni3
lAfBHOo7rTgsf40WNbosS/BMfXWpFJxBvqR2tK8t0CZlkOeKtsffQz6PO6rQ09hiVhsMF+jOLfHa
Kmc41w9B5zyMPgL37mfLXgX5jXaGtVLDcl/ix1MJIrevGjp0ccrX0p/1GpJrvUQNWvEeAFVeuQel
DfpdG4uvhIElPpdtlTAHn+cQ53IR6vbNDbT3mv+PLdTmy2tRrcL3gW/TMZ4B05WFJS1OMoxVlsDl
uo6j7mTzyyJBcDlbKr82fHVxTwfZpuXdFUxKBcgrIAmSPxpCLGN3RC28O0gMD2mTRWolNrCNfG/Z
VAtPbBvwkssFQveQRA6AglYmMT42kbqIvredX+/Br6NtMqFzQ4c5zrgIYYdc8P15ocSzDHjdx5Cp
+MkIuNzEr0016XjQWmXt3Tdb9pv4Y3EWP/Ixw3MPzpChr7PZVEQCSdeb8XBFKERcU2w2dtGpM+0i
O8k4jMALd8MbyyO+fhwRh2Yd4bb6hKvgsaFUlrk1m7WfFr50wgM/7lPuaTOdMBL/orRqPyQ3tDHc
Sgsek7GevVczLuVgeSvsxeqRUDoaHj7J9N1X9DstA52P14ZrYpyKdrJLaaKWMs0eRhESm9EGlava
f+NsWXW1i7iexM/M2XQROkhbOJJ2bwuo/O4riGpaIjG2GbKeDNwGqW8+7bKHr31Ym75JhEpnBpkI
8GPtBjgaw1jbvjm1hz+myf/rgeo+OLmMilykG/GNrYTqLYR1ofPNDd62eaubhqIZdJVPTLmPh8b7
vB5RUxJJG2At2GKyt3ZooOPLiPHA/plw+97VjRzsoJFECcxnWX732v+xFRIp2mbeY3TSxlnLEpl9
Ip2HvYsR9aOjMcZoxOeIRKFi6czrS77O90uVTlpLv5CUUqSjD9Ii+m5w0YXKfm0IuKWpPG+nwoic
SmjFK1yvKx/buXNf8VZ1BLuEKUj2f6HmO3hFOG8Dy8J+XWZItWqRPFHKQfnfcxXLQJ2csl+HVZ9p
Zu4kXwedGY/MluZR4D31UOMaif4LyFdf0RPw3XqeZPgUon4g9V+BjLbVnxpJYHevVOX3Iht2xsFi
NZg4uMxrEGAUU1CoV7qqHaVHEviiDzVZnUE1Z/386O22itOx/HvP3xaC58ZABaOmroOF19tTLMIf
RbwDEdht5cPhgejju4jbLwpfIZR/w12lUH+lGdiGgoh+4gk+dFMYwCARONTpZizzqpnsk4jp7fHn
HzDQU4pyNRZ/j7SoM4uNA1NSXlXDDb9+xfhqRIDUhovTlE+6MXcE6Ff8Ar7BZiapUZ+A/JAGminz
F20Xt0P1YtURapDwJCvKnCazh7irAAHAliRh6JTkUnIG9eI8otC4VB869e5NxRENXAgnnI56RIW8
y5Y6IuCXK6IbntNfGzrCImC9q29RngKT2VYPU5iEdEhLNkjhyRGkP4asq9ja3D9tNtkqiX+KcLTE
8Z5FSIlc4P+ZCibnDdPunWjHoQhLg3/oAXPWiby6kCHDKoCyDzj7SI+gpxWJw1jratkRmJq5JoV2
oDugvM8mIPxXWJZlhJm7Yqso+g7F0QPIDM6B84D8BUBGCT3jazlYXhvaXzkcf4wT+vxScsI8YQQM
7tTN7QF1gSsNg/8qzVaEhfUoCDyICG9BPfQLx8XQlWNX78eFkZ1k5ofd8vQULwSpDDCnNkzIIVND
XYtxsxJ4rvMyhL+wBliQzWd/3NyHcDzsO5pt40v3ttGk8OlKu3jaVUmEzEexHtUZb0BEkwo/i+1o
UG8sfb3iQc4MyFsZFxpJGpXYhHzxde8sZ98lJIRjqfKz9P4YhxAOUSPsPhsS28/n5z5sUeYIxyvX
zWJorNeDVuINxT8jBGvlnK5o28KQGyF0/9ypPx9ih+PlDVmJk4fq61ac69sHvlukr7Qkp95ZRjuS
x9CIXxWS9gUjFOuRvIPhzaZ23cr3JQch2fUCojMMgF8joiF1jpKrrZm1Wx147ToWlLW5lR0f2DJM
aB+ScK3WmIrneAquxYq4eNBe0H39BmZfk7VDMCHSmqZI7IdGj7gXGtFM5sHPNwb3an4SoZDNJN2g
JVv9eIuvUCm80rAJGUDplaSvzGno5PardA5hneRXU1qqN9H2jwvnwDjMhYj57I4a2S/RQY113uek
a63wQq/RBakqxdLn2IFkCZR62V7Ks9hgmlJdNdV137+JHKXTuM2HdBx5Vpvul3ClIMmvs0bfG+2f
Cyf6hivRVDZ7eVW56wn49maZt3CFwfuhjbymrj3JJzBr2hgc3LD3P2ih9aq0OISMx3e31h9U30r6
qYIBOiA9Am4pW0lnWc8M950xb2lrflnOJKkBeSx4CVYo8aYcmsPa+hx3ntUiiHdAD7Ba4ALHKV6Z
9Y9la2A/DfE8UlCWErAZomy/X/9LjOd+iNENpV+fcJufxhL5IPPN24Z/C8VS/QCkmmBMB2MV+X51
1Ni8t13pQ2geTQUIjPUgIwnmRvZloMCykNtbey6M9RQsDc75ikpxCoh3GwPGaOtgkIZpeVf5exav
BaGe3ixeEHL786hAKrYMungR3YT8i1+YzQZeO2ldmMRKLIWWa+Kzd02c2Cm/O7L2UA9Xbm3zu7Sc
l4c7SOtLxOpaaT55Bqmjk1b+SsPxJTjhup4QlNQWD6rQdJiZyw8SbTpLZM+r7C9ADAhlOJxTMQ==
`protect end_protected
