��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$Rx�y�<��wA�*;�x���@�̦�W�X�fa�M-$u����n~�%���P�$��W��kYَ���P7�?UMfT��q�6�U��k�>����~�\N�(�����X�e���/6U|)�X2pF�]$h���d.���9E��WG��L�X"]�Ad����ľS���8od����e�GT?y	7�������ݵ�^��R�q^]�鍦�����s�ae���h��L��P_���ާ��YЭF���'\��68�b�[����w8�[X��V�F�0͘3����q諵�uW� �h�u\V�?@��_6G�_�*�G���B�絉�f������[�G��U&�����~�F��AׯK1�`c��[<��FY���4I� �#�G��x[X�=�Q1��`��R>(�w����R�O�?����7�,(�H\�#h(W�EH=�������yq��Ѿ��aF����:�U~m<|��.��0=�P/���4ǆ���T(�����wKi1�U]ETW�
�C��ΆW�� d^�;{���<S�;6ٔF[��[�ʼ�D[�������M���2^:�!'vޒԭ��B����'i�X��N�"�0�{jm2������|m�F�m�{�����3^�B������]6i���3��=i&�v?�[��S��0��M(V�f���&aBh��.��q|���WG���Lɛq�-"e�F.c�~��\���L���$���N����p�?�c%�vX�\RUT�L���L1�yU�j�t;~��f �����q�HS�P��R.��8��O����	JRv�/�G��l��{�Xf��I����nz��u�^��h#]^�B䢼כ��l���Sp�#�������	x.p[�Wً�®��e�?�f�w��kU�����S�O����
���+h�wȣ壴����Y�5�:��T�*X�C�o?�� N�#MDb�Yͷ�fA��$Mٱ��HT��YX�%"�Я������)`Y��}���s��c� �]������l�:aEd�b�q�iS���A�8������B�d�u��LK�S�Wbc:��?v�<�s�s�:ֳ[���Fgnu!
��	�*0/��o��%�CpU0�3t�{j}��l�n�Vz�7*����[;H��qkiBF�H8�6��66�S�&�����,��X8`;X
�q�h@�a=J�`���4Z�E�WE-�z`�¥߸��ĤB�?����%_5C�ܞ����
X53��U?3=gɎ<1v��Y��W>t�����H�u���%��s�Re�4:�U-�i�{{���J(_�s �Eg6��+��`]��!�P{L$�g��Fk�q�7��V~Bf|&Р��v��jʂ�-�ա��M�D4y����hj?&
-�p� ���2�ʠ2y���D��kM�1�h(�zTNl�Z�P<�SAv��%��P- ��l[{�	o�K֬ v�n��qbs�m
�%��P^o�v��,~o����C-s�˙����'vBF`�J�sU�������e�X�YV�oA�%�A��Q���
�g�hT�+�&6��+x�hP<���s"?^T��'����4��)��KW�}_�L����.l��6�YR)>������5��dQ���6_��Z��X6%i�k��ىE7�y�\p�����!xT��9�������7�krf?:�:Q&�"l�5����mm,�{
���,̹<#pί4��GO��U��'G4i�1�ɒ�]�ה�����k����m=3���	�I ����ڗ�*�f!� ;��{ɛV���֏4�Qԕ���Oϕ�{��u�Y��W�Z���|Y6��a�)�o���,ۡI$G�&y<#y�����I���9�*�Au���I�V#.
�0/Y�M@�s�.��i�Ŕ?uO��@t�k� �(+�AWě+m�>�K����n��'�bm�k$�\2wƏ��9�ݼb_v�X^&2��js����]4���I$0#��
?�Q�J�� ~�{�r��'T!�0�q�y��M�;N5\렣��� ��1
TU�ξ�; �:�䋖��t��-7G��c�z!�wG�S���P+�wl����l�����ۥ��+�H):8�*��ޔ���`F���`�SNqa9�z{�0�Ĝ2[{�ol���5��TV<��F�KV�5&&�!#�|{�[20�ցpM_�J!�����m��?a8ͥN�j� [�E�<Stv���M���J�}���7dVD�iz6�0a�Krp�sg�٫��(j�����Hk�j(��g�QU`zP�<9�5�J��M���!�UFE����}�w���]�K������x�u��\I@*��4Q�ƕ��m �۶r��������9��mC��J�ԍ���A`>$Ѹ�a���Spӭh������Xx����s"�з7	B��ơ�K��"t��\��;c�y����b���s}vD��u���߈nMŊ$�.k#�S�/8��R �V�������|'63L2�D��N��p�,�~6�Ejz���ۜ:J�fwMZ&T�b�{iگ/i�����?E���p�����
�%K\߫���Ͷ��Y��Nռq;@�SA�)t�#$S����� \��������q��*��U�
�W"�æ<���GQ����RN� 7��M��_g����<�E��",Y�+;�h.�� N*Եh�K1��(�k���� ^�LާE��x� 2s��ڧ�n$�����ʦ��=�y7#K���`[����:.����`,�!�N|9l3� Ai�rDY���X���c
��W�رOp��iV�������i92�D���p��CC��A�3�eB_1�7��*r��ܪ#�R}C��`�G!����@��a{�/�7��>����y=Xx��qJp!~�X"Ľ�z�䯡cI#� �d�*B1��zƌJ[�,M��x�����d��E��b������X�0�
�5�!Q)W3�"HDw�:E/�l[e�A�� &�������N���HlC�����dჀpp��c����_)8?�+�x=�QDQK�/� w��ip�wɬ/H�-+�:�\O�H��C.1�&��N�)T_l���J�ap4(�X�f�s$rQtB@P��m����"b:�����-q2/7��#a+T}9$O`�dCY1�B;�$2��T���&������q9oDB�N��ؚ,�WAX�'b �y�/�����	<�)�����4$�K��N�*��b0&үVT,]�g�o�W��yk.
� � �h��WK{B!sŉ�Ah�T�b�2d�2+v;R���!�'��u�9�-���c�&�n�U�.� �S��a�8A)��W ���"�<��ގ��>��rLo)��O��<Vim���'��Aɗ!xDm��c���H�T����l�XMڅ|����´���=(jx
	o C-C�3h�0K�L-�{�Ӧ�9��dK�� ��}OLy�j���%�",�@p�A�Ԧ~������q15����6W�� ۹̃M=U���C��m���0������e� �3*�pR� ���m[E��+j�3���M���5��ۅ�pA��Dۂ�s�`~_S]Zͻ9�KsN@Ҁ���8�6t8�6��-��:Z�;.i-�AEk�.Vt ~�˄��Y*1�p�����^�o���
t9�����ܙ�1�]6\��Z�W*K���q�3�3v-�-�������ӊ�T�߿,������n��A<E��K��צ���5�o���pU���A^}n�"�aM��c�S'l�׏P�ܻ�*�l��5j�vC)gA6�Y��FJ?� ��T��:Fh{����(����&B�'�f#+�����؂C(c_q��:*3�M�dmpmԐ��R��(�A���t�g��b!��`�C���I\B�?�vRYf�a�G��%t��'�BW���ɺK��Ɍ�\{{����$�Ϸ��!_���#+H\D
l�#�0˹?�;�X�|��lp���5<�{���5�,U��HVȊ�]r���0TT��x�^"�I�%�qG��lh0jޜ���evt�A!ג�m��*��+��h��0O����~Ѱ�L�	;���v�F�"G�H�6z��fc���e��'9$^1�u� sv����e�aJ����JY����FWdl�4�(��[�;������j��w>�>9�'�6��zU	Z�g������dkp���p��u�5�{=�s���2���`��tkB�&�>/��BY�&J�B���%��O _�Y0Q�R�$����_�
�	�	�����=O����Mٸ|�-9"����]����ID=o�o���t��BS��YO<��w8,)�p��y�"���LuXO�,I�Ұ<J(.2L��B�c��kG����(�mY<8�����Mn�|�:�w(��z��L���+���2R��/)���|ly���,�Y���K��N��q�$u�vXd�(=�\�9-�^6�?��E�i�:"���;
������Z~<e�F���љ!�Or&�"Q�Cih���"J�Ⱦ7�Y��`2�l���Yv�0i|"0~��;+��A}N�D��'
n�ͨ�Z�]ݼ���$mjt�	>��1-��:�*f�E��w����2�1��.8��c�W�ݽ&p��]��j4"/��z4�z
)�u�"�~�V��Aϲ��8�k�[�M��~v/쁵P ;��a"Q�����^���T��O�=W�C���$kp���v���RѶq�D���R���XJ�)/�j>W���nV5Ne�D����Ů��Y$쮅�ϙ�ښ�1k�r�K�/U�n��@�z�v�����rY�y��FO���EI��c��D(60�{J��S�`l������mq#��P�u"u4�SF�����b�{"��z�@��O����*����}�q9���O� �4�p ��*-�t���Z�6���SL�얃CaHޢ _���<a����6�/��� �E� 7Rە������i�� Ծ�2W�	Uᶃ}��*b������_�g��(�8o9+R�O�i�4jz�ty#G�S���@���6%�'�Ap`=�q�&����x��~�zEv1�O`�l��NLÕA�\��B��\����,�.Ϊ���w;�AG��F!���=-.�Vp�Kã�w�*��q�t��d�|~�狄��}���7�e�jx��F�9���i���| ��
� ���e��L�=�G����y�x���I��=47����L���I�݂�$k�O� �,��~���@	Cn.J���8*}�z`?S��]lM�.H�7K�4��~$��	��Rt��y�*��rJ�{-Z߆p�){�FZ3ʓX9B �E��]��_q�����!�[��4*�y��&�����5�Q�pnQ+ǜ�6U*����DtpH �'�M`w��S��L�R����N%�Q��0j�{��Nh�De�h��d�����6蔥L��Q���{L蝆��VPx&�K�k(<�zo���-k� `L�޻�$U�z�k�MH�]֛�w�枣5s��Ϝ�N�+2�p�M���Oբ%��ذ��*�u�q�e��ڴ�ƭ�aDjO��*���+Sqh�&ȳ�-��̒ ���M��Y��$z+qu��f�l�		;��N�)=Y�
؟��`d�?߹w�r��x�&�`�SR�:^.2��\��6<)���ቄV��$����g�W7���DCIm���7c�+�^��*��N\�ء 5NԚN���QT1I[��S(%9��T��+��bSX=��n)}'���y�@�S���K�KB.tw�&'�(a�R�%@�ي�e������T���)w��3l�+�g&�'�ٻX͕�
1��;q�kĜV�Srh�<��F�"��'E�z�%X���8�E#˦��������� ���	V1�H�P8&�uV2��+W_[Jg�6�A��O���Zf��4ڱf��"U��,'�>��W�����uc���J�_D���w���7L�S�Z{�E@`����Ӕ�Iؽ�`j��-Q�ƍ�\�^���VE��X�>��Vy,��Oؔ�i��Ugj����ɯ�wd�%s�X��\˻�T�G�ӛ����΁1�rOqi�{���Ģ��U�����Kz2*����'EǈsR1�D��p��|�v��\2�&i���,�rܞ��P�gC�-y!1��c+q����Fw��i������T��im�K� o�ݥ��8x?D{�a��4X��~!�DEg[�@8!�=Ƹ��&�c���i�`�(N4�t�����V��8�k[��Z��D��n�;F�hAڦc�W�� G�(�lE�:�z(�R9�"�.��*��'��0���X�|��&p������])���߯�:T�,��q�%y��-�����6�����&=�����{]Q$��O�P�Ϯ��"@w���5�_���⺑��j��T]!�*"��w2�m����Y�e����v)��&輳+�"9�&�:M}�F�D������<�ْ���Q�;��� �t�ǵP���.]Q��.6�GL���W�W-�tp� Ӧ�"}5~����>әy��_�ewO��U�
a5���f�K�s�`4��L��n�0�o���=p.�*�	�KI�n�~�pF�V���lIµ���;ڹ7t�#`��h"�t�DߚH���A��0	̧��?b��L��P��~����l�&0ñ}�-W�����S>�����ʠُYk��u��02��Hō�~Q1�x��+���Bj��O!��'M&tѳ�[bk_"b���1o��ӵ������V��@��I4������^3���"欕�>}D���Wj��Ic'H��q���sƩ�%)�5N��+���^��|г����K��uo�W�#�,�����*�%"� �d�^�ԈB��_rcS�!o��59J�_�e�+e�2��׿X�q��VF�2�XX!l��=_��宰��.�F��<�O���.�۷\ A�	D,xG>f;(lz:K��`/���!��9QV�"�����`u�aJc���^�w����Ch��F_�j��L4�t�N�U@�Ʊ>��>��פS=���<�6�wһ�'��އ�UzK��c�y���n,��u4H�is�܏���Dm��0g=L[�{-�+��|�zCl��������a�g��0�1%�ң�H|�0q?'d��24Jz�Ɛz%ˀP�X-��Z'i��/���)5�7n��ɸ�|U����M�Һ� �t<L� �;�`x�����N��Q����9./�Q��Z�J��q�:�n�xg�
�-��hPB�<z��Q�;n�k{a���X�Ch�b��]��`"�3'jy+"�ȫ!*�:�#)E�<g�k�D)b�-y巴��+�ڲR�댼�2��8.���(K�J��-�����FZ7��v�I`o�Ѥ�P�m'G��[!X��X��Z�eY��T�����T��X]֦mZ?K�Zf�jW�sS���KK�(3e/��G�儋ה*�L5 ª��ù���80-�Ջ�ᢜj/��Ӫ�,�֝py�x���%U�e~�E1~q�����W㼤}ş|��'�|������H�L3[���:<�&�l�&��qt7FeLcqz�s��k��4eo0'g�#�{ج���1�s���xvm�nOR�:�4����%�G���SM%쨄|��
��SӛL1 f�X���ɧe��	g]PZ�ď] �q*s�,`"��ؤc�G����L��2h�	��A�ϒ,�c�B�}���N���{q�?c�<"�ݬ&���̮l��CA�E*��b æcZ��|��n���~��/�v-��ѓ�d��$SJ�u쇼��_&�Ǳ>y��� �FȷWT�!���r6Hyh�Ɠ�����3` ��&6L1`��Y~a]�l'YJc��Bȭh;���_�PЏ���tt����
�M3�Z�,`�!�U9j?0�y:';b/- 'а��V:��"��d�0���o�.	0P����=W��b�N��2�;�hA;m�tcT��a��oo����Kp��ȩ��Er������v���u���c��.���w �z<��Xg?-_�8�Y%	��/B��92ƺqz�|�Q�����,h[~���	��0|���@ G$��y��U���q��3u�*)��t�]�n�BTv���G��	[垮h�N۶�����"�=�~��ő�qV�p�Ɓ��r��P7+�N�օ�z���t�]T�:�S�r��QP]�s�xc����RО`�a=�O>�h�J�n]�;n��m߶�H��<�`X`Ɉ���5���N-���92̩v����?����P�˞�Z��@@߂�{9R�a���QQ����~�rָ�CG�����T��'�z�� 6�ޞB�CO ���7ٔ	���X�a���޾����62�Y��P�g����^�ZE�����C�ӊV�<*�{�@t%�iС.�HV�E��h����g���r�א�{�f@��qRG����Q�N������4��w��^B�"���,�9H���!�#��S�����^<��~����WeC�d���Dd0Adh��w�̓k�+�������=]�3�u�\1D�
�%O�6?�/�lV 5�8f⩰��P����Q�E�7r`a��䵋�cY���|<���-(&��K�E�P��z���vX�Xtn�6�>A5��0��O|�u���a��Eo�DEkmMmƪ����09<��G����Eݖ�h�b{��vM�0���LƠ��U]�z���6ѫ���#t�p��Ĺ(�W7�z�/�nR��z@@�Q�%��B�5��|~�E�|ˬ�����O��B��|�����q�ݞğ����Y����J�+(p��C����@iӃ��l,�/��Ñ�M(��� �[Y�Y[�3Z{8"��J��)H=�"#�Z�W+
�γ�!w�]�D-���۔�1�P�Ts���ߎ�J���m�1��r�DJ�{��-��O�:f��͊?Y`9�N�{��꿮~_��L=��+S�_�2&��+��@�vh�9N ��Mc�>�-��$Lt�fW�B1+��zt��V�8�/S��v�5w^����X��N\0�[�\��M1*�8��r�a��Z��_r�gsp��R�|72>1��_V�éa�+|4�q��8[	�����W�4�{K�GщFq���	6��m`�v��{U�O�G'��z��F2�H�h�0�xԼ��0]d�z3Y90잆7	w���^�\���&!���;u������<G9�熎]̆�,RY�o��F矡#�tWD�7N<'�'/݂�"���{���� "�
������H��\�	�(Ғ	!�5Oی�8�M6��)���\�o��eA��!�W��ᓼLT̴�"��{*��$4:����#5_uU�c��!�2%�� &T
=�Ѣ�|�ea�a���~�a�$��d�x*ǿ?�R،��Q�VI���B��[��<���Rmsg��v/Y�[�q/����L[��V��抮0HGN�� �k��n�k`�������c�бo� ��0�a7~Xz97V�{�V��_^"dAR\��*���@�����/Ғ�J��E)�#2EwHCf�n)��OCu���E��]�z�-�F���c��F6YvYE��q�%�bn�����|���������o=��+����8�o��[>.@Ӛ��(���h̢%�e�@v��!LO?審���<J<au5�W��	^T��c���Vv2��3����.t�]��V�<�4r)n��բp=��w;���8��"���̘�ճ����O
0�� ��]�]a�`�gj�p��JWS���1�50�_���*	�艅{���eD��7Nf�^�^7���?�SG�|�yʡ�g�Qz�	�Ӫ��~fP],��j��4�+Â���í����o]W$k�1��<]dLɦ6&J,~�O8ʋU����+��U��[��礬tÅ��?J�t��3���%ֈ�fۂ[C@#V
p�Y�������x.��P�(ݲ1���m���ٍ��s���5�k`z�)�� &�~� 4��r��2$��{�I�%Í������~�1�!��I6��(Ay� &�`�ْܲ��������TǼ�I��z%G� ����}��z�?@��,��9T�<�U�J��s���
���0�JN1����޺��.�B��	���q�	��G�8�7�V��&B�oh�A�YiW�:-�y��Y�I�\��;f�(�/�]���Ԣ͂�M�֫\j�8�vʍ�!�=�BU��A�O����<X��s�����#�`K��޸z&�x��-�Ý�2��O?��>O� laz�wteH�(������FQ��]X�މ �%#B�\�H�h�0�*�q���9�>Mvs~�������t���}�?���#�
�M~	���@ �Kیd������-	Qq�&Z��ޡ4���DF��MmE����R�����cc$�Ѹ嘩���}lT�����'����@��/L��!s����>1˳5]*:p3ӆ�l�����#��i�GLv� V\;��Ϯ�*�_�9Ӹ_~��آ%X�O@N�¨�H����s�ݛ���+�ĺ�<�p�����`��(��ީ�,�Vg�W1
_������l��;y���WD���w�mCA����;>�s3�j).���h�y3J�>���
�y��ݥB��;�4�8��D��ш�I�QF�a���_r�_h��-N��u�Mv(b�C��'���v�z	߷��y��vT��� Mf�V��y
�#����U�9Bǀ�2��Jc#�"Z$<e���%ˢ�ʺK+D�2Z(����m���>�� ���y�i�\'�tYPk��Kq؊����{=�?�F9HP6%��ʠ)y/懷�Az0W���ɨ�ܦ���brGǇ���`��;���<��3;G�Yǌ���O H	a���������&���
~�1�4��|Z9	���1T�A�e�`���c�˝��Z1t�{A`�1q,�m'N	�|����#����<��~i4.�f���B	T�{�6�Y���Aޡt�[03_���bEB�P�Q }���
�w(�]a�$~�m)ɡ��H�CDW_EJ[B׳�T|5D�K#&�<�8��
�!`�{�(�:f@.�JU��QLu�V��,WOr,�j�У�-���׆C��u���oHϜ�N��0��nP�����K�0[�X����+U	�&�3�/��63��i�4$N�XV~�q2�Ψ������c2c�S{���~vG�Z�6�a�x�å�g��B�����b����G�_����6E�B�G`2�\9� �	׻�TR(_\��5���!�G�����	Gq^dU� c�A��|'��jj����@�={�W�,;��� �� 2^��E=�W��x��9�J�MVƢmsh+^�۫)Z><
�B����G�Η>��i�nK�j��[+�q�*�/n��%��#s��K�{�即�(��_Tp!�=���<�u��P˱�����g�12�?�V*���x&#�}ZoHt�H�h#>��Z ��K{ȼ ���gyh�Z�Z�G7]-o�X7���Q��N��ug��r�k4�݋S;�T'��m7��:,
�m������bx��/C@q�t���+���k# ��o��[f7�G����q�=���uND�z:�Oo���FeI�k�4=,��%�QBp[x��� ��1�%]oo�"���ޙ����3a�Ƹ`����{�$��[!!�����c�5��M�#`�@-���Dz���ƵJ�p�̀�~�N���?��e!n�`��!xE���術M #o.֓�D��J��e�Ņ<GO��{	.�?������<53;�;�6j��T����X>��h���FJ�S�;۝tH�A�F��5�����T j�A���|*�w����d�ǎ��޺׻��{,�a@^.��6���?=�u�AA�qz��!s8���*`�D���A���͊�v�?w�"S	g�D^�a=�~�A�tm������x�Aъ4���j�lhr�
�ڿ@�o�"nНs˩Wy%�&�]�A����k*�F�B�|�ч'n&���\֠ `UTW�i��;o�P����"���������P�$,��{|53���(c(6�g`���v�/Ly:X�6��9a���5���.埊��T���Y?#��I���A�
3˳lШZ�h�����
:-[Us�-�{��Z��D�ǵ����&�G�sN�N�P�vZ$�5�t� �bd1B��Q^7\�Gd�$$*�f�A�z�G�~�#b9]��� �ᝳY+-jG�&�ں����?�;�2$'^��f{�e�!8v�T��ˡ��w3`�c�v.ň7�G`��.��o�x�S<L�ғ���{7���A[����Ya��?w����s.� ���m%eԿH�
u�	��<P��t�l>��j����Y����w0w�J�	zu[�{3�+Nl��0���u7P]�'r�G}��c�O|�o����m�J��ũ�|��Ѕ3+?�{�n�*����P�ռ�09:�`B���9Tp���~4@�ogN�J|h���/����_�σ����-�ҕ�`���Q[��Wxm)���/"���%��4o�7�y�v΢7�������2�8�sӦ��{j��Pز[R�޻�U�^l��H,K�5p;�7���6*{�b�(�̕���;&����C�HT��4.O��;�e���]�j�3��lB�k�3(Oj��VM��e��]y~�iA�ԋ��M-��2H���\;�'9�!9f[r�i�pO�$�d{G���*�W�]L��rJn^kҎx��})BL��V8�J��,�cŰ!���jj��i�;3[mK����!
;=h:jT�*<6{��4�o�h��铄��g�����^ #U�E��M�2��$
�`F��ԧV����D���^����`�ol�@�=3\�[�N2Q	�[0v�Q(���KV�&�
)̍�N�/��%��q� �\�b:��,`LPd�`"��t���A���f�z��o�s��A'!����Лz��J�N�<�p=m�%̛,c91�X�j�;>�3�>��˔���وc�֫�;���N'Gc���a�-@O�^���a�4Ӿ�<M4�A�����6/�jg�:����ˤC�%������K �N}��� 9Ϝ���٧��Ȅ���ӷ�^����~�h�QsJ�+l|���T��	׎�*�mZ�.�������P��_�%иk�A���x{)	�,U	�aN��r���U�^{M��e�W�#�p�cq����Ft6����X���AfD7GX���A�����u=�~��abi'Z~8���^[m]��~�V7�QQ-�'�t~� )^�-��P�x(�C	�&��ƥY��#tt�j�z��F�q�ӦM�ҁe���yVPj͇~�}Hm̀�|�� T)���T���G�7[���mg�swTԶ2�%+K�M0I��/�j�2��as�4��D>�®@(&uk��N�l�p��������fv��B�I�}�-������5�x�6��W���c~B����e��M�N���ߏ�H�z/�)����{r&e��j�xTe��M,$TY�g���P�Z�V��2�������'�_�����>v��Z�n��=�¬���LL�	�k�|�,�2�nV>擾�W�ct����< n���j|�ߔ@_�2���ɹ����p�3�f�*�N�߂��Ǫd/\��'��qEF����o'��9��r9����E���Av3(���ͬZ�Ş�=��s�� Z�T�;��-h[���X�(�+��K1y�2f�t��z=.�F�#v-�����MO.<��>��ȋ[��!/�v�",����K��'���|����������[��-��B�'��?<S�s�X[���S�˙�/��Ëw���=���L��nRZ�ٲ˫�Y}dթ/PI��'��l���C��́,ZN�-ظ_�g���QU�ڰ֠��?Ok��c6H�;���d#yBG��vp��6X�,a����,��*�Q����I�;m��f�rPttK�H��PC�x���x���������֓�Gf�Z���;S @}S��`sGS���#h&���$���W
�:c��Ĝwg�ş/�:uJ����I����➠�m�]RL&ݷG¸}�V13�>U�`�_z�A��ܸ��;NT�S�*��$t��hG	<1��Xb�@t��^��5������D�֗;�2� >��UHI{`ד_ع�D��K���"��Ĕ�RX����l�li�-��n��b�t\������v_0���g�*�V��V6�_��(2#�BS���oƥ�h}
)�>�j��I�#��ʘ�2�f��� �1�w=������?��6�ǉ���y����KE�X�T�N�żd�WNoh��}�1� � ^{ήI�K�S��RAr��l�3
�R�
�ʟ j4Dk�שEW������5e�����-adz�����û;�̲��de��r�|E�N|E<@�Ą�P�j�S=��}׏����9!��Q���{��s�(����qI8�br���ľ����0� U�"_`���ؕ�ޒۗ��K�j$��OC�>&�(#�Ū��0�o/�*��%�ot��T�[����͢�[4�`�vel�x̂����w���Bݜ��r�I�&2؁8|�aW�,)"�mI��w��&K6�$c~6C���8��Xeu�5u�K6<3�j�6�X�7� \�!�|����HŎ�4�dY����_.��̸�����	*[��/��Ð���5Ϣ���B-�`����7	B<�8�� ��>:�9��`�֣bP+bp$�f����cm��sK!/�*��U�"�]su��)��}�s���7�"V�N��b�f��!��+�{�`W��-����� �1LX��I҃�n����9L�mt߅�`�Ee��]��!=#�>�H7e�����n�mi8��|XG��"�B]bP��d2y�ε����l<�u_`��8E�	�v(jC����t1:��V���%D�raU���G�v<|�ߜ6�n�t��	K_�����
Չsk�q7ImPu.�P]Ϗ��X3�a��R�P��e�h��S}0}�!-�1H\�������,�D�i�
�����(J�n �I�/P��a��G���O��6͠^kO[����'[���v!�1��~�Qꅺ����4)��9 �)���e��e@1�X����\�����2�3.;{瓯��\cH����Y��F�K���Њ��j�N9KKZ?꾻kl/ V��a�����ύ��K�;%gY�߷�g���#K��V��.*���ƥ�I�g������8�8=!p-	Du)mvi	���l-�aX�AL��nd����·��q�<"��Ĉ��aW�8�q��(��m�2MJ_w� �	�B�l��l�B�b���Ҵ�e�a�X����y�r.�(պ�%�z�oP{H@��OrQ���E�8�f��$ۗ걸�ۛ�	���L���`�ENC���'P:����G	@���D�c^��\x�a��ı�(�	B�-Vt-�oq����1Y����p���l?���>�D�VQU��M[*�[�u%���W4���c"\�prDn��[�8ĝ�m�+�Mh�����ǯ��PW��c{-����L�K�arX�^�k�|��7U-m��3�W�������t^/�B-�Q4����gWi		�,(�r��&��$Lfݺ܎B�0��rP��`�v�&Ou�xҬ$(%	WЪ5Y\��O�Ø�nR�wʍ��U�V�e1�+g|�d��׫Z��5_��!�Wꚅ�7Tv�T���+��A.4b�ve-�<���T3l{_�lw�_a������ v�^ ���Ԩ���C-PV*���Ƃ��J������-1�,���LW>Y�y0����4+�ﴌK��$��tؼ��t���IF	�*�)�N���g�Q��n�.qԈE�x�-Br�wG�!1�䢶W!g�O�)��_~�EY��6	�6��_�g��H��b3�:>Go�M�� mwƉ#z�2�p�U��]�.����l�n.Tl��ƜmT�,�Gܲ�4rH���HU�C����a������k���3^��Y&/M�	�(G���2e���1�(�����j�iH|�����e	������*I��
g'���5 
���|~��?�{�y�5���~4B ���@�\�TB��(���)F'8�	�n����i���z������T���0hq��Q`�L7E�����g<��o��N�-R�����Tӄ�^��}Y�����&!}q"�����$�I$V�z�r0/Mv@��O��Po�C�u��
����z��~ʷ-G��3�۫�&��[�};�Zs2m�=��H����PJ��{B���=�j�@�"�Z��t ���:7Y��n���5�F�U�쳘0E+��FL-�Gӯ�m�p�ά��Lim�����4�Q�{�F(�G �%��h������@��Z��)1-s��Q�vF�+����|i�3�u(a����M#	]���K��V�&r��~�Y�KE{�ab)�f�H���
���ܕ-�a�}���ʞ,Y��T��Z�Ni��E%{uA��(��1#��A#��l3ﱙT{�uÃo�6���XQ<x'��� k�g�(��H:
n�6�k�������a9�d{al��d����y��'��ލkb�8.��s%I�s����~g<�:�|��`���[��GH�>�Z��f/�t�H�p��E� �I*�\����\[x�9�R�%X�H��Xzi��V�IрE��Zۣ=�[�Z'I>jD�ϨZ��!�Ŵ�k�U�N�)eL���� ���/,im-t�0���D����~D�~��|��(F�1%U�]wf�Ӫ^`p���~�H��lZ�>^v4R:�Q�y��� �������.�W�(�:���:�񻻢ᴠ�����\C3m=9�ᣧ�^H��w7h9��A�����n��=�l�&�<��&�OAC����.�WJ��Af��e��J΀�k��3����@_�Q����.�66:[�K΢��������-�'�'�E��w���gޱd�h�Av^�q�$�>�ȴ7'����c���@��+�JD�b�u�r��bX���`'������,�!lKWb�0�c�^�A��JW�a����~���LU�A�T�4��〫���w�Q��Xr��,	����W�~?�ނ�j��'�J^?]��r�親B�\+��T�~���Z��v~�A��s�����/FWx�$讆�QCT&k�s�Et/O��� �T,6��ɽusP��,��.\��l����	9[u!�e��K�N�wz���	����MZ�?(���nt.��I˝k�v6��CV�c�<|��0s)�z|���QDO9�1��;5��{Z�b�{�h��V�9��8��G]����0�UAl��VW`��x�:=5L�Ĉ �7��ۋ�	��(Ū��Ո,�?R���.��q[g�͓wh����0<>8(�[-J
��nU��{Y��<e5p�Y.�(��П�'&зr$��^�4l}�$%f�V*�oKɶ��!J�⠉�PC��*�{�C�^s��:�x�w#��DE63l�g��tMe��� ���a���cX)E8��`o�l��g}/K�F/7�"+E'!<�Z�%�k�W����p��3\G(� ��_0��]�0b��� g{}�pxǻ�ե��ᦃ�("_,B%��箁)��ycMИ�i<�}ߥb�ޚU��S��b�)��N���z�ӵ΄������Ik\!�V���@؅�B�̷>��̽-Py�i)d�Xqfʗ /���"�=����۲��Ӻ P_3%R��<y�A�w9�:�~5�"Q��Q{����Y�Q3���K������W�\f�k�WaXǣc^�c�ϘFG	L��P�e��~�g���(V;ɥ�O�Ph�u6(���;�|��U�L+��BX�&����<�:�X���6I@7�\=�]r��
���WI������b����3�$(��5$/Z$���xLtv5�B�b9�;�)u���{s;���1��l�tZ*Ԝ^9���f��/|��"i0�t"�
�s�?�o�}���b����*��K ��Lk�s�F>��z�y?dj��	�HFh�o�"]5��oY�� &���'ci�OI�4�p_��ң���ߴ:vf/2=Y��q�߁�����`&����K��������r�KᏁ���^@R��#W^�dYꘞ8l��G��8e�
��7�Us����7;����ȏ3�$�+])M=\���5�%%ؤ������;M/���*�ܱiaw�`{1h,��
�d�������i�\d�T�����br��a�?��{��qgyz'�|ME��&ftg|���2���$�v�k��:<�!h���੦�ȟ���Ĝ���f�@�!��Q�h_���|a�F�����OT��0.��z���m���4A��BR���z����pT|�K�.�̘�M���{<7����J	��Ќ#�v�m�Ap�	��XGDL�!�bIA����f�Ɠ����P99oX�V $c�Y�B^+?�.�19�r��w�Ѡ�)�ꙧ��Eb��yU������Ӯ�����i���C^��ɸ4�eόH�-=zi#�E����c��QMgҜe�=>M�z��2�?����t�;IT)= 4~�>�}ژCǃ6��BuG����Ǹ������h+Н��tİ8��s����R;�~��S}m�?�綡'��)m8I�.�dŠl幘�3㩚�iH�����^`[�Ŧ�4(z���Qd�=�e٪��"���D���O	��E��{xܗ�J#����� r+�{����~�W\1��Ī~�z��=����.&B��s��*�6X�����G�:�B;F�:�f�J�E{�C\�����{A���;����w��S��)��M7Dh�>۟}G
�L�R�K}��?��,͊�n�=�">w�-���zp1y>��Gk��qEò���ӽ�ҏ݀x������0;!Mn� /f���i��P�>���s�!�8�R�H�(n���}ć �x.BU��#�un0��:��Q'D�E;L�����W�i����fR���'ˬTG\��<1«f����j�+4Pʯ!=�A�t��/q�������zѪ��fU�<�тi����N����z@��m�����ǖ���}�p����A�R����V��
����3|RPLT�p���]�hcbZؓ~��k��Q��p���w �S�����k���&Ｖΰ09���
�IQB�����x\�wڪ���6�2pS� �o�s�֭��B�) �ax�j@�W���fqχ+�`�{� �l����\�2�zT�q%ŋ���պz��3�'�$�BS8�^Rٱ��P�X�p_N���4�M��|��a9���%���z�E�M�KHX2/��E�{������.֟D��ƍ&	FB�Q�����H�]�	$J���� `���j�X����$�l���?�hө�#q#7X:*��'��������{<���_PB���8�F �%s�{=��;���WD`k(�x�V��\�7���Ud�ƗM��;����NM�ҟ�/���B��F`N9��A����� �-k1�I3 �[OHbˌ�()a�(��\����Iv�k��Y�1���$��!&G��£݂q��ˈ/J�O�y`����K.��f�F����*�&��썽��"u��Pajr�1 ̆ڪ�^v���o��t~��t��7� Hϳ�)��כ�뺌-���[�ST�"Q)�T�/�fI�*�/P
�3'����k.���Dx�~BB�[S.tʅYD���*}��2��0�̗�R�nzE����mj�R��Ļ�K���8&���#$L�WF�pg륩��S�)�fú�xg��\Ң~���RZ2G�h�6qkg]��$e�M;/6K��bf0l�TnX�VM+ ��S����ܭ����Ƿ�� �J�:��>���m	.�v�GV����)rҿ�'�!����x&`t��(Gn�q>�񒞶V�#|�4�,���D~v'~��-L�υDY���\�ۛQ>��ar���J�u�����{{<9�����L< r]�$ճ]J�⊴��5u���C{=4J�����'%@�b�]r�Qqr"D�D��`��녻꿲*5Y�*��t��\�˟Kc���-����b{W�8#*��γ8���>I�LB^O�B���F�$�Ԭ��ȓj����=a�A�{ƷdTy�L릝$�M�YZͧ��\��ehU��.�_`��Ӯ? ��f����.h5�μ�����Bj��B c�j�V�pC$��`���n���W��,��8$�uf���Td���_�\�q~�A��J]�ű�=tQA4g��T�'Qkxnp�8~g4	c�W�G^<�	n@����'��.��I2�jl)V�z�ER!c\oĠ�;�t��6��!�;�?<l }j������&�!U��w7�҆����M���S5�駿Rq��ժƪ�-���?}8	DH�ˍe�f�VXӳ[����@_�����-��a��*��e@mG�;��W,kR�{�e{��+�*��:]��g����R���W2Cnf�$��lv�R�	8�Qaf|�'�%�61e5�n �OP��æ�G$XG%\�C�� :ţHXy�_�;���6��Չ���d��Qi�L^��V��&���>͍N�m"�x�y(�m���D/f'ׁ@�4�3/<��!ʗ|C�kP��2��c�|� �h��{�������bU��y��#
��VO��2����^3%O��(3^{N�Bm�L��)�@�4�ՃA;�6����{!�|����@\����K磪b�°�ϸ).�hJmN#_s��j���Ϧ:��.����
�t=�@�Z��l݄5�&؍�U��6�.g���I:aĨq(��Cv��XVR�5��I�'��e}�sM�P������"pr�a�^�W�=���z*�u�L<��7Pf�t�dAI�S9���3���l��Kٴ����֎�O�Nq�#��JB��Y������.�v���;s�}�!��1P��{a��f�t�}]
���C���{���N��%��@��G�uF T	k46i-�[�q��ZK�54J�����Og�G�vI��]�����a��0߂�l$]|n�\����(R���a��#�Jߪ�u(U���A#A^�o(e����\�c�jV{�#��ԏtV��q��>���Đ�D@���[�{����}"�T ���"�/�{��:�W�Ýl����[z�g)��n�])v�
;�֤�����߱<dD�V=���<��%��WĠ��E}���C3���E~��%C��uo�Z���k�9GT����V���5����F�!ui����9�L˲�ik�3�L�:����8-�:�%@���+���7������~ǧc/mV�Ƙ)(����(-°��QG���� ��5�kCt�?�Z�|~K"
������w<E��9Ӄ��wCn���#x����mTO�]d�m�����闁A{���)9&�o.�Ԟk8.�o)���@. �Ξ�4�O8�*?"B���8���(��z�-N}?�Ox3ǂ9�%��߮��x��,c~Y��+8Oi�1~�� M*�f�V45�J�W_��V�� ��g�`���ҽ�$�p�b�!���0���ӖD��=���({m���ct��^�>����f��1�J%�|�C�i��i�g���$��V�363���RC1E��FDRfi����3���$��_�p�E��1?��7�?���V[���+�����������H����D�k举O[;�_�"�5f_�/�Ф>���h��zT�Z�xe̔�S.$��nRYjU9
 bY��rZ#�EL�hn�2�s�ɸ�V߈�8φP�(���T��WOVc>*`.ܮ����a^N<ᔀě���u�nU��H�'�rc*�V:_)`����t=GG5�Z�W�$��Fߵ��rw�^��C���w�4����+�{��5>҂�n{����;O�9�\��͒D�TH��ڇ�b��A��*���T��Y�
t6�.>,�N���%Q���d����A�o���r��H�� �<��GK�E����wı�:�>�y�h��w��P� �(��T!��#����Tyߞ�(Sm'�P���f!�_�~�u�cѧ� O�@�}��i%[�IaLS���6�W.�$2��5Q� 5W�4�J;r	������(����7�L��g��J���e>��v��Kx��	ަ���0���F\�~Dӑ�@��(����cͮ�2�^Zf+�{���=��3s] _����� �ź�Y�$ �I��bSɻa�dD���V�鈢��W%�FT��u����|NDX�}8����88���8m$u�);�����c(�qD�U���ub;5���ȝ�XOӮX����M�WƜ'�rD$�D����X[�>y0A	��Y��'\l�>E��+��t���|��3��;qg=�9�Lm��i>�0�� ��<��Ѱrr��W?�H�?3c�g{0����V��ڲ:v�p�k�U�I>� xmX�w����0�Q"��sz�z�Y��m�+,Y��A��� :���]�>�z�7�g���],1U��gJ6:�♆\�t'�6��Ǭ�yh9�$��w��O�Ӿ�V��5�t;��Uː�������崯��(=01��
���������7�_�D�q��V,�*.�v�2��M���vR��DI"�����)��C0�nā����i|�D�2�1pee?�z�+���*G����mO���%�T�c��OC�&�<}U�(oB�{�=�/h2 ��߇CD���O�� Ű�ܤW^��2�-����,,S<���w�Ԓ���+q5��Q~P�� ��e�g�N��/\���l��e�2M�L&7�sF���b�����q?�) `���
3��5��g����5� b����Sթ�\ ¼߄Qf3+*6�1b�0&ٸ�����8�M%ɊLl�z.��(h$g��+N'�����a��hV�����&p%f�/ �6O0Te�O''N6�	�:D�ky�gr�t��eoE^�E&�ЧgBF��@�#���Z� !�'B��G<!�E�*�-���� :�oRhӈ��[�`�:���Ν��1鄬&"�?�b�^an`���Q�[kAh��^�^P0
���3}�f��n�Yׯ�K�Q�]�����X��=��X�)������m7G�I���e���J��ÿ�av��/R�,]�K�o����@ZQA�,�.D���e�*���,�E�k���d���NB������7,��ix��L������ㄋ� Eև�zt�,�����ز7���οS8�5˗1vj ���2�u��о�� &4�A��tz�0&y<\�x-1=A��`�h��On#��M�&L5L��~���]�����������.�k���U��1q�>����־�Y���4�.b�������o��Ze���L�\HQ��W.r���=�T����z4ZHWi9Ǒ�y���]��h��R�u�o���3�b�s��{J��h���i岍��FX�B���}'I;����ϫ?�F���; �-4$ŧ^rO�PQ��zb_h64��2Jc�(���Ԛ���/�j
�61�KT@�Y �jJ�����V�r
f�;J0��.�ùG����i'D�삀m�'t�9�.�YV����t&K����w_�i����AM�4�F��
�T�D�5�}����V7BC��ժ����0����?;V.�M�n'���!�O8.{����J��۴��k�v�47���k�^ƕI�=w�i"�W�rk�-ma�"�l�KX�P�������/ 
1�>U�AVya���*�GȆ�0�W����6sҡE
ֲS
[�����3�;�}`ܢ���s�>Z��V@Y�>�pC��&@B�H��� �)H��=t*O�T&���M!A5y�M�-��d�tqtz��S���<�u-��R:�K�lC@���Z����(ĩC��9���W���/1z�n�W�ZZ��b���;'��#-pä�"�қ6�+�܆��0Pd �FJ1��*b.J5ɭ"��j�uk�މ�fı1�(�F��8���R�#T	�r�����&:-��ᾗY\�`ЏAsX����z\�`��.E�N�%H �(�"3	�)"?�I	�Z^n0��9juX�����[�%�rp
�^!�t�X6���XS�Y����t������l^�@rG���`���y�20�������N����b�9sE���x*�`p����^����<� �@�.e�@�'��<J�s.��:��}��]�uD�W�K%�-<�����ِ�_]�KJo�b�a5�eϚ�Tn_��-��^�د��y�����m��\�zu��7�7mCx㵴�jRG0�fY@L�`F�w����Rɀ����{;5�[xz*�=���Yx��*@�*k��x6���|g�`���Ѥ������|D@.�n3�V4)�'^�3��{]�q�'��ԛW�����6��7*[ĵ�_e��澁k��2b�U����o-��e��TzqY�9cX]n�H�b#� �nA��w��!l�0D��^�ٵ����3�xN�T���r
��01�B(�s�G�T��b ��P%�T��;,�*�`������|�v�)�U?t��Oג�!V�nU��N�h0�?���� S�LE��u�J�K�~è��.�)����1�m�zM�NPg��H.U;7
�Lo�s=lB���*�//�8��Fjgl�[����ZKm���=K��r�A~����;x��O�xZ�>H�ჲ��`Ao������9���Ϳ��x���;��߮h�u��6�M�J�X�������I.3����hēr=��\1}�g ���[{wJ"t�=��������������?9��B�؛v�}o��U�.�R�*��f�g`��6J�}���T��Q�tlo�k� h8�������h\o2�m�~"���.t��hΨ����!������Pɗ� 0*8ǲVJa�n�؁
��z=a���
�|��;$�VcglL�<��f�A��B�-�JY��*]��B��hN�bD��xuY ���I+B,4')-�aBx�S�X���ӷ�iCpl/@L@����G\ww)�-�_�k��� a��UY��zWq�/ "���i��%vF��j���~�e}u�ֲI0d/�paJ�^��h]�)T�`�ZK�,W�,A_�k�Bi��-l�0C9�1��F O&X��2U.3EW�0'C3��H�x��Z ?��;Y�'m�.ڢ-y��Bon�?�[�Tێ]҃*I@n;#�KA�櫏Vu�S{���I�q�n[<��pX��(��"�k�Ǘ8KQt�������Ñ�_��v��|��W��D�c����&D��R�����藶=]�fК�Ɉ�� �����D6W�� Ԥ�0�%6�f]�|�M���aY�E�����u򲴁P'~��. ��1�o^�M��n�p~����05Q'�$ש0��|� I6M�<���^YxIt�$
urV:�����J��RlW`�Ӗ� \�
� ��\��+.A7�j�� �n���b��
�U��ߕ�#��|�2R��Ꭵ؅��Z�xp9�F�dpx��sY������2h.�`������D����9y�է,���()R2v�\N�y����<�j�w�C]�"=�4x$��9����"LL;
��Xk�B���D9���`����?�D���D�����	���5���<����D\-�G㈹����ϲ�J��Q���]h�L�`���>&#�8�"��;T�:�E|�sؿA�e�zG�TPD���zP'79�N��Guu~ko�fk$�d���YzKm7Φ�f0��Y�Z����0�QQ���'��"�wۍ���dg�K�%qGl���\UarW�X���4�R�/4y]2g�/Zo��ΐf�t�Er�IB��"�Pq�;@�5��>�"Ts�mE׊�;���E;(QG ����1��3w|\�,w�M	��0����T4�a���e�]�a�Q+_��$�Po�������r5��C:i�=��#I����[P�EH3b�a�����G�C>��M�ٜy�V��o��a��^�Y�e�*W�\��ck$�w��y*~��|�	�*>c�6��:&���3?+B�$x�BHy����r$�N��"(�2!!{W{7�n�b�i[�t�C�(6�LzrB���
�� ��-�_���m��Rh��4l/g��_��ӽ�N*©i�5�(�y�c��Ji�w������z)��T�h�t�U7i��1 ����и�������uP!�ݐ�f,bR �k߰���E���T�a�"�Po����Ch�,���S�?�b��,<X��D�aP䤩��/*�\���6X�"��.�B���ǡ7ݸ1
�&o)�<�4g�3���[��6���ޮ�&�)�F�v�3NP���q(����r-�<��M�@����[U�S,t� �����ߨ�8�Ox-9djq-P�z���د(1E}�G���r�-g�t��H�v�O�E<��ɑ�d\v��*�"Q��-'D�h�@"�n�'�~�5��ʶ,^l���}m��Y]jŗ�|�U^�}�W�6��)�$ƩE�J��ҙ�� a-��	����� �D�W��8Л�՟y�u�?����(�m�i�����-�.1^�(���?����R=[��z�T=�'���$if�-�gٹN�:�A:� �pr�o�zn�YIg��E����~��!�V�d�p\�o!�Z�ɓ��Rh��J��"2��LO�mV_~O0׌~��-j�Ǒ�m�żD�E����jV�Ƚé;�����)��/���e� .�я"�aGY�-��+v%�nDOv��IS�d��L�q��ڰ��}}#�����"P��~��.;@�*n���I��E9g�����:���C�
��k?�4��Z�+���.ĳY"��KCf�B����9MH���u�H(�c�(@~0,|)"��g䉶�&�0��tť3�ȈI�TM�*]%�K��'	-�jbvL�A'���E7�T�s�(�r[���"=zK�;:i�
@1ړ5_��֙�dD���<��v޵�ޠ=݁Ľ�����n��Z���#v�	�b���	�t�R(*��(k�ºQ� �By«�W�J�]�˙�Nk����eQ��{i+��!^b� ����N��<�g�M�˓�s�v#���G�9�8W�h�Gı�2�.�)hb^b#���[L1��bL-%Ti������L��~ψRv��aΖ��A*��o��h�`�I3z�9��1~�q�y��L�%UB	H��	�0Z��Y#����߾�Y���z��iV�}s��)�@(go�[�w��L���D�����h�����F̬ ��q)�X�ibă?����]�*���<����j��s��+���q27��Y�"v
Ss���b�fp��{bj^����}���1Ȍ���r���*��K���+�*����A�_6q:�	�n�V2L.�Y��j�M��R��<9��|��%sf�U���� ܩ��bx��<e�G�>�@�W@[�#����b�	�x�<l�-�JP�L$���[���Yx�:�-�x�F�m�6_�[�T��3��������6sjP�>m�p2Kn���8�F:z�eߨ�2�Y�Xx3��G���H*]�/��=�^V��0�OԮ�~�I4�CAjF�O�knQ&%o�h���=g|�#��V4�8������`32f9����׵"i��3�G5�.΋m�'�E��ضfXكS�׃��1K����|"���ۇ{ʸ\�xh��X4(����,��Q	һ60L �!�g�~� j
��Rv�t��SlC<�3[aZ���`J��M�r�s��L�;�d.l�\\imq��5.�����2�F@�w���G>e��c�%�ԡĥ�/�9�D?6t���	̠E{�U==���3��b�tT���=+��x�b���IW��e�D�"^��B���tz�3Ok#�)��Q���桴��1M�x���1�:O�{��"}-dF��L�E�V.B&I�h;xk�o�j�5x��6���ٴ�5Q�ʈvOWE틱eB�����c;e�-�&���)y �D^?��wҙ�V<Ą��7�+��$����;�<��"x�v3Ȇc��_�(9V�u��<`⁀WQ;�3�s��xk7�U���/�V�����C�-���?�(��b`H胰bw%l���Q(/�EZ���O��^%�=2�ɩ㢷E�o��:D9���v�c=������NM��
�UEy/�R�"�
G��B��"�#&˖��h�:�D���~LoU��@��4㯔nC$ ���
�SN?���E4�Դ�gs��Z�с"��S�ts��S�:k,Y��b�k��ؐ�	p�&�y��G*,¯���{�hQ[�V�u� eE.t����{�������v��0�/����G?ifv�Yl��~	�͹�i)���tq�J�ܬ�yH���K���f��#)���/h���)>_��Z�N2�!\�|�P0����\Kvo?�>q�fwY�6#9"�<cI!��"6-����G�<�R9�S���jĄ�	�2�3G�Oi��M�֭�>��Ja�����W$I�Tq>��t|�'��-���U�ݵ��ը$Y'���{i����"���L�[�|6�4q�e�>ʒ9,c#(���OU�����A>�Pd ������}SU��~~���z���Tn0@?�k�{�Cp��)���Y �p̆��WI��� �#�j�wB�=�j})�6`4���xKY��f)�H�@����d�����H�Zm�Wt��&E4+��<w+�/��W�I� k�{�n�f~X���`�v�o�*�dhdk4�S�"Ꞁך�W�C�U~9����V�KP�!�~���
m@����l�	���n�r�_?�cr)�Oc@�L'άO$�ə��V�c��`?��T���3z�^������1}_ٯ����\h�Y4(4�QvJ�:��kB��x�݊���Ŋp-DQp>�<�d��`k��R� *�9jDafM �k'�����[��Ƙ��.���T�<i�.|��?y����[=����!�Ex��|6!h@����Z
���ᷢOp�������������~�4?.H�q]+R75\uԈ_`>3�����2� �0����\�Q4 �4���c7��#����v�G��&��f�r}Z7)r��m�$}М=�[�+��\I�G�Wȱ�bRE4����u<B��^�e�
b��`R�H���?��iyte�d��
���!Y�����,��s4���!�%f ���*��9
��/��~���7>F�;���`H��ڮ84�yDl�l��z=\��kd�o�HP��gKR��D��!�l�l�8����kb�v����´�7��E�5�42�����s�!�|�D�6�C���浽�²��i������|��Ec�v;�+��vk j�[�.�s�ѫو��A����U��ؚ��r���|��G�x����ZF��g�P����ZA��^����ȫo,�?��a�;�ƸBw��/w�'b! &�kT�hHz3<�+J���t`+PN)��L�nRc򀉥W���t�j13E&��	�)�f@�^Y�ͰnPc^lkL�q�X����h$��p�K�3�b3�hL@�B�e~�JsŪ�\�x�Pi4o\�
�5� .LA�Q;f]h[u�t�o�J1	��{��rOiJ�i�"�(�",�f���5˛��͘��&����G�'��3���2��������;�H�gم �I0]���]���9;K���M�F����L�3Zg���m�3��u0�����q�y����%t�'�X��[�a,�@�l�9T��:�	7:�nO�Ғ�)�x\���&��$��������@����!8���P�_O��%�#�J�zr%�Q��sB��E�uM9h�Q���HWE�*�مT�LX1�('��ifտx��9��Y�`8,�M@�Bq�7��h�,�dԿ����DI[���]�ze\�����fY��l���2�#�s�u�P�W6��������Q�x`��`����@"����p
�0��͡F�6�}H(e"�"��^��H����z/���o�-�,#a�MZ����y
f"�o�Ma��0�yK�0QM�N�!�m'j�{���0~m�4�����N (I�\� ��߆ؒ�'�����KWS�7ZV����"��ވI|zd��1�/(�?b�ZfDJFdX�8��<?+gOz)`��4��m�̶��[k?��N?;aR��h�<$�m��b����M�
�ә����e��s�AF�Ѫ��s�R����N��? �d��U[]I���\�k{w/<$���$�Ꮯ{$='��K�������2�Fb���^k�w��R3�6�`W�p��e�!��k� �7��
�E��;��뉂[�XP���F{�-��&G��G�d�c��Rc9A���s�p�ޫ|��,��|שw���Nvr;s�7�c��9���1Js����b�Pe�u2Nd}���
W:�E[���j'����6p�͇� ���Q�p�Jqyc�B����eu�"�LZ�߸���ݷ��+�w�\��Ih�L�^�bN6�Ը�U��M� ו�wɖ����p�1�u#��4���a8 �>r�S�V��\(1�͋�-�-y�
��'���)�ɍ��z��Rp%��aG��s7��m4s�uLT�Oy��0J����#��k��#�\���^����u@�J�36 +�[z k�g�g�UW�D#x�/�Ohd>n�(	��Q�P,��QyBY���ǒ?z�[�����+�
�I.2�q���FX�`�y�K�s���I�4��oK$�fD_t��㔔�U�c�4V"\��K�2����x�tq�wl��>�3xk[�
L�%�K��(��.�.��wO4�Ql:<���=���ʏ�fN�*��Z���>��N2�Q�f��RJ��#��:� h�OI�����m^�m�G�Y:���b{^oIg\�^�QXT�cT�s��B�~���h4� wh�bp�����e��>��:����j�5���$�P5i@�����.�%�c��u\cb��\�VƥC�6�t���7Y�ľY�v�ad��9�v�e�42���L��g����zSDἯ�6Uŵ������(��Up=C�b�5��U�a�������"Hm�D�y���=�_l������]}JP��h��!�.?9v�ƃ�����ݪ��u`u��!\�� Jߎ���Cڳ~���kר�H4+�`E����{�K��!uӻ�E���P�:pn�le	��$�-�ͣn�� �@0m��.�Ɏ�8H� C�D� ڸ7o��G.H���1!&se�c�e��'H$ԣ���lE��=�!Msr ;3�zM��~�hO��D�mw���)�*��U3Cy�[�F���T��Y*��T#6¨���7P��\6�U��]�7՜��1�w��G���2�*J���u�^�䮯8bT�`~��ASף�@wR�W߽�M�9�����?�FX�hss��5&䷲A@$��b������\=%��8��]sJ����Lg�;6�jo+/?Hu�Y*�4��>�M܉w+ܩt�� zA[��0b��8��H(��x��	P��x������)ȃ��	�}J �5ꟑPX��Vu�6FK0����n;��z^��U����fx�2��Wu��3dju��"�s���NA�U�:ѝò�e].G��ݘ���눹��}�r��oXK��w ��-�,l_�ϧ���x��Ǧ�6�l���.!�T;4Hf��R����Y��>�/��k��_q��j�ks��T�7�PBh}.pw��A�����`o�̝&_�0܌
�h$q�JI]�z?���E���s�Z(�w�N��G�f�a�|B��iF;���lY��?�ˢ v��Eo_J��~�t�$�����ei��(^�|2]棛Wa�E_���ʢ�}"�R0C�����WK�K������!�C�|��K%�	�a3`�뛮�6���0U�`�`�\v1	���2�A00K�m�,�p��������F�c�h��Ѧw�Y���X���r�TDFJ�e��Ӽ����Xl��&�Y!��ӟ�:S�Y�Q�]�3T���8��ve\�E'ȕ�Fjo��m�'�O��'�Ǖ�f��I�`]Ї����g����hu�&<�όnF@���ddyQݣ
�Y8�2�^�R{�2O��Zh���2��U?��kC4s��5���v���B�aW�xd�m$6H�l4�Y�|��j�LW}(q$2����B.�/:$�y���
�ca b���d2t�G9�?1k��N&API@x����0g��1tm.$>~PR!�e�|w`?��"�\ *����G$�~�C�/{͘�+�# �BI2�B_�~�Y{;���=?�7[�z����rbh�`�wAo����}N���n:�4���[���Ҟj���d�rF)T��0��9��,���+\��^���f�I�حY��hbJC�L��iXw'����;�'q����zX�J팄M��h����5�^L�"���
�����K������ń�2������C����s�8�<ik��Wꊛ���o�TM������/j%��U��e_ -w�xT�p��61":����gnɆRc�Ms(�ϙ����s�����%`���F���}���\ך����@�V�LY�>�=�"a*�^�ָ�IP��na�В� 35/'(��Ζ��"�1=Q��S-��6V�V�mb(���YD�U�[bĉ��˟g�Z�M2��+�z�@���u��B�����Y��̞������UT�-νPIтn@�F:���:kڰ	G^}���hh��xA!D�T݆1��$���jOKqhɾ ��������J��w�9C�|�H���m*�[0�\�M����Շ��1�u���������i[��a��h��������=Z��K�=G���%���*��0!��Z��5�� �+�� ����.0�}�%������:h��&�'��ߙ�=��A_�����ֻ��j_���#r��:�=K~�
L?cn���axȪ1V���0�C˅�Ч�Q�:L0��*���!�� "����M� ��l�#>�V��!���Ӎ^ܓ@�Nݡ˓R��nxj�Ƶ�Fɏ*ir�=d��l5��V�$ε�!ׄ"�~�A�^^�5X��Tƶ_鋼�z�z�J#4��Ũ��r�(�73��hE^J����L*�"Ĳ�S;x[��B���d��Ŋ�mW�(d�Ⱥ���tI&��M��\&�W�Y��F�/�~3v�^�ڰ�	 �=�]y=������j�UKS	�����l��Ac�9U��8�⪏�� p�],& �D7D��)Tm�����N"KT��J6-2u��^� )��c���
ߟ�O2B$��9q�?g�e�.i���~�-��7�'�Drsilq�q�e���+{�Z�EM%@n�MIl-L�̷���rTkY;��?䧿��_`��N�dpu�%�eͲ�ʨ�x�*���!�!��c��w򘙑����߇L�����l��x�B�ʡ`ï��F��D�x���ol	e,6GxH���MiNŸ_�!gs��L��p��
L����a	��+���{ǖ,MP*4Ev��ݵ�+���������J�w�Ҥ��_
8k�pȦ�K��N�i� �������,,J/�E%,&�*F������s�$�EFo&��EWϕ�>�/�h���{.�IN��UjC��ЋsK���!iUnm��2�P'����m���a�J�M`�#R4w��^����	��+"� &��C��D��8����>lU�hhU��;:��܁�¦����ת���e1���#�}t�!z\N=���1<G�����x\:�ز��b�LaS���1�C>��k݇=���H����ɇ)��It.؏��R��{�����qhVwȵ����3�^-�q+P�U:�*��?\�S����] ��n�gS��u�XRx���b/��g�a�ﴻ�Y�,���-k�9���L��k��W^�$���G��r�W^k���q�4�+&+w��'	׃=L�>��͂���`[ nd���kN�]����Hp�#��sj0=-����r�p�o��TG/��>|m	$UN)l�����/gۚN��)nm:�\g�̾�7=܍�P����Z���MB�V8<p�2VE �~~V-oJ�D Uo�n��'�/���U�HΛ&'7J���}q�E�@B6C�w��jw����������Q��^�u3��0�r�y�KJ};{?u�ѫ�[VBx�{�l*��_$�m^w��e�#v��M<4�-��
R��X�!��g�� ������_���y�l��6��u�$N��Pa�"j�f��i�K���'hn�V��/$��'�����n��U�N׵	�R���%��D3;�����5v T����T�����.'!&�U��rB6���>Ƣ�4E�C���R��.)��	��<=f���x��B�|�����,�!TQy�����5��n���jkcP����㻤��5Գ�k�n^��Z�8�
Cw�!���'r�ڿ���I�ޔiQH��"��s���I�q �!��4{8��8o��`����ҷ�3���Vƕc��6/��Ǟ�2��5���jF(� �<T�6j�a�i��S'�>u����D�'@D�rMT^��������VvP7E�o�狢�L�kz3�୲^��\�A�Eh���%C��V�vD��	�<���<g�o͠�a���7����|X\��1L�^z���e#'�������2<%L��; �wf[C�-��F�\Kz�ؔe��I�+�w�<�Y2)��|�_?񸆛y�ZjNkh���K������Y�xTpѷB��}�54v�NǨֱ?��[NAu,zT�S'�3~��/G>����z�$�/*lة��b���Fdl�#l}����$�X�҄`P�[�w�LXѧ��#�d��I ��������4�{7�����V�Phk"��� ���Y�so���N�p
�ʇ{�>3~����`E%"������7��,gfs���zO�<�x;G}��m]�?j�Agn�f���(�[q���g�VcQ#!�?+ �
� �`8��9҂Ip9�]0�6�*i�����A�@*��x�Z\C����<"ڈ�
Ыu5#B�	*;���o��r"C���T.y鎸�Iy����Tf�
+;�4k@;6c���S�E7��V&OϷ2t��e/�5��ɽ;D��H�.zڒ�"-��� ��ˈ��eA�',��w�-�>M��$��;�������N\��$�mxtr���>��.��7�<2
�J�?mrޝ�n�e ��.�r�u��C� ��Eؔv�iK�@Q�?��$H� l�_9$�'�o���D�j����?G`�I_l�!m��j�1�V2	 Aп��ڈ�Т%�6}��5�_U�?��Y_TFc\Rz/LlB4�J���\�R���s>DI9��댜@yt �Z��rA��1��������sV��,�+ȯ)�P��_[�h���)4.g�����D]M����joj6�17��L��"��g�gެ��o�y����0e-�:?'7'z��īf��\�wC�}O��K���Z��������$�����R�� /�.������8�fF�>OR���Ek^9���̧ʅ/�:*��ak�M䳤�ƊR�S{���t�́oq:+',���N}�Ѹ �������N5�
5��!�?��P9��H�U���$+|"���f�����*��H�䕜*tQ5�=va�QX�٬��:0�5Z��8��fb�N��A���X&ZG�{�k
�ۺ�lV��X��;vO�9{z�A��Σ��!G#	¤3J��Yt�Oʶ� ��a��������	�����-�#�����%���6Y��g��jq��eRW�AȦU�PX��ۙ��n>��x��CvӬ(~
ms�(�(rޢ�����6`��;��kI![�#��jO�}��/8i�aw�}��'caYDP����F<y�?X���tu�����:@��Ad''*�W�w&�sqԞS^/��,W���u@��_� �a&��]�]��>� P��]у�uz>
�N�>?2K5\g��!P�\�����`��7�p�eb����e�)�UQ (rU�G|�[���/%U��'$�K<���޷+9@�B�5��]�1K�~�H��F��4���1�����ţ�q��'�K���[̞٪ԡ�G�p�XгN��� �[�J��9���2�*7}kv�`P�B�^�:6��$��w����f�p/5��x��,����t�h�l1*���Lh�,��3X(�����WG��"�������k��TEc!g�l�����κc�Mwݘ�����G@$�/?�Y�]��Ս��!O���K���b�V��g(�dsT��op�ux>���q&�d�N����|*?�`������nl}ҋx������:��~�K�*W��c�?D��}P���Jm�,��cʶ������%�۩-��n���2��5�V :�D�Ci�3�w[Y<��p8�$lݭJ܌ ���T��th��Kb�Y=x-��S;	i��%�÷�I�n���[�'�����H�m/����Dm��f�a\g���=Hc8����-y���j(S�����D^.&t�N��y�h��N�2E����Y1x9�l�.�^Z��ֺ.<���"�Q���%%]���-Qν�i�XŽft]�����XU%�g�?qPg��'�~���j����N0���Ϣ���J���aU���Ȏ�5n��u�sz��u'�3z��x��Y9Մ��n<A(��'�{�/1����-�noJ����
�^���<k����SW�ŶQ�kE��h�z��K����mTn'h~�T�@�}e�ozJ/�>Ĝ<�6QR��<a�[��A��s�dql�\f�r׌;n��^&�V��e@�ݝj/i��ƪHo� 9���)�t���ϝ=��� [�C_��T�̚a�Q�S#��y��+`Wb�����a��&��D�ݸ]�	[�>�H��0��s:�c�������]�K�>X�,e�L����KX+�'M���U?���L�:�������0U��d�:�T�f/F��J������H��첌�O�T���~^��l4i�;�qHR �tU�m��]�-��o�j�s�X��afڿ���\�.���o����yp�&G�����T�Ͳr��ͣC؁��IO�6G��V�9> K2��ot�,� �w���݄�[]�{�=I�;x؄r&U)�r�<����T�D��O �h�9�����ח?B�x����)p���O��/ۉV��{UbF�p-�#F9��Ѳ��{m�}�e�L�_G�y��7f$�2�A������ˊ�$�\�<il��Y��O��(�>w�	Q�6<�G��ɯ:���1+�ghg����ץ�SՍ��tQ���}�|����+=d��y<�Lr�a��S�7UUؽw6-䔔5������e�&�����0�A}�F+W�##(��#�h7��:�s{��4�d�eyC��y|%P��Ԉm?O30��Mz{_(��L
Mv/�V
R���C�̰'�{	5�E4�y|��6�]mp����\qb����7�0X%�?��&AI��|�J�uU�\�ʹ�5`�Ǧ�����5O���
��V$bs����?G��h�%�����[i8����ᗦN�Czo~t>�=�R|*�9�.� %i��?p$� ]�o��;A�hb�L��G��� N�.K��<����ͻυ]��Jf�w�/�dφ�d�$�K�~�c�Yj��?s����nQ����:����c��Smi*㟜�%9H쬤�K8 v��-eY\�֠����tq��OpyE-�q��W�@������	��?~b��]����>���욠¥(�t x�Q�C�l�?D9sI��&�[�SL��4���1z�NW)�s�mf�\�&UX�pW+P�c�:��@|�u%�q.)/�K��AL�7�G���w	 ��
��L���2F�e�v4������\�*xoŒe��s��-t#�nvc��~��f4h����#7*T���s1��¸�,r��-r��H��>"��/:T��(�왡��(G�G������l���Ѹ�k�#���̑�~�A�*��Zvp��Udm��p�;��b|L& ��z&t%8�v�'��Z�j;@7�C'�NGܷS�5`%JU��Y�^���m2�����L+ѵ'p�Aga�+�+-e�%y8�{sc��,��	2S�Ɔh����$�(�`x��A	\��D���+a1���/b����!�ظ6�5���L�~ҍi�ʝ����Y[�άg�a��WX"��D�I�	�x�EƦD��P*��wuqmg�������J��m�CXF�� ��
�ѱns#��aQdw���hȗ-��h3����oR&�D�@�kUB�J��t��B��
��h������#lT)��ǿ�-+I�xox����#�%2��"�X���~��C���Y%���ξ1�ʮ�_�e.>y�>�+G���Lߴ8�SJ(������l���j�AD�s�����23����{�]IJ|�
�A�þ(0�J�<��M�ۤ��P�n�T^g�Bj���2�ű���}���b#�\���)"_ tW��6�T�y���H�ȄJ��!�*t��V�#���ڃ޷�3B���FIkhc���6�����-�mWk�x	��xi�x�����Y�w{��WƏp	���A,�+�7���$�ak��ݧ � C�b�2�����$g��`{�t�08�Z66�v%����:�T"6��˝�P�+	�F��S7����f��U?]��� ���Hk�uAV&�߿(��WuT���v��`��Q�8%����6ᯬ���>]�$�s���l���^h�V�z��K�M��8��"���Z����V0]����"N��5ʝ�Il�	[G��B�/ �R��"�ݶyp.�fl=�bp���.%���ķܛQF�h>@G,�A8]���͉k��B�z�@��+�hJ̷�����^�_n��&�/!(4�s�7��<U!?/aX��������#D���s�X��Ci{��f�>���*�3
[D����	�W�&"+����[Q�u�9~�U��Q���<��f�� `u33��T�_���&$�?����,%�cX��0D�|kR!	�U�7H���+3�*��J��-��*�B�d]Ǧ�4�W� �x�z�����[�p|8�h��\q>]:lM����l�4|Tu_��*ӟ!rd��O�7��(?�G.C�2Fh�d�.*���O���'f=�R����*�
�Hݕ��e����P�*lja�~�hzq�����<�Ja�����&�C!�lj���l5�-dS8D�%��h7�8O�#��GZ�'Đ!`��b��鏇��ߦ"_�9^��7#y�r�����P!+���/5���Ԫ�%�c�ʚ,�iU�kB�ל���@y�y�u{+[lL[14��7��*��t2c�@�2��X����g�C��Hf}`4���_�n��].��rs@_E������AOg=<�?T���7��Uu�X�>�9������iY����/z����5�A������gVWˀ9�}9�L�Mz��3���N�p� m�20&u�'�~dn���?>�	��ڌ�X�g֍D4�viz����e�.7t�+ڹ�A�H?��q��w�X5�`#4Q�}ac���9~7bQ1{\]j��Y2�eQ��>���T�qWk�n30��HS���!F����Э3�Z̫(7�#4&������j�%�1pƝSA���/���d��J&�Y���K͔c��h�l��%��_؈� ��K��!�nNp o�e�!�	�n&�A�V��"�7�7����@�阶�祧R�@���v�b���ԗ�j���Ȃ��+����yg���"S-�D�s{}�j��������0~��KU��*j<K��Tc7��܌��Me���ƃ�2��-v9�<8:�L���к@!�`�L/�ܡ�1> }Io<bl����pَ�ٹ�SJI�@赹���2}� ���*�/�'�������r0!#}=[C�׌60[��ӟC��S�%���{�U=���\?%��<D�snqmT�k����+���ۛ�M������l��Q��s�x�X�mo)�
�&<�ne�<�j�1m�m	_&�L�]��EXFԥ����6Qe|�.�hU]��X�6�}�T�6���X���"F�M�IQ�(Ȕ��O&�����5�Ux���?B�n�_�<'$!_�-cL���Ө��PA� �k@�gܛ1\�U}8�eFtr�q�J�U��`�4Ԅ�z�"MP�>��B~9
k{��Qi2�o�rÌ�+F
:�SX�!�,����j�� wu@Z�\5��ϏYh�؅�PI����A�PV��8����a4'&@kLD%��`�H�=��d�?-���1�z�bH�{΅�e��6|Aג�o-�PL˸��ɼ�Bc� ��!VO��q��X#�������2)i������*�oV��|o�;F�#�����S��?�Xb�1�6�
���
�e�TƊ_���!���7�Њ���ˣ�I<�Έ%��z8c�`�f�C�ӡ����N;{Q��֞��ᦲ�H �����$��"~�YX�G��*v�t�9��~/w����ۍ���a����*r��-I�(W�\*孇0<�s�G�@�@h�vR����ՠ�o��2�8��)�6[����RQ""G	�r���5B���O��>�E��b�K�ޡ|b����d�1ϱDY̏�6��G���1&͛�����ib�(`\�e�9��5�L�R�����8�J)�7E8Q�ѭ}�M ��`�����`J{�j$���1��=�y�������=r��K�j�O��\�G{�(�����4h�t^����Z�~kPȄE���A�_8�6���HH�)�N�
0`Y[�Z}|*Q�Z{h�	D:�)넨Z#B���];U�gM��(w�E<ߓ1aS�]8/���'�j$�+Z���0),c%S�.;������Z��F~��W;�uԸٹ+�j�h8���S�M�&�!ʁ о�+�o����g�m��c�#p�xQI�s��2��jxL��r@�Lʵ�Ҭyt0��쳁o��"���P֋�a��]���AA�Ju�Vݔ�*M�b��"�#�02�"((�y�a>)�&
ⅇ ��;מ�����sLA��r��q\(�t�{w'����)f�[�Y�b�ͼ��~���-5w%ǯQf�n�Z-��=F�p{��2U��ڽb���#r>�:���o)3
��7����5�Q��
<�R�_�1����送�}2\6پ�(�=ʦ�b�c�@��ܵ��֩8+��0M��������a�w�a��6�C���h���9�S�P�� 1��@4B��_}~�^��W�m�|��Μa�&#=���ձh�w�u[[��Y�e\yn����w�r�0e�E��I�X�K��u��1�[^�!stU���㣐��V��4:�gJFpѶ����^2L��Xx��c\�s�+�/Q��eX�A	t�k76/��('!J5�#�1d��7:��eD����O��KU����z�����R߫�(le8���d�x&�oe����L%DL/��K|}��3�C�u���be�1}��\�
E6��5!Z���{Q�G�|���5�́ck�
߯���94s��NҊ��C�Y�L��4Nk�N�2���F�0`R������!z3���j0-�u���d�ޕa}�x�NS�"�&�kn����P������	�/������P���`o��GB�X 5�ڌ���Y����ٓ�r<d��V�v'ʹ ����r�s0Y�ס'�S�Dٺ��DI�*[kQHb���M�ke�Wc����.���aWN�ǰ=�b���Èɿ��c���W����v��%�#�D@	�,�{#e9�%G���\ѯ�4�j�,v��S+-
wT^��&�A��ۛ`o��U�Z�%Ae�j��m`�λ[��#��M̨;O������z\Z)������w>�[��(�xh��$�������3L�JW��a��ҝܟ�U�9��+3��B�*�Σ���0�
Qt�X����(9'8�;�y|�����F(jo�~fuk���g`��㩋r���*|����6��]�g�F��Mx�
���i]̩
�]B��zU��a�2�O�\���ʋ$%J�k�ؔ|>]HEy(������r`!
�I�c鞝�y�ݫ�8�p��@'�艽X�D����@�ߍ4��з�DdcS��K�{)�㘦2�r�X�[�rd�Su�<D�3�)�J�_�E���aO�e��&�ԥF+DY�����0�2iA�&IY�pVQZwفڇ��h���7s	̉��J�O�-�b~�-��\��D����J�XU��%`"�]��C}�ʼ�D�uV3h��#xN�)��U�bH����3���y��G[v��C��.�l1�ڊ&qJ?�I����?�9��O����m�Ϙ�%���K�~$t�yߚ��g@o�GB0����%Ky
��Ř�H[�)C��.U!C��a��2ױ��lVl�˲���O=B��=�d�IN��8d�0�ӏ�D�Ez��HoY���f�c�!6]�4�í�y��D�B�Mph�i�{j��O�����,y@d(S�N5�͕���➍p$���˼@Y����ËI��V|����,��A�G�P`�44 ���\1�*Q����|�KsN�f���3"�� )��-���S���r��h�1.s8�����c[���X"&_x�n����R���kQ dyQH��sL��T����5��EFEh�1%�Z��,�l,�[)s{�7C��$vz楖~���&6��]>�+�m�-ӈZ��L�x��AW6�F>�̣�5^���h�v�i�2U?/��q	b�5�H	�{|>���Ṭ�DU�[��y
b�<�R���dZ�v�^Ug�Q��.ܱ�a[���!v��"���G�u{�F��H디�fO�>7{.H>�4���I:�ܘ�Q�z/#cS|��?�w�\ӈ ��݉�T{�O����I���=���c͐��*���槱�#��m&��C��)g�-� EN�����fPV���.�9� �A;�9��Ϸ���ط�	�?
l�;�z|DD���1+1�ߗE�a�m1WQ�;�Q����}"�r��
<��Vy;l�N�D;VKu�q,`���6NO}6�73
´��<�7K�D�zx�Q}�~Z���G�rR%�!t��L���ǵ�����"3T��oW-��'υ�E��M�B�=)3�����Ѵä͏أ7\���?���.��N��.�F�GVq �����U]���Qה�|��w6u�@m�BܵRv��+e����7?�K��V�L���:~p��xLw�jy@Q�ݒV׼��{%
N/��U�����\;���WO��+s���\������A�~X8wj���v�MJxlZRj���
�{�;[[��UNB��f�;�D�-�>?����� ttN��zO���tፆ�	nM7y��H<��R�7�u�Jwj��Q���Y'���:�r���F�x��q��;��X��g#�H�h�NH����TF@QYɮѼN��)�a�'J���)�#���V�IG�7�k{&�u�]�׉,��+�C	]�t|$
r˗I��ݔ�����;���}M��vȾ3������ρ����4P�>�g�O��� ���%[��#����ՀUȱ��������)���-Df������yV�����!*<�qX܉�R�ny<._J�IvHy��!B���ʲ�JT+g�H1kS��kPB$Xn����h���	���+��&�0�2���0�Z���<p#T'�<���10ߘ����������*�J����%Ao1z5��f)��-H���f�-2���p�n�[[ߊUC��bkz��x��h@����]��A����P3����À0���Я�zi�����^`��}�'ۍ_��Z�ؿ��Dߌ)ֈ}0�iu�8�{�@�[�E:"���u��Jq>�>��	٭������~�yӍ5�k�X���"PFs;�jXtm�GZ.���;RB��"��,�IÀ�I�}g����~��~�L��y ��j��.RT��֎��<��"�#�93.� ���ڱz̯ TY��V��"Fݟp�N�_Bk]$]\�Iwy]د�u��7�H&Ę�.�e�<{|)�1��A)�����^5���� ��i3�]>z�*�$j���8K]��"�X���X�����!"��~VK0����R�%z����T���QKl��o�A)gZ���B��3�z��?���
��Dw.�9��|�ݜG�8�V9Fbk�a�!`t��.u���Uy4���L!��\�T�Ϥ��p��~뾅��v�\�Y���z)/��o��Э�mbž����kH��xD����D��r�َ#?�	"L�|T?ʇ�Q߃�a�(*�u&�Ծ�n��vM�p���xa.��>�4�,�f/�'�nEbՈA� ��
��m����m�2{Ō0I�H�!��v"��~�V��,e���V�.4y�f����r�ĭ���J\��)��:��� �W��=)���s��[)��EJ�=�:���mk�ߛW��עz��mJ��]ذM�%�OхV3g`����6������ �Wy&+!�P��7�ŧ-Wε9!��C���[�I�0��j�,	y�%�G�W����0�0�u ݬ���/�/�;����D�>���\챳ݑIXy��8�R�>�}���N^��c���1X�Q���BI�ۜU�
��T@������M;�}�h�A��߃�%UY��p�w��;e��Ĝm���SAJ6�_���s�]9m���d�g�o�om�ǬW6���W�M$�ueo��;��x#��FTY���)��]����Oʦ/�G��g���i���4��<3�S�4k�z��X�m`�J���7/&]5���;x(?�0f3��22�J�+��X�����g�2,�n.u�n3���i�X$ӥi��h�Cg6S�0�E ��\�tv˟2HQ�_��H��O6����"Л�ɦ��,[OsiVZ�Dl��|�F�ہ�:x� A�?�mӡ�r�0����9[_����g��TW&r��*Ps����Ԁ�����\�_"���I�w���)1)�3N����pNɑ 3��y����{��Ě��������֬���� ��5�!��g����t��	�Z~R�{7�'�����yG���k�Y*(�w�ɠ���A]S�@��:�/�CTj�QX��mI�O2��jf�'Lyf{eU/���C,�!a}i��a�q�RI����_����X��T��$x5���T�9���N�E9��JIf8¢��B�[��	�Xc�O�����\��L���S���D�ɒ,@�%��j���If��vq�>�s�'��XW��pے��TI��9jx��!1�a�\�˗Dh:{�P$��~�b�:}�_# �ف�ު�l���EI��~�r�	���vOb�V�|�4�*�=U��i�&n��r�\z�V�8M\'O�/� 恩�n}Y�O�!�"z�W���6��w~Q�ěB�%\�da�)���~�:��&���I��y�#��/x�ȶJ~X��}�xz�0��ʣ�{�Ǜ����(ȗ��l��<�2��ױ�y��:q֫�V��W�W&�>S��݅��͕�.N��?r0k�����g f>�NA�I�V���^������o� f�H&��J��F�
'�ݴ���Tn?�BC�
n���pZ�d�Y ɝ���t��R�ڀ��G#���m��G	� ؂�y6|��v�`/cvXo�Oz���<��śn����(Q�)(W!�r�b�==h�s3dӵ���M]vb*(�q:���TR�	(cE�{8O�|8�Ҏ�/���P�w"�����@ܶ�0]/��%;���(`a�D��`7 _v�v�2{�v��>k��E_�����X�t��	1�p��<�J��6�"E+��pQ|*񤧸���+?��c�Q��Ԙ���a�`"�&e�K�Fm+�db�զ����	r��0������;��Pײ}ߠK�X����[fY��ゟW�/�b�/{�Vj
��O��/�S�N�7�q���C9ג�+����PbL�e�smW�Mt%c����"}.�f���.��W�d�A��d!N[��N�&$q�2�GW�A�U�`3�_0ٹ����E=��u���F��z�i���FxS��UKn���\t߂����'�.����3I/���|g�=x}�x�����3#V��(m5�yM	Vfu]��.�b^Dl�w�rf�֠�� /$:d���V�J-���6�v`����f�	+��B`Sܸ4*��e6z[�qY�5k�ke�_��C����@d:�w�Y�q�lp����Քt6����U�c7�$%�$������Y����k����-?r��=~����B5�$�?;<^���F4�ά���-��]�7��"n��U����7�H���p�M�}�-�,0r0%�l��_K�G���]�'΅��A,��y�/i�<�y�R��Ѿ�����r�������д�����Qr��K�S�!������UX��!1m��;�Y��^����]�T���=i�~L�990)��ɔP���؇-})���\2��/�lF&QdYs5@I�l�'�4@U�Udв��N��j4h
��G�:h��;(5���eK���	~��t�Q!Z�z�2�w�#��i	m���,WX]�Yl���ñJN)o��:��i��է�v2LT&
���%��tj|O�q�����9u$8G��sl��y�6	��=��φ����|#$�Z�&��.�*���)��s�ş�37�V/Ӳz��c����9�Bܺ���(��Sh�mM���5��InQ��
YͭN��a����C2�\��% f|�����:i�b����5ǎXoW�GqrN0���/ԫ���\Y���r�)t���2t5�sX���n!�W�B*;�k��vV��;�奛��A�K(;%t
FV�,������i?'ɋ�BT��$}tWW�4f�!%�+۸@�7�ƀi��7�/�M����/�7o��O��p���/�ܱo$�/����*�ħ��20WJ��j'xV��Fj�~I%�;�TO�Q�i'S� "����f��V��5�sy���%�1ǚ�!"��9\�+�ħr�� ؆��S-5�`B��v�O�������D#"kU���:����'Ih�8 ���%�!}�+�&��_+���zF�;�z�wN���������X���^��c��pv��[*�ve^ς�
���J�)�w�\ܡ���;{ï��f�R�~.�N��W]@����c�3�/���oɤ�	c?	���A}����~j	업�%�6F	�8����7=mH�j�b��^�.��h&��W��M������!����n���⁽ОuG��o�J�è�;|�-\��m�e��d��ntO�u�PLg]�@ �2^W��>�����0k�[Б�j���P��V�s_L�z�9�>������YÊ�0\�>��~���]�(��4�Ӟ��c�M��?FG1iO�9M����v�*%r��F�d�e}�'��>�>�?�(~���ĉIJ;���������҃��N�*�ћI�(�8�vQ��k -O��o�A O��8��ꛨ�u�����6��rk�����ܭ����U_U�8�4����X(	�IM��O1����Z#��V"���y_�7c*�꾨����|Au�EQ���'�P�Z���$�Rs@�T�i],B����^��!^A�e��C6r���cnJ�ST���׫U%<���z1!h�p�R�����	)���~��t˩Z���GG'�ܦ�k��	�^���L�1щ��^F$���x��=H;�Y\^��+�8�=N��Ka#�]`�t+l�y=���Y��Oa=�k�e4�)�G�?!r�d?jK��E�q�w_�u����7�r�W�ŧj�ܟ3�V�IL�F��� 	}�<ف+ށw��|@>b���>���o�u��{�4�3}Q'�@"����Ľ��~�g�d��L�|���!k����v5u���!ȀvSL�o���S���??@\��~xf��x0Gf͡�"Z�Ogm����@8�	��\�k+�Tk����f}�]c��,�K��r���IG){հ�!���#h5��]��1�D��s���t5��S.��o�P.�f85��S�hw3\�j� y*!{��d��ڬ�.k�G�j�9=�P�XR'��ݼ�H�	���@l�y3$�J����X��c�AF)7ͬZ{:�5���<ņ�C&[�]vl�����w'������&B��"�ۚ΅�t��2b0r`f3l-U�����&���q�1zr(�6N�T���4RaG:��!��Lߜ־د��tD����_ �)�&�����Գ,6�ĪM!"��SלuD wb��o�u˚$>@��5�����TG����!Y�ͱ;�i�#s.�YҔ�hCy����i䰡�N������z�}� �l��<����)����>��<p��4��Fp�����Ϳ�>ip���-3��M��%p]v�"0�� ��t��7߸ae1m^,�Iu�NKVs@z�(�$�c���j�ѝ�so��|a�.��w%��{�a
�w�1�l�:5���Pά��}��j�軅�k:��Ȗjo09�Z-oAn�Q�Xk82WVq�7�����aqnj鬃��i����F��AM)�����X�	k�
b� B���J��3A���<Oa�	�l�eDR�8�~�U��J��J
�������5�{:[�y����A���������8�&e�t;6�ՁsT��~G�4���#W<���W6q%2�1mW3�G�J�鳳�Ü	c)e9i�<�W	q��DB�o�^X낳w�?�B�����q�->��<�������(���v�9��+�>�G�#��}��p��.˄��Ɋg���.@n�ϔ��Y��(�q_�� �\�R�ro����F(
�=ꄻL?N$��s��o�RӄS�e9a%�.M�c+6��DL��5����&��/_gfI�P�ڜ�:�I�+�,s' ��#������qUVΗ ��e(	aE�ڲbM�8]�0o�3��UY��n��&rp�V^�4��Un���̹Y2|�i)�<���ީ�-$̍ol�h�J~K�r���Q{�N;Yk�PG*���E�7ǫU��>l�h �� ܵN���Yl��6�_ڀ���R~��wy��=�0%�̣\��9��3@�HQP�dF/� ��g{AB/d^tq��/�|���p�8	$�[]��air��+T7���8�pE��8�`�f.#b�>���Q��j���Ͽ?[�� e7բ�$�b��;2j���f��M��A�He����eO�W�Uk�a/Al�L�LNٹ�SƓ4%��՘#F�Fb���������z@c�w\/�:L\@sz0 }�UJKs��E@��>�G��7�w���淀'L���t�'�6IH2��G��� ��|�t���qۋ���������c49���z)�>�_� ���<p�[�[^b�&���^@���ץ� 9��F�.�`5�ڟ�)�Mk�{t4}��k9n�\�n�Cj����D�q2�2���>�s��Ux{�|!�?�b*}ы�;�#��[��Zs��rv]о
h�R��J���෕ג�0�,�{�n��|�8j�h�V�@�����Q@�[���(�{W�G! �<h^�vtD)J��e��յ��+�̀���Е=�Y�چ������0;�j�O-�}���$�@&�b�Yr���G������ �Qd�K�q��Pï��xo�FN�Bۥ/�#�2�43 cY��!"a�U�b
VŒ�c"��i-zÕ�61��Y�j�a��_J1m��2����g(����.��$<�g���W&1Z���}j�̀�H�d�k|�x��OE�V�A�;k��Q�mOhI�OY��&���l]��8��$���[�ea���&��F��6�'�$6?{���֎s��<Ő(��C�d�A7�o�E5���f$�P����h�<���G�܀�M=��'���x7v��*�>p� ����	r�z'"Y_��IO�6��Q������'����K9��i�"�����+���Ʀ����y(a&ݸ� ^0���5�&�����t�V���1�7�U �h���)���	�yaF��eʋp��z��T��ze�O�e��%��(�qu~N���K�z��}��Y���L�5L��Dj�4���\��W�����&�ӡ��|���BS��V����=�L*\=4_��#������,��Ee��Le'X{���Z��&�;����R�?sj���+��R��u<��kИ~ gU���a�gفj��=J����MiO~_`D:����3�B��[�������`�4�{�� �a�l[`ܫ�b�r�o�[���"0�m��6�H0��Ia�C,LQ��q�X��@K�7�����*�F�������S�:v�����R7�fsn� ��1׃t|Y��ߢ�f~&�̤7W��Y$�RX���#��{RnO's��fm�>5D>ʽC7�B(�t����s��ЂC�U_[=�-���E:�-ēX}��-��|��v��7a)���M�����c�u��l�'��OoJ9��Dsi�e�{��'��
�m��\���u?l&U7rY��yc��b���9��dyY�S��.�<
���9�߷�P�:�zyw��
Ĥ�	b���>ܜ�D��8���_����mcy�� *��#�Nc=�r���J˯:�$O4bHV�Z4֠��m$M��6"�
[����k5�~ck�J�\?�a> �"�D �JYJ���%�uA�#��d�~$]U������9�"�
1��>�ꢜƁ�Oec6"E�]@�E�\�{�=�Ȃ߿Z��,�P��v��5����i'H]��·��D�ݐw/&!�;���K	G>���8�kkE��˭�!�t�e���?�}�3"@11�,�F�0��.�k���9\͚�r,I�b�y^���A֑r�S�V+It�c��/��`@��d2�T�2��������W�Ʊ\:��0���S)�#T�W��pe���2�d���L�U�=������@ަe��j(GAc�IGz.�J�@z��U�rsm�:�fy9t��Q�+[��p�l���|�%�����Y�@�Zx�N��!c_)!Hۄ�}�@tf�5
v�޼j-1������P2�tN���
��2�Z��F�qtLU�WH"]���+�Lfz�W{X�_Jj2���&[!��'˂X�	+/h���T� k9�&��k�A
v��B�f��R���ޓS:|_3:#V�]�e�$f�E���������bQqˣB�U���W���m��j�����sH�L�!����8N�"x{!?�B���*)@�"wh��X���>����:�R7U��-�HC���Y��a����^�޾[�?s��}ƴ�� ��Fj1\b�R�	e`w�[S�ky[�g��x��0
��'�\��Ϥ��A��w��xn�G?mE%���=�D�� ��O][Rr��e9U��r� B[(6�:N`�By8�)�F����N��S(S��\�A@V�yC/K�e�{��`M�>�!;��+�R��~�A_>�˚�w��_�UK��n�y���&Ơ�w\&	
�������=�E�Έ���$Yx�������O��P�H�[�H��Yܾ���l��A�j�%����D�6�O^sX�ݙsC�T ������M@Z��b���"�D�°A���22�%�<NT�*�|���i�&�P�u���NN���!u���ܷ:&�i1�jk(Yn�Oh�i��
��U��;U�X1�ʌ�lצ$1d�0�pzt,������U � �����;.��#+�{*��/��mi2��	+���j�M���p�mқpN!엀H��3ST6�>nB`���J����0�,e{�����W���U�Ey��v�M��+]9�vO�!��/{k|:��?�ww$�`!gw����S�u�o�>�FN�����dR&[	�ئ	��Z�����p2N�@I�{�#Y�<Bhѩ��'R�G���Kʧ쥞�G�ј�gPYdIK�Ϣw8���7�~�E �@+�I����h

�v<�~��C�l?���o+ վII��{�M��鴻��X��S8�h�	�8BsyN�l�%�5>.�Q�]���!��T�>ڼU���߯�di91[�q$r�����B�3���ё�k\\�tP*):	�z��F�??��Ò��)\p峼��Z���
}�F#h��{���!0V@�}o�҄B}
0�&��]�fp� Q7��zw"�0S��0��m���2�rnU("��@#6��֕??�
6xݪ��f��V͞骗d�,��M��t�]����V�D�R:�� ��L����0�Mŝ��sD7����ܨ�����\N{Q���=�f1�
�_��~�P� �aK�\�l�=R,5�-�����Ț<o����(���!�w����I�O�=-d���GH���%��l�ص����h�.���zv������^�#q�:������K��ʹ���̊=��O�޾洈�
�w܂~�I��_'(���AG�~�S7�+�$�O
d]qq}S���℀�-��t����+��(���/G������u��pG��E|���6��y�i��l�<�v��x`_aLXa3�\�gkN3���<��n�ݵ�!+�#9�[����=�c��<����Rߏ^�(��Z�3����GW�a�������tB�o����:D����%���'����h���t:&�̝�/K|�@iI�cv���gW�ݐR̸)���cql��a(\�F�+
?�:U��{���;�X7���B��Ɲ����*8[�����M���nÂ�Hh�Fs#�0��K�B�Hߡ���r_�e��*Q�j���/2��x:����c=�m�F�ȟ���H_�G�z��*��*B��]!Ff1�uX
���Oo>�6ݏޔ�0_O}��/:+G��`���5OFY�5
U�Ɉ�;@M���� *�b�mY��*�:����ԩ�i�9F��?p��m���n����-�e[��N~��Q�B�9���;���=�N�;q
�d��2�K*
n���t�\��v��`H���2�V$�Vq:�a�(��E/ɵ�����|�L��&��	.{�����aW�������|��C�O��&>5Աc@��^nI��9
1�8LGZ���j���p��Q�􊁓?莧B�o���G{�:�E���|�75=`Z���XMڠ��ӀZ
7\|�ߡ3�2sq�#E���*���X�<�8�(���
�;eInS��s\��Ή͎o���<����K�tf�E�V�HO�i:C�(lT��e�
�6�W�~����*tB�W���G��߃k�-�`E*�}pB�#"NvK&��b��5>���d�lӖ�P`��c���^��8��3���� �yF�J�Cաȫ��j��;S�����Uj���ɿ$����7�LF��s����}���\���#p�KRȑ���g�X,$h����}}������P��RW��IE�b�"x�^ʿ�,D��i��M���;����F-�-�aÈ�d$Yh�����1zl���Z��M�Z��|�,��]��Ov^Q��f����s��GYyFF��[�2�z�hA�8�����6�5�������a�U��A�����Wu�@}���Z6��g*��԰�9"����&I,�'�g��(��"i
0���k��?��ʬ�J�#:� $��h��uj�6Rd�.nL
vB��E�"U�����l?ER��X?���qc�1���m �ؕ�N$FO�J�$�O�N����۫&WT�k��aئ1U�"�8n�7d:���?�j�����Q��}��$����r�ɭw$���L�f��!��ܟ�s	6M���h���o����CdI�5���V)�;����z�m�3�Y	]�
8�% �,�Oӳ��{<���L0���P�^2�U�zhaZ,C-�YyW�6GU�l�!����R~�8�a�WGO;'�hh�����C����˓��n�T\�-�2T�MÖ��n`Ш����{������Ƨ�iI�ȃ��>�+i�}��Ȩ��Lg{y�C�5�����H����*�!��T�ή�p�� ��6V%ѻ�m�*{	*��1���/j�]Ya�1:�\��_{��{9�&�'�M�:��7����L��t�� `�3��֑2@j�6䡻��K��0�RE�?!���a�F�A�P4��Пus�-�ݶ#�R�G��pL+�־U��,�Y�j�tR+v�-tI�"��܏::K��)\��~�f�K�Ե]�ٹϟ骎�93aqUw+�ؕ�Q�R�t���w��Ⱥ�̌ߔ�ͼe�0j���>��|%���������R�:Z�;.��5a�����?��박R�r)KU�ߴ�Kט�w�x]����?�i�U����Rvfq4�z�#��~�|\Q1?�фi��Q!q:@'E�]�O���>On��s�O�T�y��'o5@
�A��m��@�(�|�KL���Ӱ��?ݏn��/���d4L0Y(�y+vc�����Ϯ� �Y�t��C�-���`3���}\!��{nK��Zq��A:ߟ�V���H�[]���&D��)��-��`�U��D��I��4swYx*��Ⰺ�k�S""*�'c@��'�y ӯ�u�	쫤�ώ� :ew-)mT)��~КYS�������>��N�#��N�N�]����Z`��9����Z�5�tL�8���.p�N��X����ۚ�{h���6<H4��"�\��u+UHԛA�p������O����X��[���VT�X�,�wh�o����,PΕ ԙ�獣����f�
�����<'Q�^��%6&���jR)YU(N��s�UF��5>�xi���Pyj�=�w_�q!�����z&�~���辞�����M�Y�2�C�0/
<�K���;Dҝ���W�&���~�@.�n=m}#��wňH	ۤ�ڔ�羑���7�i.O���[��u��6�y�7t��}�x1{� ��n~T��!F�svO�h7���2��҂����j5�Ʋ�ļ�I8����1������?��/�O�q�C{;�ǅU��]Q�� ӌkY�f]X��	�56 A�A�o���#h"GeZ�[�-D��݅�J7�4�Q��1Z7�;��q�O�{,D�(�*~�{�Duz���]b���c�U ENE�S�p�D4b_����h&*N�Ш�t?���.V���ɏ���{�/ˮ6�%w+-G5��bt���-1f ���l�oW�>���D���k��@g�����`'o�9�˂�J3д/NǙ� "]}
��{�_��kq�ey�}���:0�D��V���c�l��a�p��e���%�yJ}�g�B��_F$ʲd�c�!��)��S���v�IHt�΢��M
p/��0�K�!�ٙ������Uk�O��Y���{����<��Bceu��r��'
,����x� ���1k/?���4�����l�|+�7A�]Y��7�!O�ۮ���5샿�(�@N$���#1��^�F/}M��<Nc����Һ�4�>yp���ͺ�������-fZM�������Όğ�o�����f��h:�;�C(h�k[�����X@��AK����:3�2���Ŀ��Z�)I�q��s�4�!��Qm7�;�0;l.}�qYiy^T�Q�1�$=Wi����L��Y��T$ظ#����;�Z���E?��<t��i'������*�G����Dvx�
�v�c�7B�v�^7��"}�Y>H��Xl��+�'*M�fJ���b���j-ɵ\vn)��NC�y'1b��	��D 1���c�U������-ȏ!��X��f�|~[-6)p�)�Z�]�H�F���~��p���:_��Xi�%�"�#	�rUb�m�u��r9�cm.�H���w��O�~y��/�46�ޅl�>�F1A��( 6O�b��k7F���ґ#�GWQں��sW��8�o�r��V9#&1�0C��^��Kqp\uك=�s�=��1�Lm��-&s�*���xAǦ����r�	EO����x���起�����~��e��c�"l���E��hUY�*�W�ٕ�AW3P]�tyQb,�+2iXF|��=Ⴜ
D�[��8�z��M/g���hU�[)Y+���h&^W���o��uW]�-֙s��l(�|eM�t���W鈥���K)p#�I�����t��N!q���'�G��/�~,�--V�7Q�`\M�ҷkJ�s�$:�T�	ӄb�
�C��~�x-�`�����B/o3772u�l����׻�;[�T|�@_�~�>��3��%Y�s�_J���+<(�tA�)h��*�Z����,9p�2�"S�sf*4@�Q�����`����2�LG���D �Er�d�	���Y��+�ew�5���/�;�9����1q���l�/�8����<v���>(M-]6��4#�t��V�OC����bۈa�,JIS5��dxI�,2���'OI<��L*��_\31���%L)�+9�.�����]ߟ�s.�L0Z{���� o��l���b���3\D�2�$��ڃ���10ֱ��U�f���9�G�D�J�_�#�o_���>�47��5�|&�h|?�e��G�9��Ȋ�@Brky#����xbXS��������,q�^��E��OB���鸎L��]���p{U_m�4���N�����7_��<d�Y-�#kb�P�w@[S#�@�[����"��z,MR�\.dv �j�0��9�n��Z��R�8�ɲÓ�a*V�`�]&��V��y�e�?� ��xƲ4�(Vx�1vn�"�����$
 B��1u��_��vF���};��F�̈́6�^bdY<_db[���G��V��b[��/!'�<��^�~�����\��FeL����ư����}�ɾ��sţ��W����(����˔8CJE����9�2�=tJ�ȍ��d����]�?��V9b������0�aVW��<��,Yg��z<������	�����ʱ���Eh���'i'��]�6��������`�{p�rv� ��H�1m6CD��U�HNj�P�3��,,�h��\�e�;�7�GH��_u�_f\W �_�hm �#Ee���
s{�|
>����t,����0y2�s��Ԑ��*IW����kF���9ZEb�&�R������O?G+M�^w!���l�� @�:�M�8��h�Y���W��~�4��ņH��s��+���?
����J�0�d�Vfk�=n؄~gH���M�ƿ�*�+# �<Ͷu����C�ZF��%Ԥ�M�$���[���M�0K;�0��1��Q��i/� ��=5����]C|��|<�>8ҧQ��Z�ζc�E��)F\>��V�7���")���r�$���dn�)Ɖz'du���${r�1�ʘ�.4���)
��&�B�"e�ntD_)Vw`$���a��
74��%D�4eކ��zH�Y�)�ɳ�Q�E3r���C}���H�ّ�uvj֘l�)�VR#��C�e�9o~N�s5'�U�A�,*�v<�UǄ
��@�����2�m;��Q�u|���s0ִ���R�ʚ1�A�sl1����@	�Uӝ�P��۪=~	�!h{�Sq��3��L�31�hP� |�aH��	�&�:�I�ES�Xq�$��	�F%&���IN\����	$���\��9YJ�}�G
湜��h��#�yfD��Q)��Gw;���!�
��r�É6H:�G�Վij�}����AH��|�����z���nG�ɺ�x}\m��M{�_�2B�t�E�^s���P0k�@���z�O	ǷwV�^���~J|D�vpZ`xa�;�HÖ�XCՉՈѤ\v�v�"!~lKȉw���4���'�8��<��]p�;
"�w>e�1(>�U ;8��B�E��p`W�[�S�x
Q�Q��mϏ��N����鹇���A��ǔR���1���ŁA�Ѽr��3	�S���W#_x>��&����,�H|�Eޯ݉˰�w��}X)�O
�H\S?�f钷騮���~M6��sB�	�ʘ y\=ȉ��$�n���(� �
�U��x#��a�G�~!��ܻS[l�2�B}�U�x�R�����w�&����.����)�6��u2���fUS��Q��J�*�,�$���6Qc��(��
čW.��Ϋ�ޢVLl�A�N(ю� O
��p�����Ȭc;>��&jzך�����A��p�:jԭF�;i���(�jl�bM�Y�⪲�9|{R �kݑ"�iL+_��r.W"���j�r��q=�����B@-��r.�j��3�zF�a�=6�$��5�>�`.Wv��x�aP������7=r1c����Hs���E�b`�M�E^D;o���щ�j��#�ft)�=;�C�1�ԃPȨ2ݳ�������4O�@���xC�� (_���X�t����v��)��~�9���զ�lK�ʢ<�G]‴�i��eϪ�&�<���T$�^�J>ͥ�~�����s����ߨ���&P����)v��+� o[���8��2�v�J�i�UR_k�Zu�4�U-#�-M���u7�Aؾ�A�P����B�H���<�0Q&�K���j���s���%��k��k)����=��g1=16��rny��.>{j=�oW2�U�Z� z�t���j���ҍ{Bx�JW��,[b\>$7��u"�{%��Cfҽ��̇��D����ՎA\�q�ۥ�r:����N��h���ti�f�=�-���J�,w@ݐAQ��I����K�3�iS�u7�t)��m ��W$��C�ˌ���hG1{�j�:�a����ھL�P;Fd*�,ӿ\c JH6p����AsI�AH���~�i���A\�|b��c�fd3|JV�U��f��Hǆ,A���װM�zX-t=�m!L;A�ؤx�)��8��w��3�(��[�g�݉�I]y��p.F.ِ�N-۠�����H��x�NpVp�6�	"�"��^Vq�ܚ�5t�	�K���R�eM��ӸԒ���{lҵV�i�?�a���,��XYE����P�`���9o��x�Y4}�\&�^Ȅ����ŷ�F#=���	���,��jA�d-Q�P�$���zٮ7 �-о��ko/US�Rg�=	�ze!��ts��T���������[k���5o�/�کU���(��:Cj�n���n�z�
���ݶ�1=�8�?��r%C����Q�i�`�O�%�qY���ι�о�2�&+���s��!�M�-~m3���/���\"��'�4uq��������
��1��;������������uIP�pp�����{SM����`��7��c��d}��J,0M�=��N;�us��x�!%���T��͂_SM�1p 8�CJ��Gs517 ����hr��7Z�]�$������P�h�[��q��ș�sR�V� ZLVvLS�RT����6��A�i�8�ge�4/���v�[�ѓ���l)�i�Ԭ݊�64w���aA�L����`���&W�m�O�T��G��˴/gcnf4�7���pr^-p߈������D_9 aq�8Ͼ�@}��Ѷ�- ��B)��1!3i>=����6�ES�����j;:B�e�z'��1d�
'�tj3T�eȞ�m�#��x� K)���>�]��!�12}�@��)��'�li��V.Zu��
#�b�f���J�c�;`�Iv|Q�x��V@�~��0%�o��'��=�{	�[m�mw�C*�������'���G�I% ���{9qM�Wc��(Vj&M��mK��vx�X�B��0���N�x�ly�aV��0ޱw�F`��p�>�%��4����(/4��>�$dK���eb������p�/ ���v�䔶f�s�:��b%<G�Y�����Y�EtUZ���q�bAfkdK�R�ů�9�߃0�U"�W/M���Ku����/���V,�"��W�^^��k�u�cy�A����:QIO���N�6�;ّ�ۜ���[����L<(� &q� w���"��8ic�v(���f��$�eB��D�_�I~B���Z�#�j�[M�
TVU��A�}~m\8��+8I-/V�?�aE��%����^Px�'���8dM�&}C���m�GT��;�S��k�,�>��+��Ĳ��	6o� X�U��c��y�:�L]ur'��o��;���͏�!ޖr���/��c�3m�;���A,�y���6"������%{���pT�C5b��$ �|]3$�z�-v�$�vEŔ%�x��O��}OD��ᗶ�O�m�Y~)��l�z;B���V��KE�Uv ���J�hF�e͓鿐�,�}|	"ΪH2�l���\C�Z��tZ�#<�̣�)�o|�=�1ɘ���DHQr�f��w�-��0#�mm<�k2l����%��z*S�FI���L��x�Xz<fS�>Nǯ�g�i�D��m�Nv�L���e���Nw k�����&ȱ��°1c��#'?���3D�w��j^Y@�����CZ�=a��e �洬{���������\��fC��X�f�Jǋ�m�k��rr���|�wc�0�{�aZ��d�8��Ɍs�l��&���x�G�ڋxk�,n^9�������1�����-�qc�Z�ZR�~e9o�yUd��é-;�A�m�S�������褉Y�O��V�o�y����� �q'����E����Si���*U����������f����;�X��c������Y�j�{���*�����z��_��A�i�\VD�iY���v���|�LB#��5�����&�
�ҭ�Ԃ��I�5?�k	F�&a�^e���w���m����d����'�����1���� w$�#-�D����V]M,ٙ�\���*���і� �fow�:�k�vk��q�H$��?�����{�$IΉO��a�[�l��i˫ә���������83T)R0i�m��������(��"����~��*{��=�ݓ�K/� �㸔�@ۙ�V����>��<"Ж��s-����s!Уv�wq� ��0�Q�N�d�~p?"�!@4]I�� �ıg��y(��/�i(#Z%���y�٨4���^*�R���D�Xڒ�K����e�v>#S=��a恋q����������h���>>�P��
*p��z�෴Q �����7/��r��B
387@^ʇ��:��Dg{�D6�oS8�կbv9�0m��vQG��<�xX;��{l�oA7���{rہ����� � ���+�Up'��d���n��"��=�r�*O�Q��YX��ݣvG�<^��ڼ�R�?S8����3�2�O"0�����S~�?����8Dg 
��mr�9:���ZO��G]5�5Q�'�<��(z�a����4=y��7�4���5�^���M�9N<�fF�N�|�H�]�p�����䌶��Җ9��	�[U�]x����8(MmV1QC��|Q��(o�52|nZ�g�����{Ip�]Oi�+�iV�r�-�>1Ѳ~I�U�A�f�d��<0H�S��Vnŵ5G����Pz4o�����b�������bz@?AC��'u��%�Q'������v_[z�\�#�N�� �'��� �� а:>K�!O}����=K�K��D]@��vC�c�=9U'�4�YZa���]qWE�-eKR77��N�	��M�<���ydP/N���h�8F�9p։U��T�΃��&��\�T҂X�u4�xnA"��"~^���W�j�txGU�������m�l�m��sHȂ'������Q/��0I\�������%(o�����̚.�$�F��c��0�S��Dj������O�X��=A��|����a{d�>�SQ_4���]c���gv E�D���z�b/N W�b� �o*M+����ʈ�e���u]���F�j�
� ��m�d;Ð9��%砚�ѿ�@|�Lj��aL��*��c�2Z��:>�6�D�D�Y�T|w�Ј���Bg8�5���ֶ� ��?d�����>|��sߪ���;�,���I�e��X�KE>�/�Kz�ľ���P�� �p�f��hcTE!�2W"۬����O��eo*�]�=Q�o�vȃח/9��y[t�#�7�w,�l&[��u��"@����-
ّ|�&C��V�o��w+��
�s��ӧ���U�y �gSu&���B24�U{�[��K��<p
���e$��/k��6���L}��U"H�c�x� RB=�K&��t��_�Ŋ�ģ֓?~�,�j�K��n�<��ٸ����2ٟ|��&|��:Ѐ^X���+���LR6����t�(>gp��e�a֙��b�J���x��sTb4e!���n�+�+��������:�E6��̜4�4!��{�K�,�I�Mî�Ǻ8���¦;*f�=�����nx	�z��]B�`y��`��e�
��K6~qj�������Q���e����ΘരBQ�MďF,S����ڒ��ܺ)	��y����7Q�-K�jE������gDT��`��X7��l�&H�ϗ~����!�pFWk������4H9Y>�3dx�yk�LӐ�;l�?�$���E؂w�gn��ʹR��bw�&���<��B䬰��	��|�&�8/B�-������˚zDo\ݎc�b� ��B��p�!&i�u�!q��#��D[�I��+�g�XG��+�Ow��[�5���QA�p$���`_Q��v�3`�tRy�<b�#���t�JY\�� ħ�+�v�`��BVe,�!x_�-��(��y�~��W�T���3g�v������VHzG��T%H� 7 I��o����-J�� ����}�q�q[�;V��R�ת�''��؄@4�7!6��A�$��� GL�b���ʎ�T��Yk۔��#�Y�&���T��B8VL�0��7̕���i���C�X�������1(|n0�+/�~tL���H1���J�L�:n��'o9A�s�O�_8�rݫY��J�����pe�Kq�➉4���6���L�Ab5�w���!�f(�/�d^����_˺��������ԃ���UM:4Vq��r�"�U��H	z��q���c_h.��VC�&����1���L���ްJ���#~ƺA����"Z8������V�� �=\D�+���(C��ỏ��<�����Z�֏��b��U��ln���x/�|�f G��O��q�L���3��^V����o�X�Uw�F�*��L�<V$�
ЭQ���<�/��a��y!n�@j[�Ү쭺���{	e�H�S��Xe�AѬp|��j��:��M�-��J\���G��zű��g�}�9Y�^v�_;�>_П�،�m�EӉ���M�dɴDh�oE�UI�u���q�2�mG�`d��Ki�X�_��M�8�A�XR�a���]N�56G�E[G8�Υ�������(+_����wXhND\G|�(�S�_h&j6W)��Xv-A�DE�ݗu�đ�Opϴa���$J��ё)�+�QpB��`�r��XӪ3D\r8QFΓ�Q�����aT���&�=8_u
��B
���wU�jRć�0�:sҚ2 r70�Sn������۴{�����p4����z2�zI���[!
��"�b[����Tp,�:���*�����\�IZ�#�ڔt�6�Y`T��$ά5��LB]�r�R��l�o>�� !��|'K�xPzDb�Zy`�(e`ä�}]z��Dn�������3i�[&�rEA�P�,�������ג���(b!�v�~@���"7��2�C���BL�~�c����v�і9��>������CC��5lBz
���3�b���E���J �:��y�\�E}4LM��i��C��j4^M�g��9]�jR'�����	�THJ�N}�Mz� D|�|j��>[���"Pg|���sѓ�yV"��ء��	��%X)� ��Zz%����ֵ]*3�i�R)'yC)�.�S^iN�Wߝa0����.'`N�l�O��[R��7K,T�F�� k}�w���Nh��y��ba����W���O!���J��%Gȸ]ˡ�l�GI`qR鼛���w�R�-�|�dI�������H[�sՓ�%'��@Q�`�W���"�Z	}Z�����d�:.#��(�v#N<�}�A ���(!�'��HS/��zx0���G�m\���m�A�.�F?�[���A���.��h9gX��֖��da`?Q�"71.f-�΅;��i���O�u�]�DN3C�j �a{	�
�~�24>�Cf�<� k���T}�����U \ ���~�-�����^R��0t�g��H^�Ğ��<���fj��C&�p�#���*r�����:�x�H;��w�,���Q���L��_���竢��ί����ٲ���C�|U6t����;dS%�7p����uwj�8��M�,}�L�oe$�-U8mE'I��Q@%�9Ưkz6468�-��e�^��G�SН��=a�$пZ1���v��ʲ?��I]�Xf��	'X�B>�@pK;!�����w���d/�G�A�E�b��?��~�z`�����\��ȻO���'�#[����@NL0���g�yY�,�!!SԝS�=������<��P'�j8�[5��	��D4t9o�> g�[�'��68� #�OrǺ���ڃ����+<�����w2]^9��@�N�\�<�|��x,d�Ð�H#XY�F�	RHi�*�R%���{F�T����t�$J�������u�� 2��1^����`��3J9����մ�=��R$O5񬋊{ck(5���n�uе*S<�B���Q���8�}*�^��Z(��	6��q4t��GN)���Q3�셄T�����hւ�~G3/}���/K����w%��[zT�͗V��]����r�{���Uw:{P>���>�	�㤕�/g��,X�b�l"FZ��a�?������&"�xk�abJ_�X��nҼ����t��f��`����s����6���D(�	K�Ⓥ.m5�)�̢�,�_̯A���Y��4�D���f]�Ԭ�LawG���Ʀ�EeM-�A\5��n�oH�-�
M�>N�a������	�Ɲj~Ѩ�y��R��$��nЀ�\����錸u�s�)�L˯�����O�E�#j�Xm����Z�_� jN@"�@���V��7��i�t��~2N�n�M-�B�]3�$ڜ�Y��v�>j�t���JSK�n�����;Rt�d�	!�=C��ݽ��9�p������jP��8N��A���Ac�9>r��Zd���^u*��9��kxw��BL%:�纄��Ĉ�k�ա��*(m�ܾim��>��(MD!�P��B��\�>��Wò���-�ۓ�\amS%�r�Ŵ�������l��tw ��Rq"�@C��oq�nX����������>5$`�f��G̹�K��m3y�V;o��$��>�#�2��م�A����+_�`{-H$�+�M�C�'�x.�r8\�[����z��E����!W{3�Li�L�FT��1M`�+��-I�{?���3�7�pߍ�C/��1�J�U���B7i�*��-�߭q��?�q��p�d��p:fP��]��9���4+t��E�b)���	�.�'bR���8>��`ш��U�S:��fh.�h9�!3\� �/ƙj�{������=k�����j8�N�r>.��N$�!�x�Q�ɵ���;&���:�P��u ���/��蜯۹��?lUa=2t�S��;1�R�F] 4/*���r-$��Ǣ_.�m������:E�Gq����D����Aw.T%����C����M�Z�>�u)u������$S�-\�Sc�|q:7)#�N����['�\�~|�����Y+V:0�Ss��2b��>�����"C�l~me��i������I�.�d�������r@;oC�,Jow*b�qQΏ���M�,�����׏[R��w����:I��@�B��'�[����~��e��U$MO�hI�)Q���{:�(��*�(ˆ��� �����K���H�7:ZҮX���FL6E���g[2(��=(`��{��N|��%G�V��E��1���#�Z�`����X�#�=����3|#�c����g:�k�e��=wp�<i9;����v�i&CQR,* |`���F�.��\].ܞA]�b_ޱ+�ȇyO���SY��c��*-�I ���i�g8�o�Dk�͉�����O��$� &���gh '8ù�Y���J�T�8V�aQ\��Q��<�԰"������Y����`�)?R�{A���ZNj�p!�cfTG�m&�8��dl*��>� �/ ��o�?c��y.գ��(�S�=t��Ŏ<����^��!��B�O�x:[O0�v�6���j�8�^{�Y�r����1FCӓѩ�f�>�q�8��P��?큡���$mDwN8*�f��>�E� �N{�P���ӈ�a�K����o�JJ�/s�.g�qx�A��AT�!9��m��R����n�<~�す-����F��,����b��~K{����d����F�TI"��n}K�"�aYz5T�Q�1�g�X���*\�[��0]]
�T��e�f�����"��ꤞ���i��I��od�
1�50��~��A�Մ�޾�n?��;Đ�
��kv��[�U�vR��k��}�<1:v��A�k����[zt29&�d�xr��F1][C�0ɜX��-<d��-�ٔ�~�c�5�Z4g��&|�H�̮=o�Ps�����*�=�&����2[TAWR� dWS��f����3�1o�U�q��_c�6"���:���X� �vA@�^�|�8����ڮ�MX�������S��N��PZ��z��@W��,��	υ��0���l<Y�`	��a(�ӜD�����R*H8[�7�����qypF�a�nz��u,��ԫ�z>�B���C���_)�ߺl`�Ӎ_nhvZ�ߑW؍q��-�@�7V�}3,w��.�����k�Zڕ���?� �6�6�p7���������X�8��1G���|�?n�զy"i;�$A#���a�_>o�ZI�m馾�'��/0g][���\E�������� ����d�����G�R	)��-��~�\C]�|5e���ǆ����t���P����#���aA���;�U[@[[?{,%����@;b��0kАF�|'&ȷؖȫS8�&+X:��x�7�b��$�% �l<��`EM�z2F������Ӽ�&��4��<�F�D�T�C�:����׽��=����Ҏ�<7(�[�3���)���"j���J�z��.+8q1U��s��R]5g��Kˁ�D���O�v�.�<�=����GZ9z�߼��1W���8�ތ� "A��Z��Q�B�:�ާ��ߓǉ|�F�6����A�E�6J�c�<�æ^�OR�U�%wg&�,�=o(�)h��[vj��fN%�ֳ��!٦"�ty>��(�)J��/�=
E=�G<���xh�[���g.G��*�4D�^|��:<k,wɬYu>��S��G+��0�}ܡ?�Aӏ���`׾�^�jK�&ws�����c�|w�l�	�쑏%5N��p��
�/��rM~	�����<0��i��6xE��!�EWFvj���tj&1_e��e�����rgާ�Z�/t�N�k�C3=��#~揱�F�,�o�x�y�as��*Wr��X,!I`~�Ϯ̾�2�l��V�� ���ɕ�L�F��N���g3�N��D�DGu0|�{C�v"fcL�G����%�vz*����NmY����A+�k�<��?9������I�"YahP��E8H;�)�{�hr~�F.��G�mC5`�����vu��QډĬݡbx�J�ڪ�	X��KI��	�Hۃ��[�O��vWN��:o�j��y���G[îk{��)#�f���8�h��`�Nw�u�[�o�
��V����K�1\��12��a�1��ֆ�&s<?�~)����-�aF��A��]�����V�݀,�s���'2}�]�9Q9dȞ}������ӎx|��	u�<��������|msN�U���~�_-��͵+�F�+K�y�I#Q�p��`��İ혒�13?��?���b�?��t�[���JA,�R���/�a�)��+����sY�Җc�.��lqj����FȮ���p%4��Ϋo|�,�K59�h��K��e�������G`�j���>h�LL�;c4�$��e�h�s
z}��:���ǡDS�Zhu�{kI��_�NS��[���s��Q��O-5_�;׳i]��6s�"����k7��ρb^uֻ>���I ��{w�z�rog�P�r[*�&�Ǭ�ڍ�Xn0��b�Ƹ��:���x.��{_�� �����:�����fЙ&��5D}��t�j�N��=6P��μo�I��>��)�t��$�*�^��B�<}h�z]2<�O.�����RUU����"���|� g�� ߂1W����k/@C��p��(�)��61,�4��
k�?�h7���{\$
�n�0�D�`A���������/٣h�@#©P \'Xby�Wβ���ri�J����-䒱2�1�¡� ñĳ!�4V�u�����
��WR�z����������ιhK�wY[q�c�`�
����d(�m��.��FBV�w��]���'�n#�ck�1&j~7Qgt��I�ľ=�d��X凳u�YS6Vxl�`ڠ*B���t��0�!|<i���}Bd-@Ɓu���)�-P�R��k��(��a%��e��!R3P���I	:AEؕ@�����<О<�Ya����h��E�X�� .֥��S�*��V���Ǘ�:��X��pz������X�H���u-`M��V��T�gg(=�t�x^�U��ou�J�)�3�"��b3�"gs��O��t>(�BE����d�5�q��9z��+U\�`q���O���/�l�MN����/��eR2���9�$P�Dz�Äg��D �lq�JBW��3(xf�Rx&�{Sxl4`I��z'��H��
ڔ�چ�#7�D�4��6'n�LD����|("jG ��hfvыc~�fu1X�}::nkDy2q`�d]&XJ�#H�kb�Sҗ���.r����e�ӇѺ:Z���-%�5Do��;�e��d����5�)����{gT\^�㾠8���~���aN�A�z2@��mp��FaH��,L��Y`�=��"������kh=:c1)f�����E˾�X��ǵ_�R)NU�簔��Μ��/5�!�߱C�5le��<��9�v�D�<�W��.�j@2!&%;s���RbH����Z��P�sh�[����6�FA�\f�E�F�{�[gi@�v�������!���u�4,�$�&P��cs�8�vYl�C�ܐp�n���		7.��fA'M��^�v@����*;�;Қn�ζ��a���GF x����i<D�3�k咔��]��*�؂thx���{~�uj��٣��v���&%PVE_=%ql`�s��$ӐA鉛S�G=�t�_�-�%�d��1�/���g`�I���,�w��O�<�=|:��H�%	Т#L�}�(9�,	����$�gM5�G��&�N~Ft���O���3�Ϡ�	ѫq����KkXU��[�2�Z,���� 5}X�j(���?���j�&26�_j���xN-��zv<��P�a�>=7e˓0�&�>�Ȟ�����,���n"/;lթ��4�L���>�<�d�AR��#F����j�1�6�����m��h�xJ���M�8�T�8He���9�%hR.ۮ+���~�M
f�d� n8]�q�d�>��Mi6Az@>�۞R��	/W�ipѷ�~���՘IG��\�Xf�VfՆy5�-����� @��7h@Fۜ4:?U͞�S�"`P@�������}v�a��(��y������x`��0 ����,�������\A�s�L�'<MtE����&0�.Xr!s(�C��j�*�'�h��3���Λ�Ī��1��∑,`o(��˥�P����GpZ[���U
��6���6��]G�-�%�K���58	$`����8��}f��H�����G���`u4�,��nB�,C�G9C��0��:]]�`p���zs���_"goŷ�ڗ@ ��Ujh�=tN�����Q!DAש���d�z�?�`1��*̆m$	;��[��� ����bַ����sX8/a�d#)�3fLg �;0Tm�(���r?[���O���w:��,���q�;<�����H��.y��� ���M�$��}��Y�B�/}(U��ީO �Xd+	�<���oݖ��I&ԏ�����GD7�y�A�	���Xoܸ-W���JeS��`v�5{yʊ��.���p��>Q���fI��Dr2e�e>
����@�}��~�EQ�P��U���F�U��?�b^�|筤�53�2�Q�1�:�c��˴dT49��ezxz�#�q���1Y���+1,�蕝��|u�f^�t|�'�����������u�A&��V�u���ԥ�aV.{�_xv��${�a7���������¯&)&o�ն�[�U�AU\�T�$��\��[}���zPpu_�#�'ï[�s��Wր�5��~,�� �3ET��X&F�֗tvRa�ܓdʨ�hI{�G;��P�Oݏ� ��s���Z�:z��I�U�qͻEWrlasBh����|//rMx��B'Goba�y�����x�ۊÃ��Bh}�c^��g�)1��p��o��R7�SN�*t�sJ!��-,s�@�E�j\"Yi=��;z��o�1f�u��>���A��\���o/�0�\(��ed��'`��K�eBl�:x'W���A�0�̆x�������Q1��DFü_�'���8�_n�u[̌:�7!�u�:6B�*��A"X#�\9�^v6���X����V�Mu��\:�${��> 7�հ�]�Ō��h�m?�}nߴ�#J0�Ƥ���^��Zơ��!�*�,���!�驽��Ӡa��¹��O Y��o8`�������~x���L���94��������]���*C�X����~ٛ�Q=����R��Z����oau�l�@bT�1
�	#	��{y���,�.��N�g�^M`����_;��wvѝ'�k�toxqp*雜�p����%�I�����Ou a��I��JSÐ��1h-��^4�S�����6.F��
b���$6�n;֥��ɩ��� �R��l�D��X��h>�c��OX���.O9+�s�K+�3f��̇����|m�Mืa{:��d�Ǟ�����V�aw�#h�N���r	{�}#�cW�Z�Gjw�~����z���;|���sNM�}�=ǘ(�H�����^ߥ����24���%c��s��̈�`�KQՃ�n*�Ϳ��t�֌��t<���t�bWv���5@@�w]�'����Zۨ�$
��VQZP�D��M��6����E?� 0}U��Ľ	`C]�-�S�ӻGM��[�	����m�������#����A̹҄�����v��V��_��#+�GƂ>��f�>�#���Jr�������F��c8�r-r�:g���͓����Kusl�K���sXleD�@�����5%�:R��ڄqפ����~���l�#�NƧ�7�c^��=O�ޫ�_�t��*Mu{������=ޕ�H��s�X���6���<N���@��%��<M���Q��d�sV|/��%��2-�I�^eE�8�e�.�x�iG�j��{G3��}��|Hٌ�`fJ���b]��'���`����ð&�������l�l%��XL�ƅ�;�m��]��^�ę%^��qhla�"m�~ngw�[�S� նZ4�&��v0�c3!�Ȝ��'�Rf+GT"(���F�YN�x��y�Z1Z���OeP�$V�s��8/M()��Ԡ�>y][E҅�IF���T�mt��t�	:ft)=��s��P�;�"Lq��U���"�(�)p�����e�0A�;?�A��9PD���P�ح�w�3=�ԓt{�4o�|0�[�y8#7c	Tk'�	�bނ�tQ���	4ć|���x�C9��f5"�S�L	�ȕ�	Sz�ԙc���E���~�s�������)չx̴[|~���+Tv¹����	��l���'+�m~�*Bw��� �����Sſ7�V�0��S��;���8�S��b5����>��ë�Ry!|=��tH����P�ڔ.C�"�����`���S�7@T䦉g}m\ 4~;�x%H�k>u�8H�Kc-�0�b�hOЎ���s��x�u��r{��af^z��{6tz���н�9n�z��\�_�2�b�I�8�$ R�0zR��J{KB��6��Y�=�`vi,������<�a�����x
Է2ʓ�ѩx9D<Ѯ0��& z;r��o���]�e+���c?�A���*��b��\9O��L�.h��K% ���ҳ�؟o�= S؂
͠��?^9~�5U QT��[d
�I�r��-�2#� �VWR
 �97EV���F^�m�gR�IL~��x�Q��DgQge5iB�Yf�V62fx�SH���n��[�m�	S�-/l�G��a�V��%�@�kǙ�=AS�5?b���E�����<�'�O�7"��:<�$d/m��)�uBw�X4�v�?7	��	�詄{_�OP�~
�a�@����ӧK^����$�|TO���%
�	��^b��	e��{��'��M% 7u�#Jf� ��l���'��w���!�Ә�	��6l���>ν��
�eW���=���_��"Sl�8⧔�%D��D9�/��6�%6�v�%4s&�4��Җ�/-t!9󯖪��RD�څ�CW�z��Դ�X5�F響����#�
!3�j;E-�F�8V�}Aan����������9�K��8c�n�f������$������ԝ�h520����Ԕ7V�fr+i+(L�94!J���Ӌ�F7�d�hR���r�
�!������.Z��iI9��E�P�ǈ���܎fr�v�J�������3|�j^t&��]�f�i��A$%����r]���(�����6w��e3^Q�+7r�G�#	�������ks�3_�Y���޻s�	�ۉ\FPC���Z��;�Q�"������>�Xτd��1��ײe@m/�U�\����z\� 7`u|�9�.��;:�7�<֗�Rc��_SQ�����q�X?�y*�iua����8 ��ʯ��ȊCٕX���8V.��JE;���"V2�'�4M��W�c]�;7�K�UhL�y�q#����f�����E����~g_=��� 2�N��\N�^�H��͠%�p�5��S�@ss3jR9�����^�8>$��*d{(le��V��	�x"c�2}a��%���J�C�:e׃�7g<ӧh�����?�[�hǏ��>z!::�P](���KR ��ze��"7��x~}��XkX� ̋���Y
̎{�����l6����-w[T@�t��Yf��M�1��y��Q����P�SY�C&�ْ��Σ� �Hy���
���8n�5(,��X�A�nv�
�ׅ-�K{{�E{LM�\�ψ�p�����P=铼{�v,�*� ���78&�.��j�h:�!`�(�ýw�����u|%���H+xucK�6{�V7���_�[���mE
���逼�czx�pT����n2bq����܈�xk~��Hn$*a��������_=Ef)l��ZOk���W~E�qt��K">����02˵a�;Z��_Ksמּm���%��'��²U�Iaʪu��F�t�$j���f�*��I�ܼ�J�siB2mH�}^���ǹh��/�Wy)���&��L�i&(�l�ʄܰ�A���䚀`����P���H�z~UI�H��
������@���'"����������d��+l��횩[v{9�Ha#Y.��T�$����n.����E��2�n��=�vϜ�=*gK��m�BϹ�	�i�1��[v�U(��9����y�C��7�`�a��:�'�Qd�ؘzĹ�X{�M�Mf��ltL��T'Fٺ���^���P�
Y�P��οqA�#搈�̶ ��4d���B��,h��ϒ�רd���t��tG��޽����ǲY!KoFs�>��q�&X��r*�c8=�p�Q������klӊO�z�4��������&8-��t�ʊ�5�k>�vq�5�[�%"��ܠy߈�f�\������$�� !һ2�,wޗY����ZH���(EO�nBI��|b�P�iLa�4�5g���A�-��Im�j�-@�7��41F��Jݵ�f�.P���)�ʃB�� ����=,\�.Xq��w�3��3	��7�-Ԓ�?M"�#�9���������}^n�S��>Ft�,$�Ax��d"�bQ���^M�������-��$�U�A���O�o��\�������5�f��uǎ�M��<����o�{���p�:�X��jZ ƘZo�Ҹ,2N��8F�k�Q=���d�������t.|S!`�xZ�s��{��/���3�%o�J��Ft��4ҭ-�z����m��^:�|��`�vr����{$����1�(��~>���
�cR�7��j�/8��ry�j���;�[�ђnI4�f���E��W�Uc�*�7�~4�y-lMw�>���ghͨ5���>��q-�ǅ(|Ԡ\���&�R%{��m�(�`�^�\Xʾ*���ʿ�9Q�����E���t6t`��2�5��j���D��5�8���u��{x�^T3ֹ�kΊp��u�W<z�����1 }�^���ޙA#v�Y���1K���'�0�lm�a�ú�
��E6ې/?�R�'`�#�	�����	X��B@�!n�&^����HK�S�ʳ����5c��GY�}ej�ǯ Ȝߌ���7P��D?+}&R�a�)������й�nب0n
��d[&@�k��ȉ�v=���q�@V#"��&�͂*����.� ��n�S�&n_�=z�Ӳd����j�h��gA����4��o�Q�M�>;������v�w�OU�=/p�^�eطo�l��%�#aLxsqьB�� �P��n\��Aq�Te;�D��,`�֍{�yi�'ښN������G�����R��uE�81o���>Q��0�w��h���Ƕt���h�f����"�Ԏ�&*�;:lZ+�g�yߦ`!A]l�41�O�HR���[�j@���jd��� ~����4tH�?����N2�U��(*��aW�uf�-6���Y�7���]�4H;9��f�1�&餖�V���WOѩ�q�)�� ���W٥�
sO�U����؁���K���,ް�4��R^V��a��5��|2S�tW��uϞ~�>Tc���.���=�H�j�(:�3Ah�N�c�p���]	��� V���Z�?Fu 3�x�Ǔ\<���,M�(�v2���Q�e�80���ktJ̷�~R��K9�~�V}gfA!�Y�3�؀���Yq��1=z^�ۯ���������\i6��gED�L�S{G�&qrwxEb��v�N]z�!4=!%��.�\1-L�C1�o��+1�<��c�g��r>�&4������ �Y�f�F�Ko�`����c�� ���b##ɮ9>2����bo�%*-�TZ�	����2O����k~�o�&����B(��Y��dmb�rC��3�2�����
ъ;�6��b��O�%�g���g2���!r�ן�`ȅH�y�b�������y|�~y�����f���C&���3pSxn���ۂ���b��K�?ښֳ�oѓ��`rwGn�:(�6���OH-�/��x��Ԍ����P�ۖBE��T�p�f�#�Y�S�en��g�ͽ+�J*%o���U�M��	����{��,�f�dha��/?�@�Y˵���;�DkEh�rw�;T�`�k��s��4ځ�R@��~O�]8���*xz��x��Dnd�B4��5%<�W��՛猴�U�a��Z;b�a�i?�ٴ��ڱSF{*{�r�c������#3�?n}�_r�I�_<R�܅n[
�H�h��<>{Ue%F�$:�^YN#-Im-�5�r��[�Ex��uup����`n
�� ����֜��9�.�H	F{ 4�(���q��ts@Z?�;J�J�s�Q~}��}��������L�s�h?,�_��h=���B�N>��&�̇֙�.����$�$�L4��*��@���~��(	�T$@�	���Ϫ�KP��8)6��M���/��H
�	!1@n҃�� �E�^4�W�-+���0_"%�� q�b� ����Bμ��$�7����u)i��42BC�:��͇�敬9����Q�BӍT��Qᒢ���<Gk��������y��H�gĉ�2�|<�5:�V���e����dP�ﲮ�NiD�`h�nbd�Nm$�w�'�1w��0�^F�D�٢�c��� @�� Ԛ�
�vX�!�9����a��Oy.�K���!^#w��{�h4S�bskCH�s��096����
MU +=�!��0(i�(?X�cJz����"�Wo�"��t��5��+�]�]���4#��R'P|����5�?��ᵺD�*[������C	�4��B)Ȭ؛�br�$�^2��]"vF����}�ͬ�����"�׷wE��T��
�}��E��2�rV�	шب[i�H��%G��o�|=knk�������׹n�rIm_=uL0K{�U�1T������Z&�������Q���(Dھ]�}���W�d�x�(}��Q߄�ˁ
v�5�_�����Ln�e_$Rƌ���
'v�HB�^����]N����!p��*b��Y����ybrKHB.���kR|q�iYF3¥�f���~������1��k*	��ԓ7�e��?�8�/�r���K��\^-��Î�ON�f>q�:�\+	<�4i}H�Uc��{78��܀BaQG������G�hk�zo��&'�fY2�TK���
�KpʪV�䏨N��~����gk��ⲈW;
�S��;����Ρm���<w�lW3'm+��=J
�9�cǦ�CD�5���*��YD���pl>�!�X�ο7P����֤�8כ�V�WE������u����.���ЀkN��D"1��;�)0q-�>/{!��Z_A~�������4V�����,��U���P�(�CJ\����C�9yM�~��'�m~��W�R�x�ӍB�n:��U�dh�=��&y}.1Z&V�f*�+�f��l������kP�@|��rC�ߢ�H^�so�+�)�t����Qᕔ�3��_MN�U���'QG�kTy���<t�2Q-��X���3�6 �/y��ï	ݠ?�����b�ԁ3�UQQQ���	K�#�l&X��^�m� ���-�;�r�}el��Cc�j����:����~�I�dd�P��knT,��G�]�̉Iz�:>|��IБ�w�g2[j�c�~pP�4.�Dg#>�[�)��p�d���|�|A-�=���Xyk�Wv5+��M�ab��t�vv�z���(�n�@����_*k�/G�\�J��Q/�P�TG_����U>𶢵�(�;J������6�n؜�)F�%��l�p�iLz�aU�с�F�n�Pۑ1m�u�5����{�m"?L���1��}e��r�)L LkɞH&���׵pcT�y���ۖ�u1G� �Ew����M��JC�jЙ��<,<���ea!l����F�
�r�Z����P��?��D~rV�a�0T����t��vQ|���+
��V5u
د�1�ɉf4-��<C�:
=�r[FA�"�IJ1��9��3��"��b�$����i��5��Nb���N�x�Xh����;x�aA�N.@����5)
nV�!��p��F[hz���P��h�4�e��#���Z�xѰ�oGA��'Y1�A����"	D���Ɯ;X���vr�^�&VVǝ��g�d�Ԏ?����Eu�2p���-���-I[�3-�&/B3�����ɳ�jW��d����\-�_�k��u1Q !�A�=ri��h>
�X�s۵Je���b����Ic�$�d����H����r�Z}�ݔKs�m-&�[%_.\-(�>�+�����u2�2�h��_�	�.��(�/���5l)����M��o>�����R��J\]�sr��
xeڛ�x�)�9A~.oM���O���D~w@t�:�d� �Aɹa���B����n�S53����� ͻ�.�y�=��ƣ\)w���2O�<}��o���4 �j��S�*S3�*=�Gg���n �H�0�KA�Kѥ���-i�UԚ�D�Ƚ�r�U*7Ah࿽�����V��6B�l|��ʱʍ�R�I(��7d���Y=t��|1t}�6� �J�,pJD�9�0���y�H8B�{���"LT���T������+$f �|�Gqؑ��&��4@�Gٙ�f�^��� �Q�L���<��&X��񗆸����7 &5۩1�$4��l�d*>��6�Pk(S��vd�c�		�g�*bW���saS3�*˗�0��ʶ4�&n�NC]n�Q�â�
�$.`z����k���\����07'��ǣ�)L��l V��gW��ߞ�$�F|���ߵ��nhP�+`�!�:�C_�a酌/-ws���f��l����^l�;̘����]�;�1��?\���"Ƒ�Ê#��yj���Y�s)�3L�*L�Ckz������w�*]Ɵ�b�� Q�	�A#�?�Y[�i��蜒"�sd��Q��ۑ�(�k�ѭXr5�֥�g^�b���n'<��F�{��P[e
�⿜iSt׋��語�-jq9��j߅3Ƣ4[����"+���u��;���B�ҙR�*q��2 �_2�Qb�@ۀQ:�&��sBq(�:E�ռ���WWπ��M$�.����v����$O�I��i��`��#�#Dُ�uI�c_��T�]1Ƿ�Zu�8wF�Ʉ�w�Ȍ���	��(\�O����k�"���=�$��vP��Y�ҵ|a*dI����Pq�.����<��X�At����,"�c�T���WllI�#�L��:i����`��i��<��6u�s�/�X��H�C^�w�����Hd��ALE�k*�eQ#�uP��@|�H�9 [�ӣ׻�;�8�In��Ʋz��8�)m���cA�H��9���Μ5�i{�����34����PI�_�9�Y���$�sZ��e���en	���Oc�)PJ�^�����b�c*��4���k�<t�9�N��$}9̅u~��u���(��2Ss{oO�'�Z huA�UY��
� �J�IS��W�&��I�U�^O}���F][��_�A�^X��W��=%E����ǰP��c��²�$\]�sv]�%Qf�N�� :Ol��YD��|�O^��`���Q��!��eY������"���52���l��p	P:kSтA*p���n��e��Mد9pW8q���P�Xn��ږs����}v��g�@��M�]"~��qYη�o��N�����I���4�e��R��V�� f�\W��Q��3�����N�f�A$UBG�Ya�s�Z�b>���C�
Ž��3�a9���V'�q���5oma3<�4s,ƚ"��&�C��kO:W��C�Ih��iXx���1�
�y�rL��~���8�I[���4d��2P��!����{A|���$���&�
�ˬp���D��~��j�HR飐c���27W�b��o�4�#��i��	J���oO�v҅x)�{���P�Xı��l�=2��@�
�y�y�_�_1\$�cɛ��}�DB����Z��?�l�TI�m*hZӏ!����U��E��f�l܎<O��"\8-Y!��W��'&��ZZ�ܤ��:�ZX�T��PL��3��i�U�����"��,���2T��Z�	/�0��%W���V���5��i����)~���.b&��xEL8�rLbgh!8��49'�.��f��ѼN~��!W|<㻉ۿ6��H1�!��Smb��G���Zq("i6%d�����ze�b=	�@R���^�r�Ls2Hb��| >����&��o(7�I�Q���O�'=�+9��y�xz�=�<���D���?Z��������;}��_����IY�B�wΚ��Sj�� *Ƀx#~&0Rf��8�fcjE{F��Yݻ���d���ܕFQmH�1D���#A[��|��ה���J�{�T�ò�Cq��
V�g�F![��	w���m�f�R�W��a(v�_��J���|n� #�)��=1�8lǼ"�y�H|U���ui:�9`{�����W�߬�83��!�K�y~W���,��Aިe�U���\�;(fh���9F��K(�
�>:AQGR�n��� ���f ��!�iM�>�T5��F6##��D֌>Ԓj�?�%E�b��ظ[6������f�b����6��R	�m�3��������=�]%��M���b;Wb����H�	�������"�����mN@�Z ��2էe�&��޸�(y�J;��n7�k�I���sS�^ֻV���k��rk��\hWԘ<�����pF;cx�?����G��G��"%\-�& ���՜í�r�#Pu��(I��h*i��V�1e�C���q��P혂h��0u:�
;��e�G�I{���ҟB0�W�+���|�(LW!!5g��������J�$�אe(����k(��© C�x�@�3����)��s%=u���t��2��#;s�\H�Kf��l�c�@�����W�P��8A��OL��L�hzǓ�!ɀ*ĸ�怓L )K�^m�s�}�I�.�+��SeڗMH�<S�R��,Z��&&EU_H�FO�N�:�OGa� }ry5�v�D�W��#;#���䳫A���l�@�K������'�W65|#՜OCe�!�^�i�]�.�Nߌ,܇�u�^��9�7��b�?)��Ļ��~_Q0T
6�5r���Պ�a��l�S�SQ	�F�kR�+��ݡy�H��^�Z��3ޚ������������ۖgg�';��g�j�G}'�\}O;ZB�yԤ�Ť	�6n,���{ /���u0�)Ko�k��x��&p�u�Ŵ�M��(&?��ڽ��E8$�r\���yG�E*o� o�B����ݩUѩ&T����۽���Y��QGg%�������"�����MH�I���o���hZ�;�≍�H����`� �yeE�؁���Ĝ7��}d��D�&��p�/fY}T���zF�I��6�ȖiQJ�%��Yʍ��ņ.���"��q6�,�����	�� /��N}x �Rz��2�L��"�J���5& ���e>�.��yʠ�#���)�`���~�O�v�g_�V����*ߖ���qe�l��_�HS�̗1����X�N)7g��>(��l�q׀��x�Ԉ��6[������z"���^L�F�Һ���G���
���2O���X���q��Z���9� ��h[S�L�(��@L�؞g��M�����C|�� �k|��IY�1��e�ũ�B0��J�]���h�Ub���A���|�<I1s3��U<~/�,�Tؾ��F�m�?v�m=aJf�m�0�s�b�(��ծ-����9u�f���"Hތ?��=��) ���qN�����~�W�t�	�P�� �PQ��~��Z���^ߍZ�kf"���e��
��~h�et�~M�� xu�"�QKi�W+��1�:�=��c\@+�vg{_� /���k�5b�GK����}���Xb�~�9���Gң�X�}�}���ɡ��~t��h�l6*ʄ�G�b>�~� T�c��)`�y{�mE6��٘�X��G�:�$~�&w!k�7 g�ix�V�p1�85\�!�����W�1�N�I�}�3��w���,�	`�a�5E5vuk���:M��q�h�=ֈ�?h5�9u#ǏD L��������Ho̧?�[����e��x��:#�ń~���F��">/�/��e%�� �D�#Qi�A����H��8���h���fH�3��fgJcV�P2$nL0���͊�Z�Yî9P�����F�P8I��2/���h���%���%�p�V�Y�{�T:�s�Q�P�#�`�[���\d��j{�� q�2f��J���6���٘�&�:���| "�qr���k����/H��5�L��T�8�.�1��t�~ʪ$2Ƃ��hh�x� R���R�A;cSt�}��`\���P����vU!_ذͶu���9M3�x�s�!B�J�;��pd�[�Aq��H���q�:R�
H�v���?pZF���L�j��(o LK���tF�5ڦ�.�����a{���M�K��	c��KW[��3�Ǻ/���>�BD�O�����~W��49�k��g���i����
b�p���et��F�B�0�"�O\���7z%�"sru�gAcv��6W)T "���W�؃��; @�p�Y��R�r��1^~��a�m�NF���5s%����RngP��.	A�����rDԢ�Pߎ���X`����GC�$���>�}�o���� ���β��W�y5P"��V�7˔4�g(I�s["�@�xr���!����Ks$a�ܭY��E�Gs���{<�yg�ƅ::;��@������Ӂ�(5)]�q����%*�}n4�� �Nk�B��@[��/����*5J@p���+�i�3�ͫ��馞/Y�Ge�A�G+�I���2��]%sf���9�_1*�A�:XX`�@�2/ڠl�6�~�����PT���# �2�%��I�S��Q@��a������H$�ץmo���˭����$��� E�U�~ؼ4���u��V�r��J�# =`m�	�z-�ݒ�3�C��NU):!�2�o����-T���B?ō,�5��T΄�V�t�-��=4v�7C&�S���.�N��# ��YԘi�jML�a(�T�u���{���Nljv�n-V��u�/a�e�k�b��]�xnE�pߑDi9HS@�}Ƥݠ����u� H�紽��g��Ϳ�aC���t]-�Hg��A��=uԃ��+��=�Ҁ/����Zn�t���唡��w��8�����TR��dت`T�dU���
Љ1hP�8uPm���z+�g�Z�/��<&vq��&��_���7��L:��g�_ۮ�!�K�j�n�,�o���M�o=5���I~?���P�a6�Z�E�.��#�[���k�g�fX�xe��kk�����e�gK�xo�K���N(�:X���?�-�M��x�nUcs��:����q(ݐ���_0��fn�=ݪ��6�^��%d{�"��==2J�en���5��䂞ʲh�a�z�^��0�; g�!:����p�44��3i��Y�b|���g�T��ֆ��'��4��>s�,^����Gfm�q(:S^��D��&)n2P�Gk�bAы̐�{T���%�t;���/*���*=�s:��{�5��2��AN��qj�ㄺ�Vʡ�ai3MvpN�K��{o���oŰ|Gh6�l�M�*︠��+���"��O����v�ш%^�k� pO�!;�N;@'��xT$���:�Se<�Z�:���j{f��fZ��S��@��6;�8���P�_�����Tfܡn��Zy"_�ȫ�g���ѿՎ|�>@� B�Gѵ":�A��oh���^㌒`'$?��AXN_��x A;T���Eȸ�$��i��:���)}��Y]�pH@;Z��Cb��MWioŲ �۞1]�l��`
�ujr�J����y0T�7n~��:�y3�*|��J7��քU�%#}D.��G��L3H��b��#:���I�#�NIT�,B����A����!�/Nf���f#}˳_�}T�o�l�D�)~|\���N,�?�u�����Eސ��g����-u��_Xb\����TuR�x��o�/s�alDE�w�~SXX�K��^�ve �,�ኽ;�y4�^�c%�8��&��Q��áV�ϫ2~bߡR���Lt�oiӳ��@�b��_8��S�b��ظi&&�E6@���j�E�x����@姅ُsx~��v�����c���-m��n�`�0���ʮ�b��͞��}��O��H�wŹuR�y�Չ��n'��&(4�GC��%1��G8�Q��+�4/	�s-u��_��ތ�pR�����!��_�<\	u?��.��e�T%���Eµ���Ҭ>��d1s����P��q��NS�`ʤw��u�͋f7�򾾡����g�,҆Jh��%pޜz�÷5���ɗu/T�hZ�]%
^(�fBծW:p�	�	���Wv�
�q��]��j������bP�����=J<��H��'F#�򿉘#�0*r�ҧ]{�m�9��'�@�4׽���$�Hp�	��Q�� +�x$N��2��yU]��I�4�:w�D������KTh�]+g$>}��D�`�=tw�5'�H��?S�zd=~J���喳�K.%�6�	Jg������4�V��s�1�%�H]��8h�ŞJ��(_[(M�{F�r6��A
��D2�M�.����v\lg}�aӕ�qkd��fM��ϖ|��;���RL��$�u���L����;��HD��ǲv��9����XW�tN;;>W��zEf���Ϟ�Z�v��=Å)���T?��K=�㿎�|�O����ݳ��R�X�=1Q��#k@�>�5yQ1L�J}���c��Ls���-��+{�j��}g8��J,W�]�2
Yh�E?�q����^7������W��g_'�2F^Nly�U�5/��A|��ǁ��TJj+�[�\�d׋�O�{�vA�=�4Ϩ�b(Ip�b9�~�Mc�l�wъ���l;�oN4$��y8W#2�6��*��s��R	t�C�(�.,�L�(�R!�D�cr����!"���&��*|ˣg�fyd��3�����o��b���T�_Z����F�Rv(~ކ�V!0RB�_�� ���� ��wv�ɳ��^MN�Rv],�ݱ�����h�?���<ƛ`�4y��u=��Px��Τ
M�ڻ�[�d��/� �'~�����|����<�I�@���������ǅ���rA��x�+�:�4	lڝ�H`��M����(�N��8��'���4��Ұp����SA�A$���/����U�ѠfX1Fd!���8������{#�Y"�Y���ޅ[����LC��ύ���l�k#B�''q�K\����>:�FH9=���j"�u��M|K��ZBZh����y/;'��ݔN�3z���☛+��Kj	F�$�Q�8�q��v�Њ��_>���-Ə���;,��L��3�����xY�m��Cg"�k��"�4�!��V����'�ϵ�T�'�s�hI>�T��V������WR7�5��{���&T����D��J{���!��U�P�cR��?-�m��E	��r� �\[�*�"��ܣ8b�s�>S�[�<�༄��M�ٹ	j���$��� ���x�q��nH#Z� �����[�]g��H�5��t/�W��EY�u��ݴ�,7�wӣ���MZ2PC@E�±O�ε�e7ԎP%���tA�^�G��U�6�5��k�|��B����J`e��2eC��Q���#�BYz[CFԔ�՗��Q;9�Í�$�31�[�i�E�7e�XpU�8w��t���d�p�����A.�[�z���JD�qŽ���J�^|��q�$�E�s���D�dZ�������I�P�v�x����.z9b���P��~�oRK����ݾ�=�9v�:�c��אt6ʩ�4�!Ɬ;�>�̔�O`A�O	!��
X�8z^�����p�x��H����8#P՝�jZp7�#�k ��_��Ǭ���O�-�ڮ��<m�u<Hzd�&��'�%���o�ە�u���j8]�?H�	\= �u0���~�տ���r���@j�E��a�@��p�m�I5I,v�qG�����!����x_�۰�H裼a�UM��1��f%�N�T5�Sb��ԏ�|�;�'��?�6	���>���g}�� �c^}��^J]�+���S3a2��{
7j�vp#�@E)����4zq���^G�|���bz����L��۲���7����#����9s�uS�2�"�d�Ng�L�(���O��Z�V%���В��[U@@�Mh��)W�kЙ2��ƌX:	't�βT��t2����si���QD�e:�~�c?c�#���=\��<t�2��	Jki� AX+\�F �/��A�5�B�2�쯑�j�0�����n�/�g�i��*}�1�{�{�s2�\Ѽu���Y�ѭ�j�hSF�t*���8�C�|�h4���b�o��z��|"�?���Hs��6Y��)<������	U���V�����g��尠&��NO�ԣ�"WX�J�x�ȑ~����/��:�G�!�T1�l2����Is��F~�o_�F�Ƽ�?�
h_qLC������|��P$��M'Xt�Mg�JȬV��K�̡�B�3�ޣJda��X.�gƵn��lw%��>�Xs V�ޚo�b�'h��ڣ�س�4��碁	�(���ȭ(�r�U/s�=����0?�0N�$ �<co��2��ܲ���Q�4�X�`��}6΁�Rn%P����0��&��y��]ΰ(�B�2ibPw��c�M�t�n��s�@���Y���y��u��u��kH_���]�(��;Bc�U��@�E�Y����$s�_M���Δ�����k�>$5L^��+�,�rw�e$���iUC��G5m	�vu�?S�N%���@�1�]!RP��OE�0�����<�ݺ��gU���o��:�Ń�Si�&ܛ�ң?�L�ˊ@���րo;�Z��=-�ɝ�p;�1�@��Yp�&��}��"5iZ��J����0������V����%�|'��aY3�I���'q��}7qu��s��,��m�l8���N�f����Q�0Q̥�9�F�Q!O��i�X	�RO�����-�n�E�%92�F���{ڱҤ���a�C�"��P�"DY�����̦�~��kpX(�Z˥*��\6��	�T��g�S��E;��@��Z�3�ڢ,-_�xOL�W�t.ih�qu���Kᨌ��R.R�5�5k�\I�UˉA����A�3�;���=�O�ɏ�U8�2�g�WτZh��_�1�hYW��v&��L`��<���r�'�P�w�Se��.�t��\c[t��%�m�8T�?�]2�,|i�dB�d�`B��[]���)�
�,�Xls��= OX�����^\�orɚ��ɡ���#V
�X��ҙ�D�K�scq=<��n<������}{#���W�&k[:�lR|���Sx�o�`/�I�!>e��|���e�%�:1�E��=I~���9M��e&6��s�UE�9#�c�e�,���?d�kӎ�c���82zVEcU_k��׉Ϧ�%�-��z&�BB���,ެ?��b+��Y�@����y���������h���1}��4vR>��Jx�l��zˌњͳ�t�Ԝ��N���#W��?;��I��AQD'�(c���V]�1��ǅ|��[�A&���X��O�ƃS��9@��ɺϣ])��XW��}4J�d+ev���.Qu�U�vD�ڰ�v@���I6 	v��;[� ����p*��0�q�ʯ�)���"΂�P� �E�^淫�8�"��� �����˝�J�!�;["=����窺�m�Hr��mPDK@<��P��_X[��?�X�je�u�n�eL�%���������|9x�.�^�埼-�U�Z��lkw(�^�R`^|�	_��ᾐ�O4W[���R𿫱b������J�e���kҸ5�"��`�#��1�i^2������L6�3�c���1C�?�V��yT�	E����x�Wظ �a��E�!LB2�eI��I��+*�����'&�tJΎ�Z�d�?�z3���ǋ�`l��Ҵ@�ۦ��' �{X�z+<�Rl��A�� R-�F�%�����T��mα_w]u�~�֖�ďۘU�L�92�����u�ˠQ�Y�ex
�dPR�W_RD���ߦ�d�pb�=6x���fK����%�y��řD\K૲�hCQ�t�����w�`zC�����1��ZR�e�'3�ÍB�BH��"2_�SO+�ߖjI�Ա�=D(b��%%�¨���QX
��������Wc$�}	�6��q��V�R�.;��S�ϨrYo�պjH���)@���eOo�s���iԑ�5��~"�*��T}�ӆ����;�`�@�@B��S�s��_�����>��\)'��>�f����(u�D0�V}���KQ��fo����*�bda�x���`S�j�����ÿP�]L7պ��-
�*K������w���.�����1�ƛ�(sA&�6���xZ�@�G��^J�#C��c�Zg���U�`?=L����Y�ONQ�@ǸP�JY%�~����ҥ�T�y���
�-Yj�2B ��ՌN��>%57v����>��c��>�UBjx�;2��f�1K�KV[h�H��+ v|��84N�r��ewU��H�S�S���#g��8$r�˃� �˲B'��ZB�ݎ	�x�t��^�:h|1/sp4�w\�XU���P�<Bo�l\:7����?��m52tX�!�k��kY^��l�����rд�	�qS��O#�dv��֥��m��_��_�=2�wd��Rr�K���[���Ȗ�nX��k��Y�Xh�E����`de���(��;��&rL9���p�y����v����5<��S!;�j4����x�u�YY�w���*_L�3�4X/&��f�7<*���+B�����P0#*���3#A�^�޽�;&RA���}}2��e��0�'������,��v}z�2���4%���A�]�kBag>w�uJ8���i�D��`vv�T��=d���)7xU��Bo�T�&8�~��M�m#����'s�MɁ�^r5��<�8C��S�����~i���>T�^�h,ˀ�w�o[�l�}N�'�mUj�J
	���61{����Q��U�Y0J/;�tn��7n�X�f%��-%b�-ԓ����vZ]��$'���R�}0(pe��tF�K�%�t�-������Eh)& 6�V�3�;�Y)"����)����B�#XH�	I�KN����/DV��"N�u|�v�&F m�ql��ռ@��G4FP<^�CZ~�����8�DW	XY�F�/�����t1�n�&�oR����TX�kV�h,z�V�#�*������7�F���a�ɽ��P)�����G%w�W����;�����Vo���Y�˦��<���	'�܅` ���m��mBl�ǉH������GR�5f@���pfM�uY�.�Ɇ�s�7��|�`��Ҵ�_��h~�}G�iZC7�����&ߗ_�.3��)g��!�:?�+�I{3����I���x@D{RC�� �5T�[�@1���})N'{4��jj�5�3�1��bɩ��Vk洝�NV�s���+���eO,���˛���Xb�[��µ��I�UVV�_I5ƞ����O;���oS��� ���F���mBˢ�V͊D���#7z�-�fؠ��1&�G\�pOxc���9��y���j���"Ұr�����S�ɚ=��mJh�t���<��ۗ�����<7�wp�a��{y��v����ǾZ��Q*���X��*q:���go&����%��}q.=)�N3�����n�p/�iE �Z.�k���+u�<� }$�\4�]\\����a���T^:(4/@�V�ǋC�>�k{J�K�[�s)r�)�z`�d������Y^v����&�Ђ&g8l �����S���[[̼���Zb��q�g��29��9 �E���g��J���Ү,e���@�nU�u��9,��b����vr�+�oڷk
�����(SP�Ӄ�V�i�H��}>C��\xՄ];-^�2�����bɈR��|���%�mx���*�������(�?�v>&ٳe��=L�}�'��u7��j����y��.�Nn��!\���	���v萈� xAծ�.`�=R���<����Q�%'���>y��@�ɈW�L�d��� �;	: q��'@dd��t8�&�崯Z���wS�Ҡ�J����#x���o�o�c���eO��(�D��G��W��1[��,#N���;�[�ll��&�*�1�:c�8�ͣJ��0����*=�|����3�?K�Eu��uH��!�R��ԋ�Rwnn���y�B�,�W�,y ��T�˪��$r��Vb� o,pheE��Ձ��JT�쐋�$�I�\�]x�'�ϵ��@� h+�N��O�w���y��FZ��`[A��D%i�ֹ�<J��K�{wK+x����,����J7�|�j�l~)K/H��D08>=br��O���;Ku����eX���.Ad�eS��cڍ&Jd5;����帕�O3���3�b����ߓ��x0]s��3�,�f�6�?H줉��:�L`����J]r_����,#�-P��2������c����W�O6��Ʈ�&q@��A�K�`�@�k�HĔZ��.uü0���qlhPpgn�PÆ��F�_g���P�U6�z�v��G���JI��b����:�A_h=#�)��΅�H 67K�V�u}xh@b�R�f���`���o<	;d�QX<�I�f�������~oAʿ�.OW���e��[�6��� ��=�w�9��IN7Z(�a�����o�""�7���+X�I�B��p�'/�1�:w�� �dŜˉ�U��찎EIt �a�,������9���!V4�"jҽDK�@9Gnd�14�Q�kW�)�I
�c�jb��t���罸vc(Ekl>n;gV:#eI��ˠ�:i�OqPy�̃��Ȥ�a!*@�sηT*7Yc����GE��f���	��۝�O�]�{�?<��ܴ�����U��x�N #q{���ق���V�����!kAkk�����	Ϫ����L�q���y��{+!|�n�fo)x�������|W)��7F�x_�����/��(h\�?#:w�p��y��į��N�6g�1�y=�����;RZ���ɔF���jpQ��e4FmilZ�/+48���VE�L�٨=��D[ `���+j"*gq񪼤a�ЧON��\������&�����;5�C:A���t�<nDe�~���g��>�܏��:Q�u�+,��fv��Pv�W����2��y;��:8����;(׍�+Հ��\'ɒ~ ����S��LW��у��}��Ǒ�z�ޅ2۴���6�~�TR	3�C�	��,��w���w}��K6��?��6�@��'��^{=����N{�b��7�7��SdV?�R���0���x|���w{$Q�lg���1>�ݤq ��oxO	��ӎB(-�r�E_f�&{:aE�\�'o��Eύ��nޕ�]k�N���1R{C���7S�cV�iF~XOa@�<a=Y�Z�*T�����ݛ�M���!=ٶ���?Sɕ��h.R_j�'Q��N,����6`]S�+}��z�>�m��=����-qqb��r�� �Щ֖'Ełn��p��S�+4���]8��w� U�P������* 5`��J�K��������U�����/��yǋ�'qV�sm�W��f1��^�b�$�i�]\&��=��=�������K�'	�~�����l?K��+v*f��s �`X�� �0�NhB>|֓h��-�_ω -�d<b�b�]�t�3S�F�6�|_��53��Hx	���4�W��oHre@��N���
�}�g�K�W�q�,���|�q2l;5��F�hӪ��L����͖�"9�g�6��MH�-�͟�����?Y�����&��^E��~�����#� �&���ܟ֧��c���1��p��
7?dj����p	~7���;���{�������T)�r�t�g��cy>ey�p�o��W�P�ܼ0֒��%��ٯi�b��׽��Ŋ�S���o �K�I�J����<���Hqق��%I�-H):�_FU�>V�����%`�-�m-�A��i���Ef��V������6�(�7����C"�Vl=�x��GxK?]�0��pb&�H���to��bi�<�A��'���X� }��M��:j�������F�����`�{P	ʻr�^�Y(r��mY�)!��پ��&���;���G)^ �������S�������t4SVD���cMHMkf�[/K��_�B�2Qʝ=ۧ'�`���p�:
�DH�G�j�>�w�F1�?Ĩ�d
Յi��y�$��J$�(�!�$�� [����Fi/��a�+�;�W�K� )+���{m�U�����F4��Z�}�Л� �h����%�y��V�D�^���~ĳ��r�t{7�������%E��]@�1
�}\Y,����*��{� +���L��XW7�S�N�P��+���1�3$�-�#�z2%d�Jp�M彔6��t��r �+?���^ԐFm��8V��G�����G� ;c�,��a�5����t#w	�&�.E�+"�t��TgԄ�H ��e W�5����� �.nux�3�۸I�b��I�T�ى�;�p-�A��/Ȓ�.��%^2��N��9P��X*��i��4���rˤM�]���g]+<+)<�����O�𰴲�zN����)�:��T��äN��&4X��f�����\KalT�烪N�L�Q�0~ņ�i��:�%|����PM����%����/}TG���e._ �ٛS[�g�T��m���b�7"�Z>�����۶�0�U���\�|@���C��:�̽ۋj5��ch(펻Vr�B~����vEbm�;g���r���ڳ��0�+A�b�e���L�5i�`ΧY�:[��܂�g�Imi߾����~e�^�L�����Rn�7`��4�{�툫��(xk�"�1+j��K[�cBn�[ha��x�m:xЈu:�9{��KK��(59�ݚr`'���G�
Cx��&���[�D)�����|�c��:pt1����ފ;3�c�S��;�(99fv��JhHx��3Ր^��hd�(8@����S��~"F1�=]�*��v])�X�|a'�Yp�([z)V9��b<\Pso[�x��9�E�6N�L�NU�r��ބ���%t(w,��Z��N�2_Z�']X.c������r�j��m8 ��?u�y����%�������/�,ꇽx޷���co$��UNK���A�%�)�7�fL��g���L�0��m}a�2�MB:|4y�x4#��ՌD}�#?�0��ߵ��-�ǉO��^5d�]Ho��^�rT��ߵ�0q8`U�r���۩�DHu�E�9��xѝnH�~�����ҙ��ɴy=��J�E��+�?#�k{ U9g�m2��!W[(�-l�:k�'�y7b7P�˗�k_�A�.�j1|QZ�nF�Cs��I��؆_�^�TS�������R��״�p�P���[X������0�$����&ҬaM�mZx?
(ݷX��7�H���L��/9�D~}�d�'W�C��.أv����-5�q�xgy[�9����Ց��ʻнׄv�6ʜ.o�XMBa}A�yur$<]���J�h#�3>���ߧ�J�gBx%w��N��� ��Y��c-Fi].i�K�H�O�e�T���V�o�0�jW�r�b�v⧛~JIR���,�ɟUE�	*�/DAST^�.�G�r!��"	y��ե�v�E'�-�������n�9팵廞�e%�Qd6�%���v-1��f��<.�!K�Y�{�s>��=aI+k��y���Icv�N-�E����+��a����G
w����y��;2�u	�D`3‭3t�ꄿ�*^Yߋ�}�v�7��b,��T���7��W��t}��[��
��3�{��k �&��^dG�3�՜:�d=gϐ����o��q����znD���[�Ɯ.1� ���JE�:�7���خ�7��7R���_��j�-��T��@��+�s��l��j⺚���7�����d�Փ��4�(hJ���3pm���5�;��z\�p�g��و�=W�zE�F�D�G�ȁ�j��A��#�cg�넯Nc���U�-1����V���ްy��	!E^&�Q�����%=_iэ]D�9�`a����>���g�Nο�:�w��e�^�+����>�\!Z�f�U���I�%?��_�nBԊ�O�D�����������F�V2eU���$����f��ۘX�kZڤ��7V���Rhx�Q��d�1�9�]>^�^�Ņ����0ݖi�;	��;|�2q�)a�AƵ2@���Տ�]8��*������������h�/^�1���A+��~J׮F��V"rq�fػ�2-s���+ձ����� �@r��4I[eM������Lim�k�J�p�~ɿ-�f�Q�b��k\��|ǩ��Q�6�(�%o��7��h+��|����/Ǩ,��}�]Pڳ�zgA�Jh����法a�=��Xߠ���H}�E�6��6Y��dρ�DBc�����5Z@��	N�����W�|n���+< ��J��y#�v���oK�x18(�Z�o���zz�x�?�"��gO�r�
��׏�E��b&t�YX�h�����]gw>��
u�=����p�$#��"yKC�8�G�	�5"��p�
+L�;ၧZ����@