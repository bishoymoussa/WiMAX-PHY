-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
x0PhW56nh9U9xqas+FpBmSjLqA3F/kr6h5W76PMQD5flELntTQ9cKEYuxJSt9BgV70w5cGXz8gmm
PuJwmBKrPQrb+feSmOQllKsiiqJN1t8Fb51EEHWacXQmWwK+6ctgzLv+EaUXYqU9cqoE2SZQ82NX
P/OiwI9bo2D0yIrrW7Lms/WD4PNfZnsPAFny8UsgCpJEJ1nprVWmiXr3dtKhq4r+Ux1geIxZarNk
2QYwIYayHdpIEM1/JwZr+msl/z2xdZd0cJyeQ6YWnlFXgFpt2Y/UpYWXa/MR4M43v5RGPly6na0a
m9dmr3L/L0YS9MK1efJCY7hUBgQJktFqFUVR3A==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 7712)
`protect data_block
fdaVhcBw/rCs9k1BMylgbMaygHS9GOXCrd7NiDrFPJyqzRnw7zjawJIu7df51RhSDi7CcAPFPGjk
wzF7hfG8emBJNyVy8c4IqLIXHtmeLuPGEEYChMy0mKnzxJPByS9XdR7Rwim7FqhId+ByzIPlH38+
uDEi7FpWz/JP6cCvxpo2bqhvKsrfe+jL9mXWp2V5FePvXyEjSqxSXsqbM0qNLzoxRIsAo0BETlRp
ZJO+1c6sXLX0550zyvUwT8uJDWlYegWudJRFpi2x7ZQB7qQcsBVynssP8JZsmvKXk2a9Mb1nZmJF
m07nh+AZVWdWhlOh7OTlkX7MIMB/pEiUV8Ck8PVU36rZJg9dF9TzC7tTeJd5PLEKmGOUXRStFZHa
Yqq0WZGLLj6118cMnbSZmeIW1Q2+tjrAApxIPa7aj8rnrrFbp/XkmZRVg83TJkYMVpDutncpFL3J
Rb1/QpYgCS93UyyjMEYVyFTw7v8A7Ie2UH/90FlDuh6rRTjysBQRBRAqZs3U6OwDemjW/czu9erc
KJ7oa5k2+5eTuTQSl4yAi3jWo2Y9Rt88zaql0Xg1jPr/Pa14OZBHQM1PwOkqh2hfX5R4NOk46K6N
7qv8kWtx3PDUJO01YaAhgEg8QAnb9cSqhhSnTpFwJGMqxcVg0dTQTqFGgT5a2SGmF+6V+lIainQU
UHc7g2ekLUpnX4iCs+V24U/bsTUSdB8UmelX+lpnIAMRtw0csAl/vWBhriwVz6SH9+W0HpBifOaH
xbqjL2Wi88ZAd1Qvcb6fKQYI0X+fGSTCfod/Md31wY1P+Ar81UGP4ZDL8H3RCMj3qdi6oAEixhfL
+vd7c4577cAJqcpq64Qps2NadQNZQsDZ0Keafhv9Ig28J++nHRKBV8TR8il8wzK7JSwxzm0N96kD
FOIpccbj6lzXTgOgi5F2ZMQOLeDRQsXwaQtd9G1zrVO7DGJ7n98ZzUSnEtaDhclQE+xU9pd6m7cb
nHJpKYk15z5NATaesm7nViq6yPiJrUPbRJ+pOlwK2uoHFzcVpBa5X1jY0nS9Dn/NVSTK0Q7xob4k
2mmiggkEnfhnbilLHBoeW++3cPO/lxMKq7ZxOJcdDpogWwEMcrGWwuH+RlijV24zsyAFjrldbx4J
1UqLm2IcM0fvCHVC013bFY9aVzLNuCSx7ysaDKRlRlNJWTbtpze3HVlgH3C02/owe5kl3Ac644n1
tDCdoyRxGaQD2gLhtipwHgWVUmgt/IDrjsuyEMyjxjN79dcsBZ3u+QkYg/y3ar0pxKZz299ePbTc
Ih7EJAb7M/56TnjmMUK0gcTQfHqj+EWgizktn1t5qyRXAgVRZk7LRExCcY840BkE9rJSfSqiLjKB
0SzLv7/Ap9gIMpO1yCn1entgmag6MaWAr1eipLzEOSMxmRn/3avHM8oJ9VZRYc2D/rYX4zIuCdcr
jACNDnkwwng/CE6soEKPlD5XEVVpuOQuIi9k2h8K9SUaSwyVMa79ijSPljzrj6Qpslti6TrvPlY6
AT61SdW9GLIXJvmQ97Or0DMZTYcBCZ/EGp61fLQkMUSQ/rxyK74IASSXt1ffLqK3zHAhxVbMu6Sg
eQzffQ4eaTL+Vj6JxZoocDxXgNsSbdslXJ9sNzr4wAAuPXp9VJcA5JlhhWMewtcVnCeSGmFUnOX0
cCoMbb6myoTB00u+IJTsIrK7Hn6bAfSxNX/Hpf3L+obl1NYqFLFCrDS5m/+IodWGJwfBBQxIq3e2
UyJoCv8JZf1FWTVhkYEidF1AgEYXjrJj7MazSa/SrrkQGHElOp6Wm4S/dJSmTFNGGF0nlp409wjP
W5c77H5YmoIAT9ejbjcf8oAhA+tNKSvs3cj4mMkhvWdC+e+woEIgB+dxcn8wO+4PWQptbhv3qoW9
d+X774hdtd+qCBKXFHlhkxN938q4TH0btR5cL+h6wWkP6FAwrZxEuiZAr9E87ptqRdRsgzf27YjV
oQkrYnxiAHOaKSuIUadwcOwkvCYFuzZ/8KR38/QglYaBvr89FBJIO88CMU16sNRadUBjerXwH7y/
4BDbRVDbMQmWQHJ+kQTPE2tjXTzAso3fbVN5SHyzlhAzNgtGrHBeR8k4gwFR49uyf2G97Cdobk9s
oQDS1fWgyTbRE9ELRFeiuc/l225rcEeG5dSuOkY3Jj4Uls4yKFPmWkl/VKTKRcqytZA9rNVrkbrq
I6ZFcXkn+/0VvtpehdLPQYSODUiQD4o7NJaRtYvizwxi/Hlu1SyhnyL4FH8L7eM6qFiHvZ6fjBXu
8czBVvZ13RTpzkpFPEf4GVSmfWuo2QVHVPONu8ClVTuIBzZelAwV5NrFoT/00yDJhon26ZSdATij
hCe65IGnPGsOWAiiC2zl3FEk9+yYcN6424jfkkbByA9pBF2xMs4JJAHR+Uyp5kKpkp8AvrM4pGLv
RD+LanK1GxD7pHbUavFaWEPOCVuJnGm4XKz/MnQp0TfbNNA0Q8iX6UtG3wBdd7uelr3bpBqjbBng
/tkHThPPCXTWHzA/t/f2/HhsuIQ5q7zHeRdHqtxuswewtINcqfuEXXrMxKDkzjs75X4ggQMTWtbQ
ki256pnvBM24UMBUJQYO7HrfeqGNmUQctY6qB9yyD3eRPHiMQVF4pw+BJtnkIvflM1Stuo+FmiS5
8m235Y0qdV2+ZYg+iUPV3H6TLTCRBwQqlYS9FxW+AYs4tTEV415XWRQ85N5I4lplYDmldgDjcMbR
hPEDbKo0S2zFATXAJoPqj4Wwv8W8u+m+UdW6FqwOPEaYvTlqZykhTd1mZwu8LRNUUk2370fcJm3t
hI7ujAqTZpZiGOMGSzv9irjJSxpWnl6FMGMBkkupqiAgqchIYHTZOFkkkoXuNlxKhmykUCDnhVbH
/ksjjxW9bfRVPg5qtIwiuZVgZm9HWvQ37WDgicQnomQZZCTEck3dQceajEHyu4ljl5eai9+XIgFV
mYuX2yQveUDOYIcWtdK9T+kUcDwPdl67YBOHaF2gbTzjl3bJKJO7IL+VCLTRvSSPwXPa8TzJLBK7
MW+DKU3CQ0KsgI0iDPXBJ5ceE2iyimyLQuJkbvISj2IhCpIA21EKpit0HNc3LzbU6uwcRUNcbPbI
nhJoNWw9Ecj6rBhFbssPbJRaKTvFszO26dHxIahwrPv6/E2a1apUslYHhC5jCB1ueCKli2SEE+eX
U3vFVZDUBsqpfEj2feCitDe6jQ9ekja3gOmwPm5lGRLHFlehK7ll05Ai9/qRhD++94GgnOekTDY+
Z1WOoukyEnVOldpHtUK/Pl6s0zoDjW1a7kQnkfesZLluoaO3JTZqE5/twp4cCmHiA1HOlrWTj7Nf
SRtNdJERh4zwDD486mpRwbpCGXtpXmcseRnHNdWPnU8Lt0KhL0olYPD5qtCR9Ow2QcVRDYCiRlYy
buZZ+wmDVr3xDQSyVXHoP6Cpphn94dx7hgFXBfJ4MIwBSDVXTxno58bemjNIzp/Yrp/KaqnZUtye
11AjMSZA5J8AiiPQ8fDScj/sUAf7KXYMYYEhdduFkR6J/8kRF3KnZFoRdlb59wV7ny6z6lsBjte6
Treu/GbVQ3nR4+uAE/pb2fznJno4gQFV6TejH9DkVz/W4EfYLigre/KJZsztMk0EUa/9Fl8aYVFJ
RO5VEFQuv+7+S1eewWHZxN90uVpdsCzu01DWSEbc7Sg5+Gx0+JUYxveVf/YSz3OjVFCMYk/uc45Q
xschqLPRm2QUD5mc9+KIOGEgPHi6jqfjzj93QFjveygJ/iuhe1qVKNpEkxz5kQB6U1HI5l+JTSLh
yCO5W2/OlMc5CX+QukF7h4aaLoJ7CYI0pzl//eGm5YdBoRopXJNielkVWCVBM57inRqzR9GxgL+s
DSTRHOBFWIULMCcmm+21d2FHrAnGd2VcAbbcCdHIugeT/mrsEEHc6z+p2efx4ziVV479Jd/yV6sr
gdxpYokK/Q8Oldhw4QFE3hLIFskIRXsiMdOkiqA+K1H0ftjIpotf/JwRqq/xJ1tFX/EbSoasWl7k
G+MoIVGPlKDsK+jdgbT+jgO9oqJEKPFjxcuc2+B85LkODBd/EKNBN72c+eNTWs5YV2du65KOD2IV
3II63Te83OBgRv4rTWHBx//32VQ/mze2OwPYXvxjCbAoQi3/ummETpBZs4GbfisDkjac89mvrtee
bScxccrVmvku5qIAqDnNa97iRtdUQI+VS7ziJFwXQL8ypYWujy4/xGGlXm0qonZl0NOtEjgx6uFr
rQN3CHIlqWnJfDtEiIlJpYZzoXvY4CmkSlXoK3axdsCUvM5LDRR9ZWcV0QwcnVpjzOcQcglCyE/P
aOyt5JR2mIFUEIA4Pmp/hsbL8m+v5h5CzhO+gRYERIO5cXW46HQThwi0ij0bLyT6XJg7BuZfLLiy
2ect1dtd1LMdXmN017zjeZoa8revm5eCwW5rxV1lf98PxpX+totGCqmJRs3cCOR/YnWNxsVdSVie
ceZ1BTF71rJd1OO25MIh6j1LcJIv8jb+YrmX566FkrRWqh+BOy5OvvBEQADPnpUEvh76CN2xwMVb
QYhZ1pxXNeclfEYFUeMUWNaLapMtQYKAbOhtaVSzIlfNYodYPluQUW9XrmkBrbEPO4B0lHKtmUJy
hyP//MHnA5e+b7l80MKRlaLJCcrGusgKHwKFOxB5PH6xU5juYEIeELXFxGYzxrHmyijqmyZFiRVw
o8CJP/2ZFQTZwKKe7+WGv55CZ0OT4/zXC0xd7PDbiTUNezh9ug46aQmeg7ZadM/z/n3L4Y2Ylfm2
Ht+77MdMWGI/asTymjuWgLpW/WUPuVRgMM80jEHESzH6Lc9VhPKOxmkZWa4spfoF5f6Kli4s4Tc8
ER3x/WPLpQHZNy8vibQ89vtQywKz/bvKEH3wPlIo6NpwFxCz7/ECgxXWguWfQOyXzihA39tUlL5p
omNDrYoMIL8xjrXyUGPY9IWAiwv2xpeh5zxQDaM8/OGGOAP4wcc79z59MJrcwYeTlMspVI9MdKhs
zJ4Fn5sH3pv5ZMDnJYfXYZXYXLntpBtNgdLp3qpFwgBmYYG4FlNCsO1/WWf/TQSHbLwUHA5w2l24
NnJZVSn7S0G6IQUsaxydCGqr09bUtefMVNTGliZSrhptlGcijBGTJ9bULHBBkldmJW5PlmWeTIbV
x/47rtZvxPIDn9tfOzK+BX2DdpDhVFIAbmQnyaLTWhjYF4wIsbZ+qANzjoUkpIWujSbFo+m47/Xa
a+29qUCNRKwNXc+R+DP1sY8BcxL2VD3XHDKggGqlw75fLB23O66qJ/Qw7ko/nb8oaaapwjqL5Lqx
DBKvuwYpIBbwKOE+fllAq4xoKj8lDLWA0IX/1Sk9oLln4NjBorert5q8fdxR3FFicZi1Cz3TAR/a
wjRhIGA9m01mFjBgl42HxwJUWSVqcMPuXZNuo4xs525QS/CDnHsdWVkvbGKGeBly/sQIGHZCWZPo
WcIl6oAD8p6XJKBjb+Cpm8NcED1KC8JG9an4u9mYKF9/OiczM/dDO1wlmOK7o8kyiE4JulLFPLr+
kpaWpE8UXxWTGCW8GA55M3ST1YDXMWNZmv+kbFphC9IybMR0Hx4qqTPNnGwHRBgzfXOewW36h0tj
uFtUwi0lhVBsLzscSlia+Wgt2hLP77zdsXMcYJPjiTGkxWxOWkKY5+p7eheQcJaPg3h9FUfREKuj
9UNYYWG1xqVdsUaw7oEYKo2YjYfZm3shdMUfG1scjIUcoMULWaIReEP3OpgtI9DD/o7lGt6JtZZ4
I4+6BZ6Ce/ZzW5vtywbxyHzfyiOH+K/rluXfBcrMT05JAIKMKlb54QflP7rUESeC6isn1UP4uMTK
lV26Sys65vTonP6Z4elDkOLzCUkiY4StyrCRA8R0jqP55dlsXJO5hWtTe4fjGbdbYSjvZaxcMEM/
+wsGzdr02GnLMZfvDCdkZ862L5bSNG/Jd6BPC2Vus6HT4nD1oKOqoz+zTJ498CwHSaP1a0/LAG/L
JUu9Bkp4QFqDYP0bCLu9d0SxGIApKgqaCES3nFdT519HDeEn9pkpdld4d7gESGr8uMLNEt8Qxp1b
LadGpIgehUJ1yGXrBR973Kymd4aPKalM99ISGNK9qgiaE+IQ5FxWkO30HWxeKspQyGG/pntatmQS
uywBvovuLLN4mhDtU5/fw9IqGlEDCUwOr5ht5lXR+6Oal8GlG5Ql07joKDULKdDz/hOgQHg756o/
bPKJdoSSvhi4/4WKc3Mg0rZtpLY1fg6PlpLMALGcPWOitMh/zSdfiZwd9TL6Hfp8PmQQa1QiCkeJ
tAAJY7A9QDd6GHD2lVlcDhWoqCSnlxbKywTjItD5R1OM83tZStNc8U8lPohxKFqAUljjDBqwFZWM
o/nLEt9Cfv0AUMFQGs3WFI2ApJbHBmh8rkq2ajtJr9Pxd1/SBmXXETI6rTWTqxs1fQFgC+1x5rAt
htQ2FC2oF3adeSyfVc7YvWWwTDb3DK/s4Wc60Y6BkGHuB20Cyvw1AtI4Tyu/oteeCSxi2xDw8zAZ
qPf+pJPKa0i41uWca36jmrNjulIuJOZaMwYROAgUuSHLs9bxDs/94RAP1VAGPTp8OGkDaVVWhkSD
5YTm3ZK4ZvYTjm/9LqLlPUIojPcHGByMqHsI696FqLMf1LLD1t5JrsN53iuofIs8Ro7TOEBoQD+s
D9jgNu2dMOp5je+O3BXKENXvLtCIkPuTYtyVeEvdlYm/udiBLvluz8h9YQup0e30TZQy018/EjsT
EAHK1wsBUdW5nenC5oUZWgMVEDp3O4TH3EFxK1dcm7RQAtjeSDbicPSNi78R2oJ0XCXWztXSs00I
GDgyuOIirPK3BQKo6fKjOX1ta18l5488WxnGqdeR+ds4pLNcr+9csfyDNOxRQmN1aBfvG58LP4Oa
+hZhta8ztmTcVXLoh7aBxI1TbDZCgGXwqeG1DrbPkTbuPIzwj5f5s0rllKfPRI2SJyaoPGsGOcrZ
RxjO6ge6Ah/Ks0EfLEQM48LrzAkMxxrgl7g1MCLCi8qAHu9lT7BbGcBldPFsAUMfVeIjk76DKcUx
J3HAyNaE3IQzg1+yLM+pnOe/IEdY8T2vQjyCHLDAXeyFXBomD8u18lJLhqT8FYXZynELSm7FJPCb
z7XGMdx1O6c+akyvRqLcG3ZIRLAUFMEQ3pY/djEQlD3N0NsE5nSIUEAvwKz4nxulRHnqOdyrhojm
0pBCxTCMWJhuv8ssxuWqGS5v0MEI6J/FHj4v5VvU++4vp+5KPDpPeOYV82tTNYZQfHz8GOvbjBrm
0h7RDpN0i9FchIroipshrvqYy2FGRxvzigpS3mxwZTLNY7+Q/T9/N4yJ008u4Ij7FWT0icO4xVV9
IUydtjXsIE0hY3JLgA6l7UsyFFf1lZqkundP4BlSKsisoDLEshPrnm7RRXJNvSOsa/FW8hbm2MP4
lwjeZPP16+gO1STWrarjxs26Zkax4gnj2eLGyh513/FyYBRSVkNR/+c8A3IZSrxX2kxF4eKmFqdG
qjibynrxpQP23ZWwmseRgH2nxm4LexrO6ixXfki3XSWIYOWN/5P81xTL03DvQXxvDYFbj9YYyitt
kVKI/js05MN7isdhz64ligX63egKy6ZRe4wx8sYhPBs/RD20zobXL3MqM0IfaZ303bE2nyl1fwY6
nKliXlB4kwMAdKBaNjYxCJARdeOhTLscCby/jhzHOLmL1qryJWYxZyP1e9SnkTOy7kemJ1DTnlce
jAs6pe0FrQcDYR/uSh3hVTzCcuSvlD8eH0p9i6+SJ4CzoSqA+uZ0iZe6nrSTQntenVFBS/n2U9xa
cF/vn/ql220+OPRlLjAHIiuPX7ZU6IhsCmJAFmwfXm4rc1p1My++8U/BbYuYo7SSXkjlQOtC5q5y
o7K2phbvb27exTMtLLxWSTM/c4sZt6jM0xh0pZR/NqosbWRlGvIfL7FYDwJSHMkSOLUBNbC/Dbdp
GND00UcLwzuXy/UVfrLmJ/L0WWqYWIzw6xbi3zw7Rc4sV6xVnV3WnVovAUUiz8eQ+cQcyrUBeI74
Hx4KYlHX0DoSQfTuCkxImuCrMUeM8YrXsdXAoIdzyA6tTQDLu4gUPvhEwSkPyeLKhcc0h0zUiLxp
3vUUbUPjr84liNSlR2ZrrT2+Adw2HXwEwog1y6M1woMrvuBKWZPXFpYagCc1QCclJfmBuIzKutS4
pFLrdKUDg7PcSTC3eC8zfR6VtE2fNE0ax49ahvhlm6XF2GlHXdS73+hMrpXQs7EBMGoyJ2GJgS8n
xEzhwDaMvRARQc1qcocnwdBEgvNVIdHoAC/gp4a/fu97ha8JNQpkEaKi+ud+qRqzNb/2VC6paY5n
2F4gkEBJNEuNHN12dcX0cheFOGtTLGDLmm1LwK+LrFG4n1R2T3g9cmbAUG5twhjTtjEzwOSmHLhz
ceULIvgfr2ZNlN2NSTM0OsvMI6i5/vT0Nt4NNnFSESC/+XkCMFOBH/hixtIkIRIrwkKC00HM54sV
3DLDkE8n8y1e4Jtt0nLG4JFDSnCrQFjDEzVQd/D+j8cuPlHLbgs5wzirHEQlIuNUhf9oVK2q/n1M
O4yI9hAunoFq2kqeJprmQxJsWaOpBsg4dO9u7lawWFxleaK9uIuuOvgPsktck1S0rdGAme4wrTjC
c/rXe78P2ahtJExJGIggYYeXXpQ8TDo+9J+dMAZoAl0ddgTi60JS3uBrAnhmrmdjUuotLhK+3MvS
czMq3iIhs2tnObQSqnEPYez+dJnriKGi0x6FD605n8Z0iAqZf/OT44sesUKCeYVuv8Dx0vSfS6xL
nuyTSVUHOS3k57MAf04o58tGoBYyhtGtzwnTzVT87WIhKSXgaml/eAUbdD4IGFe9ZnBjX1Mr2ztS
Gb9+1lQpTxH8Hr1CimnPyRMocEyXwOyjTQENlZGZ1oQLNkoEQX0iWUvwFwPXBiK04DMkr/U+GzpP
alBs1h5iMK31TsR8GNIrQhOx2EmlIFkUbA84jBjeNJLl2frcCfxQhIJg9BpfMKwqMT5kzEzjpZDz
kMAVyPVCKw0E3XwSJKHHlZCQITOCol/Oc4gmalYpJ/h+RS2MkZabrIDh9mrevRJcqOBPGghkXUZn
9Lese3OGdRS4ly1nCrIuv6OY9vcWcpurGs0JhfUtWV1V3Khj4yuGIPIy9jbHqIFS9vJi8UbWwOgu
p4+FN1uUL7QKHEZBrU4v5FFg4+Mpr5N17Rt3fbnlwlozrvabh/QU7+j77SIA+XrCeXL7hWdNoHqB
jUHZdCLvB/ZlaG7nd9e6rBb2HBWqV12uEWOIpsHJVgCIj78KtmxzRS1pQEQqq9jZoS/EFtLE4R4C
tBaov5+k1q5f4KCiqjjhis26PN5A94j3ktcOHmRwqhJcC3XfRTHJnrobTy6DwzhqD66cJRXcEKMP
CSbQlqjH7L0uLKkDFPNqgXI7QwiCrNPz+M3ZdKiDugDWX/bxbmnQA5UYhr4zh0CiBwIpnRIWx/w0
qmQHJQ+QxJ3smY6b6qsgODH7B5WVitlqDqQ+pq+JM/fcTukuaVAKgOr8I29cMAiFzrRlhRXTvc9/
jYI8wocTeeorWc8z+tBaCnQqdMVGSG0atc8jIM4kZ4vmIOPhx2ZC85UUfO35bCoBZUkpG2sswGVy
WELGEgel0McJMX8xKEY8q5WSSXHoaoSugOvfCTeb/gxyQra4YpbjhbRp+l2O1am8tTSDfPpEZbC2
SF59o2uqbDiKvA67ISGZM2lj0OHwrw4axwQ9U3wuprJpWr9NAonUM/3mdz53+kdvtmmepM9ymxUn
dcKeoWA7jeFUNSTiUVklc+YCh4zDt8QC0DE9K9G1FpQm0+7wOxj5wf2WEb4nFWfrDGdZHeYSntar
Txj5ZnvDXQ2FbE00OSsVM7ry5udrF3KZNx2UwwXExMcKxXXrw73mawMHJQ5NMlf5QHdK6FJO8plK
E5uqHVdcAKSJuv5tlvmIWT34ADrVVPSWzT3MtrrIiGpzMUeCmMvAhBMZ+BlePwaqt5+odlZnKRef
Tmj24o75G+B8s0CdQCjipNHSUQqHSme3aF+r8jDFtf8ajUSYRzZ0dZlFiJWXKvWyMaXPy3BQOAir
r7tI6pgUl0mi2anVQ+x0kL6j/N8UqD99x6bJ4nm737O1LS1EAjKGh6Wnb9qOk5SOSadRsO0olBpN
8O0eGFcNvadoEHVd/ZuCzyapZy5zVCKAlpqAxFuloc82MZZUL6/nz12H25TSXCotcxtpWAImYLvN
LyK/k+tZgqfg3l3adstLOS8=
`protect end_protected
