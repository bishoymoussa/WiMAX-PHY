-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
wWMhjqe0/2FtVDjX7wSsnx+11qpnkcCHNF5h9yEok3OMJFQtFqXB0HS+EIPIWfz5MxcuSelbjdsH
5oCXK7PoJ0foBm4+8HRGTjUDceB/gnUV2DH1BecitJa+vTHAXLmtNL30F2LxC8ESMwgKhp2PH767
PW8gvPpgNrRR6u0eHZAWMHNqLvf46W0wWLJYjukTEOP17YjeRrvLQT0IhB9gCnWeLFAeofubCh5O
GBAW0InZTly204MzjhQg1KP8axjt21IOaKeHNsT5wzXM40+k1likQ2FcAXFKOFe9Q4mjZyD6vV3o
f6d0hjOXYOAgs0VfR3e2t0BqdyRxPI5Jw7FNQA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 30096)
`protect data_block
GMC8jUBZTBNCnKg1q9MjdSYVJXq1kXrH0SDZUB3zncjz0f9RQhuaXgVFGqtmiHIQIL+C5rtrPHXC
zxz8ksJfOw5Lpt6UtQmfLfaOpuO4HoXp2eTQO7IF4prwzxhnF0Ew4pEmSSUNZFycuPmvLV9sjiMa
ih26TTtHcdi+wi0dj7INaSSdE1AQLyxyIa8+jvMDjH+eEkMH3JqR8YkrBTJuZduefvUd1TG00NIa
Xyn06xV81PolsZgFfkFFgKy+33oOHT7DugQ528a7rCqcT54Rpg91dOMsc93JXtFVaVSYhMoB77rP
9ZwsN9yjl6t3yQ1tFSmbVipWnB8FoixChqF9WKn4mfI0BZhxO+i6PisyOq4BfjVfbtyv0Yvp3krv
zwzY+mhy5JQbnrHaqxKc87uP/4qrWRZgGYocZsv2kiGO1/N5r/M2DkUSKDpA7ie7mW3NZKFht6fM
TSM3HDwUxtGSXT+q/2fjdoO7NbVhIfFjlNwZ/foqnVhYOqZ19WrQyqQwtLz7JvEOIv37mRRHCFv5
YTqicVpv2qW2ouY36piCFwqJqSLUBkWwQcvAECJALst5+23m/hXpyrTlhmFltpsH8Ku7FiBAyOic
Vy/uHqApclhdjAz/1COxdk5adgLGhPZAxrOAtzCAxOYR+1mrjPyz8XYY1XK+uncbYhAWbGIQcOFK
4bZU+61wvTZzYeUC39sh4Rwqaa3TTZfdw8rrfXVC1nYhmkTpAbViu07OcEDAkBr4VzAG/Ygb4ajs
uG2ZtVZcKa2kvXFiy0n39i3cQ8GAUl1I1roP0ug9YITMS0Y1mj4xbO6rroLnraDInol1A4k2Fopf
xvYS25todgHBvItfGUUjUD1VRqoTtzk502vwhchaleM1p7TkW4VAX2SagOAULlP/P3akXKzdzZwH
pzUp1/CGqhteFSNH1CO6XebuEjsSddwGyITEOVW4tqXL3ByfhlayOg52CtEG0d+SCISppvcSy9+f
8gQ+AKm3uL+BHzls6lcB7AemrrIHoXG5wGMYSJJ4em/lk+D17CzAZXjnxkrpQ/u8xoABzZXsSJ49
CuSpVqOo0voqejTr4vnKSmKOXnz990U7wp2p3d+zZ881/VePKkcWSCwUnioO5LCmsfWt7KdcPfij
ZL8y6KfbXNLE/cq9vFwbhiERyKt5IU7f6lZCu1eL/KopRjYAZZjmIsi9AR3V2RIeC/Zf9ivzTaDJ
KO5Nxba+fTkITy/BB1CEe+BPWfMgGjpsUFHUj2cO/VqWqbySA1SOvktHcQ8I0Z1hS+AgFFxY9jas
qRGL15ooME8O10Qpt9p5SBSBO8v5x2FDYT8hl+9UKzLHxize71FeIpytGHJWAyfnWIOzzoCEmRmp
SIjuFhTCEcdwS/0VJaqovULZNQzrJ+bTiUZRj3U6B5ZSRIAIRrKD4SDGcgc+qTI9l3TqQLHO0+6n
/tj0YXaQUbtFTzk0zdjf91efymODYcMKGmTDfj3euOsGrz4rzt0jfIxrHlsDxjGwVf/TjqIg1MPI
MOMTaqUC0q/XJRq5hm8ie7gvjcZoTRaJZlXGxJvpTG+tSZkMDy9ugCVZK5PpH++kUyUzdtdGZgg7
aBHR3KB7JiKHagSPAAuqu/CTXN5Uf9sZmyF5DY9RdjqhBV1VSO9pURrsvwFEjfOXfF0P9YPVzye3
L9/UBEXvKAAjgkRw30AhJb81hURFfNE/yhtKlAU4g06URbKkPpmarXliGfTx7dO1nYtZyw7rFMOu
g0Mbmgyt5kC35oV5NTPRshCqDtpGXx/aOlHEFp3CkbBf/wSF3/VWWJ/u8I+4xvK5SQQ80MbtgZoD
YQMDd0sPazr00B+QrbxL4YvIa7yTJ5pgP9aMWotUVsvvY2V7cUP62WCHWS7M6RaHfsj39b4ni/w4
Q9aIuiohi0forSHoZTCZmXugQ9ct5rKFsSqI7GtAvoxXX0Hh63Ui9ZwUpow1TBhy/5Fe9FJ1Sh+v
MK+chrfNidmvFszI6xLYnkMnoAE7u+2kW756PLEuZ5b9nFvUkliYn+uj2DvSTWLSZoKYKxJAiXh9
c5lgpkh3gEVIMyNEx7/lnltwY6Qlx8Al57KvQd1P/yrJ2iCgVX94zoraJXL81HcQjpIDeN3In0Oo
uxq07nRpgQcpqcJmzEFAmZUgJbDmPlzpZrDWh8TaCduxJWGU5rmEVosaHuNoESLwRHT2LyxQVsrC
bq2UcX6oz16Oh55Z7/zBUFBat1QTlmULKzVKEncy1EqEaA+dzpQVijjxiGIUuMcIUgCbv1Ldw6R5
cPlzMntLE+siPuvh2yP65jl5o92ru5EF+LsAPDZDLDRmscGDJgeQcTUNkq/dtKkElWDr3P3MluWB
xjpz2Tw0vSp7S97jH8RO20N6tI1WexDjZuP+9ovs/yvgmcDS2ra7EVj3uVXYL5RjpIto/ilU85/j
vOnwbHHLzrOObMkIaQNiMdksrQLZR7DDFpDUjw3qBau+6hW3B+Z0wCooriDjN1TpLwSFpZLEe3yw
/vdKFogIvf674dzt/XBwyVyqB1gmmJcftqHu9DNMDp+/oWUgik1UVOoIr14nRaMWuhFm9hAxN96L
IUGWUR1wYL1rAl6SImoOhi5cQRG5//ALdZvS/b7sdGQc91gWqwhe3YYZU1oojwA7fFwYznN5fNfb
FbXYcGFsyo946jxrvhFHO88kPzXBcpDnT1hgB2mAbEWKazcJEkDnXddmT6bpgxnmAJfvp84HwhKv
OtZqlBrwzJVY3aHki5Qv+DSDuQ7SHjsgEkoKHVMVn4g0y3IlLwr7a5f7abyFWK8h4tLva+9vFL/F
WgZDcKC3WmXiWhBA9uCvrxCXn78rJc8tSEEx7mtPACsFXq7AG7bthCzW9Gfw6fotBo0wV4K+Pm5C
3AmUEcILEp3xVewGKziWxUT7Xk5AJEuEtOlKgq+O3Dr8JSoNBS/C8EGaRxwFsxfB+xB3Y3beWX36
huISFwuyE//Ss0I/M398ve1lzJjeDnAvS5KXGdQ27f4eDyWtpo96jfa2lT3BVq+spmBm7mH36yEx
Em6K8mXPYEKXOLRzltu4ZJFsP+TVOP4URctcI/QPP8tSCR1zQo8hQQpJaaSQ7Mdq/QFfkSADQoUu
L2a6aEcUrgvRHgZt7s8wY5FoEO0+UCh+GUYzMMR8BsJeNIth7yb+nr2W+ghT9vsJ6tKaJeKcE1Ft
z67gsuUL03l3C4e4MnTKUjoZPR+9sUiLQ4kBwCPUT9Y0Z9UhIeJixKSwVpGHOFhxIdRu4y2g6QgQ
B4830c4B8lO+b6RbUJPMs306SGlgNrkQWBo5+TwjUoEzC++rMJrSxL+F23hESMGMKuXj5EOE3kll
F0vCkXKCL2x/R64nWWXl7WoGF0Vps1UX26SY3O3wVOAARnTs2grF/Rk4SghCByZ6tYTV146qs0zC
o8nMIjFiKFUDQs3d339+Ny67AZIhUJN/a/lKqHMNS0nwYEMNl7Rvqt7nF++5aUxnLakvhwd71ZJZ
2cURGOr2sJBJRe59Bw+HYx0NIH7LGI3Trz5Ub5gXW3sbtve8Ty2cMDdXLE84EY+/1/Yxw8+33D8X
G/puAh7yAjmhxTisJFcfebZrQlUeqy1/VdCUo+bBNUlM41VZ8BPP01ULiLC4lBnWz6nvrfvjnpse
038sTaMbEyYCMFeaLfW65vU3ePJL4688I+A7gxeqN/cfv58gyiCWIJR6dOk4iIZ+tux6xbvsTQ9I
szYykH9p1P6qO/AWg0vOhiHl14C2f/WdsqRmN5DPmQ8sLxp82LpAyOo1k4udryC+VU91+ERaJq6M
4WCV+9MFkXPZVoxoXmR4QN3RK6lF8V5irdiMWe1hSXCBFlJDgyZ9x4tl+SlfV1EdW0LIazKAhiTr
fwVcMSPV0Qnbb6nxezuDW0IXbASXAV9I5g06BT5TpMU18Z3cLoTyEKqYK2HVis5XI2ldlQuhdJGc
sXXZvv3hrnaaaGMr2rVvJvWTDnXnZY29Pkcmrr5r4qwn+mm2o7slRupq/gaADfJ4lhEpghp6RhQb
rIeNVO+JRdLrceQpm94SiVh3DslKjlz4z1Tl2D+zcs+o1NT+8Ian0/WqDvIQPtuYddMJ1l8hqcf4
lGneha6TG7AmSIFa+4Fw34cxm+hKpX3Runv+Opx0NoWYhJCUhe5r+/4DM2qQBkzF3n/nb9NuN663
DgmmaCOxrxJSjOW5B9nb4HHNXKzjERwnzKFBG6S77STtGLY9AzAmYrL8oVzCvVA9ckLfNkSnFTiu
aKYclaFijaVOs7GyR19OxRde2KvhZ+laae3D+BY0Cldor5iSe+OPHzKXu81Kyadfszfs2I7xmQMi
meXjN92Oam8/QLnA+GT6DS0DausuUhyrarfb7cuGjJxZT3aUVULaBZ7sw7tI+JdzdA5PX5ol8RrI
XKCgoAbOF4RFYNIpa4GSQy6V9vtrw3Bv8a1vx0Atfhq2yz2+SKi66OO74XOLeYRO9lkfBrf8jlMA
dDwnEoyEpokEZE99EgHDlRbtoJOQsQm29JwnDrVbp3aLE0h4aZb8UErwsg0eAZ2V2u4sxA00TwYS
dWaTQIC/EE/LB31L5qG4cXlV34CMRh9+FMEwZSR7kvLzsCAO12ZN/AmvTD/vN1Ecf5AT7xCZMOUb
DCE0GOlYWlEPMQNy2nOiIMVb3OF8/0MEqm9qSJH8ESs6vsTB85QT2Elv/ZryEFRHlmXpBXQXCbLR
/a4FvGGxfZZkQgFf6LQgl18ayNpk509BCtctoXpa2rZ4D8cnWDft3WagnkWlnxVy79nUvCo209c4
7tQPkyIf+NGRF4cX5VJ8Cws+4FnosoiCocWNueX7dtqvnKwHd2To3nhLPairUVIv4PAqnYq0ejlD
2QSe7m4PUElcwwT1J7/pcTyfXQ3/q0/sroYxQD732Ci3ezQWzgFTtpHbrhvOhDQ6G28Nz6kEl/Xi
Zsr5d3rA1vOfYzaVK3OIxkqa3DyF06nKe2lp7919+uicEoM0ATiBVjqq1QlARcz087vl/vBc9RTq
WcrdFKHplgN59rb0dJULRWf3iw/ORmqfrXOI0ZAiefxv+e/DxvNaijInxCAo5YfMVKQb9jH5TZqV
5VcsfQwT6gvHq/MhEFUfwJWF2tbeD7Uw5s2csVhZIjsquSGQPSS9zLQt9gyPb8V87SAs9X234gX7
h922pyfIMicaGw5utMBGxGyfPn8LEsg4ujf+voq1MCYPHfGtlNW6KFhnFQw8wF7E10IAg3UHsuaf
x0XP/hb5xgxyZfusMUEwqJ+9PiDjAV9G8AQEJIrx2wKSU16E+le7dTFd9+uhwbT+FDOF1O3JeSuK
7ASuE4Iv9LMdAvrldqzwu3KCgzzZctlVa3Wat/asgtLGAqDn7yAD6lybPVQJxNXe7bvRH14UiUWC
B+WhdiyFPUJwtGqh0qAdJuQLNCYQx39Rv1/lCxAfpYNqfTyDT4yLAn3BUjEW87v7YUHopXCAFtu1
4pDgw+unNKF4nHYzhZFge7d+jXr8hlevGwuLUOwu0slpKtupt/EwtPmHktY8ShhK2wSVf2m92fUp
x1us14n/eHgvDC2qqrgpsv8yUh5e2xCuIyKwudB2Of8w83jzjft4jhThZ+S7nrNWXMs6wr3rd+a1
1k2Hp2NMwXa0svQ39SUVhVB7dv255KR+87bij2B8aQBWr1HerZrtXpQjcQ0+JGpmDKF47V+7KnRz
62hAdx/M1wjv7pqbCBHcg62GllLUtNRpcEK8NGLopyKFo7nzTIWz3RfDvsxAYLntwV5yf97DLJee
ae087Jakoa65Y33gmH8PDYmQh7ezwQ9wIzyOJsZMXo6Yjmi9BVV7Jyuz4Awh7TlOn/qUbeZc+Cuy
HiqsfTzy+oDg3G9rzjJAmT3qmXrQZM4BJKl9qJlQ997DUUqBczXyYwR0wbAXwXgocVFLYu4ajUYM
ttBHkeib2Du+Ayo4YPF74HEd4IUTVXWhX5U/uKOgp5Hlj0ANQ6Yn+6BZTOh4wUJtzKp/AXhSq+79
xNH7GwnxPVClEANo/cd6PUquB3KNVgKLHE3w5BpID+GBY39UVqsyT16ryCjmWLQQh8smVqf2G4lq
kGgavASaHCccvM7pB6692BCihSyomqqyyOJ1c10tCObO0luSncmSHLoD6Bl6A7KyTgxhhGiOApes
pOOktxIRb72EOWOUVjzHkB9/l5AOmPLkwYe5zdvvzxRzky7hFhOIvqmU5eG5rS/jj6B+3Zy4H1b1
TAjW2Gr+5x/3PHXtyaR0aONeVina+rcVjLU9nknkWk4Gx3mjl6uc/Ibtv6x+trbxnajiia1pwn/I
V2Ze66aQw8pgM0ENlYqbUsJPI/AorvoxaFSDfoUvKimiWvkcXKh6kFIJrxu3iPy3R8ZpnJLQIonA
6kxFoQfCegK0mIho51WN7z8vvyZ3gpqO8aR7Yedg/RLVZrFqSmKGjhLpDVQqFnQXB1gJDli7GIjc
Mv0JcMNoZHDzbNFQqjlmZXyFbyydWYp9AvPQF/yHI2OuSJLxOqLa/zWK3/y85saDkPwioJjCPYbg
flNE8NafjgieV6shZuPJdg7wMpfsrNGoU7xqRHxt7TAV2ANWIcplbi6bwgVBMIqxbaqdQiM0pLtV
chQndDkravIMm6pE8UQh0DCOoEtF43VMRy15EjX1Ieu71jk9KZT98tvhQAXoFdcJ7nnhjUJuOFEF
6dE0IOTlRJTDYwA2GokhDbPmL8KjUz9PpG/s+B7m28qgiZTq9sGzpRYgFqlJt3TeulorBPCMCCbe
NVfGVwhKGtsNz2Mg1jiPmiT/Uv9pgiXQq+BnEuv5Tiamqn4buMbEw8nuXextt+TJg1/45M6dNXu/
1oc7XDPe9d1EDi0wqtCgZdkoJEjV2HiZPd7t1tX33q2VMYOjJOkx10xO77Oc9wSvrLGJ02OttzsZ
PqF6DmdNxPZfr2WgGhHXFZ5vFNRGl8pED1ew8pdyaJIMiBozKGOfiqhux/JQnDnoHXGO9mW0Oe+2
0JJZxs2wDeo9nvVhsjB8XucQziIxcLqb53RQ9JZYYc77nUP1V6I0Q3Ht7VohQUhveGJogGRMYCTj
VdxteKLqa8H+DLQGv7vRfIJZtZrW3Ulbol+eJ/Cm5zFu6w7Vo7mfUlqOVZq8HGlUpSyfc82Jyyj/
Vfbk67XQ0xwOlv2AlZkYQa+xxi0wczO+vsHpgNsWFSTP5vGh+LX4UZa7JqlCE0zq3OtyXqOSZxmc
OenS4CC5+rHug/F2t8rUlX0zpHkI1KjMF6nLkDJnRwutk4nBjDbpXMhvYrJS3NDNSqXXdlmVwVKu
a8m4ux9BlnLR4zAjGcf4zyO4pYf4Ts0/N/fv4Ahk6yNfZZhqono9qTpJU3VNB9y9QfqZE+Yir3n8
dqjnDuydPxSDwaaqsEJqyKgBGVBXNCnV+u5Fwryiw2DOmj/cp7DAmGfIJfJTnypJw1TYeEF2e/W0
bZwVx0xqMXiBi7tHqhMaSB+Ur6u8A0a3iJQNI+9J2HOd/xSjcKOhyapJOYBZKYjZYhdW2nG5BJyq
rudgcIGNZSgb7XWnl0YYSrdN5QWAR+RHlP41G3Ula2Zn1xT1ERzHxqDPGICKqv4ojcRPBnFJNplZ
tOEwqDHgwNTbc0IRkKe3I+vOuHDcF2uAYGkKn8bnf/Ut++hNDftXUCq0HUGdj3Mb2Z9v5O8xfYNz
nCagOUIEMZvrErtvGxACAgTJS4Tp26/W5ErkxKlw1JtIShKnzfTDZ1WFtS83qgRpg/o4Pzdt3TyU
ITf1ARziqzbpEl0T+2Xw67rW2miTAC+b0U5o2tQK39X//V5JO2sEdG74fC9qyqUIhoTGtTcBkphC
S9VIA3JjPBblr2n2R9mu5e+UoCgE1ktJv0SZNC421CgAfRyuMRYukmJ7ebCGlaZFNOqIydp9Z5yT
YfR99ZzIAZr/UbnUi5ROMPopEYcozrSgyQsbqa4UpvNTfyDFSxNpR4nLaOsFLDdnzerr5UzAP/gI
4WvKCOWJ7XYWDdf2bpDa+VGjA3iL9PzYzyWgeMhqivY2xkO5EGZpja1Ii77NiksJjlLgKifqTviE
mUODBvkjP6Zl6ZlzGXkoIg2qvPdQ7BgJ8avKAmb8fEjudsaeHveVAS9ah0RJt3Z6rNzvcq5t8A7a
l9NI7rxHULi8p7H+TwIcWPGbdgGy0TTo0phKhOKgyT4Sr3uPwv9R7c/uTe9Kd26JAf0EZVSVRElu
UrMRGQwryC+C3GaIhw2TiKwGSIjGE9So1WGOWXg2+GpmuRv7v+l1bY/jly6rj61Cq/ZxTjNu/7Gs
DdaT7GcvOh0yKUd5KYi03kxuNwbyEyEWKXI2VDCgw9meO1MefYsQIY7ixPZbGhXMv1ZrV0qAHvaB
8V588dbAPstqzaZlT2tusf8CVDhcHj4m7nQ+BK5wsK9BqUtNxrYswLcd03pRyXeFszRRqTvqR1nV
2/znsdjngWDoa9njqJyoKQJzj0viOmlcQ10edr0hNKyK4uuQF/a814geGmDZEjJObpUiB+vTtWmN
SKxuf4+jTPAo4k/agBdIbTvt3m1UAmfJJHs23J2lKNMUQZjOsuZvDjjYcZhhmsl80ofJf6C8TAPg
nhT+EAMhnyiu8hKY7Sp3mnaU7JfgRNzmdMoMVfaGRBQbYjyBMaWNh0XoUpAcyyRpZmIiGRWvm0Ty
rtQVzA46x2yemY+VvF+3bGEIaATfXvJUJ3n1zt2Rjul2rE8QemGuw26DJgbWSafWuaySv+BJ3rYd
b4b6pdTh4LCZOlmYc7o16iPQTMdyyll1fs+xGOJFeI21v5UFJmoWrCrCuqCPsuVqsK6HtK3VmriN
80rDt4QEeYDVJTChZnzb82baNT9HOjtz8jd/ArBDyoZMe6Acnme1EWO8ZqtVescGL12OL5yqEQbM
OG5OxIK2tYJRYMF/WQWdC6+wKVuVRM0aeA+C3O3NePGDckKN5rfZpes3Ao7yD3ztbSLRhZ4nztxL
EZKoQ2EnW261uwJ34e5HzQJYKa5vds0BvN6hIwi5SOzOHuo4Eeszqzx+qSAcG1hMaIbqX43XA8ub
x0Wqpz+KXjYklFkH+z7WprwspjPf7DarrMDeHu/VwikqY05p67e0mdOrVwbytG9FblamzruuXdZJ
r1b8D+6lyK4SCMKJS4JM5toSMgb0z2zUEaKmeWhuDFWBJrCJfCj7oqnPTrwpuGG6uR06NNSuWDvY
BR+kM3jXY3ORxPYtpt/eqgdEQ8HrrtqoSuIOe8VSC6VhU8Iej9mRjacwWJ1sefo6Z5XykvZe0a+g
RVPYPbyuaV1lxpzBdk7vTWbTeg9/E2no/RgZCNs3knzHcLchUN6ep7+BA3bKHx3XbBMIfDc4fZ0x
N2fU3k04aUo6T2VwfEQG9SfZGCJDOs3X+rintDavjfYb6/EQzx1N1HFQj+oL0ExDHqTJyxxOdXnF
ypmQ2OxheUpTnoriCjU48P9NG8d4i/fdTbagcMCGGnzWLBa7mIIKMVBwsBk9KHAYbQFvNIg0/bL4
c9aqHSxse7vEdhtj0GbhAt43cKub05zt4R37JchGI/SXTGiuZndGHvStaB+Ryo9edE2OInP56Lf2
uJmE5MHSdPmtRfIXEColxLN9JhCCw+a1zgLvV3EPhKWLVqbw/6C4P42M92oPqnTawnY13PX3cmNW
zeMIMj8v65yMzMExqWAc4IKxN6PDSNyAzAZhLhEXhkz8Umz8Fcda4dp38W3OyZujXLalx09CivUI
e9koVOsQXTIhgQICWUG5ByrSM/JE5BwSpMSIh4Z4NnS7jVgXLI33uQ7NrhDB0gsEAN7ZI1ipuunH
2G/4m0uNt0+CJYEQuFTcl0QR7vUAESNvG/btd9ovwsF6j8/PglOIoIJ25W8U6YbE3m/sFqPknRKu
dcXbXQdCHo5h4UY2SqKe6JfD6Wc3m5vXHep98p6fxpqE7O1oHp208nrT008v2t5Muy0eutv/QUWU
OcYV3lXvTYc0tey93nwcrJZ/Gs7dGkOUevAXXvJH7XwQh7bufX6AhEo5AKIdSN3ywxs5pULJjwJO
LMvmZk6odfLwxTkWM1qU8tmCm65FqozDZOb3aZgYmi1PffiUF2qnwMNudWNvgtCdQXH47cSH50zW
QKw8Up4eeGBmQQLHvsXluZGZ5bjbMhBuoxMQCjZALiDti0w73oHlB12WAdKAmkHhJ4gwZ1XZz55t
sGcT451JezBTOb8O7r/ol3eDBvzXSeczy13F4tbfKN+m7r6w7cBmPrjONU4KvHucEBxDZ5koA58v
CpJ+MBJlgvcHE6zsX0WSaAG/H89eE0lQJYKYisVR4LP3qJiDEgpmUUdZNj+m2Gdt3WlldhZMXomv
wOWqjSuZ/mSPcp4M8Ro2lXhHmdqrySB7QduBE8zy8tj8RAefQrud7R1c11xbJmhB3f0/jLNKWaQo
wkAfUxjv33rlBKDVk2/vuJrB+eUik1LaROO26o9800ekTEfu+3UzoEI6Kp85HTkOg/eVeo+4f0RH
TDlzwdQ8edfn53SbRAHx3tw4exu+VvGwXxC59FDexXcle5jXbiJdU8D/kxOL02DYioNASh7nLj3Z
rP/iNWMHnJNzYm+4pLE+IgC/jqdPvZQMRxqilEhQqFv+zoDzQS4Sbm3RLJwn8aAykQXmJfmFlBuS
YzL7Z9Q7flV2FeFMLXk1NhkVO9nNxRzLAa2+ArA2oOW7fxe5VPp0J0EdINcjIAOTfu8lIftp1yLS
1tABF9XuqG/2o6JXz/2s145xoV4gcbGijw6DXTqwDGCqT1xR8tSV7lwrjnFETAFQA0/dVzMhccCe
VWFwGMMIEHHvWA4dNLcWdLSszOBxgpCtg32hWVcQiS2/NKUFFSDg5X3A4mMGqoSUgjL2+b523Cn9
OMu5SBlY//WU2jNYR0Q1hnonHD/0c43exC9WImG+HjYb6agz2awnG9wBsxcrHSHQljKYMBLKUQzj
KV3FG4CTMDsm1ZItCkZQ1c940DMXXY6S9V2E2xoV5WH4iX2c85kCg4p8YTZlgsgJcqndv/qZfTkx
MbP2Hk0BNmAdrAI6p1sx1aljN3WF6BA/wLGY98+aPq6FfV4jFlGAxptrTakDK+C3WUStnZkLHRvM
478UD6aw79aOR3ufk6/xRsOvN6YPNgG4LUHZkIbUfOhXOp1JSqYZYMYi+t0ajGWovJa+Ftsqoqcj
+UPzAyO3IeuXxWKBnkdvXDwYKkUFLngqWRyzfDfPuZcOJCUUWKpJA7f8Mn4ivjO/1TvxkZc7s/Uu
cH/XsVdTu5WgG7okAqHGoQBAuncs30wx/MdkQbDAHBAoUWp8zYyA7qQSCtBax80ca8cDtlu8onsD
KVIboikW8roY+7D2CuhI6p+ibQVhw3vMBJOTue7THK+Rmt6g/z0s1XY+60bZnJ78tKiWbNtziZZZ
+GRlcsjI7MAIbEXMhBdV9jyK4TJLzkXHYZ+T/Jy/WgrhI/8o5OdlBb5cED5EDKHEh8nh3E6c6Cap
P3e+CGPUaSb9mmysn88bO4UsXJHwiwRj9FFFsBOYZcuvqbCWTZjlqOFYa+IkpxAqqheiZxxjDJ5V
OwmPhYPSeVQ+OcoYHfdWNAeH6p6/xFfJhaA+VDD6q4ttSrV9ug3JMe+somjusgZX3e2/r1/xfyFC
D0Mphue2TFoe28eET3NrX1zqlvI7ETuMZY6hSKR9Tpqn/4uqqge6p05XrTgEvR68MjbrbxQ8JHxL
KMjowvCbsG9M9je9q+J6lYd7L6XU6S1OxK58qNEW19cx5tKueQfa0YkbmoX4eM88rSPWlbrzQG59
PG65xQ8zWUNzJqFreBlC7HyRtSNXs54pvkaFzlCfhIKeAbqzyOrA5lsrw42dBPk+MZ7GJMl9jpQI
oQd84uZ/orieGdXNOzP558+y/kUG4lty8l8vrPTMOQRKWhhQR2G68ZLSvCqy9C6OKZyHVL6jw9FN
usv+f71QLF32+iSr/AqNM+jOf8mHkiOwrxhVZUtpC8O3Od0s13OBtE/DwPRDrxLcktK2mxntB1+A
eO8ALzAgfcgMKpzPJNu1Bfezucvl9YqzOz5TYePBa6NxJ0YPglOp7/Mq+N/xN0A07w8vxNSReHS5
lOoj0eDXaR9paMLyE+N/GUnDTSblq53tkZLuGD55glJqDOZ+l97zCm1o75iR0Umi4NjS44JmnImW
vo0W2cnsxMPv1NiJpfxyxRLvcTB75XlpPegK4U0vzZQW/JsBTdDaaUZloGwTUU/6QVz49p47B/O+
dK5FiqBDG4prdYe/YsGehtRzWKoOOKkKXGq+wdyso9xPAE5JCUuEwCzH2WKtyaPAj6msZ0rHzMrR
SFeta8EuAKrsXnjHCL7ouDLTy9LtzHBxcwp/uNQNNHblJinpDLjZig0zAKMDZ1FBO7ZFVsLUrZGk
XnU2N7Cq/rWD6C9tBoWWFaXKJ09iJBb5CxScJMnrnoa2HxKljdhYQW4SlAgysi4J6+RGcHzHpV2C
uUb7TbV6o8I/JK7yDgGx2hB/GP/Yr3Z/NIbUe/Bn8FswtkHMR5xPJI+5eAmSRCHFOAL7bvv+wwXJ
xS9Un5cFgNt7TCVJnW7Kuh2aSFW0/U/+QGg5W0hz3YEsUs0kAK+K+WBpbn8qewwhAcwFALES0mgK
mOmTDdrTuPquCC+CQTjjTnt4ti0bI/w4HZEDTaFigX20qCSmPdVQB92py4yi7aox5oLlMNCfFMCa
FyydEqrZAXPmu/6pYY0OtClX03rzu0wfGuMMsA5pglYIY7yLBCkIT1SgiLXHwyB81rW/3RthNcBI
+gufh1OmB4YT4uWHqcCzQSDzoSmP7Rydcpc2mPt5STTe4DQMx9IIYbgYalOCWnAF/MLxJVKp7hNk
27eSYCne24AJjlHIpAdC3vZjCIEdq150ct61WRjPPJy5swg8Ut1loQ9zeGa7qBpX9wIZSlXv4LMj
5/qVGrm0QAJDQgkX4zRucpQ/FIqtPXUYCCot4r5P63Y0aI4CuGMwLW/PkszRU6+NnciE+FPcKKSo
MfuPE47hmQkJIT+muO/iZ9hIBt/9xIzaWdg73xKrh56d4gKqcmFBbxmBsmnlEUt8oNExipIw5+YT
IpbTkmlD+vrAY8xgx9KV23K07zbKTjsaCmuWl1whZ25Ny+gYdyoiA/+4/J4ApmdRjED910hz96Zu
ZBLi/30tXtgRHh2HvFC9AfxcmoMy6uSKsQf7YNWhqSp9X6WPhuk+vz0VtdPoFWo0GRh6wjRyiP4N
BkY99LwxKwsQ2IUCkUPkJmEfiYgHr0Xao4GUEwspjdRUkagjHh2685/fx1rklNqFXsBaNPiYDM9I
TOsBHG65DwFPjaNeH+UWkTV9whtjWW0hkSf/635uMB8xZ20Er55NhPQbRnFym2xRynbWSlsuXWHz
cmeXnG0q49lLw3VDjsN+BFKsO48zNlpfPrpnE6KU1oovYdGyYQoDc/9c1Z1AueFPb7MzLrw8Q6JN
jUEhgx3Tnp0fRW2jfcZlojk8Puw10thDkTaEeEPF7TQ4xrsWyiEMy8+7VTdZAcOTSQEnjNm7zy1F
a0RTdGcPIww2kpxW8F93DR2EXHlbFBQ/i+VznD2a+6qMvIuVykqLrFJFUYZBLH4N17jW4oWI1OX/
i8VwR7DIJhX05ZGJJlK9T5HqVL4G9EkUsiZY4UtYgMf7WJ2PY+zYEyph7Xx49kKJLU0nZYmHGaAb
hwRxzQyWzo/YbzhHV5K8ZyrGdgzw66O7GeMjwTnzvonD9c6vqBYP3c0eJvf8rosimwcH5j5I3u5W
VzAUIn7VRTvr73f9Av/yFp1SmnDqXwo9amUmHEN83VBwd6ztFW6KktI+miqQrPViGEW0dlugF1gH
L1TqsTMM4MWiL3QgvXLQVN1XvgKn/KnSCWLo1+GvMANA9EztteXNxEpDgLcTHMtpdISUPo6jB622
jR3TnLjmsuEGIr3HHGsjCbo4gnlKWCTOQJsF5WmtwVVOIudgjFTlCPpJOCIPvji+3nJgFWB/w9vY
ZJgfEFuf3DYZmDpirqdR/FYI/62xwEb+SBMTmP9bXDvlYTtItT8PotwAaaKiU0ysXFMfhn7vdudY
nymBxKemoNbrKpv9YbfCFKnM3d4lSoDzHb720uofSDzXBqnPp7I1VHMhk38um1JMj9HbWRoEKqP3
spnpYHz1b6fMxybhNGF6xweh/BYlq8XbqEZs/eCJ8aCte4vU98aM/Vmbnw14cmhwQ0ZGvH1ELjEs
7lgo4FsbNKHo1AKxrBJLxs9niZPgPxwlupryLBL8jWnu2ftT4jwRTJLLZx44PxYEvN0w3Q8eJdNi
+bKjzNyZ+8tlSkiQwdP5i3ouQtu4Uz4t5WGeUGxYhHL1AJ7I0GesJY25HJu6J8mRYNbyocKJ5HBn
cShpxZAkCf8QgU30OChJ7KwDdrxSGJ+DaoSw5j0AQBYNVi9LfXxKqxBs6oLTKbUmgeYBmUOzNANT
5RGbX5Y2HqzF9jDjvKXDflRb57vGfAUX8AH2TeYLoTAHG6YcOVLOuGUe7SNTNym7vdvJt3CPiIfw
z+rvhA935aTZpNBqsj1yEai/2+fm/jScY+G1lx1qz1U59SzbOFogelrU270DuBQtrpcc2FVI0qsu
6ExN/nwsq+XYed5bbXUWpSPEiqRkv7br4UArbklVm5TXWBCin8Qqzv4+6wSBS160nlh2r3S2jkX3
ZOIL6trvNJWldvD1xgxDVudlE4aNZceWOnrXuJ7EyKuSlufIlbpUSWVvgm3a6Kneil6k+7Lrdepz
/QQGcPJUweyovHjo5/hG8WBSE4srfh2XyFr2BnLZh0+KKqyrQ5VyiBOYVpy/HavsGDabBobdOukT
rF64EzqwXFS+3rBq6G0rElTcPdExmsLcqfs3ODQGoHtzwm/aGE5X5CxE7s3q7d76kIXDU89+3y4/
2et8n3NEAPEN80h4gCPHU2tGytdtT5QKPlg+kqLs3wbx87HTINIqhJ9zmSWXfvOB0qA/6BF2l7Kl
oIlktMMBdZrit1GoV5Ww/z2ATZ0VTOZgLySKZDRpnnK1wpdCIDIqC7lyKNRX856DqXBbCIP9hPN6
tUtlR/veQiZqahspngZxnywXdlh5cCfi5n4To17ea14aPpMZcCk9Q+5vEalkb1seJ+lsno+iUPxy
2rqPo70ldycmPm/YTDrEpN0SjW7NlJ0oQW9asxyP3DC3xPRTmAvZxroCOAxQSfDCXhFdBFZJQDE6
wkC8UC6pebmZ9CSpNgH596ivQfVYxKwhBhf+rhQ/UWVddnR+7qDeItPOaXmwmKig+fgmIB1O/rzZ
Xo3jgRAYwkuw153k81DS5xgoXvXbYiO0PqvK2pD4d0aLOEkWcsZ08I4fg/Q0q+OxXT7h6EKnEXVu
WYXrPuqITo6S01CZwe6HXcW2odEzFS3DwRkPF23gxs3iewOOncJ6GbyMw5/P4hjZXvu+7hnCFKT1
VdnV+qlm1cUAKqFN+0BSzPWDfoKuTX5Pe40uRSnbjO7Qks5XDIfBK4S80xywO/HqKiRbiSJ3RTPS
T7c6M1ObXhHB/P7mTPW4SPA7GmfW8RjdxjpdN/Qf7gzkX3h72I9VK9V1+8IbPbgkFC1yB1r7BJSr
8101QVZ2gJ/up6DFyMuEKYJJL4IsPVDgP7xUxLemYfBYLFrRkyUXdtCjm3lrg3nOFwJEs3ZG1Uv2
cPPzzV8DM0X0fA8FjtSIOHC1TXjR2nL/o9hp+FQCqUS7c+7S9PKFWzMAMMfSTxSmZAwJF5LwLLqH
yHwWjdtNUL6B6ubHANmYM6rCaG6PyeAJWxwrH0LzDVfaS1RyZ3gv3VBDHyuZvtMyj88OhZaoMhHF
a4DMJV7vcNsuCfH0Gv0/b2QVDPQjSa3F5iFKsuQDA3Dbh84gBXe99GEkoITP+qB9mlmpuC/E45Ok
jXN+wWzg6dR5YF3lZ4gJ1cf/uEp9XW5wvKMvZZy+2aLAsFNLn31bwmxWqYlaC2t3N4hmWgmgH9j4
C7eZSRhzoAEYOIC4mJO4zHYF8K0HNv7Jg+159MWnKxMj6x7NGC+b7SI0cazOF6vewWw1mrabqc8T
bkBTG1UpUmYWznif3FtMZPe86F1lp3Mj/YD92PbgnqUnS+/2LOAlV9qUJqLU/WlGTOE6zUybiQOx
+bv9PlCpIJb8199/hWHyk5T8pp44pq7VyxAyrYY99PzWlOMUkN0q5S7FEXRKZWEilXxt60wLwa5p
eb03WrAPWFMQRGAFtZOz04lUwjdGWCFTw/xSftst7ixHpSKMl4M5dYruq+5D0Ny58YCLWinidqXJ
SQWqvhFkgVWKpEZjH/K9q0qD7wucygy+9cOYSjH3vdcSz1A5RzUMr7np43OlqUkSuLzQN04lA91e
Y94gu1kcB+qt0STGPQvDKiixor7/IJubSD6mkZAMS9ZHqH32J4RYZ2f90dtRKi8BwUc70P6e+0Aj
b0KUbDmY4A4E/Rmp0TKNu5b6qHKHgKd3IN3Lmc8X/vZIwnPkDSAyyoB18TdiOqxxAozsj7kgbplz
fNuPJnIPZHk3wpa7Lhp2OQl2JI5EmVcKeOMO2sk0G/R3iBMDkd4s+iQs9iiH/t7NkAv+IKiJCKye
6YWERV8OXOy2Nl8fBxmiS+LcjDr6MWLz/iujUNqL0kV4kTl4klN87RlTaj/alb+IZTFUIhxoIB+o
CYk060JT3/643LeiMp7XoybsuOxMysBeEJ3XnPDCOvmv4yBf2I5LMSOWaYm0faLmJvqx/dEVY8e5
pSFZLTgV3HVSFfBrQ5bxsInc2b/6C6kPYPh1dNP3DIK1fd4LwU1xC7PvUwwh4jWdngg3oN/F3Xrn
dy6sNF+zshD2xNtpnKoda66SbLrEsHL4TH7nrXePNEvUD2+D+7TotDrxIPB2cXxYYGwMlSXWWzIv
RUW1DVoShkEAhGnL9VwdYcnkDUrfJIkuT3DuiizxHRNBrO6Iorw/h1Hc+PbS+God+78v3q6Yi1oV
yYXSFoOqWgCeEhQN8JFofMowxK/LfshintbTLkE0ENdBNPdI7WLa5SKfZONvmqxzrxMaSqOz9Bpn
X43+i485ocaDTPYU1hFuz4eVnjG9s/Y/gEXWzIqFnY7GUMEgK5+AygcJNCKGnp7aNTuX6ZsM8Ss+
LUsThgpIEQnFA0saxbSdxco9lt2bpK8p0YCxzup2OG9q+b/gBOl1UDh+l2cMxEt+lskTACzobeep
yIwWep1aHGL3oEf4VU0UC2O3JJ1g1KRNtc1/eWTwWNQsA8wst3EguscZsEUGhHWJh1xz+WHl8Rgf
7qmYYWooYucKRE88nNwP7cEVshzvoXkmgg1cYjDv5f1vS/C1p19HCd7ouUQmey2XJ1Nzzx00J58D
Wy77/SpR7d2cU22pfHMETbdrn5G9GWBYEvMOICkD4NTiwIl4WPQaIj7321lBG9kfE4Rfx9GUdBvc
bn2imqVG4XfKKhlHt5nlzyxSId6/0qDMMKO8e1FlkgfYmEwa88odp0lnTfDZWV5PULu6Wk3GGux/
xO99rDZNkVBZ9exM2oUMO/+2xGnWomBstYhDQc93ffICZu7gMWIOwg61zNStzBBfBuvAIEmxWEjb
W/jXIZ/bc3RwNO4txqGCxEE/KSxuPU6jlahD7PGmWW915gcXnINcYHJMBtLFtaRAYMw2aSmzE+DH
zSpPRtqLYyYmuBAJntUt5t5vBNb3fhWVgw/oQld3yNHpvIJzplC9QhgAWHE39uZxJWlYYyTHYb8k
aqT3z4AeswYpuqjb85U4jY/ilvlLlyTDQjpRR+U3uGof74YGEIiRHkhvWr+wVKjXnl8gt1hRyzTj
Rfh6aLcgN1R+ku78/6zH13xVA/4sBmpcSGrbiQOzXYQWmVrSlVlM2jKrV1FVneACO47oOUOjE3cY
0ossditw0hxfE6sfhtgONWQS6ueSKPbz2PaIYBKpOh4BtO06YRVrHi1HOrcPI2/VWAm1b4wbZc5L
ReSepUNd5WJScklGUrKTJXzDigq5xmicYx0VFKI14rjB4bQwg7u/VfqvNEp1QumlVXFfBbK2UqUU
fb8Ud99tV6cpRxceSX7AH9WpazPl7afy2KirwNO6EC2YTuMXsH2YM97g3eyGg/Rf4pi+0XiUSEpw
MeSBQqYbulUFV/C/usfibF6GTGB0iG1Zdjd9InTOz9dwn1bpi+g0iUwaFO6L6KO/9S8q3oX46S8O
jFu36EAURdtsxA8MCsYXr7Bp/F1bjb9Jzfonni1104jM2/valgWLLZw8VpaRZiycj4CH//iUfodq
4vhhF1odzElfOJoasFPT9SE42av7w9ZecGDJjLBOCr56HFupkm7awCGwrbc3mkmolWzpjeNzIJBm
J9qwufOVw20sa2hOMDka2XhQMtAFO4Kj6c4DA8ppWJgpHxl2vjp1b+aZOQ7D4AF6i9OkrHViE/ch
EnKsJg7sEE6jyW8n70wNAjNzzpAnTmf5On++3IjuLVYlGQN3pzHNwQa5baRgh9+jScfVu404jebC
IUAgIKIIcK3DYXvBzllBLS/5uHa4sbNnZ/k8knZHXheKk7Trj1S/erHLRMJ5voAkml0wrZK3UiR5
wwgMgt0KrgojbRzgacE5lhZqYMpV8rMilOiCC1oQs2udw3LitlrO/XMEfKzmKxFM4pUG2W8nmZ/E
KBcYWsmkDIYzDHneHy+ljeq+hYQFNzNHLyi2x6g1obfhRCPPNR8yfZdnA14jUR0VuwraODdHtsdW
ZUuuRq/e+LhlnANuHFI6kmXOAhZBqFurART9zIamgHKAdgtoYFYESUeajqkdcMPR9daNFWbuoQyl
TUeKZWa9mkz6SaRtDAqsImoeB+SqynvPNC2eNYU/5VgNv63MeCiGLfC5twyHrulmI6GIZh1bCv0I
xrpmKy7ifNbOLZxX4TFwudXxmoJN0EkyXCbfxcu0cY2oKPBW1LSmCTZcw2q/vNK2AUYzfhJ/PGiS
q0OD2LJyT4+hpSZ6FrzRN3d9fyAQby2vNJmEym40Is15+6ww9MFvF3IbQfCbodQ9QlJvdD0swSJo
6TdJPBcJ+9EBHwzfIhgpZZDOCfuidcpP7Lr15EC0JA31mlyP9JHt/BAcuoitH58G6JBt4/B1A1r+
PFxseUvIPlKT3Gn31ucpxeHM3S66h2Su1BTdfK6sIUsXRYfOUHRz3ZFC2N8LnMsQlXGQ7JM1zjUf
3JxwYI/wqhtbPjtUKoNFEFQPp5QNAaS59UVnPlJ3iW2u6H4LSL7gd+tn+EzrIGNite6MYA3pQPCh
mHvo+O31BAONJIA3VRRIZnI+w8Y+tLdPtTT+l9hW6U/7SbsoxIPXfTDe3Q3eapzcr8j7GGKMjvDq
F60CEicfOVhy0CEWmKapb3UpPxl7oDADXcsfrfSfvLvI+TYYm3tyQnX/6SAL5HLLHo3PUS7Wf2qS
50tXD88CekZ3fBabs+QDEIciHTceFOOZzEnR2Uv+XNb9BYuxcqLAiGWiTvX0KkUUaoe/+v+081wn
3CVJgAvu52O2B93UYj1FdEvEMFcH99dVjqKuPWoBNl1941XYshQ+9QJeA4dCfcp9rSvHjM+5GWrC
Q5wNoOz4YfWOqnOlX8Q8KD+o8qnnfOePF2xLLztz6irl8aMjw0k30Q9FtcQ4OHeOIyEuCdhKizax
ldAj6tK1EFEGTV8gNGZP4p+f/VazE3hhJ2Tpn07pRmsgdJ8G6y4gsB3roIFYQTxk2ZjdaCxz6v08
EafnYL0b/60ew9AgJKVkMuuqKkWHcSoyqNC3RVz0e7DdliznGKg1yZhevFmMI+vKkgPfBtHe3bnr
GrEOUnpdjnfgYeVkh7bR4NHjXq1UNEA1KTF+G0HgazGGuS6Vf76Wr//Rt9/BS5/MKF2UQ5W3VFDb
6rEhP51AIFowvX0BG+GO/IfGTAYm8VRyMsr6jcfZ/2LHYEClrg8wfqiF+917HZfY8scTyS9OhKph
hVLFRlYXxssFCQiQyZk30D16gne7JTk7YC74R1+GmNWfn6oALJgyyr6cZAkGyLof6gojnNjFYHtD
lENgohM6rbvwxmC0jZsTX5i0wkYSgO8Ou6YtAeWHa4Wh3Lj4fOPJ6dQqmBRnd+TjRupgvFyq54me
NoG2Lm0trGHVoyAUIy1r3UWOWHO7dynEs946maMZe0hhmEPHD89QV4bBOAERaOIni2RM+8Z9bpIS
8FXxAlVOhL6QCF1eE5YN1RYZf4FqTMjCeJLzJNiMkzU4a1O1EZLdoHMYriK3Og4W4KzHshIm0Abm
CRa9yxGSK32hk5vryLoOaKJbZX6iS4q0gY3PTomrVq8eeZ3WwfwZ9MJU4x28r4bgc8ofDl5c2ABv
tViTee1oR8Z8+J0Q7WUvABSk2mVxorE7Be1VEn6x5LC570FZ/7B+HK/fTuUokd0vdCZLhYFVb474
x0xlw5mje/lrTIEy+5QufZ7fLQjyVKaninpx2xespp3zI2MU4kkigOOt3yz8+r8eG/SHYy9cGHUm
QtSQhvwY7VXnaOm63y++yASHrLw5nHT+f6XOKeH/NEzxXG7t08lw6vAeN0WFWZCKkQ8I3ygRvk+w
p/hvxb/RPzepDMr8HpAqwWhHhLFU5wtKbzedzCm9k2bpE0ED6Jd//Tdt7WXYqX9P7loAaBU9Cwy5
5N1mgvm8chZi4LEq0gI5w8bncsMzKfNV+iujVLuujGCBhkIMuHBO+9OFirpjdD39hf/p5lDxYpOi
IkUZU9v0szYitnR+y4klI/eDROgCtSwGnfs/KwLR5pOkQQalul0b3RbsFe6SKJYeghPO9Er+4UPs
+scwTUUfMRTiRAzhZU6fgZCcyjbRJ00EWiqr4i126Iogfa57TwDj0vf8aDojefc+FUX9zix72oLm
8dJGTjbA4GG5nWbzfGxwFZVjRe1si4groFV+UkGlZxcsLy1wpYqywiTXfGhDEL9LdicpH29T43f5
J0ZBL+NAdzA6+fArvHwHQZbLMav6zbOZFBYaKOtzQK4e+sCISTI2cOC354h+oO3nh+MebBCpqGCA
QcTaEcGnnFpYw/eBLKzyp4z7C6KSIBAyps//iM1Zt7l8gvWOFTxtIodXnlBb8kWcbyiLEVadSHJo
lcgYol3NLCO+xAKRvJjMoya6+OcWnQJtWsU24a3j+aF2VOdfaXEdj1RXwcnPoYY9sU2uEr84yQ6O
IOS8OWrIeiysafx4g5v1HdY7PSwXXjylPrsMBoVDssQqQ/NXwlnJ5rvExvSb/obCHOXPbGghacbR
9gcgky/oJ8dLEbjjyXZihWFa/dTYYGNkjZ5LnLrXiB0yx8FX0qPFeqPlngbNCXk9ALznxYjYApxl
IxO+hB2q396PZQltt9Nt38aWAsuhGsTzhf0pDQX+WJWAFunn0gnNrPJBz+O9UDmRLIT0zaLZY0w4
uwlVJhmQgJdKqrPgyf7xn5u2GR26bIlvS7SnJZ7R/qdpSERY7FGs0u63irf/745uHgWzUSi0aYM6
Ci4oiIpWwGANLsCMXqnywEZ7nfXyJvR1s3fQofncYTeI1/3IvSu9FORX2SX/DsE3s1Et/llMF76c
/LsXIkhJe6xftG1W5KiTHsN4YJnREHUZOYHpKtawx0kcgKUtaRJeoA64ewcrqQvyaD/t7jcKLLa+
/LxlRaghZeteSew2nPkJqpn1kOCtBgdUxH1r5DBY7FYoPOlb9826Rm8jBLKo/gYoBHnjNVAMb6xJ
3ddTbe4NGlBJhk6VcFT/Tqzf8CmrmNuq98iUTSJkt92CHmTKQJ6wW+bfS53tDsDQNRlix9sCaxVS
hx598LNyGXLu7z5SYiu11EM2r5tqDH/7Fw/garQg2j4ncw4mKr9LhDZDwtgxnLK8g+twFnkqqVoF
57K8majVPnVzDu6R9guuAhcTBQ6tTVSFgXHQ83sa5zR/FvKCWwd1T+HXrlZvhuzYmp0/GIxygWvk
rJIWbt9Qcntx837rQjPSDyLeo7vxsMERK1mlJ1IBOX0r9Z1Yc3JOPhu8IjQzsm8OpGWi12cVpsXK
blDERKYJViDU1Gh1La+DXmlGFWXmemgMMgyij5dXqjeHIwTAzKigeP35wxL/CT9OSv8u0sk8qjjP
wYEZV2+Cu5uBNpmf3I1vXg8RuFYgd1ExCrwUnvPk9ypMSTg2c4b5fRXGugbeoGkwdra5lIT198tP
RtZ/ZpC/ImqLYR/W5JnBgNt4SJsXiUziAfi1VZMfdAvPLjs7k/xRt7dQeVIkhR6wv4dsXj+Q86+K
m5wYsWcddSjtbnmfmJdeMGUglU415r22f5dafqq34dw5uW2yeGh7eyHqnPC/iIdtH53m9ffqgVMm
JDpMgAdd9tH9jYAVTiH3wnxA9JASjoQyXgYRa+XcTXKxjVjP/1KD1SGR1JF7NpOpxYkaZCV1gXjk
Lqq6RZA3Ro64hu9Pz2lXVWRgQ/hIuz5fXlB132ZUDscMVOX0eOpv2rIVEtfnTFaRiyHdYdKN1zXx
NSCRqD98IrTAWFFqZ5ZCHpPMqGdTLTmBUqL7y6DvDB8P/8goU0wZLErWN9T+LRt1zhovjEMzgmWK
RJEMIFia4/YMOA1XCmLDDGd9HYBtewQq7Vh41s1EopzpjuUnFb2oHahaM+V2PGDn+LdolLkmu+BG
eqb/gJpncDdp4JNac0ho0py08fKfxOldfDPXAtrKsgIArRqoqnn8Monb2Dq13tD/ar3swmlPZ0m3
7tgYOksuuJBM8koNB5AIRx1ZpuX8S/xt2UO0MxXm1guwUhiosKek5BrAUJ7E1aVNyh3RwP1LFnxH
awnHg8Mzep+xa9PACLB2yw3OxoeoiBPiMko5N+XV50jU0/q2g/JibgTlxrmRya+d9M5+SjPknI1j
k7Q0Zlzi1zlV0SvMHCU3KyrIU6uFCx3NYVIuOZO8VRkvBYWEZZXIi1SwkMrfcIWI06hUNZAXjPgo
icbpg1sawo3u32HPiUZ1QHYa5UmQNyfVhDI/A+vRBlxAf/DgZxT7Vi+CtNs1mRbL7xUnSh2jPWmE
NRiFN2x1P+rHr3hDly0rhz/zB4jLSWHfKMxAuOOI7ByL3eMXug5WZu/Lfzn5uK2J6p3tVI+dZ2Ew
kSTuJzP8qn3A/YlCxsyC2keUO/YwuGKCpefd7qLtt7kOE5umjoOANw82XAbumi0zavvF49snVGIT
Hiu+GFVaxaP0DeHQrWhkINI6MhIT1hQ72iIPJCUPXeptB2vjfWBPCp3/JCbE4i+IV7PfqY0Gk8P4
H327Y4i7+7rwUMbjJ5TbiHSuIobNDkOUzpmYIEqrQu8yS/3ceGQKkEaoJbISacAdZEp8VXwuRhhv
kforPIFQvGa/JkScazkl2dVY38hz7Go+mdqY5Jd96o0BgxlUapr4FawHz3plzGZpttiphUQJMgxj
mA7S+vs9IQSTV555z99JBD1U3y65PeyztUbPlmzMM9VD7ARvu6ItK1Z3Fx6Qra9s2Qk4MpQV2+pG
P1P0/bbXkU1ZpyhyxCQopONDISqa1HvRB3KiMZyG2Rm8woSOZA8wedlH/HF9tzrC6eQDg2H8mX1S
KoTP225ns6zVD6j/jY4mJB7HVYoCgKQRVqRVXI7yuFrYvzD18GM2MVO02sjK0z/4FFvwyTN2NJHY
juIe/xAstaYXXNwlAlnhMDf/yHRxPb2pwTfB6RPjVXoYtMKuHxyO4cNBxcXgSGFoPP+cqd3Oxhzw
UyFSMHZk3RZl08QCEpZufOeKJyimsNKVMNcJ6aHSIXW9PgLfdysJ53Zd0upVKU6TP7/16aLh9Cy5
DesJTqGqDG/21gPlo3qQJMzd8UThWOErzun5ktqBfJ6UDn8wmG7ArnuChDgl+xRvQEAk6+U1B3Sn
fuLxdWYIHfVvmz+wgUvTrm2r6LXK85ta2DTlYSJQYB4cnHHZ/LGqNW0TjCAm5uHrxz+35OggKmeq
OsSCeRADcpylMaLbmckHbq91RwR5xbvQnaL6bNO1C1bCav65qxXkX+fiTt3OgKnpknfIbJRYu6WD
mF+gf6z+VMYAra94ncC2xP7VGXaa77PVjoMdCxI8oHlJnCrB6pyCCedfP46h/fh4JzcngaSlT07z
SrofdrXkCizfwj3Mxo0pp9zQVpQWD2wYrtQN/SVny6a0Hm6JD+LP6ilb8gbNStSIlz76/JyqHNxq
e8LFNd+5qhDiNGfEJzX84TZY6Ku59lBQktEaBlWm6PAv4rSi/TUgIkITiUFjivjXM/auvOzcu7JL
0F/XPvTYT9hnhokKT2zhMUzD+ycXxQbAGBNiHgAax/kUmfeM24OlHh5XeGt6dgHO2QN+erhEWws5
b+Y01hl/m7yZxg2TkN5xXuMPKQW3YOpWUqWZ2GHmETT5d/DkbESHxb9IHRvDsm068zyLO2Fqb8OU
55tB8nz/IfO/+/4n7wJ/tsZiPWBPj++Y47CDeLJfamQIfOsYjCg4P6Z55ohc7Gc3tZ0mFu9KVCXL
IM4DzsiWvQs0blrovi7mI3KeLBBWc5YQraIgr5o/MRY8jLYgg3d2A+pe1zxeLcm8Vwr1dW4IECff
E08lVd4SspafEXJcCrwOiSY+J+Fmf+R3smiMf99XByTgRGRZ730PIuYG5URvxbrHYJ0MLK0Zt3Pj
dnJcApIj3SgTvzEPhmiHNBHPVtsL2vAellp+/GWLAlcgLwsi5Px+gvMROxnPP2FjQtViacIUAree
zZcQoX6Dvv+AiFKYvk1zJ4ImDWQTEMteX7QVxu5vz/bT6xQqEoADNVgSPqjsutoyLGNN51Cyj95N
7gngRiQdyYFX8MaV/wiOxijl/dMhfRCW0tqsb/MDSLwUz3jehJqhB0IcrIVLahQkblICLAn37VSw
8MqNDvaBnZ+I7INqQIoo1iNyvAjvuthJejlyIY47bBSsJomUOOVjkCPf0zV4xwRcctmPXACqO/XJ
BpaFUrhinyJPvKL1mxx4rGzW4QucDLxReYh7r1Ml5QDyDBR7HBeCh3PvCVqrfoNN4NjYwLFXG5kw
MVQqD3Am57DGoUWJGA/75dwMTkjAzmIHKBqHBvR+gaL108kvmrySiDW+wj2dZFXprSkpXew7WDgz
M09p+929rzGSJOPOD2eigNrF8C+cSphuCgfj9QcAPOdrCKlHIIEkkIOdtjJvHv/oW6r1FR3Jf+Vc
9X9eYtIqTmIozEPGETdFKi4NochsQ+Vv0l4mf/TosUlPEFuhD3xJucTxO66pvhw/7uhPYr+uSOT5
ljwbs2rC1se0boHBNheSZVvzz3eWtB3/fNf6RajP3CNJidhvmPbwAtxiDD0JFJBZxNwG/ALkjSb2
2ny48Uoy/IVspJYPXRNfqfVin8PKqRbr5S/6XO2iwnvONvNlaThRHaWCcNMElQ3Xnc1b6ZRAug3v
xM/exBSrM+1bZymUKNfKmcfZQx3e+qylzSDJCO+mPekJhxN7jYyoEypNZdJ/CV+pE6Yin3GffG/B
FrimfYobnlahV1jJZyjZ9UQtVWfGiE0wiZjWTFCwdqRTvo/02ln230thZ8rudEhLlBmX0Rcvy2rr
VzDH3CIjIqMxHQnmou1S+CsqNPOtNNJDGvYa9YkxMhdeoD+zB578BCl1BQ4W4mCvG0UzIF2r2dRM
jaW0ts3OHhXmX84wPxh2mEtC9towcP3IrGnAUAuoS52GDzK/DCZLWHNIjHPgvBMpFLLIPHJT10lo
TBgk4fnv0dtzzbFKU0PzNxMRplJdV618+SPMzW6JRA7t/fg63l1MWcDVxsxa3wHjiEF3sKcO0wZB
tHgVWFZA6hGWPd4hdi03YmKP9mnsHGeK3hKDuBWV89jSRskn+oONGhINzPWNHX3u0+ObL8Cm+EIu
uCMdn6ja4E/BFC0sYWeFlAqDt0GBKCrfwPImuPVV/jRDCIFWeRIhHfX+Fw59g40B6rWP6rXd/KuH
kokpTRxkiPGUWjtbifu6Wi/CM+nsLT/KqIgKvRdIYFCdsvivGCsSzwOGi7JTXv7Lnf4pbzs/FZIw
6YUY/fnxUXxHWO2MEFVlfI7iSy/tT8hRHfoyFgMKHOt3vxzT+v/tcKJdOoN+2sZCReeanpbz0lPX
ybl9tmsOJJ48k4hqUjZ++qaIWDbWL94HlBrpBtvwIQ1vT5TWYYevIvJc0PHp0Tgzc84A+Osibcyq
fEzcoPkI/BCE49EENH8xMoQdKMSy6ZbOJ7XOu/GSOYhl1AVc8VDE5dOZAFFxmsyKQN4OrU4RUG5o
HCIfHdfaN357hBRHcWeZNolb35xaXUesj1FuRPnMqph8ArwheWrD91cEMB+a9c9xKKnMOJJluUNZ
AP4QCEoMEVlljpfn9UF3KZKVteD8rC/v2Cw6tCJpCo1hD7qAE4BqjPPMDWU49PAvhOqiR0ARC5Fz
s0vz54b5UPAitWmZMZriFVH4ShVXMveI/9nVVz6bcqSAggQpQEdpXvIG3tUCj2QQKH34VYn0CY7r
pdtoHSWICG8afl/i9QCDWc049KZq/5QoXgBRMnsO2w60eItLD2nOPbBNDBR8+EQwwIWf+YbXf1ez
R/U7JGROvdMDLwwQ8HZsaDquSIahca+DtUiNn7QUVkUrNw5JbLPXEk8P/Fl+O5QS9icPvsHTgGs9
O+9YfxEfqYNZ2MUhCinEQQVZU54CyGgXDRpzASzKyeQyy7WCgp2XoNEKBaYyoPGTT8SNKab/38RM
ralL/4nnwK5cVOVusBVFTQ7G7Kwxiy0OwtLLEILR4N22gATVsjRZXN4zrJLf2kFdgc3z7ZbhemSM
X4m5nN9DhSfWuGNgCsApIEFQYyHyEox1gLxi/hJjvLP1GYP9uIpOZG/4eZLVJvFbe0lCVICvwdYl
855ZHhYLPwvpDhXXSxZGqW0eLQZ2YV+W42LS8gR4J91Ev+EkEo0tgyQNjwdzNlBElpC3cVgdWECT
quu4ZbsKguTviaywC8I+XGKNv/NFL9or/lPZN79sTYdreNZk7jCiLcAk7b24R+ung4biqWjk13BM
jZYEpF0p6cZdGExNQjr9ZOZvUJ/j2gPIHDX9j2QCMFPhumKwRziUve8Fv28wL+vfuMDGdFQfz9/+
y+zBcKq5uI4rOg5Nn1ycmrkr+eQWaB7XX2Gp44bl1SBFiyMMgVu2Hls4TvHmprPe4CXFPd6fQ7Bq
7zHvW9sIQiJVJPsSIzIc1pZnaXTzvC1F54BRMLThK/MUbtcpXL0uaaNo4fB7DFg+r9HqUX4z7tsA
nbiNub5xdu2QkvoEgc0+wj32nRWahjpf7E8kkgVNqtHa/tEVCabtxYdAjxM5eqS6tXPZNoT/bTaX
d5vjt17YFAe7WZ06Iaqg4/OwkekOPuzeh6YBv47PmsmAc9kjkjSOtU4AIqcg0sk2P3eoDg1aNyRE
orLiWZ7hbNWG/dNZ0ji9YcEgdQykiu9WwTniB6mE4Zb3znrDdNJadQLWZ2Wu1tNmqFxFU2a3a/WG
NfZ7HU0yot/KyVxg2tiYfSgN0hpXc4zLiV7mHKBa7fxJyG3l7wJ4dorR63VAKjDio5aAwntQfvp/
10iFLNgecpu0YZJYBCT5dbR6UdwbRlCMhY8NUJ3uyO8mNge2PzQhpAnKNxEfV1j1uti8TFsVFQcQ
6z6e2viWmo3ZlHOxFFAevWFwENDfjXwQx3gUUJpNmqIIbgpYjXcLtd4cwy+go0XAo5zzungG+iVk
TadGacWPL08kcKWS5cWkSzCf6rRAncOzzI2L3v+MbjJaib9BJZY/nlmHCRUdtN4RVuSYMWzfruYh
U4prPjfjGgo6wQ1FWVHMBYN7tEX4xND81EmCKeowU6rDrV8ZmzwxzS50CStHCrcF00Ppti2EurZb
vgfWMy6acT4cc673Agwy0P64MXfMQyRIbxYUlTErmyHPu1bVSuAz7QqHxHpopbcn5q41HefLSWf6
sVnnBmaHjgqNNIGUspKBuMf0tqM+mEnSOKzaZb/2rH4kceSekb3Czl0szmt3RIACbBXrDAZ+GKDB
XuyyIxW7K9ETxAlXlibjwEssnD0X3a1Gb5jrRppGvx4nd7O7vmYyfSaAqKbEwJRoNipfj/EkJTM+
TvmwjvDWYk+0AfeU1aIPyiKD2VQOJ+8vOE0tDKdRYfYXfmxFoaKiyXqe0Y6tm4rG679FQt6psGZ8
IKI93+pmVrNxbMZVBbH6sTyCG5feWDeiVLC34SLogr87wiOy3uaGnl2i4PhInOwIaqOwLPZXyLA2
CnlCrJAXVBVvysnWvSykKss11SoRrwQ/J/DvLNxCnoe+WxjIPRo35sleVSa7fSZSCaxP+uXjvyjm
2vxgxZQo3ISdjPdZ4uE042VmQ+XaPo52jYo4bfEQV268GmkZNoL0xdQGYpAhOjZs0vJOmMFd/og3
e+PXuZjuswa5oKfblKs3miiBiSqFtniErn7q3WjrkUds2ufHDO5uzzYR3x5fmDFULvzW7guIdnK+
XhBwi6pv4lRdKyySfti3ysMIXZMnfz73HT5pkOAkPxvzl0VQaoejQTC2of5Lm25U3u0UJgwJQ6eX
pulKyHhL/8Pv796AmYYV1+GcFo/D4NfjwdGnCeznbZOViRlSiyamUTkEGeYgYuyHw793N4opdIkK
FmAFfLCIP5VyEzsHDwucZLqjfwbjZ47sChhWdPZB3QBiGpGIY1iwiKjt/bXxkKdyNxERDK51r7T5
sckdMEAU+1GMlJXSfPz1/wVUxMxInE4JDaTaTYi5GaV5ffv77A75EBNnr3bJbF3jfuO+F/99WojN
7ByNhy62vWPfT5t4BSM+aRb/B3KD3lZq+EUkwx3IvJp7Ij/2OJQkyq2pdNCIRHPJz9Ro9T75WC2O
alniokF+3GuZxzRSnPhJD8L642W2hLIJGLIYzZIaxuw18KStyUDOKNc7TqeIbH7ExDV3m8VCSaFd
ZA2seXOnjOEQ4Q+akWn7M9lQpQmHH95cw/RDBDEgb7Y/j2LZygVKq9u1l0MHSVV89mU/39WGU58b
5K1HjM3WCKvreXUjsADTp7DLMmrxD6oRc7Plzil/ONJKBlaq4qTNQdSk1DKPNAZZl1GoQbquGJed
uIT1wTjRCFTPQ/ddkWSf+t40TD5diCoahlHg68i/EbC+nm3cWusLRVFYAaNqbijV7thSO7wQ1umi
yn2gCTpcCgqwhB+axO6+Vl41kvXpFRJJadZ97rCCxvNu+fg5LTRp+rDNZnNbSUqV2G7Ug1nDBG+k
CsaOTly7b058YG7MFlZKp3b7C00NbSBq2m+C3J/k3MIKDEByqlNukTwcXBv9n+YjNYsEpvXeBrnM
8awLWCLUYjiBhRxp0Hsd9ARqTZMpr3kh81BUYDCwnFkd3yOYBSh7y8QYa587fQhPqtWmEHBKn8w8
wzShOmsWa4K2EM0/mzjjCtzwKmZqmxcy8CuSOBQw9VqjL/hXeRwuFmTxEl6OYice9xEj/yM2Um/q
PRpQadaFO3TOHcqDm1qpOPiKV4LnvcRQB8GQ6pWwWdbg6wic5jntF3Eam9FT/jkDmtPv0QXdO4w+
YXDi/jyA0rdSs2f1kUhnMpJ202cCPRlRVwWllQvikU9UTDE8IS/dx3HW8zdmOvFWgzsTPFu/1hmq
+VSO5ZE43QnBv4KIijkCgHNkMIGZ6uokJr6ZDnaRLGI/k8WBQ9EGB/eigiHC+uvbzLsIe8vW3XJD
jlBH7I8gqdOBNC2wMkXZWI6i7VC3TOmU7mqM5YShfhi8kYlzUPynNS9D5EjP5O5QtKOj3bG2qYw6
89qmP6kOd8yrZYPMLI9pJF2dXLRvI5l4+ABjWSotv9M0omDCdn/kuWLWlRkLMiM0lsnXJ288jl7M
yyJtR5BuT1CWRXLdgh6F8Uglx59BrJLfAbC9V3Vk5r/YUAtfL18a84EwrMHn02Aj8NIHVARhE09w
4RbLREaecfYG0x5SSLSTK4OEETLYsjVQpXV3YS76Ak3jylhV/WAlwZBBQdbWSz0LbDsFdjRElK66
dPRFgYfXz7bByiH+YvEKSo+U7lznh7khgnKuRfxcuoABxpQp3oXYwK4GluST0LoHubKf9wV8+qTK
E5i9yk3sVv5UY9B6l/a24sGja8pxxWcpwtASlXOQiRx4u5MYaulWBbdmK6OQFYTWMBzvq+j2cyB1
JmeErnudWSOeO5WQ7ahwiFpFVs4XWHcPRl5FWP4AH8dsl142Hk0mdHc4MKpruuOlqwin7Tm0kwyP
UqCltQYLuFLbL80o1umniBomS767rO56GfKdmmvC030q0AnhsmrM+ewI2EGJLfHBpWy+Bl+ytvDE
fW3AAeUJ6iGku24GRAMidyiOsl+lqkIUgWXVz8FddsLNJNwgBAR/vRJzbIFrIdWJjJ/GQpFFUmbp
Q9rL2R+IE3OixbhdkbUypmvg3pYdFQAaqHG2mKgLI2Prm8f7wYG6TfEI36uhdTSN1gHrYJ2i2sgB
qipRPOZEYVhmo/Mk77P6J6dbqf8cacIn/CSlk7Qw65r8mbpny6F5tjesRosmPTlqyF7JAwpfY0OW
mcsZLZ65O2DG7kbEnxKsC6VTiWhlFfk6CCinwFFLrb6aYnS3NbCqNMadfADaVnKFQVawqgCV/ySS
rzSrGWkx2vLEJry5KSW34+lNxGWourQYVM6k1fVs2fK7Tr5Gb5P3hnIDtPiq/fZiueN7OZpmVeLq
x/A9t7ciAQQNteAYibuLIfnRe3iA8dFWSUN3+bOZy0IbPgdjl8+T5+egrcJ3CNJCWfyJTSKD0LEb
45hG5U5KIy5YXMALOM+rPRE33AAWExdSYVXWlVL9OgsTpb/tUs4CPCoFWX/n3Zj6HbQRhDFC5lPS
ItrhOJVfIUWF/m9X2FjHQhoSe5Nyf6zVr2qUzHin9y3xRJbjWiSPvCvQ2IFLoYW8yp3quO2WxOfK
Pcu4I2trY2XRYtoezL+0vNGTUQgx09gUodCSGrn2uDqfiQGQkC81C8Kl4OP50DQ+shpU91BiQM7O
cRneiFkMSNimgZjWEbAJXUUPRyO4TUOFWCWTqLTDqs2PcTZibzU2cCflxrVPcYQ4BbFkBLbiYixr
uuUU41Wk60Q2T7Q4lmb+M3ae1xLKwD8erMc4cN1LXPny7dvhHDGA9wsoE1ZnVsJq7lcrwxmZ3r+o
dR2UnmW9M8zu1Gc5SeNLu5dXNSGdWLrD0ED2lcrMhw5rrUbHMWTLGNr4Ydw1OkPaHjQrw944ZP9+
bLhKzgwhwqBBc1vlMtwtVHl4/uu9uDh5pOSPmSXmcOnYdkU28OCRj5+NcNr6jT+hi+ptZJtdACTi
zzoAFr1V+eSqdw3+sjLJ8VivddDRTKMeC0SEXMNnr1rmTINZ43lxtWExohAxWfc5z0h3hoxgqLaH
Avex4wLSi04BQgPFy7gLcSFCvF+GlZZhsA92UrhbgJD/usYp60hiyZ8eMrVi945Iz86kT+UlBwpD
DvOqZVq/dj3atjyyf1dIh5mJbKZ0xyBTeuScuEN/Zehyw/GsxwV7RPMOXgdw7CQNFyzeN5WHg8mG
o+qOFDbbh1Rtg/b2aShJlpnig0ocu8N1E/yQYT8rQN4zSVF8URHVCX6FV6HCj0OFhNqVroebbOMM
r+17rrFhi0Sq+sgQzeXHdcpLl2I5kTaw3fspA52wlGmXFwdFM0X68Tomd+NVFPMtEYUtsY2LDcg5
cjKGEqbmRcsM8YQnhGaMGfBYNGCMqCIWKgL6sLY2cUynCYnPcGR/HewhBmZa98Ddd3wUPImlwTPA
QJinci45ND63k6uADWC8yf+hB/tMvTrhIKeKxq8LmbRwUnv7MK64ze9gFY01wE+ba6BxJDM2ppt6
sdrCwJyH9TpIR9082cEZPuVa0mhFOpwZ0uRdu+/XrS6HAF5jNv7astm2B8btSrwLs+GrHX/kccxX
8gK8/FuYsVS0k3eP/qAq1RDEV/fByFWEcr3c7VOFAXGTdjBOMS4K84Oc/w/Y6Sf46ARNKdHGSJBv
P0bRzxBBb3ksmeykl89KE6GZc/a0M5CQ9PNUbOBuR4KTRrx8PLGPuGuhV1A9KWbTPzwp0jilMJW3
YdKpY/zcz/SElgWehQIN5/6lvKBKFD7gth+fr5LidJ0dX3yqwEy/gtNyzRRybdq4GtvutcI9pVVb
IgpyIymUBhVzbZTHkCRiFgC5AxpQ81XVxcpr9RYQ77+hTlhShbRU1ONGlRYRrze8inhOJJz3yvE5
yml6usgOeYbRcp0Ts1Lqpfm2mLPYmfyseFZy6Io6t4GSMsRWPWDPzrp5/hq8c56s0GzoPeUJnQd8
pZekut3PQnUKjwMpR4cMEy9hMuQC3sbPHR0sglY+A0Ch5vMw89KC7vzNGnKNDJu2JtCuxKhfNNfm
aZlHwnSHo6rVQvuE5S3LVcMBXjyXAV6j4ztkQu28o8mHEDE4HEW56eNSXXX4fkGuvqSNmLj90eFY
VwgPV9CRxPZftzkbhfqsCpepDziuTme0Dy7Ma+wa/qgBHhUymEbep4V6eUSx1gSxmNn/4Dv9v70E
KXB5TdYvDZhPjbnMCAdUoJKjKNBQMvb2ywEKDvVgLRcV3FZou9pYj/v47bMCBEL7uyuVIE6zyNuU
SlC0VQpzbQQbvfB3J9R0w2d7IvkHybhofQwtoCECkpODsHPRhCu/jIuE81DncO34nrsu5Jsx4UPK
acSxd7DlLgOpHgiE5JYM8R/AtbQCXDPlyrm3Of+jE7nlPiVki8I6Ch6jYXdEOGFkOPrc6Z69Huc0
SszFcGkX9QPEWdqyzNpBXACM3bo73SqBGZCSSUpMAV/oJ1bxy7L7LxPRT6uNyBcmehdaDuwW4bbb
D6X0QNH+ig038eiV3UomnmuiHhWhT06dSjlx2k7eopZv7AZzq1o9dBfUGVs1odR1oprzGb5nSzWP
KPESeEyn91TWJRCKf3WnTGSY7YcfifYhprFwwLO77VL5ff4x+x+OGybCoHRQITCgxrUCQ/q+nu9A
uFqL8MP0/wWs/d5CH2RrXnKP7cmJxMINABeJYzakrRbloGAWM/WeuaCxzExjF7ZbAUPu7ADfBPBD
fRwLpCBhqYR1tGO17Msrkp1hTkqJ3qgMFiKF8BXaJnh9y5pBfQay07Jq71Mapk8bkBCmWnlR7zXZ
39uZTHdzGoMuMQJhebc9HdNMsbifKNg1MldmIBQndHelHogun+IV6ovds1xypyyuuZH2u8InPQf4
mpCKvuhn1ePnoiMF/1pC1t8tE2GPFyYTVXSC3tcYELhj1n+MVzrL+iVaxVtdb1XE3+7VIDL6JLI6
nznFMkVZLvW3ZkGH8phLBgeHoyTZl9WT6bU8dSmcZq41rPfUxFj5z5UHreh7lfEIEwVyelXM4cjn
j4J+HhEKmJowBcfaBIyHnyLDdDcWBW6WZ6PD8Y1cQ42KdNI/wdx/UVhQXt3ccO/QCztlqpTQSMPO
GyCxoKj47mrjfRSRP74e9axpxJS7jn+yNVwOY4ZMXK75PJc+DiLhNQqSHp9tfqgekLKZDqOSmHYl
Ibk4NeA2FuRkgo+uLiaAR7xCj+f283lIMWo8f2xqElK8G3NcKZWMumNBFSoPFt+yvgCvcLEhSWPm
V9A4VTB3taoYyQBKfC4eia3M7B/VJnFi4YJEGxI2w8PiSgOfWmSd4pCe90ZhnSfUYhNOa+kFm3IL
wpeylm1KSJhdTlCy4g4qEucg8yqDfq1GXr64IZRMPqTYmHh0NpXsiNT+UItrFaI1knnWsV3kOlxg
DCW3TfPV/BQdDGkiYcaXpz/S6VxI1XKWVuHGkJeEBeiZMGS9wOQ5TYENakENwMfYlghyAb8LvpXS
Laep3ZiZcOkMvlRBpPwIMfOOy0fgK7sS/1Eu6dM5xIq1mjQu4u13LdxHrAoP2FTChEjKfl/rCQBe
jaGJX7TrJIiJQpw6NYqr9ULnBhnc21jUR6w3mv8law2Ji01g34J7Nz4R9ZLjYONtvzRJv9ilH6Th
VAwIogji7uR4Jh6qTg/SOaKHPQEeCTmW9OJwq5SdbQkYxtc5T9oNb3X1pxfF0x6AkPnz+FgwRhZo
FqKKm8KIGUcrtgAMTA6Zywtge6pj6A0/HNq79D2pm6S4LhIeuDonqn0ALrgL5unYWMjQoe9AcC7R
pA6faeyRWyvbqGGPKUHB+bHR+naJIBJjAcXtivu4mqX7rAO7DOSOUfqUZmlBuTaH5wFUmZ39QfN6
oqS59E/JkQTyh/CrE/z9k3R42zs99rf+hf2QGwPZi8vBmb4ney6V4nKVpPCXoPSdM6hkA5URlOrl
Lzv6RRCHL+3infQEdPeTG1Nx4ck1yGoGYRVqyMtvQ7WhMAa7BBsjY/XebEHkuZoQkeQwFVaLvGhK
lgywwbjovGSq2BR3vh4M8SJ3ykg/qfShd+QIFUU7u+Y2Wl6LkUW71zxuBDHgim59Thb+jHa8KUQ+
cPZOISJ6Ks8I+ELy66lEL14Grbj2rHbtKukdQDQ7oOpBcWoNgwWN1s1cyFAhOFmD/XFO582R6AVH
pGpVMjsQXMn+Z7oSd+nxBUJ+yZO1Iw4yBag6mXPv/7BCShfn+gauH9J1rp02mzLP8vYIeVPdbmkv
+b5HCwGZPkgqXG7bsV/3KEKaLdBNyH9+iwrDVBUZNmOfhhMR5L/p9FRGletReSg/NtgqT7D4PFDk
TG8q+JX+5g+Ybf3wPYEEJ3eWs0/ITol++2hf1L7qqpxRPZY+nX+qNregIP+7XF2KYYdf2P+8TP2K
ohRSA3V9wODblVSF+b1o47UWId60n5IW5FWwP18ytfasHNPWZNw/bKnq0jcmlTzJt5epb1G79cs6
w7Kz75IY892YNcOn55QhguVVVMEs1YSQPmR52XkOHdbek4I1SLBvkviCzcRuVVSo24CKSzvZB5Rt
r3iSQqSuu8ZesPkWsdomfX7JcvTCTa4RosDmUlH5DUvaMrWagwJPn4GbAeAmrzJ9uSJtDiSGAL71
rXuKLZGFzzWH+/f3ij6n9yIhsbmhV3rapFDSugJgHIa7gbuZCHPC2N1bZNKw7ylM85JmeACQodXv
8CO4MxQ1fhCJ2phfyqYZtoj6Wy7WL9JM3wCM3AgJrLZhiPDXqKHnaTEdbi97yoLeUY6wOwVC1P5B
wZemc94UZ2GaHqwr24pJRgfSiE8UTcgqG1YK3aYQwFB5WTuL7z6+23cBWJ9YjQWLOaC4A9vteiux
X/utdpo7g/pZ+H3+Y7udVKCjJ00bE6DZqbfzXMJYosmhrdXMdaAfJi6gXFw8CVvoR/eLqxNieoLX
8VBgzbrJNgYA9VpBf+2OC0sa76X5+6C7eGyosTI+pffd0WkxsXFYjLy7ZsMr8/QT4vWVUFCZ9MUd
CsgtCKDa2DDYarEtq9WfRWsZonX1E8yB2TfprUTqTDQk+Y7VUktAgZw0XajPAzKfnOgz0izjQqYQ
mr0E8yLYMG+4UUqxEs7WqcWaWkYOkJqn7970ERtP7dhHhCoQAi9uXJjjrdkDQHt8pSoMzgvk3fDp
WrHThJrob+FU+rEKcUBLSpndv1qNgUmtFqvoCzv2L24MtUZTKqWJmvJAaV2tcEgwyWeBFcHHz71N
wbMTeUEP201uO+q2+9tpsI6hmTUzwdoB5wlTid9jm8xZ5/It1HAjsC+7CSv/wR36S637P/Ep5JtD
guSu9+KGTqoGZ2RKa5u/c1Pe1kNoeW/e87iMQZpDs6B4ioNW9v68hsDOuInsrIHvVJ3UR8URzUYf
Cxct/c3/5kW4JvN9936/UKTFy7j4NB+YIHMJyX6igiuS39qmNuZbsWHnKJALjMjYS/kLvICmI8L/
tUUy5rkKD8lWqR12knq477WK0KbhbWgAhMtRmGQ2bjl4fV0Pu69o3WWh4LuFbfXQxEh9ULY5sXjx
n/4slcQz0uWpOIyuQkx/MfDDjqtKgH+41HmTkVHMp3Rip30wv0Xx7LtkEWYGdgmzNevrpPLgLib4
8spK5r3TGE6X8rMPcB1IQ9Se3RlazRh5CpkWtFDWka8uP+z4I0XFCyh1QdkyyHBytcmYc3nIDT34
5T6E7bqMS6QpNrQQYwp+j3kcTN83ol2dNMrhDr4MDCd+EdrxdYXBe7rGIkBQXBuf4UjoBcM9hRgi
PbgY5QrA7xqOOLIxVlH4LCnjfh3lTtfiKV9im30nUlvIzyBHUC6VkpMiLk6+UjDkIMm27s/attLI
9myL9iF41OTOQeO8TI8Bjd/fBRz2BdeOqOWteXUtory4ZQFchnCnztKeIvuBiepO+mj20LMtAGBN
XClLM7OY+2S3CnPnjWQ2nKHfq3uEGPIVHVSBh0wRQuKd/KhDswwH34gRMBSEb7oKOhX9RbOEH9aL
iEckR1SAq7JuXlp+/IagdJUH55q9G+7GM5T/JaVxmXY+77ACFz2MmJ7Pq6Vq7QHGkM65qKXpUMsG
dcx+CGIhwOTptv/8ZRoslosywQcwa6ED83MhPS4b0+IO8LCozobQz31toUzrO/Frm4jdpySHRh9k
h74CyhnpnM/JjncebltVn0nww7Jbl/oshd5UDoSpw/KV0rg98uHp9k6RvmAtbOYf62e9tK0F0/NE
6PRMeOTlysVDIHn8N05geYoIbj7ea1dxYmkxIXh5no/Tvzq9A9R0uz5H6sb+s5bMGH3e/LfBN9bB
G/oSh5Vd1bMlMxTtyvB7uDM75MhRJxLX6RRsXOX+3zcaCRGW/ReYF6Bkf0kskRvKt9JxTpqUvqRX
9hvna5+Nt1Id+PCt2wnqU1HbZPZIKGNGv43jAHgdVyjSf1mvZtejFz8g6sQpE/5acEobH0JdU6d2
3Ca4rIEcMNtqLgIpsrXKGItomBSUn/M55efsf9wQtcP96BPNkRtx4qQ/zPPW+b+y2qpNyUHlMlK7
IsYjlgvJNKO6O6EePYLqACwanTMDqW3mH4+xOim4eHL276+EMqBrwYZ8LKIjZidURbX6pBUew851
25rZ5F5Vu+WxjpvnAs7PhNKlz+yFPaGs6aJnQPhfDt7Fl502KuMAci3pSzSrBJ0YYJRz2am6R6Kg
lWCyFqrVfPe8WVDa6E6BtzJ4wKQ9q2VyOdyFC4e/LlyP1WbwXcuASO97AdolHjg8w5EC8oDOiRzj
DznOEanrr6saMX9nQXHlaCkt9ndPqQOpGh/JdrAQoXwc5JQ7IHffnV+/QRB11S4mpXmaTPuWgXYC
v7lidMpF62RH9aKGGKo1NdGgVplXakE4Rr6cWfZLPa2OcI+6mSEg8mo0NsonDsqvaVA6MSES87mY
DXLiHphDRdRuEYn1ty4z+v6Q3VhHklqMmg06CCL9IWG6KIxm0/RtCi1WfzWqbTF6TNNgEfZJAVv8
3HvnddpwajNJrfB9Z820esDpvbJpria8CQGCM2ABFfJ/WGZ1C/7+5Y4/JM6JJbYUZyF5VsNZhvru
TLTVvcBUf6xRdyKxGyQjIyuHMhYA8RwVhmXbxd7BP4dmSiYkQk8+47UkHBsWWjH9L4/3FAJh3ORb
hGZbmAa61DH1LaumgTIuLv1RQE4DbHYl6Ig/xwhrqYWNgBEQPWExRJk9ccT8EvPiQ6G4kGsU3GEZ
oo9x+2A818IL444B7x5ZJNEfr+3KDqq0/9OhzmGC3/uizCKfLj/Er6xHAojFDV7yjZ+Xs16GhPcq
5ewkpVJCSFHYQ4Tpu95nKBIcNrwTZNPv24dLxgc2Y/uBf5cFt8j7jNhTlQjDZQ9kOZ2QPm1rsrPB
7htrYdk+JqXdh/L2LuuKR5GWiHIaULRK5KzAIQ3Bdh3lOGvqqDAlc/CzHDPDCPl1VxzR4OHFmQR4
fZXqnqAWPOGBtJZKj752EdokN1S64fLTq05l0DAK+cmxt6FXZRJ2+10MaoXqhqCQvmrKMu1GLvgR
IMj4y/uKxPrteUHNHDb5dwupS93pm1modZD0HuKRCrJh7zQLxuiSwydn705tPuhqGvkfY4czYOOj
5zqjwxideSx1Lev5XEuEduxDuIhj0Gi0BYjT0QLeXMKiLZUlFEOz4ab0zkz6/QlJrKb+PhH6MPig
vCa1Y0oRSQudDn7i+oVpXDGCGQxT0EHFxZbYJRqqyQPYn4TTPs6dDKo5Z7ddaiboswehY2wcg723
5fYogRv8Pw0Aj81mQHpIHwXkHNIhHU/pAJ0/NwRL7NR+FVrw0dG3OmwCjZ2YihLPGvAuYJ/sBrgu
in3iR8wXMsRPTDDL/dpXvVcpzl2XFyDPZseLviLQUi1QXGW8pivrTDNtFHLjCmsudHKl0U1tSdx7
HRc9Xgd9n6jouZLXMt8kqBFFWOZu+s/37Dbj/0wab/ilE/oIrEnhTONBAs+uCVAQRIH6fszzUnrJ
cQ/j4pjljK09vAPNow6S0/Vox3Qrk19heehtVqvSykcRl6bgaJkaF8kpT0sow2DEvm2Xzx2uYtK0
rlBKpWbYaqNeT4m2SU/hL7u1FK12OONsC6T7vfdZMyWTLrULFc5RUH8wxprQx7T5TSr+H7uXe/uY
O0f6ufYf3YucvjLVbyxtuNNaLCp9NeKbkJ7B1KRv87DtWM1QqjodPU/vvOj9trr3ZmiVIm/ASOwn
3mruglGcxBwZk16a0amNJzWJg1TJU0bp+YWWvg7WaiH5iytui8ympMXs11O27XapQ10sNWP0Otn1
xQ91RwGql0dmQqdkfW7h5AJOvdtUsGAU86kR7LJwfX03/d+sYVOSjXjQZmM4OG3SnaINGylMU+iX
wpZNyM6ILm86JC7gwSS5LDAdEuOTDCrkczKa+137NesQCW26Q9k2ALtk0Ajt9Vn18ZSLrmFi2im6
frr8UdS8p25G+E9iCcJSSF8q3UDiiALGIjUMPrQhesJxfnBtRl/OwH9+ZHEYcrr59me91yKNuL15
/As9niMyQkLBV1IyGZPW48T2dc9W3L1jSC10d0fhbDzuOn+BnLEWrlHDskZ0xoWNquHdSgjPpuui
w+GZAkt921rn8hyFD53FMWFXFPnpWbJFQS3TvPWvoqvrxDwCag9cGlqf/p29TF2izWC7ljZWn7sD
bT8LtyBrwqCYL6R31UHdVve66sAh7eFUYW4zwpe6jTI6oX4xHh6J1jpWvXhkZghYoieVwXVvghgR
WKuRfzVz10ho4d4kJ+TZILUj85d1K6YFK487NneTRHe5S6lSFH4tV/opD+4PGx/iOodQyvJA08iL
L6A6hteo/MFqe6OUVpCsRh0DPDW4oVn4RT7mwDx+1wUpDH1HoRFITVijrznOjbbKBiBdmoQFbFSA
FhX3g4LRf/8RKEokNI7PkjYcWIbNEh15AuKCBKE3bQfDwjIn3mrTzFldXKds1+bPN7l6YVyqU4Wd
XjAhATVYmxvKUYLkj/QhrokilUl2Dzdgug6NHlb5lOaAfS0Ylr8VRMD9RXKIoqL9GwcePNmbOFvN
fbnfmzx7zAL2zwRH0+fPWF1v86IejcwFEClf8nImpwzatodwbxYrEhoeVLuUO4ygQ8UDY05S9+Fo
kAA5P0fy47CDf/v+9jfHN4t5pu4GY2IF3DtqNt1yPJM4z9NHqUGmDbKqYd2DkTMhhkntBqfw5e0I
Dtsh79slrLCK1Ymu0/Y+pToJgIMoiYu2thQyK0qD5fB0PfkGl4rTL/iC2u0Cs8bzll80+pllu1uS
Rp5Qj4E4tIS41ikRN1uAp/4LzZGrfU/YnkVWQxA17CTyXFsfB9jTkpPPSvqSraVL6UImU/Jb9Btc
JRAjHxpWjM6qkFIjj9J6H8rBA9XkdWfSwsN+X0uJX6kZPkDk4jvrIpnrjpAGZvTxiwoXpHHOvRpz
oG6k9M0bN62dFZnCqfmDAiRdL2KtWNRDDACDFOr0QbxIlvneghMlL5X6S1YyxQ2T8oEC5uYGnk0E
+UUK8xDHbK1rx9Js1WFubAYIF1l4gQolXS/4Mc8mvj3+BAi9uD0KaWrqOJ5137zQOz5l03/+VwpF
/udDQBvBWbofDg0vr8LrPCPj6JQuwmVmcMvqIBQMe1ARBwyG8y2CTKaKgJCWVoNGnMWwFA9gs128
iV1atCX/FAlth2E3BfLimqApjTfIIrHvTyUF1hRKArAHjwR5pQWu+AOurDuBjyeTae2rYYKDnOSk
EY8+8/Fq6mqh2I9qeMz2pQ4FJxpWelSmcobzHk+ud8GIf3DYRHvp6OFf4GEuwryK3uw56IhfX7Bl
hNHwyBHcVub+43ac0Be+aObhCpQyZQ5NnvhTwMAxY9lejFFrt+PDVTv6CQqw0V20I3pNdNE8WBkb
HEi034soubkhxpzZf65AYX2XCbkraNbwI1tyMTKn6whzWgwmpjcgjk2+1ZkBdHCslmvQp0I5yvQb
`protect end_protected
