-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
A5JHqw0hKhjbt6iGZHdn6DR5AatxvtXgamKlukWHz2ns6t5BOP2vUcwZvXsUm3mdkfM8/2Re/00L
CJPZNhQbMadx+o1lRvE6ELoQudBOUDIy0JtKfgWsOi+K7M1ufXg7dDZVoA/CuFPtAAFMHpMbhk53
Z6V8WgjftH6GMeudJXcbhIDfzNrljyO6ebarEQ7+WbxphKysx4qAHlGMZT4KlhwCcZMHvRbCgsi7
k3mW3+q11UL6yTzvynWuO5Nu61VStMdRYlcNjYu4Lg6x0RiOEcsLhTthQvyhQ6HGd+WryTodceJi
kC1Y051I++jo0PWdpk+pAPv5aK7Y4NVvccPTuw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 35728)
`protect data_block
i2hYt/XjJBieaTuJh6qmyUkXk0JEy40SC2Vu9Vh6sWJo4L6LN7u8pCgKch6WnXnp7lpC1fi9VH1+
ZzuiYn2QmWeMgy+mJ3Sl7JYTLQwKjZomktwBrRa5TNSSWibNAACAQFT7BWuMUf6I2lYRaaZQxlO3
x5DkIMNXzUCZXAF+XlMOxnoxbIUC8czM+2bTNTTVMNeVwWctgpubTMzLLu8wgvhYrIy4p+OLmfXw
rvjbQjDqkvYmCTY5MLik65Axp6SfrQ4jluQWKKXcrrxbb9CDnFKwQ9QLYJ7WCIXjVwxZgaTlvDRk
Imqkd+iR50nXMIJ+2qFZ+K8Tpzh5/XYZc8BB413yHJKeTKsMCng3ZxvXCKrJxn6fDQldKsiSvS//
QLcrXu1rC+OrNpQMLggvK7/8aaUtFk8uWOVQvaMThPmcUUjmXGanwATdxFwLpMFS5+XTloLLqBjq
T7gaZWRfbfHYY4ITW1iP/tKCuge6tL9/SkqYm3GNjmqDLcaLKR9yEBt3oPbp4Wklhqv0H0V7/yVn
33c7ZRJgiM991ZFnhHG5er7z3CIMgQLUm8nDdyjwEPSH+BenK4PcKocSzIkByeYcTcc09sw+f2WG
QAiDoqltI+OHcOzprnnMNazpDSgljFFljK7Q0HpkAQNdzF3QxGFuE3WnpjLNZZ3B+kMmxXi1fOU0
ZW3hXEeW5gUkc4koZsVk27RLsTp9eqF8oC2hzFcGJcQUgBfEEXot5uF0zXr+KchNvt4BNKHD+rgL
IMUfaABEsC8F5FXNuCQC6HfGERYaa6+8hWs2sAl3hObLHvki1nLeNaj84SILiNUeM4DQDa3RLTFw
2xLQV4nqmEA5vsHbPAqlk6MGheVnFRY9CDhk/7J1g9GFm/ezg3xnESxGUVPNWz59Mf+cmXqLyP9D
MjS3Ud/HFmE3MJ8pWlqsqoL3zfdyxRPLhbsrjYiuq/Pf3dVx4BJECv1S7dxHcahHgRzXEg8qwkHU
KzKEtkaXesCXi6jk4VndGNSeu5kPbEhEOhkGfGD1NjUwzX752UiY/6RoYEKm5UySRCQZvrNT6FoH
Mr1dIyYuF8EKwHLOFqKBF08QxYcHIzR4jupKN3jNZuvvAuYdubfdA3qbJJlMi+hVJyAU2tmTx+EO
g9udmF1LVhYHRT23DIDPDzWY8NeRD4DzM1rE0PMdhSdInkK8tBP/4ZoeJ9KDKsSvrY4Mic64iI8X
1ml7nPuBnWQL9/7IOeGPMD1/fMVkuuWFr+ISTGNWH24RwRgP0RpUDegF7WZUymviLAo+ZWsAB/lR
TqlJJQUnURHbGCv/Xi8AWyJBedXfeCFyKNLzWAhLOZ/5DN2ZaQUjlq/8vk4BpRl2xvtW2O13FKTu
US82heXKEGvEoHObsPbv6L+wkLi8TQtSh3ITlS/JRFbkVLLdVhtkkCN29vp1jU6nL49sqcrx1R3T
u8g3zFNI99jz2iQ7pUYgHRn0iHMFL79V3vzLCwGKe6sPMUdnTgmECKtTgjgWdo7w8wAIXjtYsGZP
VkIf6qGOSPbsfWvZ4zo30U+6wdLB3cIdkWBpsoF7Wm3xMCcq/fGsWQNDdBbzZ1oKJ+NuH2zd+ZIP
hXU4FL7TkszOsSW8lYEQFfUzuNF78GBjf+M349zgyZq6qvRxvFoZi0hHy3YGMlIfTCwENvgwM8gj
sGZ7l2ZTj/zDo9RJEaY8KhZNW1paD2I8ITrypgwGiy0+o26bII0QTV/5Uy1dcr/lilOgMJaUOYGW
/R1E1nuuvn7OsRqiNjKwN0xd1GlXcmUB9pkDOMLy6Zw8rPok9ouV93fem0t/QVVJiCQtzJrjp1p8
U7KtQyEnk2pmSKdIQbN+lINMXH3f1wN3UPL8nSWOPwMLLBMYpi2dLj8/nUOa1hjn0qrSvys+Vix3
x+c27iaFt81zK+sBWMFUaHo5ISZZ2NtdhgziPhN95WMPzEzKT7dHfTJIqGx8CYrG7VJ8jgpxnnkV
QrlPUPEqlyQPGeQgQg3hXlCsF+J4+sPrcKGyRL1TXbnQpJbCzsQUYzlZzmpOpJ0wteqQNFdSqTOd
HBvLjFBIxspO1gHxvaa3XvUy2smYK+7r+s6PzMOR+FfbPVPJ8efSQXuIlEVUIOT7RV5cCoJCQ31/
BplL8GOgxJQYA0DB1aewE64SAjE/t/fK6VqHnilXMvI5YBTkzLJgYPBeUTDftO3ikzFZ9yzykSZ8
1z8iWGYRUrJTMiUcktqmuAHYo2Zfm0VQxCf08/Vr06M+U6Q9Or5EhMfMcH+cEFn75ybQqYAbT2t1
6Hoz/ccQw33z6ryB+gOeU6EzPXoPGCCJIlcC1IgIh/njFn0+pbkTnaotX0nJQ2SRfHttmROfL3Gv
tVwS58IUhFiOWhBu1eqqpcchXDVHp20YK8PDn0CBeBxZF95u9zP6DqZfNKeTeLSOdyADKUCOcGok
jkacBjJBUCrT+KtK+pKgr4pQpA+mo4qk7dwHXTi7SeMi/lU//7vsfnjjg4WrReV19cZx5LAQ+HPT
aYS0UaMVtjAbIHIr/7EwStNF4r1cP4TvcvXx10kMJqPnTAH074KeweAbb0MqLBjfPySiAmTszei3
WGO6uCHP8ZnFltBe46q5QtIlcKkNfPkGTrbO0hGCe7rUg/akJlsro3GUK/AQOxGZFbhBDYqRJQn5
ekRtXzRKdYdC8m86p3rIuEmZ0hRQSLH8ISII6Hd9P5b6Cm/kgIexV6Rxf8xKcbYV369tp1FGZl09
r9SKzGfZT/RWzo8H4lXo1NkKU24jQG61IMsg+RqlUJcAUnvdfcRr353WV091KjNOPQp7vQXZ2nE8
M9THTrAqsmaGHqUap48iuZY83A7bUkvtaiM1aCgQYdBjhEgxeyhVMFnd8sNpFzoh4TgIgiw6nBWj
sc8DIgcJPz7WoCBQPeczhFSWIcc6rcWhFqyQpnyFtReBS8YEfUgInZKo4HmafirTdQ1dq3d7ndBz
ppEd/T8XbnA4nFiQxnc99bwJRh+NPkzCwK4VDR6ANKD/rF83RlfZKiUsoDTCvlrPswL4I5o8CERn
zHzSBXTiinJWZ/bRu61ZBmcijgnhKXUvIl+tzfu6UtaJolWzb0scFTUj4CUNYPpfAH8VExvBfATI
6eb/o+nRp3vZnv5y5DkD16Ld/KREEn5xXsop6FO/afBgI4Doi3c9OoArha1Oy9Q6SxMbDu1kEHP+
osyCn36VayBADPikKe/CCtiLAQ1cPBeArCx1y+PmulIdL627po/OCLKRE/VawcxrDNOTSfppn4p5
9pf4yYQIMIN9z9vMqKaZpHbJ5F5pfowwdOQmJZ0aIOhv3q856g2Y5/SZKtjhnTAgFJ597Isl3wez
CXIWDsGTxPyyNtLHvjsUwTW1n89cd1LU8XfT+OJsw4Gp0eQ2oSmGpZigO1kq9Y9AQHvwZc9Dq0EY
2Hcs6uTZO+P/P645/XztOdVAoF2cquTsvqvZg5HQWUDNlBrMAO6jan//LsmAR4p2h4cuRkg/A8Iy
B2Nv4rTtG8o+2rVkCQbG0AWnrBbw0uZnkNWV7RM/T7sJeIwg2ewwhdXFlInw/Tn4otX4XhML9OYY
9WHMD0CUmUj+Aj2429TzdHuVM5BQ0V1bl4EFSKvG/J4NRWksUmndsBTpCNxx2yATlQHlUXZSTyRB
GHNqahWn069hVVMZ7yAkGay2B61FbA1bVo//utYO+KRaQ5WvQIjbehaGuGBsv9rp+ZUzy3KnzHgb
/oINlTRlklLKIaDxADrkh4XLPJ8ByWLuCZbUHA/b0McmbzpLWhLbnmsiMf0+pJDUEAStMCH/3301
18tElKurEcNTEC5Pnn4W/I5WGJw+SEpZEJqwFohDLVKzk+8PX78CPDWcu2CRpCkf0OPoeWw+xv8f
LDr2csx+VVRtKGeSIlmqjsJx7MDpKWnce2ukdEJeRHHgAHCACl/cbbW85KCnA2nu60eJk9FEvn0J
4L8Ees2sFMier6xRiQu4lq4SaCecfLC6AtPrmqhrrF9FW7iJGAGoK+QxOdNsGY59Hf9Qyk1VvyK9
5PcSd0KkunYncxm0u1+9jVai9Zwq4MXEuoe6PkcB4tNNxFl8pKNXuAt97KG1JyM/kRbbqhUwJKkN
2a04XnSoNo2jPbMyS55e5vdjEo8taMOcZMBPF6JIbTi58XecT+y//m/UCuSKuXxIPqKGMbFKsIp3
EuO00Sxj2oLNRWQU2XZw4ckoXgnrVVqvwtN7guLaAzeTMhLdB/4hhVKJXud4ttJN073MCcqz5ecc
BcRyXTroXeIV4Y4zU4bRX8XRdAha+cGglpsMppsNsuM9AHinAd859dmuQx9zN1FJsDb1OM3rGXnf
gL7vALJ0dfNQVjT17n/rC+hA3EOM8e+V4pHlonFO/0IOB0YQD1h2mrHstOjwiHJwkvpBpOIFkvv1
QSaG45dpBJQQueMaY/2zd8PH4kt3FtPjrCgGG5VrocrkJtQmCmxW7PxOPv7FMa1Cxnl+mG2VjTwK
KQoL0JnLViz5I26I1QRzOTnw8q/Egyt6qp5FsjsSAYk8vGfXhzYPBqwYN1gfcM1W9ZPy5cLyL95o
0xKGCptobUaed6nCrwaaXZ82x9guKpzCN+ULnfjZjDeDfpsbeiNq0K9z1UAaVPg5GXOczL8Zx+Ki
+LumNnMne2ZxTADxbpHUtJ9YQiYv4bT8AvT4Ug2s9/iQcq5AmAb4qH3m2QqLRORd0CNMMKycg8Pe
y9JbivgYZwEkCl+/4SXyKoHSxRQDB8OBTp+Yl7DbElso2GrEFbPqko13uLvFKaYKCOmejrAAEF6u
R610FGc1mWGi+DXrNIU5/peJ4M6EJBp3Ux8XGSY7bErLsuq3nMNgKSpPqLZmpBFp2S+j3n4FRrsO
z81uzhAGxTRCnzRFyEjKLNTah2S91m9B3NnV6zGEIUJ9+v7j3TzPAVBIdHKYn3DUE7Ma2s4ec/Ju
s+Si8PmiQH8IRogw4kf4b43IgH71WHIC0LfUzFxha7WrhOsGhSEslDyNBtiTXJzsmW1M/XznapFv
bZSpgBrpSybSew5Q+Y0gWmoByY0cdS4hA4lQuJSPsHNSODhqwmkYxeiHtcxRrWebMIECNdiIMm8Q
gRb6yVPLne8F3Lf1gzq5dfcHYtRL5RYf3/zaueIQXMQhzg1D7EsK4dVnZp/tojV8xPXQAdsZOZMs
3cEmF63ykJH7Z56H1P0X5tI0nZEI5YyeS8cDha2yPvzG2oDIZ434ZMWeuBWhjC1p84y5rP6RuQ8E
tjnwqLQuM7G/rcxTetvSyZd9WuKjz/03NsFTkt7rSH7pFn53+GTo7h2h8N6Y/n79kS1OVKk2+k6E
WOEwWrCyP5xgwGzCMEelUb6VjJfNVgWVdvFnWlGM7oN4OEKqg82B/fm3sVcb4yPJnnzzPOVeo8Sg
UdZqsHcZ9kq/GeT8W2XW/AIbtzbBWAYOwrCPeHK1vXPr7hOfIRovKkJ2aCkHDPT+wqCVb8qrZ9xp
U7W9xszSOfME+5TT7dFhfBexJSkxNvair4yFFaB2R64SxCkAQM+AyxWHaJiYJ+arZVENjfiK1Rm/
xlRmngN2Hk4PucSj6hlXYkIlb7KVxc1P/mCo+G33j/KbNjwIQ6QdLnIISKHl+jL8nI3PCIlTg99c
FRkfkSAgVEpTzrqMVLT1Sw5L9AYix1KLJqW0X32RP9BihIo6aNnRdPsJqiecuPUwQPHGIag5a/Pz
GlxPeROKGlpICtwaBnzLq1bsls4j/wOX4SvqpxFeeL/0J8BIJeDptVydf9f5YMNtKuxxn1KYrVpO
76U4ZzG1me7NG9bH7DCvWbpxPGwX19eEveWBu3D8Hng2W58pnxpokWWSH4QhhyTv/xI+eA7RH2q4
w5ERU4hz2oPuflk5b3INAjIccuTMyAWsAsddHUowfDAXw3zSmahhl7TCtL6A/rZIHpzkNgbldO2N
JwsTat8z9EkrC+gt9hqhoRemZinBjjsEaxnqxT9MCbD6+9l4U2L/vRk+AMDPGo1E/ffhDc43CY/M
kYSLe9s7EyqQw/+67SDLUQoB1v+YT9XutPyDviVLoCLZFcNUBrr018uCqhTawMKQ5i3F+ePvp7+b
NLf9eBrfxcYyRymbl+6b193265gV+qD6QlPFPzFAo6g7PPed6biGxHoybR9z6I0CuHou0Gr3qH+3
x30KKA0hif7eToQz0kr6nsFvr0Zz0CTvxsBb8GO0VzT9fPq772YtARj87wVf+ng5vueJ8VOQnH0x
kPaJNGXAm4rUXnVGfm6v3vnLzoYZCQhoX0SD9lNsmJoOwln74K0v17r2cU0h2R4Lbf5FmY+sd0OJ
lpDsvj+CGmLM4p1aXn0L++HaUJiuulZAmRM2aV5JBQqZZqkoe3ZsWQdJ1SI47bAzN0vpuxJfGQMC
jki5yXdy/FOn47ThjE03hcTEd65POZLru4RwfG7xSIGmDqZjqahBbKB4qBBoiFMGR74dL1Lr2cO4
/7ugYm8DaPaKXI+fpS/yRIf4N6DhNlgs1dUXWClwChFtV3ALfaXN8L4ZTbeBY9e05ai9ByNeDEtA
pXBOxi7aHXKhSN5rQrI2apGBolb7jl8oGjrBMHLol3R9k/Ub3/w90QadbKprlOY80xKol8oWCBb9
UjC9WLgKhDbUATBNHgBP1NxNoLF2vhmmDmJRtIUqZhe9sR/Kin+4UoFVHvCDMp/I/LrccVcnLtxn
Kevf2o7h7uh+w4QLBqmSvm++y27nsaxO9LCldeKJR6ixTr93Ef+uG8HIT6lh3nnaEfOUdpQKFkIg
AU7wN3VidzWUnmD5CvSmNEuO/OyUOrvoTE8mKhEL/Qj905XkoRFspjN5RNy+Ws7kvv3XSmyCRRm6
ouzeJdbgYQ8HbrPruLfmjK4Gz1C8lDtc70XXhfm0D4i9dgpbAOxKHVY6mvaQZHiu3bXExvAmRgE3
U0FpiSm5Q8Q1usVBv0STHvrzEoP2JcgN3gj6iXWooajA9m+xkVmdq09Jokjwkl3GikwGTZXrmc3e
+zaKp+gTu9ZyxxO2HyNXY3zGS9KWwr2WA4bWisgOCdTsgRLqWEGyA6UsOCr3cAls9vjiGJgkXh3J
c9ryNwWWvR31wUg9+Jbsn9hsYbedWphfWPa8c6e1Xibn/yiDSinEvMnr+o7avRG7XHjsNBL4pUOX
JNEuTq6TkclFgnu/3JpX1VbIgWURRvfaHTV5kawNR7d6EQYryAGa5+lTQqRvbV7hSSDmRTtzeZHU
ggIg5rvNtcOgq1hgBgk7oEYByk+Zb/Tw1pYaMAiBKUfugJ7IVD4pG04lyLY1FPuhJL98ytu7+8Hu
Iu1TiPmw5dQsrCxIazoueDlxYYalo2fmxh0bSa34yydSVqidM0A+qrsjRYPM0GbECnDpOlNrsoAd
BBJ37BIwWIkbF7EcL4zlq0VjUIa7tQjjZR7+1JB2SMpB8wh7/0cN0WfvQ4icTCQnxZBpjp1zpoDc
7c5BFgdEr0qYogePQJFYHzknmFGkehU+kok7EzQsZPGI750/jixxwd2WfoHkZrdNyOjoHKQ7Ea+I
oLtCcTdPdmFYzgrQ6pAxSWjj3hdHJDy4TacdpewA7JlWkqh7CHit4m9GuPd+txYJTR/3vUzrG2Aq
CkZ1oLHpGpjkBVxYnLjiLZtxROKBdl5sn4HHe7JPF7VX2Nkk1EkQsdGs25hJ1d0bDNeDevTTbtUf
YlXGvQhUq83ODT2RiKBD5jXUTG+KcjIhP/uedMepiD3zm/RvI6m6XexV2sMCG0cJlhqcf42iJ0kW
17nzYZS6CzWQwhjKp7RBFvchw+DhhS9jNHYQPd100iTZtoSKRLcKGMHpHg2mobn0fcUKh9z6J0em
rby0AMGVW/3C/+aZtp2m8bed1RbILC7uPiLDFYlQCrju023LJ/KtngZGITW0dnDM+1rs3XYFvYJq
Y5QzlNnjOz711E6eQSZU6jDfNL48MziLtGkze8bAGmrOfqjSBOzrH/jeXUKCZImUe9wcxa6kHy1/
MvNxT1e2rMMIi8ygDYPvhuCMvlM4HlnPqEZmkAa1+BHnxDTQEt+0K+Kn5/HIEhjpCg6rMWnEWLQC
WCMH+JrjWOX0gDxDK8NVhBf+12weIoBe5IXH7w1y/zS1PYhCR5fVIofoSMNC5QIv4krsBbIp2Y8T
YvCMR5pXzjzPipBnnfDSAvLAwdb6nHTzgZjOiryQbBQ958IbCBrBHiuJoaycLqOLOPF2Ss3ckYtp
Cr0oOfydn/yDM8lH7zcwEEdvOmwzU+UcN/7eYqXffPrDp2B3/nF/TdZ5b0okeuzD0UcHFuEnYKgY
Gp5DyWhqrh3T3K5eqylfzn2BZ0dxtQNnUZyPYO40GVrml1+kSE8jM2C8+Rlr2uzp1hC0gswlkT9Q
QLDOHoRDJxT3S2XU/IYvVIXPq0KyFhwnJWYEkxogRm9pJdocxluJOBffWonYUIsMIzdX7H3qMmKd
IZzYASotEVYk/NuAPOcE5e5nOWHYdbymtleL3DJxicQ3YstWfOEvP0LW1tAmjiDWwNi0ABUHpF9q
3XlTPJLsM0I2ePerkVAxihfYM7k1PT4j05qz741V135Xy+Rygo8tw511v1VhEL4WBKccLdnbOdVk
+DZS5gciDaDh6VKk3bUBke6IuzHXAXT+eOCTWsC3FdJCp0pjycAs8uFZEkYLgKPL14aPEC7f6QL3
D3i3L0BDRS6TJbuLkety7ibp+3f0s1utH+quF4CCCpzur7fwsdQ9DtGs44yaaZuUDMmz09ac0gyc
VcgBHPOt7lBBxG+U/HQRbOEYXkQsGSaGU3+/Ps2X5D4DWJGpmwAWQRKVEQ6mRpAGNdsD5y7JThHe
mbO2FewtfvvCTpgp+nnsLXxhkRQIQzJLwZSKRWqwYT1MSIlAmptJd+CXJ0OGOIi59o21SLF+9VHm
3uqAdxlJvVxix6wIr6fqZOCLIoe4/nODxL3G8eDG95YgfEq30mzLomIQ2kE4FBZs0d/BS8D9wrRX
J1OX3s9yAO7AmRxgLl8lu1PZxLoRFPDLIZ+epI2hOOMEUl2uKU0Psv8tFALtwtjK8Zoj6A+kn6Sa
QO9J5NDftc85Pg/QyPvTCNAGPOmmlHUbfcEv01RLEYYrrqiMT9aCmrqV1MMqnH7b5//6z1SuMP1c
EsTCiy3EMft8ppNqToGzKxL/L+mmFlnjNwGHdbHIXQ8KJVo0HnPjWavoWXt/w127aN5KXbi18ulS
DLkeiAr9c1x1m17zaF6mDhzsveZIEqHwNW1UtuGsk3yPE2WEYE+z7U487pdlfL/PLWSyEouns4fe
WpgCTWcw5FN+RDp2HJ/3f4xnRr1kH32O0YjGfS/z1pZjSE4hmfbTbwj88fMB5z32aIEVms06XfC2
3foOhmHlpYLpH8qRF8dxcsezPk/Vs7zzzsiXe75l9ogN2KSHzXiDb4RMBTglDhh1mDk1nBizj54K
Oq8HWPasUiyvqujnR7uq3oWOH11HIYlJ+giKqTjvHCylQK3PWaZ3PKTqDCbcu2E7CZwfajiojtHr
/O7kiwuo2DaMR1lW0prTGjXVO1zNdo3WUcms7KztNc0ekqtcEhfZcg0pzE/YNdoYp9ICSRn56jS9
cf8nRXbSuyspdAZymEU+7WHPA4HXlBPCsLNZv1t4jqzRCFvhO3/nL8GVH8OSIirS3g3XjdstEe0m
HUWW8uw+uy77T9GdV7wA+DA4+oLxVMNEiE1f3QY8tuMSOsEEQrsnvcUOLQTM6nl1y7sWLwl0QsKu
MHb20K3cvlA7ZAOgY4AlAzgVC5TTFe+QKZJdxtxirHEtverOiE00f7osrFXLhhEBbPNBqpdE1Gwx
v6WT4aUB/jddCIz2/HlBuppq04seP0eWojkbMDoct/Vj05XPc+swcjEojsdIutu6Kl5KiAN3PG5l
RfUrwfXkl9k0wtu2Fy/JfuqEtx1tZR3LUDv3nhR6Dx3md77zyfOuedkixdv4mLBn2Kq8Byw9eTdA
Y1ziNWp33DAKzp8DOHRhfdSurEcLwYKO6giJ3CiENRXU0ZCcEovV02DLfmxFAkSLj6SEHaCBS2/8
4YfI02lOotrn/rRDvYTS5PxN3YjkCP/5YhUsQnIiqofU4kMn6kEUwITVKLzaZq6UK7cv6PsIHbme
t/ff6Ji1bRho3q2mmM9Ok0Lo4jn4+l7qdFkU24pKiK4kVv6pwpayi4eT9bDqBtX8GuE+BzLYhJxw
ScvIL3aoWN8dg7sAQri68Qx0l+cKrM6fmNVDuAvUnBlHODbOsdnIIvhFEKGhN1rCPtpdXoYS6RI7
qNwolex+pL8TUNtf+k5uHB/qeCrBv3nsS/THNsBY6WwElVt7aBL70ppEC33bC0jbYlLecUdzNjY9
yov0qnThKSgevmnQ7mJHcz/C/SfHuIkRBJuX6y1uhM8PD2mFfSniH1kbTMveSh7W7k6VSeIY+KqP
WCqJmoNEWNAQw+qqY93QkTsisJDj5F59LJXfu5mkvQ58nRJqykqIPvHonUdBvRXiNWQG2zhPicG8
FX0Tn6Zo2Ubd/z8wViLA4VeYhGCWR3PPDom1sXFCHjHjFBg58tXJNSCfXI2ZcvIqNOOjDgW75Dxa
YB1l1DBei74FFUqE5n6lxAN01diosYBk4n14MCdPwVP9nT5KPi3MAnhYZtY0xp1+ae34t06cPulM
g+4GqQfl/rqngAQqnlMaWnfcybxUAjqf+Kf1z2Ea+4TcD2ebtw/J7TXJcCa2MuarQbtq35UjKYK5
pdYgUNEwsaUMq5GfTqdEuzrwuSo1NYeBLOg4wu9Y2hryzXg2fKaXSTF0RTRsNJ0bhug75Hs8+qAy
7GSfU/ERwuzK+c9+X6uOSKn/llbujTVtDRY8ewt6Ksf6rtprPSg4t58gorzrmbIKl0O3+xslISKk
A7EzzIkoO/Kf5bpzO24ntwEi/18+yjfkR+Hni5ooarxf8o1v2JKT7jSY5j+6RUq4X94o7U0NtYFd
qSMVUhWGm7Fm6E0omngEgg2+uE0odwNMZ8k7SAe2qZxj0kaoyLrNLOaIf0ksrbOxuSt/LmkHCcBV
R1XPIgYEw+d0WSxxD7n/VUEu9vSbjLs0xE9PoWEXCGJbFpE647gL9Kl3hpHfvk6lzBrQ6gbvIj08
Coz94Nq3JSP44aQGA3DwGW5MXZdhs/muOqbTgIuCd89dUeUA+XfxlBwH71hQr2wj3/UaOoMVW2QW
0MCta7lC8Yq2k1r5sd7M12d28Br0FwdzRNbA2L/2NBh9kWwPIFfFxc8oIoXMjYEyv/cQDb6xqeJ9
c6bKDOACwuXTwSuvwpvs7kcwccoCITQxiP842fB0WjNNLrot8AlNYMKhzWPZM2AUm/QG/6po0YIx
wGbag3hRAFRuVVKkRYuHwOjHybyIk87TEbNJJ7KLslpxd4iRqhoSKUB/kEVD7hJE9fEcNH0AzbIA
ttZUwG/H2DSGx75OfX4OWKmK7u/Eatwj9PLh26Lic0ZYbad634yQdTI/kL0Ac9XzmYFum9VD+spZ
at04eDco6k4WVP+1EiPnYwWL1hVFE3TlU2whX8VCVRzFGGk40JE0yZwVa81vkD2mZ98Dlnsb/gzZ
hwTiYc01w2CyDPBdn7n3fnPDcOxTEmxcqHU+HE1rRwPpLnGy8T0XocDe+UExaactdUots7Q457Sl
48T5Ft5qLAvXvgF5KxOrv8N+zwUThzWv/F9sjTXOtiPHDpf3v3Ap0hbBmjcKeoUD1NsZLRy2L0lo
Z8BTtB0w18q/ZeY1uijEg3X+Uhg/6Zx8PbQ8vyseCTs1TQicc8v1LrLNhor5RwfNRhymQJYY317/
AN6cwz920Xf/OZPry3LpAm1SZ6p29RXOeVHdlRge/ZNHfAk5TPPTXsAnDO9GdBI1yXR80OY7CEXf
nst/s7GL9W258vPQowp9J9xZuiQanud1C4uCHiZmhHpaX/QcgXeHBBp+SYOtlskmcRz15TBBS85E
UvEZfMHy/t5tjxfz9p9hO3IibiuEsQCCD91TFIDjjchYgg3cLKTyOuSk5iR5K6N7TwBivfuldfzD
CIvcu+vFnmVld7DWFQErBQwb3ew1LESgdgy70eIh4frM0rTQK0ZW2kEYogqOjfY8wQaIY9UPb/Gn
X6ES0I/9xVpxhfUz7EfkamGPbnXNSNx5WU05C4MbJJefYqAG9WmRY2oIhwjty/J9hIweqNcGRiyN
qxZN14jS4CA71yQ6CZrdG4rjCnkKYxGqW6ZsppdFDLWl3K8a2Dkm/G1IPpInReRwcpnd33bk9FHQ
J0TlsBW3O3DuBQi7uCs1zqWGpFYCjzNic71wF9Cw4RJvrlmkpCN8nA12bQqsBK5kJEOiOxcvdaqd
y17hZtDuNJ8mQEtk+GGh5Lz9TnCuMxpDkmbgL7pG4iARgJ1cm0TqEctYpgIbaZQjY3nTNL0Pnoyw
bvCmy4p3JazR98hjSPz+WaiUMuXUFjq9KcN1fYJYP+K89ZjGjK0lusdCk6quUYZvkDZxAFEMzm9J
Ozpn/0sMnfLot4Ro6wl/ecxq8B/0PrbPE2a6guAGgYNDnpEuqT1AwnhoTuKAM3dp3vgeMVQPa/PI
yqob1xNAb54wldp4f9XWI86UfcvPFkxDsf3TIu4Lb0qrpkMmroj65hI3Sk22Mrm+YC6CbzjW8UOD
inVvynxoA0mBXUPZsG1yL8BL5eqJkR4zP+KJoX4neboYIhbYQj20GOOETcOMJ+lW+a5D+AcquSm9
NblcVzbOyDkjAotpVMvvMsNUfCFHfKVfqnsjmdkNiTeZ26BdmyMnOghjnI5x81PmRb98quVN/DYp
HuViut1CPzd1YSgoJibsNAvt8VslixihGtcGEPMHb47hv7d2lQMoLd1QYfe2lUMY9zLiDbqFCUqe
oHLS3gGsFzOFbF3pQOHfGBgjw1ljdApb8eb7fn2N42OeDvZeUi+E362x4c1Fv2I8NU/safYdMUfT
3k6O5sSx5GK+y8jVohPJssGIToHUZu9tyrNywI8Q7ZuAtMAm3jOmP4c/zM6HWAAIzUyV/BIANb3q
uHF+BnjvY+nM0ACHGfkP5riZM25UXHLs6E8KguRSYANPoxhbLXTp66RjrgEhP5sG0yuviPHyP0SO
xmrDjLFU+m4pBpmYfwWNwuuI7jRsfV33C48XVbxctUWepjXAWDDDgsbDzyXzPI5sMLf2Z7geejEk
cqCn/xuMdQi184NHpceetEY1+ECKQ06KY9Fb6afYB8sAcXrFOCvmw+d+R33obLs3mBqBfQ98QMrs
qRdYwNOPqbJXK7pGutF8MWwiEJ25ndwgbmjPNoUn8qR7jIMf7llkVT1wfwXGFQ4OWUOUSlYYYV38
bLGc2Yh0ZOoIFomsRSFCUHKB6Gkwya3qE2aZMARNQP13x+t4mxo6wXZi0HKjOtGMCt0kQN36Zu9q
4P34AlsoD0QttGS+MR+1cEoDTXwQEO99L3iI3YLjBGDJgK+lEO5zUqUjoqbzNTwuM7tRpGshMLeT
POfHBe7cSngmgNxGxnT2x9j7RXVvJnDhhhaziGic6zjK60wycGeebl2PJZpgCuaEApL7bx8sm3qs
kpdo1nOOJVA0ewhn+4vl7yTCGwgmmUABmZjKZk+S2nV6xtBj8DOKAHTKw4wowAXbuH2ItkE4LsvW
3/iV+DrCLXdrgbW2ajO+RTHMDia+B2jOo67C972wa+zwxmMUqg++G+aKN36bH/FkBKlkpyQSzjFp
Bo/pR7LGmqyuqhrORnr5rMpvlKF69up7mGAauIMvmrL6J+dkzVrQrCHg2p+wH4G6hJR4uPQ6PJVU
aN1I0lPYF9Yf5wy0csAWgHazhyDWWSAH4KZvC6UBbzIvOD1Y+nrm+TyMw/kMzyWMWHfUIw/90hgC
qRJ49dDMLfHmCmzCsunH129PQvmOB4aeqQ3qGgfgpVQqsl7bOTfhdZ+A9pXRgp0xd+f9r38ZesR6
Krwo4YLbTwwNg8yMH8WzPVPA7/59ZoKFYA0gkibgBqmGTh0g40KKlRV49sejqRMEo3lqMBPrzOjK
zrq8IiDnVpdypOj1gFW5+1UxZX4jvay78jyHduBFUdmACicoG7UT69hT74t++ioJYeQR/tGjyvkj
xqbjJcB1zSmJqgpFL3hDsU5lmrNAmm7Ekgsm/HEaV0HrP/oZtp7iKNLWS/RWQ3w1DaK0cOX1uDSj
6Nd1DJaRBkB24nOTWU+2xDiF/8/Yp3d1UKyty/HsfC/qmg2uwSZv4eLdUVqEBFmNztyqxu/N90KQ
8vfgx/k2Ftwl7elK0iytdTi93/RWH3JwkVjLx+JnrOd+KGeWMZ7Y8rwd6DfIsoXdu8HdO/bxuYiT
r/L+w378v7U5qxb60ZYbMx+v1cLm9hfQB5Pv2paTsmU6uXUPmVA9xFriBbbUOSMINPX+isrHOy3H
Ow1M9E3TlqJxAvTKLnPEjap6iAzF61idpiCogfnARzL5aB9m2pqEbWzKX4kjoeVSK2elfStrCDbI
EVa20utqGKtOyJ1/Qj5HWZdRyAAqlXWydaqKR9iOv/VjVBNeYvy9La67Z1usGCWWkktRCMxBRWw1
bLmMbZwBZ1J1JMOE86GmxGnRm2TOCVKmrc6bEtOzqrILUJu/4IneofZBiEZLNcu6IfUuVJMVlw4d
Ew9MigBYLyPlmt8CbMypN6/Gq9qQncuwn7ku8iNlqtNKxoIhm7Tb77baw0B9cEz4V48CDn47ZA+A
+H+LhIJqlCchDnLvdk2M/FuymZ/Vl/jZGDVB/o9Fs4OCMeSj+xkzVbwjCtq+Gk3MP8znXmBC1g5T
wpnYkL3J+mZbWiK8+ayKlaDm/MS5644P7fPYxojoMZ+4XQmuFLQM4t4a04Ov4F0NKgvBoOWxg553
XTJd5NaIjW/PjCshCgCumDUWqWQwpMwrHUIU+46GaYKPv7VRzI6rK9cTMJXGK9q0L9/AKgHrXEd1
Az7TnNu6mXCjWxmsreNV3KUpAxK+/XhOunEbm5XGPaJr5kre4SW31FoEsR2Fg/AbAqChHm1uMinm
jnHBsZqTR/z3bg36KCYPuQxuD225R2XN/LGf9ZEHvam0xckyB5dayNpfONFGsYzU7GNuZIQJpdqs
7DCC4M7QrYs5tSlsDUVGkfVIEVsR+9AawMXKo1RjYtPbWWiOzpJ1OtNrurkLXd6HsQ6u0GYdmwqc
ybdk6Z4LzRNRCWgZmb/prwhqntfIrCyMgBz88dsmiWI7GZBLsZZi13sIUu/3J/1lnRlHmSm1dwgT
2s1FF+Kn2FFVGOjgR452FhTp4OfvIUZKcFvZ9JaRjmDcTCG5wXQMcXTsHOBYS1kLyr4JfF22tDiU
VsonPJ0kYkq6lqfrqI0UQx5LiJaWnQL3masDsC2xX48moCuMxpxg0z723MhXN+ceN7joZo1l6OFu
eD36uSdwHYdSX0IRvYmeWkcIKxONyEVP95hza8i6L+PcjJ2OdINi4onbv7HqydMPfk4wmsUf6PKd
VagSiI9XdPmdeC5VMfzmsMWU8I6gHDaysZ+t60LRUzge0Ii3Nk6kAmc6v3TEUKfQKqYAIzyX4lFH
qnyzRIVUQHKzKe7XUjgc1maSko+17gQK6+BkEKspqzOqge38eiu67V2syVzvAcikZGUnZbwdQCYw
SHBz5zmAaysaqi3K81X3Uny8zSqwimiTq5NL5lJYuD0JfjeoxmsxuttMbkuCMKhcDkJ2ePdJxU0B
yKpw3srLsKUwhYjv1zy0bZk3vpyVyMCBr/t6hHnXbkIIzFLvahKUn70cp6nBcCudCDtiV8msb8fT
yRSWQzcqFklU96dQ2sY4+kgyE+gUQomx7lKMuYf8yv/zeySE1T/30vgKHrZNl07/k8oupU53CENi
kQEZXfDD8/SQqbVJ+AhEH0737v7Fex59nS4DWoKbk/t29XWxPFiDP6u44NoYdcwaYvMIaDvrdCrT
KktQtejtGkBwqcNM+pHJisS2WyopzjzUuxwHjz9fb7SrJnkk8/Qi8tlizeNN6M4/74b9p1i97TZ1
+SKCoTeaCBih5PkZwt6MVgjdFKLRELqRyTUlFXdg62cuCbw1W7levZZz6BJOtl7Y7A3gHz/4R4+p
z1EuTy8+6z05CXxJomMXA8uZ8hW11pQ1yAS6voUjVtq9BpPULSyHrZTmZQjpN/h0coDvqXbG10RT
AY9cArDg5dKRArr1v1BALb958pqLcSqiAc2JVxwCBTKo+hBHMgmsXhvHSQvZWQOqwlRgT0NGe3EK
dqvJlW+l5M9PaeyRVHMaA2qk3RRmOOGuT2lYJ0TOLBdFnC+X3nn2cVVv3xl5TINctJU4ufGj6dGv
rDJhzfxzRcffSVtE0fMRMkuBGQnH7MsD52sKkP6HnolKNUF2ABJGd61VfuBFa+hsCl6fwVmOn2pb
L8VLDbxItk5333Go/hyH4UKcRWfLr6AmbcmVRmyN5+Hg6ute+hWaV/opOT6QPu/k7u7f5RCQmBaK
aa7r2rBTaA1+yvN0CMVCkP+ExaYqM9DhX52JxFIRCC9uzfXflSjO8PTxcvTS0LiIa1VMMzLVZ58j
i20FWjlSJHDfUlVZGvYLY+50g8BO082XozGyxBQoUZooJGU6TRQ/NvTSb+bLZBSZuoWYjsugKZm/
Khw509neiMgdXcfNljU9mMudezJP/5n+J3f+6JkYj2hfR9MT9AjAlvNePMOpQ96Z0GxU6SZF8Yja
kwvmttf92OVn2BhuT+JM+kZR6VLtwQxsHVHjtjsBurjJ/XFMVeML4GZt3MYIsSAMtP0xPgrtdG90
PqHobKgZVweO67CXyIOwRqn0AOrK7qoDUQC1QkJFGPUFwZntwQCBAH6VyMNv2bvsUnxjFgy/IY6P
p5iCjQI4b7wUCGJQF9bWv2bvoerLfip+HG90W6Lu1TKV90/SBE7hbJmKIVJRzTE7VhlKlcZwffg1
2jqGNnG8Gd5Rz5hwM7wF32GMi/30KPCB1wvrEdvpXS0Vk1jG2r75NLAFg09rYlPyaSk6MZVk7u3m
2IWcTHpjvjcckjGhBp78yWbK4YzBidTyfuBhAJxO8cfeQqNXKcJcktogXVYHSy6IYX5xuU6HzgDY
1EAlqYK2OCaOfc3VCKC04LOixSHvhAEWdadUN3pc2uGOQro3UgVTxHAfdwafI8NcXnEbTqlXHd0E
4wyRAbTBwU3pJOcWfCvI4TgQ0OdX7ysimYjk9uTz0RiB5K0EARjAlh2lR1/EmwqCOPn4JG+/FsGH
jp4EQjinfZbtD2oqnZ+eAC/m3fbsJcc0yt2GwE9nnyOU6kuTYHMdNgZ1CqIFUCRct9GuSFbA78ST
0/gHgJhzBvJItzZlCpqDyvvf8xkPnhQ68VbylCqUtAy7z8a8/mSTnoyGe2cb/zyi9CycOiGordfp
DLnVV88qiRz1+12u6iIJ0WPQSC8eibIw1LoXk+jR2jEJN+taMWkbJ197DlMh6xZD4FnypoQuaZC/
FxnQ+ghBCOjY91WvjFW9RcrAsYziMaB3MM7tZYdMVHZsTOOkQL6G+94v46qZB80mFbYLqe+z8wAm
2YlqelDYuMBmF2fJlVJS/v1SPAShzOBw8qJoraOF5pfQBAxi6iHag5BblRln3UESBBBs620o5+4M
t6D3ycgMakqZp4EbK67PWdQN9vjNRBhTsQbcCzLDUEBWuUSdT3DPi0X2DB8qAIalyre96tPmw5QY
jEJUaHkXh3TH320LcZHWgRUJnxuPNXx/ey3SrQQE+7bc7MdJTTWjKSmfqLk8OrdB4tDh05ZbnBif
0/J6Lyt40HvS7X4F9dvhJVxOey99mTRweimLvJARt8IfRpA2csWhS0ETpctAWmYFD9C1VGSWlhji
eymO5Xdl8zjElvOyFv+l+p7GYwUbFeJiZaj2pihblJMb+Ko/cnbsKxHVukHsSrF88wjEHS/rEJFR
wgpuF9L6+KdZuG3PAcfFUwrUKcfbv9+qlm4B+QOtBjmTH062GnBapR4ZwRo7TZYkVkSuYHwWID+7
HD87uu+0C7Bsm9IckuwlCz6jGIkPbwTDZAflZ0dbNOXscBlz4hSCh9jcNfy/pFkIPepzqRwCv54p
7Q6afg3421xK0tjgl44mR0jryKewX9PrtF9k0iKD2FSbAuy4TzrmUPGLn0W9cNXe0RAUz++Bq7Kl
AKQailuopbc1+gG88wBxIXcd+taxCtw4OVVRqshiP4ImiI/ObFRH2kD+uRrPnAdSe9jcyQ/P9aDs
Sks4TNa+7tNckA0kUpSk8uwJ0q2b+tIV0cUXrgvKwKLPIouLIK//Blz6c23FePeSXZUs+Ny4jbzB
NxbSvXlFyWdI7R8qqIce3S1m7DESGfLo2JMXzlch6ZTjKLxGEogfSNp0E7VGTJESQ3K8hR2i2frB
GDbeAvflHJylZqbAr+mHGQGmQfQ8LqKOrwTzvfc+amrPmhPnijFSrK9qkTSvoFoum00+6c9tKiQG
aV5/x02UipbzDBzCcWUj3E3aCuNtkA5ilSrcofL1a0GCdJHtnHQqPb+q7IfWEaGQem8ef2n/dGNk
C4Sd2DZ46e0w6Lcow2pudP4cg+W7+I+SDNPxOmKkfQ1X9xFelA6LqFUp2EJuW0LWR0puTpzQ/h4M
IrOi/jPnqz732HLmGZ9p5jOO/TSzRslm4EuQgoOYGqP6Lf0aZPq09odTFsP4iQU8VA1t1WZPpKQP
dEe4XXOVxS2BQW+TtaG4S7xjRPkmBM6dLTsf92ENhq7mHuAvCo/txEinleI6wpWLhEOc1Vx/wTES
pyrpkirvJWXE3+K8mpoU+jb7Ktj2TfpPzNdsp6qRa5EspHc/lliE7sRBoDF5cWBPJIsu/AoI8Rol
qdBm0VScNe4XsZB8HwwKVpbLiUXr1R8omxG0IGOTRwTGOGs0gaTMzsH6YbpPQda0PRX0xb4mfNLV
QMfi24Y19fhlfSJEAERGEc6C3Qze/grWO+MuPTSeWDbs9NR9HMYYSIKaOVNSeHUqTtcbaW5/u0ak
qx8RjU8T4k9wYv9jkJ9KKND1qKvbz+bQ/kQLtFp9NNsXAERxMVWre5bsPNnMNPDf9gHtmggjxBVr
j4sWUI4m2vYLJEBbjs3/jmQqODZb1SscBnZGbY7kLkxIZZXdDzILEuGzGt7nnaanlS0KQ339aZTZ
yZ7crH0GhGn0Vq6sCsyo7+aPkUu3FTUCCTWPiN29os6q+D60OCuKHiQoI7zZTlVNWLWaWU8Gf6d+
rxoF0PzkG3j9DGkOESO8kOdEBMuoocSL8LRUuE7YBTtQxQLctyXJqaD0a0AChsDEPf0xBfnoLurt
jGAe7P1cUQx0/NqVueRo0CnfI2WUe0XBFJn+55pLqYvheOCzAFFHL/tg2xsVOx5TPPEKxeWT++U+
ZUashPsPQWxzAHVAOHuJLhbrFmKl/sWcrGwJBWhn1w0+qWuDR9GruqYL/l0Lw9WVvvZQI6qnQg9z
pKuCyc5U4GdEzc6/5+hq/Cm2KbxGwBnETaO+ywLrNuiSq9s/tIMECdrgCifX6TqKYm3uJTvHal0q
3815m/iPTe/nxP5lhJ7gHmpdyMY9r180XvGUyZ9QnbTa0fO2MYSsFv1LImDmzgQfkssOezQTtN52
W4eRuNPXNHo2EX1+qYZDiD0PNZTwkPNbQo3M43rdwO4rmyaf/YkL+eScUj/DNj9cSjnapO4NFqym
8gNirLahuNEW7a9YYrPcgC4FAAErK0MrH0LmtasjJlPIeSzWXEitQn6nCrgdzNdfL5GSTG+BdRb2
LOcaUw57TOecLa3MAKaD1xX0X2S/Yhl0oD0Y7XRxqoaE63njx5tSerjGmspVey6Nf+SdQe5oykpH
fU57e1IzAFffjPsNibQfAihm7JiPkuBE2vTBhIPIKHti+FEP3J6k3pN9qnRLg5okMOikHhjO+kxL
vfzWzEd5o8qRREDMZKRFQEWh2me/Wd+C4EwdtHwJk51R+RL4a0JhMpmICc7dIJiKNq39H79znVtS
BpSYWMBN6x41EjNsKqHO7wZC8PUqmxKBajOx3kaMUgB8Ic00Z1ut+vc7K7DWS2F4CXwGV/UiJpI6
ShCpXWSoMZdqQ983azRqE8sL3gdOGNCkOMkL4qmuQSOKZrBoDd8l4ZjD3y5uIx0/C+dp6yipYykA
VPsQKa419OqKat8e3cr+pnRuYn9eoH7wGvGWGDbs8/qXONtCfVK0ViPw8qRbHkSIHSadoWIUjZAy
MVB8z8DHTdsgxxM3O9eOtg3Gex9bvgXNyX+ID6tSpcRuFQB205lzKp3uDLrd0f9h3Kc3FhiooPRp
asFpkla0l5jSsabWekw0zXDhtTJF4yE1ozWQpV6BvtGjVCidmKTkfuIgIjL/wZIoo0eCVE8tMMCW
257WaalK83mSzmVvIp9bz3U3Y7xApVf1uLZwOD1HtQhvXaiT1GpoaTTKzS9G/cY24g9+vhy/1Dw8
R3axb/nDXmkPIXPsDs7S0FXu0nxVbBgiKGxiEAt8Pxtm8L/uXBuMN+b+8jNQMEP0TYVmy8U7HGy/
pY8ayPFPSNEKj8MoiObf1/0KvA8eaMmqpM1QyQdCAfGGuq+7LKZhHgbcsmdaCBmeTEkhTJjKoA0u
Deo4Qy2WyxM/wEi6P41GNtvi7EP3kqAlew1brMaNskSsTTZGqRwfgtgjumD8jrf0lccsRtYPBOI9
/7xnXIyG5vjzy/qh94BMi3ltKeiHQaN5tYYl6NB7LMEVaXmNZCQxq2wyk67OHfCoCnq7YFp/9eLH
NfHyfNaMr50k04hzT7pzASBCIuh2SNgMV0JwfZeTYdHuM5ytTF89jxVAsJAQDm85ajLH2IO5kk9s
w3CAcuAKDeqZV0naIQ7iAlbKwFQbrJwX++6ahn6MbpTVi+tF2H4KeNA+V7FRUivy0ZQBR19LK7uk
G643QbaBhBb1cr7aiZSAPyeUshfhDVNJg+Pco+bpZkcbhA39plF465zn9ALr1NhNgNlwhOuvBdXK
oChNXteI49op3biC67zYiOQf1koeJUdzHryyzPIK2Nw/v/tMpzhq7e5V1xnUtY89ztHZcs8oVq8L
bNiPvdTNyv/wmksIlnGcLVvZAzCf4b2eWBXsn8la1MurYCp3pXwsKDSbYVwMZv7nyeRACRU4CFfg
1ghyv9hVTSqjDOdJi9vSw87q5R03dgRCwLjItf9AH5LSEOuSwQsi7gyCiakltF6Uee84/iI7W0UQ
T+2TXsQMhxZS9sUF+RSuTmurPR8yF5ctcLUpesZlnTaCoJKREJd+J/tsjEqF3uRXgxqwD3HRhLZs
iBdZT2bSjZvrmXbOefCDck9ur4mmzDZ5PBFa0Bn50KKXxIxpHZ2HoSJmfuBbYYI5zPNVeutMeE6j
2sj4b5djMbQAntyg8eEhABhg6WcdpyL0edR2JrOt7e1NHMH3dvS2/3ilqKYn/9/2PJX3i3APNO9a
MS0XEeN8ImWDYj8KCFBeK4JKnVC1IzxwxL1P8MTyw8RGwuR6r6ACp/tOB9OCEpmMsmoc8XJ54R/y
VnQEaNGVoPZuNUfYxe8jDfiyyI2/Dfi9yVTFN9H6fqpLsH5DeNVSnKJvgw/xlGUncyjQTCVbrPjy
0xRPZsMHBTWUrRZB92l2Snjpnp3pd0b+S+7w64Kc9labTjc6GsHgAqW+QFiM/bOSGjmdDdwUXDkK
US4JuI8lGk8OTPdEOmLS3umV6Er3cBVbTwymI6yvxFMyFmEhXAkEHM3zZdC42zyMByU7LxL+89UQ
IEQcJYwKOFzmvLxLAaY0S8yal7Bpt8ysgXE7k8s6ue8iY63EaN98LtpAN2NfmWaj4qyR+BZsl28m
nHQR4rSiHcppE1km5IeEo4A5HqMhaHdPXbE/RIpJ8sywqpyH+MA5aHvuNZ42qOEoERplpvFupbLf
cHS8HSwtaMEiNVIEt5RRGFFZQ+mrtYuMeeFTJOYXTgOlZL/XMHyN4nEKWvd8TpNx1zMg5OdKnrKi
8X6LGlvl2yjqr17fzAg/qST8YPqmoqdkrMfbXPlEM2rt4QoGIb+/x3GE64mEW7R6wkmPM2LP4Plz
uZ+5WRpiL1K5wpi94p40vGnCGSMIekO9c/4duckOydjtbkgRJ6HjI3XdYPsY7nxrlLnjkWNamsrq
TyzQWtmvXfysA8v/xemLb5zRqMs+J2vyamomFwLVxJECZD7+Ej80CWYWU1kjODzaGvxkEbbyu91Z
068dKhoZGaicaGsLGANM+0kG4e6ZwbZYX7jWo1/jyVyr6+95/+y6GSRZengjS0fQsMrpASJOFHzd
ulIpQ7mtot24WIurwttH4K0SqAuYnfgx3z6HKqc7kxmQalmJN58mIA0ySR+GKopEKInSh0axfquE
cGRliTFOPOI2o3t6IVD8R/0tsqF3sl85w04c9endhR9nwXTm0GyYNK29E3UCslHUw3oDwnXVu4Ny
QQ4XhYjDjsGNVc2ybQmqhcAhI3vGkvp9NaahHmfvFHQqNycULgmocnSmBWZP0R05iRhdI9Un2vV0
2lTX/DrGoxSpfwyvdRVW8MAH3qhdWxEIzjMsAHwHCgdF25izs/TvaMttwJZWQp5qlH/g7Tl3eOG3
9lPXlNwGLSya1OroULc2n8xOaxUPFX8f2w2RSPWWCc2BXfnv00yl73zAwXnq21F3FjxdG7X3XmZo
+kLpt6tpZf5w3SFSMtYx1iwtVogtogWgs51sPdeyneoeRRgNd2VapN+A/b3moCbQG0400UC+8Fy5
sfwVW5mWWfmfiq2O3Ey94fSQmXlAU8SbrHJdVv1xCywC4TH4ZxhInSb/rtxDQHOdBiKmJqlR1KIB
p1Y4GSESg1hpArzZyyItgv8M6QiY67ka5RH9cxgfvzrfztcx/WMYPZAp+9olpkwAPGHC3+FrC7W5
22VhH+v/zZVtxZ9RB8PYi8AuyAEkiVlCpDieI+fb44CQmMjpCtYbglB9dw8EVWndYPOIAa7wiuJK
+v+nL6Euk2cO7/xWJWMpHPvQ6o6FJZ4Ti/NfgeD9Ta7JifTQiNXzevDTigNPZCekLXt7s34nFYhQ
m/iQFYNdlJGfrIopzF/Dk7VA7G4yq1XsSbbUh2gkjOCt4EyzmqA2tVZX6juw+ZIx4OV6/pdQFOTp
8UbuL1Nx6121CxBA9RA3ExIDqmkXraQftR9RY1g8mNxNpRpBtldbAVWu8M9CgWoNaoEq52Kd5ZmR
6ubuFY+KDLj45zvpC+cbeJedYiM+s9k22EMdo36/gnVf37xJrfCTA2a/x4STqPFVeSiSwKg/fpps
sw6sArVnT1xfu7wHxcreSA/6lFCF/1408naWGhLOpxwZQVIe8GcT84I9TBX6TW4lV1cjqkG4l7lO
K6dy0kwdhtpJAE2KrbR7E5qOTZ6Ovb83L/wHHlqKxBQnDDmGDQ0J2q8f21bwXRLmn3ag5L9G+hZ5
ESp+s3/HvMFwHArXQ8Vcg1+wSrBAmlebz63fuCF5mc2nMT8D+W5kV78X4qPIJ6zRsJZ2ISTrRxsa
xB/Vp+7e1m0WmQIQ08YaEP3dNHYAmo+P4p3QDnrBEAhw5iHP/XZuUKl1d9VcQRzTMYwhgEFLStPP
K89J5V+6NZjlTHh11Nde97c8nDjetIt2r3ABKD/bQ0OpasDx22i8+TGy3IdWKPJauDlMoteoapPG
f1kL51u4iSzK0fgIjGqO5V0a+rVL41e4a+LES3hirwrwk7dkiO8Svv/ApaZmdYANb5qgKomW01yH
1ZuWSyDdQKfGGoDOGsvmmKkhraAZplM1Fnq25gzmKvGrB7XsPfHZqOtcLp+A/vXHWxQzj/GA1/KD
elqoMEwU3kSwS5VVQa6hVT1Ehj0v8pj5JZuIhdBFavNJChMq93UOgorb/pVaReJnibv1jCtT+yh/
RyhCPvPXEqSG12mnZdNdx9gf/ymlnCF8iVYDBAoPfO+WBtlt4BINmd+nQo1Zi7h/+WjTSN4UZARw
PD0yIQNkRDzx9DYJJoUo0KBe8NZe12IH466Y6t4YuD/4euXAq/cTDD/Ibg4tHq/zoVLpQu7AlNit
E6qND+OmPdfGSEzC8SS1q1dReKI8AvdYw6uZb8CkEPM9r+fwuntoJGBjIZx1xnDFpNhfdu63p8Kz
RRjU9EUf8DIcjlXZwuop3UDQloWT1GItY55IUVLR0Hgd0igOu2KzZNTxNUZLnn81eBPebTV8SG7I
m22TSHTXSyX9RWO7dmEUzbLOvqW0I1ne2DQngw7+Tz+LhRoSGREDsFemc1CBwXcz7r9QwUeZ4JMQ
JYLgZQ4gdjvfmruA8Vx+1ymhG0JdOtH06ZrACQEPFFXcAxmSkKup7DC/J+OES9J3GDC9srxf65jD
8fSi9Z+C7Tf8aCuF0p7ZLN7swrJPJx7wKJOo1EFNYm+4yy7TLMPnnvdnsDNtb/TurZlwn0IjeQ8Q
OWUqp3lGYt3UH2yN00wOdf4YG+T5VrdvXfr9i43sWChmhSPGrSJJ2cbTbFMwDsgNNs8yJ9iUo/vI
fPDLc4rLILtbGGGceninCyVvqnd5KtLFy4zCHOTkkPrZiL/Xyfl3yHtKgy3f+vF2VjtM2YOOEq/m
UYFainJmtFWL4CVPLY9nBWpqtq5sQwAnJ/xOr/KNXCezAGXGEjFaTUoRo06L75TEKO9sSAH7aZkC
VUFO/vfc9dtLjtdnVepLjhlbLrAAh50YObsGwnR9Uvah4/Cuaj4ltAAmrfpc2WeGwqssTIMW48//
QmMWzxwhBnSvXSMxtgjVXPsBNeIoG3Y9k9qFg8JHXH4vTsvmnk0Rb21RvKhxaHvqzjhe36JVAWxt
4PL7TlS90ItEV1JjYBnIG1+BPvLtzjyQ9vTOaLfOWs2JdMjcg1hyfgsn1PYMxGU8wm7Du6oBi48z
cpMsV8zMO/I6SjAnQn9DazmN2X70kF9fLVCcjZzDN+FCsCe+G5GxjB7kQAMnc5J4SVc0xZY9otJ8
IQsBuJUywtCqBdWdONjOnNL5YOX2yfojyaWjMEBk1DrqiUKmgAG1rI3+hASX2gCrVrFhRSSornmt
rTpByZvCavIUpSY/vkYJkCGsHcFkElVNTySpA2b+eyG6Go4xE/WH64OzK3DZ7g3KT5A1JFLtML9y
kqJCIvEhZw2zdoeNi2S5MKMq9GdzkS7dxnGc8M4etjKiv7vutX2Gm8aFCi7xgFy6acPRzINhQHm9
DCPlifCh351wrE+JEL6RJ6KV/HRuoggfTsB1n0fGQ7W5GWZ7/JaaRLRPsogrIz5u/DGZZ/sLk32m
2FvvlWukmKxN22sEZOeo/ztxOQ5yulpkMvkxhcL6P5sGdjJN7ND7hEE80PFtRGqzO6s48tqSy2Ka
gjosAMlTDbr5x3nww0Ks6Dp3yZMkSgdUJEl/jUnin2lmYgfapRa61TLYAUfI6xDCT2LOILnVc+0z
IIk1qjAgFg56Znji9LYBzoF4f8nwmWVGj4CAs6kmrSClUcmk45is98II3aABWESJ+lqYjsC7o6eX
GQ28dnbLYWAU84+7DAylXNDUmNLQGW/o5ZN3Deg7w/8EoXpXz81IS7YYGD/IPhJWkyTNisMAh4Sh
rmnHbLWaDy+arjYoAAjmjqWAMP0Rv5ex+NYbsf8/CStXmk6/2nBtRXFF8757DX01Ub5NYgiOBh3S
3W+Yd2vFw9zdGEnj0EaWXiKbBdd7Gqn7O+/WAithZvxxSEKLW+OpCTPIBSnEcjnE5cTGCQt/AQw5
r8Gu9/uL3COI2sOKtd4Zezmg/RkLK2zH/MwU5JD9P7Q2u1exn5NBx24F+bNCteKKbosqbl24QTi2
JmsD1EtY2JFAjuCfDtyRRAXQbEQyGienkPdX4WYWNZjBMt+L1CMDx7kWjY0dCVxTrM0i+NtUhhel
d2DUdTMjkGQxvoZAjAyOo6HLYA0E+Pm4HklIacYxc0bP34iBm6BnfsMumPS1wWeFtoYfT93vIY9+
9BhtgjE/ebTGxKoz2gtmNBfGpOtG1l5ZdWZPIDDdI7SAsK0+Zxc+ymcHoaXHNur/z1XUC4Ksunsq
XUGjXD5JziDbs7epNCn6O3cbAymngMUB7n3zqvQQNIlwVFG7GhQzlC1eq9tbNT79Y+TR/ss259Ke
edHTaZT71NTYA3EUakhh3xWR1RPsOROEK+yS53HL/j1e4A2GH//07gtRJDaWAHMBBgCM7xPNzRWL
1fZ0Z6zsN1cp7SP3Ozb+F6t+mLLT8k6hLGNOVp0mi3y8sZ03Ru7JuqbcSnsR9sTumqoVTyStDHt7
RKjJH6Kho1uUTNLHDhvuKizGLZFDXxdOrMD0NZfay+fa9liVFRCj6P4mZygAUJf6zx2olg3uD9RQ
QZpxgYS4iknyx5ouDBTJ040G86twf/qnd57j91/z9s8k8X7U4gkdeEsznlMv1drmbEYOe3aWieJY
tejPhDSZ+fyiotK6gVixzFRa+deC/3+KX4k39/TfT/RfOFgXyEhr+co2o7e42wM10MQyd3w0KLu8
ae9+3/l+6VHF0KqFuN4PMSThYrkkzgz4pNoxmsIbMJsISZYMQe8bF7kG7bKDOdlUlyrdBt107mi2
sy8Di0VpoApPR2iU13k3zQHirZ1RYg12DAyUakWG9Cu1Au50BkGGCB6vOKX4YcCWHlpcHhIMUys0
5CIucN8hT49w5AF0WUl0ulAjldGsH6EMtDcNQnb3c7ehjdk43P/Lvtk1SVd6Oq6vTAkef8HZ/vz8
Qf/aD16NoRjmzV+shv+jW0ur48Gzh4peZ5uI+oPhiEvtAuVA+UeNjm0M0X/VPZUvpnxp5413VaCu
hy0gbrBB5myjX9Xn93oDY07rpJHGDY37J6vUTwZ6IIxjGUgvuWfJn0qx9rJN6qQG7H0lQXXRfe2n
WVP6jsTjdxYm02TkUR4P5OE0ZL647uYhBuZmFKKVY6039r69Lc4ixYXYnUmX5MR3qKDoO2s09MBh
Y5XdRzOaCuAr4VPOoywKcq/DCOYsJEAOnvDjgTVKZROBQOSkcKA6t7Ap3+3dDNDG6jfRzYlCL2wC
6bGjGbRZdov/i0iNNknrFs+WXJ5C7LLlMn6dRj+GwPdf8J0wmj3LYTupAy3jylpccrvfYsaJ6T55
WWAfaCLBIgjq83bC1fZCtXnyyd6NRAf7Qi1vrD/jLtyFCFaxRoKrWA8qSDuZJRz+Er86zWDTpHWA
MQ4y3Klwb9hiIXt53BBEveJCl789nr8z+Hf0QcBitrEILWtpTslK7mM1szG/YuAAD+DXXNmsGRYX
oaPWbEPnCKXPqSvyjV7VKN8l2E6FZutdHSYqW7CTbCBDJIu6V8ZFXLUYMAXilqj2LiZLMRKPSDLD
ISNX5EOlHh9D6sr6UDsNbVlPnmrEieDuKZvsndiU2rhz9BKfiir6u5+JPh07OI4MIzGphRgc+1np
RJryLZo5n2bWURj9D84psNDevm1LdEzqtgjAHOEzk1s2m41A48AdCOZIet3SRl7JW66o2JZyc0Ey
ivuYmC2N/P06dylOwTSm798EjwZ7OD/RrzVEB5aJmMp1OWhsHaDsmK0Lc5jAPcZleq7+A2pxt/Ui
70U20fesvHkdahvRmGT/07Kvo9U4dVM6rDojk9lF6IOatdRIAasOlE68r5Jge84+BmiwGqJkTFw6
dm9Kl+im6SUPVRaEEffH6K6gUQb/DuV8OCgfcQmXdwCVvFVAx6aJhUeUY6MALX91eYoRbhFI4Imu
j+rmOapzpaT+C9O/8//FUdq8RRe5Or5urVQ5EYmjHQ4wjR2hvk2v9k2p0U5wtqnKX6M0wWlEdI57
lcRWqqAMs3tThBLaKfmdJNu7RSjwglzreYiwuCSEWS2DvE9CIFMJQb5pfmPOFnt1FcfdwzIzSlRf
EEXG6XFjf52vI/tud0/kGOjPiGwKb0lXX3gMr89eqR2imALoehNwxwV+ABTmLnZIj/QeEeohoIpj
3FG/HydQ4vkWmcIu9W91OXmPHC9bn+CNmeR1Zz+fKDP76cwVV4hNqLuD01LmyJmXuL75Ih4a3JIm
VSOL/lZKeaEfFpo7D/w7Y5j1P99YuMQZqE/dRFTfBy57alw9qfCRdxsPoBHqg0zEgHCVwHJ+9qn/
y35W29Au14kRBdTo+7fKEz8tWHjxoUS3VpG45AE+hIpNxThImCY7WH6zhVse2Mp4HFmsFP3QYIPo
4UbDIX4agLjrM61t3DO0e5kHPXUJ/pX0gT+4hFlBdgw5zrw1cPz8IscgYIBOAWx9bKW8pOR2gC/A
A8JwvquhHmPdVsAC8zzwhSbhimxQa1jpaD2WcmnWftSv30HWg5yRZh4Zm/rgiVym782+QNyfdYHR
eJgr0FiWw9lZ33Tm9FHV6zXGny8DYXcpdoQWG71/QNoGDgEZxr1bNBwAJMW/ZvdumzlZH70ksvCQ
1QeGxZREm7z7RSNYGRTWTOmqEfrZlXEBltq/PoO4a2YkK7UQjoM8fiRpKcq0jkXbZdlmffi7v4DP
54Uuq6dXjdMAoMK/jM5HqzVBCi4n6CGzvDbwyyENGPopfP8WHmprtzQ2TbA0x2Z2Rh+CcIA+ImKp
cPnwrs6lqIbNaz5OoTpSLEahQrKY+iDANMjfDEgSRE/NMh83WbnID5rxndHsyaxiHnV3OZPCom0W
Wpn3HyFXcRIMIb2ztbIuJogdpTCH0Xq1lYJvpfnoVgW09Kq/wHEf+msyHDtUsTAYAWhN+5NQnol1
IYVlLZ5ccuaNJawoO7CM5v3EayWyn9ixOlMLPQqlK8Ygu4YHK9GlMQZepTkdMe/KBnZE/LGr2M0q
L5JDyLVFGsFvxzIdlHa49NlkXIRUM3AAXch/yEy2KKN+5BMt6ZqqnpJfcPobkKB01MF4ORu1Tkaa
AiwSGY8X0NocLECzQE28SIS3+aWzYvD/i27HYezW4ES+M6f97/ylbhcYuvngH+zKbtWUc5feI0EQ
Iu9vZkr/Wp8v/DaNtL6gr42HxKtCZX/aregab0/ngYIyKL3of0IgflokgKG35s4Gg6nMjafgKAwQ
/QIemQS/SkhHUvZZWY9ix8SxXQ/264u66jaaOqD2ctFVviezqspqZ/F8WCa/SwwoTVLf0UtUwP4O
+3J9Tm4MNf0iJmqiuTrludl/Vj9qJhwPRiK4mqXgwdOYunA6FhiDvQS2aByIV6N7h/UibNmH3Ury
8j2dU1zzhhOYa1/jZoQkPUTKydREIkbYlJTbzzkrGFehkiU4aW5fS0FI9b+K6pES7KhGK8AJTsIp
L6puwORsAC5BZ4kQLVgngU/4pEQG9VEx0OJnYSpt7bPNQeKoBaCWUdLOK8UY4Dqt1g9za9Lyk9Dz
lmLHF+7j1ISObrkeYhOPCT9geYVORvkUUPWETy0lLrRlU4Bv3aXTV3+Vg1TnLgb0WcKNvU2XMMTo
b3Yvmfn80BAc5ukEqG0vKSg1fmbLjTirgRvTwATpU3v+0z6YxZfwvV+Aa0ZPr1UtQ5izcuKZfo+k
UdAkKsNEi6npgWBfmj2r40/1F1tcmH/EuRQVFf6BeG+9BdSbqzaZkxRAaYJFNlng5ilNCoZOGfZE
M30DGikRMONXtgTqfMp0rQGkVpMtX2O0SVTkhfVGfcp6Hb/GF6Mnsaa0q9/ML9rhiYfYsMEMOZak
k5plmfZyUBrIIEQ0ZcLU7iIHOilpUvX83BPUFUQiEt9FbrJI0RVgSXACIX/GjgsHk3M128wp2msN
s2wrjS6m4b6vYalFQ4w5Pbb24e9hIudWYBbIGwqP/I8z4mWJ1BiPtvsakoQbLljRMlvIVaoHeYun
LLv7GJC4BkfdVBQZ5QpY4erN97rxUbBMnGWGRaJ75V9eWbc4yKnfs/wrGM0lL+QC0BmSAKn5911e
0izmbyR7j2Yk5j9MxQTBJZPiaMiOgE6+yedliPYdUaXCOGPfJpoUnilXn52XvZAiDXe3vpYn8c/u
uzkX638cKNvA6yJPPbOqFu0cUiow2MQ9YbtesY4aa7o03I48AcvFzHGgiDr1VcxTo+M+bJISJH0L
tial5NmvmZXRnAvMP3dz5Wu9HmaoIpfBn1cVd9l2GbCJ/DjmI5ITc6c1k95JBcownHfJJ2hkxyDd
PephBhjNNd/3VdspLHySeppKEPRPK+DZXeIFKyPTKwdrB+UFAInGsTCc3NC3D1R4l+iXmGGj3QRv
6tXR+0uSo1jFajxs4VDhHzX3c7I4zQXubIKwkxfB3V8dmcAZyjpuyPVqrY1jewJxeMlN784KMFJa
HRv0VI6HX12zi5ADjy1iQaqWTXGLHQqHIc4bNeBSIn5oCV8EPI6wJA+Bhyqmrtampi+EKpbi1QMG
h/yNUZpT2+jaccsxK8nzUOZa7BZ5Owia3cXxxSZpnlLlold4Zi6cWWdUvd3r3EN12/KV0/EiPz5K
wOraKpcNu945Ti+TqRfCIv9bUafQTwiSpPbv52AYWrv/qjScQZxoi4YU3lsiRRl2dLOCeZFljTZp
Sax+MIta1M8u83sBRcO/mFZ1v9n9Lvoj1uzHDiag4BF7ZJpQ8V7TGbU2kgTge9sUokduKp/VA3cB
L72YxFEWWb8fKSqP23X/PdWakt9K/R2DHl0r5Hjqn7a7ZA/xiX8k3ocqNDvhC18P/Z/Gghsh37qJ
EiwCajuBNqDDLhAHJg8Un48BzUjHH+pZ8eJ8Ak1PAJRSNAgorEZTyzz0Ft1E+UOQvBcB5rHUVXln
VSr+9nv3TafZ1Az8GMvKeZ10W4Ef40gU9+7jVt71KDMW+SZqiYGHq9WvrK8wvPF+mbMoc+4M3tTi
lCaA0PAthKZaJHAbcrZ6sxmiVjGBrLyrn4R38S8EErGO4uXZma+AKf31Y9qYpntqqDjIlKnsxW65
2W9DgzoZNsGgtF+v8TjsaNdnEHNaG49H04Nt+s1n49cKS/J1io4TlZOWbEjV9cbL0ndtWk7JAXnb
m9rDv+TPEH+KTUE6qF5dFoHPtrlnX/85rLK7ftZOGC+BLE3R49xZ6Sgp58BmOwjZXtjTwfRQcVAH
LT8nawArjm2Kdzbg9tCCFeKqLg7LMdkhywnAVGFj1zbUoESwX6RA9hmXX/K9vjVQAXhGo/+N93/l
CZC1SvdtYaz+379IXAcRA6+JfcRTEfzLoywMoKOWPXSG317NlG+Ayvbv026y9LbxsEXXFCzqwJAn
wLvq7GocUIvPKDD8cLlE1CXZ4vNeYnt/O0edjtSLaKZ86LzCEkqsNiEOwc29jYlYOC1rTkfqaExw
PVflK/spSegTp/5x+Wu8NUaLtJbvOLIqAyEk22QPwZmQdJv2HChCR/yxTXs4HHcEx1g90FtZUyRw
VnTHltuFV9hDFM3AP3NKFnADBPgsVWnBLNoYBXmYgl+yK4vdeOrXrayxvBe/SLu6cM6zfYQeP4cJ
gXHLl/8dZUKB3gL3kWoKk1xDDcBGihgd6R+lb+ZzQwvVm2SWmsZBhZIEVHVTrqyegwW9pyplnSis
AYWAi/4YTjqeIG33xww6sslTrcFGI5apItD+8PpIokzJHaTocqKpXOuhiCDI5C4IKq08X2yUBUB9
QZrjikilo/IVRoQtq+6ypLbrNQ4PYIl4DLMhvTGd9cHYM3APgtUjG0cpZrvWkCXfvUqglnmDTsDR
YxRRaw8i5DRKrlM4Qs2DaLNFkRjF5OB2yrO8k5iawXrXoB9RYYt/S7BnfpqNqFkmQDM5qY75RfqH
mGNWT1+9EfFaBolBDem58dsmuav9trwlgU5CL541nOq+WGo8zsGGMz+6sWtqrdoEE839V/6+RS+z
wJXc5ZozyfbF3AdWsamxYHPma1V8sB1JAMWd6wvVdrpDnKbyk9fJaZ3ja09v0QjgSUq6+CepOLtf
b/35YWwiHtK/Sg6xu8mC0kBxSgapYZ1Hk1IjJruVMOAmPt0LOO3lhKIcsGvRQNer26SGA5BUnV3t
Kh4Hn7IzFHOqhUpuNhcpnBlgA/MqfRjeJ7zkb+wGqX+GbxpNZpgTjJ32WUSTq//dF79x/H6ky0n/
YopYsGAbpFn1btlFgW4eO3a+dxl88tcfGWvj8PA7mBjdw4EjbpxCcPGHVhiqZAiQWe6vIHa5cMzS
sYV+tRJ8niUmYuf7NmHdjFKft4lR7GZ3YihcIAdu4cpl8h64M0kmY/lxohL8+aRzzyIYsqqEx/+b
VnSFjP4J4IBUkzUUrodhsy84qSRa+BLKY+ickJr2cWS4ukINqUJXyQ6hzRdfiILiET4iy0dFB1gH
vv89yv62h8BE8WPWvlEhaq0pjoni+nFzFRbZu4I3xywnywO/K0d5Ihcee1C5JOiPfnRhlbXjMrNq
ZxzDyuRSZ9lEtya/f6ND/6Iy1dhpUSqMwfcQ5DXT/oF8VZ4I9ZRYqZFwZ1Fo+Zrn0/+ViwfrhAmV
4lDx8N6WmjHoGKVK/sw7ToysTDp7Xjqt64LiX749ajyLxkKJyLeL8DkzQ9gS4UYqDkerm5Ia9M5L
LuizdsKtroxXNvgMtG4kVEU3dprfKiQxsmt5Z/hwKYEWs0vaw8T+lvX8kIULfDiHvleVYzbX98F2
MlzPQk8MLDIgRt+2CpZGuJhROyYSEvdpNyCuzmMythC7HUoovsNAe6fd9EHv57btU7bbxLfK+P0t
2awTSYAivHddRlLEU35Xm4Xb39T0OH78GK6H9518ZUoFwn1JZikb3onWJN97t2qsSRKsc1lsZPGP
hBCvHHj7J0+0UPCZfoDEy54PCRdrbgcCyRpEZSM6RFyi+KwEQucM7Bl6cigVMkoU3TQLeSH7fTYS
KCd6Ap3I0ETnlgbyvTlaqNBh6igv7ASZEx6PmzI8xfUSwTgl5H4kU4PQ1y5zP4APK4sJOniJ85RP
kO54/tMjg8vuLP8cS4n1stOfLwZLr+48zAFtOZc9i2vu7XdZhwcsXTRq+21gyQTh3aw6zXcjQGYA
qXeLcUFn3jw3NYiwNStZMQgik8hVhyppY2cI+9I7Obfk+/zzypVPs3bAtYG6ou6aJcWAOekgQqVu
h9av0bOFA2dNL7pWE8paTqnkuN+gtDeqtRAvMubArZi+ekYC6V/rKYLiCkiyg8W3kcNG0yzUWc1I
6fiuo022IX3yvoYg1rqeBe1QfuVbgPGHymzFIiZ3eKQnxtuaBCb0Tv5xB4yR+so/znfucCnE5uSU
qUgueHrwWJcu3AK4MgRJ7rNcByM7pLXAVjXfJBOVRcfywmQKsQ8eusMUeAa5+cU3WSXktr1KIFIV
n94s7ZcH7/HBDdMjg9CVrcqT7KrsRZOSpKSeuHxqow2S49xSIAamUhJqC1z9ESna8lSIHadKwuUM
5qSriTVgCFj40rKH4YuLgbh7PQqqyIsLO2JFGfNXvmn9p/FTkAtS0QSemgCRO50Obuit9xbJzGBi
Xx47UFL5oDdHi6UxKlFqv4IQxSidrsUouakp0VQMZBli1k7fjStAqFLAZ2wtghnQN3WNdwSJDVmT
8uR8yWkdCPXUjYb459kE8ROQaWq35VJ2ug7yBtaYDpbHpSF1ImUsNnX0YyNPWyLpRVn9C7nPiVjN
Q0c3uuFqw5yLZ4YkMgsD1tFaINJmrxiZ6KRs8bR7Kdlgjzp0TEAn/y076Q+lgJzpPbAHjv55Dfha
SYGIghNDgSaLgRrXFuXw9aTfhYJ9W9c/5GoRZoPuhTU5FjIEHJ8edeJn3XLoKvNvEE5v96s5MFW+
zkQLIsZSWkOcRlwTpU8XcPkFhzN/baPTPT2LSOp82F9SITM3C5aQTuqXkn6lvVfDTvtvyUWpmsbT
1bQWO9wf4YW1TUQrvj7yhJ0jrpVtHgTRxfWD2hXeR23e8hCyzUsy1479ljQEbaUoooUm1YBFNYeh
ABw7boqNzgmPyKlfQ6MP4BFlxZHrhqonRmqsBDVIvcSfM6VT0xuzTZcg7BGZvDE9ASIh9Zk2hZj9
rctbWrd2DdlPRj9oGXlX16JsbHfOyGFrYfXcK1abcwd8qRK1kkgQ++4NAN8A3wHEFWf+bp352AKD
CalIBYb3wce8HERhqMfQnnBaalqm9H4OEHh8v5abEUu/UdH1VDVgYTWJTK94ItHzki/D4aJVMPXn
VHTgVnrv2ALjq3IISnSwcBOzCi2LzN82ARj5RkO/WlUCS88KhAjKzRCXiaGQB9eFTFzoXO73nN+b
2ePtUQkXOo9swUgNf0gyN/3gAMwxgsHCQzmEvDxbmjx54aMhiy1lldNPCO6hmJOMfzPrBN4oOU8Z
LrutH+KoX5W9YJXky2oh19s9bEb+HPZHqXTcrz/i2WNT1Vw+q73cS4i7e8Js/sLyFXxO2jaAbksJ
25g7oH3haHkNuvEXJv3oidzgONiKJsM13KQHxE6bn5U7S+BrIQCTZtkVxnMMfSSOQdklJVJnWtz/
o8jqHDTQD3H3lhxzZ9ECQ/7UY1+rqZj7idpi/VKzOTKwV3fnGTenYn3lhksDpPTtv77t/gMu5boW
eIW6gdXCCsUP+fR+iJEesIEahmQa8oHA0pPpTUqnaxDasaq1Ko7dW/mUQFFvkd8mtbPs4/Zswvhz
RTtgCfFXR5ACgEggAvRkRWjnFJKGp5j6kVecmy//R2aEBXNgIgJqzgFW1StZoqQDPZg9i4masQXe
mdvViFihngTm2uODm+RE0MXhQqF5HU/jUjOFdE22JeN4QR4wnv3LcFqhgBJq/d1ngggu6ZnPciSE
Ev73qGhKZR82lEnzm8pmuu2Ms9Ifq0exLsK0xu5oSWnqI/LO13nmgjuwIVJjJN2grHDGHC5Y0jnB
RHMmp+obkX/deaC4hpvubSfO5jy4JAN9XkCl1QVEt2L7/ga4HPCZLsEz5FD1pTyDwrOU+CHYNazm
7HoP2oeW0avTD0+zguXEpfmiFrB7l7RcqSpC3wLfMSNgRnb3zATyr7Vq/8H2EesnDNdud7fqqYZZ
gzfAFmlkjGxwBdRoJPpgMtQs/xc/NkUX9YmeiXFgsMZ1cKQY3ZzWs7vhXELcakNlfr2NMT4k4mws
KHdtCi2jn/DsRIRkSN6fxBmXbirLnxVR7QjHlkRLrCMe6MaV1ZOIIq2cw9ScfR1WQ9NtvCGipB7/
Y9K+2mEMYKJ7q4D4e6otnD4aYsLEtErABQo2f4WVr6xVGpU3V2HfylOeZ4VAkpiapdaFkELsPw+7
qLNHR+eqr0y9eHgXOW/OTUbN/GYXPKGu0GcMgc9wA7kL8zwJtwfGl4CVHlXI9lgK9nR48Az9Buug
7/BYHQr0O3dQT3ps+B7yA9WclRNF8a+U9sJ/hYvR8S9wGG6FUflXNCtZTmN26Ou4MMknppCRkGR1
j9VaD4dK/ONOdmYFndzxrseqJVNZvDxd6+wxWOl7PwQKSJgkGiOBW0CmVTLN2X3Zff9nNh+m5Wpi
ppRuZijBSUIXnmI0d2JfbBXe9qyHjm8DBuXDQv0JH9B1C+gnDUFlUMrVssZucgrCg87cq+/v7LWO
npNaUmomswpcTn91p5fN1zkekOwL1CkvnO2L2DhkCnUjvUvtxa51AofSYEGBGWTeTQmrS+3wvqzf
DIKNqLgxa9v6CKxUaIRuGp8z5ITOP5DM3HzcEho9w8lsObkUYXbMJad1d92padCbht5L4nt2cYZG
dSLQoPe+u9pEDk1Y92j7T8Y7rslVbalL4YlwFPKOKec9FA08ekxa0KjqXZgR1KLqPu3a9vRKqDCu
/Xr6rBKDyM7JpTDrAqzFp96uJ3OMygyqDAHwCuOpiYOjs6P2359OFF7+r/ArKd4fdzDcYC8PBF5q
mAWb+OzKxYub3cZgUvjEMUtBnkoYmZoGZvgQYOdDUQmaYRgCo9ghfGAORWnygbtI5RPCaebfCYzd
J73aIvyqvHXNnp2XNqq72UtaRkumolGB9PXD+HVKREWfj2w0izwXLFXwqPJTibfMPxGtJoYHWWPO
qKavUV6ZaGoThq8l171s1t/EkXaajEQwRCxmmXd90nEy4IynwymRrVaGWRoDHQ8mH4/C5edYaeGw
iWlYsXFInwGUGXiq6ZDU0jXGnCawLVSMNrLMqOBUg8mO+BNiA/Tsav9WzwOxrTrZY0Ynrk8PfQml
LDPiwR6uqyNg1/y4VW/3hUAP8Exk66JH4cgDFl1BDTnBo/gc0vbNW/qagymgiG1brWSId6JZbbsw
0DI71fXWYRUiS9U1g5uA75ebBIMolbZZcoEcXBXT2WKaDSG0lZ8gfByRALlDCkU+NARP3WOW8zNi
VbdXhfdOrqt4p8dIxcMMoK7h1LxI7CEVO9T8XTNXxVJmdoyOcnNvHoSfTvAF4NvLH2WICAR7IlXr
1BRbKqPzS2VPVSgX1/8XT9peDuOzGppl472f+vmH2e3GrUwKLU9iYQ0kGhj1ksLWHjUqEL4AQOkg
63nYVvSoqAZYJBtnW//xnX7fMld4pamKMYh/rTMPB5R7To+pihUQcoyckkEc6LRRSCb++pJM1hh9
a1m/JhCrzQC8TTEp7aN7wMZo1w445RLfLDKwgJd1gkqrUucSaAwRDYnlomY0iDZwiCG7L1SJTbPE
o+6nLAmlWj2b+VXNfshON1p4lFzyqn2nZ/1ENcy6SYl94bj0dGjBJZ3G4EHjEy1mhUYpSCVH8iR4
6+rpIoQTWz9QvmQ0McdikIC2JVIHvbzrsqIk3RVVeN83OHGutrbffO9/0bPCyWAPeJfmGOiV2TpD
noRc5x+8FP0ZaXOJzYJU/IAWd/83TdUXVEJyeaE7tmAMHgfB71R2bwAdiAxEv6FinVtPYbZFKicX
raAUsFxAmr5Eq7weVp4h8TRKtYNHH1+l5emXNl5+t+2vxNrkL+skEGiTHWJvGlw7U/+xC7Ew7cP/
IPKg3hyZF68a41eK7SiWDRYijVvkQkQ845BkQ+811TxAIHtEPEM9UL0LnHHnIfN/VNDye7XZpDES
pbVEDF2xyCoWcnRCx0vaWG4uWL1u9tLDv1SUnv+SSv9KFNF5eFI3CbxT9oVMG7L/vL8gD6NUB0P/
+WIbImTL27rHc7aW3nvkcY6Kc9aq42NJlYlaZ06/vguaooZQD+4gCxnjsMGPnRQ809KHjaAHXFdX
rsydZsltt7ad5MAbioUt+wkcfyHWPDAkpdvOpxYyFoZl+JFHfF+L040y+8TcDNwpBPuAWJHOtldw
NdYX8q/AkzUIrz61hCisizV9pzwKL7IJ7ca7cViftGzAKwKaxCEKFX/iAMpUPuCFb3W0mQ5nAXeq
XDft3oUmoN24foP5d4Bs/d7OXAiKrQs+uyxbJQgebm38Fk3KLfzM1x1PrGXKqUJ8OInUywELB4ux
Flt3C6qGL/6t3CZ8Kfmedxq26ahUnxs3I7ZtbiJ/YpIKAq220aMFFZWMgSCqSbf2cokV5AMYzYo1
XIBNO5d62kP5Hxo9YD/gEon5P6CxKKA5BZKRw4uS8YgIxxPWGOViv0EN0jBr292PC9EU4w7fX4Ki
BYadGyvKN9rHbBCQxvV/YhNw51nu/ad6Eo9wLLtZtJ5S1JcZaepRLGbLRuS3POsGIz95N7vyDtvg
KJF49fkQ57ApxQvmJsnZutMpohluzcgycDHT/EbM3ssd8t6aZbGSAOEgfacBu53kxG8mDIBXzson
PVk0SYEfa36Yjhj7hU2qcc574IAdS4zy3nJWnAZ0foRGWJazF1OJP/7H3lWIfHEOIELzL4cVnh0u
1GdBU+ZaSmTldXRE6xlP32SkkJ5jd8anoVn95wYi76yAi6BtNTh/AL4wdQmDv02q9RD5Mub94Oej
VF2DsghhqB9nzHTjIm0cBcbQ/TsX9Fb1ibz1oTVeupk/UGZInDuwFpS2B5fIy64IezM3X3zW2yLY
PZx1c7fqOdrh2rRCgGHvPOpFu5w3JqCkZYcuvVtQgxcYnkOuYN5EWfUJyb5o2sk6w5ANTX99UiRG
FWNC88dop+y8auY1beFM+q/p0DlLv9/KOw6HugOZ89QTzDG+CRHUe7zErKHlXLnx5yQwRidbJQOf
KAtYRLZIzTT1ASs7OlZAP/yIZwAF6Fk8jH4ALlOuSR1T6URXnoZTYdJEi6M3+L/hdEUQRvEAZAwI
T9YwNuNSmbkslJKTNMzpufqvE+fbhnmy+BMvNEZTYaHCW470RhociaNGAPvWUOR2gMbonqt1glO0
f99NBdiArIoxvhfUD7TO2gYTiPFAOIFlCYc5OLcljcNRHnjP3i/NuuyPOElkjrFXWmq32flnjot1
W9Ew6a+Ymn/LnTfCmXXGF4YtmFIHkzv+ApQGjcFKOBDYc4cnlbI2H5PifcyjFY53V8mAvN/KAi6u
m3GozYi5rRjz1GacfplWiDajpePXU6QAZExj6uMkBZrHtyG/2KWh/+eMoI/oMP96oxtk+1MLGo03
l1mFc9K6Jpoa92xKxnGsa/FL0U8iQ0UuegW46DKtNYBYDL0Qlrh5GjKV2NkNIRugyig9TSeJLD3u
Jl/jH8CMSvJZDojCWXCl96sUfF6bgS+CR9OtVqQ9z4vCrSenG8L7CuJfrc20vg7uNwkrfLPHOZ4X
0TQCQ6LymDBVlsMUlftYKPD4Bt3mo1zHKXGoVFwer0n4LTxH5dfjPSWPw89G+6xlqzLS66IIU2yp
LMwfstAP4v48oES/5qEYQSx/nF2CIzl3WV7czllPX+g0xaNtA+DVnpCcreO0lLq+287MTKrhe21E
VGcoPQRb2l/cwwcZDCnSLaalM7Ig+kVf68YwAqKbTXcoftb6ea02IYEf3OBXn6wewSkT9nhqFHiY
FQI2BuzBVHSfkGNc1OLghMu+xByqk8cmwyOZl/cWu+iNJIUtGG0YrfT3WcCYw7OzMFzzVUC7AZMK
4lX83Y8tAlsD2GYJQw2hxq5GXYEGYRlGDq+wtXJxi43ozszxTF3x25Rz+Zr8q113Afya/ImxHmLr
7Ng0HwpB6vJEfAu6AYgtrcumlE06yDALKJafcjPbIsq1u5GzqPYEcQeg+G9HgdMcyCdxcbYsfQ37
Vb2Qy40SRW/brYmvsS/Ct4IsF1O/AcfdHNFSSOTTq19lwsTUfFJhM+jawnZmEeDWjwGgytvprFyo
A7PY/jJj12B1GBwPSZ8U7v/SNbiE+aNEVLfOAdf+ZlNkUkmT+0Zn2BjvGTWSm8pLLA7B7Dxrr51H
V/1T45cQbtZfSBWo51D9FyCL0SwoALJk+0oU9+P9WIVjaleKyTGIc3InhVmTxo8TugLym/HEklFb
q8ltnvDfpk+DG25VidK046xcvHaum5zJRb1ExFBAAeT1ixA6qge8RyhVgeMdvAIti13zEhDiZU4P
RA/Skr4V/NQ3uXuOXdsuiM0/KsSDl+VjZDU3U2pBPXqSrt4dntY3dfYbck/Qivv5hBr0HYzEZLCT
5oSko9Z1L4UkmGwD8BtZhYEcStH+RLnMuRwqq3aXisMPCTIcnge+ePy6A0/SzRloAYLYklvNSuie
WG7NWfu3gfUVOy4w+Gz/hh8apKtY87I+hpzEQchQQvr96cJCxtP3z3dVv2h/RJX80ReiuVK/MV8v
1usdon4lOCACgcLPWA2J7gQXFutebAd1ea9xiE7YC7nzL4cbp9PH6CHSRUA+yRaeKJnoNcd7T+tq
RB/g9nGRHpv371S0NQ/JEFbqO3Y5TlHSB1gKQQPt+ENLEbfUxMHFVL4T3l+mdUzjOZpyD0P9KES1
LfXt6i9QyYdwVpI4eEB72iNPRDOnfUyozTXTQN9OdKeI9eZ8zxcnVB0bahk9LNK7CQvst3kXi4pE
8hAW2cfbPo2m4UaUigzkkQx35Ab9LN1T3GxijnpyoCWoXbfklHPJNDIDmHtPz6HcL5G1bkpicJIX
ppAbm/YFp/aw+TLozFH4zGyPGNjFXG0CafnkLLIf8wCbu7yXX4qpGVtreCMrd1wzUMLXB7JfYJs5
trEAETAQp9riuxGrIvevSEpoi4DUK0wjP6/KIcVYPqVG3FbeV4h9pgj0kAlWekR4ClZeCzB84E4x
86UG4v5B2ZdiHfJFdppXrKPCWakEfTm5ytahhb9MS6bNK+tvCHmcogYXvSOXqRnKXTmjvwIfa5RW
obsdA/MF5pblCDmqVK5aJ0ONWE5z7ub5S6HjQmWxh6M5LJsUW/LtpYPxEyRbtpHLVzkIlGrkkiP0
kb6pGSJMUnGQcRbWdJYBv4FdC1xXoMLnsj/PqJ+2kYGT7cj6yQMUI0WOkkMk6ehI/W4prNwJBcn5
/+gpDfMo3mMQ7M+hQR0SXbISeR2sfS6Vv0+XfymeqL0dNVDFwAE8dNrH4FB1J8IIf2m2x/3GndU7
BT87ZvrKt+ufvwqTDd8op1pjTz/23wuWCiqsL+//IzMRIFuSCLj0Ew/57rlUm7HEHMIOv2zT33f7
1/ZwHTS4WuTDRXZ5kAEYjVLAPamoBRDGq1JokOTqhp8UDCh7eIfdk3GYoCKt3ymtncZG8/lo37W7
QonjIynhPKlNDSXxkstUCa/kqRIPXvbDvXu6ZHsy19ykoGvrVVcuuC2YmYre45ue3eON6S8t3Khv
DTFHM8niBRih/nMwFraKGP7EoeaParkw08CKrNeR85SJ0wOF/8+SmIm59rWDhbPPj5dRZywLolCd
JjC9kivZS75VoIRc9SOifeDgCgQDcxLF2A8EXpjLtnTXt/8MBfFlXiJJS+m6+GjvCSIhVSA/l1LQ
ixHGtbkdaU+iHKLyn8RfZGcaSRr24Taa43ciDmjBU1lGEKgPdp0/vDA8uTblbrJnCxxbne9ZuE5N
DDcuoUebfTO7ly7yRt/uOYqQS3/MfFmcB4dMcTwgKJyUeRX8NLjckODImGPzHplRst6p+NLOOmNV
SwBTIBSylmig+W2eJYSIfZcbisi9oZmHTXIVBZwQKPwmPAvohP2k7zVl9NIMydPhHjtNdjR5V3Wa
aX5pKrNlDW52rlU8OCT13OdykSV2f+07Y8N9ja41M85h2lwNqTNRKZ0PBxTFtqOZ3Sv0LjaHVWim
5n4huWvxLUINk7pRhMiJJuPShCsSs7jCgk3qu9dRviAjSicMCecM0bNq6yBHYSZC7aTGM1sJ2KKt
DiwWxn0LVrQvPiTQs1McNzwx9Vj7tmBzkFCECKQbaPpZ64oHTzfp1Sd/mPTIbPAarjKirRV4NRhC
TKEHn98R23hu8fthatVYnmDwPAtRUPiSyV/CdeG/lZ9N1Bg81wY6pQIDaHCQ3/PbgAoT4i5P2bku
7xGItURtQuCQdnmvO48ilANsbh5+zZuHdfZPguBY7QFw8PI3MGbBAzifOT2MTiT85vvrwyE9se78
5qK6iP3XtfHyTKiciALMrEm5lXzpYnPWE+ENaJNf27Hezqk8wk00Io1cTfQ22nAzk/KObdonTIwq
sfgSIpafT/MSUEWzOtmrpL0Yg/ISd9RPsFGrTYTREO/2pH+aWCqKFmsYhE7L9LpWb56OpIzd3JVe
KEvjd6jUoI30EyqADIy3XL03kk/KUWBZQbaLpZ/NF1eQaedK/ivvoF+3nYAo9eLlwj/C1kK2mFrU
3s2/oZtjmqch20UzFvkc/R7PJZKAKv8/hNcSnLZXkLcfcVZR+gJmwGDZ+AOGFK/kd2tKh2FMKTfW
/XuF0zM/5xrmBkNg0aHPnus3B3rKi/BkKPw+yazS5fZnFrObB9dtM7yOyfdjSmpAgImhGTgMU8MJ
zWHznvE1UN+yvGeTC6fjcekxsIgjpbCyomF28h9NcyA+oLbjeOeAcQlfomaCTp0of8FuvOE666hc
TAfNHGOYKNdth0I0ubvsRmn2SS2MHi/cVO45GfdHokBR6vAWOfRzsSCIUvqhQGIkHVbaCA6lImz2
tzXeRJ4nlWJQPD8hjduss9UI9tmlkJOOKtcWA0Mpu/MYfr9RqLHaISouC0O88WWS7mFRHuAVmcLK
Rd+2L6lEESg+n4ciP4Au8hCE8LgWBFT9cy7YX3345+tpoJAAGvL56KKHuDIAczkB7SXdI/jgTwMW
W/u83PTO+PFAQZ2QtayoIdYtN9NaKq+MDr3LeE6TPJL+UHIWBy9Jdcp6lAimW8D/Ep67wHAQEbuq
rOuhWl8UjBPIC56opIqcpde/GbIVhXTR1pE6wvJIOvisxYdradsOhrKhp22nVYZ+GP/4c69CwUOl
R2i3Wfgza9pisdlZJ8xt5JtxAs2mRypl5XNcSRXPBjzN7A4+VqSDpEj3nVp7g5HgZO7x5zz75IAo
kpWsFYx4lF+0Lah+L2YilrRDXCbNnI/lxvVRCEewVVeAK0NqT2NNfFBJNyZcFd131SqKQXNiEyDD
07EXy9tT8kxADHj13uL/Skp870W+36UaZJaQB+nnsfVwNOBEUvHYEj75jh+Hc2j44J4ObBodZ7f2
wfCrOhXjTTNETGAFloTKTdQRt9D8cAjkhnTrXZZRM/PO3f8eSUkLxd0QrRJXjGnhkxtoLaP8Y2oi
cAbNbDuvxnfcAINYAyzNJTW+A2MV+uj29ouAKJSOK1SRAkaNQXaxd4c32b3qZ8t8LFoM5assOKMs
lzn2L4t0qW6xZyKnyRKPe8/77tSwK9FeEmnFYKbajaDB3TvbGy8wpXV0Af2amE8Gs2bslPy8Lwmq
YFUm+7QvCkv40fh9/RR4q7yUKgYmGmthLH0ViGygJLyXSAc7TUhIWQ+l/js9Iay/jwSmlclMVUOp
niGL0tA/Ci7M02U83/D3Fi/hiP+yBjYCx/9Fa4OopSL0IVLz4zQdjhJ7FwXZwTQUzikVlX3yAK46
FTYH9PrL6VUSPAP38/k1obCCV4GWEG2xVWIOLYtD7WQbhcuB0rWrOPmCsD2VZZJzrvG2UhLAo9eY
TsddnI2alUzrDaEd8UgMrZXaD7cfUzXepa4LBTBUKl7JRgUGFrGPuKwLxB/iSBe5WLc6DvvIZ7Hj
98C5NiIJ6RD40dmA5WIk6nCegRkYiCGY9XUt0SwuMVLrttSSfeawfQxe872SxQy1ZQRbaS7j/Fml
okaoGCK+2TEbu2dRaYie1CcyLmpvrsAKd77RtU9cDjwfITLBqhO3nc0PCA4EBIaNkKF849tgwVga
naAYG/tgXtMEvLlJWJoHofwIHkOV4YZi6c2gCQ9tSAn3m2Vyp4MySqXjEBT7WQy9LXrUMhG+OPel
3AarOMuZ96gqq7dTR+3FK3UEX/wGv47rZDysTmayjmp7kCSu9INej8jBoEhG+5yjz1Gw3Yj/8Hn9
5B9rJ/XSLU1d0xHxmoZj7r9u6onhn+bAFHrxTEm5eHAvw+bAzth20X3NMRRE0B4sZAiplstfGGmM
Zp3tol3UfmDVIEJH5eKe9HBbdLd1CinxXleXHURgjtAN6tSBCJx46MgJxftYG+ad2q7nmYuiWRVT
X2Xf4WDMTc+Ae+bJOq3Pif41/0hccuiN0FE4pj28oKKxZr71sZpFEgVXICM3vCghCIepmvnxybl+
mOHHTfqrSj32PXvoPOLNTHLWcGoleOTUAMisU7xAr0ShkZD4gVjP8XKep1V9g05Z4RZSI9vGm+Y7
/5dSJFKu5knPrtdw4biJDf2iVcdYjZOPBtyxpef9O4pjWv32h+SL9oSeG4R8ZB7/AxJA9vIZHJbu
82YR173zZFIJMWvbm+jtl4BiKv7CLz3I0Ho4wWPSvEI/tJXVyY2ZFEQeCuB2l5L7QYJbV+p5KYDA
YdI9JJxBIoDSv6AJFhrOLrHI1zYRuPURzFyeO6r4gFxZHAkzJi7tA8bmyB1kTfe/ZfbmuzuPE0i6
HijV4kDCyB4DJgd5mERP5+psewU0BUnx6YLvoQZ2METIADjizlRtlRnS5KJktV0LNw1N5DtZbTg+
26Y6phUXkBcMvLRI7xO4Aw1qx04AqHHTyEn5yrfHoD5JIA5sX74xhAz8tX2AITXXFe/7HRi75XZu
8y7Ap6EKmw1TD9wvRZGA3s9b+M+RewF+m3fcmyMsPLlP6ji36L8q2NiRwCAeb64LTWeQvfUpp0WQ
mcMnIxxVh3A10uppRYKJi/wr8ATafpnkMBGrN6fzYS1kC2ZWxUOa+VcTfuSzkTHX5glQkaHu6RNB
eZ3l93uhhcNV/s0my0J9Iz1cUbh+JDqHjDCjwpqoEcG+b375YX/wFySpv7FGp+VLRzBaIUvnOpLc
CroILse+D9iFbH8q9p3X+KDeWtUTjVtGtuJAZ1og5Kzh/8Jb1JAUtvzBI4uwKvj1GZ4rniCMk1lc
oUvECumcqMl38KPqJn2eoJYCWIJStdPf/6MyVuGamC6Q/i/ARmLqVqyqM/qMo0QZ2WuTzzzwyeJd
lGGEZCaM2TZVcP2n7p07rW4bw3meTUgIz6x+gXeaeGN6b0nrzzJ1SGvYDi7OMKx8A0TQntuZ0lgb
EdbArrjW8BTkuzRCJRC5fuM3pQ8uE5KZXwSw1Lo0IyZCIqgT58TlEm8OkwRmXhPUIeUE3n5ut/40
VZWCdPrbnPj0tfOVN3mHMEWWC2Jf3udt/scXrpMVZ76VPvnY8meKTpp8lU6vKznJurPf0aNLUk8p
3bQUxnTqIclFvXuUI2OQNMI5W4Oxig4++upNe2mCTBYMBNiw8dQC17M3Ohi6i7A/2T4Otbmv28Uf
RQrwz1fK3vyc8G02PnWv9Xb1zf9vadsjR63WOvPgXmJAhbPWeXZ45eRz0hSUp/FfwS8kkZGIyOKI
FK0RN0Xk47t+pzUsj1/IB+C/Iod7Es2wE6NJnjELJ4nRQQgutxmbDndSl+QCfpbOhCyS79qxxhDZ
mJJM43VvGN+mr4g7iEEs5jidCob3VCMzaQGJpucsqb1Zb1PLldlOwipnGVbuvd5bdN0ysbPRIH3a
J+bin+wSQhDkHCbueO1x+O3aQeq5SkUl2gTEP276yFNIT9Oqjrxch/XXU7yWYwmuatdCniRlggOE
4SiQWAauahlflx+wUSaGsgDaIOap9CYmkskOSadx08NEFGsbyoHvm33/ZscnTR3GeaWAhm2WBhcm
+CdwUnLg2cVnmv+eNHxJZEykx21K+sFr+86qbba42KxcUWVZPi1174x5ZkjW75rEA4wF43sFCaDL
HKo8+TsqC1kESlJhA5W856EMCVYL23OG782vt6tfGlzIcmyVbjtcHZT1BVW+myx5zLkkyer83izm
q7vI/hpg5xD8wl/KZm+QdwIK8/B4MU54V9G1aeJYCSNs88UycCOB6wDXroRQDW8BPGbnXIdm6gyB
TOWfMMJjO9L5Ee2K/HxO9kwOp1kCpLDYj5ZE2CKv89zAbLAbqNOruvcoi50laERFLMjyQfemxZvj
lmSjNTfHsCaUyeKAJcf8HWZFkqVy2Ff62fJxByBPJr/3IqB8/RuGp7nDYfWIiPTMnhmRWuMxotPY
4QCAaBDDOp3fb8Bm7rWey/8KcMFDUHDmTI+T5Uma9vTzP+A2d9b7XP5OqzKXsRA7sCquSml9H/R3
h3B9iR0muVeQlnZdAlXAOywFf/W2OXaTkqPNBi/eEcHaECViSNfyYl/rLi1wuj3nsCCRfjCOQnfz
oX3Fs+kjS3uMDpbNW4FK+XaYYZ+ucclk266YJ2hFyExK909djb6RnInAHKIUZOiYfTZpUYLhMw5F
+UftEzO3b8hsuQiSSgOFSGUouHvzs5H0Iy26UXrKtmNQYELtVx2N5pnXGp3l5CV0vCPvOvbWKJxt
MxuGxRpHmH/d0v4/xo5BEA1auPUi8iMSQycHgs0rp7H6JyOSU3cdNizfEPRZdgnMsMvJSQf6v9y+
/f6lHRrHlPJIC1QoMC3xbeG0REX3rl4577aXMxYWJmQ633cPWaMisEB5iZ9B9Slho5Uc84/Y+/QL
y376TiWR0INbGTpoT/f1fQjcv44dEItZMxGaQ2G+8HwLwq+iE7Cr964a2w7B59mOaMD5qHzICY4v
TMJGZbBohf3A2uP9LYvks1NfcPF9Wmy4n82Gj3aIEgVqnekaP3ekAIRylbHZEC1AI+gb8l3sVDtA
YIzIuftX/UqAl6w1DEvFMnSg0czLVxYY8Uk8gDVgqE5Yy8J2xSRAFRj96noMdwLV/fkcnyoMovOA
rx5dUOkGUJ/rUWQmuYtP+gbIMDDQfVMP8JLUEGrp1h1aqUmJtmVnnk9Pls5CQsUGtDeOpty1/9Vk
8jMlFPwxpyzXRj/6p46zVWpxLGUtcmVKVWN22Jgqy20N4C5j9YtpvZrmZJOXNUr49ELw+0YCjHgh
a4fRCtbjryEB6pb1+bj2fqMq/uP5NV2pq+wmRrj6Ibcn3mcrhchusWuEFr2mP3WBacdXcKI8mLbC
YRACq4vfg+QGzR3QF3hGHylnwcHfZovuWO8EDIQhzkttd/W06mfEuryunGZD3LzDpnsCdLPTm45l
D1h6/H9UtsFgCGgp4Mlrzt7LOHx1LL+7sfii4PTiYIwQ/KzXju4xK7FkwaFlqwUp3j8UjpS89d+9
QFhtzY35G/zKisoy/rNFC3chDjtaYXTHWFusggqfhQpSw5S/nzlnpjaW29GqQKXhFU8Y1HjVwwtu
/LOAnpcGBfwPBJiIyr6bBMWJEYNmif+ikkCU4i206iU7snMopvH+jNWzUTKaaIeVxR3TDkTzelRf
0jdpyqhc9q7qhiMx6pk77a8XVWip9uLf/23fn7QY9KTuWvd0Yhd2CWzYOjnz/Zq4MXB/h7NLCl45
NGk+0gjSpBAFxRTAUUcKmLcWWayjR4Js2JHmaM0rl5pkiZQDMmCKWtAbgjgZ8GHnFhXQjZVGHrAq
F2kdESg/fsrVM1fGx9hulsyUaQHhJlIY9nKUyIvmsWkPHPHDZCEzMZbvBsQK3Dn8sL/TIQqW6jcB
HN7/MMi/aXYTo0Gu21BFC37N6sz2DqLEnFV2eSys8wHU/O1R1JmYH2AfjMcomRWHEhYqj8MhdzIa
VD/BC1AeLRrDqrVqRyBbF+d+2ConSm5dsci71zivLf8O2//FYpqZNSHfJuNMrAC3RsMkfk0VZ2h6
AoPh0g0KqgWUFogu0ud54y4adVZrb6NE+n011E/bbBFlBo8BqoJhKOMy8wqOPHKIQdywKxs5uH61
aglroJKMMcVISAQez6PQFFZgk4JksxWJhVbwan3bCdLfjn0AHD/h8kmj+AeC73Fc/Q/YfFO40iB/
mh7SIsAeRPTXX9yUuyoAPJyYdcZgAbnJXFtLclvpImFkkEfwwUWrp2O96L+uV7Ck+W1pJWVBv/RC
GTS06t7rLhh/+++Xio0RvGqJfkScDnutPNzMaJl2DQKqrDVTP6qejnzt9LBH2tvaBCXed8bzUuyC
VnJBZkzhLR/sUdM9Xalz9qsaMQkeStFPNgaQy8jrlFm1g3wvAupzEh6EEDWkQUTnOPAsKd3YArzZ
unmdI9LVovIkcSCMonboWNlIHO5M3CcY0fP+fzdLjJlFie+3r2iGem5GB9eWS6SxiAnbJwNaaNTa
CKmKW4xo73vnF/Xf94qUc4Iqo8anQoqXNDtr3nWXjqEdzqNT2vykL8li7cSU8WXR+Zno0cZ5JNP0
ZcNLJCcLl5vRhjIrcMo7+OCCr+VZ4CL/FF5oF9X4eKxJIG/Ja4BCFwCsCaZyjEZM1lNZa/OWmsCj
6O5LIVJbWm3gjJ8Daiu7q4aSQtVlp4xuofFtSG9uqkWIYRW3eQNsBElqj+E1BFBzUQz/Cf7Hy62y
QQVJVwfVU35I/w5462/ZFBVdsxwteaBET5jOMxmYJPLrxwQocCZ4IbD5C3OHwkvVGo+fIZxwk0yv
Hb6GQHljlNNzO+LbKNiwvO94IRGCWIEqt65k5kMPQ3HTBxFviBJAQ6n4U0NyP0ItYcr/rYeC1eKc
0IizZBqc8vISrU6LaBX0pR5NwypubSuIDyIXOWhYmAN3eIX9bm9ZLIpQGtO1+awuS23TBKqMDeiD
sSK41oZU0r9QMLaNZ/x5wwE3mderPGRJQRAbi8nY/MY/AmrIVq9NW1tDth6SgA==
`protect end_protected
