��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$Rx�y�<��wA�*;�x���@�̦�W�X�fa�M-$u����n~�%���P�$��W��kYَ���P7�?UMfT��q�6�U��k�>����~�\N�(�����X�e���/6U|)�X2pF�]6x�793�w.�'J���wP������;��y���k*��u��D�ED��8�|߹�G,B
�<]&C�~H�~��4J�*E��N�$)�Nq��J-�l�$vgZ]��X����B�1���0�m�ܡ3��T�00�S��(deR�r�Y�C�6%Q)z6�i҈4O�ם���*�j#9�C�L���a�[�0�P3���7��s�X�~%Q"gd�.k�W���G�Ԙ�t�����e;�S�x����A����9����H,*��U�>D���������l���nT3�g�&�17w�&T���~�#���P��O�B|&��Φ4��V�_3� ��p�ͼD��� �c�[�;8�
�Lu��\_�_?�G.l[�����1�w�=�"��B.�J]s�|FaR.r�e�P��l���ߕƀ��p��b��l��[�/�ot�ك�:u����3�>�y���ԧ
��#8H��bS��/4#0�Tv|�����T�`/p��vks�K�ה��d�l+!b���ES��������yl��R(=(�����d�^�6�);Y��^�:����5󴭣S���oT�8�P _p./v{.�4���S�������*�Yn@���?�0�6Üz)F�ŵa�.;he��e�iit�)BT#��j�	�����:`ê3[����	5kVu��6uƱ��#����Piߐt?�+)�! �K��CT����)z�Z�9�T�x%�i,T[��M����S��E�f�q��&��7��+��J%�� ��Q�^c/f0��Q�f�'(�18�5wE�!��"E�M�Jܳ^���5�����8�K/I�v�	�+Ì�6���cG��;8��D�~qCC!�o���qO*6 YF��FT�5�`%�������UT]��!�j~�jpRWJz>}jb�/qW ���;�Q��ް�m@�ҥ� C��,q��O�2s��v�3{^Hf0N��-"��FPSa=�evԝ��{Zne���7��3�G����5R����Z� ��iޜ*x�����"�O`|��qSs.d���4"�iy���~b!�u,H��+8a&i�!	j˒�"�}n'_�}�q$��'�6�7���r&�8�&e���Z+�=_��l��Pw���>1�br�3�Xd�6=����
�O��b����9	�X0��"�$����{J��(VpT�O0�i�a*�2�6,��C�@W����w|D�ty�"����6�Fu������pfG7���$�US\��C�z�8O�����Սn��<:F��Ġ����T�L�¯w�ܩ#��Zm8�jA�pa��vM�nq�aE'Ӛ]٬�8�V�.j1&Z��	Hp��0��#�l]��:����m�K��	�A�2Q�F�p��^[ޡ�Qe�N������ y���H��U��Ҳ��#�
����eIX=F4�����Լ9�M�0SS���c[�h����H�eZr�`��>����ʙ�G�)�^#xk�)��%�&� &��-:�Jx�����dM�z��)�{��"RW�A��	�77�|$�o�~���c�=;��j�`<q6�p�y8o��F1�6oj��f{�\Z��n'�v�k��i���(����GG�X�y��/�5��<���Z ��w�n�����
���2H�򖝔��E]"�ړ"�3^��k��E4c�\��<����YA�x�:#
��|~�Bz�?���!&���>�3�Pb�n���}�O;ق�*J�#6c�{n}"�޷�V����\��w�Y�.U)�[���]��B��'s����i_��[���f�rQ:S���@���%��<k�X�N��!}��׺+5�R��m�(��W��K��h�gZp,�-5���o�-qW!`���j(��!b���A5���پB�!h/�jO�R7�E�S�:G�(e��p��~�5��@��aRVخ���3��m�W�p��~�D��/1c�ƪl"����iw�%;lX�q����?m�.A�h�mx���9AtK@�=��^mF���?BU�epsR��B��Pc�e�4��T:s�9/[݄�����T�<�%�A?�ѷ�4�"�ƴ�`��q�`�#���/�1k=�/����ONj�"(GE���˪���R$�g����1JjlA��V/�J͐��A������>˖�tX@&�o���I����P.�*�l<����wԘZʝ:���.�}��|,�k����G�~5C�(���3��nr��[n����Ԁ�n8�l[�^���Ɨ#�,�S�W4�H�O �ΧCǱ�6re��<����`Ť�{���23�}0�����7��u��F��_a^̾޴�|������*?"��p�̯q����ϭ �q<)۲�������Vb_zX�p�|��L��E�x��B�_G�jG�k�	���pj�ߧn޽p��F�菍Q�W���I��?�@@����@�pʖv[{0\� �/�n���8��+J�Ű��@�ȫ偲��]��z)�ڊ8�03��N~��C���핒�U<T��q�i`����:�d�{�;d�}l�60|�!����UT�._���~G�s�%���3$Ae2�e�
�;M��	���"�yo�:�|+����hbP���iX�Ef�\jT�W�,=�o�|`�kA�y���Q��A9<=:C�v%GĈx\��/�K6z��o#���je���$Օ ��CC���y�	���cd�D���I�Yڜ�
��
m��8�[3��I�½Շ9�giw�{����`s��x�ם���'=���:XV�^x��t���G��Ԅ�> }.�!�լF���֟HT)��%�� �t~'Z�����R[Hi��e'�x���H�I�v�d�䓺�(ݢm��;��)��@����_��Ž��ͺ������r�.�]n&��6J�����wT/N�eҢ�x�+/5A-�;kp���ߤ��z�{��S������񞶺����f����9J]�=�6izTS��A���A�Fhy�2^��p\|&)6I�Yr�Zp�&�S?/DS�����w�V<��K��ŜG�
m܅�ٖ���ƣ�1b3Ij��`�'g9�t$E��I�r�
*������\SnJo����6f��a���W�(�i�J�(kZ�
�g�y�	#VJ��������ד��]b�BJ%��/@"A���Ԉ[���h�\��y�8,P<�����:��T+g�!Dy=g7��)H�#Y� ���܊{y��:����J�����b�t�H�;����s�/�g(���B�T�$dkt��RŞ����Mv's$��4��}u�,�qY��R��I5A�Oma���0S�;�ތK�2k1��p��	ux�&�$��#�f?�4�$NS���_*Y�Q	�S�7%]J�Q!�Wm�9�gn�_� "ښ bv��5����a�t-5��!(�4F	�I�S"GS�Ù%�6� �50��9Q�_�5e2ǊYSb���bŠ�
�Hz}�=���i�qVQ3/N;���Q�jA7����).^#L�erý�uU��h-V�h�gS �%�w�Ȯ��}�GA�F����nz+0���yz֢;�IW��}X�W��:4�Z�{ew���PoW��[�7yb8� � WeX\�sa� �O+���Ε�c�pG��i����;�j �d3�b��������`"Eƴ"����+��¼��8�j�B\��#�WRd]@<z���-������I2
L��ӿP^��ᐃ����L�(�g�5Z� 6c�R�b�۫���B��E-�X0��k�����~g{����xG�)rT8�T��Z�2(GS�&�o���`�ٽ2ň�V"a������>i��4�����ڧCT8������iLN=�_`Ny����`�)%����h[_�����,�z%�"ٻ3�5�'�@8� R?؏��ɦ��-����q	�A����מ��P���V�t?[�����\�B7�T�A�f.�d���zHBu8����!�4	��@��<���aWhFW��?�3�ԡ0`Db�o�@��S���aR+����X��4��>�^J�+�V	C,(!r�ɝ���K{5i��8S5%��&�T��Z�/�)�����*mnÛoh����@���ݖ�`�_ȶ4��&  2"��:���@��U�RU�Hzv�d�+I���ӆ(�_�&��
nϊ�A���/�:Ց�Fq���"�~��ֵO7��k)%��&��g��Ѐ�D�Xq��ei�, dGc�����)z��%���*�;{��bub������=]v{�x�Z�n�?I����s�\sLO������s��Q5�|�Y���u����*م�i�2	��,B�3��_;�S����%���S�Yn]\;f���N�ۆ:�n�F����G��0M�+��|��i��!���e��ˡ��N�ێ�j�ۇњ������H��������8���H;����/u~��Ԏ\�#f����R�7���y�	^�RZ��>�wc!#h��l��m�K�Ȉa�G�z��d��Q1'�(o	g�)p�cؘeg�u[� �i��Y`(��!�c���`E>���m�K���IDgT4bJ����/��}	���^D�̬��Z�u���:�saB2�ry�v����C���4Z��{?�q�S1f�d L1t�����&$�H�O�/�U.�������=�&�=Fռ2s�xcog���\��[p��w�����ܙ~{	;��u�o[�aO��<m;N��l��YG4oVb�B 7� 9�!����mhZ�x���XA��4C�R��DU���W�f� ����n��"�/���s�p�!�\�D��?�yp�~&v�BDIP�Q/5�h�����C�G������`c�=��7-����ڏ���qIr�B\����4�G`��`�2���ʄ ���� �8�VN�
�]����wQ��͕d	+�&�*y	,�����Y	�Oּ��k���
 �i�U�y�Ƽ���K2.�o4�	|9{]����.����� a�ɱڜ�W�-WKh�2U׉�(�9Ч��9
A�I��# �یp!��LO%��Z���=�7�B9�@��	�P��C��7S/�l:���jez�
|�8��f
:����U�w���4Pؒ�:!�>^���FI�< c�Ǵ&�"��6���x*$�m��"��X��(�KN��sx���󁿺��Ǿ4@�!�p�{���)/�l1�N�_$��w%�����G���|!��D����U��Oe5jH)�B�_�
�!o�C����A�p���ª�E}ʑ�������e�̰P��i<cV�ܢ�o��kp�AМp���fÌ9?�q�2��'M�kᅳ�d{��˿U��Zّg��Ե�� ��$˥���1�溠�0�a<�#�q� �ܒ;��xVK�p���W���{8s��fV�Қ�{*��b��9h��܀�i+Ğ����p�J�d`w;E7�o�Ӣ� ����$e�HI�8lk^���FZ%5hla<� !q��v0�W�5b���F1����ߨ��j��<$�=�(���Ύ]6ڷ˃1��ҋ�q���k%�'o�^1�Qsi3�7֖�T#�J��'hΏ��z��]zͯ��Ҏ������%Ί�3+K8�(Y�!��ƇC��\�M-a�,��b�5O��{�ٴl���P�b�����;b�Gϵbqo�B��g
+��\@��h�p�&����ڜ����n"���yH;wP
�� ��5��l�D\��n��W��I���&����պ+��v���l�qt��/v��U����96Ls��g����|�#r|�L�����4����P�UvQ��ʹ�7X	�J}$�7@��7w�W������T��Ĺ�\��8���0�|m���*i-+��^7�'޻l����(��I���j�l=t���/o�&jHS7wΡ/M��v ����B+8HN>Xl��KX�#�<�9�%h�����~+ :k{�a�#���,��m8h��Zh�!`@��(����D��pP�U��i���<F~�2&x�kУ󩳵�����'�Y0�h��8)V�h��UN6�]���k���F�U%���E�n��E� �s]b����aǖi�I�J,�7�>�����u�1yY�+\�ś���	VJ�7��9m�ƿ)�K��0Vkt�Ѩ��U�|�]8��!|9f��<�G�6&�����"\�D�>?�<� �[�.+�ot��
�ז6�r�ZCT��ĩ�^]݇3o����j���e^W�c��u��ͧ;�[ �z���Վ���H���ԃ�j���^����`_^8H��ȯ�<�Z���|�+�t
�>�����>FET����:f�)h8���(��u�[m��\�Y���O �FM��X��޳>���F��H������XɊj3�7���_���ڿ|P��	w��/�l���{�kzu��8�Kǎ��n����?�P���sQ���Bw�Ȭif�9ԑ�_�Ju��%�{�R]���B_�l�;J�_�6ெ�0P�Q
���Y�O�^�&�� ���	s��^���kN����OIq0�n�pV����T��a�d ��f@���jٹ#^�y���a� 99m��9q̷,Q�K(�s�}�$����k��(�	0���z�+� s��S�i �M�:C.+����&����¡F�0ų=Xf�h����B�#�T������J��PQ�5.>��5GBj��C�h!Hz/����Z����Z�x�����H�?%P�z��cV�rWq�<[n�jV��2~��(gJ�.��=%�"녑F��3j�Nh%/,���LK�������N[�e=%��e8��p��!���x�C�����I��^����j��\�>��&�b��'U�T�2��!�I��/��q�=�!Q�01km]-r�@<4L ��r9��,]�%5�Q��68T�.}�)�#�G��@P��i��*�;
FVS���d���{YN"v��K��d.hBv�%͉���(u��e���~�O�gT��|s�{ �NY/���vj��x���k�,|��O�A�k��?�j�Be��o��>�a�F֜h�	�w�q#�t�g��ݷ�#�5�Dx\�h�J�pV;Z�S��y���Fh��da�dv7�ɶV�a�Òtl�&R{Rxs4C�U���d�l�I�Ti��t���<M��T�K��F�Xz�_��42ӄ�a�sm��A�b�,*Ӵ�-Z[���8����Z}}�c2�����[�z��� 2��)yàb��nX��{��q_c�$�ɨ�I�;J��h�|0�5?�2�^�0�$�?k�`,F�t�:w9D��7g5<���j�k��K?5HP�����6�7A���M4���S;5���۟��z4��q��6�U+����A�O��!u�7�,�N�+'�: ��龳l�2�uh>�������\��!��H�'�:���'Hzd@��?��W�<,�|fYS�&��;emZ�X���7k
�%��W�g������D���+���={�h����b���H\��E���� /|@��K��}ӡ�$̓�Tt�����$!&a�2�7m3)�'5����������,5�O؝�]�L����Q�fT*����	�[�Qr�h7��Rܙ��uD��uɝ�]�}m�5z ��ٚ����?�$J#�ؙ�h�&N���LI*0�a�bZ*�8K�K^���@� �w�<ā����t@dO4g�/#���v.֡8\��\��9qiO�i+{D �6���T1�)�j��j�(������C�-9= ��8}���!@3�#��@9���{>�����;�ղ�9_��M�mپ	h� ��!�6bzq��#-��iAH�u��?�,C��BQ�cx��p��ߤWN��f@���Ê�!�#W�=�p�i*w�2������ݠ�dY�$��{�4�ZuȧQ݈�|��h|���ϰ��q�� 2���Q|yt��,�k\I�h�l����DhZ��<9r�Jm-C�9��,��&��p�xi|&�\����������U����8"�mi�F,2 P����J_Dq����
"C�����Y�!r��-���@�6��P�ԋC):=�;Z�%�Դ�K�dn5���H�$��U;��N��G�n+ڥ���Q��v�Ͳ�!�}��R7S��o����x:��6�R𹆐� Mԉ;V�p�%s/��QIcӔ�.Ґ�[���>\ҫ�o~��t̵嚾 C嬸d���U^�G��aB*�u[rG��%U�n���c���]%���B�����t(�j�I3�3kp��uj˷�}Q3Ŏ�s��;�HOꓩ�/S FUޜ�W5$x
E�����M!�uJrظ�ѮzAc}L�9�c�+o@�Q��M���UͧR�C6CK�T�_F����E�V4(eZ*3��N�;�0���C�N�j�X�b@�����4�¾�_�ߢ�f��� J����Er�W�r��W��*�=2[��j҇&{ʭk��<��y�%���͜Q�j?�U��)�=�����(KX�1�[������rf���жYU������=�$X�X�N1 �)�:fH����s��av�o$:�_�L����S>q_SM�N�ԧ�f%�8�p�j�Y!���|
��LS�)1�͕�ʓ6���1��H��]Ww&��h�