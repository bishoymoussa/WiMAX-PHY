-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
ru8aw8+QSCV5LKlhsVhIIJHxoNc70lSfiwV0Rt7vDYsATqjB5TbSXOZO7sI0t4DtKsUgLXnQasiU
EEl6709P4rH0WZfUhe6B41nD1S+GjxuX6c73W3h8ks4f6h0MESTVtHhAXXWYTCtQ9bc6e8iZMmPg
Tsri9oEswXuPc3FcSD/1XLN5Ok/0LdsvJ+J9Mx+psK82KfQ93zQy6Rt+BBd2WTjz1dTXX9x6CmJs
KvHWcuN+P4xlcPIpJte+vLFrbhEsXa/hTTibaGb4Nzcd1gdzIOLn+drZ39ur4p556SByhNlOfdT8
RQCAGm6BEnNiBkkaURQipK4Mx1641lCfns5NkA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 114400)
`protect data_block
WPFcPGNnZTlIdaGq0G4TVNIotBV3USclJ+sjrIdt3HyyQaBcNJtSpzD/vft+DEOYmGc0pKNma49t
i6uU2o2l7MIF6I5P0J4rGGVjUvx2Cvy2XR/GZIUGT7IlwA/+Sd/DggbeLy1T+Z/va4m97HOWTeEm
eQDAfYBEhjfibYRFdWBHax0te9qWT/7gE3M9RgH4psvbkEULzhfi17pxEAzdO9Nkd3Z+JanEHsVj
Dr6H/suEuQcWKB8z8nQrPCcaGmowIykyuSQWzxXQHf6+0AcgueYn50UZFaYLlEQqVJ9ITQSJu4Fa
mWiA3ImA3Z/yvaozpC/UVmOXmVG9Sl6JLHWKsekCVlOuTsg7urgkCvKOhqQThcPYRGktOcvYqHsB
JWxzuGvOf7WiNVOT35uOYr34EO9ZfotZdFc4Md20q4qIYvOCZreJQOYnpqs8mJaC4vXE498kczm8
h6sXpCvASfgYQ5k3kyPodSNH32SlyGFx5LTEX+Vh2MM9K2rfWeQFfXZOmvsPJNYD4zPp96efZZbP
Z5Pt7pkAjxLACAg5HRUgKBj1swWBIJ/AJXp4EvSoDsN2+KUwvbWJrnaJ/wYGwUKItOjlo/nW0Fbx
mP4OFNkDy0Cac1y+pnzTttvaYr6NKN2oMM6H78Psgf1ou66oWzNxf+49+UB/cm+PCdA9CSUTBCS2
UhXu3KqtTMMonyWQpy4uQPe8X5JQELPL2CRn04oCMYxHp+yF6hXCP+NzCVV3ifUEx9niggAlLxGw
UhTCcs3J+UxLdvlwCDrA56jekQguNHeE7Y0zIpC4ev7VIli4iBol0MAv5V1NmN+xtCY+qiB1HSo9
PqEjcQsqLicpKNEYruyMVn2ERQ6ExH2RT+50AbiOH4o56gxf9zA3JYvmXhcPukJVdzDOcFQ72P9u
YdYZOoQEQvTvv+AbLoirzJTUlA3h6+M1pkRrhb2bfBIVuYBxa1ZX+Y6U0hxo+Gx9dzMRW5KMIAyt
Fw6FiMjfr6SPZWdCKdaGEt+0J+hukCnSf8fdlFRD5IPHNHxPdzMwsdoFsHRjcVSaWy/7EditdWVK
iaDcFpAlO1CfVUWo9o49hBLV7EbMiWQ+1buCHuS/tKMA7ya3ss8T1ZVJCUfray0SDOc46cjR4X4A
qcrCdHWyabsEw/tXLmfqwJQ0+BBB38uI7ubLkJf2qh8SKDxMB0JGU03OuX4vD85P1lkGC28ouS1f
p6hXnH6W6tVRlyE7Zbd6oISiWrwc1gs/FOZR0ZUSuEMO+kms0pt1EirPbs8QEAvqRMeC5rq9CRQh
kgAQOnfcO9A8TXKEq/4ylSr1tFSHAb/wPqK4zpuflgD0f5xvD7KjmJXhyLSJwBI1bHjx8w2teAhx
AOOVGvF6DeDwhL71Qpp+g/UlElfqg4Rsw0RJtbQazY6nuaY4t0FzEHZDQSZshR2HEZjyl/7oF2KB
IvhB01TZ68IZk/HDjgCK3C6TQbpBVZcc99o2DQ/ssKHUSJw3p36AezEjIyl6MQxCJywVqcFLn1oO
uOFtvPHfsikuMGy/+E3Ew6T3CLJBQaRg6xq1XRywS/w1oRuQxTCI8ywmwZUdls0YPo3H+6h8psP9
1frit0MySej4FQwrFQ3L+8Vslr/BMKxggSHUf5eqiA+ikjyoj8RgShAwnZp/yBydu3EsvCx+yhdn
b5m+EOEbIAzWtUQmoojzC3+36Diq8k4+B9lftb8E0O4zD6cOUxG5d2IuwO2fQgjUAUCULn9bORa6
JTYEHNnPF8DlyqdLfHHpdMCeCIAipnR382egk/WT2z/S5uT0Dm/Ck00mVUgM/z/8fEJZ/JfkaC/6
9gL2t7ijtMVmTYdXHkN6fJoxCjhecBv5soN+5zy0htS6XlQH6TrmBXa5fFISaeBUD1JEdrYvG27b
b02+kBs47qNqLKI5Bt2HbNn+nZkic61crWP/uzeSWU/knb4tygMJuTw/YXfWUb0apYybXt7/3kqj
MIWbJShDlCTdog+AH4BKpESYEqxWA1KaIIX3YG8vc1phSOQ+40oy94SEzfoRmanuprjcrMrWg6LN
uMBlR6P1kwRJ2y0K4JpL5VKKkldEP5hm/hcxD4Ns4GYuYgxwIVxZGScY3pLuH7VC18FvmAqM/6xI
6d9PcrA2/wcekYzZzcfN3CkCcTffhukYqOropdVkKun0Op9502iH+6znpdoseqzV+RqD+l/asdBf
q6VPJsoCu4BKFdhfcsiMPHqsofVBKi8KjIwN4pU1U6VpZlsvkOMZ+zA/vIXxSaXEbp37IvCE5vJb
yeaL4Nbydl4naYMBXNUR0ix0+WuEklvGRXPKnMJ9TjU0jKuNq/Y9jAvooSOgKZQeXgd+/KaHwnNH
y46kjD2j/n4FTHxx1/PpdyKNLqZEaPcwri9G5TOGH0kEcoiREUAYI9XsJQKOOn/Aj8csTHxXPPjy
0POG2G05hUl5pL0BD+vpmYRDF1ly5gvhWtzl71ZieHDp0hTCZ4HU4GO7CNSSGbr6hfB8P34qqNS8
+GLaxLvP8TZSZSVOORAqmuQcsysHl9RaNCvCb5vDp/fkixoSQXTsmG6AKuddOp3GD4eTOlXJcNIV
gy+eA+AK0PcOw12s4vA7Fx1zqDqCOqFoma98oJpwKHtSngt4sTUEnFLU2vqKU91x5gDVQ6VkzJIf
dpAhiB2/vTh3PC6d5WKyWigwa7D6l9rTWgLmVMRYq/FGYHwR+4mR7as5oK3Thf91Iuu4hw7ADD/N
Y6svd6+cHqTzZza/RNXK3H3hjOlxW7c7wNJclbNNIa9MVURqUUewetAd2/CjurGtB1OVqF4fa+VH
xCDhQRFwKu3kiKdji1Rl3181TG+RcfcI5tG+0CQaRlH7qEacLwdh+vi4KnsBLq01bS2gm2p8/dwV
lQg1xCsiE9aTm9WWqE9DDixGGWyikvMNMxLuAQIwWqyy5En5OrLEBOE7fp0BqDhcqMgzFFgaaSrb
zxoUuguCFI0KFZZoDYsWTEbCV5LejiVqF/5AWjOGY8IuVZCdw10vVNOyr9Jr4355zZrwHSobJvZz
FvgT2iHIv4r4+GY5AvovzcJobY8lQbQ01g0ywcONn3xuXZCJ1FH+R9GWIOisZuZKJ+bJ8sUOOD3e
GbuUYeIrxkkdONK73uWT+3gyXdZDF3iy55g1NICKnmttighouxCbdTzHBDfqQ7ZqkZO3y5Ju7tEY
cQoiwNKoCBKZkCczw/Wl7LCmtuSToF4d45kaIqY9F+tYpjYo0cVGrUnqR+VBnGxv1Ntq97CJ9cve
pdT6YIi09FDeCqGJJKC4xitMBdjxu940uR/mmlYtGKIEFr3TjNOYY3NVUQRY/DruHWEz8mckQtVa
flGJHo/eC6BABmRqJ3OxaaxElblTEaXRQyjvuJt028j1JSaGyIIyDadG6rzXQMnyeNIbIOYQ80WA
eccBr9hG7zeQvkGIW7sfbVSpVUuwqCcjvdCOsakjiWjqCXJhz4CqDiv+b99EhXVPv9INZixT/FIw
GTpBv0/jpomlax+c7tsPWC04WK4sX5mrdGfokGBSJ2CTGymgqXJnZGwSa2AWKy/V62pX4hufyQL9
U+MTnxHXgegHelN0jxuyD246NIlZ53YmZT73+qb30ydYqEQPDQL00Xe7edE3RxaMLbzoBMrG2sob
Rg/XzK5gllJln6GFR4iNKBvXQ79y05XBw8JDfh49ebcuRiAkvYJsYdp+6XM5fYn5O1zjHrV9gROl
XXwg4t2ER2MFAL8mIAmxmD6ftiksopeIl9UUdxN88We4CUGgInzxXUt4mm3S70rQ7zplT6vWGOeU
aEbFu9Gladc7jxZvdgEK1pXkqlo1yM60FlIFncGT4kOUFJJtNqiIWA0V9XBzApkkfAy8lPORyjR3
qGjqfXanNwJBz4fv5STXlueFfiTIc8YJSjP+Z5dCuRn8rbiA9CP3UetSA4vnmamu/9QuC3YHTILI
J1MJ6NxHMhyVF7BNP04OHvj0UqwM/RIPDiqFjO9QwmhRHwd3QD0Dn/5FRGlYhUUYHveEqkBkRRMw
6cfL6Gz3KSnjBZIgHIIxqZkR4SWe6EkhXsukKIHKllTuvNMnPpOCiqr8qNkHUxxv4OvoWGGfg5nY
B6nz8IXJDnydqPYJ5PqiJBojXxZzmQGpacEJq5gu/+aD8fqSSST57+sh18nuvW6pFbNAzFShaIDk
oDEXgaNNkCdHg3JKZNCZ4TvonMjTwKWqF0aMmJlFGWkzv7S1q87NPBCrDOP+mJXhT3ZIQFjOEnOO
vRJTsr4/sJ3y7Umvy0wPg+cw4/5nlAhXN+0SqhHhqlsIxrs7Az0fp2tdHAd/BJmPRqfTRKryVygh
uTVtJXYg79JNLnEynZMTbAGdWacmaD0vjpsUfz9hVm2uWQ8PkSKItmAHMN/9CKh+cQGFYxcnXsKd
HVMFdnYEaCo4hqm/2s7c32pMxhE8Gx5jdxRq1LPUUQqjQPS+Ldg3Ncp9XFtYhd0MnaoJgNQz/Axr
LIv5Gzydc56LGuF8+T95lTGBfzDHrh9HGZ9GZ35vs96FYwF7r/buFIl94UxzAGAOWk46qOxJ0MuQ
vtkF9KT2JIvTFC/UDTxdvfFP/TEa7Qr6KrJyGWOepCx1VdvxzooJiIADvRNyMk6YZCaan0laIsnA
Nk1K0Jy6Fteb49caPV+3dbN433jO9DsRmsyLBTM8EH1ENeNRTbRVdyGcISNDpWLIWrj4dD9Ib7N1
c1lH6mHMFYYkurYgALHFfy9hWIRGggKnFCGvdrT0s/ei3Cda/QKo9tgCz4nUz+hPvbeY/Rb88eWy
quptUv1NMDVibXEYJpDENPYDiBlDAXRgvwh9q5Pb0iSUIdebJqrfwrHIWkVsJyMG+7BWoC83bTMh
HfkZnKSPJdHsoIt26phHRetteCcPZDx/7jlIHzTQu02rDwkDj6BeEF4xc4cx73WRSfVcMBd6Qf6V
iwCE/BaD+LfqTX87XR3TIhzNGY46Jw732avDE9A/hzL8iIeZbmKZKvO8Khte3VcnrjbV08bB/K7U
l4uRklZ3DzVt9dGvt6JvPSmNAssc+Oge8IUIe97gN+oolLDqC0gmIunEZ5CJFfKWEw6h7yq9FH23
V2NujKUJ+X7VOd3AlxLoTIN8Wrte3u/jBY1meLYDIqP0kIWUBCZvzlSGUqKjCjeTQIOmjRqRbHaq
vobRdEur1M05I8LaCO5X1es1KlmqPSwNzg5b7fT7ZJuWBeg7RrLAkUC+oJSUJVGe+uHuR3gXxtD3
M6/PoQVei0/OinqmS3E+KHWs5uBTDfhrRatLRrgh0lN8ClfD8XYuTBAb2xZZ/j+CygLK4gSPDEqW
JTSmsI63cRYO6sbfofgKeM706FBkMNvyPOmtb7BacicYtZa/6/ShBKJUZ7/gslZ1/SiDC57UbvlJ
NWzpTdC/hOBnPoypOKhUTaOHAeLmUHANX0T9OcPPLXmrj8v8wmzYDw4sp8FKbyquNXBGZa7T3E4K
yz2qmSPkSt0hcx2QuPeUR9UV3lOVxFLyOMWXctMuvu2AeamXbAF0kXuuFl60gP6hpd/coAifdaKU
GHKjk+jQ4yI15ysalnKUG8P2d52dVk8Jy8r9dkQD7xt/naQDNwKZUu6METsQXkDzkGmu74G4WGoY
AJ2r7OtntHnvUvPZtuSa8hA0P2nvsPqyWxg0QCFhOvzV+0JxPNEpJr6+DPVcYiU8ryb6lEIDK2lH
fvFVbKbntEEucFMWRzSd4mYarFPmTO49cXXFro7mUi5nELypHNxm1losSUD1g3Bhnl/ex4wxpWMI
rCuGzlXf9Eh0WNWO/wA7CLbZO9gEZyyXbvmaOW2v75XOpoCvefpW/d7wiHSG5TVYbOmVUx2PYJZF
zpBSQRFqY4Q4n3jNAVNreD3yTzUBcqdW9w3nTpnMGUrpDbnicxZt+5i5re34JA02hlVf2LQxrdLA
bIC2JBFwlcEExsXLW8Pf4acZduJJH803NKQsHLpRcstWAv5Dx3rcHRwqK4ZjMQeP/z0ZJIH6z7ow
NOVpLME9OqDz6pob9rryJVuzO5EXOcW1Nsawk+DP6y8ykJmGOsfOIMaSIZugQj9qN+KqnA799Ij9
LBwYJbuE4kHLwmngzWgPtEmIFRcTMH4+KyprjRb0D8E7LE+McT+hM2wVtu8lctnwj6RS2bnZoNwL
6Mwo3qUfopi1A0l9NMCi8sEUJdpUDZjQSJb6UqGf+/syrVf/EzAujc3WBLNnO+vlOXk0TexKAdO4
4V3eGuaTX0VTP7z1grEpK58g1rXHESwtnO90kwAcjhOWo4fVZCdtnfVmzi18DmghcnHqgGEwMnDT
448PRXZ2+Qd6KYUeRUMjQvDKe2yjn/g1iDoAG5/TEGDdqdmKUhWbo6AybkYlzyX8xi+z5udPilb2
xhb0qUfwR9pXmq2eOZiH2Gox5O59RsiIhOgtdzqPJvd4+3elKrQvvfZwdhHOnSnmS/Kt7LRPsdKh
t7k/fnt5Qsyi6Xf0mawcOUI7Gas6lT3Dz5ONp3hOOPGcCBvqMsyj6Pe0rdpz4cRZteZWsSLO8IEe
0icTKpSj4YvFDZPI27oXuNR466zlBvQLZATfLrWjIiL3xjI1uDDPJSTBgmHFRoVgBMvCcVwauGBz
R4+tE8j7EmRCPYOojti+NMFiKSeO6FA/x9sEiVM8K7xq6XBbday3TpMYjmn+xJk8OhFc6RQgftXy
zXuM7t7qnWGFVErD4dQHckCdBKT8G2jUkhw8BS6n+YcWvxK8SOqx1TsDztPZFDs7eU3Ed9s+zJ+9
s+HHEFkTSQ5At3M3DDgbybbtim8joAtX+AH2iqBt+MoPjTQ9weEJxztEoYA3BPradN2+OwQpNMdP
wS6VJdPLpzph0g6d4lKMPpx62v/LvMLpOXDa/I3ikygyMjLpyq961alKVQruz6Tkual2huMMx6hc
BQ/bGSqMwsTQlf7SB3ZJiItPlidl5El1xzKhVybC/rK5gwuIAkd7GvaBj0RvYxYtwfWDGdCCpLGj
c6RKIHp2v6z94ut8lBAxM6jtsjcK2+4ReMkRcPyT5ubmPXQEu10InGX1Oa5Z6j0N+c5Whi6rOSbH
llYdnq6GG3354w7dIe19U4TsP0af69xs6hhdPtmgIxcKYj9n9OLO6M+QK54eUhPWiFVesWU/q5qi
jIN/naWK7o5qlVE1SLJxxfUpMge/PFQuSDWgDDbfRojdSIda54N12DOxCXCV6d9I+pyqw1B6ONFa
WMrFeO1Nx22h6GArMwWz7aX+PJQPcFEoG15Vvh/wgh39YYwS43Ttqd3XU++y6jqD9NO/7WwiCPp9
HdKqFz+qjmO2W6BWL9s3BlktqzljG5w9b0ekELa5Bwa/E2ul4AyH5MthiOAg7PIfjCDjE8YYl77k
wYTtghAtBWYGpI58iETx2W6v/cV93KffCIEeRcLWSOqHTXmBzESDCkGeChqDBevCXYBbY7lCMLk4
K4Sr1hZP6bYgNA5JdismtafCluC/yfur37o+VdAwgiRAQyFX2xAgpekwU9Uujc5b/z1M+gTDs42f
OwcRTHMv4UGRAg5WSsTbbPmDLcBLNpT3NnYBFaWBit8978XvR7KBPgGJLePkW8ba6bxvq5SnBKVK
3X3bZlYWVEl4Du3KdhsKwx9cuXFz1936+HTrk1yr63DpJZoAyE46pkuzpXhmPO/ImVZnfImveSBo
PoVfG8vsgKYmBwL0N4pQgwoK7t43bT/bTjC1NWugcE/SbAgyOVGqlb5Xesc7rdbXwie2vTc91aUk
ij6zZqkZXYyT552qLum5Z0vnUur705KA2yXwUIjYK4OV+MrXPZj3Xc9YH6h7idx6y7tmFp3vKQ3I
B+q0b86VoQaL2i909lvYqwgwf6B5CI6vss/BFPNKirknsYtzLyOYinQ3OTRXtFAZnaCFg7h80KC2
3oNjtEJ0QSJ6+d0mo4xwPD60A1Wh33yUo91W0pa0lR0Vap41djm9EOjEv9H21ckrHUJjs5f2m2Sv
5lXOPTb1nr/aqioxhXprToCd0k8MoCeSZ5jdfBArRnoy5sNTsikRsjRQUoc2QO4xOgTATCds9oqc
h4jj0dOeEpbvvCZg4SG47AOQlr8RkRe1Jvsdf8fCA2Ts9cPcLbEY4p+q9vamLGg16bdK/mt/G4F+
lBQ1ugRnNsdndL/Z/hut5SZCz4KPcRNnT2yO4a5TXauqEuekuNq+tOpdCfsGrGhDi+RUAFvTDcvn
dhIm4a3F8G3mVbvTL6+xL4S2FmyIfCk1VTnAtPF1sGivpdS0RsA+e/bRuM/xzV8M/1OHHNO8EfVy
ez5YpbBh0sGfUE/lpoOx3E2geKpFDXptQklnsc5nvfB2yOFGs99u+X2zA5Qp1qODrlsH9HiLZX3o
zF3LkdcQkjONyH+rSfDqlliozYy6scpozi/CQkTIVhT7hqtxI6Vd3WDoKX2Vj4RId2U4XCYPEaxm
N2IQWwcOChJHi6XOsJga4iOAAcxXOkwp0nPq+hdLaDVShZuzf2U1wg9zgQUuDjOUZHuKoTkVYPDE
srpFBb7OmjlxDxp8BDZtvjhJXQTmsZ9RAd80e2A5pSiL7DINc5aA10gzglc1QeUaeK8jaWdRiqv3
4geFMG0P4Z9LJxKUQfEYbTwUdXK8O5K7nsvG09zcuIBXnCWN66OQyPbvdij6//iel/QyQQPMxJMr
GwpYPrKeSJdzN0SHhPpDeL7BbdLjv1EaunXtHMTeeX3fdeb1/cnRWeNJWjstMPU8Bzz7zcZrPCVC
oDLQtasOS/O4AZ6lUdcxdSrA5Q88f2dCremUsjEpNyFnvlgjedapLZYFUluswosyfcDVpiHsQgK3
LJBGrvCpXWUrD0wEiTSat1RSQIMVANiOSaG1rnxXqD5kI7hhPv/Xlg3Pw9/7MyY+DPebI1QwkOPN
vRXwU1FbJM0BOxS2K7Plhzk4+FwInnNyn5IMp259B9hyvUkHLTF3lqK6yZqcoY8SDNlMevMQCGLz
Owuk0BOkoSzoDoqsynbqZw2x1U+QPEDpa0c3qe51mLqja9GmQ0aKYIW54/xE4fBmaOV8y+RLEXXo
F0n3dPEsybG6A94IeCgxuLIYvKVkFKVJHNwTMHJFQi6Ar/Ia7wvP4pIAcSo9Z9s5ROD15oIZnI5H
f5r0oXwYYgV9GXc1XM55a2ElQikI3t73zd8CqUe/0bbSkvx2Pzo8otYk3gxlyV213pda0uCNBgM1
1ALKM3KsIBD6Xr3ve7NknQ9bf2S6bQMpopYVjGVDPY4n8MGE0ew+NfjtoK9mZLOMEBVonW+rlhiC
cAXjKVieOdiqJD+t6DHImKZQ3TLN2mt1qRW5wbpVRPCSShPqD02RIddnHFoh9teZRFpWw1x+Jbco
6HabWz1X3LNt/IuEjoD9P1ngi7C22pmd//JRQIxUyrkwmrKX0HuES9BswwP8eS54kusWVsJV9HXr
5w4Yn5MdC8jVztPdooC3FqCKlIRCQZQXZi7XhsNctJtnKhoM3lWLpkj3jhEsTM9Stfuuu7+4trVm
wKDLh0R7+SGPo7QHPKKfr3wYU9xnMCgBxWH7EIAaU3s9nT5Qls2qUdr8L+I4wItxtRaJK7E1FZMp
C1HHWco8pAr6TOVBG+n/GFFH5ALWOLsA5Nr1xA4G6i8RwSUl1RGut7LzkilE4i/1tlPiiETOjzoe
jcz5G6b97wEZU9yaAslslDbTksNxnDApDLjUfUfdUQ4rDMVY9P5NSouTBDNfevTrCCOVUiaOYKTE
0KyZ2Y6KnpjDEX09foz9NqBmvAehIFJ9f1hXErEGkRLcddwPFdrMRUYzbzdAj5a8vNqQjPUxCPti
BpPM0PWB/iq6nlQdUc6Uans4Xios9fhoYRNwm/0WoYrEuv3RZhoQ62RlrXssw+g8pFEDW6jCIZG+
HmTpsoyRx/fixjpyAOBsjEPjfJUTWzYJotbqOZSZT230cKjsvprLFnHAPOTYPlY/+zDJYY93j6HR
FX7NoJFocE5z4cfxEfQmhZDr3Kl3w9XeJi9esP4H5wE9QlOjs6Myn8HXuxulddlYkqlGo/UXPZmm
1IwvdjaOuGks1oy9ZlP09oLDXvC7vG8Ugv9RshFHWsKbhLQsJlvbwvy0j2FNFnBtmhZT3UMfdA5D
X4UAl+BEe3Z7aERX2Mh5gD7OmbxJ3vphSSMVywaguMAykcuT1X1103xmsLHff6QLXkBrlMt/ig3z
rjIUv8QVJu+NX4RUB4STVcvt/5qT2XgkC2hJAmh/Fdl0Cd6NK0I1oeY0ceu6L4K5AgsmCu320S5i
ztU7gFIgRfXkhAHH3zBehyK7wC9hsfwZwjYrfkLQ93jiD13/yGM/e786AtNjbiV8SPpsckhWK2wh
CFSZ5ude2T19xNi7Dln/bPJiTuFLN3hdbfBmXduTNsTeaS4nH0DEjcobSak+hVcVxgYobse3Bceq
is8UXh/v3oeSqyHbnpse8AFxSkibcvth5Onsqe2dyXmDuyQxGp2w3T6HdB0UJUgORz+PwPUpYBdv
fLeO25DNoE8jBLDoLLAe8a886//ykcfMXsNb84+Jh7TP0YRrjW7BpZnTkvzKioSA9R1yF0up4fTK
kGV0xzIT8hj/uhupwKX8cQ0VHJgKTJpKcecn3IztSqzHW9Kwp5R/rWjKcYI/bTmtkSkw5LleAEkE
/DxX4MzDDtVWmFBzJN85fyC/Ek76nb4Czvu5PNh/i9AJBjQB8uFvDKHiQ1KitDaWycRkBd9V3RHV
UiMYPvVye+L8mRcZtdB6Kn7HhTCJWsPkpcYhZVPVwWoAL9R2GVgHdXDhVsN6/FAbg4YIl/d0vKRt
BxsIDBph2+UJ4lMy+F7ceUbcY2N9A/+ftaw2bCzlUnEjEti99gLPliIaCYr0h//e6lVPykMiiqZ9
Q6pNqqQ4lVX0RQDpqB98aH0A0nHlxRDJq74Pdgdcj+22RluFHIclRZg3zbNJ2fcU5tD6X1jqqCua
rHiu3uYsO3DM4lQhnOLbbYTRe4GuXcf3P1Fvp9Gr0QVtwXHoncWlxTRvFcWYzpkeBdlcrE1qLshs
KbcLA/U/oTbof0vK1uc+9u32EA6Dp31E0/ZYimtbYltiTV32nCWZytOt+g6fVJEHuMmFItcsEpS/
OG1vCsPpLIyvyMoAnc6wL+snXYtaisTaLsMEOHtYFEPMQZHTioSH8v1Xbkv0WM0I9tpaVAfFfzCg
QTdGkbfrnS1x4ZpXtQjMP3zSx3QODTzVEZXnjBpDwMwM5V6hIRMa5NbO+Rjn7pionO3QXCAaNyNl
7BnTxuEd7G5IiDQnN7hyFNPxdLMUoY3rS59YJ9TnOpO8eA9k5+RBehT5k6Ma0QfS8IgG4vbDSp3V
egWBEckUywpuXmd5RjwZP6cRss/C111TWQbqgDpasJbTSQO/H3h6V7h9InPHsatdBxcMxiH8L6/R
hDKiV7bZltMUtSibvbCCV+5fzXxjyzO8jY0gAP6ajIxmlYnAynchzjx0kYrgagHthscuinIQGTss
Wm1GyF33mSQ+7SFC2aGvaaliAzjAlN0Z3SQtp7vGOF8C+RluOJ7CLpX6J78BtfN6kIcn57VfaqhF
BG6tfKF5vikDacTkDWceZowws1hCynZF4gyVfqQvYfoNishJucxCow2GFJyUaKcn6CoHFy0AAkI1
W+aXc5ZYuRqI7OTVpUkT8DFum6wPxr99Qjof7+OqYaqHjDP6UFKCBqtZSmyjeDXZGs/83QmKWtQb
ejg8WK7v28oTANgFkB+8sjkkb0pEsofaCkpnQCk6bPSmUvhGsHZOy2L/LoQpun0Uout8fAnvEwUC
Gp6Zk8WIqhkKdTAN/8anCu3i8DptMHE6BOQuUJE6xLcRDXYViCSFNCMt4AxOBqz4IdoYQFCgoHq9
W4HN1edQFl4zGt4AYYKgkVVLXdjmbDCUqBOxftph1stSBMxesO1h1Afe4j6So53cVarPdLo7MlqA
Pw9A+ed6Kpwz/5uUbH3aRGJiguNKphER2ir3OeGoD+TkTQbmgYBaMEuqn7qBe3Tgh6kbG7NkWr/u
gToN1Xk+Y1kjxTHMJ40mNabMV2cTMl3HbtQ0OIiyQZp0f3dRjSoitCw1BkXyYfLxW7sUHlT6Bqpy
2aURfI4+QHRofkeIZ2PEQgBu5sje8xgxPnfCerVgbrs6VUbRA7o2CDdKQ+QqrXoLvOkkXA5FcUAc
ZOK0u9iqXes8sn3YMytYn2LQFlivEwYiXr7ulXNC2lDKSrQTOIwrW6xkPk4kNwaclbnA/PGdRWb9
nUef2kU6bRNDIG+negL92gLNFOIGVoJ/h4BtrB+kRp+4sPVeaJaAsuSm7SVfMAFS66qVTlcBcwHb
WD4jYzjbaAHMUAhy6174ZaQEiv0KBDksKQls+5kKemJxF6tIx2a2TZDpbBJY/v4Gfq3oWNAmVUDB
S3V9az1MJLezgakp50X5sB/X8lwmXZmDpANJDXoyN8ej2UhZhah4jS/lq0gZwvZ7EOpCGU6AMvd6
hLOA9GC6/jG/cujdGUdD2NGomPuscT5yPSbolHMtdD6y4yCW1GXX1VN2+RZKNZCrLN+JQMKgek6X
9hfBMksIFhpuNMu3KVcpoDYF1pBgLnq2nv8agHscjzclmxbr0I5dHumY3dddev7kZBlmB03MCjlX
BB9PW4UknitLenPlDdq3cGvJJxXnIltfkO1rUKbTwp7p9Gu1DFFRpZB4jnL4XhTj3d3mX6Z4Y59m
aZQ2CJtAsMsS+Emg0iRKK/THcmRvi1SBTf24JDhX+dhX7/NpVKkMHwUkkS2FgvlKiH7p77zVyxor
UYMvVYkPKlGOu2zyfYLHMWHf/g38tFWYhmoa84raqkSE5nmwdN0CP3pxjkM+89TPQwA+lZhlH7mJ
OhN6UItqoSnm/D57lma6CQ3uafPRbfVJzHsnx/vsWFATFGyCHmJYV8p9CEX0LkwzOe11nk1Ymsl6
PoIiqSdiSz1AQP35HJjLxvfaYDJIMtFuaFQ3tEj76YnFLkqGb9oemJG5aNa2ljWP4Xr2o+xUNibO
R2jrCyKHCSJSCjLOik3GaRUY/lIWaAalxcvUsrMlgLmvby48kragKZz2rJV3T+KOQp0MdrXaNfY5
SP7FJo/zNnXsPUEZIueMVY12p7YkAUpNpINtgU/veXqaUKhuvII09PLBG3bly4JzMsgbCogPT4ip
E4ad5qD6MXA/UXVp0wP3L/Dx56Pd8+P6XT+mXbMIusmx2PZquJH05pWGL60Ji885w9AiU9EmknMy
1dQUNUSV44IJnUSELxzMQ5GHpNbqwvNh6Z2wWXZxaqJ2rJHkHJp+qsmFdkOO42Pkkf4jDARaJhZi
RYbpSOfWF0BeLuvja+LB3Eh9fO1wxEmNsrGaXSxHIBXV37k7EOWs9le4uKiNT8Cy59i09vqQh7Cz
fAya1tHsMA/Mth1rRbgRYVcmkCuRBp9bQkkd2tMChPYOCI8wgN+di5NoQvVTLnj0ABcXPo2JYhvT
pTuFEXdybuwUisXAuRXwYVLA0f5I5xWZmyp7TyzGPEOIaKHasMbzoDAcPFrWBkEQHlY5FhwnyK+S
ha1YygMdHODoIJWDViiIglKPJSJiwFjP77Zpv8E5PPjJQ7btrqgHu1m6k1IF7AN2V3Nt4IiihPb4
38YbNcvxwarxEAn+oAehijxayYgTb9xsz0tzDy2qPqQCZPSF1kE+qF8elHQN3DspV38IwDfPkuy9
wemS4Vr3u93qrF+Qphem/yMWrIM9kGKQjnGYACLuAvsI7b0FT1/CR35lCarJZI6ZqC7ZPqBsotNV
m14MlxpAXPOnDy3fNtDS04BJafdmpoRV0Z+Om+lY9yEp5UtKOHyKu/fWtSNDHSPAjyRSLBQtVOci
8CCsUF/xpNFLAnaC0hFzkhe4bIqQC8/rouE8XyjLBPfzTIW5OfFz/ZAqchvcuplPkJWu4s+MjuaQ
z+bYZ/LbOCoZ336cVfPZy7xOJ9sqv6ffFdm9XQ8l/ztAXcMZ7kRvVDUTHRJ0gGer4D1yEHP6NGah
JSykLbJ4v4ubw0cd9Hawv9bIHd9E8PL7Yo6waUGiSL4GTrL4cBXUd1/JMx4C6JfbgnhygfoP86F1
mKMczCHYzFTg+t8a1MsQp8+1lQlXSQJDfix8PwNky5aJKMy1LfCvvwK3gVcsfP/aCiCFpgthBJWD
Us5j0W79HDqO/tfAgHpVOt6C9DMUx1X2+3eQ37FBeFpjK+AeHzNQ0kurYlOgBWGFm+m7IDgZRnmA
O2ZbIJ8ZJQa6wf/xsYaufnp2ujndzv0adzfaNNLxnIUggKWTZ6u1/gCC/5AThgT3sZPzK42woS2G
CbSbKa1FgLAnITXsShIcAcwLBRg9NXx5/iHoosjfqRF8xMn4rPr91F28Xvsma5f8cj1U0lo8eAQ+
n/09EvoPf/dAoP51oXJBQssMfSwZbE3DR3mhRHpBt1mqbpQRBJncQSwvvmAJ2Fkr2VssxO7GVDwg
upEi3PNta73UXaji+UoMNpo+eszL1FM3eNnuDCJ5NoXUN2trgMRAXjscddiGubj8NBGpmFnZ6GsK
K6T1Nr3ciCA5rp4bekDy1PU9EcI6vrqli71hdPb3WTJRmdzf/MxWWwNwUBwrihPXt1R74XnHuqPI
a++tVge/WGU6MSYJzbbnYpJUuX8s8cSf6Z7lr2CVhwouUyc6QEsTofIjcYJ9l2Bpn7HsEeFB/KS4
QszFdA3PnSmYqzg8tvnKF2r0qr08sv4xi6h3Usx74s9itZT/Ks4kwUznuIIkJPsIlBn6cxiM5/gc
brEgZFubBCvcC5ZGUIKIo92y9Spgi2PrQYvL3LTwCrerNl2wIBYnxa1YHGtd8hEbELoRbehKiO6m
/wbI04MOVN5TPDrPT5/y2REgJCB61GYTTf3cRxU16RDtjXnFE/AgbXeWoF2pYzEA3m0aoOITS2t6
31AWVTK05VxqcdLDwzTMHiPjj1Vn21rVngHOXinXkO4Ad6KNiwVmm3jLd5eU5SBXLITmC71Hf6uV
Z+3ipCtjD5p7VwPzkErU0LUZuaJxzRCFXQDW0hrTcgV2OveQpzts7jIabaa/+vqjdq4/0ahpg2TP
WzGCGUEjcHDvV1a5l+4sS2cU8DQpWyp5jHNF8xkDX0ek+jii+PoXlp8ImqONqc2CjnXDlbJSRWeI
G1iVR2dm3zLlAK+6J54YrOjDsJffsnMy5DIeFoPGj/G+JgV1tN6HFgxLUYBrYv/o93FexTdjLm+c
HU1/tV7CkuDmA+j+bcBY67uxeXpvO4vllsD1NC9JFuHls2lJ6GqPePy34KjpA/SjSZZatUs+DPlD
0iYU8TvazUN7wXD3iGiioBoyB7LJEZv4aQroh/2unqU5i9WmgG+UPjxthj9ti7y2AP67+IETaTc5
eUCxIFfSMsYqnbrdoyu+lWE+4QOVXZ5VJWOmG7Op5JJ8/QPtstcV6wBxWndWprNUtVnYd2FRVlrY
EiPtvLi8pt84lUehVERD1gbEZX2bZDlJTY5uioHCNVjXZthQpcwCFBBX5z+ZnyazPtfOH4F9fMiO
U9+l8UfdeHwMV4XRa5x9GJdWbBCr0MKRaE/6uZuSdHtLe+mC5dua2Euz7s8hQvrjSd4Cn8dOD1HR
Q5llPEN7kcQW7IKdx7kUYfYDef0KG7aBVS9bj91Qepf96Hr/aSQ2VmJguqL2VqzrXHQcT82rlGiZ
Op1vR8rmGEBt4wcj9r5R4hksCqJg4RvZX92bkIi/KsCXeaxdKkJoYLt5RPBBh3AqVUP5ik8qkNNd
Rp6T7ddEUDEHueA+8ENLLFtXpH01nSAuCGOTgqKTtHOc79iVmQ7G9gG+6ttCakgiqMjIARaEWDeT
vHCE4KognLuqGkO1s1cS025VsA0A2CRSAKqGoW1jtRuIgdKzB50olu6f9PBCus4x5aYJkl/4Rx96
MdEva+8q0vHf5ssBwyNwbGIfSE6ymfXPikycn+SuzOBchIuu/X5LyYTeO971gRJ0ScOkBvQNLEyu
dg658RIocY/M2yvTeJNvWsQkFD/ELoVM81EECZ3Nq5BCL6oea56iVo4Y+SZfay5djMXEuDZB8mdL
u9FB1KGAaq/g94Diz+PhbgFg4LgzXglk4nX/+axmtdIiyQTWypbfUuaoLjNMsMwskio6cC0OK4kT
SIEXc5yP0e6pDUXsVd+jTMuZNcv4G4b9UDNffyPI3UlFl7/oi6SPHsaVUX90DQt25tF4r4tWHzgS
iEoUgEWNqf8bCP5MogN7NxwPWSu1WAyXc4Ra3yzJkJP4neFW4lvGXsQPk1ad9tVZXRlXKN7tr/Fw
47SBbvWggodMa4u32ho4xH2gG9g+2SP1qcqDNOFTA3I0rav1zXVLCkUW9UhLUlSg06l3NcXiHdhk
f7krAaE58iarogeudjPkYqICWs8/vdhE59mv8XEVmUS4y9/YnUP3foCO//KIZA0hU0kF8m+5QFOq
16IbS46uEzl9Ihj+S5vXkPW+SavDiP7/XoARFk5WAhiUramw6BEobrBj8yM8RnNMMYo1Ca53wHur
pWJU9Bg4Pvpraswo06WX/6n1WUsaspnaus2pXJfVF+KSrSCDJ35zVtnWtnXQgbIlM/VV4I9d7jSB
+e9acu7LbtJMl9cxCnPH+EQehQzuKcm7KIZ3EDXWdCLUe3IjPzv+M1/ultBRyj35lPvcwOX3Jt8T
XZVp9xy+oOOQ+f7DaBppyZh/YWYq0itUEUYsGneeC/J7p/d0c8s3Cp4AvgGBMGUMBWGpy8PT3TfD
Af1VET3TLJ0x32pPxP3VplqJUOuAv9d+6MT7ayP+CXBnBeDXBIqV1+kHO5Vahs2EgpYCZstL/BxZ
KGw7FQd3+Kg60s8DdQXniS6JQOJXKI0LfLvrRtjHdbR/h5yXLVyLU28e0/5cOobDRTVJ1thPDCWH
eMUqRMaosbJXuksFrCrZWE6GHRw/T/JbaO4Jd6RfslN4tlAF4PyiqgB/rlNlDFa7igS/Ghs9nZPz
DJ/u7DLdrkBtGpz6Xpbo/S/efCgyhZrxOd6En3DT5Jpw2ST5U0yOVe4sfhnFCHbyPcpG7BsjifE6
0phKeupp2hBttNGLrze0QKMBJJuFPWdKjBZR8VaUF+ZA4psVbx89N86BQ5zBl9p8W95SRgtLGrW6
/0BU2G4Qg/r5UIMoud3SRBgKe6dXXJIi1XoOGDBMI1XFffvMIbxY/7fb9aZmD9AHKdNbLdM0ya72
pccuAKhXSmGFCbNL2nEGDzvDxiL9coGRFzdinldadsgso4TsJjZl8h05xaNb1d1Rk2uWm/T0SKz1
BmzrTlALmxMoUkaE6Rjf7Bs7hvyDLvT0LVdA6QoMMjWTTkDyOaZcUixxlIQ6KBhKt6cWdRf3c2tt
SgD5HAbqlElWJA3LoYoJMBfUf+9p22PAADpLlvLN4ppFd75VpkTilg0tN+33FxIREBByquW+v/Pe
w8gdCm3QR2qXw+1+PzFst4IT17U7c2FsUv4/0dxhB6NXALRhVroyrcCGplRt8d+rhADQ8/Yym4Do
OnJLbVsfH+0etblKRYxumJlSPKRjR7RTlsxtVXgfHi39FshIHO1/qpw+oT76ZyCps6F8Z15k7j+e
wIGjN9RPiOG1HSKyXOfQo4mXt4GmJ4z0hrMUUY+lLHdcK+O3DhqNI96dPOIqam6xKpdi5Ks36gRH
VPuRqrElo40Jam8H8suStqELxZQxjx/xOUXMB/C9Qatei3F8bZt/PiUY9V+bDIcEDbKbdGMN661W
DJ2Gve071iXsG0xaGiHoSQSPmseHL9CxNRe32c9tvgTF6y/cRxqY7wM833Sa4V8j57tmVK5Kj6K7
sJzfudApQi+LgpWRfziH6C0/CqU9njkkcwvX5EVRf1gY6dVs1bidYe07u2455C5HJbZx4RnW9laQ
m4Bv03ofwzAiFWPeqUttbkJraFu3aMe+DIwi54OGxYIzn96h7DDPZhLJOM1k2g6TQWNJmkTvQo2g
jJGKoPsASE20lr9Qa298pvFIISb8coJC8C9F2RvgeJvIuJdscag7XY4Gdg9FA4jYEHUgrc5+4DxD
i5FmkmlklIkBZhy2A7HXifdv+vheNECAmr0MI0p3mcZAEFpR86Oe1hGZnMBgWUQrhN7vcVnblH7b
8o66mi1Zaz/qWDK3neAkq5sV4y7O5E/g18mR4fVpDItKtSB36ejOGQqVpnBBmIB/+Oi7Tg1aN5sQ
O9mRSTh+2NRIyYrKhvhKCMo9EqWkU1dQUh2jZ+zXycYhkmSCwjt3gpKc/7HHC15UwFLluqbyShI6
a6HPIkwkh8gNipeRMP49cmZZQe8VdGxGMU4oJWkW0iG4GPRaDoUalG9sZhamLIrEbKETMTojliHd
M4mq1p+L9fifCImbw2D+IuTFg39ZmcnCwmuBfsC3SHjsDpcnm8FjYb0YkGj3uJbT3/VZRW13P81M
2bVN+Rw5RwuoUknPu63Tph5PuI+wVFDNLJbJGqnqJ/Y4iHWImtg3JyVundKBx8XbbEWGaVcH/4d7
cDlKcoskbAsSjhSEx/RP6F3tEL7fay8lDrfnjziKrWcmkLiSdrdNlfxqdAM+HKCk3kEbfPdijr7u
vMJtLWLIn/E7euipBdzKK/9Gicdf3PEwRg1xOoswAaPZgyfL+1Bqn7c1mNvhRI9j+8Yucf74HbWf
n8KM9h614OglATTE1dkXKsqyo0Yeuf7b/T00+Hzrxz7tEPrMMYMU8vOswLvtBfSriR2hLQfZUM6N
O8r2+Y9NTWng9CqtJw/m7oSy+bDWvW0i5cK7jRGnIVhL79VRyIxq75vO8vAiL/JhuWae+arJVTeP
GjYTbTrfg/NOoZ/RGKZau1uO28N4IC7srYXm++cHL+UODvJyAz9vamyPoqUi9/Sn/3qa16qm0YBA
btrLDDLKn3bV0mvoc1UH2bkuKTcovbhBXlUAHuENu2oBwplMFUFwYECQs4PRQhCKxXX48KYbQKOG
2caE7gp51m20XF8w4jw3BWF06v6fmJpl/2wxZw/6UtCv3mf3yOviSGFYwIZKjbyFHg70S1diLDlr
PwBXfHTk+MSN16jCkaUEXa9raOcwBew6yPSErKJaEKccQ/rK1Pi3/kUYqnbtTFF6wtA5ZW1hbWd4
+bpnmCmg3bm2lT3SgLy+JYv1RtrulvunMXnG/g3Fe0WVrdBrLPhnCmO8rwaxPOcfen/SCaH+OfI0
jQ4/E8foeHwuppZgGunCr3A6AAjtX/1Fjm3cpk222CnC0svJCTbarMn2R33J1fmVzFtg7pHMdYsG
AMAeZ8g/Gkat16eWDGkxN49v0RLjHxgF8PfZQIJbnhwlSLpKzr61soP0CLdqO56niLxjQoQfZQye
8oVaB5nf/LlxzkcKQXQEkvLCUQBDGfnvLcg3OpjdazmR050tdVaTMa6+g1R1Vx4/EvrPDHGrDgpC
R7n+9NItHJQrf8BrXpJRYLLVfAQKCwN37SxLRG3LyeYLkT6r2SxF9+RWA2ic6pWWfthNE8dk801W
TDKr10u/JdGuY2wCJ3hR++E/XTDSOdZqAI+lOk3IuF476G2jT4/oiigtz5pDKA0EVGwvZ364rOz2
pIhOrYrr+TNb0w3HhKaHkzlprMpdWG2SVqhW/4GPqRN8uSEzY8aFZ++YhHN+Rd80HKWeKiDAkphy
vQvimyJqjPnhY9EVNlu+rwBjwp2r2VMB5NUKCNX3l5BzUMEG++fqSjwDfJKgdTmPPV7fdMUm1HqR
/9rRK/O+s847yTOKozcKsVE65AlkIVBA+hdmwH5D3VJxoof5AR+UwgjG4LhrGPiVzBK5yEIzKmdC
meb477kFBoCrmNljnQTAAYuaXDi4/iixWV2ckYD3Qxmdwrz+8kR+EV6lE0P7nXD/ymr6wW6N6jRV
qdkamw2xpwi6TwtQkn9uYNQqLIhVBpCWEI17jwnaa7zQ0SsKEuyaCckxzGjxJgM6jnWpXNIFmvXu
El+CP25jJaX/dNa3bddFPA2/vmAZwQP7TYecHeK+mi9LcwO6VvvuvE9HLBaFJLKT5Tiqro5jMx0d
SllosiLw2/pYrKjzUFWt1jDfQIalqLCGwY8kbMy76sY1LfQLImOilGBM0Bw/kl6tgwqOAkNSd2Nj
hBio1lNfXeOP++ATrTryOpklNW1yqFjx3EI1U2VO04ULb8WTDIzz6NFu7RSALv24jx3b0S6l6eLw
008aYwrIyluXjtkxCGQIjfCCtzSzjv8j/8WRa5RPrpjdYprPt1+mllMPgAPKXYaflp5MpO8raKsD
V3/UR5x2xConYx7FAIlCUvAEmar6MHn1cCKbUXy6R9WhTBjYdtwSsgCfCJBjSlhvkgw1wdnihlmr
zr/1GbozViAh65z+pc++I6M48JPJxx0q+FpJlBcLsvw20ZjnJe0G+hy98ETxIPs0Yc2PeqeZiJss
C3/HQNWmOe5HYWWae2R0GxnZQkw0vIebrFOfbuLy3bvr51jNBTYzhsd7gfC2X7i768QSduDV3idI
U7vNkMzd59BBvbejh4FsnNiWkd0lUFijOsZWvxdtLg36ggd2VCBAy4RjVYz5qSSK0gOLCCfTjyUw
XgsfadnwngZGLbEiC+E1mlmx7wMZQo6uU4oy9IGKA7ftK1CmL8IlE+zp3yRFymfyTJbrk59U6IvU
1jLsGhwmkEGZU0ScsRYD2KTcr4VKUZ8z0SqaGjda1u+D/JK7yumc13XSGfDvTLsSWu6B0v+TAmLM
t4SAJnnS2LNzyYCzHZr+a8SYvtAgNgGrSo5pTL1KHjY08rrW/Gs2TWBrQ2/KFKG4qCJtlgHyzUXI
wgQj46I0EafVb4zvj/yTRM8i+H51mqlaB2CD98ExZYcGwrSKIXHiBSZdm515tdFGNY4JFEROa86O
8P/oQvyP0NuA+iA/PumuJSp4y1HuHlOQsUg5DKIZYQDtFLJidJc593paPytu1GB3zPC13RqdQYn3
lg9S1QSfHftQCzikEe5YWl6cKLbFMH+StcL1zRRqVEVRExfgb/VxuQ8v9rdFa9PpQzIsbHux8tEy
Wyskwmi0FHGu2sTVt6N6mhvXsj0UDhq7QNnSL1wOv7kHn2qhcZrGrWMb3T1HDBoUoVG1IVFHItBO
R5cAs7VdKhK8cmUjQikcuz81g2doRgrcim9JfFQMGI1e9lQJ/z3YffOy1ssAqDZ7lC6qzz2lzzuF
i1jYb1ecOg7i7I5MyBqaB4cgZeK9uFtN0J6W/MCiPwsMvWNoxaV11cKxkNucREcEIekZjsTfxpJ9
QxmE4Dm1hp9z/m4jdGgGR72uXa3gdUgNXYyNc7ISCXKjdQUUTy2jQIx4arwRHxdzd3hRgOqyL1av
I+MNj+SuCSzvObcWCJ4odooC11qgG0/SYQjju2h/6YdxSY6Q5B/P79NHApAibZWj/hhmR5cVzaO5
ckFC35WKPpj3PofBN0z/FukpiQULODk/x2GcE/gvWXllo+ES8dganidgnJqGWvkaeHI1neWaT6d4
fdbCqRajNxvV+pN+LEpqDX29tR5O4xea6QJmO9xWgrGvW3uCEDO2Jt8cogQw4a5PDb0kJ61rxWRb
5wfsawoNV+xn2WiPfEb2lg6YSgMYe2wtJ2sMiJCKd9EhpW1vXzSkSWWohnQc2TmJEIBvXRE44TJk
3WL74XMYikC3k/+JYN+a6Aco5SnMQWkwQQlK8PMTlykb26RUH3CKxuJRY2mVbocAsMhLujTm0/4e
l1gtx3Zw81Xuwg9g1yKg+T3oOOHQ5x/32++DQkfjsNDW97GGuyDHKsHyAs0L9TIQ9nyzynnQpgHh
nSeQVgqNK8l68iKO/w1e2hHYPCWndFDikurqrSQ35KowMRbxQAEG8MgkkubbXWGkM3hoZAZEs0o4
K1W+U9bj7l58ZjWybJcg1OrLrZbOB88TfHaFq6+OkoF8IlG8oHguvdYguBQVGOt2hWWwdddZPl6X
QzLvfSxAlpF6EoljeCMIgNBGiIq90RjoDZYjCn/YcgYAifNKMk6+YvI0K4nK8BI+idDtdnksKMfm
SSYQmSNZFbnSrixlBF2HcQ76c+S4SNOP1iDVKWSqQabEqOr3XfJQobgGcEG3azNO32ZdVh8y0NrQ
DdWUKSNV0H5CgrEFKte/dos15XkfKPIgVyJf10DRRRbYs8YzjICyliAmLiXV9dHKJbjVxtKX9/1R
OZUsGZ0AWR/jHq9INxG3Txom8deIX1loEmBiqVz7OyoVNTU4hVxcT5pmONFpJvAvgoXDMVINmWs3
noC/AJ/2R4lWlF1l9ZNAuCj+O+tZo4dGBIFW5OXYVDLZxkq7m7verGtKejuCyxBqFwn5iTYuz6NW
8rL6+qPvS355hZVQ5JnKtPvMku16WOrz/HiEQquMrAoqN7+2xbYqScE1WInuedit+JfN7voVxQ+M
7VSFz0CnfocrIyG92oMkGqebczVEsrhjfG0AXHiAxvdzvmwmLDqvaAibS8gUVxvgLKK/73Rjf1pJ
G45wepUsRRb51xWyjUvCvUdSOGqvpsYx14nZfPLlOzuL4+EjAGh0+yFwu1OevP18pVqe7IET4hEM
sc5/BEz2yEibAJQsLVfCB29DMUke4VC9KVABp2GXefquxHqp+OUYLEpH6v92P/L/aHWJB8PqPz/8
t/jtRvelOi5yOdkeVWrXDpCu1FJgpgiQ48jIsgpzmLva9fIw6RPaQs2C9M5Zpf1hx3UVDAwng9oh
C9U5zSuTubu83Azb1zyFwbzGgTBZaqkf3PVd60WxrD0jyFOs0xkMzccu1XiR0yhYVC6lA/3WRAV2
qQdMyLKXnjHMh4d8IHCGoKz0cQO7qj7HbfvKNNqrp2GVW0cIYXNQNUCWpBn6z0+tRrzsdqWJ1Yow
cu0VkFTuT4Gsi/r5NhmgJoVATLJuyQvM1M2fb6u15aptA/5n04xDSLuNK38Q70pSoFLNJ+hhyIma
cwS/o4CuKjdzBFpFdwwS4AVVHht1OXUXgTV5D53LiPKgZJwbrci/PNjkaaOJwzTCD6dUTjCfUXYM
vFfG6D9iz7JqCz/rL1WGuAJa+V+SB0D3Cm2r6lTv0k7OoZEqMpBoEYIJk+DBQBfYMiTQVXzFMF/I
A31isDZrSGccncyU3InWvQkPCtYHJWcFN2kU/vV3jYOYqpV9YjPLdSVz4sZy2U4t8iBAZOa8xNRh
e+1nVv+/lzXCW7qBM3B+owUGkEnp9ojfAh2ZDIgQm1Csl61gQqQPyg9L1F8LsHwLpZlPtVwAPwzi
eY20b/Wb1US4IlJiutCNVU+JmDYE23Q+G5o8c/LlexyBJUi1zuea6jpYXh4Eo/2jKb+30lU87LZU
5TJtsS2ql28e0KYc71lodC4nxnq2qWv0QDJ/pwbQmwwNrG1BaAP+yj5LcdwyipVSZ530ao/+beL0
zIJyi4E6P15Ym8t4O6I6Gi1MmYPgU107u756NEtaCEBCr2zQ4TE7angBBUnMNH5/mPvgqcyRkvWq
GX4KQWD67NrKm20iWnqzteEun/bMyHbtYEN+cUUmyE+TsCLyag41k3TYuvLl3NpIrhRxSJ3wpg0W
1rzhniOVnt4ivYprOgxjUGLRYBX4+fs1oXfaeWxzmryJQgPjrzmEOBZz+U6XCid7duszb5afHa0Q
A6/lD3Jgmx87G3bgF0e9S9nkb58PLGhMPlSbdGKFRMJo8TUPUjQSn8bMWkZ++qPiaAxE9wBGIqU4
RReg3bKVVVfUOvENXI5UKwsacXVoXSy7nEJfT4TQzIkoeZrlV0bnqC5Wqg4QwuBMZEsopX3Vn6iW
SE+Etjdb9bcsChqoce2viBkGWZX4aQcDVdo1mESfEsT3us/S/pJ8sPIl7LRpF2sGgDvOLX3JqNFQ
XEuGBQQ393tXofjxSTix0R6h0JIb3gOS6S1AcAqkKDpY15S3LZfIfEaH2aHpJx1zc5hf2+wOsWoj
Rcjs71inoGph9js4yskGCtALAfFLPKWv1vVY0/fdqt2LOHlsVwhNwp+BJthgqZ6xRhgA8urytCbF
nJjH8aFyTWbVQ10BVzGLQiWUKs4b/+QNjEkkYCNzxgbQMKLqKX68JdnVie8TpUYeZHXZ656EegT8
sCsuvBFc7zy1XXEiDS2GW/dDinwLpqLBUALqzrvZiQ9azCoTUQ15aHt/A5LboMdg0/oUKugCaMDm
/KvRM//N+oa8tApSyYLGbkMt3Wm9DmoKeQQlKscdKjTvNMpcK28Ut5GAUT+VaMFvm/+xccLhNqCY
TtfzrEekDkhkmH7047SZEm3xiFhEN0q8WT5UsKz2CfxIX0ZGTc97gH0s5AdZR6Pifr5ZSoZWNAL7
h2szqiRgP62v4HHpdtPlidBpTrcNn3jBCU2jyLtI0q8sYSUg6H19kA//thPk3u+60joA8fUN/uVH
ofcQml6R04uwNWJkrlrFY96lWvOccfPO09agn3mNL6sM5MSIXL3yStY51V+BaTLMpBYz5XT+2oKu
SAeeYzeHXydTSqUVVbuP60ziy0VrPOkEGAe3y/GP259N5HoO9lPnfoj2gR1brg/EwPQXiRP0Ri7o
+S/kWSDktcCC+0zpLaE6DmJXqNr5OWJizqSJXMproOUpYcLDXlWobntFJBBtIu08poVwo8E5nDeH
utaozxGl3LKBqEAcsqIcze3CekpXOkCI19jDqLuEsBZ3CT+zA8xjueGhWUUvCnHhlvZpf/Vmr/BJ
0Mvs3Tstc342ITkVDoXhMIYoXBZpRap2gD5A8dJkTSHoTUERNU8rh3llH8fzSJq3ud/3Nl0U7+Na
inByHrTkH5GGA8zYsxA3y/tQwnEUVVcQ+Nt+qp2nD0SKe7efCMwEZjh2Gfdw6jlTaJF8CfDrlxaB
hvywbZdD4VNkBLYCoDmn4mw53m4dtA0yvNmmEAusfZE6XdUrhen3BArUp0tDLhy+Xy79NytJHYey
ZUiUZa5gYbRpXzC0HhC06z0hKddp395MvcniEFshN7qmbUZUp0McmcvkTLGAEXZ0YTgBqr0svh80
RvC7qydWGlJxOMWXyO115rG4psLApCZxEyt9MvtVOkwhoZsX6T8LWPrpUTLZ2v916kTSvAUYTLUe
mj0Knd9km3SJvHGeDNehOH7CJG52o4kr7GOnF69Wlo9Y1EEsneGG/7FwZhGlw6RYDqmpyXPi8jAO
QTURtQwqRx89KBcVaN3EL1NV1e8AZsYoHSMuYH12ec3jrq6GdqYXuF96KEoh82HneiX9c0S9JLfO
IIKecnZB1NJrg52TmdWDIqL50kkpgPc9dUVYxU/MoKlr7+75xp6XnDjQdSmfeDpLSO8QvpvreznN
9R+BIZDX8+U0CRzSHUnUxvl1/WUnJhVLqfyM0k/stIxfoLPKUztTBeqoY0FpYqDaHerzi1/gwQWH
dRpy6tvUWkUP82zaDClDyr/ASGuoYd4/XVDLob4AGEtQl8m89D6sjxjEoIqam3UB4F6ee/6xBmKO
htECn4JmgP3CIy/PW3ELJIx/Prz1zz05YXj1DzEMlPszkYnEQ2O44gLDuDFMnTzXuVre3eNxIDRn
BdiQ7xf4w7o/zpxMymyXV3CqJ9i8PXhZVN24FVFIo03SaDWg5GpYrKxV0ro3i8TE0x36hs9+KiDN
tZyTSSlCTVLnHZoChepyQJXe7fAYcKfLOVnkVa1w7KLDHbsD47XfVohrYsttE2DCbY0P5POgJpGw
Dadjxdj3W/GZs/G95xkquU/dXN5W2F4M62FYlGCG247jzCbzKW6x5yVQHX16Pov+Q9N+gjcDCQcm
h0YpG5gNUJ9UftkUR5ZQDd7/SFidC5/0Wbvygh6G02htO1bmYObp6lYuYxoP9yw73g9jxPrimOi5
+HkJduxatynBHZFC/zvkiw9bTW12/h4fBIPkMs/+N/aIO5T6CsHB+qDR0uipGomrvZTdVFbW+iMj
WmrnZd/MdOeY8+cJ4KGPI4GRWD5w6C3nCbhtRyQ3wkn6fTEaK5uHjFDowW9NBgciV52EDtggImiR
iN1DCvIyKbfoXD4W5vCL/bfo+zeAHZvOhscHsIJr/9Eite4I8j/PjLcl1FaOYAYF9hWmzZaaW/+9
v6A9MiMn8Nc0O95wssxH/+TGP2aInSn0TA28eFToGcgFuh4Jv0dfkF/APz8Gk/RPh/KPW463EhWe
CKwjBY5ZbCTia2VgEqgOURFySJSWJhIozFyQcT34t8aoXAUsX2A/g1P9MkOq4T06z87xr/ULACuh
t1NvoLECpyieFZ8MgEJtkMM0Puvy50iO69FJ/IFxKXCC6vcnPyKlHrLAHE13/uTrLd0wFqIt3f3A
ASrcNwprCBbYluBRQQRt2VAkJXILXuPlpFPGdeIGKuNuVKyxiVP2gfLACwDMguod9Rr+AJNvwStD
NvrwOP+uWErslOi0yynvg7xZAs3E5pL2wMvvyAzeWtTa9AJmi2+WbEn4pVxk3bw02GRH9yi+kJHy
lQmMTY85vg+PEKQorvZGwhEdVX5cbxGoSWiScxx++pL6yLRZ28Pmtzs+3mtLl6om/bubiyvD++1n
4lvTIxMWWDVNZ70PBPdTlZqn5Ddm7Gujb2NIFUIRhiHtP/FJWstOAyrMULglULdrr4/ED3tI/Q9F
tQJGEp9bEd2rhaNeVqcyFYx99+JlKej1B2l1eVgYuv8gp1UcDvXMT9rngepmPou5TRMTY2ROW3UU
5elFQvSe1qYn6Mv1lPbgqe6dnJQFAHXEYMapH14hbeGI6YyVda37EjwFAa7xm0KYBMl8cnBIrfiB
GnrmTY7opJ1hEW7orx71cv3CrojumA/9Q5gLueC52nbjf2wydabhVssatrkQt79XdBJ6nsOOTXYo
0g6eMIJGYAArje0N6cK3r7xBA44ACr88FqdTTwX6R2JwVlWV9+SGLbtjrgBrH9edXtgjmTQVOJGp
EsVqBA45w0BwTE4XvaeFDxb/Ew27PP4zLrHrr8aED/moGgEh9nS7hmE5CbOI/x7SGtUY8CpikWmy
RvxGe5iJsgP9qbii02gJEby8U5fPGJ9Eu06vWSM/GUUK9lnscCXIqI+Uug0+0Qw7D+mT2K0rmSjF
iA0x2AaoB923bfq3LcOT5xtLD/ZzYCeN6ImuHE6u12M1p7ZpMlAZRKWi6A4e2itkVFuTjuaCy5/B
NrqRhjwxcH2Itgu3qiqlFY8qwk8g9BnIXngTdzRkjRTu4ZSCoonj33SHTm8mijk+FBuuacNssFtj
x2zRSE53rqOghSyMOklgEEUuN0T4JiJrPyTUcL1Ccz2oabJ4NPHwnEuJnx9nGY9E725YTxQ9CuSv
jHmf1bBB2frTcOREFLMpCgdOcwTEsBsE1/q8yCGRenvneRo3FlG3gGiH9GXd/3fRzOWo+ZZO+NqE
EmnE6GubXGQ27p8vJUaMtfPtFmXY588kgUkqhtCaf4hxpe0mqi+Xal5bjHF0kJP94t5UfWSDyJvo
DREP/DpWn7CzGCPYlFiFaQDkSuRZlvxc/sTZLqyR9zeqZyJUmT1jQYj/WxNVX7XbwO3xSw92faI4
PZSbtQqtT4V2jtSzEKocbnGjO7ONj8MrUWYvgce77aqUWJjvizkc028Qtdh/QHwdJBqHTlbHQfku
n7CFl1WE6A2Vb2/o07S5cHZ/TkhFzTQ2W7esPACcCjzLB/SW84wzqPXbYMxKxajnbvEBXCQXDSzZ
/TMy8WRe/j5r21oMpEgLSIvZIf/Z5x56rnOsMF/xxaL7wCSuVRT4PKK2RI5S4Z0JYrJ+/GqdsB1G
x0WhSVQdQ+xyoh/+Pxkd1Jx9L8EmxLUw/61AGLvFrCvMmn+TjDbvpb8ka5wg5Dn1R6BebXxWmuFM
3tH9uLL7mH2zcHeCXt/GViajJbRyZwSSEoRsSnCRIyRq3wHO4Oadn5brsiiDQy8VeifMLS1mu/np
b69icrh+TJLXamnO9xlZAdXMPQ0Xrz5nH43y/9JGqHLvxhb07PikY+9oI6y8Q3zj8KC9HWKsZphD
VHJeGp/UokcsOy7d9bOyvPZexKp1gdhIMerlji2znIPRYCfN0lKAM6uj7G6uJhHMdLi85Lz7wOFJ
QGxiR/HfVwecuFMr4OXPBRVo1ntPs6DHeg5vzIjMhHdN7dIBq2MdklEGNP2cKjB+Tsmqj5Osc5qG
AtfJJXSfpBmwSwKhYXhE9zIU+Z6+TBp2TmMk5M4kR6YRh3D/NlMqKtJG9d3UVw2z8WLL+tb2X6Yb
Ai7g99TbsQIa2Kc3Qz3yhY/I4yxdPwVNoisFYNaY4V/XZFU94Yz0vYki51IUIfaz3aPn/LN8P2qp
Ncd5F8zGqQ4f2FB59Ojw7mO2ohaJXO7Pi4KanZKIl8KaF1RRqHwRapQgjNF2vYA4rEir9ox9Qr1l
Qc/kHEkbMwfrwxHG5nUlw/AZkKPv2JS22dv7Y3X2DjtRN6YWaN0OjvbI2LBPlBT21gARs9WQGsu/
cKW2msAVXSfyqJruMU0HdOYAt9ptHrGY3vrgYCPkhHDoQPvNGqRp9N9gw7Dj1PXLWP+AV6zd55ip
BXy6Rmy9o6wZ1/ryyR+zmT+X1LQ4azqSErr+bFKPIvQlsa8uk7i4IPIgc7BuMY/kqSqiVgsVY2pa
JpRqUKun8v/py8THzosGLcaUgQ5PyHJPUIVqJxIcWpPgvpNZ94pA3E2kUuQ3rOzfSkVBnCnw6xK4
+HM4BDGvsN+OyvhRzshFunkXHhp2dbMQc/A7tJdOSIuOgQNIpSrD/485ymFpsn248xs8ZKINWdXS
4LqceLPAzHEQb5Wgvj7Hie3VxZdnUFi/k4dcVUNo7bHJ+Y5XdgiNffFMPl/SLhhAvjOU8h1fJu2I
rKUHFhtLP5FP0XVSASkd4tre1rrP01j6M6jBK7erSKgDjcUMbX4K8Nx6Ws/0aG9Sc5YoCkPnzr3O
MikNGkpO75CikmakNYwmmEQMHqlhvUyFTlyn+82ShxTK69lVAm8aAch3lr4W29QSOkO+vKPvlCGF
gkRS8MRHPqhmx4RhUVB3yrWtaqwfNE7daIpouFqtst4fLkCXRX0+4VWtx1Tol16mpd9Xgw3xCVZp
Y41kvriB+ZYsrKyyajPlZw3sYM7jVm1DMYVf3ZzzZsXWEg34GH0byqu41kQhRzvUI35RNNZNk7Fd
wB/HUVJdvtKrCXo59vkq4yqODRvOKtAUX5LQLafiFjBzN0PNAUpRHpKSVvS8ROR88rv4m+wwLSse
4MMFPLFHm8N/CdpduVibkVcjJ2cfmOtzv4zio4lnKEVmnvTswzRqEoE+JlOYnlWHzxe+ZKgLo5RZ
+Ci++1Z7vFGdHBIJ1A+mcL8bwVXsqdRS1epbrVYGGE2V6LeMBUU212oHsNl64kgPw4hIawUmpEzt
oPtWIrabbXInlKgvjj0RMIOEslROVErSsHMYEh6ZT5e2EGsSw3fgqKKn6L1ue9/lkPu9bdQf8y8l
c4el3HzzoI1O5r5KOC2CPb3v7UAdLBTzqsfG5/0m4mUPa7YsBq/h8t7kFHckqafjsZ/P/1UuNT1j
k2BXrfBAJuYow6hRU2vrcHonBXJmrlUtlH49FKXz0sIyX967dWAUTskieOsKIYO3fOKrFIclwt0u
VlQXK4HI65/KukwJU7isf0WUpAHzaaVQtN4wieUa0XXx/OcXzrhZd7EHN9GKpNW6WA8oaMlr8LRm
7DhBSp9iG9XEKB6mQCaupx3c1+M1CINzV3X/9fVXsyzkxZ7Cxk6dBN9Qusgx6YQSrjYwV2ypWX0p
DlQFGYqHAaMkguAqjdat2ZXxgohzT7XQfobfTPlTcJABDcqHaaKR5ZyhXNU8tAhxkp7jP7V826ZL
18+zIBJEF2RMgeOGtJZwhTb+uAioTGxg5Q7JtvQd2yQH4a3i/LgY2ecfAXkoCX8uL1pY1h3JEYqr
wztE8tsEu3/D6zslQCReMISnbjjyiOeHPhlgCql6jFEPF9M1g/GrEHyi3cN8K9cFEyvAGc7AALv8
tpdDSbMF3wcB2dbe+CC40Js0uPtTSzoIRZEUfbUxOqDR+4hf2NbmtL32Bb4xhlYHg8BcDaBPVINy
Yljd/FsKZk1ZqdvhjMoN0ZYwC31/TKRNp+cODlY7Zdks0a9j3fyvAzFiJKFu+jkLkC3X2jr0qUoO
Pc+6ki1D/HDWDEMvRgVbnm9ebG7CV28uNYjl3fwkNLfW5m9UTNHywd1YNgQEHh7DFlKprICFFPDw
UbWR9o5iphAEOVlO0dnxB3CA+WN41xDUuAlgjuqxXwCI7NEky6RVXwPXybq9QI8T/NgdFtR6vtfA
xH2m3kDuTgi1CsCKsRsKkxrx1mi1wZW6AxtRnFA1kjGGwNp4wO6zURr/n5KVCtIxRL7CktIiXDuH
TjdWpsuFbi3TauER45WgjMMQgEjlL2GN/+PM6r7P4DCB+Rq2iFNXnOrQMiDxrKxkM4xIzLHRWNPh
0rQr7xoSqVOYIBXGbCp4Imhii0WBW1spQ+p7RfYwojDKC97/zAKdcUenjCacl/S2uMd0PnCzp5iT
G1u0fi9cB8djWmQb2iPCHz2lLItTUczk899ydCtGpxuD9Ui9uKLEp+KwXnLFOtjH0WIU42Sttwk4
odjxICuT4rnKKjJKAaldsT6IE1m/BHrAba87eAz3eDoctxs+STEZzeZdKJpQbAQ0j4w1cXf1wzks
WkxP/q6NaSuAxqBUS/Mk/+Y5RxrUJdOsKVVtpEmwukT0ntBmEqIsmj8HbFCF3jh9xlkRLybTh1ns
dc40O4/7iISXTRQYjTNZ7pu/ixvZHXfkzXRFwoSi/SDqA/CBNAliCcDRow9WmiYa6GQRBS2WS7TM
tJ/N4Ry/I1nrZhIi+jonVXSZygLF6ydWJPmF72MGvmA6HroBRRbHuf/pWZ8Nz0qjJuQKmSTnPKtl
/q1YyRoxDiA7WeFlfM91KXGM6J5qkMiI/Yi0pejqsuesTd3ZAHhfRx27kOSgTPEDln2/bTlgi+b2
nppnOBh83wuyaQMm45tSV9M3uRMtH8U9HKRHtlPQpwodJEE37EtA+CBHHfcH6dhwfYqVMqhHY3pP
CPCyj++fXYmB9qDHEyI4m3Jv4IqIF0RKLmGN/AOwYg2uyPBaT2L+398V0qlEbTm0CcvxjZ+ySkpG
xGxEC0+ZZO9w+DX84qxXuK2tBzogHG3jTaXJAay/tnp/0ubr8GCm+VR4D9hqBybx4fV1xCqzu3I4
/4nz27PzDT7bVguBNBebNy4GaCjOm1GSlGp+yNy5LYgDlfteZbdIq3zZG7tfoKI4toWkCapJJ3/h
Q0Sc7DP+f/R2w8ivMsemnE23JsgakeFxeAjswk4T4jImbfSCIHbOm2Xl2j3X5YLZxdN29w+0j1V8
qML11ncWqo45Xoxf4U0egjDP8cqjqaYpM5sKZTwEXYr1SzOzimTpyJeAiOvaKdGf30w/Jw7Dct23
QuLNZIU5gh4b1JHRCvn6Z6gLf1IvO8vOq+SP/RLOXWGTtAZsYDIIyvgpuYpF/FYanmgSfWwUGNqa
1KtkgBMavqhT/Kn44jSro/lJrzsT6Z3vtpZsJeaTjJYffKyM2rHkh7AmMYYxEG1nLZgh7K3biRxj
R+zx4OtZpFebwdIZbyBsoou+ULXd1EtBhWW+GZ88nyZqbbfFSIzvQgus9TasabcKXl8a5QP2OAxS
M1N/ReMZFz7BpUF9rscPEVPCLIUEacmwxgmC3uBzj69UW/0MSX+475trxsjwH9faabPZbl91O78e
8eminPp/bI7FuENJnySZX6Wl1NZADjHtA8waV7QpAcZa5ogaRMFfQKaIZhs+ShtezfdL49Lvh6k4
vInomWLmPSy4FirPpXvK4hWMUFR5nPlXlZAPh3N87Tspld3FsJ18oArRpumbphHmzLBWSv6Z00Sc
5jy6sMOSYjVE7o5YgeFX2ciuJXZUxFaLijX0qWa92FMx7UVSmvcBSxQOC5NGKbP599VD/MU5CIgU
A0NXziFFSDvWJoRJ8SMAa9ikZQ3+8PlaYIDh/rcN69eL+Ig/Fxd3z6axq7ar3OFhodj4/NL2hXdh
pNby+b3jG9q516Jf0grd9M+K/kXjRa+cSXUYtvAQoLPzL9cXU0XlBYtnyqUXi6t2QqrC4m9ChXMa
/nfVlDL6H3vTp9W9LUsZIPOlyATPZyLJAtq8e/fhB1bwLdIu4AtNUfUJROnBbpanwcfNp2R1e4ZN
BpBP6/uM+6ba/VwntxSEXi6CjkKx/sTy3TNw3SrufeyubbvhJ8SobNDaE7cF541wsU5QdsODQmTw
9ehyzl8IqEME1x3gVoB1de9Uth8UbdMJ377JEYTJLHrX4N6tYUQakVB3ZlzHNt+aU53YsM1KAMye
5BAAG8m8p0blYGTsjnHu8M9Tk7u8WgJWOmA7lDvaPoJufzq+9h/KzkVL53aLQ5MX+yBUVN3E69Lw
y8Pp4in8LrVZBIEithOElG+rZsNDCXLPvxlTILjmqdWGfinLNP2Ey4EiG0/TWDSc3NMGfy24hfbB
TKXtSr9r277dFGTsYOfne+Ii3wpB/PPHHrVpXnCUVEJgwfJ/YajIDZvCl7yPiC/7TYGyDxIoY2O7
Bo27Dt5lLxKoJM86y4Y2MxsdsGf3h/QO+LzwZkG4qmzS1bvDpj+l1Op3AWnUcnmocI0iOCzq8yqd
MznrTW2ML7LiOpaHqfKX1ZXFHPXMwc6jHqBo5ChiWAXsxZfISzrAFwu9Y13O7AAlVY2At17MdYuw
mapbfU5EFYk7SAJ+0zTDS7o2o9BySGoUCg9ZtdY5VU/o327vqyLmiY06aOM2qCQeXUtgX0KtnN3e
f0kxsfWyS20v5QH0OAdCB1JK88ZTdu7ziRToaFACxPlv+56Vz/d+UjdQntdWCQh9thiJQBt9xAhi
e2FEPTo3mcJ6ANaSplps1wJUDx6Oe2J60FF+xGI9L0iJ2izcJ+UvbZyijzzykX2efIUEF7qnKBny
I5tOrLmOTfSwQdhofcDqMmR8ESFEwEgxaKpU7/+lIonVovT5JP2uWzZkhAuAWqmh3T/3M9W615Wq
4FpM0oSz+b6qTC7WktchqIHdi8PZ0bU9d85XMozegiqokvnMTzVqIcpE1NLGS9pljSKHkA722HSW
HHRME18cd+oZvK3JQeLAK6xS7HtdNkgMjqjJxFf+9wq+OyjcTM0ZfdR6tFVMfErOt404re5LnkiT
EL7TWz8djpJMvtAKBxtUzKw9ebs7//SGjgspDb0GWyxIKFXYobBmfOhOJK7GCV18bgxCP6tOGCcm
6IyyKmEctPQ2b86igjCPDkbrOWKZTALWT5ANOWKr9GWyAKsC3Y3YQ/GSNflkTOnkU+3SAyATUiUq
bCX50Ic0kFjL6MNDQy4VoYxTFFHm7kTfF8psEeX48/Y0VCJ9isz/oxwuLc9oa/rT62V1ymrCbKXu
pzxhII9MEt9EwknRFIKv+YqXm7xgv7R70NfA5U3266ZEYVqzeGkjO8KoCuet+OE/HqSFB960ixa+
OWBr7C+NzBb5/EmqyMNTD7CtlHTgjouxVvWBsgvH0GeHEHMF5OvApzIQCJXvKOBrbOKWEcWPUWfX
npfQ2sT6DyOnrpPgE1weqar767eoc/c0VWJRo89G6uWMcds8Hy0qivCPDHsDu5n765gVWkd/W2i1
rGk64RGbbevogwsE3xCFyjLNqAGvwap9BILP+vC3/HAbFm4+80IHL7FSu7L/C/t0eVvDzJF4E63F
FCKVdrK5ac6I98vXFAG+grX+0eNfzY76BULfTBKNWw6zbo8y3AeyFGLmoNn1F3e9/2tYUYRmidmA
Xrxx5pgZHo5ka9QRjze4wdAyv95GdU8lSIBV9bJ2nzXzXPOaCtltSyP/vvaPwVLv8bH1hd3F7Kq2
J1C+OZdFryBb3ZjhE1qOR7akBNqWrOGL7/3o/tttF3E6j+JDD8YAPteOd3BLJ1c8STHMQEeQj4D7
SJ2BZe/T2kikqUxUXZt9AJOpYJdAQauREod9/iLsaN9UjuHS1Yw180LOScDgE6mOltOwjoEaGteY
+xGKcLqx9Tmc0kmrCsZmBNQ/51ZEk7F9cCWQAoMe0FjHRqKj52kWzKy5bABOZ5U0nQRxiN28iyQv
dxe7ZV3Aijbhpxk0X1VSKB17u1P2Shkjixb7iSzjSoC9mpt3IDdFnkG3Kig18Xv46fa5xwtNqJVt
BzU5d2v++Duje/OSNdYSKXP/qSQTcr1Se+GktbmiJbdyiCq2ldbabIU0pwqFjNfFS3xjDzmafUB3
L1kn20IlnACT5A13Ax0aUPPq8KrP4P+6SOuP8kAU2MUyVPlZYV15YX8xodno78OjmIZQZOXxQWyb
GkZN7dfa0SnDbgbheRvBlfv5e1l7tTWboa/Ec71BOVmUHxevYV3+iERzx0L9ezkFZi90+I+7a1at
4229BmwXfBfZ7VAuXkzy38C0usIkNcmrgl4k3E+ySk5n/MvjFPTR/26kmIFIyxlfud/rCfAcz35y
fnYb5Ttawqb/ebSOX3yFJgRJUeNAO/mP9NN4q+GauNJ+zpkTLicwf3Q7qzhl0kOUlibLx3w04PMN
lFOQq8ypWofgChgsAYuaSMYUfR1wGXP9X1m8MrE8MM5R0lYN0Rd83JhTPS0DZoNtoMfUb6BDf6GD
ybJjDbN/epB6+J8m9bMJrUIfl5ZFTRfY39uXjd25466n7/1oUWYV98RRYBX/Lf0Vb2LbOn9zFlZY
tqucb5428em1lQvqQS+GOoWXrnHjMcqdAVmtormhEETlFPn75wlRRh6HDEd6kCwHMPL2nwPc/epp
3y5VERozMEj5N3WRKAaz0DeDuHVOfQW0ljfAHLj2dsxpQgmG7V8n8Z9CJRI0BNvmVz14IYxP0gLI
0R9MPOSpUQH8AVelaynuy+aZ5UIK0MiRkP7y2+uGmaauDpOM2lQ+3eeHcZtIy/rSYt8zB8OWtHCf
pEmBhPSTcXNBEfuNnv5yrMm59L+xuf7zXXdZtSSKjLK+H9lb15RYuxpWM4+NlwljY7O9mgOMfjn7
iV3zvO1Njxylp8fR8MV00rxQ4a9z7viL/OpY8oktkzPS5Ui8R2njqiZdurnV5yyf7ax43lnsOurI
Brjnj24IM0lKGSXajIYxnUilmkcsqEehRcJOyG+xL3DihugWzVkAW9U/80BotHUoc2tEtme17vAA
h0LY+lQ7xVdy2X60igjmZPU9f5Bn6KmFZieZVfno4A3yrPDImfxvqvM5jZX6hoWNy9CBbyDzxGbi
S/KiZFgC8z/67rFepnbGmIbyIP4ICQR0XldpageIADCzl/eA05J63He0c5ZFyIHg/l48jUmNw7CP
hx/cHRLyRlWat8bRuW8uPxn9V0I+1drXBq++Fi9Vz+V93Te+mWOQ9svSNKzFXPAj9Prqaqp8Xom+
2KhC/3QM/AsxeIJ9iKP9EVgK9/TpFQJzm5Ct+jQlNk2hqTdgRNPhNFDo/RNsQNw3rk/oxmy/Gmr6
pnq2HzQzwY6a8Q4r0C21ec79IZqbMWd14ZKS8eXkYlTDAvDGVq5hsKh17akkMmrCjLVk1Dw0wlSP
mVUphMhFI51VRioE+9g6xqK55fcLqLkuMnar3E/l2lz3vZRuIEyMP8e8dKhshNDZYGPwXUkzF7A0
8llMngF8oiVdCK0WBUWSg3M641JL8mVr3Nu/SbI6bxq0gviCPbiqajYTjm/bpjdQzmLVR/Xsuk0t
TBBjH6MOq0CB36vfI28sEuQqg/ATMeQUm9h6K6zwydnj3JmKy2nWUWRHCu1DWWX9sOchbzlMNkbK
bZdVN3i1/eOqgbvooE3hBU6qxX7zCfOz07QqLag1Zgs9gY+25tVZIbqgArU0u/ffESnvrPljWQsL
xnfIp+VVEFeGwLGEFOCPfV0MTsnci70N7dTjdCgI7U9q603Z17JAoi6iZCOEtih97y9ebLRY21JT
jRYWX3Woxum6s0uA0XxCmYumzWihmrax4RUycJvDaAOdUTDFA0oFN34gS9oxmtKxrXViihsSdoml
r9anh32E3jaQcCwA754sVki5cL+sU36wQpKAfgULHalaWNXHAr4qlqzkclwB8tAhn+GCCks5eRgh
eKM+/bjRu86iJRSwq2vuDc82wQHr4e7S0oP3GGPHR+gQYH0lWZOv5irMOz/aKAA1iSJlJJ8gXoUn
1ika2Nu+1SYPLBnGZ8MgKu+skEXnTl2YxxiV/bV01cjcs7LFfMQ6kNzvRjLc7SwXdx+nbkG90u3M
7NY3GXrSA/6Wp0/3Kzh5nlOsxDZaLwrSgquRZ69/bO+BjzOXplt2XLjdfO6KshkAM5Kho70bCPvv
CrZ8w2qn2L5Ltg59Q2fF/of9zAD1+e+16iIi3+t2JLa1PuHsI5RZgKkdNMwyZ1N5qBe5mLZw7Qw6
76O6yMXBcNRSHmLlAETPdERAurn/cTUfeFxx4IlTPpVkRZKopK3998DHxA25l0duNhpHmGHxq7C5
a5EhD+eJ6HWAEfK7hR2tlMe4peLFiPE6tJFrqaX17FSBz4JsvMqFWh2Z64VKzIvQHinGWvb7ucMv
hfUHRunSOLTj4SHezoIoPWLPNAGvtngW9xX18Te9mGpFX9PkXy0opVNBrJO90RrdJj8b0AD20Q5m
7mGzePG/n1nKa46CrU93oowknDruEvmBtAv2uhzJIhsOEkVysyNi70vowOWBXL1V/Q7oKdNM4vvQ
HEfqblGl3eQHFAc8FzS6tvoorjBu8TNIsddZtzPlrM9np9Lb2IpxII7f443svo9ytbssPLq1aaMU
b20QAmoSbEdL7qrNh61gaih+DzhTLHetnFEzY1nblQabE6kmayiK0hQ58KQnC4oNkoo7mlSHPbWH
Y5NzZf0pW+He8JHcFDjLH4Qn4uAEGDXWMgVl343d1zvc6lFcXiw3+osIAn5o7+M8jxJAOwSLqGkg
kuZwtokecv979qrKN9+SVy0eOgOBfs7fcQ8HDVfj0+IuevGmwRsH7VeeTp7Aiol4eeBFqq+KiHLf
eXb6yCbHVQ3Y92ljOwCPTcqde4LHwurX1MIZ9ydo0ArxJkSKRLa2P/97pj79veHR9206P2yLDf+e
wjIOhn4TO0MzNoF9vrRwpGysRRR209ZM0VIumqrVqwwxXDqEzLOM9d/F3BO2vNYM0G1riskRGrwV
vYxKk7HUKaFFmQhfuNzG1d3V+TupaEtyLQmoaieTq7r8RYgk4ZPD4qRNVKjnxzOZI/l/fFJM6WX0
+03xwkSM/Alp4ZPmtoPEXdGsFNyMguSrMWn5XTCRwujGkeiaQUnOdmZuXLEH7RJksk2l2aOwhQmz
j5tbksAsWjNqZhP2L1bv8mITuZTZ3v7L9f4m0OO+/W00QxmW8pxtuH0yHLTB4mn+qdJ2PKApLzFt
KJnyC4A6LVi2uQzXNDWX4eNmBGXjskzdcR8PpFpNt4NEjQzN1KHFxBbmf9S/YtjB1Ng5rYxVAc7q
8d/3sSrb8O1YVJuAFUsotQQLtUuSpkxsV8STPq+GxxD166FHjUVPWcYoPNM8r1PlvJCvqj+4pq3o
DeaTZqSk3SkZyqAZw4mIZYMOoriqx3qXyBjqHuNHS2nPkIHnWqUl9WhGlHfkKNiKK2qx2R+EzgfA
ble265wTFfMNuxqYG/dyhzFfYATnufYmVYlRWkic+V/kj4eXhHb+QWVRoO2tbprEGifCFLz+9wDx
vtvvzvU7AKOVXl1hZfoOgoUMLWZY6pWA1oqXMf8isLWaB+Ftyrn0cgqjmoC/y3NbNkRW8/7oNk7U
sL8ub0EyAJ1ccdZ9FLCqBvPH+qU+EzLFo/12bnagjQQePws6PMRt+TJeJjWVZL/qLKVsSFqBnUCW
WtcylHLPaJwGzlX0Y6pcqmyNnEgtv7i2ctzIXQPOVh/uSGOTg6Bkyq9uWnUwahqNDpnC6LiSnf2x
SzKgWE/HO89C9mJRIpTRPwHq8YZllk4cq6psr3ZZqaiQrfmfqBBO6ml5Fwc+KrnBqiJaFNF6uG/j
J9oRCZnW8ZyDgHbxl7qQEKoWhSjQkjq4YFzKrNYHTL6hBfT6OroWohwB8rGfUoq3106Yixt+cxED
o5DhXI6d7uFv5uJMSQ87YdSL6RzL0B7bEWqFW4JxbE3KO2u2K2+ibtOID/0IJgn8uS13r6kJwbOi
3YGaLAwoUyMXKM1Xu9kDnmiDyq5lmknIWOO5N6a010bklNhfB4tbFp2LaleWsLtyQjUboP+rxtv5
z3Qs89gpYcDCclSnpI+mcffnwnyU8n6ibPnN6r/SlzxQOZPQJoWK6m0tWoXtpW03XjVYHG9zbYiR
fzm+/TZvbxercoXVWPQCCJe7i2KAlgyYJNIpnEKBos3zPmYkb+Bnn5AYD7Ye0EiqGwUpvtypc6pw
am3+ZlBQm24gQ0k3ugHm3iGD8J8IHX0hvjUw4MJ+sCt6blqxIyyEQuk92QNA41z/+xUkOJzR0n7K
4h8gYIlbLhmbst+ASoIa7i7gl528Kyg4VCD+amX9mX27W7cyir7Wn2oyE+qwkoNCP2Iqc5xAaLm3
NyZjACFSjy4BAZGw6MPISEnm/H0h4DpcQa0oebRknmuK7j3kPFqTE1lOcQx5YbdfFVQlX5jhGO67
bur2OjxQQzYH5bxPNt+xkAbJmqt7MVTqA6VM2MAOyPL69pL3kx5Lsfqq53qzRAHlADGJ4y7FavdF
nCkbq79SysrU24Dl9TmZgJPN64i/s6B4ukkh8mTTI+BX9RJkVMjpGYbVDly25p/n3Us00QL5OZaZ
Wu85ph2WvPt47x7vCG3sI4sZXkerD1ttJTbrAGYqxRpkDIelKj4Jml2vpTbgjO9Xh8Jz/3ZDvIJn
WInccWeb+Yx8YAhkd7xFWnKw4G1AXS//ilCs49YPo64+2dc1veANH6uYXkkUFym3fIUdeJNKOsy7
VkHsXA/yLU15poqXbKNAfmkm1Fkhwtg/xl1f8fZoHO60d1NDUChz73b/Hbk7a6sRc9v2glOTd5v6
W7S9omO4N0NDPJEYwvucAh0J1rwlwJ7j+QrnLoN24x+wcSrvxPa+SWcul8B5fuU4hUTkKj8Be6PR
Hf4lWWWsWmfGGxScG1UfmmiI19fiS6otJpYHUhOq5Cp7qkfeoEWBPY6UUEm48U78OvipKyJQH6mW
FOcQuH5Z04IwuUj4GTrQc0tK2v21PVrkUWOjf1BQCO1lAyIpMQyAY/PBaIZpvQnGUy2rYWvWYlI4
O82UVFclNtWrfhov/EWvn3nNEpS8aqLRsaxqaZUTGTTZI8WNkyWu93uBXDj4CL6V23JHM2nhUVc8
4FGz5G5Phvns6LQqeWE7sacAF+J09Xpw/B9k65HGZnx4aD5OiTi+l7o3f4I1xGOa5tdcPQ/JsXbL
AjHjP9d9eJkR0kxJz1mWIA20BegJxTGF4NrFqV30QZ4O1156z+2e6plw41I5mNx9TMOq84kzFsI+
HsXM4XIn9zQgl8N9n6Cs95fljFrUivTrDGzphY8HqhFnqF5Xl8laFLfecVk/g9QxACeJr5kArVSF
dfUgGkeCf6D8R7EqVyLOAChgGiG2/K9Xbo98t0+ROZRPh79XwO9TjMsa7oAuRkHXGzivlj32TYoE
rcsUG3o1KdWWsOFfEXKbOfqcKiZW3aeZIYloq+duWdSfDoGjTf9E9WBg64SmsQC8sY6SBYbjWuAj
bdo+pkmwwBo8jOSCPbMSxP4Tvuq2pfYWe8xFvN0KqwWv0+g9q9xGxuOvhpoy7wYSA7eWxq+oMMLu
3wITRclKa9+r4N5IJtCI2llzpSGO4mt76uL81dF/375PeDMMgoa6G9XEO67x9RFiSwn4eWSHR3FW
M0pSpT6tYbRrAOACTW6jkwZ0rroDMuXcKluX00jgV5ZzkcUe5q532/6sq3E1uildmpNkm7M8EYzJ
3aKL0fE9GzNHRqcNQT+067o51UULijxau9j0Jg+XfIn18p1CCEzD0qgFkjrlb42obCtx6sxREyTb
AecNzbhRcHE4yyXzoDdWiqyrY5syYcKKIAuXcj9QJr+kpog+A3+rzLqeTDb6iDq/RurafAbOLR5U
E+cpWMw9lapuGTeRs+JBnn6b1nOTP6sW6riuZoDmZ69sn9cWgK8GM4tN7r2iz/eABbkgfPm3gg6q
wNozivlQvbDwFhbKphHfYQz8R9M8eXeI24kHPwWAewhAMJf9TuMZcMzppEoBg9eynDWZrqPlyOfr
L5IVnzgS3iSJF/CCyHWUPLnJpugSxJfG1pAaFkqmZFIyKDNH+2i7yhzu9ut+ocdqEBw+340uuWOB
N2X6czM+y4OAeiUNaez4OMBXNWPTXipXZSvzUm847xQ8UvXO8oZixmfUsIGnPWOub0FXSjZsZz7U
gwGce7r4rvj0xYDQ5mlsO7NMDsoBiuaIuL7x9HQ6oUDg4/6LRuEhORlyP1CmgZKwLfLWYpOGqkZc
IKCjEPvwP4C9e9VnrCkSMrom9hj1oizJic0XJw09diOPOynAMSwf2LCzPd/YVvunrZLK+C7WCL4i
EoUxX/fPJvFQ1fTMTI0AIoHK3SkaWoBw2xfgbuYYSssr0+jPe8x6VClsmXcpbd/uZDqYyr9h3GkW
38+m4WOzQoUOUm2hbj+okoTEUaelKuFX2Z5U0kBdUFEb/mX/Aa7rP4scir8suk7G9ahNJlc9plPE
toD2UKSXExJlX12IiQVt2nQF5WYXHLFOOKbd0S1yRrker+jOSxTZsYHO60NdLdpHXG9svEa3qaxs
fBzZos9PqmD8hkmBZ3JBsDsgTq0V2POjlvw4F1bTqE2SpnycSjGrq6NmUp4z4RhNaq5bpYe+wfwb
HlvsqxOd1qv/tAlCUhg8s1fpgQ0X7d4QgNHLkCZzoyvU1BBqKla2sNixYL3mRwXEyZHEHFIcyLFT
5P1YshBoDrD/cjIckyb0xk2r3zqn1mMJ3HXdLb+I2OgnnTyIC4aLWQKZzs5J8AzH2B0OTkmJ4a8/
hy7yEmBikJRkaY5A53r1kbwlf0pQDHvLBsJiCP5eKMgNeIXVMcqA0qk9anlskd+sqMlAKtFqlLzt
2jMum0JHMqNLby2uDtMSTmWUqyQM3nhmpbwB0J7clQyY09qzL3yU8qmpbjTnccsqUtPrN7XBmnzJ
Vrm9wtuf/SWlD9KO4thrZfhi3fR+cLtZXobuL+wsOpU++S6f89k/pSskorILcBoLW5NHWAdpu4yt
s1hc3sNx0pOUWBu5DV8YyKxZeibEuRUJJ9ayCiWBRBEO5FF2A/G2G4c7eM7uJsw3/a2p+/teCk1R
WGyVvE5dugmFnczUjzDylURWzdsQYCDLZiGOBcPMfzI2LUHvlf4+up+2mdBALG5U/bsrC4K5qLPS
eEctujFj2Jv50tJAWaO9KyUCA2JREhUJ+lyntrt0al86feNWVLl/dPvaLC/oJjvBIGJBowUB2+5u
k2slDvEAWOok9eWcLgxa/dxfRPTl9ORJa0VRCD3HyPwtPcefjR5H2vomD06Qvh59315Q/IDjVZ/d
P9lYvjoBMd9MddbNfX9i1QHVx/R1GxEEehn79m0IO9ElynENGSBFoEMMX4uRogXUYy3DpSLRLH08
NUQXBeurqYSxH+IFxBzI9AWzgS5kcbeEPAG+5A8WID6BI2K6wMshzOvDDbv64ixDpriDx8QgBVhL
/G8tH4TXdfsAo2j+MhFMHAOIRAMamCZuJDz2E2DthQ8Cos8eJYZ3rtVjEajjic+vykTxVy1Nk/xN
9bdjdlEFW34EC6LcAucNhXe1E3ne7yJt5nP6T7hdZRNg9VxEmCo5zLhM7uD3WuADp7AKdGDebwOa
l/gMMPfZpeOJbzZ7Gj1gIk3wgcH99N9Xc288aFHW4BI8tkx+53BVSG9rM5PumaFp5d3z+i6HuqjT
Yb10D4Qz97j8yXNxZIcZCioFCZQUWIFjZcT3ypzNFUA3Z3Dar3i/cIEX48iZkB5DJY/LdYi55ws7
nDYPuUOc8mvIT/TZfOrU2WNM8Wm9mIhFiJI7lZL0PSMoj+3y0MLeDhjL91TzyXyRqjen889MFcF6
/2Cw9+I4AKzofQ24+7lJxV0VoXvuNxir4dsx9Nsk24q5stAuFxv2vaYfKXE9AN6YDXBWZ5QPfRrL
gBGjR4FRkQk3K40yr/cxUaSZ6q7r1wEjyQ610V3wkfNDAsyRpQFhfUs38JIOHMnBQUM6inawvMYr
G7rVDWF/JhHN2KReVOwMPHQxkmIUFQ6mCvD05B0mLHUIzQ7YxbSuJIRlULagMyk1VRgbQnREeFoY
z63MkuCUHPmvR4Awj+zI/kPRYhUBxwtLCVs+oQLOUZ1ChDMgUn3QudxEP817hq1viMSdeqk94Cwx
9HsyXeYLjwpPhSnPpxXHvHwvBOpRbjBbsmiuw3Ru9eOJiAZGBhFUq+V66UHjPzQ8EsIJCVA3QcFn
yKQRY2yKhahqlcIwofvQvFLyzHV5McOcCNj4MLgLPaQKuMAmCUjLbq9jDaN9szqz9WfEb1RqCF5/
Hz84rn4gWh6n03OKhd2vVuEvWbGaZHRVFeRnG0whYvE5k5Wh4jX8jkM21tW3lq2iZyCuCPVS0WmT
sPbK6y7N2yLJ//dH9jfNMVHJpzz/pZMujLf3NSu/gkuvcCOgkfi7acUO81ZQ6vdMsgAfsp4xQePU
JV24zBC8XHxgPht6vRu30z8qJVWF4pq66HrEupgzjntZRu5/i2NFVa3zsxAfmltmtPW0qd0ZUid/
Jay/d3reMZci3uWUDCQWTnJhRs+9H52UxNuz4xpMV6J+7dySxiNvNZXkSqkqo1tmpLH9iLAycjEB
mhRMsbddbR4Oo9u1UBqI0wJpczTOKLc24FXPDwf8n6wY2xC5RWHzGlH0n/8NtlgYCt0uKlQMQFcm
z0KahM2ztiGlMJBUzJ5nTB4+K40f5MAwbwmM4mooN0Ca1PSKL6y42ojd/rI7o6pEMf823KVjVdDg
uPYYB94z2LnZ5b9kdL+tYqAJtTPD9gjM99SCw/SRIZVDhR69DU2b0s4LhitgjQVDmM1yYn9zbh7G
SxNpEzC6+n8fflB630TB1YFJ/UM62wretiUFmmTYRxxSfdvc0EdbduRWzM6dW11t5ZYO2NjGNxUe
KoRZk3Jdzs0TRUGBY/mF+hpWNjcVxHWRbBdJ5aIpT+xqjFkCOu27nwpH3JCHtdRWCAx2hhl2gdPd
gxPhhnB0vf/0q/yGXxq9psRETU8t0pBmImQ4/35n/YUXq1IVdj7xpj3Zq9/IyWzTH2v9yJRYCnGP
4jq85V/MjNsI+B4q2YTjSaYPGe7xjBGzSNUYeRdsxtQ4xLTHB73AaTotwKkfS94oulGvEqkx+CF0
hRUlyMlEqToiDF8GhRWiYOHG54kDFx0eWq+ia44pm71n9SvLrnWHRWFa3wfBvOhva6XwDo2gL9ti
od7Xx3BPrB/iECpnsScEPrk6P0Ny3pThFjMdB5yJ1PYC7HbDQmbCKX/nCj9p/S776ZPUeoPy0MTa
TyR42I/YwrpN2OAhGJLshGds4H3zNxPEmRoganzAxTN80ioMdFiJkYlSkLz+oRq59gBGQCvsbzJt
zwaNqhMdHoPpGajp1beiU3dfytsyNXQTXooGfPTzNBh3fmFSe87dh+CIpGjYsC5k6qBgUp1L+v8q
rb3Pl3AV3n9vRq0EkVcO/F4r65O0v8zxO/U8/v3dXzlYVQZqaOKbY3M3mjuyUgfj8L1OyYhK4+Dc
mon6BfzDQJv3qvvxscKYh2I97jDsavW+6jvvG+pJdqqZpHA4rACucWW8wpgSYrCTLPPX38oGmvea
Q58EYDeOpntyCnyX4rU371WdttkecNee1fZ8I/NAWg+6vhWPwFqcq8qfvm8IETx33D7sZh8I/fmK
Dp0cqg58CornDfGgswwYRcXyytWBYlAOFP6u94w8gFNhxWhsxLM0tZ72ZP9pZQXnFL2vG7fBv6QW
zAhJw0GQmKGGFSMJXEwUCPjttXwBklTJFtmdGCWynUVr+kpqETVfNB+5GwMN1qkrQ3N3hG5+orCB
eV7pzle1qrlmYEoRRS/wFoOBvM5bhnbpaYBgxO31FRpRDi3ScwOfBSS7Y/ngjh1bQWO6uy54Z67U
zxRA4G4hy42xPqGfq8LSsIct28qIS71PlXC0xWXZP0ymgDvNpMR1QLFF/FUTD8lzSZPu7G3uwsD4
vyUfPQLgJ5FUAFTPBSqgA+KT6QxvLakV2xjGlbVr0z685nTCPddRveHA7+DugGXQ35gbp9bUADki
G6XG9qb5Pd1pK75e4L1Ud9XYuKKC6owY4pOCbVL4nhD5pXutK7/+3dXB8w2wc6b03PxFnJnh2yau
s5leyI+CEePKO5y0cdvYKY/c8U2Rsq3yGERyBEuJKsTrPJ3tkR9l53EekfHb+PELnU1bN/bv+5yn
Q4exIOBnjuXEI3ANX9iohH3uWNVCnT7yN9a2T14qPCJT9mCyEt4tvKtUKwnEYX04A86i1xWFJTyL
k3uy3dttXgK99PxRCiO8H1rYjyfnS0LFqCmO3ifV2FkV0Cu9V0dSHUycOSd6T6BmRewDxhrTKG/1
pKT70lyUhYUqa45W6gIhyp8J7k2WKLqJRgQnAzpthJzKtJ75VVEMuRe/nwI5Kf9R7LaPl3fGF5Ax
5NAgo6POTmoglYfbYL5aY79JzJkwuQ878yxhFshFFzhvlPvzGNyNvMP2OT11qpdtc0OuVhR04hzw
fyCgjJ5naW5YwaESvshYKt2cwh/0yWxK7KhMQopclTSgqx4vAqpWoenBYQy4wb0byCxZYT+pGlKx
1Eyt4QAuW9xU20xYbEz8+s5wT2eGZHZf+EE7trR3TfTpWBDrWv3Qm8SqetHCOiAaRW3mA18+Vk0/
uFo9+o1CHtaLV36LNg2LP4t6b9nQXiAHJMBrc2qIpv/raljtsITaZHW6J9BnygaDVBJ3Ma7i7R49
lOtQI3L5miGlEzvI6XcJSPQhA/wFSMIkpI9CikiZd0q08ppUni8TKA7RXJxBk/GUEFGQLXSolmNf
ZhpYfMjXEBoJcftPowYVh6PTABoMKQ95DkF1FMAS9I1a/KBtq1LTwiYVpGcBT/wxvXNK7GeyvhlA
AJLSPSIEsKi9kjvj7kUG1A20lSVUD80VXWVbunYsoc5KWA9cUeXPIJgaX9rMXoqzVUu/MeOCD+3f
BBtk7CJ9nQGlteOIFlgXzocXGn5GvsodS67LcYg+AxX0SYMhUNK77dJBqY/g3Ibo9vDenfg9QRak
l4Mc0+lHKmWdutI3T9kY0A+MUD9F5fuNcVt5ffgkqsl1FJCTs3cBlQbShtIh4XmTYdUs3aSNlXpg
nUSnrgS/b/dRrx3msL9FhdLIrrPNz2RAqsnkBspgTeryjFig+ZZ/23KiFJEf2MZJeoqj2bO6ds56
oJOpekK+59e0a/cC5VlG4p9lUrLuE7vH88lB0WJQhtgHzzVRQR46mKixaXurs4nsSJ3tr2fIq7v2
e+/KSzu5+YAt1Kh+HwiQrzM1dIQ+UkeldRZBzClQ5C9xJt3weXSPZmlpmcZSNBc62fHGj1CHkiT+
sW/1gH+gOEadsnEZhi8g4yOICvB6iRNvtgaEsiPWPyZa7twFb0IZu6BI8XcZXH2Xa8Y+YX8wEkn7
uSAqbzLzP0oCwN9hCgMDrP/xdgM/A1h8oA1b21ACVrkm5qi3VEnyYP7jM0jqnM4vWcBwqrbT/Xu0
/nQlaKWEHqhK3v2wZKzL+vbzKuXx/cuz3lh+TwY7UOXvuTRDN3tnnW+z4YOrwDxuFSBjUq7YSR0n
CDJgWN3ot/h27cMMmcWAmfeC7k5sczkSNd3bIDaw9mxsv1hFBN7DL2C/7gMeqgLl7GZAZcipzCrQ
Ya6Xs7MVR1eGwYTrPnt69ymUMRFqN5uvu3LvzMzYhO82d+yhVpLRE0GQa+OmC+ny+8IvuO2pet3W
Ct5o0lx2yKh25njFOP7NouzdBk/lOV1CUFl6uCttmXOEovzT5JM9YtyfRXLV1A17TE6tIZjOTX3U
9ELbizs/I+U8GAqNDFTiMcOhTCYFgrzrDXkDB+DZCUuxlKLNx3LtEcaLTNAVS5ZJY8E0QyseJhcM
K/DH6+qwpCUfl72vtDJzck3WKc1ugaUracm9uDajm6FoB1laq6ngP9/N6De/zMsX4O/es3s0STu5
L6JBEj8i8LoAim5lgucr1YLwrH5d1XtZcrlCdCuCP02ngE5MQhecJBiKl/A0KjFD3IWqAWU4OcQX
aO0EZRb7FxLAR7zM06NqUSLk88KdwSKNeqjgeogB9p0ogjywL8qsh39Pq9dYSXMB9UF9MrkQIaRW
r+I+qnDev9oFZhWs1a+13CA+5/NWeQexM2nVWXyHuga2Awz2mH5Q3LDwkcolJy25eY0O1TW1q9fE
2bbejYkPuKdh+zko1LXCVp1lVPtHdp4GxjSdxVe2ebD4N+hlX2BFnWpn/ilUhBk+/R6RCsd9iTCv
+qb+fN/s43Um6tVVe9eSCy9MVhf3v7eYaON8Dn8OeVL1eEpfiTjYa6upGkDfwOkpWRlUAI5HcEpx
Dg+alGKj8HZhO3EjGRReIyTSMfxIBbG86C58MO8a/H8+y3l8OiWhEdVSGCzhS8TqqvzcxdpHmW6F
htPcllttQk6jt6KN3QYRevlGSeIrEijcDHJEq+JZvEKpMv4Ylj12a83yeyZwY6IMGlfnd6VXDgpz
Ndv1msKRzydHddW2AtemNmsc1Ick2gi4gpthNPBZYRlN0v+t9PcovMy21gWveP4mnemDREpdPT2z
ZuYx+i9gtRft+oC+4LPbInFFHQE00WmHAG/HkZJhW8HdrjqcJK09HajF6inAq/z3iBH2JeqQyHrb
DXG61+aEtFH/hapTTU3Pf3pNCOjjGfV0ph5cyPnFHubnoXVGnnk182ukJtkrK3nuvedKFJae0+3V
y+bTIAsm/7I0440nFnlVFs7VjO4nq6odYxu6Al1Pif7di2InlNKf6zgFi/f7ixDBmnHsmuHL2oTm
zw1l5y8uCoC0jyD3kUN6CA4dci4ye9yS5lEnX+/ZRor5/gbiO1N9uFAtj09195ppYtwkiNFbiXF5
mxfvlhCiB/RFVx//6xsVeARskHGDe351HKzSpj+/oyHJb0M/FKkYb+iGbJAA3Z6Z7Xee0UzdFSKL
QQmU5PX+NW+mgl91JWtYdFY7d5HZB133IUZQskE/ixhmirVxEsksqU2xdb/l66CeTzXhembYKdHk
JV9kV0qOcUHcwXwyRmYo7vEc4DdphtbIakmw6QOADeuX0hlDINQtzPWcv44GX6xgsH7FQo/vucuK
d7YgE07/sYCoFYmheA2f6e2ogcfGvVlkDvDg4MqynH4a40uOWIv/uJq6Ai2b5RPGdfuW3h0FaiNy
OJ46mGT2mpUUXseXIkmaOJbpCOf/K+kTdHPqwAumUCR55eRSB/aii9Xeafy85p0dghIHV4PFoUfq
llOx9D2KId4SIP/eMoUzbhhnbx3TbuFXSZhme5/GKEM0uMZQqBa/3QSxhJOKalJ+2FZA7dvNFA/O
LexY78Ud3N+WAdyNuzT4WGVvz6foL79xk7w2OQ5FZGyMadwdZiEdT2rN1uTgbUa7iPbJUXRrg3cb
3zKkmfn9eFviuRl0mgqd+ma4k48BPrCvvGLsgScU9LNSPY6sTl6D+BmzzMhjNGAq146IZA7EkgN/
S/daeSKuonaIx8GmWbzIQnTjojtjA1Fncg/qBuHj6p+CIsmSYkcjRlXNadxCYz6TLeJp2BdT4W0g
7gkkzFqAOJ1FwGoFaig4xYGlZEyFQb8c2kaVHk6Hkt6qXPCWN9I780O6JjXYc/kuonf91LxRlO49
ItPFpDHIUmfgy1c015eT1SlUNmf/iYFYL5/3FATL0oJU5bcTh8m0tccZ9cTwY2Qd5X19XZbbm5MZ
1/Gh7sVh7poxqFuT5y6IigNTWPGnh4bwdU1XhmkH5MCOShVZZa7KMALlAfXJLlgTZKIeRVf25nSv
5+oh+nyE7roCYIJGbbDMC50ilc4NRqXjcVSPeg2urU2kT4gUXuiH8RafbJTXWTlZ+Odp3WYy32P6
CaBSltyAGyIPZb+NgtuSJJGPyr4Hk91iXIEFmBL+oK8EkYXUDzpJ0cgQHl7D5uuR4vGMTCybyZ2J
9DHZdcOTRoabYF4BZ61BgwKyUV8aNebQzI1qWP0AE4C6MRJE+sBiCJ8Uf4SiVAIqO5hZm+QXlUXG
4Dvzt4c1xDfvrHIoEO7Ooi/47ixgzffPGkcqXokNvC0bsLzq7eLxzi52GlPY+jYpHtuY8Kqu1PyY
CJgt4YO2RVJVObjDTX1NW7/eICa4vzeywV9myja81CkjYkfFiXPeyJRkeL1S/C7ZG3pZ80ok+WRr
Q6SjKLfd04uXoJKWUc/TvOMsOngQ4cojD6/PD8aXo+0BPehKFtktDvLj5PZX5i4Jma82yTWObHWn
xVGtTmQW1TG3TcHrhAgh1ejc+PK4lGZKjfn1NqQNSsnMBHo9xXdJ9+r5knBbMAqiSY2ejKA+vfcE
MkDAZcmNeTpS58tgwFUuLkAphPqjBW5ozoG5AC2qHc4S6Um00jgE4/QU9zvu1FYGauL1JSMJFa7H
Z8IzkFUsEeQbXGQeeu/nLAiYY/p3EEAZEHRmDii9+BbY5PlYFMwk0NJQELtDWMe7+/2gkvj/FgP/
eFmNON/+yrS6bBJh0KlGLYxDApRtLksIh1Pmu8A0Kp+OyPymJhyN1Oy65o+tLR5yXg/6dvqdMZU0
+7fLMM9b/QrGVIFn/ysQMieBIkS4kTGj9A5hrNoXjq3b5gIVLB0tB3gKg8zfwqPL7E6a/06zNE3D
7kWE6sPKiagcNISGjnXfXBrWZhO3T2b4JzY0gxAlccCZQv4gjKMcpCX0c8ebX4BGnYDiKHg9ieqR
sLKq4QcUYaXxniZ/Yq9QnRO1y4U46yid19VN3y6IItj4HQggSrEZCqbx3WYWCwsPP2NV3isnD29y
990VQcfD7z8ooizvNd5NYwQ9RZ2jlmmQ9LIdQ0JwwMQDz/3e7FwrUNMg2OAimQCyPfKiEMoQl6YJ
tSbU5lmYnZy5+CaMHBA2+vfZdV+f3Vdlh+m2hjVd4n/vhdi7hTzaOdwhq3LaHnkPneYI2Hv01gat
stbgacki7th9VU047yYsFs8DVICfzSWMeRY0MBqCC46hS29tsxxbHS0p5k5TmEjsa0yveTzkL8fd
cQ4AgGsN+BcJIE573LBZY2viHswJbNFVnGkOAuvtC1oxf9YL+fUzB1zbOMxnl7eYfRwc+GRGSZ6q
6nZs4Fvsk6DFoOXgcmHHhBynfW7Tb86feOUZ+moqXlVPLpTDgUg8P38q7Svvqz/KX4L2Rerd3RG3
Rbb9WsSwOpYom7RYZ2mEbp2t4FHxs0z00RaniSDdeqxZmQVHrVAfKVLxLYHimfCHvIe6VRbUmcCA
JReciIteAiInIdZe6GpUm+DEwY6haVuHuO1U1wGDUlYCpjckkR73tuu7kY5cNbtk/eUsKifZ5IPi
1f/YgZa8i43v05VfVI4kBX25A8viGb3mvccVkFweJjYjwPgoqSweRxb+HpnLgxcmgGN8CXF1HuJb
wabOzESH3ahhOlSL3IE1Htz83CmS+ZFWA3y3jFUCRabWqpH4R8kTxluyHamyFuJF/tJZofxV0zGe
OI2o+EyQ9EpetNO1hYFpMH984G8gp9kUGVjnQ7o0HLQMjGkP/vng7ZTtF6BBQ+iXiLQHMyOBlp8R
ifItu/RewXn48QiYBjWB3/rwvyZ2B3FEtgwrcWu6GPFR9KM0/VtKNdqzLdgRFpXZ8J1HHzyuzOwz
ebiy2826CvnwgR6PqRHHlhMN/bW3Zyur20DTytOsNYc+y8V3pAx7+JyCu294wG7Yl82xuJKc57M7
h1N/1n6TL9bshHAQLZ1t6h2i/iEsyaONVCAubGdWyeRDf99suhAQNWZeOB8TcmOYrFLNwtx3Uqsb
AFeMeP6m4Y2XJMJvd5Y2cyQp+tF+XkHPBeCuX88ErQleJ96y9vzXmW9RofdzFqFlCjHIeoVPe1mL
9Q0EdjtdJ+AyWzMbQGw18u7Gs4X8CGcINbP1+sfi43c+zT4SDFxG5YOe3R6qEPykojuSGjVGpOS3
MoIXeDsevTzVJKrS9nB3NWhp+H4Mxjq1L8km+FD7MSvU4T8/q2GhZOpkGBDKhk5LJift42Wx0rHk
/WC/xOHqeAWRtIn794Uume4Dz9HaFhpS3TgP7++8zM97l3DEoEjAfWF42BzuEd9UJrWp0Iyl9ipr
4lnkNk3MEt2NfaCnYBrDb7O0rX9eismjvaFsR1JkEbAyacDJwTPpr6ir1z3H70+RY8byl+Teg287
3cNLd5LWEazYlkJa96Gf+im6UC+hWICllszDhM9hXMDuKBUKWa7LxuLyqDgEAV7R+rD2pObXOAwq
wrUh54w5s8nCwFlYnc5+vl8yrJZXpqkc4JuVUiFSubIlzetpL9pm/t893mwreFgGUj4qbNeBJVMS
q2X6O2WLwj4uuYPEwcxoj1jjXXJDcLMJ+kS1km9e2Sw+QO3gkAeRFk4NnTfY8vUc25Au4kf0KL1t
FuhuG84h4iL7GkDhE17+gxJTi4FeDugbRr3atg83cajgeVwbUWB2oZAZXRd/qADURVD2NWZvCV3g
lRtwPHF/ophkojFGfBo0E4gDbYQUNF2VQ9FK/Fui8YL0nJDNmPEWzuuFqG9AhaFSo/5jQ1dHcd6x
bfmmoy0uS5VrkBwjRAppB1od7YUEdxEuzHBhy+BBcePcMt6NqJmmkyGJgM2e0qcglD2ehSdIjcZy
fh6DzvQrsuxpro5Lky08aoFA+DJGify20pXSs20hnxmcvBnjIfTj1+g8HgFfx3UotdJt0VXQ+1cI
VlOAFJFFR2pZ8oInEKPeOmKeNMOMy0MwjTrMbd7BazskV36tU6Vtb16hWSKuCOLChPeSnE1gyKkH
alLiXmt2iER4ZnNUCyHYXXPh2Xf2LQ4zDyg6LNlAlpfhY5ISEheprorqgk6imiVrrOyciwHp3p4x
YWTypPT6ljaBO+jSCU1DZyfHUzXI7wCcHEzenMHR/lCg14OSR7RrSXiueducWEHdQkG3BYmACZAb
z4T/ASJeQjGQjjbm+h+daC4zSEDhslnOy53Dn5kX3in3GSBPrr3h6PBUFAPaF6QD5eAxvDYSa8nM
aDCX+tLoX6pIGckRoQkDYI6scT+La4y5htk3jgjvpeL+kHNPcKAMgI3+O9kYI7LgktglVegcdslg
pTShvRRmbNxNIUCivuG6N669pi8wcOJPQQpIyoztJRV++Rl8lWhXAAn9oFWnEF/yS0GhC3/8kv6I
3OhV8PTk7AKGZiNdW2N/UrH7ZPAAiriAyEGdlvI8xOS7YkfCAuJsNBBJzC2f244ympIXI7l0g34P
dSM0GsBrIMfiuQLSndXIbgajYe5ldZmyrvZCktiLnD88rI90W0qJz8QcHFXZd1HTjE2M4uK043QD
Bn4m+fqfNOU69PJ9J68IfcrRwrvfyt3TlZIEnmUkRvhN4W0Fl1GM2ZuEGScEiDQ/qRSa9gcRrH8q
mWn0bT+ITsHukVaF8BBUnzLwgIWGyVAc0MVMYeygttDviJ0G5+UkL7QpVmymaMIrI6c5+NLsF5e3
iKaf0ynHoGz787abgacFXQKcJ2reXpLOYPAZCs5iEe6EvuD7Otjw9NtN7rXne6DotQTw8pJGVX4B
cQKbY7NSeKyYUDgai0teJc9tGjtfuqohP9aTtV3bqgH77GVrxRxQAzt/zd/SbSS9aAGgKUjGZ/1J
/3m7v9BzEPkopCopzHJY+naD9xzludHy1+Vz+FWHzlwLUb0nJ654fBF8bdN1Z562BqAc10SDd9fF
No/7EMUj/HHL5Yqp8Lls6hSY50gN2As2CiLgkfICxYynQEG8pmFkPCf+2Wl4oa4UUtbd8JbGpsbr
w2dZn72UIMkfngz5ehzVjH+08A37vVaZIbMxmPfn94n7lHQ67teHg/kyVJUOADFbmxE+lZX42oGZ
sIWgA4j8oNZ9SPEVhjJ7IsUzmabfgsdrpKf9+jxh7sq2rvAnlGIHjgF4TxhpQ7mFUFGQU+U/aepX
hOdqLOCa1sH0G7grxI2hMa4qsmlTArp22CMLY1A3EaM0XOOOaTCCumZTaOrWZznIMqI8975XwGBK
O9imEDu7+/etyS+nA23XZeK8KERdxZuE6Bnd2aU45tlP4vBVstLIHHzZd2fk52uTgxJfQUfvGAMb
tcoQgXSljxS5Osszr+1/+laUGrGoKTnQGzjLqf7lWvI3zsw4llL26o3sgH6aGbkIBkjZtGFEYMfL
qad+feWleqDAG+v6DpMlt6AIxjkHZqLtYG4HbLj9/Hq1WLG5HB7vJZ7fwBwxAwMARDw4uy4myRW0
aSaKowqm3rvcOLXl1khY1YobMmpG/eKt15jR10ssZldIb2bi2HFkcAybcRha65SXOUmE/PEOQawo
XctG8SnGsLIIbQWZq7qOhxp8jkWBtBc6TGqn9aJzMpic4XnY/xgxW5EG+fKkzRrhXVASeySJmOrZ
TzgMZECMbpS16IMMLwB9qLF126BhENlOgPzKIYfNV/jJpL5kF4gZw50Wm6VE3lUwr1pVJq7oRS5o
qImP/OpvWun6eJpcy+s+8XoMtYWDInLpMnQKCfjx6dnDW8c9SYGrvliaOwxYNH+iUDuuk3QzovkF
5I5vstqYcbqZRBmEXYor9tuCfg03kLUDEALHPXGw0cSd5lBclzvaextTRzR5pOzYwmG52P0ZAcjK
P15enqlHb4IsHB4sujP9qM0q3+aQc4mIYMfMSefcUZSX3TCOSSl1LUb8yFHFNsfd2TkSd0AC3VC2
gb3E9zt/amaLOBFizGN5w9UN2oG+22Da+RjxvAGPmWcmnMOhe8DBM5r7Hw6/vJf3Zr51be+xTlQL
332O0Ihe9Bj02VoNfWunTBRks2HuN+i1NsrOq+rKDeR/t1t+Csy1vUCCYQzQXkPy8PiY523YRKts
xW0tMG4x2/D2dJr0lnE3oiWWRihCVNJfh6kXyEtnZvd5pelEQmpztuaZRHsQttcdfbaE7bdEk2wB
G7/PyzuIi90nHhQkit1YIyESxZ0yGeunIA+iXVR8mko9YPm8HyTVYodxh1mwEAnHYdhZ7qYPf+2k
N2KoB4awaMi+t5zvUFe7hWiFFqYtdSSXuwWOCj+GS5FU7Fivoeqw6Q74v/GRufQJcXktcC0g1+av
d1blWtcUQPyQvA5W97DHAiD5nNPE++yEi+B3UKrxv9B8b2WMTqApuzI7VQTlPuClN88a+a6XDYho
a6Bx6+C0kXrIgF2gwZmfbyXL/Biudso30AsvFRJnO0LnVr7Yi5qs6WmpvAV2fMRD9zynVGLjGmcY
Ic4R5u3VVT+M2XBv24VT2v5vYb6AfTKkHMiQxcEZDJyExsV9wbtJK2eGhC3GadJ+Vt/9txokm+pf
85S1DQzpV4SotouhpEnVwZR/abwcUYp1wdhLHMv8cJKx4RBJ3VlKS441lFQb6shUiakLLajyJE3U
4P/YL/4DZSDejGI6Wu9K8aorSLnGcxvqlwQN5OxdB9VHf8zqkR9MTR2kRB5vpc53LpHFGm3zWVsc
cSCKDICRb0xlvd4eceZzwwRvu8YvMzjkkw13DoI0t4yspE51p0g9XeS11ydP4+D0p2rNL+6CMmif
Ya7Dac4jw0Xwui/49WtmuOmW6qXiQVRaq9APie6H9K03TV6W/VS0kPXiZ9t0LZlOznmbyapxMkX5
97NjCNboLTFVh201W/Gt5te80uRVo/x1qjRIzXrtrM+63oBnyzD5jM38piDW90H6hxSDQEDhT87/
k+haoGZkIdI3fIcp7oryBaPD1y1hrZw+1OMactQSRNQAU6XfypLGK/3oFTcfHmzfw6QZ6yUQhi9l
a0tVrryoorsuOe18Rzwf16fwcKvOVYB6PKJfciG6GP3zrZsNv9clneAer/hGVjGJMaIXZElYK4EA
WO2qua9BzsZhcgRj/xMVYDKeNbAY8pDvEebnxvENqgVbglQAOBu4dNUe2HjQJRrmOO2uY4kuPnF3
zbULr5DegWHloJtXAHeNM1KMsAtYmbmVtCG4g2Ni2wXE0yqAj3i97a9cEm8AGNBk710lQk5qqgf0
aibgpIUZkLimKs07hJaHado4cu9aJtVfWmMRNK/5vtcdedi7hf1wiQmfT/KErgIxezHqSLaVqlQB
J/uT5XfnyYFrvRCW/CeivjVVM1w6+OFDPg+b+R0cwu/MasA5ZSIa+g7LT4koac5TElZaUTOg9EnN
nhpHTUkpD3471k5teMBxWseHSYu1ugBa5sb3rYv2X+VDFjLaB5tuh74cCGHUMArqLTntf5+fvE7m
W1pg8nsCL3ExIkZO1K5fhcEfWEhI4xIS2rUPAgqp36jkSo22GGtkrsOJ8i+icTpz3n3puTec6LQI
DcAvUW/lY5/MsoY2v88WjMGm0AV/DxQjO/P1F3qnD6lzLVv+6LyDvM24zcYaGafiCedUgb9Ny0Z3
cFYlDCrdsxvxjxnvkbhR6ZQXiieNNBNmaqsoqnz9kefOxs/yPGCh+wvNnT3jcKgFQot+sGu5e9Oo
O6iQor+tyrBTLI40EqSqXjMA+s81f4VX80ykVrqmOJQVTHdb4lsEZ1nyVFuL1C3GQFnSCzqqDaJ0
B90d9MjvXkXocU2k1KCAg2vjnrLpqd4+atuC96Z8rXZRqYkPktBG+ru1YbhtLhynP3lm6KYz0AmX
TW3a9QPYodVw+xFBoMlAYK1FvsYr49wM3o9ZkHPatS8+nPNH5M5Td86A0y4p/2dgM4Re1FyDKGPN
yo8jx06cscFiFg+BAkuEMEMyR3zYvUVG5gzwsg2fKAur7TYohD1U1MjpW0HuB5UTGbQxs4I6HGXp
VT8tSqnA4GoDDKoa2PVGTx59taHgFwH1CXYZRKyobI+3+Z4/Ip+dCNhiAfy4TsB2Iyb4sj0e+URE
vdkIQXmpHJfProSlROFBjatvI9lkRi4ill6A+qSAeMUXGyC/8J4HeKaru1M8JW2fYsSB+rsNpO4O
OCREZWnbqs3za7LJG/K0tLQYNAJDyKtNsrsgDYFCUm17h+bHuy/zhWqfI2rs5tYAJ0RCvH+e+n+h
/3t9iTokBcEsAUfATy+YUw/SgttZ191Kia8IB3Ek0yY9zdi2T7txysiQKUY5e3+HvY7813ZMAdos
7LAVIEeO3qdRRJkP7jnNNOmg2KCRSYvBU6FjgBqbuv70Vn5FYjzAGXHVcXXftPAjUyPjPQwWyGa+
FK9oiz6IvQSIgmeiihZEPohXLJwO4hczmpIWIIxJYnQUwU6XNEqbiBj31XIuZg1oi7hYyK/A+2iV
v2H8nwSIuLrAOfshGCuo46HkUm/lg6kjpFEbpCJbf0dAkatRqWSfHyt3F2M+4P6OATp28MaAQZiX
jbeksXfymJMtm4TIccWaOAb9sByzp2/sTBJTDA2ImZ2qK3U/lrBKVXYwLnfeSlEuN4TSpNT6ALXa
M2V8JnJfiIm7r4q1MNtp4E5N+WU4AU/JEOBlBXAx/t5wT6HS0+t7INw39rprI9fNuvcfOUT2mQkQ
WOYC/l3JzYrm/kjvOkIcnff/hRQ14pH4Jt/74+VpuYgAhcWsNTT7aTDrlu/DiNJAI9CFuDRH0ice
zkxJBKmC/Kj7ub4AtCgoYLiDvO9f6avncLRa3rdH4luKrtEb2A9iKwO4+BpHt01pnO7IdZ/JQQij
flsYXeD2V68LVuLWKCmNSxhlKuZEUgAN+UVK9fl6UG1Sb3Bsgv65JB2HqWizTxhB2XCz7A35dQGx
kH9HmWD7QehoFLxO8GSDr25avJZXNC1JzjHn/XRwlPR8xMDkKdxpdldOnHBJQ6RsDKf0d8Ii3spE
Uca4bOIicOs70viR76cks/Er4jKCH+oQPkI7EsKuGSGGuT0OwJh+k6CbgP5v6z9ATC5daSoxSygs
QoAMI/ifIOnzAZL9NNHNRmH1KvIw0IVQ7w0nUNVgNk6/9Otd6mD/iinzHgXTJPOnkUcXTfLxCsxk
gG47rsB5VHiqx0g4cm+qS+2SmSeGA0bexVeLd1lAy7oryyWe3kJ4smlQekXF7z4auR5EyXLYnXO8
DOfKyuRzGlMxEGWm+QH0ZzQ8xMMEB9/E9NEftlMI3ROHbV8nNIw30j6GUoemME7t5vayWhpnvnFF
1qWxrCkFoP+1veuj0/iiNBobw8az+B7YuHjv2Cqq8y6pJnHY0T1VEl38dnBjymJxRvUVJ8qwBF3L
YzGU/2Jd2msrkN0ljcVe6NFu5POMBvlPeG0s6tgn7YXxudSwatiK6mTn1E+66RTN3Tg7bOtdGkq7
G/EaC6INjcbh3QofxSWB69UMy0aIIqIeuEgS5b3rdNDbRsfWeuBio8UN2AMUeIWznz+Wz5NOiuBT
T45NSBa6eIPj7g/+UAP2a3FVOBEKSge0ivRQhavbs+Bum2P1axhB99SCWCnk8Pqqst9iSNBq8D9C
1eJ2bT0TvKPh33+MGUg9MD1ZO1jZ4MsT6Z/eU5Ym77kTQ4XmZgYtZ/ku0miBPg3Tq9hWAKGt2r3N
NQhTCak2aVU2PifPI2nV8ZWSDZYBNfACx3a4wPcq2Av4Kf9nq7HRoA4VAlJ3vH9cOKsqM+Bri0WJ
vf+20YfQ7jruA782CBP30YQMoveB3+i/zjuWf8Ns43RSTWv4E4TL7G3l3q1T1aFepPahPB2voP/a
EF4hktZUHeUf+8Vaza2fPBrdn8bEo1Zx5DrA9oZeyATApA6Q7wXM7baCznGppAja485yiBiTdNSE
VKXLTJPPg9qXW3g7QGjH4pyhLLi1Tgqd3zIrc52VT0RVs/BRBB1qRiKWl1C+MHRYsAfng+RzEfee
USZ8Xte7ATUE5Cxb+vNg5ZX3FUQz9C1wi5tD5hbCIk7zMId2CtVt1x5qDNHNoZVY6PzHdu+8zHyB
FEo6dlKlIuRS50K8UyzvWWF9Z5QMBnDgSAwM6J28CcYk5m7JY1swT2tbAerOiML91eSaDunzRr18
4NnKCEPQQkrimx4Li+mntg6tZK4obEIH3QHb02nK7rJ/27AuBlgnN2M6GvBzRrSdhe2nXNg/9EJA
FszbsHfsc0t7Vp8HXlWjJnhtQkgSiWrYh4aNZaehDyrX0fjCSVBr5h9puAP+tBTZX933awDiCZ1t
ISHKm4Wb9mXhRnBXX8CRKFF4gL+VradqVPre5bPv1TIOSVbPRJdpky15MXpEJ27iABDNgFiDpDQ+
WmRci+rQek1aC/nJUiM87azJtoG5vgFhGzBQLohKfKL5ZCsiw6Ryy438Xyb5IHk0tlKDR9nX1rdk
8DGzO5O7/J6h7nLCDmZRV6WqJ280MLRJLDdIwiPK5WPz236hpVr+krUi0fQkkE7v3RVfNRSFiCjl
Ph1fZBNs2Pyt45qQcwVEWXuEgZdURtCXRyJWEKw9GimjICbwgt1Wr1aHZUkXJ/sO5+99JiGlt4r1
uV5o8OhVAcNabtAXlV9YctZ/YfNAiXBQPGjZy4GFB+8V6G9guOUpFc5EgNSq/QmGnsnx4ZZQ7UCV
+vXUcVmu86LD9A3TRlNGwWvIW+Xp3xhJGZ1/XrjgBZlaU2uP1aG0Eg3MoNDdQUeahWkWtFugfGV0
2mCSZuAjC8frskyKILp5/rRbv28t4abNJFPBDUI3cTZKrmMTze40zkkZMOeFrlWzveCJwktghKSC
JXNr/KiHpMF45JGOIZ4J4pdAgEHx8+vbgL//urvcWcA105lr9QOyYmcYyjEwCbtzZ5EdS6UmjdjX
NhaYLecCdhgdrrWZp4jdq2TuIY3XmfOr09E9vcMJD5zORlZaXW/F9zv0G7LQKRQiYHsIsTQPQbAX
DKoftHC3bvQr6QjGYVnWOmHh6OVcLfaYaYCCRXroTce/v2tbd+MWpPEURJFddkQh27WSQNHSTyz8
j80lrOpMWbgwUEMGjJ0knhOVIxk367kBYhDpN7NtzdwM0KfEvUh4ieqFmAZn4Fh41WbKkACjDQN3
HcnL+eGQql8PUQ1dAI19EE3kM3XuOG4o+w21on9UkV+EFYjntV9V+44z88Z96AdHyq1OldDZUI1A
Eb8PL0KFKhJQfA8AUeSzGAQm5nB4BTNkCcxjYH1b2m0nYQm2Sn8TJBINVGC+oDMhz1ISMfMosuIh
5X3Qu87W0oomsa4scautKNwUBgoAPHwVZr0/pDIlKdhDLYOyMU+7s6Fd46S9YmDUu/jI0Vl4xPVG
/lX42wzUF0SRlltYbVnyI91kEi/Ad5XQp2JtLVL3j1zARLY+bkfULXqN8IKGLTnJywTBdSs+TzFf
5ZP78img7E/xuH6QzGE7c+ud27qGjEiDANuITBIEUF+Nafn7peSWwUOScqQEL3qu4rRXinnfH68y
S4jTSBGcbqyPCpxU/oME+ldnDyVbAF+Qw5O+0l44PndVZr3hHFpS9sf9qRtfgG246ck0kEqfc39H
MMuAH4plIJI/it1/w6XW8GIGkd/X4shf28wJY/ZYEB4LGjeR8V5Nr5YgocikSpD0CdDSu6OexA93
IYHzuPY9eypoa2yf372hsuXv+K+Y2/XUMJAo91UfDj31TNUziIq414WS/jPI4Dj3ZCtrxACnmWGr
VC0OEzbAdUdWIvxTLKC0IJUe5wS2lPdiKvJC8gr0mjNl51EBR+j0qOM0nbjkk20nymGVEeEt/+0G
WUTdSTg1ycfUoxfgt4yWHcZaRLiO97NQ64v/N1suvoKsmwkC0ps9eRyao3eaWyD5GZudYKwMw6RN
J630+SU5OLdrB/aCmSqHxiSpxJm6lX9ZCtBtdhzSn04PhkopYq1vVPkhmZHyz1eUCOc5SnxJaRQM
NP7JKZtgRdy31A+fyA1rWN1tzMtX7hkn8D/4LxZEAp/9K/FX2aljYSg4mZPZu8JDdZr4xyeZPnbC
HP5Zsr3/j2xcS7mTdA2HDDwmCuHkYB91uAcQaSjrZuXkHfilEPOTDjlZXksh5Z+yGHB0aWCagml9
c1ZtfaPq+2+n1/dzaNt0JnC3pxj1xK7vRo7pXu09fiS44PWPFkyPmvHeuxQ59j8fbIQePdNtp93p
PgrwLa9e7hvyYpp58KeHTPw3hOj8Wz6lSsle/Pch9CDOkL9L4Zztr0Fh4wRg/RNrMZrbjU6ZO5nb
rEK2DAVovy36r9mA5nhGMOIxxBEj/XXR2iSs+HrEDRG+/aP4d+IPUL2tAObwKuHzVf05iuI92sjr
1GxZBGTT8i+gU8Oe07Fpe0+VUb1TcRgOBap9e1bOvdCQDUgxmbmxLqKmjnphY9IfZ/8hO3ItHO6o
tGbAtTS4h9jlHBAeJ5xaqQIzlnDW+65eh5UGQoI0sZeTACTMrjUI2yrCKhhMsydmz4L/fLXxUsuP
oD6i+oj3Bk1NQUfs6Iax0uaXVIfO3fB67detOqO6pohwcXYUfGbBYFHXQhCmkXVSEIq9tt9yKy18
PW3ps73EY41bF68tGBqnuZbbY1xQqsfsVzHQw0CsxVXHL7rW9n2lRCJs7DCw+p2N3LQ/RtPpswiF
QXZsuSrYvbhA+NoR5gxN6KLq3N8v9xyhdWBo6UK1Q+TZXk9EYLfeA9acmCgLYsehXCXyzgoSgtZS
PFCA3rXiBsonekSV4qXVuONC0ThCjk7E2I7CCn+ip4rgRYmmmSjLjVdfXcW8SiSoNZH7YPCbDOc8
5qftn1mocuPX+H3UQL6jMvgLkom+GR+o3Od+bl5Y+mN7qf6WSapBDj1qdG7FvQS2Hxg0qwXvO9YY
UBginIXr7SjpKgZ9leLfgz3vh/9373W6eF8dF154iklDbBfvYimv3BYEiP24Flt7yqA0Dq+8wBug
Y3pyGo0p++t3/mMoxG1jW0f/cIRZmllKoQt2KzH9baxt1OuabWse4Iq89ZRTN17qX4glgFJR7O9C
SsYdK12WG2n6wnsqwldztTw/oOwJ7SCaOwmjjTuJ9xa2MnV8P66O4tmg3VyGNM4cFc2OLfiekNEX
or05Cq+YZKuNjIB3rV5Jh3kcuc6CC0NkGjN07UDlqXFS9VEByi+Tr3Q/b0aCadqQYzpT3gnEG/e0
g6txf/U1A5cXLIhx0MI9himntptnpBhkEIC7V01D++n//jAkQThJVUeB5OSSjahOqhT/3PUiaF3Z
HWnCbvry3bzOhQe0elUR66eLIWyYmW9sFMG4jQ3M0VWh8ZxhDeGGtJeNUspLkUZ9/vMTcRKlCki/
eKfZl5UpgCDLUZ6ofg08BJ7wkC8sAnCXDtiS4U+Y+FIUpntF7WaZKiJwMAe9WFvL8NXlxMMiATG6
zXuKCa6j1sNum+6ARmhbjEqVCzLSsB2vVs4PgdRC9/M54y/KQ3AVdKL+rsN7o0ieB3BVmSUaHB/Y
rsWKfrXDqwhL+Aw7ZNRxeS/vdLIAV0qOKD8xm8MIeJjd9yZrLlu+f68obYGjc/xekv50TZlQ9VXk
U/XqbNf3dkkcOqmOaN+5ZXYGc7D6mjxIQl5LAxVAsHzIytOGbMhns+AE5X1OVoBmaot5XlPLfW6d
qFGJV+eE4HvWlrXhItUzDKhpLuNdUQ1K7MIe1aYd37oRIfYZUCClxxy4v+p9hsV5Af2VZyeegFQN
YIXsf3I5WMSVCX36ZJiC4Yv/UTq4OOHxB7O/VJJF092SAUkpUCMMOk0Blkt+uKYqdjDW/mqPgS2b
MR7SybN6fjnAJsXEJz+yeVCLOR1GMd/ow5qHYdu3ZENXn7LcKMgyfWA3jRSa7xfQpOu8akUNaQi7
bIoSSHSA0NTv+OGDWgoc+XGREeyYfgud6X+9vln+txDXK5kg8+cLp/wfLQdWae03Wxp8f4i0JiIa
hcfPW0GKyLxBspxwyg5bRRzj1LQ7mTDcUS98CyE+36xKLiToM5fGD5SSItOzOLnZcSCDzKO0sadB
JRjWfI3WRUpaAqdBEV2nykDI/ZLihj2IWiT7etissMDkRNLNtqNVjHWAH6oT8bx3rnB+64NZxo3H
3bpiZxBPjCIR/es3QmXMdZzr7fJ/0mRPmN8qv2rKt5SuuZCezm6s8l77Iw/0uThM3Pb0ik/6QcgY
M+mkBIHM8XnrckZ3DuDZnjUp7629viPFnROGvJKdNLhXh9JQ6+Z8PKqr24QZ1vXHay6KSnE5wona
sXzn8shYioFgiTZLwh//gEAOZekPD8hrpm4OpT/6y1G7ksR6DpOb2B8NUtpv/j2JK6vzkO26wEHM
QYCmy4aT5gc++y9104qd7r5wNzXrREEyYbuqfVCkLxxAp5irVEijrgGjrBhY3/+hAq9EhQ0Q+mRL
WqFMn1lVP6Wh30j7pth8rymMVgkO3GSrArAyq92yOZ9AhVNZn5vQ4ZaPRRoicq4rXmaOHIeL++oz
c8cb473L1eInrHNeriUpeBIh5Tel4RF5pcc3/Suyajgp+UuXkgjMHci714hUTYDrhjzjHh1bPQQW
WQtdhz9jkFWVD3IUNNsBXsQdryvLsZ6s57k+xWXELNwkmyDPzaDnRuxUeGwUDQZfHHXb/WMY6eaV
tAMDF1VGqyUWOgaVX2iA2LkxP8ZouidR28I47ruS1manAWwCB8nlTfcUkEPsgPsqhQEkf9rWrjdZ
0Lvbz/eokbZYG5GR4ivPSgsWdIj8jGeEWOnhA4tTgRr9FDFRe9totUPc9xAEkms+RFcez5Bkuvq8
CNhsfNUmcR+YiUXSMBdLpt5nWj09bCIC9sSL/CezWbjLob4IoL7k+30C8XTj/AJCwHcF2/s4Y37h
6xKopB58cD+OkfAsXY1GjYSQho2DsxIh1yFKwjI9u78d4i3oub3dBrd6O1cZAF10IWU6V4GA+Jww
dM+C0R/IMvXXfig5knKjfvaTWHL9K0cL68GzTQC0Po3vJRhiWQizcWbkNct0IJpnn7DrQgNy7wZA
X4/GWLWfg1zp59p9ZTw/mv3yEb1SEgmEiv6KQiemWMzawfeTH60OatUymN/5OqNovGd8WQn+xfix
EiS3G9l1ynn+L0JHfZll3ly68FQb3J3CwDOHPJpakZIoQxY/PxAAvNe6fRS8TeZBHWFU0b2HVX5z
AyEllgvr0kaD/2IqeH7A8BL7h5iKdmIKPtsfnXMxShEck0ZB2TRV4JAjJHuPxHg1JjOcXy5y0gX3
KrQpasb9vydKVr1w7X+tPlBVo3v3ShM4Yhnn29JJ0yU8JoBiE7eSPOiZQSaOFC6nJGf5EtaT7AMy
FA+/zaIs/E7tsnKL7DXXEdlA+gjiS+6tQZKNfa/3/gmTmo8R5E723jUxNN+a8LQHVbbLdXsWhqoH
DrAkjNyHjp79MeKRvT21jPwpE6NVJHI++3X1Gezvp5wluCtFWCRnyHaoqLwDSya0NYoyBfEfUoFG
rRolKdIDWiCY1wE2l7XvuU3/ls45gEiJLCc6IXr6gNnz2uYTENxV6F1bhbtSSpQq+2MnJjNEVkWC
TLozvxab8oAzt463cjrUCHNYiN9MQ0iABCxxMwy2pDTV3FMmaKGtsLbSNgtPuvOBmkzoBOAPWPyZ
2jheXQ19tFpbg6OPCWxpDxzbXp8WqX4xE80Oa3Ux6V4oiXTw3widyycATPA4hlnIY1XSD2YAjJA5
4xnhaD9q9iDZV88lNM98jyco/zYTSWYU4QTkz1dtmmGHNrCXqWARVU5BV8cSkSmXfD5hwy+pu4f4
qQpGd1F/r8W0Vz5Ofv5UIWw/R3rOUGMokza4nNJvD6p0b7ug+iNNmv2N1DmEDIN+QQ4vMvszHacP
k7bHNPnmbPbmAaCBFvLJaX/eRGwHKB54SShz4OaLkLQlkBzYwUgbBWWHthFrwcy00FUm23BxZM6Q
Nf6u2QTE7O6FktwFpaNq0JuDJprnc8e9GuWBQWEmzJCOOS1IHP5cH0feMl1VtqnXVbCKCK42Jz73
xuW6SxeDFiWwXPlx5KG7DV1Sf1nsE4cpOnmJY6verfgconwydnxDHcJWKfUPIUdWiKFhDmg7VghO
6qEtw3RnsuDee7VZFfnpDBtuAw626+udLSH+HIDBiDQU7B/9Q1CoxVHynBsasSdBK2oPh0Le9nTN
Yy57rsRou5FxgZRyT98u7wsjOtCfqcNb/N0lX6NFSmjV255Yo5NTY0XcKgKXMaDeQG0GIPHtLcZ/
wu464UVhaTtuf+GihsbnfdacJ9bEf3Y4PPn9hzJJOy9aSEUMpOwtuJNwCH0pbVYJ+OaF90dBsWfE
rQgpufd89LOHYlOOLyt6hMIXmow2VRJPZqCDRwHdKss3kuv97n8WbGJ9Dcw2oJxp+tkJvh4GOdIj
Oc5hoSho5kwrnGhjUx/zlwNg4kGD5jduAu98JhZNCGMv8/B/JZGuwntwsmWLmMYJ5lJ+w/PKRXP2
ej6uOcHdHu/KDRKs/lvyMw7PtNPPJScQi9d+WzkNl/5YxjigQh+yswX1mPZ9I7l1lmRpuHwhcyHg
w5LEx7cBtAcYPMYAv+n3+NETNZ5g1iimQSxz7WKKRzdtIpQrnKn78QQsSeJsJCiKhaM7LeUCtGHX
DnTeSfpOvwoiukpoiscNaPxSd27Cz5SI8mbOmYx5Iyycccx32/LmZTrzsF6+oD3PWYfs3rdXMqPB
ilyHd3LvuErabL8dy5uRGx+YeEp3HnQQ8ebdeic0oT18Xl7DclgfpUsfaJwLmxqfXfHwoiAcLj7m
hY9vC0qZp+dCHGTxbMPdqLRmgB2eWudR/h73Q5/XrKUTd2vr490Ac+sWn+a1g51cfEQ+Cu706bb0
RP7SXXbaL7YsLhzvCfHu+wo7K5P96+laij74lvaJ54rs9gfCgzwo0KLBf0062weqybYzsC+zHCtc
lTtksc784Bdf5A+Vo9fGmTyoMU94fccSkjthfwY1KkYZ8ASgwLUZd8yg0jx68H4cmArlcesQRslp
gc2oG4Bq8f5EmuGzIUbiSvLH5/UPZH7piUxl2WF/focL7rSv0oupd3Xok5aNl1Z5Pl9VxpimRzmL
eNdbvS/5iKdEajBZnIuMnJl/oqV8EpR0Xp+CZ3V0kqGaLtsIlKjwiaZbm8wzmr2BV7Uf0Pxg0rtK
hOO65bG3W1pIYbRvUumOwX59VJVO7oPSeicnZYafpjbamK3uwkFkqiNvy6ihD+45EKltuspyBIUk
dEjsDNq1LW8dFdfAJ4bSFX3xS6dYdTDuBN4qo2eePTG1EvFsM+zaSV4sGuYQKxhIGmBhJU4sgwBK
AlC1GyPqX2Hrh0g3Pa6/Necn+SpJusD39kqMH6t3lzlLzWtLIt50yVda5yuGJRBtG69QM2JeEQhc
BSk+TFEfuT53iOIVFVUhtZN7FUuED74WosNWp9b8+ikR5YZsiBMaWXYbfWVrYsPPn5AZCfOYPeMQ
MbmiLv9vXsdVVqT5myKckLn0hzunppbMkGFgRe7Mbg+C4tQLTCyYWhP2CKXwugjdGWamDwBG2tma
eIEYjmHIBAlDPuFAQ3sLb4M23A6U1mIpQZH2uK+Cq/jimOGLdn7zs5+ZZzmKOV8mXAgBfxP89bo9
2b+ph+pe/KH/z/NUe1VaPiCw8L302skV6tKegATMPYejVbr1H1G5n2/lxJyrFWhE+UtCc03azcKs
cMZyBZ6J3nbDRowntnjiEmvuZr0QXWL8tRA75AqjNHXGFaGNzgr3/+W49jbxpnxmg9m3paI+Ou33
+eUtjlipHbrGl3cVI7Fy+uIBokyydHkbwg18p1cQthJUFS1yEo7qpJs6TI2u5U3OcbS1YJvnAYFk
evIb5snTErH7jgUM0uBdPOJS72LE4nashe+P3H1hHgvJa4+MGnWV/79Q98CN8pYFXW07ALmM4sk2
Ejjq/Z/EhiQ1SIW9fRlOz6EeNP6gaS5cPzJPOLIYw7LO1BmJ7yxDbeE4jWuZjAerBIHIwDm2lMQ3
GOm35yZjS7OzyQQYocSNOMz973j2Pm8oeIhds/+FICfqtduxuraOk5W/klq1mZgRF99g7Fpo7zmY
SyU0ltb0gZiBpSrodE/NSDTeLsuaUXCCCLscz5pnmDod5UXbyGhy0brohreKCteRJn0dbvwtABEb
g9T6NZWX0p+eb1iNM3tuaoD6kYYnE9GTUNH7VANKirujfnr+iiMe19iOOXbxCsuYBAThYIiTdxK7
laqXiixrHH96VroTK+q10DirKYeotkZetfYXGiPzLif7uQx/7PLcqUUeoSKz9mlA84eiMCo8Aucm
+uXVGcfvwAtm/o/8Bw0uFfwWBKQnQBvVBfmCKYafB8/dYV1ERG+YtLTteVJnuxxnwQFVwtEGEaXg
Q70XqWveTFiiixODkMnCKL3pHq52Ed51s12RGwYYBLckoew7OS7Hb1FNRGPRaAMCzt20mrl03eMM
/AjoPxOqNwz0Cu4yZD8Bz/uXLM5x/oB3eJ+v9pBao6Myjmj/a54G2/1lb2xJYhGg2ETSutmgXmgi
WeMIvr/Me6118HELo/vcE8s9SHEWZ3mTepwNjmRl7pz/XkM3SG5+yMji5Kvk7d2B7xQ3TinuLEzE
4WO7hnZCC+ZVQTPv0qxZvCr1b1MaZ0g4V9qNd/A2pEEJhJf55yIlR1AzEDizqxOf+fPChvkt2l4g
gw9jmFmifeEqULq6hTMlG7T5MI370XCswSkWGZtt79QkEHngUlsNjO8pBC0wEaCwNritHhi5R4YR
DMESnn95M3iX4bIFeUoZVhENS4Pxm+jN7gKVt5W1ZNyPgl/wN4jmrSt6DtIg61KkloA6ERc0BcRe
upWy1fJneD+wCazKO/w9UGxxziLy1ai8knqilegNPftcwLZkVvLAZEod+o7DzLmwWzq2UmKKbJ6h
8A3GvmNbhXUy+/u1rcFYrkEOAAWqRzGfhW2Jm4Ni0eElQBukxBcPBAgnpvzaDeyij9X84EhzzuYO
r5u9NqGWE8uCrI2aAH5ltDYr5opLhS+DuplLPXyT3QVnH1TrIeRfvF7umziF2A1Vzoqocn6K72Za
beF6xFbJjmJvaVlynCbJF4j0nZWUm+h3MlU9r7PZwlZD4vhZNj/juRFLGHoLP7wmO9eQPSMsMm9/
AROcJekGg+TST0xtlyIMGW4YzwNqWUdy6FZYa2BD58oHLkMBbvclnWS/n6Qitb8U6MWgF5D3Iq6o
TV6ssi2KQ8ntdVcSXrUedaWJnO0UAyY4Cx2u1615c2o6sd8fyf1Z4tO/+nDBWupj+PYuP2aOgEne
Ks4DZleR+6n+o5XtGeMSqCz5U5DVvKmVz4vNfj72l4XmtwosdEE07bOEdBhMdLgsRRNBdWxRRIFi
1FS1xws5cYXZZOogHsIIOx2ZjvRwitgk7uVeOfpmZa+xnJp35+2ZzJTSUQqAjyoPn81GfRhWNFbS
CXSyNk08fSNac0X9nHgc20SdRymf/9Bvm6jAWwuYPBjwqj7klBUQDG80codnnLL92sE+MT5yJMKB
anBBMhbqqnVnM7KpuqixyD/2OmBGDgxFpSrtUVob1d6zn/5/BvIYjUzPy1f6eu2I7w4Wgq18TzO5
ql0F+eOdBf5/lhdKY8Y8xgKZtO4BGaJQR4vowxa2gvghKzKsUaVAqZUFpsKnwrm1ACGDVrrYP5xg
pRpLPiLDo87VeCccmwprCYsM24RsxKu5X0vUMIhWtRPro9kzRbODp+oeFKvq6gLulObFimmZvEkN
L09f2qL4fhrey70lPVRECuOegtLgkdaoZf00+7jMHhRPf7FdOWjKaO1Ox5EWJx1FYXiJRkmEdyxl
Itx5Lm0xu3eI38ZsS7fgSyexRggjuyvK5vxXO2Foixpw1KBXkZ760X4x0jM1vAR7IHXdSjcECT0b
SY2i+5q11F/Md7YkdKXWZw6M1gGEir69Cl4lmFsHYacDvBCLb1OeVJ1nLukSIwk1krArlkv/MjVe
guTPOXUgFJHmT7htEc3HWPVjuWdkQ6jUhoQ55UUxvMBrqarV6IYd45KKmpshs4rVwshO9QoO7QIy
Lc40RWrZyUzBvVydW+TQUrp4PktkXNto+UqCgw3xwbDtvkq//p9gYD3yJtGaxAzUIlaM6YR1WUQV
+QJbsFldkDENyBm2oX1S/dvVG+3qC0PwmKLv6TXs5SQO6k1oFMLEObOAAXy1pzlnsnmCfoTOBwuI
SLCfp4cWWjeQWfJEdoigCoZWomCi3E3k/31gXcdiMw+e8tYkCEyZ0q8yGWEiCduqXbmvff+UpLvC
p40FI7mbJaP23jhDBUb6EBuQJpYH6BqcNL9Lwe6OyEuR7Pkk3HJj+Pi1+Cb4PS9hLsbf1RJilG9b
7SM+XC+s0G0ZiiwNUKK0LK5Vl7XlGt6G6FXvfUids6uEqwBfNRVCT3BLG8U6lnpQ01iB3Z/uFH6t
qwdt/rDoMtTJQj0N2wIBTdZvD6QbL3G2Bfwbw1i68itMc2kk91WozP5cpPAvKh1WQj6VX3AKOHSI
Y3T5KyjHu8Cn1+RoAfH5ZBTnyd3QE6kNXT/+F8EZ+MoZuMmaiuqXVtsUjQaF9EHLHmUxO7XpaDjp
4z9R5EnkX9uKuDoddjFu1ui3FujkcsZYY88gss/9dLPwOjgN7xR0lac2wfnvJEuzcIR1V2Q3Q8xG
A2DOH8q2fCeD0AuHbFFkcfWFPi9YRQZLrWGWiSI+K95f/oAlal1XJFKAvvUIzqhvc5kjOKweu4/A
VQYz4eBVMrEGgJjKeVkaY+KZ36kVvBFnurBmvEDZrfVjBolxSHoFGHQ9s5TkM+c5fbsodaivvLjs
RWAg+BQoM5OGnlGYWsGgLYWn4x5/hV4eG23OhyMz/EHSu4bdhP3uzhArxfN5vrfsS1YW9UZl0YSY
YUBh0QqOk1btHxwEnudbnUCRAK3gHs+gvPZ5kqv6lAkqFpW00fA3evYf3YJ2v76U5Hc3xpm3HMLH
h+XL+8pVaZlMSyKmvNcAwS9eI3cM4tB5oK34yYNt2SiEB9JaBbKmkgHjfhEy0Xxs2NKU3lR5JGBH
n+iX6laBBIzQkvkc+YbLcIAkWge/3McYUtZ0LQdXX2Rf0FMHKPEqFTCPXb5hCog8qWEz4NZOGJtk
738k1FfmdJQqGnmJdK/Xjm7GGKrZ80myE/tvTDoUQd0ZAsxvjIoUF7sUdw5BJj1Vz6mswH3lrmUI
sI1D/x4zL1OXOUEnBgycGXlhbErYHyUA1IIkAEWLAa+7Ip9spMFQ4Pfi+jiotJVPABzsjOqugSgb
I9dqDoG3T7V3wHfgZIG/+59Buoh4EIslUUyLfUkNhbqj16BgLS33Pid8DWxwLr5ueLoD42clUXHr
ZhdtoasJmPwGZohHf/Lc7zlBeD5SGaEFhQ0kAw2l9q9cInW/VeifecNfMd4WnO8jmqSDv0WGskrb
IeMfIiH05D+ZIqlweFGKbmNoUC9VdF3tH+c8y23V0S0VgGQpUIK5ey2ZyC3WvxsL0UAg0njzQcjP
XtOVZo15ZHAGh4TPB0jhKR+7oQR0vrE7RFISMFwZzTatDacQ4ClQtetrP20ChAi5nhXFNIUCdEqy
ouEYOo4HEYkGbF9Tf2LDPLZSyBSi/BZGmB+3LeZgvjq8rBoS5LCVoxrgJzQ3noEmUjdVYWBc5cy+
Y80iFrPeaT41Ve4GbwPaQtBXAlf+xbWCFFFUIuv8Tr1eJf6yEoxo84YfLVn9ZDWwz63uu4htVH4g
TgxCjOmcdGuQ9oWg5NUJ4qFN+VbUwuQHeyjW6Y6vLrMiKV1Ad6aW6Cckdc31RUIag8m4BbGontZH
CJZ8sIbJ6Cq7TabDE8+FeZXO9Vg61k8LOjANHwCiDcPtd2d2uvrzd3zz2uOaacipa8NqOy1dbEQ4
VnKgtmC8LvJu7XCtGPGkeg+6vEeKIKqRyVQV3NeFDG2g/ZWUs/5RbiXmkAQSGwj7lhJ/pb+/grKe
n2LFEsDUShv1xvuzTp9zzUR9q1dqlOtWowSpCegnhCj06+8Q3rt8EsQ9OrtzVUwnt2wWLt8i50Su
z/dyaOVXmUaL3JX0cJoXBwGXHscuUDNkHLU8CUpMgydWYCs5F1IrGaK/Vr1p8ldYutEz+pevGoLU
ae4wvfvfrSf4EO3nveOIFLiViZ4wu3hCt5BLs1v7wpyy8kTWJLHAtqXxVPxCUeOIW89XIxTl78IQ
81BLMEasxZGqFVOuTCvJq5dbPX3dzvgN68QHu4GVlu2TnLzUKTD3ccwZbU84zkBExWj2h5dSHu7Z
rKOg9h3MU8EnSNuhjHUOWtZdZxV0Nw8KAVUOtQ/ytqGf7Tvgbcx0vEiGNI1c0IjOHvPUb0dLraGD
Irzgzv18eTTKS7xNpK/e0iXkdN5OIL8lK1fIByTkw0V6mN9mCAUSU+5AZyWYTFJqkU8G6Z7imTif
oPqqGdWEF76n3oWzBi7oat7vh8QY7WOCAd+JRsrZl6hCzJ/otNLxXx7wTQfyBi1+mFDMn7ZzDY6k
b6O6NPCi5KM2rESM3YerlxfW5QveH89pV5r2byXc6oeP4BFbx8OQub30VIa84HTW6EGZN/lWrDTM
0JejqBhoGRT2rJGRLpX24lAK/WpB860EjbJLR2Ket5XMCXo8gWArFiLfTGQCJfvKtSvg1y0SjzU1
OQN+JEEStqXo2QOgD5CVTH3nQz1kDCp+uFs1a+wkQKl2J/yLiPnYvXc/CvZ8PNZl4AKqkRJOkqD1
yZd6lJ42h+dPLJMI50pe9XBswoKfN+qu//2gwoqww6mIflQZDVgaT5fsa9eqW7eGaoSH+BcEJ1qW
iGEpVIZNFFq6TNS/kOwkZynohwTDfYa5e5qOUYp3gwlWF1gNw6GHvMPcsR6itwkYQP5IHjKDn1uD
uMWub1s5PVM2tQWfW1+bx1lJr8EK07K9wShGV8CMulAAuw2XSqNq1G8wBfoQ9AiJiPiaTEvf2XM5
oqbmoG9ClGIirKzMKlUjYTq8ebykSzsJuvlMvRVVeujTaI8gPoIvyi+DPIHZHXPyQNgjtXDjpUIH
5ylG5WHPrwaLaX3VbP32QSzD4VyeJvaV2njx3LG/J/4RUYG16bJMCBMrTtv1RCVfJuosFevmBtAD
QkAMWCWu7uHU/8yFEl6I3RcIl+zZ0AEWDoS0UxAdgMlJQRU34dEg2HjDB5LEwWySZr8NEW7Eqa0W
2qvEpO8gVxEFCowrCjHjSBeqYP6Yn3jwtSqnQDanDHwbOmhRz7bqyW8HIj+ob8VRBNpHjVZ57blp
Rbx83vQwpsKZl5yY0fpHI598cOTY6NDOmFTrjvDnC54MYU3Q6oxNV1TyCdrlgbyYUCCnB89dwQvY
GdN9g9K7zlJH1txrCo2h32BKiMA83U95THlVLR3Zuf0MLlk7fVPd0vDqfoZuI1s2DzI0e4mB6/eC
+dgehcS5zteZOin5hCw8A8MuRhtgE/WefTJpoi2kMF1qlVQgr1mzL5GxKLS5179IK2Jgva/e4cs/
kqOEf1TibTdWMNBN6mQQLJ4UUl/eN+zBCQs+PmAkVk9N4w8zV9jDlEN5sOnR8FDvtnF2Aryf0Lhn
s/rpogg8icYqhVdqFhKFfeOquF0eH8xsvRpER8LzkWugA9SOtPz9p48FqSzjnPzfZDoQZGKZhSz9
p8v0D8RldamLuDFsRmEwK/n3a2P4k8clNO/umhhz9aYnLgvM7QJyaIuj6hxX0Al+jjxqUmGKg0oG
zo92PhEnYVPMJDxr4eISCse4XnB62alrYJVxObqgSnlYHYylyzfkb71RYoIZjLkMRJf1jY0pyJ+R
pwKYNWyuL9t19/JKlWqHaBMwXsjgToYM5Lmjq3rvyTqkdEqCk/HCHtmUgwYNyVESmgQPQQGjrwsW
bR6XwVMwmq8Q9d8nbf2tOaKP0IBXSds/QeFQH9OcrMnvpNXZOruoX0cfaJyxmhK5lqD6J7y0lAyk
eoEz/e8jB/SlFyyWq9p2M/3wc8ISevbtgPXtQ+bTZCOdULxw5cuFZ0/CPokSK7XUCMJYs+ulQsmN
tTl8oa7InILucAwRQqmjoy209H+U/EXOmA//IZPddpVJ07Z/+ShnpTn8F3TY/xFGjcHSowA5ZRN5
IS1d/+Oqa2l3ovhuatuzP9Aq2c4x9OgYuzTsOowN49epLf4B+WwUA3P1aQEnbJ3UGBun4M9hzVFj
Swmj5FGFBY+yp598aqedtki9eFsM2IsLXlgmvJlGwksdTZ/yhwtLkHuWnqjgUvW/gjWcysFhS1Qm
5yxoH+P+QYTuHUETi83Pi3i2QS4Xmh2Ccyk+4bertwV4MhkZPebXIdNeOMy5jE0xVq0cQcicrHVr
GzNTgLujcvF4MPypp4qJO26yebal90dSqAh0XYa6lhzAZhRfsMM21QoZoROSLGIasJwOUiCwC0j8
724td0zkj8hzZb2lYiHaJHGIKeYiSY1ST+9lYwMjV9X7dEo0fHXqoyAViMEmsckqtN9JgEJpY2SB
QKFYV20/dipS6v+u7i9ARKMH1rJ4TCniMzxwUZ313veITVN72XNnQKHHZbzjjQM85ZK2ypxqTJK3
VVLzmIWOQOWHP7FqzzH3wz6iYHdM3OByR1FOAWpzDLK4k1LZ7LDuJN4wQ7lavTC/IMi4W5kS4jcb
DAUeLwNMnOa9ZkJc60EGxTU3CXEZbzUovohiS4Wk2Km9R4OA+euSKVX40EoWbVJjqWVQGG8kREdr
xWb8/GMMWG1XdsLVd1wafrew/CBipRcwXoWgdUqE9QTr+tPjdeMuvkAKWe0jR/LKyMcJhFj+qutK
amJUz/nKzpkskMiz3owh++iDtDWQ0AoJJtve1TBFa8kWN8mYeOdCA2AgTugqqUzk5aeeefibntBd
fxByXnN7CP6KAsipijgy484x0nyq6pPadlhbq19bgFfifeEGzVwPDSu9ECHsyMbOKVOEVzLet3hv
gwFcrXv1VB2/EivoRZlZSE8Vh41eYiWTga63pv81J6VVQSyO0kWzfVdT1NirqnRAt0dspFZWTvZw
4smTqvVTP8XKeqVnct6NiPvANnePNRph8k0grNFxa+IL2AcL+ojdIbSDg+6XQlOus3jop+Z3uNNB
b/STnB52k89ggwRnTTvlZ6J4d3rtR7e7swEXr1hQPu6i0Q9u/l3CgY4xNPMkw76LsPP23QlEojkl
+HUMVN/8HlvEAxRGq3iOxRRuAvUMsupMJr42rYj19ZGoAYLu/G7vW9SPl3j+Vlh9SzmjJ8R9L8T9
IqWi9Ytxrftx2iJEDkSvQFAJmifVCqZ2ZclIMqvxmPrrPFT9Q0qSCRaXPfMEylPiAcuV9ygqgFIH
H+4Qcucco+uyU5682QrcUdr2aIRqyHiSNizO90q7CGl99WB4HJEkohAdLXnv3+Pe8VkgU13BAcJa
BTUKZu+RoPDCTyc9FM1StbQwPwmP2Q510lK8vYZ21DJGx8rxwumnYpLK7kep/Wz4+6E6s5SG1+Oi
F/N0gv+N/z/YyxCSPRrSD0UbxFdGQKi9JgWNZHS/AE1+hdMRDgnZXWY2/J24CY3swnIJeNeuNano
WiedYBdeusuMtHylK7OvRnnvQuy3Ue+Z7JeAQMMerrVj4GnkayYG0DR1SmPX7ix+0KPE9ya4RFV5
ScPYpWKRMMapIVICbJnZVHQSt/p2+7jyMpTXaah+b3BczelSsgP5ucrVtePQpvUOQwq2QcilIrC8
I02amEnSK6cHOJlZxMAyZRl9dFld5uePqYXyYOKD0f0NOlVRoJdPu7Jj2XTozaaSBt18+eBoRAk2
z/bWpl6gsBHxXm4Pdq2UzzqjAA+zQqXheEc+8J7mMLsk/W2j4oUnVLYmG93QbvCGW1NOF8kLAFjk
VNgFndQ+apD+5RcRsO2g6n7vblDwZi+YCqeCs+0F5AzbDiOQrfwXLxLH9LEbrUsPdYOX++cHGnMt
QHmkDDHq/9D2LBATHbR/U1CxEj6jVQN5N4S1Byq9shw3DLpbb+6nt6eYaYaTwBGkmTIpTmXjqEKg
vYeBtem7Fbgt9zvdFvUTlUS/f8VZ/ezXXMHNZYWQTD+CtNJK4V5fa+omByX3qReQvNRpReIPvojv
fIednBgBTlLK584I20t1OWWZ2K+tz/FpYacbBWUhzWaqq5DF5/vjWsSlJpn/5rwZGx8muiKJdxzY
Ri962pYYJAzlmYVcqfbWwVpiYK5qISssPTUBnVc1jmaV8cv8rsdggUh3m7SrxPCBxTgci6c2gc3f
RfWdQXyHsQRJm3120LPqLKl//f/dAEOu58tAO3HSHTZa1yn6Hv2XnkZlnupImlmQ+u6N9aKm8Yq8
SEmoRNE8Dh4oWPGyR9aVJrKeITsm/m3OEQhL6A7+Dg3kCKOWvRY07Yi/JpC2htoCH+ly4E2IW7Xk
27ZcNF2Btp1w/qynqVrwe00YLZkH5RiIqHyfKBsa+MqX11mxbfhpf/crAL5yoXCAisJuhKghBGbG
zruM22y4RAkSVbt4VOLXYicvA0b3abdcPWZai2Wr7oeF4YfAw6cIjVDzNYR8NR3ez5S0iaSycBOd
owqAOV8XFgJ4jMDbcUoLqul6lwmAs4sXH4Dw9iJ0+QZ7bytcw47lxyFG8gf6VTA0LGQQhzbuTnzB
A1lOdn88iOjZPTSX5RsSWx8S7xptH/BRxe4gQBgE994RnQGkSEIVhhJtbq3eKflIHh6glQ9EUkWY
iv5aoGXIt2HSTQHZ7p0W2jTUrAde/Wa5Xb7vYDrAA6EB/jckWYnbTMzaZooKfH0qqTjzMUQmLgIB
chm6Mudu38gQ9iCWI4kTMvbVWiwueuIC1CRNv6iTkL/0HIqMVXRH24Dhl3vrwuBViWrvIMR6lIm4
2IbmDUyJnYF4iUiUUocMUr1Zs5AJ9iIUXg+W4ZVGfYI5E7+F1qRtLPCpWLntX1sorUNV8mzyQqw8
6LhJdfxibccVG31imh9pZ7IkYsgY+fm75N7RKaWyYW2xAe1KnGW0CtA5g3dWo0xhXBkXAKSY5iOY
+Zmk4MnSNN+Vm9xWS4utc/HJNOLQVhvvz2yFb8ZqOOPi+k3IIVIbINA7GPudoGFXmiUxD1yv3dUg
YWeXIUPCP+CuvcQkHK/rTs+BTishJEBsRrl42yP2OrqII3O59kpOEucAv/cmi/brtZ0DX4/6qa67
R+4yY46+j4AQ6FsRZ5TJLdA0eUAzJGBF4IwBr+YO5FlKI/LH9xlWnFpkiwtdcGA9nzY0tVYgen8B
4whSrjkiqwWw/AkZ7iak5Cw+g79ui6DpLoxDXEOPaGPZFZwh/z6uF0pkpy1MS/PJ7garXpkT5bp9
gP6fUaJssPAzHO6Lm+po/pQuoxVWO5NnbN9QLpgZRDf0jaOhrDYaB/B7qiZdQTDSnR3NFuq5eV1T
u5uzignGE4d8+UcGEow7RDGMDlaZ3ltO3DClmtF65glau+o4h9XaA2m/h3Wtgp8ogcBjqb1a1OGk
De6C1Bq3VnixxDNmpNjnkmO0bRXuY57UMlW9FWuQz10vA6IUgOwn1yCprrNKSZlHnPKRNl5nEZ2B
5CLEJXXs0C0ROTnnjpLQcRWZ1VBhJGACzp6x67Q2FRj+1zwpCdvr40F4KJBA2P7SNhtxosGMzeFO
P8rnHQHIRd/hVBxF46T+FTOiUALK3mMNSJsJh8DCcGIt6tcQX0qzdK8xaoBKLGoS/5T3pAR1+DLP
AoRA2UyzewwUHPXDYnb0SYq6e9rEvkpPecahjtmWcMxIW7mC4EceN/aBjOJspXeU6aiZE9Q96wRy
RPDXcC9DqtYEXxApWSFBe4BzlNFSeYevfrC4eRvwQKz7nq2XhMOEP5dinCnUCYFZCL4rRJag0Cy/
oBy+amCMxLe+w/djTo/tJncNQAlFqAE1MFM4tVbNAUaZMRVY015z2IZOUi0MxqDm+Jn30XqOLK7W
5xpGjv0syYAuq/cWPoLL/5xo7wU3GPZz+Ay/in9xDfU/UG2W6fEfd3humTLAtVke+MwnGyOxbJQ8
WshSg+PHvIo1dv/Fa/v9fD0aWmvB5MTEJJvk0ScwflDeKuCi2d3t/V45iA19/nAz6sZ3RSJf3V0J
XNvD9x8dkbC7qC3NDqphbA7agsh5v/93tedi5t6uWymGqpAwND2HK9qzw6TJFKbWGjVxilycX1xZ
ZzjhYjaYs6ACFCz86nnamj8MubzBGlPsIKIvJvvnBKeyb7n4+faupcyvDzJUKdag7wvdEuypvXx2
YB8Rl7NzDCVgdu8+8pCp0geOQeCTfVqJ3708QCSx+FoYjhIJq9wooP334lG7RRHUCxrlNWccnZ+7
Kcnh5HvdGrXUyYFuos1HzPwUVlKY5SrhCJb0RNZj1TK9K677vH8c8TlpuAPTesUUsPE8rKM5GcKh
8OKrJttLLIHty6ry/rmZS02w7Zsb14djYPteBu07anu3zj2f3qhaTgYJ6pxI4KjaNL0u0/vCGgdg
QiAEHA2IVAvnihdtADDFy/sDW0pQNzxNiiPi7/vprcqXVTaGAZQrgDYgPTg/87IIKWpv6//o2+Ye
Kfb4dlr5JHQNjcHrD7cGg0gZFnHqHLYlBsF8dpjHy3MHoN2EeaaTFyTvTFNCS8RYAYGu1GOY3iNY
BaoGYIMxVYIFu2+fl1rZZlK2Qjnn5PWWlbhbqpgKlmEyS7cV0N8dMtJHoX3/aasllILEDrEoyf9k
X0gFFRzIbNexhqZhQLFsYTy8xhFAxIP8Ta3HbfIt4lPMDNNmxava7g0dDEDj1M6Pp7neZ+eVPaFY
Og6xJP7IkOfnyQ8mZ+7J9+A64E3GbGNnFtEDzix7HNTTY9kD2+uoDEBkotxkQEFhIXSBmKx9yAed
aq+kALXoYMl55wpN8CHG0Tkb92WMQgqh3UHogJLjGUZ7HNEx3JGwIUMCarsLY1FfVMEAZEBdnoOR
so6+bfkVDIWmzo5ap2sbdP31N71dMDSKxCPjDnpqBQ1s+/LJkYREFfxkZj4HuMg6sDU10YF/JdxN
LKL4xXCbfM7VDB2cqmNYzSbu2fDqUidi14UabhffXRr3Q7Wz7i6/6ySPXi2prpybmytpnlM4BhSK
O/yfpU3SnKmz6WpRHxy1wZ3zl/WnYy6ZFizDyhAmcFvI7gIZRJIDGfzQ1nwDG+xPzUq4U9fOGVMm
fFUsYLP4luxlqk3TglUWdGa8kzMBIysMTXUsna+MhHs6mVs2CHSEMcYwUUpb4kJ8NwkSI8fOX5CP
uKd2+Y+eMHVAvknCrKT4XKPlWWq5RFMM9+nzCZQUTRXLtTYZ0/k7wUfZXT+cctzCbyr6W9yShTnp
aOT/jG6RSNyoV8EjdsjSHT85KrJmueT7dWMnLC+FIBnr5Exnp1RAbRy4ZhgUTFBn1Oa6b0+QmUgf
3CEhjcMAfinSukTcgJFa7M7l1KJxXJikDpXVPvWve+3BtIIxMWPy90K3FPeDPCsrc9s3i8lCFcb/
pG15WT6e7N74pYwEe6s9XVqFqBak09IfrhPbZ3Nnrw5t9EIn33NtTWySSQyAkg3CHHXXkE+m/AeI
5FR9lLOPLW+2Op2Rdv4DdEUmD8O9vY+bGgk0x3OSvW6mO3TGass2Gxy8c40QUb/Y9HEtM/sCNLQB
i79U4PAx/8O/HuWZxcttHdt1Ul1NfaBwc0OqBttMqpr8hauosr94jf9wMhu6MxdRO2zbvmHvQDbd
vB0mkC1XtwNsFLyXj5/y6ZfNoDt3rHx/55ptSWXmDLZp8Wmr+qReBOazh6V1gNJNgxmnC+aOU4YG
EcAGR6m8+EjSlorZnlw8kOR4AUxJfwDxPe9Dk52b7taBgGtdiEwpONs/lzaSna9YSCzg604uQj/X
4N5RJU6X5I7ogwZ5TlZbbvDt+yeLt/4RYUPnYdVpxEusJvFMxGu03C8m5sX0I73ISxeGv+NefmPV
cR0pR4bXXzavBWGERKPQw8cYqzWvEPtm6TG1X+YQjVuMDvpMzM+vXSFJikJCo0/aaOEtd9zOdXRB
/2NYopLF+d8uWXkeVajDxpb0B+BUAoDg0jJ43mwygWF7nQkuxBVwX05auQEPkUjO5ek7aZhlzbIL
e7L5GVCU7GGP/r+ULk5KDPafZhkVxLORiRpaqFbbKWz4N6ODDK6EoLBsmSmmnRHzF9IaFwSq9DWp
5ltHQnft/fKT+e4VIXVae3QBHg5Iove0R47t92q630REt81Q3eoIaZhZ8SevHKZPJjrqAAy7uxQg
pWMas0BMpxt3pprRNDcteS+i3jWxcGeu+oLzWXJciwY++QAO2DnL/6Hg7wlWzH1sDfCLvOi7N/80
sx5spYrDJ+Pz/cEgmRfreLgpSPVSARxSAfsqzB2eKeRRpIzfCA0xzILhAcyvbaMGG5YPNPNzY4bZ
CaUnTWTX4FIe9n3O35BfSS6ML6PX3gKVFSylYxJsoaw86l9rpmqb6FChggT4GSvqdMLh2Ddu5Gyb
x7sZHce5/95aZhr+1MW/dHv1VJtQ0+wI6Yf9QW6a9uxJBKBnbUXVeX3b4ouqydz1fjBacl01PYGs
fUtp002Wf53OHoNzxeBmS3pcydIL49tO5gIHbwdHBrqtuzRJcz2jypv7pcC7cH6nRNqnQxAAuzll
ES0v00VhOwWDrurSi+GhYaa7yqZlRqj1w1A870/fr/nJqGX/7N/MThSo7HfGSEwQV+112TciwUBm
8GVcavrINjjggabQtknRJUHLqlHQh9YViWTQqa+ZpRitHkz6pgEq0i3w69Oq4tOz5Sp0DXA/P1gB
bceYbCT0FRddJTCc1kco9Cy/RwqCYt2FIDguf+xuKvj6zl5p6w0oHURFF2D30BmM6d3G9aUDdkD7
58YkLO6yQavS5/VtkEaDzj13FcwbEUhuOBnlk88CYlPtJJk3NXGtcw00PrTptBri3MJ8Z5EeegQr
3r/JKW+9qohX6RBAK7emOVYMaOLAUkhaDfxN65bukvN1LNRRuR689p0ZI8QiSZ7bgl+WInZjq5MK
Cl7dymelOG7a5TXvjjFVBOeEFaoSpiehj9AyucbCohfNZl/9vL6X7Iqq7syVNq6PsDxyUHW3ZExA
P6wr5SwTWMSATZ8ppNU2zxV27vdvwQ99KLVFpYNej4kF1QaI0/NgANyTPvYrZPBP8NXLbwlyacOS
4z/oXN4vY8DjxccmurJLLEPVPcsjmAAZR2ab6TQOU2XiGAZdC2fPF9VUVZH4vC3elzE/02CTz0sK
TnxIxJESnpNwn7Jybjy4Au/x8CojSsyxlFU5am8IV3sRLFXdU2zqMNfHeDa8VxkGPi7cqAulK1NY
rJIDwFxiyJXET7QZgCBv54LGPq1WGJlty9DcSH+nSCnHIzn4MUkPxYRxww03Rplz3TS2I92jcEKv
73AtamC+tm4jvpINZ/WDcohmu9IxZWSqoN2ZrPu2aAADZebOOt7fyqra4J2G1efN9EpmLAS3X+CW
pYFyn8XgnXMiimdIFj7TaNAZSVTws1MG7Xi/4Ec0iJVp+oQ9nhE6/0RRv9RPoZeYh6vSECwwUpWt
9f5j808XXzsPLgOdgne053AN/Jv0v7jc/SqjUt7lRP3z00/0rPo++9mWtH9uF/+XaDwUkEf0IWBX
B7R33dMeT03bbYlfIUvaAlSD9swDC89qK0McdbqBLSDafuxAnqizVcjyZbHv4FAoJFXp7HniKtol
fkv6NB30C5pLzqwwKhqTdOXjhP3mUvmm4oyPCs22QyBtoS4VuLexFVvDKfiuXS5uV/qbKwyyfqpr
lQfN2STfXUaaqdqt507Xyu01edXyyCXughQJIt7+UBy0DhUk/xojyaag4LQNoAJfy8EVsuxHZ7i9
SxpzkCbxUCnpPE78KOVf6YMKQf5PajClduGCp9IoPExeZ6BTw6SSh4WClakIl8z8RY3GHaSTuK2Y
qAD7IEn9dmsldOx6r9ffRAwmqpbWIs+dU6yNZfg1erk2XxKYBselawrrjK+NwqWmJH9Z7s3h/NwA
jNGdlx8pnQN3DhRoRRPE+mN2S3wT0T+pmNMsMKbhouG2IS02tRFa5aVe54JhIcfu2SYYli8HYXqK
cnc/hTGBxApRS1gU9NzCN2jx+Wfj2F0ZepYtCMCKi/KwQp0CZSnJtJz4BDlSUf0EOgCOFgYeDWtm
RfoEeGrDdK/OjdGstiWmw4Aw9xytVPj9KfecGSVI3osJugHJk5IBYtQvKSBqqI0pk4es61B2KTXo
8h4W7xsXXlYUbNZOH3GdEFEK7ydVAd9fMVYa9+LsNQwqT4WRnhmY06ZXoCoL/GWQSlnCjbCdRC5l
ODtAFb0GfuVUbtB7wMebNUyM/BGC7bMtTHlCQjcn1jskdUWe1wDosT3yl48c+FgEaJN3dhbrpiwS
VhFVkBkYZg2BKSrtLkO48g8N5U4a0lBK57hqzXHW7nQ6HTFeVFHppHeWmLKj0Y1UQHyuDy08P7R5
hZwsnN0LcyuOAwAlj1FAHiFuqisK6O17Y0xqRsSp6jWIWJVV44QN8u6ULgYY0UvVf3qsXPL0YUVu
p6YL+fdNZV6kae9P+FZgNwxOXKWBEosK9w3R61FxAIMMAEswFZjZ2OOyHXm3a1zVYwTO+qyt54Ve
0Rtzq7+a9R9CUQujO0+e8EfEvn3UcRIdlPpXGytjU+igs5w2IhmyACE/DZjXrbFcP0alVpDcVrfV
3M3UPFbobBAJZq16rm2zKeGFQnzuBp1u/see7vgQqMWvbVGwEKCwQPgu5l4u7uuQ7/NoSid9r7gS
1PpzCdZjWbENP/bRQs5e+SeOPTz77yngdQLczmUwcpYratoN8atlCunQanuPMsaEfQEI5wOYjNGf
8bXdFF+CE/cORO7RIl3P3s3EWEHLUJrLxCkm0hlYk6Iwn7x5x3sExLoqmb0ax6u9SascQxOf9NjO
T6H9ajUH+G9gd4W84+xv9IsoYqVx9w6oQ7VDwnhLn3izXce1NI/K7/dp36c8IVETino1ScF1PQXg
pUqBZoSXk/aoVgk1BT0EjwiRW0/tmuB+uJvu/cYvBbmoEiT1rRIv6plH7ZHL4ZgxQN5ZvhmzyIpD
j5ObQJldPn9aIZxSFncJwBnOdMPmFb9FWnCF3JKc1dafkSGktEymW5TQ2EnZDOKoVkdR/r+pcJL1
7Kra4vgxdNcwe7hpOlUsgWMuNlf04SdSeVmkvhUK6WmC409Df3ii4ZpORCRLW9doryW59TWcJMmx
ATbeY7TzJqowLWyYj9kPSwvkH2xKoQWjikmHIKD6NXSQwz4sOVpyDvhbzbQy+6wjNl+l8p747+LM
s2A1U6NU/eCS0wWKqCWZsPjCN4H63vAuIfFYGeEdrvZdZqyhJuQn5cGPHIOQnILf7pqbjgdeBC6x
p0SyeTfwiz91H5nnG+wrF7EdZxDgIejx3NZIeGEaPERdqKqq37ur0lTWLk9puVnBmC/0Q4Ejb0HR
PoyuIJp/NWeOQ3ALtr5bVCm/Ue+1d5w61wGb1YcQJHIL75R7Pp/wtnyEsqSUU1oPB5IDTRGfcPgY
q1by3ATNtrpO0vfqXbTlstW9nOUPItZV6wB+ZKEBztrsc8XszaqEnHequwPA7tjkShxRA+Y9a0Cn
toLHyl0kM5Cn5LYLWmTjPkW+diNMm3Pm/Q72HFoJvzDe0hU1TfFdCqW7/yRtmoIqQH4i3wO84bKz
oESo8/FVSAZchYW7DeAOkLt7fIqbbtA4PlLEuzu8RM/wx49HcuW4vQn0czGjleSkGfGflCZiGcRy
D7yPCBLjj4wlPj3rfiWxr4Wq+60BQl4Xyiv+1tiKSuVmgfSxuhvWztx0U64Qged6j1Z0rAIpJwSk
LbUpQoJgjPTVb7GXAh5aH+4AVZBELOQOS+MoGO3aKzpWBRE5q1eAtoQFnBUPzvmEklE+N/F3gUix
LcCFdeQNAbXPMrtUJYqOjFWbr/bUg5GnUIFMYhcfaKfDToODdWeBWwhVYbzZiUGLyZvA2FIhZh12
zbJGsWryU80WMQ278GzQfh3TWh59hvJ6cOreG1fwMPo8QvyuQdsdRHnt/Bp+mCRHVI6KtcbkA+LK
4jOQdbzwzq/UpQSfPxYn6Wet4G6P+dStZctTP36h6Zj27oytCmOYRwgcfQ4OXGMJ3pSn8tnUyVo2
v5f6GtgUno9dnYyvD5eRfVxajWMM0RRrA8Yw1qUjEeCTl+3O99qaEPYojjjFj7Lji7prNm6tiPYL
wNEqAMynLx1PACv7N9PJu+0HbhfWfouOOCG/nh3Dq0a8xhBNowJALqulnYTyVfOu5Fy/edA7mUr8
yw87vT9zBtl1jESqmMP8Qo26rpY2jdeVyXgHq9tp1g/E/54lW7luRRbCPPeqwCxAmCQn/xFiHRWu
EOyt/M82QvN2jgQOnP2LQw4RSyQ8OaHnwtYE/9VJukxeJuhHvG/alEBOMCAULIQjKYnHAB8rcT0U
ZeeHLDb6rRftQarbsqOf9PvFb+aWlKR28CcvcLFAO24x7QZ/tMaBvJEiqc9IjPwgOwRwawFuemDX
NJYJGk5nsOWOGPBZ7dcEW1rARVbqlQIRbI+0oTdyX/qraMYsf7sG04+/1s16kbtZ/EDCWRj5kSIO
qVzTes3hcyRAF6OXPYwOUzWo4BuweCrcr3VqwtC+0DxcqoTK3cR7sTfN76yjbQ0auBi7y8IxNcUe
mSfdwOT6vY1I2ihDAyQwlYGJRtWcBUJB5Q1kB7YOmtjm0ZaudShQlTKXTHrt71rHXeFBxx59kLxX
wK4K1z10gUmbKLgjVE+eXRZxRKKSGInKHu8h656hNiMkuDVDHfp/8raTnbO0sbrHMGn6TzHpU1b9
JaXsAkFDkae63jUyavM0eqkOkbn9bomjw2+TYogVAVYw5JZgdSbzSVYm94Qu7nB4R5nwRX1zuZ/W
YmxMvf2qTtDDxOBSwO92DboEjOy2TkwcdiyDA/0RYvXHa21eRrsB3qpzx7Eub52byMyFhYTl8hif
GXCuaGt/NGKiqTv9iw1G9Zw1lR4sYG2qbT4nW3nuMFL6c0UoESBrHfB9EZ/+m1GLMmP+KJSdszXo
cx7OE+z0LjmDqITPFpeFZEd/9Ap547tH/BRn+dH+GZ/O3JbsxitTT6J94VgGGSd2DCVuUhPnMU98
ceLu7CrBzNXPMEP/YgCye2saxcCUR7lNi0u6mkJlUvbmUlPqk3EluH3RgS7MM1rBSGq3UFUWB0Py
Eg9GNfKvci0+wX5fU4GCozp4sOQS/FClioFgjAEp7CIt+ZKaZU+rxFrCEpEUA6F/kw+Hp/AZUe9k
ZtQLamsj4Q+vfN3X32AwlHnndHg/Est57moo2cOXfaR+iT6tOerR7i9rKFcoll1CIyaADqXbDzBu
BVXC1bE2Iw77snzw9dNNodZeDQgIZlguHmWgdpwF8e+JI5tTH7sU1V0x52oYyBycQE1MnZC7/Qgi
g1u35imIheOq2TVeOAoWhdo7v3CK/X4xYZixsbB4rdcNv1jieaAMPVLMHCaBbyN/4OJLZ2utPDJC
UBYB7qbh0VL54244sqCCrGiEcWii0hjCNK6jnuI7OqpWfzDjKzdCvyKRJlc54QYPliEY4buM+d6r
7gvRYCF0WnAF0WYz2f3Q8Mf0b1Hhy3HcmKrhNKmyY4exVyi7sNelvgIso5Btf0ma98zHBwgeUzQz
upyzrDH3BsMvhQOxdfRL35ssDvFSGVtowjnQ6rlI3NUoTZjrGpXaDiFpIeFhudulF/+GePDYEH6m
IsFowPJByHFLNLkkwIEnFctuI+bUdHoHc7ndsaqu/7LgcNGQXY4bqEC8kf+OkPLlYMNjo9DVi1fV
RFmVJ50Gh/h1RIBRq1GtDzwrWRNvW1yB8a1iAU52nKyUSa9mWUTMEUg3ozmFcjDWG7BSfKnU9KNe
oJVIIM/NhmONohkC3yhkPsr50BBcmwdlZcKg3Ii9OjHKhA6D20GfAAGMKQjwzJLq69SFd1QiShKd
gbad1oc0k9QKu05y50SoS3OJ49Jqz4aPIM9/Tl5A5cc+YV84eFgpQP3MWkZEPgFcQbijwCUhQtNY
YrhwlN8NVVnOUi1rKsvcIsXXkFPGdGhx+7Nre4YDovk0fW3HT4aSfcktxBPEaP9Dmpg2Ljpe0NsL
10allRymNHZJrBciSvmjnoJdGf1xTJop7tYOaxSQdcoYUZfRluHFulRP90ewsosBB8/aT4ZvVShE
lP2O6U0I9oLFoNuUXu8saqHaqYfuOQ8BpYZFUL8ZiWSPfM5FO5nHqRdWfUBYNPo2SZw/7W2aTAm8
Ly40amwE2f+8C8RSvAKSMq+EXX3Aey3Wj87GymZ/3d8knAxqBcnN9TxruUG4X0KAHNEiMiMIQPju
hSJU8jiXyRZNUyAadoJcMEv28Rq6fDjOuowurt63hmPo4UsYI7MVpaBuUUmv0tFqBR4bzWyYnEWQ
EO0kkbSvi/1+5Cp25r8Aa2Wr0t5agG1chgq7AVAwcgaTD6lo8hm3A9kPu+56g3racI+UVy96Yl5Q
OblUAuBKr7D9V9OfDMDumMqv1rNRdweEFzE69pjXmH2uc8OwxkiOD6cfjDNmYFwvpNfOxI6zu8/S
7YkaUoW9dMyL8vt/UDdYFhlLMN012Teo+WO4nFd+MvglguoMcG6iqRSFHX4gRwJHc+bF1PjffHpS
y2cG1eA1Qxfrd4lnIJ4HNvU4lTAywDNo7nM2nxNNh8wEL3kabyEK3vqAJlpmGDXQNAWPRlI45/nC
6z7rcqJW6wjf4mWr6ZUow2TrpE8RFSTW7Wf0hb+4BykqwHIznkbXhRORFGhHLQf+KkQOKHN2VESb
kSmDFLDQLwqiM6rvnuUhqYOV1y/NMmFCqQL5ggMtCD7UnhrDVS43CSJ+MPyxL7nYvvZ7yzNziDRP
+0+nVSdXHAY6Vs5t5ipGx4e3DGX4KhZewOgiWHwSLwTAJUZuVZCejIQvtAuGbZPTkdxIYGMBxEK0
8UEKi04JSxQgja09tr7641rF9Q6j+2u/WoHI1OnHexdwu96wjGckc0hTx3WtYzxv3HEmKcPqubG3
di0Qf0+RDW22SyjMOJWOCefBh4JJoMOjtlpSMN2KLbmlVhBBlrzQfwvQbQJdkhz/fjWwzTIVQf3D
2toMOPXil2QmEtKroXWJO966BTK2MQ+jpeDpfV1AQbfB14Sx/KCu2UIRghHH4TIa71UeM0TrSltR
nnywnQlQrCzqll0+SQJcWtcuEIKdUrYa6Rd74bUHSYn7/aRi/c6dx+iQUMG9Xj82iZyUP8FQhlPc
NBG66gPkqCk4Lg4ABHkZyQ3O1b1D7rzBm5bQKJj6rymWjkR5Zrl3hVhuYilsCgb8gLdxnT393Kfo
K3R2SIsJFSvdSpvCQXdVLPTM1rOlyuqeaTdRnnMeNlJimAH7yAU4QHWZTUKnap2SdeK0kv10FGHG
a30G5HL/7Esj7IaflTKC5RSF6PpH803s7shN8tehhRrolVs09lEV8OUyRSMa6AToqbN5xC4pfMYl
LaPnIIyRM/BkJSnVNw0pWhGOpK0tuM1js92SNNmtQKxnNolSCpCNl6U/zIWHqgOyvyCBhhPw33nW
LtL96UWw/1vC1HJu0zVtK3A4vEFNahXU3Y9AnpvGQR278apDcGPvDmhnNP5V0Vdy8mexbOeyXoYt
i2U7RaK9TKsSgoi119a4MChdSA4PKNFXskPEiTLNwXPbZ1iqLsaz5yAsazATjrp5Uo6i7xVgtoXw
YWEkENhIMDbXuks2d+F0v3yOt4b9kpqplfg3VNzuoq4OpOQIf8UFsrMi9Vwvq8jx7TkQU9rSM8Wz
j8PNH+Y4c3b5LqQUi7TzS5ngD8RklSBZ8OSA3kWxo8tKe+usT/YGWOaFdR/6ojjRD/m3+vv9ar7G
ltlPa/WszvKlNu/NMbdYlxLJcBw5f8TEg2UlRyetsFhYDe9Ca+Hj2C2oZ6EZPafgdjzz9WTM2Ppd
A82RUqQPu7G2GYJSQutaUtT5l8Azjm9Z8YYK4nQuaHHnn5quH0EQf1e3DcUu9J9bj2s/CfTWeuH6
DPzxh/gjlRE4rTGNlCZ+yhATn4e0QQkASRnLTcqRCttg/v1MpCDv9C6T1ZRCNXXXdliAzjD8JALB
M4KXFksBoHkGZbkWMMbQ0+9wXGunzMmFg/5g7t/TUNlzfVyDg6tRY2UGLr6New1o8AFDAcv9cv36
rjFNrkX7ePBSbbEyvHhstopgNn/RWmJ+YyDrMLcUylGt12FrNJDh0Q39/mCypEzmVUEZhx9eb8jX
7gttBbKTmjTpgnh6Z8M1XdMdS8MMOjIxhHM1z0pHm99ScBBEPDXql2CUWCk23s8zS/OPqZK4CeZW
aGRR2gwibE6ZzPvHqmpLsrHPOa1oGR+/FG+Mot0XVaIjygaMZkunzhDGcqxlVLapoEU7icOMvG1m
Fs5RHdtWWTueuHIh0A8ROpCB/sJVU+ZD95Q4u2gjMiuYFZXiR0m/w/Ga4JsIuXW4KUmOmWVqYg5Y
nB/AzK67OvPzDp/JsJtOd2TFrrRwkyp666LMEYILXpaM85cfq2sOF+SjsBoHV/vMeSofiKqB6ghu
MM99YLm+dSezqqT7BQaZeKqperIQAVLfSGVCzls+fPdDyRK1dklTtsj8whxAb+7Y+c02QMSS/lm9
uk/2bkam9gKzCBf/JaaIJAoLa7rpX2ymXE+XsPcsZ/mfb5GBezmuNE2jCiSG5H8G+B5Ed/uhZIyY
r12lbinSmWP7/zj8KJY0JsJ/fl9asgKP8f+1Ky5k/mlTIwkFyonraoTCyHQyIQU5uQmPrci7BTQo
idgkP7uHNBjuYyaOm7dSKIc1skHJGCJrKA62hprNHrmFOA0PUva4DTQYDWORA1Yjjj8IGqQxX5BS
+G2BU5o+/hCqDiAtfxRFKDI+7zZTCqilSfG4Tr3PrTFO+sOmJurBGj2K+sxr+8lWvshdPffZXRq6
0YPr7KB0ENWpqXMxPbe87uZ37YJwGUrYqjfrr39eUNe6OmJxV+vWEwo7GaXwI8Yek5eGLshzy0h5
yctjJYvKVUVWjACGtuvcRYBde9SGdAPIiiYdcMjG2jkK66CW3Pal0IZKiW2qxmiDYh8SKLw5gl8g
YSpZ+evFVwKs+ScYTpESg3pUidLgjlF2MpYfna0T0g48bzu5vsHKuMhakNGGKoLFohJ2gPbvasVq
8/Vd1ZJQS7dxo/TEOe/I+M008MyoPpi86DnFv7EQQhPXYtydyCxjqN/Uc50Ac9myc4og3Bxo8YKP
+cQfUAeuGmnZ00rQZTNAzvfcQAmG1noZq0DTMiQ1nCMar1Yr03r+BOmLcJtqaf2EYCrESCXM6/2U
AviWkwvptpVw2a4dHagwIf+P0UqDf2FR0wQYG8tnchFUBBVGR1p2Vhq5ifiX3nKH1zYjr7qkq4sV
oe9D0x3R5O9mBUlRdO6uptsALUqfzZxoXejPRer5uoRliDnye1cvhRRYLfzdAETg3EIgKoE+CErr
En6GWpRYrGvrBF5LJ3gs4J6hOmhJOq3P+Mbam2JckyNVobDM1q0WBfVSK3s8dtS2ZjSBVg/V2iAM
062IayVxrLZPGKMSha8BrBDHhjpBlT1pgZiuCksx2DZ3F12H+E+fVbvCm0T33+bDZdPUGEnA/iKd
sb4d1U42bkqpE75gwpeS47q45bplNLQG6/qUk/7nGRshLKSBBTq0zo/gKd6xl3DxauZvEsbdEHMs
8oml3omje7dKj8WGFQqjdC5zjWxrFnOgCZQefKmnPeEDQtEGkD4VD4eyzYeH/U49vPcHd6k0nDE7
hOxGoX/H2wjWyCdT70vbYDS1rMmBbo3ezJh9c1wIuzXsS+2jM71XPZI4kEpxw0cJpC8JN4qEZ4xC
MKhUAwa3P824Vg5WRKOj7adLvrQua0utodQ55RQa50M1NE/r2kabit80rP5d/L4Bcp6bQZQjigEt
o4Dzpb4+anvrMCUpdQ85V1BvKXsYPBepRoDRZaYxaTUG+AOoz+P8Rmn7ZxeFJm9uppTg1ao9w9RQ
Y7fWMNvt6aULgrPYvmmZH7PT6fXv7gEVAN5HOiokeXzwfHs4AMGYzJOvMusKfpfR2DlMub62h6fV
wkWAdo6SIOnVbPPAVNxlaUFHMsHGKIWn0TLZlIU3K0U6PG4QVdR3yb7Lzml2HZ4ew5cGZTuEdvCK
J1283XW6RwBttwk4uKaXTegO87HT0vMBtYLTAfj5WPBto5yImai4tv5ruwjC0n+8OsAQupR30hAF
N3kcFT96uxZgVhfZ2zcqx16y09VfnOnr0wTFZBo2bf82fSXtX/w99SVHdjTxVapAWYGhZ/6tod9R
gvkc1pGLkt6xOdYE5O16iSsdLHWKOcAyRs0+1IIxlNmC9+Hx1eRC2VQyZ0e/yfhoev3HrVDGZl4H
aQxCI1J+WEZ7uMKN/RYyPQj1tMggLHuvRkoXkkwM/YJSqFQ2LdlRU7qbHphIBLcqwBP/WUurIX6O
lKzpeo/bu0duzWAFVeoI7FLbsG46H1GvBP4iSYvtq2nhakn7ksuBuIdu6HO121ngT8lfnCEm0rSl
l2pkBJMbF8cH4zmDR18PgTz8dqfguFpY16BOaUwlFMpPO9xcbQrkKzJRnIeWxD7ViGwN48/X/pKJ
2/NfKHks6GHvv38s3b2RbSmCsiWWQYwH2mNUfkEinPqw/oGM2IKtJb2oBYFnvTgcl5TpXs6jXhz9
yi4GcI23EFJirMjp4kDlcdBkiaDf3UlitpMc7YQZZ3FeN8+T3/fMQ7sdo5++6+Z60LcY+vFeVuAD
TsCoEbY7uuixTrROkIGfPG+Kj+9DIOZ2NwJsw46hw7aoIoCycfWJqRc2GYCkx317NGWXEeLm6QAq
14zq3XxHpdIr59Y8a6kdtxHMwui6WpdAxrv/ML0TKvyhqSBFa/eVytcegpv1itPXjbOlKfrCdds8
Cmn4WwFPu5idprmrCCQBzPJxwev0HUV0VIg768TfvyuTdijuLUz1Sg5eSdUH3X2MBbyS47ik88Sx
ozaQhSPSjWQAQKlmnG/rev3EQ4fRFnEb/TnIGkTTqJysF+mlD1ywCHIySVihoAVHYQ47BpF7ECpR
egmq4+xEwuMEZm6w3Li8qfPja0gA8cli5bS6ZGTL1Qs4Eq9/4lvlXCdfRFm9bZFyCIaf2u/kYi3M
H+dVAhbtVlSDJJdv/UlqwDI8j8NyqleaIqBmneu0nHTkqC1d+ORQ1ONMABbBDcM/oIsavPiynq9J
mEa/lHfwggMts6bHxEr3GlKjqAIOZAaKVcAispIsoOgr3YK9rjs54qSJ1El0yeqvfp0q0ltSH+Ex
cLtHSJcKHch3LOEi70tKy54mKF1G6cT+bmo/2hspPJk6Bx5CKmS3F9zD5WY8CZ001zQxBmXjbi5o
e8b6XgM436heNc/p3teK1CxB3Y+LwF+JQOu8a/c/lWhZealotjkZRZauv++KQpsUaJZFkM0z1mMn
W3D42Sl5w8Bu65Y7btApvjcEpJtFSmLkjaJxrpAvSSJN61xXXvKUwWStvLGnC8CZunoWnDM8BGvg
kQgyYblzXrrfcaYCrRqRM4cO66l0bczwOI3O+yWNc+R039nU1+vrN05XXHSVb68xgqTNyNG5Xg02
st+94KtIYkLlIH1cTLj8JJfxwcXwNunGy8pX0ryeBZqSEbdopgL3cILB8s/VcP55CgL4/+Q4BZDM
3AqMmUE2sGEX3s8zYq2M0hZBVQsU+EL571WzKVA1c3DldkUyz9QZOo6hJSFSJhfQkoEPxZTtkinq
hnW+SO7RN/s4J+0fXvAX8sYypjoVXHmmKQ9pUo+VcW2bMmtHYjEc0gdWXLfjzBjosGjrSTV1yR7y
rH5nd+eF+2XaMRUKbpv2qMErPWEcwqIjVSCpicXfPcrs0We6SAzS0f5tp6lJNfyfPgFMXKkH7Aqf
a5d7z6HTox8jQotWmeEiY1wKFAvDVKBKCqTo/RTMMju7lkB6HGjBfxKI/ohHoIJ1xqJ9S/aX1q7V
kV6BgortLJhACRWBY8piSdkpxHa9FjIV6BYeYGJKvh0bFCVk7CawP1suwmGnj7sTph/XIAQfY+U3
Az90wRkzrBl2ya4FjecXBZeqlbxunuNfnN++5qRQLiC+YmI4MIBQuTnavlaTYuDeD8v8ZabynahP
j1Ul66yY7LOVARWnm8+JuxLvfnlVD9VTnQyn7CqZeRyYEWm1OAzk9n+ia1GlxjS7ystrklBOknys
BmxXBg9EbNp+ejmGYziYq6Dfhn5t1NqY5akvs4vhjAXZ8+iLqHgTEU3r33sOsnOAscwAAcCN2Rt/
Naj+m/blvzD2ohIxhSXf15pMwAOvFz9AZ2p4gN11/V/VESrzFYeVt5mMfWqhN5gI2rSYBMTiCtib
r6iRATAe92Y8Wy8V3N5pOpW3J8Q3gLVXfKpWizKDjCkhR2WUonDehuyBpoG0QkFnaSxawpGt5BR+
WkyuSUi77ayaN24QoovCC8ciOUc/HBBbrIKxttmuU5mW3NKxjQOXsowYiPbPrbX58M/e1r0psHQb
kORS7Mw2moWvea9pOyiPaEwnIqI469843Rv3fV/roVG7z2aewxGx+PGx62g716aIhjugtfQuLY4h
fH+Z3Rogze+uSYvCy6VTNqchwWWkG9aWOaFeqj49vY9gQOqSCvCUoOkGdt/PD49J1m19vnxTTLqe
X5U+4y+FstIXXw6HKMTRBWfmoYZOr463DGN5FaJ94kSSnJmVotAvXn6USHFhn3TPBgr2yPP+yq7u
LMdI6j178v2BFtIXujRYxoSeS7IeCPadbuZDdu6pVqM6VDoseVslND5O2YrHMM9UJLKMMlyay856
VON7xlB3c5zYtOJWF5djQtsYg4lHSFeOPleoM7TvFxc82IY1bn1nhdUkycwpN60GnSWiB6aoaorc
JX9Fpx9f/ggiDUq1dwFrbsfSLKl1BfEjwPcOctLAkQuBb7JkJ6NRlqmhdZUJ4jDTV5KcJXjJrDyl
TnZ4E45ZX+DqVU3igWYaVqhERMRXWSYg5Slm4JaTaU+vEasbgjpyTvxFMZRpyGZbpoT+uIYKpdHe
eGYgRXrayFIAKzz3fo46BPLVJptwLCmvZBHhq1uJIKVNLaVSSFEhbcgz4HQdalThA9SPJqPApqB0
nM21IuaO5jydDdr+Jc360MYx6HRJjBiGNtAyLMNKPwVyiU4tH7KWG/oB5h+GybRFJJuTTNbcTPXk
z88bUFRL5buSaMURyaWugHFc+aGFVBoCeAfP/Tu0sMZbtlQ5X/eZkJlSxhhYWB7MshEp852ukhwA
4QujomkgmXRCfKOM59sFUEDOYDxOI7KV1aXIQHdviyBf6ZRykqSG5k0XzlF/eaYjnoVGsn2EXCH3
O9DBvvuQqPa6GnZt8dEbuEqDMGtmTb+qHjuo/piHEoOlkQjyPibjOEC2RmzTXRGBLMW1vEUhBmwj
TjwECx6VyjcHwjlEzOPQdsKL0l1aXm86JaE6MSEf8tfbRHncXx8bcgJGKNcB/wFC4Vtw3iVq5eRA
WEEy6FrlCRf1hCLtf5VhsAIWlpDTmlm/5qcvrnFaytpoiWSCGDHWmOKK/bDhGCkwMmkILf0wo45R
Uwdyn4r82DoFRxWAGBIR0Js6bQltQSbkP26f4EIbY8aYrZMqxWfgyI7X0C+vH2qGTi6HZPbegGsO
ttrnPRKhqQUHR5jC27bhPpRlGTUdFPpxM7Nc3nuTo3tRPiN3ym3OFnxg56TMwDcZNhuIny6Gk3pq
6e0xYweSp5bPNuv8fnhmP1VVFktEXcws0U3huOhSBmEfhJ3Id3Zr4lOYrSbTa+rlEOWDWezrY7I0
GpMMQAjOUY06BEhBOZK1KEcpmHLjrJxAr09s0o7/JT6/EdGDftswg6KtSQfq5u9nz44mS0KdUDnw
nlXdOHepK34yjMsmupFvxNC1ZqMbzej96SzfWjTX8b9136E/3wG1DQD27h3TmyEkwS/lRpEId4sv
0SP6EJd0ZdWqCMT1zk4IqXe/Q7Mfu2L4eOBIfbaOgU62wNhQQM6e2yTHNx0fF9SVUhU237j+fOrQ
5EkPSd/c+oHLgC7xD5lFyhuzjDhCxK3RY6j95D3wGIQOjKZDc+B1xrdQXPPl0TH4EPNs6n6SOkeJ
Dh1Xx3lD0PjZml1005v+1rM5SO3raMQ64BS8IOmS7Z4RGYqVGakDxMuqAOPpIhl13o2AvbVN8r7R
SkBy5FpQ6uHElP2i+8MIjnFP9OWRbt0rHdPGj+cKR+aD8Xjop4KkRpDmJzXSvNhZcJW1FYrip2/j
vAAP/fZZbRFEvO1DpmD7TDck5+wRQPwxtP6D4eg/6zOXGz8MPznaTIpMbzho9y/5fqLZqUhfPb8U
0tTRL4i/TF5a+jZCpn/VUErizRM1/7bdSIEtx6oicnzcsJS8iFLbw9YyRjLFl/OydGeDVMiOSAZ+
1EtcR5Sg3jZoClSJ9uxSSd1YYVJDm5e3gk5AJItEHoN2HLTWbPGRHdvfAj/kE6Bt69u4jYPH23sB
/Sa0ld9+p/OXT+8XDEsg7nXpcVjNsyj4m/OnNwkxFW1qi6aKPohPVbqUzRaRHzb1Ybq4iokz+DJP
Uqm66i9hUduybTE9CjKRO6Rbw5JY5AzfoatBMJ9+xMZXil4IIcMNvYNaqPSRb8BRgVhM+GOZ48LU
xq8RVESShPUd+CBASXc3yEL2ghLFr3VBYDu14CKbasU3o2h9lqgSjaUdttidR1AClA92vGODG/YO
/mDct2eOZO7qI9+QXGOpyUWbSPfNcMJFk91WSEb7OGeafseClpMfOktra+k+UkqZsg5RSxIU9IuX
d4YT/i42mjYuBvBfRtABEMJv0jVgcswL/DSV77uWWnW/Wy599vzAtpzE0iLIAdtN3Tg5suzdBCnQ
DPTGeVzR6kmzFz6Rn6GFcpHlI6Axxiusomf/YCiAsPm+dBBcYLwWhd8q+6NDpssywACmMijjDKhq
M/0ouceqkawBGPYKKbb2JwL7JY3OJKG4561HJOESJOuk77nYG0rU4Y9jr2ARqNhyyaj8pbttZOTH
BSfvit0vE/gthDRn6i/Lpuxt2QBlWiezqWXVSKMEsHpyypIBGTRrxRCN6jxkR2owz8skjDKVdaTE
uYRCraScgCxSp//ks0p93KJ2iRDel25shXowfdm1KJnVuKgmKx3CxEwW02veCaqkntLjtYXUPcxb
x9eCEhmHY2OixUotolqOxyUpZHevoDrnvnZLOSQSyZG6FcjSuVRmPoLkWSLPKS68aL660vluN9DO
E2f4DZ0gaT0GdYu331wwD0sML5P0biDA96gSP39b1XSAmVKrFI70xn0aXo/Qx/91OeXo7Er6jBl5
dF7NarowYNhhhfQyxXLX5n2AZpgf3nb3mz/kVmgHDPLrdUvpMHkIRseJGGNTu8OmN62Tt0igf2cR
JgCewPano6OSzKWupuj9mEeU9H2PmB0DTL7Ez3jAzRa3S5REhOELYcbsWpXW2Fx/f4MXS8iR+5gK
90S21yW9LMdALWP1slG3tVeToDnZXXtxXkHD4Wmwr8sUXR/w3++cHIpIOoMScxpS1XP35DLkAbdd
5AmHD0ZfwZpIqYLlNZ5o9BUsCEG/sePh/0qp19A/yIUkChg812erPPzMbtcNCyBkd3wKDk2CSETU
9lTS1PozsdnZ/WMv8/XNr4wuGgFNFvirWQwUrALAjgJud8oyvR5BZemhrSw8O+elVuN0uXE0ssHk
o8dy5pa8uwVuhHtVRXeDFE9yCqAUkhUgPnCZeSewEWJY1qRdrGG0xA7VE4qvWu4FvHJQvI5ebgb9
nFWim2S1+NUtxDRiktFNklIqQjjDPu7rejXgW3YxLbuZyXGYwICe7xp6DZzT9VozjRxGpXUBXPWZ
ydKp2KmkMbv79fUb8E4oT/JxObb06v6IRMAahT7x2UK7IMhHFldwQYYcvV5lnNo3XpAwaXQhoJkT
sLtYikIQTuVPVNXpUKBwqSDfSkvZjYpoUZwavMwXVR2uR3uzUxardJfhBkxEcfSvEQkBDFEwtQUa
/pjrNZAOO/LqiCpD4nd+JBLo0a2tYcojeHHH6CruycziPyfRfSIyR/1N5CKp0R5UfZK1G1nKQ0MS
0vEkeFGPzRiEjG8gbdz9SPxuGEDkKDnjJt+uL1PkonLmVREJbW4CyOi0vH2BlIH+TlHL4rKyYis4
guF0GXcfAFMHSMj9gmwd5QwcSbEQb2j1KqTMouQkvR8/1i+/n2WgJ4AbO+r62ZYhUp83rKqZO1Mu
36zMZZObaToImv3ic1/SRD6cysEGOc/mtYSbvPJqjuXoneDybaiXgYcNXzqtjwZV9dbVfmJHL4+l
MrYYwXd1pP8lz0mKRMTm3LjrN/fXLAhQSwhV9hNJGDKkI4qvd70HTr7Mfp7AyOybBdf1o9fevptN
4h18BXSONTbPqX3Ifq0Js00anHst8hSbVp3S9RjJ8AjsFdGnUg35/VtvzU1Qu5scJxUgIW76WNMG
3BY6DvUkka72/DtKH0h5u/dKS+uXlU97RNVa2SPEq7Cj5IFZrTJF35QVEYRE7StatA7y0NPQdDqn
9KIHu6PpQtLWmYzFv6O6XNNoT6KJz5eEFy5MvWNXWPAzFaioL0bHBSVNFgBThuFShlp7+NnKY15B
+wLH5AWPdUpmhRkYxBBzvff2xUhoQIdEB7/1tyyvt08kaZ8RAmfrOPGLQRTn5dBhFzY5dKTPm3LD
5V8R92JKY40UlsIUSzzQZpm/vOi7WDQfKalA4rgtGHld81xfuOzbrpOJPTJ+LB3p12EsV/Dj4W8J
IANhZ5I+3LpV95f6H+pjc2faP4lpILvlyudy4w78fx+pr0P6w2fdraV5RT6Px+TRxxBCRk+d+DCw
Q80gnohXGO5WZBQQCL2YEEDqDVXEK/3z8L1fKMOyWbulQURKcAhcvHzMZitX3udXXw0W9dhanLAq
5rPYMgnYIc2YhlQdkXb9JP/37KjnI3cEEkO8JM6YDoY3x0ZZH39Hq2SMbRf2cbQm/aI2xIya/SJF
BpoD7F1kE3XTkOuh7+x4QEOXxdTzqteDnA0bBAQA0WooMDcmSXBdafXPYDtiVQS+8edHr1LGuocQ
OZpHF3eqnQEj3BOyGnKaOIpzwntPNd+axoYXemXHGcpvAdo5OokHbP8SiKzJXxQMckaP7/afwV/O
IiHbEw1LhflR/zM0MOQJZ3CzA5ghtw5HOjmkLeWX4siNLfnj/HbIUkFG6VaPgTuoICyI9sNAYMmC
2xlX/2SLLmFTwrZTu09MntY+dvh+A4whjJk60fcNuE/7Nh7YG2Ob9buYnHMwivvgy7nIjeLRU+cz
bMhLaAjbhhrmT+7iDPj9DLpQk0+B3KGMrb+TooKaAjATfQOp4Okbv/3X2snJ3VyIuuAFYLCxUOuv
hLOZZprAAToc6+NGaWWNEm46l3G+/7Tz6hpgi8DyVkXYymTJiYnYK6z1i4HJObqK6oC7sFubKZlM
L9aJCXOMPuL2I014C5Z3Q2gEHSLcC0PulVxJ3zE3LtSu9Ul9LBVXvk+p+pSRgdm422uItM1mN+yZ
jCR75c+QHz4Ak3gxcE37/pgBk9bg6wITc6irPUS+4PdssYx+KVBFC6VDoMdLucczro1bm2IxCl0G
r4dPaDcZkuLNia7zfQszz1938Bt9ojQJpCd2kvQiOwSWGlf8GinKnfG0CsJxpzhBeBXY8bZ4PJBo
EKX7cyjwemcyzWmboVpTBBydecpeDRvvPkvbslDd5ehgemT9Nm7WfnZr5z8IFGQHc/J6byIGc/A4
1H1mrp9gAUkoWhprifc0fCKhd2hjU7SNDIGV+AAbV5xVeZDX+DyMTRkJE8zib+4FhuaMZU9utDyE
/OzgeNRQgX8IC5abNym5NQ3CP9LYZlWV9zyDFMNeHfhzINOjqH2uvBOYiBUrIhFxuMrG3Fkn2HJ5
s8S6RWSl1vlr4bUMkweLDuLG00N1qyJK10ZO17ioMfmbLQ/h6RjhPLT3Wb2p4STcrzVwJ42m6reM
HdpOSz8ELSFxx7PNnb0o7COc4Lf8aDcJsd0FD/lt0Ax9vm++waf6ubYgOg3GAzhKE/PK/b8ZTSoK
J0FEy1w9NiVrCFjT6rlmNNCHkrwvUsuWy4/QnTdFkBZk5hky9Jn5nhFN3UbONbRiN6dNbvgQ/yz9
XN+SNOOw8sQoJV0/btSlxeb3FDZhvvsmkyzv0BOQERNwK5xDFIemq14uj9ejS79nESTZrNJO1w89
N98/NTFXWRvdW+5FTPJRoVSVY1rfpaCx0mynYna0ZG3Y7w5xmiyAQ5b7mcgMhKP3IfyxkJ6mWz7f
I4iFFOEfBr8HXdpltxN8IXw8gyQmvXw9dxOqbWFGmdMst0hpOc9rmWxPTVcbKfNcOkWD8mG6D1Xk
iJO+AfYDf3ZyqjxYuXBR0GQTlkOeYSG2GeEvUZSocF/aRY355x4Gb8mqtXlS2eiugLODvN3gHW4K
u+B1INcul5x5FM9s/botGPvz27pz0DZ8T3fFd+SgtIE9zTDzCeZu9LZHC4rzpzixl3yqYlQYlrSM
gRqbdt8O9ugxKJfzJAA24IV564QOr4XHNdq+HD4YLZBgDaFp75lFxmZRAnP6uVUTe/rOp6vPpSY2
v9UpyiG7wQUTwRyn4CYbmZ/wivML7TeUBR2GaJh6YQudtGQF3ag7wATy7YFTwil5jNMjMUMpVm2X
9wUa6bsp0K96gRYvh7v0lQG6gXvM5xJZ+QRoy3/Q/MQdIL7lJP06AV9tuPatqtmhSvv5xu0z9n1V
RThArQjRW7ScZejI2EReQtYZjcuuEvK86J7u7iD9GZZHiqxEldjH2wkEysZlwMavX4aD/Xt5tnf9
7AsTZTXG896yxrcaisaDmPt4hLEAusOvKpeJkzrsMWT0BcW9zygI+OIImJYF8UtLtX0VPbdWxDy9
CXfPaQcTXnFjfpHkZOHVLuMPFj2R2ueJgw6T1He7FAYiysBu9970QI9xvAOgpQCkUfJNp/K0RTrS
JcL5IKyeesnMz5zxrzTcWRSR5GVBFLcfvGeUfAA5cufJshU7Cbjq3TI+lsbTlUW7WSj7BJj8SCqK
EF78sm4+GMKNvwsS7R1Y8HctH6vmiRKfytBf4udpZvw7fiadbsSTh4wyvtS0uA1RmKOqFE7cQmJW
fsfRi2Fu1WKb7XIOtf0AGZlwlHAKH8eXNjCOKqrGTsE/L7EgXOGvVqddoPUsQIBKwtnswHdOqgqI
H3IK/vGN+FBH8PZoqrs4boJB0UPObI21N3HDgAi1sxhzLbjVAfyVkA9ho2KLCbpBhHhVUeIMtiUI
Y8Yf2JPhw0War+ufPQI538ku+ZDvASZ37bKqUWTqmsCf9Kl7dWlPz2+nw7m+RTYnRubKyM5mccrD
Z7+LdvBVTjJuvrM5t9U5F1zNhlN5Px+H8imnzT8wFD9FBAvwL6gPaODUOhRyDkHYL1NCvjfgGTtk
Xw2wlIwk8y28nDjiJ4jd1UK889xohM6GVcRVlUGN5/KOOAzLvr1dloBrQek16HD1QhtSWSmxJfxV
/2R05ROPFIexVTSllghqCq1TRoeO96Hit5Awj/cLTwzX1o64ZRY7EhYcBZ6B3+ToTc+9+arFejr8
hGobiSgKe0KeU3E8om7iXfmjI7uPXwXhv8aruvIjlcVbwEByPr8hq3RJAXEN81T7jWvIFr66Jsxg
HocnPG4dH0p8ddBXtIEY+JdNoYichApo2sv7BMEOzAtzrJGto99J/SaCKNtWZ8M+e7ZjLU8kkW3t
vxleNmpDm+U5IC44t7+VaZiW2m2JufsclMcNsDRYtzm6DPryxWPhGjvg37foeFHD1o/AYd+yHyfA
H9ME2CfkibqpVB9OJBKh03PE88RNdLNFMk2aZMdUIECbfC9zLR0AdA1aHueLHNUw0j26zMJC6v7C
+M+TxCYuOVYotA4Qhnew98AxB0nRObt+jLJL/JN3sq4YijYeqQL93xcdgZE+UcUphwGAUwk8tZbf
SeRYLsMRvUzqXQEFTHs8ERoKpqlb9C9nXUtk0RqICCioJm7K3Im35m4Z1llfaDEJ+S84gM1WVZUp
MZzMyQTC1+94Fjji6sZXmux4YT7yuy3cJHtKMGMIHgFH5CDOQ5bEjSLbI0PeuxuMlD/5adNYsSn/
fwlWoBXIPKI52vZQAmAi7ngagrGSsotZIfbsX3m1JJrWuLcgiYfQeUkrE8q/AEogVdpzhz7EJDRw
w961UnyZzOtlDQBRIBAIgU/ggDkzO+/FeV5glGgyMnl+ffs3FeKQLyyi6NbvUTHwuab+X6Kx634s
wjbnMK6fkw+X5NvSRBgSFW+/VbC3ltpd1a1oODgDA9TuZNoBfHCOFMwHmAeVIRZFGPOwzKASM7QO
LSemnjCggHijM90akUlnRJ09nnui+8NCbgkwhFdw86kNl7oyeDXpjEisR06ELudMOqMzLV7bq/Ph
oybzIxN/hpcurwFroXzvAm/9RWbcUZTbXt0g5wMURxkAwUbvHrVddkKQcwVCO5AX2HyjjWZgQQBg
JDloIc+4kL/3+TOdrOp50sMQR1wR8ynnSjoMhe+vO+P7dYJWk1EiVg8I+vuN30DODHb4etULE4hK
+XQNtBIEZiQb6Mz/iWs1Fz90LK6HBfyBZxmcCdzVKMQBvd1yKRz/O9WB3ES4hf7OKIXCglsy8XRf
g5h6001HnJ9LlnZNo9pqGYbNXVZ+kFhRQf9mSM09PQ59IVtxrVaNq9sBKbpgQdP5lMZP3YtOIzBS
RwU9+loAUXWJVa4O6fcuJHg4q/gNjSCXRGmJyskAGCJ0YemGgWGzNdobkL37CDSeHmf1plGJGjpC
5NtcBh71wLG3IWjxECb2zdRKMKvwl39Ynt7AKIipC+hCUidk6iirwsEjQk/gRulSgeOKBI+vrEMt
KTon/xOGX5+oarkhJ08rFggZbuoyQTf4t9WJtEkVFxVG442hJpnhOS1bmK5uNI1DZBOGr/4DEOFV
aWLKCjXmecAKJah5upsXgxYAcNCRC1ZgNg9FZ7pomCqzUfvrY0BX6kpGOCcecxRjvSTVcbW88DOh
ZG4EqjZtmT/9seod/sewW5EkF1OKbyNl+9gbw9HATLyKFgnNZWbJ6ihQmCxTr95CWqGQ4HyPNlvw
GBsXaTh9TZ+tzYgzAjQdnDKdOI1rvgQX1NbrqY90DwwzwGPKzPE8B6O5fooaPju0xX6Nrx+lLtki
UDcx9uLYDsx3H425IA0qtUQxEkGluf2ILTo1mCZRxbV0QvHV+NSYGbkt84v9yj15gJ3aNEt153dn
Yv7eG2moaG2sOXMzrq1chY/3o1l+7PE3peJe4RBKUCDULD/BYvPQhyKj49FQFTnm7FYhqgqiLBhk
/dARnkzvCcqJgx0nyYi81qt6sAZu1NjzANBYg1X3w7HMHKlpHjCmQzTfKv1cBraNybIJtbUGIA7R
18CyW22NUSZNcJ4st9nMWrNm+Bbr1U77F7uHPrQaRAEHCBjZcR3JEr81xGsgkg2vbhjJOdUUdUyF
Sc7yppLkel7+3IonLWS0l/UAAzEXdkLpn7nIiJUt6Mc1bKi2qYAdJU/prJy++DQfJeQV3quUsuse
Zwp705WqC4chQc0CeRMpLSeJrMjNB6dli1I7ONnYFdBcMLUbEgUuFyXuaZ32XA0roNEreOhBXI+D
mWA4BLrv8FmL13bq/ZxugiCgHNYRBF6Pk23V8lFHBb42qYHErqGNvUaXKqe9SxJ5OsM0NrEmEih9
zkrw+myM5OAL66xJu7lUK3b62ZAk4lPQFkDCCQ00SuBf7BODdi3P+u5rdbHspo1vIIxKANqvh/1Z
dauETJoJlp9AjfqqkCc95bpwraG/BTFVYzQ4JauorQCQyHBBiAhF8xFcz05ew8oj8CyHPCG14iWt
aBfIMxDHUxnPFFkwhNwsjZM9NFZmiaA+UshxN7k79BZ2ws4J/VdEpNweGHPXP0U0Shm6OAvqszcI
avgEqJ/mZYgGCMcLwtfFASIQdcc9P94Bu6+oOhMs7ZUzFAdCYCYBb1VUOF8VFCrV5DgI0ayPQG8C
w5uWEXjGIqyAjr6nbq7ZLyWPbYbYkGaGzNpsKdGeCUkFF8MGpMw+jbrwM0UaLKGepnIqPe3Aa43v
KVmjSqlAqZxYLyaVZQcgykqHmW63JcUpaCBsaYNL4oUKixLxSbM3sCr8PUnotIF4Z/70HriDLZ9t
PyKFzbehoS/lykAHhUvjPpn5Fpnpytw2ngoyIndLNQ0+Ds8Lh8K6vjIR6oeGp+b5in7TiY3jH9ke
GQGFWdgPOffBWE1sgK/S1C1x+mx7axzeyfpRbTJb+7lC08uHIg6z1vQ1TXEE9Bbh6OtZ6cV4rPOS
1GTfDuiMqGk1DTGWuGmV8x1xTBCLio4CeOqHtQHq88+jPsoEr7gGc92mhmB8yGG3zzABIf2AA6BJ
6o3FsBfRsIc1kJ+kilNKhdBiisZgVuY5rYXllJ8Ix92QwMet4TuR8v61mQm2JJQqAc9e38nDuVBJ
oYm/C+Q4OJzF9HHKOa2PjUMoFngoPiqNVYiqRDWx+I13zrZuuKruEdYTC6tFyQRzVczPSE9ctISp
X5vtq50aDEU4aELP955nXgpMFZrJcLD23mrCtartd/0EStRS2gNx9e/CKJ4v/P0HJa3xUCjFAtqb
91S6wdZDVOhhq3bW5ciVWnSLoAuHU1c8erF2ghj8OEu4DWbCcYepoVndtIM8n5t+rfpZ2cpSEf65
FMzSZyT50iN4Diga/5BE1uX8Kb9c1dc7gfkCsQufCLdKPeZ4A8ZX156yFwSVBNAz3VpAku9jFHM+
EjkMI8bFAGk1F6gwppyipm7KAc4Dd9fYPcAkcZwoQH9LW6qMXN0Y2aGdGPWerYJ0dy7qHW8KImo9
HLJi+hWBbOtTopGcQRGkGOYmlp5zxNAJpD/gMDQZO23Jg6YSIhFl2tjgPNZJ+1QFYWa76kB32+tM
O4PJlPDj5YtIdm82ydgY24AY3JIIuZ6tSFicKGzIcE4l0lHZIfX8T1LB6xcNiOAcJFg+PXomspNP
7+wzNKzlibTHhMkgnEAg9VN+aWldeBRAIHkrWJ791rE0nIA6pcRsoluPi/EO7X+L/q1u4aj/nRlA
NHpmJMnWbMRYYzh1/uvBzYbz4OMdtfmKwA/ZeQjaqUD7zt0dpr7JHiWw8RI805KNlxeehDbVSWuf
kxuBlx6fmapbW7JVSjTSQ3EhhnnJh6Rv1JfLPX15pz8yz8NdtXMSUYx4Sxc6w4AxBt9jkvc7fGy6
f8HyhAbQdl/LmzryoOTwwV7/m5OFrbQiYvYIcmR2CXdV8wW4LHy2lWT+otrBFkmUBpBgMRluxMB4
MMQ6lYE4LFXnOU0c8KxCq+xtq0ZCinOxPQAs2hPE0CGWX/VA4e/gkCrwqEN7bw3sa6TIyX/2wX+M
7KxkbRZfbcM/CSgUTqBsMiL3tC6ewxI/w/oeUzL623NZu0AiraZdPCY5ZMay0R2ZCiySV87Yf8ee
o63IhSqfiEuCWuj28XDLoNZNM4Fef0ncDCpPD3LJYxymloriebi0K+YdzMVc3ryzXqJ2KJ6uIjOF
Qyg/6YH8hUHhgrauZsrAUqcEUQJZ8P2vDH33V8FkuwKIaKa9wmQSOA7lq8hVD0wKPDiEVfMtPAWo
o2QDXkxu56olmCjfCzWSJ0chlz1EIQ8Pzbt5U2Kw7ld5LtCfvTzMuW0HsyMbBtluC/WU3gSuLtnS
wxWXVdfeDPCe2mTPhVBXD7h11mIMOCRyxL3O1AIYY8BLlCVzG7IfslaXaSmE7VsM5UMgLZnP23Ph
ZNTjIGytRJgqSYIrywG3h1Nmp64xKHVQGi48jXYmpWicHCw4S9HZyR1tw3D/QYee5ei2hejHuqhn
WpSELduUemd/yCWJpt1DTjwZ5C4slq8JPEINC0AVvr+5411vO0kBK/HwO511e3LbFBXg9gQGXeBD
HgAJMyS3EmorVOiNvMwiTuS4gxZQkustt661yzlss9U+pF8c2uXhKVxk4W+AyE3HASHCZkBIceDZ
CPje/LD3Ba4Lpwpn06NNc1wh/siGspPiqitiItn5A2zGWgnJ6R+eaLhH/kCJMuo/cAts1yNsxLMm
shKLU+RPULtwq4QLRYMQQmhoBN1pGOF3qVCda1LgZXDNUFTpV1H/yd26ddd5bXgNkI7GgJtX4Lvw
o2e/9lv5DuqYXnwfbHlJPcWzt8rMZU0G6lDVYBctZSIooeiCF9mn+hYFmbf8imWG7ceKHnG9HcB6
+kk6TJVs7kfW8KvJN+8i9zTCP5D0NJC4LcrYE3UKwWKqU/Mp/yHgSh2eFZ/u/zQLZzPltuoBKsNp
V2JtmCg7nqIUL+FL+RqZDj6I871yWbIt12MNz97hjNYbitPLgmnWbxnHKZnPIqytllqY+2cSoWva
yBLo+9oIsvsgg5IX3qww6Gpjx/2Y9kyTQp/eT6Ra8lhASBVklAip3ZIdxyWgwDVpGoyVBnUQathc
Mtz/hchiS+ggscxQI5VzPieaV8rDGObpSFcIXP59Gq9QDzMfZoht651G2SpIZEjTLcrJF87m7D2F
sat5+0sI84pePQECLvzL6tdqnkWX69tOQYIqefajQx+dDz5kChR3QtRLPJFofUkhOOVVCPqU1mc2
1iod8k5ldsjcHuNo3Q4akuhvuk0YJrsyKANQjSZ880pOqjv+AJO/7/ZZDpV+OFGhaMfJ9IqyXbmi
BUwS5byU+kEfd4myXu1CzrVOL8erIkxjRPfD+P5MGpmA6YaKtZcre3s8KC6+rGR/93p89QffJVtN
5GgRstVHMBa2imDO2tZVYVKeBYwuBV5Qst2YhpccrmC1unL9VW6aiUQMtzAxoIXtQfV0Mk85P0G1
q0u3siw+ZkfHrSTArfirrQHwkQGJxKFq7KoEGiPQQaLwDIHissOsj0w0VRl5TM3PQoK76UZ6hVwm
tDIEmnHCMG5TWGMJxGmmexP8s0sFjOANfpKmCfXKpSckP6nOcYv2baHO5wUQcCAoFkiET77bnoTU
LTVeI0ZTDiKMsodGOtIdK8NzKNpOmbchCnAztYibvuIiC3+Tc5U7skEHUSGHkh6pWXeAd6LPKuwD
EDMagQrs0KnyRavZyaGrMnJDcU610VHBOz5D8n/x1MJUVG+OjMLJFgUT91qmwmmJU9kOHG7S11fP
aJZrg26s5N98jdHZh4q0TV/eNQkjL5aFEDMdM207C88NecN6wd8YWn0PDHwuPrefBY6qH6V66pfU
dFogN/0HeUHxyXX+Dplyjp5e6Hcry7heCC38gK5LjkcRXodWgx0lm3CKB4pz+Qf0sCu0TeEvVog6
Drvkh3Y+ZfHsTlRDy4/dKAuWjdNVstvSObTBtpXaJU8TwkLBY5I7QvVBa8/nvHcvxQFnrMAcdegc
bXEf1Pzn1nFkwScdjrAV4ALfsveaQ3GakpfvYlYg09wf5RQBSbtzlJp/8akhaBCgP7DCX5BLwwgE
dZJ+jz1eWVd7gtInHILuiMBchbuqhQRKzVD7uvUPDKfpWewi0Sp4AokN1WDkpZ9U+fw+memrdLNl
2jq3oPKEbM7/85l7+vH00CpOdsTKFJaYL2oNeTSSa+xx9d6jtdj+IiHI/t3bPGzevsRBO2EVUA0m
wuQc9HvST7qsWPydqbJ4RW2jO9XOB8ACsxJbiBZdtmlejSQUZ3YPXwpNIZ9MoMCOVhW2zbObpAsY
0HFCVsxAjJg2Lg7jbZcJEawCPSqi0cMBA01nBJ3zLDDRz99BTvih7VdSteHlo86mFloSW8KsoE1Y
ZLH6+kiPvyYjd19CtUCcYaY03oFPQzFYuhN8Vtxet6InZYDGzgGjuSzmMfsfHQ4uqWYUlznad/9I
2gtyTS8HhgHUk+UucvK2GQ7vMwAZowFqEjigRayKQvJ1zYx6enNCR/1C2Q/zorAteNDhnU3Gz97r
jOUMpXisBjpU4y+Vi1xqa7sEpTsCr8eQ5TBvQh4DgKsCnb7v5WdajHvNYzcTZbHj/OStO4GKq8d1
7QEKdryh7j6cJQZZ+ouIS5wrTxigxm7dFoc4ifT9572O9w2M7VYy2eP/wIXXRqmiu2B8l46rZb5b
U8eb61BhQ9qAe8P0VpsDG2KaabAfARhIPK03KmJgvEe9vgqUyQM8WpwE8DGhLd8UWs3RTj1f/sUl
8EzQoYkHuYfpzQH/5CKZfaWyhILlQaTDY6/rKGZYIpxhrGD7/oRPaO3SRwf2L2bl48K1j8utmuM9
GWsi+dfpZ8HhpFEMQrPNGsWTqY1xXULBBJ+a1H5RuLKRKYjNERoInkx18n7MFGY8XM1mVETKcR7S
wZRSR7bpv9MUxCn5EVkloeDQwSLaGoXSvEZWqbtfT1enBqA9vp/3K8IgsEuNjBkxplqsOGLUDq1R
0s8qqVdf54VrVd2qvFiy2uZAyPqzKqqEJxb3bWszuwB7sEsaT5gs6zizB23mCrSzVineftXR4BWC
1qfeDTmCbfOUZnNlSde2dJyGlMBKtTQETWeqtmmuGmo6Fojrz56N9IJOV/4q47aZhusNKhugzfj6
Rc3Rk+80Z1w0dlkpqA/iKIqbM5I5VK7edDsEr60pvjnMcaFhygbOXZaa5WO3bTf07aHenqSPV8W6
Z/cIm4hIlgT8WG9SxTskuw1HbiRehAgW0MuBM/D8b5EI1mrn+c92PZzbkJGFPmgTJzw0M0eOZORR
B56BBoO8qctiW+duZ9nbhppVVmljZE4cdmmHEMinHBc6sUudz0/vw5MLWGvGHMq7oweE2Ti9MdC/
TJb+oxHrgAVEPBUPjWjOdSikthPH0Os1sljQe+1KQu1ke80otVgwVUfkwYc2yyo2IDiEmP0kx1kG
Y5m1EPK4UMMQeQ5mrM2D7cXK1kImOp0noTK6FMlQyviEAe924xeCG6NHVU9Ud72seBQrFz1t6Mis
qvk+nAXmnEMIl0L0QYjOPS0+tKXzWyBvPlMlOGw8CLxiQ9BXPGWb1EQ8M3+anxIcZE6KnRImfVl0
OjERtKILDzzcwPs/2ulnCElzlwM+qMfAcoH27XEsiKKNpDmLDx0ZWq/leiAZMorSxcbHpw0UXpdx
Q0mFtQT+aiUCCqXpgziMWbmJ5MY0471Eh/x4nUu8wErhBOJQpotSdgJM757jMyVIhViZD5uPteaN
xYAO+yJkU7Sf4ujvDYayU1O5LhwGZ4LZ+d2cpyu3w64+HpJQ8VHEZ2n/5uDCNhgnqwRlSXQl9VC/
2pIsHcSIDAHUNeplowdEKGbYroR1lu869+SppTxe+66RkwuMzb/LiSYDIl7wtxk6ucL0MALpkUTu
OFm87blLpSHdo26SkPWYxWL9IhPEYJ4tq5krdEXlkHFi1kyirF03WCnuvPrPkxsTNuOfmk8ezUB7
GClmbVRJebkCkkPZevRlw3xw4w8w4w7o/kPC318FTr+KvjnVyH4EaBKSHPrIKNWJtUysWVjgRXou
374J5ZdxTo9DJH/y9XVOEPPyUDBAv0TsGXsSxYW9vQzlohwYtSifYXWSTLTSBCoPbD0uV4HqNnOQ
AsJAglbhJs7CAQGsw3gPlIdoKfdEW9Rf+WvZ+3DMHGYVSngY/4DcYIxO29M19WBLsEOP6GwuDILU
pDyWD3Bby3mkAVXn5zOkuEEA7g3nxWb0/F4MSWvSfMvoUVzWb+b+YhhrmkeofhTpDkWWuhp1D592
/CAu48AYNDz/M3+I2daYr0Yk6/8eY08ZAdGQdcVCwmOVDqV/G5UcsYCie9KsvxSAt3z+g0S81YG8
9Fj5fBGSqkvojl9sjRBydzyBYoSvbE8lQsiNoAhUWLy0btkeWMVnBMFdf2JzFrCHlPxXLwR4wG02
ALPjhe1EMI1lnE6bVgsoL544iZ4HN4c0Jp+MIfsFMinHczUwOVf362CEPN/GoW726BUQcH5QOPZt
o6THs+MERdGVl5B8PfxDOeZLNnBVGZDRwHD++HTMSq718q+TIjCTG/yTfOmN+/cgIakPNQq65m0R
KbR7eJiiYqj+NHkEUweD8h0N4IW6C3BusrRkVub0x2AGxblCNhUxgXR02dCzowDMYXE15BgOtU14
RCPp7ym7vjHv4XPXP/N37BGVVojdyep9TBlBcX7g8WK7ZzQTuHa2Ah5nJ2Y8eQSkIYV6zqqbsfb/
QUTAWxp1gZPlWlxBvmnDhNMHBncSCvxSFs8xXYO0qyfNM3cQHCsqCAGy3i3SrtXWAwmeHodjAPCb
/n2pS5GuGcOmEU85FRkKH13e4T+mThcCDLUvcrD2B5kmFiBwCb5iTZFA+/gL6/8INersm2o97v4C
z8dpbIebABSTHfjTEdBpM2SYZKPS/+FBFIcGsuVBrPIUqSYgPkzSHUmoFpU1wShxfqU23/+KKlep
M2Jezh7vBtT1wyZOr5kFKjExtz3NQvL9TjczZUzqTFflxIaq2//0N0f9bIvMpUo9GdgZnyl3Xu3q
CFv7FGvS/nhqeaAV08VkErBLRYt5/sU8cQl95RiBsXWgc2qp+6PGtsH3p3wet7PdbwWjf2JGUTf6
nH5eh20k7gLLYcNCnCgQY/FZhIyUlc5ovtmZzp9UOkt3QhnXSpmupSH0gzi3LufFOvAKXpwmahEI
JQtDoViXMVhPxSFyzhgNz3nrr6mAhCKfUtIBD0eLFbQ1HIFULjJNzvsp5/pYg/PCaYM7vy0UEH5f
aJ7ObovJ0cpOFwBTc6ajKlGNKp5cUTKwKo08WSShOnT0540N+SWHH8N/ZExEzqW6/uk+mDaa/ix+
68Ot7ymZ+sNPYeTiW0IRqnYMDUZNk2QQu7L9EV9D8s1pAfT9rsqRT9TBmowkNEtNSxFDBWOF5psH
ZNf7akMXWYGskx+MKQH0XXEgQ7VvkMXTlnfqgkWU79WVQMmP646PD6V+Ojl6bXbs6HW2UzwJMN+y
dSCWLuuNqylCwMIhJf5jVoKpf3Z0jaiIPWfcK6bhaL1rB8+Kl6KCS46LP3Ws1TqlKFrytBM1mMCs
H/HoiJOdUIshJK88OARvcyP5Tl2SZ4udc9GQpWX9cyxlE9GOXG1ipQv73pFezvMpeInK3U6uj65h
hyRAwleGDhgrD37VTmrjJyj9e/RKO2ABi/0aplOEtAAcBzZE95hkGHcl9DvLN0emlLOBNufcpdEy
tZh4hq3GCwLd/hm3Wl4RK+PBfQdQPU6iJ/7gL7+KUBSNCn9dyeVWP5mlzooW7KIDhxN1G+oQr1Aw
Pz6A0DqSLzAee997C9Hn1k2mBJfyoUqIwcsNdn2z9KZSo7C2SKZyxMY4P3KdW8EC4+e8UwTQot8f
OkJAcULaI6/l1uiyrWPvqIAfPfUc6yj1qvP+veHT5FFBiaeH9h3EaAbvNMF0zApCy07QdhZND+M8
V0UnLhFC1DCBQhAhBDgIbaESSl1FCWFfEjKIWeodptoxsZtNRYawHCNfRBjj1TSyFRvf/Jhoi1Ry
oyPNX8QTv5Jej5T+sFzRrEDlGUs3WMvQWWX78xaYsCLDEJDMG3NMLuJYuEVJnR64S/rHtdtYqZ9J
t90opoq08WndptCdjq8aAJbpyN7PPI3YA06xJEihVwkrFkhGr4pQOz+N/AAJzIIWxh7dt+EF23MG
oGVDtaFofne/D8plikZAVEspiwDWAI1K5Fw+FUdzl0f3rjsy2+RNfbBphBXNdbqEgq/IAFuW6z6J
3/TEL4Hfs4ZoW4wQlyEr0V9qp3qftIarmYX27X2A+oo1NZ5YtwIZa2rApc607ceUvI0fLFBy/AK4
IFxk4RnWlik67dSEAddNQxSpo2FKgHZSJnxITq/4ATuqq2Lq2pPNjdQz9mBxFoWZaUM5T8kk0QfS
6eMjHthDrcJGhQxs35g10wnsOcD2qZb/1a5DB62pRYMB4VcR1UcCNKJKBzkkRk2sfzYLS0HwGYjF
OF3INVxyN20ldUlXGS25k3UuGOXuiE4CTorzgpQroZY3bgBP6KnRWihZX/I5j22ptua4BT9jf4MD
9hpWPLWD5OFpMHVAhVOR32B7UcSV/9GRn6u683IFV981hynw0lQj94KlC6NdJGh/pIIK5ZT2UXBg
hHCHACOvtbdY+YJp7bu+Xip5vMR72JgvHGVxbhtjc1KOyxfvOwMrVXbir2lCYD0gTztLNiW5Um40
kNgz1nXedoUmN0pmKzkuUT6CsSigS6lc4ul1/+TizzNEhNdEs0nuWApWBHOMh+tUMbUhQ8ser5tj
7MUQFGYKUGGJTm2mFlW9oumakrRqrd3Ym5Nu7BPReRywlGdxtyLHBh2l0nXYNdpz7F7ZE8Q6AyBr
0eI01dmkzem1x10h0Qjk77JEo/Wp1mBETnNkWAb7jQHtA0EM3UXGl5CqJzVM3F/831hVeSyQolj3
/I4E9aZU6bQH053yGIUtaD/oAWssOv5O+gIKJIxyj71vUpH5ncX36X99lDwDpJWaTMRIlKhLeFVV
G+ycCoYHul9Y2VHiS18RwsTyq8tHDNymkAtx52lAzVbpxf1a5qVGntJiG/kbmmxlfAj5aYQZcua/
NpRIDhGiP6bNGM70Rk5N1ycZ0KLXki2YShlQ+VVwYQgFU41VEq3WdB8XhSmgJXq/ErfdTGmBnX1J
YDVWIvfUGakPg1PyZ6MMi4LTpjcBt5Fh3PcF2zwojg8lFZ5eIibZlWwEJmoGroyIR521qrn9yPwd
Tn6dFqdxEi3uN86bLe4jmhm6aITPvPsu1rYakmrh3Gq8fqdbjmWlbjzcPIFrS+6pnStobrd8tf0Y
jFZrt3+kLEV5sbbZ23lBWrUw54786i6R5TyWmrzmWzzglCprsYOyrlzMD1lfU9hpgC4aAPDw5ysS
Sr418qjKNbZxMX8uqbs45icy+mdVojbtUuDMDQ8kC/cd8HOHyL2zFUiqHOcTSTBly8pJkGVZRAwE
Omh3RAJIE3RJI42aswF6D4N/f6cAOLqKuHhS9d13HHMRzQwKu59x4kaYb9JGQjBg5TKlV1m6qYLN
fCokDYsrR5kFHVdECF+BaM13bXWuWR0bP8e6k2z9FnvBLs+q7QIhz37O27xf3Jmbf2a/mfOvljFr
nR4vXFuz9E6YGPLiOhFBuE54DHGfIcJfVZ426dD1MAhVtIQoW1gfLUI8Ce3FnJCTYhMme+zJUHI1
LRvq2U9qrGFU6r6o4OSlNk7th0NeIQx3DjLiS/HZqGGbxitZdB0Qwmt/b+bt7p+waCsI93U0egQ1
kKE0ZvjHaW+LefUNlXnGWq0N66AFZac05IVMEQtTwlAVcfvsWi68SMHq16QMUnttoffO2hEGdzgm
/twSyv4or0lFuL1816Wn4XUHM2wApI+s+L4/mD2Nq7p2UcFdFjsuyLPZwpQXzm6puf8Tx4aGQVPA
CPFq38MhPjaz912I0XitlOP/iZt6OKERRSluXG0XU6ny0G1+rJm2o7cDBxka6YDTG4qO2KqI9LIf
mw2TMJyEUThrllyE4dlYMaLI+0Dv61ndcXo6zzxouStw4kpIZ340lcYC3PPMishp0v5XTaI/c4xl
/WodPJ9PyI5Zeq5SfSe73AvOowMIY2mWZ/yJKDFy1uG71dVJCnS5gcA6XWIUpNq2NqNzRf1udB/U
OsGkERU4btWvYpcUn5kI0p8mqzTON95LFEjuRCBHlJthPizON2BLkMyjfrbeWM91c1yWorLsmNmI
aTMx8DdDD2+YDlXupkOG/AmNZLx8zWKr1pXHIWjkQ2qSeBVBJi2uzCrlzvSYDwJQguzsKf4zkLj1
5ty6uoQ7Jwi9vOu5EJGPVj2wi3tGVxdFjSufBsytQ/w6hnr1rMsSl+I3yDV4kwbTWpxfnC5NBVwg
BOXAohCLSmj/4/iGYC1lJVx8pAzZA/ewWwwiiM/+TCBXGo9DeKu6B6tzTOh17XajKFcj+CbObgVl
yP03AgOqVS1sk653KLRItqbz7IZDY3Z+gUbUCp+G5+eGjRqT9G40+yU2X4KEHBjJ0u7Cl25y20pK
lup7z1LmXwonyEYxhVoUiZjhY86z40ErSrI7SJua2EIe6JO2Rvs1ltE1eI2/pLuVAzlxAoqFG/Is
L88RSeSwyetzmpSBt+2Jo4A4qQKhn5sg7mmoHlsUDyy4CPpvbCF423i3xf8bfj/hSD3XjVo/7gWO
rx4ouiY5ydZEsxd2CU1EeJ4rBN7LjyiC2bBy3tlsdZFnY6AKKYPHn9ij7Mke3OIFSMAK/MAkECE+
BdFJx2I2WHqeQrfQdrE3NYuco72ug7ROams7mGV3h+PdlXLJeQ9YGnEamyIOC3XyKtdHABJmpI/J
q9BGFEge4583B7sM3szEs+BN4Gv+y2SCKlpm8rMmaGa8a+gXEvueNzN0gG9nJ+XFD1QfbTDQrZQi
YhzKo17WcVW50xitCxN2nikanYFVSWO0GdYs63+j9VPGcto7UPcBzpiCdE4bfzpjV0KscSrU2Ril
7MUhPDj4UPoQC1/1HHd1w67m6m4zojProP8dgiVBUcu+NwOUtkWYxnaf3lqf67eEg7h7a7DtZ8gy
yQK3H0JwJRbwS/tSeaHkyAKqmVDWt1hIoh5xAsaD0TLTztoS8Iuj64hsdVQ3Gn7JCEStInJIiUQ1
qhBZuCmK1tWg94g5IVA00+ZsxNpycjeaPaC4icgzXVDfUmrPB0YOyciSh6FtuvxGaac1AL4YHSp9
J5IgqlfOzWq15wKqH2puNRXNuq9/8F9OX3vMDhWWw3DCVlWSBOXo461AIqPn36B5m/HdMUuGRM9V
Rot2IB0mg9McKR/qfaNqCxogWAcDoqxKfVuEp0Qv3CH8vMJMYdpobWxFzBkAe2QKdHS/U+E2wXiP
1wm+kafiQEQWCdRh6XB5XKlwfO4xLRtYYyn0owTCNrDoLlYusqawmmYUlguYYCi7TxfHUD7UGNHB
R+W9C6jdbA95trnyOdaH/hAolkU3hY7iZ63PQvvt1yHsMo3bpVH2n4LwBlTQ7mVurX4aklk2oDFK
H+Gjfm5wWxVoNsV4J1rafU5PV2D1bkL+uPpPKeGsKAZHu6kr5EIF5Ks9lvUC6X0jXsdYWKmpilor
P/9ugnwMIyOhLwnlUowc5vjVqlTMCvK2pRSpezKHmYc7VsQQbIDDEM1VPU7CybhNd3Tv4EnBtTA5
Ofq8y4asecBiCJ70XqsB6TVhAIH1qpGsBZWJzOI8e6YzK+G92/gVQffNXfk6JfjEXHtOXyRry34y
lvu++pVizw5GPvjsSDx6mWSVreM2dbYC54+8poVGkcqy/7zRo1KZK3YAeHiX+uERA1fgUPsErObE
05BJI+eQ1e1bPCpYmEAF1m1C2mLNE51Fxz8VOS0ZcVg1Nku4vANBv8tElf/INVYB+Oa08NtQak6g
85vjh4knGxXcvqTEhiT6uJLUBQpIHzc0MbiU5QEhuBaG2+6/rlJYiX7waBNlLcftJUNKL2br5iBv
/+xTpgTZ2LzRsQNJj9347T4rIwh/WNHJyOlXOYlVA6Kb4SBY1LPV2MRvwytIueciPWkM1WHICDyY
IRhK0DWkNM1y8+PrEtBAaFNCWAe0WwjplZj98whL5K9X5mKgQZqoHZeNaaGYE6ajPGTl01FQ+lYS
Xo7YuMEvneulpQg4jD8GeP37yGphp38i+YqlOI0i+jt7V9k36Iu2AF4zDaR6cv5uJuC2dJyisUBD
zgqHYN7k1BCaXTwTkQ5MAJ6Md1JuOC18PUVY2SLfDOebT47tL7k/SZF5FMpnvNztXkoVqXMTMPYI
ReBQf8R0I8F4XYghSZPJMqGrXW/k0ZQMJ6LE3V8gm2BK44dwmlEQJlpgPgm2prtvkANEXWO3CQDZ
4fbcoqDDc2Q1j2haVzhH6qo/wr7olyKVGC6DSR5yswZ6wTWDF+Xi9hREqrTp3w+JIT2Egmhk5RcI
+Dy3u0bvnenoh98WHuxiUKImKe/drvJmF7ufZKY2/5QTxH9Q5aOaTMwGEsbmrkY8naZwdwBTagnb
JwbFTzzJMu/WgHY/URIkEWJmDtt/v6Thmh/NVGjZbzZYpvz1Bxcd4XjaAGTQLW4fQVOtIR0rGxZ9
dnitDhzwPCazCefAp+doVF/6uH/Rm2bHbmGuVYpKCdNcP/ABpNkMoKe4G1Yg0XMge1GFUpGNxKPb
ozC/OGpt/JWho6KNEfO4VisAWz8fRAkLownzvp6Z//qUarX5A4hIYr2kZTD+3sKNtnmc04T3dl5R
TbnoW+euO13mfiYDV8El2c3bF4F2bc2vwemE4HKINzk23Z2D0N+Nzn+KbxLfMMrDksnIQaV2d7x2
2Ptfzzu/bYL6EkMUnQLWRPOfPPXU5jm0KuYoNmvhfE1nRlzSu3NFv/l3/R6ttfagbcG32S+VBVcK
F4qCv7SKIEJITqKfEcDcwvkOd50OSZhnDnNjehAzW4fvYViqdgDAbxEA7pdmw6GygPQS/W/zxqEg
QFikjyiI7ULIRNXK4t6OtRY2GikyXMYqs8sK/6OrUQ90N4myV6LP0j5bpdDlb9m7UuOFjCN+zPkW
L3KTze+EEvHYQCl/UVGB6NrIzMB0uWT8OS0NKzE7TsF0QBxTv312Hu5AW2N/nK+4nfC5tkj4+qOb
E1kx1nbSjfW3o4/ud7ZVnb9g53d42v6Sn2g5g/mR8fpZZVdy57UUjcIURW8rDSuglGMjUnmczztW
vL5kHDCnmWVyqti8N0p/ytjkF+RZQg9+qdw0i3pNAFd6O7wDziPgi66IBNxBgDQGcVbO138E68ja
rMUjvEqUWaU894wZLJldWiYrbpBtfDQbHQNL6HcwdaP6HRkkfIhCi2vRaeEz8mmF/nYb53MHVWhh
Zeswbc9fW4Pdt4dcUgYQ6Ky5qcRym3nR3jVWY0QfbnCqBSV4cXasgdwfgRbMwGVFU0wXpO4ridHU
SspXQ0VXAM+sb7t0ckA/gmZK/HePtM7NHV8jKptvopIVY6r3lretWZw7OapOfBIETFxHhjLXWbSX
RyKYxsoo/TfYTOEa5Ye7ze3NuJlByc9wWWTiU0Es46U8nIOE1690FBzAUGe6LkbpWRmBvgaNa5W3
dUkSqSykPdvHEvvDOFMSiWMGbSZJoeIW+wdGq/syRoFJ2iFGUYZrwIM+vKeSYzAY7G91mYIgbg8s
aa615OdZgy3DKPt9/X223VvjR9qo+SnCgByMHx9DsA3sWMRf8I4bfOzAVPRC5QVldRvfoy20hlW6
RUyxhesdypn8cEHxU/L0RP6J94rUBi99rdk2XjwtzrtmmQSF2K+0pxVSSQ+1Xk0RNO/Qu92cnxxi
hCz+5eSf0ncqQRlECyojQwDCYzyG2IZxLvdUUZGtbsqammkc9neKPns32StE+x3poSdN9S2goI4p
Jrxf8JRI0mU40Gzi6+9sV4Edcykq+S+TXmtUh0SCxmP6pRe9Detp64QLALlJClga5qi6tZBEMVEO
hIb/LVm13d2O7PIAGFFJs3DeNXLsAm78GFIgsj2IZBJtsaq5VEiE7TcN0FiP4ikbdsvV03762n7y
BnHOyhJG8RapL/PkNFJha96TKro78NGPzaI3q22lI1taEufo6+pbrBH8VmSs1l9AfrOMsqVeeBGE
RSvuco3fHp8/1KIdOTMBv1DJuJAgovivDhXQGVfdBqcWGBEbPvNyjSJvirRLukx/CoSIEKByv+Ab
/ymaG37OkeweX5sihzF4WIhcpBFhUkt7AGSYGdKqiERiSnYQLZif5AvD823lzA0HxsUdYYV1JQFY
W3uU6aFc7q0unVOHMnjmK9wOEaytn2jTjxqB2hr3YiB/VVaVDjHBzStaoj/Ji7earEinwqkzv9Yr
UEbwJ7i57U/T5zq7G5zKoQ2bP2YdkqWfbS8GXaxXZ62/mQasIlBVHfrdxkOb9zEVbw+2BmDCVAGD
H3liHHvSJs8XzRHYyHCMhWF8OdKYiESbcyDGluF314mMWK/0MMC/GL8ufk1B++3M3ZIYoc3Uaslo
aBk9CmagJeF4bibnOQNGy/XApfo794wlEuDL1KgO0IxJe4OA4E0MnGOph6oSmhbXnjjYD4ollIkZ
zKCegdj05qt8bmVBxyMwNJhv2kwttGTarCdlcUShM8TETpBtpyNW9RhaZP9Gbu+hmqO1TxByG3yc
MUNiATS1r6vGh8hxUKwYglkOGoHGcf2o8FiwBQD8ysv6r0ERa3qH0chBTBIhX506QOq6qQOga3CH
hdikkxRDMH2G3P0uf4PLwvAHA4e/YCeiTr2bVGdTB0lQ+OkXOC4ezD2j1ZGoNawaljjv2FDofW+D
hDzeYXnoagsc5AjjGKgjKV6Rk6E+iqy3XfHyyDgfDaKnHHtynpB49s/M3iRGxxgCz0JFYlVwU2nj
iA0LQ6BYOBxnmC4YrMv+eWA0UVh04x0a1KhQCMrH99GYLDXe5eZh63B0rWTqZH/Scl7r5QZoB5pa
J+ov65fN/5aZQSSyz4LSy6hhl2IIvU1zxJfUgfsbuVlghnmaoRyy27auDy4pHTHPfDJrC/KcJpAe
FMuDAVo8zDtal2jmNTQAVVJAogqk71SnsmfXH8x+wYoJPu9y/tF9n91dGopmUtOf4STJkgfo0btr
yZZ32Fvd033+vesqvvhf0NhFdqlYC4+iI044H6RyuN05XgiiaD4c0JwjUR9keS3d2xcdwHSk7gWp
JKEOLXmorYNst/wmccPHDC5aw4+IAS8Dbc/AP1LhUVFp2dzr209ScJ3sbq5aae/Zzoczh62oe5C3
atm5eLXjlfpZuCddOZOgSSOwlnb2V6dOWznFtfGeOzSnFMaAjWpIR95eou8nlz6yRfz39tLIvzh1
jmYups4Qc1J/U3UHln8ifE4LXkLc1qigAwxCJGvS30LR1uUfFZcJB9pzQh5VJjQd1NvS0LlToQqM
pR+isuI/hNIdVFAlJ31+7s0JaEQ6vEG67LjKxGXiaFicBbfi8JBAFtkr8fbSvArRwlpvO7zOk3yi
YpkWbz2Txbn+lF/2hzreRALF/LiBI4AOKpMbs+V8l3yIX4SEuDqYEn8LI4CvryCJICPE5q2Z6oJ2
AgBzbJVz6HH5b0zJWBzOR9KnJA8VZwfYt7jm6R17ZhJLJT38EfQQagFKXCtvaIURB1q6gV/gQYc7
7iN5jowGdgIWLfSdSdMobkdaopWsO9Yms3HEb2RfJjfOxyICmqMwf+viKQ0Hplq9S3ufu8EN5wJ5
xDcbrea876bKy7w3153WVCU8YhdLnm8iX8xT2mKhw+9kfMXhWwjiknGDUbTtdqpeDDZTUuSYUGDh
xRLdnZ2EqQm3dEHpawLqkB82Z2vYQhVOUY9mpQDuH0058b9+KYahBMv5C2P7MNKNh4bZMcBMwiEO
VKCIO847be/QdjtAgmQnGf1Ry/Nx5KjnSr+ni6TcnC5QDY3YklZOvmfKHuIbxfLPof7aCSSE9DI0
LZO/0lYw84V35hJs9t5T4dC4i6hZYLah0akBtM197p1/BWI20Bz+PW6oTQn2xKzhW6aamCJLg8Jh
3iTnPqVjswYmAjTqJsB+npI8PxpfXRW6bYfseuyqxGXBl/2XpuzBGo2xW9SCZOmsvSftCPSrY1Yz
OQN28hbevhHneWvPp4dihLddrCbo86KWfVJCYWbOEtp/2tTtPwfWL/0s0X745WjbwZogZVsMc2nB
y47qbwk+og8yTG9DHaa4jyiKStYXAlq/n973lZg/cRE3yLDe2URVXKaJ8N0dgbkzO/rNDKy3TgVT
Kr+jVsa2Klt24f9HrjuAcLQNgmiNSAcQix91oqY6/aP3gNIRDsJMF4OB8Hy9znYL3PsiX5S6goVd
0SDNKU8h3A+FyWKO13IxjTB3n395cYifz3GsaZkNtZRCQ/n9w2FvgW2GT0nrtZ/jzcDtYpqnpF2o
f8n9K8actW4YOgTQu9g6WQxKk177NCLrm5PseNoyvSz5hM/E3UmhqIG5NT1yIHOaGM7FH8OTxGOA
+vrZoikDo1HgON4WBGWEYRKxqual+2hjHdloRMt6QD2b9wA14xHgeZBqsV6ohgikU4+mBKVbpqF/
XMoMMQ3YuVAA/n5St/qidFBC4amzdZaVURmEI0YmgKG13bvGJN55JRRpn1+5PC5lzWafeEu/YfqN
IOyE0AIbGq4W1mMDkv2bOBp4I+I+TJF9G0/AOzhiCnqoL4RyxapJqcC/e+oo4e3F/DY30Zm2WtEQ
ybRPmx5hp3HQyL8PADgqdj2PPOsd0PuBYy0KozzJWKlYvtlDZWtuUWw86K9Ff2MduPW3IEfH+dnV
x9E22Oj85EmcTNttMs1tF2KYkLdcHSCZy2rdTulMZj/DkvOMAFjwNBVc61kttCHp+fg5aS6gqLfx
HCBk+PhLIqnb2VmF7lB1ImDSlmHupPpQ2B1SUTRUU3DxVOUxK8EnLqOP+eh1Pu4OXMijTbaKVYOx
el4ssf8+vB/BlfJzk08xc4c5jvMw4J2DRBxaqEK3PIaOYrfGryzg14QJRGmYOP9fqIk15XnpVqWp
3yvgCz31aQaNgUrD6Hx3n5G6yU1kMNM7GsZkd3KHnzN8IBvEwNACUByeZ7HXpNulq6SofDHnTFoZ
AIEvvnocTRMYZQrJuMAVLIbIveq5ktwB7TmnMOJJksZcwBy/3Vy0IgUXtEANKt9U1mRHAC1c3WET
r+LqtugeTSKF9NPI7YJK772BNNDF4SqqmzysaQct1gzhO9mIKhOIW8DnE9OP6Cr86h/beDXsvB46
yOpMtS674X3b8vMfPRRUDe2xQXf8mkHvKm/4NXlUyYx9fMl2HJvl8Ox4Gy+pgi7RKXrMHD09TXwH
ONxzfdv8JkNhaANjtIjX+gG+JR8e0ZHnCzNqtiZhJDtDHzem6yXPoaIwcWpEACmNfdvpMo57IxjC
AeSB0yA6V3RUfkfnjnEQi8aGlJv1E87yTqxOG7+d0qyFcwaijpBtpFUYNPELVGs0y8AS8FRPBSLZ
Y6J2xd4/BlYu+SSnxwlBlWAZiY9BReeLfd5zdaOOlcq2r4/wn5BiyNXLa/uZeAwyhflhmuSKC/z9
UciLKZ+OSMovmZwtesh4stx7BnsOHHJjOeTsAwscbRvUCLVFD+SdG9PQLVXuQL2IAhlpAC7La4Wj
8HySLL1pY76S3+KPiLRRVriDLS3JFPTux53zaaofF68qKvaILya0wI/hFJix6xHCcvOO4p6gXU+h
/NdboOvarMsd99WVd2NZa1u4EEIGqnrs6n4n0Qhq4DrhZ/zSlV8vx8q1qetjDfYtA1nAyfGQ7t4b
IMn50wdnkJ2OEpRoQabjEkSt7dK3xpEHoBpOGV1wEnenlkZsiBnn7xomnZL0agh5BQCCtbqBN48K
7pHOra4ozmWpvVZ0ZX2Ic0/p5DnZKti2zCVDY7rzmnz4td2yeFEYsgTfSG3HqpoCfNJuBkOCLnkI
pbt8duWmhAqCT6skYt3re3fEt9uh66khnrAECFO4k33Pfl2zzAXJtNnDiA+HKTDH9mB5dCwUCAoO
YGFzMQPxinpwJH/MqDRdtbfyzpy/MdjXltv/q0z6RtZQ+eNs5JFBxHh1xc0tOAAhLrfrfPt538BI
DdqYZUV14yt0rndQ6NiBKJUAEEzDuxsVZwLUS6uokVTf6x3SHk3ZsZMh35qJHN4sBe14bPJeLk2Q
opVlmkgm0VWGxVdzcyPaEq1GYE2/Ji26IohS++hB14VzPQ557SqbYiGhHBp7Vvm86z3RHQNbUc6X
K7SGYRq/P1GEmNl6B2CcpnqRvHRZ3oXEhNw/eT9x2rmMIFOraJ/HBJeObkfMmDGcrOJItaHns6PV
o4/35iwy8npY/8zqGsNNbOB5/V/0vAXO2YNuUqjW/zgdgcHd4x2JqoE6Hfj8e4l54tx2In+IDNTa
m+t7I+Zl4DNlKFcU+kLxu4ZMRzy8FOxTMwV25P6crnZh7bZ12+kkrZEMRHtZY2rwfX8HJJ6IF8NP
VgCSrJvmGTDxlrTblgIIuHwBilFIAdmOHiIUM6MURcaYjMA/6k41mYJyjYrYeFsP1ipPlGcSOhDj
zSMv8Cmgn4SIX9YO8J75lc+BTdPRSdOaMQVLDKoymGDICIIFdJNEroeALwVyEsMx0SD30AQ7pADU
n5U6uREPKB5iX2f8MWxJvvXx8Y2MyafN0PZAcEJDNgbLng1cNMqbKBJegqdqiHDftZEHHx6gMOJF
SK1wiPGgt0NzzsLqssyY+EyNi4fivOyjRgf4ivZyMu8L9hrUHFitLQDGyo+IFAL6rHRw2TqWrlGx
zKKvaMwVxt4YOF+hGH8CiAq1qcylD4QICcPiMiij1jJtp9uNFS2S0d3Ms/K37N4VzVGYw6ErDajG
fWQnz5xcWTx4YRiIAoqJFF5H2AnVpnYQkS6Jpb/YqTs0+UcPoLiwUdXTvENRgPfc/yfBsgm1Nb6d
IhoRtEyWUSX8cBCPCl0Qc+mGvKBasY3d7pejr6QvloSarfVGr+K+Un61DGHUulv4WU7zizyDWnaM
84kyEMz6XeIVXAnU4axRgxuJsIPYITCc6phsyH2d7A7Hf8w3f5KBL7TwerBq5GFteIiVI6lhb/+Q
NoLGSgQqqCQKpKgMGBY8VVrtAVRHMvmRWstIQQcwXX4LryryPC6B/eB+PiNcVkTqz48HAL8m0SUK
YIg2RRKYPYN7tkH1FPMGc422xFfIs/KLceuN2cv8XOc29PCT540cvQr9o9Rh6NdWjS1B6QgPUGYm
heXHWzmbw4lQd+MSPswVUVTyep6naa3b+NwSJmb6f2gnyTFlfqfZZURrdZIF41gYN32KcR00LDhr
SpjGHGxE6Mkp6lV/8hQ43s/6wP1I7vZwhEZtvpUwqxYmrWemQG/z6gDl6jw5CHy3mxuGGx78sF5W
a/5RNA3lqzblkqskfEfcVBGveB0wppUBbY8u0px9/JO4/GgCfRVgcqnL9zCF0s7HM7XdCUq6dhdp
Pk/Rhc3rPqRTWb+lZw/1xPrQ5tswfTuCUM0pndeIcH1an/Pug9nOyY+fHgw1d1ET4yzaZiK+TAIn
2p9E2rCk9sDi0VvEH6b0T3WgHyR6CA3OwXJB9oFBgg8gi4jeDz0WhLPFho5+w09D9U7pSuhLv7lI
qBX0m6rt84ynpDDefRP9+bSXdSaRIj/BKqhfwydxNrZs71LJflEOW0JvB9yr79f+k5UcDe3E35Rw
e7KP6E0/M5mZ/RNbPSr/XfhgLd7pb6eYD4aksc6oEu23pliprtBGZ/9B38e2++ewwnCFjuEGk2cg
XneYyh4s6Tm0NhJCGMc/rL2Luy3+9ilICSi9lNT6NAAuru4SDbaCNub8bThQDN9j4ggqWcZcgp/s
ZhKofTCKAOzJwxx0f1ALBASGsetjLuiTimCMcAmLTtfIG6UNeSZe04bnlZJUAyhH+PIH5z7mxUgo
jse3+ZISWwZZLw5YwU5MJmdWHsYvnGyAJjm+QIBsvY90ClO+OUqqXiS5ZpYXbNxfCXRlG1ELjQ+m
b31rhGUowco/xwH29m5ZYmXxpAf+L/CbgTzoHNH6XUe+e4vybUir8TbPHEVbRr0fKbtauLh08AvQ
VkiZdebsuWKMn2h6JnVVA7dR3vxwBx1KhU3qiYoRDRU/sL6lXZB6jg/CrrXUrAjFoi1uL0k5IVkP
iMQwjTLqHyLoEavTzco8t0Ci3zAr89hC2VYiCg40eHNT7S42EAvNh127i9V/RHRnAYRJVjJMpZty
8b0aIiTwRqF7DjZFsR/VVWJjEqXsJ9rVHegOt2rcXbBtlHOVzBC1NNFuu2755Y3jjPN3OsvkmCeW
B4wZb6BjuYlx3jBezo2e3zL/w+jzy/Gl4WNbvxMalCJhYv2mfjZjsUFrot9eKGzbCKvqVMggqanQ
2Llo8+gAI88nGTgHNpHfb8gIixwZ7s1KWeEwJ6sOziowAihMTw0h3mgOkk+ltJWgCtoT/4JuUjf9
jihvBriU6N+L2cbJSebyaEf2fN+sf4Mz+OI8pIlPKqtSknMR2NUHfrIOtEg+s9c8SdTE7GgM3cCq
pXYjLOSB9wTkIlJyvTWoX18KlUDu6xYIwpEbTmKO/1mS6SyIOxRmSBbpnQXo+WY1rcDg+61roKMU
o7aoFNW40/pCxLJgJ7kejSrqedF2QvOQd7TLpqEI5lZ5PjZbiuFB+8JTvLZBG9pKrIotkXVWU4GI
6Iz91IliET55jvwHZ4Sq4qJtSHcw+80lCXy97ErSoJor0FXjtlkVDMRHGp4DJwqz/T3TrlNuidEn
efqRkS/0PwBVitYzlK4OXHEJR+c8On5JcRIv3EtrXHscp7eD6sAK3R9G+tWeb+ABz1FH/R0GgK5i
YHOG9m0o6T9WaQ532rwRhY/qARlhYMSEsUGUqcLIEPeR1/8j4jkQEsuKjuV0/Ww+sUonFRbyuvaD
KvXpopbXl7LQ025MJE+RbAG4UOVf8qpjEwDuXN5WluOgI2jwPecCf1PBeb3XVxhKzawv2N+udq7q
3A8lHuQjDieCt4PWFuxvX8IWXXa4cvw7/TLFAbMI6uI8uQUD1s+jWXXma2fygCrv5x+hTCwnRp8z
hu5IH59UfC05tfFkOGwh+SQvX2uhjEFFGqt2un9DpUkdNpdwGRafAF8QyuwILtrdg+8EOUKBleXv
piG99Tj+41M/zRnHDgAIjCaZyP33I7aQpd00c+J82RX9OPUKfahWEHH7DyFFKqUYLfeg907+7r7y
TVXmjYsyXDTQL91+1EKAjGhnAfeGCjmbJqNxF4E7P58cibDJUF+VL7uD3GOoKC95UZ/6PweARCNM
4/mvZwerrBofr7EiSQyp8lrt2LffCI9Udt/RJu5nFdqJaIzXYihy5Vt8oF+CZKrMBygci6kYr4Eg
NEuSXU2oLrj3NA94kRyvD0g7v5X68mC07sOxrTJxZv5lcIX7qD62Yz9a/6dNfU/4PbijsZIMQzGF
B1YKbQHYenNt8OUcruYywu5vUYacOTywo2Dkr88bsgFXQxAPwo+ozdehlNFdBiAoFSvc06eMcW8i
pUEmR2FdisPSGxzGVlkv31j9OlrfXms/9hxLFNQiDsz4nrrqXvQqzDpmJzvW19NsFlOpkDXnEwWU
IgI6QRgYIgI4ASBUG5er7llWjuu8383hE6Yocij9aHXf7blX+/GdAcUQSJ2CO5OngdwfltdJDoMo
YKAPniBCQ95Usf7gpXt3jVTr2gXGsCMR3k+HSeB1QgrzBzLMSnxN0DI4AH0WVMrH5T4qDMaT/lmv
iw6F6VKr9UH4cxKdz1OwfpULff9bQU/96i8qwt1zv39LrYCD8GzNizFObOxdhNAjYJLgAKpTiYnU
K+CTK+RtRKvBXGyW9CZDbJys06vTOxA+8m6oVAJMsfng4QVobqB9ZFFswvArKGCbdWNLuZfyW3y3
YDT4dLkRNXmAMq0weCObyxzgJg04D5b4XRo6LruAKeKb/RkE63jWMDjNBAsVexqoaY/oeTHCEtbr
Of8p1okDbV/z+T8oXz0YA9CynCYeTk73ZZOorvffTfKlKnBmoCpVvMXtunSFXglNaPkFzwiA0ezI
L7fmddIwIy/njT9hM0pi43WZnuUdQVlGFhzMON/zWV1Gh/FLIMtvM38jPJNE6nAdC+DC/hk8QSRU
j1miIuwAqS9NVtkYXzV53d4owUUzMzSUymOfR/n1iBxQ4zPOHTYghajM5/CmIM+5JYhVQhkkYiqL
a9xYk4KnYlj8xRbBV+nkjaRPCmAkAh1lgXXoSS4VyDn59fkKpBbAMY0bOiF+hjemPpg+58OCd9Ts
zKbB8Ao/mEo1NKue8TbYh+AiSs+JAlDRslhuaOl3jYCz5UKGGOoyStjv25RTkc2Wb3LIKY6CTMFg
sQUsRwfZmjXS2xKWFUQ5qsnWopb3g//S6JOrKPsIienfbzntLbRghWHGW9taH9z6/mNuGegYMjb+
Q9lyaoy7MAzTLHer/ACFqWBYXgA8+Uqhraxwt1fn0RYW21E7UP2zHseMqBko5jU2YzV6qdkb0fRF
+XS4Sg8XnszuttPc9qX+nPDPZrp+tR1eomly+ZVI8veCWXbAfIH4CcGF1XC9KehKtAvBvvfjcEGd
opNj3oJJ3o2IhyFCymxJ1t/aFrG3rm1RZ9a1x5zeulHo+TUvsLawiUxTIN7j3mZ+mK+sDo25W68D
QziQwu71q5/4vP1TGgyVYrrpXICDoJtebOLvzQdiiLLDkSEl2zPzk6p7pLIO2qeA9KQ2qnCgaOzr
lCF1MmWp/ztMk2BegAPCfIr7L4NLk5i4MSp3++2FsJRWG0TwsB8rt6eRtywxCHaB+amE28qvhFX6
Jy6SvjzqIPAja3VebJT6d3nv/kxBMyxRWeHpqB6RJHrjNolkKSabTthPLq+7m1IystMDkFONV/w5
zBG+BTSFi+o0uMPbqXRmuLaaBMLRtPcTlfmDGTQb33m8hPcY+UuElJTE3c7DGLA/3jjVYC/RzZo5
qpzDrUMPnck3iv1DwXnMNk7ciBNFPC3Bw+1CieITfKW3lKspOSUtItK4J7yrqL5s6A6aC7bRDHmO
ms0uf8Y7Xhj9WcO3H8ybGnqnO/QyGhemVzXwc5dlf/5fx0BFcbRJRlWM3XVnTsFZvQcPt9n83jIW
kUcgQCFzh9c/dPZE1V+hITgSXQIBsX5SlOrxIn8V2MmPna5QhZTwRlncOLmAqUvLqrWC3kp3zUI/
Cgc+9g/XbbBVNRc5OJpEfJ23OGfqysUm2C6fhqDwemZ9qx5scihQw8Ex7lLHlNYcykz6s9j4RYyQ
YxECe9P5wU7b35WGRI5uxW/JZWEDZSTvcXBWReIcQ0Dvx5lpGMRbdEpIOp42ZUc3/xvrCdZxeZCl
eD4LXramHdeozeX2EhYie7sAkVtErDcJ+KDIjahTk2WFjJadBsTsifzerj0YpIMmsE9aDiQxh7vl
Xc/jQAB3bP04/3CIy/5xrUHzTlz/TBaL9AaoDENC+1Ox5NxB/W+8LAD590u/KMY11nxkA43RPB67
TI5CCSf8Io6yIyjcem18YRhUZ5kp3WCGrm5fw+DeGwTHUpCY67RQjFxmELbRhu3BRG4SNEQ1WTqW
o8W5wR9dCTFE07fn2i4MYhfnxvr+Ig4aQvH3jhp57Ahn+aQ8WQgDgtDVrXghljG/a04LuCC+OYkO
dw7dmqQyjDiYjyhAde6Od95WpfMyHTmRNmy3sdgpkRqbkC9pIpJYMEHgkFlGI31G8UmJ9pEo0W7+
5wpIVLZEK27mCB93xejxhbdhhQJ/89G4y/rts49+aKAAown+3H7Ht0FdsfgRu+EpYpDnnSYAdHiY
WjGX9ta4TARYZY1xNAW0b66N4+eVsr886CKd9gmM0NxOyJTfHDbjRNpOkjGB6BwyQbL1fWi5KQNi
OJV7YbYBNY4cDa6qr9Wox7R7fzq9GoCs/Oj5Dz1RXkWQBgg4K67bY3c0QTJz+AumSIBKknnQcc5V
394/uCnQBbSSbmTIi2qZi+O/rMv8D7qrI5vDbrK09Id/guE66i62RdJgm17i67H1kXdzhFBOIII+
gkOhNqrKnmHFUMQg5cXmAAC8ZbHNMmv6+mbM798UER68hDQsDN82ewcKE/3tuzhRJWOKCwOW8NzA
sU7bVF0pNVysGkMEHwYTOuwWhIARqTedymg8U7c01N773JogVY1d7rdyh4EMECDhvt/h0irwIYWW
LDlr8eSbZAU76K+rL7ktT/xOSZdwmW13ML8+JZf/K0Mj6Js4xpOcClCKkya4iE+eqZbhafMH71Fq
8GrTsJxeWshh7SxvP/yuVGChgYnnSaFDF4YvulSSZOwO8myuE90n43sj6nUqvhMJAmmOy67aUsL4
tuMC28xFoF2ESydsvbxV3jc9usV2PO4JJ6MquqpA4ShdHuTJmJo6DrD1nWdfB1Bjuc+gvVVroNCz
6472YGNoN+QGxlh7t1HmuPOrIfTZu9WCK6v5D0QztKydtxXJmFJ+aPto/vI2Tg5JtXUpPw2QOWSk
cohTFj3LuokllECY1CVAOh6pnHCxqXqSyN0555FFXcnOXS42/h4ECtEiN+1nr4u8kBccYiQrE+JI
WvpDHiZKf4dAhNkpFq7COd/wvvTxjxiLZBtlVuBoKO2bE8VgkNhZmKkA+e3HpD+0odMYI4nYkOS6
0pq+dxtK+jBeBFNDxIdw9vf8EsBAO+VEy/kR/F5LjcNC+eAGiAekaXQjqj5wNeBAn1k15nyLUBJ1
GWgws3D271EMhDfwzgAIp7LGC6Rs4EoQZxAXsv31oZ8S75uEd+NZm1xd22PUO48gOcuOUAMu9cjK
MvWNSg/hozboZgA/N2BCgQFE+eOT27en3fi46BZEW7YZ2JqS/aj72wh5iDHK2FXeKrucGm/yN3YU
0X4SeZ7KpE0uVrCSqDJ4FYYjTpIHGVUMt0jbe8M7N53tcJq6TBgLQWAO7dVIYVuprd8T8jObDS2K
YoBrbOgPKB1A5xmYkFPEIw/h1yIlQz69SGRH8ppVnqDP5hOBo3WWOgQ0/UPa/VgbbAYkYwhj5mzi
9ID0pdyiStTWGiQu8ua1pHuvfgfnrvDSIvJFuUpdrQy853UBA2mOKxM1XxnKbjtMYT/iRq96WyUX
1E8MxTuB7XU6Dh5qxKcto52Be5THAiSqQQLRxJQuLnIMG4kY/1yKLLVSLIk+8x97tqK3bxNcmeOx
m/L2urHCWNV/tMNjOrVZIRo1/3xZKegcy02Axeb1cCxwDmbnvvF3ybssMQDT9WreBsrFowCDPmc5
1QnjQl6am6tGlrdu7lGNK1XblZfLD+XFiO0rbcmVVm2+3Y/HUOHCaSeEut7r5swwQuQxpD8Khm0O
mQJyVQCJ8Wqo+vQccBCkDolYDtwfng+oDxeuUQB6rD0pTEhCO7aqL3r90oVRhe4GxmvGiJTc+Kjf
FefnYfmAW9Hw9dHR6dgE8Vy/Uip/Yg8hfKjyqAvHyyGnye3PqxNo7AAQei4s4Kgv9197KyPkAs1C
XehcFLZ2h3EkDD1JI58FeQJBIxT6sEnTabk63z7IthAqc98jEZEANEEkIQbUn9zSch6C/guzJvsr
CoItZuUl4tnyj2BfN5u3Hkw3dwIzBQrl7cjIvt0vMWQdGxYd+unOcppiOVCmShGDbtUaNV5xmfEE
0eBWBD2+7rxtmtAd9pvNB14Zp/VaLV2RyD1xCQVPHNUOULjZzOTlbQjgrUkKhV84k9zYcGOUOhKR
JDIyKb/UMYfsUXtxawzEDlX3K0DD16wKX/XHd+7sovQ5YAWErf+9GFHFYxq/+k1l6Y6juexa+mnV
JG6oNwYZy00vErUcyjX4n0JTTxaoR437EtyzuqFpBsGKLiCwIwBwYM920yrM2FHdOW+6F8YFhahD
oiiQMsLyV6cSIXDKPCar3LqijLl6Rog2fhUqbCuFIrBwTOMui3EdOqsvTKNt6ORrg/xI6SeNNXFI
vBOYOT6DxqCC6QCoiWB4MGoooMEYby+eb5Dkh17aR9qq+t93x5lssCXGEVULq1dDJUkL9FDoViNl
b7fVrzi9DbzazZsaKiKQ1DNaQA7zmXMOt5WQiQzX2h1pGAaLWhzitO1YL+H4jAqVQw3Us8ng+mJd
9aC2YweWYdbxL38Ggfnw/QAg1xZr2xbpY9pZSbSV18JScCWqvDowHWkTrPpsMP4hzoAlbj8G6qVq
25MXuikBWjbI7Y2E1SdnIORnC4uDUF3OV3LHzAvWiGGSQTAccNnxm+6/NUCIleyILbfJHcqv/jU8
DGd3DTOdGrGLamJMe3f3ug2ycG0OiKlHsf1GJYxf3K1R+FDPHdaYP+L8NLVkLrQhpet+huov/u7q
xaazFzJ1Bg+xwIwypo2CzKHpv4t5EWCww9PB1qhsWgbMCAJucdkvLno+mhCQCyz39uebrjYeyVBA
+Ao/O7wbhkx4DJkpYxTfQzM6Ce4vTh2jFoW1/pIPnVe5Dnf4omNYOerJaRNMB4LnTd7Xi246a53V
jzgAmG7Xe1VDAptpFpWRJy0S2hTMiGkmXput1d629qsM6utWnfmskwh4Nsi9FXXbwRTwr+jlB7Zc
i1YDPPFaRWEiZfZahwrW9teTZgm5TsIhW2xMfDM0w/55ciXjk2TtG4AryV22AhIp/OtI1c6oYO0x
ZKummMy7lTixjRuDFXxRpgfguptAh2jOBckS5EsTFMDrhvvph027koRcNidOJYx+kyWABtZ4Mp8Q
PG+GO/1I9BsSNJRhlUrSeXh1XbxX5K6QvfiW024GETvapeFoQQuIYAJkap/KHqj6lUNVufHeETUt
F85C+8fTxjPPKJXEkrlLZlteTcxErhm0N1C98InRSOMoV+APWK9k6f8/bWOBKclEzhriSged+CdJ
feJIbT8qxrOzcYhQwuYd0DvAAa51k6a/TTxR7phES/5hVH0ecYBzRxkRxyxQhJTgn0KvOlPiUuGc
oUJSA1JLBLdVYv3lIRko1AQXUt/pqjtbma52LVbRRJk+LzFkKGax5z02TG41pyoR5XXcFdB3CQqx
0kjJjA3XELk4tmlSrERYfhF33KYJSYlBPMRrrRp/gXpvdN35wH07+Rl0NSFKcJh0rMQjsaBvi7iv
O3zqbP6Mr7p7SrP0WxwUZZxzkjoK6XK0tTJ8Cz7motrrWFJTQaMLgF5RlxE48qWntH34hZZ1kpKq
IHpnRxj+32BCpjY56R7Cd5SDGVycTA7qaCrZ7BEMRjeTpROcLDcxzXkHNQdMvQA/TWzaDmwVkAm4
YTJ0uKrT9qxOtqos2iQXKrzR7s2c+8YfyROE0cID8iK0Q4Yx8/sOyoBmieEIfgIJTjebFM6CkEf3
GLsqzkL8ij3op/kVxwdGKmnX1CS4OdlpOBUzdccJEHVEI9dQMt+65s6lSN1GYYIKAFqooOhUHipj
1O2p36mi818rM78SjCLlO/jKjsz6H23cAZnRwzeABfy+V8yEmSBPvlK48xSwCP7MY8m2zC6kMc2+
3b3y1BPm3gkbmtMj9Wa/B0CIe6/VwBPqXipC8qjFpvmSZBeTF7YYG/uplhdRfx7+7B124QgBVrae
u42fc6z0dbbyJNx0ScRQo8RXX0FxhzZxsMcDWXo65ojISkb/HqyAXgoRhdnIoAtm8U2Fo1ZoZf/u
YxZIOlD7c2+yN/BwNFoFmBNc5cnqlIE26eQ+kq68ECFTN9c1MjHRAizhKeB51Q3wlqKvFTLQ0YfZ
LIb1f4TQmw29vgE/DHvgpcFJbMFKIYS/QkC6UYGe/IoZxL/yPbsSaDIgINSJxSm5Z2ROpQgGWVjI
JvRLtfPvED4WbgEMLdotfFejksQpVbiac085TGLe65X10iGipQAyf/RVsj2dMaCMFqRe7iiJgXHE
V3k4iInuoRlPOrg7Uvckn8ffpEfhaazw5imjR8YRf5KWSWQqxEvK/m8NMcoTZnjRymCSOZfstr/2
LyKh0F8tsEu+ofEJ3yRoKSr5SYOq58aBy1Lx9Y+tfFmnR5aQH8l0behzlXoPiwSI+qyD8W3/U88t
ufNNUV5IbGJ1ASOFOlQmgoH1EQuLSypwlGKMQ2MOOicW/0N0adKSObDY/TwggQgrRl3b3Sl26Lf+
2OPS2LijW2AIkLEIcbZhQKYOMiGOekNzd4zWxNu9JB7UGKWQmLGfMq86y5tCt6tQ2qSBHZu5yAJ1
ZgY6Ju6CU/zNpOoj8/ztt3i7aePTIDyr5+hqO9+s3yL5usoN4wIk523e6Yl/S9bHzoE+E3VXEnf7
aDu3LpzAF19NpHi/dtnXK/19c4Jb2iVxCYr5/4UpRWenxC+JQMCUnZASWpx0IXg+l5/m+QSND5Ke
5bgN42emL8L0IMvTyjC2emp1JO91bz3YcLyxqNZjWirMBBhP8V5XI8INj9OrABU9IZZTDEwPiGth
BijbRXL+E/PJOuaT/wEg+Dx8pBl18i+gEu1zwImsJKOw9iXcoJ6MvwElk0Ds8rWDDuItpRApHZq4
eZ1U2+Ua6k4BJKGpeG7Rr4CORb6WDsL+Rh/Ik8FRt2OGsNTWQUMgqgXP9t54pxMyfHKgXtdUrMdp
GKQZosBZ6LtiTrOlAlmxHSl5FMU0yUaTdd+0DZf01GgKPjAQhCx5f06yBUebiPofG5a4ho+awhue
gvb64Ez5nDJfDC/PtO5JQumtiO8ELbtak4hSNL2lwJ3VvM82/OclUG7UPnwoXySl4MevpZhM5xcx
quTCjPmsCyB05qjq6XHcmskQred64jaPhePiBMtris4fuJPdGzxO3YNaPvb/6wYYWvq8bRS/mlfK
YZCccTvcNgDM0u3DvLV1sxJKq0S+bb13ONnFM8T+goEIPOQXQagBAazTfz+PS7FbPpDUEIdBqFEd
YPcgyj/1oYJDhsMmxp8YQuUwrUqXlAp+IgzMOOuJnQzpeagvfK+0v0e8XVWxs4wNBni7EXTqVqEp
SeMSnXTC/+GffqaYF6zTZt4leyOO4Bb52Gg5PmxxCHgwbW5r8baJUwKQr8laQPN+hilJu1Wj4Pv8
88nPaH2aCbDE7v5QU91YP36Y5OpcTPEneBgNNFUZ+5z+TytzA2kwFxJQSQqof4IY8HDWSb8OPD3f
O4gFYSRSW59ikTwRxc+6bqOJzpQrCkX5X9TOl9DE2fdFZoM5E7kcn1WqCleBFNpuocx29+gTZmk0
NlJEJMpXr0qneW9c8NoXh1hmTLCnsmHYjg8Wcod4SP6lb8YOQGXU1Mn44eQNCkhGGNA2jYxydSMF
COCkJORuM5caO8w88rm+t3mgKaxxDhNZA1194Ui/onUcaDgepZflI/4aCy/gi1N46KxxJZKIkpO4
laBet7zmc5Ju+ok9izdcOA7oX+COPutI1+XxhMbWKHoSwYxXSf/N7fzR1uCGS6oLuIXeq91oEyFn
jdomjDb5U+yPa8dgsfqWs4h3d37A83RRWTjQMU9juqoNtOGSqA6niPE+2o7gj/vJTfLVQCPlI1D4
ALZ5yn1n4znLMRprjmJD5KjI1WvsGCILUwzwkafYNj7zA9WCk3JUmn5me16W5M6pCw7I++CIT/mN
g/58mPvt/i6JURcaFSp0AG5A2KtSUhE0fhgRAPhNFVURAnaZRMD/TBjc7XKlo4djMCCqKo+xvTC6
zABMbHUYGnlsJ01k4zkR0fPAulRGPqP/J4fjAH7aI3QBG6RUHS/w2UDi0l0u75Q+nzwcNbM7Pdc5
6XyNpXmloj9G0zKVNosuDuybwByv54+x+2sTOUHXSXVKdefJUTz97k46Mn7MPZlARcvxAwmklOj2
PkxvMZq+tYS/vePMVC+FSsSIEcv6CZf1gSQb6QftNf/0AuReyYVfZM2nBEPmUcN94LfvlBEKEWAp
j2elALOC41pMnhJlHwSxr8OuKt4QYUsdf55Uc6vKUFgKmbkMURNIgaf0JHTeZh9i7CKJo3tpExBh
cof6GE48kZxNwNimBt3/LgadC887Z1yd9KlWoWuzgIr1ToadF5Ea3X6cBiF4yPcNrv34W3OXPR55
FxEw97xnLNXVgpug4Rneo3fXhBlLrx8V2noCZJ+Re/V7Z7TNb2YZTEaigimYtqdhZu61Kkj1VoYt
kYhq//hVWFM4qHQ3FlmFzAKbEm+C6AtN+vVcpdw4FXwqyfDBIO6AAOLhG1WhCoqr9au7CgPbE4HC
uhQhXVdL2jr3NCt4ZRJFQx5N40cM0Y88lAqd0B6Bb3mXp3WAF0T0cBa3vEjDRW+FlvrL2OIey4rC
5nxGxWk9j6exqiFI3EvK1L5bN52dGjieKQYXm3cCOr1gqs9xAIE9fnnDJ5t7Kg79EoKLH5NOia9F
0NG9mZpwsYBjBhF0sHCOUOLon+01QIIZlob8iNxZa4njzZls31VMvqTB1VTB2Gni6Y+Haeq8VUn6
TUvC7jSXIwqJo4hyaNXWxieeaDdRrcu+tzUubs10Ks8ZBAuecw5X8LJtDLpKr7o9uweoNT1waHbv
r7d4vPRM2XkAApva4VscpbbsEOs2pWO3sobJbQFfCgVnhtBeioOuug4Vh6Se7YIrfGKTTfLxKwxy
0Oz3SkYpBJl2cPPaU6rbSLxM06iNyAe9/iJS1NZc7wOyOsnLq5mxw0QAH18EeGhg1mRsyUFR2xpD
m2zY9A1d5aWuq8LTvrpMmiyijNedKK7V34mfnmsg+2SxnftW+8XoqfCM09Udnz7HY12I1ymXsPjP
GFShQ3qnvExBkDLywlyuYHSkmTCk5WbcpbXJf7FMeczJp1SILv0/uv/e/z/gcnXs+MHrbwcE1aEK
kQnUySmQ9cVqFjqZfWBMTGAvatRfnWA01v/pL1ejwuacWfb92GtrOt+HqmFFLIHnOF2iBH4XyOeY
d6C+OqiXeG8pQfbGKPZrAZm8svWA6ZjIqfU06UyKaNM4Qi5V84ROwPR+uGPXpHKbXnLlYOTGVNUu
M5Djm5YEjsXPDiMOq0W5lNH4JC+5nm0ryPE3lMeEbyIE/iQejSjVyyGSO0NbduUb3c/h+uScXvkE
GGX4+fqm5q1M8gMZzRh2mkOG+uUZW9wxpQzpnOOOGwm1vQP9bCq0TP54VRU0AfFx1GGOW0aeRxlP
c7RWGJFasjB1VPNpBJjIA0KJYeyWLZZ82hw108imCyQWl5jkvGsjxZKtbuyEwTt1lBXzsaQsRX0M
jl1fjPXOMgbDB1+E8rAjvkyrMzpVZ5JvzeMEwfOf7xLh/gsXuR0M0EkTp3vvt1PAsedS1YnLvreV
ZgoZEN1BFj3rHqUPak00oFUfax9uPoefsdVJYtYTCHI1QEung+Z3fcczmPsRVFP15pQxu+YElMTo
HZsP/l6LvILZoD/e/1eUtZrzYOAeRqo2BmoV98yaJGDJUvLVSdI6kg0FxflHUEKFfFUEXGsm9Mj5
zHIZxFqwBmKqVeJpboHCSwDtmkgDQ2ddWMPtNMKsitynnbu6FldSWh1JUMmBIgILQmihYaE/nx9o
XRK1A8klXM/Zj3NGfAeHWjMxspb4Pr6BEhjgRYwa5mHW60alEdTdxQXrHVaEMu1RJV2JIhnSLwsd
e1xeiN7hhwqRaxmW/e4xfuAqOtzODAwNupPmVa/9sU+PsPtC63l1aawkYVnR/BpUEhTBWqZ24Vgc
GUlCtKnn93L2Imen++3v+fYfqA8JSbF1YojxB4+VVnuWYj9HapwdiAPy8s5FwsrKtohIi83sRs9o
+hwyQx71cghInP/daCf3kyp4f/uGfB0gJnYqG/PjGi5FR0dJPOYaJgN+ftlG8dwINh5uVa8//86W
EYTkZecz5ooXzhnI62oSiBfxeZX7hIbY6bOQcYU5S4w43uT97oV9MJvjw29uY6Xo5cnSlehDQxe4
Ws9J+ZMRXFBmPfeORzYMicIw2xVVe2tinilWNCcwaMKn1zVJGrRaRfAXyT1QReK8lPxNfiTe2wVS
MCtPSAzWuyN2bgLq17XEV7FPgxa+GnWZUtKEdujhasNgu0CH8269r8y81VtrGUaLQ5P2rGC6Pu8h
TOOgpy1zWCG8gHfNxiMrteRbw3Vyes30HK2q31tE+osbvzbIhVAG13c6A9SgI5sTh4EetJWGTaGK
47DrWXAdMBOcO0rVGBnXGOsToC36agoGJOByddZ9ItcDgh1Exd9vCiz6+L4owYuW+3KhxlKKSZQR
oNhHYbZys/6kQa84hLZxMfN1x0wao2qL04WIboX3BOwFtuLimpmBzuizoiUiLS/AxZidoU5o5aFk
jdHvHPdyydkrDc2ih3tVwa82Xho2ffboPPLcJl41SeCScDgt1Qe5wZXj/PrRYowlLw9/teW7fGs3
czRcnloDUNAUNhjmgA3pS9t7oxZ9qQLWOPv+9iRJFB3KvgDjtqRFnn/+1Y0G01+QeVgL+GVtM/MR
zoJn0tww0yWSXnxlS4+1x8Qo6WjNkpagb7KLSlcRuIcmZuL2J5Hrs0laZIHzGuvx9OemPCkUCekD
7C9O8H95Qq5OloFQRyRDpzjqNQoqdOLMaC/7MA/JoM34ZjROs3GVSls3cqqsI5yAkyMHgmjH6XwC
lrazc6wueRaPlTSwzmQdZ1R+tiFB+CTcwxKB1VidxVVacjMDXYNbaNKbiVWg0wmZW8GP6KKG0c5o
+oAbGE2sadIqCiI3fEb7JY4vXb8AdwkcYwlJFnKh6Z6Mm0UBDaH1ZxV+XPGalFypx0iAUXuV+7bt
7utYdatGDYNt5MRHg1SEgApG29iFAn5W/qkadZmGH/oy8AfKJ+Kbv9fhqMmvb15Yq9kFIwZ3/QUu
awf+8YftIKKJbPa/QXcmHOMK3qMmNtqt2KrjWofL0CbUyZTZ34lYznovDD00fh0pQdkU+pb6z6yD
dYVUK88I57Q44CwdfPcHt4OGowOWiaias+kVb0a0NlHrRI5bBO/eWmMCHeLXQTJ9DtXY0fZUm1dO
ofbqSi3PTHLWtsLrq4BZlvklHxiGEurCCHIsIi85r9nVyRncpFTD5qy9H6ftElzEGPpDKDA1LIz3
6X8Oudi90gJQsl4WWrzVlxLsX0mv4i0gDN+lUObQQJsBUuy3w1R2OniabN3jXxI36eEeGs/FQOT3
6F2fTlDRu/IHJY/IFtLsu2MyhhtK8CSEtEva+z9BCBoWlp6m8ZJgCUd1AW+c4WYIewNRlAku3mCh
iP/ygxsZeC0ZuSBZKQBAloyutYXOQHU5j2cmRtvBuQxBD5KctD2kQA23XWedRz2Xe1A1HMs8gSic
tCgI26HNyAYOJ2a82Jsq7uI/fMEuF9lirsDmWvX+SCQXe05rIPICV6OVhWjKyNrY+1oDDVvVyjfi
aAT6Y3EXCh8ZfnVL8vLR3+dYBuO8DVIZgdn1h1eKcw94kE0G4vjPR2Qu9MQFMCxaanIUX7xbLI+e
yhBxGrF6b8/EtPDGi6H59hydbw3Ekio5n15kJX6GUJT++KacgfdiUXxYOXz5K1R0WEmm4QyoCgqX
6/tcy29TjfncwcPsqVhhegQkySpHR/UmUamW25JhHc/J0Kev2QHVtuW/fGiiQRJGme2v1CoSLtU5
k03sv5gqE5yG0WuhH2IPzoV4Zjc7PKHOXFA7jepEW3Y1Aa9jWKrMM6DdD0KxW9cQ5n0e1SeD3ucS
E/HiD2cPPzkc9hNCF0D3wSBw0qMnGTMfQuM1IWJh3vzlAqiM1qoDS334PS2yES1vpLGtjIrN8A3h
1y4ru7RK7JMgNMM2MW3P+T9vumNezrfl1IuE6tCboO4FPn8xoId+9E/MovpcyQHxUvCVZY4RplHH
b+6YMrSa5YwKs0a0BNqgZZHDBZTRqqxW83OqOs7bW7fn6g7iPNhw8bSjVXhsCYYPKv7vRM2G3tyx
JdUgpt8YiliD+PF4vbL02Q0lC5BAbb4ClPVmLKB3wXiyZIIUk81PFgndQaFukei9DQJKJJ2gz/00
PUyPyhDEItAAHioP8lW/bW7jBsf+Lllp7ikyHpdWRrTiUcKWPfeB/X0X3ChV1ioND4GR8PQOFWIx
Zd+UWnmfg6q7BAqB5nnBCsNc7v+zhVfC0Mgyc/ILOUGlK1FlRj8E0EV9XMLSULCLTw6Oq8kF77d+
ekp8tIeehv8I14ASKMk0x02whfzYEph8Gbzh+EyZCJubvjL38fmL7tZfESnpLZ14IAFk4pJ0o4Jq
eDWLossPc8hOAvkSWiVJB5NQI8+AR/bmomUE3uda8Sf82rtrADPm6jifjGiYet4IE9re1k3Imvde
8WnVa8JINv6kvkPniKjposeeKSg3G5bbDeQdJ69eTM1MORmud408ReayZgSfQizUZVFqBnZHfIFl
0Xz1BiOvjD2nJqiTz5TNbaHsP2d6tykbpaIb+UHu3wy+OvimlfskxXZUt7SWIb2aZf8hzOXLQ5kW
344CQ4PhCbGL0ksVQJrM02iLSAzuqMqsiBFja6fyq466QdpxaliNsf5J09uHjhnRcKBt7EulpXz+
JUIYU2mgiux757MAPRb4B4P9Q7PvNqO4OkZ08dOhfjQHedgg4AJRL+PvbCKPJvdppKvd2wX+pZNZ
qB/ZQqNm9KzX06S4wMf0wcW3/GNDY9rsq8vobqgsd0gjQwAZ5Er5PJGNuxq7R5JorVsqGrhzTnM0
xhNoGEw4mULWRBsPt1/j+6wmxA0sVmMMfGeH33H2y7kcgif8UyhqWk17MZvujbX/bVlqZUFZ44y0
RZjZcULtVkYZ4tUZlHUK83+INRGZ52KLJsOt+iRu1czGigP1TL3dmPYPCcaDVOrYyb9L8K3VHG2h
Hd1fXlUtsN6uPGD+qHTzg8f9/5Cp6682D3sj6Gmek1Op3RkdqvNEZSgFdrPlEpGZ7GohPOIEpQq8
FagAoeyHZ5tBdK7CzCQd1AL4M+6rLUQDMrzR6eazm0IFvffmAUrLUMnuxL3gLX+Ws1Buk/P9YGIR
vjoCyUO7EWHCdaGJYF6hQJxNsy7ruNCUNAMMRY4z6le1aYQuq1fb4w5Xkq99UHbhZ9/NmCwHkpf2
/sgy0MVQzV0LXO0IAWxUaPwS/ZJIqSRrdNLWQPY+D7i1OXYSDJYsfcbduT0GEKCdKgHEOY303VPX
7oqRUx9pvMjjzrHRFk7DWBKQGYQwL/Qdb4UaCqtaW3tHbnvHn96f/z7eMdZak8vZxhGvjPzigtB8
m2qveb1F+5UEF1nDBZ/mLFFX+xOFYe+sHAwQGeFhJNE0BepPtus00ce4msGd8eSqfvelCQ13kE6l
s6Dcq4sCagZg/G9MRaj+GIUPeHlKKsmJtU6tlgltCqZjslpyoibTffVsZ575YhlWGW8E8dxi+pho
qvqv/XI4xWHeM5VL17bmEQrSc6AnQe5LBZHls1Iw5ZNK3JpfXeS9J7wocmcr4MUWQJWoAeWhze/g
Y9YZbIaKq9J74WBhg9nSYCmaov0RzddBOsdL/78guqsQSmT3XQdNIiTRXGGiFGGfAurxMo475R7W
Sg97RMsFCZNhvkuyG1xrlrXG7TfSf5Bo6Xa2llt5cEFR3wFaHxlc08LCP23NPDfOkg36LV2t7tcD
cg6S322SUOeBqEifnQg8DIP6xR3DPuT+iW15xGGcXkL7+MdByms3ClFeLo5RNMwZGs3ZSoCINIf4
s9VJs6NnlyE6eHwYQ0+7JB8lDBUPLv6EuNWiBF/Lr7+JqyIMJc+6j5vYPmsoZswBMgW4rJD1ymzJ
7/oWYIW2b7u1wWClb0NVMq6GsRXqwbMOu6GOgLj+A1csuIsQbVD+XgZ/v8ieixfN8AZgoj/tqo11
sNQveRRubPz8ax5XfDJ91llnUGvQtTsY6ll/cpTR8bBfeTVDSWQWadvtwdh6cByj7/TskVEtvCU6
Z92Ls1EOTQXAKaxpWMLuKoaCKRHPFERkP+5In/qaS6sl/r6iQFEutDvv/ftGrhKGBSv31rbUOAuf
nWL2wuNxeZerqUqhtalr3m5J80o6dc/P8PvNm4Z4ixW1HVRaJPUGLgFgs+BeOLI7mkXzAiaioTQ8
NxjqOq5nWmkca68tT769hsTHdOpUYz5n6sTpiM5f7Y9Y7iKTroWEtj+zqMjyNWclCYdVDggOlEzl
Y5H2eV5ukCjjaTTiJVQhobbwh3+KGfizWPf3MCkrup1jf7UsRUmJ1w0mKStsOawN1nnnIF/TFD4+
yE1IxiXfuTt6Z7YuuptA+Gfqoqxfp3JBoINgcs67NH0er/qF4TyGs+J7/VHp98wTzwlZCMa8gOzB
GXcVWsOqgC8TyriFbDhDPOniYwp1zDUAZesJQ+soeDTVPwLc9Hi0c90qnO//txFwo0/HDoQe9Ovu
R8oOmAghJ1gR92ve/icLTj5WEMd7MZXD1SXFzyHRbY7cjBLWXQFLuXC/tT7l2eSK1KGyFd+w9jE2
SJ/RHM5duxzhTtzZVQfINZpEYHORT/b4qh+nY0s/eIF/rCouWFzXojd8VcypS7Nc7wmsiJ7Mw2Rg
LeX7+sjA0nANjvgD4sJfT6+vscbbhnfGV1MjB7YSfGjwQjgkNsH48QzBdZRXKI6CT/DJJQ7K0ESP
yF05f4jKw7eyBgCpe6YzMss0yc1cqsKm4qlUwAcG1DVAC6vd814BDvd3P0xc97YtQj/TXZ0X072P
TRvHaR7HjNLaOVpfBPKWn+BuymsZW5Ou1lXePQJJOyzuaRjS6DCPGFkxuZKmN9lcFKqpAtmDIGjb
zwlQGXhOhpTDynXHSr25zNAeca++EbV1hdxoYi318WfL3qsj+8pUJcpYu4FatTS8rsnqxdTN/8Fq
6gRR9LOaj/ylod9Cg7hC97STjHcTimeet9vAK3W7c2siseiBRaUHp8dihFtwWOB/ffM1R38PSREw
OyYnIlSGEvOyaKxqFPrt7oWMS4Ymg8jNwsydZgcCVSipPKy0ZNNwKeS+rCfswZ7pA/WAPKCpfUXQ
s8unTE1XEbN/gNt0cBkskeoU5SadFNIYAXSAWI/vCeWtOav4Xy0X8K5lfnpW5I0ZnuktK14Y3Jdu
LMWsaBpSbpmn8MvnPOtUzw5+Yp90AbbZK0YSJ2Zxay6mSp/tMu++fqHsMtP0bo0NtTYjp4Kh1syx
tpEtFRITaP1QZ5+SMhvItxE94vz9MjZXiS0hPMM/ohaNRC5YVX1tVsqTTB0TFCbnWu8mi7SV67zJ
W8AAwdu+dqVks5u0lQz4OVUBdmv1x6T7eTTedAn6l4/nj3YsyxESqGWlRKgp8DQI/2yo52VvyAYa
UIEXdEm9to5NKUyoWh3kO7D8GoKNPTqJZBS36bzolBKZt7C51fWRvSn7Ia23Hm/EkUi1mS5CLDAn
y/wujRfiTXVKj7E6cF5dv5H1aMi+i9f3TWrPFu38zlPj8PWsWIk30T/ggBELjhHv4jYZ7UPxblIN
zzu9a19sG0GJ5SK8yd0led2DZt1eznAGD53w2SfCZeTMI6L1ijNLYKULCLKyfAvMN4PErAv2wBCa
QDWceXubMJkv1oCT0EPhEDHV7UtutcRb9s6C4pOFOfEqQRPCv5kC1Ks0t/BIl3DqQn3+psS+wl8X
r5+aQyqNf6QmLLAXI840CwmSpKp3DTejAcIqUOL7/kN5Ie0TfnGmBpCBwAwNNB4K7RSCRd+1UI8q
1jlAUCRqHQIPzMaQDmdYareXcZS0sQ868ktls3XyMS1RfL+uLOvnI6UUkOL8FyPwo1fI5PG+kE5h
cb+4gj6cYDTMEc9vpX7UzzzX5aOD7yfwumutFqNTLHOgAKigWu5DeCVjndO+HgADzBLH2KVMjWlA
MMe7UQqTRhRH+jN92iPJa91mThu+OrlcJKiaFbeO8UWtb+V3bZ0H7jGvvmBdAFCIikFoPrSTCxPh
cKgyC14W4QEPDLHKGrz0irUuITNp1XLK4MomxkvKWrsGmeu8QVYXvgjB3iJa//+AzV3SwT2fsCuo
jlu1wQ8SycTIspHmeO1N34TQu8hTkK27EoHzeG+Muv2hh+dz6dDCpKggP9JV1T0PKmcNrQbIHE1F
lXvgBNWvb8bp1HvDClyDZb2j+xasOTjMME6uFpAxmZw/EJ+aOqodsmqBQb9wkRyDx+as8Kk/hyRU
ZbR9mYB4Vo70w1FmRddl7L8XSvbgljtw4ojl7lZWADnvPolkZ5lvl+gdCbTiCt7H7YKGCdwjxMdd
TfuMDuwpPzFvJzhkKWZSiid5nXzT+LO0jugSCMZ99h9lxZxSUWvzf22seStcDUxGskHHssKPDKAB
qOl+Ul1pFZYGWrRY9Sw4TGe5uxMZngnnV3zccjyjSNHrrOmKyFn88Dysu7FarluWpdKoVMytl1gA
KdN8YLYMpg7invCR0NWx+SYPbY4e725tHV6Wr1yztCv2/fMW+JqImMEV2f8rDSjunx8fVzZj3APV
0bQizYkFg14sWqGRW4oeteKecua97Ldqejnbpyasybbxwm3Av6sEzjVaHo4B0/KB9pYfPPQBacZn
xh1IzQnofAXKNoAbkVlDmk3HMdIVQ51ZSDyiK6naq5Nj2Lbi+MFfzeAWjqC6DQJ6+KI/NfKXLaF4
qpGaScgMMsA0ATFgucEIF4yLz47xFpEKKi4M/cm882jg11gYW7B7Goa5ta9zt99FzAwJoFauoXEk
Dsbgcza0AKBCXdhH3fZEQWthZoR3lIaW48WUVMk0e9hjBAhfBok/EamsE5h+X2R/O+jcWR2C+93k
j3LLLb6XkkHtnO0LEVM3Syb8lPiDHVnsx3eXNNijIcClhzH3UhSZRQuLPHj6kSb236hnH2TIGk3J
FzVreKStwELaooO3qZZARgKdZBQV/642T7w8BmQve6/n5YeBMXOnbzY1MrhYW/FKrwGxhEQG5BCn
oHuPngQGzgYwVo7SO69vKZ+hvu/nddcukkraj1ehZFbIUiCMhetO8Ma8hm8KGjC7esM1shWF/ReS
eGKJlimyMHwmkm98997xQjwEEjsoyU/o/T9zF2K+up2LcdfimEIb0tp+AZSDHQz73Ie03ihGSrhS
g9Z5sXbb/AuaS8FNvfMhqwzH8pEX3m3fG0beci9e6anomMZG5vjUcwNNukZhIILRD/G7yu3YCXbo
NWIngcKP9om/OzT5xDXMV+H5oVCGe3W+PEojuTieN4fHQ+sCkTqdH9B5QmXzTA+85fr9rDAGWLz0
EDDQW0DdclY6Lu4pvibCRPEUIcmk0INflJsDuDhMcnsb7+n8ULWVUCEMicX+CfsOiP2+2tjKXujM
1z/e4bV44AHcebcRkchLKL6ajRVPBEAcjJDc+wLCrKgjDXUzoAp1OeMuZRqfTletHJxqd+H9XhNP
VMcGkBoX4yUeg3DVTidN3SiFz3/HwNqpMh8CN4hNgFamRdsfQLyZe9rGCE9YQnNJ6H/2Kf2evY05
YbARg4UrjFVc0Xr3aiOqbP6LOMeisnHVc6NDj5SWsqPM6DJKOkGvhwZaV9GfcYTdcv96WEdEsenS
bD8EQGxLMTT4tHghRU6zwlowLcc8GvpMDCrMwLee7VXNYyEE/c50VAfyFfvedoOUdpfisIxeaRcQ
ziksmDsLaC2icwPqXOmeq6kTgMt3VNGhPdQWx9flt8PeaRWGhExzF9l4lL3UREokbZrRL0rzGvnl
W/bNEBJQeHSc8TFYiSjkjRgJ7R40NAytCJdbqwwrJooGU2OK7nhNWoCVA+9FBWkPosFoXkgPQmSc
PIlZcan9CjSVsbhxfjybUMOVff74CWDZAxvrXXjsUEtvfgDxd0WK1pVqUNDKe23el1EAySEYxYoR
iJcNneBl0HRfepOlC+tv/W1L66XHImdNM0V8JW1Zb7Z0uZtVGUovA3fihIcUkn9RXSmkyb9dbvPK
0oB+dpto6B1VgiOeC0MOMBwDU2eQ76ALUH0PUrHN+rD36XBBfNYbzJUEps+3G5bOgyFHNe35SuHf
RuuJsjhoBRf4i+ISz5NdU2wsmCnK76nngg2gGGeVIzUx3/6ppkZz+oqwcx7tx5uQPMPsj4yK9JOO
o/NwgICq44GmUGm4jhFUpzVCb0LIVAC+HtAI8PH1vINdPdmE7retteAjaRpXUUqhsUd1iWkRjr2G
BoaktV6FpgaRZbFpJAXcayqFZ9CBZwWT2Tw0XU64I8hiRQzzd1c9eN5insmkHSw9bI1mb65GnUo5
uYEj9Qb9HHxaw0+yZXG+9kfYmPVcqYZcInAAY2SpemzJvB7eGIxCzBCxiHYsnEcq4VLEytNPtntd
ndcz44TAKfd1uwsE8QAU1RZUdXs1pR0KRFGjGfWq4hduWQAGUbW18aA6nZXoymxAh1e5A/4Ap8Zt
26rwt02Nfp9pe6IaLwkTVktk0AHVvpGwst1MErF8hTBa+3R8hPvmTfVs3ZvSmjhGawdPu/jy046Z
10NlJ9AfWIEx5xndgZ3rXwa3rYQOcu9TaTEyRaxyaNYLa1PlrrLCj5uRN1XcpT79oHVz6bhSKhBF
Usq8vLSgOHMi61FW/bwuHi48SJe/5G5JIfZyi9R/doBg7VvXEK8Yka3sWoqjGR+iAHk6NLO8I4Eb
4R3aKtNFQE/lXZhNiMfdkEpMUKUN7vsSRexdQAuyqTqo4832nDBRYVvmMBnOkeyQjHvqohzjQWYV
vsgvjHVgLMa8MU+21aF0Ce4rZLmYtQ/TgREwg5M+oKWPgjItVWqerJfnktuevE4i7xhB8QRjg4X7
F/rKNFXLQM0dzcq1Do0FG2dGoTQkCNMovJZGnmQr2ggAK2Xyx9VSfeJbdvc9vTQNJXXSkhEinIOa
bqtjgaVzfYYIR3IzZ34hJpZDvijs+fQNUvnhbRlw/AztJGx2w92DzaKQMoG0meehKnfB0PmWBKlS
Vb47nfwToCgDcGVzxi6mDTnkj4OQVSu509ftpe2XQeel6B/LIbf0Dgv5LSAB0LcvFr8nKXS8wrOb
MJnepCjm41VA3bNsRsfqjjL7yuMLlsjZyFuGyJgQ6BcYNWtKSvvZ2pHnuExAOW2Zq73xdQa/bEaa
bAZtMXJfRM8OxABfhImU1jpkkO/CIhplyQj6o7/JXCfdn9TERIORR3wKKSRoqcfS4SnCt1jKyIb4
L/KY1HB+uUAJWbwTTIG2M09mYLR75VurXXiuuHvW+SKKHzot7RuUDT7POAHpPb9yj6nO/yrLoLSy
gRbJDoXJkoSVIJqZWvYYgwm27Ly6R5M4IBBRXD0NBcymvYUS2vAKEecenLcrbszRCfLZvzdGZjBY
eoTUH6glVHLamQMUBTI4k3xRS7DRHqiQzr1qDWKGhz7lkKBOa+jnUlhVW5bdd1HTabAKb8eTQtn7
CeSfzTJG1U8voZduhq6oX4xsGKZXUk5Q0NdDQ3ckIWdyDXC6F04rzwj8qqU7pcjn2pe0VGpeZ2mT
m5+y7NrvcuAJzoubEBe9Sfe7MLlF9b+zqVmrA+UkSCv2Wv46jQ09bVN3fOuutL26H0FiGU5p7ZX6
njkXBu2U80svvtQrk/imsxNp5jFF3z4Rq+514XTeNojDDC7StMDfXLCa+wV8VxFIz2bMpVRfADww
WoNVboi9wF7zEMpzXy97xBp3Xsg4nNs1mf7ieL8yNfCYbSza53iYnMptidlo5DewdCDVPeKeowO+
M72qkJxhIwAjRS17onHJiMQRRu1lMvddGBGYZBEpmlwsqnKAe4QHlkYzRni3TYRHJTCemNm9N6Jv
fpKT/UoVMqcPCqQfwZa75Y6FDYf5yT6J7YTuFqixn36BTcm+wpS4b8Mq/m6MXGXd7KqDAaiJOBt8
z5kjpbGeoOvs/fwUMK5Cpqs6g1JJf3gly2MsrJgYoK+0KgzQnnKoAOsuABO49lRkr34mvZDwZ9lx
UKGpU0/a3sfvke7wRnnmk0HuTnRU6tL/73JgkpWGlve4gJEDkdKllJ49GSBLQ6XoKQR0HJqLAkzi
b5ecXmhySTRui0dGmrEgi/im1Yp0K70SsxnADjmsjS06cUCmycdtekaYfs+bbTqzHBuwZDWvlusF
kRDl3jw8Kd9gllArSIaoLd0h75NblDit1fWnwYbJPKjiGUingP1FyxFAmtxNhGSlnVmn7V2EJhBL
RuTjE4YHNSUocpAt/ZAQYTUhm2CcTofeYMTZR2v1sGl1UeSXBWTCKl52go5UzjSFg/mlrTilNsCp
80bf81VFIIXRZGVsYTYzbocXhNm5HWieoec+hIFITha2bxecLQjF/BwZojvfyNwWiOJTMKpkLhKE
PsYFXGGn2jtUMQfCrYUDcCwQyx1QhjTp6+MZ0agc1HEvUsJQZbuIzh80PGn2Vm4xN4s4gJsNsEvk
cTPzBC3TWVGZvl0y1C4jqpj/hR7x+wYwiQGxTxoEq01olFBKwiZFHaU/yHa/arq646D2gApmahHH
SiH7XvnZkmuFcK3Le95VNiVe/y15gHQGZVN7V7CrIkGv95A9jObc46nru1cm71JeSnU60VHdv2SB
+cNuiS2zyxlMUixqh8A30DPB57JBvggtTWFM/1pRF8JuUIvY/HWXh/itVIU4vcwD1sMGikdm2MkS
eqP5tr8qwqHwVUsSGpOc2o2XWg7cAsThGk371W9rr5q+EYCOFkwwyXtwIH3VqwjrvMiucgVKRNJn
aeOfvtWO0t3vDT+i4tnRKbKZtPYTb4IZb5qyZ7VVxtf1M9HcG9/jGqHSUM0CpMpKcIc9ahX+hCPl
Q/ltQlUIRp1DbMOTZTXt9dtJWdc5/vJ4OYC4DIyVRxd03A0FVAh5O/rYtTaVOSXfzuv7dXfmcd4j
mYBXUrSY1Bh0GpKIQAvP55QZgHqnKrIAfXhIDF1PGofDQkfD2sIDLoR9vLvEGskCVb3vrTixEcQR
grSis5htHANEhOW6sCVPB+IysgpWZSwaRwFMVO45ztvdqMbF66/K/T0NHyKrXuuiH4YVjj2kXJN7
/gDbhkO1n5mBoLDVHzVMRIcsr66rNMzA9a20FpXGo/l5d0tGSvLBcnerS4YiG5wq7sh9a12DjrXU
rC/7gm6/mjVQqe6RLZc4w4cFV5MkUy8VkkcgmknHVD5+pTvGOYcIeWM02mEFoU/c09wIQ2q75+Ys
NPou6xuZSddNChIDEVlAxD0QQVnmc8P5HTmd1O2HbIIqb8cgXboo+e4HCQ5KtlsJaLvoopgX/Bww
DNSdkJze5eixhP29dHxBaCbTf9WNvC3iBdGn30EfyNZZ2qHPhjH9wLbecX6h7Et6Uww1mIqqBXge
nusVGG8EOCQuCT3l/04fiV/pDyFF3DtWsIDVuAXpVbt60t/QUZqhzSCHxNnjotv6bmSXoapM9NB3
vVVKc3vY6+SIw1uBxCK9+9ZziQJxmsFRCsUADvkBlpIso/E+d5RmBc6/WvPIzsA/J3KleAK6mp/I
0TeDR1Q7OMyzIxifFT43dqlnavElQZ3wTCxclVj9UFLQIXJVrH0C2LklXuQqpLEAdQSEnl0XiNvt
RXIKjDpSYj5uqHqH4RvA9Pqw2TrHHzS+kFGgcIdCp7nu4BlvaqO+iU/vTtiKpjT6Frisyg60h6u/
2kXCxgZPYwGazQ9N4FiW0DJmd+2ZkgHagEfPk4/EBws+1+XL1KQo0t5nrDLqr4kSZqgMCcL/J/BF
Yx+DwZToQNqkLiBP389/tLCcMQfet8MKYvOA7lojY1NH3p6LjxTP0fXbTaGZy07hC7nPj5kKP6fi
NX1xXJZL99/OQOhHK7e0BqwDe9EJLWoSSxj3bEryVebN3JwfuC6jWHKC1+SRl1TYmq0lIdu93Vh/
hWfgzHiOc70FVq9ix0gipk+A8i9wTLm95+rgY7jz4Hk3CIFiMThBqC8At0/nnjZwtDz+zzQ5SJLy
kQS4QQITFDUJ98IRk35VCl80lyw65XemTMWB9521Q8e1qwrsnVfZxzmpE6x4J1HZpMcRp2EG7Whm
trCtJ/fYudzGQk1fForSbs+7rQPXBDv1MZ55U+u1wVSzpe+0W+2JJjgDs8QDZZnTqfxWruoIrLkP
bK9dvAA96jZEGBYS5d4PEjo0zxloX5tqn1zcuGM0f1ghjFvGMuZXl2dvzyP7ilsXDcqwknRCHwLE
eFUOgMCUY9Fe0n1vMCoJN/3VWtOLdNAFlGj2ImcrmxdBJ2glcEzdkkZ/M85HdC1YAuTO0Sq7qd2a
bguJCpZelPV9wKFM4LWjGzWy9fOn88CPYRDIdHabW/Yq3BTKbTz0CzmacXiVgSzcGWwDzKgQWFLf
f9j7QzboI2+BCjjyjf3ZifYupJVqMi+kQ4yo2slbsE8y0JPLlgl0uQoStXpcVLnG1xSTxTcNXhqR
k6d0XY3T9wuNQdTyjuOfFcRz7kHZWWIYCeQMqson2VkAzJ3yem6/IQLh5vBNKuGkiLZ0aIDaVE6L
/m0hcTmWuLODMXRgjsCGdefBd1/s1Zg1JoljOu1pZAYHbA2fl6x8gT0oHlZ5VghXa7MnTMIiK2Xh
LveiajPj8BIUluEF9IZOx7LTDNGorUuDdpEFSSH8lZp5V9trc8ZoYQjihvln55RK5fgj8LOVVyQf
f8VCrGk0PvnrypEHuV0u8J/XKXkOUkOOfZ0blBxNb+S6wPoC7jlbDXl/DUVQS5fW/BJ8E4BZeFpn
98Tvojks5bRWzfq+YgRm2fUZ7cvGDpAb+bQ+nuwt6TLg4Q7DxGU41Zv4OfLnRcDG4xbFQVgI2xOp
fX4/POT78P+far1NfcwPKuOD10aUuS7tj7teCanYXFAIXwIJ34mpOO2+dkdhYvtaNTonl4ff2Rst
Kjm/efL8eoOjgB1CW92kUjAY4I7JfLx4/Fa31xWddug5qJRUT6DAULDDqSLM9DW7EODXwd6h/p9T
yRVa3X6qEN8BndqkbJmv0ilBdqXBX0C39B7VKMOjYU8f8i+/W6iLAlx44+l0oay8UydJWlXEAy8x
QpO3kSPi8+HQW1/LSjRaA18MHiqWprr+UUJV+vWP/2RQwpG86YH3NTbE8pMlMpvV1RYIHa0GBtXC
xgnx1h6OSIUU8tiBPmQNCkwDwM8CPI2/9dTWoctV2SsZ9oUpsruxmrFvz3sj6Y2ZXwaQX3GXBVEv
biQVPfpKgKHiZedrRwiwmI7vGdv9afhsflisAl1HHz/S4CVgSvAG3bQ9naNOsswIl+tSgAurOEHM
mEDFgVNqemqc1t3b/RTYQ/mtCy7lkYMsloJeA8MxwOo8lDU/NugNrUHckRhrJ2oxum8QjmOYWRn1
R1SYnPMZn8zFFjAkr7F4Mzoo/dHntfb6i/fXVya1prYHS28tvzLnt0SVocEW8CQSYJG0r4abFqOd
EwGFQ8mA1f4mqiUyw2jZGdzdRz4N/AwPjxriOSInQ6pdn5aZPlNX4YFUqJeUOm+4CTcK0Wl7ulC6
U9wyfvzS69l04QUPS6TS/U3YVb2Llzf8VJEPwp4VMe/wEmlwSlUCXal5fx+0RDpaKLnWFOsgeEpG
7CaaQV2QI+2fDtAxTQKmGS+EofrSVBk7jo1CkWTcBIEfqjbUCm2SCAZDE4ySefH6zlUVLIJXTNji
7AAaGvJ9RM97rsvverJXPlL9niF/hUXZE7SRLp+4wszdpxssWR3pRcOviT5pCyJUu5jyZFC8nzEH
U9EsyR732pfZZLO6dLRYeq1q027bhJOHYg4XDRV9tXG1Rd1hV0dFg45kncMyyD6lh2Ze1FFHNxcz
/gCoDJCviq2NTLdirFZrnVK44+RFUCECiQLAoKcn7LQzt1NNDhwKY0I+VEOfkpzt0/cjBhxaMZVW
CvmRMbh4Pa6AQGFRD4qpQS29iF1bUA3XxxywJVsQKgn8mvv1AJk5YOh2gup4ZAmB83zJVk6SMUok
FXWINKVPBZ13TZLGr287MgdESv/mCQUNhhwnvWg1V2Ln3k5Pe6NQQ47jJmtAJzTmEpyCNKvHmk69
0uHzbCe1rT/WMfJ9EEkQxzro39NwLH2STUhAm5kLr8M/n18nv1EamtmmgRh+T2pVz06/io9pkvo0
wkboLq7PyBjfeCQvVyu1UXDwXtELv00+nJ3opNT/Hbo5bAQh9fZFd6yYVFrnkluF0ef+nPidq2mQ
tdP6e09DS2wrZ9lQssc4vIvFUQDRGgyssbd03344CeDnO08lf+rXGVxXCo2qKWzRENS4d0nxuBYH
Iy0ImSlAfrc7E4X35NIpsUcz1s/VAV9OyHKjNmZFA3DNW+pAeUZZ9XU9S5G7+w5ZC+8uiW9HZeTi
3FBANWiLAaYc4XF9DRNtb3LpfYzxBg7+AUvWAl6G2gZDQ4eyZ6wSVjfFrRyHoJCDDGVUCX9/HlvW
6rDU1luIqLBFCZZclmk4F/7BTOVLBE6j9MdVcL3SybUqR2EpVU9aYbHQqH3Z3/oySwybVlYoo0yt
lPD8CxbuZfnvAbKviUXCdUBb+ohGByfQt1q+60tfJdhFKAQ2CW1CbEpvLk085XhQU0DDHy5IAel8
LxUZDZiRdyYuvtgBMRKE1VVTjV39fNx4kjrF8a836aZJxEAa2SlH4WablWIO0S89+ixrup84xtUp
6af727jTB4/1PM/K8GfvJxELthvSxGD8m1UHAK9gyNuZbaJanDbznG7LoDRYoFMAxUu2B9bfqQay
ZoftUm0yqGp281ypWnaUe9j/hiOaidZ6S5YnVTmpmRC6GcPXbPy4jwwxzNihvgrevQkyBxOFgMJG
e2c9eL3suaKNdFfVMpnhHlelN8ascewxSOx7pIn7HJ/73sk1tobOhc4Gez1bY4rdKdEpGeJuNbgK
oJdhpRdi/U1PPT8ra+oE0FhukPMzOl+VPbYRdKXvavEGR+6Z4z0PxE6Nv59nZqOBr5VgR5+9sg+I
iYVWXQLAT2BhAkE/0tQW0hKZ1bMafNLuOVbNuDOj1oMSAHSHO0msJdkLEVsQfIe8N2UveehxKaUR
blmvO4BxiB0hdBldG93SP1Zli/sAzSu0Mlofjy/YlKKdGd4sn06kCNIUgW1KpcKpiqW8/hfSQW1w
XFybSdBcZuKWq4438CcJhJaV6gsiKwMn+/pYlDujee4aHTPkSMpnsBEvZBTwGpeE7IHIInMzcnk3
LJUpCj+C/3pBHxBdSmifKKlMF2Hgs6KdmkwAUraG81I3jS086WnZhVyPMeZ9LjmOAd5WjGI4DONc
LrDXiGQ6benuwiZRSGyq3wYjkCFpw0Rrsm08H4ofj40UbhRL+xE1wufecQgnaVT0yYwQMQ4L6vEq
OlfvtUxwkz+NBwRPNfIMZfYjojASRNUBPbZOY2ceChzpFGED3YSkenPHT2JE1/wGn0s9EUFPG/a5
clpQW7EbUGg6ncxkMTx07Jxch/nKaIv6srwtQ26+760XOV0B4cS9prKBXVAzZsOvjC6J2clOmY2Z
CI89tYuJnpC/jnvsZ0zErMJfXGuq6+fdT1EcfbywtZikIAAm8JH71NAqIgROrAm/c/m1qsXtoENV
9sR0OUTvpjn5Fb7d4OjDWK5SKmBQWidsD6zJBI8he5tCnt5fvdSqnNtsijm9Kl6Zlx0DOknXP1JY
Fup6IW2+i/P4Vs4rtrGzmxx66GfsuWKBKMGs7vwzC0p+GqO1fcEW6LavqafEHl28581SRu/gsAaU
4swiJm3SOlGnx3I9tg9iGwC3MtO8xL+GgUTkJxi0WF1Z7627eN6AQp5A3KFgPMGyOTIQxp469dau
jkVo5bP4AOpxSBkZ7oGCN8HoWZVE8kpMmftp5CV8EdsnFEJKU30aXltb7DDU3Agtgo8DGyTpezLX
eLmniXIt8X+rUnbGVbThrmZVy//3NDX0Obe1j4yVma1avSTLRpjWJvLrBiDEMZnTPtiZnReACpxI
LNqijZy0g/XoGy3AHZe6jkyg4jbjm076qkSVAiZKeTYs1z2dw/mP+vUbL9jM3BaM/7QabS1O96/p
3xgOg856/OaOAWHGGkEMdrWuORSXCfXiHGjr0DUldYZxNOdpav/MRMJtn8hzGTXd87hpcg5FniSM
QpZk1erzuamrJnSNEEfDrn0ihuB1bINMwFwiIXvdRAJ9rH38xkr9/PX1f6QDacCGvr0DxF8eOQAz
geIOVA9fkHKKsIPYaPW93gnwGDb3ZQ4761ofhy28M9bgTXJEuC1nsgUn0weWyDb9O06cN/l7meyt
zl83YYNQjrNxgRlPGhMUtkK+R+v6WhjalEYM7jDBXAs6WfAyzezXeOgFG2uPhhvqYGc7gpcJXw0l
58t5yv0DAgOdJWsJA6n1V7lg3RWrrGbA2drB0D+26tc2cway+M7/HZvtKt7Fv96S7pOlGxd9U0Ky
k3CtyRG4HHljuYlAkilw43EACpf74QyBXOenoUCRjzoqSLpCLfgwnTr528v03d3KTj5AwikP7i+J
+2fqNL6ROs+2Yibm6FSfreTIGFDjbKr0qI0TcHfClArYcvkL2HprWNlEZfu3EBXf/KpmbTvOv+Hq
zoeeG++c3uHiHsQ7x93HCxRlZY9MlGLLj0nNlSww4nE6gzBOGSPhq6zF7Ko47EYKvj+kFWLslkP/
oklLbXdpzbZ5zrTFYLmbpOAhR2+eql0+PQXzBkH3sB3AEmL5TPkBcZ0gve86gmkHV5OTGrWAj9WS
baw0tvLLcEq+R9PNQ2HnvX98RSscASK4ly35bvttWr/7Z7zZbtwkjp7L7Hzj9RzSe+t7ZOsAktA+
tbAfMkE91jQp1UeLes2BDPUzfGdA1MedVg8o8vEd28gZddZz6Ha/j3777QudWVn22pIO53tZ5Vya
ukUz37wP79vI8wVWeSpARmXbiOF1jN4WY+f5gH3SEpaTfrwgnsKeh9SNwtLFx8vHsRH5S8q97QOm
auMxiNI53EXb6HOhDPWrENWYrJfWjWjwNNT7E74gz23qUOKJtvCtdBC5Cu2WGktBj7PYsKcmdU4S
uaOISLPsnC7E8J+XwaWNq4G5ZShfrJP8BIVRRqSfoj19Dl6qMD+YGW5L8poAvXWN/tVkqjPmErjV
IcgpF8D+m2L42lQpFz0RF+uyhrNpwM1ZgjfraBajzEHjcea2j/sLH+Gd/UlNwmnHlcbVHVmePO3c
rqLdcTtINyXkj0YHfn1M9VXwMnUL0qzdgyBCo4kNtfsGRetoO0ntFp3Jc5QsVwQpXRL7fv7cLQr1
mSS/RtZtjU+gYghdQ5QPCLYMCysd/JH9OWMwbzunqGJuEiZL9usUHZzA70DkpG4bN8eR+d8uyO6S
PtqZoMpvlb46gjXtXlfyjWGGIcFPXZaN/OdZDA3Szdk7LKSInZP8ZYunjY73dMBbGoqYLmCMJQ0X
WOPpOsuI2lh2gc8uM9YYSQX36jsVKPpyTpwj4VXXGhy/cOeg+N6hc+KtnXzryR12+NjsSwrAE7Mm
ROP6KV38rEJter6Mu5yEPVjiLXh6iliKnjiQhKry+7JD7BGHcXfzO0J58m6mBbPYS162V+ItJbqN
mjov266BWlA8FLzhWJKwnoypjHG0Bce/g0q4iIknX+lZUe+bROQEZlb2YwVQOkBd/+E3/yp3cOuh
8vLa/zjUYLyNPmueFPKvXE9p1Da5/VWj7CBUKFZrVDIt3GL222sOGucEQwXiNqxUUDTsRHUzADV1
n1d8PdBth2ugy9wOOeUgB8jTFvGzf4Oepj5cfh381A6XE1FcexBS8rKviKoHlXnIbl47VzxQZR5/
EzztPUplXvRxOsjaxqcFtkBCRfS6sfScLpzYkMeu1CiZtkPVGZEWPMjrrpVGNl2oxV+58WJBQeGF
gCqDnalUaZwEq7Mof57apA58nmaqVcbpFJyJTMxfI7rClHq0CBccxtUDRNpxLWhWKIq0zUTUX+Jj
PzJHqWwQRS628WUqaxXP8SWDESh/6L2hBr0qDxdb2q8M3e8wi52EkHvBRGvo2jrh2a6OOYqz3tC3
e1OXhViGYqBw8Vl4E/OoCMPsCWLIQQNEswmIaqr6x21y6/Or5lXwBdP38SN0JjXC8ah1l/4byYQF
QF6oe0KrhtpXeIH1XQ40NdrJZW3SoTdx7m1DNgh14zm9PoUnTfMkw1NZZ2TN70jpdFz8FnKyAC/T
Zyd57MWLjI2+GLeTN6RbfbJevwgziZapcMGkrhPXNexDNJboW805uyACciGCjiqaqrF35qIaowRo
hRiQgJ4MNJC9f49AC/KVUzY357J9a3zxxdxj5FX07Y4Osa6CEZFQox65T3622tyi8jqMMjlCuL+P
hJk7gTewzbrVBHookcdhjGueJIq6oW6eY2z6lXjKhHfM9uaPIa0ZjWdA/4cSaEuzg69/Y8FCGduB
5u5zi4lKR2xJIlfApUEXhzRZELotJO69jKPws11QST0QPW0sr6xwYesHC7W1wyx59MsLSpFmuPH/
t75QKDu/6l0CTPl0An/iHfLaol7/aNiWOh6ENJrboatJhbasTSKcY/Zi8pY8L0zKkJDM6QUcKnLv
6tBNP8aYU+J7XuczGYaIeS0abiApodk9Oxnm8dM/Eo1/knisBZJE5N/LR/5jiINclSoNiYd9uNl2
oOwLi1T3v8zJxq73zHIpJCVKX35GxUPRdOvYQJ5RTfDO/fV6vKPQ/AeuP0bUx2T+515gqssvhRI1
1r23WDpr5cVtjTGG9Khz67P66LAG5ZR64zVZfF3kWWTL6VmrbcWHJYnuO4kaoyZWpzYgCu0jhrnj
2Xi8G4fT5Karf+BJxIDOg3ZQGU4pIxkzxCZc5rkBXYgxL2+fUbk0P6L8mlLWGaXNyiaMiFnmsJFZ
MvtKiHjj6wZ3SoHfUbw1RYnGOXPVdo6Z9mjIzNNbBiCN5DSfHG79MI1C4W0zgbQfTp2nZ9draOxo
tX7QocNBU9qyjns0GnlA3bewpQxlX9FsRdsvl9nutRg/ZbUQ2aZ028p9q+m4+VzMYHj+R78Gl7yo
4H0Tqq/TARUs+SmhARcM2jL8Jlo7dqJdYYpDgmYxiOH2DDMhBEYKf6VXxFpEM0ErJkax7dZLjxHB
tzmYU1y0h2GhYdLe5Ls1PrPzoJ8DP3EceAecozqTGZy/enNrnRhKX8PRznN8+HxkZgRW23CLa8Hy
C/nSHD1oWIrsj9zdDM//aq9SIDfn42JA4cXuMcofyXX0Du16R8c9VP62PL6GL7CK+4Xawe7RlpXB
C2Flx+Voz6HEwhE54EWfeAjAc+rhgz0ttj9JLSwDWqDwEX4fyUjEnmoCgSML/V38SY94eYeP6qOJ
YnQrqkfRDwN95rWPf/UllrGKLQ2Nyf1hGZld2mscQNcJ589jwK87ZrZvOtVyQinibUsi2ZapObCC
8zysX9sRonVlXPyXKBlb0OAqZdJhbbXRH/aKyF4Pc5rZRsx9UETRdjN5tsYwym2BYB6OaxN61VMv
97d7q+7kRi4yEI9upUyowPK4+y8z4bG6Oivdt3rXUZm8vjfDCuU+m2zkblOrFUuJLALuSlY8S+zg
8BdjcQnuRNYLWNEfpNRmXsZOVgT/EsFlPnD0s6eeiXMpr5jafKqUKfz/W/+vZ0WelwNU+9xhMuCo
kS7wqHEj8+ez16FQ7CfA/Az2rbL6mpjtCKpW3NBT8IED4bG8asxzRsUPOxo7fwthfAr/45rYiRw8
2x2FTeB9ySvouiFhTWQvvmqBvxbA3YSw5h+rg/0paKpElF2tBSAAChlHih7q+kIYE4FVWAO2Fmyx
XUB4lQMdNKm6VqX/Q5xFlZu+OsbollVSZ3lr6X9t/IhkLH4ZgMo8ALkaozLATIgx2jeO/TYQEt2n
aqObkQiVSfD1YbjjujRot598JxLOtSZ+CawkuTqGn8/tQjCL2cdgfAnEPzZh3DOI4GfpTy9hJBf5
5gdk+zKFE3BpVOPyKDkVtQMifufl3sYncGPOLJK6sh/foWMgdFpOyt3OyOG/bjjKDyvjjBSuXHMA
rqbEoRo7jEQGvedh9Z011vakpsN4BZxyxzn7dX0mRKO0HYpTzz1u0zlkkZ+TTGc2aiQd7ykUt0ro
OyM37l0qYRqCP803DZTMVPA1rqhOKGOWyy5q4VegYXNXBHpItdm436bZnKj+t4dnBOCwel7gMu0o
29JnClAEz08LPpADPCdHzNa/GM2T8Mtj6UkTmHvaZJ62c1vc1Eu5r2YE2SEdz9jU0FUksAca2Wro
r+PQvqFqWaijb08as2++FlnMCGCHxSKEFcncvA+iNQov3xzWpSvZPSlH8USgInr4IPUOg/DA6dxI
eZf4zps/343QzHETlMu+3tvMgTqNbIqGm8/7uPQ+oy68v01nqP6lMCbfeVQGZz4+6/Ztw2FsmM5R
VNd8apTzrD+AUNLJrpDPJmrZUOG1dl9saIwYc+GN+AlaNNKYmhmiEkvuED0VJNOUuzdRwvxMCNed
tRmyofSOxbpAL4Qh1/Qn+h7PCrtImcSnMiRq3QwfzVaKnX16tEnqm52GNdNohwxdnG/d9PKFvOiU
O6xxjomZq4VB7CJ7zKQzb1ltLtxiKkl4iLgH7f8gIJYU1n+NEkibXm8g5UnEVGhh6yLEDujdcP3Y
SdtF13F9iPagCH21LDExpPkUxBvbMn+DMldXnd233/lsz6kRPjkJP63vKEWI8edx14pGnhUx5L9P
PhcPyFSNf1oUkFLjofYzIP629DjWfxbOmnPrhCg5WS64qvJtFf1t2qTNHvRWvrZSiGuXMAWS2Mjz
2++/C/DAM3teC5/aybJX8BNiy02Dj5l9tAgIOijKTfEg7j/B132S7xNAkhxljr7nJvp5wa63WabG
g5BBfq3WDOxAJKPJX98z0tlSCyHY7K/NZo2wtAV5TbSneWgzwDryhrGyl9BNLYgzrz6o2HmSaAu6
GsuN+iCseNEl2/qMvZsgVoNbuTWqRfn5dFNQiwHULkJa8+HS5OOJ0KZxuMgVE6jsi5lfsKW3paUL
Cj/GcQiQpZRcdnejF1VpGPNZ2Z+JrhdcPGMCLni+HYGngm73uQ/LAiCG1Y2eDLzvicMv1g2RvQul
Pd90iAM4EGPkLrDu4SpOg7l+QIIdobMp9QbeWrz3qhDjxOxJMDQRop/zSSLWtn9dPzxPIVSFRYIh
pNqmQ1BsQDTDGITv7XxTavfN3pOn61xntPRx9Bh+lO8oYSEDf8V/rZZcrVk3ZJpfzl3iDMGw1B5s
/O2gy9KAuKBpfh3u9SlUACOS44abvf7VP2zlq6MlHvY+6K8tKLKHGY7OHsJ7wXt6QziShpw6DlQU
fTUXS56uekwp4cFfZv2fcbuMUCIFSjYEuFuQ2g08KO/G4sKketKeCa/2tzdIbaNnBEFaFboXyjWY
6G1B7glayCh4/KeifKCBwE9KRkwYUs3V+N1l2fxoyYA/nT/6/E6/XBBgWID/ZHwrcmSNQAjf4hDA
25ZgqP312pJTlXrfKOuo3PxmOa6IQquyOKFFK+rdohK1s63RnEyGtn+5ok5nLHR5nf2L3ehDaOsL
ChlJP7HCSKzsL1v4Mjm9dL6FtPlCKGtI7h4uKS/DTtr9TeuTWtzmGpppi2Dz5ZqY/dSEYi/6a+27
rKwZuQELX3X5EaU0+jUd5FJGOGNVZQ0epSIa6Dk/Hz6OrcnCDNis38cF9dfqW4ECu4oMx2dX2H8s
45VF7dkt9pjycNRVW8EZp145H/VBckpSKAYLmcwtY8no4zahOw3vdQZDEgykHMW7UXhancJ6hKU/
u9xZRqoRc33ozY1uxBVg9vak40MT+Q5gIDZ3ri7gBG4niTEAas0osr4FsAdR3f0vqr2gZ1DFoVtD
1Ls+3WjH6V3KwaFlCctPRhsaD982ByINwaTR2RwheTN2a3K6BtLkQrz0d6kJj015CPZq6/Aenat1
q768b0AABjpb9B03dkwrg5t5JZ2ft01oUiBQ3QaMEIOgCofhmt8IFfVpEutZtqZFwejSlC/8XS8G
kYiaDKJ0KXjx0ZdxJ1EEpM/3O1P4zaXjDdHfoCs2OGm0qYSKtWJQW6X4Wz6DldG6iH/FRZO81S9i
QkoyQrscua/jTmz2vrqL+Sr7iTzhNLWo7cXaKPSkVVOIWL0edl9qyEnd+VUw0BVmspTlWhkp4z6D
Zx+oSpkQ8BERvtU1Bb7tVw64a0i2DUxs6uEQi7krtbYx9brmCnrd1YSTRMFr1Kxm73/uY4fft27M
V2wq88NW5zlDH/qnfBfgmL7ucanfhGPmZLAMkScysH1/2tNHly6RLlqXsUdwUGzsSr27xHbtpLi/
E2gxMvVyDPWK02gS+gbl/7jwhSwPwJZYfYQfAzHIhXvTB89dN2qCBTKsRIaRrHFkqxiku8922A3T
Mqg4fvH+Ar98CqB/la/l6Uoizg4f149QamBrXJ8Gu6vHpzMEZSEAKWn3tmpPKsQWSp59AR1mkxO7
z92KmmxdLIEkQtnLBjptnoPyfCoPz8J9veAXFUZ29LB1ff984pyJe2dVYE3bUL8uxjQRz7TwYoUo
gZVcfJIz28569XmPNRkfKIcHW6t2zD0oJGO7LjZdbb4DiWaiMcwuAukCxE/c6TqZTjY8kWax77sw
j3vIC6BxhDlZ/WuCIiHd80iywH0a536fcqfaYJYPP6ELuv7u98YIQCS+BXTQLvF+5/iBUwlPFm4R
WVbN3QHg6NdN8b5/mVwRDsNzaXjc+Y+M4vJARLag2t321GU+77zM8v6heSFY3UvuJInag999MTt1
GmNiXzo3Ju52qv6QXwWQWiLv+gdeysAK3W0t6EcUzlJnGbVJOF2JPx63/ziU5In7ntLP60rBwTej
nvwWOlmqhAMaVgCbjYyf7trhRacPOue+tVIoqNSj484r2S8H/LEviCTBGYONWhlM4wh/IPm8Db+c
D/rFF6BIgq2KKBMAx9wJTigo/6NXdmuNWx+/tSSdGJBpQwmzeTrRqRSL5tnMQ5WKqW+H3NOVWk5H
lERmfwQmKA1q8b7bi/l4hONoW85ZLTTANcnxErQTBtz3ZwN0F1H3IRvE2XswqH9Um4Uysp4+dxi7
NA==
`protect end_protected
