-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
K/B8r+b0Tbszd+2pVci2Y2993b2ygcuV/OVFVwC5ytyIQeMyDPe0ibsXOX2zoNo0GtcL+cYRdvgD
W21W9PpfI/j5Z0ez4/6px3kphYt0HaKgJZSTrMwU5TzzeamzgK/oZ9V1JwoFQWYuNsh4ZjcBWazJ
lR9fi0EFb0Cznl97TAWXAZ/HM2mx681ehCENbWM0pGPjAITuqaFDJGy1UwSK5jWIXGlFtfoTfV0y
IOHM3jdF/KtTSAHu6SHWH78icXn/rpvmk6sm1C3xgCpmOS18bWimqnMJPqKaIqpIV8w9UpJaP02a
wKh3arkEIHLanKzZTaN8P5eBSzNifR4ychpe3w==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 12848)
`protect data_block
8R9IyjfiXxjD8wv+pkxqfzBBwqC2o7HOkRm21woLnSyw0dUwGdinBWSpkyXGcOYKdREDZyAa8uKc
NlP/IKQIxtkTa1HVgeYXsB3OLBQrxFwob5U2YtZ1EyncaEovTc6NkzvnUhDsHqa2ZqQhbriqwGUr
WpyWHcZOY2GJlM47DhkAO/b8zjDYZW93e5rcX9cG95IyZ7h4uL82/Lczwn9raTdcW8YYo/bVH5YZ
xDqn5C1xgpzPrpQqqQYy1WXR8fFs8pHpGGKzWc8OWR0dpoVaLBeVg0qYHIvlWLHqhCyH3FxNZsw3
6fbVcCe+YWpmxbLRtYRZvovIyW06qNXSkB6S2oX9mvW+6vsyMuPzpYhpt1mft+zqbEQZSavO2Cb3
TfZxADsrOBUrCAXICx+i2bNwIAcQ/W1/nGvyqEUda5Pn9FHG2PSLyLFfFfKJ8K+1gLPS1KNjLyRh
4VyZIivzlZSl81NQoJyTB5PRcB0F9m8CANGRSNwikk/+3RqgJY2M9Jazks+4cKLPPhmw3ozxZHDC
rk3lKTHW451VyM6N8xgxtJMyPMncEcYotW+EBe+JXqa6ZrJVPu3eiiQtmi7OcLqtxGRoTzWZ2rDE
of3llu1q24saM+BVJj6Y3QjkiAbZM/uMZqYLeZKTzHZuVCMmrXy+uO+rKZzQvsUkq6M/fGs/4MoC
m1dWHQm4pW0IThklDNlo0UQRfjsUvTe+Go1fNS3j7J5lQHssCV8JT2P1ERyzXg9+jK54IKaKzgE2
8bc5RO8/753Afp/dekzPL+sZxlt/jqMqBvmT2alT/3vOisfaZ0K3GLynIzqm3voeYdY7DVUesNn4
26YFwQ9mt3YmvWNz1xvGXpIJd8OAJXMARwnv3LxNAgk0TSwPwIIXearyLcYVKDCgScOdyyqb1EQU
7gIkRwNt5Vjsq4mhGUYXdD30z7BlqkOtDD1YdBIApmaZKxUpGpwfpWbq0xt4wDJlI0eX52T+jVNv
osxVfIvb+EZG7x//b1xZ14koPlAeKOyE4SGnMyT0jL85S3dCacF1gQjAeWqsJ3pPChHJkAmkYwA5
HBxaGl25uAbai7EquUyZJi/tea3qD5Bff+citEbnummFEOlqILfhEdLOaDkrPA2SH7D5raIJ6r/B
9BwXAMtcSsz7ngF2PthRxzIjx47kZXBrVsnCn2wCK+1HvG07kjK3/oiNJ1tvYl73Vb8e7rkpN4hd
gj5qQskiAOmIocMzV6mGnqvG1vKqis6WOT0Ukr9i4qjald21rPmHDbnwVgLr0lfUnUI+QELobupy
JwnUk8XSAUWG1iaAoVq2+5zM+xY47ZwKCGzPmyuLPzd8/LDf70XUwz7ftIqXWIBOjjuLI6+pUb32
V9oT7aUjP1gMIjGsVJQD5uu/Jh17mputf1ZDPWkWqgdROdezcGhBCDyXOoEG4yRHixAWWNaIXs7M
+cba3FlFo97ekqqLjh8Xd5Ii1p+6XfpoHFh7dlCOETejMSj3dHeWz5R2tdt5bYbG8ZwcshL1qHZJ
IeihpAu3sBO7miLqSZ1AKolU1GEsRnKYrZ3RCVfax7VjsHzoWAEvo9QQ01Fn6IPwW12k0AGSD0lc
ToTQ4gYpFcize1x7pqH81/qBf4/s4/VjhOMMEqsFh6yVFhHdcxZ0niwHA/xhO7HgFNc7goti0tpk
gxMsy/J0eyKBXdurO+M5fDYVbEQIjuXlxOMhr/zhVeDMuc4fSM9TZ0prz2j5OHr2oRnh/eL4I8sO
Cdd1u5+6ayI+lu2jCvnRU/ZWRdIXYXgJ34eYi7Ak5bi1rqnRNN1Obk9STbIX4DWX/GOQjE5wCyJk
63I7EvEA0Pb4IdNQ/ivBoK4ZauC29g1rb3jvAWOsh1NJtBVStRvxoNS/8fIJ5l71lkKj4HzBtQAE
0h23ef9OPBG4R7uYJEWrGtU5ACnFuIVZKJPPqJiMrnSLOGppL3AytrOX+EfnfqVfyHx439WQ3dPX
0a1HOJFJPg3qaG4xs1X+A32qfXgtT79MIUrXJflgGI/71kYlRgMdrNFx+ZoFaVM9IpJ5J+9MqdIt
949gF8AePdvUf6kuWYSWvJuAcn/bQdLjaExOlk8c+ox5b4uOHK9X5apMz2llejVhGCRVKX5NEzAw
B199xZx9Y7KvFV+Wxd2cBewCQ7lQaVYUgy9TIMKIpukvFUdnmaim5+TEN+i6AbBLQcWkF170Vkk2
t13tdcWJ3t1Mi/ahI/jBhR7rrQuVcJHM/A62G7FG/QMb87Y6nwBbG/+ZRc61mPGTCexNxt+zO4mH
TbzcDfqFELGH7Zbwvdj2yk4EuZQZXcFvKL8hVXdJcA0IbqX/X3vPdP/+jdAiwGkh2QcrgsDVusMq
dLprQEaxiPRV7DqRQ6tE1nvzF6Zh6iANJZRvSoYlFN0Cxe6ampaSgCQuXPA1V2VJqcOtjLCUd686
3iKCV0EwlNypfkUuvaIlQqChuc55nvWbzKYa0SVzf019+fAi/3HSpkOnD3A/KOUmDNlg3Oebqmfk
gBE3dBu+rAxXwEkAnmwvkr6TN0HYUP5h4cmhZ6rpgP35HcW7o4Tj7sCjcAUvPDVgaKBMcaPg7OWx
RvO6ObJFYesWZSQQh2NJlgV6RsL+KfLnhtotNc23FDEXghP8EWUeh/Xp5zxDnRCMJOyPv3fEvCAO
e2g9q8UxM5GRIlzcVjrmosQqoFAUq0SsHRmQ1QznEo2NDvtT3kFlO9+iXk19nSWpNxaI3ViPyg3C
eD1Jsqhhr3CQk4PCYWWrvXapObwr1e0kZXGNUwQjrWOl7yKLjIFVyXW15uAkkHWDYwwGB4S6FafU
VGYhr4vyDJeqVBUt27IGKaaZSNpRA7l89IX69svO0A140Lv36leFEB51MRID5uULpILKGvKgJSmM
U/QJnZ8JwolvVTyfqnktWwfPLEPrLLPWIIY1Gx42P5VNKUv5LtiJTu+wNT3m754QZD3b/nZCv15g
fB80SvG72FeQ3BcMEbjLwwaKu6ltsObUGKpXMlv54k6oNRzYnbVaeSglGuUGmvD/zgk0Hziv0eAg
F7k7jQKhS3UCgm8GHk6ogS6Y++0NXi7cZ3cTrfLBrFPTzEt8jMVUKMivC0cJixgEUQABDdHhxXRJ
CeXQLeS5zSBkWWumgUPr66BBZoKiWsnaw/TGGmopIoPMyWuC+d8KUnWRBPWtmZyFiTp3Dq68lOUf
zQ0ocnBDj/m4y9sLd7JxFD7FZGRMMA35M9SoLPiTIbPJ++t7v6+IBRiuBx/rYc1GmqJRa28Jo/eu
OmpRoXpPmgv4/9jJGDIfZO8sUMoOYSP0rJ5mV5u2qBDGWEPF+MM7DEFXYfTKlkR2O80aZhBlNgY6
HDyDDlINwUHeCp7y3jyfEsoHgr7lfTIU4TX4GKsGeN4yo5B59i3YoO7LerdXPEoiqVq9XJK1jh+p
rFvg74lza1/HJRG18nYFhoiVjQUQfVvU+SFwWzTV70XLYSdn8fAA9D4pz/mQZeLojm7RehBos+8S
ebnj1SKuDQTWvjkOVR+FLs4mXeSgW8FSLE6h2qpOXya1XoglTrNHac6JXX6y1Bws3wcyiXrJ3TEV
45+w6lMl5Qa/y73Paj3Wzc/T3/89rlGHEtKbwFbLmoMpFO72WLROE9NKN0m7agmFg6RdDZeDF9y4
7m9ggKVHdHjTL4At3Rwwa9ZThP724i65/cFZV4V1o0t7w1jh7pGzeFQEjE2X97gmOBlBURfji04K
6nzDA4LMdiSyF2jF/dn3d4oPJugJr77MvBLpTynyne3H/oHL6CTQjlihsk6DsGWlTjxTfuMBveMo
ONtmMgZLsXhrWL5SkK+lTq9fCV7UzdCDjwhsOAQ39FXeEfaBPr3thoREeK0P8koXCipTJishMeJ+
B4A8uQK2i7bYagaEKbOioimD84nYZJVeE5FCCuoW6G2S95B8Z03DeZySNOtVCIkDE+IzD53+MjhB
ZbZUrC8R/fO5oaIAfE8dXq7Hrc61rOHi2OK8PX0wlkR5a5FF6qqO9s3jB1LA/OadeCUN3Ow6V8Lt
kumJmzE1oeCdwHaNDky4mH5bpNdPrtTPA7C/JoTz8N+C08RicYHCgFeC0iKsFGWI0R3poWxyUEXu
qhhxWIHsjJNs9HEiA+kqb882GW7BO0GlEB1PxYYDTpkHtEPpsPOyhioahxquHiLOWQGc7COo5LrA
hPlb3/Zz/eOnmiDQzZ1HIvBgfO+GX6a7YToRZaGKbbjaRkVnmBaiONOpWJqaak5ovw4uvUz8kBZ/
FD21aE40/RD+ytKJrcG+PYVf7l8gvRUFUNq4RhHFUGVuw2eKnbxxnLGOltIU1EhGskgOwAhg71rh
gjD40wTnxDwlk166nmaKVazCrbWc4WZyudFt5l+KLehCZgYpZ/p9ntzGH/PyOBiK7Y87rcDctgxn
K/7JpUFMCSaIUuwXlCzs9zKUA7rMGw+BdeGWv6v3/tQIgU2a+656FvwsHc2T8kk1uwAvrEIGWnlw
jkS9+7uoPIcRCVekpVHLlcCPk4aKdz/kIeAtFM9hpS7ORKpL/NoUFjrEwtkaZRvrtPxVZM3ezqsT
4afCYO6PEDzlALyXj5LNxx0WJ39jH3IceqLMBonInGnC5X1oZhomX2wG5VHblrmAheay85Y+M+LJ
IhhUlUkU+AbxwsJ6tOfJK78UCgAJ8vJVWKundQ5WSJV0eTDzcgMu8aho4t0Vdhtq3cMVjkihhvBr
4tCuvucPwI2H/xl1GhdcMYvY2XBg/TdBTBcIobtP7pSgv1L3kE6/Qc0+F65qRhLc9fu4U605x5pw
SbMynujV48MASdSwcphb6tebH1jfq9SAqpyL6IZw3TNSugqkfyC90TWP3YkMOmHIv8Q1YNpZBzyt
M7JqdJqck9xEIHIWWwj9H5+QYBjLqN7Q9PhrPIakY5BBUXVu4wKc7ceoF1+Zr9wcIVFNR6WP5Pox
yE26FGOeYwZorVmOvMrRLmOExCN4pdLhoO1vMv+wpn5YUZX1Zvg+iROXzgsluFRqh3+URTjSNO+1
wCpE+EQfsUOjgJBQNYtpHzpNboqJrKMCIY+sAXGrQUs5RCkFNJ4mf4OvUNzR9G9k6ikSm6Tj3qxx
ZWbRoQ00gmvVHJCexun2bPDUjooTmuyDR3JySanmSDsLgooeGEi8xX0xE3MIC6pKFm3j7VfTEWF5
ms/No+nmITocS+dx3EnKrobIOAS6uYx7SPYKcNg7LIfJprfVxCz5PznGAhXXtG/C13qWsloE2VGx
MnD5koAIDUx8DtuCp2IOP+IgD3pvpIDyPYIh50lh3qC7e+fzRZGvP2KWJE5NznhaQvdRVexY9h3m
XxqJxfiVWUrIP7uIE437jKGuIqAgHHo7lLISvmB4zIuz3krr/IIYKei89Q2UCO3k8gWJNA6TQtBK
zFElIaiSw3Bzt8QzA76PfJHjcdl0UxVGrQObgA08jw/lVN5Q5aTGp0bHGdBi5ZgAv0tcv8Si9HB6
WH12tW/3px4wXJo9ejVnm5Tt7Z3MAKhmPJ1UPrd55Bd8n0q2m3lUAOykxVawqbC4bUIXY39kI51y
8Malfv3+eY5IJNzLifZ+QZsbfvxh/Kjb/pGOME0mjFX5RpkpaWYgb0GJZexJ/tAHEEsSmzMLloT7
XhnQVUeNyy85rS2ZHOz1iHezGOhgsynPTZ26njadG+XlCfo0RuI7gXVO6cjt+IQipbK8UHtpwuAG
WtHQK5o8rJo63C3EPIoNAXzxx+eW5LOQz9R78Sqrrd94OvGgFnbQIN2xakCb4p0O5sIVZfIZjW8i
C6Gsm+n4BS7NfjXy+lN0zxWIU7icoPXn3RqNDETW4Ds0sFtx0y/X0mYjwlbyB5oMHwTYLbxkRIi8
6NzljPYjq6zuslFqQfhXk8tqGEgN1NWB6F+GXWQLykOD3q95Q6bQOKhDYR+zxmcYWp/fpBd7Hl8V
Jig+EON7LYcZIBfyzfuJo63xCIxryLP9Maelr1Bt0BHqViqlGxAm939TefiS0n2SlBgjG3lRApqp
0qrqpDW6+FOcy45+Hf3I9S3JPGZ5b9+2YEougLPpV7+zssqLCxWnoeNgPWGUwRGTdLC0wI42A29r
5WO1biOcJ9yKutC1vD6KTLIGo1DMW1Rg0jR3pGeyXNpuj2uFTqflVYBf3+nPYjn/kUUUFESuZrun
kvgz1bOh+rMhN0REL/HGkXRla6A/QzzMl6Jh8pwHL1RrMWuVUy+1Q9PTVNqU+GoLGrSsJswGGvkj
vcgWNMhg9ul71Xp4TQYaJVkP9bHyLenHmwaaAlbNXa7jnp38g4+AcZwlXHgXSKsgGQtgsPxtLrSC
lQLkR3ybZyqKGdtIym56bGIayR9FFeWEsgp7HGabH2zV/cLIpzWZ7RaBwUJuQTy8mOVYbQM2RKzK
T1V6B4VR+ul2ttpJgQIMHBjlUr+5vXqvaLg9BwHY1ywUD/UTw2NZBmFiEZK6mX4wewd/rPgjgaks
9y9Wxw1VZ+vM4DoOsqqKa6GUqETzIG4BUqn5bDLFNmkV6BqWh4W2SHf63Om5adMjibQAW5yCMBSI
7YOIVaqXN9ggqJrinY+Uq6c3OoDcuekcY4Z5YJKcGEKtK6W32/Vwv4U4e6QbTqJWeYpVivQfqv7P
egBmAsX/p0sGJfDcLT+FlnbztiNZlrDf7AB4wan5pbeRgh28mj3yhP7qH4ItZo8iajNbHDSV6kH1
MuvN5qv8Fm/nLI8XRewbaFcQVfs0mTVBgt0SuMKbFIYxRcUW35bYVUQeytvyfsQ6utuyw4hfJZX4
75Kg1f75XeTwCnc10BykN9BLyaxIjbZOKp7BJ5UDn12C6fZC+KX4uPOgDyZISr6j0VDuORiG3OQO
YakqDHoI3nFjhp+hZVM3H/r5vlk7cBL5UGpDTKI7FIPtBuLUNKfyF1e56oMRDiktEOJ9jPv0l9Z2
WSy89tix6eABPLsyTxEsfOgzyL4Rhq9/eve0m4L4+cHNgUTIHQTHLM8aqMevb98m18VKJwuT1PFM
Qt3pnZZMy6cpLjQxmpZR7PGrBYtBL33NC4FRwOP1gY6diFi8gPSkZBa7k4BMdTmoaSATDiFONsn2
8wC+f1f4PzWpPQRFLuyJB7pRU1S926TVnAEGMKsUHbMEJBGFFixHX5KhK/vxU1rH3R9CRx5zQEG5
TK1GxxLMx54YqAn0ycaynCKqeMdYBtyC/sMer06GpT7hakigZfAab7ovxc3P+Yebk/dRVciY8Pkl
S9EyQfI2711WVO3USUEhAe3V+DvPpuR9PE5DTYmKZozw34y84VKGo+PCPmwqm+gtOEyN6TseKEBq
XSpA5viZJ/w86AQdf/EYcC3VKl0c7/8JzRJ4cjBRAlDsCmHU/IazI25CSGhG5Mel+fIdevWKuND4
l+aVXAtQgHfwlkpF8JxKLaWn8GBJHzSOh30/rfqKxPvDUDFKM6HUoFmoAvKns06cnmk6odTIo8ac
0mLbJqxzoQI/L8u+Nf87RGKz03E9IGrIFtSZp4ghC5IR85lv7WicmpJMH20PtOfc7iydDoIjxaLH
ew/upKjETEUX9sDsGky4Y1NBNygxcP6EEc+K/9ng4ZFlU9QuBGfS4FMnUlHVDpHTlbAa8dC5kSbu
SU6AHXCOTteGRvpljqUf8wgATBkssYonFbkAMAF8/WRjgFBA2Dn/rhmS3L9+g2Knaa83qaqwEedX
4zRHWiSk1noNrieQ/+8Fy0pZt54nvk/eahshaxPIluxrk4KXLFfbmrOKJj9Hd8c4P5SqqhMNZCsD
VYDQMQb/3jZimTyuu5lAp1ptGPJ20KBDT30QOvLwrSvzxadzzai6MiCuoNNg8q80k1HACYIln1y9
YDADXyd8407eZzD3JR/DYE7bGudtc0lstf2r8tBuBSQnu/D5+cJZO9LQXIeMTu8JoBfr8Q6b7OUW
7mm7fuvgNWrfD54J5712JqHdTDYC/h9f59K/MsrcAZlCoSFVGKbwz81FJqReR7DPo6max+nmGoHO
t2PqkB0zPI1qldJoIuCCNdboBHyqdBfSUAf4F6eHQHuEJHICgQcoP3albPu9RMIhcL/F/DeUGhnd
0iDJ5IB/cBBSqyCD0sPg8o/TzfRbrPX9mP2cjx+TyUVRLoSJ4UQDdUDTYD/ny1QEifTeeXyGT7iM
N9ozjBy/XDiw7LTLa6367J13HyXi+Dk/BOCxgUTeTMf0eYllG8JgMH5oQdaApRPRzI7A7L+KqYrA
SYOXES/1N3W6d2pIZBiG0teZkVmqxVOY4zYD4aQCRuAX/+f8oLy7a7bbh92/youu1nTRvXyMWrbg
h+XNfpkeYCvfz/fOS+pZV59EXq3TxqnclZqb1dAtCJ3UJ3rpCTxW8dl5KApYSt7KZaE4yJYDx/f1
leCrhB4tR2BQFOkYr4oPeEsDIsqgUa8lJq7/yg4cXQkb93ApqpyYXC/o+wkMcvva0hXM0nZl93UX
yQVeGRh/hGQMM6y7AZFgwJcSDXt5BzvWvQIvoljA79YUFL2Kym0dq9QDogZiTocapROK/TpfJVW3
Qm5D/tKIlFv/Rqik/DaqXYVPV4ZNjZKodqx0scE99LmW19TU4Vv+SqZp2la9BD3ihpeHW+icb955
dmzNx7TtxB1hGfH5IubGIs31QwQAmdngsGaM3IqRi/1uj7vnw17f9SAlx4K5Sw+wSoVPLrBXDZ6u
B0UWnslpZfzf+lhmE3nSuwxxSMZqjWf5cvAQ89CZoFaB0sU5en/aAiz/2BPfOS18mezKtEuEGM6U
UZtndoUGrfc1UVPQ8MLjUMmkg4FTpvlQFtEBZ4eOT9x+CyApX5sBrTo1CQ248QLHoJudBM8GEPfz
xi4AkgLNkrlxwVUR5HHuxAT7PJPW03EH2L/AS+xGVp7XmiejeoejU4C2tz0AE3NFwhvh0m31UT86
aH8T52KWtEHdOpjmnYmFEfV0z36kPPt1aVbmPoH/yRLzJ3p7emtLfeT49jSFX6p4DK9qOGUb6Mr3
1K4ZL+l7aFKYhohlapz9o97EsEHvadwGD097/8D6BSynJxg2r3FtZx6AQPCrPLnANTIMrgiOEF/B
i0/QD7b5qjpR4wnnB+k4rQcwZCMMeTycEk5XZFPTF/MwWh2VAd3yTzuX8CbUB1AWT0IwDLCG/6Qn
cyl02lXscpfiUqhMQsV2jZbD3BTbI9rOslAjowNPgauyWQecp80x+foCclPKNl4wTJcJVqfvadbk
YbVCZCtkC4tnZAJFMBnYYWY4dkyz5S5UWM9E1SdHzwOIlmMm2655gMSycIGIR502uP2XuBvSqzxV
rpJCHCYcFvSJh2qunbUw+Q0Ey97AvhRXSzWwY+K5kq3muk7jXTjcFJGZ1ZEPi2ltZv2Tg1l9kBaM
KBvuhIDSdhGC/LZ2lq/EyVVVvWZYZv/GrBcjaCwrtk1UeG/aJrc3T9A8lXq/e/Oz6ZmrRHHOyij9
Pw7PnL2VjKiC/IFG1xb5f5wXd7Zshm0eWfQve77HfS+zwGNkKUqWQnm/SAV+kflp8OJCNwEIpusa
NMW7S0VszrvHzvrh+nAmWv02ipKC+xhAwSb9QlPZJ86fnBfvYRfRSDcV8wZGTc7JInFezDJYx+2R
aDfox4HP+KtGkGLLWuoTzUgIkq0fkX0iw1aBrrn/0vTHA/AAlTx6PSFMn2VNZ2wtbxHc/Algc8GB
S7RfubUJu04iWGcahtvtvkpv3HbQuOOz7LQ5+ZIGZvxmVVNnfS1840rv0Te7VuP0By50fb3dgam9
n9Hj+459gfNfnoUQUwKgIGhJFF7R8zmwJcwuThxWuZpLVUmIBXNrjTvKYC6s5i2SjREDFHF9AYAv
dwRnYJq8WRPrr4dRyWxRXz1qjKNrhXcgo6aU4BuWhJwKvQIZsH0nPrk2voRTVrOzh81d4qDruugh
3GDf64+cIDND6AzPXOZJvOkVAVB7ODAA5zEAth/cK6rlDxtcgirv/JWfMQ04gmd6EUAFglkmTgG9
pEc8kKfEASs/JC9faoOOpRQiR8a3m8ErcFvt2C/tysq3EP6JDy3+HFXumjhoqPA8wkI+38NFrnj7
pN6pD41ZrvxYGT1AX8lkyCPbPCBlLarOuUS4XKkU6lIH9Mro71FrKATI0H9bw5fNE+MwF5d+Pyko
ja+RmfytbrfcW1maEpB06xQRhdOrlnDKCyH6476ops8kTdQvUKMNkVX9vsRdg+h2JtBeEnzzH04R
DgzN36Qy/Iukm9P5AxoCuyhRAvofw+vyTLLiO7hh5D3uGtqamdC/s4fijOdraNMMLYeurpD8XN3Y
w8+gEmqBHNGxd8jqqoT9aTveobTOoqf5xOCDCMl6uHSa8eXfJZkV9LSIKuqf+ehfycm53Xvyl+Gq
MQE5ww/ORy20ZiMeiw05c5gkWKmRdyxpjMJciCpskm7Ra5dpfLkUUg2kz9kentR+5J/OdtLOrr10
dmZmGmk8RNGAz+LiwzradR80NVKjgbLdh32+rBkio2b6KEmHw/DdJyWUh5/erAlvJ/RNOzgzrQOQ
i3AfGrFt938XiTnNXReoJNGKaueMnuZLJ7K0nkv+Aes7B+W00qtogEtUY3mmaqXtc16EOvF/zWvN
oR/OMNiRU6PePEd7PBsjhr6XmxtjavHhuafw+yTdkW0LrrNk8UoGdRNkNtxf5+xm+Cuaac8gLy0F
j3bcMI5Vl7AzPWR0ZghI9XaiqLYf2z6oPwtot0Vx0RLHaZ1gscIkIMjn4AMsunCQpHvmcJN2p8w+
CCvRLV9SrBSlvplEZ1wG1o7I/pDnRIP4hodBrrQ1TJ9Rf+ug+v2Lv1fpmPWCZczBP7c3BGmh7bTe
CjfvKQDXAJJIeB+sHUK0w/bLIuWX9gWSqM0OH9Gpdm4aEiO6Fuf5QsnB2S2jkNqg5eN+L0rzW5VH
PV51Datv9zST4fOlo0syma7wRid3ZFkxbo2+X8FfIlGnA3axS/OEppwj2ns3p7VHRPe2qkSM9lOO
cTIIRxkrO11uTYQqOT+iMRwNwqueba11d7jSFroBmZr8Hv5I+Xa5nEx+2iaDhaBEjMK4EDCw431C
jFSLpUgRczbMQxg4Ej8xQb1gd7O6KPB1KPwIbc5BsIFGESkh8ABTfKPb9Pk7FcXWnY4JOIS5oIfJ
1fi/U2OUZFA/5otEStcyAzX6fUIKnBBRd2jfayLTe+1ARjPklID6OvMlQm/t7/y6YTGCrgHh8QAP
OT7+tqNQOh585b9Y9fmENFHBezmvkHnyWE69/tcxopbpJBRCPBNcz/vcx1HMvut3o2dI3TE1i087
rzgidfIaBag5J96u1UljRbv2kvkIicbGrBpr/+H/6vaIGB7+CPnX9B59UBQH572cvQ6MJHFMNOtE
9dQPia/BLjXtOKJsmGF+i6PmjlzDDmcoiaCzKcNL8sIOE0/mD1Fokr6fCjao4jUmoiIw/1M5cCcD
TKjJP4gFSj5z5Inddd+jgkzw4Mo9OO7gqFIU5QOwnil7sWBoCxshYtbG6qBs8H99nqo69L1g96FO
HTrQ+WjbBMhed/oGWv4yT9qjpx7xlAjkJ7Cb49So24E2Yr/chqpruoTCwogmsz6xnbzjNigrxWQT
QTmsbVYNpLi5Ni6nFUdyQiBqOQ6kSbqY+TidA7Ih4tahiubgF/mw7mS8tdKUGZrev9Sn6it7pSDU
TBzHxucfR/e+V49Wn6XThjJmQnK8w0vm0UCKFqI+lxqR4cQ9+mtc/2Gd26VVV2tNFk6uv2LLY/T/
yjZZUjbWYj4IyOlzPY6g+TgPUEcTDUol7fPaqxut7bpiDyM5sHAAI8P5qIo6a5qHuiNPC/Vzeq1q
Iz4eadbBiBqZbH2E3G1w7/lXIRloXzOVy7+Pq4CDlOdaEWHiSllkgEdjsNuulPR1JAfwZbYfcE2H
pvRdHNh+vBRuChv/xkr2yjUA66S6hmkdRhs8g9ydYs5WCJVHX0HE1Flcetr8DQrh+2DmE3nxh7q0
8zTiCeUrc8WVjmP1LsyZ46dp4g1G4UVu6tWXfaPjvXW+C8pTIKRa4m5PvF7NP1xUyp2Ue1OdXn8N
Rfz5AVowL14oivnfovqEXFxp8bZLha8mkG6zbT38aRKV+UP3Wu1Z5p3RCcwCMILLa7NiBW/uYkL8
UyxqXkgf6esqq/vXllBlIVMzH3vQh4vzcZ5uJuk62aE67Rie1I4ELjKYSTn0vFQsEMFO1hORW3Ch
Ypz3SufsdGyNiIaWhSzwKCR6oW6vEU+2V2JtQyH6387mNGbYw3unVd5KLwPwkIBaDL/p38+j0/+v
/2/+CQXYGN4uh9QyZB5lnFe8GVx/OTMQnmeWBUp2WRCcQF6ukZMeDMzDqtVz7OM/pY7TvT1eQnse
91V6nKpH1uacLiC1pBfKR3GiTERnp/UyXhzN2A3k674srOBXzGTWEQS6PatzE69uu91yrY7r/ELz
x9rPSdo3u33xeLJAD0hYHgjMUQF4We6Wz2AcUoPKQO+YUFstIbIruQt+wXSSiBe+nHg8Fgc2GOsj
aSCNwZrBooAuNjt6tC3EF4iyC3YA/O/gyRAjmpMNKe2dLpBshCsX5ndGLzZgumojEF9/M17tFmhM
2EWKRcj5p722qr4XKTtcxnhKcTgIhUW2OQ+h8IEO6Fi24kA/wPUILh8Se9Lps+CvN87eokdGK98+
jPZQhLZKHOLCWgYFZPCEKKUCa0CSXOTDMBYpTFfiLmJZMT4lAkvTLUihNyepnQ+fWUlp5nRT3ZIL
/Tw0TX1n1kTi98xSDRHReXFG5kTWEuUeWVYuAapjZMFDWm77/Q+SKHhBee1vGy8FFklsAPoTMxvL
4HL0XPQV8AvgLlyK35NhFingzorZNCwF75K/ZtFIc06HnW3ajd8zderxZTVAXk90hmODpxExpqkQ
hgB06EZZi804MCKj2UQmB/F3K7FH3RvTX3greqzqxZUv3Ru67Uep5QKduGoq5yOrt/57ynAqPJkD
V1ZEIyT5A4bXQrRnOIKYskrgtkFxnvSQXoxALntD5exFJhRo+qva3NfQIRs2pHbdTpkKHpEsrIne
z7KTFujuTYz179I7kMXHD1dqFXXXfHhm+6T9wyHGOPUIiTQmBwh44AilZ9P+ZNL4faMYxxeXVNfT
rpLHZOPv5o7ZmPfMGlfAITBPhRJY112sKBBj0YoJ4l27XZJk6yVWrxZ68mudUWTDqfbYUR0fYser
4WxYTel3hcb7P/upp1111X5DlSZTWz8XR2F8TmxHebN0AVSgYjy8UBSast/pc97wfAtb6LfXKzDh
IG6DdtG+xAouplL3sxA+DmwkGwYEotjOXmgynPT8e4w0Qhfs/rv4WpYXxtegoktKhVpwh+3sCKsc
Ik/Kg73uRJ9Cz5u1MPFyslhBbJcJstHfx7BlJCGUD5IDbJYznenL60d/2+1kalDiWgZ9X7XCdZBM
HplsfRM81Zit1GIQBu4KkdKPQ/6nGNsKhj1Y8zcw5MErpuboNawmrgZumw3EjKvh8Y3oL2I5o9D+
FfLk8RX8cQ0dBPWd7nwBqU4lruj4/HyVsAuhZy2iy0XnHviaOTnlw2LPkVPJ8Z63Zp/SnN4Dl+Gr
5aKeRhhPkZJY62esWG09MzrJUwHhGqCLCz94PHgQNQQi5JJhxp/GIAzLRpqnHkDXhTOG981d/Pn0
mdec2G55mcjv0AZml6iMYYNXwrVFbEn+cOXUqQAO+Ng2l/K0t/HJT4aum225i8SHFrVjxjWTriG7
jz8Ija/jZAsMOQi7QYTMYCvhJjzVPxz0S43Uau86wYex0Wi+3RefQq7hbyDTe/shTxKw7bWYeVzL
yErriaDkCOgl+/SIwTFPVTe30J8wj21kb7KmSPlVZUOyv2P7qE5MZ0pl0DWV2mC9B8cns7RwkSEx
ysT/89lIKNoVQz5wKeausbITjExc8gZLUBikXtU5LhvhCDMG6DYnYm27VUKWYkDq4PtibxzjHPvU
ZX4thsL/E7/wqMGlxP56O+LvQa/ikCK0p7iqNiHYYJOOvyAoinNL7DVDT5UFCkC5a2/a+M8AM3/1
MM0DkJrfzOmQfUdn1HwE+L5SITe7wu3Q8fLERTF8hP2bRZpZvnFbFbDVN/S0aJQhkF/s5s8QaFbL
BUWv9yIJt6q3rdq2SAaUyVTh1UdL0zLzGMizziQD3cBiC6tODEX4TezFE7hHNik9LJGZHk/BSJdZ
Aq3wwLxzVJRXg7a+/3qQxQbMEQS8XXfxbc6nWuYQ4vYkfy4ZeoY/ZnMum8F6XDmO4NqzWGZMf00q
fJK1W1DXAVFLUFuOg2r7TYYYDBBsowCgXY9a1L4dl6ORnN9vXnkWq7jl5mgcTftdexr8J/n4MCWN
ND59R/OcwjG9koskWVZ26R00wNUbJVN25mYB3MfoQyBKfOy6hoNHQSf9mSpn93Mju3I6hsAhKBNh
3fihFh9pNlZt6/W44HCsZ9RKzSs0FWtRSpyrvvj2hLZDttZGZUGm2o+NrB5S1sDxPQZQgzWcLwhb
cmn3aEn8j96jXnCyi2sKIzDm7EloQ6OVakmrDRu3nOcv3Itd61qu8OmnreI9dQ22ZxQBkHirMP8n
VqtGfYAkmIc+SyApbLrlSZWO5jxRpbxFkoou0yePUdiKbDEJTXFpPSXGsXfsjEvrX5X0iGPU72Md
oqoE3PQxojB0Xcqc/ovy03XoSJdm6eIJU1z013XcbqpQI4+qSdrXi4B5k8WyDSv5iS1averiwUxY
rb2fOIeRD6WaaTznQoqqtHFid0hi2ZAVMDf/UPnSDWvu3yOZPDOxWrwMm9QUbVgEXfXo1O9HEFg5
bHiEYvPl0SwEvR/nCqQxZdevwXWqQgaxYZnQKjxEfFlGQkdXc77M6/6WTizIjcA4FztcCTadmau2
Aq5aIf1JOSnSL3wmSrmYvHHGVyU/8nHr4xCaJ/OLz+Z3NdbyuNfidhYzM2C+i/C6XhEUFV6qLFY1
/z6vx63YrUd51ZoN48OwHT/z7+v+g9495afXkccI/CqMJg0Xcp/9L90X101p/Kk7ax+Clzci1Kkl
Em0BLEXKriqkwjRPWC8dpOkLl84Lwv0prx2E0FZdb1xbc+4dnStgYjWBdejRLUzEc1Vgfw3ekv/O
ubOJ55yljk9ciOM4ENUA8gYocx6G0hrwUuvAFqJd9uwelTEK+zl5f94CeuzxUMObOwUY7qlzpslp
uD0eyFO/eT0LNuofn9xld2pmkhohoxwHcOgxpdeAzGKR5dMpx0V3BYZ2ubtilVtoHLynfx3XEL/q
KWlZzYBGx6ornReWQk8gBCCjyJxPqt9sknCWG/cvm1nWM/t+fpMn4TagiU73JEJqP2jRUTqmJ+JM
KDwMk8jXchGgiDeOCbrmJ5Wc+mIBXpDrg+CBoerZCLnttg6uqOia3taG5nsvxeppyNRlJ+5+P37j
5otUdfTijUPnBytdX0O6Oz1n8vUM/dlVOtoOy5DcR+5qYq/3tYLbFgnohyy6OZwvHhWsGp1WX5Xx
sK9Vl2FcgFLClz6qYaloB7tAwQzRkKzz0IjO3e6veKU4sEuZsx9x1I/rlpl80zvM4f355f/q3jHZ
pZ+fGZYGNDVJP+FwHnQ5oy/uvYa8ZLyYm8M3qVcjCT0clN8IhCyu+lS0GPqPPE2eMaWFml6WhYp5
U3ZnlkpXoKQemmQKbyaht6oYFOTlLtx/sQTCyW28DXJwmQABuo+36dr78wIK0A3m6w1L7EXXSX2N
uzOEhHfphJHb8D1fX980uDKWCnThJ61I7mYJfvjVEQ09s8yGkYcas81CLnH2diMmVrbia3gSfNDM
GGL+FBK/JL59/GSPaXd5DhdUoubStaObGf94OQu3VVeXDBiUqThClili63RtOV/l+i/9IJTDYHkE
1cFqiVmI+H3sACPlVT9HT0VbZ0L2exTwzo4/RA5FQyN7KZD++a3ZvkMaYEeYqXrFfEebSyhz14zY
6CHSDaW6NCp9p3Fl9CFwCZIqlS3ylwumWLrLwmClYRpCUXdYLBwHoGs+2Z1OfWSaL7Nx9GnUJdVY
/SNqznDrOC+d8Lafhcb4f2V+swNTAL722T4bAJIHiB8N76tazoR6ZaC5RhouPdXjV1O1nzZSGPR7
A8iSJrB9OqfHFCcvOh4pqnC0gKH/liDwnvCpA1J3qCLZAm3zA358le3kelEvZnwyTxbbni9FZXul
2XZjzDX2OvKRronGunv01oBGm8Vr1sbNcRN6MHAaFtsCTgVYIWVba5VxZXTu1Cy+3usvbsTRmRxp
2t5sD9jX5PjDG8ETy9WYJfbLZ72LgL+z1RJXkEXqzXqKVZTH9nEJEeHDqOVESeQml94RDw2lKssW
Jv6wt2unj1LU6+q0iBFj1LX7fVyI4NTiC+lXfzwtlccyURJtRvxJO43UXUwjtCGGCgg0HNLxGWEu
hegqWpXC9yJeN4KIRDJguuA4JRSnq1KRXjImf+Eay5jQ011V6DaIkHRt+XB3M6pmVPgzl2zvpLXi
BhDgHtTsF+O+Oz3nR63yOcWAuC3xVu4o4ArsZ3ORoK5QON9e+Pn4U2HSB4fLyuT6bnefh5PqjCea
xA9ZMUIRYXqbinHyShKNyj1tNXFJzH6t8fGGRvHl1+aFVe75kvl+zwg1nskzm5ly3FURwrL/7s/8
GqQBaQ5BYq3L0dZ/rHw0Cbn0AbNWyzeCsGgl4e6ONLLJV7FFDgNT98o9v2tyW8DUzb3EGGGL1zHz
SK9xzq9x/YymLXkql+JBMSL/t/j4jR4mJcX4Sj8sUxoJTydHWHegSAE15pNDCFyriuikjHtMOrxl
dA3StqdSDeyt74ssYAjS0WcvJfJ1LMWLaaZGQ1y0uXauz0/vmF7S+uObe0sHVFBWLBW1RPs6ESyw
pZxaIwolwmRhK50msoGCCKf39qCNLPVHxgFFiVz0XJvww+2yaWKDG8dqCthbGyYdMXukL6Rjun9n
WqAn+T7+nLjjgrnlQhWwCSSUwt3FpOjmdQc5227oxUOQLEudts+2ElXUYMvUurueIG+Kx9UiZdxJ
Nvb9ekI+P1C3/66YUC+QkUgbmobGyofLMWdI0jUiDbAJJkz8XAEw1jzXXlayxT89RrpYIa7y+okn
N6Otd6ad87eoWieKypXBOcrvO5b/4jaoSLsv2WQ9NU7YPAln3HiedC8Cm2PFY7v0TGrlZDySAode
g0Acb775gRM3qywVYCYUDDOHVbSckGo=
`protect end_protected
