-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
xH0JkV7BzuFQ8kLBREVVjvokI2ufsn9u8eoAUyNsGf9mcZLv7+aBv0gCdPq4nyEWgYnE8wsOkoIt
XjvK+Hy/jDwE6nwjE3UUJSkXEQERpRAV5IIfkSoH+9yQjQIDj5eW/jcXJ8BOObNeP1ZFAx/FjmcV
iq+NP9xMRVimfeiR2ijDUQu/1VNV+E1u1HT7KZVxlC9WuQTlTf6dCGhvqo41tNWpL3fi+d4fOuhj
0WxXNupbxgGaDXBNPEg8uSfpKvxuEOH2NyjNw0cFi/S9JX1RU0BcZDbyiOaEc/kn42UiG4+nm7Aq
f9NRCw0U+twoH9gik1Fn4KgptfJOIsMQrnBd/g==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 72832)
`protect data_block
MYfzhbyuS2VDPh3K+jakHzi/2rdxAXOioaMZHHy7Whkc585kFPoKEF/fIwiFu7i6iJ+93s2k+2T2
/+sgv/a75kv18XycaDHt0pm9Kl+j0TSpYihL/j5VZG+IJKLwvCanWHbkyqW2vrWza33xRhahJCz7
m55nVbidMAM9ys8s6FNotU6fkF8pKAkhRWF5BoF9DySt16P6jFj5Rf5e83DrL3ZSmxUN5Bw8fR5i
fH3WsuRg48xNVS5Ol8Xp7zJHMM9FdsVyWfi1qyqrzaHc3p25god/E0pM3RipCFh6wgsOelcFUGjl
wPc2AkuoGtn1lXQqWl8nQ9YKawPgbsdYRnX4w0TiMgnUS9Q4CBb2O965PtIGik7fnIsWVDWWzcFi
vpuR5Wq2JilwoGwWxJyXiSmSslxc1IdJ8/oaKnPNQ1eXfaOTpkIfby2NwZWExaVPEs0i5hBLHkBV
ytF8BLjhpWyfQM8PmzUc4q5dKvbMukxMfcy8XX886XsBJIQqAVB/D/m9WGERzg4hQSeJIFZARfe1
hdmHdCL3CxBYHrNbt1yH1nmH3ZAn3g+Lm8RQcOi92uF0J+yp9wensfsmiuKIHgOrjg4hk2JeJ/88
BPIEldEy8CRr6HJmt2FO2vUdLPdQkczREm2RZreatxuojnpkzIgVQ/oTiVqepFObScmpC8FaQ4Ad
3HHptyP5TK4H44uePSrVQpMlgl1BKEnH4gTkwauCdrG/9gC0PeJ0cnKQlqwCtAdIlHWyYz9nVsJC
d/er5JMHN4u1JXK9HvH8qO2ZVxeNMKcajO0LrwYWfSoFrir70HQmC/T1+vwedpjfrOB+xR72vJmS
Xw+3/OIG82aZMdMcesC7h0DqMnjYgt0fQkYiludGXT5Z4Z6es33/aiuRGa3ys7i/g4fEPWDQxho9
OuOqlV0O9ooAG38mCQSr4ksYsqxq49siUPnulqR0SUAgfJTEJ3Qh4dtooXmk2s2jKozsXnk1SeaI
Jf5dIY5wg+KxmQbyzdrkTDj6x+zUVIc40FPXCCTQm0kN2B5eAom7m7Je+DC/L8euWp8HDQ0Pvqqx
OASOOrlgwhAxe3Ui2AYUTr1qB0YFT7PyIDtwF7YnZpPcBOYga4ajE94MuiNIL166MEHnl0a3IHuT
pagSDH3VVUxmsO14virnDDOucV6/ThzbH3u733wxbYp1MV04k/Q784yD6LwbszmZpl8bscsq6ZAn
mG56envdGkGfPaXmbM/1eU/I020CuicmMHchPlVvfxh0kzcdDwiW24Ao6LA6AY0EaXafKCCRYHo0
a4h3O5xi/ZqQlEek2svv9MiIdQBdEL8+QSGav/sF+QFgf5vMA8rf9RGPIV825UT6LhDYWMzsCYYY
n4q6PD+nGVD+YCDabfZT+4ybxeDAUSUSnf6QWeCbQhhNUuic3EFM07r9Wtxt9J4EjDZMaqlYpHEB
xhP4DCyMqnSZ38tF6iPxeQO4EQIA8M23Av3cYJVUWOWmZikyEtSr63UUKgrxls/lsuTvBR4UcOpJ
TPAaZ0YrzpGpJZiU2o5acQ80yVsayBLvsWAo6RLOJeNNubRlaT7oSN9BiW9YhG8MUPR5CCWQd66r
CkkLrgPAUpPE0PVCNU4o7g/8rF3tutUfBKtkduUIZiWzewTLLfAkLUlnqbylE370ub72uJqrYtBO
7Yn0W1y09yK3KPvOJzkhBehI11jWxF33JEiq8mstDhQn73awI5/SqqAhxVFnBapGR1tdVdd1u+y/
NHw3CsaN4WWyW97DUr7jldMk1Tz8oMtZgZypHjvdBLGjdJ7qj9EnBENXEaTNGObrrAo+DKbGNwfX
UAzMI0y3pba3IiAZNMnYeAR3ZN3Qq6R0h0sMi6CLgRUi8C06t09H6+/81oFKtyJgBh6J4QOXh90D
62EwVCTOUmwrlWumG5Pr6He22Wdpna+zhnuBeREIuy3KNCTc4V7taT1u9YYl0WtTenVZTyRjBwUM
Ebk8GHO8a8BigmQoFjcsE/6zVZFrbR8/cJMDgUhkvuVB4FwmuburzBPk0yp05LCNw0MifjNUfoi4
XfOgvU8V148EEKPHoOF1pjncECv4njV90mWsEfla2CYv0uniwYP3TPtssIcA2XpOjRtJr5p5wgtk
KVJw3Vwsjw9eK1AaggxR3F9JLoq1Vir6Ts8rS25PDTAbbExKgkaENmKGl2mAmd2FEVfp8JUjKWZd
NoPvHakVSAUgOTJDmjYIMkadMBiGzRacKzmH3sdcekmA2OsygM8vtPZ26msyKSb1Qvbe4y18kGfk
2HIwJjeYlqHzrwe8kGAy47rHtktrc+k503u9eUqxzy3n1Xme1MdruItBSas0Or5mnme2E1olKVFc
M2nYKBKj4K3dLIudYj5WCscT71vta76pwQyCVaOCcsF5Y6dFL1CKCZPnyOLd4j731mWIrMMpTWmw
pQDhWAU3YEyR28E3O1UC9rJbveB0PfK+/GQGFm2j+v4cYyzSUVhl/M3ZkRgJ0tfSWsCNQyeZycY1
kx3Kgk8d2Xx1/28SI2olagbyV5L1svG8NcEdILT0JQN78fcHWoxeosHTGCd1VtF0Dw4Vno43gBv/
tdL5jmIZNj5H5nApuPt/l+EIDWgqQ7eOGYB0btOL9AVmg1gUv00LQCXpSqQ1/33cjP6nPNtCDYwx
zCBhsUn7tBPXgZRfqTu9DNjap6pqz5y2MN0j0+P57jkKCCcZ17fhZ2HQFQtouWubG8mF3jojrjt8
qHzoy7yFs3hhoit8WW3k1/jcQrw6kokvivkfyZym80CCuzkQBZ5RD6iI+ViP1XE0ATnT0RbqWkWi
+OKrrNkTILGHvl51HxeRkMAQHH8PLQCCcra5L2UX+lJpKfGZ8rJQHggwoUaIGBy5jbaLC+A0PNkA
qxigdiopiRoWpqi9oifkmU/P6Y5vNcnimb1GrlC9U22S4iFmbEew5Vyglvvh4BsOb/3Z8ad+PFn8
TjqAw/ZYlyEy5d3I/hP9gw1vXGmKHzWyhQXHxxOhD/4PxnWw7ojT/K0hSrF5F+z8D4/GqBHfAdoV
/zQ4WQg/6nt+FokaxVe1R6qWqdqvfSBJS2qgs8SKJIPh2/0ZTBGj3eBFNOrEDz1QG6qKpl1+pSnl
dxDQLDTPuYFHY57XfrNL5aG8iWY+wpOHvAk8/viu3AUumhHnvwqpIzhbN9FxUqhFTVm+/65jm+Hm
IG/GoPDRF2kH06kdDwxE2YQHU+TJLAplgAr/zATEy45AnYqCsEhxfSKXQSKv73GGIk6ZXSS9bl9g
hCFEg501arqzRoXyxKKneeX+e/U29/D5kkoOeX+IBRrXu4mH/oisKdkpyheke7k5KqNoKA5qHGAs
VKP5uGtNWs2vGhS1gGgiZCqmbbpPq5vivR/ntwquZzRPYM/GMfwWhn/r3Kgiwrca+iCkkXS8YXps
y84fqCqoBsklpvmDy+fv31HwsfhyvzUt5Fat/ARP+xOaZoXxYJ+nCqgFlRUDPPoLh9pt8m9xWLO1
M5kS7Ue34L8XZczCkKRj0Zsz2msidtqH6ljZLJm6KacG8iRh5Aki1gSmWc68V+1S0F0CpEVGfJak
ASFQk+aa/l0IPQdpkZzgJbBUo7wd4ut4NJK2QK5quDO4ri27u9up5CQkaJ6D/FxUW6s+Cao4ft70
TdoJ8kJdeQzzCIKp2G9e1I3heNCxtf8k3B84h8fedgCN3E8IYSbi1YtNb89wXkEu4rp6V/C5KW7+
kXNDWav8swrhxGChYCF/T1Nbomcgi0D4Bu5PJLPGhIRoyBIWjU64lxA9WsPGnbkLtkiAZ/6RHuwJ
NTAcbSuc/PqY6GIDkHVssZWYUEE0kfYkJaFk1QFbhcep0Fnbai1knI6dueUwUYo4IXGSNWS55LqX
n30+qcjp64PwTIDPHfh4y4D12NfNBN01+JHFcZSox4uQA2804qVwrXSqqL+bdzc0KINc4QE883/T
/3DSkAvcPL/5D2U65vOwQMfz3bC3grSA+oMUF17l/VBGOdNCK1OVZNCOq9i/fvpcj8NE7iahQZkT
pmMR9tFx7G7DRSjMT7w1RzLCYvYLMVHHfNzhYII5vGAjUYdY96Y2mwH1xTuCCWWSDgKeEkXTshNj
PCA7N/ryWBrzuP5eOMFkrkIcECULmLbr1fwTXngMSUGu8RijA6Qzmegu5+fT47+W1/RWcGnrNQ28
5LyNIGP3JEnlm+wO5g5jkBvG/JAuGFgCfvACVXQzq6ZgjpR7IzQlcpfflLyIVqywSfOg1j7xRG3S
fMMQxkWEU009p5WAuU9Yo32YblxlRkUHsKwdOj+B7RN3GKBzWjEx0iHsCuIBKuJ4LP9p3ucPJUmf
mDaspfsD8+NgRWAFgeBtWx2T6/KCbX3aFVapD1tnmv35RK8+26arBBqcJvM+ya/4gcNSbUvjChiu
8iTKc9IiCsZWDc3OJrEum+GFGRaVVF5DpgenTVLd0ZHYSpe0oJ6aR+QL362LWDwsj94bMC7bHoyO
VyhYsFIawnwUSaEqFIcj3I+tIpcdINDsSyUWubhX1a/t1Ojnmax5V64Rs2uep5rNHNlP1frWij8/
UHNijxYqfbfqm/EgxlErRR7zAaVDph6iXHV9KpA7f9eCN2BHRvcUSG6zF3c3fWI1j0gutQKjgeeb
LgqZI+3tOap7DuBqLFLpiIozoF+k6pRzcUSyjdvJtD1JW+/V+SY6JYnmKNc8mS22TACbcPF4Yx22
3YlOUtlqZUaMjgV4ZBi3c2uXwo9ksyv0NcdNb0f1EWMGsWWah1dYd95nYM4rJ+tsAOqBhv+pBwUf
PKFHMR8ZXnmEPJ5e1ds/WKonsx4mT/z3+qCaw+uDimfpVrAilfiftixOslNCpDrCD4jMAeiiTCwI
UCSotS1iquKxl7MGUCDYMq3ecw6DXMLI1uogTtlm0y3Z7gmlTruLgTzoRZXvw5/OkYwDOStTnxMf
rWpJMg/8LP4xG41m+Py8Fz7iudQxRpnexgQCUYkkBnE7+OOSdeiOmdGWyQdyhWMiG370lQ5EPVM/
0gPFWleScFc8x+twHdHbXBZJ2jqh23yk1ZiGRUxHiFrKQTsfjSQQU1BIPuRMU14s5aFH3zeoKAHg
bg853KqYnYQCg2ojNtvIAHd+usBXp6DgJcgqbGpzSVFppIdpe5nFZb5hRdCszwyvdLkkNvrYADJU
PclWnLToSc04hk0iTGE3pi5AxxZJmhwgv2SIcVw5G4LdOZiVuuFE7TjYy4dL77hGQ5kpfNAYJUVy
JpGuvNc2roZH+OLCpiA6YzyT9UloVwz0Wbys+AychTTMTY8ggW1V0hxdnccJwORBtWlSvmIwhzB2
Dhi99m/x7nCW42lp4OqcKUZTG4I/8u1w7yjR9wpgHzMcoERfYc8QEP8Tn0dcmcvNS5uj18Kdb/f/
wpiO9FN8LdzUXFF7zDffPkewcxuq6cYbXvTuWra8LZkNiQuRDuEGEaIoXGm371YTkJWs0SOflHX1
aadVILvcNZke7g1PLOmW5RDqIQqIe00bWLmixHVPurqzOeZDY/bEBngYWuS/UIBNYodvrqtjsHOC
KGck9ZzzaHr0wuDl2SOgN9M/mlLO/8eBVn8w+PphykXG3Eb/vYfQNpnVk3Dc4DlkKagj/yiYWQWE
on/rd0g4as8sSZk1fxXxJKoOelyu5Y4AgEUKRqf2gzp55k7ppI2gFF3jTHobWQqc2G3/9FCNiAdR
Wn37ilPViHEVtsha9BK18Os9bHdv9TN6itx9Gd6taQ4F79LPy7biKyKihXxImsyBv/xF7QUnt17o
OzHVwInw2UHcLGs83aZXxnlDVJSDzfzixM6311cFsbWHbRKxafYcZSX1aDZeBQMFWVvzNKuIoZ/8
bRgyEdpajq7GvOgVoGA7Un78A9fxnr6dGYM1H8SFifq9c6bicYAL55uPHylIpynbiNN5BxNfQxQj
yEp0wwC3o5QF4fEQw/lt26392gTaMkqKMdm7Jnth2E9soqagi1ZnVwq6E5f1pyupwenlucbGoMdT
UkNm7hboQAjvyPcLWWJv1+eixmAv8I4uCbiiMQds0ExDEkuk3pLNccktzEcFQLGk2dhqIS9Xa5bj
zm2rr93n5BVBqniKkmWoaAWQU2X5+LlipAIlWMNEMRUw7HWSfFCkjcS+23or45Da8jq3VY7PUIO2
hMcz50HDKQ6Boe+LmC/+OEtlCXkipuWJBC22T4UsKjwrv0bcjrqzltTEiZ6cNU9HAu5fet5HDqkI
5gFivqrvsvO47kOIDsPcBP4G67tWEp4xcbYyC47Dqd8itCTwmMp1NDFsz43wZDAnsbQvo/BXr82T
W8Jy3W5WCIotMJIDmnKjVxFMplp6qXZtLFrx8X2GU6+n/eqqkI5cgAxazqPRbkLQSlJHjbpUauE7
+R+6+/YLdd8GC7Fj4nLfO6jDZS9ikDifJavamv8tUDRV2gr2tdyn49qsIBP9GtavzEYJtKnRH83V
g35IS8MeO4IlYzhh4RqjRJz6l17aPK+jNE7i3i7OJzbHwX2eWV5ps6//Fm21niEqx0YVivbjox+f
ep9Kr/6C9QYWPnahsZyYtOvR1E3bgH3WP2rAXb6a6EmKFVZuugdgRJD8hJS4zySwqKLVUOMs/yWc
CDZTKcRmyU01f1+qhrBdmfvNNb/X0DlWXqziTKny95msEYxSPXkfiQ+hjbb+pz4X6+gx5b4jsrtX
Wj9wolUyr6tywXNLHM1pKumvQIQRhX0SPGn33RFS/7DdP1inRwhi3m/mP1ZlYTnFnEMt2IegybOA
M1a8X2rT3Z+Jw5aySgAvnrgeamZf8WzQXWbVJ4DSbI4Svg9yE9B2IHGz8dvItz7fvE2U4mC8qVgB
SKVKuEN6sIf0CQMhHfPs66fNQhUwRlRj/x8l7oS1NxT0yCxxspxqCLVDSlkALjN4llA4dXHk4iAF
/lqbXBce9EDEa6f2CbU+YXoINOcn5CJDjhFnY6BL0aj9tJzYqX5KiB3ZvEpzPiiigt4mj9kSXHmf
ZqnVBPsnE3itpJz1v3EP1enM9O3OxHt6LliGNOtfpJra2hy73SgeOUKha9867OL1vnoCAkUtlsDz
tP66fXs1AMMHM2YaItaYR/Wim5Utg6+aWTkY9mNhQagEPt4fovFA73UodZrZEoI5z4lBQnDS4c4x
xei7xAalni343S0RBnSCGs87febQck1X8MEq8eirFQZeTexdqnNAAzjvHc0LYsJwBjtgnH1FsW1J
XBW2h6+Gk3StdAolout4LJHf8kHUhAtZZVMlZFvdcqWokzP8cWWccjxF+qZBgRWpT02Aq368KE+W
kuRjBHzVtxsMnMFHftG32jC5OBwL9B435WxeQRgUY174woClqOJRxFTusnRNrc4DWLDzcJwMx8YJ
8zbeuyoBCtLx9/fe8hYZvVlXoJ1NKsoF/qAsVsGnm5AnRUJUjy/9kzKPEG4BZWJUUxRDA2lKXxBD
D424JkcVuHLOPFCPhRo9w2h5O1K+xw7Z/Qnqjw2iPlsOrikXTnSFBKwKmIyXEAej/3+AtizbClkh
OW5HTEqAvWTSGHTtaCUBbNnoEOuwZH3RIC+NujY3+DpVTSILRT2cUo/U99h0/ZXXigMeeuCxKHab
+7s/5Fmgk6Qbdgr3ihRP9NVscLlD+ufZ9mJ/3giGnv7VbVdMocymwbY9c+A10LjJFczWA6+iWMb4
1sDOJScQFZQ/Kn13aigez5wGmB6OmEh6h4/UpaQsQzzWk5mUteBlEGLAEsOIkLX0NOP2t9vNv5Wm
5g4zkwRdetbuThpu7JZiqqjyDoo1BGdjUvo1s2h6FL3MMbymTMn/RRiwZT3496bUtSs+S7nlMNPL
YKPUoCrawAvlz/BDbsLgtm2GX4u3AaqWl4BWCGYmmQCtEUs2Adt4XvsNot3V6DBG2SunuG6BtbBL
Y8pLrIR0CxJUv6Lf+8MnkrsklYQeItmP3P/vMOaa0u7o0pPs7pKRz3XJNLHC3jqNBmPAJEbZVtMG
KhRhusPw+hpxrJVEsHclDTR96HT76XGj2V2BJwPwL9cgunDYz4zkNc9mq0s1/SFQdLO0HHTqbaST
Tu9Q4mOkPjuv4R4e6kzQugRQKsBBPkO+N0myZnm2Ru2GM86fdCkzG9l5vhAbtG1OokxdL3P2m9FM
keNLT3xhCJGh8gau6Y+25Lyb6BHEH+lGBK1lIsEbOZ4VTcqv0U9Je+0lOoNIraUV+qKRq7hVbi3y
pfp2QPCh+xi9nK3CYRAYcJ2ydTQu+BSYmBhVdu26KDhrCpT79Pg6JeGx16RxjEq64Au595O8DvWL
Ph0DKitHPd1eGqRyIZBAmTh+x7I/kuom6Oc4Tpa42iy6JZjRLvafhGj+KjsI3ZEO4frMfYL/ZmA7
5ewxcuSCtTf94RJOWyjiyS0cWGtHkKSX8YbdAEJEpZbFB0TCtowyyU5gl9+DoNhjix7VHgYXCTfh
ekPgno3XIJ2k4MDtOzk9oDjydljp0tloaH2MBRj6YzR58etTeEAWlJGOARc7XZShKELIdLuLccYk
YNRbCONG5BT7auZGcJ/AUXvgh+jslXcds4Y3z2/IjrMDqtKSnMcMUJvVABgpuPcKOwoWRyIagK7E
RzALkiZgqBnXb4SGcd5rTZN7uLDclzu7lKTfJaoeHCn9qoGSVtJydVLd4s70m4vo3+zMZyIJmlZB
wMYXnzpG3YKJnkjKDFiLH/FnoRfbts70r3JgkkX+hsKBt6bZkqvb4k+b7bzZ9h3y5OznmnxsDZFD
e9Zt7qhplXvXHzKGL8D5PCkCnXuy5ieX0g8jiQfrL1BLfgAhlqK7uiOg+AXoXIkmJt/xJERkMKYD
7uhY/DzVz+hnxrYBezl0YjqorJYbQLWeOVIFhxD9+jeq7o89gFbFX/f4AYa0W0amqVtd8p3AKO3+
V2FI0wrmI/4KRQ8k6wjXdJavLpO7zuf0agnVCWVGqdurFvPFLhI8cS7WYKOgrKsGRzszsgl7XpFE
RkGxwUJxQCBH6apOESgqQ1ZKtOXQlEVvhewG4KgqFm9/kAZnTgaXY+vIArXb8BRDxzwYOMBq3J7A
f553r1efeKP5uSVBEEqGwt/iKCj4lV8UZnUDhKL+Y/fOdL37XFY1LXyD7vjot4Ztf4U2Qbcm3AQo
gKE8u5SNBAYNoG+xaILCbTiUN+cpEVVpDNpua+8HU/+YjBGOxNtNQXLVFhuKwmlzvoxpQSrcbsoE
J5zJLWMUIytDrTfexXQI03a5kkDByxCOJaoo8GEx+5vTwL9aJTZhZUmQHSYrLSC1l/UOzgY7yIoL
6gUaT3gC8e/uC3FEs5pztoriOPDZLIMrKtaz0nwzXplPOgH6aMWmXmlCMkyRI17dO/v14zyIrf0Q
0PlRqGSbBQBeDvuMCd+732voJaFHS0NjoeSCi9Fv+vAM3mRkK/lrTYhBX1LafamL8qF2nyPfzwzm
6wc5RmLSd7u4jsfy1U+/bPDTH3/Qrs01QNQZJzp5BpsMQWUo6EEVyoGBCPRA2ffd1/4MIz8oypVP
JVlQpRUGliIapyjAwMK9XsN5biCeNx+1cJwYNVOFYeXqhiwbFTRM4Z3oGvYFZ5szv/blve1208wi
TeAAOOfEP9uP+oIICVQH0L6JZhJ48yDPawxlvki40vKtqP1X7koNdS/VbiiP/saon5IJQax5i3eZ
bumAJyHflBeKxVUJzpdI0E9yA9NSTSF6Ms7VrAHQu9x7KmfTpBsCpspcELM5XSB4o3iJkw9tkaH3
abOolsgDfch3r7eHyksI+Lo4N4H4hpbMaEavtkO4JJ4fllkrdePreattbG7KKI6Sjpr3ALuHPh+E
LsywlV280HfnczL+A0pe67weWY/fNKa43+G8vz5Uqd0b/vbgHaihdS4a9kWyF5hwlL1jbblxDsuP
7pEmLPLrNj/kleYSz1vi/wteCr/bzRWDrR+RH9UKKfLr1AUVJJlBkEuJZJ4gZeICbYBgaPmx2hf+
xb+/6iVoqte+F6quay/oCO0q6p+3p6elbM8cKs+zV3xJwdf7uWubMnpek0CD8CL5Xz9wk7HNYjlK
+xK4kXOQkhpftftAxBxQ4vwVh+hayrwDHEk0sJ/Ha6DGI924AhKtEYlJBV5kTdH+5mn7Tc8uScPV
L8n9OSuxwT/3PhV086fyhhTwnGt09tYxU7DRT5Xv3zo/u3iGRd1rZ9sralSFfZSqndMBuIDHvA08
x1gujtb5PqArVzC5pFmFNart0pEOVX6yn55sx/wF1/ErcoYdqWi98xjJ4C/PKWgVwSw2E7IUoc0j
2ENCUoxuD3LayAvOkN+jigk7G6hZJxMlat52BUEMK3eda5Mv7trHmqFMBlsjH4pyzBgVAF5x73Nl
1dMf4dbQNt56J31Kax2/o98qqYxNovGbodnFDjQj6oGoldpyIs+/wZOo8H1f844olBFd7qQhu1Cf
FIyIs8xEohb888+gliUEkkB2YPykO+6D5yAH4kT0/d5PeOVXiyipw0WMi0TctnjIqfGj4CudkVfW
RPj8ZW4GY0YWEKzpUhw2sX77idcRgKNGet4zXjw4se+NYC6cVGPb4cyIPswHRyTmonfGEP9Q/qnW
BFpfOo0CuiwzmGGbfXM0gg5CSE60YqLkT33n8VB32Qs86qy50UG4XoWo8gxZ/Hi6ZxeZTOPKJxyz
p8e2e5PK0VEJEwKdJslL2OpZ8pwarbsxLy9juo8hGVTwPJOHxBkLW8JJwqS7w07bJTUqhMV7lsA/
Bmrsk9ixSjmHZPPv8scDPuag6VQ1zBIxoTZUFxTciu6ehDM9CCsJZCUgos+kmeFwTlWJYFJ8n9Dl
uU286u1iTp3dvG4H+k+Hw27fvoAXG7V/suJINZOuhd5pcKaojLiqwUt64WHZHDx54OmZ8o0im1sC
gPk5FcvxTtEFTWoyeELvlVG5vpk+aPFX/+T7uXn2eCIml2lqixX2KWjlQtwj35uu11HiBUB4Mc4x
WUxMqRItgA/RHbaB7C6x+Y9WLPZEIFpZHG0KxjUlCr0/1SvON/INtq00sMfjkuUJP1nfO2Xypw4l
S+VGBs8/8AP5zbuUImWmJ9oYpCpP8KfSVSvURWG50uyWVSmzY93obgWe22jHPTbJcoppo+DMWjaO
eidUvBWFSXiBHMiAjSX7P3ZvqOC2nmGZrUt24FO+sJoFQjDREKxN2uSjZ5qDzG67UfxA9aMsGO8I
lxbor/p31lsG0wuc9wUmXOL13b0MKgUZhCN2k7vlQ1qkvdGsER4GpBChoUS4MpUSJX5du2cxFYQ5
nMLw8cPBjjkrVeArFyPSukHAToLx+QsF5WIGeVAHhT6Y2U2+6C+F43KBCOBtqPlwyziGrDWslI5i
C5MRZV9yTZoghYc0fMKpwh69r5VioSN2mYpiozapnZjqK6VcYQWxTQEvQtIpuAfdZmy5nkuThQN1
8Ofh4WqcFCEgny9pJ1mhhey+Xn6OKHATHGiIgNzugc/DDD3MeXaKgsbHReszNbnNf+tQFiZni5pt
/saJp/9loNaP4seMZAVlX0nO3x+R81qK/RMFXU1YV8y/gZlzoXNT3zSVWAH0mvrfdZjX7zh9nVeQ
TJVd+LjFTBESL+HQEXBYIFkQBW07zoEVXLtw5mbmt66P6t6SAplI7TVx+pSI/kReB0gUa4d6aCte
n6Vi5KWJJ+lcrFQGgDu/X6VrXQcncs49Q3qLVw7onIhYpNE5WlyHK+d3Fdojca+MwaHi5F7c9SNL
2Y9bYn+t4EHmkq0RD8bO+P1udRuQpoR65iTkN93K5e5Si2OLBiiZaekR5mm6vvDZjtk04BE48a5G
GLVaQIOztVEtBJxUr5lexYCW4gO6wGcedo1EzgMKQ+WXRa5bHRJ5OtG0jZ5xGAoTBv9AzR6avji5
A+m/hGj5Lulo+CCXrTlGWpqCVIQpDggcQE/2bTDTQXBAaNrjSHOgK9q05aXvEv5ipkIqvcLeZqOx
2gPpP5g9TCjlwu/fWoQ93sNxRS8aDXP6Ch49PcssA07wbHI777/2kyTGh8u7Ir2+u+UdKLLA4PaL
7UZDfL0UD9I1r0BR+SgFXDrY7z2ztW+8juwaMSZ/UtgmFHDPEZ8uLwCxWXcaLC3zmyQvTZ9/U7+4
NrcsY7HPy+fxY6IiDMkSNhGfskUYvkanD0Mva9LUcnKIxpjcICsoNF6qwD3fwRAs7vO+1+sOdJi7
MCYEJQ1yjphMuLVHewxVD86wtOcAX6Wz15gP5IoP7m/ZnJJtBNDTMDSqqhT3PY2EgOvpIG2i5sKR
x5nc/Grbt0pFkCbTrwOsFZqy1qR0yE7aRZNLRpNRffVIxas4H0tgXH9i7TlIoydu7j+7ncY5lis7
Y14TFZK997klneEfKz3xkdfXetCO1gU2bxGpJpDxMLmf0J2GDqCuuABY9ilussLKH/q8D8caZc+p
oCHa91W3UiV1u8inEdNr2lv5/47hpv4eOVR8bweAWPqwqk0G2KhXMq9+cA6lAvQhxhukOpP0X/E9
AkcF6Wh1O41BzgzTk9JK3QwcKnitYizJj4QdkBPq4nCVN97inq2Pq2lXLlvaH79uVQ61tdk2OHa4
VssYsxKjKn21vnBG65H87C41IrsC13q5JcQAbPs7Rxam++wYAry3dLuafZiQadYO1bunsfsJD7gT
4KxwULR7UiM0V5ONlbouYJtbICjlWGOQv6OPZlkiA9j4EZK8SlCa5OIbvP/l5VmhJW0ixENdiKfC
zo4BPXyqmRtMMj5y7nGnF4pCMB9dKBS1YfBMk2Ik2P4L4r0s4X0HwmM7IDl7I8UHACGytbuS/bD3
t+olPFXMHE/SnZIP31j9rtV7ArbQd9LuaJgaRKD28+5RJLehKOOh97WOr/+PhvMIjFNyrp9BOAi6
QX3vlh5UxKWNmNtob8FqCNFiwCMW+H/vRWTRYB7oym2kdD/6YWMUya6lWJOVoylf7MWf4rXOxwn1
ir9JHeRTXR6l605oe82CTdHRyshMoj6NShJyH0NPg3VWjJVijpeCKBGZznsuxKDxENMf9QLCNN7o
M+14l9BT2+dBD5X8BgcopSGL4PKbJ0pUvBLaKuIbn8dPVVbCAiLBa+bEynXePXVbFWmiOznOtulw
a4OSPcFf/Y7JqgsmYEQNnLrUEPOTWOZPAnId3vf4upxHZWH63zgZtSVPtY7PsxnBe/PFgeIKK6or
D548Qxy6aZSdeNDx+1JgX8bYDr0ON3dtj6gYRscvBlQf4VO0mFH102RiueoXMS47SA5H822WfBjy
BTHqsiUCCRH7pzCE5KHJdKhaIMXrspJWbDZ/fCeO6q+vPY8IeLHP9hH9OcMyiKeJBuKQh1/3kLSN
nnSJA9gK0jMZqYr413twhJ2AbOBWdU8EHHPeOsmLlrSel8knZ8z94HRXgJ6B123inG/B14p+gysI
LYbJbc0Na4hT042lJif5+BqMC/IYC4h3jo8Cw7WIWljjenrQ0guCKv64IFuzJG+54cGckLyzbfHv
8EfwrXr37A3M3TGxco4wY01IizHuf5xJc+HRhwIAmxm//hwIhPe+2YwO2F1o6irW62nZWJmCp/4B
zH8cBVuroMckN6keqxxchoNSIldffuVVWWJjs91tj2kfWsLN3e2DcpY9b3woQAtJxGaDVlYjTq7d
ofiwTaqbA7+58QYQzFRhXjG7salnc75EJZXzTofJJK1X1Lry1JM8nJTpmtk7X8kJRmqDoplPQelB
6q1/octwaTR5u61sEBtNQFC7ag31Q2ziyRnEBLclHrUCx6tmUe0N2NgrIntbk0EgEnKz1vhKRLXm
qhTH2qggfUgYaiHPDkp3A5ojPC7FKvDV4hDGVxLUUzwqpVZDyjQuvnIdAgFnGmy92W9jZRNV6KqC
fXI9l3VYgnpQ3ctL4RV1BgAp3b2vPqnIr/sEfdWvINA6axJHzyM2LRJxArv3wORsd5vWn6xmJNQk
WZautDl5dpL6GKRBkesk3Po27dE3FUhBmMzWiSov7hyjgoYOutUX6ycFtoIRdgG3PiMUPt5255sm
5Clxs3KGT/+fdXyTEzNMqTJg5kvImQau47yGWP8/gVxpRPeuyWd7o4bVXEoQ7RkiTCXG63CtSSuQ
HiEqiIYpzj/7BVCCL8XRva8xg+7NcvWULCkT551KZfO3Py34IZeXtzhHc3LQdACGsum/OYB3jR9H
EH0DeY7WwPvqcdLPn6bT/UTb85xSmKoei2cCzbeTbig0S3qaUDLQxkxthxfiKMYTnpz9hEcRB/LJ
itfqbbEiiBwaxVzYGSHr14wYrwWWkTXObEGqZ8/9RVtJYaXmvyi4NprZewj0QTYSXyQMPsba7va3
prU4/6DszsWP/f1GmheAmLiCkYZdzdPb/gVYkgajlf34cpaYzoS7meJY+hLz601uME5GdMzAQewC
7iYvFd6q4wIC7DIPu/Gjy1twMet3tTH2MYfzPZGP6fAItsUB9fpvMHvVr5154W3P0x1i0qsugelp
l9D8s6uzvrOxDr4gky9QiMnrq0G8dmYSHYG9tXMP3iaHpbAYRqz7VK5WCPvbNPwKzdBP8ew6mWyF
b3IyZBXDWlEOYlphTwifZMXgkCOxBtlRJDkmD1HmlTm50a+BSZGQNvxG6g2AYiWEV+e24qHigpRB
Bm5cDnbwRrPl9PQzrmnzsK5okqZ2Qj1woNYqQbjR2OoHf7+dqT06cPt0xo7Piu0bpJSEAgAy2ztW
OrHPBPpukTUTSso2WxFks4e8Cxe5qRdo2o2Sakxfmv0TC4/0YZnB8UHEda17h1bKVhmDJRE9HBGS
0E3vIfaHN2nl5MLKhUZizJs9cos7iK63zI54jXGfdCvXh6lr3Bm6/zHdz3FL2RUuU5gIDKMnFtXj
axY97/hVMoBPkbL4NHbFL9R70TvYe6PVvdjZj/IJ1hnJZ4DMHIIAVBy03kjq8AE0pSiDFrtiTNxv
ZUAAcK9IdDJe9jsEH/SYL8VdMph/2xKzg12sO29/Lz4QO1cyyNopGr2x3dgitRDWAGovdd9fP0AQ
te2IcM6I5HdRgIVIVN+hVmUE/vdAf1HDet1P7B6ptCGGbEYNgwwn9WDi1P37iRIf7QMYhHS6Xkjz
//UoxR2WW5EgWIhbpNEUqHq3qH91i57UG7FLpR+a9UqdCJDBS+BlTwGZ56dsfodMO60q8FMdxaRf
dWR9qQWTalHxlB4Vq86gEl5AmQ0nIarG05DC+r1hQGVzbwelFvzM9AFoq58xG+iAKhwpzlNUx/9N
UJXheKwjs8EPI1y0TWYwKcKonmPuFu3HDYl7EMdJOuiTisu0k2Inl7sXm2hUAUVUrdvaP3TpJspR
ywxFJRc0pF4zg1j+gHjBN/1Prt2krNmKxnvZCkH83jkJUY4x7AdFKWw1ynj8KFDq/SnHr78+iwyF
a/oVlOM37dQdQIr6vxOoU2A2bmjoygbZOmPIhnGEiu3rkpEtnAhWkG28NCsy1M5eRfKfH1je/oWk
NWVQDxcz/OKxZWwUIXoenDzHgafBQEp/Ui4vL+9Fqm6HmKvA4ThWS8PJEVQXfjizQ2DNmulGi/wc
1t9bx5wwQsOtol0pjVOziw1UgQMcBH7IScxIKhpEeoXeuyDVClZjq2Gg90sDipDHF6Gpup3N/WhC
FKUPiiM6jqb3Z4bIYZTTnyu8LaNX2koIZvPeEDue1YXwREOqLdMtFNNq7fBMBApnBXvskz75MVgT
sgf0TSiI/lS4TsX5xnfwLgpccYjTXIuO0Fro1jLDhHGKIRfbAj6KQTTO2OwIFl19EJukbnTWHUwW
glVUlS2P0aZ+TFNrBHHXoo8ayok/jpSyJ3N96EDHgm4+XLIgix7uOLmH0Sz+JMOY4/2dAmFX2aNW
TfrXvi4jVYgvafvhm5M/7MNF2UsJs3jBWdeJhOBLhUr2NkQlOvcqgj4xpbZvv4wJJ1GnGTRPR6gx
i8AsXmoR4ANZtm9Gggf8yUXxTcpuDqZ1JIdb7GdyKbUxTKJBsInse6IDFroZcmVw+zypmhCEqiI9
cSjyqdVQA+ibvnaJO1+quQn+HqWifV6WYukNd0HhIRvIBd1oNN2jkucUxFDcqPWDR1sRjGZCFrw5
wcN0k///NuBwcT3Aev28kRrU8pAKI4tD8AxRm9nViY/UUANLJXdujpKUM/Rw3t+3FuM4OWK/LgR0
jVZhUPpwqPvi1OzMIgHxvveIy3tNlk4CxlcmIWCXMznrgHATKICgVIeB9sEgimu3dq5+zk4aJ/p/
tin/1YEoIO90BXa37XXVyB09Pox20Urje5tE781uMgFC/zOXyKseVOBN60e+V4/U4N5KQtQq8qrV
8jXRENA0AzssvybnfDNXzjDp+EqDPN2xZu1xdyLR4WV8nAOQ+GZsTpi0R6roOLYGagzFrxKelORR
WOvxUR08Mbg7BcoNg/i6gP+v01Bl8VMwvjUF4pzedh8153b7+H526848pc2iJnOX0IEJs8BTJEN9
gMT3PXho/Ge7d1kui2axHzK1gKhYZT5D3yt+bV3ph0cim3i625ecDFXa7RBBQHl/66Nbqi62KFi5
G291HZCxN23xg/H3TUaQaJzTz+u/OJ0mdiad++lhKWjteDTrkEg1LOxJDiJUeMYhFwWfMHbSSaPM
ZhfejFPq3/zVeYEKE9lPaFZYopPKadyj2KmiS3+P/LuklBUwPuDWE4M3ZY8bjQZ0frdh3Z5FI/z4
8xKlL4aUVyV/JCsbuUuJWossj1N+oJJ8eRWvU9DKoytj74aL+btdk3x+c5cxxHBr7PrR2IjXcjxa
sRBnJ8UJKwsHmkMpiPd2ZREZcbyC/8q4t2zSC9elFATkv4UxYtYb/BaULrsfuDzvJnETIOVENOTF
YyGwWBiJsP6hCj/yYulkWLoLZPSFw0R6yxkKYMNXH9E2xe1XQffzM7xrGYTbAuPeaYDnlDJM/YFi
D81hmFitmu/eGVLrnS8imz1gG4b+PW57SSuIk9coM4QWNPVU9664qt3ZRDvW02Kl9WPQVjy2J1B7
cxZrOGBq9T0dJJqcqrnLgaYrcO0NIzp18nrCvzqFbbYiagW2to6779sOpqmM20ZEJIx89jKoL5bk
6hjeAYurDtTPKQ2xUPKaGiM5Gi96wsnqHM9il/CYeTu9VMKPJ3Wy8Mrtz83SaBG7rrLVKjcfz5g8
V0PujRQbHfP8n84Xtxs8GbHGkuxUEr6IAyk1LwNgAVa7xnMmdfdxBIA8WHqno30Blflsb7IIW3+2
EPXais1Y0NmlRr8qDsfKCJkcye84Oz940k27xrhVItBWdJwbOF7zO/VltSPb7Um9YLZXYSobH4+G
OXFfmcuEkywCK/zBC2E0a4+Qp4YOjt85gFUq1sPOGj5t6UWe3Dinoyivxk7+A24Nr09vnrGJyznP
8RJKDcQJSly0czvVcpy9+ZVWcsmwRedmTOdfugoXjHCHynNFerWGP0Mk342GJl5AZYNJgyaiXCSz
mjNMFsnQN4QcuaTO+kCYBWg6StBg/9jYqqrsL8zLX7JiUjoqLS+iOxKi2Zgou2gY1a/v6WobxtI7
HQreWtmhQ2pkJdMB/+YrL2hP7bqtDYXVMrUsEhEBcKqCAdUfL4IT9icBz9yjoNK3blmIzyTcASWw
zQUUMvNzaNo8nAlIYvSlXFDFTSacz+HVDLpaEPqR3HAeAKZo0T1DDmt3vBW/qeEdL/jl4r8Bytu3
ky82KaitI5LnKjm1CYuOdLGpmmdL2qZROs3IYtA5ui67Yq/pvYOy1gf1OdwMYBQ9RZTqxCC4hQOD
JK8f/LnGCu51o0Uo7BQsR9wDVfXcOYGasZiG5ZhiV/PcabUNKbc+7oiGsV9Fpnmwt5RdxsRyQxj9
dSG/cvmvoCyQKaIwyDqDXLrdyniEmySeiDLy6TgO/xz5/B1kVQlBoBNbeEFG/biunFuuw0brBbnc
boyRcEt5m0IViNZYDFVFQAJvIfA0Fy6hd99TKwqXy2JkSM5yvqslyZuSzML7tVmqKqyOLU9z14/A
p1gBCvnVW2x6LqFXEayaA11G05MSACEMWDKbw8psel+UqG04+r70JqJqvTPb0XKwDHCWWiwOs2ml
t92f1FBgQ7kLhxKZaLazTQG4lF0XXX0RSjG6ZwdMCICxmyvMbuRnwvi1hpomS7A62+jZ5d/1D1PG
NclvF98lZut6Brxe9qkW2sCWL1T0NCC0uO2Ew/en1MGhHmeJbQ5zPQAJoWlK1BHo/bRRYngCFX9T
btWQQI9DYMGTP/uoOQLz3gwXikb+5OmbUl4rKJggvyF54tu00rAf9d+HgD0tvgbh8OnA1aQmQV0k
c7qW53gfYxCrD0zjbjLEx3PoNhBoOo0ClKGMFrxo8g9DZRGMGFi5+L1vYHr1CJtfLwwWNTAJEGzr
HI/iU7IyJRBVpkbcsVjzIcghUVEtjKyfhWIMu9vQCQbFNKTG6vlwmbbjhJII3hQlz3jsBRakQSxC
pkkGkkZaGT6lxXsgYW9nrQa+xALyExSyCFMG9H315BcAS/zm9PI+Y8Ha5L7hYkivRD/tR6DX7OAN
vlzxG7z8xBuhrqXjMLy+W1063UUnqiWQz0U8To9nlPJrp2mKl/wIMaQ4zgm0Th9lB6xcaPJDDckD
mKaj3tciCGNA074cKVZJ0bL1yMfS9GjeiTyZBw+EaiO4Ozwr0TT3CnDSHvAI3WwuuZWqATOxr/MV
DZxgpkkzmmMLG0EHNuBGo2oj2pcuSietMPr8C66XW8NlB3uBlnf9jWWZHKwx5s8HVIEgU5bHj9CM
YYuKdmulUcnyunmg54BKAkRmLr8zx/DBOazpDZEsO/OgHTwmDdXYeopM/dXwVd6SBxLibr1Y39Z6
WNPGlYF6XUE/ZSssJJd8W2HMiLnBS24H8vfUqHQektQ7c56f4F586026Gf419AA+jnwiPAedOvTy
05FBh4pbj7wLezSqtpU1e2cdw3hFB43+LyvV1lIT3T717kx8P9ShWWX/V33Oq2GUIATyfAfHWSTt
lP99hQvmjDcVrW+pnB0deoWXevr+7moLkJxrKYG5cWVX4LnUVVFKThtn6yc7B9mwCNhDhs0XZDtN
S9QLgGw208GhWtzs2h+3AeK8KGfjyGAHtNogVASaT97g/ktvEXuBRTz0pG9ZUGWIDuS5Vp89NTXE
ipAZ1grK5S6qfFdarJr1i9y6AP0HpMk1j+gfO3uOumzqdYUNbgJ/L4NKFQ8RWgV8CyLapSynyxn7
DNUHx72MVx/ZbqwohA+tE3BUi37GUwXdE+/3Ma3K3aBCBn20kTB5yS9vtq1rK74bO31DXpwEA0eb
sje0Vq223PFaZjFoNecIlG3DrZf8szzgkMBbRAQpRsnHaxN3pgq4peCMKxp5/thrt81N3Vh78Hko
8wcAfhsqyO1ATJmYXQKvrw0G8Ndb8hwJty0xXtZDuuUd79SJI5KZnkmKRvEq3niv8L/u2gpq0CeU
brhev5spgsx7SIwf9L31MqkbrM/z4B2R8NQ/gSJW/n6e21z3KyTPClSWRQof9SNKkl0JHZTsfEcI
iR0WGAPyxnnBEMZAKr5B6h+QPhqPOoBQ1k6AKstraZNp5yeuLZlwGA3pH6uEYqcOXYW5jq+20Xr7
/uufRdlf6vrHTXwSJ/tJyRSdFXpnei2LmZjbhrVc7g+K/qUVYn0hLJAm+iHOEJPBPep7Xxp/CYEd
MKSHO6I3HPGzPLxOkgT9hvIkSPrH0kALDjKJx9EvOpUTP6HiApn93kcEIt6fPLJ661ZtVu+1R+Oi
lFmR6Euy6EoWazY974DwjVB+M2G+lVSyMtQrVPIKENaKtp+ngyyBgjJsSyL7i8pbFPkorQgheyB/
MIJiGgn2na106h4Y/cFraJr+rglS/LJ/1qcergEYO4c03MiX3L5Dc6Mvvubyv61zUW5QFwjeaBam
OAsG0s0FO7QbwwYIvEgQFrIGejsy70mPqLmtnwPkek1fDzDrrphbXwpPn8B1bBqAV/BY83xHZB93
RTraiFtEsKWPaAZaBM99prQIty6uOaML++LDX71vm9/nx84t0VU1JGermrGAdW/dYJMWVLPGXzT7
8//J/OLDEdJ9PUgMFLIxE7sIkt8X/7+gVUju/EnWWM7m9VD8erNQVTFFZkfFwQqY+nNi89BDOsH+
30a5cKbBfvVEJinaa8N5puj8E6esIF8D6uSCG+CSXZhMUFH9NoCHAYtv2CJgdxEqYQ1B4ZvoN4so
aJa2FRhAd1TbnTdg4mnKA9IoDzO3c80oBhrBUoRXGrb495TJjQ7Sm/B/Pp9R/RDDGwd4Dmlbqlj3
27FMoutExfkVOcfTa4KGx/5dtrm+TZ6vSOQuvYnzTHqbSnV2dq46KBMiMY19mitH7R8fVS0QAmqm
mh+EY/NSJxe5ELdSmlZZBzqtAjLjsUrWpDwv+apwSFkRUoKq2pm9cwnhFFCxp5+XXfJJyLJpIYoa
FEvMNH17/zTb7CtD4MymRvHszNj+0+VDrk3KqPtjdxY3PVk0cEpNvvGvRPF4Q38Ge1yQavC90dLz
BU1ZmErq39JMwZxSJHeaQnBtMD7wrqr+8llawQEKf5yuYm49Q12GVZxfdoASkcZBRpoZiS5kRviU
u9fWVZFrWF5FEBJMaQKTIfxYPZ5VKlueMi+q7hwTam7ygM9YcEKbs1uCqj14KOlHJn62NVT19qTZ
f9BnN82++a3ZLxL1BNSCFBZUE9WoxcDEAM73eFQa8mAScCv8FWASDnVNYSb7uZMPhlEj+P5Vjg82
idthpOSBVkRj8+JFGrYF3oyK1a3cMbrxVhQco6inLOWFXp2XkEiVj6lO0xa3t5naJI59wiLk5cYb
/L4bGcsqIvDLR/aVnaHL8fz3KB4lCP5hDNgzyqvzrMZ3JtniF+IX0qFrFqsHJqPgdcHWC79C1YQq
bxI5ZTa7X6d5FwRk2hofE2mcQ2NjbDtfcr9cJtKCL7AvSBfce7nzX4BWSkkboq+uCfGlmtbJ686J
pK32ya6onsDg55MUkzssdMVz90+qIDIGUW8a5WZ4ZLnjmJpLC2u58nSqgxGK0g3pX1Jin4cvseUj
6Kmt+Okz3fm/q7mIEWC6AnBwUaN7KP8gLlAytJAHRUbIIA3Psh4GRBiZoNBV/kiIXqg5mrTFeXrX
vNPTE+WCmhGhr1iY/6WDJYe9GJaLUT8mKXy7JYY4jDlmcTGGbQ73Z1KysYmWvti35zx3W+SbzkLF
cLLTFdmffz2Dfc51e3Qgn33P0p5f+HWOJyH+6EZ+3W3yEOnYFTZ0rFToRIFpCMFqNqGqy6J4YS6w
rTEMA/YNzH5vTsyd77ecZEVNjwARxT+r6HaOOwwyk1K9YHHuMyZRrN7/n8a8xg6tAju5Zb5EEG6a
uSJSXgzRfIuxZBBDExh7gdk0qcdOUz1rkTeUjDY86EQcZl54jAZ+3NqO6Mta4Lv7YxCtLgqv1mr/
TdZGje01uyPNkEF3QmpOasHX/UmgcW8jvoKZO0nxuYcfohQP1oA+TT5GvviHNmJmmS8cJBIpAC4R
iJcn+oljTwfzlY6/PBnBaUYQ4fjgbFfR+W1X44Xs3oAPQ+e1L/yYLewBYTaNG2TWecVwTDlO7YaX
wo3K/o4JMnEflBIdjmdaRR4wlmzMsiusZbeL7gG3jESSjNVt6CFXykHZGYH17tcYGxvKw4E5fA5F
OL0WuoJEfBPta6Q3QskcvMhdNCk8P1MSZbtomGkh5A/J+YLB0dl/BOfWIQBK0/b1bGPx/j+hBwDt
A0WlCeSSecFMPJJwwN12bsglBN/33vzq/bFlBIDsXYRp9VE7SZbnnMmtLWqCfa4FFIRWhDHLxCe/
331C5KjrOMMEvBxNT3QZSVFv52+y0GJj9ZvY/CqI0Mi0CRqlf9tHQn1JjOqBDsxg4lj789LOiIon
2J1BqCTgWmb54eZh2ZJC1BJYXt5posJrCM9O3LJ5lr0NQjcchmMjYiaI2rIFO+ELy90Or1frQIDf
o6k1XxHRbXy9qwc0uSoAQKLIZvm7rOkwrw1WxhRw15UzVHPLCsNyaugQ+x2FNEakbF6KsPs6I2Ct
v4wVXl2v146sjKTqVp6Z7fV0EpUzctiynZNLioAkrcDt+Jp0eCwsncXfcRD+b1CWIHxhvyeAzUn7
hQO86nNJKBlAeXpLrfqKLpaIoKo/9bg93ZAKufIUO46aAyhhq8HtZWFjyJSGtbPu4MfjMiN757g7
7/QmdrersUUlNJSySvxb04LzMuWK6PIM8cdh/2fJHIDNUEVivukmCZW87jkAPCdXjTPSprDbV460
/AUmRC6koef560XylsOnWS+wZA8H9TYJw5bXq1yKhbcmUXySPNic9UMHqvtr7Y4/S3cjeQik4gMO
XBF5gq5LAi9YLNI2FWbztEqTN+zBipTfyJECQ9oBYEFwHsArE0m0iMOl5VIM9zkq9+jVhaPN7OoU
ZqAjo3R7tcImVQ+vZ20M6cWNxdPI7S+Ga2pzWpeiB0c/F6G9gvhWG6NeccN9rYD5mKjGLR6spwiQ
npGVOgjGbkj3MyNM2FM3hwVvGGGgKC77ERigJ5l/zi18S/tZXqspi0zaI3mwiVNluCMTKs/1Ab6m
Zi5/iFly17MZv8ffRXQK9YGS24HNsYChO9ujK9l/p4Gl7T92M6dPWL/PB6Hjm2ufmSP6Gl3iEDFd
Pl4Ucaiy4OLosVxPXxmvJC2F3LheyOabUpl/XvATpEklBxGhsCD3FG4s54kVmnzVekecHESPYyeP
j3L+pbb16BUOR7Qf0M16WvR6OzUQEzV1rle6d/mQ0YP25odoBysxhPdIGqWcVGFBYdmnr9BigBlE
EctQ2d2HN08cwPqToDM7L9rKp50GA9DeQYU4Fvp3Szou9OTB+TWnFvi5lFl1FYObEvKY6MiBw1oF
aNN9r4qAsCaMewGEE9zOA4yN9lcqBfkEA36Lj71vjTDNOq8Cl7Je2SfNbbaYgfREwaANaU4SeTuv
8tDotdXBlY6LAN8hJZwLlTLkaz+j70yB+mdOX+PrRb6fr6e9lHvGuvx3BTycQ3wycx6obCToE7bL
n+QXv/OX/zN8fXlbGsHpFStP+kt4WGQyhFVGM/83UUdmyrz6vJHfi2A3RwKcAcP/PHNRSxcW4NC1
SM6onKrTbnhzidmimtsYoZVST3850N/dqhItKXAOXxA0GaqVVmiu9Ix2SX0auXmWIR3t/ACt1fsx
pk/COBMswE3rQqBKc1ziCoTHzCC+9lbgrfQN6bLRuO4p2mB7OAL1uVrHt534LiRzya9EZWF868gk
J1nla2qNhZHs+R1SnLTzNMBvPZRRuSC6nD1dc+bpEyHFZ+dEXAgKUkRhUG7sfF4cJzvFTAKpPWGJ
UIpyNkqOeu7bfa8ps/JNz24DLNulHqPaGVW3QhU29NUYK6TnHdj3s4W0X+vpGreqEVQ1HA3lza/C
pxOrMaMtSUyyIWOy2nnGwNQ/IIIo1XRQRFwxUSggGUeuuUK6notAgRym17wIR2Hdl74dlvgstMXu
zk4BfnZJYCuCEWOOFdkbZ/XbmLLwKr/HpOyDZV8+EGiq6D0FoI6S+Gm5kDQLNBvdbBkrZ0fbwl5n
1J9ubTeoN3hmRYltZvr8EreM5J7cSm/ZOAOiGIHA2lZ9hNvDIrRA8nIG1L60aN1qHFsZMY4tdrvV
Uzp2+Fsl8ul8belmDhfQLNFmjAaoZcVDenquqAjH2fu1Er4Ec5YIRWZjfZyeoZtqlt5sE67svGQR
b1w4rbh+92aIi6yoVx3DH+iCLnSVjLi2OTrCXAT2ArHydHel/3Fu+S2GfXGps+VzMt4fORVY+wSm
FJJZiXAUMjKg1JR73IviUpgUMHC/a6/h1VXTvqym/52rAooVNKfPanA3Pl3RnrLxiqT3Q+DWr82P
9DZ7rXfVN8g8Loq8u+r92HQyR2XsgZk758GE4jWg5AussQd7FJWKm7lVrsxSYjbOc43XwH8Olb71
CZiLXP4UgkvfjaD8loQ/P5FXpl+sCGiOBWNePpSQbHKLJo4insWj5kR9o6NE8UMuRZthFs6GJAvG
U/opGlk+6tu7WHLqG8nTIjQorH5NnvrAUPv+R7h/9Zamcb0LBW4akRHCESTKnaL+YGMB6l8q6uHF
EoFKDBSAa9sgitNPnQDH85v3BrW8KYb+1ljV2pbkjrIDSM7ceSkFTKepzc6Ac2jdZs5g4IQwmmmo
y9ys6azwte1KlBf2lKKzwqBkUsLdpR2nMRP/M28IQ67d7Lk3a9VUhNTkjZqPQxutcuN8UWRivc1f
WNS6ZkEUNN2IRs6Dqom4rfWjoVlY18GQrUceXfEDw19wH5AbivD0qkFezvgNSlkBLU9vBnt+gtTS
JFounFRZ/z0HEn7X3/qKCqLJOoS3J0IIg2BLQgt9GMD1JZMdUQrTw05nVyW8J8bNYjL6LRTFuFlq
1QC3IuTEKNfKBTR3i+gmFWWxN+W/p7/C42IQtW8EAWCBmw206G5WUydLAOF/ikncQtCxFmxWgkco
YDU+7KNDkFES/380hekoqaux5NJsGYE9RaybHGTDM+L/JqR35jEz4XsvPOI1kb/yBb9INH+JGjiS
wFojD60PzaSHAbWYuvixz8dL+8Hmp8M3nsevi1vWeNf9/Itnkiqzw2ry2KfN7eJ5yYOSWeQp6zos
Ng4mMAIe8MDy1qEfecHCUyLFd5jO4TdOKS+N6VFlXpTbHxcyeL0czw2K30Cq/vXDAQYUrk/ewzhC
Kd3WWN2abp6hh/kG0UTg1cbjK9zlJdjDstVART6yk3Q690HCyk+RgtHw/Cg0zueN7n2g3BwVGlly
7Xm6lhCkJciGE4Dwx/QN0fVRG/zhpumokhug33PfWv4R7wJP7eiw1Oz7LkqrHv8B0mlbA08mZ/Zp
p8qB43VIeroEstYLUXVT/wAofUTaas+OspgZTVTYMtQYTUvouMdmQyTKk9vsahdzcQZTn5AVNHeP
v1rzw3s8jzT0V6LYyaPn91RVrLblShCxX3QNoESbnnDeWVPGiq34FCFRdej3HYkS/SFLneOMGFg3
dvccHpRQsZfGckvkLsYzMqHYEFluFl2Hwn+yKgPaeoqrSvkXjWWBjTYdv8me/ir3psEbEKXGQdBK
qwqXgNYb/9bD10mgnk1YxuBrx99Ul3Pe7ZMphDr7vqUSAWa/+eaaE3YlAE00TdjexZnFkjQ2/SpC
4P3VOYh/XNL3iKouHYDd4xYXtDTwf1n+BxtwZfDq+7xd9YjR9LbXqKmThY5AFDpI7WD9zibfBZra
ip2w7qSKFx+EMJXB0nQiaN/O2mB1bsXwvub3j6jUP8rKY46t7C35AKL0jP8hZgc27qIbJ50i5ETG
kYAqkdELalBq54Vc48yuYqdgavFz4+9pw7SMUGKaHNO7aJfqZuQF7kZwXfBdj9g3s7nbHkICGuy8
T+QciBI+fEgFpfgRXExLoxMbiZsiFTqKc6ZnnTYOaC3nRfmL3Qnx/G8oZKNN87ebkHTz3UxVELdk
oRzH7MlyGw9ApdmtUr9zF2JRid8M6TgPPX7McnRXo8uYVUIVrNRVpFf5zXN2o3aNsnd2LN/iGZ/5
27cOAFLlPImDYHiy+FtSFlu41ZIwka9BNzKf+05Fnf9d45HrQpHc16F6pzbAsDDr0yiIX4x+J8Ki
7J0xYS7dfBPa0av9B1FkBpfJskMTjIC545Kk6jfhTC4S8gUOAGIJQ5M2nXOebsBsg4yxjGB/dLUu
SUWgHgDdpHy6g7Bq6pYXXvg/ulzYY2JOcps+XSHHapGPh/s/vAuEsIqHQ8Rp6GFzaaE/+7q1uhaY
Insne5tt0e3NWMUsd1kLpGPtnpmQKErhWpQmTrGOdzfzbaWlc3X0Y1U1PbpYoGGlToJPYRm7VEbI
KOmCB+pSctVWVkaMJlDIaXB5l6rOsOj3nvAhSL6V3Gb6icahqFCvupEWElgAo4d6WUEXq+MaZyeL
frqj1wk8FPuSgSHulwCGiBWaPOrB3JSJM0tGz/55Hi7Ljdh9K8vzNitYZ98xgxrE/+IijFCgY9ar
dwZXCbT7Aez9EkerxEKIauYYef3/9u6hjRNCyXKhbdBWc+O00gogkBKwYIA2+YYnjBAYpjAZKYt6
9dFUdFw1XI9WoUa2pBEwcWy0K0m9haMCM+eLhWc2/iTkj9OIs22rYtB3ecvPUGeP/GKxPbX1Ztay
j86V7dqG6R5Ke0ZuCmAEyZl/+jb4M/H1YV7hvN4sY7h42eC4Bah2IepfA8Ql+iKoIMl+EOLb+t3i
d0cU+b2vDSLwfZLgv2ayCDS3O2CqTMBJGSVh8OSMiOy11tP1FRfHANIV5AdC/eMwZQzHh3qrJCqk
glCa43rX2PgSubibmMtfx4DulL9vUgd/FKxtn5VhO5E2I5A9DC7poduhoF0wNL+CV7ECeBeLrdSp
NkphrLh3D80vu/z5h0mzxuzmEaQ3Bt5j7SnbwDhqeEDgtc+QZNRgPdCUssXyGMm9lkhDVX8SoOg+
8wjvncD5e2Zx6z1c8x7daIR3SzQX/DnNeQ9R0vRpemzrl8mi1evgyt6o5TlfK3s7KBdR8cuKxrlZ
XIMn+uNUvNlrmlxAZ9oUhJbcWestcuJU9nvv+ANlAdWQtknhe3IgkmhR77EtA0gMDHqvj1pmHOnZ
ZtI/K34kMtGEPaIY96TKQDaHgvvgmJEazYfXSkyDkGOuP1I/vHsHpMB9WbLlFuf4Ze6Oa1O5qNuW
2YhssG8+7zTQ/7bcafp32xEZszjhTVEdiJf1uFAW+Mz3h6qnLNemio3v/Gjt6xbYvYBVbAilth8n
5U9JyCXfWg9qusyjnKgT92pbkBosdIV+cCATef3XoG9yZBfsfickTYbo7VOAm6j0J+ywxLeBv2BY
lAKJzHPcLmsXO9MKyUxLejHb+VDT+oyNM0b+f/ecWwNtaLEGDxAmyelwYkxfWFYnPbDuZF/e/H7U
eizyvmf37tldLTduUHreWSl2HjwA5zvqAQKG2fM92T81VISPqi78De0fhoTVjCsz8NyVxEgIcpTD
X/YGmt7pUSi2tWN0CHCFCFFCbHmlGwCYaZDrb9YjsguhzFTeQBwAdQO6piz3pN+mMQf6+ZA+TbGS
O5Au4pBP4Mbr7uUyKukUfzu+Ve/yjXtEUxZasxLqcBtxeyQi6gecUedUGsivcfO4jzp+VsvlwYFC
kUXVh6IVH5a5AezbeCmJeIiWaw2Qe28n6Y1rKhpFrBLY9gtWPCVYusyleNwDwaPK+F8iVYiNuR0a
qVuDK80MNfi27ibk37MDgP029lGeAotDpn/P6jjhNnSMQcp5mi6ykbtEZ6F4UQnn8+uUeImfBSbS
IGj6WaclwiCHyrNb/TnM1uyBHeStuAGCdlGJbNZ3t8OQxNHKMFIdUrz+XfRMBXgJwDF4tVqknf9B
QP73cfCpJEBv8b9M7eQA/qMg2T8ZNXLBBcSMsENiB2cvKmcKKiXRIHzr+w7PtroUFCIe08eMIffI
9AFC/kzxnbWOvC6BXcnRb8agl3Pp5yBVXc9wsIjQfAoFPZqAxVh7LlMsYJlPqNO/e3n8G39NcfSG
rIK10+pRFz5aEoj/qJ2Qj4Ly1UQ8QDksjkHkw5m3FNCQmK1ZuryaVmLthE6JAYCV/FrO8zvE1v0B
EgTRlhkhpRd3eBdnm5IBtDEI7rkf+Uon/dbJGupiWlR3ot4PnQXbCFxP9Ac9mTLPXHWPPptyVB5E
HbXZa4VLA5ND2vve8lJ369oDU+s792Xjd7LS9QYHsM/Q9nUeFBruFeNcbqX4DeixD+l4tE4SDel5
vC2X/6K2Kq/BI5ql/frYAzOCMhqY1voE6YrZhBCawLWEdLm7MI/f8gq/FaaIrHz9S8UhcDEE72tn
zNq7TNGavOZPlvXqnN8TlI1WGNXKlwtsKOTmrsK0b7iLXg1apdH8+QKGq7XI1WMrio6Jskt0eXho
RF+Nu+eHX+2OYHpzz2NScxAh4rxdLmKIDj4npb7R3TafYwQF+nE3Y/0OiKyELgMddORM0fcqvO7h
laK4vvoUACMbFeHD+P7kcYfYzwuxd5N68enQ2ZQUgRAldWwPkl05yITwJDjKpVrbPiaRRgVxwudj
mVIYd0R5FgRrwuBJ1HUvPCX93bhEHlBWEOC74JdWO/gAkfV1NswpIYYIX5yFGOOrhH33/MFF3Oc2
oVh+nBgVaW4ygTfYDaA+paNxlZ8xGfyxthxAZNEHCA7qVl8Dk953OYMzeeAASM+xJs3HhbSp5E+s
yg3ek9FuERm0/LTs+uW8gmW3W+SvzSbVxYhtGwY+3ShITEXyRD048PU2Kuddq4SmSC5Wqsi4z6pB
FXsIa3dKhpcN8tXQAKs0e8TRVa+lv8jaSnflOm0NlWbBB+o4EsPe5z9AW+UAT/aNKieRO7z/wQ2b
P0N+epE5dwtZr3/PTV0NwST3EkCPae19ODJYWzq/fYjqOmDkKYkQ+O/RBO/Wlnwo5aH3wNA1wAK4
2L/3D26NMjLj3g5+4wM9Fh5sYRAWxjOoL7OQ4UK60WuaAxIMt6MKNKfWpcoU1lF9nj4yJRstuXi8
ljiVX6PyGYwZ6UPK9i49sqm6NVtmlKysP+zMAPUkHSbKJvGbeIt4VQwHQjeiO6fJdll3ATED/yIV
cTxcEa7uRhovTH411Sai7JjwfUoFGn21Od8VyZsboWKulHCzr/0wKLJMubXMvbrqUVeMr9wCJ0xf
Jv/yHhlnVbWvXutuqdsADRdDWGJcfnGFryQQgVFg0Wv1sn+WLDm4niKM1y1A+Va/flakGxlP//DE
ZbG3z0KK1yO5qNQsZBhy1Ipd63koZyF8wzaOsObOVC9z0oREk9icIPGmnLZT0hb7sY3vPUiB2d8Z
JzKg+LXzhjK7m25m5FfQRt1Z3EeNG+OTPrxhK77A8avJCDFoQC4oqwn3NYnGGLsCEp4K5Fpf0KjD
eMBoWx9SsDRCcB1gl3JS14QSP7vSk2yTOaS2KrKsgnw9UsS+OA0SO8K0CVIaY4OaAfMck/3S3aWj
luFisJn6SsXwJ6a2h1Rmo3H7qz5hAPxBdwwDWCFP2HbtN3H+I61tPlFbj8Lz0fIDY5vGK92upJSe
5LQlyvm2B4TQ/Sb54KatE66Wd176k2zLUnalQY/PF+dan+hSjA3BkXiINZtG8m4Di56q5IJsfLva
gFhNJGXS7fVx17mnMYVFL3b17jH8OYm2k6FnFifh5h1MUB34t/Z7nrsnEfjHwIlD1p302+TiEgAD
fzzsRFEEQm8KpO9nDe7OzIfALDDmjNOuWTp7TvVi4QhcY/etvTZciNTs28SiGC9d71TDYRy0zW1f
TSDn87lgktEqoyI1z2V3J1S7rW6JfXSeGQN5/gLSJj2A0JTG1C7dspQF+7u0BE+W4jyyRtgkZ9ch
iFNEbVriYFFkfzlRMYksEMrDieRMmqhNls3Rq4iSssrtOoJutT9wlNcwgrgbfyjScoGgV5+6hgUv
sXyLffnR8i0+zKqpiQkun2qPGUi0uWrnItANR+gtOn+RU0kOjL1I5si4cc84XrIMRJelVQrg9qwq
xlpvXh5EvI24DOdXjhojgSzu4BU1GrxAbqIXzK6x6zeivCAbOucvrAvoJt5NsvOqitvkp2eQMohj
2s/6EAWaocRVZQ1VkXmQLPx1+qV37Y7FnLfGKShLzNwo9oi1zNmcNQnzh0/MnfSv3nCIshvnQBsf
hcykn8J7dhSYgVH59ntgp0knCvyrOwjrpWKQsUSXEs8ACqYhbRuQRuyUTboXcRxpS9WcKB1CT0O4
3RU8h8D1pkEW0JRn2PTGVZfEgU/z2t1VNuk/aXw5W/LCchMtHETPpZTQmWDqO9Ursdt5RcxdKGFj
yfZEH1TMgObrKcu1jro79F9D4yX0dIjSGBe+qp6nul7NeLorSWOfz7eLGyT4ut2tR85ZuUEVG9iF
MXDnKGKkvKo6AnSYWXmlSVuasOk+crLUs1Jdi6/leXuaSZ6J1L4FBWuXriEXubWa5wSSu9foI+CF
G5PSQIcCtp7HQkOBUnxSebBMtMneK75ITt6JJrGjlUILzQve8djmxb2M6fZwqJNLZ7ddm8BWro/E
7BNJIu1NbgB6eprd7DtH7zuj/cNo16yzTVItVSODUyJ6HxoE5gQgUM7af6Ml9fBjd21gb2foVrsD
6ZZ7S36E252FrdXFU0r0GwkmpFOd4f25pze+a3S00Cx4W4USjDdjn9OgoUOBpJ3cM+UXDMQfBVup
XkUebt7JbqYW+ONbx2TsZHBa3py0jOfBFM/VEB6wPgOiMmHWzqyVDWKA84B5CCkT65RbR1iO4nYG
iJZeeVTLWAwwv5ivuzxx3/fi2qZZZSh5snQSZ6C4wSs/VqXGS38rWuf9RekAUmKbM6lD0qHcnFL+
r9f2qRlc5KjXw/jD6tUVxuUV6YswEhPsdSXxT1FeV7bReyqbXT0a9EskabIyY0RIcnRdyWAwbxxy
f/ojvip9ATMieB6FbZvs+W0DY7jJDz9ypAyTzBHgYTJblJaJFx333bkPGADOXSnNrVJyMDVY2t0n
N5t4p/HapUX0BWnLoBbVlUzObeDpp3P+tPKBweFaE8voQDgO9+L/KXj1zCW1GNdXdp32KjltG7BX
86xoBc2l+Fq9yC+qn87wIhN8AIXCTyIs0N0n87gSuUkZKFZ3CaPg8hSnxQtIQ5Ijw0oFUrFW4wHi
YTBjO+qVN7y4KjW0QCwPgozGdtyKmL1dw33qAt269IUfXuAsxtCIHNhzaEI9iZzXAN7DHgLKPRAv
lQ0jMLhnVV4HNdyRRKsyV8IsmhpIUzs9jigCN/Tau+sCw8fMZ1PTM75YYNlXUJHjA5d/GqpKCGRS
FmHZ4nkGRh0F8g9hXb0RTyTXqgOCiJprjW/5arOnoqAiHLTYvuEheT7iYGDpxl61WIW2+C6rKqJM
J/HN0XMioii16UJTrk57tTEI7ggyBoCCO7Z42tb1S7nqN2dmHDS0lqEia9yhx4qfeSB8WlldBk6X
rSKHnHezJMZeeKXYdEYU+tZ+/FKBWdlUgDXCdF5bZ2U6bGrwJrziELXXuGn8UlVCKA6szBzq92+3
uaA/IIY5TO5sd1I/V9aXcvENypQwaXMmCK6tAX/43D3smNN4CiWCoX6Ckr99fO8N0AZlwq0hfyNK
a/35zlx9BV8Mh+wy2tgHJlCFatBmA+sUVDkAoCJ4Z8z7dLhC1xwrdJrLzZ8ea704TinLcMrn0Gxe
iVJUTSkb6gDF0DAuBnP+nh52BRXGlbO+FLn9hl7miZSw3jKNwHGO/CCuYwirkKVaWTMLcqsyNnCQ
FRfSAxe7F5/OiWD7SFM8dU9bA13ElYtoBbG6vlSfjE9p4TAqYnqmov1Sa90VaZMyZW9BD1bkNeTv
7sTSHkCFj4FmdtjPo5fUWqRNy0ZeAXXhTEOq13ipVESqzsLuAt2NGSe1hjYJuFX+lozF6HlE++MZ
tB1WBfqvnxwSF0XN5Ac36zva11WXLyf2zsjNc8Xot8y7TdxPvgGiA+JARPh5JDrigRcW1rEg3pjb
8UaTs+w8d33f+AnhkBoDyGmEgF6xc2R3a3+jE9iTzLuLFfIWqcleZ7hIwsD3QybS0ciAGT+derBS
M6J6eLGn9pDfD+HS2kag4+uVlY7MFf+tk1akIe3q8XMbS7OoyB/oAumUHJQUcsdBi6IhbVVrYcX4
IaerKOhEDMMcOS+ZC/37LnasCLPTiV3chZMbTjsa2u0rEznP3CrU5cpism5VtFUi6vhxBosNdRaR
0h8KXqyJ0UmqgbuMHoW1oKu/YosDpfgxgvL+lBLvB0NN0LC7BXQUx6ncPc9KMZYQKTvJYuh6wydD
10hSS7HIFDZcBa5ebjIaBesMbTOXp5bblNzlrbqVhOAgPQabIsCS87Jh9lq2ivC6wsAUjHeixYXJ
mjVhEuKnyYuKhJk260rstkV4CeyEl095SEVsDXmAx3Bf4hbdq7uwWYA4E3Qd4lZhXjYrY3QnVVE+
+GrrUsiq/Hewt37KiURyTHGr+e0Jx7hskwO25AIucZNLj4stXPNcsgCXF9AU9yFZr7gWwCV09646
Tn9LCMOYRiM+TPWIeyUcc46tQFVUU12/k72EdmMx7W8OuXaO29mN2Elsk0Yp4u9fBM8tg1KNJpVc
R07zV8xLth0UljqIWpNrHnwDZxG+D6J2z8dP5arfnkFlZwUxwVeiH22OK2dmGRSeTwA5DuCF7TJz
pIJ8DSyeJOkMyRYe08TpyqDU75mv7D++9hYCWOlENwAtr/Qe8YcYz14lLCZtuBqBSDkektHatMgI
RAcokTCKNkXCeEde1XBXWaJKqhPHoXbk7w7cGdJZp4I5eo6V/krQSrlkPzAxOfM1GHkKC1VCyb6j
zplNPWBg31dDB2hN0TBZvfI3tn/NqcSItSmz/w1A8CLBYaxzsbQNai7Iv2RyYqCFxpT3NaP4K8Pv
tsGVa3HOmi9PCBLIKshzSRn6YOR2Iab+NvhxAe3PrlBq0BWdwzn1Hlya2nu+DuvrhDwerGQ+maNz
NcaeGnxuHkibgB/mqQ7d0OxhYizwtwiSGImbXuI77Mx9XA02gnNJ1ZV/s4kSQciB+QRk5dfkjSNv
meniOOOZ4aJltaEwVtF908qo3/67H17anHPUwa1Bj4H4VVIQhoJ9jBQ0UrJBFUHRh9OE0ez08cAb
F//GbeeIOQiBi1mh+TPVIhk3brDAkkN1sbPtwUDmFja5uZTO7v+DJtQerMAdQ0HkE2SsHzMkXC8f
srx6mEvsbyjRv1Dyv+Ww8oI7mbN6dKRIXDf06gnirkMXbR6D63zGSHpARfAFgxK06Nrw49AbrmWV
XCqKrGKGo00EGgVrov8MY2bdaFz8uVjJ0UhPnMA/bGN1VtrkNkzlHA5umoritlTIWoNSYWJBWSeo
tp3KF6Wqhzk+Gg930njPIz/qknmn/tLOIMXQsx2xH1RxClqWUvvW61kRqy4LE0pHMLa0iJKYq1io
H9Y7MXkXeLrpKKXg294+EUsNwDsg0C01Raq/WvroL2Xi64rbsXb+PyFDbFAW1ms902hItVOdv5gr
rx6R0a9kSEJuNUxSh+9z1iMsq5SLbrleX+yuSuT8SP1F0to2rQNZRjOu8oCj37XdlndFrJHDKJlh
6LE49YCBUjOarA2+xkPNOSfau063zBfLt7woBk4hs8FT4RhOL9egRY/KAYpu247LHU33eRgbT5s8
yuIWGe3wkO80E8ymCpzY3DBBMxa/PZ0AlW51wNO2HtW6/pkFNhAhe7RQYsZwUaLDE0j3slY+vX6F
vjJQspYxaXmR0qIQU3JHCMsrk4N2f8RXiSxSIJAnnSy6haw3GEMGMUx0jToFlQCw17KRhmXbrOln
HNCMQwSaXdcpbY0n2tJUIS+46FpgG9ZxXmdy5NUhemyp7d28xGvU6GuBLR81MbcLxLAD8UiIUpgD
X0MO0ZzkY2M+exXLbLQOyWjZ4iJkOl6fgpFbxnnl8ktqYOzg44uJstEkBtQl6t8vPPcXHMUARZKO
9UCUt78j7Z01WV8LZAwYZUxmkVsgB8VUSuxXptPBJaHIVoecKcX7SDnrzrg07B3xFD/g5sL9h1E4
7Bn+yec0NscltymO6En0Ssee/JTXTM53gWDUHTXvL17xhCZrUR92Sm8DevM/vgkYZYfZqX8M2pvo
67Jpy0T+FJRDLg/OiLKyfMG9l8RErNyIzMgLLWRPG2cfOKV3BuXT1KeYd7X+6uwSJzfzOeFf+fGG
/N4H25/cysLsDYDwRuKSdug7ny8KMpO/mJGKTR827AA3vAESo9T/+GEJHU3HNXLu+5Frh3ICeHSx
O6f7uUrhx6jDzYzz0hb58+haUk6sv94SPmT3w9wv8CZ9zvCIpA68zepjPgcbNZ72wowfqqvwlZke
nWG9HPzkPIrixPSjmYcTkaGpKr3Dv+/LrJ17Zra5yEMgVLrXF11YLFFERr2ZwLJHg25l6hmQNk3b
OuWl3jN4WaYXdxETq3gzBIVAvTtgFbJbLVqHd3GQGf5ET1J1y2V4Qod33Mm0v7H/TEd0GsCzdyhn
u1JiRVhrJ85uNmkPJqo8UHy5f/RuNaPp88ZuVg/ckq8AWVV62fcTqSDxgdFcgyPoVrcLc5SBL3XT
JRziPBNIzGzvmfLp45HcR5GjtCgIUTScvMn6a8qC4ZzpCN50ETDRbeU4WxxKEExFrd8zhG8ZN03m
JD1IgIepqe8/nqOIzDrBkYN8TstkythV80Pk3V1qUkbHCG1Nx74YeMm6NgsdnFgyfi7NzDuq8hT4
yOwxdSWmhsb8yzfmJrIsyhA+qUlchJe+X/MOtiXkTQlqBZ5s+AMuJLt+vx0BXIwMsfmOgh1PKTLB
h+1oZjZDhz4sR06ZkGzH8e11syj/igbcUjeIvN42DrgHe/K9T9vwUxQYS6B5uMk8vZ/L/GfiAgr0
F3D+P00SKzSqGPpc33xP0yApkiQD+5PMBUXJ0yfpbKeVsXrX9gyoGyrL6Ar133Y+ftpNnIP8T9hK
ilatyoYaUeMa4ODh/q9IYx8BAR68yjCS40YiGovWI7tYI4zD6MBE0KNEnXPUtrm6L4MgS835+v56
cyFRNNXyMniLeP2ixyh0q9Ns8QKNwIawibiiT4Q6KXebaP9jhHO3cNiBVJU0ktU+4iZLs1MB1QxL
dRdzWDbBhCs2mBddWms7+emDnZte6NsRu+/5KnkKNskARghaAr8jcqYVoxbzWmGAMLsSWcrWcwvz
hUmIFV39IeP3lTNAKbqpBHeNa9+AsmSam8+Og98xenlEAj2IYbMyQGaXoLub8AIA3q27R/ykg4to
V89TmAwrnOXgnT9USdxZr1/EXsxCZNEGPmQH/1p3YivRYAY49HpcIasOVrnOxzllVCWlWwBttyZS
Q/55kR65MH+O6OGhR48oVtPvMzsywt3S7S7GUg/qGjBSC1n1Arp7MJSARXF7AGoSl/jIrHdAgCoJ
j6b5syACoMdSzhjQ7MjYFJT1SJBYzPiX/DMXGY0dZdW99Kr6qY6ZTRFCZkjMkCrJX2uwdkJFIcSJ
cbinXgOkyShTgGQj/z382Mn08DXhydLCxxLZSw924uSwhY0sNYeZpKHigbgV4Eo55KQR3uccBhBO
2Dc245Aj8u2WhMZwuvqEPId3zY56FgZFtTQec8kIlzM2k+JCCGRuwrHUY1vM7dNuQIMFGzWQCV+m
cJviChifKN7gPmTZUqAxTLwnBalN6umrJvGs91JmT6q6hvOTjkYr85qT1zuARg0Bjz+PjjqTMB35
FQaWGklnh2uIjRCFoXtVmNWJ4CU2V68/RJK5uSmnuix5NeZyU4Dr1Ux9UtGLbejVPW+Ck/z/HZ2s
Ugvb5AdcU9SSYUK7AytKsY5/l8rfLEK6DHbo1ESzqp2Xxz4859+nr0A8twS6Y3kRDu68LgSKdJ+5
4jcevnD0BdKVJv+Vptlo0ZE5zyGQEiijKeP84LQxkf4/FF//+TouwmVwJcK7uHwVkzoG7p/wWKuU
+aSJWsPFiaevbOgAwT5O4naydGTd9Bph//hdaQuBIoX9hDEjKD+m/0gN5yBDARCps+ZRknl+Of0b
RIcs4QLh9Vti5fpaD16CPcLaENEzP65K39XxhRp483SIPP70OUeB2gcpxWpVvyFA5lH3+3NEzLnO
YlUyoubNxTfYksYRU8HWuYZcBOTuEOFmSdJonq/s+ZOQwmHkU7zSrpvqButyzVDMXTVXtyg5hVwS
sD6XljALD9LEYWqVMdSX6oG/nVTq43Kl0a2WLdQA93yRaO9iMZvKGbxo2nFm/XCxAKN/5Y3mimy/
5wJjKxelvor5qa+zhLR1L5w5Fxl1w7/vQIfuk0Rkdz8V31EfvrxR1WrDbh+4/I5t+gsI+FNXbWTX
WXMN7gySuv4KILHDp8mL56gt2n6I2z8d/Bc8h8+HWyMRxPtGU45jeDZ8PTAF+IgN68Lvc6OoA+2I
oJafVOv7OfY24VaVe8ftlK+rg4KvFLHgDXoXw+eJCEFi85RLPsfsNodRu5FWqVubM2MjeOlTWbii
ChaYnrQI5XHrN0ZYFfq5tKcCQuPGVeDPRIazJvW3uSVP2AVkGGhm0NH1YbNPWE+NIh6Prs4AhDPU
QoqIT/uW3ePBtQfUIZ8jTTuafmUahwNhqlboQGpMIyjMCVbfg0NYZm80eziFIht8SNDVAxfQZBSN
910ZrJ6MA9IuvwV3yuAab9pmnZl/yTP+1CgY8nsE1yvq1LUlgOsBjy5HN9hVwTjODgdClE4DdhoH
0iJe4vupZJSHvzVcsh/vaXJvGHv/Hkn/qtfu/zUFyKVFVhKlze+qk3YuQMY6LkvnkE8MrlgU0DhO
HCDNDNNYHAQ4GvZlHmeG9Apw7Eo6+rjJMMdhDLqmP5Z9c6RQIrRoZSPtVMNRJ9ny1owgpp7LmckN
19lLjQajrkzFKXENebxizcJQhOanmAGszQ05gP/k54MXOTmFoKGmJOMX/Zj8XzERHm9ttBp4U4bN
dO6zrkkcnywXppVUaXS5REXI/EaC0sa/bE5zxVbABmlQ50Q0elpCZyVzFbwvVXop1tHGPqKOwHIW
BsK9oqLx3NjMen8vlTKwQYYjZ7dyJVF5lMRbThCRzKB3GZM34/0Qs1wJaKDo6sU2UGpby5xMl6ON
nDnihQG9ZxhwqWCrmc2P7RLshZwx0h52rIorXHS+l1INWPVUFtBfY4Blk/HbKc7Yclscjy2fPlIT
DxV5Xc4wyVoJIHcD1UlTlaiDslKEjK2k3EmNPGEHrI5Oh5NAozday7644+ildkxNjFAP6hxZWgzv
3PuMYxBQA0TDkskc3XYAoFgmmLIERCU/9EKpGBTxfcdfNpuatwGioYVrP5p8lOwxEfE11TsdrPOX
wkRqbm6sNNCUW1UU51F6S+ylk9455l+++uMX0Ds8GbTeZUXvRpYbot8UZtGQfbarMfLcwcPmoW6t
8dqmOQB4E8pMesIqbAvGMArJ0t12lNkVFP9q18f3Wj3oDiYJiTMIzvlHXciEpTtZ757OaodyTMFe
4t/u4DD2FlYRKVkiedPFuSfGPosHht50T2+s3Z7rMXmM/S29L0TUkNl3DSjpfalZUJ9xx75lbopF
/lLKaOs+dLrebNOFCw3i5k29hIvF8nqHwazilfV3tEGEEolJPfgcuc3OWNDtmzHgmDwrwI4V9VL1
venjjmdeSmGIf62Gg6Fda341SKw4IePXRPrNMyP0ultwbX07qdXTYYnQx0KQBInnocwL3BaXO8Hq
bOlYpItpPHpFqEW3VqA0E/r3+EVKi8YsxC6lrFJjWx+huLLxZ5E3Br5QWJFU5S/WRk39j2EpCgZm
oqg5sdol542ZefHZpKK6uqHKjzGTlcr82RUvFeBhZ7NGdPofDqguuSWmlpXWV8PM3H51Nqmsmngu
b0V2F4WQAOhPeXUj2c/WW/YTcRuPS1zAT20og7K0M0C9yAfcC5NjSGJwX7S2cE3Ge0I9VZpDWbvg
Kr01+PHDgppXVq2cwh01pmKC2iHMtvvQ77iI6bBfxFZqW1PULYlTGTGf0bgzVfJuxvFnUC+1H5lQ
oHsXGwLEF24TTGE1PjpX/FTOa79tvKUphQB0XPW3fsDP99dzt9ZY/WRVdA5/ABwm1S0r5l6nu3hz
b/ErgT/HJWEHBdyprGpI7kXzS/elXGpPi7fHP4PGpVwpZu+S9lve870qBBMqjnpvu7afiHeSFyf3
94P5Y948WMDQWD6aV6vKaLzKFTajnKCL8vjk5D/zOCzbVYjSVz/lxc4nZE7PkX78mOCehhriYCoi
ShaexhgjKbt4Uz17J8udY5oIDoXXax4MMYJ7hwQqtYB2V0adm1aye0/bv0chkuf1+hVIDCeFIjb5
IBPEjGaY/P53AASt7Uv2pVTL4B5XsRMq21CU+rsGY5DjvrdQVHGOOXQ5wI/SYWmlXKAOXktLlF+X
vK0rPQpjwD6/8vxJJcxGvYE7XVBI/JN2o4jSykVmb/VMizRXSxbQSW52DUQrkHsJHBq+3CYuw5Q9
ZBOoIu404cU1HYL6FYy7knwreZ+IARHZiPpUjpb249oLuMoUVfm6MrimTmTziFveK4w2g5idBzmv
2zRcfYdaG3y4YlSY0Uw4kGX/GsPYrSjA4nsEvyHOfm/EMtNGmX4ys2HcuZCKORl+Uqus1avqQAgP
4nNovC5CtgzbBBVwRHk0SD+KSbULbt8SbDVBsWnvtR6omVgp3MXArFR/Oeuybq6WVB65cRFsRr9F
jnkTz9z6L0cEfJ9CXQpnWpZ8+7xYEMIgsidduHKeh8SrrmIfqL9jfwB8PTYlo2cppDOW7qyc9tDD
Y/g0TBUMAg6BY89lCNlWjbQvqRDIq6btXvtxmPy6XBYl7rwC8keZgHxYtD3rOjw756tt9QTUilEc
U0Xg4I301nsSpHMb1l0V9dXyHb1ZcNrlTlsFq9p9y4RSsW54bBvrP4x5w6ZM2H2k55y+iJpx/OHW
CIpgyZXjSBrY+W4NcIJg6twyOzlMIYbg9EXitQ5Vm6aYafAfi/6A5jD4WDZ+X0FMZ5flW4pFOMHa
8SpPGbNYwMD2H6OcJQDPthTPu1/C9rPddH8WXh/qAUxpfbJdiempXMMw07ARb7lE95bCGH4n2kWU
9Hq8Zs1WQ9KbU+ItQNgG0S0t9QCWrinwjZj9zFsiHg1YHfwttULZMSqKV23/RiQJYNm39LNFCOoH
B7UzN9A0dLAzdAbj6FTdKoh4f7bNTfp1J/9bU3Z0enV5EfVAD6U6XcnMf4J+TTG1J69ubr39mK7l
gWV5Av0kylW/wqCgFUtgwMhpyWDXcqafXoSAwzhGWF1L28Atsm89TRt0SBklFVXe2yrenfZBBO/D
MqMiTWLGJipdKo0aQ9OdwqAS/IyUQNGinqKKfYwcBuh8+MaMSjV12pPbp4ioJv1rD3YfL0p06XYs
mZReKiX5qmynBd7lIaRJMQonmAc2jNe54YnroTECLJCeNqsnGctXTrubvSvek9rfDLhCGnVlGQ8c
xXQ02SAIPTm76fa6F9TNrp+umKcXoKeqVrnrLgu8Zk+oZfx6p7Pjh7RBAemh/+F9WgdQ7JUv5gQL
h57U7DyZoatGEneXQVCAWE0LQlyOIz5aO+YwZCHafbJHZZAlLwV1r7LzFf/uUUEc+i+bCniEkpEx
LiQPlDyyHmXnmj7O6nVTx3dW5f9pdRiPvgflRgBx2pjOx7eHBG4p752MQsEofppRrhCm4paW3qEH
3iR3NvSQt+Kh91ilgClYd6ptu2qipkhZeehqn3YQMhkNiy8e1zuxHF6iZgtBhz7mRVixzwEKGFVF
Edhgz/9Htj2oLFZOxLBLsGhURrdzeVB1NbUWNUp6w63Az1rLDHPUfwk3zZfNoVfa2kiugNLu8fI5
90aXRtAu7lZ4112+buYUXNnio2cjZzVtDJUs08GiMq1f9DSzIPH1kuWkuu1Da6vYQIa5eHaVyIMq
zzQ6qCktPUo6+cGTrrdVE81sNO+Oo3rPfCNQ7uQNkXppOvIBiRQXJurXEXrDMu/MsgjCuX+TY3lB
V1Hl3Gft/BfLJ+4MM+xh27jDp6ONbtQ7uxpoauyaoIvicj73qRbKWHOt3KNBlx/WZjiNQudTwzHm
US3fcCUPbdUNfd8AdxL6Qjx2YofSjoRUi2zwzhx8oejTtI89P90Ny9rwvE9GaqI5riNFoSab62K+
/k5eTFU366FQ4uqzn9X0RT4rj7v+eMrep2HEvSOQMtZAf1CYs2DU1mLLo62zZhra+IE4zt7OZ2CN
Q1zKI7tMdPpPdpnb4fp0O6ZWNkriigwEQdaqT/BgJaqSyNZUoJ8nRIYRzizJxoWLJicTcmi00tt+
5dchvATSFSbFRHTR0Ji5nvpLaB5kozH2kGy49K3b+YZrGqTFJ0qwMUVg/DWiFjmoZn/sBb2tQJwF
eGUCaqZRYUxFAEKAJblLtIwDLGCLhO95+P6rQ/xIXX8YQ9enGAX+bzV0R7iFbRKKPWRpddcXMmwu
DHoWYAa6l+9XJplKtnk7+GUB0DC5RDTkBJ3hWWJtQyS+FHhswfg2pRnfFhc9juNstV50o3Rh4vFp
1L49coOjyeoOdZyl+A6mbz7aU8CnE5d05a29vAsLa9Rh8tcd0Hoy3U4jtMwjY0Y1J6U/0yHbEjk6
HoPNCQ4/s3amnoV66qEXuJr0WvbHmVxXq6C4NeD1ahEgbLC1Ape5/6HhfEy6bd72ty10ZAFa6hZV
LMIUtIjls+pi8A/lykvKMRTxjx16I73pqAquMnPxy3ZF1EHh9yJ0ldCSsDitVadC1RxoiZAIvjfc
lyBkVxTIrHaSNU1RkaY3DsBweppeJ5xVG0GZ21aLAp3UaTkBGhMTZ0uk336TOEBz3rRcG02JwMen
fhytRC1iIGBWBhzv22u1ir0HZ0MrygGaWyeG0a8vJhhfqsBAEz9lVOy6Qkto+g75ZwvCVZquqjUf
nVEv4oQsfXziSgSZkgp6V4xzq/UpUOkNSpjE4v/wNciz2z5tPXuGscqAFUxk1KCTzwzlU3vbk775
5zbFIVAiXrI07lk625aswIVEfVmwcydWIIPOGwaO6+0To0yK22eugV2NHJgaB8nOyMosplXXpEnn
S0mHa1SnEr+2gCcHTO9lx9oeQn6Uq37pkoSaVYIO/IrScxAdmn2MYyhHOIzKc4GscMgs322hcbjN
ulgidnRgYw070437jIcc9O2ucxiqxmU4Bg76xALIG5jNQwZso1mnfu3265BX2otK8yTWqqA31ifN
uBf2oWUM8YGiJRXMWMSrEEBZZfpQw8sleCGNhTNAVyZBXd4E3n9956Iudo16nbFLhSSIwi1iwSO1
EasYRfCdgefPa3fWT26nfop+9QQQ+U3AqI6+32dK+tMlaveBP5I1LQOPjztlU6Nx/pqA/iq8hJfb
XwDApMH2zSwqK/G4xJGnYq+yYZtzJpk/JHwTQmFgX2JJfOH0cfn7Oyjxzx7ASF8lRxBLDSmBtgAo
4AmPaI4KWQ92tDe74ebcYr6y6nsiVjRAjVAyIQRNEiwbHarnuZD1z4qXx41rvnqqht7NIHPQRCVn
89HeFlkDqWbqCuii8vUETXwbVtI+vRi3pLmJWgeSdKmvGc8Wimxnhrho0P92p0sFGyvx8yK+lzkN
9cHNLzEHk/QKWjTWIGRnSxOjv5bkhmX8xZWl8pzOToSCO/RVihiZHiXUh2Q+2JDitQDci4+MXjDN
OvZp0yXKG5amnJiuCICtAgPs7r/1qareb6I6xYquRFMy/NQu6Q7rcgQsv7UqxoMr0+P4bkkRYDq2
AZdLqYkwa8Hr5uK4cAfmLRAyB54GSo/js0NAQd34ZNaOb8h10GdyEwJ3Gz4/7pQMjmlsOs/IZ+9z
3qcULBHyI4IJEtP5RFgW1eBk274GtUruQtUcK1LxfxfXfcSzYaKqqYIXDFktbL5We2pb6/QWWLMf
z9YSZi69oyhvg3SLM/yLGvg6KQLYnKmtMBxZMzNO+A3eI5UMp4C/tk11XL989g6+9BqKuncAxQtx
c2i30queyb+43iO7YbQ5qSCmRzs2nUy/sKa+zcA+m8KVpwspOzndHZhfgccEWu2wb7Sj9t8+g0wm
MlZ2nywHv4nxpxBkIJOcJBrIrsHQ7owlrrhCNAP84qVfvFOJnjlQdfLstXLkgwreV6hcFU8cAO6n
NtUGhbV25kfxhPi9Yjn3LDXe+lFE24t6fgg14eBtOz7KukVlP1IBdkbLLjVokb8BG0ya+74Hvgbl
bgQw13Xyk6fd5BaygYidtf1IGScWn/kvcWjqgbJIcpdogpusPTdXCcavM+3F28Aeld14Gj6d0IAG
C6M4NCq6eZhgc5bZ2tOcTeeE0ucKzeJImrhB2g7J++SLdBJuuhKnxpGN7Sz2wPnCMur9rGYHAmYn
5tBd7siJXDWYnuq7K7oAjMEO0L9TKeD9+pXP/p3vfpypft3hvsiw1iun03L+IKzdCRzTMR7FTDJj
s2plWjJNrFkX00i9bTkUKGIyzAxkSFlEr70P5FkqlNAx6mspRsc394CGCH6nIHIe9I3pAl7+ua/j
OpEsWS3R5allwCsk2+758eOhw1/uA3+B8Y7kVtfpIzLlSTI0CvPj8ATIq26G0SS+5LZbS3mVKGcY
81QzJKZD0CuCWGa3rNKTA4rHEaylmFkK9B6jJlrQNjtZiDNtoHmZKZV5hIodqL0hI2jnhwzZgWC2
FDywgP5gkUrAW9aenkB9aVO+gDAXO99yvJk68A4WDICXcYhOfO7OKLJuQI74dE3R8TgxZsEP2QYB
wTQsPLUuwIx9Ic46Y9XoDA/PirH842SOozwg3oaw5DT/AtzHqkNOnLsyLwQ8iHBNGIU0e5Y0MFor
9zzSBmxyd4eUC3RDHU827HVPYpL80X0QJGsrNtf9NXilQnMR4HAR1dnpAxP0HEOQngHuQi1Tjxgs
vd9Yp2MmKZ8ZX4EyBjgd1qJ5gx1VG0R+Ym0IHhrzItzyAR1M2kKqyomo6qzlN1H8rna6tushXkp/
4ZV8Mwkf2LKHgCzeziMvKvrwdej+CUl7b+UibQ2wJ970qAI70yKMM5H0xuSVhUGsY7vzq2X6rXM8
BkacK13D1wuFnbOK9BVgz8qmYt4lK0lmRkFtE9C+20zPoldZt5DOMiyNdZWeI0F1ceSTwnvzQudq
wole0T8e8c/z5NRaPHdQiw4LByPjATrZVGaizsBrJTC+fl5L8CSf4LqYyBgdq4WQ1dt3O+HTKCwo
skzeKS8mQBlmj6sOcIeiWYHjTwuZ4gmEgKEHyojUnno7euXCi75Zm9mCdahiuP5EHZJxPvZzLHen
4m9hc/PyAxAvOZwsQ2OJkRLNnuHyxcwNCHcs9lD63nd1JC0zGUImlfl+WGbVYP7KKG3c2WBBvJtD
hd9vO8CbWAf0j+5razdz05Ts4AFlN86rBGDnvzwLAI26zSzNocW6tNmhpF/RTGtc7rzIDISESWrq
mJ/uATeg0lQzKcC5FzFvBIWYWx/Dlrwe/SAKIMbI0MH0l8Sv+QTZuofN1VncGWJxNaNIC10GN7ui
JB13DG2JtB5ictvRsEMmblkjYJ767PHj4ryHBFZ/06oxefp/PTR61p+Ck76lHsk659Ie2IlN0XaT
AWTiVZgieU3jF7ZfjzWwQNldxf1DxRJmi8/rcEb82+gwqs5Ot8UFjTsnniZSh967XvkFtA2lZBnN
2cen2ftCT7I31zr9d0qJdJr7F72uN/Ko+lh3hb7+7v3HcfzpjYit2aonPmxXYqjXF0Es7umg7bBs
A8D4kyaqcP9ysJU+eDz92Un29sMDk+vpwslUP134KgHDo1yx0GISaC00G7wQjxSpDMBOjJ+ZXmin
qJmVRyAACeCMDBwosW4Fo3+LRGFP3usmbShG3VEXN3ayzjYI/ALjP4UwVm0UUAmxny9V+OqD9kzn
Mg7e5hVBTBWsfgP2wUJeJk/5bYg2FRD2w/Opl17L7yavzYbqv+7M90ecdhgt8IDZGJEXsKXBt+nu
C9UBL3e6SZoxtCHvQ2yI98LVH51Ef/F6KncNz8Y9UAVxy8CDwolRm53KENoidyr/Yh6iIo7gN7TF
v4ZFcQ16xLQLAdODtXvE4mbu/ZWmPrsy45FF93YZUxkviuNrMLSuFWWuJMAZNJXF3YjlUeZttqxh
zm/tiJwqRmUxs8YVstzcI9khuWowGhgbg7lYjLrDTHvB5LlOA8obmwm2/vOw1eQm0RDxs8lvkuuh
tw2jI09Rzy2o4uEg0txVeLlIXb0lgtH1JVarg8SoNnwkRjVeTGvXeOR/wl5kRNpvqHKuhV07RRdJ
ydnLgqBxCcEiosbUAj6V5mkbtiS2Jm+m3SFnx0EOKVDgsEdAm4rfn3QOSB9rlKnDB7qBE3kFE3xM
YT/D4tOCG2XcFKu2SlYeBB53KA2CbjlQkj01nc3+6BhjQGNm8lyZEJQx9BB/Dh1YArkCnDYsyHze
Q20GWa7a8QygRiokcMf9pCDqmRaxsY/NcSQWJQ1t76ZfGrt00QnMX1/KoqoDcOOc/FyYG0TcICKp
QPTSSDLL848wvHmwCJXL3siMECscmfhZugaohHipLhqN4E0B+qgA+adU7z8+OIFAEE4i1Nh5UUpx
NWyroKeHRdNztsLjxL42jkCNgygFxH6OgoZ2cYiJ/O+SVC+X1N2hopsP2NkxPBPIu6ihUfXfi0l2
an9AVXyqSa7teH2CHjmFpOrsDbBHSG4gzzCY9Je9/l6KISy+jpXwuuCCNuRpatDtF6NCj6JwYQOe
ADLnxT1jKDnCfc+F4fKSiZHwVsgZb+i1VoZFDNuCzU0R9Hw2rlsh3SVYwJY2kQVEMElOMECW+rZC
EvTXZre8qJVlhQk603j/h2IquaIpaMF7CuhfOACnQYoj2vK6dg8A6ti2MrFiRzj+4Nmp7pVttBPE
fpwPW4F9ik1Qd1to58vIXZua94HZRiFmqIiG3BJuqOrlWJg1BxBGOLAQcocPrqUTDB2FCRlhGKs5
IDATEfmx2KB4+NzacHvJKyY1jB9Jz7FOUTsIulvp0LKieaNCrkzLp3LxkX6p4kV9IgyYqJNemePn
6yjB7b4qpys2KN1zZIkApz7IyDcW2ccvZ4bmm23/KkhSLmSDXvtJhRIAx0J9nLsPD0t9oED4HxHY
bPaKeQYI3nRzpBPtX3tifupMm+9o+DXhre5GArICw5cRh1V6gccMoHlMVDqK7LXOcQndmclrFtje
uGudbY2nBW4/I+BoVtvI2xWO7lkXJ98FmoNhTloqZ0Yd2imgUsbBePJFEZL57hScoHOQi62mdVl6
g5n2GC6GO6zSgm+Q9L1/8Bvo90I/1aTl4im4rn9mSLs7uQB5xJTjFwqG82UhUiTzp1LN3Nn0EbWW
Lwkpjg8thD5A2dzas5dSGzSMwNG5SpAYUMYZAiZoCsQPf7tTYSGneNp7fBFOvoWf3L1WdIwGkzKQ
Q60CssTu1v9MGHW9bXjhUSX0IV3PNLlTe2yavN5OdyHu+M99vKBXTCLYF3fdrFLwbRrHRlhXxsn0
PGWe33h0PnMJwL60Ifo4hNOTvp8DIoFtvhobvxP+NHQEzUn38Vtg1DKW5pOUU4sDeAuWfq5bg13f
MubhxUjT+DM5TF61TkISbFx+PqrRuC3Ofoh8OBSAAFe6sRvhYICaKxSfwSu6Sx9gRSqqtWjyb4VT
g3iM+/spGBe+GNXe/h+0Ir3HGQZyMUHQ1BWHuMb85/FwPxe7pNYQd4IJzZKrBRRNMwOWDDKGqW1E
vTmGYrbajyYZ6zcjFcRxZN5Kxrx+neLKcof/mVaoEHhwrwDpNmi3NxC8RpE8kKKwA0UPAJsxz+nH
5+YuYC1ledMyaeRr2h8Plwhuz0UhJMTV0G9dGTEtmxQynuXQupCEG96hIyiOzUFJofOunqhpcs2x
hgQnWF4Qup+OF4HB8nXdys1EDC9+3OPFsPiAAsqMI+GYexaSrdSYRFp3uwRlQdkFi8gnCBL9deEM
19175YZ8FeHdeNRG6IFyE02EmafHte48QcHtpq2eohzLIkNDQyk/JcCOUppyZtw4s51lTXLPTPkg
38dIkOiAGp47HsobPl22/Aqq7kHIlmnG4lKveE+a2ZWTblchXmGYjlajd9Z33mPvTHRG/rKP1C9u
eKLdGUvDjjMphq9EijZoR3acW/n2WKFyJqS57LoPpBuHeJG952vsHdZP8HyiqBmTKKfOAu+RZFej
21vmbC5OOVRslD9loX9A7/RJX8MjEHnHs9QxzaUUYSrbL1ocyrM4M5TTO7o7qrMMJyt8qgiOFDh3
iV9lzZINZOlD5Vkc99faCDE0n5/Vk7wzWN85QMaugy+WlaGFzDsbgfPHY7VcHD8cV1l6U11qXqjU
HwgLAHBY8Me+TIhuj9prK3cxmKQnpWzpf0/2aWa5KCQNZbqQVekOvEn6oowdVE4PNSCLth0Hqhz8
h2wiYooxlQunZz5AIY//+J0JWP4gSshBNeg7u4uXzT+7/0c21/8KPKlJAUukLx5q7iPfMwoKI67a
4/cTzj4IQowJrGpbLgjE5/E8NxXtwJe/DVmwSlFptHvXfxFWD3gXAQlsI0j1H5EoiKc+ioRoNXoa
baWRdooISvJKL6YtW+wIBDwqUV56CHxF7lZeDpR+hjS4SGn9im+sJ3Ompm6X8gRehGRSbWMlS8qe
tRgS/OPP7qEDuLcu2VcLVynIf8BbzmZq6urdH4z4egKDhkhmAflQcN4F29qiwKiQXxNN0jvid1iB
ZhkMQegdF7Us6zAaTp2bGvww6aoY6wcrUrv6nMT2Lk9WlAzLEbjiND8c21WFv0Cl9/K4W0P1LJny
HfAoMcQPyvu+mFOwEPZdQFUYdGaF91ZcRdBxnL/BCa1TsD9DrHQ88aw3SuQqFBBxQ8MQ50SLMu+V
Yiw7CjAbbClwwSeZKzPDH0PQu348IJ32CjOW/AXbUrc2es+It6xAd4FL+nLkPShgwcjFAqxdXN0b
bI1Lwome0djJ0hR8ePm94ZH051ZSfXzdQrkA6sdyN6I4I7R2PtO8Dau/3RslrRbW+d8l7zVVCeWT
5bhGjYOV5ypl86hE0LpKjm+ILa0MaRWX6R2TZuzEZ8aYrxBzgNDwZPBmP8I2f1tQIZqhP20qrJVU
++8qGCdDbg0txEJxJ7hMpqXoIy/RH8t0eQZfdnCcPJzgkKU5e8VI44jcrp33M1Ucbl8dejCh9fz+
jhDXwsnj07rtJQQx667yn3kWjo9DZe01fJTebK0G0zZ++p7NhELHl1YGt/YSovYiPM/Y9jnH8oln
e6mk2UFIODKin1aM8U2vHecYOcuzURqo0jK5G5WceIxy4XIAzrDxtrZs/i5ewOlcvGRdPWDPg3IP
XbauEvXE4+jDrxm3PFaJy/ioWDkE1aFTuFEDLfBVuOcNJCXZZuxWdVn0dgxRNHhavNTdqQhvYoe/
L9cpXBp+EOoZtYP2n0tA/1EBNOCui8Pp/L1JHqe3blrs66nCJpIUh/qoh4HM9kld6xjsiEBA9le6
vSyTiC3A4M7a2KXwlxbHG/f3ONuSKATQeNtuwUImefuKn+nim13n0C8qloBdB2S6TQTc4bXvXgAT
1Hidsqpze71BTXuqeC+0Oja77QbkTdP+024pjZo3jgMUEAw+haom53O4ndfIOdwFySVjcq9XK6Yo
+lJfmX+ev8Gt1qI3hA83C0dRYV6u3q3YZVs5tgOwZV33hXPC27ypvDNf0WhX0awqNhcyt5XSamFM
n+/qQXoOOBa1ML4nmy4u6LaCj4+ogkNYesCZrn3EVBIRS/Gzp/60Yf4zbut2OuZNuXFkWD5dS73L
uuihYj9LWEdjjEAXUSnD5AvLAl6cROSGw8sE3P9aOzJYagBBEe8e03fGF+oVouaaXjVPUDm5DOXC
/XAsOKc/LpAmlYG/4NbER9N1fQfGGSmQixDpG2JAN0tDZDKGpENjmwPltHXhu6nLlBupiJD74usB
vPl3sNvym8wiylrHZLJIw9wz/vHYSFCENi1K5OP8IWGTZi3Kj5TGtAVfdcwuYO6yRBCNvb8AOK0n
QGCPzJFM26ptEuRNrlTIQvepHRYu02duCZPE6NMmrRWh9IkIU+4H3W8izNOhofF904TGTeJ8l1zX
M9esBkrmATHH2SVG9XBPkel7iUE3z6iJ/f8huc3oZFoUSKu7bYOYE3jRrL8UAtlULilT20cGJQf3
/Wbvi54MTmTIRoc5aARM1mpxOdcbDnGeWw+ThstKzRB5Idl9TABRbWqI15ZvCWSLQ7LxD5nay2Kv
+wrO+Ryl/AgJPivljrdPQueQ9fEPuqsCmFrO2vX8s35NGyzgncbg147fvG6sPX7LH53MulfP5E3g
9c23WqOGCKtDI1eiK723U8mTbIIAmOaqsObm+uwEGguyy+6nYfsVgyY3oc6Eovheea94zZeEtMaj
qAluLg73Xlm7SR/uwN6BwM53sUkpgdDDrp/wkd9FzVmiOUjSFBaNvP2kMVE4wuFgQ45jvCu2v0KJ
f/VyuFJZI1c6rZs45x2/BVKsC3XlKxkv13POP8RJ6gbV/yTC/BMEaimXBCL4gOIsewC4NM6HLeUs
eKkbYNB/GJC9wzEB51KtTcnxpThJoxKVzioXGnFKx44ZQi5X4S/xweVypNZaZZJc7CFBVYOVigmB
wjQC4oWrUUUUvwAM9P9SOmr6JZ1PGMfH5HEC/YDMa2cZacN+lt6TDMlMHFVsWKh42hKGxSIioK88
zpccCRkDFytOAPnRYla+xOBOvBfOmf8b3WWRUMDt4/+T6LvVvnS0ZR+zETiyoJK77eHNCtqRFibO
/wmh2TVse/WPC2OCD/YTtjmGsmxKn/7hH2kqska8FAY5GhC/kFk9HMAMKl3ELvt0HKFPEhrjXoAA
V1qKHy8R4cVJfkR5P1LUSfGjISnBcubKmRI2sS4GAT2OKO7fly8/7AtcMtS8H7GTAkYfMVXYfHzA
iw1RyCFPEmKHxu1lRkLhapFhhtGSbJtlk7qj8ubG7NYuPZwGfB6WR5kkVA/uZgacpiE7QTyuqVcU
UijPOXY4O+7aQb01u7j4hgLul8Cp7px1VrodFJ/iWx9w55LzpZRzWFAjLzEtst/y7Rbwiq6YMA4Z
VJT9roYJkhtSEtaaM8u6WIoQnJE8bMikVyiXZPAxtUwRCgUBxz0yQihu73kxFKSWmi+g10oThSgI
DP+33oHi8Ised2C4v41bslnW+8C8UCQ1VqnFRry2lL1+T0/vBhapkxSUdkeBE3hX1fJKzb96y9Ag
JqR0AHdHdnSV2RD6wb6ZI2iCKtScqavQkap865Hg8EI+SyD35sd1eoCt0x4PhFpip2ufl7ycnd+E
PGJ2LRb6IGNWhAh3sJF3kJP9mhEcdS2PvrlktsY+g8Tgr4GIl0FULnNkUoZNcYJNgwQ1p7xTm5gP
8xLrQBxJ93OkHH1woDI2oTq160EhP3ez90W04p3tPnGa85Hne0t9HQiQsm7Yh4Em+A8fSxQ9zv/+
zusRuCebP5L1cnbjsHFQ/XKiD1EOFNpDsSkD0rpXVytT5HWWPKDcXzevOglL9pT2i+Ixt5TDzA85
GUu2ns28TwgrID/lm/tw/O5OH4a2QWVcpC6lHXoqP8ysseDHmydvE20UJYA0jetgBl2WqD04opwz
19Gj7JpQQW1hjLhAMjkMdk7C5xoCbVjnoh22ohA16mdBkse82Cu/1wMFdMT2T9BWiJaYpEW/V9W3
PGXhPcllANuP8O5dj5K23cijXZKyDs/tiM+HRwK+12wsTcZUGETlpedFKApLf+yRoKq5ZOOyW55O
BpG8o6g2FitNhWdVYZBXgFgMtyCINeRHpwnQon7WxPxFOvYPBWbffjmlipmb5k+8LKDJaUmfPQe+
xAfbwP6+743gLGhNc3HTvBxzyWbhEDVnLw4uILVn38QQ/+E8fuO7kAhfGP4CXhHvlkFsvwpvIeH/
b7qN/WG0nSnm7TeuVdTDkTbMHo7ZXhhQAmxnHU8rRuGW0bdaf0FPhZ06pIoB2yFfq08yiUSiKCGe
nQ9GteuRIL5n5eg/w3ENe08Gl33hGe6xJIEfT0G85izdBft2J3gnaZwnlo9wbqlT9aVxnO7sGbbS
NVKTwwupOnSrVA3qyAA6iTFWveCEN2xb1bLctdjdtb3fryxJL/E/bN3LyQvj0Jj7R/iK585w9FSw
74DI5DCkb7nf3bMq2WIDbO3bkP1H5DQW2is6s8QIU8FS1ZdjjM9D5trvgSFlR8TIEC4tW4LjN28d
MqIDYT69ZT1Tvbyx3T+SvTeoYu830txwnRKBbiBW8iJEEycQhrjOYvP1AwWg87+AEBT2h6Qrp1gi
6YyXFcwKhULWqKmaG3yKVhCKfBwqraUXMtOjU2gqtUHtZVIVJC2av/VFnlH9pjWyKDVonCkTgRCz
HCi7k4SwzLyOUYxAOWNQWuZVZ89eKM4UaGvDRmoDWCiXZx7HiWR5A6DESBajx5PGclEq4jwPrhRc
2O83pChvTj6GI0HqDM00kYNVMNEtGqlQ56+acsDE6qsoYqDUbRLG/aZMFZ45U0e1NnDXmxqRD6Fq
7Y9NWqjWtk+GCKtI03pHE9yX3yjhj1dY7E2nFZdkeUAr01LBKEuv6zpR7LUEs6Zal1payxg2xBLi
v4tNxWbdQFKCZGntLCMMpvFIb+V+uV4ZCZvP76c70oOIjDeB0xhhDjS24/gyQstZ42kwhNXXc9ui
j9vw2L7+FlKAYL5ZSqhRnq0Dhvgz+/LNxvUwL/PBkfjTHGXM52nmOgje0YaFTWcKbO6UG7v39h10
e0fST367rcC5Z+artAoYqHTbwsXPHmgjLdAi8v4jtVHeTPSd43lveSIVaiuMB4SovkJTRGFdAsuc
z46k98vKfAAEUMWaVuoPUdqeRXoZ4K4q3Mj91a4RkoaDlrADS4iC6V2m2VZp2t5JlAfNQ1EziVY6
3CFOSOrqN7JkdnxtZzHiQ5tqJXUQO3optYGcStdjncvjmrygYuh/ppDrjvOCAtfgnFZecrwqazY0
Eq41ux4p/BZxLSWNtCC6VvHfnMYYvnJga18YmeRPrXi2L5XgPPlxxori8XWwnIAtOIcuFQiZdtAe
YQOT2auTkwO4gosJVGOQMnnhKkn3od6AaWSKtxV9uDwCoqBqZTWuKW4QpDn4q2uaE9CsuktLT+cB
gx4fK119gcmselO8TefSfacwdoefCjTlLvIUZD5NcqNeHIINxr8vm/7Jy+xxA3kQ/piJWzDkCc8i
mzpxeqmaTOc8+eHngucVFV4h99UZ2yt8mnfxMyP2Xm7sVHDWSd9107ZbodXEZaEqaA4Aw8Ikqcqc
kXVTz2OEwtBL9sCAQ/wO/f3nYk819Fa6mSN3CbUXSXK8SuRO/em5iY7PaY14aNL0SJfFKNUjWR4i
Z6WG2gNOv9nvgvYjbKLu46mq6WEO8W5CyIbeAjjNLg0VtuWGMFkiNwuwjhOiJv0ZQ1YlcSYPiWPh
iTRMeq+DvkGSb0mOP7d6Ot+bOIOw44tS9ydb1/8tTQGtBhM74cpCTwQtzTvAScsFnmlbiuXvVoKA
O6Ld+wCpKpoELto+WZe0qtY1nfLX7uRY1yWNBwZC4lUkIxHpfNzwUk94iBdQfzXU+qVCWIKc9oCw
/1XeO2Ef/QIZm3PCrwObawX4t0EdK/wmllUkRafgdpvHruGk6HiU2NRB59zDoSlB9BeCwVjRYQnx
bk+VoxG/SejnY/vzle0ncYx+mUAVPvQlXhqpJKHABIfKlH1AWnVg5TK/VjcCfzgSE1rX4FtVRub8
RR3WJtQZbvD9WsAnsgV0Q4iWrvWz6hUEhqzYgj8luCm6b5bDbB7O+I/aPfiELvsaCQllAe8SpboL
g6IymGAgmkAhDWCflG/h5z1i2D/GVWLy7P1Hatt0/jRhAcGkc+/t7V53ADAGuIocn3aeAKvVg/s/
6z6mkb1woLjqe+uw/WcdHKoZ8hlhoUlYZyEvjMD44AeIbdVPiWuVgCdw2ET6zD5ZwJznFzMoNUfm
V9X++iln5A10u6tsEQjTJfhKObTJ1Ns5aqSqG67IQNvopekwRAIbMpFXLJvz1gbF2+DCWOmu2zMv
g37Y6abXvtR42LmJgAMv1FoZj/3+pA2/Hww2B64c2P+3Kw2wUJzfMO6+/rfsFpHrJkzdeJt1KVac
dhwcJvHdPJeN1vfb8IZgczfClwLG+WgqugDHVLb7MXfbRM8lqzffmlR61kZxJQpgt3nmEkah/KzW
ZVU2PaUlgtWYPVV1Px8AyriInH714tir7cR+XhOxhbMOcfz1kVr8qs0KgmdZrtQdtUTwof8ngAgi
Xy1fDCc9UbGa3jJ2JGiyhvUg/lDzvmcuuAdzRCf2buO/kK/rbsZYl2okSDEtfe3+vlCSqET2rTQ8
+L60zqBvBbDHiNY5ktmIQbD8VIHZUWOxh1DSqPsdWHAI/Q/OLWf8ZGNJqoa7nBrWJjUEELO8WxaV
RgeQGB6483R97AcpqgmKudF1ByTrqxf7OYrMK9+8zxmjEqPG7+IZs7jcpkZ9346zIW+KEmomNm8D
jVbyuv8ovzXyAA2+aWYtRQePXyf1qmrrZVcVkwosodqFne13Nkl665LcwOa5myDXw8mTPw+8rxNd
lGuaJU8nzeThmYpQI1IYJjWBVFzf50X/HHs5Mkv5OVAn7z+ogglQ+7ou/p7aprRB5knoZK9Bz9q2
CKXtRG+QTz3zLstLGFJfabZRKjK/w+njMKe0xXjH/gDf2dJKI7XxxPPyYRQDzRSLN2pZRFsgEgl8
wT4txhejhFbfomOzuHs2E2W7bp+xCEiRLmuDVWVo0rscaYkJ1d8VdkuwTa/FDnl8Czz7mvks6zpa
xV0+WWiaN67LRvLsG6HIAwWCzpmZqF9Wamt6cZVG1SAjxPQqRQiPZKVgWw5Gra2qS374ekfqMNDo
x0uQzj6bWO4VSFcdNDkG8uuVH5xOhFOTJDCgZuynt52gwQxaKalHhZ4ZgoKOq158WkxZJNMzyKF9
FiTPSBaXl9hcAEAkgvj6xPS/BVBn6VOUUE4uqyg59ArsXEs5PfHi9LN41pKSbErywJ7JhLnLyLLe
TyNUcwYY0juMz2mSRpSLPnZEPjXDSKHjgYMyPXjPf77cU2XYFzm5N0IBygFqtkVXphegK/puLAlo
4QQ15bdBJ4UHerVv6guzixs4C3t2P8encBHQpMvY8r3ui8MNRpsqKjt9JpyglWA6oXQ08KyVL+m9
AcavLOu/J3bIadNbTnh1gqbJMNQRkMcpz1sonyzN8nTx162FbqBzsCEh+mhL1mLrAVjq3fKkzR6O
/0l3skmflfJThsCP4QirwiyA7Mt8wPrlQTjSf1IODQqEcfWIyi3XdYw3AMTFv6PGcy+9ybmX6Yx6
A32U0W7PfM68lTFQiLmKYwoErdE8UJzqkfeqPuw8yPv5Txyw/qxpdiikI/cZ6cAGt/TPe5ALRa/U
KZ+TUyy1+W787YapjGWS14gkocjzc5ESTjMmQ73KR/A6XNWniRfIe79MamklKhhEVeKv3AMcGVyu
2Hsh4Sbpj/HBcbbguU3nVXovhYWbdkrXUmpA9xDxVHyUyW79RWCsDPoMEUkChTLENOYsYPNbz38h
TCG3dh11y9bs1L136D6i+CD6c3B9Crg3Kk5hQJ6mHGHmkA68zU9PMhVB4cdK+8nG/8U5eGewbfll
7sivFQXZxgERHMJCgd1np3HMPmdtV24dZhS8QxtsaWe5r2pYkzfccupaWtWvMpMxah2c1zMJgHgV
pXuiA1uZ4TysM6Yeeo684XF8KwbU6W1vdhoSPUyvMwC7c11T3Z6PFUtNyus95EGMcyeKM5FiGIVV
q1cc9UoaI5xjIpkVmt7pX6vuzjOHUU9Jtx7G+oAKqM+414uc2CacWjituG34vl1r2m+LZbCnKW/0
+fJvStbmMpEqMX4ONjKQJ0RcM+HgbMLJKRuZMDODQ6q270Z9qXgm3X5v1nWfMI2hZgUOJXmGYBuv
9qW3swbGJudnKy/JHusnBhOxAMCqdRK7oysglEWL/le5P7z7DhGODuiTJJ0ZT0aEGXWabZP4bisf
goyu7Ayqm96ycqhN5rC9FgGG6nmQqaYIlU89RsGsk/f2pSuybfC6csQwQhp+NtgRPED/J+vXWvUH
utOxYgM+t00g2u5yeKu9RLbIEBg9xxQvjbalirgjKSyoHz1sGOZhUa+fyUsG8Wiu6sblb92M5+Qx
BAB1SROUt9h1khBUdb39wQVGmEVSw45gnMmHtMp11jfsne9aw+KCx/G8QuQFzNx6NeePek8K/xmd
HCaDt5LdmDffGPwVF26qmdvTrq09280p+wAU3kqQcZkxSQOqUqpovTP+Kbm0lwiu0XdliYV4WlWx
H7EVMQ3Mk3au6D97CfTtZnk2Aqp/MuIqpmlXnquTucs1ghRIkwZ2bRzeDkMaDSeUC/h6ExkbZhpA
BOOCa5wV14Xpn0rwy6NxqefxNnNY4saOHJm2xZfLMoVPnzQEiZPz6dVZPRgq25JCzpZgQb5TnE3N
4hHzL88M+tmlPQOfeTZugWYNFfLuOYUqbSYSUxcloE1/D1v7JhpH/1lLu0mO3X7p4TXrO8w0tzox
oAP5W39My/MlrsHJB/JJKGNli5Ef3ndoIVJR2PTH1VX9zXSpUZEKIP0dbLovXsiPJNNRTTQGBC+o
CEPykr60v8Jjh0K5HGPjVZEnO4OeVy/lHZKQuZugkmiEllg5BOOfiSr0Dj3/wYeWIIiqTyM+qLP4
POcgOvOv2jRgyrauCExf0YZcT9x7ZUWwdxO26GrWHsRzYUVbuU8BLX0ee4MpFcrmteRaCKOANnnN
6eqSbYE745I6aYXeTobDPBSPVdAVGqM4W/lbAM1rMZlFTcn4MVqaR8opAFcfrla+EDHLNWZdVjsD
l9L0zI5k0H07PPn8iBKHpPSUuwdl8jieD36UsKZsyKQJvh71FqqMI6Dt2JsdPqGNflm4wMu+hMEm
cQEiv2T6/le05AzwlTkHXOCJmJAntGnnOuO296QotfHSqnQIUSHjFfVjc4n98+SRFSJOVX6AvFvn
K4j0FKTT1AXcCZCz37OdJIbuIAjPr8iI07rRPKByb/74ZFnmez0ZMLeSdUjZqhor1FQoqeqd4BOT
G6S2KrGJulj4KxuKx2f54D2n+Sj8+Eew70KcGumMJpXEQSX8hQplwARKICDQieANwjAy+7R0N4Bw
Z+MqYOH3kZmX41sfv79x0GkoDONx3XpIkc57dtxFYfyvnMYMQkPEPdYH3EDb/LSoGUXOwdlExM9i
XolVfUQBbkwrryX7Ef45Pl2gXo6LsweVAjT+bFWXROslOrlTiBLLismf77spr4w/p1sT43QrEHXg
BxJT9d/faiqzyerNUCTNkgMzOXOBPtHHZ8eW6+w/R+EvydbaMf61paHrgvEonLb1CbJjmvkwd317
Ka7GvdC9o13eGgJ7D/cTjGrHu8Gjys1l9ybaz6gm7uyV1lcD2l0CFUCBvCUbjGJeETcO+Hs+pB+l
dIKwUqgzsHxIc2Mp06jWT6fq0WVulbzPTuLTl/cmu5hF9bOkJX/DurHjnzSczPCp6o6vX7n1hdQh
91w/F4EmKk9UDIdx5pW7Tn9Z5fVTP9elHirIzLHLeHjrcr3XkyGpGgmUdUk3LPVVTYS8cMsKIpXz
nEwZ6znH3uyEwMRhFZj1o+o/hzYgfIIlu/YSdzIkxqpuR41ZCw8KOXlgj0NXSaGfduiSuHBG8pGR
1RI53RaT4vICRk/gZdIjh2QZxJglhkx279w9LqQOOzVfI/q1KMEbjgrH4Ww75UtPuULbDO7tTMPF
VC51EU+LUgY2uOj+To3l8t049084iYVs73Nf7YKUWuWicryNRwkL/xVzRbH09fHs3iS/kR2UzN1V
i9kz/2cUrDHCuTf+tAvWPKNdZVEUzHDvMN3TT+zZPV8KmJzldUGYAa3nH4XjSL8coPM4ZBgdmre3
RynE6fjVgWYbHF14WeJVn4MD0BDO//mdqE/ZDp59FfcPq2Q6sS0KxOemvXd095RinZOKpDewiR76
VYnUXQAFBi7Er8eyi15Mebo9tFnpD47ByrozV5kvzEfoWpDU3xELg44KW+l5NncSwmkB+T855I45
WtXtRucuPEYPmzhL0lMf1FIhKcw/ki2hYNWFLRgwow5ldG68MdvgVvBbRm8TfeZWPT6nzuz75dMV
053R05wKCQoE/5CodcRQAo+jeLelrZpEUbfQnxswLxu1tLqg2tKRju+WCzrxI83rtpEi8iudmbGA
n7ePygY73mCsOz9k0rd/1lOpIAYfTGI6CJyidE5IkiapLpiQ6XspKNNuI9kQdFWfwp/nwQK1Ubt6
ZRlxxKqGpOZRCezBushdyvM426dCWuWzKLx7msDarpdp7qL08thA76RMeG2IMz2OWHp4wJq84Dt2
HdH33ntmxBCdY6Tfj1uTfl0NuATm5Nnc9JBiNm2JeM/KX6F2uheOtcs/51wGd/5STys/8q92+TRe
4wj1TvxM1ewrOjpEHO8kKwWpPT72LJ4uDBH2RHBEqFGe7EDbB3HG+sRiQNYrlS1oqQCzpF8F+b2p
8UhdgdmFw85qQ7I1SjJJA+Ym1BjUEdR0mKN2C83PlRMVkgObMArI7sWp4qDoDObcThsRvnfOwj3G
CgH7oflDZDq2nJSpCAfQ3XL5Mx5eYgrlpnU+RRlpqgOwOfrCYQqR8EyJSaWyq/66zQFvWeGEjyHd
NL8dIRE525oTxaglhwpqLYSpW5YqH8HfPdOxQDNu0sgoty4VYwFNgSBgYFrqrefX7xnbgKtx36p4
5FjoDuRQkQ+JWmSbhdDl4eFoh7/41YVs5JqvI/jff8aH2BVLCAfYaCcSVOGWbf4kMZIRIOkitq9H
1Kqheg7HAb6E7aF+PqOGxV2SGx9424/fuL0yW7fyOcebc6pvhh5im+ACRSaLmSvuIbP98SJJYxL4
uDjmMWrk/aVI2Xj93lHraR4L6Ib4acAX8xMWNGlXV26WazC96PAEiX71/GcQXpcxKfd/xFqsqM4h
JW03LGfVu3Z5XjduOVTuNg5lB1gruMJ1JwiKzgM0eOTBGWZi2cmWv53C8jHqNxip3Bv2PK6FiaA8
0ywvD6bKG+YK6W5itq574sLVsvFze7MEHMgnczFEN4cHwMsXZqMHnqctBWdazZ+uVJjhbUxBmGAR
tfTG7oD2LZJEIb8qMi/MAi+QRnrUkQiOBbdblTx2Gw6cEn0QP2QdPdZn3iwklY68jmfieuyNE46z
cM3Rr7OIouvO0MPWOcjsXf2FoEvgeVRrTX8uYK20Sm/9w9JlhWHA1nFZwnFi2x1zeHGBwaMjq6Fk
UozcelNq8BbTu6ROYXgClbtxY9m9ZG8hs57mIb0GcEa5HxQQsHmtrvivELWuoBLwHW014rfXyNg6
mayDuBfA/aluw79ILu/ys9xmTfIG4XpsB5OET0WPWF9jrKJh51CYX0ovyfzGY9Zru2pk2tNX6Srk
6+Ym4Dmv8iH/mzit/9IU8KYqvy625tCrhnfBC6TLaxMCXZS8D/2UHyzhm8EEwAjv9+URV81WZ5yS
WSoL+ZsMjLiSAy2vj/mpUiuUTG5AE+gJSKg4dE/UC+92h60NaiGwNt5z1CuycMpOiuXtY6f2RGgr
kvrbz4pdZhGYt0s47JmvlWTy2ZngMeTjajJAgP3q8lAt8vn1czWu6Te0gU+C/89tDg2ulPlLcMO6
S/n5wRkrndEQXxS3q1hWvpyl6OjHZiY/sFZa4OAH2Pk/g9Xp2NjWkxF177qeETMRSvPUCOmzrEmf
6x822d6jrId9uHQfRsaz3BBykpW9hVxhzq4lREet0POF6uD7tQAosbJeFIo7HIM0OhX9YRaW8v/5
UvxKm+1LBuVYu9KiQpyAtTd2h/tTjQuUPmebcwOJhB51A4s536TeW6CLtHWctrK2Jmk8f02tHSjM
EGft+mE8EjiRcxMJRrXny6pYruAuV/zD7XtaZiMrcCuilV1GjjzrG6cVQkDrWV+S4BSPSklBrHo+
6xxcUpQKAJavx/qlehn+lPL9TpTxILg2fvKBvBGx2Sr3937uJOilP9GMgGcs0bQ8oEOCC1y3FbSe
juMKqTqlFDOzIWRifLlzPbi8WdKjnr8BcDmBGHhAsfdunCnjFGaAHoB/mcZxYO8buB4lkwYojYcw
EnJfAsGw5QlX+nhtCJgp3R3AOOUoJ+8PZna6d7n8gt9e+RINm+/KhkPZCFAemt5BHOlgOWZUU8uf
3dOwxPFD6i0OV1Z3xM1nVHodiUQNwKI8beIRAgiJIrUE/mDRqQDg/VvRW13CrGQxvYtRSYhi6/EZ
YCsj+IG6iXbyKcFSymzu51Ag/YeQenEnIJ96L14a999fmaVvRa36ASAZ4PRufWhH78Y3ZHfgfldN
1KRqycCVmjJvlYSuZfbdXDl6UUfhS9XPHy4mycXrd4UX1RLavRtZFx9RrYdBxwjXnm8M5D3QZfKR
koAmOaXwTU1o69qLvSJZL+/0kNoQitN9eFH3getTXGuQyfJeZxbcBqE2dnmbHWfnMHB8FCbzUs34
fvLb1ED8TxQlbVDthDghwZTwPGNTXvZcJqLUxqpXUvN/SBEZPYzi8WsWYxTPOUcn8fvIuxgUxXLP
vy93KJjzspSGCaFqqR1TPJeSCHds/89hmLQ3uvjF040Z6+6UOHjca9bORUZJ0UKPc8w5rEdpv1cz
ikSDJYbIUjSdsznpHmY9NxA8QA3UyWO/NOyLRZe9X/Ij3vDzPTVHLe8G+PRBpzhFkCefFKp8Cdhx
Ir3t2IYMVO3e/D76QxPacCgetJBDwXVdVeo/h6QbWsO6+Vm1tl6P0yMWW/0EqOFKEPBIxq9rXTum
zhYdh2KnuyWbJ6RnM8vZitPDZZQGXgXD4wXhnJcPhpDT3Fo9QX4wGpVXknT7BtzY2XA9+my8QP/1
z2SDh0NkuVFJHQBg+RC9sm8zeFId5PtAHk9TnBQLVRm1ZQ6/byTra5mLY9DeLC3I/WgaqueMo5uN
HQkeFNK5uNPDfE8NXUpE7QDwGBUQ0y5WAUiti7TzghWNAWAKHEDGXTn76TeFZIISUTxArC+8fboP
wz0ku/07ce0PejoDq5HYb2jHAD+GuvdhFEPXUdtKG0aoiassFNRAsw24CADfi6qlHoj6OoCwSo88
XR+SuUOiXQaANXqZC8xtclcwjTJud4uiPL8JyWZ0pwvEtPzm2OEwKX/w7O9GrrpXK3GxhWxgqPUq
aHVodO29MlN9vnouAeHu9PGo2KSKD3AgG4o58r1nbo7ILjiQtEYpovuYM6rifLMDvzDHQklE1uSd
ERfE0Y4mRodMgENMOt+b6RtHiR9le/uWUX+ZcmtOcf3SNexHWm+nu/J1puaw03xZcus6D8RTk95M
fcwwF4HemLi4kUx8m3NacxZqMi1YoFEylTnYlOc3aDNmDNPL3sjqhCgUqDpVCMyTJVFxtvAlWXFF
yeSb4m8S1rHtBJFdx6ks1EvrAPmCy+GiYaXqrZhpLPKR9QVdK6Fu45TjGE60LW8Et0g8YG45poSi
wn+1dZHnysn3qrgjrhmOv+egzCgc/Y1yR/xx9i+I1dD3STan9Y8EgNvFIfXZexAW58gEpIFRF5P6
CL6Lbuc1WViJN1cpTrmBNuJn3QAcPHFWCXi8CJkW3b8yL2HIwsEaiEIcRQVvqyePcPIX6zjIVgtM
nfzBH79wKPyOFLz7SmgIfzCcoSytFzMox74squ3aaNbvG7e7cC42QpvQfp9PsmD3BNF9dXP4NuXm
PIT6cu3AZwdNmlviLLwdHq1PaTIXgFDd9UphdivV0t1HwP2kTMSIERWqtsniFRwZMw8gU4IwlseP
gF96JyuBN+qj6/gO8jMxOaYMIPSJu1bQ+yXoGIg9JkrDh4Jo/0ZMF1Fa71IKCynqf/D8Ahh/wt9Z
UWNIRXpq+B1VpeW8m1pr0DsJyJOjM8mr7208s2zumH9Q7RHji9tPy3wfGlTW7zDgyGPii2mjioew
Se8J9+U5VsvFPlqw8E+prSGXL9qO0OySvAToAnGod+N9nBAy/j63SBLPpXdGXjWdj6stK2xM57ji
9SoDQx8INfDHMdt7dA07pF9uFV6E0A3pHMd6FyD2105g/LFrw8zxmwGCMDnqp5d4pCTf76+NJ3Au
ia43n4TX3bAy3kpwVL4MdWyVobRjNjth8MdZPMWepr3oR2E+DAwb/pLbSN2PcgZ6k1Cv7UuvnQFd
JVlFaKSPMCy3WGE9owqPNBwcUAu2LgNgeeLXHJciURtx5Cai6CSv2R2xYqpZFgsZgcdrLUZ7g6Qv
3X5BOyR3/DgkW14pcjPbNJQOYOoTIWOFHw5TGKyT6ZAgVQZIFwondZu0M1amFXH2pDc4Wx3VwGSW
iyIoG/o6XIr2ijYA+af9jeVMARulyJitwckCYVOdizOzVcAXElKrp0Iqjc6EVtg5pv7J9+wXkK4F
No6F4Dpj/Aw3rZGQQb22ZHmthT4DX9cxz5ceWUrIBDFsoWlE1UNHOY4dDlQeniSEh+hrnbSbdkE/
mETHAuPyzJxSOg+JATuPLbkYSwx/vtveCnx7gfiVpBn5GCu8CdGtkykdKBf+b+7nGMalU8a3/MdQ
Ln0Xa/bZvD0yVqzfau8JFqWDEc0+ZjmVRvr1iR5UxJmFq6SnLqouS4HXIyaDbbL7AZ3uRZXJJC94
IkV3VaICgJODmIdrHXGPNBul4JQ4X0GPHpBnO1DeTmSwsK1Q7nz+3q6leEgJVySDsMfrsgbKlqth
pjmQcMOkVXpnWiaNY2Ycn9OTtuToQQPpo+Cj62LJf6qm4mNqgeSwBUYn+soVqafDlL1auHQA+G3Q
w6DmX2Cejy2kL3ZpQ3U/F7iP1dTngQD7P9oxBLKZXr6XHZV4Pdjmc2fb+p6c6F24t7pBpcH2OWU1
rbVzwQ6YAqCsfE3mB7eyR44JE+QaM3WLUWcmgi3H6CQ+bdvqZzlJUGwGKoVyv3vxUVWMHivvNBX9
BeqcWrXFevIDALUBYH/nMsDixkbfLGW73MynOSUUfExqM8pf9/xv9wgOyqOilsbYwa7CnZxyxFl5
LMyJwKsVoI0bs8ILnACrW/hfL8ImanQTnFwlzHzmWAjeVctlYLxQGHgWkPdoQYOaBuen0WYfSHLK
kZFWpmerRXF33niyOGjOTuh/tAK6bqJMaCznjy51WjY36mCZ2pqv9KbxdgA63QTTIPCHNrC690tm
P/M4jRTBpbSZe0n2GpsDT3kC1qSenZgQZkngjW9yr7GAd5Dj1pTPy39GVqOX5bjWlonZ3347dYfY
pQXYUm43klY40GMj0CVQWd8oA9R5oWwKP5KMnsaAKGX+yHjoDaZFujNwHElgpGEvSFvtDUXHMqpZ
VvRDIi8n210lWA8wwmUTtVUkBZitZa6tA17KCWmBccUlMXqWp4igRnPsy8uMlVCOVtsMEH+Jc2qK
IA7k3bqijHXdrKqqrLSN3MbcjAeFpB5dNxLrZie466vXtoM4AKYv/9/l1L22OaowL83ToDJQJCjW
qNaaWhRNcl3kdnf1tsMbvAMdiT1aXY/Xl1MI4rmgTTkpLtiyNSCMT4Lft4IKGb1Ht1uDZ7z6piLa
cOXztawCzsv2z4qkMYiXuSyH3QozA9TT2M+SqVAq68lax4cneCVR2KqjuszBGXA3M52LlkMX3bbh
aP8RXDZfeKXQTDYaCEeChJCc9K3D3PhF8W3Ciq7b40uyHSRmBSNwzkJZfV/GSMNYM46wq2yL7r+9
nZLm0Ct+ThRZMjv1IinO0gK5VSDELUFltHl0UNfVOmhfHBJtxxN7GybQJJqdnuGhFnJZlBlUP9AN
BfBMot93w/rDbPW6S6qpbSstiMIfvFp3L5wojFptDBPbmMuIFBmEwZHTFr67bn2pz2oM+34cn4QD
myiCpU6inJQwGGGq1Jwq+T+8AgM/cuHE2GyglhCgNKtPSBj+c9fJmqws+zfIgGU9KuPBS1aaOW9L
JLXnbirTXpUeHs8N7Pi1Gk1GKaysXjpPmYY7vKbnMrjYHxGJuf08QwTVPSv6BYXUPevDVBbsyZuw
SsWf2TsZJpYxYGCcn+/AQGgS7mF5mR2dZRaaZpqGkyRIPJm15/4hALamgXieNQQ2AcC3m9Amrw2G
m8QUZ1Hf8UXrfhJclfg/tf0deW6sMOqdp58W69luXIgMOPaWi2bUt4+W60MmvDD+KVTt4Q6yVGA4
11ozmX0n1r1CJfelVtsmiNVsjVw9np/8AS5QnWkVy9+XNssDjnjzfByMqgqVPzMW/ukizt4VjvEm
E2gTYmosgj0Sm02CRWvSlWsqyqobrWsUmTltzjUUX4xhau1H2wM0uyjWmfIggqZeCP+cgu/SLsu2
QnQp4qUzeNGhm5qnunfO1eq0C2Q+fHYoWz41CloVKzTQJ7w3D2wPgt0a7HRcfw9FmQU70QHEm7E5
XlPFSHUpeIWaV7GKB0/KL9AxEOoSNqgG1EndRz54Q/+xexHYtY2rNm86/AWJ0GPcM/GxyG8Gkuh1
QKbt5UJ09srcjWqcqIbNgKwkFLgJzqoo9Dk6GMbxhaD6P6C9v62rPU5F73nwB8VL4ejZY2CjUkyS
A/hV/uWvWc6rw6fcJP/fw+M/d/Bc6Ev4yogKMU2nwf1IIROVCqJsKiwb9ufOtPXUn1LuIFualkva
+1TPqTDzU02IF+lExgVns5QexT/EWMRyA2IwmCRkT8d9vIqLcItXQiV3n8NU7JvBTZbMQ/sBYg4T
pg5vdtyVJh0r39rNk4KIbmJH2vhODbL77vuMRB3pkJCUkQQhoJvpyj94Sj7LhreBjb+ScvFPSAhf
B2KLq0yWjdpZS0eiN0GGPq7dC3t/LUrgsoVqSbYYkfrt3ocgUyPH+HRZOTGu7xz4pxazUbD3oksk
h0K+9eGB2utDp73WmEycnVk8zbsEeJNdnNe64l1tfLWVpmJoGuM9fYdG4veaeMaD2tiJUQBRe0ze
O60EtQwjWuqEb7+ZPevXvzm6gDcv8NM6w6eachvJTVrDNIwTlE/VkH4V63bPiaGX7j+7KxHaUAyg
z9CEGirYLhpxjooL4OdQeqXidOv8a/vbKB8Gncqv+WXvzeC7Eg1jagiScv481W04LKtnnd9Q5Q+W
L3BrGupw8fBenA2e2mph71sAmhQ4tBz0wbTveTDBYYwJdj1elA496o9472IWk27Exqjo8rFBG4XZ
oh/XFjz0ZTZbTVlyXK5sEDSGEAX6scPOdQeXgrX/syJvNp53DWrq4Fsn/nYTRDr2YDCoVFr5ycFB
GBRb/Wv7VdA/qGEQHmYE5bUo+ctGUiQL7fwbgQprWhot7e0+C4uFAjNlU/xhpm7yNDhkYbv273KU
AjAs3VEyl/ctnF7XKsOzJ9k+J5z1r/Mit4yuyw9ckuD/8U0Xx2k/oqtbaMxglaV4+DB1YUY41Voj
68PuD9SsNAfFnKAORdidBye/q9KuAxB3AD4sReMG3Q1wwPp1S04UhOqHa/MZGom/CLYKN2zquLt0
nHxi4XlfOst2xWOQbe1XE3IYLMD9ItwcWmnliqHbP9NXSXCru6vT1n333rIcsouHh/QBZ4nsurR2
CpmnqBtEY7Kqq33guuDu7qaBxTfw8apQcatc5ave51YGfchmb5f9c+I9tQhDFIiCo2P7/qntJFhI
H3OnQ4sL4TF7eCt88rwpWn8rm1yRWiSb7jvsmVzI0sXn9wJhZ5drNahPdRJyURFYjqYzPoQvp4O5
Nhu0TY/0wkxN0sjK3+LbDY8RT1ATSS4Jm7+nDVPtbPKK05aXnGveDVZT5s9bBF4JlGJf2OWRfUPl
jeduewAWZ0eiCwEZrNbuLEJDO2RHm1qTpolQZFMvyER9V/rJvDx9TxH563dCpDnw6y0gXMnH037j
7zv87cQYcWoRHO55fFERd3SmK/kKfyEViFXq99GZkDY0w/hRIOS7xz8KSQqkjAxX6CeIMEea04JX
wTLDn3Hq7WNMzTgEMvfgAoI4mmaaizm9svbk+6fupVG8805J4hW9ZVW5yt6K1LM3bygOwMhQs65A
E3KTtTGCHZ6HcJohS/8ZSmArCTVwBlnehiAXNoRF1aKGHfsqDfu+3Rc2QgBWnnG2ifIgGDymzLAX
K1LGf6R7dPgri5m/Vf18havWop/sOt/GOGifZF1IchV5d5FaX4N8+0kbU5cXgxBOfRY26jH0J4ea
45y1xaweBZSKr9AGcmbkHm3AuAPbxVlUCBBoGsRrg4PH4QXu49iQfwRPhuaiupljwo5hOMpG7R25
2DXS9zCPSwsE3T01cXzgPYvsDRLUEFz4xysase7a4+/EV2dNLUX7g6Vc61bSvjYoUy6gOitPa4LK
FuhmAbormOcThqQURdERD/2DOQMdwy5rXH6e3Hd3fs+nwPFfib+E0zsMlqJt14xd1z3whGcyNrM7
BYpxkq22awU9VTIKzY+d/fszAuyZeSQs5hplWcMeMAKhltzC3zbV1wNxJW1e80ss85mhQg3UKZUE
2dY5+ygNvjLzvwUyXL8FIaL8ZKnaC/hsrAM5oNB2vyD3kc40BRu4zhuVhOH/IfzQs68nKQ47Sl0B
16n/QeyrVOi4wXng0W9adOM68cKyK49JXkWgfTEfNseJ1aVY6zsEtgeXYIq97+WrWHQJ3IowjCjh
Bg67xbQyoErf8xqalV1oJoK/dJRsVrMzvJauvOV0WFRocweLKxZkt2Xf5UXPtYwh6QUkQGZfNDr5
2B+g36iF+Cx9hI2Vs+orlojp8QyOWpNsG+pTMkn3Vj+BDqP5Ux6vRvycJ3YiMaNnWrfTXlN2jxId
uYIr1bcrlLRDyj+6DLmYqkIf2S4B0LQ08I055A7KKbAuWqXFhvSP763EqQQvd+8b2RurRzdkcJg8
Ss+swxCfOIN9Zx+qht6O5TJhY1ZythyP4/e6L/7y2jZB/Riw0oz8L5W+VVAz0V+s4lQcWnKTKwwy
cczud3RRCVFts9GuIi0A1qbkZEE04YQKNneTEyUKUeqRwqhIrCjYluppKQYqYZISBt5OURCwpUnl
N/t0VjvI3ONOUY6NQQLQzHiV3J2hP/v8xA88Q07KWt43dGVaThc5okHCgjDJsv3AzX2lpP3aPAjR
0nhQlzjFuXogEgyFE127+LIU1H9HP89JAInYbXKD4RHUgMnS8+eRRIU0dml+FuN5nt3IV34EpU+x
XxVlhH90gSzOuHOZqKae7j5rrl42ZIqQRYe22qDzmndp0/XuCeToAcAOZ5WaRGD84JM6KqdBYUSB
GtxI/cIjh6XBSnciIuBhKPeDRjHFCmx6ZueL2sMSQMfPt0auIpE5NhGQIk6Jp8sOJb7wKFJXpM8J
Zh6RsT0ozx2QBJgXjF+CgkMICy7qEn3upjPKNTUyUJqOZ4vlht8T5hHqwS41/E+BqI3Psf/oay/G
dDxqbVtc/0G/h98JAJHdZgn8Klp51cspk8qbr/JYwN/6if7wRKNzot6/JWVss2sbv1wJ9cFKvQwU
ATrUYcZwqYniR76j5wzgG9fTyHm/Gtm1MZrBSJ+SmW0hUTcLc8T9guqIW/UnA6wpfd4FG/Pa9rfu
e5pI91OZM3w3tBPcjuUfqbnhvkfektm295elrsSjHvfNZzmc2yTisc6ZLz2ksYvJEid5phPsuCdP
oG5uT+IfTa4U9pdOw9lcEPx7IgCYd3PuNx2xFUEWGJBFCf/ly3eRYJf5muD8icSISkz+l0ehzL3W
mtJMLl+afNWVdF+vSljzr6VoV65TIdhy3tNDUU86pdAMcYCsiRfu/r3LNhUogzIcTH14eMHTB/mp
x9GHR/gslqu4uQ7jyJNgUAxE4/HvhhM9CkT22xhIPkUKEAAYJRWPA5IGTmEUp84wX6o6lOs2BP8n
BFOYM9MhfkvLcoiUTe1QtW5D8RTE+QYHiF9aRq/Go1K162DzDxv9A0qV34mhK/DJxxrHtO7HvnHU
5H2QXk7GrHrAHZkM19sALHRlcqUgZFLmvYB2lnoSYsFE8DJf7mGkkcjpjbkBOgWfSzZf3pd8lAw6
kqsSM6uO6Vg7082XVFsg+WVDjhAqi9NDYZwfxE+mjLjUJfrbh3IwFv5m/A9eCcXFVWRhFMfe8/AK
R83B3rf84Fxqme1+0J7BWuftClmo/RtJpNF+7DFvldc/8qfFcGn3jpdO/fscCNwsRlAe8Swa1jaI
Y6qH5pHMZMPN/sCrZJ840UrKv6jLQ60bq1wlImsofkZR71eUfWI0KK2cSa/AqjR/9Q4rLRI6M9a7
hGGUkb+o/5gPhUORoq5dvyD30O56wJV7Qsr0sCSUbsImML1bXVEkNXGlXD4/egKJEB6YOLTF2CLZ
Wg9AJ6hrJK/SGISIV7x1QHl1YubnwAHnkHX9HGaP8GR415SwdGkTxkzci8ltkdim3S3XbkvGK4gj
5zYTM4NPFgtIK7Umob/DdVdzYA8Q72KITiLexkTKLuKJuW2/OvknbMwEXjvB99AP8iQEwrgR4Tms
qJI88ygn4Zh5Y5q7g04nkXarlNatEVtBuXwgQXpDfaYMv+DLc1sfwn2oJrP0BPKqYoyDKgx8kJYG
w2ppDC2p8dB4qoczIIAFWmuIxQAxDEJ+deercZORJBjrDTpBNb7kf2XxgpWx0+tcUDW/I4m9q2o7
DSdhe184gPUFWGJZjwinMcVPEIhYNWkedjwiL3uED+EJgS0oMq/fY375OaITKzM2b+p7QnqSKXWZ
TBeTsxZ1LdTf+3Uhu+LZJ31I2ifi/RLSh+JfMhgXg/XNne+9VH2WUdx9BoQRLB1yCHCkPUpY836C
mlNfZNeP4SUodaEKqjFaKy7e9rXGtXrB8mc48m81fUYXcl6WEu3YKd0dTsKL0O4HgDkrf2I1sJZK
HmxMGQZFhrmk5ic0qWwnCtELoutYxjfO0OIkZpGN2uxH8VHMiagtnUVIAOpd2g8uuqqkajmE1czj
AdmuojLdf2UUDzFyFWoNtAsymh5zhKOhYgh8u3q8OE+uflQcXiL18QV3qrJJoWX5yxy//agFyT2d
QQSipOMyw5qH9KkJb+HAaco0AWz8xk4Ovzjo0xeNATsICClh+0RSlSiBpv7fCh2x6lIbQv/b4Xrd
RA482wUtsUkvTjFAoOS8e9kbFgCiNDLys3ufoLSeaUvQc/yqjWlGjW0/ZIb8WWVjc+QIxcycz/Nf
Bw08EEJK4LLg3AehrxU3XF6daIV+lnEm+aJ8e9I6HGPIo6sBrKusRBCApW8gOJ9xKqj9gbavyvEm
BHqfmLPqA3z1HBslGurfmrS/Fyr3pUtrtU5MvdBaGL9neglUcOvo1//IDZh57UOPsGRUTrOfPr4x
GKsc5XR942HP2EM4DZiCIyQ6zNQC5FzEFvsMOMolLAbz7KdxrjfJqIbl8V0X4a/78DflqN2Pjfp1
3zh3dKkuhMBOBmoZt6g6DheghiHO6pR+TCp82IoamocEZ5dO/O0qbpXlFAKafgVMkXvtR5Vdv2lC
vuv/MqqIe1CYk+yhshA3gcioRGyRd4T7/MDT7fE44TGkwSRn+gVAfOcEsPDVP6DIuQiw7HbLZBBa
xSVnhYwhLdKUxtQ/jbh6anN9Pw3c/L9AvpRlbJYxj4Pgv7B72/OYoxJg1OMxhc9XfWEmlX/kSZQB
bdoJGqHCpBClwTZg5lZMFVe1SLeoRs4puwbknXP1xFw1IK6dlkY7dRehxifw70/MOYbiDNu/9R6V
x8KjGBLKeC0HinRa2FfIrwIeU+gwV9+18vZpjgOg/NgGFYNmttM5LfYKV8zk3Kdc71fiLNEHzrvI
84LDLcbiAJc5oO3M/2UWnibpgccOLkHvI+oCIG5TKJUFZied1/N+W9TEwiZzJTDE+XLfUTxQiLWf
DTL7tixcQDe2lduR/SQynEHMXcVI+hHOj2GCfyzznGFXBLWBy+jdNQmpC3jPVfrbLl1nNn1JDhrs
1kZ5jbHonF3/uTiXNAhcHP0Emjrfk4P2w2bRPNNICEngeztD4tJzY81Ax6cn98uN+SeVO6IFcJRU
uBOScVgerlJS7l2urtKsEyIcV87qYiBf7OLUPK5lzKThQVgVJDnsE/I3BG5bQGfULEeLsitNcjOC
eTZ2AwmH+gecsSgvKxGBRT7VXRLVx2sKRpSxHXASR+XKZ+AFEIiXCaGjah7WO4DfsA6X1F5AWOUL
8GbrL7AM9NEIJMv92dKKtFnolhKrXmkQyqIaejvrdEJHNqiDf9LqCuGbIjSSSWRO9kAG5VImyzyQ
cdl3FYIxmKCfyk2Xn7lqNC1AnOD5mXKJrtxgwp68uYOd9cxe25rpx+UbCjQYOvYKQUlilqwZLR5I
7OtUn01xY5pa+cbOQKkboP+7gPFLs9HfdtVGzveLigDb7zXEdephWtVk+AUClJQ5dPNTf0HsVLJT
JjU5r/xV6wYsyYdnxzE58421+3BTDJq9hoU0eGT3mSBlEs3Gj738Mc5cEY5FbBy0DHZM4tjZA2Qu
1qP1+vdoVERn7yL9GNs+Nj3I0/Xyc5Hk3ZA+Xm7HIGTNX1zLTjmYPgnVf37+LlqZsmdKprzTu5s4
uxvyWfeSQB2fisqggpeANraHKhe5+RBXRZ1JDrDmrfLHLdzHKcTNIzknT4zFHn74KIeg9zwOL/PB
XX8qTaCwHb35kNSR20GJatF7K+gGxZWoT0kNJ6KOWSYlmJFuiXB8JG8v+QtYZ/pnRdOVGG78Px2R
3GrxHa7bVKfaxBmJGuqAdQtUWXxMdV/kxT/zr55pYBXAMrmpSatKiqPob7HMWpU/ceOFmgSBsOfX
6aVrqpdR+OFpvpLd2BpgV2PkNI+9zcxJnsSJh8/skRzFYFbvJRfawC9oTbPkh+LStCfv3y+y+BVw
Yp9os24OCtLy7D9CY1BRK3MECOKL1o07ZyUUCiRntTGl16infp046DKATipMgdFIJuyhylszvy9C
PTg1nax1IbGMEUZO1bZl4KL1o9Uivcv1gPcanaRkr5KuFpIOI7aQ+3HXecVcc/7QamjYixKBtdTF
g5xAinz3kkdrQEO473daPfjKPwaaKfFm2owTCjiHPMEC325cuosHauwpHjj0gYI/p7O3z22fsNBt
FMRP+6mjEuH9oX8BiPwx0y8B5HXQ7eIZYKiaCcQnItK/wJ0oZEg2QivpQ7u9yoz/Coh/8Bs2Fbua
B4zq0G/ILo/W0FKuA7PZSi3bAoFbK9pU2nKuh7VN9pdrJ1o7OVqRICBkj+mWINt9v0MSJxoOPdJX
tqcsvFIPMxDXYJwkke31pmdkh1rzssV5yh0kA3IMfkmeKf++FNQp0oFY618kyIDIOdI9Bom/wgXZ
xoc91FJvCcn+YIznlG6NDiCpcq1fap5iKaT4NbCM4kKRXcBb9xeMg5nJMpZujlYnAgZ274TDFELu
lwg/4GkIHokNZIjgIJzUDNt3WvTfEMsprGUbe1kpTiPDBgLnmFKjdlERqp7TKsW8oZSR9BJPvsOU
owePqRyIlniOzX60wcrbIHQoO6EmSJOW7K3S0Vfpar7puec0zhCN0rZZbrFqMMx+ugFFVf7eMuCC
yhTYqpEP3qsyO92odcJff+tsJ4Oej5WQYEgE3s8e/rZGxy8SDkMtjXfAmC2Ky3ANhf+s//pTilbs
nC11lcPQXrtlOzEG8FuFSOaLmYxaGlm4fb5JD1mwVSR8NKGvWYhJMY1RxfucSw7CDj2AeS/5Pa8N
nSABhZyRhf5i8C4zeMYucMFAnh2BvyO1O+ZgcMkfM/QV8beQZA1ZrXwmtR5iISXWSO7qYoiIf/uz
aQwdMOuCU+YD9ADcfaF8B6d0fcvw/u23Ts5T1xrLMOB3/rmal97/942Hgj9A/BG+ISamAs0KwS0l
2II5q7zUhJkYDlhYeqlrvly7foVqipQHlkhCkb9+NNDjGsNvxoTN42XRsqjrY3FReVa2G2U83TEI
CCHFcZcnFZQHmaTd+FUN9fA2djBroU5LsLYr/c1UYNzHaAIX0sLwtBatNGREZ+8BxgmDjeufD+7l
t9/LHgaVjQdmKI7N7ujb7r/Lq/SaU2hcPC9u1QIEYojH7g/DGCDz7Ibw6qA6Fts1cSz70cZpn0Oq
4saOUU5MqW/Wfvrz6CzyNUdXQx9vGr1k+BXYu600xJ7RZkjCj+dexRtDgWlhFv81CVrmuCA5l+Yd
OtLBExF/Jw29V6pMC1elddcRhbwIafoNx8yTENYNR+dfkebKaBMKfZReo3o+8AP3p8jPt5ONJHP0
OhvGRVkrWASsfJ8fMZw6Gkc2oFojMjD97JoQVpdQEzwfv9/05d/auzNlp1024kMwD8QjWXhs4tYr
DAh04x2OqmRZDtiSc4MKPU8YRqY/RthM/+TTeJKNpreUjFqhTOSkhiOsdWX3IwlHVfOcFbJtzNSM
UjZ1pnOsKjoczHCIRuxI7AppDFZ+K+z3abEVvS8ZE8BUyP4AV2lv3a8tY/ugFn3EpLgX0FrORk7M
ucZ4S4eAC6h9jymFhtR3ryfhC0yEP34mi0j1lmFUHzS7KKFZZV7GtfB8+XlX968o54W1LcWKQN+j
ZMtghUxb3aUaUw11TghUAB6K7gSDdDqorXptYxP8NnsdOTdgrnBiyWaQYwSCFk29hfqE4iyyZ31p
UJXq+njt1v/wZS2Rk0mH9bmqrzLB9do5rLb8UyZiQjUy68aeQSZnCfj1J3ISxGzvcNDQ5tHkwdD7
mMj3npKD0jEo3EFhi5xIlJ6CGpS9P26NAQWdkHdb/pQwABWl7sSR1fQUC0jF01HE9iVaGTEERI6I
pqlYKW9t2V6SkipJCwl4R96h7+KRBbdrV3gBG+0YB1eEsqhEmWjlQlGyl+xaMipvqJGHv5oIfXlL
k02gEIWG/xOVHgnHd5qD4z1xxgJ6odJOW/FA2w2DqgY0zlVdmA2joKdBxX+dpl/EH++wR/O9Rtqu
dO6smH2XUR/Lqt7mV8Sh+T872dDDAPpESxCbEotJ4cEKxuATJxI2aFfR/JeoUQqoT1RidSgyMVXz
mE+pwCI4heaHvtMOHRTClDvwyTpqjGEHoGBX8KFnwTtd083ofTWVzme+J12yXsWY6ayuz1d/SGea
nKvNvTRgy8Krds8ZDnJGFH6vBZPlcGtG5v5Ipk/JBi/JWJI9tXCsTkTVbwDq857cIqI/DIpZGXi0
CQ0wflXgcRjnz8+Taj565USgjb+UWU6EC4dqAAJ3g0js6m9vjtuN1cX/P94plp0Fse+DwZBf6aiB
5K91T406T9tkEtMfikKCPorXRjS1D4cfTM8cAhc1PHtW7XBkVEEcj6BrYuMb44SmLc+x4FkvnvI1
yrwmpNi2kelc/AHmtrpOFCEI27mp/S7hF7waq+ZK7EWQI/VzGSW5jCo+BMw9Ly31L+yjbJjkyvER
WwDd8bu6ZdkN+rTRzT+yrstOzzDmpodPTl/RRAkDIeaeDLJE60AUajgcXYBLzGP4/dJm4zwMlQl0
WOK1sS4lhZbirI9QPRX2HPf919TWLaJADZZ6hUhdNlQdgjyza77VgdwlnNCFy9lbPLatLcxZvblF
58E8yRlBZx/Zj/Zx9BpEJQWlHaimsGETw5FkKWsgnq45iVyhgmC0clDOYblYZosAKpqPP2uhOk8o
RbggsCkduDBUoNe2W/wdksfMqFLuXUFDjfOnfzTIqgUvvbsJJmrYz3eb/2jDpDAG8wvW76yohvLX
pBYphxBBGUrW00cn4vXqdd3CDJg3alfgO72B9x+3fiXWf4WSMF3l+NhCYtrn3OC7qYuhjIXrcGQn
eloXmaXORzcFyP2pxXJUjU0YVuwOz8oVmXf+pmWecIuiYfhT/rIkpmq19iBNZCjYrOnF+WynyohC
rvhrbNQoXCpeaRFKdqdU1uuv98xniZqvrf6Bh1adk6kgqt9X3YcqotgsSuOHPXnNrdii2mcod2oD
lRZDc7X768UX3DgUlANajjTFDHim68scoezTkGjVz+DkodOwPdq5TpraoNglnbGUbtkLdQmtbqPA
2XrKvDFdwNNwCPv293eGF+VClVzJrV1Ly20xZnGpV33XWeTZBHEWhMEKiaK8qdOxmHpFHAVO9R4X
tTJHOohAUYHy7cQDK9IWW2NCQ4A8x+zRHLTNlN7bl9siG6iV9LmtdFn3koADFih+DyCD6Aj39kYg
ee/m3nU61Zn9xO1hgcTxy7t9y5L1oV8/OYCs5C89x6klq2GtTusuEW/3vTZKWF/BbqBCreBK//X6
ePGwrXe/ZSVpikCg1AF8R3d9AmtGvdOw0rz4coMF8BpUx6nP1zLLFrY7c7qQDu+dRY8MnuevZYzp
Hcl5/ufRVyI2z2jKni7y7W0BeGxrRWB3kTPXfYbzewYc1y1j2ZqdDNBWnFOpVFObdItcO3CdWAmp
Cj9/eTo3mOW5OhGaqB7BHN1ckcUmBu6nS5iaxOkp3a9gk2rEnWxYmL9af40aT/95uW5+a5jc3ifd
DnvKuFMM5qa9GeN8nGceY6/G/RuAJuBh9cCofcJIhPULVKuKdjqCTu9sCiLW0c0qJQP4OJM7+S+y
q9xRuesMzWCrXmQgOLuqPYPbAbo0pBzim7710w49B4H1hZZmG8Y+dMZoZYwtoaX6qUgCmCcqydWY
erfsm5FC6VPNhhoL4APqKp57kwKVJ4Gl9nExet1iXF/rDMoQHEfccuYGesIqk5rIufGDZO1Qptaz
C2v8US3jdAr6zOEGXgtuSzmQ2IbncQ5Zrn3vvuxeq0k/CNMivZdYT3hvu7PBZpRa7HhZ0uN+zFUJ
o3imQihAp8X/05Mzx40GnUspnk3cahKWuJxiYf9TpM0ENFM0MM4Go02vQJqDjO2HhYHsHuT5jx43
EPeXUJLdgs1GV5p+FpqyfwkFfr/SDsLK4j1M9aeADaSl4x8l5fUWLAcRjp4yjhdAEr9o/N508WLL
7hYAv28wGtLdG2na7c7q4NSakN0d1zTruxzrUHTByNKk50xRJsQm90bD9sskp2qXfNS6EQxX0bwS
yZc8IvzijcGlNBPrfF2Aq05y5UaHlkv6WSTtMfbsaLBSwyUTywEgwfs5rZVIIk5C+CemyLBTNHyd
8V+yTLvup3zk8PfyWBeV4EDQLNGQpr5HZ5PosnkPtot0I26a7+1VcMaNA9PipsAIqeSaQclSEuv+
Zr//gqxQ6cKnWGgQh1BvwI6IkL3o+KD+JKLlwp5FS5a9TOqouM91UWJoAwpvPR75paNLrkoyviZ0
9mTgggtwnzB2Qarn0KiRfeESfhKpo0cNV03fK9ntPqdlf02SyF0DJXHQs5P8UwhDkTABgaBNIL2c
ibjbvRr3wp8bLuazzw5KiiyR10Dey2jIjiqoZG08jlGWY8q4wCTXXye5+r9t33XsdRt+Bt+BSxsc
J2eEPq7m8bCizFrrG7f4baeD8NMNAChRdczIARuocrQLr9+9NSEE8a33SX0e2jsMuEZSso1UwtAM
N4nVe+V1e4s7UnlvD5hCZV8bQDVwdFznhqva78tl47ImvYombBdTBY69zFrj/z+6dHv4R+AvEDYV
yNmL9h5xbh5r79xBv3mMMlIeyjtnUy7mcEJUHVyf8BKJytvCUbjhb1Zwqv7nmbVzCBv7+owf5JrY
PBFOiXC0qcS4y60KLNlZJ9kn0yJbPZ6Ji/qUzWPqMe9ARj2F4BPV/NRP7wVw0ubIfIqKDrI/Gqj+
3Y4qnCPP3QKC0fFmXE2/LB1RSAQ3jdsn0HdBn6rFFNk6faowS7I6Y6fd4O5CyQkwLlU3IW8lfUH3
Cf3TSNqC7xrRjcRjMaupSyPKBMSM8G1jgF4dYfWqDY8WqSJ3Y3IW9n/W7myKWb5KGT1H3KWEFibt
xSJbxqLWwaNcYTNhJUnKJCjJE1RV9oDx1XXEDoB9fXpJpP36elpdfMgJ73HU7zgLUoLDYHt3FjyY
fsQaaBAZKyelO/5hW/NccybIdWooPC5pNVaq6X995IIYRxTUPNfop1FtfRL3LIvJh9ds6/NMouLT
+PaH/eKMAWJ9blW6SPoSBrgpdGJ38p5UywaEm7mSNpPPkrEwhRYKGn3KXuRsBtmLrc7u3ZuuyRrT
0VK0ONAFDFg7ERPpC/PHUtClohFXLuu32rTz6f6xOQ+NqPyeoypPEJjUNUhcoNBxDTLoHdGgbs2F
SFkv9EGZqfJmT0czv/k5S/yiOfV+aNn5j56dcw0b0xYweuUKLk+R/rik44BT9IGW4g2zlooehXJC
kRGNDz3sf+69/kAHNc4ios7kxtDkDp4q7ASI5n2tyKhR8gUQ9L2vIkm+caGkWoSStD7yzpAAEoZa
jlTN4nGYuiSQ4NsqRpuv5bZmgqUIrFWBEMVhl/Idjk33wcno8tQT86nvN7Uabs/EXRg7wnvybzmA
KiquzTFzUCweZol0d1KWh/pHQhgWzpGWbXbH5W4X4BVKhZ3mWFcKluDa81ZS//hZIgVZ3pkC3vp2
0nIoISGMdxSkeNsUBqXe2pMswpJe9rR9HYQluI5j7D5GnRODRGHxF/zafi9csdbZuXfd2Owa9Yec
mslMms08gIMCcnFKFqVkVPULcco5YXDomNBG52iWWpMUFxa937NE6PtlMoOWzuOT0330til4P9gy
MqzettqbvpzO1kTBqCi5QCN9nSqh6wXYagtPpc9hdsmKmnyvG2YGPYdzRVL5f+795h/yyfq7bDGB
IbvKZLTzbVO/OMdQkdzHWsrjvhBhrqo0SzTwPBIYtWaolatx3AwIM0RqIZ8/VbDien1tEFDLcYRK
9Wgi7YXAtef9PlMRaviEH9H28by6vUirGLPDf6V/GFhN/a9vRCvXk1pfx2ZStDTMFoMub04IQHV5
ynCp2QX1QqrBuiGvKFQy78rMd1bOaNMUyEjB8bx9qaypzOUwA8b7E+Oymtp6hrFCOnMYSZzFtm2N
PSzXSkDepuLnvnjwfIF9Z65Kfg8XEJqMNVDUaS6Fl+KAPioKvfa8VpYkGfMeYmi3J0YxdUcv5IlN
K3wahiORQEOAdzAyoy2wGpnMGGk2pERwRDa9+bQbEbsURs3imUnty0hh+REFj35GmEdTP8DN4wOU
BeluR91la98N7FujB/7UFxBtgVvnB/3hYwePP2BQxl5u2S7nijO79BBq9BRx/Uv6QEg1Y/SlhC9l
WDab/r9AwkbZOWnglce8aiyBaEuZnGMIbnNbIx92PRjSnv23q93VH3rn44cvMg7Wfku9Fa1rvHIi
yK97QfAbwtUXVdteVKP3jHdjyGZPdyiBlNwUMaKEVTIZj0vKzOP+gHcIakfMYUPq3gu7ppImXx9/
fZCK44H3bvAyS6CZfg8volqyCUgZbzIP4tExWMvae712yQyX9yfG7Eb/zewtGy40qeOAbp2FA/Ch
M4HILvhuOOhfg+EkFtwmeH1yRrVVd1z9ITvo+hcPTI/FJgduoj56HChYpHz3GOmWtyFMIdlgxYTe
O4X7MLUXUt43MIAwDFBLZtY5C1KNdFHXmD09762XUCQzur04FY827HxdZ9+fsqekxwnKA8gxKCOd
eBJxCvlQgUBv2RxIUVFQ98QKuKA5aHq2wD7h33QQPIHZYffIYc//T1qcM39jjC/vSUt0nLIdLsl8
trlTIJTtAbXvWt8c9GUk0Rg3Eq9LGsx8R6euRT0Zym8qjSHonphFtTeu2Bk1+6PxFQnq8ra6J+SX
y8M0EfILO3p6FVFwgmyvIquAhBuVNB09pMrnGKt1y7ppyJH97f/89sifY8NO3k3N+Ogidq8J3cg4
Wfrz0sBBzMsWfP68nGbA90bbOOk0U9SxZB3A4P/ixIdhsPzy3O/n50hFlsHIo4wBiHN75XaTRsg2
al7ckxCOkVGRDFFvDoFY3CJC3+c792OYcM/j1T2NKf1P/jyL5cNbx5cOwRvfY4NLXuXVmqmHHvSr
x9iwezngSpNo0c7C36DEy+Qbfs1EoR5SOiBOxZBLtN6Ir21JL+PIgbruTQ7XkNhuMtKflIfPNuVV
7yoTf8dZplNke9HGBENB+t3aV7JYWde8YsWb5OhRw0RS2eAuBNcxVS5zwNldqkxkEROUpvuOqm//
INMO2VZSqiuYXwk05PzsjTlrW+jOiH6eK3b5gDoT7YSyKEe2+tn2PzIB83zpphO8xMQP7/MKLN9P
lvc6dHmVUo47XmXv08DNbyicma1sr3mHOjlIkD5mHgoP+KDmHDkLqIFtTfm9gigUhjjmfvvR3GSl
1syZQ7ppBE7QVIjg2UDdlop9f1H2xp2ZYkHfPxE4zHr489XGdGd/BmrDzHDYbqeNOO86QMc/w9t+
ImylNHKwvyHPKWAZ/R4qRRcbBgodA7KQ8un4GMBVVp6xCzwcg+IEGEjJOZepMn6E0Do/eMAuYfrq
oQo2nD25EXhVD1fZ+xINtH4/usbtAidccV3u92oWEcZkcJ1t4xMD9qsxvtFW477H4XOyGc28pXhV
cXQsXcbybmmD7nSRqzgrYFVyDryTUkw1nR5jq0kF1739o6muXrTX/YmV/Nme+ft423bQ2hvnUnMV
UlcLyjkOqQzaiZzODCmRG8wK27yZYY90Use59Fbi5362rfrHIAzYYK/HHci1L8C8L47VbRDjrosZ
DMi7W4swE4eEhN+cSQOv1djiT61hoF+g0Ww+MrKLQrrMOm7NM1AeGMeiZ2fhtXP6HuV8OG1aPJma
LhYuzKuiTeJuNBvAy3vnXwFO3QaCJEn762mbdJO3sVZ//R0wEtwI4kwZTOIB0t8Ji2wSJTdissq4
M/RmSLKZYxV/U9Cb4FAGfgkafWUPUfvZ7zRtXyFFdW5Z/CNYWBDjqIFTxkBhzWfeb3MT6/54ZSY4
2cDtCjdoZdWt/ky11PX1WxghrToG3EMKmTj880pyX+99uI8fqDTEyWWfaaVievX/P8yrNNKqudCn
4H623aS3ssKBk2Z8CQrwH3J2FZxHWkh0P5YBpDhQrJV6hdtqQxbAbiHNMjPvWdaDLMFCEqcuIpBk
s0IwcEDPwtKvL2TMxW0JhVQ87NuOKgPG5swMyUJ+Af8gkXL+UbFCUqawIzYglxvsOmH3pOKfeUfx
tEjmGgdDhUy4F0PR/iS40ms25GEd4sCh0sSMqTEnfRg23bxlwf6pL5HU0I0vC2fKUkzIZ7eoAg8V
FfxjvnNspDF72FMkApf8OlJ5fDObSrsoLJ4raCyPOcV/t7lbCStN+L/guxVGXxOOQW9qq3rdVV/G
edETXLSqndYxE/WRhn3uZEVQU6L1HgB5o3dmKc+svi2UKJaeLTMoyXTIygS2HemTEqmOidCcruTd
9LKAbrYit6xnaN58SroY8i2vp37/zREPZ4TkJ57V/ZO1Qs91s0xmMXp9q/UAUpGWJYCOYpitlOW8
ioIAumbxAcDoLJ1NFsm7BZb7Kxqz8SKvfuVPhl6eIjuu6JAQRfv30tkDgChlxMDxkU6N33aSbBjq
tdAJd9doyQhdrqIwtHcDRaNfCOKvKhTD+/nwlPnhdmIz+l7FcPKm8k5ZPpKJymsAP7kDJwE/98el
GxojWcRQTdoxqcY94nm/7g8+P8tWmBjh3GNaLP3yzlk+VQK2r1cDsv2QQvhlPVSZzmcOJYFtZUmf
EwnXL6maAQiqZzMgAI51YtD/DM9TKQvY4IAne6oz2i3kUCCEhAioy2NFieOgP9/T5YMhgiBEn22W
oPXH2SBo//zEHn8ZP6SJx9fC+2fNVKrYz/FJMfhq4zTF0dLwHrSU9t0Z2oOm82BrCklh5NR/5Srm
FkWDTfa0CdsSeKmVb+tl/WCK4Ph0CEUf0czhw+ZarPN0Nrut4YDRxAjhQZpR+6b5loSiefRCwBZM
82+lXCHjdFufoCn1nGCKxPTETw1erVqJHrhQKrrcjPteEasjDemOiWH2cCMshNWReBJs9Akmlitc
kUXNLujdbYWRK5fBKtH/JzSAjg3P7D7Av5pREEI8hUHruuRB7813+8jmSn0We8ic0SJZp0nMbleS
Ab+APch4dAJbdVKcly6oXIbfk+BGLWSErGYJCCB1YFD0RYIBvsUwI8X+hvY8019b5vULR5me5DYJ
+ZHqvyyKcRrhnRgKFD/82rO+mzwYnbjdYf6f4deVUpYfnGpo61GmNY3RqVdgSeAECMLllm8ZCHur
72ToCK23AtI7OxUhOny+Vk+aS8/g9ADiyPFCJnk7wWma3t5kiOjpApMEmue7yVoW444jNPuppJlS
K/SF5Rj4ZqELVLzrFeG2v+EPIvV7CSSVkeECoKKawdcnN0S3sUmDolg8yUJTnhIUSJS9QeECx2Ru
4vu674JAs3Cnh9NlF9U0KdChElK/bYEjDqParwVLpYsFuKM2jo0X4AeLY2BR8qsDWvO1cGmAWHXl
PnqHUoamn8e9A6qljFwirLQ8cdTnG+BGf3UOPECxB/d+x0tTDD718eYt/dj4/8vX/wfAoWWPuZ//
XOGBKDezZuDwM0yp6JKg4hLErMH0jKUp5kaKTAXqpBO1Rigzh2GutHDPT1WOK54ZBbtounSyOq87
e+lsGUzHerya9iae8Mv/2l2vqzDRWqjIkU1VG7ul378ovmsdIQb87FzfKQtTgYGKGwLdNG8PSuy3
bfxjogTL1bJVtKzvwDlSdXcfixIV8rRvPi/I0QeWIRl4SDghYR+H+vCkwl60Vn0YfQdlOMrgYoSU
3hC8qQgzwUhx6b6Q7KfhxUinNpGUGp0HX+vmO5rJ8IZdqCmgeCblLAxKBhhKEVsea/2MBhL80nEX
iMRZHWZZZQOr+yQDrV5jCV5vK+Pczu7vGKTsYLXOu1wqINfk7pgQOq6nt3o14i2VTT8MVlziOObj
wu5BMb65cVxFODS4aZe11XkcUArMztZh0glEvnBn6q690ScCp5GVFEV8yTigZhXbMdSjjt2FGNwl
BtNbOqUAnQeSWskWG9n8dbbdp5PWLnDtuWLHEHGnUpd5w6uzsRdfB6y17QjHs+uommLctOoTv8oG
qRupiAhtRziks2ChDc8CgGRo9LsLAcVTfWppdNkn3iJGWEynFoXVNnOgKbP0I309QYY5KJkD7gAV
rZLOU9oE+nY57y08DGpFo7aooa8K+DtL4rRvqyF5aWkNu2yOgDuhWh2KfbD6/IidWOk4coMi6lKL
/WVLb3OQwt3r+Uun8NC1ZmQCT0oDW65cHQgsnTCVrJywv69VWCxG/Vn/pSKzvC1YKWQ7k9TaKPh3
MaYrUKCow511mK4arYENd2QdJoCRn4kt+x97YZfBCHXIQIdVAQLkTKeD/3MwtHIYsihkd8lN0FQ6
GS6Riraqgu9ZaI+o1FdTW0vrKvjzaPf7xvIa9/ybxrifq/rzxCNBEfTvFHW9VPt0Ku3pGag4MZyb
Edj1SI6yk4qrWrjL8FgjghK5R2ipFd8a3adVQys/nsSWUSQfdqNCS75Khy4tN1KY6sDOuHwRWgHH
wglQpSUUHgiCI3loxNot3Afwpm00oL5G8LWiKRU/gfakpimzZ4kRDUZM09EGjIfCgTuzi/X/Py8X
4TwEVKb91+sv09ZrD47Pe2prpLL584z5G8sMzXbcchn23oAakQLiqe+uVIZci4En71VR2WvtxEtd
nZ2LOAJA/7zVove7HnF/NXHByGRApaQKHkyaFYdMh02XzTTFIs2+DbWe8ofas0o79xqARCx+aCYX
R01Mp7sRZ6NnnCCBTEGYJkVuUDmo+FWBrRDpZ5NSbSnNBNzJLNwaoXgG96GPSSt9I6dWrG7EjmkW
MVU6ThwuOrP2CSxGOnzvkS4LjuV9PVD/mHurmv3IH+0gh29Z3PMyRCMm/+NZ83Ple8HUmfwc1GFv
P80wLa5O/MavWkOSjFr/iY1Cja2VIKRiW/mX3MpoBQa/yOt9T6QbrblF7NCEecAeAIOLlihKpOUG
hIkMmPXRY+NYE37zQ60pldy4VLK5DBpRz2KrLEvV4QIJ3WMzy8iwF/ln4I1waURlgqtBIYJs+8Q2
ZNYJhWC+3MfJskFjyWRUxGQSnmeByaCf+flEUHU8pnbrO+T842vyfCwxMi2JhFASVSObji90tPFw
PdSsA3bu9DZMlgMWt3H3rxHZoFwUe6/zPwCF8gWLDlH12bfi0hcCkv8M2Wd+lLuRBHFn6AC3gGgV
aArMMi7x67R0iP9TZs2hUVbEJJOsbvgxOwukcAIQEHh0hAnEj1uJZ56fHc6KR/JQTbCBdx36gXS8
RC1n1BM+DfbTa0EWj5aogcd9DuaK3rNjdrvky10zcPuxKME/kw50GL5NvAbGr2gEq7nmc6xXei8m
oRe0Hv5ZBpK3h8xmrq1SEI/zTU7jNc5OVDLrCX7sURsgnxUebp0zO3iiegSJadeIGviR08LvUt9P
uDQertXfRjQfy4yAMqpkTUHjJUZzu2jFfK+4FdxqE9oNv62wWiYqr/kdOsk9HLmV5sNB+sYmR9ot
4pNQPSekfxJHlXtxYVjY63IGuH356EMebgHQYIXhUxYXpFV5t254TjlzwLJ5DIv6Ic9zul2/cOUI
2if5ZeJRII2O6/jAv+6U/be9RrSIfg7vYofiwgtJJenkh6ePrVhmuFtv7OpdVopKvvItC2NVMasz
EZKh0mzAXWfO8nPhCl5X7mlnqBlW9AUvbE81PF1AmlAV6zMxYCt3+u9IBmKhgU7FQE7RVyCMqJml
91x5dTfsVFgOV6kv4ds//fjEcyDdHIVn/lqPsy8xnCBGYxYJ7vk9sQHyhcJqpoGYNPjlOx0B+AJK
QrEWj1mBpM1Kapget2jf21dBFbAeKIDPT82VbeEeSnLep7PSP96GFvfW/lJ/UiqfnlPboGAt36P5
H/O2n4Gf8y6HUyfY6+e2nsQgkRGCuSJdr+pQ25/yx77KDf+M4qVliHdoO0hxaesKXEi401vQ+4N2
Mho/YZiUzMw0GYX57FAKUfZSDTTF1M/CS6q0Dxj7YXceNwHRjNJ8VLp4DrfLnkyMm1W4fSLw/Kdw
wuOkhm7jMHGJyrmng2sYvolqf2M0jRTEX96Z+bEUp0BJRp4TS6TaS0nPevl65nXG7EHi/U0UkFLk
aQQZ4rlRrFNdV2+cUqixvLq3XJhdSZxws9X6n428cPS1VNN5ybDtckikWinFqkOt1vkUREDDYz4w
o7an/mvabSiza4cTvNGEN61Yfx9hqEncmM9OLd6gsKHS2zNesPofzbH4uP2auVE5yQYqYCJNb90b
PoZnWHXf+40t/icPJe6xzp+ArUyAFY3zYvB5ufMcUCZ3qTi50eTbbUDP1GKbn62U9denCLyqaQOv
YLra4m+XgGD8bTkLhrqRNWc0FkdOOfgkWt9uXO0k3ZwgTzvwGFdA/JvmLfI+W7xIukIzcVlwoxPM
LGr6alfXo5ohDaaqVRua/18SLcjmwccflT9Xd7nt4bZHVFLiClsbZUZmttYFRAaYXj7u4YiW0+Vx
Lkr6ZY1g2vg/wWcDPV5KW2MZ92xIFATzlAxrsfNOw6vMennmpbljDrLYibF6B1c4Th7Km6YV39xl
XcM3rsWt2pjwapQYVWr/vBVBvQ6zfTLVxrjOs32tel3NS2RBxjEpR8tPcXZtQQGv1+iqU0ZDaWQL
WGMjadB5YglCwvJpZW4SsdbPt+smLnLw7Jg58GAC88bOchdcOaxlNlvZ6mGBv8nMuoQW4kD5P4ZP
fHDODSvGItLD6MTWe5HzC5arcLAqhD/kIOHtnhuQ8PT6qncczHyQBK+RctPI3al0EmT84LSKHi7f
UWlStegDdyCvR2VYpSM+FdLqNLp2tpbvfCJjzz6cjkLYpmRnbfSvmJUI+D1MinOdxPg7dVngqkye
0mq4Wddjwma6NuwQUHUTw8pSadwpcBS50jrTYwlszQ2jnzBCVaJhiOvd6ILgvazEXfor+QxK7pKS
x0HEvK1AXLXsYqRFZdNWCoPF2WE8GeGlyMrcfToy+RlYfASD3Bc7JgYl1TR3oU+9QvhJb//4Bhp7
aB1MAUrfv5trzYM/NGXUW1JDR37sTw8hbPysreAbb3oGWX8EK0WR8TKvcanGOYpcNpeal0r4cxRG
UJFUaIBBwZk9AFpY6ZcZy+ZXd9F5i6N9XE7mMWxDmdbuA3NVMHy/UdjjExwvXPT0N2Z91GBXWI9e
sJTxUTIsMMo4LaHWd/1tskI6c0WvZ9XpzjRcPTx0erEMfaGoSHsbX+YnLG9viH6zUD4iacLDPyh6
IgGy9KtcGLT9ivooonqEp/Jljb5xOG9zNWtFKfiZ+AdEWEleuB28mnPx1iNecCbxLWGU91iZoyAA
orXck/Ia8ZrCfT0OvcLdUXw2DTDFpzV5hlBkgRnZOPW5gucz538aUPUPPIumMi6nU80+QUwQUDx5
AH8ZZdWbNCNAlX20zp5rnkFCleAc0BdfybzXgR2OXeMfktYETWyOydeWpT9XCCEmIvWL+tPyKJjp
TuTxDAns0nSv0AAKxoW4B4ZRCAS8MxDVpRc9yQDnL1KQciglYy0n2PJsp2++wlhNt0lKl9+1sfOX
6Ih6fcSkHdQKrI8mDCaYJZDX8Q5xJhribDxYYuPTi1pnmX/w6RW3ZrftnxlZJX1p1tKPtrlmUzlg
vMnuUoAelvNllvPtUA9zsb7SGjgf3agVf4jmhlKd3Lai4YuHty9GIOu8peWLedB5/yWjrH+YKIpc
Y4SXrR0vru6o6fL3F4+OjYe3SqP+CZ0ri969P3VGBmxeWripQtNT3VkCStkcB1mHWe1tHVTanpaD
Np4cnJ354FA0EEqGPjyA1az/miZagqZnd85rBeha8EE2iQ/gOI1ybax3ZLyo6zzcQjnSZD4LxyZO
zPNcWKtZC+10pI1hJtrnYTK69OBqkI9Gn2W6e3PRwgL+eOPb44KRWopPclMKGIE09HoHt06Kwf4U
ucRUU2SNkxLxBj7Qu3C7KcCFmsB1/+fFF3eT9JyWAtvOd5nCxYFvAx7xrnoGApeVZXGwNTJmbUNe
AJkh967QNyE1JD8GFPIihR/60ISK/+t0E2emnknTk6T4RCSYR1Ogl2mDQ9U0nQ/PTOGmbvU0aMsA
ybjxk2s+xKltmVNMVxEq972udPg/r3wZnL0EhKk+omwF5Yg8OcPjbfL51ckG5E+bI+08njFfy9hK
KTPKAd1wEHSuLJxENxZfbBlWwyoNUZDBYmL8ZQp8W8rFafNvyKfjeSVOZeetPQyhJKsL1NANlpgY
qR3m9URCJEISpLAvv0nGB9yDK7cIpfjQos5JpT709vzIjshYIflMmJSAjxXAxwkjYP33nWj5p15s
YQjifHBPGbfHFhxZjUz2Lyk6HcIodegKqi9WQdXksV4wTS4r9us8APUgw4+NjBnH58jdA+0nOlpw
7W9aOFenjm8uTlauNctFFn0bySL2XC9x48yx4+rnAnMUlhILtrW70QLGFwgt067DhcVH0L/H4A6S
+hwDfu0nP5Xns8eNSlwBztf+R0saA0IEV2A95sVYptk7sqSvfc0JwvbStRSiVjcYRcDxGG5iQ94X
qYSTfWiTYLCHEK/bA66b++1R4r6iUJKBevstuBY4u+zhuY8yuEwhH/SnIr8V5P7n13vsxtAZnNh1
EweJW4kyFQiFv5RChoSazX8ubWCABWq7nyEmlKcDN8Iu4kBSt8FuhhBDXDMK8Vz79KjAM4M8KvXw
Q7XRNg7Wnih2bs2v0XXGEX7ZyIBz/jDffRpMf58isFC4kk9TQ5KqYq7cBrg0WyefzyeRJlASl/Oe
8h7i4bQF3TqWo0npb5EptOUEhVdl7VotT+Mj3h7ngSWVv6QwNzJTv/F+RgpvHYZCItdJLE8yw1wT
FbQd77o1qF1kJ7QfYo5p7UZzpx0eWpKZi/LOQO8/AS851A40WvLq3qjuxh+VP2iPvcCl7Nc3xufz
sWk6DFUp5Gwn8niWyddWB9yoQAaIxiv7GWdRFGh2oYduln16Q66hRbfnJFbnbjuTg7qDMmnDMD5r
IVOclSmDq9lmntThNTlQpY7C9xbCGUL6Daox+2h8gFkCG2ymWxCFxDg6vf4/FtYSdto1TFSTFW5U
vcZ6KfBAVbKBVvJDgyvAxUL6mbAPMnmqR18WBmVpmmcYuAzQ/A8L+NXYNtzd8yeVGokuck5cHXKW
R1Yti18B4IkjHqIIlxhdXjkhJY0LyvIt4v8NY/SsLRN2tpMhiANrtDapDBugKowQfrC4CQgtseyL
z9FFntGODfi08j80RCtpeSIBaa5CL8dV6Gsna1XByG3JFsjnCsQJhuWt1GUMqCzN3dMd8LDsoPHT
XgVQVr8p/OOu4Ahp4GFWwtzi/uiMZhz0gQIX31ptMpzWtMhgpF+ArjnWrHN3DIr5rjGQUPbe7iVn
ryb+NN3A/gTvBdzugANR5S/3z0rJ2tF0f4EH1tVZyQzRGcocnicWCgh19713DKdJHVbsqWv/qbOw
oM+IGOUTfn+rhBLWw3KBDFM+WUWA3XG40fjrDbx0TmxWjHS6Kz6F/x4h/nT28cg+xJDWUsmAt8NH
l3hnSGmAqF8cLylOjVs23X+6BYEY5DsERmkt7QDeJqpZNMARjNAAwZnc+CLn0hwjwylx/Pdd7zXm
SPBxFRhTwG8x0jsTDX6C9YGRelOXwQT9u1SYLGuwiwfHPujqNwOEoNACQrrL91CVYCoaKphN3wuJ
mlpiGBbTAT+waDfKpx+JbgBzXEVHhmPKW8lpTFht83lFvtwESpQmri8d0mmK5TSLW5tkLHaJEWi8
qsmZzrsqBBGdjtthATeLLXu28NptLLcJENCTzpQ58AUt/ansOmtHErKb/8SKuSKXYIu/+HFQYSdd
KxnaUYNv0CU5P/ZjwgkKUOLr67i4YEn1d0wQne+cJ2FVe5vPBGk1xXSPz6nWxfujjDo+XJ94EECY
x52e5vyAXJTn34NrmZw8hVs1FfVJtmTwfwC9eKdIT0wU8FfbjCu0y64H27JpbJuPsPWIkpbCXfOv
aNFUN4iMre3yPq+xqvJSP3uhcLBcRv30c4TddPSGX16cH3qkXZHg5ia2UHz8H3XER7x+0QAchbJB
Htd2ZPyQ28FSA0RwqTP7r0lvIHiGKF1b04b+92PAlE1tkcW/bO1PUIYvfYJkm7RD2+Wg7VWZttn0
X4vhWMftOIUKMtkqudZ8ICDA0mCSCr7Se4u9G4rNgsT5zCZGDC+KFM9dsmrwO0qSuUf+nA6kYURH
+62rQHGZsF0LPzvfQBsKPU1iXtoEboHwhVeQ8cqtEqXOiYS12OTcpXiCRxo8Gz0BIqKLo58ASZh+
9lw2D8IG07taUMqWsf2omHbO7SuAWEsZoPQQwXCGbuSV/cCBTabyhBDz4+Nx9q56dXbNWwnqX7qC
LuPPH+xD5ran0i9HR6aMmL53EtNdot2zn5P54cWaVGd3Mqvfx2Sh0A0SHAA+1/Msb2OaZtBzmw1c
hMqrOyBiOmEgAcFfnUY4tZVDCFcArc1XloHQ+Rn5a6Jqgc0z25GLUpooHsKjrBrMjuTol5H+mj9c
ruQcaO3INUMBPbotM0Ux7iaUPONafC60dz3JA2IJFPuQMmEIGj0WpDRB6ykd5d2C3NnJrqOMojwo
10hy0rFT0/g/VIPbHZbBXqV7rgL8nRWICsTaA8+57Qnugl5UH9Vrv449pnEs4+5aoem9FH8DoUum
HYVA67AVzWjIEPSBBm0IepzS38z5GI4a+ONs5Qc/QwkK6YVvtm4dZO/9EkmUXl7gyOaEap5XFOQX
/8yg3rO5OgAVRiWwbTx/ApNa0tHTko0TcjBiCJw2k/62+l3+zOPr/5oJSOy7fDsWNzWcYDPsAnCe
K389V7f95brloPdtPznNuwyszScf/3c1SdDVrWYYyIqTT8wRtuw0LJz++fOy735Yehgy9RkDGWII
2vlQTTgr+45F/VxInzjTC0b6uO+PsFph3ZHo2hpIVeSI2PCHrguiwhZ1wYV8ixJ/GtEr8YugiFu9
l1VQbxJcFr+LG+Cv73ICmCnAGY0q9HDW7eUjZq30iMm17gO6Ho56HbXjrc0JlXQ1Y3A+qfY2pZu7
xI0f6/KnwDxSu8Ivk5NpPQqNn9WX/uQaAEY08kWFpEhx8TPIobDhGEsFzD7LFbdRzldHQVLlj2XR
0sPRtmC/cAx1tMAXlHONmIPFS0eOZxqzqYU85fx32ecoMITCx6DP9GP8GOR7op8gUYhrmPEju8zr
MGHCNY9ifRZrJAINWGKeA12LgSSDbpNWAFuqk9YdbF2yXdZD3+BEm+iiKtbJteA10VtUkD4AUGbh
ag2eY9d9ktWLLnqc8Lj7Uqx8jgSWIxBRVXl86dhUvjG0NZSrdbpXnriU6kVUZpW99LG6byYthztL
p9ALTwLC3TYFq52v9ihESl4Az4PWORoBLSEO3up/Ied4PxduXduxdLeMpd0xp3+cz/EfZ/Y2KAFi
Ddyk+WIyhfMZlVyyVLsAkeZoricJNPYCc5Vxi1PTok4rHAt/ERcdmMgwaqpiD7m7whGhMce1LUqy
Yv+3gxlm+I74HKQnbh2mp4PJE4CiXkUECLAiBLWZE9BoH+GmCNH4ZdfCGDjzMItWtqKSI63uVA86
O4HZiu/A7fmWzOfK1dXXsig8xdN3rpj4EgaSfEHOqnzUQFWtM0VRKx9J+64jiZDTt1/5Dxiqco+b
T5mqfD0IJ1ETrrTGEuFJnqlFo9v7kQmsugf8w1Q7XX16d2lqUtFNQcolAYsCLYmPxO4lxWZdf9Zg
8K9G43TvgECMTj24gq8zWcaCRZQr/dcKVnAlXGqHpbwdX8dbjv9iVUPu4GNhD/TbWAAA6YQvpu+M
CHwysZwOwpQtJRqNYr8T5uiJ+D4G/LQcIdVNgQBOx2fSm0Lcc4/v3U4+BF6BIgmp7cG45ypAZfc2
04xSD/CP2iSeMiQLwet4lFywRnmtO3dNCsa/eT2M9bJmARttJ/jYN3/qFPxkpwGKZizGUcRmFERD
KGHfA1C22JIMDwWtRNQz88hangvc6XbqoVs3tFfR7IbKiYD9e1Yd6iFRMTP1SrSgMucV+21FaZtu
oapTOp9KVK862W2OfUGI8dRoL94ZRArb651t4LSl8mplVhI7gMJ/miJbxU13FYWBpyqew7Ool61O
vDuNqeWA70jhecSy8UoUXLLzrV3CScGa4XJD0ak6u1uvpPK1CflZavMKdBN0n59aUV47UOh+DBtq
w60igT4NFh38CbGkgnV5GE0P4UVPh1e7wgJv5zsWimY5UyhMwq53ISC3uvJ6PjRj0mJat/409lRK
HRkfN5sTr/3Qn4u+euggmWntQ4feKkS+WzdLNMyUg7jTvSn8cZljd1OXOEOrK2NwjbX6J8mMcqBj
C+wX0bv4EETjr9tOrHujpltDYp7y2YvzMlpwAXaRjneMnDu8w0R/wMBq9WGyAychM1hgGTda9ijG
NI6gPwLk1yKui4sZ6tJpqU5fw6K7aFvgRZRKfA6gVXvRGeYxgaOB6VdDR+mdH6p2w/sKfytYSfTm
p2ML1Fuq+XJDnm1+P60Hk2n+/w+D+fbBodgmNnCt9bq72wamCnDoIgSsNUgrtaoMUeNhS+NpFOyo
CtsamQIsPjFTWI0Bu0O1uwCMUfv/WVUGPv2MVMiGpUrmq0KLunP4HKcul8/xi3EkGsJDljVLuNum
7gl85OwO2VGkMLjE8kXzdizSm3vWiQIKB2jDspNrOJCIZixGSyzFwB6UGCYAZKIuon4d5DC0ohmE
rLdNSXxsYaIQqV2G5z6JINj7clbmehjT2YCh3L/TX5duE9BbCtFQjlwNlR39hPY1ovFmvBUfhosC
Jt1HRYFxadUiSkQK6huL90JFIGAScvEElIAX4qAVg6rMo86QTlJgNSkEhit56XCpqmnH+WeUG5Qj
15YAXHBc5i4cQH29sgOVsScJcvW/YKarFdYn9OgCyns2+FFUshCcH0xKYoD2dn0gYmYTmUMhAXRY
njHx9vN5R8MenFissPbeaRfZAM9dJ3aIlYJ5V3HzSPabSkS157/KPFaDV5XpsCxYSHOQ2tItNcFY
HZ2V2VZ0kDgIMno/VHYxGXEMxTs2e0YlwzBnyWNiWb2F1c15XyZzKjOKXzWqU3vE1pmNtGsN2loP
ZIS+jFz/WJn4sb6eIzTJ+/oDYg9lDKQ+WIicCafV8rr7KsCq5pqVVBZqgdcGWXbP+Wzt2xV4TlJR
5t1C9Nt9D5GM6PLgbqQT3wUAa5YYWVXdMoSaucRuefo2D2AFk3+cyqQklHujLUpy9CttpyWXWlrG
UZatMGRC6gzAJkjwCZ26XBSqjQdytu/dyaOiEhXsEzp9e3T+HLlneX1Z7QYgtXZQ9dT2r2Or/z+A
y1TCBKdl4svnJMu0ETNz2FORza1nQ902MEQdZJlmuRpG99PlLFIg4cz2oY8yjByx5gMvTb4E8Apy
3OZ2QHgKjiEwn3JRZbcyoJ7mRr/TDiJRXPqsvH7dL8Aoy+SaUmceyz69y+xP64Uz27O4rogApGB4
YKmK0U8fpwM+w1qAq5Gm4v5b8zW7YFhgLXNJOv5Q99CbUG1Ic+5A9qkRSvadjMC+moNTLz4wVvLX
QGdKojN7SEsYAFX5ewhYMSIbZ8jINt09X7deg8I5pa3Bhd7aNtiZOVuxNr1poK6IuPCA+wuytMpN
Y7yYegApDxkO3DuU4b4IvKQRegIgkWifZJU22KdB0Jkrhlkn1YEMwMWG1zXDhrrTATlNAoJMQEwu
Ovyx/XOPf7w+vnjqBfXoBwwdL7azJpdSuvTXLXU2UJuZSIxGFmfCdM4kV1JdQLD0U41lGNrLoz8p
MYW0Q4nZJWXv9WTNsHEHJ9N1g4M/lHTXXgrjioB0/5323CPuhA7QyXtNO85XGN564hD8issGV2/r
a8muNU5V/U0OAvbsgQ1dznAmc1LxAP8uVE0cjzs4OWnnMlHopXcB0/HKToUd2Gi2hlDxmNqYkKbP
JpJXJrQeEE2nkLhd996HaFskMT7wimWalShHjWJVhOmjWqFY5Ph4tlP/xX5IeSxBTeXGIePwccHZ
wm1be8vksVpY9v8VJSpdh/tMhL3w8ipXMcoj6fmW7Y/g4lVArxjSPFHO/GfhDiIoE/eTAIBIBRaY
B4Ch7h73N9JRz/stOOt2pnuciIwuHg6HmIVYvQEiaLPxHLaoSBBBvfDTqEWBP8B3L5A45xq0dlS/
2eyt09zdOGgoYZI5y3BhHebX/pSsOwAHxrqDDCyt26rqJbY0Cc/vT8OjOA4QQ/J4OB+rl3o1w9hr
jbVshiN7bYER41q65VtMTw3yvco23VTnDOY6b2y9AtSz0eSjkRMR9xl11sVgVZWnIRiFeBjQ5iLI
3daV3bz5+lR9AhIWto0VongyCPmfzV5VwNxpObHz6X5FwMAUnDgVkQFf0Irmiz2zArLYsILn9UE3
JhhM5q38ibsDmGOWX7x9MVeu6D9Jm3ESwv9LOhD3Cp8jR4rpG2uGJC29MLG8Um00rVNbyvJTPYs9
56kw1ymP6juL4VqsE7qqYtc9EfffD13GNuAylfvVzhtVyuCgfLUzfb3Xm6YhuHHrFIhPNE2l40uK
n+jZtgCi5+XbFH0L+bU1CD3siNZk8+3WDIJFqmbY5qD800EJG7NLvocQ2f6HKDjyN+RvcUFVhM9d
VT8xvrrxNAcpUqUoHZ0aL1pIiqgoy1YHBN03WOQ1DiFx6jA/UdINJjTDMnSooKoT/Cbji/Ua8ecs
qbe4+a5ipMudIks/9FTEXJXqyBWdfFXd6ThXjCOmjPMy2wLSkJhcNOCLAnjOjG9bb16mQSoKPimh
e2zLrPvNq7TNqIUH+QwxS1d82Bw7IAm4a4IQ7NZYixChSE90e74Prpq8IRyM+mIrnn1oWpIpOfcV
G01xRpcvCEwwAqc0Bs7SHGJMKG8JvLaD9mmU6Uh4++1JUrLFsrnNHe+VV9K4cl9mZHmbnd8oroa8
VQpLVwb7WogbC3D5PRdcY9bSpOoGOJoEgAh9Q3ebPlKxXFjK1HJXQ2erQLWLO04Le1DuLpy/w5kW
RzGn8vwiz/AXLrwb6TNz0lLbqrwbfjEBz33/xPk8805E6bfhsF28ebH7z/hRw5jZvrKgdGBWxNlZ
Fid/qEbSX+vHHATx1w1aYIk7UH2dRI1W4YV/i4dXmv2+TRx+mK20/A99yfB1tAoNwVTc3blDiEPO
0zlK9YR0q18t2aoopylTqthG1qNS72NIHxEWNVZMH+xdVKyz5TkSXjar+SaLknJXewu57bkg4BkM
qcY+TolBCNj5SfrMJq/5KMCy/QmgHmRk43NUI82bX7kBj2ZtmoNVMKjK6fe5H1hJuZpTE3vCiXU2
GoxmbVgose1n3Q9MS/ipR2ZjMNjh+noN8OSkVcEsqK/D3BZDIXkCX9TWWzNQenRSdfX/1gux/1Np
fX/wSv/bIhBPusX6sZhlysBrBHb2OrDdM+0tDkMyjShQ310htesx57YKkUCMtY+6e+NI8mEqQz1M
JgnXZjFUYNgoommukDtLWZiaNFmc2g6wG/TgSxeHsO7uJYWjhGZGebncY8+im9m/Ci7DjE/Ckn96
AcIb/wwDa6ZJN2QU4sRt2yBQN2D4lPTLJuHuml30h3nBkbtgD8My0NtgJPOnQhDfLu9TobeXvVdL
Sg2HCv+cWcIiicLA93uPqxEa3vIbYwJ2Z5j/Vw8Ux7ClXXPnM7c5mfj02Qf84m5DJp1qklc+gAnM
lgJ7lUmzZBgsaTse7nZqrW+5ufuMBDaCcznV6eciaE6e54PZp4VhpG4qr3qz0AtGGjDQhJnmri4w
iLW7vEYr1p1ielNjYghDlUNqtLZv+or7h4lqzuYv3kpC0AFKVAmDMAlbtGYnKX/Pzz7rpDhpHFJ7
6/Cv38xzqdwifpginw4Wz2E0w6YHWQgcxTt7HifyMlfaUvZdxFLM5Y3C/A1JHxm48Cl1B7vnFB6i
J1U91iBeEQJ0zJOig8OAYNh/3IrO1VG4QJY9aqHDy0zT09NA6hNSqnqp25XoEAwdwNPjoh6YAvy+
7hK0oJJijtguhiR+tpFGBL0F1TSpBBlGw9VmNppqFs2iJlIW52XSxUTszCWoeZsi+USsGc609fsl
IiCy5LLw1yuemT544SP6W0cCPtWAaxOTHVmBHZk4PuVL1tESFlmII4GNZf1l/QuAK1Dn7L/JV0kj
Rk9XBZVFlX8+Wnfom79p5XJlltqcUJw7PZOA+UfeBqmPD2gcQAxmBpCKcIGo/WpkQm3z+Rx7cXQO
ctsIBUH2HX0GVP81gMFkTR/A7+4qNAPJljKeAgjww82/DJ5Nk9thRwI1WxOfK5w3ls9AedSf7kP+
LNQBE8C6eKyCz0K9YdxAHxKYgRhieGeV64aBTBqJRo+J1apbpAOtgxnHg4PSKGkP6CjSPYK3mQ3k
GVBxyRdVZKj4otsiltPKfdY+r+zGW8OtD0Zup0rm6FlQy5BW26cCCM7Vgf58GNhGH/mc7k9SqwsQ
OtLs49L5uaRon1f88Zuk5oQQWEIgo3nCL/KhwRkWcNFvFAIiqHCojOK+B6yCC1RO9d/X6KKObDre
mE02mz6CogdomNl25OGCYcEXAN5mSK3fjkhJrRA3cjr5Tq31EA7oTF92I1mu+TteF5In6jTaXyOb
60DSoeer0BcOpJM2txET8ox0HEcsTpM8PtPSngWcay7AzhXAon1D9N2tma6BqpbHZCd/5jS2Xwpb
NGeBX35XHA9VN0ZnnY3NnOIZuELKbI7DpJ4cx7ZjUVfsO0YJhZ+cWDHw6ruMtI4gZcLIRc+Eb4n5
WcGb0Xg2+N11yCcih1UCQ/QD7O99BkW6se5D8eqFWKQrug7EjJTFSrlVRfyx4oMLaVcgaZqoVUmb
OT8/XEBYR9Yt5iD+8Zm//Q28HfYofqEtIlB1C2ylAvUL0Nf022+NCAkI4BXWOnrNxDlGXpXHLRdw
ejFq/GQ5fODvCscKBs1wZSDCEYGhNxTALnVEcb1ZhHbUjzfSg521fHdDOStCsX+oR7imWSRpued6
jm3I5Z2PGwZSHHrUNDajogzIhmzxgtmpVT58niltsm2PIZTiZ460S20i+h9F5g72MSk5ayPNJX3A
PZ5YOIcgqlzbTZNsQRlEipyKeEaww2ionyLoDoHomZ+gHFHYw7GXwTDLVmhNokUvvYnrDfSLbxBr
VT0c8NcBkK0B7ho8B2OOSBihZxwCkXMg11i9z5Drag0ICh10O3Ss0C/rAtXkd6KwSR28abgq6OR8
2kcqH41bz9MqsNOVbdesVE14cAPOsJx5JI/CpOxt6UYEP3Ehy68nTsVQunhBjbNPAJkxr2xEpwQD
bIdbad0iLgh9xlbw20SAWxKV0RDad0IMojCIuQCvBTwO+mApFeCWXYfEYyK1fYGJ+rZRHR+2ksQq
MZMD5Lc/ovIsWLJL+AYCYhm6Tkp52STgshtgAbyWpYkp3q8xI9Hr5bndfucMIVbH8cr62jfiEfwy
ju/jeFTAh1C5mfAAef2csYQNJqBbZ/Af2KCH4ErYOXm8roNZ+CotwjvwguQWTc9YpPvjovlmY2Gc
tnEcl6Ye7iCnVSLlfEocXXq2weqMWFAF/bL0tsb/dV1lbh6Df0vuFG0LEkLRQESiP1uUisTdT+KX
Vhvc4zUV/Qjk9IVVs9aN0ELYprJFYJ3gHhlEgLbc8sLvtK+czadxAgwRvkyffxhukRrc5QRrDXQY
v2YrLdzAEgO7CfsUV6QRfRAykpq9y0T1jQxrYbQs4H1DtTceoN1xRQ8LV8XbtUSL7jiskMtkbE14
oOMjN+rBlz79UHDShs2dNq+xKXhOKvv3+ZCvwOjZjf5N9e5adHMBMFauLacBq+rfks4Wx445EuD/
j7hazf3PUiEnh8Y868+BB81abtfz6RI7xiFZE4REtXHNuC7svSAiOFJVuxmPfwk+plOBO1tzsjca
ufk5q4L936B7XBhReXAZCOMW6kyMJc6soU8F+RORiyWs2eonUSsL5m9YfTrClGImEy1lo+nMacxN
hjPYXOSM44Fe08taqdXCTgnOMkmoWHuVSNkrzBzMjf/ogmflsD/EUdulgk/E67eG06PhpMufBqIi
P3K07Fr0cwgTGgQj+hz1MrGvaQO6Bhkyg/x+NfuqmV4s+eFtZQ4DSGeu66oGt7OxuzqPrX7GAyb+
Jx4hCBeqreYgFZPMR72+gUUadKntiDy8Yz0ntNngjzPIUcOLUN6vmyEYuaw04/nSvXWB8QUbaWN0
ER3g4fVTUB/+sJToeEG0YoiAVoblykidJe9WBasfA+9DYG0MTQJXur3jnlcVbnZqgkvLohRGYtoT
1Ouw+ZyqZG8MK8n3+tAQEwaXua1KoHmg+YaKncYDBZFwBOWjJRwD9i21ICgj2dxoSvZSYfrDSGlO
t7A6zKIsGWCAF7VoWBvrs2iq+OkixC3d8mK1XWGH4gyaXrjV2c7X5BrrXEapHH5Js+m3hq8UfqMG
0UtXg2ztvtS1SN78TANB9Dk5sNMpQDTN3/kyxJWcEqC2W6JYSVA3JRdVzkgNk3uhNmuLggWm9R2Y
1teCsiMCagGSSz/NnZ2ze1es+VT/OWnOK9b/nKxtEvaa8xxcp9tL3bjaCMxAHgfzFdT03gg/28sr
2/S6dMh2HiI/k0KPx85SFWfrfSMaHaFvlCFzB/XHKmVVmFjHx5W1kvYksoaKMYV38zoRzi/v8XcM
+UASzGz2YN9hCJoFakql3vd9yIl+4KKhhZ5oSOz1vRIFBs+rzjEJrPir7IcmbOYxa9SLcwjEAZl2
/1qqu+p/9PI5qRB5XymVI5A3qC7YK0T9jtPn76auIi4GK9C41rQiVKcR0WiDXTsUOg7qY7dzbk6r
vqsXOWwz0W0zNsqWGJR8O80m4H6Wg96cYmq8KsLjIXYwbXoyyX13V5ZG37IKTR2P2t/gcnti8WvB
2u92qG/x6xBOmBLPlLsIGRkC6GGYyTwLzZ292D1WJpBvdlxAxX37KFU+moD48gr7a2go7vuN4Qu1
t8+mptMvd3kl/EU11TXiF48D/N3uow9U5HFQFtGlUZNOHZXnse6YwroPLS4q5YxN+5JUfKZCn0d9
9npFZUMW8eapUwOTDl+trK3X57yxLeaSD8K875+NUJULAV0hkmpzYlZbhn60TKqfIWb/C78VK+Le
3ojumdImoeYcbzwRGx3xg9US5z0peMS8WGWpaAmkYNTq+x76/28NPqcoL/l4pmu1PuPh+9OXxP56
zUzbGAZhdaIMWrv8Wqb8UUPnqqPkgS5znmWkPCXscykFJ68qLoCkQPfW9W2q/ddeDslGu3uY72jE
eijvgbNG5Zrp7rbAFGotrf3It9ldmhlp3bDMi5/x1xpyorNOAFVdvj96UF/BCE4mLVA5ZIGqTF94
RkYsZqXujVOwrZwOgtlof5JhAjEUV/GjNc6EYTkjKj70wf1QNJCYxclwnLw93SQ6tcS3fCTgwfk1
1cIu/7axDpOrfOCmPSWFWFdFos/xn1hUs8Jz8k3SNufyxLpiyW/AVXAbV8HoFrrf+vYCPG3kqyAv
iPMoz+1nbYLQ5f5Y23/zBrs78xiLJAR1Y31AXmXQbnkVcyGT7Zcnd0h5LePdFbFPHiGNYW6+PSpM
oB8mq0pXRAafgSc1uo+zF7zk2DtMpHZtIhX1vLh/Xs5JLPotx3efJzKj+s+AmRUNouDUF8D5pQjB
NmAwlgCRGeHLj8KPvIhciO/A7GdXE5VZI68yEo80/l6aUTQgnGjxufhVRRt72qdwCV9beMQ1NRdD
WN0UgElr1Gz21own35yGrYiogbWQ+UeL+wqof+77g6iXbH5nlLPlKcY3KaXdA5+Gr6BzQEC3Nnv7
5UzEVBX/E2juRVwdTIqqd7w+x5tGHKDgybqaw3ceiwijqcCSfTbM2JlFnElzSVzt/ASoyBu0YklD
urEjQlKwrBK5QASpZHLuix1JP6eWk44zOD5AJQd9LxIq2UAE9V0z70CzI6k11MNOfmqnQAG5LZO5
sG+XH5yHjKEfOpT8FTEjEmyaOc0zF0rf7USXoxLNrHtkoBGfIxzcngcbMPaFw6mq/nssMZavBi7d
fwcNfP76nvBsarr6nMA4oNKKmjP/FjkWmy3680CvtBHgXHFBn9kdlKlqehw3QulpBww1JQS0VFFZ
OkKWgZEXFpyRZFgjTwyYCjA7RQ60PmFioi623GftBJbZTzX+atsksfmJjFnAo/wA0k2rMTCBPehS
VwrNayZbC6E0vpnbUnyxg4ToZh6jCSQqpZSA/cIcez7QYCeQGu5eeUbC3UO4Bh6eOmr/17uqqPnS
x/D5iqyuI7DcuK8VZR/znYhmmyoo4mI2p+/4fRhJKBjVSXcmGYI7nndIBcsY3iIpqQGqbMo8YAX3
UFiX/PfFMBHj3G2yFDoTuYhOXE6mXg4hepaCeCXWUNi3JAZm2lR8pevE8reY7J2oi4hXmT24rTF0
3VJORe19DsZpHW6SAcpLB+qO7HuqzVFRMbd9In47Zf43mvL8Ge78eKBHke9pK6Ug8DAopr1wkW9/
WBw7xsk1DggqIbfA/p2QnomXsEmk40/5RRJUFR4r6UXfAqj81XRZjkGHwrZMsNxxDgnEVtGKn/2O
VW/+UhS8C7MCBf/FU+JNNZzZcYhvvOf2LW5XYOeIhuNpy/ITzjX4/yv0ckaEWciprtqW218SIIJK
Pzb4P4EcMGdPvefXMDzduI3jtXn41BENE2oznSpCmWkHWXiUa5vFcDif0pH8Jt/KPWfcmQyRVUiH
jkxYG93phYO98iBxzlXnwK+ZhoEWg8mROG7Knd5cwyZ2tQzQq6V0iIkGEmQf2eOvE7n1Z6iDzizm
1C/xOCtWIJaNbU0bbfa47u31dBEgfwDCnvtDC6hIUbaVkgWPTrS6ZCAfDHKm5qCdotpl9v/Rcjfn
tz1iotz1863eckBpesgr4oFwlG+BpTe5/1jabCSNGXTyfsCyVdGSFxGvYmq38E3WgzjISbZ1y3Hu
qVR0pWOLNHJnXbmnP4giZ+PUt0QsJtVE6wrbTrowAE48pUPTfahFxYtWcnqCVRtsl9/AXiMWW2Wr
nYD6tdqGNDBYgqHLPQi0jZtBjEsBm1afl8fFSakf8IMAfEcSuWr5b3hclsmAHbsxZhM+JP9IRfUc
TIzLH1zBvMrl2m01ugkhnYN9qG7BGxn04EDKPs3xuS0UdScYm4KHjlfYlBTq5WTrCLJXTnJrUg+Q
qL+1JyR8TO8mypTdl1frh3HAKZPR5gCKGheP3zgeWnE6uv3Trtdsg0vluxo3IOl8rdhi9rc6c476
EmCAA46mc0zpRBBcqqqOF57Aq94XEEla7bUOWm/+ES6QlEtUVecfPLE6yr9WGQR9itt0JKvzj84S
rNtho9T8InbzXzv54Omv/2KHmIhcC0a2ad/52B4CmlVlHaW+3aRooAabjpk0+QgKvrR3dyCn8zm7
hOEmS7Z0UAe/4NNKq+b9+DF4qeFDXSRRW1DTcfJupOc3VafoJHBUS8ct4tzuye58vlv/hWmBMgzE
jgTIsSCInF7SDINrkrkYYFiYodaNCbypIEbM2e77GzPcA9MAs2QIB6o9SUJjoHm9SPcJi5a+UsCb
bi41JWl96zC0AHlL+N+Cz0o/tU1ATRJyv+VfO/O7P2oJzIACU7OE4hm7T6nGkZkurJXBgz0cjtHd
0inNNDNnCTTPIKgGFxd4WFlg6xQa5+k7BW2Q7UU7/6L6+8Ac4LrevT28AgH/FpN6JMFeUnE8yvON
fOHc27sTeQia9pY3QNpnUrRQt+8T/lNHS9IEnZDE8PnHmHn+fUPCKmwZDg87Ht8g1RK9YLjagsnD
QMXCFOVD04BHozacCtJuVeJbwV+EtN9kkxSwLlb9LZjy5OPZ02WraZ40kS66nntkFFr4E4ImjjX4
hdbfvINV/aRrQnyFWDOlmd1lffAcmu0zXn415ucbtABRYpDKhoqQtpCHN00MsOgl+LbRKPZsY+eg
ROWhK5hnRdgQvuXZ0cVl0l4SBgx0XRWn1Yj+hbjvopIFDBQGSIQP6PqCFwvL2Eq5hHrlzHlY4tmq
HXjPdTLENmQZs6ClG8g+lzNyjd7YQzEs6vciMWREQIuZm718CFO6Gp7suKrfv54zbya1Y7BPv/7n
HiByvAS7e4sqO8oghmXnYXjZ6AggGM6md0Dd/bEnzwTOzZNV1R6odt6TJygE1Tp2lITLJnrhNJlU
5luppLrFWeTcqVncW/seaBmUeKDuxlwDT0AeMrGD0PSbSqOVyToAqTXfW3mayMs9vPc8BvynfLRN
l3eKbHe+uZrSbQRevt7p+b2NMIm9GouhcsyH+75phohYGKq83lCCf6bcvq08COy5rOgvggJhg3JZ
k1CyVXqo7k1G6VPXqcccb8nDpiGhr8YcTPTJBF1mdozo7Ae8A5zD4cl6plisp7e0tCEHgSdRSjtp
uSwyhAmIYjdsoFYbK0G/O3xXnREyaczZgK009WgoK/dKEjam+Kl4chAZQjRisUbk6af+zkTpdzRX
SAcZKJoQBCL62Xh8T8SHJElOfW4n3rILbrmpVx/YQN5MqD4cJKYyNIBikZws49UBR2J/+zlXh6fG
x43w/CiKGFCSjm9RVEsVuPUUP5wBUQ8SjouPZGnE6LnrPIUKlZX5+ZlX+kzWhra0UE6ywgiwITmm
bEutX0g5+49Wdsy3txzm+PzMXFJ8BPN6NqZZI1btXV0mPK5O2Nt4hatfleQXBqAvwa2kSfoIlOkd
hHiZ+4vFs+0BuOvQ8Z9GNqY+f/5OaMSnL1p7ymeTUBAz7a0koDARnk9vCYVyA44p53JRLZ8GQ85I
FuNLXIOzK/VeVREClRCWcQgXbpQa0kD2bLsEvecsszrENrIGymZb14q0IoJ3UQmOLGVXyUrg7hq+
fIfeUn9Tv9w65nfuSYHGLFZrzurtrGRC568FnDA+vOY2/tSUYGATGLNQBm3t1pWKilMXkeK4pWYx
gq/YBtjCvm+YGh1M46rzez6eYpeWxKgc+1UuEUeqO4fHCac/luNqU0lLjHiJ3F7E84/8PPTc32xA
QVRZ+VN+kXL5C4GsMF1pNrmSXOrQSWCGSk974wdZ/T+Ws8uBX8nQtD/XAw==
`protect end_protected
