-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
v3Ip/oxBKttrK/3tzyscUJH0T7z3rYmUZGi9mxGOKlVDC/l8PrIgS+UH1cij8s2/FM64SgnjWCRJ
94RVCB9bUGE+9KTgkbf6eM+9qqSmeHmRuHbuIcU214V4dKMFrSFo/DklePkN4x9APs3tjUrUDA4z
OcL9SCNhtjAKx7ulBbtsRNqkBXzzcH2ww1dv0T2YZRlbKqcqTSFNQqXdVW4+TzT4zLpfa37kS1hy
3+LnULFbJmjYv84AExg8v2N0pJuN1cInEuvtG7iLxxwiCtZ1t07qBPj3fmujnM8TWcVyijgEoKNg
lYEpeEG+3YXOB28cqKx/nroDZTgH0UKPqyTBxw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 20864)
`protect data_block
ohS14saQiuAzL+54hdzAQpJhdA5LSFAFQ/kMVQaqpLLkPSyJUvglCY3bW+sqffh0CaRKz8nCZ3xb
k6c5owD4lWvhRKjLhIGYiZr1901qJWPQxBk7GVNhEdrR/w85v6NRv6TTjeaUJBZ0y6lNy1mB254q
AZ4aR7cYYfWaWcqIshYPLDcL4GavC/WFzEGxhKbkW9q7WCcv3rwpyhaj87UnV7s6Am1+DeeWhO84
08nGR3AhBnsvA86xsKP3nQKEznHmiM5JiFz+7+Ub8n3q9x+fpSvS4YPBcIsEz8hrkccWekjAIMoW
wCxnWsqjhZTeignScKgTBjr5N9Um18snVW8EeSVU/bQUBxBhdbwVvdRDZdEFSOonrj4o5vou88zT
6LXGZlhI0LJq5wsXzRQ5FCP9KGRAgR2Cv0ZCF/eUa8Xi36lB9Ckw0g7K/NT1ar53jHDi9JDd9DG2
GVuKQkRSH1eIgtmbVV0pgdiGv2l16uXXIPl2r+awTu5xuuxyE65SX2jTpg4mnVSwKMF9DVhC7EQ2
ESKexCRfM4A5IzyDb22d0B59zqWDbc5p1edPsRG+RMSDmA05/awJ42gVz7YZe6sLzc6fot30yF3K
/g4pehC7+UdXNofLENjk9zCwb3Qye/UeHDnZMNOX6YDNk5xH6fj6ZmOPQNKfXkqzQL9whhfVEbsu
ypplnBdCn/EuyybZ1wMoLVwcZSzCLydA+1mM73WkH+ApTq9FUFFGyWl09PumuEPMwdqhHvaG+zSL
rwotsC939HNics7mM4Ppbeg+til2/f8jU2ZZ8vDOqSbjoyMaw24hfu8xG9JKs3KeIAeEmUFyjzJq
ko/ariexYTsPg4kUkcKKx2ptPJ/fFSsm347TMn13lWhWf6JNEn3DiI/oB0IYz72hzCKG+ArGL1Fn
6J9Zk/rVGQomrQzFzXiLmq7asVonssUa/Dszsc7HCPuCakjEYw9f8nDbzJg3Jqfh3p0sqmL+kH1r
kxzWTh1JT79mmEzkgFHhxb3RfEVNJTr4e2YPR0Ja0YtaXjCm9c41gjtHbWiN/Kauve9MV5ZbXmDT
G9CFRbiywYMCPW8uOTSRbOKT/CmPD0GSi5nv7Co4Jn972uDyJzDRIlEWeyl5SzbOE8lG3XdY1v5g
xJFs1Zt8Al/Tdsh7LUbZ+UULyzOYyWbPY0yawbyqVRmw2kF1rBKqLZkYPOeoTnha5mS2bhGPZee/
k1GfzZHNn8Fb7g2bo5evd/Y7QBJJX7gebcyU7j1oxQFi289uqMLgJEadK3Kxf02z/SKCsWlu9RqE
j+DJI3qFIYaytDwWJ48I6SPko/6q6cfIspoAQUdmRPZYwAWGF+o3k1seplkBHPB2S0rphqJ6d41t
GLy4lK7JiJd44262TAHCJz62Aobb9Pb/AGj8ifw8JcLKMCzjDllz/uEqLZa4DwYerz0vCn04i9q5
9FxXCjj0ijuR50CwQ1tucpBtEo9by/hEK7ypfshZNy6tbouoPcnsf5z64RjATXtIFylOjrwMy3UR
okP9x6V4KsObwRoZySg5Szqw5XglG80C95IbCc+iXtU1GnRd9Yg+x/b2eib8znpNqfAaoBvYXUmX
2w8Lq+Gplr9S994pvgZVkUuy2uaRVXerXQKUu5oB1LPyz5mbtaNAh/XvpMgmgdXPL2x2bsY6WT9p
MSrnppGWVKOkC/ZvV7xgdpafy04tun7m+3iKSjOWkeOY3IZ72oExKYfcxp/4PdfcGtAgQl6IwRZc
9LcktUw/ENnx+l35l4nTyt81+l4leOlH+5db9fG183hBS1huaAmvUFfSUnNZn0VLv0PTa4tGNv3s
NIvSA73GWEsJkwQ0Nx3zcGwnqqAa3gv2xo/LL2co3gUTu67xQYeDU3Ub8eo0eVpBOQftwrrfs/xB
Tw8e4ygrOkDE0ssC0DZNuAcDv5g4i0ttIZTVDTyrXZg7rqM+2XXX5EUrWuS8Kkq37haN4Zi3UFE6
byD/3lp/Y4eptNw3rBkaHQjgmuDvd0TKpdKYkOvrAZsSGzlS3iQFf6YitrWq0a85yuBFW7qoAOkV
GnQnD2VRFdY8dN2gAbgWmsZpjITlgEkRbnfdjKS2WcqL07PaR4RJd7jGrIZdiG5rHINxVLcq77ZT
FWhkStMlNIuqLseCLi2rKw0hzdBECGCSL++YDVmODUkqvALmh00Aehsm3wBrKYeAt43HWdZZKVa/
zZmvoY4PTO2m2KQRzCQsBzCSQxLEhpasjUoU/tYoF7qpoWXp0lAUnV5zEE+LSkpKRf+RgrcrMpG4
qJtYruQQXLojHJKTvQuZrrL9vqHCw0EC8urEaGX04SykJRwc7YO6BXQ3LoN/W61D783/ACJYVX4k
eT5oZuZLjEshfakZ5GOwFPyb1PVAq8d+Z8INiPMlcvOJO/jyVC7ZlAz8+M9/Vcl0IUhl7WJE0jm6
/4HF9/jGji9+qVz5tGqngSg8nXIfVAt/QzJ5Eg5PbvHl6a4iPV4Jfwo8Y0Y0soKgWTYCo6hQKDy1
Nn1ehV5jR9w6QxM1v824iTskF9kvJqQOGJWZ2d/y+TZJsTQSveBvpw/EZSWNsLqqQ3J8Ms3ossHp
oCi05P0Ud3+vjuUgbE0NO94MPNluhybygn4yeXVn+8KVptt2UUbC/Qa6MmeOD37C/68nt3+JMyXf
vudb8I/T8+i1xlqPzqP3FpM9saAxMO0BoeXHXEw6Fo6Bt55n1st5ZlMfeXJ77AEqgTic5mAQcFqq
uuiUqPhLaB+iOQmHc8+PPLS8ldufVGrbTlnmuaFyuJcmd7io8wyAzurrsuyCeRQK/xvMvkXcXdKQ
69AulyYLcgTBRMGC56lqo8VarwJSVWZ3E/JyryEfAFirpmaUZPnSot1wPFs7WRkJ8n/6R9Gd/X9E
i4K7jbDZqd8vdwMd+ixDTugjoogyNZJLNF4DGbaxsIKZa3bL9XT4hEmQ7Zj18Fkn7l0C8CjWGjek
F2HgR+CAyZkItoFo+zAKu6Ad0I/NHYXwtSSPB4c7SD7tiJPFO7i1+bgFlKWLvyZTF5E4Ad/66DKW
khkl1PLXHP9/wXym8QpSkUhfk0nKJQ38J56uiWhELrswjU9HWc/lRAf8grwU8jfMQ357u5/tsmfq
kDiToOG0KDIyN4moA4GJ0DXZLNlDFyBRiAjjRd2XtBgDJNDL1HzyVQJJ+iDuMXOKgvnvjt8gCKMC
OMQP/pwdqwNQRmLCPkP2p5L+wfuqwNajGPjuf6+J3wpHc0SzM9FLSh1XZ2x2273GQhlF7o+KYKVO
KZohDV3+7Wx7eT+B2p5M+wiww0LJIIxwj3nh34L+pQIwoxCoXAEA08BaDnkSlXQqObe4dBlHCJMf
fUxmX18ELAsm01pTn/GP/fbBbjo4k8DFhJbM5bd0ohABV3653QYepz/E5j6UO24JfV9xGyxdq/M1
E3QPr/ciuQvckH2lCpXPtjj/gptW6kGVg96C2JiXhGKx7GBPC/cNUmmU1E41Fw7WD7yL5rIHm4Q7
2xlRCBM6UYu5thRQqjD4MOwVGqnk0DqF9Equ1KV3swRp1uywY/hK0U51ehP4LyMTwWnjMSm37ezk
AexYQ0Fd6P4tfS0NTwdD1XBkPXOySgWpWm0xiPT/HwW/l6zy+NgNZV/yAM4VIN9H3pPIDEeDH7mp
PKyS88+i/lCqOqdZW3HHMXKA12Mylitc64iQi1OvD+iFbj9FylKfyEfRsRsRyBghwDikodDv4ID+
ZvA/TefvzYm0CWeZSC4t5sOO6d5vhO9OvRy0G7/h1n/cFKup5YcL+lkOq3iQP9zh0NEY3gzYfedK
pImFYbBEbJDfCJr9DcJ8GBi+x8NThXjDTIMGQOg3z/67rr4b7Qmnd2lT29FaavJTopqSR0E7m1LE
KaAdjGWy3ylTgPX+tyofrOEOaTWRcFw3crNVR0g7XpvLqJAsTA6OKvA8zH1IiTgotIIZFfw1Uyl1
+EtoRIEhPPubjO/2oa6EfNZKzTEptIYFWjwsuFH0XDnaYFQOrLMFDeMUz8CDCGy9t0q0q2U3WUXs
wKAY/6CQY5/nebGLRkj8ezT1aMdyrpjA4PoSwLf0Ij6c09oJhp6jlOVzU2N5JwgELM0LaXbyugXC
K+QeqcOhyCsXPh+3avN+UG9niuv/5H2qubmuJe7mZlCI4JAdkEvF9ojftJm9HNo8g85e1GaLskaE
WXx4soJaRRIoblbfm2Gi87a/669kkymoge8QCMai+9hQS5moCkDtXdBV4v1OWMBBgVOsq0dNSkY4
df94147JvnNkTTrug3PhK5JZVcfPaaxt9vDSy6IrZYoUPOsILDQoAV60TZrCV0U8QOpeXvLAwlZm
Wy0OOfW6Yq0V5LH8L+LS8G6pxR0LTeX0NLWdeYjcxJ2GrhrXcdNn2uS3KBv48o0oOFf7+cZ+syoe
LhueL97c2G0ZlEp+m8Yu4cz68UdKKxEkhRR4vYFckcZpQD7csPVzyz6DVpmCmosQe4k/xyKwZpey
fvgffxRPrVkyvuBuNOqTmU2IWpks9c6WiSMyBxqVmVbsN3XNv6b98QZjuXZ+h3cpHdGz6wcRn85d
PHMcvVHsio6/hFI5OAOFbs9inc3XUKZjZtr8ateAeL+1op3eac9MqenGTeQGyzCaiwRBABAIUtlx
WkegkHm6S58hbBMZljrBC1cMV1hT42ykzrKls/q3oDJ2MWtveg6PdVVJriIGsfkGx8wUEwdn5CpS
s5IZEw0N77iZ3uHagW/yJ4qXePWicQw4Coink/qyarezEDex0E/f7139zeM0ZfYKYt+B9zEX8Jgk
gjfDPj3XxX68285IXT97zzipjucgXmi53E0Pk2Yzv2+PKtsCKmH61M5HSIXoNMcnH7TLBU0fKk9g
/nWMcr3obxqUj6uJBurpxJy0cIyoMJhU2w9FQzOjbGWgyTlWvxmqW9wozo1OpJsoU4Hs3sIbtn3r
slG0a199Au4sONdZssA/rW/haBwPPlGwhvNJzCPcFszK6gKvk+gLGYPMu3Ie3mK8qA6CMqZDVo5S
FJ+eYbIm4DBAf+SsYd+eN3B0ZxnOHEelH29AyL6MvyaY6P+R3r7SxN7rFFyReO61hUTXN4RgG+Fv
90oW/Y2DGrI2xYf2GzRqMa6+1KSFP45gy8/iH/IU5DIVajCePUmtc0oY/SXe6n9eMrG5y/d7n7Wc
j1ObTbq6zS2Oj/6TqfXaOof0+oizmEP3RuWoHIZ0aglNRRNIh7aWO/TsFTYxpX0mXOZKNCHQ+aA5
+kHEBZRNWdj7C/SsIWb+jiyeLvoE7btV7aGpgdYcqDdoBy8EDe/pAxItz/unYaL7e4IW78xUJv7a
//OzqG+HOF446uaRCIS8fZ+6r4xWFRfI7tlNNa7v/4f9D2AjHYjufiOZWNJauMGWSf1bVwv0Xp+z
NmsUahL2bS9JpAY4HPc4lYTxwJ70R4AQG0J2hPWj5fuQTgg/eCbvygkon5Y1mycT6gGFDqK24RjP
buykEoQ+5+bqn0HfpbvnozfXpXCfpuL9lCv6iOivx7UiI0N+W/PfxYMdF22arqNmsI367ET5RZ+d
8YG9jVWpuC/56jGptiLomXpPZxnDBz8gC5Bah0ng3kuFs/zzLYVmRXgHAMDmsn8u9q8Z2cZL9+O4
n7t+PZyL43yu+0jSjMVFfYt4hRSjOxIivx6lfUP4XHcFrUXYX8OulhgRmSkqLwCHdfb/ahLhAWOS
1tWYw63CzhXCXBW7Yur/BO6V0GHNHWcRh8IKCpkey9ER1sCJVKdRAArr4SGWYyjkqzB85+D47tGA
Lx31jjSrqqaGEX4GEXImCPDXRXDucHVqQXu8bXIfVBMsfvvWwTU93VTy//wMM9Nu4/pn8t9QOFRO
JaHAV1/69IR9zrBmL8RcTkubauU9x3AuwlK3UEFqmo6GEcDJKfD+UzC2ROLpNw7w025+79gUJn5y
RtQa2l33z0HtBlSMFXGyLsx+pTa8P7k/F7Lg1HSNA7JoR9WMx0q+z7X1kViL/SiLUc52F8Md+uVl
mhUolbzWw48Rac4Cr9hsSl/A5DRbtzJGFKoU9SAqZsuUCuWqkFItPgV3LZ+JhdZUrDhm3EchbbwE
7LhzAUagMwK5/79Unat+jUGEb3lRPBOluZpayWwBbdWmN+leKTstmj/FjQZPSoFBqc9OGwKXC5/n
CHfx6jKZCLOuFuzgw9a2a/r1TOKiPmecmgx4BZ+JzcOrg8ncl2rayNJJeAz6oLiFlRSasJRyni59
am7V2fc+8vZarLgpM/y9U5LBnCqKoduAIlSc8W9Ahlae4Zm+efNzTte7/AwlXmcAMBP//sNNkacb
4NCfzHH9dFxaegcBFj5SWjRSaeSKVNoLMkBh+dLwmFrqAd7CzlAYs5IUk8nbCb/jOZ7/Lo5R9bay
yWHHNovFr6gWuW0Eob5olerovvAf2GEfUmGnu/6ur//lOm+tB9GNn6fsQnBBXKKzvnX8QxsX4Xlr
/oTRfluJylxlUjjm00wCyAnaxd28AJVIC2FQ/B5FZT/Zu3Z9kcwmJxKBOTpHaWTuRN8gz/jh6N5p
pKGt43czthzaPRsQofX1q0GZVAz+gWnKZCTAiGfK6alaOJ8JWxuTd4VuhKG+TF6HJDmF01MTqc2D
70GsGrPZyG/8n6J0Z4lYfJHyQjc8vcouChMqP8AdXZ82Nab5uOJelLpriYUEj4b7n5cI7vRDWQx9
ST6NMEmHJjoz5rTNXRtbX6hQMGpewyMToERwR0clHzlRfiW9cQ7hvvGPDqodzj5uJnxOBT3hhr6+
pac4LXZiVn0FuFTxCO9KFI0mSba0XzaX2at0jVweZvqkWE3mVtYoTF/k/Xy/ru2wk2T6kp2HEZ7z
SqcuPJRNyWPeFzeQODi9epeAtzEkAikhEt95rz7NHdSOrEIeeH6jnZj3sQ22RPRVcpAvjsjAlyvc
CdmwcSyFaoPonaKDc3mw9q/6KmNNPm3/4yPW8foJv+y3qlj1QpJg931t56eUR7er/4bPi7Iol/Iw
oFX3y72enjXJm5Eh+8tuiF8nxcLnp8lNVYkEairKq5ESYUcT+Wg1236g32SF1yAj9DgQMXRz1eaL
0CxgMFV1JcBWN/6WdWWZSZIOHfxBAd1euezXIAAkr22b+esQgWy3TRSJ4Z8/mBYlomJKXrNjx72x
BeGMJBwA9gzAI0BsOj/lMH/U7EvR8e+Z6/LLutlNHo6XOW/GiKuYhX4Q3bkXLUxEQZ2NN7NbiOMZ
kVj7rcZJK7hW0GXeO3Ft32FyBMbAeKxlyX0j17p2Lff3WA/FPGN5OgwYN5Cj2aCbfdqltNaUFh2b
bdmN1FFCFjsvDPUQipvhO8zrV+HQRVBfJIHDn/ZF4dijpw5SJ5FfLcOSeluUSriSeCuzP2Xk+Gfm
8S2wN8SUFVUdtXL8Xovv4npgcLmOpRSs/NHJNni1D7NYXi2iLTaXlQt588hU27QebRQZrcVg6/W5
cJT22TT4WmB/bNNYRdCD2iSxEn0bTZlMgUG81pBVBrJV4oxw9/fd79C6ZGz+w7K/HmuKKL+GG/Gq
swMXx7L4iblKmoULzWmyHNKgJ2fqFnAIsSzvDfVHKMwOTdE/D6koYfwzeWzcDSSQlRyZPSESFRpo
+2rrjpEsi4fMNmAOymLNBjEQGTt1fLWCYrjQGb5orfNuyufdgVnmfNbuI/IsbFtC6hbqK5P98CUf
uE+bxI7tXNvIm4zf7k1zjE34Mtev6JfPAnEDyMJ2L3warPjhM29VHX1/SHpQodVekSh4BXIKj8zP
TNJgYXV/fOsfTSa/kAl6gZybGOHMk5bCwgF7BVPeRXsX7eNXjDa2EvbUkoQybLKiqkc85nmKuad2
kmJaXIwgtRdDngqgCTSc3mSWS3Kx1RLqxT6feBUuUNEcM8RgsU1hompHZW3UYsHdhujypu6wJQQ3
35N4QKkaeikaNJvNl69Tplb76yQCAmXxEi7QDN0l8N3rx207C8cvm+ge2AWWPLhheMS2MoajVnY9
NJiZeQ8IXN1k136ywpymDzF107PzxefuMSBN9EAUrvm33f0aJQFYvcn8k+nhr58k4RcGBJ0LSvLS
P6MjSU6IYCnCJXgMDqEOberV+wQn4bQJVc9tR2EqhIUXmxXw/a3iPB3z6F3Dp/kxzsSuQKjCkQGn
6YAO2vkDx232lcVr5uKWuE82MFQTkYCUYgCxstDlbjX0N8iRxXj9TWotKDBy74CDt4bj7EQ9rjWH
576wh36qycdYqI+++JauL7AsWsYiBBW05583g53wuO5X4oW7b06CLacdyjJz0ddzrz5ZA1uaJh86
EYXpDTLD3XHCQ2UcP6OMVfd3/56txvocckrZpEwb0beQ1oMBH0wPTKT7wUwJPYvoXDSPop+AXoCF
KzgkDkFQ9g6C7PxaZ/Lqyqha7GBHSqbqtiWrRwMKoJ307TJ/Je5F+etl+8nFp7Osv/PpeiNwDeM8
xb5qX31ZD5iyB3zOxFK7hBqc3TaaP9uIv95JXXGaCu4ZNaU9VJTS6RFPCCkVgwtuew50k+XPNiGA
xmMBOQBKaDVT+YgXQfJGLX36CwFVGU5t6T5LZhxac6O2xPdiAoIDAQhnyrKbO6y4tBaJrlhSaxuj
Itd57lTF+yyg15rSmlvpOyahiEdhDlcu4JFIpXJu9xdAV6T7dNPANl6AK9aBnxWZSLE3jOARGvz0
foE62C2fclZSBGwSRs/6neJjB6mH6PpLFUPUYZTGNRBH65G4AjLV9cL/XEDqae5GEGzZyCgk4lha
iv1VcpR+UV6U/Qx88LKo9WPUSjzBRY1/aEXVkEwWYriK5HCSZ2Bi74VUQNpnonjsuQSkgcVzBXlb
8oaiX1/xtMNkhXA1cAgvhyWXQlj4yf/DeSMiktowzV/7nMffQv3N7cWnATwJsmsxMUEp4zmx82XG
9fhuH+NOAaPJCNRTLwv4iQm8s+Z14eAr6lD64wYNSAWin3VFhff9tryhfW88IWI/UTUS/lW4fZIL
fXh9dkODbM2HSAKHvz8beEIEIxKr76+Pc+7yIzL6P7r7JZtpIC0MPeUO8GhchPwkhdTNx6FJzuIv
KS/erYQP0osn4DUxRAe3jagmDPoPioNTEh02ebg3H2QvKfaM1MtgD61s4tsz/KDCcQWqBk5LdVZ9
IkBQXihHsmxJS+ctRQvqRFb9q0r5Y26DEeS3IyLE0iznbbOS6gCBJv5vJQpqXH7Qsal3jdQW7Ym9
R/EgOlaA/aXknItnJMD1kaRSiU5TPZi7EQB6jzFXXAVLODQuLL4T40qK9WMNCz8+27s99zG9uwk3
qXj19sTHcoUHQAy2I4sl5DFYXldGeDB3cAIkWKAR6NIXl8IMJTBMI8zaqK92uSpeJefjNeMicI+6
BekFwXaSzew57tLpfzC/+0Iz2yfPD+jCRVbYBwUyk0vey+2UCJrhd7uR2/4XfYHOpWKLi7tqe4ho
1UEDAKC4UgLZn5gMTi2zMAJsQZ0kNWW1hlc2vHD0SlCGm0VSuf0RNiI67cUHrvrYRdUNB/H8nxnq
59mTknNGw9F4/qmIBo1zriwc/8PYe4S5RG/YtDpcqUzDQ3SMuT2xLG1m4TvmzU/7aLECFwD60Ixn
vJvS7md57YNUvbvjs2g7z2g+g/6Nu1Gqbj98yKah94AjlJvlaRdIcpJvGjispr1bXDbbd5dgnEai
pvIpXpwS0IM+Kw1AFZR0Jp7E2nANajLQ4uDYzeNo0DD18KT4VOipfZDweBsbKbrcBTWRh84LoiOn
bYsKB/ahkHKHNKdGJt+KBAVa9WCSYQrgJVj+rl9MeefXLnt/+W2e5s2UsvQkcRUeFKB2GyA2YCXZ
QC0A7EZwyhB6DCuUWVtoXWs5Zq8BkGhEJrAuqeIvQ2PirdxFnNmX9rBXorXaww7mrb6FbvrISe0T
6MLMSFKllTa+u+HlawC58jG7V4ZeuWrzwSXPOgzFtAV3gHQ1rv9kjxSzscy4FMsA8ZCJg8s4ge2w
qAYs2o/wLX6X8f69IVUrfbQDAw1iaP2sQOPOyQLuCQQEgrAoEV4CrX82nyLpx2kCgF30Co5t+q8c
oDVbUXOvxpFTtR39744vPifcS7wdkftkXhVnU1uvj+X0baVVQ4codTE9EKYA+2zrC1wvv8s63kKM
qBm0E7gg8XP561zeM2wg9li5n804yZmVrpmtJRQDSAjlbZXhRVRUnLEZEN0+7G+gYta+maeVaJRt
9UcQoLQeSUw5gsKcfvDJ6xzwDXmNJfeh+254LSC3SrI12CLLY5c2HDFuQdDalon4YiLGZCNFa2sQ
Si5Jw1A1eOcAz1RKu9L//5AOSKu1cgKRHGsAAKmopmkpYPqCrxXjn64KmbV+LxWmnLuTF6gaHjSa
1UNAW8v7ECKJLTpssY/n/zCLaJWnxGJTLihIeryBPvpMIf43BmCt6NspiMo1s6Q3Buq+CWwOlr4m
pqLsfiE9Tqz9XreGm1wZQ45n0Q23fgJWFPOpFNM8wntvfilZ4RYuK7bg22I8dXeMvsOnTzNjT8p7
dQW+MSO0rrIq2PpnynZUa4ZfKgLMGvg9W1Rdygf6ZPug/ucVVqWOzFo5KEBbSf1jorgf1znz20CW
5snB0/JjID7Cnho2/fMkpRpq7WMLN+wHVipZcYoaq2YLHk4rTU4YstSmiSWuLJ0WXw0928Mu1NV6
GBONq299o4Q1EbXaxwMMDO4ku4U7u9y8TET1mug6gHViUNKrrPnROMVDVKDhXPQoEX1jDLJjNIlJ
u31ZgJb2ZAbiLENZKvwZ/cldgZR6rHb16R1bOcM/VtdBle/RNKBYCzZwVmf/o10FuzU9q3WvOwac
voSFsio2FRNGNIhtoHqyDGgBS0lL2cN+d95SmmXenDQoB7WPzyz+RG1IcsgHSHQt093TvHdXMa6X
li0t4ezxfLbdMWgiDf1ro7tdfPcEj2mBja6Fi8AdxjdiCQJIKmdX5WsRVrqx3vvLY/UNHJqHvIWx
qOV5v3+Eb1H4oGmFi1X648mx49S/W9wPkygRKc/Gjw81wqlpAd7iA0O+5GWi6Sd5xpGG7+JeQFIv
P5CUOhALP1vFtqUW1gDanpBeCLSiY49aGpWT2QlLtvKZVbcim7H6pv0x6vZvni5P+F59V+Wc5OTD
i/nlZF0hDWvCW6TERrJNNs43zbGOtq5uT0WjHTjXh9xGcMBjfVQgPX1jW763MbiJ+IRCJDmUAHGi
SAiFAzxRYyBbJEzuWrGwdEgNGGGWGABckcYqvqhgnvoWwiKu0gOui7xrzfczGJBK6r0+vvGttvkJ
q/HZWk6xBGfGwM+Gm1Agb6KF30I0j59z9BMNqvckJbyvyHMwFCeaBEwth5lPi04o3NlKACTeFGNW
YORRS9H/d3NRkatj3kylfVU7lJteJBcqk5+jWkJC8RrWeWPujT2jL7l7R9KQcCQdfUyY7eo1ie4o
cFW2a3uCWY0lExjtx0D/kLqr2FrqCPdMVvZuYIN1vXpSix+1MhwSogpbdce4VcxC8LidpZWnuLGb
T7QtgUkY1xWfJSCPuGaZvHUMATt2yMWqH29S9Pae1o5LUPik8IShhUgx3JLu+vUgaSQwD3Br1tJK
CmB2nCx6T7mv+Tn7/OM6UHxVcg2P6F4CVDIamkk8MdrMOvPmCvssIkrFv27kH4gmabMokpo4u9Px
J6B34LgmqmH1lLl6Wx//4Ssif8YPH5h6kUDp23qLyEoWVL2N5R7VBgNinYSK0CUKKWgsxgfxfruc
bsuSoaTN16IUf2FnXEcN5soAq+Vn3hEzMut9z3+51Y3jIKPI0yJeEdhss2Vbta8AXBUfK5oIvGK5
pOW0qcO9lR4xEMaqYOziRzlC8PM0IIuRGWelpHs2izFvUfwXjfpSb76Kv5q+7WY09g4qBOHZ4DQy
ROvPKV4583o9QX6ffGEbR4BhWQJcA5gzLb8Ls1ZObFCCRi0JPA2Eu1uHE2ckOW3E6flsSTfU+Z7V
k6pKA2Q6u27FVukbDmzXR7Wa117rBPPSNQUn+tHR0gHJ+AOh6m7dBL2Zi/0tRZAHlk+FHVjm7VvK
Xbe3YF/8qHlD49pHEm5qUb5y3Je4ak/OCipAPK8tyyG/DgbjosPOvpkL7pNVhFq9c41I4zrA8DK/
ZVuhr1Wq63DWEkuul+U3HNUL5Z5NGgt30iY0P7EscJ6il2UBWkMufKJPoFq/KCNmNjEb7z47mHy9
C879TAiK2h5gJA7q3xhjYibN7rKMWK7pZVDms3PZZlGuO7dljbe2U25StREt2jD5Pv/VVCAIAVWf
AoQdZXWvO8EtL5nQOTFi0hW8ZvqrQR6SCslETWnZRWNkPdSVHVUSiNBfJvFo7sYq5z1dUBaZMgNC
OU6eNhHzkrCm8raglhcXm/zBp146ikrygS8XciQAYD0t5LnnzfOq+clgsOFQP3hjjLoRAORgv+Vk
Qzgxj6E7BA4noORllH1lH/AXdM5s8qfFG1HNZkJneS1c7aBpU0CYoY0xAeCnQtMWBFBpDCxM54wB
nobNDFoWZ87UDGxcW+8ux/Qd3feXsnIPxVCrnLiIx6OcByr0P0MlkV4c+BZu/qw1qcjwZv28gwK/
b1Lc3BzQIIATtDP+srVRvrhPANfB4v+QswKSLRreWQNTR4cKyVkg+0oE7RFtRuvvkHxKrma3PbBh
bzO07go6E0BodpACsaxYmvheG3VEZ2owMsHda8kqKWh27+fPRlv8HU89zalXuwFu9YXTRux92ciO
xAqX09z2zoL/KvQF1E2+7Err2dDAnW+9lt5ikx/HdVdADqkXqB8/ZT2Qo04SCUYwimbOsKYSaxPg
c2eJenBvd2G583inin/2/oTZBbApmLSBjLrNmuPbDihMbYYRQ7Rh4/ffXFLgcHJlPb789b6XwuXl
6HMxkAdp9gujpTR0er9ZoYTXqN/J3WygRnAADUA0+nm3HwCniUgDxhgfhfUzBcDslcTFEPcLEtg9
oX67Hr+4Nqup5JjNtAxRwmut/JGVdEuUn79FDddUAByi1IlIDBeIq1VFuDhrn7DgFnfM6GHrQTLS
fnB4TbzSaupz6nwJVg+8hFGwY8esbc2QBgjQxo+BHNahqM/ruYt3oXMQsGfshMBK3U1NUAXQ6XJ+
1bTXcL0hD/QEJ/q4yzuECUqMChjBS08swodzQ5OTooM7YH2ghUKOHYZHEp45CaxiQ2D4lPmjJgDM
AIV4Iqndom2d8c05qLFjSqlCMvj0bS4wS3rmka7aKYQsO7blPSMR4Bxyte1OfQdEpuewNHKRV9TY
KkEIMICf5XDg75wAVSCW61L/NA4vXafRdlewbQAUVGcjMhqnXLDqAxBX3R567NYmq+JNTxanVl+Y
UH7+3zqpe89SsbbkzBJfgvAOCuhwuntvGQQuCP29LM68rLHQfXqm30eWHjiyy8GWzTHeUXaS4qP6
EJE1Qs5tzxcNF2aly1FXe2V4fOMfCFDFspU/3WTDzPZTzvDUxLbyv2p+bFlrVnPh3KhuSDAT5+tr
2MIV+ZPK2k5t/U306UMBEbI0elGDAALKLRioGfEXjS1kQ5zDKTMIJljHOKoDR1aBvGAc+RfcMjOL
4Uvi8XtTvt/Azbcbf2Wqq4e5bF5kqnGxhiVwwKdF0ZvVsCmoccyyy9K2pbcBFjdox0WojeKCNtJS
USCWVAFzDKld4GynsZmYOQMGF93AeH1nAJZkl7Oe1UInmWdcI9v225p9ADRrLsW9is2SFqkCZY15
w4DoXRirPKPy9WtULAMftK0EB1A/xdww/cQmTzisXY8AZaUt1iMs+WAS5Tq/5xROZHhNxO++ifMU
meokta/7W67I3hG0f5f5UBw3/kCCdToGyrmmDPKJOT0sCgz6CTUUaHkx2xbOYOotVZhMD/uVklT9
taaz+HY3wcpI+vKw3RdmDXij6kNMeqOq95ZZDQ7oO04h7R/OrSbGxMvffxIgO7qQvUUTnysAZ/ms
/hPIIQ6cUV1rfdpPVqng4Bi93u4c+sWzzvnegqUav8Vsw9tQNFEHYBeWx2Tgr2tCG36O5IEFYi/j
kCSeu/cOkoi5h+coTmKWEc+iKFnkDH509MoqoWmaA7eP7t3EUrVc9FvniYDx64scoVBGMH/ffaZz
aui/9jWsRDd3UR69016gchCDj0/+5fWA9NdVb76IGtMUn1I45tmEq3PHPcjiJrhwCnZo3q5l7C8g
NtBFemiS7G4KLxi9312G1uRQOQAzCgmltQx5P1WpHYyxBi1QQYzjDP+F5qRGvcvtyoW39IoyimN6
Tb35iKAY8SmOaCaGmxxlVggdz+Jcs62yAgOmcDJD8stz6oJb3UoJ5PogdQ82z9QrvUazkDVd7eA8
lokmIVIpvaJl0vNWySjIXr9ilgUJjNyqLgVJfX8L66mhlOXgG/QsS3wwZYmJ/9KIRPYHf1YvZH7L
KQxzRAF5KIDOY6Stlqq1CeD4Pf2iMnEMfnW9hXbn/lIWVXLY8enb9+lioMYIIohqUJvQgBAx7PQ5
RTAVoCvb+HDwmm+ag1VLaLgVVfW0AzhuXEt4JogUQi3v3BUioZPKbbkY5B2OT04ruPhAEwlRSX6v
l3y4VYoLFgZWvctnTQAXN9+p+c0BQ2EORUEKbFANu5/49HUasvoNp6kbKwfz8b4Zw8SEslE/nkkc
m94XcoiM69MeJ2XeSERrXwrZqvvGhMufscDIA5ry4LZfKbO3hvudnLGdGyQ7KhKdIsM6z89NZotI
pQRMCMPv2F/INWc/M7Pfppc7/jWOLTOFP4Walc7MTomv7El753nOif1GFhpNGzoS4LE92qQdiksh
WVxgh7JSP3lA9LebPABaigU4yBtWTlm3Ic3LuthdIu2yoKcepEuJ3L9hyXQ4gydl3yMg3Pulf5cE
Rv949G/H+GkM1D1Zl6SgbxQw5zSAMdrSrGIKLH/wdSWdOY9cdByRaCRPwisyoctcPwHwKN+uZBe/
+5SKZoPCNsGdLBfs9zLUWuF33aECjxdBKEUaLIqny/XDdCxwLgEr22f0ZZmOOoR8vqNmmlnUx27c
W4ZhUDbhm1ZZHvUtYL42roiTIGQqzUECKRldbNDm8217i0F3llwHcckauaHDZPRRreKXx4A1c6dM
wAvnhbpvMZifCs2lD5UK1F2YHo40WqkfCWJsSGG2DDjlIQH8D5L9eRgqLk8ySTLlE9YV4zvIkDaR
+YYSS+tQFRfJ1SJKzibI79JNiQgsxaJtiLNvJAnpdwqBzZQjSK5oEkY3aj25F/1uZsxSUBfGISrs
4D0Te4raLUyasUJN+RUInGTy1Vj475w13vobOmkZ8h3Vq4lNq4/xwLw4U8yBAU9ujuqtntyNmZoJ
X/CD+EJRsbX/E3N4TI/2VdOijlqcdC+IkkRRBseoxL0mb+TZAFCMuSVjdBoQdVZHXyaAC/fGA6aJ
e6LqA4yNV0mKvDg2F9q+Q42y54k3fEfplQt05wPN4F+ujamE5fC7v5TmUkoJi9IIHDfEWiRkdmg4
dfrgW1NZLS6rCwSiFmhy4AyIPGeNdAOHwireASOruiD7bWj0CownZspJJPBkIbRJsTnwZHu0jcN9
D7qzggzYqtvRDpUmsXXiRVoEps+ArgoX3wUZ36vRMlt07DtP1YnTZ1akn61K5HVv7hBMHq5dyzqh
0rY7klMRDCo3ydeUZZD9us21BuKiCY744FD+Wk20QXrQzB1NjNmyOx0aeDIs0XDelJP+aN1sQJXx
nE7tB5mO6ROmH5eq4Qufx7zlI8rFES7wMx9bN2efHumtH/ZQwKL0twfjl5otEMWdnwJL/mm3iFNw
NfTV/UdAqDufA18ANrJQvKK/n0XP+/D78WyBqmsQNCYrFi1rKLp6KIeDoVWVvR/gdmpzZGPIBOyi
BwcyPr1nExTN5ioH1v6zcbobolvwTVxuk0ZGddurnK2v8G/14+nLSc9j5E1BCTiq2pKF2r3nYsm2
2LLXcD3vS+HC5yzJsHr7ShwvxNlIydfCZ4gKW0XIgLj564GR1VrSrv3pZ632kMU41fy2ouwNd5r9
0fkwPJzgWASfPsCfIPgnd8DNq3UkBuJwe4zDn4OLLd+3uvPZXxuk7khhad8mlXCSmS+T+Eu5XS/P
JWOvVyhKZFn8x6WSy9tOCAwaUFTZjLkisPnX7Eku0iznExjKrcCNn069aIgtoNoUa4myYBmmOoFL
W+R4GBn+PFKt6J+U6f/R8AWG2A1r764elq0nrKdsiNjap7Uf0H/BFdixF2dJ2UF+4cCUBAePsZBN
b60L3LEY4rPrtSMwPdBKUThU/FdudgW/ZNsolRwGOqx98Mc9kulstreG32eDH3o1CUHUDvWJLd5i
V/pFChz5zv6vwRslKc/SlN7mrCjSJCYmSqHR3PdSLvoCUYNIMzjtuZTJ/Ofe9EJxlDEmWTABC1+R
vqTHP+S36ngAPFpI5p3EHCKHCvzBc07WUFIYZvg5GvUkvdAKB7JqAJ1OYn69fGOJpO7oGWSVt50T
Jc83E2VZYNBvRTz06LAKFNFapg7o0+Nw8mrYrAfY/yAdRf4FzdkcbZucGlq+0S/l4dEJ5mRak6pp
exnhT3j+sBXw5vAjZviYlqyh4jbEeo8e0wmxJl3QKIW1HZiHIdv2ZTEXN7myV3TPJLSgM/lFwPh8
l8FQFV9HM25t7BNKdfmRdMdtPKYfSi1K2d64820N5m9H8M2fuvYJKPmLCK1PyuRIpIv/t6og8Gw9
WoxQuQ/sKVRXHyTBuqxRdcKySsUQVfnx8obA9voEVic05x5XuAvO9HgHcO7wyfoAOebnN20whcAv
1ZEQiiDDSZQ5s6kRgXlr1tNzmYpOi/xRAEMGxKOO/3r8PBjPBFYMMMyfFoNuMNxwFJZYK4LNw74J
JhCbqVUvOxaPQ7XmmLiIJZ1v8iV1h0xv4a3acpHhxV9lJ4eMpHde91jHfgr6IjsqTno/79yCwka2
s4VW7YxKT4f9DvNxEcIP9GXd+9TBDWrtSvSxfZE3gx9alKScSw0C4hmDXffBNelT7HWjdJf5TABG
pIg6YZ4j9VKnMJQSQNxp2ZpUOCgUsPWw1onRWmtfC7VY1VoZ/E5Q0snDky7ULRrAs/gcHGyyawmW
B3bPrMliMMDbzDAJK9TifpDYpX9F43zvVg3cfNUkS1F5BDctNx/yDq3BkbvBbm10gHrFBIt6N7lh
0TFpdwO4akTR9/JXxeACaQGtzm9jaX7UiNHvHwMKgmWRXoeYZBWGhVqSZdNAtJvd5rGUfQZovDM+
YtXJESrUw3NeN8GGBerZlxK/gv0Ev78S5FPB+ouOsLaIvSoa0gB4075TTM5EWBKx75CqvvyJ78L4
EBfPM2NZCxiZrci7DlHYO0bF8bkNHtktfJMd2jJidTjwfJtf5mB1ocC3a1tXL7hy0mjkNd4NwRA2
2W0P96i5zn12PUVlSKp5JEb6ikAewgCE5VpkUFRUQTjy1r2DRZj1FttTV04vyb74GY8KIpeAQOMu
ZtS2MEERyF3JMIBpK2IAz+C6tDGvBAv5o0gA97DWZxCFEkAq2FhKX45ybmAMHpl3BkEZpGiJSqli
tAf2+29T1cI2zQfWnPOeM9/IXR/Kwah+zlUCVgkugg1uZAlzAqM5zGyiVUBRgtrU6e/EArQVX+EU
l1GuDfCgWiCxw2JCSztRTDFl6+Utpb5sBaCs7H6YwsAI+LUjA7Uc2Uhu/aVc017kCrWCbfSoiZDG
gACuMZnRsjdlIcKwRupFko+srxZocuTQCNjRrPZ4imMxOiHZMsD2vK8wYYnZE//g6spnltunBXCB
quTsdRbKgeuobJjunx8kUmIqgX77ofyyQIwAK53IZRyoe8wYg8m7K7gurMqFet6B8sAkJjqIvkKE
imqOK9HgBpGRAmHK2PZgn5dmVLJwuBsEcvOE1zcUdgGYBOoU5uDQShQTjenCqRxhjfvEpOOstBUB
X1Qt21yycwoGD/N69A7jyojNwVzCu4Cp5KV6fL0lBWjqUWY+N8o++HwghEMQYuiW1/Y25wGXRgCx
VwbdG3UBhRwgAd7tdBNwIuPBJh3V7EpjwI/LMbi35xiZkzR9GYnZw0JbgZUPXYK0dReOCn0jCejg
pU0kccs10FH7VRsedPQdXcXXppz2ROchHs0bLKcFo/kEDv1k1rB5ZcZXI+wolPCWYM1IzqQCw9eA
4E1dSlnjvJtPa0XM/ey+u3vkT5MFzI64zdtznOkNpktw0hDDw9m4ilqP3YS3tDllD6O4k6Y/FzXe
TJEkiC8u01dnuxbmWak9WtHZvZiBDinOiFE5hLl9iEgbnOqI7Z2Mj1wIs+4bMr8YahMbiouT65Sf
+FtX51W9GOcP/REOHDgdY2ghvFnOI5b+K1UoRDEUqRrEUjZBxlVYKCqVDW3eaMvqBXSpGoDtgW2o
6cMkn0nfPV2sy/NkBeZoUgn1Dh1XDeM3U3a6CBBuAkBYV1qXq2vzXmOQpvXtDzKRl6PYisV5p9vx
sE697QywpjdLlqdaprTDHNqu9rcuWoRB6E65HF3WekMoa58eM1DkrnQ7gpQPngnb5357ACpKUjt8
D0ua6lqjv2m3lh0nopMIARPyaNbbnCSVzBGlAcuR0xEjEjiBfl3dQOyLi7Y72LXyPIHzoUD+VIuH
vvNm9Xoi4lzjSkdxBLZeuRZ8eLK6eezcQWkLrMvRgWkw0lNnq3TR/p90ovr62FnCuncCw+42t141
LjSb5fZCI8fmk26FEKKbIRJrP36/EQDfmbzKoZdgumgUbaYfWkO/fcs962AA2cvGu2NxvU6OPir6
ZNREFNq+Kei57Fa9s73bSbkSaeas2k4oIkckHzO1pdKq20Spoi/cWtecjypdkV3awFZG4z4VgeYV
zK4Fiq8t9aimtUII+iOp4vztQFWLEKcTunJNjbL62leucA0ajaH9NooWd+dQWGaBg8WipO/w0ovY
CEe/zfBIvXVMMIKM/TCKCzVXxmGYbkKQrsPMeVWuWtAPWpYSA/7MmovzMEwwLF/WDRC23brvc6Sl
Lt7dhy7/ZDBKb/q+vQsdhDnhcFzQyESuHYzCcexV5xXtpOu74pRI2OEbm94QChe3YB1bbrAw/ePs
AJjDcMINExHunODCBIo99rf1a7BktJ/5h//2N9eM55gYto0ounTGBr1cMYA4OUyMfsljLBclWvL5
V7+9bMacQgxeE3Odz2u3cHKtk/67okoVwcb+H+8/9mgJkqe99AY19JFk+2Zw2JXt0kPnk5Q6Bv0J
5ZcN5Yxa19TG5/ArYwaxBlX4tK6XH5l7SX4qy+69gS8qg93zWTaa3qLcmmBsY4RlQYQFUK4g9Y5Y
NIALNq3KQXEV31UAQV2VMf5qSxhHYGXcyB+Mo6AS3NAGblpWbGdQtIdAW8xB6K6ZruFcml+vDGTY
WwUKsU7OfEENjAcGLwnm1IcMFoo6dDmN9ZtFYWb+zhmbb+AraXdozRsxP89QPz1t/yyrD+HKw76K
7gf/rEg1keeRz1NkpiIpdehBske5RTYnsNxi84hk+1AQAOukJ6cJ3Vjs19qypcdFsDBmpCTRuhbi
DBpeSDltuuYIrEb7jhX6GDNPVx4msRm8KMoxcHoPgw8davdJ2hyH1/1AlNHqyEhepugsuNS5XCQZ
GgdBtepfKSp88Lwyk+lHg3UXw7e6EfYcY9/obrXQhnv5/QLblg0yfEmJ7o4W6FZ4WP8UY495wNmH
RYRWjq6eXErVFQWJpQhYkib73ns/Umn4QwuBI4OQ8W9COC4XSrmc+wQQedmUncwwpfyXZbuObxgs
lzLI6ZsLD26p+ELyu5hoDId5Wwfyua5OqO0rQMI29d9yFkN19fp1440ZaajR5x2RoUTYAQJzJaFh
SvnaqEJEVRGHRK3p1JhW/wfFNdzcID6x1DuMVzbs1mt0e7meEOtgn5Y0eu4YmBkssc72npnMLOyy
EP3uPDlaG7eNXI9tdRkqUuVpxSzgWyxOrWeknWsKgPOkHsj3zVqg8N3p/hoLPYd0CUMOU2KQpzz8
b9j681XjWhtUxEjoyFz0/M2epkUpONJ8WpL+VtMeGdsuCcVCxBDcQlrLkGFyP8o25yHIFTI9LHxa
5gUyl3NCbRTL+wgXE35TWQZ6K79otKdwBlp8kX6TZR8vi33ACRTb+D5fpgFcQ6FUN+9xCY0lVrG3
kMW7ADeBNGwuLHTC+58IkzPib27vDIgiSLYPvAtl5nwMv8CcWTLpdPS7P0M5GfuprMzOtAtpXj/+
Cya2N8eJumevnCFBhOFjZiWwlnLHDOoI53YAAwCz9SuMT1fIaKpmeXiIoukeuwl6mU3RjB4hSSWL
6wWCuUfqTgf3ov389EBWbcu7vOCNAIHsLoj0aU6HbK4G1pYuxIFvErbJROfEHW6vdpVYKT2S4q7x
n/ashJv6nPKI/5+JNmhEKdKzzbUK2YwSBJhgfqtZeSQH6YqsPSFp9fhXdDJuiiqXW/TDrLqjjKDz
tr+Ma1nitLHja8Mw4JRk3NUYZUDk9KhiCgSPikVRu7qh+h2ifnCRslPHlzbyQN+ECOqCyPaBi13y
euTIBNfPwmgLfoB2+geSueOA9GJXtgS5KgZLoIYaCX48yND7vuPDsO9/vSfzrfU4zRcwpCuoS7LP
cZHzWaxfCAHCW4pcx2DOke4ZbIhrd+XuSC9zc+r84jIw9CfmT31Zm2ani2YqAEEo+0sRoSEcJNKt
n4r7PnnK2CvUVRJWttbp2t/kw8hdwJcsuVnWXjWe/rgK84lAh3HVGGnr6SMyYiw5pnoLY51DdpWZ
MlRUBTZs+2WsXSQzZM6AOQnG7tJnXmpSy7u3z66PpHmb8lZUz9HOmyjOoRI46kHB79CdSsNc0T2f
8IYnv6DGaEuIcJaGuT5QFLtDTTgzeVw3vS2XXNMbuzYrZldOyrWYAD63W3t2X1YKY9o/RnGTuby5
mm2jJ28LU3tkWhsgNtyr67vmDRE6CS9xsGIz1Qt4IF96UYRrdUK3A7VsYP0fEapt2AElLhByjT7/
mSmUnE6Y+lEv/AsZRTblrqd2Vmm4JfiSo4vwt7zYaJe1UOYV7gX59am5rm6ICgDhpbgLWwgVrOEN
a9478zf2QT8SrHM3M4wGkSs8jn6Eqqub50MwcKigeVceWN4hDWQItnMoK5NVIeSoU01DYWehTuo9
Fp6ZAwWK0G7P4MHdOAe7c6E8/l47JeEZTvtvXtZlOsKAZFuUD3YPoiDuqZNI3NQrdC+uoe4yUZ02
VxBGmLBk+yZxEvk0icCFq2yuyYv8ne3susouQYae3RdEbYAyrucS8WphXwAmq9kk7v3Z7R7LYDES
hY4cWvqQOetCsRpqOGs5VKd8bMBHrvRWdDxjg0wDTMvarCRWx4ppplxvsIeZGosD5CPD/2SeLR+R
VCxisSqEBbY+F1+zkGGjM+b50Ot/xaU/W+7ba0HTboioUXepzLQb6/LsNbJVUcUBeiBDgEX/5OFr
OuopzzjXCZoI2aViDgeJF87WFTzacvHkhWvlCPpFNXsUvyOd6ZUcOiBVOTvYmD3kHUuwJQN2t/vc
uFoay7xK8pSBcNPli9Bd6UHrtV9xV42RlkIYX+IA4T9+BWZ6jX9qluyjjWaBuMGCec5+9KabxrS7
6yLBnglbxXVnlJrOz+ncrwQl5k8MLNGjFaHDR3qHDsE6MXwKjwG+6lHpK/2VtKDQbEbayNjTu2RM
9Ayt0fm/CQkF0QwWAgUoxcAuXa3gn2rYHW1y4AGKArtlgSLAZuhmdXe4ztHiyFXQg3p5yAjFH/X+
O6pGFP7EiYtYoYJA1WkFITQb+IVHWshv+819vHTyjtpatDZFRcmEhZWGqwRvKxwUVoLLBZ8n9jsu
iABfnb4EybGkbdz5ru6/30jVsM0b/y7teQsPiaYC36OJytX+9l0sO9krUeok6yTo22Uzx2jSjDYK
Bm+ptPNsLsQN0j1WgZlTv7txKLRujFrWKkQXKC+n3KC8vc3GIhAqNH7WE28psZAM1FyvG173PF2I
fFDf5cyh/TntRsA1B1ENGYeDVd3PKtBoiv4bIqfW2eBt4TxdpdmXwX8SdvcxcfY88eSKD7gpsihT
Foi6/xWLgKiNm1YwhORd7+WFUG0hfOdd9UaqVFdbCrrulhPZYq+l1JN6fuYWJRFAA1/iVdAgpzDU
iut+I21BV1GC//iwhsUqQvpxa01sXr+zxC8KcUs6lF8xvtNM2sKXosMScsjAEqzXh7vugyJPKSZd
ltJn1gBQpiA5ULTO1ay8+UrXvTP4zTibtGcNHdvmC7E1pJGc5OauDaFY73TX1bSYjsDvpg+RkVKz
QP7Q/l8LYL0c5omF9Gy9nZZjo06emwd357/QJXCQ0BrUGkBt4Nm9drjsJZN8KeO8BV9kbWTE8izM
1JZcOATfL8AIlgpxlqIU2O/Tq0Irg/R261xHyRflgSKzw6ksyIDhV2DvISqEylviXkjyEoNCyGzS
GdZKyntspYyBAelOn/iDqQ8lu+qZf31VnNdlo1suu04UxbnQmDUQhZGa6pQc37+uh01UWtCwByvr
hc+NTXypLhD6aMOjq8DLDcxsvi4a9fdfiZyphvNwoR5Y17ar2DBpvNuh4UVcM/8CWoM6K25SJAQD
fsY/CDuHY1bIoAzeMjWSWeX0x6x5UlnGliZ/HOw2FoSr41qhT/fF87T/2zfsA/QUNpqswCDLELF+
I4nu1iId7kDXkLG6YdeC6thEahFB2YHg7B1D6a47y9A38Sw/T03WBl5UTLsvQkVw+0aIafm0kWe1
Bp+laEpjmV3EhAp7sn+NFg5fgfqcjDMaG28514xEJS1oSYjIU0d2LKYzteVFwO3Czyq67y9hD87L
lIu0fVjIzR/wk5eB9/VnTX9pBkUtkdqNxHElh9ZTR68bfmttLvBAbkc1g4+hAmoAz93YsA1V1BmI
sg+SuWkskTVWMfBrGn3cdOWcecfdfZeG7l5E3IP3a5CNdWLysRduHDPx8zE0pAI/ZX3TdSCNrNkD
ahHdfihInJoZLJcQfbQbjuOCWZDy3mtgUZP0rdPA4vH+f66Rac9h3S6qEaKlQ55CsLrmZuEwkGaq
2xFVDF17ioeiDak7eKg8hZjUhF9GFaXVeTMz+0wzNVQlGFiCvXEnTJmcOzK7oUXq+9kLn9fPwShd
9OKW4Nl80jfHkgpA/qONhbp7ExUArALlAoaAiwnKx/AjZY7UCeGaRsnJ1QLFfI8qGNEJed/7F+bS
MBgaHZ783rHpC4w/vTWCdlHARcWsh7fxOoGlvBuWaAV4yRs6gyfB17xvnkUTmvNZI1qL/LEd5Qjf
7nqgcb59864R7J0r+I+qz41A34eqSmRJhUNF8fVx4paG9Mi205Jzlurkbc++PbWootvjJO6OUvPZ
mBFm5CdKNOdLtpi/ayOwdqRzS4h7/oih5GgMgv2RzI46wv+vHcbVN8BGOD93HBU+JDKDYxWd1jXn
qHLNGty4Gza+m19W9VJ6+EVt/U2wDij0s1UeJPRd0lSGZKgNe+YIaLf2jFj20LLpi2JYwvl7zhY5
RYsVD6HIQH2V05LMkIEvN68LbTf+CEp7ifPXh95ixyCjpJca+um8grhAuQ1tuNkrHp8dBufC2lOT
r61/eoxP4AOK97F65lUWCnJn+7r4IDnCkieyCXgSjkCFyyBnsX5bQX6CT6JjfTdaZraN3xusx5Gm
97TST+AFq35hdYG2P4ZeO7ttw55ekl7sLWQZ8Q6ye1MeYiYhwS1hb1wDk++NQyV+I2YsrUyPeugd
aKa5qUkG2ar3yq2UQfmuSXiJxABPvSPqv+MNO25luZSjf3NFG9umOQhNSwEVyseEHRy2SkfDkEVZ
8gYB8QBQLycu2sKibkAPIP5x1bn1raBQ03Fcy5lj7cn1Q90Rb2plJrV8a8atGPYZ7UsuOWZSBL//
7ydjPuRcS4yOfBpXk1Tf5zOb6YLWAtClS2nCjOWZtuzc+sxe7o8apPT0pwE1tI6ToX5sJ8xw+/bT
KnXTpstU4URNLPv9/CB7ctg/9hyTSKViILhNGSlhQHKODSSLeZ/nPBynCFqx23QsDAu8hSdP2YBf
X1ofGbVBBK63QSE7hcS6dsbq3peXCbd80+Gp2dfuiWhS+kq6Xfyx97P/5Zb+knvYeSusz/LXmlK/
H+e6mqssExQxgOfXl/o9JXMPRoEjWfjVVN+M6YOr0bCqh++Q+0JlIkSMqoyGRyTp1NlCy1Htkpwr
MZzW2QN/hBtVH3m4A+KqfRbYRzkxjXkHR1nDdLXePo45MY5S+BCDmTlAqABGJRs055PcGBlQkFhP
o0D04liMHPINr7m2FYLmMeu9Dh9y3xGWAyzkOlOBERGpP8m0KGwmg2GWEzx9F6Ad+oG+t47ZFNEO
jpsetcl3iBUOqUoaGUmL43DQJ1t9ruL5McDYYmy4GbJNtzPgPVp2b7am/RO6bk/jDso5lY1WLmNc
2XN4iQdBW+x0jASzXophiievPcKpqS4PHBhY5saQAXbRHWIrhqZidZIxEIfNEE8ecrOMi3HlpUfH
cQrh+AR+Wn51OkFXHEGNF8sdDzXkuC/BI5wXWLCuad5SmenEt07gKy8ziziVkkIwiWNgKfrOA2rh
TVq+TbN4Fg9vf+R3t0Bgo1IGR989PJXj2YbzHzvTXf+ZPK4NMwKhQPvJAzz8uitwaryxVV41/ELm
23UIjHzoK9AlBW7LCrKDW23z3XmWeFqbFrcytk7BudkdVuM0FiSjsR/pD45xMulY4ft+Z14fn1p8
s+YkWtwsy8YrB4lOPni/ilYblLS5OdHFw5GOqldY+l/FumQv57BRdsCM7Odbve7wbS2kwkRScQIj
x5lYQkZzG4bfFAX6t6xUss6cY2zdl4yW01W1QqGc3in9KNM6bwQFmDBL316Ph7erw1DEgdnNhZZ2
JmYq7hN1fvnRMVCnpE3IMnpOCLBoaWQoJyUXwnyKX83Dv7xcQZ33RQ/i3vi+s8j3Pz1rdlDjDf0x
0297F0ah2QNdIzp6RpGeutvGvy08Xf9yYiwIDsaw/rjq/UZVPcbqZkUMg2LJ5slQUUzSn4u+uaj5
55Gm6tT9AZTwBVR51c6pc8nqUKmGxfA2D/YBU3TftEk8Gdu8DNCLNSJDsl0+crCNFTqXpAkPSciM
1DASSwCUtmyJuHk4iRp3suj6Vf9ilVnuqLmzmZRHMoCh16SJfJ1gSy20EUovngVJPEzMHJHQ0B72
5K8wVHi2uC4n55SET6ohHThrKta0dgX6aW2NEsxDPUKPzyMk3rbBt/rC+3+OiVWJGXkMidvCfEnG
HqQYFbzNAFKNWgXlBsTJA3gkh5MKwZSpTazUReBgSVUTUUBXj+6XYSZTh31odwNT80MyoCAYm1lt
4A9yhFTRxc/qDYDTpyZS/n3Bcwh4l0hHim6fP1MTd7xvkigPab3mXQa2t+ih8I4WaST9mlFc8CNQ
lWZMv6lBzve5dTi9orup0IfepgEGgAHnjHMMwcZoBCHov9Tkq3xRRU4DDKlx3bdbC3sAhdkg23jp
U6vEz5pjGRBKnv7oQS+v0EnWKz+XAqg4Yr5pIpKUFU2LTovkGRs06PHTcw2Bpd4etZpFxnyXtGMD
nsUW3ReCrqQYLZiZp83tQRSileum6q2YDkL9ofUeiapGQ4qW5beddJQGd3azuFuId3PKT+mlMMjc
BvsEr+xNj/BvGJO12jrkHvoM2XwoA/rUNRv9H2JBvdJSWC4DvEqAN34heEZJ8vlDrXRIltmTEuxC
U7rVQQyzcDL8umKh9sMF9fUbt8m/t/vF9kVC2ljtCc9L9Hh9oHEuP9oafKOGe06AgdS+EIGl5zCI
gYnyrIDoLcsels0+tLFuj9NM1iZSdCpqJRyMsi2JheMfjH8M8B/66VgRkHXnuqTLFmz8/7gszjNd
1Wob1vQWvCkYVyvUR6Z80zM2XyhFX3HW76SUJKHos4YPkfUQNyupF/q9nIFsV0C6znstRqYcne9H
pkiFqIGaaC3kTK/sTnq3u4yyotGX2PYebQHzwKEGpvurtoQFDrKbqqHe65Za+6Zz7HIF+cIlOA/Q
lo50iMQfbElFNH7VGafZ7Up8nbWqe3ncZtjZNR0SxwTo8V9cn5oplOMuau+NNMs0/CWFthlI/kTq
EkVGviMI73THYXaUQ8W+CiBPDwiXUG8VWWO0SM2xir4uABY8q7ewJtvg71pyLDMBPLqzagPW0jYX
W8g1Akd/C5Gy4L7Dd9IVkafO8kKazbGf3827akn5SYp8UExrvRmeV4FRRXrXx269iLpY16xcHdH7
TVvSQs9VuaOuGf2cUPaZ5sanFOdEQVeL1Y8jvuq3enM3QPVO/0QsyMXIeFkjBPhdakF90gi312ah
yECHoH4VtwIs7MrEyQMlklDsJxJdBnNEDaUXaSja4ucEdxnkT/af7094s1FYUkDAKAwwhN4vnkt3
n+9Bq7yFeW34XFTU9yejvJcshrXlzzUyMs9n4Dfqc2hDquczzeWaEdnmo3e5GznABbF6L2YrStIU
z6O3jS1178Xc3IlvBhmkztNsO7XLXHiLwU3XHXcg5kUtUCCIUnnsgYVU9qbTxCTP2F/2lfeM0IDE
Uw6kqQcS073vBiaBljC/62AQCPl+4abHTP+aEEiZKDbzzquUMgiRLOXsb/oX1BbZgoItmc0BBDBP
3a2dO/NxNd9d2V9qSgdmYvYxpHm72AeR7CK3CtKDWAUkROJrzFblQf5N+9Ic8HpvUL9TiwKYfmv3
vnxnqy+sQyektD4z/90bGr/CE8KwJJaGmxiI1jxj+B3smyYKpBzzA6e51N+sUfAJtYJ0NpTsKYnG
WlzbO8YJPgd1CMlIAErcCS68RwQ5f15Ssb3sMW1rqARetMoQXEWBrHYdJ1S1epz5H0TFPEQoqyrD
EIYoYtx3I7ww80hsSQAtVrfMZdWfCo8z79h8wkV+gX+dWKXp3y1ncdhU3ZVL7YRyjvg2bPu1Z7R4
iUJ9/qm7+nN64s08oeN6K3R8mLksjx2bcxkElLaojcdOGNITbxgAfX9rJLZuYF86ZAG9xcn1j94/
ZoqTGdIZFL1Oowgpzk47HNT70padf2RbptZsYmnROOQhqyG8ru9SaeUbIXqRMI+67l9lxzwcpQkr
Q1dh1nGSST2rxmIjIcmZSyp5N7vfd+T0lr+/mD2FPn745ykut+xWYP89I93/0TSns6bhkNhit87D
33o7oWQbpnjzb0b8PbYH4+wQQoXMgAdRs0kUXRkSHUUbZbMPPDLtlngJtfsoydIcHWqj+TwoblQe
CEEhFaebYOe5fNrTYz8kZs9erCR4kheqYBk35NVckez7OzcZq4gwJd7Oi3Bsl7ucpeuCNM6yl/jl
CvOtpsZrQ9/5XJp95Yw6n8oVZCuDAfhbHVNBHg1DCFEn6y+tdK9ldv+WIu1qWy1xvz76rCMISlT5
8AOoNwdlZ9xEjrM3Mo8kM4nk8Jz81+SpEvoCOl8wMyLmS8Gjkk1fFe6UqeRb+QSqV9bQCOMi+m4f
+dq6mq4XxiZxfLSqlUzMoc4f6OAHYjVgM8OGALB5FVc0/FtZFk3xR3Wd00Kx8Ak1Nh5naFXIgpOb
P1AQVmLnE82p4KBW3wG6meRydTTPrPYoxj4yIQPDy0m4VpN6JtrZRsCtULpV8b1MOzopJYnBYr8w
4UtzlIsGKgZi2fdMkKD6NAYONoSXdZSKcXb34Cuo2XrCZ7j5PX3dqYxAfsKQS4SEhM2y2xVDoBT6
P+/Um780Tr5oJoN6jsG9jeTeEfkMfKxgP9TS2KZqkT6ZJVLz+0dIOfCA69dxh69S976Np6jMktMP
UG/3xQdrPpHOiiayR107v5PQsWaHB1k70faSvIhn8FExk+HuxSUsbfw4inBanrC9sIpu6lgUScQ8
GQSpuFQJ7Jair9bGjOM06N+nYhcZmZUE8D9ocJAegfSTWr3ccGxbqLgaMimUr0CpG8Gp1KzEGLlW
3cw=
`protect end_protected
