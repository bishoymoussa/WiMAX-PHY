-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
s9SzKyMRF5NkRvrpmzcHGmS8fiBghchTRCexQxZXGLwSNTjUsaNVkzQrjlVU6zDHzsibmlZT+kGX
Rnoe3mBarIR0jSRScltrDrJ4Gi/joW8ehswgBrABb98GIwpvRuJJ+ZtGnTzwzSBnIihbP+ih8bST
oWi8zCZccjuqE56XPYCMEQPK8xUe/FuvXDi2Kfks6G/QRrB/XbTFrGGTQCchtuP7XLW1U+HMHBiV
Ag3ed32co9UbbMroff0X6K2DbUyJAmzvSF4GU+8en1I9SJo78B9V+eq3WJ+IBgEUqG5sSKsbqVV1
Ql/1OTsPPbYTogUipkOiYZiLV1qPOyg4OmWHTQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 90624)
`protect data_block
bqPpxJjDlgJ+YqytLq4YMOwWMHYPfOVj5XQYhQiQH9TEZrCB+qZbUGwVLXzwVHoSH3+pU9sYCyTw
nyPRtZR7/5Bv0QPVj3MwInRk9xur/4ObPDnDME5E34/RuLL8qwsrguTctSoF/ZVfAtr808LkDk+Q
4VfSZayKxZWgcmiLk8Ln2TP1qZOafFzONbei2hQx/kKW089O21mGA/nlEsWMVFYvT8138JcsUtai
LN9tJaD/sguNUUM7m4HarzNcjGH74Kja7Qdc9DN/ArGIIs9qBXIsf9sauaoPBW81rle9gZqigTOf
1U7KPa/VpJkLJufMk2/NCrxeQIZQg70ET/Y1uFawou3iBU2c7XhdRURDym6w66Y8BB35LCPovzWy
T0PSJkkgFjfakrK5XO2rV06mbJPgOXcPtOu2gJQIfi93jpgnpSRisUYRVAEDuREelOz7Zhntpaw9
VZ4ZUAxGcNNM7kYhRCu98vKAFgpxs6HSyNWYemWKbNdX7vWAtf5tFTZZ/pt3wjuIM+zmboK/IQng
oTQ72c13Wy82fRNWIEQG97lNA7bGtxzsHG1GV+/Ocka/Pz/jnpgsnVbcj9OoEwaVvBZ648m2MNR7
j83rzfmLpxrEGVpBuqvz86lAFvkw20Gin/kIM9QpZyMLMA4+hs+UXqjKunebfBf6Cte5P+dXm6NL
xDzWs5ycZSih8jTNvrK6tcekMRhnUkujVkc9S2IxSolK2PpOgy5N0thXJIVK9ytBc4FjXGUkaZxd
oohW6PV4qobNgcJ2a8vB36UpJqj7cMzq4sbqSWocrAitlEoPgSyGW1QuDhOyoa355IMlLvwz7pEk
PavZUDmR/Dul3df+pbly1rRyXfCFSRIsLMKvodf3nduoO1O0s0sxLI4WF6WmMa2VXTjyPwXaq/xv
ikY29nNa4b5iMmLIAH2eGM6gH1Jh12NJrgV9LGP0xtcpxfTXyx0fN40r9e+pARGzUjsdAqDF63sL
eAG5WjMtrZ/25L8d0o3bUveNZ55Czd3ksfU2egRMQBQZA0BOCaqTZfmbHRMS/ZC3vicB1IWRpjPB
0ST/CUpK6qV7kBLmjRy5/TQ4DyWeIP1NSSuQmlgfmPIZMK7GtVu7P3UDZS4Qid38LrIJyvPBP31/
b6Mb/AYgNNwF5fUideU8KcXY3+i9MGtIA2ufyPK9jC/YtUQgHbSoLUHW7X0SqIeml8XF+HqZQEw/
13Psqs9d4sQhFh7BzwKrHrY6bEN4xWpgO4rl3z9L6Yzi8V9Pwy4VCLiaKshnzN+g+74azy3KnSz2
DR8TdrFJZakQ8+xuUNNQJAqFQEvUj53dZIf6KTmP4SftjACSSUWiXphriZEkzzVXIoxJ+5Et0y73
zsUAjvYx1Nab99dV45YDJjBgWaxEL7oBuB3fuyxNQNQKFjZSglUTvp7qiNLQgZQG7eBbXd8/hBbg
gQltNBsURxST2cS2DaDwX0ZDht4xLyPHWKnz/VSqyXzGa7XxMw5VQliJ95r6sHNpyeWpyU+auRA6
FlKGi9cyRxYC1MIEFq4qvFIMte09PH7DFz5LqZXps98xqsJ3llYgL8fD+nohlh4gBHxxMHVXmzAk
zIRAxagkFW/fpeQA+Y+j5j0AUYALvc0aLpfFdQHD887M6E6XmKq9FImmi0Zwg7ylVQPZUsInxcOw
2PV/XxF7wt52WAITvH3U1k0CkU6Fj2Cn21xw7tiZRJJpP7e+yZnJElwCuwnK3nuGHsGyEGEeE7ZO
dX58kza9hWbbzqiPeqoOTbCo0hT114hjOBeHWXUggarTCSpsE5OEK0LYY0Kmd2qNmdAj6/XmUAyh
ntLTrP0COLOCwyksqcP8rHPZditB6aOUbVxF6qZ3HFZDP6za6+gLDP0O7E7IT3Ar6kYU7boet/aW
yV9xlS8LDN6WiM8YYn3I7/YvRv+SvLv4YaSE/hz7DRzKRMQumDclRDFCTLZu1K113x5WqJxB2jZi
2pL25KVx96hYEhUIXMvr2aVwbuHXDkm0xnQFMi0qtGJFjjYAxxgGUy5x56E93yxSrrMq1UhQEsKt
H6aHZcbENgUu55RBEKIiuMGqhc0ehPj+8czsk+q0jkPDX2oO49T2HGp5yQPXKx1ZEtQ3gFn/1LqS
a3n0aIG9x3ZzMhp67R3g9shnelIuFWoqSCnebNeYrOiauCK94qLsoFDyo4RppaOzVfIO9/TXluru
q561vR4uS6Df4xIVIrVOtmtfgCZvyfdTxT5sf0gi9fAdOKlTbdln7qzE+zVFAgiEWLCDoK33ivNF
F9dzJhuAcGkBy6JTUGjkLOD19jayiL5UzbtKqkZSGVoVLPu4s3GJc6DU9MdhtGkaLfAx4+Rtfrb8
MhdNvZPZi6DPmDcz5kpCm1zH44GKRt4QFX6POteH75Bgq9ndDMmYcVj/RUhhyto5B7cCp9N21okG
6msIsiVRi7dq28OAfl4x7pnx3jbkOIHobv1umxZpnAOER0w1fhbgDPcSZ762GkyWB4oMCYQqKWKB
IMcuC/27FpaoKEYBNOP78eXyW5WpI5N91Wt5DmnxR6mW3NOppHj2IlHBrRvVrxK9qlzT2hH7ximA
rGZQ210XeSmk+cU1xlVm36/wECIzeXqYVIaZyc8In60X2mKs8Zd/eBpbiE7fhIkQUcZJvqI6pZQD
6rfXPyfZahNp86FrOP1JARxt0j8/XzIu9NoNa2YKCRJ95sfcYWdloSJozt7G7fvi6yAHXhqooNJV
CZGQFiG405TRO8jDa7adIvEnvUfgHDhXNRnXQnTSiIRpCIDaaRyk9Tx8VaYNSi4l9/j02B0frm9K
OlUSGLXMzLz8QnUmgHOY32JoJeRo0tJyMI0vP1U+pzJC7JlHLyd+yYXnuhA0TJuwkStKsdoxLgoY
3I5n9Y/hwSDXnaRSE2M7tLHVm1wOBZNch6jTYdprq+yhL6LNMfUWrNaDUPZXthFopcN4iVyqAwWM
ewLqytD1XDPGxGz/rS4dOpQoqTQ9VQVEnmbnps60SPs6vY4kvYbNpdgxo4guQrR5RdjaYDjqMgfd
vGP9wQDucBxXEB6iE5rNrx5698vCss6VFaamQiu0t3Df9ZLjkbK3SNAxmO8IE0E0uZ126Td42/xE
pbLxWESmpW/HPTQGP/j5Kag8R06Mxchzw/+ojE75j6W/5nC/+5h8soso8L+YceRna41tSuM75A7B
fIuzP6aD29p+AqCpslVx0hehlNywje9lr+fIJ9o9ja1uuZkzpNFP3+nJkBoJmCpC1c+4JsAkM6vs
f+NHzL1fU8VToLUbqdUz3zEB69o0RAHJGUygyxoTxh77WkDFWGBaPs+qWF/vcFSegViuniaKlszV
Ty0uhRmeIxRf7KtxxgfYYvtL5X24o9ehgc5xCbQaJPhAkC43YUBP+vsUv0tfTFal0bJaSXdDzvmg
rOy9BDEFUmFpbzsvWd1f6eESg+onExFDDGCHv9Q//45R7LF99EtSB3Z56TgQdVq7hkOvsnrgC0dn
AA0r/wWbM7/dHcyA0EzUWlFOG8woLpcpqbILrlcbBAxBLfyFpfCOtYyCf6htaYm26xiXzi7EAjFg
egsBQN9DKzEQfSZcMV2H6kneDuRrjpNElqNDuTpmvfGBEJCYBTLKhoovPAPSMkBvNmJl32DKtxFr
I/CyH3lHMkuj+dpcUVyuz6bARkIgDyeHpq5WIrWWMvAB9f11dBwDibD86JtR55gu/NUkUAm4GPol
UU1dqXsG93DClVf2lthM8JDZ9iZjFKS/3Jex2RhOL3xPHAp/+4o3m9vWOKTy0GEHTJPIfUhyyMgX
P6KZmRfmJDPhNlCWGxMdLq9Ry6frV8ljB5kRgnpMyhf/0FQ5Um6gRfIXvceC9j761q8o12eSzDvq
MhQU0Jek1piD0Q0d5VNf2xSnMJqmT95xj7lyfihaGml2ExWu2NTdWdcUjFxduJAekB+LkYiKPPhJ
F+n2aVTC5snqnmnTBSGT9FwBmnEaH3t4RCSa175kiET3LCRDh4TlpSprLbuUJYAhNVcFUKaRLpW9
ALagu+vM5U3cpdvGcJb/1dMycJJRTfhiRJT0PnKEXGNmwV/YbbZivClPY9vzXPpPyGO7OwTvQfwa
gO6N0oYeanw5sRUKvpIPcJYJH6gFuGHWaAmE79NIqydCWmYOApiP0x75XhBmeDxAacQ/dTEW9Wbw
pcsJPDTycOQgdBCJN5opyX9HBZi0ZbNlsOAOTPczN4IVZyebLub4Cl3de9rTu1tnBiEuu/Ap86KA
h7bjCxEE2nFMWaAsPfdRusTf5uLXGaMGWh+WEO2SvV9G9VCjGU7VF0ex+pKOD0KUj3vo0ZJkkT6X
4ICSVeh1TkEGTpJh10uXKJ9fADV9VFOhFoBLlOj3h9BsnngHsVt9Lcf2cylKnNzdhMF0zXxgnBYR
v5oo4axf25o8ExNUPBhdhaA80QgxClF55iSwwupk/FAnt7mQlBC804l96xgY/E7bYh2b01Ggw82l
C8hf8r7PAEbnVofmOQGs+CjcmHa8GHuMeiolkSb/U+v2Kv1yTY7s8Z8c9jBDEer9dheR0nWelvKe
yd5Oro3Vill45TC76CSkmwuiG3jENitRx6NNJBnW6BSbuNKtiTexVKp79wu3loVGkYB3mqtbwsSY
NznM7p23gTLiNEUznKobvhnGY6s1e9YGtflgQA6IzGXAoazCl5TsWJFIcCJzg8nqkoy4CXEaosh7
bRGP4PDVV6jNn4NmNSDojNxYq+emN1KGywWzkkiLafssV/Xys5TO4O1kIgUbnIeyA8O4GQc3gIDL
THnomocCJQDZJ+HioB5zPbHKZW+/jr7HI4xPMEmMGaliHGPZBDa02j35JSE5cdT98Ngvz4AJD90w
wXnOwRLaIA/7xHwhRZDemaJV5hhSImfc4tU6UX7gPJLwUeD2aMBmf9sXHFvgi1DDiN/syMrPIcNI
pdz8yyg/wrj5FV3jufk0OFcYB3DlhAM81vjtkGzyceq9EErqzwA9ScaMv3/rCeHzEQFqTq6t1e7J
HyKXy/uAilmuQOFl2l0UpcTKGoI/iJTiiGP18QGe9mLW2f5oArmXm5BOeXgC+e2SVmL2Y89a6q+C
X2BFQq3zGw5pR1r2i76ocCiBBW2aK+aojrfHppxLoQLtmM+F+Qdaaa5h67TsZRzJQBN1q9Yc9bhn
2ESgL/7A1awiw7MjDOD2tesLgXXuDcEP6YGch4RDqy4VLgfUUl3kWesgblr3txvp3NGx7e7z2xSd
8s0EuI2gasEqb/mAKphtSHRaumeQJzPyhuo7u5PJSUB2EuDIRSZlh3lXKimMgdemgZ6TJSEisaz4
CKprBeUz6XT2Wfd02kdHD8etUUp0oSnzMXSPv9px5sODd3yHrDLLSJHyjyDIKl/4WuSLQx/PNHsu
BMZlFHvddT8xQu9+2NwTO/bDNB6C/RuHY6L3fzw6nIya3mvBjbwSbo9Om6BXnFu5bkNaVuIw5sEf
hX+4ah00fSBysb10Xq+AP5S//bGwzcpfR4+9WDDu4LDunuUiCHNbr4D4+MkIZW+ufzFt/nI19OGB
WzYnqB+1KkRSWgvmLnZH8D3qP+t/Nb7OeLG7kuNRpfBAl65GEnbfVJBnYZMb9ySiLWg/9XmBWdqd
TieCSFkUbSWVOGHrtbl0plwCqkCQdftHBRkkQn1lG6uqTAB/y/6hq1YxV4PQvVibB5835H3H01E6
qw+fvY7x277dEPfyB/E2bLjVlxPCNR4eLHDAMwgNS+KqZkdMvmQYcGJcF/IfkmSyPW02PiDTZvmC
5Qtz680cjKlcd6nwFatvIKAcODaKYDRKWZHyp/P6Hf4U7R6nKuXLLlaZhv7dvl2sskuyHIHfbO1p
wrjR2YZBrvEhLRe05FRvbaGiB+ivt/23nS5AXgWsSCGBB14yK4IK1yHPcB4hEPSdpu/8HfJjjUBX
vEa4YosAVg28xE0dozrIv1brQnVuiWVIN3ne8UtfhA76aeulw/+eOOX4jLw0USGRnmvOkwtXyhJp
tbFC+udpLU5swzMpRaxXQhFJVQzhgnuUKV1QQ7ZgiFhI+Nc51cb1zGm3W6b9E7bVvVoqwCALPiCv
WRdx16OT6ASK4ugjDDhQekN4vBghyUlY/hD8OMafxgztmh0VZaAaC4ezJ2zAEF4qrzoqXn3wbx5n
n+tG9ljCqz6XGf/4c5tNS7yfPnxo8msjPFx+/y+hccTwOWuebZmZ9Wdfh5sB9+hUe7p5nAEl3Bxe
vqZUvGW25HKlmUixDwlyuqSlb4+VgjSLdAA9PiixJ88vLeQW2MHeG/99TG6TYCLzUE0JDHdCMBFg
0a7h7YQkQy8HRW+7mGhQxCN9fPXUmab3TAq89CCramyXEsMwxLkZu66e8sIkKV3aSS9KTbEeKCaL
X5u40P8qQphH1SJ+X+5fB/PDZdeYlTup2yP5nF5vsdRFlgn6w/Ivi/rAlEJbFay2DpB5XO48nfjt
TnPmIclBzg5c1BTEVqsSlVm+FBsfi+OCc0q0yHWP1X8hPv2Ze8PAwYR54rG1kcLCpWd1I+La2Mfw
ULGt9Emo09E/99/Y+RslWulheIt+5SB/YEbozLXxfa8rZrIr+kva7UyrfVL0pVwDPVSSEjoD8mr3
TWx/JIZSdrVCvYBpDs/yOuDBhaR3qCuiNfywuqTjnZQT3/Mrm2eX7U4phx5FvXKMfBPLTN7qLSYs
rdHQXIy9jHqnI3sqOc2vyhfLRtwyoIwfrUSroKkNx//DTgwEC9swG+GG0nQfOYB/H34qb4uO9k+d
PdYuzuG1iwEzNgLC8ao7eiNPPjaBHlA8Hf+T+4pPg9OZJEXqOR5Qz9IOIVaDxzEZKrLi6x2WKfZ1
T1qPHgUkroO52jbPiQlclmd5AWyw60kRqEOK9Sgnb9rmiCWvYmsz2PIfLp7UjPnoqM22kE1bI/BF
nmC7yLHAcSHlN+fgfOkbPG40PNV88BW0YoxdYtsmQWXemvMlrSTt2h52j0fefF9DJrSgfmB0PNO3
AaF4rUfKONWLLFg4GZN6MD5pkqjqdg8JNDRfp/k6m2/yp5z3Rc1t40G45MZ9/jkgw/xADnGODZjT
rKhbJ3qB/lbd5uhEDwwuYScDuTMLCifmSxlozps6bShWxXwZUtoWfd2oQWnJoMptfy3PZRPX69cR
tSZItCoGCzRsGkRTU2pAs4YdeaJ9pMOndjc3qcnoJHuUc9qco8c0T1rUk/ipK7T6352X9rhC5fFQ
gROZ3yVWD0svmIvvn+3zu9R1iUTuGC5kamwiJLdEEcbO9hDAT7kReoBfvAu6WrqXGOUQ3WFgDFFP
hlyroxJCxMufnC2He2sYTfWHUQbq7PuRFkA0DEcBgZPKEi3Ae9/7mdVE149lwHkIm8Ku8zvuCUbq
Ac8Ze+kNLCYk5u61fQY2K0bYMytoAvzSWlfSYPa3BSLtt23GfEbPKrxewz+ih6yQAyfXg14PModq
IG/vCnGAhqjfwTMHiJBq8VebIYtfyo4ShIsSykdehP9OhVYhbyX1T0AvTRf0c+q1Ag7DUmC4OaHw
4NUO39RfVP+U0beYmMvTrdta7jheGlIghi3EKgCR6hm3mxNgOdaDwifrzqISS3VfgZ5nJlfQ/Lk9
SC1e7KhDT5U6UjIBGualHa1SLS9EaydG70B0G8ZejtfiXSCQnlmWwtZlySdQdvGLTRG7397gIHVG
oj7lnWcFaNeHbrskGsQ/QvZM8pV3+m82LaSh9jU54j36P6hJpO5cDVuKL3DaX+hr6yaxx1PNzqsQ
uzkiDwNHPIXBhnw7IyCuqSshTFRQyDSto7NF7NRThHrr+6yqUhWzMczOLiM4if8HrR4y57reNl3K
iK9U9VLdPzwSlJij44So5zoahAKCdwjBT/GpmBt8tB551d88DfI1mhAgLcisJ7TOoqi019isFGji
npEMZc7UzwurxUIs079LyPo+6VLLj3Jg9LI6jZs92/YicW3O4iDJtgagXWGn/lUl1XopWNqJG1Vi
h+Tf/EOQh3P7HCL1+268HehMpZC++8QYsDMbCLlMNsFlOlo12sufnuHOBAFgR5Rum1qSez7U3B7A
Momp3FRgrn1OV3RfbV3EHV/M3EYedbj4BLwfHUr+JVSsXSTez54KqqqHIhYrhGSsgTpm+SKnpcc3
/O6WgRuCC+SRI9bpCpu2sj9a+lgPdgo3vWMzg9XjWZyFnpuHfexfc6c7w5dYGnECHOBY55gRwxwJ
aFlFZ/zbomgSLgdqnJQrfdT5L1BOH3vs5Mj1E+LQH13aGotGBMCIKD3w+XzjBTF7lLLZq1V9GzYD
chEznEu95MhqW1oEvA5ReRG2KHLzGSRDWqwRoMZc2uvP0GbWayOqmv10adiu8Lv/aMJ8TPe+wt+8
nRrwc3ixbso4kVCcaewLA4laJy8jaIHIHHErCu+M3WrPqwVD1l5RFpdTp7UDXk3kVbarFtdvWm8H
rnaQ6bc10BHWr6W1to/f5/IHK4pjjQvfQ/vzDsyB00NVDtFtI9es7cPFXW3wDn3KaBvefMuHW84+
8ltljOmeWwdw5Zb55YXPivCq9MGeuNzU3+ox5C7fhjkxsIaXu+7/JZgJ2igUlfeLEOLiFPA5gpdH
8UX+FZnhIk5WA5KA8Bm9vgtyLqhFsrwELuiFJrTdK0+0gnDdqL2RsgT5JR9CIvU72jKY780SaZnE
UOcQSafIbTvz5OPrWL3CJNaEqmnNL8w9Xs0rfhqDDthEkAWnx9i4w2ayPFQUvefKFd806yjtAd1B
yxlRM2bATFfJiW57+8bVYRTX99C4+HgGzdwfeIeBVpGi2ElDCT6TvRtgXx/ICq3uG8IaFspT20zp
2OBgHnz8+e2TiAR5+xfgrOxIZYQXtK9xUcWYe6zT6uRVsBhZenNxmBL1lxSUIigIl3P95pBFum9s
gTPMqLqOiY9I3SWJdKfJWyMBnznFusq4Ed1+7iT160ehWweKX2sNHNSLIJO0HeYL9rEzuu4+PIpe
EmIegejUsIwau3p/OnhxlVTW4Kr1oZpk6qUq0N+ffooaiw3WOwwCY0ZadkYKQfZ0U9eAAj5p/ouu
hOtiJkwL2d4cpqpmENozgGbQfcZKBLTWYzEZcytaz+cHQvyucbMxZXeaN/14ciHZ/l7f7ldpk0DB
l4HtIsxLBJyIwRw50h0q4HIH5sJureaU9V6s0tqcPW5841VYgy7UxIcVjeztQGD3E6w8oywfCq6I
qF7DTJRa/Fi2AKBTnqRqSB5qKyxBVLIrgcpJDXbh1uK4zpOsFySgAL2jXILSAOOMeg/DXxs4yMI2
/QoWhA9TRqCcEVvQ2tibiYZirOLj28fnalqfH3q5yTm2k19rNSGBeaIkrtVrERv+d8t+5uagKxvU
v+c3QRKTzG8wEdVgrfW/aqeUl/lHKXpMW4CCvqkeF+5EcfVRN4jYVYAYyT1pA4516wLo1feaxk6P
DRWR/DUIkXQQbpjGOJYECf8EldvnzRUiGFqlQ1W1/D5DuB96UEFuHHBhOWHSqBJoiUfA6LaUyaA6
jwT2PptwjbSpba/uHgn53rTA/iBZ1BR9iMzM4RvKcREelf3Ff9NIWhmCUX1a5IE0bH9OF7niWEHP
wsir1M+7STA9/j9PwyIafQAC4/7ZO+6+ySFn+MkgoZbMgkQZyG3Rte8jK9w26Uuy+jiI9aV6J92t
NkCCj7V/fhh1ifCipY41TdA6wQEZsQHilx4kvJxZAs5KS1coXfanPlWeKwbc/SN7K4NQMAND6wqu
9jG6Y62GVfzWtXgYecui/JYaKDbb3pxICLckALNierRk/7aiZkWUVhluT1ZEnO+aJpd2v3C5oi6Z
7+LQHSbxLaKWclfWyck/c/d4dNAgGZe4j1Z4626biV86VNjXt6cSfJrK9wroJkQlAIWG97g+ZDLN
+X48W2bHbT3+LtvK3LSarwTzoyIYkVt3bzAqihvhK1WbeeSpjuUqmZ4lY+56dllRYEElJ86gmH+T
3Txul1zRRtfIfVymr3II4itQ66gHuTvETQLsYsPHTTAIDb8rSA/O3Vls3+8eGapWOqCNr158ZLuX
s8e5jStEydnkVms8KJQ8R0b97pYORwD5FZBg3OPo8gVubGr3947l1tsrRw4yVP5oWOaHfI1/FrsP
ZBIxsl/S8niuB3DHV7dPERrVDRWW1FyPEc0BU0DGfl44ikTipF2654GA3YjamGp5SFkrZkoMT3Lz
PezGlloPPRpMzVaeGSS4NfC0Xrjc1o3TBLBm3OkjJ95GzJLdu31zh6EYATY8vKoPCb4Y+qyUjTpR
CacqA9dmvm53/0En6Z/ZIZGXbZk30E3i/NFCCMlrQ7qKnS2HKSYqkDDllqjVErS2cgnifMBUa8Df
yt3r1HXLYAiLGpvl6r2QM1Idu44m2HYrwEMQBijdWt8sULXebesPFexC7Bokxt6rbdq3i+aL5MAJ
WiU5S2bowJNT/0TUr4/MgdKooIiA4F25rmReA4TVdMhcE4XpxgO0wvxDMy8cITvSeyolTEGUyzR2
mYyP2LAyJewUubpkdWfAXY6TP+Bc6AWwyOltrqmtmxSN8RMQ+JQKATtjkUXUX2GFRpKua8LQZjsD
H8O46xp191MrWNOi/x8NAuwiYb+xcO5WmfjmWi2FoZUnYa9w8Tzb6MJ7Nc9wycQvVREEOWKuzrS+
0PyvbfUJBhFQnn39sR5C61zwZlR2vO07zZJ4VxmFYSpagqEWMIMvgvfl7xp/Ciw52Zer0YWbhi6k
YY65Xz7wHXaTi9luUCTCLYLEHJeq02GlAijsboQphakJ5ukkikNPMW7gH/+aCszo6h//inQJ0iym
MnLRQFof6VduQzfOgvxYrAjsWbY33DIrH0ghkF0dtOFtrf6zFeNOw/8gKq+Nx3r6tyx86cj6OOq0
hwKDVt1tQ+FlmflMSkXL5w2gisZrmWz4T8IIDLmKfl9vDsIkwVai1m93EB3KJK0k2uvUyrW+7Xwi
s+WzeYc2Fg2KQyzqhvyFUuS7kLKw/yTU1Tq2wXmSGYCUVP85zSrucVudE31funo+j2KRceVjyLbe
8iDdtjiVfxL5gwKUf7B/6fsw5vBdME/LT0msl7Kt7wmr/HgR2BiKYm8a+ZcDIhobUv7ovKaSiZlD
cwPa6elOgoGlhPRmWzjvmCwLEm9RsDsP8UWjPIeFAmOvlhh6XMngXBMAXSo4QcDmUBNLpV42eJF0
pZinmpI7LXctwa3bSKDVhIcB4jWXc5fscW4KKim6X0AKl7fltVwxtPfDJWOcH7CN6FjCQjQZavFA
CAEJwRIX9dOK4PUD27APJ51Tmrgh7RcIE6JypSZLTz/lqwVwKFb4Uk6pUkkMoB3+buEuuZ2rj3YX
R1pMs9BrXEm0H2Z8IC9xVHWpcXx+fFxY29CCsk2tapCosWFSF4vHdCakSyTB3L+KvDkEww5uHMf6
/FVi2RrzEJfNW2w4wLIsvGZIpm3qhjZL/MkrnnBOKsbOMOh3eiZWg9ZjJddsxaPT5g9aHaLtL9V6
0g5QiF3Q1CCeesl4LQorJ5JglUB5Hwp1TKUAicuSBL4y385jKE8/KucyrPXxnIHF+yc//V9d38M0
5AVF5OknE2s1kdbfGpzTXA/sxHfRbhjFV/rv7Bqk5gvOvw2K2ImkK76kKjhZvLKhdSUFdITtoG3b
SlunINZJ0whNsl5Cb1VMP7EbjsSiJtcS2f/NpOwvxQmrzav62jSTMO1k5gdn/28fm98SiioZN+Bs
VV11zS7myW5eKtw6kmUsXr9sGRMiFKKvo/Z0nwo/TtrPmq4nUxiEWLcWMRX5O4OmIJYcO6+n9Dt1
5wjMKv27eKaE0qalsX1v9d7f+DxDvGZLExEaZCJQE6NmgoOJuof7HlbZ+2ETCnv2ZrwJuS0AdaJQ
tOPSfYvsIBq1yhbD8OkHAdoHDKHwkTaW/BELJeGItz6aNWbXWqT/Fq5BkOlqiUaM586rq08ytG2B
rDGA0PvIFBhzDAa62JsUdo2z6kzPdGdUnCPCU7KSx0lk6ngNo3j0Yq6P0w7kLGJDoqg8snthurZe
PDa77R1PPU7Uod16hrpikrLqZN72kxsA/ePty1G+AIg+61yPxRNf/fQN9TtGjeo97GLB+tu6IXsT
vDJLAW0Tea7OEmgN9vdElbcJTXqxbEVzSLxn4wG3FWr4GPmdEpu1KvfNpGJkoNR+E8Zf5SbRiLoS
Ahgdrvxv/51JFVP+oVmFoq+6Ix7vVtAyf10VUiLohvpvjcT/uAdM08aCRkFfrxF0V5uli/wIOxbf
lPDWyE0msXwuj2CTYojtM6TxY2p1lC4Ugv2LOqZwVKV/raKO6jbF7uYJDUyu+bElQu1SIETuqp/H
nblF4Hvmox2M53mBY3i4OPaL4Lm0su24f1uEL9U6biPa4ZmgzSLCeLq9pGIBGyURh8i4+j3g52Kj
dcOyfEmi6vRiN1bbWW59VY5lFJhCiVX4VJ/sU7zmn9zUvAc5+Zyv7obD5+gFtpeFLEH/uzdNeiMj
PIvnkQEfmt7mWbid4vLKiULDb/nuXwzfCR2CzyNo6jdnTqnmA0m9tMACRmoFxcnQY51CcgDXmX67
maAi6W0yD+1pCYS2srPRFmsFc1DRWfo1Y/V8G45gTU4aSUc1IZf0WY21aKz/tS2madyvEhAaoCtV
7hDygE6v84ES0Aykn3Yj980enSBVA/dnbr/qsWie7NwN6SZxBvfCJtQYHNuyI7GsVcNgk/UsFlpQ
RcnQ26Vv4iGzBg3KeFbVO95BMPheauHBgt83z+WPa0nFjNS5Qj0NU3/xPphq6l36TnjoQJReCoYL
uSoJZRMukIKnvMa7vYbae/MO0KhwCi9PaOg75sRT53HpQbOn7gPVmsUzTflVMnXwgzHUYxM7FEXj
jCYIVSz7aU8qOOR3lkbyq+zzA9JeO/46ZFJUuGjQZB+Kd4DH3cGCUjLBkxPBoUNAOxXOMQu36yVh
+u3CbNLBcjYcE7j+NX5Y2NXm5lP5RpaqhXuKToOg/D/PjAkBPu6hSVaKiq7a3aIIxuSuwYOov+7m
JUmjUPP43f5cnueUgL/mndCPVBIIBRZi5ewF2ZNCXqCiIe2Ks23kmwUq71p4usNRMR0iVrNH4DRp
KwDCi5Wp07rgpD6Ip6DA5bk2t+hMtzlaEhNDCqFbs3EmaqKGDDC6gHKrCGICVMCBOW83y2gwA91c
DVcIp9HtW6zIigpbGZLU7OG90f9/ESBiAzH57q07yrsIRFmOvoaAEFQXlZ+KkF+7DTtLcpVNaky6
DS9ZmjE7MD3sD+/WeYRW7gQuOk27XRygovs0eVy1JsXO2fDXSGXA02vaLzBIJNt7ktE2SFi6zVDH
HCAJh35wCiGP5vexZmKvF3qCeT1w7+COp/vP6JoypiiY+Cdn844wzVcdorowSkQQ+B0mVzwVjnaM
0XX8CMx6i1rev0eFEAzepRIc2+J1eTlbOOB2Y0bvzFH6IdDk+tqefn3irO8gQJ5tsgsu1d6m3FwQ
HcPCNfoB4/GIPI7Anz5EuFNMl86HANKRprVd0D+EI8w/hKOtJI/iFi0I3rI7Vh8bc8xonAMc6NIm
kB/uIkZ5a5RaQJUuV9Ypq1lM74EVsY/np/umAjOf6/oR4VWaoE1ux7QJCfOFEowJIN5KXDl/1Xw5
P3VxN0NT0UzvjzWRTOFGF3SPL/pYvrUPRzEIbu6wKfs5+bHLU8s34zwCCqbHdIA1qNeKY70Z7iW2
f8PXmkg/TcdNm5fIOtGk/VuCCxULCPukqcaYhhUWXhES2itjyLjnImttQZqx1F6lTOgcuLJesD78
0Uv9TVSRcYf85gsh71a1ZWzbxz7wpbAEblBWJgB+eGlZBnfpk0/97KUXJsuS4SOx0WDH4MA2+70d
FIHSz0v4KE98Pzcq9OrpdUq666quVaKBm14CI48Y6xHrYW+j3BgIiQ3WjQBOjz3xNI7K4dNn3f8p
QhSjx2j10yNtcFh1+l5nYqEuyTDN5R1t/FZpnOLhUHNKpZzAA00v4nQDqYNWxnpSQCpiNdUx1jhQ
CMYMASldc9OjSE8Dkv/TmzapPC7mfFi3mYRU7WxgHDFIvLVxVn+R936JfechYb/RO/fwW+ggNE2g
F/izw5n7Bp66MQcKLJP5LsTsuPrmZI0uAgen1gxdWQ7WS50iMogUKpqu2GGCdB+M82a+AwcZe6Ts
LMnZRoiI39OSrL7QxQFoN5kH50SbFDZm81uq9Kx/nQgoqGZWccL57XSi4zSPxQ7EKBq6I9pqL27q
F7Soiq1s5TGt5KSLTFCQcqflJHVuM2BD9w68iQYbJX0IndQk3IVlqM9QnFpqksIsLzP6NLg/lM2B
SbymMSKsFy2AqToKPBYnXUD3PaZg3fBtCniD9cqVbsbtj1yF9qC+cS+Ul54F/056V9CkxKDl3N3S
s2S4EocISYHxaeQKxLExkRkmtW/TS0DeL6U8O2DHWBS96g/bYc01iuRsTjyMSDsgmnXQGku0oOYT
cm2ZBq5BR98TUvCswKFIJtkRQl3/DtkR0zmgyRZcMnlE2q/VaJ4ZivGwpeoo03ySGr5SoI+bKzFv
qz2VrOXpUy0MOeUaY4rCsDtYQnYdeuPlIfdptRais0rEkXYi54/Rmmgs1XCuYqqJgbhg5784sqOO
KejyXbwd9Hj7EN3rX1i8RIS/Qv8NZAfZNUuX8acxFNVvJMMywRMn1xdOLIpkdOaVs+LZfjcNGNGD
toI7AvJrcZ+odcJe9McWqbR870pUqA1x9i9qN0XVEKzADv7pl3e5PO6Sh47hOKjdABQoJxDJnoos
FO049fERVQ6raAsruyE34BgY4j4pP1qWXkRAlAbgZ6+92aHXjX0f4F1n6PHDBTpSxhf7SwiTno/d
JMGiDs7imclzDKNCK3UmU6aDaabsS0gz1CpSlLJnyPV6mRknSmZWMdPTiS/dbfMOW38It9aFclGw
e5y6+cQcE4jR/+h6rmQQ+AfYkAUzstKq7S87Vl49cytnWrTCXVnmr6YxWUoE1MxwIoTSQYl3AT6X
CxMc39yiczXjvfUWESZc7fgAjin/xHZqAsiVREGsHeGCWJmuC+t6lHmaRJBwYPUCo4RhGiy6mA8J
aVySTHDz77rQYMoR+Sq8xdcgLBBhxfFu1o5Lxm89fi/10houXEYqAnkx+txXg5FojN9EErGfcsPY
EpAf6EqkFLwR9Y7G6PD19Gdoqzf8o9dLGZzJlzIG4PSO/wTgzqMnIRJZZr2F/Yn7LUKcpzYJBmdT
yQGY37cn9ffJK9ZQOt72Ikfn0kVQvpEsZ3bgi32qjX1YujNFkevUUJvCikqbcQQe1eaVA1LobqLq
8zQ8a33xdHLA1XPNPAmnH8bHuUs2gzVgqsZjuBWvdQVenJyMKNriRIoDWOcfR0cczeAp6WbhWp4H
3E5NlfHShlyBG1GFmL77t2oF0iSx+RRADVCnvvdqyPwB425oH77qu9sky0l7yYFfWl104XQ3v7lU
x4IQ9EJhvQg//gPLsZjuvW9YBgcXd/I+C2gnX353XUNlaQrqGGRTMGBrgwD9tPbdwpJld6Cv+HFG
zBl1FD+OEaRj2atBJE0j3isIndNUIrAzocf2SZcuo36DI/yZJhBpIvjiEZ4XRJYl3QRzD6JVI8c6
w7QyNBUL6edGJ+ZXcVzLfhvFVJZdHhvqrVQgHEmZ5/JiZOLtzzb+XmMT6t69Oljx+6aTNcKPpN7d
tfhEiK7bd0Mm7x1gdDAvnokO8N8G8LJFKPr6956ZSzTsZuhcM6n542J9VIFAG/sC9SqVe82cDlpW
4YUYsakCJWzfi9nL5BX/OPqCogyfEqzC9QQfX7xbxMXbuPUfDreU83qpWb3UPZD6J029eZM29Raa
BcdwLMfLSABYPMX8RXSPRowYIcEc9H0/7vxH4JWmFjd0fZw9hWWwXLImwEaVMYXrEhQckdRNOidK
sEGFKxxMR9h2bSdCHCHwuhwOsLrC2/Qp9/kbBtZCYf00f2rOYaBvXBCO80EehL6E1vf6rSNkrpN6
sTYMvGzc2sKPx4Hxz/Fl8+kfEwfH+kfI1inu6LhryDrcVLDcjDj/miV0sG+y2ZXuduWjhRKzLvbl
iV7oD9oCzeVQnj9lzIYaxdlAclTwz/bsrq6wrdyKGvU+MnOwicp49XZzG+IA1gU85SA5u2MjMn9g
3ufJZb8fb/NokK0gjGxtv5907jqToE/7qDOFJsDW9QLPJTBHBf+UcfVaeeXoF8FYl8TCXv+bN6M+
g722g38EddqFKl7Ec6U6ZN0+GKORXBkVC7JoOuK/uuA+9q7CFIfTuAcHuhl7MIqJ8W0reZfndNLr
fZkLP+G9kzQsorrhwDszfwP94JOqn5qua9Fb69vL76AzrJbeV5L9LmneZ2IPlzdHOg19P/TtIvu2
KK6FADfZXr/PquKLl3goD/SF8EWPSdT9NBnYs8ZzAl6H1KMMP3UD9OxCwyd5bmL73hyjInXFMCYY
DUtwsAkkbZl/z3Q7CSwrC1JXAcUixG9RwANURA8+4G7w50bxfscWSPwaHQuJIg6/WLlyLRXsE2yW
7oAnPGiHHPmEehHdcWFCxKfCSAirFGt/L5C7h5mMb611kOf8F0fTfQY6gmQnIHvp0XqiWquFPRfy
hZI02q7gSn3hGcEGYzTudGVsX6gCNhvdjHdMTz5UIjK9A/Cd203r6I8fURC4ax17qabI1HAGg+Al
h3Yo8wbp6eq52mEdilNseLVvPeVFYOoXwHjqlSCbU4fbqdE0XZhZ9z79SN7rzoj0BPuaDYTPsY/g
FO+Uwkvl/rK+QdIAjGHfwj8YqJK2OylGuagl1ESt8Pq1RYf3VfZ5W5xL+P3b12j9EbsK7r/5phsg
JOLB/c39EcaDzfAL/JLsfCfpucDzo7yXlUkVPjtb8C2P632aKRAP/Wh3d5X2TidhSfzCRxQ41AkH
r2LLyutytCxIrBAkOcreUNioyBOsD1/yXCoq6eohLvyk2HWgGFlGdwwK0rcoIewVtCEs/aTg2xCE
GA+nVpjVt4e+goOTJRbmGVjPONag9QBAJ9CWEPYz8X4unBIwrq0pRF2qa8FmmGCSeZcsLeunF/5e
4dGBzE/Zwj8G5pPGo/ffe3Hc6uxR2d1gfaMlDx4o1PCz8g0/V0WXszMQ6+pnNMG3L8tWSRL5fDU5
9PqkAZGmd15B1HQbzvOMGaqGQFmXf1biEH25YejEF6E5S4UqLiDcaPm4G6yallxClpK6Ut7NVDFO
W2Ebr/vajJPSQxJwqip09oE+TA39Xayq8R/LxBWifMvRrGpe4YFY8SvGmHBHjvBNkoh+C2LSqGbf
YtKoIHzcsxTUpAz9EuNA9kU3iVW+BgK+fOY7rspBADJYdwp3S9MYKPi/NLOLI8oxR5X0Q2nFfLpP
6KMnWrzUANiIGjIGL6JfpPc1IJzYwFYWwYipo2R/dBYwGobJOSPk6OiNDgB10EhBU/iqtWBdCFQl
wbDwzq7ScOErxcGHPpFyEPl8B5uihdImJTeBa3Sehj/fTeoBDGT/OnQBzldijjpiuuvOs8Mr6j5z
hKAR1++Off1GEnrhcRjx6V8mdSabMxdkEHTvBjlJwSUslmE+J33gmrnkezkGgMYsgXc1KKhXG8om
9DNlE4KQ91wTQHXSv+xBbSj4cUkAA5mPXg3b+sTT8n21pieNs7z0gLTw49y3YsAOTEqf8nrNZkjc
UtzqQgJ6T42NHmrdhAR2Lh+hIuZy8YPZKWcMj8LrHd9+3Eh7zk8pWzRA3B5BdRwKbsPGKsGNFBYw
Ozr6Aza2sufYLTwCkqxZW6j7kVCv6sESz5O6uJRzCJNVUX0nhvGYllvo7Bu+27+ISNNDZ0LnP0rZ
Y5OZfGazMiOGtmLZax7ymAGn6cUr506Y0/Q3rKIF+Ga7veXV7j7Ebi5q5HaFS677bWPWBRyD+GnY
uVhLryHAua5cxrRuv5NlJdngeWlGa3e2ML+VMizbKKQo3FlNXM7vnrMoGvvlC07xzkapnRMHgxzT
XDDPmmXpwcSPbEWRpKVZlz/Al4enVYBDNWdA9a27L+K1YOusLYtmks6CoRdcWi2vhrpOgnm+qAuQ
UcNbcSuYhis42yYZwmOk5v84dun7hrZg7IY1+pz5iImuTyZSnXTHpZIhKhKH0iLegWMZ0SkyQcCJ
U164wzEYzfXgD3f7ZPh2kXBKrDJ+WZMAEGn+SeApvO2uQb7u8SLSRnDD1oGSAorGP7lTDnmaVXmm
BhrZ89ndi45Q7EkqqFdNMHYd+dsxM2uuGubBni3XtdwgsRvway3bPqmTM81kW5Sw0TbJxEuOAPfY
ML5ATzzIMy0ZqYUScCY4txCiQiFO8JV+kyf2pVW3lMRVDxtTqqxAMRi1dG/5hqrIrbEU69WaXG4g
sTavt/jFIkEyoAdXIds1D3QCVFW9znY71Lk/Tf+3pfayi2e8IqmQdTDwQvVHNwug07dH5oJPa2gG
RLiOc4U5VkSpOOoHgA64pSHi8vmSOads27zFH2JP6c8gKUiLOrBWjhDUD6BjLQt4tdsFONH7A3t1
A7+ZSBbLxGeHaarL5XgklnSRUe5PkwLeQxmh60Od22lnHdpIQJAsCCvmzVu6xdMX02lciauGfpPJ
qa8888eNkbIwDgGBgTY8WjoBXIA33p7XzvnJS0v9+SwaUDF+C3oUMx9eSITP5wUp900KCdbJaWHp
wuk4jqaMzx6z5/54iNR7H1cZZHQ2Phzaka24ReRz9/P07jpzGRvs+ZaSrYI9BpxjfvmEHU2oRf95
OxqOSJt2OXhndy0oFrlWbopjsjudY+b5iqJPL47bg+AoP/fd9FzXzzUalPzxoR0A8C0sHV4iXsRD
6xOGpKY6YPuoGsMga+Rh3nlpZbwgVKG8BJmjVmoS3IGyZDQy4a9W1a9SWMeylMGaagwIHd073O27
i+oX1ysVWI/pcn2tW9obhp2RCGwyMmi3GkSmflQWdW6VdkhGsoov54hakYxW5iSMN4JCznIBlh2g
JT3mMM4Tpx2p6h2vnNuHiIJEuAiwG4eyVeMmsbnmfLJ8zInhknyaoBNYDXbkYeMTzJH35/BnVVZI
dQR4ajous6VUvEkWPiM52vZGW94bvxaz33AyPSKBNcZn5NvQRGC/3BJmwRO/GJeAtpt/sYcMiqQ0
nlZkIK2aZ17NgE0JLYfAVamunjZx2zZHC4QC/ImK71zzxQ8sld4OPKOtvDbVnm8dhupl139Oo1Ox
RvrUjQONssErc0oJhXpXYKrz41xUYSuV1ZNzmJkyWhAsMVpjIn7j4Ge5BW3jGpguuA1up6jDmCHC
aQ5hPCdtHIwC2O79fhPzv4kZ7Kf23UqAdHxrrEzx+g8ekHAqoZmW6rsMmd7+CKAEGXBR1tpxG0yG
E55YhESAX1Hxfu9pskfDN0tqPpg4gXGJBnsuhxV0nNFELV5ebHJismDp43MsEllXf9gv1ifc0s7m
dRwMZsr2r8NgkEHH95OZd+/Qo/S858yZ4p6b5e3uxrf89uPvIV/jRtn/8AhJT9ZTxT8TO5CvUG/2
YroBfX/uGc/XpQ1k3ohhwBiLHXx4rGZ8WPN07HcBUpFF3E5ToGEIyOc+7knV/b9CTe3bp6MUAvpC
DEl5vUms3PzRhjjv19ss2s1c5k+90Ca2C2GUHJYrKYPBzhHgo0d7E1PlF1VtxNPRW6DqtDms8Y4X
3gdVMuFOpMhcpiblucry2pGWQDhj7JefkR/Lyqu1w3nPFcbyNLdt76RiGEvHcSZXpz1cgbnSf0cD
mXuAqtxIx2rtP3ok1J4B9VaNEamh1QCtSmKSr4Xiz7eI/TTgcp84Qc3XvfM73wAWdupbTSgZ9194
EjBn67dqv1Rz2hJ//Pmnncf+v8QqNrTRG702Y4ytFqClI+Q3sUIUL83YqYFF0feeeATwcbYIPnp2
GYBS9hfE10Q91/2waSSNDI9oQ2fECBftlTlmtVXHtTkmt0HfpKmE/9gTf2YJGras9aS6iYt+z+Dq
hGC5RNLfqlehgR+twRjlIUYOnS3HycOzn8V0ntYF++5QPtYVI6VC/wdgx0zN2T0pizR0jDXqIXUh
u70OusiAXmJAybyXAzdybzPmSedxURrYPop5wKkLEVxT+M/gg3a+EubIaooONkJ2HNHSVHHuhJds
aADC6iDC1N4BeXcCYSwSjPsWnikff6Dh4o/V2Ltz55NpPPJOtoTm8S3gBxdRP1YJDalyhpwslHA+
QzqLkPmI5+dL3QDvVLFSta1gmsqE4B3QBXQAO152TSIKl4XTaOFSAO9V2Xz1fmmd45Q3jE0Xte9b
NiicrLdkX8nMGgAdxbXOpTXn2wzVz54yM/8nlaNCB7/pFHuxZtRC6TgqXUgbo6NO0+In2zRubqVi
Sg6bx8BAnRvmVtkqE9EaKTCQFViIlixFwh4IyGOqswbnHSviRUPX2Yk+5zc5p3jV7Xkliq/9QUp+
Aff0JYL9vu0p4ahLjwhrWjFmUOkHvlrnpEY2FNBZZoTOEW/D7G6wHT2cnu3O2PUcZuiynddq7bDT
gF6HZbItce7TjJ3rII/DvZ1ifq521rRsJpNHRdSQLALQq1W7ZsaQcITWa6+C4d9edslIm3EK6/ti
nRqQx2iCpzLUxScqyZcx88dj7qEmoX1BXLR5CPDxS5dhyo19MAa3TYwEwFCN7I1Pm5cEURup/Zss
J8AlXC7wCHmheZuQckc/dXu9vQX6K71tGmQqU3twKqH3rdyHsJ/gfSDm3So080eVmp6a06K9q0qW
pyWTT4CkWY8k2oQbiSn4EdMktX0X4PwjUQVl3+6eaF2KX+p00uPhdAixsp1eQEw8S9H8Rwqzg7Qr
DFYY06ubb4AAA0NZzBW/jRaQngFCZqtshQviUzqcDXJ0rDkJT6IHg4so07+KhOeJV3t1DPJGkr3V
X9xXJ9uIVbD1xyLCFvN8shVpdYMIL7WjFL//p9Aj0ffzdO+OUVCzaaKL8RT5DXV3MZlyqzeolr07
TYZrQt+XY8yRmRQntjrrWj0b0WvAibHV/uQ4PZyASTrfxrt3AkwAbTSpvCoMtUbvUerUmU6x1y20
XAvM1DFQtKRb9ceaRPW+lK3Zk/uTJHe1HGaUCk4GPrvOZflGX2WwbBnLoWh0bH7aiQIh8H5Lk+1N
giLl5fPc/fOvyJQ4pu8F46g3PkSvLFjaCbS77bYlAbOY10dSKri96Yz0nshpngiAGb0PeLdKnAnL
lh7o8gJFSq8n464UkNX9/FRB3pdTW32tAlAYXKHtTIdFfrGFyT2eNfiirUSLpS8jpUFxU29TAIyd
+bKK4vGdYGngSkYJm2OytRvZu1p/xV6M/jY6lon9m493Ok/Bo9Xq4voNGdMvsfkW52PMtUM4BCer
qkPj27QFP047j6SkNBTkMDDsCzO2SdCk93Tn5sn4fXk8393NpMmoqF0NZyaDz3Reg3TZfR5egSPQ
jM4KuQKGimPCmM071iGHaXLMWrjibnph7Z8zMNTzad2Pluqy4LkDvgVleGrtLdKi/ThL0hxkclJm
IXopHNPpkfFWHrITt1JfryHfS+2UyB5wfMcfU5+RnWkki9PQ5xBm/bv5GCa1Fdry8nWdmsrealTQ
9CYsbRvVEF5zMT1zHT4f06XwEMtTTIZgUgWsbJSw0UE7MnGIrbuQQxcKpTQKU+N4qzbDexzQjfls
IocvlQ23Nr1YHqckauqNpHQGwikbQrB+lSJabYFNbn8R9gvqAuy6eu0UaBDZsF9bZssVpSRK38lj
rIyLcAlNuUoWqEt5fqrJAAz0VSHokTlwOcA7UaEXrZ8on70XGNNgkUFFIfa9WzRmSENgv1xsqo5U
cboyw5T9VlpjoQ8bSU7skdSkGzptQrxzBFaRmm+Y1E9+6AiOXUhN2yoSwnpMN5d7Iv476iXknjSf
P9o+v51kWN72mbj+ZC0MBupz63/92kq611yqgapciRv5t8/qURE9UY8safpxarNwGR2DMOrlhtWT
eAUr5MuWrVWltjq4AHU016OqFS2GZqKzUVNCCrvHj3ehsdHfjmWxdZ77Ifd0ZTuEmOi726A+UlUi
D62bzVdCokeuObdzL9cSdEK7MXDKx46ytQSL8YLZnGyNOyggNWieitfGwisEkI14dIb4qFjdOVrD
T4+IypUSjA3zmANLUYuw2xnO4xS2U3Z98LaBK6sEJjtDM+auKnx3xuV6h1C+k+YAIwCjY5uqrLv9
GUmh4Plk+T5kubtB19HhA2bi2MVedSyFm7FG2Q3K38urhd+oR6adirbbt0xXQ5S/Pf8nq57J987D
ChsW2KEsJgpgt56jThIJpeYJQvBF/gMIrWAZ8lBjp43loWbpzhtDT4vv13ekRT+n0YcaTZ6sCk7U
R5BcbVwbX9xUw1IQZx5qvl4kNeJQtf8msouFcVeW0dhYwx2IGmBlOtUPcgHGJj6kksi9O8yFvs91
8g38f7FF+yrAH1khD5SlFZqVwaBdUYO8Dghr8n1wup1v2k/4WhAYVCWhLWf126xg5fpU4PIu0tZd
AmpDehgboryA4+PTlkA61X4c5as35Ug5CGe7WcwJsF/0OZ1LBxxAaqvkqV9dNqRCHTJiJUKd6Oha
137mRyWq3ULWWuHdHRPyPDQecbZNzaYdshwwFszY47W+wsyoO+0uti/zgfNvX72EHHmA6oxdTZaL
xRIJh/8zlIo/xY9uOeTiydPngBc2GIOLNw+ybyFYaTvpttaGbN1fhFsnhHrSOm9Q/1EjRyjy4Qva
dSFLeWJlmcV0gh9g9z3fpngwm3LWbCogfU1k9eiK0jP1x0lNjqnX4zXXsK5SSl81V8vAL89yZhDz
sToYo5yIdozdT67kQB8uTmei08uHlBu2nDhIec0jO9qxtzF6LH3EqIeKMidjf7nO6VF7SFNUgU0t
PRGspw+9+YRliL2xFSzWXriptl2DDD15c1wpkcw0qRJZoOIrQxVdOWRTFFIsBMuq4QygSa0Gasyb
DERIPlI9oSbnbGUqdhUmasrsFZV1y4Q3tcBuLvuMrDUCjz9CE3RWLGDIPZMLfqnjZaO5wVDWRDO3
sbD9JbWk5oB6LXg62kxlIT5qV4ofGv6T89CUbl0ko542qJq3OPT61c81d0iLNad7TyVAfkcQvqIb
DNNcG/+OVHDAI3dpe2yZHpvKZ6D+HLkqnB91fhh712HBsk0C5avaZDHfkyrxsI6XAsMFOv1nmUUP
7qJq1qWRtLCqAXHEE6VusQbdi5DXROsivz/fh7uIKD1A7Bodd/0rN6pXkWwSA3ra7eH67B1NSnBK
rNbQOuAmsCCMd4PZPyPvQUwxJuSNU00v6Lp8KNrzMIQf64badSRmrrhV3mJcKWvtzkmC8ZKuKQ0w
yMP5xlG0a9gQdCFxVenicftnl1svbqag2WYQDFTzmWAOvlmuViwpuyAiUTn2gCjEyxl6agwpxl+1
uNhCP3yvwGT3wzIpa4/kWnXyoqrAPI6ctdMWmc+jiyeXN/AaWmq5Fk/FMaW2tRYCi136jq6X6WTt
PfW35VUV94FQ/7bMFMQTX/HCxWQBxkFEvJ3xEKkCI3qNPYCmlYYjbZz4MeM2ybu2vDY8bavXPn8M
FEAX39Fz2/d5GuB11fim09mo+9s47LFQfdJkjsxog+b0stuzCJd7pQvscY5U9ZqSQsXBsYHvaBVV
ZO2wTxxsyqYIpadPxJvuXd5JeUwKyvljynV03oZ7cvmviE1/Q9vz4iCgT7KbIqzLGe7FGbSVCdyq
hOhhWUbmZ0iCYDHX63Ly6Kk42rJs42eh7oZA+uhKHOlW0jy2EE1bqZTmQSPVKgD0sKcxSxQ6xux9
yBCs8VZpIIFMbta/840YOaki+lHjF71p9N4bi3ZPjcQU4pX9W3k5jWuZla0yKG4KPBI1rXsGeRQa
ob5FmZyvrR/97lzaF6aQSeNmazdf3pH/YSD+0im6ZT/eaRPT7eFTEKOf/MW/vakjt9WwHSiVdIFu
rB0W8dh7gfwnuslhRHhqsYBv6EVT/X3+50MbwBAe9iaaaZOlfe+jihB9tCr4cfuU+lix3k4+dgqo
wzy1tbSqTBgYzxJujw5lHhGte9Q1onXclnnA6EtoV+D1BR1SF+i5fK+Xu4cusPxbJBxmrMy8p/xL
Pv1VkZ0uXRL8SvzroC0lj8O3WwFQesdXoc0kKeAVs2If2XSNGe21YKnZGvPYwA97pMTlXiqUE2u6
5iGUCoVI8ADhzreoL1KUd5bqZwc8jCPIREE+0KnltJ70hiprqtV6CP5LH+t+uTjZ4gO1LSDLpyhf
M24bbTU7o6c6mZ8v4wSV0kGw0Kn6ZX2r0/tBQk/hVG5n7ieMddqobroTU3d3iytvzxwdHMU7wGK8
9vpg9rtXQltpuBacBZpkGBycJx5Z0Bi/dA848QPSdOSM26SbZ+hqw1VcLuYfyidwQLYKkSCQG0O3
Gbt/pnGwUBr1aJLGZcAI1kIP+BpeUKQMhFtDe1SmOBA5Ge/wn1b1H8mOq4EJP68o6tUh5TLCPBg/
dUj2ta31DdsfePn0x+AqKjQXaNaOiMlHVvvVil1ZhJyLel86sDOGgLmgrbXLBW5xV3BtvXYYENll
I1ii9pTvIyHYeqUztjADJ8OeSWZx+dqOG/FEzBRSfEb2MVAUGsHIZMXyePV+uTAugeeGw8iIQ075
7ZRacSDL8sBtLkTK74xYTUXBKHCVxWfmRuhzvblmHx8UtuRAyYA7NeLb6SGQZCjZg7xIP2P8bQ9U
YGCpvJSs7NDv9bFa0uml3QBKEpR8AsiTXjUJrWGBtxsR+jkBERVZxIuKFpyeF5CQrA3+pFv94iI1
lh5xFoee4gPL6Kb2P4lsy5gc+nRbpLuvJW18uV1aVhv9+Lk/pI1lJnyAi4QZDL4unFanxNsYNupl
Lm+DlS5H8NJN/wcgMKNqtG5WcBob+VmfN8tMcB1Z7hzCJXAewJY5Ooxv8mmtiQ6PavMU+Ev6KunX
lympeJ79TcBt2EL7rxSDhmbI4NBf/C9mTjRp0EW6E69457LEVmtiJbmDgJ1L8bBtW35psTVAj9B8
1yHB/gYlKPQEWhwJicBC2q7/alDjzN/Fi4/J7NPmPOJ9u6vUp1y3jEztw/28sWg1JYy7MuVo3Yda
+GU4vyXDSeCKxT07clknIEZ/GiSdc/G6mlt74jW9OVsCqk+6rQaz6gnv4sneHN8+jEhRX52JkUl3
6bNm68LOGvhY3bnr6P2J4NimhmrE0wntZ5C8sNF04sBEp4kn3n6Pl29m5me6A7MNSzv8lXmzUoEV
sJg50dET2jGvo9Twj0qqE+CSzS9Nyt3WTeggf11Y5Y6smXntPomNWkwph41EwcYP2hBdXVfdkVUs
98+gvmCeXA5QXOvQOYllpE/rMLYSSKl5xNZcuyTFOAQI/AOwUJ0bwhYqmdIv8KYtPvPuQH13t5jx
6btCTSMdumj9HovnmTxVEBh1Fy5i1TMRQlcpFCdREt9hdIRD0aQ5XmU8CZSkrKGzxv/lpcTCOQTf
20DyceSxwOpvYPUggYDJjdBj+m0vLoUlS9jKo+rNHVeFHTK6Lzl+d9b6vJrXhrPX5MblVxznWU1P
vuWnswyiwNJUAcAUP2XJMu4/qKos39D1drewH/vh+D2g2PX5DQd2/1HhvroedrqZ2yd78ozXPMfp
TLI1wGEFzHYn1YqUrjSI7FfNYEiz0K/sF6aL7ObDesuQpV++PQemhRzTW++VzGVr5bLIOkUvu8zX
Yx8HEUs8bDdZhkgVckdoeuXEnAn21i88lgF404HdxaOpdzi9MaDiOT+Q1PFrebZXxKbk17YA6tFx
jRFiDk9XURq2HldF1e0SPIUrXBVmjtQ10aXl6Np1uOrfErApH7MdUHwTGL7x4S5cLsLc0RQ4WQRM
PRiye2oWTWdUUw6M3wHt5fzNVad+qdtWXB1kNk5GQoNAYVmJe3+HuxSvGXvBtDIlGiUiIrnQ+MRc
/oA3gpn75wFQllKRox+WI+mou4mjzdwXMJEcWCvonLS4ALiPaOS9cjRT2g/TxIZqJxOLPFemczLK
nvHeKaqvz50OzAwhly9DtWrKBkEG0CgA3jllG18b1wcXWmb0ImD33aio26SQ/E0wSQFJze3TUWgW
CBdaFgTzOL9HBve+eI69B9+xZE4i9peNSumo+JrrMqWDpKu5eUqeogAudjniGAQoOERfJVMdhppD
bVo+di6eUNlK5gPFJtvSfwgXyByGxFUbL50QF907HA/b6yHasJyGtZQ3mGeZ5/61eFzWfvKe47FW
ZarRuMkOscavE9dtriEUoRHRU3LaArxD/yjUq7OcS4OzgX0E2ET51ozPkS7ftVv/HA/4sImLtDNF
zJiRvsl9Ae2dj4Cmo2ZJ9fAuh+Q3vaJQzAJSurUZFonDDWosT2feeG3L5KSqJToL78Kc5/Zm7rxw
XLbiAwRRx0ANpS1eHy1fMkceBx5jrBnap3/J1Vo05Y3odhEauyOUX6QKXcCq5MASfvCBFh+Ms2cg
XQS+f4CM78vY9ylN48fwo/qm+v3u3BKr5EI6CelQOda0zI4mSkVM1QBnY6/woJRmyfF24b11GEyg
fG/9vtJm917NG/4RE3fjZ6BcwfdeUKXhwVOB3GLu8YKbvbBdNqpg2oYYcCR8TRn5NeIzFkOeQd7o
pcCVXwQAlJ2mf2Y74BQuOrRSIMgDddJGQt4brn42n16VUkriThnBYsGP7rpi4dnX47GI3JdeW1Ky
owbO7mlmwb2ubuNDfKbOijeNOFuulhv/cIKoqH66CphRN/PAKxqU7wRtLFAH+uuk9I/JukXBMH4u
o/yLU8kCo41OLYEU7Oz9Ypb60cxNkLVp/J3DrdnWPaasb47RG4vIyhTRFJjN8Pwd7o+qm+Qn3szy
6saLyDr27w8ckPIysDpJlhv+JInLrxVHKMzW5Q7zANVKLgsp2VYSt7zrnKhCkuRM/9KjZomSKCmU
IippQ7yJNg169pD7//FfgzaVOeD7+ylzPBRH1PiDZAsOn0AE5LucDt/UmQBXU62jwQnpSyDeqgc+
jGG0JHRgUOia+ITS+ZMfSYe5fpzvzyffnl+jl5gICKCcQC4/JFm2B0GgBGICNJX9ESZ90Occdbwz
sbG845EdSS+s2FiA2p9rNIlhURA2h/znkjHsXba0dAax1PRj1AwzGp1vsij4DC2S/f2g3nx8NFbJ
5XbQbS0+jnTn3ThBB437TQ/2HhmBUwGVrNdU0cJ9DEHgGkEsbsAZW7UzxkPzZ55eymg11XJevQpO
itN4pb9tWurvYhiavfgi3UUhcutGi9uHV1JNm9RkfQzytWEwPLNHF0kttub+pq4uRT9fmkJ17XnC
aLNXhPoWuRXHEv9RzwDHjqvyFZp4am0gaZll49YNIJ0PNU+8KxVPAhHzqeWRay5qTmcNH2nrzgA8
3Qi4a1sNDymUlfHpCIEmL2aX9iTuzzlz+L0ibRnxy3cHb2xxMy+HAUG0KyY+uePr2Z8Fxqh8xVUs
ZfI/i8TVkn1+N/NBCIdkl+M0S97WfXZ4/mnMKCgT2kbjCC0gAkUrNQBGEywZmcqgb0e8IA3m4bac
Ww/FWeh+W7gajPoh/n7nHNCAYMOTQjUoMuXVJ83NndVdHpD25v40Nmr3hg1anVqEVG27zPd5kkLI
D/6iidOXrpWL/iIsObRIBR83GjaP1Xj/ZZ1zJbbtbXfLVFsgQJO4STq69eW8imRbWKnr60tIywrS
A+iq/NEGm0kaiLLyPCPgD10SkXOfomr9TnCK7IcoNxzVLqYufuXcalr5Q+KegPkkg46KUuQcJ5+9
1Bp79mlTNse/TR2HEvnCPe5zcBSmF62puqaTV6Thi6fVGM48BS7Vex7efPgywsLBOxhYLoTF1SR6
d89xypAiT6zAzR1p5mTKUwOn9zneKgmQm5UVK2PvnjSs9hGYkFm2OHsc4wsX5x+7NkIPwiF6iAr8
oXX0awzzQusuHH+r+dqKXbYwFQSl8ZB+85Glw9CBIWUp2uF9VyI6Ejl1GSyi1zy5rkFjak+jx7kO
9JMQgcEcpr6Hrk/Z11uzVJE4B58nA6W31li2Zcxa2OURaDhXcmO/czRjUKRToySOz7ezk1UFUWV0
GB90+ls5+jiaVUU+GTNV5YlNdFV7A6qDNW4UqpQ+P/RSjvGlSbLTdil5T9khUTbkhmRsNzIy4g+g
ZR2lY9ptrz7AMiATpojLyvXf2fwyh41+gic8ncvr9BCxrT74DelgVfAZpToHlON1BeaBNPhPGu3S
dUorwy4kpdgdcMJU9xP7WBGbHqzrgJLJc3NnRSDgNuWnG+KVQBiiXHXkbqdmhwhaKN0K0e5t/RcS
yBHCIBEZzszXpx/6qP6aPNxcYYJ8wIT6Zx7SJphWEPepz8u7BfDpqub+3GADd7KkvZzZoLaj1xIw
V+kNjPEizEdO30xJ/JvTf/r9Kv+3oOsnG1/ZG4EGhuJ34lhf5FvzeQu5ak+Y177TLe1aP7ZCjWhJ
dvvOPUsut+3ecIqCYvVAgIyTkg1pD2aHlLYIusasnHdYbAYmOFIxMGJCMWp9Ea+wHINF8a/59CYw
MPgFHJPYhl96GzizEsQRoPhaiqF8alzrqUVY5luBjsUn4lqc8W0sJ0mxdjJBjnIGwlInexK8ugVn
8j3dMtiwFkJhMokZEim4Ha0bloGDklRcLjpwiJd5dAFBzT5iCZi4LXzyR/0PnqcoR3fQtZfwa577
X5myj5q6IZUIcFIJNMhG8aZB684hILDhRwaROmC/txPpiR0lyJeN/XDMTJXnVC3vm8gK8hu2i3hO
kA0XC8O6aLXWIqoxji8fgsDiNptYXZPEdXDUVOffQUKh554ue9OONRf0tI20dAdXQI+x+v07wL95
ZfKHdm9WD70vlYBIe5XblL4/SLajKaLSS7l4pImIvAUzdSaHdn138ZJlB3GYX5y391MMEDtZmCj9
iKOqr43xHpywRt3GG99Q0FQ8oYOfeshdE28mbin4Fhauo+Bxg2AQ7DlQFw+RPlqtMvsum+uRECep
44AVRHe/lMEEut8wvmT/iyySIqjPFEBnz+exBu0FiuSoalNNyBYDj0PYNmWsNqSoSGEwjClNinVy
YK/8giw3mZh+lqij1tb7iUARWW2MXfZL8bD9afnMSOLoPnUUBsZ5+G/MBIOKVW/D6gt5UNpmnAiz
K6Ntv+AGuE+mm9m+yoPitf+AkTfO6mzG1v1xXlaIp6sVXN7OaHFylw/60mdIUxHhMAY0TEwkC914
0DKrdy6HLkRvA68ozdbHxPBRiodtMiPADpnUtxcsHO9J+4FPX4WQwFeG88bciixVOEqtfD0MgMw9
OIFcePBtr+s4SUUuF0BfW9+Zpb+B44oK8b0FYidS2Q/donbql/LfbZuCQuLJWwDzT+uaO/dn/M08
0b3mMXAnmpYKfOt2Cs4nvrWbDyW2hrad30wYln6uxa0aw+J+ikP/JL58uDMVyu0YnK0f4hydCMIx
OB4mrVypr+0AAVUzN3D6sj9ZetyEZKyPfAFplcHk4vrP2gEw5MaINrfE7RDdV/dX7btQLHXAz9D9
54+VhTraDd55wexhSDc+sunaz+d2/s6XPSEUsnSHoULx4Nuv3KMXfEaf5Gcxb//EeC2RKYgnjr3t
VMu5GLRIS49zM1Jy2UmXPcUfSLMezTPuSgCO6MMG9w6AEPNLdPbMyCu1DcTSv8hTlfMWwDwvvuzR
2V69khD+oABYG3Ppp1p0k1lJSiuXF08t7KVOKENDfht7A1bnBUbSX8vEkihhrvArrZP06lY9r42K
AAwr+sAn1SjIapKmaB4TV2icDKY1m/MaIXOdN2c8DUB+WvFmZHyP9NWiBShJ8q09YiN6LGo0gd1E
dKPr6u7sjhZUDcoNuRfllKm/AEfn6rdY7rxMXWJd/o7hEV67r8Rfdn/2/yymTv2nX1Q3wk5B9MRr
q5cXG68QjLMe8eD78I6jCxCeKDH6ss7ecipTX+tck0yYUcA2OQMYhPZgZ53Hbzu2ZY7sGP4CQhU8
JQZPCeXLvMioV8c0rMAfy3pi8HfQwF3S6QLr9TAEju//yGKq4xTRxtNcBTwFd4RLqtUZZhn1m+he
rMMBsFUIfFgFU2ecBR6KTZhMe0fgHqxCOnTg04TrIrErfhBUnDRsWZZ6Bn+cfMgAMnQBGtlxYvJE
8iuN5wB+2LqoH63y0Ib9SrHRBtjA81bx7IBB2gQb7stBeTg0/I1UmYJUFpdp+nTXEWUQZntkwdQ6
2JHd2s4sTbIIEApF6TV/J0Cb+EtppbIR2Qqa383d9utqtAE16qouI4qhzZyKb6Jzb1dJ3l5qODuX
eawLd0S/JRSEKHliznXCOTLFQ4Vq3X3GODjsf/Z2vCI/jfh8uMslvhVFVneOAeJHBQYmyl8Yisml
rlJqs0EQC0KbIySBKHHI+OONfczH7fWFIXjNZ/6N2ZDU7W3ZIZfrWgrClEKVuWe9Iv8btH6elIJb
oIkmphCCY29hllCxsziNOKpFzFLsOy3WdlqadLDID/9prvd3czmzxM2lCY2wxtQNICY7XUL1kjYa
yVtCCwVHTPbiQ7uNwXR8Cd0SupO9JX/RgYmMQfr1aAWamtxJni58mJykSO8U6gcQhKUY+Y85A+WR
UPlJ5Fv+fT0HMPSqorAjP3BUbI9FDIP4eYP/R1dX58kpeZ6NA47etYNtc2zwTzp5qnReOg13tIxc
G2ostRMN+IIQNQjvSVgquK7pjK/iV73AFfp0aPBn78UgMueVH7/XEBvO6NpOwqUYv31tsFAdPhnW
9PsX8jfbTtDw3e10nfpHkf4k3aPSYLzSo0fhOABgCfsE/EgAwA1iQFom26oaeJDzzp83H5fwmGpp
6wdj3mtDLHdR44h4GJpa/oFcIrlisoTN7IrmtHPwJhCmv3Qnu29PH23wRehVMc9qQGOfxR3/0N/g
XCRmzmqXoUlAmtJpnYANxZTA7GnKwWfl6xBPtbzycRThhGCIlhCRVAEWv/UPDf8Wq+y8zDA09cjc
5e2BzJ+sc/W+/kGkdS85QBIkRrCX8QqL1OuLOGIgJ7MReEBIIw5nAC9FfZF/1Z3ixTqpPDP3g1B1
IL3dIdaZHEJ3HTARba2qPdCUoQAWB8g69Haq7mjUvYG5B4Z3PE1ms+mvFhTKPcao9+5DnTl7qcEJ
BkJlid67SSKcLnHllXOpZyzlkdx1DVcJodXb2xd/t1rS6o6LupnyoAKu/LT+NyH6HuZlDsSfuSRS
oAxDJxXG8aWHlc1tzXx4JmXqhUWLkEiIRZCYqU80T18rLax0O4F/HBRaVKSQGcuhJGj3dl6VJM56
FynCQzVAG0MKpRuIdGn6V5oeYVNbC1/TEeyrrTHH6bdNjAUSHOCryDFX1AM+7OOhwwlGeivNNFlI
pl95OD4Bgc6RSWqQpqgK2fWlCKMEeZ90259EpRrl9HIn1U1QgKyaku0U6goDQgYQIYu0tyO8umyK
2dFfSZRfzKBxR2XyDwNz/YlN+I370H07+3qAVzO0QuG6CBcn6hUuxrfVDhsy31B2231lkf+ULCBo
9tONmZx0Q6IMy4/zRji9JDt0txLlQhK4EnqUlv7LfgQU8rk7QtXE+DoFmLitYJMwDdmcVZT46OHE
RNERnkuasUz6xMVCgRY1rmbEw3HC136FL8ekxQha/pS8xSVMvbRJZqi9j3idFVZV4LbkFJEqYH0z
WNNUMMESqYg9xtWZ10KLN97V/84OYLvODM/nAy3IlV0kqEL9NiYiMx8EWRowwh7sAR+HozxEHFLn
kqmG8FlsK3ZGInHE0QgVAzOZTQSXrpwevxWygMRXOUwfTBXPsxkPGhfgKbaQr1EauB0cqiIEflKJ
p4gm/u80HBJt00onSDpdxfkubX8kcT58shIx9oqTnHa3H9xyW3X0++64+RZqPLOeou+v+i2ofXVV
Tv8XMeTz5C+HGJmHgzILv48K8Lvyi8X/rGBoVWf4IpEk9elQZZ0B0PhgRocleiQK/gVoUl+2JTHS
r73TlGXsJpniHRK5b48j9HfhUU/PNFjT/IG9wKdPHLoSn2YIX8CKDefmaA+vkDrxFVqH+QUPveb/
Ip//TELuc7r9G9FsRjxyl8ySbx9KDGQl5qkPymTcnQBG4OG9xAUyaZSfeyhjawRXk9crD+/Sh0PB
2KyfFSqxGRs+ZLf0auRiFVsZyS4UX9wre8Mm51eIU2zGkBWImtCwjzsuFjHT7SU0GqGLH0yYvv3P
0qxZovPmE/O2f39IDMdLIrJm6zCFlq9PTVLKAe78r6nS/B08CbYlo0kzFlnrHEmDKK3f8rm/kgCn
snIO6IQ0Su3vY7PCg77P9qCRJOj9vfDVP40c2U+TewvlwkTvlKcg+Xkly4bEpo3JhdpGylOP3lUI
i3Ix2/yCZdLw+3Ya5yuJXLSk0Rk4uAurT4ylnJwQdaxmymLrEsq8h31EKb0dhkgSgundbTAeJIsO
kV2F5Gcx5abM0PzI6ozoxzeT9DZCIlQ/0nxGCqpi0RxVJW5WxhabrTrk+yD6EOlqE7FKYZATIhwn
ijaDNv7/NAw4MQdr3u8aCDZk4IstCzEgfVKIKf81Wm4+UKm7sIQMe2WHhGU8W33/fx1fpPp0S9jf
8kt4NlI0AylgglE/VVlgJVkc62lXxwqtkn/ZcPo0g4GgI/HEFxRlEKWrf7lvQHncX0BZSfOz/U0l
OwALvgPMouzdv0cZpHApfbUd5Rgo3gKhbaoZR27A7TvXpZwz1D/YooaC7HjP08YxPPq7B4fdY99J
pyvSgbI4KX9xbLe/RrwJmlghO26rJ7fDC+q4Um2v/sINc86N2Z/R4/EYPsCJpBjhvhar/kdDpgpz
3ga81MjD+SXkzlXAjTCs1VBrZKvVdnljMI5jDG45hm4yaCp1fqesmVmgM0yc5sDTsn5ik83XeAL2
oVlxn781QQLeUkXePC+pjJcednUCkY4ZnAv5wyMHKEZDzRrlp0H5grLuI3mZhgybQ+E8IuTT8NCR
tyEIFIcv6sgTz5Xai4i2qmf+bMsgVMZpFuMX/MZopZlN2F45b4ap38xYbIPXqhdThNEMBMjj2WOm
2mGYVOc9foxs50ulCPOn07Q3WYvbhSMP9M65PdxhS8/igSeIxtEhP/d4lfdX0qif1cp2idg4BBWe
lRMuKZ1TtJPs5DBWEWPy6vuSoDhEA5rW87lwfve0qj24y4GknJvGvP8fNSM501TTMU7K3XIiKkBT
qPrJT0bNR4rI1S8w7BzZI2EQfkWKb54AmgPjesjl+7ZuUSs6OEy02SwPHKOsQp+/ZQ/x2+8RizMy
/pUtV3Vq630dK1hTaqAf2lGDZNsGoFjzHUAmYUnmVFG0d6NWuZcejPEWTi9QAAHG0VtH1KbnQM3O
FgllkLsmFBmwu0+eaU5ERHi3hfe7trquY23KJztHB/YiU8tH6Ju1VrLn75WA7gxpnSAhjLoRXYnH
OUHlaHCjEuL9Gixh6xNC1dRlbdO3+kqLjXuIF3ZUBNIDKcaOmC4RcoyBkHCpRWPlpSfzTS8zmB5C
LsHlIIBSnhnFWvcedyxDjMybzaNC7Rx94rq8t2cCaqrvc84m8YamrT7AGQXHJ3XtZrvm+vY4V+HH
LXbCsY66i6uMEI0aUIVk1qp/ixki7JZwf7xEZX/lzU0dF3fxqi1AAbe2Fy+6rR8gWHNKQjCEb+XY
DqxCC3XA9qtkjpkutSbPSS1gGM2b8MqHFo+mZn8AS78PPAoX7E9OAiF2nLJBQOZtyOBFPYUMO+nV
VGYeh3j3Xb9v9pAy+recLmxNPsI7GljhIHR4d/GaIBGu3GJz9TfGlsEQog+upi5D2w5SrrgDJY2k
Kw39ZrwsZjJJ0jcIeD9O0CLO4juh8n6l/irlgbd3ytnJtlBq+8hqF+wId3VhxvGCI2PEXrs1zpP/
1P2l4ZYxCkhMwkTtn09i5cSXgqH83LZRJVZpYTvIcnlopAFg/SrQdsS5yy6hHCC2TX6d+E1rbDZd
/id10yWdG6VCmt5GWxt8a26GsjC8puVXJDQu6+oqUoMJXi0COgxT65gI+4zHo2aiva0Hq1q9zkM1
juRdh8NsXshr838v2OagFWPtHMrdBhUOqXnG/gF4kixeAgiGNefCvqxXtrP/hnOD9fmUGoKkEBgB
vdEwapSWAh22pW3AjsFLrrudBTxAKPKAM5ygkcIig5/cO73VJbEl3fANeTp19IZVAjEQGvuTzEdv
aGiNa4EOhu2Nz1dRIpiGtmJBHCJNyMSH4fbK78gP4WtKQNgzzlIEMfR1StL7aidoFIMSEbf6mnv7
64bbC31tR3rR34Y5epSpKh0rf6Jq+BiheQ3HSJy0zYa0eWP7rB0jIQjb5Qe0UlgPrGWF+qq0hLIt
OQxRaANuVqx2BmSGRV8evGXcaGtAa1BNVkyRujOm7DboAo+gMFEcUq9BmcBbHBGl6d3XBJzLfdvs
NJUxQmQ7cM+2A0a+qzXJ/EWU90vhMLedI13HLP/R6lPYFkwMYAKo7zes/7vauNNIBoEUK835W/g9
RI2DokmXWa0HZUfz7cnjW3oRSZ5I1s5RyB+/mMJehSv/swmiOnkgaTD09FDF2Nqm/e73yThWB7w6
FKt185h75Eh9uqi25/Xdje8ka46IlgSWawMAtrllJCAR1NzLr5GqIB5Fqb5yXSODoP4oFztRfv2h
M978m4YsdrZyANrovu+GAr4f3DzHt2rT86O2OiNxagtpxdhTEVLA/FcKJfzoRTnMF/c3QOiSWXXf
UF8x9Czag+JfDLNStKMzmzvsXnyGaH48pC8XXEuY6JGDaVgypiCCR1d9G6zXgOoSK+aRkXi3AgBz
e8nFL+MoXKDbeCIVZCJARAuWuEAE3uIDNcQLFwfSZSGmpwBuFFv2P9NznhQ4UW1/UK08v7+Lwz6p
lOlr4jhWZwV7TT6d1ZvihxsSfWsXJkdXv6USuMInb93EPTY0jEV7u7IUpyR6edA/eT+5hFKexuEb
vbCFrN3azzOSt3c/Rf6qmaUXvofPrQejfmLxIVhGmgZzOS7ymsN+5PDEr5c49Hs3Xm2pb72xhPVh
i9yM9Yl0xOWPM+QZjfJwIMTZVIupmTm/RapTPMy//eWgunt+qzMIq1CyE6OdmUqxeVOeN7wSmQoL
I94jkXvtmY7X8csymmR6hdHP7Jfbx0dUZRXaajQzPAhfCbCPLWBoVl+bT75O7CvVBGEx9py1qzKO
6QSYGjT/P7p06s7UxxcPnmDz7ZD0QhNWRLPicgk83XYeMnVdpROQv/askTknj1LOb6S4A9pL0LOI
rgL9zoveKkdwJMS0Yb1/WyoPLZchxe9OJHG66h3MbnpjQUfpcJPshojdbFuToUUjze3I6yl9FT4T
8NZTeKP0U6ovRbAG6uD9X1AuuZXmL4eK4Zub8dyMpjyAGkiwLxPxb2EYxTZ0u5iM82a//DU3Kp5g
lQbi5SYvmRNoaBbsW0NsFXMSXQ8n9tK8a0M9FDE8jPQkR6uLFnrhV0i/Zv80LacGtSNv1QximfIT
Py10wjcmsNNOfbEFDEuPT42xv1LGOZqu0WCQrx4UEAU/mCG+kBrLMhGmlhtB2VZ+kiqgrYH+e+Gr
CwUM3ImCxjyrUY+Cu/uVPZNcrOf4QBTtoiZY5+01YoCBJNe3bCuUh432iTm0x8COL+pro02ViIvr
4aYrXygLsgNy6DtA4k2wvKOc4DfnZMy7KNEo8InR0ssVi6aAm6jLJxAoRYEaG3AFcIItTQ1SXCUj
Ld3Oqvoy8fhbidXcSa1yIBeKLSkk9RsFCy1NoBxyDiy9jksiDVZ47DNSVOfSM2i75iSdopt0cgHg
lgc7tCii0sYOrjCEVHcHhOmnuFDNNvHxncM7XwV/RM9994HXPWRTcAdvHrzJhnT0M6AS35b3B13f
+rkQc3lOaWe7ZgupwGayMK5UbqnifLAe082ulmdGgKkIMAENLnvGj8kNNm1OGyazNVUiCVzdXWvs
gtTxZ2WwmAVLt9ay5FuHuHVEFTgtiKPpIaUiTCqCRQ72XyBUKlq0uIvomlbN5fKOpQzQO2916LDF
SoopJEsKQkttvBsPFJxX7jTRZ4oGxXO0wyvD+1eN45tGF1CwOFuqq1/dnyzezqhAySIBc50YIEK4
jlHvsC/eDpy6Er3IPYHWLWIg4viGwUqG2632pmw6+90i/uNcB5Pk8dj9SLe2ODyy1CDJ8oqG3nEZ
28/OT/MyX1QBQtbu/jWKuZK7DtkHKAtAALOyD3PfbWgiwOpaLSveNGIGCySq5wUQTnZMu8VLBxjH
Sz+mu+ovDhr23KsRyQ4V3JtJF+EUkPxfVFB5nmeD7neEHSFJKnqVMTTqyEsUvTdY21Hitg4qzNXo
qgkFuqcRCYpb2y6zChDbBMIq9howwpUPBFlUzqQtHm/7VXKa4Tw3YPPitRD1dN5DoGeEnZZkcIT9
zBqNu5g1oc5I12EuMki1R/ABBmzNUOz2lzEcqdZejWckMW6iP7sBmSEJvg65MCFVS5+CNBFuawN/
YRjlqC6Ow2RRSUTyxHs0pY8EmLRWme/slwCMNA+3c45459xMLyOTc3tRJ05446EMo/4jbERCD/y+
o1aU+GxgjSKRjXsp8Z5YVfnnHmcwLawU0WiblQ6EL9CKlfQeGX3mOMTXOThSSBCyB5EtZv1QEMaW
/VqwrnQf/fujX06glihX6Q6nMV5j3fvsJMeskhGzd9vBKDZvEhLj2kQC590ZIqXO+mBbG5KCdJxy
K3tgEpAdD86sbZVV3jvhzqmnlFH4dlPS8z2acaknUdBKU2vIww9WoSdMY2CDPhephZK4Oxe7PPSZ
OcxT4S5dkJDTkxAt6uZa+ROPrcvAcJl/1lknDqp2EfMA2gWib87QSFMLSwbDYL7rxMwyH5Kl+ALs
uGLoIZfXCL4CFnNd9PGTzesQwoB+4nHamOijnupiz05V3NUVMGuUaC+QJyEYQUsGL6QzNDfcZcyt
u3Y/Ew0QkPUdKhKxt04BT2eKyAL+eQl/+wdZ6CxvKblzfTkHIuEUBwqpHLX1fiYAu/G1xn2w/HPo
J9KrYM0vXFryPB6rce8Am7JNqJpFVHyTrUb/5S6mvoC8hykcr9atQk+nZAIHX4c2M5GkEMeQ6eUJ
mADy9TO4WCDadfVxl2zTjTNxV9rwGVLz7+9m8QOJKveZzII8GoqeM8Xq6FNEPadTiC98iCOBJeLV
Y3NSotbJq3gLMxl66yTQvmxSnvyM8FwBJuU6jcWesDb2YUFRc0jtMvU710h45hZgLM0AigIJLpeS
HTxKFhqOMqCn1/Nv0aIAqH8UGeFrm9VBAOxzqm6cr52/y6ULnGPBBvUE7dH4C/rSxs1mgOcq4Pbn
i+ffy9KvmhYYVnDRqcdiq9S/a1bXNvs580ium2+xtJVmmI/PfTKqn7CkI6mP0lsATPFk7O+NoijW
YKtcmBj5IEKV6Z4W5lXUZysXptiP4eMINkbtrhstJ06gU70/GIYSJKmh15j7daeinWwtFYMz9dQb
hPMmLmgYPE6khGsU7IdBF7AEr7dsydDifdGXoA6UIfObhhZRS7iiGHZ2qrcAVR4lcN5+pDRZa8C5
8ySvRFe4LbOF5xfbWA901iXZDFHJDGrwt8qzfui3yx6+ObWmoIVARp/tMmz6gaYk9bVw/9IBPCOu
t9YVYFGbblv/82nuYu0LEaKxuTo9MTES8wZ6KHoEGlrnLqmVglqrcobvXHNxiRHoUdvSJ5fYo+KL
DgmYZpcv26J/3WInjsg39+2xGZBNUyd6py6kDD07piNir2sE3xEoOyYnKYVObMQyOx/JMTK92LMc
yirzJ7PLPe5Qar6R5lm2LpxSuC569WTW/lRx6EcYsWRStnYJq9FaQmnrYXusMnmUi+fvPbFppsYZ
IEejJ/p9AVYy8npOVI5qdXJvUN4ucoF1JlBg2ReznYW0G1EVRkItVjBJawcAxfvoWr37HUVTVcL2
Tk5G+iiS5S3pOefi++tapqlm1MkEJXkfkSKL/RvMWrbopfrnJCJHgXk/MMcH0ta4wKvk4ji8tTvw
bH1T1CiC7gZxUg4ohkX3rxgA57ajq/krrIDc6KrWTbSR9aXyy71XiCD8MSCPd0r8QzjuGfjQUG2A
waHD/3oxub2GALoP2XKY5E5Pd/1Wjw5UlaRDyrRnKxp5sMNVke0gpvIc52t0IvZ6EgwupteNurOk
Y42f0Jsxz+z3tBfiwC2StxvSY5VkTO75Wx30iv1hh9PJaZ7nIFTJsvlNpRvPJyFUkpMc21csypgq
apDFG0ZKdQbclGOOIU7O27veRrEwRBWghcqDmpjZ9oWmfDOtu2PmfjfUjeCZP8fLM7A0hKp6I+UQ
XgfE3Rr/xJR5Z23mnz9YKQ2sV3wMpZVRzMnZZHWVNyZCXPGV2e+Z3IsViteuSWhNgM8BoHl8XzcD
gT9OUldMqllEVII2piXjC8pCeQmtodxTpQs1vDQsd+NEuh8ckgKr4lin9VsiBkWgf93TnQIvWshh
HmgE5FN5JBjiySg4v0t3s43Es7qrvVS1BrCwxdHuD6iEJPRJIvtOklA9zgPd/Pwcep5kJL0QGNrj
W13A10p5ETzwZWDi+xLdSnZK/5lpw6kYzJWMmAvq4M2wQZGgb2heAehOVHHYiw4XxarnP1HxAat1
sG0LV6vDdp1iEFUqxHT78bavaXUHqa6kTg51YpDNf26ksgUFAGj3F04ACi4kv5WHcZxRDALj4lHp
cpZBfnJLbGVIUrsNr9IWKlGnRDiPK/Lr7wzjjcQkwLpATLYqoAxYQygfajpoIudcad8uqj4hEq0r
x+9cAIYm7mdCVD6VEPxMQBwvaPibhk69oFcw3EOgnxMxRB2nJhlKlwtu+0XQ9RlTYXngGxoP0prf
6iVmhOQzfoQHZS/E1YLm7aw8jUQTT+/FTIPwbUwRIFLZOaugc7CH5ZgXj5DO0Afa8pxaEkgz3WgX
CtAzDbfkIvqAqxRHfW6vmmS9axPGHuWaGJAZGeHaaU8GjLulp7RC+X1c+n7+uey9r/xFjcnSv3Nl
pDRA7wwMwoswm+S2O0FoXwc8db27PIdguOz15Ao2OOpFh1a1SXyHfDs4mWsOBCttBzU0VwXm7FtQ
BGbDvMeBY50GXDK32k3PUy1JZF1nKFQHKKkjDL05IRO8Tkc8SA4hPyDSvq6ZRaJvvCe2PI7H3Y7t
MdA+KyBKyEBuSAjgWuCrB9zhI6edxE/elWsL+ulnaF3/720Y/ebAO9FEf9x8DGj2DPk0tRdfgFlT
R9BrvIx4uP8xg7Q7phC6Eu4fgMvuxcHdG+xvPiiEoWjBN/fm/QBkRWAwvqMpHiVyi5bwVLDlq4VI
suhVXkqjBVfqao9tsxAB1m+z734jfHux/5Xw/R0tH3sWwvexJ+G+Og6/nMa/kZxTfApt5Fg/Luvw
0XuY+oYsSkOkQg8m3gtfHj5FjCSC8URxYBBOQWGJjOoRgyoXJB1MpzUFe5eV68AeBxfV0x/cTMMd
fw9jQlFwRZiqgNKkIbMrtDEjZnahMhBJTsKv1iZ55RkcSXxEL2Duv+bu5Q6xzA/ykk29/xA/8yoC
fmofkKO3dEFVbdzcEcH+NNDVFzUY9UVcTX60w476gX9iL1LEUks9nT2cqW9KFvYHc7xJ4ZyNy8D9
pZEB7icLNBilrhBbvMRp92AVM5Tt/Deg9UAY2k8t7ar9DnwTcbLTlWkppLYtpTzACynquDwB5OqF
6DSj3rmtzgwyeuX95vL/2dBTgbult0TTyKiay0UPyVf+B9q0N7g4o6G86r9kNeIEyPgMDI1W5hmX
MNFMMqOWUzpNHZwbG/wYSs3ldN941U+vllG/5T95B2dDShAx/mF1qC/2INA3xMbQcRodtT3OPDDz
YQRWlfH5XQGVZ/Mu8u+VwCyVMbf2aMj9uXDHiNYyIY8wHuVf72Tzf96XYz6BftTIYFYvjIEXCAdJ
QKLVQKMtXVXxu+2szPr+VabEc8JzZmHCtu1FDiKKVdhu30ck3HB750Ri/w6GC0uKPzr5NzHvPevA
FmgLaKRtPZamwpZPeMAx4JTnIaR5NxeQhbhMelIE8sdgV5dGhSM1GnAtpRokqqJ2tg89M9K43kvI
3efUzduMpg2Ghc+whoBtsxO7xEJxgjbRGOdcuPq6yXuKvPXwqnxQmRKks6NkVLlsrchDCB8oxL4g
b8mpeWrR/xZBQ+3+TL7NgmWCNNjxWGVupK3J5jKlVtwXmRbRkEBuYZu592ZEocDye0V0S4CIK2IK
XJhrOaftEVT8hkC5m3b8yQecZ8P0cXCyyUOWeKyElr7uZ1AK8xBaSTxO3zSMP9RjA0zAT0bYU+5C
gt5Hacaul2aIjd5ymHdNv4d8teOJzxVaZigNijV7OubNITV0urHhTvt1AcMend7rWa4ZwtW6I6CE
Rbg6+9+ch7+7Qa6l6hf03zZUnX85WJuWndw7XSSBprD3kt3dKG3DLxJUu47Ngbtzd8lt5qgwv3uN
ZGuvJqKMb/vEMww4vdfrQaFQ+YLg+xJYsk72MVlSOVEhqg0480uL6O6RwjiIboT7hG5r2fkVqdpY
4Fp3H5zp5Gpb7K/rdYJI9gd1k3ddRhYJqPe4S+l3/uZjdsNZoZScIAPkQCM3pYdW1EsVGHlhRSal
xRFkNgujqRJUt/SBH3CKvCT4wr4JDMEgxIeNZ4mldcCQHSRrX74W0CnEhp9+feDyuxiKiFd0NZyr
ACLz/cpM9ITFBJFG6XfRks3E2H+pRHdu7ejonEkoEvb0EOgQSYFmBRm0VeMp+Uxa1ALG0OSdm5/4
DQCZqwpxqvaky5wRlejk7mrV5fyJDWCAvevGZa2ltCVsEZg2awDpn5AFuPGRtOJSirHzzFB2Ny7L
bUJD3QZ3AOgsf1XOKnrCPmryP6/VsXeuXffZhgwJRx8hvhRKo0g+dJo+znk9bmRPHcvmThCSofe8
sTUjjhVzdIE/g2zzNo8k0OVpnbOiNP7Z3OIeUHJAp9M4O1Ktmz4w/VSaR0ELq8nMoUOMEl5CA5iX
UJNy2aTKVSTawfpoUk26CS1VHADBLhbo4Oen2gJ+H+fvb6IZYdshay6qyCeJhfra7puF5Jo/qPb9
cGiHtzUtibSDgVhSaaHl5AQZ53MjyGtxb8UWyxyweOnqeKPOL8WhUevGhl/miv/IEeJm68XoDei9
lz/tSoeEp65/HbiZ3x+os9kOKy2Hn5YwxfUOVJu+ZSTL73qPHN7ifw1eP2VckLlTRq+7hVb+Hb9j
BogHLvCO50A3+6240XrjxMSbJnSxu/t1t7VxTbRPMdf6U6BIzQAndCG2JClMoLqfCEoA17nJh2hI
hXhg1NBi3MlnbDf4XnErTwyniSQnesRVD5xVow1/VlMvdXU0P+tiqJNschmwpwgdS//xJw6LlUAN
LIndYP+0na8llpFvpvXt5sI4ri/uvrR+9Q9IUr7cfd6D+COEPp+A+F/I/EKeaMgpOvwzRISCWYNX
ZHMxyzXVyrVcpd6x6+K3kFBxf59jHNV4NN2KMS4ltHYztEusrFtjFIKhMr3rH0iCXqSaE27/ikZ1
To6vYaQLZlGbKLPTKqWSjfXBB6JA11cC2btvc/AfeKGWdjH1epsxn/zH/uQ9Vdus5AyJt6vlVY9U
/S8Onx3+gpm7XX8SDwwANOiJIwLQal0CaeIltvCRpL47zltGwyVxlzqkbigJzo2yUbdQUU83XpVv
Zek3m54MwaU5wjJYa0D0jzhDPcoYw9/+RVm6U3/HuLfxVnGBsZn6RfQS/pKoKQtE4s3Rpy497+VN
BYjW/je6IxrT9jMyzS+coCR+zwLd56JNjMNkpnnGhvI1wRP2tvfJ1vdB101ragCe46aex5yB65Vf
jZIW3i77Sn97xuYmRKDHfdz1rEyzWtBmFoJ1NUvG6r6aPsoAEflSzdD22iyPhl5ss2fcWBwP/zw8
acHFg2e9rpko8cqAkvYX3DuMWYes0Tp0agqaJLnN0GD7V8ZBLquLE2te2Cjm2ulP18ZJzwIrtUpC
PX5g+Rg5fujyRzuU1alEAUMJk22UEN/CvDhfPkyl5vuNZJKdNw1zfNNDEAyoYhv48GVnEho4O+Qj
/4yqS/RM3O+4yMnnz5Gshb9kJE4IBHdixOe+g5qJtVCwB0yihPfM2v5MW5pjjMYQdmkMaX21H7zg
1N38AZtbH6KTuYN82LZBkkRyQMzn6H1WU8Au5+L4JYVi/bUaVPSc555hM2xz9u9bU61/RFO2X8bD
RiwLVuHGuvlz0yQE2JmrrjTxVpt8v14WItOwdx2DaAR0Dh/8hdErvPcMr6JzFJtkLyx61O8vdtrJ
Xevi13gp7F9zce01RGanMxgMzAFp4bYY6kwfqO75Fnil+QrZBjX16lCHhCDP1RQraMrVHPSpO+Qn
FCkOh/TVKsqGHL/ePKEcgxLkst2zbSFm/kff031xyqVCKtUSZFKwGjl35gleyCobWlvWU0IWC23K
P3FnH78Qev8z8jo7S12fWbPDiCMmW2KJIFjXnwThd+NQW0RhLy32LP51x3XoHDpBjh/VQMXHuTZu
UwygrYlLSQFZoP8qOO17gI/MxO1PkuhxiNqXM5XXavA/HZN2wCptICKhvD0OEiCpPM7isfbzD1vf
LG9qNxewc4kgvb/cPJcycOx7sC/MT8fFnhN56dfIaV2YFxczuy/UPaMCS+sids6Kg0k1VgdqRm2a
kLYu137EtFuKNRTSbQx32uGp0/rFXXWmQLoL4RvZ70FDNSUhcL8g5RRbfT3T6v6gzLnFcYo6SOXQ
8TAK5eaFaa4ZbZTglO75qCbzc7Qyou2gFLoQj4iO5CeHAJt8DdKDIb3l26rcJPcYHj/6/BS/jHjW
96RrVCkdEMGttgTt8txGk6bFaQvX1NVWajDlxZ9PK+qkNEg2VbzrcrJ5zn7Ok2FT0kvECfCntQgp
CMXncZMOqRM0SZFyzVxinMm21bHh9CB9UB9dkLXZdANnpC8pLMcwBRT9S6LtiUjuA9objvCmVXM6
fJA85XZcRNDw4zwxzl8jtKB0Y8EMiqVHTqJduydJRlaWOFEGZL7w/hEp5ZI4fl4RbplAKbrPjMos
Wx7Db7yT+tavMJ1H+D3T7XQx2tCO0T4oxdoZj2+HFr6jJzTfSVfUrDkS2rR8Lf21bupHmIS3c8Io
ddIeWsBgiAcFE6dveDEIJJ28I2c13+iT/1aXKiGoW1Prmoz8TIfY8pag2R/vIi6NmE/lzv0JWhS/
Bce1E0/YP3ZaGFNpWk9j+At3qiZGi6EIqw8S62YhP4o8J84HVPuI2UEIwNzpkETP6I94jiSkk563
BRrRCPEg1Uga8xOwM8AyQxeFvf8U2e2G75IXeLtTddhAhCuTyp/Nbr6NT7t+ZV6UZO47sKm/JzwH
9v265wlpS+BkXcT/XQAtZ4394pncmumjW6FXvzAed5aGQ8wVXA2trMnQZLfb8DuMHqVZ+Qo/qZgp
xZLuvooxGrtuw6a6qeaWd5WVPlAuJ6VjjeRoBovH0On5308BwU26ABvafJ1M4vruIeVCY+ekv4A1
U2TAzoay3/jD2S4tMlH0jZQRS9MAbG5pfuSW07fgZh6TNwANI35PjGs7SWBOLxonUZRrQJrXVV2k
NvSGuH1cO6xHHpnPTEY7VLTVg65PrMT/95wp3BVzK04bfI1mLD9+BemnhvSUumhTIir/Q4yfLLAF
x1v8lsbGNADna2eVP1EuxDnw+d0e9P9rTxWHjVhqb3sNTKr61klS9itjS42fUvUqCU8LLt6nMkeb
dQxYBp8VmXnvLq26vYBAlAzk0kTfigivV6dLdGYT6zhj6SNm10gxKkwKevqgYbjYjkkYfR+rmEcz
tUK54tI6pddZ7fX5B4yGSp6hlhEnrJ1uRsvBBnKOVy1505dpTdJ/153gaoIIML3Z5iQGrmyXzcDM
zpGGk227t37l6FDEunepWEeExBBAilpVcFhMCQ7GJB4eAIRVD5S5JDJ/9bO4RGJetYqO3lsGvxtB
/vq1eTOVc6r+gWngTZJp49ImGWPEWIDThzxjf7+6zQSVy+e4fePhCANtKBW24iJo8ijEewJEdctI
iYT6AzqROj5A35UPlacPT4LAMxDJ+U6QQ6Jnhf9ux/o00sseT9FfHmvI51kqjLOiqVEDPD+kzzq3
uZJKDa5GmGp2BfnwJM0kDRXgtU1KKf83p71PPMMsa8euslVljDcZAb5QmOHfUW6Es9Ca+XrrEsMk
XLL+9TVHo7uzLO9c9PiXZtyGbQjKB6j6hgPWKE6MOjNpgIcEuu20E4B6LOOs5ZRXMVjPGkl1mJfz
6KURkmX5FsoI/yRd/wPoolb9Q3CXNqaNXHZAFQXork9OS85cZmvdyX+pnnUlSqXkn34+aVnJx3M1
MJHi3rtAg4jYvWaCHkqKFKe2bKnITVOYt7lZfhbDpr8qYz1Re+rs5MQE9VQXUrPfS/oliwr176HA
UMcGZc/xkSmz8UVQLNjJdpI+b2SAbHHQQ98QZptuwIZUMwZT6YR6s4MaFHtAt1P0QpBv+O31LW2v
NTjh8EqcH115SRhS4qu895ArRV/A4jHUeH77dTGQq+jAnBTTObvNaESI2DmLRWBvJRm9a54Xcvd+
e6+u/XgWFntbzIZQQBefpvRS8myYe7bZuym+WO8KGYzXYc6LPxhFkm10DjsYnKw/Y7xVt44ZY4bP
CYshMi0EZJ329qagDnZtUexGaVhY6eXcStI/VdarEtHKxJV+o+Sz2+IpjQo1nnbM2KYBoAb5d9tH
OOTIgXqnprgUh1w3hknH3ZP+NNZcUiioi9WMYL6AiP8s3toNlld+JUz87bXRaEEihrANgQx2pgJT
x2ku2fL8gsgBICi+Vz56ckMVjc00Fx10HhlpfpIMA5NrCLaiaARHTmD4BQF8WIpmMeXychicsG+z
Wyy9zAKHbuFwiyp1OXnnM5/O96xuC6r7PgcungI0hmQpzyoeQQHqZAVn5TrbeQLoYQehkGPYlj+Y
Zs9ArMI/X2sWX3UKyQ7Iey4StFscexipwr+YbSjOa8S2UAMkvW02POof8GYP04PYUGLd5tuMYbJW
U+4TfkmLLeZL/BHjZ2ovAA6a2PE8FhZPuMG9UIeSCUNpdc2doEl/AuAIMrjPwqjd1vIg5ZHAeLmh
KQnPYxYuY6N2RMpt7bttNDvHmTZGp9xRApkOgdARpqVwemhWysQN7xE1tPWJCowYKFNqwNHkYmlb
wlKLPW8Hz2Y5fwY6gWX8sFbbRT3IrWbZJzPhQxctUs8RCvqfkIsgFX6y3ePpXjComYX3DL4B+7mF
uQub9H/URm6UY1ByHx6eb5A7HOwXKzqf0WnQ23NKPpGMJ/RBRKGSE3sr98pkIf69pmqI71mHqSGx
I1QJA5+vUE8e6Y2E0De4/g/EEvUMO1zF4OfVietMdCExbsI9qk1RFg+WROnI/c9uQ2nbrH9+aFox
HfQIF/fY2RhaO1dJtUfMmcriizjGJVTp0iFkygoz0BYiQSqydWyem65ulHyXYK9azDeplqwZp9YB
Hy7eCKI/KfTx5gVHMR9N6e5r86oNbzw9UpKjJv2i8XWdiPObLaQgDb2YUI7ctKHx6cyJHAiGRcui
O1fZieMFn6xhyzikOkZkEzhhH4WFZ2zbll+mVbeK2PEIocEAwfhHPEP0azccOoi6bGXZuFGDOfGw
LuGrTvqZBm928T9ebvgCKgsSyVbDOX/cAZiWt8iiwA9O+VSMde5fHMADWaLO4b/S4d2a170Uov1r
KtQM1gSW/VyamMJs/IHUKqxdDh94Y8nLiIQ432OfQbZ8SyqiIP0vx6Eq9L27GKdbYCGDO2CGJsZt
Cv8joK6ARmBT38OQockxdQd8Q1z5PP+43HNzv80cGSI7Js7ddmmOC2JvuqEY7+ftGbqzHLBx5Of/
NNon7r2NJ0ze5BtowEcZdE74EwdKfrWXbNAoLRGrtUyindpMTRN8mAIWAeInbX4K0zaY4tn2GWdm
X3By+bC1QRxyPPE/2XyLtg4EbhQFP9UNMW6gjee5LwNTsG8GEYlHO+ihNScvTcIeNlYDpYywOIs0
vTRBaj/YSAvLfIpLlcgECAe8+Q5LpAQ1gfLSaNLJj+mj38vsKIxSqjYK517glenSsO1YmpS4Ib62
RCa3KpxVZlC74Tcg2F3hoozHy9A1OXopjgbdcOE86aGrkIwLWeZzYhpcfgoB80u8E3O9T6WmC0Jq
tkLdg280Cquwcy34lA5bsPXuAHRE1G5x7DlUNY8F0V4EQlByodJ8YFUBaMPlVxlJybNwY/V44Sw5
da+H15ExABVHrrjBSPMBX8JXXSGWw+B82M+0uYh3S6aBuON/7VbGKP19qp4z8x5/VAzVomduftW9
m8iyGYZJdwbFUnYqCsark78alYQY9IwDpSjIzugnL7zuqqcP9TBBh4G0oAuSfstH2nfZRngWpP5L
jhtAmroRwsKL/fPotCmTKkR+0t9kw9b1j/tc4KOv9JtoVzuqpVdCIvYK3l1zuyOlFv/Tf/aJMMRz
yqFkZdRSS9QnU15G6mrqcCHtljZ9NHptHqw9p8SoWvKz3EexTYr0FVV93CGSV2dQzbwb84kPSb7n
9c0l9ipbDf6ure2hhKwaSogzJJLL5oFmuORZ08C2Y5yFfCi8lKFPWj0XPo2+XbutpoFb08VrESgf
TUn6bGD4Z9GHFPK+d1/5AGNBCsalJhKOwffLso7sDnC4eqxSoKYvIcnyI8g/do6PXJdVnZAvXbmg
DRnpgM+nvduVfu7k+tx3fmuLKQZ9VAlL/H/6FBYn8B0IFZ6fQPdxIhtp9swi4nhICywiNn94Ek4r
HPGYCXUInjHlt1mxduDh6VymjbpGgZAAvoTON6Zdjr57f8BkZiScy9F40YlxbPlAOmzQns1i6L17
hxVNV2+7Xs9qS0pOZ/xFeFSKvAedHxaLinjez2Zh0KIqVvWb7vxla0xOhQvQmqPao5JWX7gZCcvV
2cz+FoeN0RjmywVfMu2O6sWSSQGdlszd3cECeS0YsUEPHpt1bqx0ZZJypWjidDZtBurMAlAXvYvs
3TwWSMYBxaAhwi3CRFdeXuWOkSoRves+MFxZgm39je9D1uPAl2My+dkHnzDx7xh9ze64A4hOojaz
QgwAwpQj4QGL1goZADSoNCu+56GfYOpvbGlwBfsUP4hlG6UHZ/wsb6LTC63d1XleBuCrAFJ4hMnJ
2bkTLxNyzi5Q/bDHpysP+PVYxUgLT97pbfx3S8ZnDCXiMHGLuiyivChdHrNfCJFwJ0YXoayAdYiB
6InGCSLwLfTWo9fSbJllBQBt5zHKcchHoNeT+Qz/O00al505r7jO7tNhBkr/TUzKV27KGQD9Rqf6
aSoKC71xWILI8n5ZNzffL7+EHaUFdh8uOjbOqBJCUAcbuwq+HVzw9Y4hIxZibv6VFvdfyO1wX3U7
vl65OMkwF8JmSd1NAYtMrDVZiQnl9FxrJN1DbMBOwzw3iwd9GZhDewkjQ1sontXIQ5DVXN/D5ymu
GDJHGrVCL/PaQ8zOq6uAdilwLKnPiDv/f5Yo7ZBjwRHq6gdORfEPYzgnF/d3tby6/NdKCATkOYlX
r4DUHH+b8kQWR6kxPA6YnKr6UaUc+vRRozJzHMU17I+TIOOCJxlxqvps5aZOauA1deVTN5QvUv8+
msuOsHGV62iJVe/JEYVXIH97tlXecXCBWX9w9QF2avTTQOeMVp6NFH6PIrwq54qfMDwSPM+63NaY
ggaAoj/bTEa8w2FL3BLwgbw+CjuoXGyFIf2hUEOsxyImtgxwCDcWzYpwdCqcXZpsQaD70KX5YJ5O
KL5vOqVQWIS0wuA419cIiCK3MmELwKJbjxrtXJwcP5erkEvNRGGw4oP4eNsL1EC3ZOsIFg4EVIA2
dH5fSNM9hwRZO7oEPV2qICTWkC0abCEqIEzZvRBnD/cumoZMg8tq7t7jJl+D7Gxpn105DMeUGc4M
olyaMya6NC8PXXJb0HuYyNUFVJDN600GUri0hJBk7t588EOvy64AFpSSP9CidNrxuzhMXqp8fqId
n2rKitv4olxqS1Z3lnvr5iS5pmI+aTybQoeRzo8Tf7n4/igciU3/rKu/d5tcE4ggS4vhTPhDNJu5
oZ0Q172o+zdrtbamrai9GAJPlqC9bZ/oFNrumKOMCfVYdUGy0cS4hh7L0lZAN+VulG61ZDwwMCoL
f+FgGH5fUAoepmpSTPmHICTdap0RrKX8b3ujyDu6GPWiMZ8wRb0zE/iUM2kI7CNj2goaPvMtMYj9
No/TVp/HKx8WHe7D4L+1N7lx9tloDan7sxv/IOKqYE2OetjQcg9N3dbnxd077mJBGZ/zD8b2L+pI
Kb6+DnFoJwW9/evgu38djGGrp8vC6xv9usrJy0G+j7fUvX0UG4qntwv3bNfaCqvUI+VTzCl4L81x
QBxuGWsU4ootDDGATV1y2+AmiggboA26QSQQQVMwzLaQZ6RVfKH6bQJPK1GRsw1/F8S9hTb8FKyj
R0+PmuxZOSkC7Cm1XSCErVsSh/SOvnG4KlOmzadSCrj2L8gRPHGsH0IILgeoU5YR6kkoGHqiSZQ4
GviXSDFh1aThCEJGpXOfiF94g2AxyvViL4ydW+t372DRnuXHIfLExuY1HbhJU5RnNBaRqzyLoDIC
dy8A6BZ0hxXuOr3NTCTiJ8rDU3/ApGWS/jLvG/557OfsrZPHM6zg50kUNX+dcTFCPrgYRtYFZSOl
LYo+qQVLvC+dCHIlgNymURNG4oh+SceqiUwa0ZPVJRFNBdNX0d91itcOxxQuL9k50AIAk/pqO8Sj
nJdzlFCcC7IIrMHe/qKwGF4pWU28F2S4H3Y6DzhlAxerMA6h37PS2EbN/m989GVX42t4Oe9l+uY/
jaHJFqltqRX/3A6yQzvZo3fdquWkWd8xXhq4FZejwqGO90X4UDsTFf5hxDEZ0pErZZSQPLlnrQRc
n16zWihJCcZZOjhveUSpC+aT5Eujpe1OWnL/hYe1Romtebx9Qw292wB13IHXrDOk/m4/2rFRwRqf
Epm8i/NWF870AByE4xDP5Zv9RJ0wI+ft6HKyfqkvqz/HdchT+8qGveTMd1l8mD7HTnSDrJTdjIRG
5rt4XUGwLF+TsuLdIPriVYAuG87kHshzA7G0KeRQfLS1iQidCfNvK4ah05HWE65Jhg85O1NNriAt
Tw8vd1Q4ftXyT09aUyZvuVwkrgnuOikzYMJP0q7WUB8vrv+Tgd/7Bxb4DJCoHiEElhUqML2CjXma
6I4gP9GuArpbLFiCNQll7pkIvORX/0bts8llm2mg52vFzjTaiPqt2ShrlHMnDY7ZkA3TCF1aJKR8
IwtQPzUS97n6jGnWQgr230nsCSb54YPtdoa78uIARRqRh1xp3SKhTJa7CeRRPkii+bj/an7Vkp0I
WcfhMVBgBiSpe4Lp27vm3K8NnkE/TVMSDuifk1aGFv1dLCsG6bvcDmf1GaFYiPPOcJpnJX4x0c33
JE47J9C7s19vvriJLcozyVbXmRh2ODfH+yOYG80/pNr8AaU3DJn/UPBKNtHNl5/4TqIoIkEk1EPD
byF2VDtjOwIQx02uE6jJKkfoxDWbmHhp1u5y8wnHlzwVPYipsj3Vmsmm/8mBKcNRcce628LiqzAb
iqmmYoy1tqGbyCJiRj0OkjElZtAqz1rKLaNp6gbSj0XVTZH03vSe+YbW95LcZs4Ry4T2WQsrKkGv
TaxDMOSlMaWm3/SOQtX14vWdFr3Ma4bbkrE6RX1XCL4XmW36QZGrHfO+ID5+dEdQ/OXDWavDmcfB
RrsnJcqVD2yDFZUAw77CZ0t9skeEeyEMqa95MnEIe7/XRdXNkJach5PnsIi/AgMWV/3xbVAT6s1N
/7AvUEYoVh1UiIHs+PmbJyXsCwGKcDk1iR0wECsNUjYz20VuyGPKsy7ZvOxaSFIf7/m8Owr5xwqM
SmWDzfrMdNIubPZ+MmireqblAwAFCrVFPmhh9+OrEnGg7X1lfY16EttbZ08/1RsywCwyp0bFdBc2
CryOKZK9PO1l5SXZhF10SFOfIVZeQTuvdHMCLo7vu2Wzvm4ynI3i0a2UTwVBH1y7aDfy30hvPb+e
GwAwyAKE8tytSO3HjUiDTyaeqI/whJ0BRAseiiXxYOnAeVAAL3WDRWaBRQFi2Svj1lhAAPSTnBQs
D7+984nlYnCOcyuVDPS23C0icRbPJmsMgBFbslCWP05hjvdu9bC5WShWktZ0VoQXq/JJHHHFOrbl
ebPoDy1QTLxj0jedXixxuOjhKVbwAT0E8dPO/DKgmIUVfiG79b6GSxtjzJo8M7DLslpukuOHsU4z
4JIWso07EyKembsRZwl8XSwemubEzha/WExbPd/Ou1tzA1zWUVNJ6Y+/nGLjWWiIGnjR8z62REHh
6oJsC0AXkHg6SX3yhhPvRvQhvczERL6xXI8Zyne8iM0XhQIf/U0edMsie3l8pngRv1LC/CHfub7o
jMnHY/gRsr4yzns5Sb3Q4bjdJ1Hq6Itxkoa4AZG85CcGxmejElLUsHSc6+Vu+erM/K489LlhunOl
CUu71DPcf5bF2tvGttqhUFG+0ku5KqvVtGqQDH9DxYdjZBgRpa0iw6+K6B+cbkcfYOKgRyosTDCJ
aHVJPI9vye3B6VwTZAOWgZ4F8DnAefBtcfO8pqNtnsEJFuOW+PYySihHb6S9uJ04ivu7LyZks8UK
inhSrptsSSmj9/vToG59CtdsZ10+VLAY9opejGDiU2TvtRr7XY/1SK+1eeOTLl3aJtixlKAGt3w5
dqzBnuABNuZH4CVAoK+yZWy6VDjjaOPPYg8PJuG1rgzXOXQmaGowgH1UfE9MW+f+mB0k0MvBJ1Qe
dFVslKGlF713wrsAsECSNtmQ1GljXbSu1kA6bumEzvMJvTjXv9i14z9zEn273J7GaWveCupdJvEu
uQnwvRnq6gN9HU20Gf43Bmh67rqFGgQKNfxb8vENh0LGnmoSQ3wRUmXwV9NRkDQR7abKnD9b5Lan
gFr52G+UpdCBGekhq3S413I/UovssyIGMnHi6jyxQR+9HHD5mvS8NspeiX/V6kx7CpbMpqY1/Pn+
aIxCb+Bl6OX+nlc0pH1nMUuQU1PvCOeydijSeobOK7ozCA9XXv15WV0rmNXNZnQqYSUD/kSy4NlR
IPrYdZ5AubIFLnVHWI+gOfwrpnD2oFBi69EdDavhpSddfeD9jItKhZ0ueC3M12FxtuHVN5j/f7tV
YzNHgXFYO1riJVf7moL4htvH+hKsY/1c7cGt/o5JCzdJb098yTk+Dd9FCL1jlo3kY4Hp2cL0C9+L
GYv7iKnvYQGJax/w8wbt2k/muckrOfyfWZt1RIxqD61qXakc7PUGxbNTwDEK1yJxyBWfSW3AG9v0
eGNohk8EAYY4t1+Hkt4KlqDCpA58t0Ak8ZN5ZcxKBA6YlVT69NxNhDGPo8dLSVXdMs2dYWdh6n4D
9CeWU5lrLLtjTsZoWt431GYR8r5u5QNjGvkRSKiob/GC12fPRJOnZL/Q2GXbXt5QHO14efp9Nz2J
meKcGL2NEpba08WcqwFikJEdzzgOyNEZ2W29rlPBuplvMkC5lzFclg2QpFVDdAHV+Iy6EOcX7HKO
bm3mrPN5S3sVLG+cQJox4NY0b+cMLnCk7Rk9SdW/pvMKTIvRW5mfIx1s4/6saRAzn/lQaSEFrJCY
b1xnhm4cR4Iz4fcfewJCN8uLUeivBYENq8CwsP+QsKlxpGM9GWv4bvckOcWaozerRquKCowji0dS
6VMzBfItkDGTOdiKh0ErIDNNBGskFm4p1gqRAY6WTYxoy3ML1C9X8vRWFbG31Ltq/uZH1txuuSO4
coRZ4b95q15zNCGBXSqUyLO3ayIdlogIQv3tJF7pM36LUMYqApLHz4BalIf2QaXUQ5TbMgflQBtP
RQxf40ADIFcexgPQQWmJwG2gwEhqi2AKOSgGwnHVQ1sBN9joGAQAaSZ27ag1pZdxornZk9W0hyy6
9mDvy7ZnrYfVtQJ+YzdJtaQi/FFjFdvZie9BkKnrUOlTiAEUhUo2m9wV/eAzm8DitLM6rYkm66ik
8ne6gGkzZXExt0kJbvGzZiTafuCHx0g9Cty/OZM2Pei2VXHIUO8Eey+yDG7PGtu+EykqKPIBny8z
cqKtGJVMlkUCGhyN/5nBbd2kEZLGcfsjnQjohHDvy83ZmdtLviSEipT54rnoxizbs9in5zOTX9Iz
g9sXG4OB1X8EO6mq9TjOf+q1aZS4jKICNLFinIEM/xbgtv/hyybCs8V+wRt4Qk1u27DqamEjpV3a
7jQ88vH1QEjU1S+t3xl+7NxhZMcHiisbG/FZIUIrt7LABHTlIcurlFyd8rerxwwZHqOqN2G/MQzk
BugDe7bCtWiNfXrmWcyiD8B2hH/0MxJ6SYbr7MU8lf7u1sVpKPp3Uw1HOm3df0mqYNXet0qpcKe/
WpZ89YBrHEprGQo7YoBrmbRh9SRD+8JppR2VQKQ0Gruueth10dHQt0p2jYZkJPKNxDsQgvQNXIvk
iPiaN3e+/PAXWUJ49ygpjLtFBeHLs6Yvy00VlglG0orrva3sC1P0BKqsyYHayKb1008XsmoPVQcn
OQu2lOqIqy7L1hi8qQN9tdXsMRsYnHfwToUlrlWtzw1sqFha0kir2XNjh0Vwy1kE++kfT0STQ5/r
EBAdNsc8Kb8ZFjn05p2Q0DpHtX4x01p58kDAJJNm23JGNudccHSlX0D1LQxemVJUiHvi2JphAR/v
plqtK7TFqKt66FXWQo8y3KGld6SShyijiAkBwsDnN5yrbXHqQhi2w0hACa/JDqFdkJ5oGchLCRO3
qYfuEadqcqSamEg2qegZSFnxx/PIwufk9+3uv1jHmS1vH18DT9O53NUK1/mVpvusNw3W4gHn1+KB
28rkhmKvp7e1xa3/uUd7KCmXKtcjbQ0eqq3mJAkFMCKGvMAqqvD5K/heRaU9DPLUDcfQijK5DE48
rMl8GUnDkD0nut/hqVkhAEf/sw3SZwbwGyOY98QiU8pZk2pXsmKEJJaieaCFiu4i/nBDXpeY8dxZ
+j3Cnpds9gclXb2YeDppi5EyuyyX1c2wbcfIoT+vABg10+qeoN6GHNgZXzn0R0Aw+/AkvOoMKXQO
ghP1Wzh4xUzK53BzndTsY7r+kIJ8ZnUE96GU2mJqPXbvgFlbhHWctaUihlUW39jvSSFARvn6PuDQ
lHOP8u/WLDe0dJnWL/6CyfEfZYRDhhyOjbzhbcWzcCyFa3jXmZddEDcjj+SbtOuXbr0A9Wb0ynn+
l8R/Pwtx1CxUh4OA7HomDHHUzpvzhETCLFS9Mne4NTYjhEM6SCpxFEhsBmLJYHL9Ee0V3iEwpsLv
Dh2/qev4o+HB7ji+xXPcc9quXALLEPtDyPAC1KEGexVA5WuiyEEe6sKpOAtxgX8ky3w6iRvQfaO3
2DI6AKP4GhDVnj/XE3HSBnNSJm+p131o00LF3AXn8mGKLo49w9XXNMs4NAU/Q8t8oa07hh+3cLon
V65sFSIySEWwMFPMWVrzM4mX3UX3KzvelYpxdxByXJ0ZXqhFjxVUBvyR5BMddlEOmGbC6P38cuz8
Tw3jIIvThpu3LYFQLwgldjcImeAkG9Ee46fNijlfC7tATYgmWvm2VPmumgNHb6zSgnrm8NiomMi2
/hEhzIbEiAoFT1bix3FHAHSHDzo8eqaNXNpj5AY/NjzebfgtrhPrNclmyjrnqH1UpE8EBzZ46WEG
+t+ew4ciabWfxWoi6X6BaS0TYUQMy73kjuqxrO4Iwp81SKXYTCwRNAscIKTpPtsQjGFDa7Xvs1z0
tV1mGpOjLAvmAvVuL5F2hn592uJ9PgPev25kzs1WV5w9H7oOQzAQIrI9YfTaZ94nY9bj93L/yWn3
jx+flEWeYbrIVBEpv9CXUTHK5g9uZ6GJMKZpeXwWOklexPjvsulUXsfNg70CK/d9R2yWkP2yUHmZ
tVn3fuWitrBrCeD7ZiSvqpeGKSA6eO4HZQQSvichI69JCDY1R+3XoAj7mLTtTbCziDnZAQzNxZwC
KffQdyYKvz0bU8/U1EBG7forf52M45fD3jKwHAfscULT6bKivFAxWrrJSiMtEh4Hy0a7WGhGHkLo
vFbRsx/XKFky54fKaywqqUACIr+vh+dXN8N7TAebmITtIwDDmyxqPMB5wbS6NgbIYa/Cxjz1XfBN
3opMC5AKwafU7Me+qFJ1bfDmDKm+vAgmkjfr2t6XeEzwzFpr7NQWP0zmhnAcVlcV9lSzb62p57Yc
cqL6RLTlpouGwnG82vlgCQ+HF3nLIO18nHtSBWwy4v/LWWwlMacPGOeU9Y1uyEvctmr19HGVJaSM
3E8h+y3rJW+rATN9nWGgHq56yXtGoiVJbCy/RTiK8NL+A82GipS8grk6+/KVRT7BbZZaqrubTaOY
7S2rF9qrOP9JD9jPqN2FQ8jDQ8+IqllmhL1qxqc/Ht9yNd8HBkWeljHPmyItiBFs+nv2HTCiLmeP
f4UEmRjBggoYu4QC2HwdmA9uu8obKbwbpMBrV4bAYwqg9Lu2O1BgS7Iag3anSk68Qm4j5F/ay3oU
ntrozOAzV+ou2nYxcgxR9oTFbEQXiaFhr8l43jLMnhQysdrHEYrL3mw8BTpmp3pajye48GOvedAh
hBl7KpVTM83MIvivXn48mC8bE/xDhzczkkmPEvcbyApLz47wEWRr0l+ZXS9qWo85sakoIzi/Jwpf
DVN4S2gIDIYVqpZWcaUThmpopqy8SNrx/0WUxQ2NmiyU18eZpSrQfq+hJQtRPgDENkFEd4sBOBIX
TKA/ZdkHDFYs2ABtADcR6MBgAvnjPX4xlPKDSRpLfHKDFlk/xoJmf3pxetAwKlUHNBxdSkBr3u0/
3On3qBV4x0jWSZGGOqSOnQQKpASjPGk3y+WQ8IDAcDXcP8XtildLxMaJ2FOtsGMz5QapvNLUvAho
cSbwVRouIFCjE07TC7S5EfV1dnLzphw/YIp7fzIWrFR3s7O+z51EuNwdJqraSNdTbvnaJUv8rCIi
RSolo9uYPcLj9wFZX8RWhV/en59bJaSAyQXDVmQAzw5IYOujaw3gn9xfsVG8sQZu3upZ6q98lNXa
FVDQwQKjWM2/sEwKFTmifaAsxm1U/jPlt4caXVqRNi1FVXrNnym4i06N1DycHgBq7EJXczF+uqaH
TWPYgI1elnaZVwwlnxDiIrSHvJdW8YdQHOsFNSY+uPOeF8XvIgVTa2fnfEkaGRwwETN3uN70nBr6
KJxUlDcWaaqrAViYhjJnt+QiHf59rHtgXtKn5128oKKHoZFOaZtOquB5Z6BYgHhaGWsk1foqKTAA
+/pS9RQp1c3CcrD8Azhs8DQmkTsHGTEP3UCXDxZeOGIEEU6k6nr0cjP+/4TBVVeH37rZQ9Q+Pzx6
HD/H3nbRJzfAiBC0UXrKwyroySin84ZawDSCuWU1755c39jhRYn4eUIETuSmKYcHtTHPI3t3uShX
n9fMH4XjVVHP+NwJMQJzy2W8djGEbqresj5lRcbgzJ7qmhIwF4TLBHaotzKFNYvdmqMSaAp+jHBR
dw5Nk2IdHRw26XMWuuBEv8hQwiWq5tuEipd3DHRWIYsi5SNHLpuNQFjLs8MCXGc/q7cfEJru1N6V
+K1DtXAc4Bsozgt24Rxsz+WBhy7FUzqKVpnRX8Xdq2wNcSDuuVlXBr+YwEyEYffBPRuntUocGdNo
EFHcpIelS7j6EQkXE7G683Uo9NYg5PxesV9PexLZiHR9xAeRbbnTOxI6zeQbn7KmZg2Pg+3akszq
r7HkAYn3Pi2cVvb6771Id6rSl57L34bZFyfn7zxW9ayTG6Jb1HHTJqVENEFm+48oRP75B7KYdsaZ
ZQg43Lwwz03y6zkua2nVfIr7ad3yP52w/E0ONGkpjlOb7mux8+NqlUliP01x9GS1w2y3I5mw1wvL
zM40yZNHkpjwzS79Y4dlgL00VfbGW/8sCab+amJfmzkztgrOxvb+VmK+sW7Oad8mEhWA1srjkw7f
15nSHJ74yB/XOUksaLgdKyH1N2iYP1wLoxUOP32uxi+l7ZEx3JD3XNEXDzvCUNihETTYbJCPIPDC
skF+DTmnXylCbFufLpwXcyjnk7NMtlqfm3D2OyfgkjgUL1AgG4rwsr9DwB8MnT8aDIXFjMc1+4L0
vcuA2WUiqtTklzkq3XCQoF91+F54uoreTJht9td2CDQPKGDwm4QHIXF8583XWt/j7AqKz75VIZpT
B6FuzXOSllO/jU4iOw5VyrDnElZ9HtbybGOSfB0+Y9PL0Fm6titJitMLCnc3rYX7x3uHZ7CbVweW
V8gA6lmb6O8F5Unea518KdfkuJyzGbKnKL1r2wZP+k4oC+kDtSxGRM6M+6QuGaFlWVkYlRP0ldCM
6QgS4sIBHV5FSd8slkdZSchjlMjp+5Lp1X0ebkK9NmY+FD0dtDwkcxrY/CPj7nstHsD8JEbadZSH
HfFsfOpcP0xPHMO5AO9bEQk1uN/G+wUpe7lqY9Z/CFfuYd1MV5EbvbVzDQy4BsJIAl7QBG99vEx6
2hCcHhOaQ4lwz7giAiscDe4i9WZRPAGbc+jjvSLknAINROMLJ87vMh/2NqmlJyumpRGFmUVc6R/u
lEJocym9Qn+xMfRuk8JAJ7g0wfQm1XuEsCqaKCTvou57k70emsr2EvkKLs9aIw1rdDh1cnPd0Ros
Xd+Ge8KgFOr/j4r0nvlZHKxqxJkc74WlfimhBSWAQqhHra30FV3PWyHPzXxOvAEhBUidzLHKUt3B
uyioD0RR171XEjm4rLJcSwSnxwtHJe/Z4l/WkKg+9grdXkFZQKuZzyXg4fvg7tI7riIbhwxtvk5K
Er4w1zNPCnNRfyGh5yRxZma9mC+JDKdu46sn390SPN3itqNeLccI4nulufPHn9gUZEOB/XxGp8yZ
6dxvCfDd0ETEpLNtUZbl8MQUGd8FLnrqpj3xXU4bF9FDkkllCexq4wgopwrQDltpmYd//9A0ZJwd
FsZRRp35qQpSAT0m0nogIt0UGmrZGbgGGQfVhBgtyrfaYNS6uz8jzmghZMyZ/h6F/3sGBZH76NJC
Zym0DAvLPgV+9fFvm8izHoh3qZ50beMnCNXKyp9HWHUNSCL/gm13XWVSXwVNu4M9nuXHp2jdbTSw
wHVgufRP7Z5N1xCB4NvF5KYIy3oeR3C1xZPd9acnHGOtYe9YYjgS8hTB58rpKNCWILRRz3kXIb+w
Z288TkHJXxhcqCiTaLOFEy1kTsM4UdRtoE0yooo0U19RqRWFa0TedDczrcEmAoVD9MOl9YnWj1EC
0NnN9f8j6X2sTw78F/TDjkrDYLbOUC7uwudWIy7q+6oos2xkn6RtZNwY5O465xvI94dIgoumfF9h
bYrg9/do6FAkHAEZJkn5yinY7Oo8yXh7gesCDKLghmZ7UqIQeNKbhyf8KRrFWBinMqTx52W5noph
zRfG46oneUcstLfM3X5AGjjSqXBkirG1WF/UOFINKCIs9viWVX3v3Q1Zgo7A+ZEbx36cTPFi7wzp
tHZzYGfMvC/4eJTWiLdBK0+v/TtPRWEriHVZI1skmDNgiWjZvF3JwdIsGTky0oV4uSrPnRsHdBd8
qIT0YcjBKcjnBZWXJCCbNcoA+y0luMgFNcIclgjfm9u4WadoWewytGwuvjDT1D91V5qRTWsNpnx4
7DHPoa26MGkb7/KtV0Q5QoTM5HQCqdSbyIcmtHv9KldTxNfGht5qy94I0E2Rcb+gBOqxEnW62GEA
W92lxpnklUoo1SuaRWeHg0WM135OIE/pvqqHhfwozJ8OO3b0Ss7vqC5q4ry4r+Rn421oOO1kMlY0
iAXANM0KCts2iT9CkZ5QYTBWM+iQoTt7MxwP3Kirao2UcnTbdTjKTsRvcNRvKAyXbog7mIz3psHl
YWmLPPI+btJZ/wIMYChR8zE43winDHLS54T9/uamOFsv/t5e2JmdjyOv9jkT9P7fY3R/e+fVkTcO
lGL0agmJ001XWshNTgAyfNcDqu9ekC8qlLZMGdx6L0MxEtfgY0WMNJTQ3B+KOAT3HP+klYIWuiUr
0TdTP01S2jX8+kSrGVSnbtVNvxcRWVQaodDi5uXdqHfcxu7mSuO2EBT9usqdC8a7p+rT8bIqLVN+
qmRBaGBf9xMkITNAp6fYZGKWN6GxKZFwljt4rUm1q3LaH833M5wn09WLiY6sXQQMFRwd4P/KaaU4
ylFFuQDfgXQe3VNCdPOVcUiSNeU0Js0Kx7m42b9yeegtLdoz7VbEjuP7ZAXy19PtfV0e5OXDG6x2
4GYPrZMUuxeMhgqDENw3VAbz8/VyhLwUZZpCvEPGmkp3VXwx5hD3kqApJPs/lYyPGl9u2LyKEkck
0gL8x/AbELlKFW6lWRSZsJTuxEE7E0UYCJ3D2505A8Q79twxQcUkdstwX/TlsDX0Cll84cWlv+Hj
xcoa4khygZBLHstHCNyqtR5J85VJwnhAP6M2oyz7EQxM0Ih/sOEc/x+TNybASGFKA4zGM/kj34+7
qfPi+o8BkFeJXV4VGiyRW9JpNCE/14zJ0YfmsEgkIJoinNHRBV+jCTQijMuNBuuRUy7h3p7wT9O7
K41OlBJiPPpLdGV7zH82B3yJhbn68vCjh3RW5TOFtnLu5ngCw0vSmy24p7jkjLcMPVVS+hw2TYTa
cuNBHxVI5rmlJ8D99Gw6Z7i3v+gVaZh3LvXKzCm1M526nt0oKQX9CGA1mGKozga0POKt1upcs+sq
BjwbOYQNiffKZG8OQkKCmdGs8Gjr+1ILnF7IT4rkwGO7vVg0yMayGy4p66sXrrD011DWzIZPvAQ+
ldNmsvW9y2rSJ5xQyUq96CtWLRHIL2yfQmp0Fqty9nZxqZVHO3rnQKgPPHZ415AigLZQbofzMTJC
fS5MGmm2G3h4U7bw1GiVVLWgj91rpRiZhFUo5ftGC98zXVQac74VI5OJ6eyAQU4pjP6/YKWBLXSt
T1vG1yL+crVokgyP2UpFM3hQpnUFs7aqrRoj9EY/0m4Dhon2zSnaBkToy+mxSsYBimZnsV4qTwG+
coUpaQv4y+mslLMyzeYmeiaY72zZucUljg+dbIAhA2aIEGRiU/AP2ZIjjWn45U4pNMtykeYMC2Fr
eBeRq1wO6mMM70xMEgyOB+1Rx2dXpxnZag5JW7h+Xle0At4fWC8nz++uAtZyR37dGR8ifLGLRgn9
wyADwWqKT+tpW9R2HRmZdoAADtDEs019rdqFqpKL2uiKthygRbIYQAbC31Y0XNxzvguAdGJUMCNT
4oxBRFipeRwdeD6ka9Ypy3aKP8HhU9wLRrYoiDlsXhjBq52qS4ezP38Y8/1CW0omDCYZDZTuU5Qr
vngQyXboeQqojHTjSHfUmaEVZMpWgo90JHUPnKvNeaztoav/c5A4gfEoVj5NsMSpXKOYeZuuD6c5
NZse01TxQ3aRIcHJtLFbOSBqRlKT0VbKqkaxYAEYy/0MBzjDcBVnujTIgokI7BQNCISMq04O4aZd
WEmuv1wG3PWASPraXr1RtSgLfYh0xwGwMh8zfRm+4lKYIHUaF4489hj5GCDm4VweLJYqw2RId6yF
l2gwZJndRZencrc+PtjI06Xo6FQrevBgfIW+HOixXzzapQP/hxmNDkk/p46C4dXGhyM8b1kbI7xe
oQO0Qm+BX5fSvlDv4mAH2mjYmq+3LleDXJu35MRBMFYTeDUv7C3fx3FUllVcW6WjhSVU+gLxRI8v
iWIdAfPSi2db57M6bV0H0eodrX0EjyQ8o5p4QwAmhbkesr2xKctqtIQ3qdEbYe8cw245cTXI1PCn
8Hg/aXmiTota3qk9vfZw4ndJzhdAsgSWKU01KhLwXZMe4urd4BxxTSB63ZekG7aJ6YDOuhP4OS2O
GLt6WTtOvsqYtXaZXVDqrLTZ63qxcsqkePUWxE8K3kGw+sGdtTX9ckIGnaX8bXwB+qj9BAN7ids4
ocxBrACCLsyzp73nD74yQSS0W8EGIjvHtgKOXDWU0LOHl6NRX2MPb3ItoC6rpFb/9btOV6iVjDzM
jIUV0R1VX9Uof9O9DhI9IFPQTgy2yGUjP5K6K0TZ6vsWtwPiTgcqKZcrVop6k0giMKN4xylE9aFP
Lb2a3N+DHW0PIf/mIW34W81MO/mH9bXgl89V3uxhp6wSwy7tKOHKfe0zyJo6vnJpv3+ZKKLPWqWr
l3WZ+Iy9/A7YgyiwPRO86DhW2QmvbDcSfqiJx2yc9I5sDIPyZtyl5znbeOZ+1RqgzpByH+UbivdL
qe19FS0mLc2eI7rUix+degPC1vsSKIz4Ql3v3I8qlSRNuTqyRPW+7m4q62ei0kBij419Yo/WgYSb
fRDK108eBVXOBI1EP4qJoX4db0KvIookUk4jGyKAZh8wmlD0TZTLShOahMo0vE3ufQymEam6Flwv
uS7DcKtA/Etq++pz/0EdfdnHU9JLOOgQc8jX6rZxlOazCLFgr5xhHXPiBgGgV+xvcv0JTKO9igcg
E2HieBYbc5zrTlSUd0dAA7IDM5o8CkHiscDixINu0AMHEBX7euboT5uhEmyLWE1qxI+6Kt+Zj9f9
AYHkTsbOMIY+kbiP4qlL/RNk3Z6FZnrskb8gTvqZ6INcI4QzIur1/Isx1rsXRgcmIxzNEbxuZudL
vz0itmFk2rsfqqHn854HiVaiPLkrD+4yLiUMtLOkR2VSwfMSamuKsw/xR61kJjdyKaOTZNLXvgtT
Qjw7jiD4D3/Wzyx2XENosN8AEKcgXZC8mIAppojLrluOJiskp1+4s+k/Wk3Z+cp3Yaa/RGKQ+Xyn
Veqk7ZlHoUiqMQUh5miMYaX7YmAQD+QYaK/uAKI5NfnvjYDS7zlmOJb2tXuRHXfySHb/J8vbJxda
5Cnddj4oJ9/25pREyEj0hHG4jdViz1enJk52vDm+qGHf+9QzH5Q8FFYIuIO8jeg6SYcEAJQOxcXb
PuYxe+Hja/a6NXvkZIpV0xoGIg3BUUcEZlP2xv5Y40KlxVo2+EavYmkbfyiLCvFKWVZJc8xcMfhq
JZ2PACNE5GcksH3d5BxawvibN3Z5Op7UJyTcXEcvZDavNmF/SrQ4navU8dVdf0lTtPEFEy4Bkc4K
5Q9yQ5awlVVQ1NYeuePpstVyP/BPSqZzr+xGoOMnyq/gQn0PIFcU+Vl4xuLK75517Dt5F5Pz0rOg
ImRqGJK+55TdWMzHFyfrfoa8kCaFFJLKQ9FBA5Nv+t4YBaBidsgw9nxPa+BsuUEDN541wYx3ZE0d
KQ46sIChjmK8/rhDyHvq/HIgKreRGNlOoljapOR5HmbpMdQT0ERvEqAfTexKOKgBdjoa1pS10Rtf
UMGRIfBaY7NeIQUfD43wBYZgb9fT66NP4bMV3ILwtzrkHhP1DN1eAUWyNWTblJgpTYksDRpwniBF
FGXtEKpLo4nHgAn5MlZavTpv+nnqefjMWaouvWuTTHpl7cuBZigLiJ3BHA907VQ0CvA9lMac72Ip
a9qp5wrwNuNlSoMEnstlmznW1B+z2nlBE/lQ/PmbvnNjKYR+BGbbrOUQAlzVmw8PHfUfthJtaMBb
iKHaQNq5k0hHxF04I0UoPZVEx/pQ4lP3eim6d4LBacuazPC7J4LiqBIDd0a/gOhclKDeSGWOl7V0
idDzdYeDR7gNBVmrgSTqImK+RMpBE8iWHopM9wUYx85YcKqEmFMkwieAeZ17v9iXjjVL/1oDhUFw
PXqYg3pj47QPwgq3RqfAxqQSXe8XWs+Imi+5ewhi1kvEVHYDxUg/le+0qPBo4YFZHdRybj1YTt8V
yYwPyg6cvLe6B7gzzHbxPp9qphSLSGvcH8mfJVOFP70sLpkjA5hqLZsU4qjPCwu8Tue8h7ZOuWGI
c1d1SYqg8Rzqu1AGGF8Z5oiiIAd6xCHdYkVdbZPTMJDHLweVEAf/EZprXC+7Zddcj/tkOcUlvjiH
fWcZQwOUuVKY5iltwwaYBFUtDn+TDt0e7qHptI/oGtaTi24YM9G2tN7krNQgbfBzr7sfJ/tzXqHl
hZI63OYhsx0xlVMJMhH6EOjBbhJt4GVOv+/vpzyaGd2+L8WfL2ljsDFX2QDuT6YgYiCXpMyphTQH
jxST0ti2WXM54vWT3kkzloxNHXLf9DZNMlpnWvlUufYhk8zNBoWIDt67yBq1gznyQAR565AUE18/
am5CF5U6Z6CgYldVIZ8pTpsPBkZh2Cn6dOCYjrwUDNzINosHnUGHoZ3c6UrcIBP2jDQzaW+YenxE
9Icje6z2vij4d9OQIea+Nj8Zv0aVl2ie5s3Zq+0psg+JmwWr5Wgxmodz8OJhRpvLIjWo5EbBfrmU
SWqKagTN980FHHyHGrfvq1sVxaS/wgnuZ1qo80ZR8F9EDHZWez976BFwFRq5+2LyWZBwIZuxsO8c
TpXim8MGOSTJr8plHDp+g/lEhY+BaEt/p4sz7aYgOw+bvSO/HW+BycW7Zz5vwxnE5QnBZFT+z1iS
GbgXbMavK0y8bfuu6XRTTGmIzJwIN/TrwUCEsAVqvNi2wFZWnlgJl+OD/MZqv1oXrhpBiwP07dxb
7EvCy3/j94KIrBjZ0MVJaw05NmFz9Z6Nc6r7nGzTPqBaUzPLgfUgV4ookoOlc68wxUUeWxgu9ykX
kW/QMnVV1TZutYXyvQG+TNXwk0EwZZVh/YL4TRDjuF/SOHm+s+xb/VyD9m9KSvkTgxPicckOPYHC
/dWcpyzVozTlff2zstP1jfzQ2M4rJzOLGEUnFP/+Fm6QWp72o/y9N3w5BqnV6SmlEBMW4itdB0pF
63rhPjW7WSpgSkrvCpZHYED/NJ8d+dcUro/CuYD3OlY/ymY7rZafRrMrJnYGNMrboqylgFkO3H9r
TSQLWr/yhVaEQeocBYAmgqBraI81ovnuAFs8z4950kQtklXb/2M1EJNo/SXjfhfW3MqImmTfwyAh
I1LxYL5+HloQRJgAM0LRnsFzKdMLTvA7WqS5lKEzgWPew12bOhOTchQANwXxydaz2N2GX7JElGIy
jMy/BG2ICtXpqrU1n+JrIMR8g1KBZComtkG7YADmY7eE9lP5KSHhrcHBUb2dcAhZc+/kp1ppu8qk
N+VgDFs/a3nnlGcF9OGuam8AiI+IHXVS+7HFrhzrNmxJLuw8bkMgFDV+rYZr8VIXJqzlTb3ssROW
e2nIWTPmDCnMeEOORrbJ6RCKrb4T9p1yqiX9C1ot6EhXwWMH9OmptGul8KtMMMiPX+MzmIDDB+0c
sVjvWvwvmjoH3s/qyMpcND6UzOPxoFJt15+LY8lYAtU+CHIFxwglxpnQzOygEvCaimTKhTV5/QxB
WXfF4vdzGNsuAbkozqDhy+lIKqfffRi5M3Kkt3V+fb/9+J+XxGrH3DuyWLj4DfEo51vUymXYiu5s
3jHL0cgS6bI9xJ04BSUVaUcRuNDSAQ8Gy8sNbkFIgB/6mxTk8fijUcQWXi0ddaLk6GiufUvgN+0u
tVBp2gnF0h+sPfK6gbEme9oKp7RzQ/c73LOUGKr5ujybubiFW0BHUH4rU1eLn64Cd6w6HQlvS/JD
kHyFpUrozc4mSJsiA6FPhyWf+5Gqjq2R47OLPtyJZ3K1UygS1fGAGoKKvrX9vOdp8NNFmlhpql+u
V5Uk4/s+VuBXah9YUA+V2Unttm1pVLlz/3khI6RPB0EZeP/+aYaQvkKuVGxliKLe2IvofuVZqkuF
1TO7GPHVkwhsSlpF2C9yRwvdPmPWQ9kmdIcMkbj7CvzY78gmKkb44jGbdGSN0nkoDDrRDMUIz+VN
hRg1he0VoGFu+YE3W3USYrzfwrV+H0C/l7l1uuCQLZlyZdRI2Mkj6GZLEnFCCXhdKEKG9t/gM+Pi
khc1BddIsqxVMrMA48vYg+9c2p4QclqZQBB4vdZdol50UNU63jzxLia+1+lalGVPCI4dsWlrgyxG
XT+dvqhZWlbY/1dDWJ1dYs7u5/QbjpeUzoskOuBfT/Xec9fpH2sqFBl1XMDNHQi7DD8gJ20RRaNh
HxOU5rkhUqsb8XfeB9nRPMsKakCej2we8xk8omBT7TJFW5KSWDqNEBnZLk0Mhqduoj5lTgEhBivP
6GRQuDzufMepdPcP8ujHDPWKQ0oTCMcAkBedTsdRuDx0SDXB5HHT/ssYuCw3bBumh3goumBDmCzo
TJ1hmAL/L3EAQfJh1vlhbqruA7G3CId3cJKXtv8iiS7ikIqItTQfMvz39AuLM8DbsoMvozCLwfw2
KmSTcE/T9BM8TsFEUbhVWaJfbDLHVPcn03BCAD3pU2a7e3Hn+IJEx1wWvvtZsSPYOcMNYaVWIusd
9Zp7IDQ63vaK7U3ReiuHRi6ZfbAPjMRYb/LfdEkp8bdJlLhus0kvHd2c3p80Kjtp7PY4e/vligLx
Z+n/vCqFzFQEotYGySsrnCn06p9K/piKdX1SHf/AttZuqRC0Rf69rc4vwfiE2/Ama+A7SyfNDO2l
zwT2nc66T4Cgq/hTFt4Kp5JGPe3koyPI1eyVcGlH091i9wJixfEiL6NmO3FabZYuuVP7gQQETMkz
pP1dMCYL+xFl0Wio8+8OgaxufQAyPdwv5Ba0iIychehevRHLd3kBS++UBlnKYr+VAlo0psa1AdYe
SRc937Cay6MaU81Br4G3criBrrk4iIuufZVw5GsnXvpqe6ymNSOl111aMwGXnt96fNHjQEGXZgRZ
nDpsDS3hI4gxvW7nX0LSRHHcDq/zPh8a1l2cuByqVUIi1LnYb1B2owohMBy9RJnR8FYm5244k16b
L7stj0LMXTFVySNuDO1MMA8mqxlDH3mn9wpG362sU6+BirlbrKJpHIgLFTmQ+uLztBVFWVrj2lDC
p6S3qpAKZ3pPQcXKZAIYMLVoS8mFnPLkGzLHoUj/NLlLiv2dbYQqk3uU0DNOQLR4g1oIsLxYw5DE
UHWFgyUKfvXSGIQ9ZOJ0mBdsM+ZIQvtlfp8fI6Ne8VBard6VWkvAZlMApPUKf2+gEOH6DCDt9WJo
KX/IjMFhlD+2rQJ8kHZYYr1guZRlVi8wkWRVzmTh/w1gFP7Q3F0BBO3SC/CvdDPlWo/6br6tR6qJ
NYui71tTDRF0FgxDWYKheJ8J8Q+WitjCEg2so5t37Hi2rvmpQxxVV+XXV5HTBnDoaqHqgxJZdJE5
nDCP9gpaqZb4p+OfCaVIhU79sU9uHcOQYsK8SqewzTcI8rS9UhyS7uP045ymRf3rDSozIu1v7fEI
sk3prqFIAFAyx+DWcXNNN1PffQh6Kb3c1IVO2m71/qHGrdE3ixfT/mH19RcC7JKel0QJ34DFL1Zf
g7WIzz+JOQGWYLH2HVyYEc6nkSUNAL/m/G3n2bkNwWUZFB6NTFTun4A27lflhdfmookc8+2xh324
/H4z0+lAKkCPmcpKBcb8w0suOhPlyEhaca8xfVtjV5Sxj0MwLtIB4zkr77B9UlrLNxM7FDRopXOG
K2/0EpZm8uVvFtFghohrqpFjEL2GWKxx2RkVUkdNZuI7cAZuF0GfFjsduxOd02bAbqE1jUX1ynVr
bHqtsBg4Chc0v0iAP3GcIeIKRDMGzZxbop+e9na1obVp7MqfJNi2DThKsiqqGTuuNN+QTlKNaDVi
T5FiXf6myPaighm0KeoVnqB+lSnf1J4uyOlCtl85HwPaCBdN7Ws5kZy2oUC/LsEzAcvISKVt7+t2
mY2YdV6zXiiQ63agaNISgpxwUJkarmsIfBHch6Jnmt2hA5l3t0ZZuqw9ga07Bhx3XIGmt3KQT7lV
TGxCfYQ+KsZ50xWeLpFM+2ZoCdlBjhjyIwzLcetQlaz8GXqdDMUoouqIVT2oA277EoLz30zGiE5w
ddaMsfIzqzxzjc7aVAVzGl/lw+mDNQ+a3gtjFRXankfukbBFH0AndbstdYTbgZHidSXY/o3sKlQV
I6aBDehm/MdXcSsTgjDExhBIuGdITx/raQsWXKOTgskN2M2e2Ye5JeB77Epuu8Vnf1L5FODXledZ
hiMm/hzd8YueHFZhBnv24K2cq5lIeC3Mq208oDdTaYt4dauSFOkrFlmqX6/OL5xtazOKa08K5kU9
3T4FpWQuePJBuckv8KbyLhJHIpKVA36edy1FwMx+XwxxUPYFgb89j1HlD0EmeAW2ZFp1JmElZtNw
u4/TNJLaidQ9zRR/4ySY9JCMAZFtjx8Scwo3sOe0aZ0WTFiwm/1ZGP8xFo7tW6XZCr3Wb6rt4K7H
ZiLka+IcGbKMOtjFjQC/tAAHleKMv6D8k9HHXq9/t+A3XeQpLPEGWrPKZ/OdCi+SNIFniREgCce5
UBnKp2DJkctdyUazsRo6+c5kqdl9lEuEnMOGukq14X5LsyoVTElmrVb+iG+Zoytr8fGcY3gyZ2mA
WodJz0BVYdz6MdDz6380S/PCY73GAKQeduI+ElZi1sx3ImoHvhwBunSzPYrxQlfxkPImACPLTQ+i
oIRKyhqDA9QW4loi2Tqbybr7MvOvijK5QpyKdHueUHKGR6TkX2YnIrtMtDG0pME3NkQqm+e1aMC8
ukBkyPteI9pPzCxOnKg3EnMNFAoB2h0QM+nWu2A5A+RSFzNuJbu8Q6xeYH2eJ/o0KM/ZAH0MNQj4
eCwtFaaLi0kxU+7lgo47amM0JSlpC8cQHSLsTagZeBrctoGcGN5n3CZvAmt3eXSRNSzhomQ18OTo
ws/joEdCX3jUnKg+0BPf+yt0qQg2V3ltK4Va1p/c9KqnDj8qok4Ze9W1B8MteiHTpjmrHpso+8eG
It4wNPYNfFZlEWr+u7B3VkPL8YsGY4iqIjcVVWMgLuKxhIXDMmEWOcj/EQVdgt+HEr8/baobCXdj
Dm0S0raTGtbBUzBjNGyXJo1w/0Xf4eqg62HDgXUGIiKV68nyRZ2whzX4fWHevvO3fIq+f+k+DsOL
L2fMK+mFCimyhIz51ru/wY2bJWvpQOFnjL/YweWyKj6DxEAlCgiUduoxEKuuUZtXb7BCURFwWF5r
ta7m82+euPmvxhReRxcaguHZ2gDBBjRUVYUamEaAoc7BnANivwH04QqZULmvDIpnI03w8yrUNEd6
Y/s54ihT8h5m6iLZ+yswEwixQPOLDzHisXyjIBi1VEuENTZtQ4leCHKjRLZ47q5RV6Ok7RACqx+7
MPDOQOIK3tjWtkx/jN1jcOw9ZEa8/Uyyk8yfh/P4kHcztGSpanXvZQF4cs3Ztzxuos0Ii86lwQn4
04YzESnwGKP0p3afUp+smK+g+jo413uhoBofhPqUjKUtlaf1nzQWUla9NS1BRW28RypB0Vgbdzso
oQWHAxI4+rXZAQPoOHo7B7gZ4EE3bthUjuIPvvJDdh8iqgZh8ydGyE2ucrrH9+ByP14Lzx7VgvCU
7Le92DqGpFMJXQ/kFT2XJRnv8XPrAB/+lPXSf/z8NkBFMcfXcxT6IpimvauR+nZZbuQsdoTGxTM0
QkCIxKgvZ++H/mWlsBsVkRrRmMV5V1x8GtJkNWBtIe36n/cZLYR/6RoKGH1+2tVWDs4OrC2+dKyG
uWtnWNRkPRYrZwNq2og5BdMX01yA+YSZfaqF0RhCkxW4gPq4Z1fFaLWJOiHc/UyzkWR/96XTeLw3
icYxnx96oo8eNzaGfDYgVxrX8zcvPDzibGANtGOQomescpPCRMM4xmjmKi4Zolm8dt3z9vUMBI5i
5rxKjhESj92RUvcbCVfZSnM08R1QZhgq3M292wjIGJXmt9N+PZ12w7UwKThSjHekc+l3dttcyIEN
zqU3bFQ++aqNkmX/r11SdAHGVY0HJpfvMhxREBVsj2Qpx0Fa2omT3IA4HqOh8vg6NGlKJm3KDqn4
4urgAlx8rXFq62xhR3QajUooiUZj74D3/49WAfmnwI2fDQuGhY5umNOSVVR3Ky6xfCGR45hUWc/f
ndIW6242ve1yFUUj83tKNCxYN6ZMamXLPjOF0mQr8JO102rVTFaNK6OcqxACO78M9GRQJMc4KxRV
DBeSaJOXqNXRnFq7ueOJNTASWRRZn2ZleKutgZtgxi/CmATKCRNh510vh/DTCPV0KNZAygY/6vDk
VYGuFu3F/S1qMv3JmF8M7nfLCDtoPFsv5h7UXiHi8DxrnbHCS8T9qcAS9wDPT/8LA38cgXxrn+d8
vymqw/1inLAIpax3evosc9UzYcW6KubtqW2Qos4AnTdOuTk/k0FVM9+qGPm4dWWE2EjjKBxvDaNn
43n1TVQqW32zkfnzudOqKLsyV6xNH2TsYACi632sqppJHyhKSgPcioP6RdI2GhP1/fLIgWKrvXpZ
fi+SRq6lO+J5DI6P2YSvJ9ZvLhd0gzvc/+qh/x+FHo1eA8Scrnr4IHONhhjJGDS/5XoyHVUMNLlL
anBNFSKd4FXjFkqhAxkFyrOM7IwOpl0RszdOqR6EFPBGUbrMvo/iN4S4WQ7XqNn0B/DwjzTuyw4D
xYh5vaSnHX6OG1jZP17QvLkCe8D9rCqqQByZYMIc0HlzEpYeqT+W7PPynHb9hp8kFXe9JeGorlX8
FEe35J2Yw3pZKk16rivxODW0masNCAcFLjhgL1a2OZk7At8GSwneh9PRkAruxBhRKcxIM5yV0rdU
F/6Wwb2SsF7JVa+9QW1pjvqHVXHHPIW5F1zSoSKe6MSpwb4eYI9gragRC87yYhFESrlyBY6MVMms
O5J/vTsHD1Nyo61Dor9MMQUoz+4iElXosjHjdaw3fvWqU6ikPaJst7jSE0nSoR/d0dFCAdFA2oKe
HWl2+G/5VTuq033Mz4GfpDmuhYLmsXOM/VV72fJCXkUCkDuAHdvmfjzeog+MY4ii23HEkErnmaPp
FR9e/tfZmPHaqqwXoIdzn7O7UzE5E24rMliLzOBor+9oZEwG3aLVXzkMHfc5tmX62zbCHiiG8JS2
L5Gak9vJGmhLr8AD/mBrV/mwdhv61AnchJvN2k6QSazykfEvv/2G/1HUtJaMNEpu2Aw6cPjdbVTh
YSiU+jVDQwA8NDVbH+Q+qxJ4KxznOeNXYLAXlpecEam856/Px3+P+cCiqXUz2SdU08jBU2sQCG8l
1RnJ0mn2/+iBD2uaytd4N0gyr/sZg2pqUbWdBcIASDVPj78pqDEklYLOHQ+W3/JglzJdZmYsDWm5
0dmMPdhyDivOSECCupHrhv6Sittq8M+4udNfsVtHwtwT5jIkyE5yoBkO9gjTQy4Cwni2zlkP2o8o
rtuI0uuFjnJRo/a7XG1xDTKtqDUh6rPydN0i40xTOBKfERSObTUNHGGMd1bhsYWKNiXuMowObG2G
DpV/lBxu4kIZagtEBZWxYylRKFfm45ad/APF9ApBYxhNMGoFDPPL1zZdonCknDNc8lrABiDCTn9p
fcN0HCdRrHLwmDCYgCyzwAH/VMu1iW+Nf4lNVPBnD1ygYVqEV9/LW56rx/KUqyxsD+tigEfmbdr3
STguepMPdNb5VrifxOkWKMZhEkuoqVEJM05NGKYL9vIgO+c5m9v91obvTq0sO/c3NRk0x7+ORcSh
Bnomt/Dp+mlqBlLizTPe1pmSFrxtek9gVbnZy7dLb5AHPU13S0pQ8mpzZl48SiTFM33q8mzyXKod
Tx1S9H2yPpwmvHmzG6Rt/16xpo304P86DGuzMCCvKF1ZMv8BBfuqivxSs+n0GqmkVwAw3V2sBDeN
ghHsC+CG9cEBvDf49b5XbcjaKXll34RB6gFmkPTLDRMVNfUmjg3mNDk9djefSC3QkNWR5FjgSzHD
yaBvyOJZM9yW1S+lXbFGnpEvUp0kbwzJECogWOfhAqkR2VfTHJibH1XFVTMZnviCrypI1R1auYlM
C5uFLFhaxrMCfp30APIvCyG4VLCjEB31FtaeQMdHAde1z0IYVcFRZv38FhK59WWAu3NZruF0hpWg
VhCbL959YqPhPbkA36bDzrAgwFAZDhP2yMYiFWkVogaRL44V+z/z2/sJRBs9+jbU4Cplh+KX0Sal
ghPXrRcydE9wMPxvVaRk5vj0iPbV0OjzDebd2jUr9WFnGwRrT52bgB3HjznpKAoYkndHdOKR6fc2
FLB8FClNQSFogznlAoiJ0ew2akUFRwWHns1A//PTZvtEtqQsy21zuwbD5w+t8CV+ocjvRG5cK3Tj
bng4nN06SHi85SAKOeV/zdiiVvjCuWT/1WJXcgenoRB7GG83muzYjGHCwbUM8ZPRiFMn2m7kDWmN
pGWcQ2r7ssPptsN5o9e0d9l8LgIunlhvEn2e4uSoBtoIdcn/CmWusC/WysjW25Pw0Qme+SlLdE2a
yO+oOUqnUnFDr+LeEAPM7JWNpPayzoG+Nvf5XHd2TJD/PtnnPwEMaXAXoIZVk08r0OPVH/SJqOuZ
IsP74aX0/Uq9NhYDkEh16J/FtZJQ0x7+MY9N7btoRcr7VyAjgJKaIYPxI3xwjCF2aHoBApD8pd1C
myegNRFHAMLGAwpZpGBc+9iIqbjy9eaG5MnPhn8vNQ/tQF8ZYxEq1IjYHTZiqeRXBjxWIjp8Htbv
ani/Lz1WQAS0fJRi6Ln/FZAGKoWul5cdnaJACGQe3PbTQvDI3qO3ukzhqfEZ0+o+sPP9VL3O4o51
wCe8xKns8u5hnYDChZfFFU3xHZyl9vEus5Vp/IAQQeGPkUkNhqcrYtY5dO1/F21TqdxxVEms1V4x
vFgy5Ug3aD0kZJPEfGS2qVib3obxdHtq5PHiKyuEMRGAWcqRIELeRDuQFW3cBb+yo8KI69b34bPP
G+wevRxiIYvFlVJoT3MzA2d08BnxXeqokMyhXlCO283zKKS7QNIZBr3UoaqgzqYCdZjQUFuZz360
ha53yjYjhaV866tLl4DhoawW9ok1aCLhO6ZQ5tcMIEq1pAyItycahHRUgWm4RFtIpfWg58xdBd+7
rBoJERjgF064q77ZNBkmNT7wZxx03s2BLGg82TX74GW5zoCO6T+3HAtN48pelIyxXKms/uE7mVsc
STIA4WEcFeIABjqD7R5cMMjL0t+Bpn3XknJQtNg7aY7uyN2zdjkXVOs8HMnaf/R11LaPsSseut2m
hzn4mCkdT/0dIKvq0UvGsGA78nMnHDIyJ72mnu3g76QV14+NHcmrsuoLhLfUkpVwXhJ6fAKcltok
KHfz/bKp53wzLfxwQ9RRKTkLeKI+8rFF088TSoohOmAcduJOJM/XiJzOHYoIVmmbV4ucFgToiM2U
dL+Wz1eP28JPURJ1YKUzXpCiP9K3QZdsd6v0KL0SWCXmhWjMnL+NREhh6Lb5cowvF9viOLZd0vwG
6W0iR9oVAs5x1YedTadptGOiD88EbWqbsoJW4eAL8up+JwnaRrX8jKVDKwgDkKUjdrds1SreaIa7
EoK+qDOcMczkeMZA1Fvq9Uv05gjpDBuK91K8gjtzIpji6OZMss29E34bx73gBJiJffHL6iIZ61JD
ZOrzVKttb9+sLKmOMLq1qGDhm90Vp/H+9bsTRG0dN2E13rpYfZ8+ey4Zs87d/xPS8mxbKBBWvwAX
YtXGaRotZGgd0/ZB4EE0anuks6tR6AFJW8ZtFCU1IIvely0IIlQsQp8MdGvSnMbq9FlhNfgJ3uAx
jEJpaopjVyKtoedFd3/l0en9tM4E3dfvhWLUUTF37Jn5Bf7S3/d7jB6Ryrlfs9V4eFjdBJ9/lUgP
N4HA6kJDZZRyHnoHT6KQYzCZq25j+bChDrftk8o32m68+Jp1AjvbkFrFX/Bomhvbnq5gBbHCJWzX
EANgfezTbDRPyJz6L/UNhE2vD95NqlGDQGPwnP8j2WmWD7beo2cX5+6Yo0umF+voMho4RptNt38y
B4/f4p2mFplVTSji56jr6zI6TLQMByAxHp9RLWvTUpwHwsd0hR+iE5rmK68iWywGAZAvpq8Lt3EP
LDUoTnzjvKW70fuCLlioFv2X1vQsq8p+PXADEdyD1dX8LAOlTkP20/Oec3VMe2Edtq/Y49pm6igr
9nZaJjFIG6J9jMus/7tFYagCRt+uUi3Hy+txLKkjqY5M+4hSXz9g9uIj6HLBTGpHhwGg9IUIhLmZ
a+NFTvwqddWxQztgvHoWJh3G+Wvm/SfbuHum2c98opM0C/37jta6pEbtNUdXjARYCOw/mG1296T9
dbyC3gvBvZot26QX0DU5HaTzEhNSJPPo1ZBIetK0zEvqsXjf5nizUGj/a52QZnditTIEDU77xTL+
gcZY30d8lOVER+0edNNL6nZ80oybhDMN9bslCQwv4TRvbLp+bcuJAXZA2vD0pU0PgTZNOjIBNu0j
4AxdOXfcW7/w192oHSepD5x6oG41DMVIzBXyOWc6EGksGZVMQYynmRAfAEDxiTVW8a6rPTn6052l
xBGkQPTNuElaDIksIaUAOKXeLwgscBJ3QcK/xfBu8wshY1o41wClcJv4wtXjv3cIO+vpW9hCB+0w
89ecn1tMJQtHEF1hDRzqWtcGJI5v8LXKQXQC+vF5I3LKfqDVyxesch/2ZdE/BN20Z+bK2ILj2SH9
gepD2bf12t4ea037o/Ywjw/bHBx/jPy22+UOQ6MTAhQk3J0s12kTneWE07fi1b4dAUY/Qgv81Zbz
2Icl9iGEc4IHD3aqQTTxlUgkvm3yf2ISYqSdWoDlfdwUdURcS5TSZTQiArJC8kW7btpsfCF/0exe
qnHsfStIppXM2nKY+4hO6Mqr3z4UCy34q8eEQz7+lUqRRu8IzNKDDvQ4F3Qp3fdYC/+HMOC6Sjxw
a+bE/d06f/6jIqPf2camUX3AJHjBwTuUCtxrsexVo8z2mOJmSjHjo3VJ8qymJH4up6Kf6aictVNV
gh0uSAQ3sy6s/JwSK5zN55YDj5L0IASUQaPqL2ro5fhzZmFefx8cbql4sBS6fGlPMNuCoU+qc6f1
PVASk+LdcC53YcNG1ugvA0IJKMpvURVLFkpF0q2MJIUC5jtnt0zLcn2YxIyWroas2RrOgA62qy7t
W35pS1i/UrxiW+4I1NRmThk8Dvoyj7Xghdb7+2DV97FBKMLyXe7yQXdYpzNuHnsZNHB09ieYXPd1
DA9oukf0WNJq1W/8Di2Q3dgTeiGl1KKyvt5Gl023ODf24A3uh1L3WdGMIjWnUtYhIHtGwo/EGxkj
42BL2oJSG4FTZl63eF8D8o08BcOXLb/ED1/BjABH2tAOKD1kXEQY9Vm9jupMrfi02vHTGlsnNQkP
l+doMFLcJV7HfjeG45TUxmXH7o2SWdDWECg+ZinZT+TD3jOzR1aMF4AOLM7H0RIScPBMCaRYDPUg
hP3L9qQfi8OVGQhhSoqyjiMefcYF2Kq97qZQhWdoR6OlieMAwBKpBLBw9dpmhc9Al9YbknAnoA1v
k+4zayW+zWPigEwGM0JKlfBQbcpyEi6qifS5iH5jQU8zDyY7VXjyk+2tZ4dGa/DytozBSw62uQPf
B/utvfS4ea+XT0QHI+5rBocjdjlg/SBF2cHYOEECDi12NF978RkskdsUotIks9yPmImC0j0vjHhv
Mrpn2TB2oF/rIlxgQQL//JhbPN4jws0eFctffeD5OIYTHVzRFJliKkT/4RmliOCJYMhzIutNAcYZ
oSpCODdFn9mP3+NJIFxtWVuy5PfENfDhaRmk+ARCweuAKGBhN275puFcvCl+4E4/S0k7TXiKNjoX
xHFNcHwbhKauUaKzk34L6hpw6TYrpxia0iabH6eJREVUUfbGAW0lDIzagJHzhls6nFdN46zDML17
CHYyNO6r9HdYFp+Ibk/aN6cUBsDrUIk11BNoBX+PH+Esju+cC/9Naf22zWj5k3Z4S+0s85HsSkQV
vqPuXqdC9DKUNEAhlwAXDy7Y7k3p9Cu9hwUw43sC2+GX0ysqaSZTUaXYt4IVwrKpCKjxeCDq0kx5
WPaAFBdVUk+Kq1EOfgTp8nRb7pf/HstdflOKzY8htnpo1jxmkfhrd2w9UYSLE7N9XfVroG3nDLda
OX3yxkLUKl+9qNFJ6mwrKoFs+prA6Dq78VRcX6538UGEAVbspLh71C13Ui9FMt2tF/TzNEi/J8Bq
pXW2g4H5FPBpH/rw51daP19l/sU5Tv9ACfyPkOOB9mdQa9ZSVcyLr/nqVRSti3sbVFUm0RUcN9y4
VsO94cmO8Vzbpj130R3RY+ulWgX+rTGWNyN8wB0sF+OGNBWbaKVOtlZKl4MYP7e12ueeUd3AVe/r
5MQUdb86VWP2seX5isr8FeY+yCzvqFS45ZC0+PdKH2jf1QCha0lO/6qCLcbusiEzM2ZdV3NTsgE5
OL+RJZA+J4MWo8YWMvK7Hq3EuDg+fOtnZ793+zFU3r2WPtGAUWBH9BGyPjMIqJ5nSodCuobGc/Rr
SbqX8m0b0VaucNelJZgBx+n6O3tD22l3nYAeqjfX0pQy0jUyqFtfwyMYSRKqA9838P36NetErfB6
8ex0aof+0jRKwhVPI82TkajwB6TiJq9ukYBC4hz6SDsHWFDD7n9Bo6SzrTmVAn25MRKjtvYOOf6o
Fnjrj6hkukktx9KuBQR51Yg4dRcjGWH4aNJquTjmE5G0vV/ZVuhcMROGtXiJT6v5d/Rej7EPh+3G
9CfVlCgKRKSuaUkgqxAQh3f24T79hyfrSl6Rm2cRN0EdPU/U002VnDsbQZPP+ABSYpQNsih5Ie3+
eALJVGNyLoVkFRdGnxbFTamiluWduRZyZfBFz0G3rLcJrt6qG943lybjoR5y2owLX4/p71ZL1fyG
1VJhnIMNkl2P8rWZ2BEUTCPlhATeBAqXnnN6PL/g+JjgG4nagDQCd1fkGCMsRG+CjHK3+6D8GBNm
VL2C+njuHZcp8Ju3xZy8ZIRmx+oT7969D+KwrvfbOgvOwkALrO/1dgcdwy7WJJFnyxJLIxDsCBXf
XtuQaFhetkLRehCwsHxcHtakouet/voPg3++IrB61rJFasO9Uwc/1yem78QMEKed7v2xTUTIT18e
oqux6H7THQc84yctAKUwgXEaxCZjSc/0pO4DgKpd2w4HLllNzs/MShlnUPzBu4iBz1HZu9SMPh3R
SNBfnX4R2mQeF/GCGPR2GErfmv07FsAeVRsH7eekLcir6OqpIlLid8a1XG4/V+aebpuMPXSrDwO+
LapOuF8809gzbOx5jkRq07dy2FzRcOBqerTPMQBFAd26gj/yNwm5K0gtKZDoB2WZO6k083LWjgsa
+WGMe4pvk4n7JuzukFLrF7ghM7D84LQc9k8MPnw2aRuRf/3+x99PlfVqRY4xLTzK7PnKhVAfW9Id
Jjvnzjq8MyUR/w53Elpygercl6+lqycMYFVyDR4As7j9eTKX5ry4bHviBupZuj7DXzo5aO6UUJm6
a30rS1gcsXpGekQqAP4MuYzK3EY1T1gk2BFSPeotEphvhZxlCHhKyusXT0MCC8fPZWmdAUtuGi2p
PsLXW+Sija/lnLjOpbSgRYYm0lQmNTPZ1hJKESfeGsGy/VG7nN3CPxTp0dssf0eMSS4MGWwmjX2k
HZsvCxyI2oQRdzmoEpmcRovjgZqgcJ2zwi1ZZhcKiTbiV6s+XLTcCTAPb5p2O+tfHKjtGwEFjpv6
u1AG6f0lnycPGvfFzriV/uFGDHJ4RcmuhuYFePBf6fuh44g/PMtDxnGjOcWBYuq++KEgbq7UhNxV
9l1+iRPPacoF6unLr7CtjJZaxF3F7rj5SPOkg0YVfCEAtt/kr6cR32959xYBte8pIbstFKKpVfxV
qveBfm/5m06pcZbUftzfsoktVF21RAYv0HEn7riwGskAGz88d1qbXkqvudNxzDEgCPGnGPrLu8ih
rWwSY+A++5nxgJKYhDWjFTyemO+WL13geQGch9Zc3hqbSqGl84+2oc/UQ/SQg0GZR4QDq9X8xb+G
T8ligvKGGr5KfnvXi5gbastb6RKSPcVbbrlD4ThXj7Gb3MDlOlJlz0b+3+pMXKSQjIf+XRwAtJWE
G+3/zbNovlMOivmblLwkFfgMIVkqdNelMPH4N1k9/eJ6kvRy7oS3JwgQEtO+umRftTa5cHjQCz4s
8jmAQfu5QEWoLsB6X5ZjdwS+GRaOiU81dyzcl/Qpa4faX8bD9gjUP1NRzy1zfQkqA/bW0+3LrX+U
I0CQEFs5AxO7j3NpsyWNhzViwFONYfwf/HjP9oP6mPbVo/uVK33ZO0LJgqT/BYLoB9JAFnDFm5iH
8PVt1xaJM6lMxRSkENfr/jKH2vOQ+FWqQCAulvWf8ddyxqMqjGPFAYBXVOZVLPLBkiRGMgmMHeqr
1thL976yL3IUsStB2ve969AtDfJixoZVMJCHQDrUIobH57yJfnNhnLUOa7y6sPDMcyDCaLrc9enH
Dz+0IGgN9AKRoDevpmiHMsfwlSl52uHmM3CN8nw4RYEJUmLwBmn4r451PZADanfMyQKjGZSnM3DK
BjXkXQ7+UcgUbppVMmkrip5HOGj8drh89uYYVgHQYOEWnvVh1dva6cm52uWyt0vhvLHrxa7r3epN
Vv0IcxDOLTAe7AiCoOKyDSJqumJaETqpAZPE1gKaGG6F/GtjGsukyEGRr8i+zkXAFTeZEROmWt5A
BLfFLUJVhTA0PMG4Vh0g3TvEJ047uoTMTDaYNjUgleYIzi6vPiV96jsJk8ZIOK2t5o0MPoKtGUa/
CQ/HC3JIeuVinKarqslBk8848AZwrlWIF9GuD8l/N5DOLvAVts6ixQ/l6FgNkp0M5GfhZAW4ZTnr
psorZmV7YUIOEviypx1uH/Rm+9rXwx7aVg1ABQEmU211yR6cxRO6G+/vX2fRoe+gP0UdpMC5gD6e
XwaTm3UPkszuWYgKjmjNBBd8vJpTgPY475991wrvH33MEvv+0SblDUEluL2NeS9yp31FaSs9kV77
OZ2tkdAEEb3j9aO8zxl3vy8GcAv0Kah6EKrw8lxQ21M3fNK7muKMhOJ2WQTuwZcfKVNOz0K6Sh0K
oOyQ1IV57f9N7NFC7VZOqkh8vxbmTECh4yeKXuhgZT1NPYqqgNmh3NDkvBZSax/fpPXFY3ihyIAa
yDO5nMmJC5CWIpiO9Wc/unva72kudlaBtEec+qA5/A1ye4sZC/FFoVpoDTOKSWLbl4ri+XQNkIMp
zs40vjto3pdO0AYJ0VxnXMHDp/qhol7qDkHgDAi3BuGwXZ/7mxAm9z6qkkmBkxdR9j9yXYQ7Uinc
w28iuVnRv0t0pE6dBCVW1vBXAcj1f4StXMQ0inTg7MCNihIQMkT6PYzQZ75dT5sL2nuz/XTC/fPR
48lWfZsZBiE0BpBcCkkOXrLDCbaD76N0+0zKFIdexKCqqkb8fvbmwte7aOvDQ6+irswhQf8WW44I
dYFRJAZVeiwpX7Pi+eEf1gkV3wJMKs+qeoo/1cLD3jROaXhnESyU1eSP4gKvVmytSfcMiR8MSGu4
5tDoIKjnXY8TwADy+Ruo0ZVTn8pq6oZ0wNyCK3gyymzQNjqhBxAdDYItOxB4FRtXZi3hOfq8A/Er
33CnZ2Wd8M4eNxU/VAKto206LUVe38KO16CqgBYZB/v/oQa3rIuLuSXVfjwPEaH6wkUBfGqZXfht
9oeARTefy8sDx+64ZriDmoVeB75f5T/5Pjeqz/rhx2qncJJ5J+sgLYoakBhSUVQ8pt/BrRabaU3o
NdRwKWFo5p7/9mk60DPcHkjoVnB2EfNnsxeQXb09Lpk8lXMencpHVE7TcQaQuf/Rrczm34o9UIuL
smLBeeWsMRSWy5zE924qWCONaJyRvJO0b0uwz1l61PbDKzQWUvU6FvSXIXUZuRr27fIICITF+QjQ
9BwNfw3HZpNxM0waeqMUqbUEqJyANjfFntvknNePPOEXa8aPZaB8V3/+UP2kIXacUUXyouJsZZim
X5J4LJxh/oKkFJD/TchmA2KTKA99+p04HBnni5J0zNLXU2P3TKd7a1WmtMVA+dOKxX6UOA+Cqvvj
B5oBBoZSm2xzSMdzloGgwA4JANYUMYBAet8Yb0j0DSZsLqlvmj+uytB+y28R7JBSl+ilgk4yFbKD
YY1FWnIQHB0HTrnLwGqQMvBjEFdBp6dYG7+b2qZVPPbcPKc02xU67UjYza8kCsNVUEwkrNYdOc+1
TDoxP1er1EKXv/nXtxweFVrBX4V09GvAyYYDEdFeIyvGoi4V3GxVOAk7qyl9qZaXRZNSU+09anvs
h9lQgDOPqURCIyl8lNcgXHJaxYDMYa1B1oaSro/smnnUDsE9e0MqE9P/UMyr7JG28TLaEunBDLPn
uNR0X7cKnmQyP/P/oRHLmMSqu/eq6EmJvazn+q6aYQ72x14qgO0tLxxcXHRN9OpubGP4/Eko0jc9
qEsK7KvGlGqOwpp1WsvF52SmxcVT6cyJ/dWe0jdD3LC2uphyskvxwTakfxGDmgaqP10c0xd42MV8
3zMnQCXrq4kchzGKt2ifiV8SUQapDQ8LyfE/C2le8qrODjyZhwHmRAIzpSE/rYN7EsgbjwLEmOeT
7MjtqZuxlpm4qAAwSHyPAVdn70DjgEhIafrGQnbALScA2qD4Qi45wZi3goInQZowmRrd3iR0xT0O
jRskUKThChOe38OIxmEcVDMchFAB56L7p0PNMj3C1tNfgA4NPz23DkOJo5YjXGrbOm0TV3pTTYRq
HAAlnGZEHWkpUH12GiLwuUY1JyLFZsm7zgHtfoXRZivjwcHTYQcBkUmLQaX3aFKSKeQdkO0VdA8W
jtxrlbDIijyrWGyXfDFFnmBKyM8thXTgnXP5DXaLTOXUZH0f8ipi/aa1pPpXSTKF/dmH5IX2c46U
ojltsjNBGLDieb+Dn8OCT8Jnj2VFUSFdsNwILOy+40mC8DhHRsE2jPDPrMC2zAARaKxBI6qla1wU
rPbqBxJfDm43qBM3HjazrcjIJIz+9CNf+s1B0Rw5SmhoT1iB6fOaELUOgLA9ouxboeA5LHdkZo+g
OIBlrTqzzlJsr0GlpuRVWDDDza0IhuS7eIYvWTSG51pocx8JOhlHvx1VnlFQPBMHRXzRYGj4wxLF
Lyj9VBdfiScedJs2bJ9H2oFuGglcwTFUdPJp1EX7D0tmP/CMPU/kgtcEBNIrxpFQc8db3+sW7kty
bvX3uEdGGLWeKYoQqzUerbF3Bz9Pk+cQTk5E4sSNSLz8/UVwRfUUUOalabEyHL+jtL+oSGyPCVF9
PbeFX9xw/vFK2IZER9MvAB8QqE4KrsXHvjUGDQu4ExQ6go274gwUKgI/V537Lh2Be+lSYF5c1g6K
J20TXojzmH611vFeJdRRGf9+eABt3XFU4io2L8Ie/ga0ulxrAgz4N87n6OgXwSfs/dhV1V66xfn9
8vu9aXyoDVdOkrJRy6zztKZuHrCm1b3HOqGz75yk8R/LHApED53nuf8E+TJWvdF8xT2MRVQga2x9
sqhCtyPgdhrCfuRI+GN59f+YSLjrn4GFBSiB6+YxHrnd3E7TVkBkii4bPdiFh83vDh8wWRd6ch4C
zHBngVySkNua0SfmLsllnHWbNFsDRmHCbsdp1LH3KXTO8S3Ptobiti7iE3xpPjdreT2xcmmir1RP
BOIhgpMikPimS64J+Lhyml8HNFNhfFTI9EwL9B9Tw71uf+RwXX26icYilH6oPgSXFw+YdFnH1ytq
MdPIUuX85vKES2jdl9jeML3W5E+MwszQshhAEfkITPEuon8jv7DjQZZIMckZ3zXF9sTeBbGWPcGo
z276hkgzqElFkM1bg20+eD9i1UFGau9Evaic2r0m7j1xN//LMXxfA8gLqm88OsSOFQAJ9T8T+64P
SMj7Danjv27VMKSnvsGscGLH94f9CUP9Ti6uavei8mwngZHMRjWXD3n11JY+Vfz9IKvabMEUSRh3
XFt/PzJ2C68ifENWnaJptViNr4yVIKytIbfrKP2vtu7F12jz1iads6UOg0SDlhg/UJgcNHuvzg3Z
oiz82+KYOVARIWvLop4NR01+XzfMN1FHrxFzX+IFZGdnaDZcPUqFLbl/KUChXb9zHosn2p/ZQAbQ
WKfPoILORjFLvLe0+HJfgIGE5kfC6lhaO4hA1MEx2RgDa6ONcOqUXiV3CnErMtlN/dnbXiZRcEtT
v4L5KfwRJ2Bt4g8O7zeJl7Hqm1qnmuylbMCfThkLfpLBnZ8NeSqnh06tYALfUmcko4IFDg9DNcou
HeXqS8RL/wx/PRFQCnF7F5ng7y4+m5bGh8+Wj/dvdbaRAa8sWw5kN6mZViomaEyb5LCmlZpPt6WZ
s2iautsUc1MkLOuepallRgv1HYsCEaRwOF1brBVTfSoCMuaTOplRNOjmTEEhfPaljxUVMqx2BLsL
kgKgIpIjYkDYadXiyc/eLqXiq9mDwTdSzP3P/HkEBTUUy73giuOjsxsr31029lFgJmUoLGk6wAxG
Hj8RPalIAc7l8xoCYsTYjZF12T4PxEZdzV414Ltwry+dUC5ow0wmRWhuqEl5whbEKg++L+9guK8g
v3yKPjYPJOAh/vHAWoVBnKhdNCPiMeFWiLNc3D6EosIbrcIquhkOg4mpV1Pdn9EzeUiMA+zTxp+l
WhDtf5jdTK8j5EN0i87z+h1t+kRD82CHge571oHGEqVmhvI59SKSvpyQqb/U/WMZNwwRxaxQBYGV
sAfYYnFgb9WFA18nwC6w8S5vv9eLAutBqDx2Rhckwgu4H7ZBKxYKgHzJj1Mp4CvELzx4M5Q4SIEI
vD1cW/Dp8YQtq2f3xEK3i7cI+5OVok+IZodbcgm+npcg1amVyxsNa6lu7dsB9FOpLOijvoBZUr8p
/ZBz0ncRJlX1OxgVpRMwHt5T9xhKC0ovqfDBW+P6gyKYRPk4w6zbC/i2Lo0fZceGKSPJ+sXGp0rF
U1lpvj7YUrqm0SwkxbhGA1NKjb5MdxoK1IEIcg2PKnEJ/Cso0cmps9KTxGpd7ZWY6eGapmR39/Ja
qKzYx6ksyCaFkSewVjIu+fJw9JylU7cqTVz+s/vHaDiup/KbxDgCcVMJfFgDTjBjCI0MUt0Vlf06
YLBNJVh2t7aKm+jwOmaangrRoaEmGRmWYTEJP+IRLV0tktshFFPHskAGJOxT+jlTdVeB5HB6kdiE
mBVU5+N3A+AtiubUeDbISxYQeWxQJbNifeDJmzn26DPktIRJbxQDQnX5sal/SIDU+suFsOHoxHvw
UFEIZuKcXEf9KqTrsqavlygZVzilarZ2KNSmCfAsXQMfTJJomygLeuGPiS44WgUvkastjZWMJLGl
KsDVJItgN3cCfYH+ao7Htgc2kI46X4DeeiTF6I5dfux4UqlacE+KB72a035peD3DfqHStjviJMOc
NB1Ic9blZ+SBWvsB1QtMkjRnWY/ur/5EvMbOV/zFL6cYnN9qrWecraeaP0auGCR44ngmCfGHjRXO
rNQJqh9wG45aFzk22iQE795nr1vZoX/N9F8thttD1oXh4zw95XSi1d+VIG8h3x5S/kcAuYjBtw6F
Z8Pd8Vi7sTxHohsQNXR8/V3qL2TKoNDHWT3PCiPhP8J6WjIh2BnqfHCBFVjK4IvnHDNSA5ATdadu
i0a860HLkfhh7bicxDRxAqkTyaJJv9al0qXJxbZ1hOda/WLPltAGS2Ro9lY0PQUYifYmRlCrJ8KC
VPWsHJxlxOYS2GDiCAh1MNdKCFvX0sNLyfMVzSgpYysxXb3q9oty4TClIc0QTOGWMSWcSr1SMAHT
GmlZbHoYDHEymhXy2zQocfXteMJKTiWWZ0wxDIB5jRcoVBpv66qm0fqhGEAGbD8ukxFXvzMYA4kc
QoomzD0SEDufo+GPjhpdHQ2cbWh1coYyRsnrj8oWpljsCgF3QDZHWOsi+eCoFYNMMwMvHXzrbxwq
mIydyFZ0M92/napFwS3ICoWwGkpb19PxWNgj5j45uqrgg1avyoo9mok/mL1QP7s5/eXFGL6HWizu
tkxMVat/uqNP0ywziGOV4VlLtxT3SBREIVVobqRc44bBNFEHPvnNCIAczDuiTE3hhO1i2u8Jddjv
5hKMbZym+AXdSf+ahUL8RZMBlcxMZBn7Or2//xvbmZWdz1F5yvMLf1fMBy/YaGioKMLPbPf53Mi7
orTIcVcyXqTUfpLgdm192iKC02QKGWvm7UTUV/Z9fx0zduZsqQZwFVw3FgH59YuGxBkCKmo116nf
ks4sf/QZmHr5YliXagskZjnpuhHT8J7QcnWr7tzk8GqiXscdJlshQ8sUTJtbBPf3L2+K9LthoZ/Q
5EAc1beYaFzLg77huzhTbjuYyfslxT3SbTVzvrd1wXTcJ7sDa1X5L7vvESNigP5fo78jICwvZBkq
Yo6tpkDYMffeNZRdIFt5ByTG+UQr1VL87Cc3wpt3sztidiwiNdZAzbFsEGjVdMoYuN4p+BAMus+o
PInfmxqK+zlV4SWjGXqmB0ZeEvNRy+MrmPfSfu4U8ZkLJt0sVxIblbWBwesWiuQcTZCCUOBah3mB
n6N72/ZNv+d0Y9KCIMV7qMRJqyzHbJlL/vvFiDaX58681y7LUwpjxowx9Zzq9z99jGqIFTekzFf5
aAnd8iO2nidYjvGDfG12YWQvGeo2Y4yzq89L7IEn4Wk9g1lk6qVjpqAnegQMrZkiXYwBvKqg+k66
OVT/T2/YUyggRwhstXzPRoMTATnspctEmMGE2upu/F5j5VW9PWdvWcugVKvqqDpZZh7ySzn1Rqar
xYz0w2H66C6ZELBab04G5+5tdWYyjlWulQp4tWvI+KbHbXAWx4yy4j9VGu8QEa4hSuJNq6E2UUqI
DR24pzawAtPcD6TiBcSpBMzlV/p8VxT+DAV5AKl7q0D8Nq0DZ24VLaSba8eyOwovFhA5DAMVxlsX
faLGaCoIVhJVuPOKy+H8dujesdxn92hsye9H2bP5tObK11VdUCBUj+ilTN0JwVcyQlJ0rDn+c+7k
1KsKM0Ha0peGh6v/CF5WZsfvN7NZjUI3Ldrq0Nx/wfYkg1OQpKtXN/X1KeiQX9EGpEA/kAZ1+LaQ
omdsIcGrI69x+ny1whlM7z0AxaT7MmpNsIzhaQtxRG9TVVgt1/XT2xiVTjMYxWLgQuLfrNyIZSwn
7nybZxQFvO2oT/Saa7kF7yFnqI1NwWatvYLgpGXzeRTMJnUDZg9YUu5FrDYGQJs8ouFrP/2XnUNA
trsspdQXHva+B7HvuD4zgC+6gE7djE89AByUIRT8qc1/kHD7j6Tneef+qHr8MscZcBXIHE2noq9B
nETRcQpW55I5J4nnivLwspZycnG2zHK5Gj3juYHBulANsiiG8k3U5dPb7y6K84MDOmDIThH358jG
HKNWVrQApVHI1mfalGnuhZsFSJI3xt2zZwxlvxadsaXfa20yPId50KW/yWF8ow4taHaViHYbgi1d
N/tx308NfNeI3rUw15JOSeJ7hfeC442+/fKKcNNd+938Jubu6la9Apslp8ICAVzH1HRNSs4viVUg
JidzKtsxGwv+Ned50Ed4N0XAjrLLx/jPZ5+IloFo73p1kgMvb/Ij9xxJdMG1CX2cM60B1I2YrFc+
qyt8ODLH49Xw8Av9NcLmcx3qL2M8M8hTctzO8R+2q5KbZmIc6zbr0KkcFrkfmkMz9o6NZeDS4NQL
Fobw43YtqlfygiPvEbHXM31yfzWC8xhTBl/3/3+sMwn3xFAviTTRDZbngVSzmZDGG0PtJyxFpM+u
y1Mn+ddkrmb/Dl493A6hiNql00Fq22zCSDy3VyMlVGi1603hldIjMgOWuVEz7zg7oHUULbSuMODS
5O7PLLRMZeW9v0O1CJktWsS1lHvv1pZ+fvD3rJsfVjAKVwJGs9K1i0gs3iuD7FQdrcrSW6p5pZxL
/r42aWdL5zLIQb8N9quv6kHeGVMaQioUBPAoAUrbrW4pxAOtr/WRMsKCH0WKNrTQt8UxYpPyoMgo
ZGL/97tYQCrnmrq0aVcXV4cBEXF+aFBbQSRzFQEyg8S1CUHhU9mubOV97N+RlYSAnuyQefJK7d3O
IUhAR8WitvCsNOF2L0QIWawbQAZ1Sm5IHt47tyDmiIKai61t5Xnv0kVnheNulcfXRMGJoOOUmLSi
ZGOXi3Hu359n+Ggubo2Sxwl8CxeqYWafcSGeMXU6xdcKuGpUB+HDaxGMEnXwgv4uiNiuAT0VTZBx
aFXrm32JCj9dMTy7zBq1Kp1wnSj4Dc8AOCOaCq+D8EvcWVXX0bO52mqXBsl8oOhODRsA57Iz+F+B
sipJY0G2Cl/Q+SezXNESdcDsCuxSxzdpbiyXWjcneXhTY15AWgmCZR/ngdiczAYOeC+1xwQzocLU
Gt1VxRYrFP05ATCblwUvLejwrJCmkd8SHYnf1a4LDP+69iodXyQnPK9DR/aW5VzydOpRZX35Zjy7
G2Jg0EVVb5yQ3XBkvCP4OTN2IQbPpcldrCPFHfhw3IAkbAFtd9Cxhp4xhXZtRQ4TpgrUhnxGFDdz
DeUZtGalN3hFIa3JnpZt57y9oXQS2xqoP94ZF78ka5n23C0AaRvy3cnPUEV9+CJ2HnMvXBgw8Gf9
OiFv3jrFX/30kxm8CLEWqC5NFrjRrzcBXMnI+wV2TwHsbd36df93fC6U+LPxMgdNG2oeZpdubJK4
nsouWlarjtmR2pSYb/+n38PJ4nb894WheeA3RdzlTj9x8f3QteKoXIRt3hBJmVZLJApx2xjMC9tX
dp4taAwmx0f/A4Xri1tDgIqU1K0TTn6difAv3PoUoqBz7ELoBN5NaXvvi4AJ5UnK4de2oLJh2F/7
oWwdbVFMzUcl7T7fRBS2FudGUNNUnkOdRew//btXbFinOBH4ZhHDDMoTWGA0e0b3Oa1xZZYlz+of
UTRF4D9fn6NhoijQTP9at4PC97z5tR3IMB3ovRUbpJZYj4NUsvw+k1rkqM74I/Mib8QteQocfjzD
REmt1+/HyL/FL2qF8UFgH89kYOOu/H44EgJwqpFUAf68VUUvSK8fQwPWMOO0FntQlI98pL0fkcB4
29/XDDddat6/ivtO250iIfGE/I0ikVGRYCWKR0jGJ/OJfrkxvq1qrSW8oxdRSUY0b+Pi7gECdNMV
TIJ4t+Wx27UuomkvErMQbIGf0JHXnU8ehdPxp/IOxc4RvSsrWfqrdmphS34eJUgGskKEkNdnRwEE
OxdhDepn1cL0mbdyItS6rrJgdrrC1OsVcXaAZGhQGmowJ37We7Hy0oNZL8XbNpIQWR1w3AK6+5Yb
QPx1s7VjdKbaff+XTtgO0+WdHyvM2IOHZORzR7YXd6WobiPo1AdZpKld8vhpqZZDk/k2D2BTXq5M
I/LD8MX261oDhE7WCFVet10RGLbGPFMuzmuJqwxv/2mYJQvdQFHbIaUhKE4Jc41DWtuplwZWXCrJ
KHm2Ofy/5MOJ/p2dyQ04G3Aa5g4FqdN5cMkRNBIZLA9XJv0zmIgSdiCEZfb1LbbtyxEtx0QabF/y
vG8oR3NX0qAADtglj2xABqboIpiUYbKF0JmHPhSA3F1jVaYf9O0dHj6By31tLLicprxEZw8V7NRD
XToR/NdckgLgRVV+WoijqCEq6vR2ZMymMePffl5FbA1NfgIS1aHkk4rbA24XHkCc/lVsrO1Hdv+p
tnp/L9rwOk77UjJ2XJwoj1EwJdaNCxP3qUDSPirwVqWGCd3iCsDYv2WURk+gOUemJCyWzK76j0UE
ImDZ3kuKvnQj1OWYxhajZEJzbtOzFsfIYDNbxnsLpFFz5w3gQUQ9krvCwsO7Mwgg4yCseY3XJKuQ
Gcc/GLu90lRRwTeyLqZPjPqDVLJw+biq32+NQ2B4XNhkyi/8sTfjoErByOKGpv8l+qUqwZ1udGla
Y6fVVGHbmpwgt8MIjx1pXgcNwMQcI0yU1WHPEUL37s9Tax27fpIbPSTvq0DalAefJAmKpNujQETb
Abu/YIH0G2vCu/nkuoXrln70Ntt08Zmac/E0Vs2GDSa9QAg4V2932zZfeRbX7zlRHOL5KQhPA7qc
jsOR5+55WZ/Lv8t79EXLcx3vKnX/Tn/iDfABNmez729WbyhzfhWVLza8zYeUw5GmHmmclOjlSdC1
EIHUri1kDaPfdrz0pTfvYpbANylNXKpM8RFUcV7/EoTxTkPpnBzToIieXsRyslTF18dnLmFF0fW3
H4wLDZAiL9NimzvEiLbzeYPWti8uwGxtx2lcvb/R8W4TFvBvj2KEhKssmnGvmK12jTnyKZB43cjp
ROj0cgR5XS1+W+xmveWOu2cAZhIdhwW2HNgoWqG9EZlSiPcGX9eHInx5R0sMst9bZM7y0m+4dcKt
5gMJ+mdUqlQMPZpMgt7RQRFRtfCAUUtp36gGRvnVjHLXiUOeRehCYqJdD1elFOWuvq/dJminrHnB
hPs4EUY9GqxU+4LFKysD6Jid7fGcqTScAyGG8zB+Ee+CygHnEjsLwJ4r5d1l8O351qodBzqXiNgt
MUMqkDOjhepTWFLXrwnbwyEGGlQ9r2cK9vYyRMb8EGm49hQJA0A9SlEK8LOnxgFJll+ya40hR2dK
R85XjOfjp5m41FmX+Ckrn+TeIFyck/FYkB8smxc470rPISKOT7AvSkir5oGCWXUITnDNmOne1NVc
Oc289falkpIVyu3WNdgN+6Hd9+6XTXVSJuO1wkJ7/l3IY78C/ADnYpFGMi3zLoWxEobNh5Yl2119
vpzvfB4KPALdSO9rfJplTgHXR7wN+72TJB+JgZA1Ar5eIU+J4PUzRFR4zkQOVr4ofbeINvoSr4RL
RcvsvRn84m8XgaxyMVXjT+EXpphMgyjMPHiDuYUe0z7DzkCs2wrcjGY0Lk4yH2Fw63f4Tle9MQcS
4+qQAxTueX2kqoPtt5xIFBHczPbpNLvNlOdX0ffP8I3qeWQvgOtS+i15zCTWXTnfi0bQNZdxLSw1
r5fjOk3RmaxFK9C/DaHzh1cTLFd2MtUvD0rkYOIwCJqq9VLMpPo/F0VC3ZRLxMdkHfY7/sgB8RjW
67SgSqL8iDLafQOwQsVZ4EACOge+6sc0DyFCwocDG/+iu7q6Jq+/6dwWM0FICvRrfYrUJoXnu4PK
/PcxZk/7NjXSNEv7NDzNRfZ9ncC9azjW8YJBHZg0ltwPTYmSMT1RNpO9tRQKohYdMqOG0gtHInb7
yfMyK/FHwcUnvDOk6VL2Ij77sSLhMSFMeb509zu72BrvniXoYKWP0e15tT2W593gvtwNuMq0Rc5Z
2ngJzwvI4z9HVWfNwDMDqd7GreidH617816y2VkMWO8kBvqSkozPqoufDlGmmx6fICTKYSmE7IoP
8CDj96uK2C++QLOXcTwCb3u3a1GI3cdpN7mZRrHRKYey3LCQc1OnlKUir/NSUDwy2s7GfXBQUstI
XxlWZUCxurMM96dI8Y7qhrsCi+bsb4kGYzNH3pfRaBlVairLQjIfx9pMTKoIGXEZJddz2dZln3go
FFCdErJRjNu9dTD5GovRGomi4rEcIgzdCnRZo4jl3mMvE/qp/2gnMiIOW/02sRnB+iPYSm9fvKrI
6WCVa2LcNAOAnQ4V6msbmGwHAmM6T0XM5ak4SHO5lknRRn28r4vWQCdsdtypRpmO0UW1GPKlwb8t
vT0LoR4hFR+N9J16UgXL1bsKUe+9k0LR+fTDBD7cr79VUJi9aSJzZxGMJcMXjtDgJq6u/637Kwmx
07YrBJXWu8pzH8FikV/XU80VPb7YzPPE7lVbJO5UL2IXwex4cts1TTbtDPceJ6WGok4MW7xDjEn8
GJio+PJr4YAXHppp9ve4lOe0CcpMO4YVb6I0QN3RC36U99y3trhdvR8ItvuOFl6coaWuK2kk2VKx
U34JtzEYDyPa1Xcot1aTVej6JTFXYyfmS6qviWvCRJxqFs83MasLbVLHx07LXqJQjIEKRWXm088I
KfEplCkQvAj3GRSMVbLuNFwGb8pRiH6jfPSUc/CBa+PlQPxXX45w6328DUxOH3enyQwHmh8PMgyH
zOzGE0z8aIjhH+ZijsDhcYtWLdEyTVoYPzoG//oevQDiYoi2SjsnaFhZYma0Os8K4q1SI3Mm5vc3
/uIAazTPzVT9gZeApS+En9eWOoiMHmPBeNyjbpUlB0hpAPeKxGMiGMRZ91UtdR/9k1ytVgg/2Te+
TzGRuLrcc8dX9enoXcJz2wYiza7nlT/HU4um7F0rQ3Aye5/CP5PGnTpY+Mxn6BVu8mBq7QcUHbDC
edYTu3MyNRwuBtzBSWmNG75CS7GAIWBN2WH//RX0FnV8AMWUxtZ+DYq1+2qbPzwUTcMRudODF9wK
MPV/G02pP8Xdgi1h9iUw+SKk45oG3ssDybxX0wLdJjwz7/D75lSb1Ng8YY8I+49fnqDaupMFfpH8
lvdJu3nDZ7joZ3iQLh3mTwAJKnNVlMimxnHxhv9oVK45Z/GEP1/pZ7gg14oxZnyWioCjpA/iD0zU
8iTZWewkSuyNQXq5A+MVPkoP1zOHTDYvpCvWeXxcaSn18snZRF5sTNzCNJDoru3jVISvDY53Qhqa
GG/LhhVqhBksFC+GkQhQhG4uOleGQhHFz/Y1Alhrx7IWxpbk/ShpHL9TNTxMYuvw74I7IInOL/V8
NxUuYIs/vabPQdgxx17ob9HLOr644+K0wsiD4CxNdH3zz8QYSRZSeygnovetOvtgt1wG6O6RxGKf
kVVL7YaRBkKy2SYnJ9gosseWLU9o9uToipttC1vmZdxEg+r48Oh4Y9pVp/2lzs8nFCVr6d4wni3P
nAbsnk1vID1q0GH0uPPBKY+m5B8CDi5y+RGXSDEp8FdL3RDlC9Oi39RATLCE7bgDlS3Jqko/8U7m
e+sn6nn0hZjWn174J7DQQHd9by3U0Nlap7P9yPoEk9Ww23W3rsX0RlA8p1CFu40qZMGlzMwq5D0e
JwXMe0e92ZMmlEqQiJv9lQZiLkq47xuVBI8nL/ZzJWBf/4qX5qKfBxZBNbczpq2LPUNamzIO1X54
MrhrMdv1ByjxMFwioRJ/CO5OwcfTujshmrkO9x5vshjsdrLb2PPVxkJDQN0/HQo0x8NppxP586QW
ZT7/duVplgcXC2ZQviv3VgPWCZ7deTO5g3avsY4JbXHvotU3ppoJvx3Clk7Auxu0Gl4GloZCBbO1
I+O42m1J0AXD9VNG94JCllEz6pcJtaPSoS91oNp9p/xOEyz/BN1h2YB78O0QO9BnVRZGp2Aw5PEY
bjIdVaPQM5dxasAXqCAFXDgE1nNsVRL2QKFMPwHXuBNYL5L/ImVRbIIsiy83zIoOdMjtZlTYobCy
zyf645ASOdAj9y2AE9DHL4zfeXP4idU9y0LxDCw/PygtBeux9NtjwZubShPL/jutJvHbHqcU0RZ9
Wu2eqhTz9KP06SM0rGOU+3du6raONtk5FDQ7B19hRgw3meQvnjsPTqP7JE9hRKOWGhItNVc1u08z
zVCdJdFx0LtQRRGS58d7ssgZahXTwgdA7IvBA0HbPtHfpihWcQpBxQCoJ6RaKPkPRt4lw173FdgL
JmROS95+Pv+X+wG14GLlLRKLk4lD4XEwfVXm3EgSmiQPEJrfB0sYqiJv/5+Jjo69Tb3XiFwo3an/
/RAUsqn/kQqvx6vVehACBOQKZaMIY40Ygf4b/ZEHVe7l/ReDEFE3mtX7ttS20E+JQM6TZ9QdZIzu
+gK91yl/lH8SIVtcL3UxakUbKpLbaeB/u3TI91OaRCSrlOqVz5NSYms4vBYhlSO4Xxd5KWTfK/5G
FEmmQFjxMtEL0fYem4wcjeN3ZmC5c9ESmhHD47lvKFhfVHkG2zSVfxLJ3wHpNj892yPGILtNhfgN
BXtCMkUpEj+p5x2f3VcfjcXCKulyKaWsiWbG8+X2XzqhcAA0R36VgS6zjntR9UTf5LGXKmzQXj3t
wKWjRmbRHo1bAnXmCAjOhiNmO5fENqKc4/E3RMdxf/hKBuNMtnQ5d+QgN4wUlTVNibSa4jtotC6o
u9mGNgim5I67rg2UHxtTUxFJJmdcRsrosILeG9cz1fEf9M0DeEymuKTMI/LKPwdl1xABklVtxnyN
FVKJNnH7M9w0scvNZPXl017ZCbCuKPbASMp2oIfj1gwSJpqXx1/QtBRA2/5BVjGJoL1Y8SC9+JHQ
f5ApSg3wlwVcBC7mK+p2UZVL1i0owjmiAAkPDWzx1UVqv6mwRYqnXsvep9HOo/xVn5ClCyDBC+l2
fn+PXub/yPxvxI1IblpHViHt3LvCxEKtnVfnH9sKnzzsgEefcY5Yol53dPmge0DBXUiQ006H0VjF
fECQR6FUlljXChxlCBwIYdF+2f+Tj1puCZf1r011MwnxziUAOUGAO0O16LHJlLMD2zUKwuNVsRKr
SlY6hCRaBdpkKeQYeYZcyxFGgOfeT6SSQIYPN/sjgLWaCWa8HrK24Cidn45YYhvREhejR0Z3sAQx
55+PlBwk4wAaDIQtg0aMqE4tLHbq0vY7mZXMMU1xGkOguO6HAYIqQjf2d8YeyT6bLOI8gHdPLYiT
to1P8kcB88sEH7w7t8gCAptSRA+RdI06PQC2RlutfW6XScUCwS7j5UdV9QddUHGwtQNDnNhQPxp/
J4p8KFPJqcRNFPfuc3tfY/2CMVQ/lqQA2RIv/Ui0cVkOtfljGRIqBorXkSh14xwV2YEN3opRyDlw
WzdYzKYhtI18iNLVgjbvbPo2rn3KGIZD3CrwNN4z5HL2/iewNjiyllmPOKHGcdvWcDP8AB3rfbd/
fnASzAT94Fjsb0Gbf8UEtKwJeoQ4Ee8tkOd538F+24xE7AyQx/2qh8KTg/WM1JRD0rxTMz9NGYhY
EIFYqfMAEv0MvP9dZX0XC2tWfE/wD6E27439Sgg9zViH5VBvE6Ky6T79sNuQ+m/u0M1NWoh3htAH
8k7fBSvUYRgVPwITwAnih6VrPWL5cf+czQsCf29LAJx5maSWe+u+qkBALB4cISuedltSBqo56Idx
6oR7VI41PFGZNLtkvvACiEq3z0q+BIBvu5YsDDh7AnP9VOCFfYziWawqJJ1noFLIAKXfj9xB53Y4
R4LFKxaXA02Jm80ZIpuV9IK2muvqgpf8KCB1WM9oiPHVB/uvTCm2/r7LjUiqFjTdQmf1eYqds6uZ
xvuQfCLTp9cfk46AEQ6VwolY2bjkCDPISJf97CKjifTLSuLSonbT3dR6sRR2DkMnEGpOxElX31jD
rX7zWYSpX+rXteZ+36vTBW57vxd0836ZTkX9vYCWEdpX+kxl0ft1mUQ/3NQJfYXLm5lnGIeifk65
IarfVePTLz9OFtZXeWXeBMVcm1Z2+KtlvCjiwR8A+PRWm+bXRLsFM/nwRcx3/IFWfFhCUEVU5eoc
AydrVLHOmvsZTyB4tCw5srslIOfPAgQisY5qk+sDLGNzT6oGioPtxmUrqqCsN+ZOf9I9Mdg8+BG4
JM/x3jVdrcKBpiYPfBNujklm2O2V7g35Ma4zbBFM4lKctRznyr4FRouwkJOdWrS0EKwx0gHWDW9d
C0ubkSKU5BlPZpttdR1s8i5WphpXhkTY++i2nH0iBQn9bANQe79wPzfFa10ho0TIWubqIRBiWuuN
8ASUq1g5G4rkT3DcPu1qmgw6X5NJ2g84aqHmAiWuSY/G23p7s1RxBPwa0lKMm/1V8TIkwDjgu+52
RNDZqY2cpRM/QHhRtv8T58hxH+7yqPSwsQgU798hwdWxfz228jHV+oquYGnZ0802Mcz3ZBkMkpnX
oRXao4o2F/fI/IJqgTeRrN++ygxnvJBP5FGG9/12ALdyLpg46yAOKqeVGcPlmZwUKI8YTJPmBMkQ
z9LfUfsNYFcH+51tH7tt9n+X861x1tMkn9C15G8T4Ikq8LiqKTeVe0HYZtno+9cePxPfLEqII4D5
tsh5dD9NANBleD1Gtdg5VXQcEhZwzvks7G9lM+D2qH7+E+NT/vDqkhKkKtE+odrbk/cxYV8Q9i64
7/ZYkQ4wQ4Ax6UYKB9WRKRk5fu2VQuAoMcBj/+rpgadUyIRrmDCWlkcEKEXVb78HQZyFbZfs2ABo
m/4cFIEdRiIXUg57jizLbDG3EHtrjtzyl4Nx2bMoQIWtyFCL9IGa57mwF5CgYCGtjl6ZJh1vq7R4
zqxwAfpl8BEeubOWs2/8+wARNIjJ8FL63t8xMLNv5vew/gQb/Ga7fEnZFu9Dg7L1lY0Hf1+6k1Uh
KmGUG2j+Nkqov/LnB5WVR2Nkv4NHdUBtz4hFIwpiI6ViUoiOjTOGRloxYWxHU6wro/0xH1MTflrG
yPltydGJ2Y6Z/DI3h9YvqHaytXsoi0GYc3g7lHbfoNFz8VcUMZE6xHV/7FGAz8BqKEb9Fi0wDiTG
2TJL+kwh8B3ZEm2+Fo+rHrtSg3lHSRSqy7/Wf9LV1eSUL6dzSxuYsvg4X074tHqHV+R5vmsH0+ou
imXwTOnO3MZ66y0FDyHCYODMrW3eZ8yyNJ1AxCXUjSxJyzv+Z4/BMGwC3o7AEwq4F4PZkx9R3N/i
VYnMEWBMIQkJIWNg1nS4qQSJZ2fTkR7z4M0XtZIqV8OpVpP01cbzjub8zM9PMawRLm7p2Fm/euUP
VsKwOG5c9TJCB2EhFbTjf7har4C9BffUsRY9Wy+sFzEkhmPY8twTAehVwmMbIZvUoHG8F92tBo/t
Ho6GXy/i4kwW4N9pb+DhHsnfonxw6mmR9zr4XNFVct80+J+w6vZCUDbbGwxAO055JqLlthVfq7ui
O5i3E18fRsgr8SrzySDbuol4srtUBBlyDLFRyKB9ZpDdgWg9vLCwOGFGhRJweG2A6sIdalrGrCNA
957ItoTMVeYFf+a5aFanHkX8OgoAnB7i0n2gBbQcrWlZCKi1+XWVMNOO63Jx5R4DSDic0/LHeSJB
qKORWrafpcvCp2tUxnI05wL7pNvDSHdnOhuy2MizYqKEeTm1QTZWIz3cQN+h/tbQlzS7lf5zZO4W
dgJHlSX2IbkrIU2TH9pIqPKGanUtMHqx0acvgMMnbfHSgrU0adP/yPNepwE86+0fRTVVOf2BkFpx
ySmR+MMWJeAmLyJy1fNynexNTm5sD2jKqTjECzNzxJS2q4El0QkclsKvgpF35zsUsRlFDDXNdn8W
hAz0JZjCJk6WuJiK4le+J/zY04i3PB/dJ6yvOd8dtnNYjiNma6T0+odWCrEojpP205DhxfsgRyHe
/okKgExtiFugD1Tf4Laf1gv8MoU1yJMlokuapLfexj1zxmdiDxf25T4q7UlkwocXoVgZ6xt+IaIR
9ZQuzjsP84HphdS0F2vveLh8dwi2eghrEZ6cXLvMvVNZ2XHFCaC2Qz8JaDBb0u9LgFqPIGc0EPii
v5IrqJgZngNwh2K2tSrUnU0MEvrV2PDS0n7QYJGd1OX91ccN1Iy44yBCoMTmm7I4XuIJenaMQEr/
ZgXovJ9z4hT5Qcc01yXCwnonZE2Wtfj8fGFlAXCrrzUyBsht662k9lRQNtjt63ZGL6YUgmIzo8Ck
WyXWKO4fUlfXbfq1Iuy/hbnd3EGWupEfgMutnW2Cblwmz4WyWHMKls7z/GcJXskzYz5Hz7Z2ZVip
JeeS2R/m5CJkAxRXgCUh0Nk+yT93pNu1Qd38RfHCNfF1p8zK022kOWE/VMZeg0RmkJd3NT27C6qX
9JfGSVLBjuc6wVF47h60Wjdi10/dCerl0cHOeOhbqJhuxN/A+24DtAl5uhhlUJNe9aFS5Jp6V5JD
4VzU4XPpLoW62LYPu5ZO5S+yJVqGVKBbboFoMipeeN/biym2Qpl45AcfCxc6Z0Fl1KlVgIPGPCQx
BeRWYCreXSC9sD+NIrodYfgkQmJW6IJZiVizAl6LISUHea13a08kPq99abDkBMlHMe5EWS/9jNk0
UgR0JYRTBhIi9Z/aJOn6liSRSC2CSkJpTyUdFw61U6/OKiiaHoW5lLHIC1jTeALdH2X49G6ZLGFM
19Y0CPHttwfyaOOGcumU8SPwuSUioXxdOLvHbV40f/2kvxYXeomGFvLZ01zq1hUmi2XN63bFWiKP
MQl71XIWTRTRceBKVoVw/wJNzTDHcW+3+474SIo+X6WUuANu+45B4w1wHAxq18+buBY0V/k8S/pR
187JyBlwnaqdAtV2Kd+I3NO9d58CGX2DhLWJ6lJ414L+fg2pfOFtK4dmo5pGbOHb2/eUKmdtzbH3
+G+Xs5ApweKXP2o/s1+OIDxzsbx5TbbO2j4nj5nOWbkdErx+bNtsS5eugXcLFIanvgXgetSSNAVT
5Suz5nHcXGv65Ov7vFT6IiCdsRaYd1rsjLDikmbHM9rWT6nW+NWZHi4T9U3tmZPtaADz803RPboM
RDGVyExaOZVzIVjvzxMb6llaPjSNFGfvApci17yY5f/W6qal2BA8TxjwpFs6x6flkZu1l4VQUgaz
nbTowE2ApJTDDUp39+/xeQtOVaF0uRYh7zQxSm7zpAX7ql1qpHnZoMXuxRCvNNhwZ0Wz5S7jXMiK
io0bf+ca43OsQ+C2LT4oQMk4FZzqZiutceIjQmhhgspB1Fbuohq2wOlYOJKPRa0n484igJyZEUq3
ndLSZoiT2E99xyta3+ksJNFr8vzhIT+fzCq/p6xmEc4Vs2ThqRzbZ6y8JcVwOAbTJAuY9+USyOFy
bOjfkrhkeswp2ruugFsZWS947Zxg8JKOEQxeYl7w15fhYuwgt4Z/9Vxx0nmzqFFmzbr3qQClmFVV
vgmsT4c/K64Ujyq9BLNSjpLBh8l9zJADu0YJlWpQZIHp+NkOTyZcys/gknQA5RVrnKbfwe17Z4ZF
2x+66h5Bg+zG1oQGXV+kc/+BshQKKxYYruCoYjeosrK0nBhZQ9bONwjPOIA4jZSu2jqPn6QK8Oj/
UWtUJHDfa0vIxDkJVhAWlIw0mZTCZ4N0DcdvihE2eQYStGkN3yj4BFOodJP89X+zZqcGkTcumrQ3
WgGvvdMBECQ0qSrGLm6B2a95wqonygs3FYxKblCGqj8kU1G2n5FdclBpToFi2P7ww95wau7c7rKY
o0WZ+JrWM5TWmrPvdoDphciznnXEUJsoe7T4zPxs/Vh3kRek+xfsT6fwpVYHQneRthQoircP96JX
3CxU8pQz2TMCmW/lY/jqbcq+VfIxbSYprAIm/FGIaQARCVHYMwUHEu3bMoTYg1vbl3+iF+B2Lfjh
Gi09K30VFyhv1ULEo+wfl7lE/sSLTVilN5X7XukTQyRAk1HOpzmILbmOrRZ1pBlRBwa0dhSa6R6v
IhbG50wGnBv51VYGTaSky1lUGeB+EfgL2xEc39W40L4zEwdnxfK5B0cU3Dek1R0RVidF/u2hKisz
ATVMDbSEZ0f9G6i0UblAwKMZgDPW9BDJfJB5pbKqnNvKrvTw5wiHKFP8QFcKPf2VpKhjopOuT1sA
nsv/JjVPVoJBGct1rKRjV6t5v6OEEQIQ2afiHpNdWLII0dYRYjl4t74/L/ByPYxEigOlVfuINZqo
JLPejQ93QK55Sk2ADMzKUy5Ow2e+6hMcb77iXsUITMdW8Kx5Y5P2cXEVfBQX+3hY4MXxFIrPbmqs
8t9JVKhJKgdh2WDc5QllUqNvNUwxJhPs9hL68wGZ3PDvivqeYsgfMXK/z/LlUkpu0ElA/OBHbIGW
hMEjrj84Erl9dhZCuPlqKu27xUSAp7ax/+HrEFomC1/v9o6gOUuZqVsVQ5H5By+iqC+92kfgkUGb
LoEsGFk8C8Vrb6Ht1KDf+FgFJ6+bTMn3/w6CtBEB3VDdb+wpGKOyxa3zm0kibc1s4Fo7JOxbK/O4
mTPlz5Cg1tz6nQFDumT24lzCnd+NREt+NcFeHsp8+eCxJ1NMDiOnPjIvKLp+W177GeedBr0XWtzM
ZDXfYddL0gjXOHtLngcKIr6Pxut90U0LUyCIRnIo9++QKU2R8Pp5jpU8HLc1UN/6+qELWWpfJxWb
qf4Ct4xihwtW+xK7yOweo4pJ+N13D/FbbagKzpYGdSl4rV5Mw7C7jZkq5sDa2QBaMKpDt9gvCkU1
XNdicNSd8jFBP/WQd6ay/KC08pKEebrS5ea0eqbixdG4+58+TPKt8Av4fWtnchzt6rGMfc4ogLLX
TFmsujT8RChGbZB1L6Ga6CN+0+yRdJdoSEV5eJQ4gUfihjG9CPR8N6Svt1UOw598Z+FWMoJvzPpl
nUx3E6sitQdoS2nU5QpZkIfH88QiNAR4c6tSDj2YWMxEE+dw4gBXL3/JSxXLEulDAc5/acKQOYoD
/Jqr7hhFIxj8locqID3nkywe4NBq2aeLC5YaCMLGoQuqL/z1PeRIbEB4wbApd3cjiMepWzZ1bu7P
siRfEwKlJYQmuRlxmvZ2AQXPRfZtkJAa0EDQfrTQCdKiRLzB6KNi6yg0Y9X3nkMRQ1PIDRSa0Ats
JmVHf3auNCGyOFzZGtao62I0qqOyQLR67YUHpfrcPilJ5bzw5QX4i5nXRnSD06+tkVLu9NnMWkVw
097o6fYfyO+RTUiyQuaWLXP3WPMw0AeY2JX2XUhKGGUgTK9o7bDR6It0VhKMnlerWHRAGLO0tbuN
HsWhUjzCW+YIhaQsgTX/Rq/4WRCDDqVy7ZyshgZUcAXgm7S3PTBQvoFxgqSLQ1RttUFTXbYfWd0z
gE8IocVyNj53V34uwKY3nTY7tAlICWo8V4rdniRVgeqteqrdcnhFNs+RyEi6vzNccr9qoU/Z97xv
rxDb8hVwMYqy2AWdeHnCLug+/wz+WDwi1XcBH1MKn4iGqW5VP8q6T1rrrPYg7mvIXSinIFPCy+WH
sZF9MJ6pbasXO8kbFAoBmD8iBAHDiDYFYkcDDNwrJO9Gfc1AgkSzGoWx/s0P5qFZPWTEdhUYaLwU
jOnlslmi7NOqPLd3kA2km45PUT7ugukgCA3Mbzi96MnQ7CMXlXYucM9qsDCjEcYCdXg4XEJMJEdi
LFT4Qb8cFL/cHwIsYksWWUzln7suiyhR75HwZZ0DFrW3KujLXMZCYLLYd2iHIpU4kKeOuHcCNA0J
PDmIeDdr9Rkhrni93+xs1JmQ8pCxO8IzlVUrahkhZsNevx7054b4XhkIDWS/ysJ+p10DSlPqUg3F
Vsj4EyZ09OPBtBb6FychmGSf6oP9mg9bkf2yrogx0rzONrI1a3F+NeC+6frdON8gxFqxAY4nlO3M
FZzvGkJwXCBEegtAAf+VaNnvK6YXuEdXw/dRd1i59YsaVxisMJdL5XHv95RGbmagE+OaiM4XinYZ
gwruI1GYA6WhBsQ7HeXeNPqNNIo25lABy01n3Yo4D/Xkyymwp4fk2eR8RpL85j2zZ8/c7ku/yb2+
cZUMSTn5uMTs4CDYLGuSuw9aeYLntWyIjURiHw2t9bST8N2AaWX/aEiD6MUPVrOH6Y/EHvDHxRaa
lpDwBQVgcAJVqFO1Hwxcb9ksvWQpKyL8ftXK3ES8zmCB6oy8WVa7js2JNunxOKfBRUJzKaueu2WY
LLVnRXGi8BeM2Rwi2mpt0hGjVSFPpD4bR1k7Nkhu//g6m8NFOQt5aSesa8MNd2TZHVejCNbVqIgL
PZrlYuq+5LnlCImWit/qS4yo8YTEOSSj2d/MiU+PclRItX5xvdyMkp7GVaseQQul3KrbiU3RKMVc
Z/WMSulU43Uxi4JmCvmqnvU3eNKwu74uKwyoG0KsFjaRTitKMgswnSDv+a/byuNqUB3DGloveFza
L3WdVR28Yb8zOZtHXkM+C/yxLEULboqEhpv87a05P/IsSsc3zDjcKLS2759vLfGWBrjjbox4xPtH
Zf7DSUzZe6Dkf4EWBtC7zvkQbqwVuaETHWpZr1OYtKuzB6n5n95plRb6Kd4WiiQTcQKrPklrj71x
qq+2rTHhIp3G5+uDgByvFEzEhNhtb8ZpzL8ePtX94h5cIqSyY0JFXto0bFfX6HZsrEbxK0JXpV6U
kD5kEo3Zt7PyfL4ZFM+0zQuppXmW3eiqWEwspVt+60TfCs8dvpul4oR6/XdEi5O0hkWxJctOgOq7
cSfTNxEQUFQoMzZL8WhhjEXldj3IpLqMG2lOAam9Ekc16RfNrlFQxkv5XmFR2RmflwbxV+gqDTCu
iFDlGTXPOK1jmRoKVo0DpY8pf4Gbc+ne9MmP11o+N0uaVVrDYEYciUhhWFKjmzGacajOw7avfQGB
ruBXFFQTMMp7JArUBdRbrWqnCQaXgZQxCMUy/kjZv3o4OU6iTtA4j8pDbsuGmhZPjDdBimeKvUB6
e2ittGDV5h8+JkPzz9NaU+/Xr8fvDPa79aoI4jWOVBeBwnBhG0E8rGizpMXKBHjtK14hS+GdGgoW
eQdnpAjaEbDV82u2/3pkaE0CHMUl7HeZ4hY+ev//4z9Pv453h2WvPjAgor0KtnFPgsRMNpxgGHWV
JBcE0IiDpWqbLwfj16a9MMh7b2pmDP5RVodGlRbDDhKNItTzwsGbdtW2LHvUVQZHc+2KuVxUWrNi
b191l1zoIrvki1cnuEXJuS/hBoK/quX/W29YaSDv1mg8utM/qWsPkfxECibZb9FC5YLY2UukC952
jRcN/8e6WvPd+a8vtF+kVs9E6/LRLuV+h0fRjAqqk6e7sKtttVGI9sTXUvP2wy/9lrsfZDmXBfHj
ZoirXIupjvTSE2Iu3x3BAkzRVdLa2BIcmEKxQnripTL+XrwdFerzcIFkrhPhrGBJKCF1A3Rw2duE
rmH/Nyrn4vVqRMDco1LcJUA1Ez04Hu8iR2v7KFI94BWWGPL9mXCy0RynlBvZcpiFR13R3guBZtbC
u3umuwnt/Ml07jEPLjG8zIASphIFsLw9/lK4vkMHDcJT5HKdHx7algYcZyEAucRNuKQYSVXERDrv
IW4Cu85BRoraC/09avll0ipu7K9i2i97LnHgPPvhVdaiT/C9Q++EKPQuDMhiUueWSyCcTT8oGX7F
cydEgHgYowfg/ZBNI8FCwM2Z7TaFcSEQ6u9SZrBKzRSyw69AqbY/KBsD+GKrJBon3xoVXgBhGISD
sZCTX6aubUi/tyyIQrsydLCGFbxECOKnOmGIMpPvYEGfscmsZcscKEUjDtfrU2uL1XDoxOz3C9dd
qeVISm+x3m/bn5jElaFPS3d12QXjmNPNy24vZTwBmdHVOxxRW2tBnMXpy0R4H1YvfCJ8/3QACjCe
uHfBnzkILU8sQPXWtsDSsRtfoVB4v1un7wL0GDZF538eCnuADfXGBZSCS7rq3lyO8ihyJYVifEDs
G64Beezq+ptyMULSkIUIepqvvNrgwPovJCa7IrGIybP12L6MH+YOPcPbLKAH5Abwq6O57Hoazmbg
nMNAkRQ8uDTAF+PSnXyQPIy2FHire8x7BE924rQLGyVNyMnjcKovDwj2ujcVgjRz7ZHCAiGhKZSF
0CHUfCgUEY7shT4NtZcjGT2jUWnuOkJRmIdhZVkWQU1d3dzDs51/cyVbTcMPywE1u+f3vB19N4n/
JCb/azJNn1bhcdBGzMNfBU0H4TNVy5pDh1lUA6nlSa8ReHjdY7zs7TuduRC6jWuDp4DvSn2GE88h
qBD1fxqy7bOVx1DmWyZ+OGVvMltPVycCfDxtULe+AqnJ6mvpXOkA5wT3ITiSy9fR41pyg4JVb7RE
Ax4zKHa/vUJUH0B5iRUcS5LFmUJdTpLO+duicErU4qlk1PojF6NoLhlvD7pxNdqGKo67LUkPNkpn
rSRV0a1PHhTNBaask04hus+kwRqD1LxuFVNYJsLjy6PhR79AX/Ye1uIv4qCSJ8jlJYzTRFo1Qxa5
CQG1ruHxcqX1wH5mK0Q8//RxqqRtLK7YStTAbdbArfbW+3+n5wJNBNcnxlEDb5waud0P3TXuN4+7
Lo3v5vK8HpE0yHQU2el+DT+pVHQPwqaED02CHXUHVQSfZULu/B+9PkZkx7chs284iPsYkKMMsENe
foXJ/dVtWPGmGtx0zYj57FgYwQMJLUaoHRzpYl7PCVKK/aq2B+1Hj1ZVfDnH6tG4sWPM+MUUWUqA
9qw47hgudUhvx9zsAn3DQOF6Oupi3VjkMHKXxra9Ti4JxYz03NiaPlnojK/32IGP0QPpVw8zmM8H
i7x1QlyFiY6cnK20OYj/c2rUk/9qJ+6OYRaizG4oc9pa0GHmVfwpMP9xiwXbtsMKaRHY6MBCsgTP
zJ1jeg6r3lYSr05pogGMFWHAZobVztOJBmD3Nw5kryT4Pjf5llYBoOCGIcot2SuFnP7yZ9kFmcup
ObylYge2oJ73lY/Mho+m3zwHfbKESD5a2/Tg8L3umcRSeJPPIEtzfOxLQYAZmhiyNN/Mv1bQm8vm
0NbJhgoJPOijl2ab8D3ysUvnE0U4iehv/L6hqr6P5ui59u5aPGLDxmgYeYWFxWrexCxq8T1D8Vvl
LWOlYXXh8vlLiwBMCSE4o5aV07sVkHzAf9+v36m6z5We0FQ86T7LXaYe1BJ/fWG4psl7rlKvH+tW
IxV4YWC/pKnbnIzyX+c8XiVJMp2HT8GGRDWb0cKWK+AGbrHhNjJLo5MfEbzdvakstnAKWtzthvAo
bRYyaqrtSf0KsUyuRy4TdYnLv7Ub2utLE95zOKMNENNvvx6wtMGLtzzdriR1tIOIb8NFv7ShAS2O
R7dKmt8H6V3FLhxYwwf1V0RK8fZBphvT3TPA7vU+mzhJhZqCuNO4yZm7a3XbRBG0iea1wCX77guJ
7xz68sdW/M7PQYWzNjNSqRrBgBVm7Z6NgzVTfrdhGBuvR4kd/M/l4UvrRp3S6XzrMqdw3tKlDLkE
SbGzywXzpogB/SQMXexy2+ouNH3cNlc3BGb3UiUOvYYOqB8Z1+ntjD/IgX3Eo51HWhC3DE5ItI4A
c+XyC1Zy+Zsemqlbc0qKLQ7Bw1NeJZeCw3msoUAgYFu7mPGbHLeOVCyWqPvfxUNt1utPq6Ywh93j
g4NzzEwJxEWh1V5MqrcKZ+dedYOd6ePN85+oibcOEyY8fBm40q7KH08Q8xd7daXgotq0u5Warnrh
W+uvYQ2Jv3KEqdSUjk0JoWI4eTFA+M6wvMO5N4f723mw0WXBah757Cgs+6GFS4/hix5eFxrf0bXV
hfhZaticGVykOAqWX7vSRP3pfhxswJCduBOq4RlRV00rjaSFsMoN3P9zNRZdPOxitgVRTZivLWSq
EyBUMKG2cKSw/7ECKx9BnjmNsUIjuA+oaoyvZGu1QRTNK2L/lYYK/+E5mVXS1s+1nDySsUFjlZiO
cJjPs6XCaqux3oTycbdzqTz3biBf9Wbge2cpEDrN8yc8hs13lV0VS33uD9X4S3KgZTUFC07wStb8
2TivkXirq+mxAx5QlXMAX8pCkd0WQRYaEtfZIsaZnaT/IcJQISa93DDniW9z3fDywRho7InrhvPr
mmOlWULIwWCEmvc+FZwl/MPK16oBqgSP8EFTETYtBXTDxCwfDABmPgkGIAKet8Kxf+ubMGq0W1f+
nzUFSPXO2/ziStZwSOhOt//nq1FdrZ+XssZU5Vv7XfWbfAOqjtiUMgoiIyLX97M3P3et8RsvL5Gg
SVdcVznFiR+FcywDldXP18yncH0ZX8cCI8hLG9H1vYteXks1gYX8j84U2eWeDSp7J/6YDPlxjZCS
i+LaFk7Fr0qE/FjO1UoiXnHWcMNnm5ssseBxwaLOHKRrVrEJDB8HQlStV2NSYFDzHGA6Wg71999i
ljhOcZfKyect3DtOx8/PAkMFoIjfydKLvQcYzIqj7F7FTzZ14i8jcFMYV2lAj3gKvQPN0CGOqYm0
hiDT7EEQIgeJBUQqTdOgbRv3lWvWz1tH44D6eyfK308L2GNE8B6xXZOpgn52WWNyy51jhqooKUzw
SSvR0SOWP6/EkvgQx1Yq0oPbOWO413ZHFp+NDszdRUtm5N+ReMY6uLTjOjyDg3xa21o7AOiFmreO
AmuZ4omTIiffw1qtsOwlUnELf5nTkN5WWVMa7VR1phCTDQnn/trc8JG4/iOqQz2YxZlOomPTla+r
+xQgwtZjq4qyj28LcpDu96QOpVHjQu/THujjylZqZPcAsvJG2i92d4HQFfP4dboG4E09KpRZjlmf
FOpriha5nPlCYguw7lIu8/gAxB0Ofq0lXJ3SWmPzg5rso5AhKUhlmMCUa5yPNC2EgBj5v80y/tRj
/WeYxgxh/2v74hsxee4btIcuFC9QXcjlJlsy42gZFGlYXDveYwoRQekbgEWIT0SYAaThiG08PXkB
dkaAmDZsx+RMD+k9Tsu/x9+7lzfui3X0iL6oBo8CZTO4K5MFLvqr6oNUFlYoB3deOhm4hWdU5fqm
6ohj+UcYDbf3l9MBm+PC1SZAmo9ZiHV56K9vH0Esv4iDz8stHbfUgjtHGs3P31wgBjwndWVUwSIv
gH6hByYNwRxbIbAhS+V07AKs3gW9jtjCsl0d2QG0L2QO5Ig45VczHFP6yzacRBVQfDTpHgjkUUQ5
StmqAeRdDIwVsJ/BxhulEreUL/C5nOjnIPHVi3Ka5IChZRPQ2gg8K/pYXP4EbxlED8FCLVDxqz6n
BJyT/CqUBTVFMBDHp4SshZ7jEDiAqSjYjm5omixLVFreDiavc1hM4jw3tAPmd913++y6mNfJBWEw
FINODVUBnrqtdJh+Gh9KcccMyx9z5axhqoRnXTO/TK58gEOeCfGjNnNDlls3qOBAGXphozQilhRk
neopBq1KKI+0a/raOgh9c2BTL1GWbOqYDh1eIxYg4txH7QlblmPMUZ7a0+o/KTyjw3/NORfBOMd3
gZvPXLyC1tX09Ly7UJe4hbU59IDhQioMRTRS2AghEO8o2usT5ekwyZkTnelN5ok9IJuKB9HBwaM7
Uq5fGRq2qZZyK0rhd5wmWtBD4vQwFMzKCmQGQGiGzZK4NoVdqumu1XYyXFbv4PcKT/dLnPRamUuA
nV9iXwsU69lcxnOb0q95D1L1Z23hM8onZ3siRtlj4rhQdCdq9tWvDXSwG9Rg/Wb3Cbp3n2I8e8/w
D6DI9+EWKVlaeWos9Rlr6VzAApzPrPR7pHfxRkmsc6vQTcGCRLThA5ExQSn0U16fN+sXpsi3Him+
cvZxErkiwcNmVLdge2QmAodkcF4levw4UPhLZYdYNOrBOsISkxFh/gGpIyBiQUziUANg0buLTUlN
oMWtTrXsBt5Tbn/KM89st+1Vxltxijxx9glJ1K+m8I7Oek5aGcSuhCjGq7vfiUiQR+rU+Z1SmNqH
l/yVJnWWdV6u4L9lPWL8O/H91ttmI4lVYshkct4qSY0bDWa43Ikd9U+ijvAGN18w5Ro6YlbdiuvT
czDTPPjY6M7X7+eGEhW3F35pmu/1VtmjnhhEH6Z7vlICxohSaR7HTiIzXFePTcEUEkp7yS3Tm8J2
ZMKOY0aaADLtnote6fC0Gr3zMhk9ZQ06v4iu1YxqG6m4rH7H3lDw1HcOW+/UYaQRKEGs+VKybcq9
mwhZpkcUTHyE1Ef4TYvAlBPBZRpSx/L9TX6IkHACL/yn7R+HMfbv+s2XC5XjXUjmR5HWknNxkACH
el0hTqFLxFIjOgoWYjE/JgZtwxr8IAnEaaa2L/rUQzysxbI9V4yWm3f1rLBva//kOJdX2FOxAaan
MPjt7TpuCcrF+AebiWQqyNaO2EW4UM0eNFi9bMKtoqhVSTsc/7DZWH6I9svgtrqo/hDEk4fD7klL
KgB1ozZ8v9NqSTiTPkBwS2SD2E5hxwxhEIpy0i3zmd9YFOXKi0DPpDiOmSDG9BhLHNC44640xMxP
/GwZPquu1tQxkkHj8p8b1N56Z6Yi5hzrVy+a+o+6qa2QcUM1DsVK0YuKqr/4gpn/ngN+d0EbU2eO
hiD3Og1HVXh8BKzQtwhwSoBocCV8kixtMFtL+/dH0FfdSFyeSU5hKkTXifkBygO0S77Inks1E+JA
7M3YEypmoMTYwdrZVP0/D/6rXqrxjQUeqflxUq9wweJmKHo+t+jZi8XGRKtGzsS8Wc5g00NEOmar
0cLnFVrV1HXOlSBwe/UZ6AGiiygMgIrZpUZyT6AYMEshYfICSL92PIvHR8uDwVFPiRs98+xkk03d
m/G2OYSZDe+W5QEl9CMSTts4oA0vE3dPREAUcW7+Po9IkDFy1GQiVu2LQfjurcp7XBxVPrpOQbVx
UrDhxLIOpQJVWOjmwdT8uyOJdIsChSTWHCP3RyhaF9FWwwbI1WIeKzh+r8FPT7YZGZCfl5uocMVG
+dFT0181wSbuyF2eMv9yja3+O7dSQxn1Cfe/E3zhqPUN164nidL0IDBY5XzY+qcocUxKOelR7ls+
IlsuchFGQM6JLsx1RL9mM3R2qPVkug0ol6e/C/Zx0M24ZiaRyiPnlgPGM3M/Ub3lUCsO7sgV23Ht
qNYdAo0MuNVZJAJVJxAAT/MXjl4Amzsscg6bpp7PGj/ckbzmVOxZFjBBhYB2Y7y11hcm4vI+xPOD
TDOw7COPp+NbeSbj2gF1WrZWxmgT1XDE9icwI0KDw1dVZaRhY67r4kbdjgsiVvoVGogWahv1R9tQ
Ytt+hYi74yLM61ITkLwflJ953IwXdIYoNTxtYM/7MEQyHUi9O3GmB1W/ADzHatD1ugEVSRXrxJaT
fk3Mvmn9cp286xMLNnQ2iykeGQcXRNmdvSqHbOWBqFYmlmubchueFjiBR5BuhhmRmnkvWQcj4qDc
FoDAwaBt6+eTTWhO7jigyKZTjre514Ki/aK2OOW2ojsjYJeT6A5tirS0S3P/IkgjWue+ltojQay3
e5KxYHv4moZHxr4+NvUpo/MaFAVi1Sjg9s/240cE+NWcZivV+3TufaFUB4wx7Aj3NkXzs5quT/Lp
ks8ev3CaxOivn8xdfaCib5SNvNNYYdoIkF/pABDoZ1KntBIikjoaPr147S8a3E0mtLGc4C0eHh3B
1VQh45+vuPiVmwGGL6zIOR9+GkkVptGIJ7CC0DyKKIGlO4iPCG06cfUns74tuOSyfunDHERLsZNL
e0HixUEBdhhoR2Dxjy+KVyk6kmX1i1nh2Lvx5JHHLXd8vdqw7jXpanUwlaiC6ycYIPD/oA1Y+23c
uKk6M1UjtGfWpxPEUHmCTn3T9GYcc2yZLTrtOEUTf3iJzbnn3iAVOFxy0oIA/lMP8ebCX6GjixIQ
/EowihJr2D+NSh9VMB+riQ2gUQWUDkJQtchM8mo2WuFrbcqd1thkVqyD8BcIv5e7DjMH1KkKS1ds
ZNZyMRHzRpTpqxIt5GOd4kzuenfN10g+mEN7++oL/G07Zsi02HkXMt83yhQzLgM4HVEUB4KpD+Yi
1VAN+W7jsFjfW6q8lSScQGP8Uw/yRb4ds5VYOaqVd8zycQDu5O46JdAQ6oxRAL/Lv1rRnd88/cDx
WPH3VVPHh13iIf4I3RDlJE8UrlTDr1nHiaUuccnV1xL6G2v0tPFW6G4GpVBVmT93pv1wUgFKe13o
AetTkfM0hbEZjmCzE3SQ7KmfsJej58AL4ZNX5IApZEqsMd0BNIsBZbJZLeFhpt6v3iQaoN5usE9N
m65oj9mIdcsLI0DDbmXF65QVNtdfA/hFu1VOSn/M5HXfhlEBl96bSEi37N0Qnu1qeEp4kl/SROkN
RTnTtlktWoJbA+vgwDvSdsTGoRQpCDiLQIWReW5Eh81+qX6BUgKYiCvKgyi0sWBpiYHhasgX6oPy
GCrHkVSHmoHMGmrwrjthya/n44Un7d28A+JwtcubopeeAqsLT67Vkej6lE1HEc/c2NnhTivh5kf3
Vf6yEs9fSOWDDXp9IQeTGPR4J5xdEVIIDp2J8Hk5lUdlT/fx1NJQi9VP6RlQn4kcxRIHziuGLWAs
4BR3ck9pTQyCEMu1s0XsqfIwfEnE7JG+FyhS/pHBsHnFmOlN6JvSvR8o5Ukj3t2ZZbY2H9qWmZJl
jt+PNrelYGBVwKTFxlEhu4Mr7plhXmEsvytqzDDj4YJruSOsXy91rYmx32am/uyPFsxYFyOmthm2
X7cJHU2hpfIntwIpOQl32LvIJ/YUDQ6o+ZYpmnx7XbaLiAiJq7YSroJBVa6LClU3ZEwjMpTy1g9N
MWB5g785DXws44UTKi1mAiRPQOenO6vb75mNm1Jwp6j6ch/aQf9O2Gp4zMYOFf7wulemGWp4zgkj
81jzRI7fyTgM5SG7F0WCy6a6IMHhX11ZMdeDxRYEElzjTR3wHT9EfMBcjI3Q/geIMBtq/yf71kIV
Ld01QohvhhObzQRqV4fW2hrB6hILoNxjLozYdHDIDhTx4Ig6h1Y7+QMkbHSXyhxHlgVHE0ICYhNJ
U6VgK8kM5j6dbuOTMPa6B/NY0ZbZ/IJf+iewU/QnVM2Bt8Jzr54/7X5ecnJEHFabuaGqCW1gq6b/
3sqOBaAYo/94ei6qMWneQMywOS2hiQMWGmt9TggG8uYQ9nwI7InVntLeEjvGYR7Zb2DOsxPCib/d
6me8t2c80qwU2ITsbtKZHZnR0DEOSAPp4j+ni/qbdv+uk/Y4BNZH59TX+K8/XxuM/vLOTEVryIz7
zZgL2VtJDixH6JhbAAPPSySki8VPEm+ps4d1h4TPk/wzvFK7vtbCVqjQuN5NIor2+TmsujsW+Tlc
mS83ljqk5caHQOMo+VO0ZOVi9P6WeL7ZJu5Z8d2MQpbKv66py8athi2dKjwrSndCrrC/1AEHSNOt
xjMriCYxIRW+oRJelx45d/ImU507b39Gqk1QGCUZOd/X3G0PQf1r/vqONfKCleaeXsGUNTbScx4r
5tHaUSzHSdX3+xhXeA+Y1yXudo5IOlMzfs59zxLvLu+SetALr4K8/RqEqcRJiwwivzIJFwnBRfp/
Hwkl1QJyZ01NhhwNUiouF/ZG2QBhNMJOYROmC7cLl66B6ol0F9/0VXTf1Uj47sOUhXC20S7o5bLI
qqnJOl9P/hc7JOdiooineYXwX41O0jei5xPMH35bYzgJZ3m0V6rLUK3BY8OMJopeS41RQwteQS+4
JjNObGU5C5JqMSlDKsgRDYu0H9MnWaPS7RzKKXdiNQoOQd4SI2HAriyJfudSJa9uB+MNTEpyXrh4
6NLtNCVgALB3AysyD3x2C7Mb6Uf2qcONMUgPO90xprzUc0Dz/5iWglTb0WrtJzjjx7Ug2iKrHHfZ
dxc3fgWnlCet9NVJYV6gsaNnm3u2j2qHACzv/E38I/O5+r2Y4z+ebGd8jO97IgLArCLo1GFgks7Z
UUbBRukLl9zzdjDrIWLGaWxQNqYVTizXAej4WriMbMz05ui8GzCb3lTUaVuR4Fa2qpI3DXHrjN3R
eCr5Qw6OxVaM4/dZ0Hjl5X0rUsDAHwtLpZzFyl3iEBivO03PpVro6S0xJc+hyobhZ45M3zJ1OmtF
fWyNhfFVhLtXw89SL8jRgRlyJciT7Shj7M6w1mkR4QR8DVCqplDWFXoKzmfRPAZv3hMdhYTkx/K1
RMLuyuPru7EK2Ha7S9IUJXb0xD11416M83OvNQ3tJ7pbWmNMQmPCl27Ln3XbqO47QGxy9eHVvY3d
HH5W5Y1v1X2hvsLJdDbfCo2Y5Hm3q0Wujz04M21irlSiYUw9EiVs8BqulDl7RzgxlRPCnxXK5amV
DbG1l0dhtBgno2X+KX4mNF0CD4BohIkJHrvmXQ6hQ/OUujrkd0bi0Iu2TZtROQGTtVzRCYt3Ogew
jVQCuOWwzxL+zxHkyzeFpSfMktTrtO/5KWnXw/078l11pjbPkXUtOOgclzaFuMWtptevSZARx8Pp
dAA6dc2Tv1SLiMPqXERqWQonSXZmwl3LAk0jNofup5unaXWvJNYgw9s+rJC3D0puaxNqZhHQ9Xmm
imiq8yU2+Qwv6XpJgJcEnWEMvIl9H52H42z9+6fIrut34J6YR/D9AhKFWIPZ45FiqCfhLjRL7dZ+
7mE5q7Nio4gjc5cvOCqCkIM2gxlwOq56FHOUJCMqbZT9zYaxzVeGk5k8pp/BYmijW7pXaFcgUPS6
72N5ZgsTIfi9L1K2foptA3bwU1yNKn4d3wjfvc5YAx0Nw7Z+7nYXbL60aW2RVbyc6+n9dQGJh9aL
JCuAOU01NhX7GB7XWCa3Cp/GJGdvY2mQngUQs7RxtAOWwNRQn+lAgt+i7qdBHhXyRTPkD+gDIJEf
xpmhso8afSPM5BFT+VBsIBtFldYbAPZzkLf7zloKBebkv4th/hBRaHaXivKtcOdFLNkhaBLJxGJx
IMZLBQ7IQHaMWnkVuVnZGD2dVwnUpTZ/tVQl5JKbVRs2EDShB8MgzrJ1E+gdPFq0K8KJyl9Jy07d
zWxd9ZAC8BKFYCvoQp4jwPdf+Pd6QX6Y1b3xa3z2a5sfRMtxSntU7oqbSIofUEVfVbB72EALOQho
lkLZ7h3VviUtGNWHYWNKiEVWqtfdydSwXRUDRguazog+G9P/z0r9GyxrOe90TvizBq+mgps65XiO
sNLVKETV5MCOHzdIoZ3VflCMtFSFtjkJuL5FlLnljbHm2MRnadDb2E2f/pskX0Wu795u/2zQD4W8
8dN6/hpluuY1s05msI/NH1xcW/Cyf4+WySC4Rm5no6cW5kGnQoVrD1tzdhVg1dO2/qeaMZyVJ/0e
Kk4D3yIubRU6PIvu3kfWwNS5zrO4ZMZuUnTyKwhsFu2l+eX27Cs48ZDHD+iySoOTQMHjaVhYOkqA
KM6kWtpnkOT8vf0XlaqY3XXeDS4jUfoqvuOTmnndKxdW+7AKzhcVhzweaHbHwn/zU4fjuXhjRzWY
YGo+2A9fJlY7Bq0V9cgXGyi1SZrJQpmVjZDMfkfAi9jeWsbXYJO9Z9sZM+OSFK9F7n/FQgiFqhpW
GkX/PMNl99ebbsjdZMbnlBZsTojm2meqElhl6E86m2W7if5DUKtzH8hmQ+5whTTcFpc30PjJoi7q
X6swGfuyebB9xvW/7AqC8ZRJxJ+1xu2F5TT+tv9cVnh8np55EqoPapKQim+G0rxKSHM0HBIsfNM5
WfkFNTY6a42ieNp6Z1LnyUZFTR6/tY0hn0B47ClkrvWJAFPMMTZRBuAte/zo3EObom25KrqvwARU
aXqtLsYvFYTAFAxUVgIciaeD7L2awZ8zkrIPTWAqcCiSWck6Fm7A3kxAW07ixzOOass7x9wIG0iF
5VE3NN6k+uurhQMVx2Nz/5uMDNP9+YKStBqCl5JeNPxV7NcJWz5PSsgCGbXa1bRXsCDWr/zknsVK
oCZVJ8Y3YuMz0xmBGn1HColmf54V8NvD67RDh5AG8ELJ9wX2DWC2usk4lh4v+iewMm48QAn5HiqU
cUZSZZcQH7bVxavc70qIp5pjMr4nzMOO5RwUixMG8jx9OD7rNmBJ88y1qGsbpXntwEMzegrd4DOG
knCqTchVOWkmNqfoqHwWI+NXZ+ZwURgp7Xn4pDDE1PWF3yRI0hzKqql0DC378QoLpyV9V/dx+EcX
KRFTHy5HKYL6/usetIKoWr0KEyyddKIaLt0zGeoOHexApg4lLzdXLOOZwYpUkKGwjrdd0kP5nC3B
BSIeGh8NUuzQCV5vgjd4u1zWKHFoIfIWi4yrXNihdiyTBPzu3XQvocCSOLvhyC7CJ72PtMHiuMQF
qx1+g12f/wL3CCefcBc13uZDvqmAotGhBvmtAR1aIa3VhqRTq6y0PGK+uWn3wQ3UwNnalPGu5RQ5
6O/dpRnhvRAR7mrLk1tlarNRZEMO6TxUQo+cIG9bTbTENpDq0fqG7g+nBkCkt0/ai4XhJO4kwNtV
Ny73M3PmmrJClQDqaibMTGfY6Jpz+ssIRiti+7F66zgK5CFfX8l25qDoSZN3JOG4XlXekPP/VUh8
dYg411scwBw2yE/KLvhxyfrfAeg5x8Q5Wo3WQh9En4SLcbh9sIcTQbX8Dg0JHQHpuEfB5hA0sxtx
12TH+drVJ+EkkGj+yOzLYVtTcwe2keEJL0gwqdsMa4Cs1oBeaag5cA4/Zihd/aT27G5+8RsO+Qsh
Z0X3D7KWFiwrRIbxs5zXD5WF4/rffY7mkcWrR1jbuPiteQI29E/h3iuhRqxtbBLpm/RfmnCOhFgd
7U+Y5C5adp64IIvt0hPM+xa3EbaAe6abW5bev1HZ00TMpdsZEkQzoHsEVUTT70HXOckiH2scJ1B9
70xXowIhNqaeaa/N1am2D7j27Wl2kE2iD0N/+qfdxt2MP5HJ8uA+8gohrc1/3I7nULemavTO8ulR
63J7JRCTEMgyO8n7UUwIPgyUc74vmLiCr0Z5odtpX2TaBDQpdDFA2OLZS2yU67D3qdLBnZoWF94g
9S0TcGzJwYkswukrp5f2axot5jTdT96GE8PxhAMyy26YEjK98jK8uF2l4vP0cONJfDPzDsnoU7np
ABihin/Tvmm4zXXUNbLVyWXgn8gkhrYHmdzo3/BVQd1s0ZDtG3/6CLbPP5bqbsvyAvt/dC71+tbg
tZp257yPlt71UFc5E/XBWohNUpsFmhZlAPudZf4NmhFSucgyBIbxMBoz6QZBxfgM5XZVa5hv9AUw
CgGbM0P97TXE5zLLwQYh/J9PeRLI5j8wFZXjXRip5nZIJ+RJR5qxW0CTcFpE03q3iWU4mOglotBF
FMfSilq98pKMAyXtK+m8Of+rIvLSnEt3rrNuz6KlA0Fw1K+yD1RSwnR0hRQ63tQV5xnt1s7+VJH8
ECgqff1p5bNrXUYOh+9UbDLuTJ/mCrfZZm3+68ygDvV5ShJljbOn2cMnfIbCenF2uZ3eyNwTp4K2
lX1gOQk3mqGdpnWqJ5Ami6gEVG2/M6Rp0d/9XIwxiKV/okNCEgAQuSWtyotDM4/kz2u2GIkrn4sj
j2tMR35AMBW4FMsBYpWU/xzkDDdZAA2K0v4F9cRPu/0DQpENwFc+xmoj1aMf3XB7ZRXaj17zkYYK
0Fn5KYQ2spTFb+08j21pV+7Y2/u3j6BqcaXz8bEM2UVuSEKSGWkQhakdoF1PlnSwn9ZG9d0wiKdy
pHwUAb2+ROUjU451iI0h1czRzRcVvHpS8PJAWqYTG4o4VBGkrbKtZsTwddFZmEnlcqVQYOiL9j0c
uXM7OZk6MxtZD8zT2Nbrprx2+CCwNwLPNUtbqNI20hkqK2kXMOCrHegOVEcLblB3RU09DNfjzFdA
vtn7/u/07Go80KvG/NkIG3P2a8tpwpwt4UsEiEBfgcqbOEz6Iorw+JfHZoqt04FMEln20xZfoRvB
WW5PHQsGSaIBaLGFyMLKAJ20X8hYqJ5+HIVET6HOH8uFir5IPrTTbqtXvdJI+CBBdWHg6KzLfA4h
ZO9u+M65SXXOIFR2Y25bmvpsGMXusFXlLS+wkZNvwYsPJEOBR1TEmQzIHvD8qufDIKgadd5qpyIL
EeVlInUu9mFv26jvlKbzpDhT2ALOw2RhECPQDs53fBBGZ/r5UuRfeeqk+mRPMvlNG1bOcr50HB9w
unzpV05dzwrZlQjfEjVfarPc6AVTeqazj9rdNYHVAgD1gi4EErDRbF2ImDFhioLCP+I960LjLzyU
2tjohZoidH42iY/GJXSqzMNoQCq0u4Ukq09Hukj9r5igCOLPb+uKus3P9O6qoJCltpWq+JGHSD18
+pTQb8IF9pANV2+cyBh0pQbsJogwGa0QpZkzPeY9xucmjVy8Ja6+oquqNngviFXZYOuhamZgAQ7y
6H528Zbo/fqCKHcFfyH6kqAUFTwp4OL4T5k4C6SHNGdIO/f4jx3eLF5dCjlzriTRdSvHBGaeGoPn
5iGSCOMkZqllvKAbp7UaAyrLbAHriwWm43l/B9Bh4/oR9dFphN3b4lRrg5Lrfk/Rpls67vUvCbi5
CVT4AitAwY8YTht/iC/GFzmvN0wOqrHbACcw99h5ylWDu/HoOL+i5eKCK9j7EcMZmmNc9SHn4sWK
Z5h7WzKo3vbxsCZJZf9z58gJuog1P6efNWqDDdvuCPX7RerGmgxDMbmT3DcXQkk9uWHLfMg1Tb6V
EG+U7q54VhH3LnaivGKaRmunFVmJO+BybhV4MSRfOigYJT4xyoGKkoILiVoxcjCI3MoohkdRzPKt
h45frBXgXdLR7m1wmb5ITtpcoO6zbPC1B5pfcHgHTvB9Xi8j35iIVHqFg03WnLrvjlO1wkSEVtUW
fn2PBA5GYEuCguijguHeq97PSoQSPnIZUnlXI9D8LI1l44GUpKpC1cUKTIOmxMerx+i7S/5sfGWs
M3tjqxqW1b20PuvCLGssb6oGou6+LfPNEzo4TteI1bzocxj4hmqX9KtPQv3vLVOoaTD2mfQ7iUqV
dK7YR/E6jotHv0m3waAo366sKA6FYm/ZClxbWtZ10nwTTBE+DZqYMNZI8ZpTufgeHqSGG5wUB1dc
98ncjZMlwM0p8f5wSkArp2SZhY+E3SPdMaxinNLHOttdRC845c86hSY+RMtpwcdPZliFk//OsSO4
xSDdh/f3N26cJGRjMxV+tm/lYI/Oh8H6k+SfzzfavRzxXuC/i/WUCU7XdMpofFRFgj0R8nePTXPp
LcQFeU+vLPoBqLat0bdoockhYnXsQXgnwCXGv5pBVG3NZG/XCGLM/Y6ljmvUcNDQDkFo4Mj4GbDp
Qu/POWCn8Q1xLTV3uTa9K1gjgZZTVCbhwoP0LIiVpO6Og+e80SibjXvss3U9qdWPvdtlxk2GSxi/
zdpMo1AYg+lBU6MGVC3Oo6A+4jI3y7jZhp3cQrnrq9DnNnYoZaRsCh7GCjaAJiWbzVNY96CpgciJ
5TyUMfsLnEgGaqwivXSGPS10qk1qiWzoQ84gylVaqKL/gIL18Uq0LDrKXia2QzmeGbTGPqrQ5ZWx
y/WnVyQe3LD24m8rD8PaChxYq2y43B3P7mTVfPViw0MJ+hWQAyiNyGN11lS3KcW/Y3ihJloVA5zH
SEe/QZTEeszvGwvxjfiyxogqNcgEXe2MDTI1VZnDdb1V5hAvTEws5EpRVm0zMIEZKdI9A6squxQb
hgkC9K4nIVmkNZRR1mauCA9b9Bv0wZ8dXRnUCdaPOMLYPFTwyV5Ma89C4Y3UZ60l+HrFP33bi0It
3ILMsI3y9QSA8dymhrHBjIjbPxX3A1fGDk5UADY4Aq76ougU8uRrQTqBr5VZZmslKcP4LdEAtoSK
sAp8hYba1s4Wbj8tUqnaE6yaXjs7uvXJB3xnO5SYOnPftM419EKWi/TSogJqzryZg9YW3o56K/Da
FrfS9EHLtTg7jRUaArAQl/iTehSYvgN48wre7IatTZ9ddAGH09jRWZQ/+lpf+n46CeZzdbwmRsJm
jQA17BOeshJz9z2wg2cjQnZZKCBFc4hLfimBxov4lTuzO97EpbOzOjLyDK514WV2If7Gu9duvA+M
OslsUNupzupYpLRkbUcu6nGcHVYsHlfYBIkHiQnRCQBqP14n69QOUR3v4cui/ojypGOF7ezkJwJq
nyi+pz6OGyLYffQRQjc+eQETo5+EtRsWB6Kf01fZelA+5QRi3o/u5fcimn0ryxf+I4sK1hfv4+3J
oUFsuQU9jHQ3ZoIQ8GKK7NymCFgLXc5Q8XIRuORn/edfcT0qU/12oE9Z3jpv6UPorwzQnwWKvYxo
y/y6NNp9ETDUMSJga1pLWo+RTcLIYAE8w7EnAJuqfYXnlZ0oxXUQXx1pmcg/kfCtJolmt55G+n04
Hx6866OxD8K+GGHdl+tyNRNbPm+CBe6sd/LzSniug3ZolUsK3nPbFmHm5L8UR40REpGbxxQOwBc3
S2tUOmRCKxXw7pMAHAjl2mHLBeCkpoUXgZBkGwWl5vA4xsm3xjRiaCJfQOqTfKvmT1uaf/7uuefJ
DSj1LnWO/4IYSSM2myQeKx6WwNBjt3c4xE7+tq81BYrdPuDSeP7MA9wuKqRF6pcBvCCb7wKXNqpk
C1XEQ3XtWf4omiPWOu7r4U0X+ZnprMYsc0lOLcM6jzRWO251VTV9V9p9uN7I960Uqvpcpg9j8Swb
4CHH5WLvVrZ/rIkZT9CxJftq2lAuHrJMDAC0HNykyCHQaanuoT9chq7BsGPpLtgBGk3L9v2kBZ9L
U1D50bNncx4UWs/hEYcTWP7H2D8UZ1gFfVdv0kwIU3JyZIulXBY+9aoWaxHoTT+iTtIU5erUNXfu
ci6/vn2qPQPpScXqUEwYHLCWNFa3Hf8S3Qi2b6oacPMeB+/85mHJH6rTFfNYzwJvuz+30nduikuj
mxmVGAyZ3EAQ5LkW8y8QUsRirioi2XZE8BWhDbrGZhneYhJMQ+YWub3nYPPvxHayEIkFB8mjOEXS
zAj8vDX/zv8fUdkHIMBV4Jm8O1A6PfErxvcBh6JaJhX5M93oRE76YQLAm9gQ+H07jbuJ1d5pj4qz
bgzMlAZMnf/gdIjOtNKj492X92wxQk80Xabjwao4XhX5PvPEOReJuJL4m+g2naTWUpJTKJbgbFpm
nXPuaqKYELwzTA7cAEy3iZPecAV8cCWBrJ7eDiizapHPfFbaTqOIjk2gFGaIvU5YLDRkxyH3M41J
/ztwr7F8opQyr5E/ylZNX8zQU0Pllqs7Df80bvs0sW8gG9M0OnEULXyxRZLkKqY5xFO+e/sOwL0g
8N5cN3Nbx34AEPrhu1QcBXVuydo7YAStBHJfCgNv0xwAOWxVGVK0DikEN3xUyRZ6hQw7gOEr905B
LTW4NrzKURkCo6QsKu4Hk/sONU1zYpNqNccZf3RjjJdunlGCODeiDUp5L4DOAl3MMa5IvDJoaTKf
D9aFcYI1jACFdJ2i6b5BXEYBECeI35dQ6hYWDMP98AYXwebiIVO+KjsiFYpUnywY13EspkFAe7i9
yoJgtYn7JhalXf5FlVscLWb7dzC4BRsGVAbQ4sl7EoQYLH4kYT6LaEM26jMZjJZ6ysjH/1YQR3yc
OcUI09E/6Ii/qD09kSGGtM8fN48IDS3ELzupIJB5Q2JqCdGsV+rV/5rj61o2BnZ9R8FJPnZrHKaW
1kmOT0/ZvmDXnkZiEyFPTKkqHj3aRdj6Wqg19v+b9tNm3zfh+zyp+CTsdhcavAwUBdnYcspB1Igb
SfWOeW7dXWsrrNhWGqAG+61/H/CsFN1fvfI23X5oUPnWutdG0+N46qCxdqgDaKanj3NCRtmdO7DS
3DdcOP+Lil/LbndhoASadkqIYCRjC2pKqM96GpnkbIlALx3EfqkBZwkQBc03DsOWglHN7bV+26Ex
X/MbZMHKo6b5gBIywfAXzwhloSWsHAYx2DrQEnOR2XTTFf4erZoDJiQTJ0QIr6lKrT002c4bW/ig
P6zl9/fz2xPY7Y4USE6CJp3AgRjVSVIQJEQNTyDB22jEpibdBo02E+MhqCTy7Gxb6d3y4n8wzjBw
zBsfHunmtgVrOsPdit9ENCjHLR8XY+3O1VKBPGdlgM7O/Xf/aQBI8si24ghIEYg3FJw/5KXQ8ba6
ApEc/ELqS7fKEHys/Pqtga+sbAnzsyWZBU0QRv52LT11WkwaUAb0CvISsnYd4QY37bpgD5CvwUzm
N59GbPET4Uq4hrHEsF4uXCSqyUEsmUVM9uczQ/xiv51ffqH9HOv1UGKRIUOfE8dX9b4NMswYOSah
TX8VvkZQ6RW1WcJITgLvsu3zHE4DwZoFDHZM2s5KflgbkWra/8+a7LVCcP+tohjsP8IC2Y/qJOqv
TjtgezyvIIotI1euq8JGYSlPA516yGs9tEmQP4jvY83Rav0fm0HKO0wgIJNevtEZZOygOtcBGT7r
Ra0VQEH8ErDOXPYBToCLpPh0xfomf3RqmiQg561V4iXmT2BMtbA9QgUhxB9TG0lNZYS31uuZJJ0n
xtDx+mpE5hGAehuRV0jrbLdjho5+9QhvQeAKGkqQFHSBi3+vO0Ar1PbXz/HUeI9jqatdFfG4hDZe
viqVeDsD5hoXEWwLt+g2ympAfy1tUNo5dOoYilKr2RkXQuOecZJqxW+70K3W4ATGFlPv82ZRsQ+p
Trbc9BL7q4ljnJv4/EQ48dco+dk0mBTUjsFFpch9BehsAGQMFsCtXVtBfUl4/kW/LuIq6SIkTFXt
HSGPaiPcx/HtQobMhoqu6vCveQyBbCxt7fEDg2W5zRMgoHSJb3+CodFxM1GGbrHpFPXajHxz7isw
FZML+132iJSTG8EC9Z+nTjW/Stiyl6v8klyHagmT1KLwCA8BZ7X6HlrPeGCpNysA2ewrqjVBZqF4
v7+IIo4dCgNFQN/Mxij8RX6F59W/BR1eS5P/Ye+948IoXXZL9kikiSoCieCDKkOJuFGLWNBs3PxK
Y4AV3vKwTiMRFAZVWe8+N4QamJXnFeJ2vokhVXol2p/uH7lR1Qkj6kOkrX7gYCy2ChAk4CLgYz8m
9/ks8yspM6eyylmyikFauGgG0SNGb6unhIlGjIHCNbDYLkbempmqmwljIVbXDk6Z5WkVHJJUz79N
M4+ZwySwfyD4rtudUm83On2f63lfaph+OBgu7BAoWGHfHHGmC7e2XJwubpcOwQulQqyMiVErEm2M
JqwFFF72KPt0pTlhWwx8kBgTwETmG+88GQ4WnPKPQtVyXPiN29fviNcMIO6YPE7DRT4+3Wz1yPPm
JUEDK3borQD9uFpuvtLx9ZAklIqaf34u/lTbIqzRKTSINcmJlAjLQBo7N5Qp4ZINJg2DW12JoLWk
cPzUpgq7NxELePdCM/M2nv6vSpkfwRdCbwI5JHWfyg9mY7FuahiPf/PLrmzXVBvF6D1Qc08zPREy
2lVFsVyHGXLhZYjyZ/0WMUPr34q+DqzAfiYSE1dMx6aZ4NqfPe3CujoPvx3BMLJhKqz54lcU5ROo
1L0OzO2l8HbMbwNcvET9N9w5XSBh1WDT2zJ2gTpfogH80QIWmz3DrDlx27VbqT/X84BvCw1rCk5p
wiDAB2SkfAtW3RYksKX0GiQ1iRXYg8IwhmWrUX00Ez0QdXOAW3RsLxtVQR5QIFIKN9YTzTrwn2La
RrwXVxy1d0K8e4MOVFBa783AX/HBKHPJJcCNRZwUdzPsDTqgRIKMT2GypMPHmAKWZslz1NGCH1Ok
FoiIUROsHnvvxwyzVOmyu9NI5Z0h/iPuFat6TJI7ZBzEsJqDT1ABxIhvma+IKS8uCa3xq2/PD7BC
U3p82519bdN5FrW+vySFSc7w18XvIWFZi5bd21QkAjcUX5en1EEvqL/XPf311glGVne8BOmaTmYk
fN47enynC26jKkD3XOcOMOmBIOEF+JxjdxOw4FD/LJoEVhiQTFs9B1FGYiD5SVtZZy6l7kygA1uv
/qYwhYtMejh3Cq7eJfufnOtyvQ/txj8CovKdAF0/dx4BD42W85rI2LnRAA0T8NbJI+N3dHvciJI3
/13ezf6Bu+Acvs+1tmZK3nIRlaph4Og/nE5N89Alboo9K2kHX+7Us2ufI/fssD/FMKkX9hSst/SL
rzf1jX2zU36h/CcitVSxWtYAzGC5OBnxE7BJLCULWAuf9UzispmJNWmBhc/Xn4IBKz9bF6n+4CdR
JYArN46qKhDOdd6Amb+rrlgUgv50k9I8CLKMPNO6KQFTji3KDrO2bdSDNariFf8daQN8bvv5xdc+
m3T7vJplBEhP4swiFEya65tLydMoS9l0UTRgQsX+XxjzCE00NHlSpmeiDRn6TQthOsRMI48H3Td9
aksrm7UXZ7YSI7NMDjoBWc6BsNjQmq6Ya+k4zYlAth57xjWOD86uTKfg4mSTJzFjz4lZ0NZK0+x3
S0gdsCxLxXP/cnB7mUagDOGmI0djd8mCd/7OJKW8Wuk3ICgjgnWYKmpZONuUYB4jW4RFEpDL0KH0
rBinEVRhdWDbTTu2KvCvYzzV/Q1HbWsSe+bM3JMD6ny1mw0U6ESWa6s9YPfFdsCzdKsJtZLtLnXY
N0J4qNacBjwxGA3PjVVQembayS/Tw8EHs6kdr+rHt4vxaZXpthr8ipLF5+RfAIQar4i2odNl+/tM
asUl2P36tuCVmKTgxgz1Be+azJxFjmoEfKaxOl6IdrncYrFwDTKYWyvQSWbv3jkyOHJoZGDKJxn8
Q4Uu2EW1kk444yf5nLo6LrlX86WNLPZw8WY03RLD9vThawAk4O34FLYJg+Ze75nlk1C31ZDqKABi
grRp7Ua/87VqPzXLVEynPlJYOBPYjHP9SABiY1hpbBuUAdHZDlEP3J9EeRUS4PN0YbDSJNeZBbe4
EOxmrvPoreIFrxtE56ZxKE91e11UIzdiOrIDaVgDpP1QDkKkh0d4Nr+Jvv++T3EvyCmjG681EfK2
M+abPaH7VYZKoA/qtjyy6kuNXlAaOz3FOVeVq1m7/IWmnEIamEDGu5WyYn6uKbFtzeOkBxv9VBR5
JTmkvdrmfnUSMhSql3OFYL5lIpGOzMohMiHwgHJTA8bNnQs2pjSHNypVZAYYtnrqSoC8jhD8G0FO
C8f201p1IteJ2xip1pU1tCoYfWo3ukRcM8ghlSWKlEqlLNz+Lq75xxrcl/xVDQPfpmh+Q+WWAtEU
6tyEMK9xoclOhjgm1+L372iavOMj/1Oc/LRkZ/sf8TZPeCLsSY0uoRU1MXGtlxjOmA2DuzMxJmM/
dz9kE8CjYybhZ8pSsjR3UB90OjTKTzgyMDEuiho918AJmaO+mVCTsMqTbB1pEWSwxrIPWEPEOp7O
HillroppFIC2B3UVpKSuD5Gqn9lkQdkqtnc+s2k5zb/ui5q1s+B2TvRUI5L2AVbmARjDvUg0UPTP
6gxagpkOqHPKE/EWbLQ5Jarpqp3o3Mh9a04cBX3mC8NV4q3croZTOq10tFgOMcHOPcRfVeL2vE2S
rhsDxNIz5kJ9rjsoxrS3l0L3i9h6ph6JwOPSV8d1ZjZCjtILhMbHR48K/1LvzYVRgli1wVIjheX4
S14+/DNN/snIXhO7VEMFO/AjLoepi5NUl/FPxkHsR3KNmYIXd5TVws6sReEhHn/FUL2sv64KScQW
hr0a8CSvsvg+66iU4WxbcuAXo6ceUeLU0GCeluISJoyTQ3XAswFpuEgrPX8YwnrprMvpb5BJTTfe
EnsrTHQBLv7C3Mi0aRiTSmc/whZP6DKAfxF9ce3d3y/lP+C7uNzicc4wnVqRMhlqsH+OgE+ghi2A
+Bx9cQ2pQrk8aUCIrS3/ySMDl6JXpSZShaZ9pXnWLrUEL15hUHTHjquxDVlqWeJp80tqDic4ZH2x
uu75jd1WZw6pjDWmVVp/AXhRUFUvFiBWKMNf26UKsaMiXNTetNLR04FkAvj5m21tZfbU9fa84wjy
3UWv46nr8XUIQxERXtaz2limgaIYAwmm8zg8j2692AdvnyEG+rCi/HKiaEGUp+3muXaF+UuQyIwl
ISOwTYGYCbUuZIqXGN/FopOzg9C4jq9DobHZ3lar6Wd2ADOBPUjYjJrlilyJyI5JWcJwYWbjHI8K
G1GOcu22XoVBnoXw1efBnJiYhlSu4HJ0ggnJCs3P6Css9paJvnei6bsttRevZbRmTPL5oJXAJQ6/
HIE69LZ1G7rt/QJJ2z/weRorsQHXsiiuM2rxsWc7kAkghImmng7fWE2kIdDPXwKHO2j6Fxnoe+ey
OkgPfE3wyEg1Gm1Kqh1aED5Zeo6D7ig14BRa20qhBY7xwII/+sxDJWm0Hf4HRLfgrH5jZOh6AC9y
M8l/p+qnZNHIxfZugjr2RJycjHRExPDi41op7nW01psNOmp9KOy2A9Xy0BUo/F3h1nqjVhEtznrG
dUb544MoTuAZBLBRr1G/e+8XOrhF8+GwOM/2klvb8xwdC3+W/gxA6COeQYb1fDhFFQwg6qXVCEvc
Pxl/mHuj+LaD+stGFqqZqQGNEaig89KY5qzFkwzfIPepvJ6udk/uFZ/imn12bScg0Ki59RHO3zZC
qRQspAnXBviBZWK4FUtmviz7KvWGnMqpqUpykuRGpEVra/AP5oUE7zBsp8VzN3Aao9/qlI1JkjPU
hPsqc98le6eSLAGisfqtBObG5YdlcMU5hYybvwaRi93RjdHa6et3Rc25Ya/vpbWh3PrbT9NJgYA2
WhntTK1jlD1EJ8msGM4g5LqXZCp0t6O7AZ3Xz1amWkT1YdGzYKF9mlVTstupsxRVKb+6lHwpLm5f
u1d68/nO0XdVQC0jCpnKabMd/hb6eUpon5XWOZwm6duM1sefzedU+BWiOFpzZcuiZX1DhFY3QinW
bjz+fM7flj1ZKxZpoajm1iwfpUP8RwJixwDB3nEP2aHO+lxRgxnhUPFfOFhmCd5oIVkJtV0lCKR+
yiQxVr7XwxJPx9QWfVGY2/n+5Uzowxs52wlNRiGfrktp3iQGClNLe4ZJteY8hTZced6Uiy9cINaG
KiHgctR6Al/iuiU0rJL+rcLC9TIFh+z34tKHeUBJJi5/YW0/PTmu7ENznXyIUfGDsCKXjt+I/VBv
k0uooAE8+SN0UAlyrXC90cfZhuqL7Us+eOWIqv2LDVemDGAnwHxY0ZUQiXsfaMCzwGIcLqTZSR2S
XMaN2Vy2cUXZK7QOfT+uO51iU2iL41IRuyEQvt1X7fSnA7Q66MO8+S8agvMctQm94ES4B20kHWqo
08GIyU9XwY2gnhgMN6w3mK+YGaiJK64uQYnb+6SpLCPsnBYn0luvnCbpkIFzTfGPqN682whRylb+
8sdfRnMoTxf5WbBRBnUP2X+aCZJCniY1lk4pq9TA8oOMp+7VcH8Olsx6BxDXWhiJDJqVHRa0THP6
OuEe/ZH+s0ru3A+4MNBMjkBeV/xtFUOpik6axzXbX2sbfl8P7p/kcs1Z1Ii6iKscP/Cb8Pz7J/4/
t17KtMOT6/Er1SmFFJY4X+vZnwjo3I4dU6TZhBMva8PimGw/w0fHDMqlz8P9vBVwSTydq+U2thVf
bXPnpoh7wZQFNqbN5wKdrsEUz5olBzsQWnAvda92TO8gukWkEQrOxuDDKveLcLFvQVyQ688M76Cb
MLQ/KIjsxkzuKG7HOsHGblUMec3q6F+NNVtfDtHZJgxq+7lwsxzIPhMLeeoZJULbZuKuzPQrgCIk
Hn9hFX7xopL44aTYKf9cu88pVuCRbUy0NAHFZFsXeEZgGKshVcEHkPnxPPjc6UGMKzC6pysvN/a7
zIW7Axmjr4sTgXyderm1k3CoJhb6Rhz6neRQW18gKVfPYRuT6z9BPdqatMPYMv1KvrWaDqvmr5XR
jrA+TsVroYJJTAepEFh83zfI0QluQAilTstc/SiwBXL30zLRTR5k6f2mexd1rUexazbqS404iZcR
3mLdI83/1/pgVhx6dizF8QC+e6Vp7mDQOmciLLl14weSV1atb/aywoc5XgbhbUz9tWrqIrq31gne
5Fp08H+ceIADemjaOAHulXH3cQN5PuUV9Q8tjxoEjW06P+Sqvbvn0NoKuReWz/aD7ZzVm7gogf21
lfM/PKIvanL6GfGqZejERbgCjLxTCOK6Vr19Tg8PQvPBKPGVOCjdCe8cnc+nf5LXQsWdvaTlJ5fW
dmApfH3ptTLLsiEgCC54KiuThDf8MTMt/aPj/MMj1U/N2269mtORhBk03Nc2ETFiENMY
`protect end_protected
