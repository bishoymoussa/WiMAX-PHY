��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$Rx�y�<��wA�*;�x���@�̦�W�X�fa�M-$u����n~�%���P�$��W��kYَ���P7�?UMfT��q�6�U��k�>����~�\N�(�����X�e���/6U|)�X2pF�]$h���d.���9E�	�IN�f"�\��e�z�y�b�����Oo2�?�qˁ'�͜k-�K�P|����y:����3�l�d���bl��ˢ_�d���kx�rq�mh�MذM�`aS�.�DW�mS�9���Y��+�>��!��!�T�uOB���,��\L�7m�O��W���6����'���j)n_�I����2:��$�K�2�Sʫ��l ��!���{�l����.�j4�	��很�̢=�����N��s���s5���_�R�>����ТP .W;������	�"�מԫ�����]�#7@O+?�⡾�Ԫ���e�O�\A�	�ͼ���ƹ�d�	@�nQ˰��E؁Bf���|D_�%au�-�'���w�*%��"AM$w�*4���J*!���mj���U֌j%�A���m$�UL�k����s��}�0��Z�	���Hx�@�C<�k6>�7a+��&�aS�Z�Xx�n�$�eh4֘�C� ^���z��!��Fve�wZ��G��}�dDcr	rJ]4���@��Oa9yH���>���o,�6�A��xu��^��<��*�}���J�o��%�� ���	?s���Y�C��^�:ZG��X�>5;m��������Q|�İ��Q!���v޹(��)P*9��e��TR�biz^�>���Os��?���|ݲ�!��ق,m�Oy끋?Z��˦���,[Ҁ'J�W�����W�	�G(x%��:��ɇ�,���a-����#��m�g�8�ff!M+��Nq��7�<�b�l��0�Bј��r�I����?�~ALr������C)���n��W���g���U~"��^p
���o���u�.|�ƹ�J̤t�(U�K�V٬I��o2
�M��.��k�L�$������gb�e��ޝ�#��3/]�8oD�$�|uzmw����y�b�_��!P��tW�Kn���ݸ@��� �hj|�w�J��7n�l`4��X�>;��S���^�yeCC`/pI�}�#.�$`W���A�4�TF)�ɨ��I�1
��`��K���7(�+( `@v=��B�Js���~y9�KB�e��p�`޳uaxA@�|}� |#�?G>T��a-�T�X)�}#j�.K��0r{iW��ؓ��6��Pj'��g���N�-цg�#}����t�*
n�e��I�qXx�cϗh�O4�t��)����o���5	�[���w�L�R(M~��t(�k����VR����L&�$W���D]�d��B��4�;>�8<�m#�(�����ٷ�W��\Ԏ9F	�b<�f�+#�@�Rƺ��HϹ�7�O-��4��EM{���"��ʉ\�����0{d�
Y�Кg����k� 9I���bg��CR�E~��`+��V]����O�ua44� Do'���`��^tpA�� "ԀiU�c�\�.��؞0k!���,F���3����w8
�{�sag@(��k��cf����h'b�O��Ln��6�O��,5��ڳ
W�
�5A�9��4�<fwޢ�դy�ۧDfW�A�T�9W�<�5�^$�k'7U����+-��Թ�R�:�Yj0#�$v4�\�2��[X?
�T6��WV�ɟ�N��ˉ�b狆���o�=�j��P0n7z�%���m~#q\K���tAifʜ��@�:�vEn�@b��]^Z��_Ȏ�
�-{�����D
C]p�{�:�X�a��h���H-��dnV&�UPt����%�/�b.X H��ba4BHu�pA4���|�\mH���q���'E<noV�B����R �{y�9ʱ~��]a�]Lr��L9	���� �hܩ��(���(v���'	|E�)"��C�w��Hkҗq��%T9�|�=�K��@����wϸ��3��֟Ol�҃tH5%�Ҷ %/�=+�E�]���f�J$H�����ޅ��*�Nt�m���]3-�?w�F/�o3),O\^�[S�̒"�Q���58���;4�$FV���=���lAU�Μ�{#��R�� �~ �f�źy{�=�t�D� ��l��GD���s� *��0G�j� B�3�ޥ ��N/�l�϶�V�xta�7t�y�4d;,pvv ��EC�mup1z�S�*v\����;Bx�����rw���b��7:���c]�t-��T�p DQ2jQRK<��Rq��!����h0�Ƶʙ��56��kY�݆���J2�~y����o$���}M�z'�p�������u�)(��K��M]Vv�gy��xs *��x���E���?�p�۸�h�����B�&���/�S1ᣌ�0��=ŇH�Ρ��N���ŏ39����Ḯwx���FW�+�����[�h��&��td�l�0�	��!ˀ�~�b��[�c�v#Y��\�4���b&�Nc�?�um<�{x����\	��S��+R��/���R/k���Jo������J$kP�SX�s�1C>2?0����:�X40���梌eh�] ��, -v�ܙ�b�5�ӷY`�!���r�U�C��h̻��zZj�(���MFW��m#|���8�fP���Mr��~�2��\��K�����V=�c�$蛾W�+��������-��vRͿ��ˉ�􎸟�`e���\o1t���� jal�A��ٻ'���ՊΓwJS��UVzJ$����DWn��Dm����K�i�q�T�ݲ|iZqY@��f�%�V��O��/Ň	{�1ªh���糆l��\)��|&����:�HP�Ў��v���C����cHƤ��BCn(�D�"͕�E��6���@Ub���K�Pݜ�r���Y�"��rT�y0|��A���{�c	���o�)�Q���am��6�D��f@q����5o�/FB��y�i6�g� ���A�E5�'�`I������[s�A3��mY_�z׌�,%�Ii��5��2�C@r2�yk�';\�h���J������9�̑�!�J��e�#Ml`N��U�.�*��L�*�+��.J1�L��3%�S�Hߠ���J�$�c>gA��~/�{�A�&�mv�E"�.�b���4�/i��cƸ?sU�X.]���L���bH�hi����a�Q�m�\IF	��B���ppWG��D�z������v���:B��;n!+�q͚-�����	Yq__c=�j��@�Aqq������Hg=�8灯ć@h�#o�(^Dm�i��~B���z2%ɤ�%$S%C����vړy�������H���H�עmVh��2�7��8'��\���9�j��v�H��<8�V�h8��9p��U�=�g� I�(�B�P�!��|�ȘLOm��}S�'������p�&����J�O5�<�X�<O;O?Z������-��5~���9'�^5D�f�-�!��va���BW�t� ���LC ���5t�.���(�"QԺp�w ��lYmL ���ˈZ���͸i�]�a�qTs�Z�To�*z��w��pU���g�;Pv	�0�Q4.k�i�z
��57O77�~��E���9,��wK���J���֛�גph��v��F葻��ٌQ�2�ƴB��N�f\	W�pk���;�z�t��~�)Ԧ �����o�zP< ��ᇻ~���0��4��`"|v��=��;��y��ݏ�bñn�es�:^�ø��p��ҫ+a7$���&�4���F}#����砕h����)�C�a����Y�Q_�\�[.��9�t��m8�}r�\�����ht��[�e�tw�[�R�0�}D�ʇ�yD�*��%j;��P�$����IjU�ߎ����jy���B���~�E��C�A'�w�[13��ԥ�u&��c/�9������C�|u�ۯ��S\�ʈn����H��	K��<���j��E�%&��ڼ��\˺@O �e+���F;g	�\Ę� ���4��+�,6��I�޼��}\ȉ�ݫ�	��b䯦������%��vΖ�I�yPH��:A>�<V���|�:֑t��E���5�{��}���'����õf�x-ߺ�p�6r'v�JP��ճ��^�s�n�",�n��V��%�S��2�p ¨N0�?���&aj��y�_EV�j07�h�{��EVW\��վ�E�@ �d�r;�=d<=5���j3���"�=Z��'��u|{[uƋ��U��LB��^��$x�N�� pI0�����[�����̳|ɵn˕��>�n_��֕u�m��P7�o!m	�wa���h�@̺�aC&��ӻzƅDp*k��۾���:~�z '�?U)\(1�7/У�-q`P^�$�O���f$����d��TFw�̥��܊�Ņ�ٹ|[#-�#-�%���( M��m�����}�ʝH�񡤫������l�T��}�
��B��ӏ�2p�M,,�W���0C���v��V	�<���]�IF�F%�4��yZ�B�TnZQfM�����W�+�M����O�ۤm��4d$N�j�̒ �����s_��q�x��j����f��W=�'=^�U�P�:�ow�l�#�r���/��F�Y�(ة����5�|��n(���Q�W���Bt��ƚ��*�̯swD�h������`�B��b��Z���J��HXx�,�I�>Ƭ�c����0�o����8C��]�j%����EwP�'߯���b�_��V2&�`vK3�g�e�a"��3��,�|�i��m�;��s��DuWId��Y����x����oa���*tZb�Z|V6��1Z�����Yyp���%�]���_)���6俎5�f.����+�sRȐ^��J@��s�bx���v���J+��#���,%^�A����K�v���#zD��lc"ć<��p�?�Ҍ:�3}d�w�?�k��W+'G>����}���v3{�y35�"�^���h�=�=��#��<}�,$�S�Y���"X�E��C��z?
� ��#T�M�������؝���u�őx���(jQ�����D�y��e�.�>���[���wvD@6���
��8��]���>a��e��v�ֶ�M9��Q8g[�_��C��K3���r���&����#��\lT|m9���}��,���zj��p'�����:��&�@���s�^T�P(����T���
|3zltc��}� �X8���|��<l��2���E��f��z}�?�W5wl��z�0�m�l�\�S���G�[�p�ka��@���l�H�a��֔�p
�x�WU���p��qb9',��f��+]��ιDKJ|R���;�*��8Pf?A%�����B�?������#�w{����2:���.}qBi���h'����S;z2�ƀ�5wȖ&��[=:.֠@&��?��g���i'��4����ǉ��)M�����U�����K�x���ob�D���1�����r�����g�ͻXB���F�4����(Q^�����xRr����*�������ȠꚐ��������9�B	���	�.ƪ-�9~V�C7lJ�]q��[�iA���]wٜ�s�"���7��.cPr5o�v4E(�\�Bo�(�iD�w*f�����Ͽh�%e&ٞ�T� ��j<ɸF�%����t+/u(�>[*Dbh�C�8�H�JH+��?,�
-�wAiB�wW�Ou_�2I��V��Su�W�	 =ZaQ�d	h":�\$�97����x#y��3��S,	�A�^	�'5��K,v'ܲ�[02k�6Z�2�e$~z�]ݰ�i�v>�MFW������^s:�?��)W��V�ڼ�Z�'��Y�ui��|���XT��$e��9��N��p+=�Z�/<�ݔܺ5O���71�#�y�Q���|��xF>�h�!Ru��̄��i�_pλ�n�h���T%;*�dݙ_s���d(�ap�!^�L#�'��|=ჴs��C��C����:;
�n [HW(z��o�j+�wY��M����Z�	%?'\йܡ-V�̱fٯ�����|/��*m|W�׏e�'͹��l�c���;����1����@��~tџ�r��-k�߸�n��s�R�@�0�Kɬ��Q�S+E��
c�P����h��(����b8l)��(M�=���8:��ہ� ��%��qQ�\`��|"%ngԪ ��D~[�,l�rQ]8���q��Q�׷��p�7ʽ�]��d����l����7�e�fQ2�$�j!`ʗ�M44=p��k�4N��8��M�*���U����nz��<�`����Q/�k��MmC+6*:��Z��Ȱ���$�+��~�7ήy�(�c�5���͝"����y����Pd~q|��H��0f��M���;KX[l&aW�2��EIk0��멀H μYVL�1��Lg����r���w�FT2iU���_�%;p��6w�
���~;�L����L3��؀�e�%m�����wz�C�H���/��5����Ե�+��/ۇ���ly�>�0a�jsu5F+�R`�[�0O_ND��M9���~Bx1Vr�m����i���[����p�'d��Ϸ2�zH��* ���AW;�.s
f�����y��<��᜸� �ɴ��o�m��GM/���s����;k!=H[w��ݺr{��Tu}�8� H�(���ͦyAa�r�D펖��DO�}����>&��Z㙜�����ά�4����Z��f�6����jGoЁY�^jn� )�nŎ9C� ^0Q�=R��g��J�ؗ���C�S����,�a�!=4������w�&���]���p���3����^Nf�\�".
?~�����\7�?����b�CI8�g h�A�� F▗��щt���'͋aG���˃���N�d�P��mu�;�6OA��Q�%��`��;Y���~*�/�ݱ�bp_���AhI]hKEm�s%��smbd��nE ���3�Xfb\0)��e��Uh���[r$y�F�y�\�STͣ��ׇ%�����X���ۚ}��A�C��ѳ�3���r���+��}��`���y�5O/�"��I� 0Z�u��v�UV�؜+�y.�0z�G�W\��*�L�ľW�-�z�$<n���daz�&h���b���CV5�����xNh��[)J��0�q�'�s�1D}�?[���dg�����XC�rb��v�xEtk���?��)))� A�B��xVZ��	��;��܇�8*{$���*?�bn�͐���ګ����D6�lFF56��Yl7��L��_@~�7*f����{��E�ѣx�t����l�-��:��6ZQ�/|��"����ue��dւ75x�X��cy�VJ���	�p]�k��$�kW�3�[X@]�3�{{aC��8vA��� �	L�^�!�N(�y*/�S��GC
��?�������k����%������c��p;S��)f;A����d��6� ��T���S�<��X^�U�m�7CFv�y<���>j�T&���t-���>��j+������e��g(ȕT�X�|�-#a[&�Vm��#À������q�/TN�T�� �����.mj���,��X��a�v�(�-�N�M�����s��.�0ZH;�å9T��e�oMx�Nhc�ȯ)Äq���v�5����W�Ъ:Uv��	9���&6AJfL�u�+� sl�� �����	�k�T~.��M4X��Gov�o挝f�ǤYF�ק��>!�Xm^h���3J.٢�VQDȇ(t�zV�~q޲����J�?ć���"���K&v]���ޔe�m.�S��3Si�Ǝ��%<w4w���]�VM��1��_*q�{�4R2�^]}$j]�{!z纁������5{<B��*�7M�PR��1]'�I��	�&����:�/r��
�Ȇ�����剄UO�uN�%>;6M�>T^`���b�q�AT������3����87��ڿ�r0c}z+k�$ޮ�Q�Fx��r�0��s�T��CI��t�������sjx��V"SĖ���.��Rf_��FHyK4�tq�.�	.���S}��6����cz|*G<o {����\D,~2���֗$a9/��M�+`�����K8�Z��tqV �L������U��|=U6��%����h�ܣ
��W�3> ��C����9��p�`GOE^ς����n[�2:�C�,��9��HQUo��Q��[���'��@�*]aP���_z��.�H�Ձݬg��Ui�s���e���jY<����t�i^����@�f%��8JQGJ��e-7_��M-�Do��]�Ƿ��6�D��(L���
������ݵw�1�2�g�%�����<�:3m��E����$�Vwi*r��C�-]����9E�� �� �ꃘ �!�����������^�Kɿ����ڲL`}�9�$��'��u _Ё��B���ۅy?������ɍ�tr��C���stEN�
kL��<p�fn7M�V?<a;nXz\�������Ok�����"�;�ո���6� �ZY
�&�M�q��O&����j��?&7s�U�:8
a�����<P�h��
�ĺo����� 'c%
܇.kY�n�G�n'�������(�j'�;�������Ҙog��).g�B��M;� 1Z���%��,mw���b��,���$�H\��kE�WH-�����J��F{���w��,��Z��g��M�y=�>�l�<�V��y�U}C�@j$hI�1��J�t�ް�(~`=���~ �F�BB�ݝ��R!jW�{��>�ź�{�
I���x`Un�nA�L��E�A�WԵ7oo6"�1��u᦮�f
6���jv��w�����z�M
�����=��a�Og������)�eO�8xN�f�f�o��*il��$��������4"M�`��Q�x�'�iR�@s0������/�5+⼻q<��S��p����8�Kn������sT$��~��g����p��8@�Pﾛ,��:?��Ʃ�˦Xjkȵ�&h��m+Z�+(��j��gd�l��d~#}ﬧ��k!��g`=ձyA�0�d�Ө�j?���}��[�|��4~����s������.�cm�N��M�ᓻ���JSė��]腕���*_��.��;��_�	iN��k0�������ƕ����X��%<y�)m"��ܣΎ��ӑ��OjPm�{x"�y���Z���}9H�Â�.�k�" Xl��h��$k�#韓�^F����#������\K7@,�-d4
�|s����3��h0�Ne�<��k�P�������C����'Nh�ߞ;,���o�1p'w�M=��b�����d��^}�9*�?��@�9E~�e:�X��`v���=���8Z�(ŨS��ffЛ����V0:��<6/n�L,��T`ߩx-��y�Ni�&ae�����	�~��sܥ$Zʍ�c�d>ȏ� i��<���e!���	'��f8���*�$��X  (6{`xʿ��4J��,7E���\�9�sL�x��k�HR��>��v�����G��3����N�
-��o�/|����I�H]#�p���M��@g�:YK��/��X�yEh���iT葝�n9����΍Z#1Y�#�o�P�-"n�*��ÜJ�Z]���óV�$��
�7:���s�LqX^;�{�]W��p8>LppX<�Ȫ��x��d�}+�@j��FyFמB��"N)�1�/�E62��^B�g4d�$������4l[���b�d�=�T)D�ơ��dj��?�r3��}&�v��S,H�[�����=�e1r��Tt��������u_��Y�!�-�S�\.���*2����p� M�&��~�G�R�g�^�����r�b	�#t���C��/8��Dɔ��܆823�g`���T�C$��P��,o��aͰ��L�߬33f�-8ݨ1�����SS�����B"�/x#����"/k�o��m%<��Y�G�<m7�dP=0`�wŅ��yíl�Á��� ���R��!kE�9/� %��yt�g��?88�*+����ݍ>屿�Zp����Ԯ@�.�p6�n�O��(=��^*��&bB�F���L�����/���K���L�)��4!��aQ�� ��fv(��-�LM*s�հ �FW�q��/3�I���aI�;�ƌ�aᵠ�6���W��jQZ����nP@�P>Y�TI]�C2�7����0��*�%K!�`=A�ᗧ��[2��ܳL�}[���q�3���	�aK�1�2��� `e�n�}E��^��K�)�O��V+~�
���sU�A����O�z��=��t�P��,׶M��� R�ͪ�]�Ic�h|�5�%?:�K������D���9��y�В�� %��~�o�Pvn�Y�x��F�fB� f�^+�,��յ%*�	 ��rl�:���M'�\�$=�����I�/�ds��UF�I��=��VQ���]m�ԯ΃��
1Ѽ�-S�,�azn�9J�M�c|�9���+.X�������X�<N9/��v���i��~�=%��x�D�iJ�:�O|�5u��34 L�ыgp9�{_�������F}��X�U�)rK���z�Q�S+rP�FA `i��s�p1�p]�ҵq-���ke&O�1��ϖ&u��J����TЙ��8P!��D��u�L$y���6����+24���gW�{�DBr)����m��p��y��yU]z�0��m�^,��X��t�د���V�p�#L;�޼r��_δvp�Ԯ���5t�Ѓ��$�g��b&]TV����=&d�{L^T��9�.a�Պ���;������rw���3v�A���ۿ�٫��B���N^$K#&��06d��v�����gA���P��u��#�Ⱥ&6:Q'ʩ��2��ޛ �F��矐�{3Q�n�� �H�ElƼ���W4t(���z��h�X���+AeN�ϡ�t��9��t�S3����W��?�BCX����L�(4���-�xm�E�?�G����2q�8�!@'k_�J��t=h���� �+���0����u����H4Jss��m�����]�#@,,�b�P��~�D�3�r;�	g�O��O��v�U"U����$e^�C`���DP����X�A�|�H�/(���S��q @���iy�xu17�|��B"H�WJr�1�흑fY�F�î�_��+_~,�������� M/K��_9ƿ���#]�k*��N�����1����,��A��eG�/�^��e�,�-P��|�ΧG�A�X�i� �� ���k�W�k����Ɛ�<����\��"����R�o�D@u�vp���e,�?���a%¯�?��;5P��"e��1���8O�����L+ҏK��n1�_TlcY+0�z�K�^��)>����t�8�xK�����!��U�(,)	��χ�x�IJJ�<���]�6/~``�!Z ��L���U��ɥ#�f���Z<�_�(k-| �v*����&����~�|�?�,8�czz�|-�j����r�?0�����U^�|f$Ȣ ����{B�}��\��Ku�I�� fß�J-i�R"*R�TM�<�M���܈���(]f�<֡qc�Up���`<yהK���tX7�LX��[!��}MZ�U=|A��M�#w4�$Y�5%�8��H�o]]� .˪ݞ&����8��&?w����v�6��L��N~�|�ы�d���;9���W��g3:�{���8�D�9���0_��i�X���
j��0#���O�s��	��r�D�1b��
>�e��ܿ�������+��U~�n�g�s��K!��t�dj_/���D�J�Sҩ��Bt�E.�G��zbc���3?�'M�h�Ҟ!���v���Q��Kv��R�����lN��ÍH"2�ܕqR2fE�T�c@Ex�[&��L���YL�ⵡ�����0�f,@��d5��9��G%��EXg�g>�{�9׃� 閿OB�+S�5=M�p�`��[��8��Es��6���D��!2���~Н��/[h�W �JyC�"z�����`�%^�6�x��������bVj���C"���XU����oy�oN%���G��;n�ZbN�Dp1j������q�/�a`p�Gf(�������������ͳ�cř]���TP�׌{�*s4�CI&w�X�N��������z+����>@	������5Z�[Y�9&j˞M�5�y����x!T�>.���P� ���?�d��(�
�T�B�jX�{xYJβq�8]���r��H5�q����+�m���� �å�HP;�AL���ׯX�$������q���"�f�0�F���+Ha�izj�֭��%�����0���!M.2;2[�\�Z�2Hu�RCq-�A�XQuFo ���5pg��`	rf�	Ȑ���>����O�&)����b�O��f�e�}� 
��ԙ\ y	�wߊeB��#ݧX1~Ǯ���H�O�����(�6���%���H����Ķbn�1|�5#K��d�j�uܪ��{<�QВ��%ȖS-�e������2�2�C� X�̭�g�
W�y1jdgg�E���z�e�7Ҁ��-�#�^B���-�}�nT���6I�3ܓ�ȸ��Okኺ������#7i]����4��*8�麥�#)�K��0�X2�鲧V��j��J�ԵK�#�1�/#��]P3@fn
�"*�cĩ%��n�{C�}?"��=��#��J�M�T�s����X�'��*�ջ��	�U�O�o�����1����HipQ�&tJ������� 4n���[��Z���t�H�yT+��o���m�G�B�XR<	�3I9�m���cn�_Ƒɑ��	�򎰛�4N�<`��7��Z�lŇv��LƆ��j{��і���f[%wNm�r�>�<��U����Fi]���\ĳ��"G��4Aϩ%����l�h�!`�w�Ů����A�M�����ߩ�dU�HKW�����p�q���~��������:�v���.e���҂�D���o�H�7U�QWA�c���Kh�O�Z�M1�t5����ݳ���`��r?^0qXb����xuO.����f�K7�o$���y9�\��Z���׃^����J���P�s.�݅6�ï���7�).Ѐ��P�H��̿K�+~4�� ]ʗ��`�R�(���+����= �q�>����SFy��~�Fk?��寍��,[>Gv\j��d�����e%@g��n�1Nz ���Vh��u �Pm�)7U�>�� ��׀�\B��������Q%%��S�aԽ�T�D�L�%e���й�^~3G2܈h/y�T�w��P������̢iEm̺Pun����}�<7�si��&/�Ġ\���^7�@XFF��[-�5i����Φ���X=��;�HBZT�z�bO�Eif�˯�ְu!����y��B�.o���g섯��c	�>Q���k�1�ֈ���T���:��Y�g���j���4��3���^UU�4MjǕ� ��<��<��<oP>FI�,;i|<���w�޼2�u+_�����#Z�/(��`҉H[.,�_'\{�{ �="���aS`�@��mFr�����ԥ�<> _Ds|7��u"E�/�����Тh3� �E����cD1����v%��1�1�c�W��b�,H�C/�����_��x�@�|BkM��aK�ȓ�|�?(a�#�H�?;P�ŝVpq��?G�G��^h%q�>ՋP�M�-�v�.�e?���P���w=:��!�ov���%�ґ�+�V7b��̕c����ZX8���%,�#y�g
_{�#4f� ��,��0�ёP*�;I�����"y��&���Jʸ�P�*���d#�5w���V�3�+_���}~�ή=����a�Hx���j3Sm��Z?'�3�����9��h�Lƴ��U$��B��E�gq���|;$j����?#�F�=�!	�S7�s�`�y#zx%��' 	X7��_�۠A�����[�Q�\c���pA���<���j���a�����v��2�ZM�:�?'B��Q%x�k�$���|����Nv�Z�B*��8��a�F��"����d�|��7)�&��s��&<��l�QL��o����"�ր̑Պ|J�?�(B׶1�z9,��yN�;OƎ��h"5R��:��ת�֛�1w�;�OX��Ue�/��� q�t�7
{�8��Wx/�GwƘ� |"�;��`������L�Z��w���n�L}z�Ȯ�j��h1|u��("-|H:iJ0l;}�X|����MO�x��)���u�����.���)(�M���}ENdF�τ��ĕg��L��T��~�IC����4�����6�7�;�/c��f�c4lTF1����\tV&1`$�6��r�]X?��l������Cǽ��=��e������\���9?q�U�^��D��_���n#��na� xhfv��v?�	�,��A�օ.�	�3��@
ęWj�>��r�__D����	-Rx5��nG��ؙ�@(�N� �9������sVD��c ���9����a��ؖ2^ 3��7I�j }�۹Jra3ϗ���F��:s�S�z�=O�҄z����i۬�R��g�C4��[|�z~]�pm؋]jA�>=E�h��c�+�p���;��֟��M�6���9�Ò��a:�w�m���^��c^�M!�W9®d���@dp,<�[�K�JĲ#g�24�Q�zg�v3���a�SXA�?�G4�"��ՖWzHP�呤ul���K4��(iԇ�B��I޴����fKig���0��8��nȓ�"����!��h(A�E��ؘ�B�/����T��F,�C���Y�m�/�Ag3�w����38�sJ���k-�k'T�g#Gw�"�'�w��	�U�i,�&�sC��6��δ��̩O�H���z������+AU��ҩf��h�����~4K���p���6���6�K������zu�A&�'"�b��02Z��p�a!K�f�w2��>n����
���p�$GU���&��=��j��?���_秔�?~d���i�i��:�e9����u���n�I�∔)����q��u�H��*u��c��C����/�&p�ŻD*7�:�M�ń���C��"����1��_^�a��֌i���r[�Kr��H�6�x�.Kv���ˠX���hv�����r�+tw^�|2X�����%�kZ��QC��L/�	a�:�T{K���]^�,���˘-��ݸY-����'�Y���?hR<F��z�����떸)�%"�;T��/0�I�1SA8�<䛳#J��Aw&l[)�����hczE�
�����yr�K�P�oa�+@Ҟ��?�^�?�h���k�����R����k�b��`�x��!�b��,5_�#��ө:<����2� ��ƶ#a����"E��?��(�@n��� ��\WIMU��?�:�w�7�j�_�8��|�Q�ݙ ���,q�)F0C٩��6�EN���0��z�P�JD�찋�b�ź�oW>������T��&ߵ��n`n&��.�z;�� �+�㑏�x{��L8�Ur�/ �С�~St&[YWc�9}q�:82�''A���,�GϳETo|V�� :�a9v��?��d�'R�� �a�S�'��Z5�����t}>=�	~��ǔ\��N��N�<�3�AW�k�[!:�Tz�����u��|������p���
�~�ʯ�#���&��$��j�r���(!�4C�a3v�*��V���Q@e�.C�3�O0jN���O�n��Ldwׁ�É~��]46^�:�:?��:o�޽�O����;&^��M���U0� ti�_k�(n����T.B�&
=V�[�
���~g�5����(d[�]�?����ߙ�K��e��[��ݜ�x���$���R�ī�Ӎ���Yf��}%�X�M��B�XK����̣'�P����|����.��OH$\��'�N�MZ� 1/V>�e,�1s�&��83�z�;�O���m��ᨺ��`���U���%�� ����FXS��O���T��.�d����h�e������͗�N��<����P|U�b�N@���a�:)�m�ەð�i���:�#�أ%8 ���H�X��Uk�����!c06.����{��|�O��?�ȴ�٬�;ז�� ���KH_�t�Z�
���^��6��ꢽ��R6�au.�O4����;��f��X��{���ѦG#V�(��ϱ��hO�[��*��g����K�5Rl70�8�ӕ�"_?{��A�d;�=�=��T��v<����<�7_��.����ft����>ِQs�>p�0�b�w}�<\��5mO� Soos�py�V|��r�f���fHh��n��_<kQ�V�a��OM:�
q*�:�����HFHN��zu��\sw��}-�8uA9��{:ڮ\ �7��<i��Zz黎}M5�P,�n�!�a+�]�6l�JA���S�q4�qj�2�h鍁���L�r:ch Zv}��eDsC��2��:������2L�Λ����C�ǫe���cu�W�C�)H�k��8�}>������!��9A'N�eQ�0�
9H|�rM��֪�ݭ58&���Cƚ�j?i�a^8nqӝ��>��o�L(��,"B���*���*ۣ�f�`�)�������M��8#��*˂9I�:uY�=�4rm��e bZ���C�g,�ӊ�����U��N�E����֛x�@y��r�%�~J�k�4M{tt���o�涹�.F=�&�7Xr�'d��EXom�+ϯ
��e:���_.�ݰ��Nw��j\�#�m�E�:�GW-B�37,eF�-�+�D�X�1?"Ʃ����YxDU�#��+u��R�NRzsu^�zU �S���W�-'�$�u0���kì�_���$J���ݶ�E��Z9M^��د�	�/��-WIn_���M�V*��i�ы��_5�NF�#���h;����v�j��ڊGd}�q̻ퟕl�}GZ���������ѯrCO)�rLBve�/���J�����R%ZPb�G��Jo#im�M���45f�]�S�hS@e<����6\�0�^AQ�����s�,޷��y`���qI=����(�����<f*�HPz\xT	>�:B\2d���p��FN�q�ր��NYlsk���a��g�3$9��I.5�t2��gY����#�a����f�pA[Uo{N+��=&����D釨�f�J��|���)�R��v�]�����������Z�1f�V�󍽅�_ɦ*��Vw�A٣��-
0��?�����Wu�ᵫ�|����9U�_���,+˶������<�0o�7�@i���vyd�9��H՝Ҙ�l�&�Sx0�y�쇙SUD�Gt5�g�Fɪ�s�~��#z�~��Ԛ�C8�a�[�,x��Tj�i}���4�2�ru=h�G����� �-��L���\�����qy�a�+�*��ԫ��>�✛o�9����ژ�3Ӌ�+��VO�#�}�o��r"��S���O����7�)�xl�mU��#��:����k�*M�J�RK�y��c9lU��_�7�Ȳ=D���]�Uí~<^#�K� J?�p���	����?�$��/?~��ovd�:��[����>PT��w~�d�
I���/���_j@'�e�ג���ǣ�[���,�I�օ������(�k���l6���A��6+P��֯K�\�۰N|-��&��Ѩ��wVI�����ݓ�6��\�Fׄi#|�q����0����/����J��P�JP��9Xm�+�Z]�4����(z�"d�s}0��+�t~�&���/�c0p2x�3�x�7�������@���><��EE`�o^}j���ogl�i�[�c�H�97��PH�@�bE��[�v����Z!R5�u�]0���� �˾g�3�`��j���5��(����ӒY��#�~�?Kiع��~�� y����r�
��V������M��ԠVHu����Ja|� �LݮGƝ�aI���t-<�kq�iӆ�F�e82�ԙ{h�pA�����3�Z2��T�{~|�pe\��=���ڍ	Кx۩*w"�=���΃�|>�j�eͪ���G�u0�D�k/�Rj�6z�0~!�Z��%�b/���Kg
t�&��Kǒ{��Rs�tlXy|��]�[2a���W�Nvz�.Wh�P~h�{���%`u�9��}P����uB�Ƴ��O0dSLB;�k����o6c����,�is��M�W�Ǖ��8��N�rlۭ�_��fE�c�����-;~�ä�P��~�-��r'�c-�܇p�:�k��'��b�࠼��K�L���>�;����Q���bt���:�q��F�^��]��t�.���NL�~K]�E�ejW�5{�pm!�g�!� |�z��>����=��T����B������Pzmy������-�vU�*ʈ0ϣ�`O!��X�!��t����I�T�z�~f����(Ҳ��	��qn�F8|Z�	t�C[UhR�y��>&��2��S���Uoχqf=�I>�����M�Q'�j%���!o����zJ�8X��ނ�hQ|DnQ���D56����ڒRm��VJQ���G��Wto�>�iQ�Yj��Wd�]oW���${2�!����_��#$�m�K�x��a��v����V��'I��oZ�����kD�pZ�	$��*N�rx)��OW�_�E��w3���"������v�/��v8� ��1�?��̻<�}`��X������zx×ϬNh�e@�i�-��z�w��AJ�fp{�U��ON����5��5�+�Tlq)�?�=g�nVgqڊ߮oÒb��J{�[f���A�U+�&���c�OUvNev�z�S��Yí�����l��8�u�t!��l�����:��T�������R�B3MJ�w?	[��}�I�(�}g����~�����U��V:�1Ќ�rڥ-��x}�ZVb����w{�貽�_�����r��c�Z�X����3W��qSl��o'���� ��3D���
�P�7��̽�#V"r�.�Nt�Q�<~��ƫ!�8ݶu��~������TϖMCq�[(�ޮ	`�[�
x�����C�V�1�ަ��i|/3O�o͔M�!ɶ��`���^�Jx#J/�(�4aP��n�U��q��Z!"ᱨ���������WO�������T�aא����P�L@w�
ع7|+v2^G�p������.x@���غ�����\;�q�i��q(�p��c,.��{a���~Ջu�{��j�t��6�me֐�{o�����"��ƺ�]��I'IQޯk\[N:@�<S��l̾6}���`�/6eǥ�x
U3X8�w-���A��c4��5	��as-�� \eU2��c��H�ͫ����{+P�#~q�YYT?�E`�^ax9�=���p��u��큩3},S�!r0��!����Wia�W�rfp��-~5Zؽ�d�`��Շ]<`�'.C��ԑ,�c4g�������%�P�e!I?Y9@��3��̄ڹ�.�L&���`�$S$0aw̆�����c�����i��6�o�:	T�� ��/ߔS�p!�x��3��_��,�E" �<`ж��ڤˏPsS�ƹ��/w�Q�K!+�㙙ڿ	Ϯ�=��-�����#��胄��q1k��9D�^�|����/�ь�A�D��pʟM��b3�g� �j�N� [ላC�������;��щ�]�3m�4�{�P�'tmf���(|+>>���2�0!���O��_w��*_`(�.FT������"&ݜ�!�b�VkqՉ��A��}�AN��A�7@^%��0F+�m���m��P1�ù�4G�2��Vn���Ϊ�V�d=@	�Z��p�D��В���HY5Q�H�8{��^"vƶ*o�]yי:=�m}-�[�sy��\a0�]|�e�Պ��+ZkD|���O$�fr_�[�}�Vݑ,����:���X[���J�,
�!���|"�v�ˏ4����4���	�1iV��J��@�����;Q��ׯ���S=X��9/���o=������Gw�,sR�����C�w�o^���s�(���Pe��R0W�!>-=��S$����TL'��{rap�&dì���,(b0\��.����(��U��AVp]JY�CѠ���K��[f�GY���M-�\����w�TtA:�;��xә"��L�����L����~���@�	��G���'d#󠫣�*��_*˪E�男t�(�@=Q=OYW���R��������]U�%-͗�t +���iT�#��Η	.�7�� &c�����~�s�a�?�L�TD�;2:E�44ݶ�n��KP���2P�����n������ 3���
�ZS�R�	p��f��ܥ�J2C�]�)�h]��f�.?����c�|v�<~��@<�ؗ�G9�*~�-�bu���� ��[�>���D�T?�2����G�/��O	M!gjo�)��'�@�����6ilRM�&u-KvL~궠r��2�d�&�J��˿��//3�+1�,盟�_ٕ ��h�뿨ћ}�S¦>G�)�.Ot�J��!���k������w?����s��r�qi¡o%����&��L0����gJ�x�+� �M_��Q^���V>����?_����W�h� �T!!}�徇�Κ�f��1�'��C����Ų|Ȳ���p�s�C2�tʪɩ{�9��PVE��&��R���� _L^|��oi�nQ��c	�s���n���ԥ.Y%y[��W@�����t��77��YL}���=n�U}<�pr�;����Ke!��@�%���pf��TH���.B�1�c�FXV�ct���5r|��x��wH!��<��	��n	)"��\G�k&�%ۨ��I1V`cv�	�cO(iH	�2�?u@aM6�@	�{}NB~|b�Vn��n��S�!��u  R��Iۘ`�(�6�W�w��|��I/��f.v�GZ��Tc�A�K)��|��E{����ߚ�Jѧ)X��/o(�N�^}�,�0�8B�R)x��v���X�s��p�kt5�dLy��<$Ͽ�dղure=ȪQ�0	�;[������6�	E� S\���x�G$9Cm�B-�۔.{K�݆1M��ۛҰ��N�ӔW��@'yMe�d�my�-��_����WjG�uiOgumvS�:D!��4µ�Эw�7��"$���f�-���ٻѼ�^1�� �����z�*��%PI�֠[�4\C|W��0��Ǟ�o=*Pb� ��S`Q��p��t�>����%4Enr��� ;BeŹ[4�6�� �L�Fc��7K'�F2c��S*��j� ��ٶl���F�F�$6����s���LJ��� O׳ܶ���5��d��@����|���E��`�ޚ�9L-�2a�nRP�<��Q�� �~�>�~Zi}�P?&�� �������Ⱥ�UT�$�v�G�θ
HWH�>�$��Xׄ��b����i���\\�����r�`�c ��Fy= ��c�P��X�@�r� �=~�0��qG1"W��I:���2�N��pu�|m�\���$���:���
�� D�,�|g�=X�"u� �g��4a���O��#����2��,�B�C�ц�S+;؇�,6}k��'�x�8�<^!k��Mv	 *�s��jB�~p���X9���X�	�ߗ�e�SLNt��V>�;#����9�Z~���n8�������&%yؽ�ḪY�0I��}���2 VM_���6+��6��8�A���Z݊a�*6�|Y��0���&��W}��C�i�#B����;f���S�2z;8��F7@Q��������ˎ`]͏#��
f�,�F�W|��  y"�����b�W4�V5�b�oTq�,�;툺dڶ�k/>�]��"�|��]S�,�����&�1O�T��?��RhM#�?Cmj=�6�b�8^�!��$��X^�Z�b���Z�U���z��~(�eͿ����p5)��K���o�8i�]o�'yM��kTr��Gsh��o�@�.��-JZ9!���$J�H����� �{T���n{��Tܸy5���.�n�!��ӡ���ƥdw6��z��1iӮ�l�@�-Ec19W.K��@B���e�\I3�&S�l�^���B����_�Ođ�E���@M�10��A��Z�D�L���FK�T��� ۶��Ie�j?A{>3d���^��I埮j�(&ƀ��
p�l�7,���C���_���l�~��Q��[��H�xC�)<������_��#ˉ�Da<�F�9�e�5����/��AF��"��J�2B���}�[}�9�!�nI�雹���Ֆϔ2B%��l��l��h�	�H�w���1��Ӭ���UA��=;��:u_�b���x]j��<;�$+s��nG�3LFbI`��W��4E��o�Z��-f��L\'�_0�?���ނ�!�l�����6���Ap��/����l��O�=-�'k�x��)W��c�C�``"ެF:�@�v�UJ�/G���E�,w��	B�Ge}����LD�*��#'��|8Vb��D���Ufm��&P�ef��n��gUK t>'v`)�6ģ��sL�pt�=w��h6�b �n��f�e����i�
��S���n�{yT�>��w�X����e�(�,-��	6�,�}su���"��95�aA���T&�]�h8}+.!]=��y'K���"��К����^�z��h�DPhZQ�2�
G~kHv���pRd��cuqL���u�#��	���ֆL�3�C%D���y;�Ã[J�F3��]rТ��`RB���MK�2�V��l���}�+�t�1*{R>�PcH��D��Yo��B�	[T+��ǅb8gG�4��!����5�{��4��X��:W<�Q]��j�c,u��Ӄ�%1{�w>0���r�ȍf��ȵ�
ۡٽ}���~��
��=7�ZO��)�a[8 _�H��iHF�+ɅjuL׷�N��ʳz���z��r�W1��}8�����Qi���͐mNU��6ѯJ��-7����;��mآ��G�m(ӡ1��Ѐ�u�ʤ��Y�:�f�s�H�=H�c2�f�����9}W���.Na%g�k��!q~?'��P�]P�b)�(M�������hˡA��4bH�����[�%����ur'�U�K8�|`�W`�%��	�Ag�C^�{��k� {�}1�w�o_�f*9�B"��)U���F�Ʈc'mǁ�����+p�7��[_�F����_��*՜������/����Ӕ�����g��������<[��h6gTj1�LK�\�mݗе#&D�*�sJ/��Q�4�(��u��`nl��q��(ͼsR(5�w<��5-�k��ҝ�q�L�R����k_u�2j?����$�@��9<pAO�c��:'���FFF����|@�������%��Bkٕ� ��'�2�d/�?�t��=?3~��KC�3CX��t��t�?�g\�!�9��n^19�B���]�\a#��~�C��>��J�19!��QgV�׾�V1���p��̭p��Nx�N�"��9u�����F	R.����m|;�����T��%��>aJU:H%�X�_�3�J|0���d�-�xi�!I�"�.G� ڇ���ߐ��
쵇�"r�g�!"���CH��ϟ|n�O�a�EogHB0f�qC
Z��Iysy~R���
�?������o��L���d�0f�jU�	'K��@w�kR�D}��� ؿ���<�s34]HyW����=$O�`g!�r1a����>; �L����\S壃+l��zP��Ĵ%�D�����3�����S ����A���;���Ueg���<n���y�~����,e���~;����x6Pz$�1ӮS$%v��>���n.�v������Z�l}L�Z���(��JH�S�<���a���׵�e5g+_�J'��'�˵Dc��8������1P��J��6��*�Ta��O�=i��ʄ�H�FO�Rox<��,0��te�63�`ae�=��V�&������Q��_�Pg���C��j����\>ŗ�%�q�N�9\���l����4:[�徲~`�e�o y��0 �F1�A��u-��I� ���1����:�wN�w�ۿ�Ք�	t�ܠn"#R��Q�h7{x��;���e{�|8[RCT�	E��kw�e�B6}ԙ��Ir�(׼�*_�k��Mo�۰ۯ>u����ej�M9*��<΄�
��OQ\��L-8,�n�/����P���,�xn�\���١~sغՄМɃn�pR��L� �d0]��Άُ-3>]E<���8M�E՟H"���~ޝ��u_9�duҜ{V�IТS�{�2y�%bGV��2펳�M�|��"e���C�b.��`)k� ��닀�&��kौ5��6#�h�ͺ�J�۞t��ܰ��mB��*�X�,���� ~�c�XPm���!�3-��$R��x2?� �)�:S�
����Xs�s gW��<�/w0�a�[��Q, �;�p�\�F���L���� m+@S�tA`>���ߙ���Z�����,�,�/G�g@�?p�q�#@�-s d.n�e~��Cg�
���'Z�lɑ�/���Z6q-�՞�V�R�:W6,c�������$v_5
�<�^`^5�u)W�g��$�{s���Õ��;*��AԪ�[
�U��ڋ��9j��h�̉�X\��2�h��i��H|x��A�����K.���Ю$��hbD�����a�R���3s�
���ʡ��~�DY�f��Oœ�`&���N�H�~�;�Q���O7�0g�7�)X9Ѫʌ�g;� ��̜��:VH��Wp�>IHH��r�ݽb�A�����H�����no�NTn��?�H?yw,�����QF*��ȝ��ߓ��#H˸�g�t@x�����b드��C'�[��m?����穷�ێxk?�x�m��rޤ1I�cqK������M¾'{�.���G hR����U��M6<�%��Gq��C~��6-D_�pg�4�"YL[����=/dѣ�'�I�>aV���_#:��O!%��o�p
�� m� 5����l���,t��[5k����*���PB$Bzo�~PD#6�;n
��&lSK��k�^\���}���ƇKQ)����k����	-|���CL�=`�O�(����y�!�I ���ǼmeRЌ���Okn�B�H���*���	 ���`�4�K�V	&D�Į��NB��<�`�jTz�˵�~���/��.�-�DE�k^N�C�5F�8���l���Ŧ?��e��}���;}A[6��jҎ9=�oEg�����ߚ�j�	e�$��w����q��@:�����G[h��(��z��A����h?�V�9}LV���`
x/?CaG}�A1���~]G�%�v�;'�'��㇋�lUJ��!^�������R�\��W����:L� cyw��:�j��*�Ϙ �P(Oa�;��~o�Ps�3[s͈!�I[Vni��c��7�ɤr�F+�؍����<-�V�G܃�̓`/���4uw�y���2MO��{��Ӵ�)^O���HN���F�~�vO�>�jrL.*}�S�����3hb�e}*զ.79^��g��ܘ�sHX�I@9�j�2�'{�-��	�73�~2�w���3��N�a�ͬp�]iV�C�U:�w$�F��$?�*\
�F���-�6'A'-4;���r���sJt� ��:���T_@��(�՜��u�v�:��mF���je�m]̭����s�i f���0���\6�qJ�զ�0hǮn�f�
vИ���N�e����÷ؽɑc�9��.��*`��f�z���"7��ꚌK�����8=t!��� �"B��20序ň��uK�b�]h�5����s�(�������"�	]�V)��
(N�j�?7=��Qs���>㛰*Cq_'���xp�o��r*e���@Lg����h��<�U�vG4c�����\�6<
����-��Q��yu�pwX��_��6FU��m��N+(�G��`J�yw��Ƀ[N���߀�}��䯗������M3�^�Ƕ���8�Q�`n-v�sR( ���ח�Lo�į��	k�
�jȈ��*޷���0�0~�Fxw��0��S�C�:f"�h�5��ћ��6�Tإt蛁��t��ћ"'�����������	S�3�p��yur��唍�({�=�G�Ӻ`��53��5R;J�um������s-���E�a��t���PP�������;c��$���ިY�,�J�44*�V��y���Z��F��u�f ����|�MF6��S�^����!����U#g�5����lP�$t�++�s�	8�A��~T��4��C42�K�DrA��A�Il���4�MU�@Xw�J�O^8��Q���{�	���� �\�M�U%Kf(�x5h������OQG��x r	}"Jb���w��哠��TFo�MJ��d����.N3�'6Xk�!5JL�w��Q��K��$�zh?#b�9�58�} `����:!��\�I�V����|~�-{�z�/u���d���ƆW �����̫� �,�	��i�ї'.m����1%��;��Xa�@��~,���+ ָQ� xb���7�uK���AJ�I���F*�I�|N����,�Ǵ����/1��F,˘gT��p'���*�Um�+*n�3�F����6<o+<�V�n�r��4%u���0z�V� O�l*#J��U��������J�����$MU��6���<Q|���%��Lq��v�W%���ʛ���X�p�5w�sx��p6���m8�2�~8{}8�z�� Ü+�%݃�Q���mfՈs�Ŧ
KJ�FƴAm��r���Jw[K��W��i ��b��i�g^���4�݌  ��Ň;���k�� f��*��u!�|Z<��3���:]v��c�m��Ύ���m�ڰC�R�h�%�0��@:�i��L�G��D+�D�����(��$c7�N��ٻba���(�K��7��;*�P�r hÉ')�tt�k�zO�x��xˎ6������w��m�/�oB������=4�Fkkĵ{3�ac��h�퐧�y$�s��u�~>8Y�1�v[�R����pJ���i=^��Y_b�or��Y'[��Jh+����xӣWP#@�7�� ��Μ�j��o_6���J"�s\���x! �>��9�P���8^MC�eɨ	N��fIF��.e����;��ڍS|���S��?���Y�w�&R��&�+y�%]�2>(�C���`�H���G����͡PMy����%��`���Ǹ>\�=�׆�^X 21�X�g���:S�,��	����Qbᖦ[�r5.��i%,5�cD0�O�P�2��_���K0f@��N��(�k��(� ���ַ2�!l}Ho58ۤ�d�K���y�����8�����?Ώ-�	�������.
/����-�fsv�	napkm�gu�v�����<�a����G��R�C�pg0H(���������`�Ԝ�Ff+4������@�B����ʝ�t������ {Of|
��o��V���s�bSڜ?�v�?�ط"��"u)�����Y�x���P���O�ڪ��d�`㭔������|��z8�8��W�(��[���B��)�!��c1�����/�H��P~|}S�䔺��s����sꮯS�;&�0���`Y�a#�ĵw��(O4�IIH����mo�o���E�I�#	�
�m��5(��6.9���9ef���5��=񧤚��b{�c�0`=�`���T�!������߶�l-�%u�ߒy-�9٠��b!_�H[�0���j���~6�5�Uh
b!^Z�F�(�xs�s�Μ�G�J�Q����;=��v%C�8��X�`�Sm�*����)�&&��N��Q�O5ދYQ��+�2n���>>N�������o�\��Q=Y��b�t�*= �R1�0,p������ø��WC'	2@+�H�{%�����S�.��)�4��֤�Q���	��-v�8u�%�;�2�݌;����)��G�h��<T������;>l�ea~KN_�U�%��'�����R�ۺ�<�Ȧ
�;�SI��&���8W�6�5X����xܐ^��ͅ��oo�\�,�-0~*͹eL�]�y��b$���)��R A0c�5jV~�\�X�c���%�ٹ0��f���@����j������E��奣��&R����Y0Ҟ�-��,!��\ٺ=���]?��������ʈ��4,������.��t>:�7����4�i������62{��n����"$ī���qǁ�����.z���b]���F��\m��!��a��r0�3H8�q_�V (�ۥE,�g���I�������*t�=,^m��n˦��ws:>u��8zy�3�(��Z�z�}� ���AIT�������z�TR5�(t�)�k��� thv�'��q"����	~m��{�I ��,���S��hIp��Ư���d����X��v�YZ�Be�A|�m5��	}%\X	��U{��pK���	�(F`=^���瀊�	���Cb�֚d��k��&�����w��%�������^&!�p�X��2�0�C���>�!*�E?��_��Wo5�4���k�vF��ـi*��J]��MVO���i+�ˁz��k��@C�M���'pu[fb	�-���J�%��:K��1�$��p5y8�wS�?N�}�n�1���\�Q���D���W�+����;���Z��Ԯ>�$&'��$V��x���v��fS��7B�Pk%���I����ȕ�^*��k��њ�˙�����������������J�<��� &Q����A9��I��˽��B��9�~��� wD�:q��'��R���*�Rg��O�o��R=g�M��EH�8Kiz��é5M�|<���d����mJLC�&���Z����ƃ����GU��J8W����+Ǹ�����{��N���b.��K�O�ꙻ+>\C�#����"N�m�5�'P'��>��N��c�	X&�zt�,���κ/+y1E��gm�飋���/���kC���^r뤙E�ŭ���!���ق��*��=KB�~D��l������e�Vv�w%I(��Qf��j~�&P]�E`CӢUZV�4��O%DQ�v�ț後�{�*�{��1�V�;�X�<H���+�8�y��з�(A�-*.*�c�pV�S��3���㟁Ip�"#-�~�,��b��eK_�I"x��W�������HD�;}�����i@���b�b':n9��&���_D�Q:K��v�M���H&�˄	�o+�գ�+��ʡ��V���<6ɱz>m/�#��uqI@P��!HЄ�q3V����G��΃�@VX�h����ᨃ��K�(5�:4����}6+97v|`c.�cv���I�$� ^3#0o��X�+��f�y������3�;kU��;I�[E�w�j��K	'���6���R*M����ɠr�P�ȸ�|lX�q. R��h�@�	�|�(�t���7���wl"���77!Yڟ����>�e:���a�hS*��=k������L5Ɓ�%&GbXGV�E��*�(���is�.�5~�,�X/�'�U�2p�,���&�ٮ�T�[.��P�?�-w����[��6�#�a���p8�x ?���K��y ����U]��64�Ʌ�`����0k{q�A�ja�Q��Y$U�G�}qa����Χ��5a���:�`���$��4�~#����_� }0~)2"��������[+_.����#�M6�0M�
u���R�%O99{J�r�Þ��l� �>���ϧ���@aC�Aɶ��D�t-m���/��>`�dh��F��}�NI�u��#;������u�Ǽ�uR�MtW�!P2���O�[��e����A�ă��8;x_8���q�L��t��;H%x��-jҝ̕p!$/6WK5ǎ|}Lh$�p�.���'��
h��IV�k�w�^_HkbÄ���5)씡�6/�[�v���;�Gʩ�L�XtZsW���.дr`Ø�:VL�hEY��<�b�n������j��%!�8�{.^�9��H��cݨ��m]ܤ
 ��_���U���?uO���T23�i�N�&��CD����燸�2���ٕ
!R$q��D��+�P1�P�:�����A}P�9-�b>h�"�x`rhI<��mk���e���*phu�wj�ջ*�Q@"ҁ����0���#3�5�[ʰ"��J��-�b��P	�@VQa���er��	����[d�[�;%M"�3R��P�Q�O�.�jn�.H��p��$�i6$m���w�2�q�J��9r4C�+�|yQG`5��A�̡����L��ZI���:���s��M�7�LS9$ ���!5��"vF���Z�`)j_m�,_��k�tT�̚]�ʚ���[���Q�>�D�q�����~���qZ��خiX��RC���c�C?�nȂ���^SWw�R�3��|`�r��S�Rܘ�C��G���-�@I鵒������[Y�p��z�C���g�P ��}_�ҐV�Glؼ��A�kg�� ���'E�y�G��cp�S��0�hSp�0���S��6Qƒ�ڏ�p$��Η�𖣧��
w�ax���;�\e�,A���XIxn�B&>��Y0���޺0�`�Kuޟ�.e|�V�:W��\(��J,���}�9X�#���v�;U�������C�wv9����D��VdYg��G���f�Ѹ�BͲQq��j''W�}���:C���&�_������B.s� ��F�u��*����^���|���냙�;���/ݷ�8 ҽd��Uso��]��e"&�"�L�u���cALQi��~@�����'MyU�m\Ϥhet�x���qѺ���2�����cV*m��	���%�_0��ځ�g�q�w_4�;�썄ra���n��p;��8S���C�J��8��}%��GJߣ���?]RQ}�"V<�F����l�'�m"�vP�bI� 	����WC�ɠ��&@�&�Y�4�܍����� �mS[v�c��s���l^�TY7~�- �j�v�%A��-�yT���H9�2mF�p[�����Q���AA~<�+uћ��}����ND#0��P�!�N����?B�<�'�Ȕ:���e�>�_8�Q%����l�.�$K�H¿����p��R�^b?z�RQ�K�g1<+��f�Z	$x\�w\5s��?��07'����� ��h��>*���!��_;#�����~�k� ��d(01e�O���en`+ȁ��X���qsY�ŏ�B��C���D��9ϡ�HP���QV]��2 u�<Ι��H,�E\�?�VLpwr*8�G���?x5t����K�ʪ^��`��C_c�C(DQ�.��� U/��#ˆ"��U؈��C����h�g>HOGT�e�W���j��� o�D��2��X�Ž���II���P�]����ˆ���SfX2.�!�a���~;��՗�R��+9�Ż������IE�zih���@Vt�������@�?�SS"���7��I5s��nЗï*�!��vBe����ULԺc{i���N�3U$��v$v��B���b,���+a9��s5���a}�ϙ!��QQ�|��UN��+佰4�s(���
"��u�ȜH岡2�Ʌ��)M��p�$�%�;���[!����$�&?S�G������Њ`�\a��������GЭ�V4	I��ǯ0[����w��2#b���d��?��sE׫�Ҏ�z��7e�K��چXBΥ�+���e2��w��2���1����P�B,ul���m&=�����:�m�2�Yp���	��O�"%����|���{kz�Ďd��g�M��0-�u��ɮ<gl�e1�ߢ�����d�e#d�̾�B-=��=�(���������*?1�$��O_�^]_&��Жhy�V��E���Qfs��/����(
L[��5bM%q{�����H��ހ7ʨ"��d[��H�+hӁp�"#dˉ]Et�2�<����nߍ]���n���t�]+�OH������߮��=Oޫ+���1�N�-f�����Y�
Kk��{�k.Qj}���`ɰq1u9����r��U�+�{wm<��#�n�Ǵ����ti��T������v���n0���p�'Fx���9F¦�	�e��[�W�ݑG��V���K�@y�]�Ԋ!��=���7��v�߼�]�=�^O�p��RZ��ۣfsq�$���'�{[o:���a
}H-adRdV%�$/&�݌g�m��۷����=�l1[�9r����KC�y;9��O�,ߐ�c���9K����5�I��g��9,�[�u�R�H�>�,���2��:���%\�q����nF�$�>oLZl���Ik��eu5�׀�a��94$J�ަFă���es���#�X��]��x�yY�2`d.O�Q�d���ö��(
 �׀�R�ɳ	�o��Z����K)90�9Z���@K^��8oU�b�_
dQ�N�Μ$��4��"�ʃ5�*F a�e�ˉ�FS�y.tv��|z'�ج���6�'�x��9mv �`�AE�Ѳ�^���;��59��?��I�8%{�3��NϜy���D�
G�DS;֕��
@/�x����Ł���dx�^o����Sf/?�Q�>F����-?ҭɆ\X�W�/K��rf7xorV&	LṂ&����N�_Γ�pa���� Q�uhK����:w$Z1pf���Je�=��'N�O�t�'��0�C�efӐ���j��_�C���C�o5���V�+�Eu�56	�<x2/��ϓ����tj6qI}mq	^�m��Gu�	��� na��O!��+��Q,!����wQ9٢hvP�`��,���ܤ����'��(9���'�LS\�;������S�����o��U�Єoz�����v���E{�F���"����=ld��8X���;	qw@����)l��(�(�Ic�9��?
�h��sP�#VI3��|xu?`�ɚ�Dc���y��.�H��kP3#KNL�]��1U�Fٗ�����_���2<�Ɗ�}x�+jG0"�ZD�|�	��wn}S��j�3�/�[�4�I��.>�@@.��v.�W�S�)�TF�H��.޴���	�.M��R;�`�E��ߨ�hyP|9�<_�^'�J9i�B�?\"�Z6^�k�y7�!'sI�ʞ%E�$�3��X,�[ѽx���HX�����v�2}t,��cMc��'*�v3Le�/�co�o�H��a��0O�ۭGy�񔰱�ZY�hy�e0��!���L�L1:e1D�L�����h���RoCoO����{��f�?(f�K8��]]͘�D�[s�@�?�&��{z:�d�����L���V��>1t�����L��蕃��,|p���Z�1JP)�\)����U{��S�������ɝ}��]��2MS}��t��wb���/��0̩+�6���p9XT�o���Wu%���fh�(�s|-�,9�Fɻ�S��har�ت�ey�`l��\�k�W.6�t�;��a�S��^�KĔE�%5������Z����:!'�zc�:.��w�E���g14~�7ea!� Nk?���&Ah>%����;��@�e��4�zIA��>8y���pz{�����x��>!^�ZI�1}G�l��Y�Yw_HW�H�^/u[�m�Q���2�y$��#9�ꎡ&X/#n�G$4^Z��hX�m>��dV��)�?�>���S,AHo��g��2/m? �`׉�sI0o�_k�#���D��_ X`x�kN��=�P��"i^���šl/i�����g�0��	�D���>�l�
l�(�:�r��j�~�3Ը�r5�ۻ�}5��5� 5p��rׄ������y���̈ys������U5=�ԇ���]o'��0u�o�w�F�3W��n=�h�� ?H�b�e8p��5��ߖ�ܦjWI�p<5>���6�U�o�
�hWՉwk����_hRz�u�[�������R�h����Hے��:�]Rm$&�)^"���?5��RނP|l��zV�$2.�W����Y���[[�X��+�nfc�,��x��γ7��&���*���Jd�[��X����7�񰞚��"�~5D6U��lX�����)�U� �pf�����]���t(C�r��~��}��,��:�LS�|l�堏d�$���dy9~��m�p��ޠ�;U"e�9�_�-�>-CⳆ�f��(Q ��V�m4Y&II�((x/�����uBl|�VJhoO����w:�� �[s-�M�ɢ����"�!R�8*As&~�	��8v��y����\�O��l��̮V�M�-�I��P���=��G��ܢO�U�Y=��Kp5�����ʯ��8y,z4T4$x7�\���� �H���(B����� "T#ޘaͦ�n�t&�}?C�Mr"�i�0�W���Y�[�l�I^�=�?���O��X�!�9z)]��Oc�i��l�w�� �>���Z����t��/[%?ݩ]��"B����+�e���b&����w���.TM��g0��c�{.�}��bP١��W��fP����y5sDJ�A_%���/��>��Y��#8���+�-�0���7�#��'O��P%+�_��H¼��?�m@+���I�f�>a�_r�)�C�*٣؀��УעL(��.]m�q*�y�Ư�H��z3��7��1$��:;�c�n(�0O-[��O�u"��|����`�_�گ;�J��H	[�'(����>,Y��څ`����U'K	bA�);���A���ͯ����{���N�Yo�m�qC-6�P$��bQ)�M{P��r%+�`>�E��{�>��@J�ę �a0h�*jJ�U:��cjq���*��w���:�.���YemI��#>-�j��� q���1y�#,���X�!5�]��=f������L�ܻ��
yּE�ϴ�$�0 /��#��-Q������p��"�b"�E�d�c�)����cOӁڀ��ك���h2�~y5gm�;��l4⮘3����΅�7�54D�E_�p�,�19���r�:xWq�v�7�&,�G�̍?��}i�����F��.خ���~R��A�|a{
�y,y�h�����mUOe�%�8��Y�sJ�uZ0ʕx�Cb�@[������ց7�v������!\�Ͻ�-.�К�'�@_��d�"�'"D��lLg�O�`��c�t�V�r �S~�c��)�/;�A?A`>@�^?���_��9�pTn_���#8_�l�PK��:�(��.�L<��pEW��`	���q��?]�G�{'�Cq�àv#�X������@Z#z�� ��x��ό���@u���E���烰4G0y�\����o�2��¨�%ܧ��M)�:�뤞�)w'.�@�m�O
�@g&��1�Ji6�(v^
l���V��3A�d|M�ʜ��`;pz7�J�x��#GE�P �������NN����<���L������(�4�_�m���??���EL��V2x��U`)mt����g��x�IP��Ua��Pn��&d����m&��Ɂy���Ò���ba��PY�L��"l�	Sf�:d	�B'u�`��o���*���� V{R:�y����v�|[ch4 �bM��rT�:{Io_�~�\�\����k��	��	5���P1Sf
d����Ʈ����i,��I)���5_�o���gy?�?q�dr?(�["�v8M�4�p�پ.M����&��~��^ċ�;��vSPݵ�L�?;\Q-%-9�noؙ���oZoȳZ�o�ǿJ�%���%5�M���N��7(1v�Ⳋ��#� ťY��8 �[^�1wr/�I3��滳j�H�����4������hq V,�$:3�M&��3�9��}-�in>`s��Y`mR���z�k��Ӕx�X�<�a�N
t�����<��6��yf�2[�BYU<ƿbp݃:Z�Ǵ��cі�l��AAJw$�2�[{<�U\2
D�&����d�7�O;��f��֛k�>� |©�����7c|9埶ب�>\��	Kuy��zZ։�c㷨�h��y��������A�Y���o �'�/�f�t"!C�l}����^��I�!�g!�O��tԬ~�7�<C��4SJ��t�S�^��L�k��赞�dV��o�`�����nz��#�bL���Z���9]����u|����E�(#�14~���-��\m�5�F����kx�}-���J�-ꋅGW�J��i1��|�[�
�}���y�/6F�2��<a@������=��O��!�6@׭s�:�LUO�:������&:�V�_
vE�������-��&�9l�ە��yY?&R�:wy_�ąW��ڳuF�PO��ɔ�A�yPɭ�n���?���GttGU�q�V�!��Mz?n���[0��0��!^��1�~5@�Iv!�,@�D��ҭ�:��0�m��w�����iK<m���H&�RFY����]ܠ-?����6��ts��M�mj�k7%�1�~	�S�Hf�U�.�����s���{��&�֜޳�t"˵�@!`$3��09��e��0���"&��*p#��l�;��'��i��������y��᤮�H��`�Â�c�L�{�'> F�	�7�1��|�|	e!���P˸�չ���6�0��f�%�d�"$k�GHH���Z�ť�.~VL�aj�����k�����Z�R�*�C�f�p�����6���Θ��h�Xх��(�&�����n��p�R���k�)d�ٚ�����|X�(���>�}���#� ������kޡ�T�}u]�Ҧ�[�1�r̻�F@��W��G�A�9�=�C���z�»F��&�`��μh�0�V"�i���M��[���N)�V�D���>%7�]�"Rְ���p���g�43�5P <ۆVU��)2��mss��m!���X�oʈlo�ɡ'� ���5Rpy�g��C�R'����8�_�s��A�v�� ��5/Oq͓��쭶�Z���s���L���:�j�:�F��T����]��M�g`[��ZC��A�;�uKujR�썥����z�=L56((3�Y))K�]q`�Q���5�;O������H�����߆�b"�Q��Wtv+W=kV!��A%>�aY����3�V���7�rK��~D(QhX�$�(������h�+ȽM\{۷���+q��+[q�$?=�ވf&�U���=�����
��Te�lLb���=Mg>�3����b[p�ͩ�б	oy��t��!o(��i��2��Z�O�;�y�������<>3�*����ug�s|�dQ����֟���=��d"#���?�'���JKW(TEP��
�f1|�@������&Y�:p�f��,��I3Ӕ�<�"�������G2=�nqWHY��SsN�M9}q��6-�o���%7F ����U�km�� ������Jƌ3w�� ��u����3��$>�nQF��j��!�>4����t�:�XG���>��P'}��G��w���#��cޑm��x=�T܀3�'���Z��>����q�?M!]��s�y��������ҋk�{����J�y��NT��
g��(;|Iw���㡡Ȉ��n��kަ�U��Й'|���h�5.���ʸ�E�O/���~��8
8e5D��t&��S܌���lӽ��`���]��S�A�5Ľ�m�Afar��(��{�D~L�W�U}���\T�mO�I�M�c���|�����+�o_e]�T�/����Q{�G�e�_I�ń\B3z�ƭ�R�/��v.?"��*\��/G�Ev���V��v���q�O �z��V������)��u��r4�, ���#���!e��=�����=��I���Z�(�- 1ۮY��ه!5N.�V��F��������a�U�ǦnB��f(��"$|�B�KR�^N9e;Jt�q�ϙ3;-t�X�^P��9�V_�Oef@�O+?R�z�6r���I�����࣫S?���}�j�T��� �������/*s:rX�ȫ�`���l��&��ڰǩ�@��~Q���UEh.>�՜3dT��3��*�آ��R�٤�����a<�C*68�3���@%�'�Ș+%k�!/�2��r<>l�9�����T}ԟ�g?�97k�@�seD6�JYâ�]ٗs�g����ю<��U��4�!@6�(<��-�,�� ���`|���7�,i��߽��!�Ua�",*Yh�:��8�����Tk��g��a���G�����Z��i��lwj�_���ޡe�X�
K�m��a�L�2��+�O=���E�N�R~��1j��Git��nP]�mͤB����y��iߧE��ѷP������AT[�����B_V�m�Rƨ�YA�O��g!�;H���|"ؔM�b��Z�0�� M�?��A�!ɰ�%����	�3��$���i:x$��,W�u�,U��A��6Ց�h2�:ݟ��M���A�&_�F����q�����s~�'L\AG��	H,�R�����"�ߖ��װ;���Ms�������
����& ��{5��	��ѕ��,FK(궷\�3�9��5�0��/~��W�DU�]��2�B�U{� �L;ߣ댤	ښ�r�NEC-����!��2�)F�y������������¢�wҙV��?���V��WC�"��hÑÕr��ŭ�����������G�ϓ�Qw��6�+GI՞��g~��H�8����f�#;���C%s>�ht��߹����0�s?
�n���*���<�;l�)|6�T�d��Xv���i��!Wh�u���0`��iݓ�.�G�@}q�d�|��z�WIH����=�Wck	3�(
ζQۮ�C�?G�x�{>e�$	|�� �B���؉aK�����u���j��BE%�2��H3Vj��R��5�RE��B�����/ ��˰j��'!}S�-i���ӯ�>6�ʻ��X����u�K���rʚ�p�s���[�;R� Q�C���_�	BA1�˽T�FZ���q�j�\��,h=�{�ת����'�K��A
�'sQ�K�X��z�.��L�j���E)+�̳/�	��4�����˾����z�xY��霡��F#�U�:{4j���V@��������Xˆ�%�����d�9�(�XV��ӵ�	5,E@߄f�^�]�f5�C��x�{s�T�9E���Ѐd�V)�re�sq�ZnO�z#�3	���:;V@�ݶ�J�4ۤ��IEu"E�\�W�����&�;��&xgr�XI~:���iUm����Q+p�8y�;�Y�d�QN��c�6��S�m�56�7�W��k��@��@Xն;���3Z'#�T����b�j-���BXL=�l
���Q�[����
���>�!k���vϟ��g�d&/\x6��h�W2������^�M`�3Sf�>$�ꧯ=�k��x�Q8\�:��(->��6���:v*�F�&��oP_�����S��=[w$ё�zL""���1�q'�̑CA+2��
�7ʁ�+��7�y��1�)�,iy58�^�;Z����� ��A��; ��'Ve����o|�`���l�����iz&�Xo�{HhN����*��V�Y�<ɡ�u�S�����W�MAo$�rU�H/UC�d:�޲^X�-��XlL�F���m�����@FmM�ا��(�t�����z�ݓc�U��#~&�X��}���P|HS5�FM4p����'�� �FRco����W{2g��A|Mϛ�	V\;,��:�z�T���1�8��sSt��[z�G?�۫��Q7��t{�k�Ws�\~V����y�:��O�t��c���{�֗0��=2<�E5
#m����<��GY�i���^/�|�)�^�E=�7�?��`��G��� Ś�-��z�X�\O"َ���-��޳�yC8��2A��_���O�h����R�֤�����pqq=�,�*[����>m������;�9��n�֒T�0��ɠ��/�ʠJ�r�����?�Y'���;s�U9���N,�����������o�sFf-���ho���!g�I��\�U49��x�����WhO,i��"Z׸��`$pE�_oE�N$�A&����ѩ�:�!H"��JBX�-hRƙ6�t}HhC�t1��;��Y*[����6G!�}�U��cf�L���J��㐓	����3Ipv�]_ ���yd��Z[��m�����/��.�&s�*a8I�Z�`^�?��*x+�	�zB�*��m>��M��m���w��G��)�;�a��� ��[#T[?hcI�8��Oܡۮ$�8�>v�#m_x<Kw{Y��Q���S�Xk&�w��\HǢ�"���?���j��θ��$��]�lA�eh=�x�e�1�t��x��wciVms��%��+�)�?s�ūbM�� �t/$4J5����n��7ZA�$��' �繫����"��k���]0ў�$jF\D	����<n�6�t "��ɘ�ҚDc��U"Dh�U�g�La���H��n���7:5�D�	��J��o��+�*�������K�o��P��ߑM����C�lնQ��r��sD�2.��&��n�`4�g�־=����Q{hi��7[wMK�*4�>�P���@w-S`�4��xk.����Sw�/a`��4,�W����Z�4,U���M���Hn�=ˇߟ�m��1�,~��ɐh�����mQ����я
��DL��p��ԥGE��Z��`f�/�=ý�N~A<��<9�Y�����\/�����2��2QX�D�b���Dr� lD�4 ������5�X�Z�̓'�QeFBH�T05����o
S��JƝ�ܓ�)����]p��e������ ��aff妈�ݣ[�l�I�Z���F��j
\xU�]�ϑ ���&�op�z�P�L珈p�s�L�G��1��@��e�=���H2Q\3s9�+�D�W�mâ��緀,\7�dn?���%�Yh=�����H�{���r»6\4�m\�d\�7�2�X����`1H�+�4�YS��?0ZG�����k??����a\q�?��I��掇# Iݘ�lCѹZ�$�S�,[�z��`r�/$m/�Q1����^�UqķelC�Q?jf<X��>�>��z�����1����s��g���8�2d�☒�@!�V���j�҄WQ�h�ږ�v>�����M>���ݗ�o��Kd-�����&��i�^��q4R5�]{��T�Qz�E�<t��Bq0D���҇:�������e
l�����x��YF��Ü쫭?������K��$E� (%l,�ݾ��ܶ������[�v�2��PW�N����7e���N��T�acN�E�����<Ů���cs
Ӱ�n�I���Q�׃1DR<_'��o�4�v1,�7ф�x�?0��R��giŷ�t��m�ϐ��u �P1|��a4�L���.������O�\R�V��Pi�e�2ί3rN}J|ټ��M�R�r�Cl�)���Ǡ���x\B�ֿs~&�2=ў������z���|V�YAO-ZPƃ�+nG
b����$�9��b�8��1z?7��K�5���{@�TAdE�K�F��[�����#��V�I�{��G�ڀ$g�1�Q=���u��V�no8�j;���"��{�!�\���t�`�����an�k�-���PRٮ^:��9�W1R�r��A����������d�0'9��D����%)p��U0^W!�k��!b����<x{?D�o�~��˧\�H�[�Ӭ�]������w$'Ft�!�i�Y�]L3�pٺ�[i�>p\@��Ҏ?�F�?�󛛷��mW���")�J�:�"#Ԭ榤�
\D˿���H,:&�\����*T��pC����~�	[:i#M�6%6zY*=��͆�9�k��+�����4�����`����V�l���'<"�������/Z�$@f pJ��6�Ȱnµ{�0,f�K�{���D�m��Ba7	~���D;֤-�R���͔UY��'_���2tf[y�n[������>Q���Ĭ1g�b� r��ƈ�h@}�ފ�J�q*r�iG�`@���.���:�-�0�=��S��"�X�)gQ��W/�8��,����ܓ��M hQBo�ڂ+���V*�fY��>ZR�{UWо�|ۓB1�١��7�A���6�v�f���@���XM~zc��0�p!a3�� +��a�(�O@_��{�"%��)��DM��2�c�q���爙)�
���n��Z�~P����yݻf$�J�+3����S�x��2l��ƭH�i�T����m��_�X�pph?�C4N��F8��2'�&B/n5�D�"�cq[{_8��y&�B@�%�����[�I���l=H$�g�演�/j���=\�������.U9/�D��|+,L��+����h|����'��L5�sI���$`���[5c�����H4M��wj�Hv�_Y����$�Y�e�M�5ݞɼ0���5f�ނ�2{z�w)�qD>~�ף%�<������;�����9- E��CA�x	{̈��������O�����	n~��m�bp\�r���_Mo��6��j� ����I"�C�!��x.!f5����}{�O��j!���B����A��h��Cֲ����:�YKi��]��#�񺵍����+7Cȼ���:�m����-e�"���ݟ�g`O!7��&?��������J�k~^]@��M�Gؿ�/�ۛ���-zg��Ӓ�I�A@�51�V�ۦ ��:���S��VG�/������Y��^s��Z�~n?S�&c~�>��W�؈��oz���}��8?S����I���c��=����`0�Z��z	���ÿr��;'�+�,͈�n&����OM��;���&�i���zn�.���!�c�����z]�
�C,wt�B��N� k)���O�Ɏ���%(�����߅�г�XPܻ1Ѝ`Z���z̄H�sh����	}���$(�YʬD��k�����^(�P�p)%D.c�}`���&"��'k4��q��!_g-�����^pR\X��Z5Џ/�!�C�T�7�e/�m?�g��U�ڐ\��s6>�	�[2�E���xK1d2ۏ�@c91`heQ�����$�rp��jΝ���I��ewp��!3�%=Z#ےҒ/>���^.r�c)>�=�V�9O��/O��K��P�Y�F�3A̝S!�n����[���|�V��/�RjE:����ϼ�~�]���[4�5�o�
O�_[��i�.s�W�L�6�U�
�WD��Ԧ;j�E�	����ػ�$
Ĉ�(�\0N�[�cf�R�~꺖6��k�F�\fB
���Df�Q�5�0K��f���U5_չ������z��ت����t��n`���{�1�~^h��Ռww�FL�$��t�߹�P����+��
�����D�7��h�v*�O�z�H]agQ3�_HA^~3���������<�9��A�y�.�������JV&l���ɣ�(��i32��@� zN���fU������קF.թ:}�b�YX�a�By�*C	�y5������� +
�,����\~��.U=[*=j����ު��+hOd4��+�ox)�bϽ�+���wA�q��nH���$\J�0���t\<d���
*ċc5�>i\�r�(�޼e\��ܕQ/��b�j�Q£�����<O�D�*0u)�ܜ�6��-ks��1FE!�>cM( +ځ!����u8���S�oUs�r�G��-:�[KH��Q����n�fi���I2X�]���_؄��w�܋�������ă:�ghث/ڳ�#�>a|HcdX1h��5Vt0Ev���xvDɟb�H�u[Y�fB���ǎ�`�jYH�D��U�	2rk�<����&�'(�S�I:����;C8,��7��DJS$�p1��N-e���WϪ)�!�{���M�gCķ���V�sNx~8�"�i�z�#[�ԃ)��.��+��s�sC��hN��WTav�Rb�w�`x��H6yRB��:}I��Ow���A� �F�?��N��x~6L�$�oL�x-<01]C�~��#��z��U���j߻�%D�FG r��ޮ��[�|��OT��l}���)�l#����ޝz�U��f��!ZS�#D��yQ
ٌ�|^�BA])=@�\j~/�Жji�����ZV���chZ|If����u�P�����u������~L�a��d��=[^r�����>h �hNU��d�7B���ZsY_��1b����L��KTUg��t�x%�A�[%Ub�M�����k�4��:#����$a�1M:W�Y>��S�to�U�i�9�&�O��.�J+SZn2�Eب�9��,h8��x�/%���^t���5����%���7"����vK�MTP����wgq��@�����%��w�y��p{3TgM
�^�_��؞����54l�����8���2矄�ȵt�ߓ�h�라�UP���\ ���*�Y��(~L��)s����}����q/c��@b��}�!����7�<�/�#�x���g`�vp�>p�!��|a�<�����b�A����uw
�37��1?��˺� ��e;#2Tϒ����2;0�g�j��ƪF���݂^�F0	�A����H�iBA��Ԍ��`Q��-�>�r0�K�ZBw�- �U1^hq��m��O�iL0��  A^�e�_,�QD�쟖�Y?!C���Ų^G���T��P�5j�Ǹի�d��ؔg�}H��w���P>��"���P�>g�p��V�|	�PBőpq�f�2D����4!�X�1
�G��+"�X�y���S�6��o�d%��nW�s�՘9&Da���	�jr@�J��r��f�C�=�
L�4����0�8���I_�����R��
D�\��{~̈́�6�N�������aRT"�'sn_ΰ.c��P��Ed����/,�W7���*+� �9���{rx�WB����%�W:�q��2�=�� �y�'�����ӵo�,(�(0���	�5d���i6|�^��x|�|!� �+���e��5j�\��]�r'�6R@,9��a2=�@�N���J,�.��j˕J:��:u�.�ejn��v�a�:�"'jyGu�p̔�>~���8�)8�LZ�kA��I[M{> zcG(.��xZ�VKr�ǘ��%�ZoR�1 �۳�����١f�)|�,�e�k�ya�$Et9e�x���q���cU&�%�nq"��I�����o�aޙ�߉��/�����aq�)k����q��R��ʳ�wS9�Ҧ1w��e�p�Ņ�s�"�}�9&�5jV��!��J9'#
k�t�����(LF������#������f<��pJ��4���4%�
7�m���L\GtٝV	2w�u�EAʻ���{7��A�$t�Q���n��ᛦp��8�*厺�Ve��F��_�Pk�D��[�,Z�d[�w�f)��þ�2�*c���tpcq����k�C5��~��ǯ[
���ƃ�����<�~�ʗ%��KJ��N�n'�����@�)���2�.v�9��1m���	^�'���=��z�g���ѫ E)����Y�B��lL�QcY=�e����<,��Ĭ�TQ���r���'�ʙ�
˲�s����BR�0�=�d3%n@�V����E�/َW���͂}p�=1扚~w�i �}bo�L�rR�WU3dwpBR��� Z��=6E����'�@�EA����3�If�;bg=�b�RA�*lc��6�_��{��q
���IL��ft�y�CG�t�@���P���[� ��߱�Wܫ��M��5���+�H
�Ӗ��陮,�,j�O5���ÿ�i�P~�jw�)؟��f͡���)A4@�;�V���$#�u�ޯSm7��h���-	��>�5P?�����T��s�l��1s��`T����O�|��tҧ����)�=B3�5�Bn�EGȰV�u8q�x�p">|Cx�s����A^և��@��A=�����3P��k �\�H��}x���CB���S��oeR��~n7E(Q�?����c.PQ�ˏ��}���uw�2;��u��u�3Ш��0yy��3D�%8�H"D#B�^�q��b>���H|�Kz�@0�Rq���%��QBUy�h.v���Z<�K|�P29�ɍ5�̈J��D~�M�U��	�7���x�l!�XLi@�u�>5Ĩ�4K�z&��Q����S��,��M��~�]	�,YcVh-iabʢ/A;b j�"a��@	p�	O��j� ��a�)ȱ��G�dG*[.��w�!�#�ޒ����%*}�s�dN�B��0{��Aڟα�bL���:��yJ��Kh�ʙ�ӅØ+�:�&�R~~���H�:w���vmz�4�m���)�#�.�0�_>�b�h��P>��A���I�{�?r=Ux�Q����ǪO�XT�0�{���]��%��c��_�t���,޻m��ߗ�k�O��8�yj��ش��W� ���r_�ڻ6�cm�"��xĝ�;]j}�4꦳q��Ik]N�F��.�G��Bx��ck�9�����*�@�=kF���ti�������ƻWf\���O������_���O�΂:%XP�w�}���s)�-u��7P��hi��;�M���-���H��Q����c��]�o�y�R�(���A8'���!
��(nᔌI�T\���R(nQQ�~Y���WA�[۪�3�ٯhDf����ľ�S�Y���OOz��<����K5�q�t95:����6&X��Q���}9�z*=�q���$.JQ���l�ͽ����J<�?��i+*6��l�}�"�����#+@�OƓ�;�3@Ƚ�}�;���Lm��w���A�c=��CZ׈t5���~&�lP(C/%J[�V�Np�on[^]�ǆE�1� _�����p5.f��9�q��
j�����/i#��IE0���#�"ᙯ��/�v..\�(w�HВtTj�O��0 �cZ&}�B�P? �Y��9Y�7ѭT?�v�B��gG���Q��VxZpT4n�=]�p<Z�av�ۣ}�r�J3�xG���%+|�
 ����+�d��@lp?��St�Į�8*�H�}�O< �c���A��"�į[(BV~�e�Q���T��G TI�0�M�B"�N���W���ê��I�����`Jջ%�=��e��̅U��{����qb��E�(=Y��x#��P��Z@Y�]��eU}������b���˽7M�����#;ʛl�a�oN�Q��L��M-$ ��u�5�e�9L:�J�ZN(��rg����A��>��&�"�ҝ ��y������{�(�����O����Bm��"y'F	\�p��]�����c�y��x��[J��w�+��U����� ��#�_6@�
�pk�ȇ�<�H�O]�ݛ�m��������
��;�Z7=zM�p�V�G�G��nkr,E��B6��h%&~G�^SJ�c����?+�\�+j�#�i?��7+����ܿi���u������`k�P.�vPyp��S�2�7]T�W����ηzi�06��Z�ʲ �LL�6{Ӌ�g��GQ?{��0���;5�QW|k��C���"�ȨA����z�˪�Q������:� �B>KO8}C�s�r{|�hD�J��I�&��aZ �3j���wk�� %lڳ}�z���|H��'����w�3�]ra�����GN���R���Я!p���;a�3{�6�{
f\��E��O[���nH(*�b�#��TJ�ѸiO�V�|���Q�Q�,�E ně}��Su��o#���G����@�F��J%-�����E�TJ��#�$��z�����y�zW������������X���UA��7�kC7�֣��U��3HCX_�����U�89'��t�u���PwO��"
��7���^�/���x'Ȫ��:O��N�B�_�D?M&u;�:�^�E�Z�`"6�}�#dm���~�a�?����=Y#_�;��y}L{Q����C�5�XH�C��l+��H/�BJ����6�R������J������a�)���`�ܕ�teE�OwTm�$^_$�m�+ S��:�_�ox���s�@}��#p��	�����}f�AI�ܼF)8����]S#".9շ���j"�������C1��E3�<�l�����{v�弐�������ܱMo�L��n��������Jg2�<1�����k[�r�:{����nY����<�x����Wc�7:��*i�M�����B��ߛ�<�l,�f#������,��e��4��p�4��N�r6�k6{���>5D������^�%�H-�[b��+���h���2M"2��b����(�J�+���N߮T$�j�:Y��'koث���U��HkZ��v�|��ݵ���Ƒ^��.i�A�oa�����߹�1"m��M:�k�� ��Q[r�aH�\{r".L��)+J��-æ�9�%6��``6�3��=����;�tvg.��7A�N ���q���BM��re���D?�|n����HB��6�gu\L��@|,�}�1��%�rC��m��Rd���&3Ku>��%�'%���	�
O����}��[�}@w�3l�x3Ӫ�љ��	���*2����gJU�B�����%$Y	�ĭ��fq��L��.��ӿ�yz���K�������$��G�5^*R�c sieZ;d�g�� ����k�=K`�$��7�9f
@�BY���N��S�kZ��pE'hr�M�] �!�hߺ�7u��]�k �1���4t`I���Y?WX����O蕾v�&4�������ɾ'�q:���]Q��)e�W�(W�꼘��\G�w`�*�w�L�a�^����d\��j��;��X��O(+.����`�����{�xu1Z�#z��GPrK��}�D�3.!�݋&��ׄ�]�{!;q�w�AY�����%�
�hi��_E���]���Q�3��
��`�sl���Ͷk��o������:�������Q������ϼ�|�1{c��TF���T��v=����/u^v���n#��2"c����%��LzK�A7�+#����3G�cg8�vD)��v7�ǎ~�N|�����v�g(\ܿV�i:�q���8A�Ub�z]�@~�dѐ�<�/H��z��CuxǤ5�˷�(����#P����z���q�1�f�p�Ф!?�(鿔q��������}h�p?��Ϙ	N�� ���G}����!_�>���=8� �dDu��$�<�=<{�==��Z��: �E��}'xh�}�]���MP##��#��;Pď�z?u�8���_�έ�,�fx9����@�lrl�j&ć�����^��ھ_3����	=ą;XJj���s�c�K�s*���a�Ms��g#����B.��Ft:&��V���6�$�m�$\t��]�r0�j�Q�Jk��J���J�LyN�F5��<�"w�~cC��7�ZiH�� k[b�Zo����G:�/D�C��Be��L��"���*��i�c͠h[ }���[�2��[��p�l��;^���YXa�U5Y�`���v�r��a��Ӈ��}�F��r"�a/_U�w�ߺC���W���&iu��풉(�pϧ��X��aֺ�}ʡ�:@V]�Eh���η��l�;k](x�Ң��C��\����=�S*t+��n�{�� ��Xi?'���?����eWa��������4��=bY�'���!�hE��s<�-�|����+��!8j�{Q@`���p�A5`��ߞ�(��fO2��LKJBT����z@��=��Rg	�4�d�a�*�n��)�&W�7�����Jg�6��"��q+��'���v��`R �� Et޽|B	o#Nxo����29�K��$�x�;%�&^�@����7��]��e�*<�C�}�
*Ξ��Q�7�jnE���3"�j��3�.Eq�q2�:�]QI���e�I��;�2�I�!���l������V1��q�y=�z��2���
�Iv*pb�7�S�L~n?4d���8�b�7��J�v�qM�U�}/k��*�"IA=`]3�.7	5����E�bZ Z�d��ZhHJ�����L�����ռ]�r�x��Ŋ Ԣ�]�S�̍��Qg@x�y1-?�U%t�ʯ��8���]�֌�I�-*�d��T~q�o��")�r�I]�~.c���,,��%)!�m�;R ��^[5n<�޶bG���'C��\�� �~Ȱ�Oy�k��sK��+���@N���_3͡(f�"0jag7%V�sE��#v��eB˯��~�G��M0� ش�ǽ\��	y[�7ӭM R.:9�`�ZTr�1HG����LՁc�s ]��{��[S]��q�����<u߱�Qg�T��9H�^�i�����/����xٌQG;}͚qv�����J���]2����L�����>&G�PP֘7���2j=4�ԋ�ҷ�H	�*��?̳�����=�G��_Ǐ���y?y�N{����-���}6�w�6�9٭jH;��J�����0e�G��:r�zy�͐���6�\�=����n�0K�G�UzU�2���L�@{3�d���l�R�N���w�u�Cmx��1���W�*�
�K�$�5e0�ش^�E�������e�}�������"����D;�#å�h���1�jY�u�&�.�-�g�f#�z�!��zћ���������ˤ�Ӧ���<A*!R����iY	�M��~��s�C��J�����Ϭ�����Ň�Q�1�G�����;��������1��à����\��1r��L�7u�R��`Vbn�~�a��.�x���;�mo�(����t�%{H`��>~�q�A�]&nT�4N3�� #�pD����Yw��BOQ��u�>��o���>�U:�􀸹k������*�2� �7f��q�~��L������ �>%���w�o�����n����Qu���B�[�S��3����:T��j I�,����8�gg��T����;���̍�AWa�1� ;
h������e��>?�טg9yg⇬.ǹ�*G�]/���~%��UlL}b�����5��ֳ�խ���WG���tҋZ�]{!2���i�[�	ӎh5��se�������.��v���Ʃ8��nn�$��[R�f@lk79�Wy�ث������A$���C�3͍�A(����F�NP?�<��ΒY�����q�~g+X��P9��U���]�w�1ԭ'������f���`�.ָO�6p�PH�U�y%|'�@	�"}��_.7��l��K�Z�9�dĞ�^X�8�Z �� *��y��0]@�H�Ն�ȧ��?#���L��1v�`E�=M�����?�r���r��<M��zWkw�^j8��y!�����[�����+����Xc���ӊ6�aM����&=�l��_���[Z����?�;��D(o��? �)�b�V�z�����	yN�G�%��km����w�@%JǾ�xaOF�;՜U����+��Jv�}�!�g)�]t�������l!3�i2�0vI���8�^ӷ{��Àx�d�Q�4�x�sðl���A���86�Zz>]fP�G�����1��d�ϷKrWO�^J�rϞ�;,����!����Fy�*4�P߲��4�� cV+�0_A�"�e�7J� �Z���o
v��M�i��a�Gf�� ��\��9v^E�6�CHO�M�c�:���ʹ=��
e�]� N�L~�[AP������9&:{XQ��4O3�3�?Om��g��	��u���͈1Z��x�Լ�)��V0I@�VWi0Kݻ�:ѳ;�uYC�D�a��
��I�g['��p9r-\��Z ��Cp��:.H�$�a��_%�eU�+&<��zV�l{"�5�+��x��toYb��'�x��}��KR��y�q��]p5���6.A���X^��@]*Q1$_������>��V�e^ǡ{Ώ$�����/�2�;b��`���^l̤������f������/�܎�ā6�#�X�,x*Q�!$��F�8d�;ݕ�Q�:�q)W�A�K�^�ϱ�'��N7��'Bj��L�y����p��_�D�:�2oQa�S@���G�p��$��EcMB����M�)<C�� ���/֤n#�C��f�����	�~C9�ikJ�}TX�����ԁ�C=���0�J��oq;_�'�L� nn�6��c��$R_�W<�dI��mB[��#���d�����t��&�J���^R�g�qf�ڲB>Hu8��p��)�vv�>�o��^��O�u4�SO�1��,'��W��x��!��a���E���Ss?֡u3�~>���PW"��S��?�Ȼ��F�o�Q�G_l�)��׈7v�M�;�L �!�K�A�t��Q������!b�/�Z�D��tɞtn�솋�>ᵓ௱��Sʋ뇋k����oS&�5�"N�UPғ:��K ��(l�Ε�^l�@`����k��[����F�>�Y��`��7h��vO%��e%��i��#Xl�@M����Z�U��	tM�Q�o:�V�!F�I���4�#��>�;Jo�9��L$�E$]qү��8��ߛ=tV�u�1��hޡ�u�Fn�'P������P��r��䫵�b�2�n�nˮ]%^.�"�1]�bwZP
���f}��R��d� �� " ]~�0{�W$��4�W&�)�a���Qc��� �,{;A{h��\����\kq�q�R%��@`(O(�L�d͓���4�T������g/�'�����\'����-�Y��P�h\�o��7qi�2��s>X�!�Gw��'h۩�m�kF�E�y�A�z�O��`��k\�����)�?} ���4&��������I�7�ܖ�]��g��M_i�?]��Bk��C���Bg��	�}��qm���$̷}��p9�%���'NÇ�	�]ub�ќ�e&��������շ����W�Uv\<�W��B�Bp5�i��@��H1:�� V\M���#&�x�]f#���xg 3����/����Ϫ��I�������s���ug�p���F����\2��K;�F�hc�
9n̔ikh`�\k�*$��됌C��_��֧.�������:�		B��'�M,H&�n<=��9gs�<g@�w,9�v�?x���a`��^�f{T��c���}��[=���s<7/�&���%v1���(s����B8^�d�hoF��<\��y� �jfBy�/_\{�� 	\G���m0[y���ZPj�i�����w�8�
e#wp�W (�
�>~����I��ި[��<gk9LyjX��Ft�_�$���d������Q�Ak��p�F��+"0{�^I֑�q2jT�K&��%�Nt5�I�9�1�kX�̋�2*�;=N6��q{���t��̒�
j��󻷫�R�����M�����j�Z�
q_��F�]~�3��ҳb�U�mM|c[1d�a>�~����ƨ$}~����K�Tl&��x?�#�i �V�	mһK廵��H{Fͯ�}Eh�]pk����HG�y���[�1�pJ��$V������"1C�}�L{�����c�m�}��#�
��I��+��Y9�%E -�e��hh���a�Z0*ҟg%�t�P_��Φ�9�6?Rn��ٞ`��Fm�Dcؚ>��x?��;zeO�F�o����H�CSl���5/꿤$��Ё���������D@�LL�'[�@WB���C�h�ʔ	�A��I��p��6��ؔ2���|�S	Ԗ;h�Gn�LM�� ���Pv�2�CT>�A��,	a�T(��\`kc����aD�Й=�<���&��!����/�X�� k�T�e>���m��x��z�O�u��k���]����0n�nk��xb��[��S��k�J������E�\Æ�]Y��r.��ϵkv�k]?l����~��uQbF�ݦ�%���̑�̀è�9x�,�<�0$GLꏺV0^[x�~�:�.$1&=��X�Q�v�_�A��{nY)�%(.3+q��Zv�e�j �������UO��(p7���ޅn&��g�;s��D�ɔ��$ėNZ3��4\�rȻ��ĜQbսx��"��s;:cM�/T��ɲ�7����
`|g�bp�V��2��b�f2�;ԼYs��:t��(w�\]]�|����v>�WGޏ&�m��ɋ�B*�2%e�tJ}ֺ�#��wN�kCE��R���O�,b6��9���8��gH`�"Ss9^w��x�0b�a�$W�m2��%���ex ߴE��m��Qθ���̺2��v���pWz�|s���|���3����V�IZk-�9�O��ʰ������ �u�����x�P��c�*=���Y���+�<��{�d��~�da.wWd�����o����U}$lt���(���z20��B�
k��}�&c�e��c�ˮ�;
M�5�|%���$}�o�{�©P��4����� >�RR����G2x���{�oN��m�oU�Z0�L�����`��͠�0xz��]qe��X�Ku���uaΡ.p_}�+��!���r13�=(蠟m���:c����x������Y�6�ۚb"9���i�����XU�XZ�1N�"����2�r�N��\����'cY��x�խ'N�'�x��g���lb
-�L�^ Y�b������_�<�:����X�f�[&΄B���_�H�¯��x:���ҲwC�}]U��j%{eu��}�����;�Xc���/� 4T��l��I�a���AZ�dE�|Q�LK����ǩ9P��F�y��(��4�k=p:�-AE�0�kS���+NW����Q�eCy[�qm�JB�Ϥ_�B1g��;F����vt7�7�Gp5t��:�q�c�)4XR6ӄ�\�-�B��*zA,��"р%E���QN]�@��9�����P0-9�rm^%:����/h5�iX�OޢG��R5#2�D�`^��P�Eh��4���^6�Έe�h�q��75JSF���`�����?�|<+�}�g큂����@�o���<��Y����o�w#���%cDڶ0�l��]��7HSj+*v�ML_�2��'�<0b�J���N��V��c�b�k+Jf�@$54�E��)A�S�X�^T��%���E��&8Y�h�e$a��dU2��Y���D9%�9>{偓�M��T����A��p�iaLzM�n��q|��0�{���tο���"rdA/��(����0mj0����;G1�(��Ǒ���p��ɿ估"=<.�ŁV�T@�L�cH�O"��=��޾��gΈ3	��ɍY��Y��n1�T�;�V�k�� 2�;�q4��KK�>�j* ^FˠM�Hz�r��䟜��y�����3�*�0����4�*=�S:��<݈��a����gx�#�\F��f�fђ��8�Wb7���A�B�h����Vi?|`�6%.���͂:R(؉A�3�.�G�ٲ'NMƃ(z���^ӥ�s�7_	�����n������i�t�n��-	 ZB\4U�W,�S��n/���-k� �0ג?��B�-�)�G�����`�Hg�,1>J|�p���w��d:�N�����_��M�X�N2Mo���f��z�ݍ����=�!ƌ.��3�:��a�,�]��������n��\E%�J����^Pz�U�L��ژ=!��(�κ�%j�霒<�(�(���[�D��}҆�Z������t�jWAm`�Twziɏ�T�y�x�Dhf�B�No߸��&y6/�s��j9Eu(�9����Q����2��f�Kv�_�dQ�w��� �È�(]�vI�I1�I�Z��u%��4�����`�F2��SŖt��B���|U�FM�E�XK��k���w ����'*���v������\�̃Nf�(Ǫ�곖HI����
�g�R��Q�iԫ�����OQ��;ʁhv�p�e� � F��l�ŝ�.�N;v�^=X7�� �����n��b�l�DE4�$s�$�-�o�_�2I%�6���#�*+��BU"�[��RZ�
cS(�e�+W�˝�6�|����X�s�������e�9k{e3��J�
���]� y��n���p'�5��� N[�QɮZD��!j�0Q�vr�x�OE��r �8Fا9r�dڹ`����ݽ��O������/&:cdda��]�G#�Vc�G�߃�o�չ�\=y��f���,��0�g��B�]@�s��p�Q�X�&U�-�']�4ٗ�	�܍o�&�F)5�R:�$�BV:6�����b O�W��Q��g�/��N�>��z5w0U����+'
�ūgj���&�[�!��Z��Z/��Sʤ���f�9�ҕ`�FL(GG��?�):_�+�~��|��tw0c�{���+�4�x¸�y� Ruf�h������c�S5k���;�9T�z��_�G�%���,pH�Q�S��Ǵ#����0
�O[UX{%Fy�Rԟ�"�����Ҧ�������d�`J�v���2\��[��̆�����Hp�n�<���$x�\��ypr��FO�i��ɺ�U�{7�f`��<�K�~se�{�v�Yc�#-�������ʎ����R�؊� @���(��Ʉ��Z�4)t���jN���P��gYf��`�}D)��j��!+��OP�LƖAm��1������A�������9��ry���m��|��O"3E��s1٭l�ݹK/)Wڒ���s@����e��&3������4�q���̡�d���;oj�}/�/���+�'}%�����U������pM\16�i�*yx0KڪpHzI��zCۛ�z�C�]?W`V߅�E�/�Q���{�c�)�_I#�o�G����Zɚ�q��His�b�じ��Qe>nц�:��-����\1R#1V� ���l�e���ӻ� ��+
`c��l�RĜ�j�ρ��	�V\����Z����أu�(>3��g�!�g���"�GɌ�3c˴`("X/fl,<a��8 �[�,T�O4S���UǸ�+9&��n�	/���v)C�p�~fa���l�k��	v��I�4��ϐk@$�j�J�4��BmS%�?v�I9t��.��W�F-TK����?0r�U^9C������;��:%ͩ�[%��S��*�h������z���7�`�L't�
j<�F�~�/-ɻ�ԾH-�O��g���������^Yh^,u�="o�)�D߉W7�S��?�I<b5�����K���EZ��,��G���������B0���Q�#���{%:#����)@o�MАĀ{�zc�60��1W�}�Avmr�@����{wE.���_����N�_��&,��c��L��j�Y����H���o�ک�&��dQ�R���Γ�f�Y�!TWnR��7'{���<0�~�-RF�m�����#��DTn�(�I"8�E�}	}[-z#���:�r�d��x�#��,�]wp�8)��Ƿ+��@��Eج�и�eM����8���~����Pza0��5�JXOj��{]y�'/K�`G��M���%2b��Z�"Г:��q�gE[nԏ��D���a;�j���.�\����C����?x�&wr!�@M��)������ϔ�6Է��>�e���i����f~At����)"�t{��Ƙ�\��v������S�h�H�B�~V�o�F)�~�e�+:_�V��_�+5�sѣ�����r�Q}���`�=�}�.g;�����|tB�ǐ-��Y�,{�����	���������Or�/�6����X����c"�T��oL��%;�߸��1{H@�+� ��D���&�:�<���Ή[#^�t���#LT l�أ�>u���E��B�(R���>�#�%;�\|η���Ng�k�R�X�
嵸Бki�`�|��M+�H�ar�y��Z�ہ�wG־9J=lrzk���6A���J��.܍�Vu摂�`&�4L]�{5�M�$|�>XE��Ra}i0��n2��dHx���8�.|/������3��@��H�rvJ��"�8薦E�L�����ijK$�*A{6��g�{ʊ��{���P�k"��UX�ay�ԅ:t������>|1��?[�Dd�p�)�=��;������)��򿹰b5�9T(
{]HKj�+�|S'�ZFW/��|�v�j�4��]"�6{E4�K��+)y��v�����.�1 |�ҕu���$$UF��-����e�F>����X6V/gu��j3�RM�r����|���!�k"epe���nO���S��s�)]h���s����	S<���i�
�����9��$��V��Hq�V鸶T1�A���s8�_ 1���̑��6�����t]���Q��3��6�ґ�SyHl}�b-i��hJ����L���{6����>��K���\(y��Ͻie�KM���U�˜�zҲ����g=�Y�T�L��PQ!�s������w��syR�ì��|����KI�����s��;J�	��*&�+���9ؙ����ie_ݧ�xd�zK{B�u��ҋ֯Un��JYB�R����A#��Q����?�Ef���i��]=Z�17Z�#����QM4co`uǅm��ж��b��}���������A���.����p��(�s�V��/�`k2nڜ�H0�e2T�����9�0K��x@CۊV��lG��rmٲ|%�#�נ�Oq_����0�4����/�9y�&- �������g�lC{��hd=uB8�= ��nF�#������/�	�BD��ݬǛ���.�,��Y��ِU-��?�>�����������q(J.[C�jY�u'3d�Sȱ.�.I&�}�ڄ��T0�UM��*�r�4O�{��p�L�I+'vo�>xڝ�,#�IW�������^���p�p�G�;h���"M��mA[Z�򌃸��{�q|�@��a�����U��Eg���m��{�j`��a)KgV�X���=��׆AZ��q���I�Qan�5�Z�2Z��H�6�d�s&|c)������x?p��{�rV�a�uX���Z0��Ծs͌j+px�SA�:^?��g��h�1�rR�^��KLك��[��߇��sNQ�7��i�K��ٛ^ar�!o���_��E�x�m�A3���G�h��=+�Y�r�6����[_Ge8U~"`L.)V���f�E��X�t�0�A��k�;Y��ּ�����<�v'�*>�f�/�3�{�!�?V��y�6}�NY�`V��Z�T�e�'6�j�I��/��A�K	��o�'�>Dr$���.�:I]X��ͱn��2X3!�T4�D���b���ีEř���%Cڈ
�Q�T��\.�
�����-��Ld`�֞���[i�K1ci��o
t.�2|�U�ܿz�m���<�|@J?%�t{jZ�?5гvӁ���hU8pz{��$B����sĥ�w�Þ`b��6	���c�6QM.�� �q��$\S�۔���.\>��x|�刍��YuȺe $��{?cc�P�@�r@Ș�{��޽�f�^������[��p�T�JTB�Ɋ^h~?xh{C��%�v<V�B1@����U��ňzk
$ML����:Z0,����$M�b^��m�t��a�8�3��`��q&�v�n"7'�]ɔ��4B�V1��j�bvml�p�8�M��Y��C�k�
Z�X�:���N�=F�Xy���b��T]z�~Ӹ�jFoN����g~9�oo3HSl�z\��s����H������i�����TχVo&��y�eF�'x�&	�8
�hX���t��_�͉�ڭ���wb�(q/�
_l��!�
���4��\uUu�k1�rte�{��ZS/(�R6`��*���T�N�|hjY�F��<�RB�jG. FU��-�E���@a_��a2$3��3�Qtۢ 8>��_㜷?��r�O�z%�����f��;�$ 8-�y�L��ۧ�t�Ŭ�;(V*|*�q�@F�*��C�d�m,��Z&ؔ�bnL��D��K���m�?�>%poT�<��EE�&=�¨p���'j�D��m&��f Q�	U9���]G&��f�+�Nڲ��ׂ3���Z��=68�S��&�=����Iw8�,�@z�3�ܺ�:�N�e�:ܱ�Zy�1.�]3>`cwO���i|��6'1�]je��ey���= ���"��-���«���r�ڪ:��X�6[y��V�ޖq���pAf�@.�,� /�.c;���E��|�f7?�w�}�/q#�x3�	ٔ$~r�.�ʲ'ؖ�9{��Ӗ�F,^m��Hۻ��ʀ5�l��μ��q�̫�/Y��4�"�j�dOҍ"�\,�T�0�"�q �*��5k��>X/��/�'2H�g��_��v_>	����IHt�t�����`��c�[Y�&;-��3��n}��H����;Vvo֪��T�0ֲ�67��q|��L\(K�����&(���(wo���������x�)S0�Q}3ŉ\5!lj�w|�[FJg�B�W���Į���L�X��ޏO��sg�U,�
]�ԝ2�(rB�i�mOv��,����8buB��9Q���A9��;�\���@��L���5�
0��J@�@���>�c57�M.Q,��F9�rm5�,8h���:=Ė �<��k�."��g�j�L��g�?���3���c�e�y�YZE��nRҮ�e��V�����P#K�4��#�u5ϐ�u�Ah�	O&U(ʧ���ދ7%��r3꥞�a��K�=���6��	�&.�ֈ�w�J���EҔ�[�.��z��C4/��4�X*X'h��@?k���>�V�h��>�`�ʲX��J���%:�<�
�������X�ɍ�`���e9�ĽS-�@}΅�	�Rr�1�#1O�nf9�<ث�.\�7�4�(۔�	�}%��8���b9<[5ma^�3>����5a�N*P��ͩ_B5˽d�U��h�+��~8����Z�/ �M������y��iy���ʘ���skZy��ۗp8��v��r_#�}��65�#^m�U�"�2��x�%�J��\��U�*9�;����Gp�J�$�B5���&����1V�*�p?G���S��AY���#�
���xnd�0 ���C����5�W���0��"��/�9��+��ˇ��M��y8��Я<�y�2��v�d;|��W?n��qϹ�e�e�~ϝS��wpgi|�pO�n�����0L`���L)�R>:��rًJ1<$�(T�&09�ݕ�]!h�P�P,��?_��`����]܍@4�����ty���s�ݸ��:�7�{�s�(3��5ݓ#o�۴IJ�2\��H�?dv���,E'L��}��͌�[��d�M;*�z����b^ 3�/���:o�Y{Ȃ�=�Ў�5` �VC�dF�Nps{�7��d�?S��<���]I�����@[�
��u-.�N�1��]^�s���ͩ�YTOu��g٦v&[1R��pg�su����]���fK;1Y�{�i���s���)���xB�p�;#��(V�0P�b�]T�-)��|7wb�z]L"<���6�T�@;R��CT��z��j#�Z҅&.�As�E�3r�9zT`����EUGP��N�0�6�8QO<~� ��RQO�T�j�=��mņѩx�K��1eD=ږ��*F%�ô�U��csi�ZY<�Z����9��F��S����.ӏ	q��"�(m�����8RӲ���5!z8��a���� �ؗ^�t���N"�N7��7h��F�~ N�����L�W(M�Kd�v���k[�޷��i�e�	���[����z��U�3%%��dqR6G�!���t��
�k�q.�D�/�����6p`��I�Ն9�05�~�~������>�8�H)+���l��1�H����OM�by�ok�Az�H��f���r�5�^I��"�6��qy�����gH F�"��X��@��$PiɺJ�+@`�4��!��B�Z9@�a�"ŏ7�N�#0r8���
�A8;L�"��7$ƹ������7T���b��k��#��/�$d=�E��ɟ�W�	�BU�kz3��A4�|���vO&`{L�,�h�U�/��Y���S����QYx�<Z8�����\��GSFX�@ނ&���A�6��/>Ǎ�,"�"e+��EN7B�+aL��N,MC%���Z�Kl�o(�!��>ޘs���ʾ=?=^{x��~& X�ܮ�7Yζu����������y� ��Z��q@�м�n��\1��-+��ES��EH�l ��W.)t�һx���%;�7�}7V�&����椢��nP�t7A�#�j��ED�i������؄ǽ"
;�����k��{�]
a{��%18]��6��ZWy^�-'F����x��R���a"�Խ��Ŧ�u��1�B�ۍ>VIp����7�	*�s�-��W�t����������P� ��s ����F5�rKt4���x��eRM��]��b�d�D����f�a�(��.nq�$6�2�����mw ��"�;=�z���Z�w�:>x(Q�����6HO��6hS�j&;FB�T����lm��
��7��JfƆ���M�U��}����}4>z]^�'6��x���fjkCp}/7��|+��� �v����{X�8��_��T(P�������5����HNE���BN��\��w��w��h�B�h�F�s��ah����+Q$������4qūy�q�P���n,iȕ� ˱�vβ|x��(����=?�]�6�=��@³H��ViA��of6� � ���[fTW�ؚ#�bB�x � �N��Ɨ�BЛ0�+K��	�_���K��}2�X�*��/c��ة���t����!�#u��U���yȅ��\�Wc9�F���1�����v Pc�\��T��i�.e�XB��Q��m���݇C	<�&Ux��t�`��>�)�GPfU��F���� �Th$�(T�ݧ��4�t7���$�l�%��5��'�VB���I�)�;�����WH*���0C2����ẏ;@>�崪hn[ȝ.[;�<!�n��􇎼��6��	�����_�:N:�y.�7��\�oA�	�~D\t��,����ؿz`�[�^Easf�F��m_H)�9A�.��T��=Fq�5�*F�J��a�F��#��yi�����#�#�M�l� D��$+�+�̎�R2�����kYd�!O���I��X������������"|��4FʀR�9̝bҶh��E���=ñ�Զ)tA�u�5�+�E`�tI��*lj���ǳg>(�Jᒱ��͚j�؄�\�"�s���JL:���?$�<��a��Q��	8U��Ut�2"�Ha�X����sh;_��'*{�8���\+F��öB[���ܗ�^f����yF?�a����	9�~9��~`���K�C|4��r�u�CQl�~X�t�#���%�hl�*\F�Q��ZXl����tI�������\?T>���'�Ⱦ��.:j����n�-RR����*(�(����|��~8�������]��V=1�&Ta�A�s���ǛS	Б�,��z�b��ۻ�2`�V��:<�qż	k��h��� �x��,�X�[��wMt��:L����F ��<�C����SG�6h��-PJ��
�}b��6�E�'2�'�����akxd�P�Ma��7�_����"������$R
� $z����`K�hF�f�2h�c�h���b�ӏ���K�Yһ�����H��Mc����c%|�V�Ȭ-�������<���v����8r����)!nq�ld/�6}N_IԤ����ó��p��,��D&s�S9J���ڋ't&�w �5z5�,�[���S��J��\b�L��sN1��/L���ʤ�k�mC׆�|-����Xw\�3�:���W���=6g�X�SBP�|�����pfT�%��p�'�Msu�!����lf����������,2�?���Y
Z�z���R���Z!�i<�������q��������
�*����J$Nw�h�~�r�� >y�|� �% �h�<��;:�h`�iJW@�Lπ7�jI��LQ���,3My�>��_�H����c?�$�|XC�ƹ�;?�&N��	�ݤS�繉���-�3>���#|�S���X���	���,���[@����ӣu��V%'jC�7.��R�LH�ǈ)G�xc�7��Ow_���CD�#����`�e&Aj2�s�wKQJ(1��;��~Og�����p����o��I��#~��]#d��JL3�r}vp��)��kp�jfCm^�J�F��>�/��-?��_����<ƪ�}p6(�K����z	�D�}�S�����ۼh�x*�1HkGބ�K�u5]&���j������g��̂ߔ}.�|�,N�F~W�Y�h����e �M�l���z{ ��n�������Ņ���&��?f�)w$���	�r�3���TKv=�C�N�$\
�H �)��,�ŭRC��+�3։y��RM�Q������[@��X���^+=)��%���r>�l��R�.T*�))��~U�P��3[��إ�;f�
4%:�C�F��Q�� ݮ�*�J*�}�$��a�̑�{o�� "?:̥wF/��E�F,`�h3�ݫ&"�7Y<C�VU{{&�t�*�:�9'�5��@��!��@S��?J��1��ٺ2A�:��� ���H�����Ӛ���׋	�"���e��O�0>M$1z��T�>ω��A�����|��V6�⪀�;=��*<ǣ/�'�ڭ�`9V�z�$+��ڶU=[���%���'X�]qD�0�`ݤq�)��R�m�֖�&��x�Gx�+��T��]^�7�(y�xr}7�EYd��q g6��G��yn54��<���7�˟�<��Γ�liM�j퉏jYѐ��?�����g0}�N̗;W�C��x�ʷkc"Іa�bY���3���M���f��X�S�䭿�K�6��Y�x'��~��{a�g^xww���p	�՞�eWV�2*+1ɚ�̹�M=tr�5��ojs�������@��Q�a��Eq�*BO�L����V�ΤQ;��&{�D���p�-�/ dp�S˨���~�;�KrW���G(���r��y�h� Z�s�+�ߕc콻�L��_ߎB 5/��84�1�<t�	_=J�a�~�cB����+z������;s���aqf��$$���*Y�p���͑�`|���ј$s��$�����wp�c��	�z�zBlA��Q����F��W�b�d���;C��dH�ͫ����V�fy��8��=_���7��fD�������Ʈ�>��;���M^§LC���W+�$��O(刧��34c�Ҽ�q���*�u׃z#)���	;Z�M�v�h�V���k宽�@���B�♷����� Z7�����7ρ���8����J+v ���!f#��?^m
���f�ӂ�Fސ�g �Ã�ցw�0
A<��=ܧ�v���gv��m�Nr���A2�����"zh4�;����EM�J�6瓥�q%��@�ۿ�T&�V�W.���c���Ӊ��[y����;�"��iB�������K6�K�擯���q����X����vȯE�Ui�|�DëQ��t��*��X8<��F��I�	�wh�%��[<toセ�	�G��-?\���С}��}�����+b�v�7x�Arc�f�K�҆{�v����-�_�E��͞%�>�7� ��OO��v�����E��(���,���
F�%��8�������34ڔ��j�V6uj�Q�QO�5[���u�O��<Z�o9��Zs_A ��	�)��h��w`���vy�]𹶽�^m��w�q-k����	4�3����B���R��ڤ�A|S��7F����B��HD|hY�=�0&�{������'y��21W)��}qk�s�Ћ}㰎��&�5X��f�s��솶T�K����<w��t�����eth����k-?=����w�47P�ݿ�ke1�e�q�/28�E�K���ъWK�8ᗉ�?���m ����\��Ю)w��aTM}�Gk)���W�^
<��w����f|�C5��R�ɞ�/�;wN3���>k/ˈw/�Fه���Q�o�>6��m��\Ъ�gF�nU��%w#x�~2 ��'��C�\�0�LӋ&���1��ںMI���`I�@oO��C���\��!�ϛ)ז|���LV��b�Dt����kK���X
 a�&b����b�ɢ�ƵE��Ψ�>@��<�cM�2=�o48j��������H'ݸ
�<rX�[T�I�Nێ��}9���v�_�CѾ�����kDY�z=�S̏ci�ɜ4��L����2�P*��)zR(r�c4�"��z�~���5ʯH2�h���yx���l^Z"2c|������!h��M����:3�.Z�
2]�.UiI���Zݶ���n���W�'MD�Q� �I�{ �<�k�n"�+�����۹�Q%��x�;��g*h�'��}ܹpg�0����;>�P���.�6-�y�����&�5��Yb]��`�po�9m11���;�����;�E�����@�0�7��ݿ����q��כ�Uc՗ȧ/�@�jR�|�!��<f��[�-ahn-4�����R��Ha�U����:l�|5$�#o�de� �@��%�<�5�:_L�;�?mz��`2+�`�B��4��~��tx��
�u�fۺWg~ai�s4]X�R��M��TkdB�ȁ�~����ZاL���"))F���:k�Y8{%��h�0dx�$hct1�hkB��Jg\C��|.u?�0�f&"{.��AZ6�lK{�I�[��]Q3�d�`��i��� .��z�k�ɝ(R�{--A���n�2�@�~\'Hʺq�=�ۼ�İ0mt�w�QL�#�����dq��$a(}���p���l�L"�w�Cgz:�D�V
�4��LP���g�����q�:�7;)C��!S���B��Tk�+^�g|=fP%B�dB�s_�Ź��-V�[S���6�o>�O�k�D�x,�A�Ƞ,��������RNA_�\��@&^��+<�C�4!G���\�r}���){�
4 �0 /�a|���L���21A2��g���;�yn�G=��K�4����S�g�3�4�$��4׾_]E!Qߴ�Y��{����$��K���]&�L�����!��_㱪����J.���lD�a���ߍb���������͒Ѵ�44�t틪�֤'`ZV`塇�jFA�z,e`/�^�o�;1AP(��j�Z��R�0t)���2a������;��U� ~=����;a����]q�$eڔ�#�[�01?���H�������������d����z����TD���/�5*rq��-�8�3��ގPξjlE�i@�jHA�J�?togz��5C�YkI���;j���ԩ�v����,�����2u��
$���6��2���g�-�HOF X�U֚�v"��<�{��:z��u��93n�P<���ͬ��&��x@�l��Mj��/�V��i�tD�C*�Yy��؎c!��y?�q��7�3�5Ӻ	&��+�#��X����������:����U���4@�8j�¬�2o��b��o���u�e�Fua�V�0 r�לb�w2U8�;��sBc|��k�>X��0�Ȱ�J��$q�EB��ni5��\�毲@pܮ�Z��MbW~�Z�K/}lw��R�!�W=X�[�z���&fq�韙��u|y��D΀XB�.nԠ�U�|p�h���ͦlU��'kc)g�T����}mC�M6k	��m�9\�H^�R�u�o�����̃W�s�۶';��t�rX�i��ș�>[v/e�bT�j����L�� �Gw��c#θ��|j�7P�,��釽�%I*��=���-�
��<\F���'<�ܚQF̪��?o�\_�J�k_��ή�	''�3 v��������Й�N9��GU�1m��#�?t�~Κ���3��!�W5G]u�f��M��q.2/0Z�eE�ʀH�=@-��EY0�D�~�~�b���2-��������ǒ�F5��.����|y���$��Lw�JeBZ@�ޒ'I">���@�O� ���t�S��~#0�2�+ڝfu��(f%���)XK��wm�o�e3��/���"9{g���H��
�q����u,H��y�a�I�ԚKi����I�D���{������<�<���w;�����i�~͖Vk(�HLg��}\6x�)�1I���d@�|�����
g�*u+��R�Oa�8�'��G��|PU~��#�#�)�l�C�=�5YԗH���n$6��]��Y�1t^g-��l��h応��?�<�UFZx4�l�f�l�R0X8�����;z��k�%J8~c�p�?��=��:����Mn��/$gͤ�CG:�+U� f/B4u�<%+15��_���հ�S��H��3Z|^݀r-�7;cg~P�hw�Y����kƨJ�()יj��~������&�H�E?BWu�@��ū�IS\	�1�>��ω@(��l�]��/���u���e�w�(7�a����qw���:3d��!��>����غ*�@��\�{k�L�=d�nd����˪t>���v0�Y��>�߅���Sx[o��>�m�S�^;@�h�Hm�ҰP�� ��x}z6ukV���^��Lt�S�p��Ϸ��r��2��_h����������"�؋��M>�9[8���y�,��yT���4�y�i�L��˺���!黋L�H��gF1,v'`-����O����������5L�L�ԹWJ��ŗ"���_�g��6��Z��"6���(G�W#�Cwd��{�-a�O�����Ы3RU�w���h�_)K�b{��{�M��ˤ>\J�:|Y�f��O�i��V�Z��zjI[g!���/�J�Pe|u|�,%N���sh}* �U�x~��Y^[`������p��Gd�Vk� �0��\�������r�=íA��t��{t$l�!y�������^��EMr����3����2w-F��ɉhÏ�r�����W���-]���I3��P����O=Ć�y�	�}p���l$�5��MP���nr� 蹌ă��f{�R��ļs�)	K�l�v�8�޵��4�����H�9@L��� �.�fS��)_����9G�1���.j��0�*l-R^P�P���ĺ=��7(��Z��`�N<�Ѽ����QA����N5�1��W��b!(�M��Iw��5�Y��?f������ף��]|}�F�y"��\FN�}G������nu�����n�[do����0�����̽���ul61�J�&Z����:��XΘ���c"7}�W�Q��S]����|j��fp��]�Ѵ�9(���/m�9��o�u�Np8��`�F��#=��X�a�k�a1�P&4w��$wCG�x٥G�S[��<|�,JY�yY�FΠ��Zl�� Ț#^	����!�(���-f&#\�͒�'��m�=���0�#���b������>��[ݭZ��~���^i�����!(��	LA�����"�ǽB@��]H�rC�1iQ
��	�3L2`�@�������0Y	q����t����l�%x������y/���$���\��MV�ש�����<I�[��۞Pi��O�:�"u�ol�祑���"4�m�4�P>BJ =0��:����:�C��q�U&�^q��fL(Jm�g�]�?���qLm�
<Gz�h�������'3�ƪM7�y��R@n�1j�z��!�������f�ؿP�8ah�������D:R^�����r����f����ꍽ{��`�C)'�Z`[-���8���j��#�ۣx�0 L��(_`��T�S99��^��P�-�Ə�����X��q��y;������hjq
�0����bGUI� ��	1 &+�9��dp��
�8�JN�{��z�*�L�NY�ܥ��Z$p�ZHcϜ�X��[��< 8F���L�Cbs���{zB¢���1M��5p�Y�1��x��;1��bj{��u£Fr��\�h+�D�����a�T����h����yQ�!��Ѭ�,���y��v�����f���>g��<H����?c�c%7�N�j�сw�{����&g�=ĽB��'?s������C& 9@�����[�'��d���o�G%�ӌ��\T�6}�C�z��yˎy�e0�n4�,@��uqğ�Z�;=Y^��z�Ekw��A[�����{��d?�Dj���Bs`<wD�|9C��ud�(��\{D��|C�"y��^B�p�'ɞ2H��;���j����X�$یdS����Ӊ{�X��!���=����II�&����_�R�)]BzIBũz>�@�Iċق�R��M���17Vg�Dn�T,���Ǵ�A/;��{�a���H�oP��U�􃺾	]�6�-���F|����oI*Ś�ygf�}:P�C_X2��Mϊ��۾�j3�\�h���
�Z����9���������ܞ��~m�T�cs��F�$}���'��K	i��%�8J�-v��U�I�d����r�j(Ot��x)^yB!������#���c�Ҁbo��ɣ��� ��� �#?#��j�I}E.�f*����>���_�xߕ��"�4�;���='|v��U�ҼGUhH��v�㎎v���bԒ�X����"�o�"Gw�7��ֈ���c�VMݽ�.���\��/{�:)1�Q���ZW����u6�_Y+s�i����&w���%E��pK&����/�C͸.��6U���$ckT��%׼̓��oe��c�E d��o��[�wǬ�J��NV�MCdL=��:��B3�t,��[D}�D̙B��JM}G�]�_};!&��<�u,�{MͣS��>V$��C]���ȥ?�+���y[�',��X���q�>��tV%:&�w��ˆ*^�{ё���D0�~��
��"��[I�;������� B�F��� �����J�����F��{��<p��)\^��mo�����oN��0��	�&��cp� EX\��znv�aLv:4qYvP:�z �h�0�S��T�f��<�2�B���H2Մ���M��b�f���X<�gc>�nUe�'^8:���Q$�,N#�m�#	U�ꝼ0�
��E���C�RG2p��+m�-�?��pg/8���� ����P9p>��{X�-������0�3M�D@W����a3�D�y::G����8���q�{�m[iA6�\K�ξ��op#�ؑ��w�C`�����h.�)>5�)��L�(;z6�S��[v����]h�1�,�5���� De��O/a�Rʯ?lb�8���l�A�"�~qR�Ĭ
?J���R=�>��r0
��e��t �h�J}���{<���_K*|� �W�ʮ�]4��� �QU��C[�G{ �z$r��(e��vc%���Ł=�ף��9�ǹA��A�Pa�f�`��3�}��Y*ڲ<>�]���CX�*f��
J���Ԩ�{
re2L�'uAe}�^����,�Mf�������8��z]��Ʌ&T���$m.��7�逮?�;���U͈V�?ز��o$z����ڭ'�pL��'�Q&te�!��1�
;FJ����:#"w�M)4��Y�����e^��w��\�*Сx����!����'&�^�����Sd��xݣ6���~%�F�J4w�s�B~���
x�@��1����	}�qV"An�}��L
��&	`�̰85�R>}�����y��_FXj\��^$|K�H,
g.)�5�	�BH�tŪ[�h�Y���ݕ��	�P�c�d�4ǔuuSJr��ltDq�!T���y:�O�,����0��N���H����U������t{?��KtS�m�U�*�Ȯpw���j����Ȥ�	�f;��րׅ��G�\e��ek1�X�����B���i�ޚ��Vm�L�������bu��F�r��J�I�He�ù��"�����H0��;�-�NqХj	�]��\5��às��G7V���,&���8m�1h
�y����cJ<Hr3'��wa�������t̻���Ѓ��/����
R.&�~�����DK���D� �8�c�p���0��%���-��[<P�%N��Qy�_֔Fn�KX<�%�4�k�K���Lڊ�(��s���|t��2Ѱ}X�I����忮�f�.�S٫�w.x��d7"��S9��Yz���̱?���$j0N�e�'>� �e�Fs��9��5&-���F�u��Lk�n$b��͐E��{|ſ��@�e�mJ{� ��hYU�0p�s/�����+F�.��;y�N�J�13��
��",�ߣ�[���E�;̒k�_�mT�$�3�8���V�0�%�.w
`�,Z�}')����z��Dg��2��`�5�u����P�7����}K�>§u[0&��Z�×�*�����SPk�%B��[z��#�[��d��
�t�t�ې�߅����a��Q�����6R�B~�8~�ǽo���j=�Ӣ\5U�K�:$�E�{�]
Ȭ�h%ɔ��TY��)�,�O3D�wGd*��b^�G�z6]�AGtS�~��)�9>b'$i����l��V��չʴk�8a�N*7^���S��y�l<k?�Oʍ�\�]�`瘝l�����
�e
n��7;<��|��9װ��3UP.��א�F<�oL/W�4q�G�	�i�e���]^���z��4�,1W�Կ��r����
��9��'F�����N*����p�S����̚;1������i���s4�p�S8g$�y�͔b6]��^�u>�������k
�0%O�y�ӣ���M�m�N�yK w�5-��F~�f��D_-���Y�P����YDTE5���#�����C�'�� ?k�_�c�m�6��6��������;T��&'���c�
��V~$�̖�y��s�u�D`V<~n�<��+̟�K+�o[s�2��&�/�V��E�����V!=�l���yR 3�OW�]���O�iB���D$�$r���W ;��Y�`����Yp�CyLG�}�8���m>{Ek59z�ۚx�����/�\����t��$U�e�N�+��l�TVU��*% ��&_1�(��<�v�ߨ�>�QU�L���r,�`af���<1��:Wv�V;�$Z(�2�6��s[m�R=�((զ��E�����xĄ�G��_H
�Z�.vU��1)�g:%�B��k*�u�

U��\UOq�,�f�H�.�hmI���O��U�Va��u�cr���"PgP���=q� ��T�y�ꛡV��p�|���N_=������0.�Z�f|H @8��F4�:�F�`<�!���U��_:G[,�p�H/LΉѭ�"7>���Wv��M�tNť}�����sg�P�m��-1{g]ʋw�����LJ�i�����>K����V�5���NhdM!P���3ѥ�O[u�sӋAO�|js�������	]T���`]C�S���q�x��G@���e)�`�z��Y�W�6>���Q�l.��\��-�ގ�*)�U9Ժw|��f�IJ\�����D�3���-Ǻ��	*[���.�L냌�z����M!��yMq1��`���/5��>���8 $S����������(u#]�5#�3�g{��㬍����%�VDrS��=�A�?K�����o�]�e���Ѣ��=Ѥ£t���Yı.�4I^R+��k�z{���u��j1�V��>����/��,K(�qD���D&��NEO�Ss��c���f��$4�M?h��,��a���Ѷ-T��Q�EU���n5�@��p�#��V�	&�G�	�Z�HVl�oq%���U����8��~ZьG���wn�6�5ޯF8+��K��N�D)MB0�>��ՄpM�s��wDv��S�s!��tN�L�V�f������y�/�C�F�i,�5xG(���rms�v1q��H?T��/>�z�k�ՋeJ@|��Нi���Ҋ{�A�#�WE1�9�`d��'�~�g�����U�l��H���ZP��o�	��� /�����Q��e{�W�|s2������4�'���b4:� ����n�
0V/�1~��9,":�c��[=C������uj�]��2�(
[�Y*�Q��$�J�|`���dx�݀�u�̻3t[�Bw2��L`���u�s����n�YN	2u.���T�Y���� ��F�/[<���)��<� �=�*����%n/����<��S�s�Q����YU�=P��~�V��yYj'������@����p�Z���s�WX��	�猬H!ڋ��c�����P�~��M(��/.���&Z��t��bXR�Q/A8�+U��<��3��k����j%.�{�^�(����*��<.JE�S;;���r�z�V_ݹNc�s��l�\l)��i�~r��B�8'����A���i�G����;�׌�çpz�)�qg��s�$��Ɨ����$ަk�ͬ���]�#p4�8;J�BF�����$�y=�tC:�J����p����k��&#����1���� Q���55��]O�C�����V�����j஌�����]����Y������"�1Vv\<�}���&0�"9��������7�V�4q��7.�!0F�?�C���]��_���,���"qs����hm�
����\��<B�t�����?��E�W)Gzj���+GGٶ��ܼ!Y �8�B�]ѣ�1���m��5Î�˳@�:T��u��Ŧ����LGG�����O}6�#�<D��i�ev��ok�S����PP�<�Op�o��t���匓n�]@��K�z���h���~W�]��)A�)m���}0�d}A�KX�V�Y�ٝ��%��EKbP^Z��ԯ��H\��xz!3��Q�k.�;m��Oķu�
���Fۡ��)#ΝE�䌚�?�:'�kp��zF���"X`هؕ�V4<4R3��s��,����1�.��T"���	�!�����Ͽ4�Ok�sN<�����#�ǎJ���:��E���m@1��c�����}������^���n9s�-wby2�	�6��N�Z�����6��C*��i��E�r���q-��=W�'���������Oȏ�N.���	%���w����X��{JQ-���:R|�eZ�,�NP�B[�@�yQ��B���u�Y�qˡ#u�e�-�"�2������2I`q�G=@���^��R�A��.	��gF���_K���ɸ���g�Z���y*��Z���L4�~~Ŝ��v���Q��(�vH0�V(������2J�z��g|��� �V�y*����?9q���r2ލ�vkَ\�o�Y�q�^P$�<0zN�D]�V�G@�oa~ĸ%d�h⦰r��w�N�LM�`Fɇ�qU��ҵD�ל��`j�)��
���]����rY�%�T �Ts��Ė�mόk[^�O�!�r�x\���=�c:���Yj�q��O�|3k�˸���G�e#Γ�� n�k�ߗ!�tV�C=9�6=Lj�����(��K�r�y���V�K��^ޒ�[�[%ƈb@�6�� �[�o	J����n>�Z�GY��8U/|p�����
�1.�2������_ƕA�uW�%����fY-P/�+&��q�)�%=��O^���k�}����\�c?��T]r��0����0��� �]��Ƙ�3��?�'5:N1Ѓ�����nM�����U=�����*�s}�ǬB�[�5�s�_Lb@	X�TA
�گ�7��<Җe)mr���z/G�����O3�/���|9M���BU���sJ'�{Fy�!�x�49�GB��r���Y���{���M"3!z
�3I��t#-��l=��m��K}�\"y-��z��O}� c�'Ð�┩[�jH���s,�^��\�R�ǥ��`��_؋�U�V�m+��^��#�f��z����V�:��͌�,��[���#O��.�)`��݀��G���`	�����	��KA��[�i�0�W _>��O���ֵ�ȃ8�s��xBmn"�IZ$,�rU�����ܺՎ-�uu�*vjK�VG_c�ǒ\t����ysj�����>IG�� �d�u,L�O���_�A�v�)�o��|4ӜR��.vu��[Y��4��1�{�4E(:���� M�(��P��3�g�9���6���G����E��$�J ���#�I��\ȗ۹��hY=Օ��H�r���J�o�����]7%'s�^7<tG�� &e �L��f���*�%~��	��8xz���&�a�S抃p�3ip2��ζ���;����,{��7}��"�h��v���d�p��1�Q��v+�V�O�A���Rr~�=YŇ����7�b�Ȑ�[ւ�B�7u��I�o��� n��ߵ1)�3�^0NcC�݁L|Z���6/x=h�j�>s�)$:��7B��*��(�Hha"�I3������ �	�;K��=s~��o��á��� �Z�o���c/��������5��Sb�{���s�Y�rk�:3U��Q�����"��	2�Zr%G6+SE	�Ew���	b��@7f�q��S�r�N(.�q�mab�O�p�5��Y4Bc ��;��)'pL�:
k���^�G;���)J��e�{�a��x�_�L�pԖ�ig�������|0�Ԗ�|T�h�2}%:/�# �ؐC�Nh/����-��P��P��ę�V�T�s�&H����5�R���~f���\� ��NQ�rj��giF	��;;v"��==l�<V���@pA�:D{�gh�8̵���py��g)?�ĝ�,m�#�۬�Gʣ���e�pG	O��x26̻2;1)���:�B�0iI����Vy�d�쯓 �o ߄��N3��Tp|�X����S�J������wk0����N��RD���1�Dr�
���94K �A&y�Wi�P5���#����,���X��\ZC�6&��JSo�����ɰ��z��4�R&���2|ا��z�.%]b����T�!��&��M�~�<7r�^��SC�>���3H�%Doh�W8C���ic�D�z�S�>��.�<8��M A�z�.�}O!�&a�ZD�;�5Jf ���,�xI6���B�l1�ݨ��}F�R!��c�&c����a��W���Q�+:�`�io ��y_F� �$���� ̑�L%<?�GH��\)֙����zg�3m�*б�E U,I;�䓛q�(��-C�����^�.��C^��׾����a^R�~@I�ЉR���*z��Ӓ
r�.����H�
Y!\'���:��'�j�|��H�&u���A*Ec��L
��<W|b�>1�a')k��m(��C�o4+�C6��C�V����{�@��[�_�^�s*|�"F�k����@�r)f���J��~��>�1 a������>���M���� ���fg�U�t�_15��0#�⵱�E:O!X�'&ꀷ����%i�����#�H&�	�&��Gԡ�.PY���8fTŪ�T� ���ͅukx�N�^:b�OF�Zε�5Z�@�8)q��y��?���3$�_�b�	A,W�F��p��-[���^�V��أʖ=oU�=�'i&e�r�
�kt�(��|�T:����nw��=�i�@Ov�������"q�G/v>��wH�J*��)��@����y`K�3�E�؂����o����vl*�/�-iA��J�(^1��% �΍���s�	�6pRw?�x;O�L�Vh ��)�3��g�:"�E7��1���Iu��Q�T\�M�w��&�PNxߴP�]O�VO)�֌O /�����'�fZ7h�u𷾦�w�O���G*�1�o{�x3�
�$�ڵ�$�Ln���+����W,
�t�-{?���Z�"}h�>����G��u"L赕���dfO�D�"���
^S	6yA�<�+�΁��}�p��7G�X���qŢ�oUz�mP-To�ޘ����_{'�b���Z�e,!Hv��#f%�| �7J���&_�4��p��+g-�ڛHF֔�p�e�I��x#�t����:�������^��3�����a��I"y�ǴQ��o]]�wd\�1�o7B4W�H�:l=��cZ��a���+��?���;�u(���j�4x�Oχ�/[벩˵KLhY	���������D���� 	
��.�������Y�pE�8zI��8]������r�1
)�-������r�������c���5���k���~�"�-��ϡMe�X�I
Q�8����*�9�70�����r��M�d�P|#�z���f9��Gj�k�5��Wrsd�5|{ߔ�]^i%�7����m��S�*��Q�}�RO#߈��l��,E�A>�i6�u��n3T�˲�mo��L���,�f��0<�F��'�>��]C�鬍��NF� ���Si�6�}	J����Sa��J')z�[w�~�ӱ˺���V�񯛿P�vn��z� /˴�X��F��� @&AL�:�����;D[���yo�p���:�nƒ�qq"1D��ʝ~��8���I��7��9����e�):":I��2��7fKf���@!W�s����@�(��T{�oV9X�㾀��}?���2����:P���4O?y'3��&�j�����Z�����
���$$��
�����6���i���)�Ї�
����{���
+��Z�8PQinM����2JEȄ����R�'J��/J�nN�G��RS[�< )/�^�]w>e\v0�,�s�ܠв	�F������!YbP��N�*�,�1a�r\5�a��n�A�$ '�hހ���$vG�(r��~wk���Y�qd	�#����zi��V]��f��_7�� _���U6ֳ�D�pQ`/��yջȔ_����kv����`>���E�賂�l��!KV�|�Q��H��'��W�ȏ��:�1i��Hs ���B�y��7W]����+-�ё=:�C�{G����F��L4 ?0�miM$#�&;J�˴pR�9MY�������!�roBcj�20�3��!�}<\���B1Q9-�e���ys������~K��	p(U���"Û�n�*S��Da�I���(�9.�Lw��'(�}��e9[C�jǛR	�BL�=T�4y���1�{:����Z�l��[,_�ɝ=ϔ��Cc����%���<�C���vR��xp��0cҎ�Y�g	��^6����,9Eε�i���M�~)9�L��i��� 1p�Č�=���M��|��s�C��3C��硑��%-��w��8�b$#�_ځa�)�G�VV�2eZ���Hz;��%#�5UԬh�tq?j��4��	�\]��]X�!�)�k� ��w(cl����׮�$ ����K�������#���I� �>f#��#�nQ�6����Pb/��HX�sϓ�(��UlP��S�B��B��Jx{��		N�����䡄��D�5��+�P<��R o�Y=�l����������������.{�Oɕ��|d��զ� U`��6�����O5G} ^�7d�\�K�7���)�z�}��>������ݬ�_�M�#TG���j_`����J�R���*ٹ��|?�}��8��/0��[���	��B��g�Q�+X�i���Zט�R��Ӽ�9'U씕���!��1c��]C��qD�>�"�f�n
o4�(O�ض,M7|��&��!oJ�[J[<[��2�Nq*�8R
8p�3+IM��C,��eď����]>a+��������R���~b$�G6ңQ�PUb;@h4!)ZQ�_��n%�D��.K���ʯ"��_qI҈��>�s�*eҪ�a�r��Ȳ�f�����|�bYC�"�4S@�򱏇�����5K���X^ǅRb�|?N�d��
Ҩ����^�F��4��#��0!p����.��_l�k�w�p-<jͤ&� ln�Y��ʡ��r�\��c�!5�q<E�����X�*[�@��F����#���<o�4���m�ZҴ� ���&w�6�%l��Q��)E4/�âk/S�3�t�S���`��W�x4��b���C��J��X'%݂�Y�{�����t��� ���M�t��`
���x����eg|dk��bIz=I�U�����~,�Lwb��O��bXhpBƃ}��.s:Z}��:e���IS� ����*rImy�-�	�[�g���,�0�&������[�`r=���LU�$�FK/�V��Ȱґo����7^��Wް��d�EB�~��ÿ�ɒ����b�p�wOk�S�Ԍ�o�f������Î��w��5��t`2�3�Hꇱ"�����zǎ �st7�OI ɗ�Rl��E�^W�x��P���8u[����#<��W�mi�T��`�O:lPZRE[u�Ϩ�����^wo���l���Act�?'��b�©̟��vږ���c��I@Ѽ���e�q#uvѽ�'6�.(���K-�{�������Q���ߗ0���|���^�+���T�Z�M����(
����bB�Ƞ�D���F�6|����%ѷ�����y�
��'Gt�b>�<����f��g����mXm<��3c� 7���a���; �S��E�~$�I�P�e�"�n�����d�t����)����/4��!K�Y�z������TIqN�$�q~���5���Jӓ(����f���mH�_2�)WP�߫��qL﷙s��;����·i��$�1-������	W\�O�7�yظU���>��Q���0螯:g,F[x�:���mb�=��������:p5���C?��:��g@��[���U~��uF.ޖ	���d#��O���J[4	"��v�Q���O�gy�e�Cu����0�	:��/
��{ F�g�������(�.�Œd��nl1���q�Nd�ᱷ���NV�"��{&ۛ�xI�S��^�
��۝�-�`��/��@����@�5�?;���;Qmh4�^��2�q��x��,&�k[�`"Q�����uR���֚@���M䔺�)�����[��[�	��P5vwE#ۥ����#��V�g��(�ځ�8����0�aA����Ϸ�0���8]�jg��Y���d+EfE�����윋������D#H�RW2�"C�ћ�Y�D~�q��"0�:�)���6������B22��
��r��@иS1�0v��� ��=��ٱ���T�·hs��j?��2	�ԉH�����F]p��pp;�����"