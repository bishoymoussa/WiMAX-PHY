-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
1Yd4srlrxHQUsIHEyBfbxOiBv414L9ScSHXeUk6LqIS3O986nGJlRoCsZs2AjbbEc1S8fpEBaOMI
0OnlT7t2vQFmJf/gBFFXDGrJ0gKaTNPC6MoDwajWC/x3IwIblWbob5l0NGrigiSe+fWAgDd2w+Gj
pptiYfdd8NXqLdHjyNS2f9rki7D9NrcEiLtdeMP/wVOovLrQuGZbwZA8JTwgIRtpIYFOfecuGi+g
Ue+vjZDuug6DCX1uyF0SKq1Wgqn7udN6rNj4LULK/+5r+FzMsX9nc0OmUYQ7Z9di9Hn8LOzmfLBY
FvXPv3HgQkxNDUVvtVj0iN82REEDwLZJjbhA5w==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 12960)
`protect data_block
f+Mt9CEhMVhHFptP2vF6YG1kT0bexJ+IEGCXBHYyItr13VWuLzXN5VwtuiFHIV4/VmjaOOD4bCt7
/TTtz9NdaByL5RPztsP5ijxccSqC18RGB8+oFU5qJY8i3w7s7f3JWqwx9gCcZjpZZvfLJWGWpSpk
7751Egmnm84SCdhN8cRphUrDdpNZLGyGSNEvI+zfpAJT8GE2hUCU3Mk/t1dEoKc/aDpaL0xdMQwo
B4KBNwVd4ZH1Bv0rh5sgxFMnf0d7JTbUhSFXmeRDJrRB9kndkNNc3BlOfdrK2hJnE+Y9WM8TmGbi
5xuScf/esE3nMLwmkZgFLZ2dGuMkrRb408LJYwIjXBDjImhSk7NHb8AZVH+I1xv3ZOAo5rS+e3C5
m/p1Yf/KCgtAkldi52a52T7L3Xn6UYHgSw673/aoFCP+fk0Tx/gBID94/kCsIIFNnSjfUi+BcQ7E
kLMGKNEBUN9xSYDY1Ce6h220TiG30jYigaZqc5I1uQOYH5vLW4b+6uYLQX7GGPbC6IWIq0o6Fdev
bQQAz2gy/B/pq/V7RrafISBkjbIPOK2IO6MeHf/aDbgdmbw4BmGdgh2GXPuAeQf/STksbfxHuFqi
J1uozUka/lsNKaezslZLaxNPc5FlP8IrLf+r3MX047/IB8+fiehUOohxCg++pXr8iXN+snKNbgPc
13A3uw7yQepJh7g0eWSgrXY4LdyVKCUzzS/PNHI4DvErXxPu5PeqcRsOlP1rvvLKofXnfaPoy7sE
2Au/cAI1XGOPje0p9pWjkLhSYMCvaABUMWu6xo8owT1gYCgfZJZcOj5AxlTDt30G9juxs3n39yj5
lSsrqwDegp/eaPZGd93dVy5arM1f9wKZj/4IR/UlvHaTyQM9nyXlJqGebey9SvWnQ3aI/+maA0X7
iyqzD4POXCxUZDokKP+65SHKdeKzTvdyFxJOlRHPngnSxS8B6AVKs/1rAJGVhYZ1xm22klD/ikTj
dbTZeMRDbv6esHOlmFr5eEDAR3gNr1tn9dUfCBIWQOegTkyAHqo4PNt3R6GksoktWOMZ/5ePwtCn
+S91yjjXRbGeqKaS96z4i03kFY/bJY4ZeBHbgar/vaJLX/r6L63TF7mkQ8h85kIfxdPtjVv59PEF
WG2YCYoc5pYOQY6OkgVE3sNE8u0/Dniw5vrBQ/qO7N+BGKdQ48ZbYCEMyGV4PkX2DZl7ztwE35V+
0D9klnVoNge528hmPxZ5sXpqLxPZcxLklLlLusdP8kLubSAp0jGYx+0fDs8ReS8sGhFBOgkhNX0z
HrYLZ+qdr2l6elxFrueJLKcnpuXIlk/pMRw88L/OIe9WvzwxSOr7qs+L7jFcFPe2ajHfYWbkCJgy
5PZzsa0gbWZa1w0AGIvPAi5/8+o//ifw3SvNbLWgcaLAauX4lwiEg1J6VC7gHaJNrLhUm+YORrwa
3Ifg7+pnFQP6HeyftMcyRfKiMp65uuGr79SACon9Jqz6jViIr8XxgrQBf5LnwubL/pZWQ5gov62H
nsfrQkQfKoEueu0IcqTz7m+o7TFlr1NVW5tBVn64DwTps45rwuDbISzddInmFrFJUwuLdieJtNmL
I1SOtELQ5Nce/vTXNZaB6AtMvpisnqToTpQmFdHyneJsCUKghe1xMtX0ziU8cKJpYLZZM3ZlMs0v
0CzpYHCPSpPW80PTN26Tfl/QgQ4bn2bf+okzFLuzvASej5du60ORg7azVRW56Xlr3Dx5BGynBt+H
DBqMcwuNs3hRCnyqbgEM7eIysXU8utfCF5KAkYCkPP/5UnIV//ypUrf1hgbpVGIKmSBwHK/uMKQ2
bmYLof3UH+yIt/siWvao9H4zjcqROLSGmz2fXuwABYudo104wG1HvRAxbk+ZWWdV1bT53/wi7jmW
oO4fhQUg7C3+cjqFo+tZzszVUHgMs27Vl0b6Gmgq2pe+VZb6NiZ3iAxzZPnRdYB5U4l6b+ZrwOOp
WgRBUgyxzjK4mJFeXCAiX72KCCw8K+YDaWrX3MTZ99g/J1WDx2E5So8iWR+T5np7ES7ICA8sbdgw
K5fYurDDtDDJ9yvfAvyI2Avh2GUnbDE4CErQe1iAXN4snZXAbcXrslyCaeAq1N5zRZz5w7cmu6/a
Nvzn7gmBXmlvWxj9vFUZ8CLuHutMHa48MjO7ymAzm3OOHjjs9Usr2DhrsOjjBL+OK1dDKcB2RaNd
xpJh/BRF+rksWLVysWrN3wyUFiDjCfcKmyncguT+znkj84WGC/LZabwUECQKiMHGnKM/Mic6mT9U
iOMgjflb3/uaz7pBLO/3QUFoNgu7hHvos1ciMynac5mqKWZ2yiSXANJ8wBD7mLLtFbX/vCQG+rMo
P122gDh7Grp/yGWbrv3wdO76tnTohYEBqZeIeAu0teK+8F9xx3kMEGQsOQ1DXBLCgV4Q9l7ncjUj
+su0Gyp77Z/A66B7LLdDcq/N4wt3mtvj/MtK5u4kZqw/DPNw/3voeNL7A95ngBAlkdVo9j9n/C2e
uH9XGNhdHeuan0Zp8h6FAsfC9K1CW5tNawdjEy84TJnRSzT4rqYPwlXdPXFn5+18HVTEKZDl/cqp
k8ep9ML2wMJAtW0Ej17k8xiAbVhJlA46XWeBChUXvQQ4+GZHaqIH/LvFnxiwVltO3vXjkHO6j71r
0bkj+YNYfQCZPgbFaTIQHpMPz2IDAmhE83yJYqILng8R3M9bGDePpbEfLqcJ6pgmNFWJdobOB/0/
7zgADdtA9FdIx7U5nIyaGhqdWZLYTy3aRlNgObA8cVMO0NzB5d0jpxSrXSxZus2eB8MDhjXrr6wO
mAr7dwmPngDwXDNDeHXx/NvzAdcFazKhg+8fXBxPYUhch5KMcTLIyiiA6P+chdo7XpoDq2iFd9Gu
eSZPOTQBcZdreUJPjvzokQEtHZ3kqytmsCJ0cwI1z2bxk+bVhHm0IWZVbcgnQrnHr8wAsKTD1Tny
HLn16FJexox9ej1SgMeZVaHrRKoPBrKq9XbkGlsmKb7oHZ03LddDzaV7B3NJ19ctlFLbOX4woR4w
fwOaVf6rdq0v+EOIk2oOmlOG8rS90tRKZ+yDHMjGiKXxTrzoKnsvn3GZpgv+lTBd6wtYv1XYZM2D
NVcblkO66v/Iy4yPY/yVKlrK9iOh0NyiX4zmCYqqvfhZtdVQPymiV22wu92Os5JhutDk5JgOZ34g
Fit1nMf4Z580HQ9gjXU3PEA/m1++TINzkcjuahxJ50WNagZLtFQu6KkROSX7BELyU6P/8Prp660A
Vk2DnhbMAcXoMwDL5axPZF+2l0P89OxBl008niiafZzln7/553tqaNa4ITXpmsMqBH4BjR6h9iVV
+UvOb3KYBfKylVgzbt7c0FDKhSZ3ZkJ8orWNA9hJIMXfymEG6dFnRPBPOa56zmKvNqq3z1vFJRWE
DBk35V0h6MLhMyMkApzi+C0wyZWHCXgC8BmlWVkfmNfaD5xi833jQplKMzhOfI/ubxLDZmqUJ/nV
yAkQZg5Hri6k16uPv0ppD+Ag18o6L4dY2TFS0MHgLRmjjkIHLWS3JOlHDA4Amb+6ypsMajfjV55a
0SnoFZDZzwFulKMCozIZw1+9+00w1m0QnG4adXZMEPtfs1l8zFQnqCMZp0h/Ae+CEP7k7XaYjK52
piTN4gW6X7GVEsew1XX3SSI4i720xHFulpGERi62B7W9dUtby0OpDP8db1Nx5QZr+7tbg7s2ecSd
P39/GI1HL0PuzKwWyFoGX95MvvSQPS6Z4b7/pL9d3tJdO4iO02p4mnyOHB6MJ0xIkqUsT4LlHQR/
B2I7sC2Fm+4lIBrn2EkHGj+hoYA6XyFVUao0ATDJiwyn6q+UmOglACr3/gl1CgikdhfBcwTRQ1Vf
bk01u5FHnII9JYDYp5VCC+qVyfdyul+/ZaArOthn7gZSiPAQXgwnU3ifTQWJjVHnaR7uM+ZZzAWP
QdstHwQyQD3+trIj6/CvddWPYHE4yjDzY07R8iJuFv79RebKCO+Oxg5LQrzoZBM29YfaIJ6x5JC3
u6PTfzhWpsBlydwYxtPT6pXJCj0TmJ2TntjmpWcxDP2eQ/gWcx0tKzO+qSqHhHU1idVep0yzGgdL
vOPB2bX0lTkCioDfufEolfdPOlOdf2o05UzPyoEAqWD1kj4kso6SxZVJb9QRST3Rvo9F1cm5wlie
AjXzzMzg/FLknWm3euCF6PiI0lPbpMtoxEu+fX6rz0okbwHBbYi9c0Qp1jivJRs6XHqVF+xV0YSa
yWPsRfHbvyez0JcBWLcGNAuJBkc4WLfZqbYdV5vdNeMJ3iBHD5IIj0yodJGTzVatZ4yiQz//PHaa
2WvCSM21w/5mWL9auOo2arjMesn32jfvrcy71dUNzYeDuK0zsSeaeuiX60njvQm7hQvN4faoxm9m
t9JnhVPdYVjA9p4sJZN3FEau+/JDvkFOAuahjupvUjiu9WW5PYFjJ/qUUEPk0uFISE9cEf3Ui2v/
DzC8I4CmmXqh/D+3VsRzLSsesjrR5U2GVggaek+wvdDBM/gaOeYvwc999Xjp3qI3zmVegEuK+Dhr
NGN2D63XJxKK0mSWeLbSr+gCO6KUq4mSA6pvzs6i0ZZ1tH5e7Sr7pMNpnnxfdi0/QbcrjmOx4ptf
BMfpKKAxzLQPLr2If8k0ZOigyqsFHntiaVysYXg0PlfOorvqOCLA+LBNWg29g9rUJHn5s38NXXh+
mNuBoLMTvBYae7LNeYjtx4Dne0eplWkl/yijlXmJ+VvnCJT/nIllcJ8F3f1fuM1G59WQSbmAw/7P
DMNX9wbWLbDuNPgi8JPOvIzG5q8HAxoCpyMSs40bG0F5Xe2Y8v73x51kQ/knTaFxswebUPEv49fm
xXck6FBkerqC4IaCB56ItbE2nfvsG56n/6x+NcwjAQpLX6/bjeNWm5h7WHiTaVIAz3beEYL64ufk
uyL3hFWajDxJAN7Cjy+IC29lSLM72oeGWjestdc+RxhKAFscOnYwo7juImIOs23UC6EwMwWM26ZL
Y/gh5IUBZqD/mdP1rEF2uj8QWxtD0QL1MaZscW5w7+k8MSEStXQMcns3Wpe0hGxGPc49GB/ulHCd
lWiJvuzFrFu8iB8GNGcDMv7qgNw+HwJeCJ9+A+2awf/t2EMh+ZwnS9A5UhrfwYYcG6/BuPEAz0c+
hS2XxkZ7Dbn2nxoiaqGVDvjjzehRSaw+qfKm+4IKwtf7HFs7L+ak1/oYxtJklBUdE7TZsTXMeIOk
E7SyPwqUD0xx0qEPkG6k6gi8CF+80NcbfoitmxBDClQ0g1+pP4+LUTDNM2EfPA0esk3NQPYs2CsU
sugW+VfzbjnCRUJuac2LrfUoO4XiBwIPKLr8f5oYj96xsiL5ofy2SCLkbw43zQ3bXN7pSZMQHGdc
IlKpo2nwMznQ08E3tINZTYNMb1sXFgufOkAfEziiJUV387pCZPr23btvB1bQN/Qd1JQ/jvAXKX+p
/juFNG3iGAB5E1kEW8CUeIaGYYmUT7q+fDEO8j31d8M0kfXUjl+EDVFvQB3uT7hLoC/UiKGIkV+2
6Vt7MUQ+9VOkbZXvnB2+Ydm3MGGpzgMa8cL//fRdG1Xr1YdPOlsIc47S4wU7jBbEbpm+idvfPj4q
ASTP5tn+r33ZOwrb4dMrE7GWs9L6o7C0rCegWT+uT6LKH83PA10IMrlsBjEBy8CL8I3AKxzrsbA2
eQEo5TwLJ8WHwwvDa/DhTowZj9dayh9wQN5ua9U0hZXY1YLbIb4Xp83/w27qoXIKT8zMi5jPOiHK
QbNFk1mDuh8X0BIw6hA31X/D4bPKRfemV8AqY2R3Pk3qWYOs9KOHZuGS1bQMmAm4R/XoM1lA1X6h
l6L5EE0hFbGn5tpWYj0mqrDdS+goJlxsbElQl+UIaExjsg58NlKiwt+KWw72K03kqb8hlcbJnlQm
zRkEKETDEseRFRobewo8MM5O+7hJtKlSteErPu53xIVv4pfnJNWd0Y70pvlllMbUeVuMFKBe4FJi
l94KITiSXona5Np0teaMuSjSy4x0Xs0YS8HtzFpOz4B3oBqgf6KS53T8f0eRmXkR20+BBRZgxN3s
LDuao6u2FG3hTJ323QaqUn5/nwriw7T8zR47BTWhuvOdOIG64SJLjsRvcI0/5RQScHfmXKTHUta0
td6u5p/yp7uY1v/Gb26z8g+MVSqkpomuvaSQmJudxn0LrFYtCOLOB7dqXGshO6xPoov5cZkyHO8G
nHyLMhR0osxmWpcEVEU0oSBwkxFglGeBMvITDsgJmg872HxX5VWAYday8Nn2TlMMgCy+aUNVRs52
IaJzyE/ZS6YMTmZJRm+BffeNtgFXebD1jYOcyADyCjPbikSmVE8CZzYM9YYsCY55pqpdwt/C6za7
wwBldYoMxduxRrmv7BqcKPlF1aPm0k5khp5geY7a3Sa7uPa6MwdR5nesgmP5Az7t55MonuO5OJ86
vcoO5TZDG6+CjYEQRrGy0VBHi5BZQdquWnpjBU8uXzNGIcHvmt85kZ0Olyb/cm4wMCXp5pJbt9QA
Unll/oMDIi9VFKP2IJU5uQy8RrYe6kwieZsMF/lt4ryvnczprbh4gWENS5KACLnDzRzqB/KQgwO2
u1NDZWEEC2Xssxi5Q+6x4u+YhQ4H4dg5azakjJ/4HbtRPuC2nsOVlk9hGlBe9qDJhRXeazHQCIuB
Y9gz7cQeBiwHWvgKQsEFe36fYOAecWuvem+7kZO7zilbW890Q9J6YJ5bGNUQAUXV814ApaQNfcz2
txpQyqqcfdIMANAWNVxRPJMI/pbswImbGiBsjC8yCkYXJPgni5GOeFYhPEZKjsmYK5o1TXcFHZ13
5g1qVVR0Wge5RNx3+jEjYvnF7rYfdo33hwP9F63lMYYOf3kkrm5cgKJQsfIrC/7wM/hCsjDYaB4Q
BQLcOl6/eEy9KkeiQH/cWKCvpXCHP1o6Ndys6f7RWbhNpSOsRDoBfKTGgQ7Fx6Zc2IWloZ5slZ3I
B0GR/EdIDQSMBvttb8m/jJSrySOMErpFmdus9OH+yC4hWJDWQkGRLMYxVlfpAgoJcADZEeRYUwhK
Ap1Wah+BfgTkkIY7l/ODZKKSSWEnl5DJaC/gYdutytPEcIHLwlfL2jeESFvmbMoJixtCRRj8Jy/d
5NE+WSrAZvw4yC4WiskwenX8oH2NrkaUyflKCBTzsMH2NXWv14vKHkuETiYEVwImWhjK26e6ETL0
f956mSTzIAouLTzPs1E9n7X0Gd7ZKPt3Q/4gj/j48Q18Qq8rHeoVJBPYqQFA5Dwj+ik5VDf9nley
NTApjuQrxTmN8v2MlVimokRhKYDr5HogWcP30KxasSKsQzVMANNM+cC1onnsaHt2Vgdup7bGr/fs
3GR5eMlRKcadkcHVrP05rvZO1jOZdsimlavL5ivojxDkQxd2gvjn4hRN7NRTWKza9QFeU4KeoBbM
jgdvdgNJm0bmArunvoE/JsuONDg8AisOoNc0pPZDQAibaPKE6MCTUOd/iqzePssVUIUfpOEpGCkX
nnjHzwVpDuuWJQUgT75Cz17ukdKgIZwi764wI8vlRMJlddEy80cR9I58IhaDylzXcedqphYI7US3
lhoTtTHFQOP7/eE5a6jyTtuWthr8U4UTM4BGbpAJgdB3Qx1k09f2vepdjT8dzmKLgs2XhWc2/SlP
57r0HfMYBXtqzBmmxK/4Be/JLBvi1xLE7p2LOaJoDndflC2pjPPOa7SaHGSJ8gHhwrNmljAMv4uP
i4sEt4qHOi+J6kic7Sw1rcbxbJC8VCMHDluzkcnLrHamkPR0bcT9pRRlyz0y/2h4FMb35K2pRK/d
uR/GAN068WfFFZOx56zWZuji/cwqST80xw4JOm91eufY3M/bF4c7vIYY/bSQglocIlWaViB12IlE
MAncDYoVK69TpxmB514fuF40RJAXLcaKhFJTgjpSvJ/Nt7NztS7NO+hbOMSYC8CDUz7sGbnW1v0x
UaO1N2xrHsRuaPB3zA1iZ8NOV4L09f9NgM0WGu1u7foy1HYFi2wem8t/8MORe5HML/JyunTwq7Zl
DdmXzAROS/6v6nPAwrrxv4cKOqB5NqeRSpzcuRtWWQhEv3FoZXGGWVqcREF2a1SA/NlSB3jMOFKz
/Z32emr2lPhANHbQP9XpZCB+8CwOwIC2rCj23gNK2z61iFE92eWb1V1oZk8mBngQNsCd6Z7XvUPX
wM6L6Tp919smIjh/BgbkZ4WdhFny/lgxrB2e1L3qVJCDarySotKz1d6W6LVsuAk8cRMDefDNyAOB
zyoJEgD3fbg9pgFdOK+3qauNIP1zvnq9yl5L1yaymPsXVAmylBihKN9whmhKqqjJ5RdB6f2/MBS/
P3SFiSSn4CHZ+Q1wCN4W741241LFFXyreiMEflf3MfMSXVgcj3fDLgffjajw/lBEP0MG8y/Sjwwm
MnsijUyShfYCDegt4owT0G4mHp/iYC5scS1Gg7QiGAVtSfpTtm7YZ4UARQXOxeRWHXrl4Fp0vSTf
HwOn4JIvNtevpNoeCyq2tGPZW0gZ1mDO3BRQ+VhaX0tR7iFETm1eWy0TnFO3W2MBIda1qZJ4yIs5
Yko3pmCzWMlGUc5MEZysLee44JPNyOKaDOw0p3VGC1QFrUBG5tHXylVTcjIdwSf5Nv+n8v3QJ0Og
UcMJeoKT25qV8g5rjmvZzlShtvTsoBqAq+vOLa0Ecxf/xsSB/t8OwRd3cNDbHuI5GYpFcUySqhk+
wDqLHQdvP90YIITrvm7msrCKN8e1OqGhHfsx7Jm90vXpqgNwD8I5AMN1T9rhEJvBq/5qpGf+em+7
NnnaI89R1AnjmQQOI3lHiJ+ANGHkuu8mO9n81CWYHg618ZkcTtNAwtcYEE4jzkdqQKkxZNMoEOBD
A71S8WyEF9wmKfQqLf7pS0jsUxlefGoDDD+83FDsiY8MYgon3ybbZ5QfqK/EoTHia6kcmosLfUWw
rnnD6lD8Eb1atR1MrwiiRUfGcMQr85sGIHMbQAGRsYNEo+Xfij1uL8/sbw2aWz/FwPqG63jKXh1c
m2TFBWKEThqNcRoEsDIMCyRxACnyeYbXghGEn8Z6HhoVTJsukp+pyekotNIcoTr9QAkmIiMFDCSb
aJGxVkLzmQzTooDQWpaLN+scOx9PA9pi0Wj0oVpCTTsLU1KYqNQFFNn7ThobXb2o3PPOzZgtaD1k
0I+8rxRM5hX9h+3ijCNpLxFrTQ0PP5WkUMMwS9EXjDrSLHm+UffmKebJ0/hbXQdYLwI3BvsiJfko
u2hVnt7levVP4lG3LKDQS6731od8iL0ioYvxZYyQHwXt5GDhjIKtyoCJUd50m76eCk55/21gj4Zu
WrtnNoombeFFGQ3h0Y0BMM2Cw7orwJKHz7Z4w9sdK5/hHgOb10fqs0shU837k+7Jpup3eCBYuhXQ
EHRf/rYsAD36Wal/VSjmiMq0FoQyoHVObtcYftCzzrM7SrFe126NLfLboPJBu42N2LPuV/MD1jRU
h/eYAkOlHvLFl08HWUWIjoqmkL88YJMiKu7Sm0eYL+fDmVQyJJjNWPqzRM4WE28Aflvm3EQkiIE9
7bXdCzL8e0eca4FxuiksqzhmavB60vVsGVzvci0kirmtHhnqstndMIkHye4/ZOao9Eo0lihPTYwc
AXz2hfR0oYQdNyALztnwTFZbn2iocNIbBT+k29rvu1G6ixb0RBavsu0dO4ECg3X6AQV+nK3ZKP56
imIG3FUcLCf5iUSaPcUEnH5A3+SxhubQ6Sabc1UvjfQgN8RmZJJXWzBToM1pHhJ3dRY08NKla7Ts
3H7iYn8GjoBXuJX/E5FUFEVpG/SAMi8wBCAcncDngRInuh/VgBjIPur55Gjcmb27EG1X0624/QAr
nGOFEETuaBXBmj9A5krpS1F7nLfJL9h11f9mvt7G1u5+rHoyhc2sUWQK0U3E7tpLqPcLj77riBRs
u4zvY9cFcvDNPLj93FyUYZpEKcn1QSNxyiMzlh1/aEI9O2mXvf2q0FxP/4mGkDT77ydvmXyatVXa
lxb/67h9VO/Bki1VBBsWe3o1+eF72km7v+O+OqP0sWEb147XZkwOT+c5kIL3aLECv8+sAjyWcOZx
fnVOCIld8jQV5AaCegKJYXkJa7cyPnQ6gUSaUtgvg67+Nj3eVl/812AANyc2oKSUEFtBD3/e3+3g
yAWog/8uj7sVcX2NalIAGeKDWQ6RaRVAKv5IlH8pYIwdqnyHkxO6ZUvtuc9JbBBeZJosbAzcNiS3
OuusmtMshGKXqMCb8GFHE+v6ysZph2cS3+KeWRxfbBETc+9MpD6kEBU/kyn8+Ivwky6NG+nlHTba
/6G/uURbSCGB54Tz1/fIF7sCjUe2Z/2bqUHF5n2yamicPtQlYJV9LFE175mmzX6uHxogjULCtZQm
8s6WOVJkdW0UrgEvGzcMR1Czrt3I7CdVVpXCZyTSFDVDT4jB5V7gTTaB/zCZb4MKZi0YiHdea4wf
Aoe1jvGmBJcgRNaJ0oN6Pva9JXgJKc24i/8hgCteEicuaBod9UjcVc8tk9aBt3YKY1wg12Jf4Y4h
/iJ6reKs5wiUZyyZdgafF/ROycX9GCo1tsJQmD77MDqA0OmFM6L7+o/+EslFR+MAg8/e8GPizgSm
bL5lzK/VCsvyQ5qH4XMFUWZvPmthwtnbHDJmKDJqQ2Kkqbj8GNnF/XHrc+4G2xE0oPEPWAf0coFE
LiQgCZ8mWEaS+oJPpzMNC5KkAOZ3LrQ6IEfyXj+eNh9oj7nsu1WoUOeq1rUk7aoWBgYVx6QHxxqP
Ef1wkCY6Zgp3CixlNys6DJjW6XOmssRINpAlZURWqHqAxt7mH7u2drUqOTCo11jY/tnxzoSdtKmy
gwj55VeXZlcrpflwKUsYO8BaZvjtEOEdnriWlLfeF9IEd2EorGru2DXI2lID8iNY6aJ20bAuZHwK
cKkzW7zL+Mt5thKD4mm3cdPdMD0+EJql8vCfnYWwJe8KLdwFNZ1LeKiwsPuLe3OR0oaWAj4TyYY2
S1PMu5FV1y2MT8PMoCptS/DrGeoKQ4eMkEc59rMd7E4AezhUykB2tmKb1X8WCj8CjLHpy1nurLDN
ZAtuVoiIFPq3smlcmWgGOh4myYM/WsGP+dg3le3tTBixFHU84dYXK2TcUn3/HUYYdjRQTfA3778w
6LUp6kl2f74/NUCq/lCDp37H4qTbpyZFwFF4B8pnEmqw8RElRgSUKPexIHBOCT+wrvKoeG2KzBFj
Zd/CQxAz2w2UZiKsLYCQwZZqiPSeM+Gt4BklBi6BxKGizvE/dG0MpcHWJ3hGcShhcXf40I2MFHAr
+emd5nFFmCVv1Mg6LB3RrkpiFa2deKGR9l3OSJHcMnCRsUq/CVAZ2TukVvPO7xcvUVueNz8mBAvE
3x2itoWcjf8vAVOsDR9qh0XYKkF5DsQ2eAk/XkbHLTpjUreAwjDFZRYTsLnd7ZSZeSUYvPzPE5JR
BN1mZlPA+3MIBZxA7COTy6X7hu+XEQ7KqS7seVnMGmbAU5Lo7lXBQWjFYE0K0yi7kBTuM60u+z3P
vHvHsH2xG/lUv/7X1arDUX76zbi+JKMSy8Awvkzi+tzQmMRy1sC/jPig2SYM1f36n4ECfDYGz4aw
Gt5yTsM3yisru7zj1iPuotv/EeRtk4tAoEH/wh4mt7sJ5Z6dD8chRrFJVHFEVZde9uwhpMz+23Io
JgMGKBvwbuK/G499l7O9t9Qc+sjpTkgMmYOEExpUz9YSPELPnuKCydgNB85olly5tmGXQ6DdG/H8
H3hfa4LvSWiZUsLgb/u8TkX6LUQ2o3O3ktBt9P3m/KtMbfA1sV8/8XORJz/8EZ0BJUJsSkDhvjE0
lQlm4hQAkdgQJBqORT0aqDGu2sCxM9TXCacTzsRLzFf4Or3yGNnVxATLbR9r/x5NwZYjJwnI6HIW
PECjdf7tjylpthRIAW5fWy84uwFxkYUGC3A9mgNKwykg3DObkJjfYpSnWMQIzKlStuPBhamUi8mL
Jo9T53WHNntv6wGFgk4yM3T8dEtSZWNLM/8c0RT//jbKBBfU6TgBYSWijoJAl2mjZvf6ioHBSZQ3
z7LX9lopLMu5K7/wuDWkBsgECVq5//SeDr4m3CcuNmp0QXJSa52Ba7ZNBMxwRdwvQ1VKD2AmVSuW
L+SakILuo1z8pvoRlU6fOuqbfz0K6IPVMkx8/cWU9etBiefkn+gXjvFk3FOemA8BEoi5ou+7Sh7g
46KEzE0RG3abVvrC+tsGk5BxjUV6RGKTVHNnAcQMf10xppu15nGlkh/FA2FYY9NmZy1saSJsT6Ew
zloL5v/mE+WszYOgqU0NApWMinCx3i/Udc8Yzy8hgcv73bNVc2DGg90tYZkpQSRDWnHN3CxOwmzU
MBOk0VTshWpacuyatypRUt6Ld1PQqbbqZpu8iAs1+UkbdryclnSuPNB4JhDh3rVGrAj6VjmzLUmj
mEey3wbAVBqEBqxbp2to99x37u/PdLGDxSpcZW9Y4Ntw6j6xOZ7oLqgPE7E/kdZhGOlAI8LImzRx
0oY18O/e6pZuBqqLr5y8KSy8nr5ht/+eUId2IQ1NNB+j6Wko6Ko++byOBnJwZXlb3RJtFutDregl
Y56j7rgCSgdTlTn6ajxxLQWk11WpV9u/ItfBToUKemWTFS8SNF4w5vs/90WtOX6H/fclxphIe96q
4gaRsNTWJFtr+i+yD9BPIxLkYsRxza22pQBB042XC3th7mNSdGWlpq91owLFXR8cAGTbxCRX1u65
CljKJ2nR5rt7k4+0uCZLZqxDS7xSj/aPaD0x3lHoG6oW8HwifHVWZddCD2Ici/AdTMDh4dgv+RS/
FRk4LK4wXbCyXIsokKg2HT5OQmPy5exLClJF9xAsatHT7Q4YlVSKBEy+qWqBfuIY3mNvhCKtEMy6
SMP3D1v/Pg8WsOb4I6CMF2nrU49gZgHIhjlRAzSYNIK5efBw3niZEDuHsvYIo7JrKNw1aZoFgzaf
5JQzLeVIE2ZIcjBwxRSm8++WkihF8TvN1FSYPQxLI9R5JRubTiKcg1vZXh8+G9tGN5oMKkXnCUVX
QbkcmlvnWZOXiabfRUoSbALWg8mhyKWwwpb8AcA+BjH/c8NZPuPNOHpXtzmeRQcH0tUt1SUxRUti
lXOTvhUH+aNT444JoiiMb4DX3NEnDeWrAZppIkP4SVsuSYf4hpAJ6wq37vUC412kW4Nk0/D1ghnl
DHz65na2AKIQJzn4q6KtkhHJBuwfj9vkowUAF7vQYNh7uegPOCcRDtNmSV6eUi1ovCu5A2kqbtwd
/hl+BCz3pfTjucaMSaR2Nr9wJnWROgY8Iz3D3VlTYHilH57lhqAcRA3XapDhWXudki+RiY+0lvjW
VkcWbzaxua12R+t9ER2l/ZgXzKLu9ubdCaB73geGOZ66SjDa6UR7tcKabXAGmAzs9m3sbYCSsEMp
L6lWk86TA3iKHv5nu1zOmj5NJdNcWp/8pAFIFxe9OftlFYTkaOEdvhNrJF4mLR+lNY92HXQkc9Bd
Sc57YJMYU0deprECEfz/xDlBLDqaKLJM+rpgem3e5OXLM6O5hmvIkfD+TqHlVpMQl7R3/9OlcCit
ZYHRgWFjt7nGC0CGzwTxkhpvuK5DR8XFhQImnDgCxD2HFy5w56yOFppQ97tfJ/N5aErmIsfQtfHG
LuQzZYRXtOuRqjkXT3EK5/u5NK5mUy7b1Y7rmm6BWav8LVBlWAqI7V8KpTiQ9NL5kA8viDjTaoM8
8UXl68kq1/wjiEnDbVA+pM1NJM6s7AulLvaXlCulPUEGpFG1NmmbtN8s4j2Bx+mwMsGi20tRNlcI
SA4FTflHqi7yjdIlJ4s2L1R0AT5/CAFEXgcslWbpYayyurCEGYIhbDxKOATEMKGq/jHAFXix1OhP
Bgeg67yySHA1sT+WNZg+bqVPeyGADajFPaLt6c21c1h6HPchA5B9gg7Nx6Ugcf9lbXu03aMbz5Ay
/AuhShBMI6QKc7yNz1BWlOZpu0cWa3xNQ1I8KvJsqLmnHuVvvK9TlzzUjhP0k78Ot4g643x6qrxE
rZJchOTiw+5/1I8Q2O0sggN4p+9BMAxpqNPgrCd2+hT04tu0NHOqlMM9AKjk/6891C9XiVWgvMuf
Z5o72YaKKC9e5uuLeIZ/R+VaL0AkObgL6yiYIVEcMFohio9dF3MTuOxPtHHEW2OjjmgvJ+QMCfop
ov2QJggQP+uQuZYk59MDAGOsFdn0TCCYaM4IYNAoW8Ju/JI/gK8Lvd1SdyKW7WRUHN1hrd0k+em1
GD749/LLvW/pOGKzQgcjorwDesYSg4St3bm0ssAg0eygqzdS7XtW3UksbqgiL51M+ZtYIjqI5Bvy
r9B1agu9OP+ZKYdjUO/PFqzbV5vwjAgyQ0DpTTDQ5NxKguWLasc9jEBcLKbrOheZH+wEnh7uYyQz
YVDu1CfIdH7Ig2sRu0SNLjiH8Y5I1+dTPIIKLZ3mGuqq8sBkTW2lu4EH0ZdSmAWrh9pzDUBooqgF
PalDOc5x9RVMoXrXPUOfGDvn4TT9PG6R3sZKFLYh1eneJFx90i5PahyIdfFbX2TBS1zL92pn+zS6
12jwi0XjHy6Y9NWQ2D4mjKGh2ZMGNoBcAvOKKvSp+Tal4c4DfEkE+HS9opE2xc8nmGDg/WK5Dv2L
2DMgGqcR7SGb9nLwYtkAGgvIHrwxAZ2nkP/i0O3zSMy8H7CIFOPXo/GFU6k00CDo4ziQcKImHRW4
2oBcH82NVQcFjB2vMSie1mop9BLpnrrhYZqq8K/tiYdVqcc3e3qpFqKQaMeI0jPoJikIY9z1iJqg
8Qp1iDW0vpHcovPN68i4SSPA6EjA37oT5U0akcY4lIPgKsAYn6KQPqCTsRu0CX3WqwSiWIfyG0Xo
9LlTYHpujAiYVpWKMkJ0yK49HvXMgkHLdcXTuwJ/wRzK3D4eZrrwPsQyWyXy5TOcIT9gwIquyTbC
C5NroK7LBK9n+/iNOdElSV86zDLh+NUHv39ycOGgxa0YgE0q3y9w8ECcArmsQM2eoIYQcl+g9H/B
B8b0z58faD8f00BKHpnCyWlI8asy7/wGt45O49xl1L0esc+dJqsSviii2SbOAhC4bDjm+RlVvP+Z
VzMxvELOEFrAarrsSfgbnCUKh5Rtf2wnpUnIs7I2BCgS4SlDNeOlPho9G7AvjmOSpYorywhxy670
im7tiCT7vv7tQFuAmLLrSipE2qZ0zPTZzkspcG5g9e518V/VfGcEAyFQuMshA1S28xOlf3X4ByMA
hsLrrevU7FNgsJEfCIM5Dq33TF7GM3i93B89HMHFQgZHR03f9JaHkilXU0oL1pZtgPG1TqjZ75aX
DyZXb7OAXOIbZGUKES+JX9W3Uty/Koj/UNYJ9xtLO40IWMsRJGRdDpKfAbCCxK72QG6j4q2yIy/W
0jrYm1O1I1+dZuLRGUPJ8kbbguULND8yzJ0YWcNNbvqclvmsE1Z0KIugVPEKfj4uBxO00PoBDTTR
5Ed06/AJAA5jrwHFzpC4/qDiAcHOKmyXFE43ySTYNYvyrCxCjQcwd/pL7WvY4UX0fS1uMXSFtqh9
nCoOmIkzxWAIK66iJcTylTgHArLJoLfN/TW3FVbk6blczowal/f7P0Q61uXQszshGRf7Gia+ohdf
+z7gciV+RMInJ7w4dAJ95Rw5/FZ70DWLl0JjWClhLCL3cOIxnA+/HUMIvQamNI/OhWnAQphJvc2y
d2x4BRUKsR3FYoGf9nfUsjcfRef36VTixb9akc/tQu2NybV1TOkJq9V3r0uQ+jxHb07dSegC/9mn
t8SBt1VxGgdf14tELYsiPoEdXZXwiAHiep4if4xta/CYCmgYlJEpxA8Libil3NCg/B4/KrBNrFZJ
QfqZtlLO5rGsVjm8q9wAUhgxZEcCVI5N4+5YELs/yOhXZVooTTMp2g0uQz0PD10Aiq7x59lhc9iv
y5vvWJK/oU/shi1oPYTW4tZu2RHurOHV+kCaYggH5rou9eIqnPJsx8YuwKupXp4rH8SZMsLkFy7p
H1P2D1AftRukqQKye36bTDEjg5YRz99v4o9JwsqDkRbM3xIjtC4TU//CQlS5uVwX8uGuXdH119Lm
v3SsXVkjqNpksi1J+i5U5uTgBuOmCfy7wzCXF+SV1MNUmCCavUBp5dKGUCH1mT5WDEzKW7QYjBjH
PWnzML7cX8jGdNraxAThn7YB1JkrUhCq+XcsJbLwXfL6XT/0DxbApwyXg+uBH9IKbIHqhyBTVEEg
l0E1iTanMxG9YmVRYETMNRYESPK4FTi2HP10q68EWXJcOtAVu5TqL9rzE2EcjGe4X3zgeUINsXRK
M2GQt54YAD9eLZFXDB2O+TQfVT5x37wkSTBh1LjdpBNG9/Z01KgFCyk4UfFuk+YXYDiFjMY90jDP
dwpc2nxhjCuZ+3kJLxdVQLPf0DVNiHlDlmvPzUcsj5QeMEqYcFywEZFk9BdDomg3nNXXtDixmBof
ZGjBXupK758r2N3KX6ZAoFAPKgNu1S/spdMaSP4cxoEmAj8KN8ELtQKi4EwsWCh5l6inGdbNZh6r
n3PKnn1WGaAuTIZvgAynP8E7L3xoKZshXmskQBiyK9kukRLrcGGfxeTXjTIruCHQYlUR/hM/zfJq
u0BNs9CKgroY5O3u2TQPPQjbfbcl60osVATAdyHMijZ6qT235j9bIEfrIZ8dV74mze2g6ftoEH4k
r3ptSqh29wRa9ctYdCj9ghJA19JDd/uiCHxgdq4B6ElqPa4IQEqcYCBFEREJkOia+hLpN47fTyPM
xy2R6mpQjoYaDKoUgWMo6rRHRQrR2apkkMIfL7wmi6tBHPIjwCg20DmexVlUhMq5cEBMSXL1nwf/
ONPaG/DNZLaQX3ojh2Vr8yJWmcQJLhnzB/oN2czBsaf49kaelclDcRgiD94QOCe56Gl6jpWUFbXD
ZdlyZv7GfCykUyYbFWInLdFkoj3GS+oHy7pkjLhPlrn9t+GZyzk8erW0tRNc+QO6dT1TmpqfM5q4
PhFcJhPU5O1tNefAtWlEt5fYDouH8D7D+BczjKsUYrf3MnMaYEFNC1vJENFwc+PVuyjg2XS92N1x
uUhjOb9Yd/tqTBFEE3vdZG87WrFKRiTj8pKL8m1v65e9AKg2lFPjzZwEFheOhiNbc2P0UWl5neJQ
rg0a+OTqG4a/6DGt2Ulx+DPWIFZJfFodmOhE10rDtcebZQ0+7AUVC7d9OY7Mt5lVPhTQKmBLmQAP
d2edZUa+Dbf5b3HAOr6AsUXMvBGl
`protect end_protected
