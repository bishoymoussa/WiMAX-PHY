��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$Rx�y�<��wA�*;�x���@�̦�W�X�fa�M-$u����n~�%���P�$��W��kYَ���P7�?UMfT��q�6�U��k�>����~�\N�(�����X�e���/6U|)�X2pF�]$h���d.���9E��WG��L�X"]�Ad����ľS���8od����e�GT?y	7�������ݵ�^��R�q^]�鍦�����s�ae���h��L��P_���ާ��YЭF���'\��68�b�[����w8�[X��V�F�0͘3����q諵�uW� �h�u\V�?@��_6G�_�*�G���B�絉�f������[�G��U&�����~�F��AׯK1�`c��[<��FY���4I� �#�G��x[X�=�Q1��`��R>(�w����R�O�?����7�,(�H\�#h(W�EH=�������yq��Ѿ��aF����:�U~m<|��.��0=�P/���4ǆ���T(����]�┎SR6��gV��ޒ���1_��8�!t���y����cN��b�ƥyB��X���M��s]�fl��
u��G�I���__X�C>�N�5C����)$;�;[�P$�cf��/��()�#ݔE�l�_���}d1�MͬXd�l�e���?�B�Z�h�:��z�����⑇��9����Ho��~���V� DL��l�m�EZ�FT
e4��
|�c<>jD��*�i�V�����.Ku����:��o�a��ƌd�|[�2��h.���䶶��� SV��~�ŭ
U���]�rq�e�_���%�a�x]h�H�*�z�Yn$���)��ܛ�6�lc8����xl����eƓ{g��{��0*�c;�w��<'��ʇ(�E�ؒ�ʷvV��u�@���$�^�t�4�htE}h���i���	����}��n��w��એ�F���;~��>_U�\p�r-�N�M~�Z(��j��Љ#������8cn��X
�~�W�ȭ��Z�4�����<��v�Տ�ŗՙ9$
>"+Jm\�(07b�&��"�u��~G��MU�sh�"�-%��h��bXjiJ8��q�:�o��6!Vo[2�b���8o�K�z8�9��xt,_�M�r*�J�16I�������/�8����i[k�i���
x&�-������Bk��nd�^�4�M��gPXǘ��2����#�W�T�6M6N��C
�?��`R�]�u��U�4o�Ge2�pwf��|H1.�| �&��m|,�u�*p!iP#�6������� gw�E���6��17���4\��	���py�3��F�22�0��FjA��ڌ�P���e.��"��6�|�%��5�P�Y��(�Zd�h�}R9߰��Cw>}��"�5e�e���7�k�gQ>i"K��yV;��1#���[�si^Ty�-N��7ChJ�ow}�^��AO#lWkYq�x2�-r�?��ia�Wn����ROg �u�}l��a-���H@����6�W�) ��j��h��VU��\O�25%e�M)r���RħW:㿩�\�w�����N�^M���K��J�/���c�S��&�ň�n�&�]R����ó
��]�I��ܢ�ҳ�0����t)���i��V�rʘUA2�|:#���?.9�P���09��JS�x��+he�V$���L}���b�"n��
��fe)r��4��[����Q���|�������rh�¡-���農��b(̎bM����/��&���q:�{�i(����nO�Fk���7<OH�1p`��p uf������]#�����K��\?{H��~�Zu��Ȅυ�I�s��q�=��2o\�DKYrD�[�.�K7BF�5KQ�T��zv��8yM��`���ǽ�<�uZ�M��0O0���L��@�[k��2����6������}�2�����Õ]��B6sR��Ix �V�H��3$45��"�	JPr0>���E�R�',�����"�KK/�'㶫��K��4�?;C:�;N�y%�z������9
�F��s��qI��(�\�"��8E+���P�  ���6�%��LlY�UC��9%U=���3_鴲�����T�|�uf�ux����R� u(Y�KHD?�S�=S���WY�X��%~����̐��x�0�vn�i�z �Q��h�s�ᚖ�/&rW9pb5gf����[�*%�)"A�t;Sr�r�"YXT�<��l�Y6�j���E�5����_�B�6!U9"�|�'^p��|ɋ;'��l�x�zȽ�8n��=�p�]��a1^г�����-�Svlh�{=.9ca,P^�Ί��V����sƏ�';d3%3Je�?�@�<��d�ec�e'�^��H�;F�D�q�~�����#W$:2�)Q7��~���"����P@��up�Å�b"ҟ&��
�\�8Ҕ�� a-,��$�-�L��l���0A��)�<`�d�b&�D]x'E����!�
X�ԅ���&6M����W���_)
�D��Y�^�a�Pי�&j�ΛRbqh�*�W_�'��y���0G�\S~M��w�h8�lm��&'�.J�eMM�[�L(쫍�n�վELPXt��yL @��Ώ1���D���
�����m���Z��p�
S�M�'$�"����O3�\�{� ���o�;t��;�Sw�ο�`pkc�Gr� Y�B%̓�.�8�)�ܰ�䫄yn��/)zGk���<�/F,q�gP�:���u�b��X3JI8\���wyd����<H�
��R��3 0J�/޽14��A����aE��*�q1��~��#+|Ob9E�,�ņ&�U���x�W9�Q�)F�/ʔ� �P�(���ݚ��-�x'L�s{H�S?�]��4�тɇ�T���C��-\�;�0�rBE�\���\��}�����tQ�m�`�	��_s�`��r��~i<�}��. ��:�G� �p$��m�{��ٯ&����[���*��~�]
ܪ%8����n��VrL1j�fM&�1*b�5沑r�D/wb���IJu�s�V��J� U�z�R%;���z�+��������,-$�=���N�/�r`�������1�5)l��g�j3;�u�%ՖtО�k�s��h��r=��3��q���ɴ��<`�/6�A�N���ƫ�`�	_�i��:��yE����l���	�V��zV�Np�88V�;��}J�5�ʩ�u;�ɩÓ�����P�/��f����y�`$lyw:c���9h��Xc^���f~A<>
�ڼ��Z+Z���[?`H���E�Y�W)9���J)��5�j�ɯ�KFJ�_�j���NZ�9]Ą�.����K��T�No�)��S:H�8I���=Rzg��d�lo�����9�nA�60|�떸-gEj�u�U����u�I��<��B��(�xz�@�}-:�hL�9��n1p��TY2��`�O��f���9�V'i�)�n�zO�]x$�2�8W X	xx�{��c�Z�/%Uf.55�iP�9q�]�uO7�#^J�϶�2�`��f ������sL�}V<7���#�pD}��8
n܉+j���˟�2/bT(��C����Yi�oi��)<zO1g9�z�"~��uCĀ<��d�>��@�MVb�C��__d��n_w����/d��&gw��8Ho�J�trL���٘�����h�8u1X('����x���H<�P�P�U�Ub��(b�mڹ�W�`���X����
��&"���n2��� p�' 2�Sf�y�8Bz���m�2���Q�!s:��`;j3S���q�P�ˊ����un��(��f��b嗙�qv
�����2��d�{�B�Ȩ���; �iŏ�]!)0� >�L�n�e��Ҫ�)�|����sG7pS�e$��4��rH<��F��T�B�6P8�ar�����N��ٴ-~�ʾ$H���P�(����E����<p�y	H��q������#>�։���X�m3�i��I�._�fҏg�YȜ^�$;"LY��E/5���%'qR��9	��./F�ah�`��f�Ju�}!1e�_-��E�0~kĬW�k	��(z�$*��ϴƧ/�rsX��Kߪ��3���L��)|+D3tΧp�mSy��?�f�zlN�Ã��y�wtC�r��@�;}�H7f��=��nb�u�������`3���X?c_!��^��C~r��=����`S��Ja(~�gԏ���b��&��z%�S�uh�����'a�R����̶{��`5=���k���W�P����)Ѐ�{D��;kǏᨖ�-~��j������T�K��3u$�oi�D�Sx���U��w��h��,U@�`�l��'OFX��F�<��M�"�χ� t����=�<���C�&�/�]����3LV�}�� ��/���qt����Iu��
uz gJ0	4㘟��o�w���n��ª�����Ix���� �ƌ��������cT^�Uc6��e�@���<��EƗ�'�DsLK�W~؏�1
}�?NI����ْV�B��2��Pm�m��x��ן���M���WtQ5�{e��IR�8�A����`N2�~QeHJ�D���B�C��1VH���B��i�My��e%���z�2���)[��PS��O�l1��@oU�/Z؋ѣ#|I�}onoj䠾��+����z\�J�ϖ�(����YȺ-�y���JKW���S�0��u���%�hWF���=M'k��|�:�8�Y���|x2���!�o���R��CX�! V��}r*���z��4��D2��:��k��(.�A!-B}�6[� -��1n��R'vZ����.d�Gkh@���������	���#\(����,1�#T퇿�O�%�a+�O��{�O�}�<d4�����f�a���K}o�@� <P�ơ�!'ڈ9�S�@CN[^�<������[痻�M*�D���!���Y�G��Dm�ob�7�jי����$����s�ݱ�?��0����4y����d{I]���=����1huN��!