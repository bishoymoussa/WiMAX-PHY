-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
ZL94+NfcYPzG5/AJXClU49cn4J8AogzCOHWpB7URxpZJctuOYplmk7FZPWHHogXgMK3yzA9IxMAA
Sq/Vf0ac4kNTFD0j++/mxL5j4El4k9nGXEhmVOgMl/faiYO8xk5nauQf0AlObrGci7C07qHdWT5O
TxfQdE1sr3+rMs6JhqQ6x5STZf3yQSSEyuAbkl8iIq7cQ5z7nTLwsChJafs6Q1gXfcNeOAahD7H1
HMq7bHHPtN4JjtD5mxOAzgKIaPiqujJ5xLr422doUtt0bblw1JYFBT/Yr9lV1gmvcEaul3iKWzVG
4uG/0piLV3JCFvK8HOSuyW+D3J3YLh8qw1JRbw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 9728)
`protect data_block
ZiOIYXBf1pMVJ8iSJLtpDumBi3viKEmi2bsBTaWrx2zkxwQOVfz3FuZLhzRBDlfDVLoBm84CDfXQ
ozBqr7vOItmNGEuBZIdXsoGJPzmP9c00T5V19FutVD3KJYRXGfJzxrKjj10QWvLO0FHOdpex+LG2
LUbXSfKlppbT5XImbG3NFJ7qv8oU6hQfA5qTt3sIYJ+X/dn4kPxDVTISm8nGeejd+OCNprLyjHLa
iChPVNBehMcmjVpC/6A5ZcVz3lclnlc+5vsY93NmIe0AUBetSzESl6zorBLzO07O5nSuZwDGF5EZ
zq+GirFzpd2RNcgEwkqxAxSKu9K3NnNH399NDxm+NlVralU0nuUcQYFwKZ1W1JuTkeXVPCpMDrxi
dg7R0LmTUWPPdBPKQKxOLTIc2FFCRjIxHUyoShCBb/drgW5eMmax1eeX+upa7Jt/GgzQscHsFd2c
bHZa8ZZUySY0ucFHjj/IbhuExSBSkcAdQIupJrG33LCNoiI2w+fsI/j05Tefri19WISyCi1NVJPP
WQG6K2a3O2uyyyfK7m7RLvLVaFWc+88y7YLuseD+1onZpgMVHN0kjeVwiP3CH12asHyRTvBaW/Xw
qAZSsgz+ucKqTIBiWOx8czgKx6U1ZKZGl0RnHlt54ZVAc6RbwAJ9s4cBojpoCczySRNg/oyMWY34
zagk+WqTCF2g0NAX1v1w8RYDiro+JvRZSQMj5IXa5nYBnjd1FGQWHEN5H9HDzJPqPr0h64mw7rJh
nFqnKHvLt+PG9VmoZ6uBUMVMqUmtEwNtsMxirGCFdZMrPwsEmVAJhBj6OWtoVByQwOUzuULt0+yQ
xWPofaEuoanIrBj8QtoThGsM9AYeEgJvvw60AZF737Uq7C4ks/fDGb/VotqPcLTUyHbrOS5wrmGV
nXIrUoq+f3py2vupc7OOQWGSLud6SlKVsnkB0tPqLOt9yy51/X0yOfmhfsa5Y2RVAioOIf1RjM10
NOis2BehJwOKwMKnDVgk14u2qU8o2L43paWG03d6jHZO13hitct4fP418S1Kqh4+icaZOSnQ48ao
k7FAl9cv+si2AeVig4sDkAaap8Mli0bZNB7N41U3VAW02lOZcnZTLfDiV4jgK4v1pj5ugIz1wvtG
1JktMpycV96VnY4c0E/lCqaGOVBXaF+HX6sZqX4+oHUrhBsL5VB+JdOnYnFh+2JcC3+sM1oGQvkg
03ydeeOlIngq+9FlHKnPj8MIjJWo2mwfsA5bubvFONVxs9ujhQ9cyWbi/W01y8Mt1gxnDsQYnzW/
uioZP0qxh6ABeyyaB+qcTeHar5E8Y1OalVTr8i/QtSEQm5kf7Xk6A9LeklyVQJ3BcQ5YxS9G1V26
NFU+AokzxSmwiO901UikLKKwin5v7Vtwhv1CDH0348bsVpaTwO2s0HrnM/Wzlt1y8Rp7L+Uof2sm
AJ3JkqpIW+9tJN5t3haq6ItNHs6fIJuZHma5WPKjVQYl7JamFDvYWZCnyDjk3U9OqOsvKZht0Svw
wxLiYz60PAOILymGHhOiEn1b+y2Q8DWlGII/2OoeQOCgJQN8tWnQZ76HoZM2qW/FrmEcOW1VUc2Y
BLfynepO4BW2iS+TYnqzbklLO45cCi5BsFBk3xhcCnP8e9TH7nb9JKrLp67HVxuk9pYTiSkPEaFd
9MRj1GXhO0l6PwPqXGJvxEmeajlgkU+Hi8FmdrDtodno2X1hvX1xV28A2a5zQhMs13IK4QatofR4
/XuOKeo27iQRM2wX4/TGqMPXqPvVdLolyIObwlajXBCaiERHE84ySzzmB5QMVYHy7dm29NSOhB6C
ZIGn6pGcBjOzqXmprKNYo/DBbHwee8QwopQtjfxMslxcc0hAwZS2Shb5w02t9KX/NgQEG473WIeI
6MCEjknu8PBw5z0UrMGSgYEcfg+j3A7mDMzI3T5wq8gxsZg9ipO4tEdahgpArKstJ1YcygPCCoxO
UdbZhkUZid0TuzY91054S0E3fKUi0JUl1CI3voOg+g42rMuIutLsLMVt4ZnWxk7pW1d3/8N2JvB3
HKR5tf9Dc9RtMYmuFv5E99gh4JZfeAhA8urFNl6Zo2hIBaAB18yw3TNcKewJBZDEXE+GT8wJ30V4
Q+4psg8xZsNtZpqVl6g3yDGFMNuiZEZ2pHJPG3tHqUa7R1aX2WPylwQoeZB/0rCcT/WW2XNpqPTN
yAflq+3ArwvO3iqGRYwehX0sRjMkHmmslnfw0cE+FvHMkvVntcUBjR1mlM2VUr30d7j1lpa6swML
QJtjyw84X3LF8QbHgmoZsuhlLMTJLj3hin3V6msEMJvlhNMSTTMeXlT1ti4SY6ykPNZUEDg0wdIw
7Y4b2FnhjT12XGEHxpNxcqH5zxsDc/iIGVvQuoLCG/QZVgluQe3wTuMmMWahG8B7GYFUj1uyGKoF
DMP68oUYv2WrHzyP6YVh9Kr4jaRY4GDdK2HuqNQ5kKfzic7Ch74SB0J1jYreLBrKIp81eHAwV7ka
P4vwmFm03VCSoyhOxwQtrS+40z2wS08//teoJtZ9wcnV1Z0K8r4uXZbPWPB10PJ6j5ZoyH513EvP
GFUKLpmesZLOcQqroBJx/soqE+gThkSUgo30AtIilZYs+RHAaA6jT74dfg7hvTkJF4TjA2JELLwM
t/jY2nSPMb/Drjv6dmd+BwoQcmnve+EoR0j8fJaPgHutABwvMeK2zVzFOmFW1WBo0uK3Ndquxrz8
S/Dxj/ECew3KHs2Y3ml562k7LvSzXxE5gwH/m3szT08027dIUj+X/sDTI/Bbq8D+60vBukiS+ldy
F3uWzY9XChIK26ArYaajPnt7lHo0OV14Zv2oSLIgV1ePV4q1jZ+cqybUVNOJoNkx4Ws8j1Msz064
yTje8R33AYWUIfiTZeP1zwukYZJstB76b7SeK3LCpk42hQcPjskb3VecROoYgZp8+DZh5C7JIpVo
g/OCFoaSp9/nDHvflkq6GPZ/1rrX4fEStBdKTHwEbmgl/SpOndJWdmVH9h5Rw1QzpCeIzajgl9xv
2S2wZhk3v77jrkXDgLY/QnKCas0gKddtbYpvRJ9I5bKsDY+t+Jk31zIctUy+oSFDLFMopKP7Q4MF
EWVkkKiYYfkayW9SIh94J/jpM7gqcKeY8fHH3PXFvWXAtgU2UVLUmSU8ii7zNQZu/3XrT6bpai0S
YwANKd/OORMOXk1Qhi4vDM2D3HBeS9Z7sD4iXjh62hKrzGHKoADw1ceCqs9ZKTja5gC0cSgffTNc
ttYV1aG16ooCxDTgFPLVYYpVikPrVqHT1DaA4XYyw3erAsZEqiHXTifMr+6N2+ewk7g/njMi4Ewr
86AiGjF8cmgABmJeuFAuqisTWoj+GBvFOCflEEU0rhPN4M0p0gi+fKAsHGfJtiLF+mgb+YeYSo8J
vMPEqrOypDHZpcjiXywEHiclc4K57cVI3svkzmFQ3R05dQpRPgeIFUl8gFyBaXUKdCjdMYL8ONG0
jt1Iy7zTIq9UVFC/NFb6yfQy1yuwZANcHVQL4NsdlHrnBTrwv/xgXhMEhu8Sj2F1MU25Gv9s6NBJ
eMAsgHmgEkTu0oioe8q98dakgkHp5CXB3IPhe5oSBFpa97uZoI70FtrclghUfp9qfpC1bEqcJaY3
e9De8mTiysed6uTTd8v4gJ5m1Z1yyH31+Ne85gApSWxzotZl4eyNa+DAeHbvrl9h4S5Pf/gahm00
dtsKwReOseNxKP29Vt9SS+MsbABhTZH5F+fusPPoH1EFuRdQ/Gcc9yriCvr38ydW1f6kKlJssyjP
ybAxJXLLoDErE+IBd7R8cuAkH6sKBcaBZQRSwQrfypmRwGeR8r3r+qhJR5WdD2AtcxLOoyDCzfNZ
MfDnG0quNBFSMkRRnOP+St1H7HUylhRhOhlcyztJtTuFL/gJnpWqj5vpRbImsbPjkhLHsslH/4XD
OYv61zHf99YLSy/ygS8XCoKotEu2MTDGnYTQKKuSiwzSbPdr5xcbAEqyimhnqsVkBaiFiL3Mo+RV
AtBqt5kJmlI4pccHdlhXRTWOVjVe10fa4iOtzjt3OF8z7LKA+8o1L8jfN+f2G4oveNau85KfRPat
99luoVOG+FmxeozqjVmBcuM6KNYhCV72bdqR0edumbROg/hyaDAijLDgr+jWbpEcJitGhOFjFsLt
KTGIk2bMrdGbFZxdU0XrGi2k1NUTgts15giunO1b4EFr9vPgROsAeIVAbabbI7l2/DGgaSzOW2s6
B0iBUp488v88T5fAZSI0OPzRC5tqXnmBdbW0lgdqZA1Hj59wHPRboAvxXZEQUppDrP7l47JnbygE
xXt7V8w3fljAgiWwv/4XD/QGploCX+/4uEMqBwyOgvGmZZkg9DstNQUz5SkBD/Za1sXfU80NOuyx
72WFJd9npcfeEC1g+eWkk0+0cbH2rAXHNvUObS6rEEVOMPRkORJyCPDdDMm+vF2mol5EENzRdhc+
OIO4UBDOlZCmo0/b4mJIYscBjLBqM2NW+ybNZwWyVUl+zwoDsJOu4pQNuNsKTv5j0B+SP8r364T5
p2cx13MbGBLTRSwUgSAOK+SSjEQPQV8i5J2yrX+oDCHBE482DkC50OxjCVoDq0TIGfiv31j9Bevu
jnnb58CffvzrCMfSaxyYpoUNcxirPFZ7VXNCPqyq0FH/VsNCAhA9WlP2p+lTgRvU0Wd9YIRKhqnn
OhKTHwq4V8ztBiPND4h8UMXqlVU7Qk2Uj/Bpzw1dw2CTJsAXE6KyxiaOXjxiW0yZ9Tx/ttbwxQ8D
C5bxg5qIYaqxpkkKHK3ggX3385+8BKBxo/8LqbqrVBPEiWSyD56YFrZa8IofRXzCEqQA0sn10j1J
ii8JcNgeBO9GPjYRgbFXzH3/2cO7/7g+TwhNPyBT2u9dmlh1VMHMSS68vwOwxitr+v7mKw/yrFA4
RFnTXkdOSGhgrOs5qC80LlToYifu3yxX82AtUtNn6Jcv6Ny3TGDgawkWiky68o92ug7OQxJznKIr
qtr8ZpHcbON1GwJ4BKnRWlWAfUEdGaQEkuCnTU0Kt6UtmWpGr9yJNOdXE+s9980zJyzip0zeaCYg
WceprWw5zDrOuK3UCkOiPI6V+QC312/ZlPP7hL7LPL+HiODfbDm6I8mBVoTtQ73+Bwc+fdA9GFzZ
ymLpNLkO5vHQsj4SiD1JsJUADajA5iXVccftdoitdmYmOrQ2enWV4QNWnEnadawBZltH2MQcjT27
SjeTDIySJQDN6MDhp/1aZHLKiWSEiw+Z/AIZPPwD0oiVpb+w8zF9iCso0eBkQ+/fer8bAoH8g5zg
LghzHauCgDqHBw1hArLtN/CA2WLhnCiL6gJeS277Zw/6LRmEshJ//TBPG1uM1Rbzynrv10j8RhIV
5DZjtnKoznc+5o6BPpLUcU1Ka+gp6HZ8/0yllz+j5vpph/IuW9UKVJpU6V9vp+gbhUbn5aGXX4ep
NoxtqS2T4W1pTN1b2ZPvGBRRk5kFebcvClZK+a/hI5hqaFYmGP/jhUQqEVQoD7R81PvMWUFARIsi
XLw3xdTKsNA34HGLo3fRO9BP352PUsrVjkX0XrlSgKGCnsqpSdNuOW2LWBtW2AOU6a+Z1ywbJYno
n8Er1F+BeijBsq4blvSMB2MNOU5RcJmdLdhoOXSkCrEVJZAnlf2epfTg3dBZOxBAJseal8I243Cs
6iy83HzFGNnMyY+a+pMla7t446Mzs8NrsbBTLIkFQ15zUC44+8AcQm2VKcNrx/nzkfeenptTtzOV
7ZxrQiSYC/XA3rgmCUwRFbCkV808AhLBNTESRxKMRHe3P1nqNrbeaS9/QMiJt1tobziED/aO45LH
DyGLGG6XCI3Ukwiko1g8lQbaHnZ5/ziMLimxtSEveSCiUJOk4zg80VTsI1PpBHCFcAfRxoSUM0sI
+OxuIT9YOXu9HaJFdTSwRP6MPNTIA0pLjaD/UVDJsEtMsLYeQQnbm8WAwqv1AQkuWmVHGRhtae9d
Yo3BTnOea1WbYcdFR2w8uF3tYc5VSZ6fSajVANaX3IQumt8c6mg0NBaXL8Q3iESWXOgw1p8dZE2J
cLkiWfCgNX1AAqDIWGKYOV3m5yDVXMG/3unUew42E0fL4DT7NJfjmgdb1M9KRxJXOBk1H7GXRfIA
MzC+wriSjfB2qofE4M6GbkHSvBUslscchASrH+poY4hXmlWWzxKqmQvviZKFRxv9x2BRiEkrwE09
S7ksg3Xit0YPwMdf/kKYeGnnWURtC/6vuq+QY4BP5XwACdppubvrUymhoCrO1eYZhDAlESkbnNLS
jCxjWzjLJY205DXKX1OKIIVc7nV0FoMcfCcubVtVots2ymLgx53tRFT0LjOs0yzHytmXZ53tITS9
Y+2ej0oGyj3TRbuxIXedU9BlmuiEtSulf+wi+NMKzyrJVzrzX+2HL4BhOxropWouwU4DVodkumf9
CDLq1i4r7PxFX6RMQntu08zLjbJ0vxxv2O31wxFWqUySyhFyq2kOmd5qMhYXUxCawFZ7L+Rlb+y7
Uyr3lle12AhULonYpN2MZcLFG8g8Ozcba4Zld3JukVS+5NlNUmfsG50xLGp/0iomdIP4BF5IisT8
4XfvvfJWtLuZbOQDC1aA6mfdTVtACL6TJm+UcjmrBZ8N2volaVBP5OrYCMkYLSODVTyK5PxGxXVc
lC63sV33HSyRe5ZuxGMy6I/nd9vdPbkZGT6xsEJyn/EByhUZesoqPG1f/vnkYhGfc91IBhXUCOES
ZKD5XnGW3BcqHb6eJH+vIa/rWCxLYHuAEp4BpL0yMHRiGmel0F6WcmFrv3cLu4CuAaybBmcyDlqT
8PUNDihUDktW3xLmZGggCcAfjfteVAYJmkLaXX1UmRivWQj9miWXdYBd0/CMCtHFn5EpgUim7GB1
aNUgFFepyu4O5mzWHG3dbfl5hgTjSjwFYXc4LxhIsJiiK/LIjvhQVqPoP6qG97Ev5hQQEChquH59
2J1zaKHPhfou7KHeJrppHdkqLtqnRAOrAkhjHfXfGbCtSUCKFjgLjILKjWULUXHrZI245BtPlQKb
qhHVh7GtPJbREO6jWNA+Z7hN7IywSpbJ8vXhKHmiNSfyCJ221Zjg9QTrVAeG5LfvHrHMw5Q1oGZf
ZrXWbO3kKCJKSWd9trco+0qDruajUrhLTabdrMsclTldgto/BNeS2JqQMCsjWJ5dC10pUOwK5i0o
ybscsLNKc0bDr7bgc1eHI+RcV68ONPkGefgoZNW757S1WfpkSkO6KJ6rgmeiVCHL4h7p7zU8e249
uwMQwtkZDEA3A6g//HKm3ls3Lm9/d0iBVRU28B2p9RauDqVS/SwnhMTe8wVNga1cwsSXfxo7TjoV
s1FnWSIGHNbqTi7JjZMgnNr+lP7d3WT0IJF9X5Za8uxXx/9RTRjCqxCIz7ai/6wtzfc96g45m31s
u+gmFSmF2VZxZRtq5VHUCyRX4ZC2yJKpW7GmTZLrQmhhQfXGcDNhVbblDeDljZBAzpy3WzQTy9HO
+qBPPkhVZXkeejOdG6zGwNOsHD24rhpInkYW0W5QQAqr/jD2tTU0ZMquH01WvVqu/p4FQY38zEDH
ITWp3SUi3aAbA4U4Q9HeAldfZG/sy4Ity8yWtORCoIOA01wWYPdDK0iYEshnryoPxX3UWgpNlNLR
Ewxm2aCgDD0hM5XwmHj0daD7D3EVEx6jWtlaKivfNxXlufLJj7yKthhUSThmIobjVXingD+3Wu9T
xQcNY3sNOeNjKu/CujFR0NAc/jSl0K+COoKAmUmMAXjZc+KV2/SltAUap2Yp3Bzq6aeTNf/dQ9qU
TQOMpqzJkYO4uu54TOKdyxGah5eI+dlwzdl/IhnyQz2cYM9ke7d0E3ts+zGQt+Eue5tk0wLgtqNB
DvN1HbEDLyX1h6H+gXc9Vja0NJD6WZX5rDCOMd4/tt0qjAEeBc+A9LD8D9SyfXDD3Smac5mNygTi
c2PwTjxVVN7js2Ebay7Uo5DFvl4+JQ5yP0keHjXHPKmxJZkZFJzTEonJki10v6/TVhmNcJ+B/fYs
ko/XgzuMGHOUzCFjxFcjxpHv3Np+yLUqIkrjR+P43LD+GUwExorO58VdN0zZbb598fZuCeszy7B5
bfhYeQ6H95+e3oWjFC1Abu66MjdX1n9O3/HD3PhBPP/D4lagy+qJG33SBz7gA4utO3hwOR4wZr2B
QDQuaSczMokq+WWq9bIm5ED6yp5gwVOKF+Az35he0uSXTM0qNiWCtZTsl1GQt4+7P7fqnyUE74Xn
3y2X9SWGZMCN6heojp7tabik19VZxPCUh68ywIrcFttUWXipaeYiNjzrkqKi+MSLIKl1SvOpuR/v
dm7N2ZfH5e/ikbNKbkleb82lTVVRydINmvMdrsP+ZrB0e86NQzWPua2ZOVloBw09PgBHyVdWa8rv
HyWwQU1009cJOmPt5dd+CLpTp/0ZRGWnNpJPNKm+C1p7j6qISL7kGlmYm9d2VK4b933cyU8L/O3s
RkbLeog8s9TJ4IW4Qz4ti/IXU8j7BF/5XSvnQVY/vRS/oCNhC20WAJszsEOd0ija01oIOfY3BGet
bAorEtjhdWtYYyK/amuHEGwU2TT+Tz1HTZpBS3kXyveNrUWqW04Ed1br0NI9MK4TONg1/9dPv5ys
nuE69Z2FyqbgaGjTKxF3EvOERXubAXT8mo6eYZs/pcwX4VWaQQi5tWXru4HQYThsUWCal3vyeCdL
n6bzQMtRtENW88dkiV9ja8y23iPfJGLwnRXfzLA7lJK15eUB0KXkEpj7fONylno+uuiXclbGz10J
LR4ZSoeXWwvAHy2WPCT3s1SiiTu6OIz0uPECNlehYU8ojuGtMimi0FO0zyfw02z/sH5dBVi7LVWV
SKbNNA2CaiO7vrYYX6/jTeSdum6SL1RmtTArVy3Rv85eVIU/kFQWlLmxIVQu8xD7XCnVnzgONPM2
aO7skY9jXMm1PH32djZWaTwYLvH2uEjXq2taokJv6XhL/4AryfxQdMvVndVnCJfxlDsJTr8UnjXj
aPmA6O39qZ4U9mrxvXbBBW/39CQ3pixoyC6LXBLbWEHlgMXA2zKw6bPQDbkceGzwfX2e8wESww7C
pJ6pEWxwMPNRWAXnDe4O2IGQ+vjPGpVRJ4ePc8/7PtPlADVPLQCbPumo48Nf0P6t59TcFu986JVd
SZ+8doTOIMfljx/MHILiW3lOhzrYhA4uLeD84CV3wcZlQW3z1jhj0CuOD4yDOA+BCSFel5aydqFj
YEo8s8OPXkzqyBRTMRJMg7dwo6WaBOwW1OCAKBZYPH62BmPU1MsqYgCQLeCasVXr/3rV6yS3kjY7
L9x4nMGc8dgi24TkLaNz41/btVQftoQSKyiPlrWOaqB7G2ekttn92b+lDClXyMB9INmATSWULrye
4OzzQdE42Ol7ASRITVfT3sX03P6HlVQ//OWeeQOxmxGpFf/9WjAPS06CjZvQr7nkWs//fPjus2u1
iCD1B4cP0xLmM8QDdDOiS1M9WHCMLVLRG67DezaNZz7lYp9FmcMSHJshsW18ua4uoyfu24X72idG
1ekNJ0frP/XTG4vDNEHqv/E0YaZvi7W4Gpk8MXzarxfFCnhoFRjFOmLmuffKjpq9KLZP1cpd6NyV
2fZi/ctr3GAwFlHE2CjT77id3N4kLhtM8JfqR5ElAL5UlZ0rRb9ufVkbGmmBW2oqUD02C4qwvjXM
Q1YIEZ61sYrOQ4Dc7zxY6RoPBkt2rheurP4XN2sBEh2vTE5ldZSbiGMcwQaTXz3x3kusl8SbH8eD
PA1qptepOcO5L2Z8FHA/+v0Y1CdFe/z9Cxx8VS+aaSH1MjsrobK9oXq61RCn/SwfNj3/QTNjtIQq
4bLfPLrSnw2uvPQKaC1hECiDRFqxg8EFRYvDYO6tB89i30BvefUvlcpIaK34wlrL1G5DUSLOY4tF
mrOeOkm3VgxXXIYM0bGX0O8GDznJSvpUp0IhWU5UC2qT47Jciabermn+dVJ9TKcGhOZBc17rahKA
kZ2c5J83R+AHoOHLiJ2DhcFPgo52ZA5rUwm2hBaE+95z9jWhp/52IHGIo5o7hrOjMlX1ZpASNRui
erCPQChSqP6u9R/OzmDxveayOzYXAznKRTOHpvsXX1SxuyxlGuCXfgHq0uW9xIrWLw3U0EQiQ+dG
ayCzqtmhrbxBm14xJb5SDU+fk7TTNDmtHLsY18GWMSzw+VGXk5hLK5fxL+4l/QGkf3Wn5u0Ob2jf
YWXZZa9Bm6Ep36GqsV7N/Yh+WVPDgXND+h1+g6QBmsDrmBz/B243KWVMgTBgNcAp2PL+oLrrQpMU
esQ+YCINkANVA0/9mGALNQ3mfjyfT/nPQHwMtbdo7W1OS8rTNCCZ8Jn8Dnc+aSsoVqXfJNAT0CQ7
eSHv8f1Kk+j2ha1q3FH3Kdmye0gWjiajetKkwLuj0SpGqmeCWoMycFI6sdipw+4eLArBpdOArVvN
0srKwUk8EEyt5i24jedVA58HfIP0tj6HVThDOia4de8w70DdPnUgpuoMQiA4gxCsxyQlvryDDd7w
gPqSCqF3NKJKfJKnw6nsfDRleAYnYA/n1x8i4Yq+ZCwSfNRQC4OBN19Z/r06y+HSs/IIQPasVMk1
wNZ8Lv35Ov/faWBZAsyWQURzDjFiFPEiGDmmaZi9r7BX/J1Wn22SaZvSph47TjXfk6xFhoL5nv9h
YcluS2kGo7rIgXO1VKaICOsnFqtlc1EsAAu1dHiI6oHJLAB3+Q0R7epytSzGiiUa0WCJRvCQmige
PgISslxMFoVtGZgnxO80VunpXea8IEmH+0VEHB0y+tAkQTHITjmaPf8br0GYhs24bvaqz1qrNyZb
UWi8i4BFEOgR8x34JA8IoK+xDQqh/daPCs0tYgPvPWTx0g0udRVFRZOA46HlTYLIQV3/QBKnUa7E
UG3zHvWWsIQVVsyVm8BiboRgHyoEItM+bGX8d+Uz2tI8OaeaOjLGNkGuitr8Bbo3SIwwPtyHg0Py
XkW0tS4M4OBLmewDDDmouV7iJDhFSyrxRio+VuTbeUo7tpPbD8eKxYMII3Fp0//uiphTI+hJjHJR
s2TnPuR+ss4pOR+G0F/GMvCQFGajwZr6iDjCHzlAnVCyk/8ReLCCOMX8c3cDduRhE8GnxxOkbTK9
swOCm+TaHbVZoIjdwTovau5IHP0hnj9GwC1FfF8UzqGk+SyVcsa4Vsqk0LkGYMCyqm2Tv55svnlb
oedcX+xw4DQCSUyAZjiW5tWEhf+KUlg/EioqJXOvNv6vHvKpchSTjJajiqNJI86fUGNLPqf13A33
mPcpg0qy6Ux/kTadMJ0Pa4n9B0yKUc2+hYatww26x/PljdscwtqLkmtdi5iJm9UU1XVtlZsNqE6e
Z2eRtD9UzZbo+J2byfZANRz/xSs2KK7vs3lus53mc3mmi5o4cRgqPUr0QMoTTJt5S85nS7N7OLls
0TikbKD/LvYRt141QfCBKMy30ComxBFhNZYY3N+BTDCOQRbtyCH7QfXwyWyMRRKeHV72krhW566H
3hZ3xPjKtQ7o6d67gIsvASdydpKzFgb7ly2toDA6v9GY2UvYsgCDPB5yKTV57BnySf3pU4zFamP6
5Mp293KZr9tF0HmGPt/IXS07Wz7te853NAN/awcM6v46clqYLDm4m9Mr6fhJ2Ew1yHBrf7eYRN1+
8P5Q0Q0SF2LNTXJvPO6dX+GSwvWUKvvG1uvGl+0ktI+sJA5DR61zpcNJxWiPy+jr5efOVaP3VIlF
YAAX6BnD/0aAX/sB4urhZjBb/MI6KnViJ25IdcTFse25xY1U+Y+X+KNyoAV/MCNavIicI3E/4jn1
nS1tPSWDkUNm3sQV4JNqVjsyK1Td8J4BTx+BD5Hrb0hgOc9STDtYR9lLez8BqvPcGC3nfA+r7Rts
Mj1yckSmiskJ0lEjLCyrksdmwa0Cfbnj3g4F3JbJAJd+VLuNeiMT7ZdyxXwJqj/TIG32DgriP/Yf
ym3e/tDbeHjr0rra82dTAufff/mF6A+7xh0vAmnk65HlZzp33Dsl/9cpqvuChtB5KHDI52U+BqLs
rIORRP4p/Wmuurk0ePTJueMhnusvvUHKGgh2wdQZ8Q/a6uEe+oF65MmSQ7dehL3dT0Qn7L0/R+7q
VZg4z9rdxylYd6Z4PYRtxxo818RPDhIpgAMT611Ug0lodz/Bw8yXfOPiZTsG5uoa0nmKNpZ6db5i
cRMw4L7Kz0Xv6YwlQkYiGRNiiw4sIC91GqxKNUV8oEcJ746+Ha2Uq8FK9prFfy3AxkOO9vmys5wf
TibpzoBBOHvpFejxZVZygwUE0zX8s0wjW17CnYfwlPulGtzqrQ+wPMWF9oqQqdpdvg8Jl34aSsK3
ZKq+PUZUZ9KcQR5WGclgsM6cgXlOn8qG3/e/wGTsFPiZofTE8Me0F+qnD1XQZ7loVM0Fbcermfuh
ovelAgADOnZYf2R+T1j2YoAcwtkTXhQ7qyNtc/nVY/lAhDnW/HCsp41tU/euk/1qR5g16OVJtcwk
LLP8sdUiW39wPPa+DTx/AgxMM0yexfAj3PH1URw0Csc9r8sCPVLRPwT4TFBRqlabot1/NiSPC67j
S8ykmPW4Z+2+4gYO9ZxjAEoZLHBFZXMonhQqhCz2fxNbDyLWwIDRcvZS1yIw5AonZvNd4V0YC4jV
9qCrrAcLdsED3tipAQQNcz3dU9la+zbBmWGMqUTVzBPZIPx4KGvKbEhC3F49eTl9+rlW8DJz9fnC
rjXyTCp/Scb4uHYs8lOOLPePjqBSjYS1FXlaH7XVzOLBQ5b3+NMZRXPoSPC/egb54Blsp9+j/tu8
yiuU5FErgnuXQHssQm/Wbrqa6Lv80mPtzs725/IN7WLnIZSfLTCRXb0lh9UTMaATgwaF+h/+ZZqJ
lGFk3BlsFDcH7hxxe5wxzTdbeC1HoZWVUzYGaUi+X6IZBZBlPI8=
`protect end_protected
