-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
hKu4Si0xLFZR5LIWn8nzrbDWETGpHTfLQXY1ShXGaU69XStjd6A4u9+3RJszDiuWkEwo4DD93X1f
8YX8E8sSyUGZMWqrWppN34VuDxu3J93a92Rykj02FpVznNhu0wYEEoRqZbpmzLdjyKKHl+T/mnFZ
UlRUukuJ01oPSpiMnJ+5LUmQhl53qNrLfrMt1xdJfpLe4NVDwoMTcDuQGydctgU0akEFJKKQpH7Y
GfUAWO8u7QOXiEKQb+yRlXE9URXOxrXdW95uWQ5KG1yhIUUl73GdVinQjQ+bV02soNqT0AeOp7Ko
e+LZqe0YTIZa3eZTaECZdxruycMaELFzJ2708A==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6256)
`protect data_block
+wUUip8eEwdh+umJSG7c+h7HCFoIKfP4iPWz0XGWBQGSCZ8Yb0h0+eHbOCbONqXFESbrsmVpHPJd
nF5YLA1q58z/u7YLNp4Wk8pqZNQVbXvwNHea5cd9ZKFOem/yZNdcGsUBhiWdcsm0z1KaB6h7lkVR
mns74q5xZ++Lt558TR8l+s5i/MlXLb9smhDEnm84sIuWOcIJzyUi1hn1G/55uIwfcrVxluEpwOJ/
5pqEm/b3cdbYTI5PneNGQ6zxCrUsQYZ1pwJBe0NvspMYOn5SG3CWyGxmuQ8XhH+YIw2wRxlL6RtS
uqgnhFqagSeWYqISBSyfAoxwOdZHyrTrwsL0cGQZ7BszfMppWRl1BEhWYjK/p10JWi3znTKZiQ38
p+G+CvJTMVo1yPrC8He44GxuXjyMdDmybmBc72bTAUcZZ3xJ7BbSWVeP59Sc8DQNajPhPA7gkMpH
EXaRGk78qCvc497FQcI1B7eT8I9qTnCG6gJDSQ/RH6rIHR9+Ix3qkgdPd4Q8nAdrlSv7xVe7h3SE
bsF86ARcEng+/bJ9WgpS0BVaByA4En29Tk3DGwYsRn1GyNZu+en7JzmzYdiHR1dO/y8Bp01BquP1
EFop/QIbKWs4s9R0rdPA3uqBF+s5u3LF68d7/rtEBvaapL3DOI2YLN4MPhhapEN1HsCPo9wiA34Y
Tyx8cYX0jO5biP3VglqDupuBXmEsbNjhmkoz1EOb9VphLMX6qYn+bzyOPpNjAagduaJa0a3Y5mBb
8i2MchV1vHUh/riPVlljzHgkOzmgVyq7KEj+N5g8UNSJ6jhqWwnwblDf8vKOhg83HKyZ5FXOK/E7
XdCJOqNpcuNN+PIaVMyy0Luk0QwFf5uTcUM3qAdVq+jRI1PWLSkXnfaRpAk1CwVYxtBlIBX84Utl
JfxXXYTBmlAdgRT7nXGF6rBLV/1jkN2voI1OIQ7YC+nm8hUqYX1QF/YTGeMaJInDlJE47WPGSIeb
vo4cXGiJZntuabV/0uNvJduudgOEHe4eQKgru3THEfrz8NbTPC7hIaadSVqE0ruwr4SATjJvaM2R
128glaYS8X+4t1Pt8wtXZAsOZfmusbh10igzRjJTIKOaTDtkSbKdXNEGqCB5PIntyp2ucxMxj2Ij
v2LeX5Iu544E1UffgkICm66R6O0T5mBJuF244u5bumtHh73YhskCaD+SEQVjzxibh+Dy11krDVcq
ph2Q5Qr8LkVMWy6lMjmxqMC5GPwjAkKB9VThxmmpV+fQJGbjIkvkXix0sJgfqBpgAjeU1Ba0W6Y4
/ykVu/feoVOKmgurNO53v5ZxN5rR4ucmlDcSjIWCuxS4/VrrnAVhbr8bHdQ8iUb11Thx3IusNCS7
voX9NjBBmxnicHRfbsUtkM3zjM9GFQlRD+ug7mp3QV4j2pX+3hNsQvCA8+XMU8CtZwcUvqQ5o6Zk
2RkhYQqgL8ln0oBSpoYgHXsNLTO+d6TRMJPWEsnl8mYRfp/FcupsSWVM57aF8xkSMfDVsb3nA8sS
lqxsdqzEBWd/LRVTv4U+fTGrx7Q0ifSATppTTF2sSCd6q6UoG8rG7BekrMwW3mCVpnddWT3VEcD2
/2vtHjjw1jBBGECBtow3XLbXFWplb+I51oxtO6uzQAk1ZwMOl38a9zFWCYADWpuqK1hkQcRg+GPw
S0pDhkzd1y8dmlS8R8wIhh3AohH5R0Gy68LWxhbf1rl74E3qni2H3Lu+HJhZ7cSKcU+g9iuA1SfA
nyj1eWl6HPsff23zRyAP6wdlyrSuhJYzQM5bsdHJJJFsk5kB8T3fuTykdMgfqhfR6lO6Famornqy
RvSS16CkEouJoBbHOsZPklTLNs3XSSsR4OXnK2S/sJb1BeT45TBwLN5r+rUdNGYohSi4qF1S+Rjf
rhBzqcuq9Yok9I28AMgtwIetrCP+T96+1X5H57Kd3qKKUj3C6zFpic2nVrD/UBL89c8biLlvfoe4
gRbwoBzL6VYzOlK6ka8jU3PLxGfs1Bnj0WGxoomhK12LlyxT1tQDxJ+cHohOOfCNGse44YyHjtqJ
o6AMnUOulxBhlmQ5K+/542b29YJRrC8YWhwwt4/vfKIjLpiiz2mntOSA4coAYoemqYoUSwDoS1Pe
sVUfdWbFiQZIwfQjtrRJlSrgKfWgniPN1jKuNuIfa2wcNINbaGavsYw+8BKiZJePYBlUhC/1v3Sd
5zfKuEpCNYi5I0sIhDTLb+nimAvG5afg4s8ZKxS6PRATEmJ+7m6tjLKkixAkp1QTGMSqH8IwqyLM
JFkqzWwy+xlH1wBlan2zPftAbAKzCOnHJrz6Z7al6bkrhP4pZX1h2pNh3Ksos0KtaXKyBrjddObM
H8SrkPLtwmCPaQXxmObVSuYTa4ew5OOWPsBHxbElY/z9E+A4CDdzIGWHt30KQfQJzexkyA/gEr3p
8sr/Y/H31NE+MxtySodYd7p8gptXWpofYl7IRk0giGAicGJGhr5dTsA1olP5LqKwpX8DNhcBSjRq
cEvWofYpHfmR9RrABtGDxjCj+dkWPYMsPVhKQQkeY1treO7/vbATzeCkCa0TwGYuaMr/vYCU3Iad
isvDDQ0OC2hWkVuEwN8zvI9pm9NUCb1b1PnRuaSDIM3vaPvz9MbQLlJ1PyzVHcOQF0ioskS0BZ6D
2aS5ek4RdG5CtBeqnOAi+zfcfWV2b+QrnUr5uzBW20GljlsVUvtst/FMCt4UFrLwl6pPqWDo8AFh
DP9qM5x6nE5NQMlUMxpHd/lq+cHTBs22CMBPTua4r1/ERjLm21VtoRR+wnEGqyGaqTUfAEkNaznp
BWaOFqLCLjLj7ePUHBc495TBiGLGpo0W8NdkOEs7IeMpKw5MN97kkfR96Ql3UohbxKtr8OVb2rOx
G1lJ+rhrfp3ZDSLuw2ZUJ35RAqWg+URe8Lf8kasKoAUIPIFXPHb4Sbr3hzP1xeYkIsks2xH/wqtR
L0j0V4teWMB3omZvhhd473gJXWNyIxOa1DgbAI4MjlSaLR2dWIy1zjOYc3henIwZpHmNYuhNJ3CH
TrBdTx6ZUJDF2orTNc/IQcqLFxBbVOvjyQRHVC4+4CjZs88p0P+5wyd76+EY7LKj5rxH6Csz8swr
gflv5cRRUMcOW+qc3239gsyQM4Gmuw9nvOnA/ca1lAT6LMnJznmj/52Ul4EjUQdwfPMB0olKB+Nc
QOmUi6wZmGDUh6dJlzSrratRD058M33jojciIAub0NfijtZHc4urwNUyIWN9Q+1wDd2i4IMUR09s
+/mZ5N0M96scio35tnZSrKqXiRn0t2RAH413iecpcPFBSdbrNwvyN7+naUMqjckuCiXgUZCcFaFE
oWenmcD0/h0+/gnzKEvpvleXQpJ1jnlohVXaT01cWxViAcJSuez3sBu+4Jf6xVqoz984yuREkA/+
S9WuyYqGtuui5Ro3kaarSxpnCQVEMaxrTlyWxFSDITb9QFPcqC66u5qU13RQi9JqkDA8MZDq6yIf
fpYi6V0PLb+WSuVlV2UwfNehNJfvbikpQhGhW2AppO2fA07FQdK63y5NYGRLOQCRF4ji4mX1u/rM
Aedb2DK2jUasopbFzv+ceQO9nP5V/8CcGJjgdgu0SeeDwmCoryKQS6VMuf/jYYnRrP9PekKzNQ/h
v2NcZbU/F1wyXhMUrVJce66J9XQPH+WjJtGKn4wwHfo2EHVNLxOoF2A08wPI20Pi+juqgNVI5NBR
zIoSPttpBIm1fmUTygBjC/IT0W2Fgo1oDzIwTHnAPi+9QoW561G1jPQIsloWQZ0kQGHAi2dqFeZI
IHcjYAn3F7osJH0EQsNuOv8xe2pCQj8Byd6m+m2l2KQCYT/e2otqBMU73R6QgCrcbH3Z/a4vJWsH
dfuh3fReGs7ksxIXKCuWUYGoVgimlUOZxVeZtE10k81j9k3qx8AGTQ82hz7iiyTbXG6Mli2nZ7lf
EgrL3m/mODZVMJg1NRtdyRLtreYqhCKk+xQlRDXBqEouFb/yt44VBTOqCTrVRi6OGZBQqUOipoXc
2LCnVEgKlmX+RaR5kSGkrSTJWtl1/UwChxnTM2eiyqUeBP27UyXWx3oYLnAG1b7JlhFRk7uOtklA
oOEeDWob8lMy/iR3/W3md1fI4GMRH5zAB9CaXOKGzFNH49GcE76hOUzHUpryO1qP+cVXzF0vMQSn
PdjEPDOnacHHfKlqGhCTwlamlfzr4NqoJ0heQBCH8MpKk47T1K++ghyBFJR8GL8Wvoj9RYaWmUAQ
hLvzwB6Xqp0X95bNiaiNzhQNNbdYuwLPqa2tgq8JyKfSsg/E+JmGOfKsX3zy+fE6TFxt5GBlQ7zH
VbAzfo8zWnIWbk0o8KfK+bRNsZ+nmUE1ONhxJUGbc+ZZtF4hR4KAbZMxgbhGFvoWXodX8edBnynw
AaYr61ptTBdfmNh4sd0gBukMVZSbJzLE2FO+Jk/OBTS8F26L6UOqH67bCnLoJ5eVtwJ4rF1RfImg
ovKidyVhT5BrdSwquPfHR+WnAd9HCaTrys/glf3JjvIgsbutMlSO5qczWfOUAOLs9OZZbtA+wcBf
/HjP4dmXKXTFhRXPXkjOGpkmObscuMt4F7YOuDepjh2G2SjjN/I2FFzNeLGYQ1XZN3WN/Re5iChB
gpqvZMWA/lv+AAOHlNMEej40jLYpIb6wwanvOUDk61SOK8uB3n5PH//QVIWtnewTkkY6EAyboobf
lwp9un9vDs0UKgSt/BZFrO+ZKQYD3zS5b3PEGJ2ZWdo/P/VCHvwAOD8mgpP7iGk66LZuYp+NzY+n
+rLWhL3MNPSowkMxBANyIb1xRZxj6ltMkhAsfGtwS8A/wvRAfM6J0sGDEaAHQqxprkM739iOtiy5
3F+qm4d8HPCsaiAg4b9u3eFkYPA4Ifaro3A9BoBQLzgDdDCbDnRwPW4vWPXws/yeiL0PqBn4NiHu
uHoLFl81MI8TFnkzaMCJFDOAPerb/k1Zd3QvaeMrxU7ojuu5v6mX75pMu8J1IhHnDnxg3czdyGGu
AHSvF8Ano6BdvtBdM+Ba+9rEk6I8xi8yxIb+aXnitdCsr3BjgM0RaHbOOLjAoJOmsPebnpHwq5n/
691jOIyqssL9M8z071c4+Ei1Y0iSvdSa+UVFBY96yPTq7sCg57dmzhx6xI0oxrKb5/pcT3jl+bgC
FKBRF0DWUJZYDIu9SptZnLbj1c/mKgfA7Y59UowcoTByxxC7TrCEkwyK4DrahKPS9toCpnHPLMIQ
0MyI0lfdaoBYxcrHzt4EUUekWWlQSKdwXaeUVHopkRSFqYrns2RvVj0hZIW9h1stoIORQPH18Y5P
18FHBDbSItjBY8X7a7zW/IVwZtgBicuSL5p2mrFaGNCCR7yF1+q9ebXH7OowWsU8iqRzR0u+qz9O
h0EL+WmnP5opZRzGJ2ji+54Q+V3QnXfUxpvaPcdIHD7dHwJxJCEN2lGIEFns3kYCdZ3nK1ALoZ5P
WLNapSxPDYogFMffKDWv5xvAwtvQ8wmMfjw1o/NkNOfItjgh/TWdVryMHTCHRJp0Lplcw7uCog/W
dzoRNvtacswn7decA8u4+h+jl5Z1Xd6JQnlsns+SAbFNVFGS5PNauA7VgqCSU9P6LWjY2bb2zf0R
af+A8LcB7lY/gTKgkjqOKM6RL/zOP7a20uVcNi9U08Cw+qixTfrf2sNT/1uynOu7bDWajBpyqSXh
g6sVWkBR6nJx+18wIbQ2UQ6QuG5wDZnmc4Znm+Eg+hHdeReCYCIpCaWj5De9Ih+O2IO1+0HEMXEh
lBKLNP00iz4PKuXTgLFggnH+IRJbikf04aRrOUgpvYb6zqgt1XyDCUQksSBy7u2IkTGuWxcViuV2
3gnzgLKFAx6linEtl6A4g8pZB5E97lgB7xT9eDsNJu4ER/SEk4ELmpMMvRY1KEffaQ+jzYzFT11N
R5fB5hRzag9YOrALdwCNCr7o4jy7Up2/2FtWT4jlXGZk1mrkjlGMyEfga+2JRB185I87JpbyLJW6
JllxgGit+RPNGaSGbfpPjYfdE5j2wUYIteQYj6rwSc2a3Yk6q1mUBhOI78GIfYCH+2RbIUbvayer
+uxhqlqEWQtCNqnKa0QAZ5aL2BANhp+G5nIsxEhCrP0mTOhgPwALLN8HulHz+Ui4CD3BY53tanXP
21DSYU8qyV41wWjMa3oecaLbzv4XdtF+U/fX0hYiC7yYTF8KCHfFU4kgENNMrxgyTsDn8hn2hiW2
G5bOiTmmpMhmMknTCyfQ/fFBxdMpKy47ODiz6t6vhSFxIsUVcw2i7FDrCXnBYZQuzIc9zg5kxP3C
/kRU106iZU+dohRhWPz83tyWf33ZgR8/dHXgnexRNWlZy5YTJ/600T5kYIIFvkWRFhBxLEvvCJD4
FDrlY86RDGSPJbRTfdnKpEJZ6APN56QhagbBSEP187zhfvGoXBtcbF9SeCoBO0KRomWgoajfWjEF
7HbS1BBoudN87x/xXyDARtf/kWQRYLFpLGLwm/+42O+yD/iVrc6+6gneA/L1zTT2niL+YcG+g2QP
ClQOqx/NSuFRb8pJK5bbi1qYyyaaP4Y4HQntQxqvJvT9gPN0ZeYCZV5NQHpZk9AGK2lWUSyjtekn
BO/szghBICQTxjdjq9fIV6KBwoEYVFIdKkJfJf3+xFL1Ev667LCM2D6XPUCsoPOfWXcVajCyfcT9
fvNvXjqz8L1ofC26mwE0YYDhyFfR8lDEiq98J2Lgm05gR6ICULrXByxnK6RgFD74OIQ6k4KPy2Fl
5CNkldRRfSJEYuPT9LovfhN/ZdewwIgAGqB61J/F1UkagICi+OtXNsjP7JKdd7h6nj3SZqHnAXmS
TPsNO4UZMPbAfF4C3EhNxoSThPtu/pdOA3hu6RSPeC2/k8zM+y9Wa0FS/ngvC3cFcJ6Nia6ZndK3
qrytpuqSTt8hbbR6Co3Z2JkEYditI8FKvtt4PizlCgQRFECGEcSk91Ki3gt0KTrvmrVKWWXzPtUa
2m1nKq6kmXFJUEfyJA0f83B9yKIj3jhrrTcW9uz/ZPt3F/62q1hI1b0/oVpxbbzw52Gh1MOzpfgA
KqXUyjhD1Ssf7ODmYBsYdR7ZnfDXptc4DyTX9xoveek/BPHg+tKfRGmwzOEY8/+uv6njAc3q/STn
BCHxZH+MMGehA0IdSyPCgh/C7evGbsEzwekP3KGm0s+U2bcdURKgbvy9f48eshzM8uXsHDqwMyIr
k/4EWCNvImMvSKDbiyKBzmIJsKOna+lIblJv1/oxqSMKqaWsmgmCMJSLtD+6ppXgE2/0Qcnj/N1z
PSIegX4FqlTTTkdXKDokk6agXG66yatWCEngKOznS+RAeRxz1F9j1z3ynilN1iM05cIY/s9QEOxk
YIwHlBQB7FgfIIpx6YadPZZykOrdy3/2vfehEmjfaGNYmEtSOhTDjbMw94cJjq2CofOpeuth0OUY
y1dp6ovi6HX9mez6D1CCTqHhQxK9t7ruJLpJDj49XxD3f2JR5CfjoJkgEcV78T1NDY6PiyzyfzbO
JTsgtzmwanFFFKMq4npYVjjEvbT2c/B18nUjSoqi9vM/8CQX0/VRRwDHc2miZkLXdQpauS3tXEDd
RSV/qvya/bcf9WEKW73hGZYdi3pUHctVWGf7CIvuueHXj7EMV0UTgKH8dtC+Cf9Hs4dZiWA4Wnwy
F9WeUFzeJY+eUJ4XoFVNbarkzSdA27fArHbLyvrNfto/Gt7TdANb25b/WnlYcVBAmeUupGbykGD1
h2NOgeX8vEw16cKjPX0mSyNSgvWMKdiSMH8HIRE5lkmnJhfJo9h4sZKFfeEuDEcza//ppidhpU2k
uqiZEluS4n1Tw5/SfTgzeFWKYT4TZGmO20/Wv5PxEhO41ztr8B+yj4noRRHD8d0FJjA3cHaioRZu
bJt2MeIgr9R2DVC1xarIu5nXaAokttG5AOIoTD9jmDi9d3iInV3ssP2c8IpZ5NTtFKOX9amX5L67
ZQvEibIKU2UEDqQX3zuQXlQeZHi0O5h3w2o2PTK7aw4XVSIpOrQx0dec0MPlIBAVyJcKEIuqZncE
owljNv+zZXaqoxSx7HD96iO2SM92BcUnwTt5SbpqBSfNzgnnOsNd46BK9R0DJcyI6zwaVjWp8ZxC
DacdjhfTC2sf+dZnen7ECF/5qunR0E6+NKdhSEBdqASse83B3XrwjfnAH/zbCJY4DEHjkjHqxPUd
zeag4+Pq1d9JTTUltnUKtXBW6yIZaYAyinmiO+RqcD9gOylGT9UAITw+b2UrFe68tC1Z+vNvyeOo
Ybf7UGqycZLzOLu9l13w8etc4n2OBkFOh/llpIPjTsBlNdwKiy+JgxIAjg==
`protect end_protected
