��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$Rx�y�<��wA�*;�x���@�̦�W�X�fa�M-$u����n~�%���P�$��W��kYَ���P7�?UMfT��q�6�U��k�>����~�\N�(�����X�e���/6U|)�X2pF�]$h���d.���9E��WG��L�X"]�Ad����ľS���8od����e�GT?y	7�������ݵ�^��R�q^]�鍦�����s�ae���h��L��P_���ާ��YЭF���'\��68�b�[����w8�[X��V�F�0͘3����q諵�uW� �h�u\V�?@��_6G�_�*�G���B�絉�f������[�G��U&�����~�F��AׯK1�`c��[<��FY���4I� �#�G��x[X�=�Q1��`��R>(�w����R�O�?����7�,(�H\�#h(W�EH=�������yq��Ѿ��aF����:�U~m<|��.��0=�P/���4ǆ���T(������=G�چT���p��vxW�%��	������ ��v������M�;/�@?a�e�E�¬_�z�h��x."Y|�,��B��������^��g��Ux� � �T��g�ְ���A��ݦ;#VN/JN&�b:�����6�O=܄ a��xh�yYDQ=� ���nR��)��YT;���O-���4��Y3rD��n������sWý�Ǌ�*φ�) n�53����U J->%`�K~����t5j���t���Z��7��x2���ŸtH��.��������� >��)|����ގ½D2��3���G\q�U'E�I_��;�wrt)7R��zL�*���0��v$)�D��vM���(ʇ��0�I�s��:u�rߔ(>��As��"���*�g�$.JR.�����L��Jײ����ޫ�U�x�j�՚B���Z��
������:��7H�WA�`��`F��<Od�fk�ٖps��@�y��%`��~��̽�� ?����a���W�c[��alRo3���������V�b&��X�ະءĒ~)Z��AU��e`K.ʶ�1�9�$m�`��SN�4�����o�x'��/�� ���S*�h�RL�N\�־����OhW��G�j�L����Ё�oXg��G����L+����z}�_��}h��~G/�J(TD��"�Xh�%Ûf� ��v;rn�>Rn��@�>;$�]gE*"�=y�0pޥ�0�r�B�����#����3ΪZ�R�0�7銡��`��p:�"���:,�!�?A{�lo\ �䵵��������B�5�/vlhާׄ3_�.�I(�D�0�8j� 9�`�7q�9��ʰ���j$t�M�N��N|T����wΣ[]��r����'�โ�W�Q��]}wl�ٙCA�/�x��b� x�������oh�*��\�\�Oӿ�Q�x�S��]��,��T��ᇅ����F>����{�2�w� �_Mf!�<תd�;_J�zbK�
���'3�����uj�PH`��Mn������eb�`<UY �N����Y\oC�~NkU�*/Āc��Q�ac�� ���\�����e�i3v��B2��l�}ۨ��
��s�<0�t���U��q���Rj��%�S� �O=J()O8�_f�M~� ��%��\��iy����Czʍ��9=N*Ґ��Zu����	0b^�6�����y�ȅ��of̙s�9.�o�$#WZ>ȫ�Y�ξ?W�I%�c��I`��MA�9�蘚B>����E���8��O6�k;}��`��:�Z�H��y�d!�])]bh ����[l�p#��✥�Jʤ�!�_��SV�ME$��������kQ&<�z�jN�:�+;��ޔ��cIe��pD��B�_O�pYzK������K�ݏz�M���ԵJ�U���� �;~s������Q��N�ѹ7uVZ�%Y@�QN�`�h"�L���������;���_!����O��ɩ��E��$+V�E�����,��{m���5l�6a�U=A��&�caU��� �1��'�.��±��C�Խ�#���4��Վ4��sn�V�(������&5'�Z��|���\G��=I��&��� l���0[]�
q˄~د�t�R�N-�׫��[z3��RbM��7��J�3p����V��<ܼ �-��!��WR�D7�!�O(4#��Z��m��?��P6����� =|�lMS=�c�qKBͰp�t�j6��-|��[�ǹ�����!����!ܯٞ5��./���{<m� �{�,�㈠�r"��90<��