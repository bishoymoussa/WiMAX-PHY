-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
e7y/8IvruMiOtz2/f3MxHjPdm2daGGLt9yzncyJSNWtz7uqOJ80GMS6jQmXJjgAD5hzlWNj7b2T3
/L2A0M0JLie/Cw1ysa1o3/YGS97LjBvQ4/AZX0LOBmk47WUobrpV3zn6IS1qrTE1k/P9mcfn/5Rg
TjwyI6BqkFU0hh5GWpSrhRgL5xI7j0nj2LTekRBPpdbL7yFzk01HIxHxiCo79bF8DJ0CLUd923D9
vOTgdj+LF7x7SeEdChETAjwAQBP8Rrw77R8c8ZNFNaZZwIoMy/KY/umkSRvNUx8gAsmjUnw4q/Af
BoDaqpcZlTlW/9MB8arSwoQU2qT/uaBXm7mi9A==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 14656)
`protect data_block
aq9gZDauF2qyGNO/IOSoQ4F0kMdW1mq+xAJ3PZNwUerWmt9u134PZgqSecRxudrHHgb44C3f8/a8
1LqQy1YWqmKzcDE42PnCRVdOMUXOvyH4MKJmbMX0S9Yo9MLXO2GKYMBhXumjNiEWRTwueb7YBrxw
vksUlZ5iw3UXEp9zXcEO35TkOw8OzbHGaBIlu0SzjDdTfifvKuiIj6Zsqkm2vGQk4FlU0+DY/uyB
mH4E85HNjSM4MDNCiv9Ehfd7fMCX3Bi6vuWgHXFx1jckCQ/lMPaJWph4CAYYg+pM3Cjj1L7OAn2w
ttzonGL847uexwqTlQUGYpSKkeEKT1Fh20wIkCy9wPb9d4tBvmsJeS+0zvPX8ujYapFZfrM26jAX
hoJtJr12SyzhYIsWDSBRCVI7IXgqk3tckFjJO80npvzeyl8UHsXqAzAOCdFThecH5W91zWQXA4YI
iYu/BYROcK2+nGddomtnpOPylUqx8PZusv0A2ZKsD6bKdpHp0hK0SvLsv1rYemdrIkWdaJ340mYg
gv4Jxkh4dw0nhrXAz+F1pDWyFLiVBM7uZCLgNjTycI2l30ubtSb9dugCDg8aIaSMDDdqC7VpoYXO
jgFi7COugZ0LpdLXwqrfEGeEggzr944YXbji1/sEzNpW9+tMGBb9IITcW6zqsUFhlNiPXAQbsweb
xlHJ6S6knB2pG318ZlWvrAq52mYuoKYg+WA9OhFoP8CB84c50RRJ92ahYnA/h+epig1BId7MAGkp
aMyiJC+ByRr/yXyikeoDZs1D7UYVWlCmOTA2xGD4pGRyJhpelkfJMkM0qXkqzXf5HrhJdxFiVbyk
hpReUKHEdFTwzFchLDi81uSGDZM5V9aWYDS8rKW5zT0I1kYEM9O4WkvzskPe1JDJdNeUpcJy2NmV
shLGru7/zuX9RuN5bDK1QpLJZl7HCFWRqjH0KnZgQVOvBx9Wk2qn6z3Mb/dHZPcBi0oke1w4Uddq
gK21VPsjbeZzxccjwTQ+pOlsek1yymjYrakELMZEb1Vxsy+5bKi5bY4FXWZOpkxIhLzUmXKgTNoK
kIiRihXM/nrhGXW8APNoETNjlfi+Yus+a6pUwqqEUwMbZD0kT3r8J3rG1ZpmmBG1dxvwMDfovZ6I
C81uwjBwldrb4iiOPbUQufiFMSHQK0FqvuJB/jn1nl9apKQgcPgFTuCYN0rgMJeQv30lmN9K8eJJ
IGpbCKsmaDb//71o4tZE0643GSb+MPye4YdkFRaGpMPutZOdd5LdyO3ylnKxDBSTGFTPeeSAYr6u
Ih1fjvMvTrFh7rWpsBs1KB64Yb3luRinFEyNRvmIsrqoLgNIRCwA3XGn0O/pDxM4YZSUkRobw9WB
5GJHCFKOWKiQaEMSmJLhiW2obhbSSk8NgVkOcPYQgKRcHDUcfy/IMFqTAmSLAplqEPQJ9eiG/AVI
bc17YcKeKz2Xls2chQjP2eDCbzHEY1l/Iked9tB9qh37SeALveLtEDYpTX++6khKpDRADrwUZyw2
th/KcO/cjwcZKUAxDpKAXlPgakqAemKpSnJE3zNeuqPjeiucz9fNjG6PLgIXtB6p39hP1dW9uGNv
z5+J/KkWUQ93T9/CIfbkkoFEAh47jY7FmEQMRCSxuji3GyJ1f5JiPMMl8g+8QdbVxKXIQ2IDyBwq
DXZTBh58rUPIzmgdjZq7EszF3ChPPlqT6t4L3hBf7hxZRi7oBNesuJqQcVIB9NE3guQiZ6I8y7Vu
6Xc1V6TmIp+8I6Q31bVj88wxsTX7zAQ01D15QI3QDJ4UPZMVehfV3ydwudL1s+nPLotZn3IoW0y5
bdw17CY5l0Rf1NbrzFgsGzJWgMSqGoy9aKHcRSlf636q5wqKFWpNgC45FKZD/2/5foSJkkWmKhOn
2fQIu3XB/MZeWTpSrXMPSt7w127kGyFVOg63h91GNaDhij+iq9Gar8vMqZMJTPc+meoXZ7/+Ucjl
Jzs7yeum2bUBoOeFvFkvt0nDSZoHwEJ9chFqJrDzAoPKmp540hZfKglIwKOTWjyq2jtSpZFcrfKo
Ekolq3XMzYobGA8Yb7SKCS1WDTisjbEOQfQ8Mo1ZLOwc98nMf0itdLg+TssaeV5x3x9i3rOpQO0g
+PHA0os5WABfxKu0o7fvYY/P3brypqBArXHfD7FLqZJzXms3Ajy1g+GW5YcwbIHoY3KPN/kSQghV
9jN0+kpul+E2lxr14ONIKYaVwdUD28zbX290EwQ6YrH7HIo4UpHbsx5Vw8xpY/ACdvfRC5mGas2G
vXxZsXJVAikrXAF74Bi7A1Fu3QQ1bwjtekjxDs6fJ5aCpIOVcW8+1L5fbB4Y9+ZaJcOnAknx6dI/
UAhm2urd5o/3bA0dmWZel38AtR5bgpZJVmFdi+JtwMa6Us8zm4L/haXKZ0fGPfQppkWmwz5dw3JB
f0+XP8aFNoktV6n4x+vCs3JtfGICzGefKPh+XZfUIXUwC7qTj1K2sLZR1OCs43cgq7jpiTM7zcup
s2XTz3VKeXtkSZ96Q7x3W9HLz7wdTUgwqpi1uOWXR4dvc3aiyqFyfZVxe2Ghz/AJDyj8BWkBk5VH
K39TPe++cubtgYyaqsNzwR6ssgr4OT9AtA5j+xZ5iuBTj6jD4Dciar8M4qrUR9e4tSfoh5Pu3LxJ
p3dkEWhdNU0GDTbbNnd6Utzk8A6zNZG1DtAKsnLikhUvN49rlpis9PwaNc8K+XDUzWKLmYRW84TI
mMistk8WIrfC+N+YgCH3PJETQHdAKXJgSDtENC+qefRdTKhvV1nNM5O1ZspOIcX24PTPrYitQkby
O2+eFYEP8+EwuY0P2ihJmSw4N6K/XocHG4SefdgftY9VAmroWGZsTkVvtx0Xi5KXcZMLSQj0PExn
tBPaHXhi62gQPROIVTwJEghqP0ipgzGkmSfvzPzUpNRQVo5k142jgGzgtcBEHzhNjqK0WROGKLgF
iZXBUu6XhJZXLu5tdaXdbIapBTx5PtFNR/2JW+syiItXFqugomt2jIaHnYnIR1iZz89rUf0OVs4F
qlN+xsb+3KFVVJmQX+PWcG2uSDES1pKCfcJpsjAlfTUzhlF749v8Qhc77jivPuyLYZ0fGWCLf+rh
PP+uy2m2agAav7DyM5AgG8vfEvKeppAPfLO8moifCV5uGNa550d1fQiW0PFmlWCP/7MvY1h/ARJl
msVIUaH+Z9NbDdrPiiVFxKz5h5VAyQEsRC8KCLKrvlq+DR6YoNqemq+jkqdTW6uRfFoPXQecqJyc
itUo85zHA6wgJOk5MEMAB4jEo6hObAapggZLG5j7gbgZ2l6p8HjpsRTTK6v7gs7lXRT63pQOO30W
r77seUDJ50iDsX7wUcGRcleO5+Q3Up1rcIhtHwPsVywiWN7U8lLzyL+UPeiUOaHNur4/WWj3VW+T
dS7Y2CdPAoBbWQctm6gTKp5kE+CdmzxGUsRTbG/SqEe96Pw8ijkDdbkZ8hWF9ZS7CZ7y35MKZ2vB
7bL3ZJ4rZTrhfAJirYjZxANz0W+NcKaYt0k7Y6tEvIb6evNLZkE2LqvzSmgNQifp63O6R5dv97oO
oceUkK5QrcwZ/u7qlDKtnJjqFHHRlwcHnkvi2dY+OBEvgDDUI3GyAHefIKNpToCYo9JTPDf8XiIo
jVNb5r4N8ITfAb+YGZd56Zefzt4502X238UIU79DGqVXkboWZVSgst2qX9inqZULniPtfcZxLyCj
/0UPTLWISnFJAmLikGk7zSnDpWuIWbX5u68Twofl8+QtvGuRGBEDiaZdMh4aWKPAvKjg3Uf3VBoY
NcYm7fw4wol+aQwvEvW+fTYPpAk4FaHHBFYJcKBrQ+C5VACNy159mt8bWpy0Z3o6SNb5TDMoEo1B
P3ep7XMoy/FCelzATj0Z7pmGH3VDBwyXruwo7xMVGTBrCGlkHHQeaKk9GerZb2v/naQTrr0q2Twz
MXigXs75FfryRSOCTCwesXWs0s9BlfxTTqXxAUaPte6ruW+ugoKexqFGd0e0cZ4ssZQczeYISLdB
HVg2BSxyUuhzvF3I7OOkrc5eOTZk55P1pVTt+wLQKTcpL9AX6vc8DmemzTnRn0qfK1ITnFr6vDfR
lou0F2DcJCYcQIFZmtI3kQdFEYNKDAYUppSm4Q3LiW+KdGPsJEqBhxGkwL+U3l1X2Vv58sm10ab7
ZQj8Dt8EMl+kLZMmWIqiJf66YewWgiWqYhayGwRHMdiaZ+wnUh20zuI78slJyJV0M7L6FeQkS5o4
Uy7aUxsDW6ozlqjeHLYb+jObe4a9w3TeY5Vdk180t8Xmvygc/VCEA/hjOo/C5/ZdD940CoG0gn+f
aA2/+0gmuPGmf3U4Ky6ZWCd5a8vJXiJ8fmGZU8e4kjAE9+cR6cNgBGoK0df6iFEtOINExkQcJuzT
1KU+rD1n5sFVrPfLVnnykoVU5pJT5L/7fAIQkc8/Tff7/xvF3Lzkq+UZ6gKt0b3AUjN0hSpMKH1o
+RDLTM/ETjoKFF8W4xQ3A22LparF41/7Y+jKcliBaB5xw8X6gRzOoWWe9sGDDf//iM5kmJPr8Qa1
44dMY6J1JmwaWlRMP92mbhyR52GwmYJsdS0uJgHBN1qSm2xYlMIRHmuP7yBScLKzC3IWh4XofXpJ
kceZynSYjf2kFs7k3O+iLwgKvD1/krWy+Gn7FGvzNSLYsqNgs7LOaygss8BeaXRnHttrn8UyjlUe
3gmypNkq3MXbg6RlOprVSRMJfJYjt509as7k5KeeMSYl5HqWjA+JMCPLERDFmStZJjcZDIu+38Pq
bbvZP0gujkWyJzU9mCNSM3bziLwBP44gzEwJ3Tnv8E2Bk+zIgHy0O4rM/6fx0+49dnd8pIWnQeYB
yaLX70siFpPHDWxXx+8vN6I25xxnIYJWqBKKUs+nj2RQdrjMloQohYrn0FF2BKHeWtP4eVPJ1RO5
GhNtPAid4SViY/ThAN2So+Qg4GXD893cIxWfF0x3N9tzn31Aa/KlbQ2IFWXuKD70YrDn0+hbe/bA
k8MKyBliZ42iFegUxf8/wCeaBf13I4j01+nLwfRgXnmoCy5PIVFSjlpGuZ3F28vcBGP7q2+b+r/f
IHQ/5I0uUYVs4QQFVz/RQmYRa2mk0NMJl4Avb8GwKDC+93W/j4wzKQcahawevq7fwUlUD2xMFhd1
i4lMx1xUMzQdZBHwpQGna2RBpX6bIaoCDFNBvlbuHCjZpKDyK83NYiJQU3fXhU04EQU7h/52EYlR
jF+c1cn2F6OAnn16jjErdCcnlq7IJEfjD60X5vWSsNVr425tth5tyxEEPdFHZYiSZNxPpov5V9Bc
B/XsnP8tYYCylef3UJX6Wwiz5X8NCnabyKT3FY0XEc6fmcjA87zAzEniy0GLhu9p0YA4Nqdxr+E8
9C0o8GBvDDvIjp9YRb6wCKraI01pj2ub4PsVazycgdOHC8OMBobxGfWDv3LRimlTEjX8eY0NLYmK
SSLFSzqLKA7jeoe/vHwnY5bbckmtKYf31UdWrxXxdbwp78g8+Ky0T3PVoTyb+GKFfwycqt1PPrqO
YCM2xkKkKrAyNlboJyxfkT08UghVn8sTHuRBoWMrNN0dtb8lCdj66CAT7xXeIPnnkOwLBxIVxkUK
xXvS8a8hHUJt6GALCLzGQ2InC46nUbjssKEOayyk1OsJ/boEfyzeWU44Bd8xM3hLYEz+10RqzQQe
87fxA4UfteHNVaRlcxuViPI0JLld/yhYeVydyjHX4/Id98uohE8X+Bzzp5yu5O+WINwqjEe582JZ
0DjnHYkH3rhVesIxNOgvhZcE/PrlG4Mh5jV7bCQHHmjLBLSNbgglFJtbz4b4nXYnQ6ygnIzCZufS
tj9BI3mg9BLzuhJxqQuDlWIrEIbxq1TKr/sNsb1YfQPsOPD9YACq6jsWgWfgv9U3oTHEvndkxvVc
X1sQy78D2+Lxu2mn2lHkdzJ/gljPCrSPRpjfhQPf3QoYkE4GPKGQizfmICQIeqtuCwQHTiF+JyuR
EISj2toUHslbz09Z8GBxfvaHV1/1UtfBceILmj2UyPP05evQ5VS2MQBlfxV1OvRpCLP379Dws/6L
YobMVRTSw9VLtBDFx9YC4uEGw4EUfq5lXvJC+sHcX8l5wvdtr/DR12l3RlNXxgH5MGnrJbmsKw9l
IkFGRhDFC9Hb8o8td1wopB5X304nZOCuRRIV/ruH39HT/PzU4011xxJlkXww/jnXhXfTeMMK83xR
96HUX7ltl8kiFoFzf56b+npgfnSwSQgcWcQY0Kh81XaAmPo5q6Nc3sVQuBeM17ENMcsUnN9jmELk
TnXLyFd9lS9IhulwqSRv3nHYnULzq0tv4gJcKis07JgF7bRA/uarYsBSqzVGx19tYTFi/ehnAbzQ
mCdsc3MnDVsV68bLCol6QomFTFBRklC6pSXYhSkDpA7rF1csL7xpYWZ5HJKYtP6saQOB0WuoyKYx
g/K4cEQ71JAU30ULCZ0mi71tHwphx3oZE2upeLNCFn1yutSj8uM8VpHksCz7Uk9/7JdAgsjZR47f
I1LltMU7wbmbnxsuai+w7WvoxWkv7g9il5LThphdnKw9Y2F8F0t5Z8bI0hs8eGUmqrJdnQzoA4Vl
VXT4aj8Si0r5hn68q/H0MTKZDwFGaSJhk0qtaRCZlO6NOSEQppbIa0nmzzDuYun2FORkzFoZMxya
nzQZ8ZQqv33gXvZa849NonrJvtBmcD/SqqLR98P6Ia4jnozOJsAAUNZb9aROVxBvT9VQDHxquCm+
6qeNVnsdLu/uXOYjehoGjcxk/EGJaOlALMmC3jKXDdN/8y7rg23tQwHGEY9f38HVkqOLhyjieVEB
EPkhaC0UYKAU3I7mngN2P4/azitdrukRyg82LuoLUztp2G6YirM/j2d8zeGgVtFE99/fBo+Yj47C
JUwvDFLIq4JBLdYx9sA85zwQUv4oFA1+LE0WkYFXU0SRGFG+PkiRF05NHNrDo8inQVKtufKABWjR
dSpfY8qw7AOyQ7jCTCDUNG+aTsLRKqttEoaVKRVe0mKESjykzCuRwAZ+0X+7yYlLitBksRvwyLCv
l6ahgJFso6H0MMisrfAOnffJTnKImU2f1yQZOHda7vppp51z2ivjMD7ZtpUSkkSSiUgrYCJjjhNi
Lc7rvwYkdGYN+bAfOSTee3H4nObyszXjnAEkl+tSdin+p9pFTB0/snpiZCPI/zrCA9CbxBH4qJj4
bmGmxc+EwDJt1t2SrjczRg9/lmcd3nrP+23rW+k49Ka+y8lt57of7Wjpi0V7TShvNCLi5jaObdQj
HZdRzpYZPOHyUMTNW03wY4Yun47BH0rDqW3LOU5Sr3ZUljIUltKqNctlAve301EobbkOr7P9Jthd
l0ovEyTki52SW6CKgjfgwmetge4VwjPcrL98V5GHBVmnljAXXcWFEjPIHcmXFYFPGDFrFx3IWtk6
PYZfss7ESOWG78dnJVsSm48rfYCm/wk+ptxu4uOFpnMMBv8wzD0dB7zn9Byo7jmiRhhR6oq0Q5KZ
jUdSD7zN4ZjFfHk8OiD4SyE10rCq7FcQvpXypLGHc9SlOpYNBYql7oTwVvA2uk3euS7dpMZKUOK4
KXqW6nfv7BGmmtQbqzgVYI6RgZdr+ghog3X1pi/P9fI0stE9BGeTLSpOluiXKGNUFBrhxNX2GGDA
ju2gfPLEHxaaWmyQvwojEeXYck+r7K1JrjpMaiwe7GXD3UJTp7RTo5LTmlKlzAh0dYGKRZGV88Cu
ZTzphq8LQ7lA0J5A/mxAxIC7Z7QPaJxEnPFEnxdfXBPKoa6X7L+WtcBHe49UsEGh6wZdtzYNwkuM
hi2KS9iIgFy9YX2DCKEM0rXWcHQXW40QA5eoXzZljDxq5NBvCSef1yYThWZqE2mFF/kWPARECob/
pZPJxt5oGCQCtWLweZP9ClG6V2ldLC2FBJl+9KqCtOFVUfDGMSt6K5hOR5JrsmhLZbdEC4hP7eHy
Y+lFk7jplXmE13lsuttnhz3raCNgz51xIywDNBZPJ+R4dxWNtXK19jVN6QhUGAdlghRhMHUPq+Xn
UVUizCNy7P/2n8sSQEbPXHouxapu4u0Yp+SZdFpXvS2LVjk9mU/04PLsSrKIX//oHzsPpGA3KTfx
Uzfmfnk7TByl+KaB7DqwsK25ba4Mq+9TSA7IwdARcEyIT02M13jXkKyvN0fU7YEgx7WDlRy2HkEe
4YrCM67D2/hSj+A40Jy7ly4j94ApMeyYtknSg93dy8TGSSnebGjO4IRATZYgiXj4cGH9Q1MA9yku
3xILiLTmRXURKlTVSUXfWM8oSGhmo1xMgHGS9H3v7+XUvCJQKBnLgSUo/EusqFFZ0OTkxcBTbcXm
vi0T0HwiwlPSlWfps9nOcKcHWgS0PG0zsOR12ePKjsV1lE59fJFs6tl0q0iBEpg6pnt2TsE5LjpF
r0RAIuuHzBOvQOCuCNkiFu7HX2pfssL0QODCXkpIwZkeC05gqSCTiDgjwvQbmKzGC32xL4DwjEql
l6uO7YG5dlaDooPFeIoLpddpQQIcvdnvHKgbxW9Ia3++M85z9FvdLUSdNHmoeU6qIRUvmzo3vx+r
m9LbofM1aslakyDrvD1XaglVJfa4f6f+McXKuROMadwlOvEXjJoe4NRFns17/07vbrF0+jhrJBHD
kVOmRgCBTEfV8FJfc2fAMo2RKxr4XcdRV8Byq3EqgGuRGa1MdIuAWasTcMosiVtvvgGD/tPTFbHM
YvmMNKSwUYuuJ9VLHL5CLRtv7n2Clo+p+LDsK1sc7nBeoG4a/+P5GNxgjqLYUspV3UUOIAvfU+Ph
sHaMyEkNcUFtht10SwIdpnoYcA3HQbP34Fh59FtnG6/ZPThrSVPFJgPSlBvFgV2pCX8ijS0HKwsD
d3Fujz1v6lEtiphkk2Fi2PSRB1Xu6MJ1VExtqXtq7vuyQPXqc9FaMHOUHF8hui37MwlVKGqXDmri
txT49PiQ25T7wyxP11pRRnqdgCJknQ1asIudWkjrXgeX6U3+rP8MIjJMABolbaMLc15U5QEvLDYt
N0DQ5a+f1tDGiGoR7CRuMgPHWXpS/qHxhbaCCbFI9M0Xr3nwAgVP06EPZ6CyjJsrsNxa21UCch3E
haE3+3JecFZoOH7fmskRFNkAqkis8M24yhm8lLHWjLeF/uXgARAYZFwbqV/0I0Q3Db8IoXsK5v/S
JpxDxt7G1ta+3MGDOKwjynWvbhXuDBsWJOmYsI55vHLDZBvwE+0wNc77V7FMN4nKtjt2fyiAC0Zq
8iPpPe8L+P6OYv8z7nTMtvUdwZnz4OdN2cygh+K0e81iC7sR0KZNCgbvjjuun/PDq6j0Zg1etCC8
UEt80EaA38DAvQvL/hCOfSDJs8mDfeN3A8PeZirCDuCo+cr6x0K3h7z4cq9JFkBiDf3S8hyhO76g
0fjDQ1qDcdy2sdq/l6mrdCedMzRPW2DxksNDE6v1cQo0FHgx436vDAyC5AdSAuzSi9h74Hchi2CR
I4YJk5x1TTT21ZxHdKooOJGwuX905CLG+13hsJbe+EWg9eOiZ07iZqLVTl5Zc/L8X9zW2cmdZgdA
JyDJkjw6cCC9FDPgPwh4d8cZygMZg7zQq7WyM2lU3U4Kxe8dQRIXt8k1sZU8UCLi9ZmklA9JAhWO
E4YHkJKYEyzTZrmYysA2RHTuDQZX2fYFUZJAKwrRXedyO6cwrhNZKftWLk6ZZjK4PZWu9fZCOCSM
MzXQddhr6JXd1EcODy7/gIFZPjr09y1qzMmudY4+JpIpm53HoX0Vldas/1hPwmMyPX7v6IlmGTFO
Jwd3pJ92qjzrnFh3UGYDcdJlwjNHlFeZ+/rvJ2sqzQvtmCjqRZJcLFLbZ46YB/aSjRihDpTdOxhs
6/yput+4crP7fEMWgzP41tr2IQ0T6TqORVCVXVlNOIOTiu7d85P5HZTzgJtiC1VM0fPNPrCJwfY5
FE7mELq1Cevkx/e89ftzDCal0Ds9vpnkByulYCAtdrWPo5AKvhutjnLuhxLD7vW3I7yCmZMtjNs0
2/kGQjMRGUXhoV3qks0UtMvCtE8PyVMQRoSnWQ+p7mRwlDhL6MRAvyx3s295aSm5xnI+S/ipI6oV
rzK4IsJMLQVjYSP3HY6bGmTseQVi5L2R8ddvJDQl65c+lmV50niE0b/WGcmetcl0DEy631CKHWmh
vQfE6Re38LbSU7qMb1Strl1Eb9vjdVpxOzksnbF9nsFQz7Ne19ZYVJmVh+ZsNdKMsXhwEm5VvkoW
gP1MxC9VEQz9mCeKiV8XzDYwUTQZMJ7gsj+mBvBQsR5Onp6zqX3+Y+gOFZGilCk8mMx5QVda9s9+
iDxGO2+onqAjgewVTWYrWSkQrY+iteWWzGCHoWc8bns7MkrHzXNH8XV1bE068UgJymGW7Z0VkzEv
oQP8ZoN6iDUM2LL+OpBC/C7QjMCcOXCOeVEFT0wPi+3A0KrTBeAKLx1f0KjWRmemadgGKgPE6H3y
mnXZjmiP7a0GrhBu/b8CqjwNRQFeyNZGPPzJWnUrPOGNjIuH3V9FjgHCRKRG3hjUoZFSi4cyX9lM
2LirsDS0NCvp8+GnJ1M48eggtG0vt3kFuPA55L3XGVXFOgu4rmEoFw5COSsHkmyEe0swlygX+jI5
R+Oc8P/uC+FsqIg7TnjkC24W7L4dEysxxx1A2e6Raxgd95pqVDkU//pBGprEZldy9oKcLLjfB6Ml
3BUMi4paD7jfnGnnQxFV/HozNdiU5w7/CbNjNab1ofs5N1LXC8m50GfNZRCiQ8dA0Xl12dOUxhby
6Q873zRbI2pST3ZgQj6ClK/0STVkKgO/0qpLrp0Xm/A5s7eJYUjCuDpnaDkatl9FproWdORJMquY
1Bd/yqjrSMxXlHJRDSEWC/uwKvp4unqhlBkh9biTqwLqawPJGlIIQ4KhMLse4g+yNrluB6VGpPsW
bpqxKK+Pjt+gWSpbjcDkLrHW4F1gmyPkWmmXtre6uYAoO1Swr8o6pqNZVzus5e+4UnGpxq/DQMLa
BdRdawdlpXfiQMKXEh7PZnXSsG26p/jl79qTErs9OyrTvdeyPvwp1jV91jI2h2qD3WzgBOdEkrmQ
8thovvDOecbQDl5cLhe2jCzp/SAoY7pTdUlWTio9+Zy8b/52BV/k2ldLIF/eBhC+U2bkMGbUkNCl
LzkWP6IsAMwi9sntHexNMteIss2nrkF1ZkhNRTPzr3RL3g6Okt8lSGwvO4BbVrufQoCgBH2H+bBQ
JO1BXbv924iLYmKxJPEpLDUgVRt2XkqcTIWXTjBADT+abdWnT/OD8BAGt+FiPtde0VthfMBg0zCT
OBlGN/mCVkTBv+iS/IlB/IfdNObrarbOuUqowaA++YtelBOJISHUiA4GGihVSQaog5Iin/CaRr2S
7mFcNEDmEbdrCBy/TkfOLqsleNd7RZoAE5jNShygC/CGkzwae9Xy4mQVyF6IvNTgEwlYRS0b2vAr
EqN3JIrkNf5YTTzSHOalb48h4VAtTLz/rxHDx6jnvtIOExUmMGWiGkMhl1E3PhjUyPxFKEnNx+eN
c+m1v5HNDA/mLYDGTCHOmpLrZm1RhoYyP8KjnkxRh6sodfE9QseLMkfnmMLmKvWlKup0tEYlubfX
vvPSREUwe6WH/bnFF8/z7UMdN3HPZVc8YvQraZXI1Q0O1aoLQMmlysCpie4+ttie0VvFvXJoeY3h
YJSWiHzOOq83RtEGD8BmDIs7oJPMOGMIyQdLmwcQ2YQKYzV3pl0MY0WXwf7Jti7tsOcv3aktb+5d
jigjzXDakHpAU39b+jApvve2ivkZVfNzhlMiUm/MgkmMxgTYznjp7eypmYCRIIvOmmYjeXscQtGv
zjEEPVTx7TVuuoells0E/8XTWTmycbYl3hwf3Te3V7zBlXpsMNLNSq60n/3BWnOvCj60dZzzQjHs
DaSuwkSoIqgJh/GJGyB2gCIAtqMmr5F0VSeahx3ZkVDRRkcI7+JnE41FOEkYauLYIOLUDaDqoF1g
459vnG7UQoZIgace5u0636/A73F/azV5gdMG2ezIOVpNNTbufkUp1RLTwUYlfm7xP56S40l4ygNh
+9Wkl726NdU/eiJwpIJp/gQz7lSqcXYb5dXpu4q+5PX37i09MmkjFME92IZiorzkjSBuKbGOz1Wz
SpBfhHY3Nu1DrwB6GDEWIpXQIOdGbt37tqlGKL40wYUzH7HcuCSB/8tskvd9IGys/3j1wD1hKOej
HEYUi3Lxyk1PlGYVIdxNSwdDTVmyOfBvxGNo91ErsI4oom1TO4To7lVK2TwpEzHZiQNqmF64fb/x
th9lEwMjwc8O3z7v43O2/yxJctwX8URyywp/Ze9ASCuGD1+PpwX/moVUp4zxb3lIah8H87UPu8lG
8ZujXhMNNQnxrx7AER/48ACOzxEtVC3VoXSKoLTzgbQqFh4epEC8OqQXpvDap2uOGInywNFLErip
B0fXwUqVRMDZJ+0D2L+nCqNpfwwQIIXUbsn49rKIKJ5EmT+/OrdHRglC3Aer3XKSFt2zwC9rxKXY
fvJdGy8dRNhujDv+rcMn9Vb4hJUtrKHctBtWi3n71c/tpG0FTGrjnVh6c5YqMdDVSuyiILzQCahA
ieFiYnz707wBE1hWUnA1p3lrbOwBtv6uq3+ZfOkSrLf3LHdqlTnjVHm5ycX/wVHJP35I/AOYKMOC
Esu3Wg8GBpVLSo7dSLLxehKfm3smIaerxqZFT1RjOjYlFWetP/dl9vXQcCFnoxybsYUorZO9hzxs
gRZVyd4hwmRze+vxUKxqcaHIhqPNumCV3HqTIfsCnh3vgLopQCAhy5Kh59hzPAiRh8QBPD1DtRjR
8eWfxnupPSjzDBUp2T6FmvYtte9Zd7sSjcPwBjX7cBy4RDu52EkfxHLAyqXozJjpdoN0jrv4hpfj
aS10vieFl3YP/22Dl9veDqpmtZZQjkxEEYNIGyBPrAoHOOS3Vbrg2keezX0vv9Q91MxtJbuFr98V
5hyUaCvhUBY1x785qQJJqDTxFFA0nPKZ7r9hlKLgub73kCAJNmvrqSoyB1UrfQNRK/x1IRndzhRd
wHJ+joAbo5b381Kqb9haCbBDH1+738/qsY7PR2dW1wqcK+UmxPrA3v7SSVUQaOsWHRZYM7kgsJQ4
D+EWHlVLS9/19M2cSrx06HzBXweO7Nln1aLfNTVrIXfAt86kQE7tzJ5GU4hF9vnqyN5J+Hcj53Qa
zaOvKxpPkiCLBElKF+q/fTi6AUjTk1k3pADrxP+as8N9LxVB80dpAXVyRUhejju2lRggALUuQT4K
GVbzgLG1LLnRxYbfDCfUNGYUyZ57Lg7831NWISylxzcJKMz6llQuxd4genIimQGA3Ke0A+g/ZtGS
Obr4eqwekmto8PDkcjO+Dxvc+QtlRMc0SWuF0wjFRQQdUe6a8pRch92Dx5rogUoO9yO9lFTAIOX2
paGx4wtHGNERS07gMBhBJB7bwTNiGxK/TzVPCCWYOJvvarp+bwcB/c/D1xqApldJXzVZu/CmdwMV
l45DmynwBa84rKMhloKO5uZyj2TWeYyOKz46LIRCAvauELHVNuBc8kuw1G25qN1YFYAl96ra/wF3
AbkzJM/DuRqYHBlI0gd7MI17/CkssRxdqUTbDXYYpFCE93041Z0ImvQ9ijOezhj/kg0Z64lrE4/D
RTLshkfljOShMPbXM7Oh72EYMGGgv57YDJgFz+nWXAwd+qCWOrdHtdsMMwd7DL3I9SgkRshhv/c6
tWs0FrWF0pw8ylVPuuLSi9ctQZUgTjYBeMePHFFgv7/2gps/wdHuwhRjPe5xnzIbpl7Mnu6e/0rr
4kqGDbd9A/RhNS6tTTEHU/Nmcpwkgyw6Ee9UmuQ9i8wAQ+XnleDV70KrKLw0lZfTT3qyNYaq3emL
wxyz82Xsx1FVNwZHJAeMD2BHoBPLKWMQzjOCPz1TVhEd0OyyFg2Hcr69eZfBmpyc68iEWMrpe14F
SOADWGkrrwLm/Ar4IC5cA6fzCpUe6j5E4efh4FpYizrENSnPhIkRIPJvFWH11zzyIL0CpfzC0LXg
4/RsJH/EfgU7IoGLw7TvA2RNi/oXT7iFdWNNV0eXyXA7YM0OVL1w0MuMS3VPUaM+VbamWCVWAY0D
wJFMgg2FX2Uxatj687GGVELj6eoNTe6ssjXUS6dKOhQ1aG5xCJ9fTW4lkAI4UssuFCJR9qw4/z8o
tFwYEOKvgc1Bfp6eRj5xJfMIO2vTvGfewhVogRSM09VQDhWa3E7w9bCuMEsAAnzDdn3HPP2ibdrY
rE0+ZOiAQzy3Lo5dRXwIfFdkrCH3QKZwATxwCMQNU5tbnQG7qk4Z5KiInRhAywnf1v3c6js+zRGD
v+0vppRA2MsEz4nZt+4M8q0Po6ogXwDM3gZkwbbJNTNcLetosSvBU++u38/hKm7ZNOGQtEuFKDmQ
oZ+YE10CzMeSN2VyanEGLq7oWBCkm9Veumsdj2LGMSsJS5ysOQ3tOa3mi48zGsAl7fY1z7GBOuhc
PB7JUOhfxFt7hGtiRxriWBTz7NHf7IC2gwVJnz47+PUTpbZoWOx+FDProwXLbv1M97ZdNiIGy+UQ
vr64G2HOt48I59hTkafZKCdWrCneiQDWA4IIRIX817jONnj3y3kEnyDqIzpPGPpAHPAOKJpwIsR7
QHTz052jGlpmFZg5///GBRCbt1aScVTkvCZl+EpSrgttxGqAOXx5cW88LqIWFD8rywNRmDqIjpon
8L6zWi9QgQETVUgMEn+u+Uxk3y1Us9hrNAivGwj7VQTaMA+G4mSngwSyDqCnphaFDPQmj33xRNLK
8eDxHRhrxTWnOAsuPP5EuM+rjshkt+JCAjKLA8ZR7GjG1LEwkFmlwZfMxwPAbkwy7GChbFZp+mqx
CP+AOn9mEYHtrJRZsicVBN0y1WPjXPhehiSkjUL7plCC2+OruFfpjZKqq4keFUQ9lHQl33aPdRPq
jHTvnaJ5MLHh6/0P2s+1Rrlt44ZKZNRPKk6C71aaxKSSKENnBG9xVk6uOfnd/l7WD4ZgGSIa5E0e
Zf1nvLK++bZWCyQj/x/fatlIjjKFFJpovP4bBWj4BQfwq4Y8QSY+zUoQF1OqHcGfMkHEBYep5Ks/
/VnwF6vSYg2MPqOg7kXg8ofYpqAB/PSYuy3dCJdXYqaU7GpcwdUxTjXLqHKTUWtpzQ+fofHmyroq
O/lTlzi7nhzHzmbaqqll923zADZw+6kE7VEIdxmM1RijZI6HGl/pIADhDY+xsatrqaVJnkPaoHlS
frm41bEA9hgpU/pcOieri6NGhMWhZe+4fPbZzYyBO0t8OQc0hcw6e9j5opg1zNYbgWhRNEU5yy+H
44Qyxtsrv6QKxz1TJ61XR1RCy0l4I9pWCnshONqnCA9pzwKj9Ow2k3tIg9v1dNmDIC++qsDRCvvi
j6WtMisOpNvrfDThTymiy5B3V82gb4t5VbJ9UzqoM0fYUQCYzr47ehNKiQc3ui6nlvJg1GpOdYy4
0dwI1npBO4kbrLp10gB4QLo3hnPChjWfO6b7Bwv2De6iDED3juVNc/Khi0cqnALEGvt9WGB0irBp
ghZHEsMX5Oe+d2C4NMVXunFA5Qfd7IT54uU5rhW7KUlTjnvZ6W9Ub0D/py6s6s268uGx9dzVWc2c
eBdYX5HJyzzauaIZOgOtYuxM266ILdX8J5rKWa5Asj85yyiR9IxqR95CjdQrmcethIDmu1e9RlGd
PSYr2Ae7/7RJ8um4VwUelBpTmgek8tkMxmxfYiECVABaebpJAlkYkyvpKII/W9PXNI16LCMyFfbV
iiLJZZdzc7qw3U81bNOk+l3wkDWpg0WTCickekhHAR2+SPU5bgIg2vCo4lUKrDXEwAVO5ORDmGHp
DufeMUzGJZjibPAw6yuysUVZXOVznr2ThHuZCQOr5aTAmbjeyuSbevMhazpWfe7VxS2UMEQ886Sd
5ypZkrUpPYx8ncPxZI/K+hDB0EyzgDTu85W5E8j5CSK90655Lt3E23EFiRSDMIUL8cXFDwjP/snV
rtBy5Qltsuhv+94kPHptK9TlS7zDjQudOa0p5YngDmoIQwz+j+l3V6WWNrmyiURIfj/lOAUjqChZ
Z3vkggDccvP4DK71XQKaZiFABlz3IY3izxU+aGYbVZ0lVgGSqBP78RCQlvy3CUrPDxI6lSs0z13X
bVT91v+4ospINSHcxVRS88dLaj2iq9G1sj1obzfdQ458s43Ffp5ONyrz0ZxyBq08He6OHjbLflzz
3au2kkxilKETob5XYY+d9tSOksD+zzVgANyTo2PqG+peBUfgZvovgXgQYvaV19thUUjrNs5DlnIS
ZqzR4UWoplXTtXVMYIBF+l4P8HQKpv1Th+8ZQ3IUamUoV6COFW54HSOuKij40JrfMLYznOr52oRI
3jdC3mRjKsPJFJlwSky4wQ+WVRMk4zoT2J+2HU6H00Jp5Ny349llCz0/Z/aBBpJEhYedVSD79TsS
s8ROCJE/laKnkEcjil7RK+fLgqHBmJozM3ZJzkI5Wp9Y51G5kgbgetDYjbYfPyhziCJeU/v3pn6Z
t09Bw9PPO4rqd89dzUehgQA9UUTYHOX0hpXP0DNb2ZapzMMo9MdabAk14SC4skuxF2h+Tey+qsJZ
sAYlgVTPs4mp5Tjp/oTsM1jUx8oK2DKdnhsfdxl8bO2L+n3g1fx8IpMUbKAcGWl0KW9ksCB7+RQH
kI0XYuyriNo9s1rekJhEJIjwZOLja0ia21I3wLCdx+ak/VhlmrvynNVBBzyfMzhoKEpR9bPXU4a3
DvGSD/WPZ0pkDK60LNeM1Amp9tCEGvi//P3YQyCDxwPMFNxvu83PdVp3gf7QosiUfn6hvnReqbSH
wbJmPrGZy4eyTWgBvCNvRcytdL59ZJkMF6FvH+ZPBukHAQizJv3H9H4FZb0HxQFMBfjc76eB9cov
IBJd/aAdgn+CqoYVhqsZm+D8o0c50xFuj36pJ6fmc00vZcJBXaDh/RSvGCOdScIARLSLHd1j2X0t
GJuxqKqiRmCmSKbdVuN09obzm+0tPfO3aQ6pDmBKVu9PYl6fIuY7a1h3TUAlgFanCVPClQ5U/23d
YhRK8ycOjA+CjD/7xCIjBLGFL5XbcFLJj7Pahe2e0zU+6f4KDxKqZ5b3g531DcqAwzYBO7vwdWYT
LNy2WVPlF+O8WAEP8TFEOPC1SyN37WJX5UWu3dUy/gABsdm6k046APgXrPMmsPsL+HaNrvmK4Gii
AwQWJg3y6Bf1UkMN2/3iiinnFshx3Y7NdrMxSaP/gLhXCAdtN8hgar7MuXHhpKh8necwHXKMb/L6
gPxHuj4SdMM52w/8XHy6BvjuaORiBBEd0mN8/JhReeeCCQ29JaQ2mQVW8wFYAF/jWLko1vsFn0RG
4CBP/yaBymMx+gpcsNSNpgpmaPG3Q8NbFBmpUI1MdCmR+yvGRKiWQsIPq/+EdzcWVEYLlY1yNvvs
kSuYG1TNFpfL11pzJF2jyrD4Fg8lFy2Xc/Fy0ts3rBuKVcDm2HB2KjhpSNNihnRMv1a2/7rwvdt4
vWk6m1nM2/zWuPVaOnxGYzw5fjIU6Qw0TAp8VbsICpuWd9ri91PBlH2wsbOG2srw92V5XAgc1ZJn
5T5wdQsg4OHFZvylXd0dBoxca4C7Ojwhba9l3o0rhqrfVGh1Y1qUpcDvnK/Vj9wtZk7cEIh7MK+q
/Y/BylMm9dozefh7L5gH+rx/BlVYJTdXWfb7791y4oVulQ9/X5p1dySl34JLbnR0Ea4opgyvPbQ9
CczrbjgyiWqOybdJWLteQFqbQzJ6hSRNxXNQYEuRPvcaqsy9FY/paQar8ShlnjQsUxNrtkk7tTld
XiwR1XQbfb3qlldRYCziK9yW0kdvOJaxo8EeIBY+VKGkI5tGRA+PPwdnwrjCSrATWos7sjqmw8CT
WOSimi55uFTbM8U33ZRPs1+Mvtz6VUjWdHSgyU08wzufVR464Fkov7O17/TMgcJO0GYas2A4K5VW
+ewKP+Qz/RjS6fQW80S6zZi7QscL06GA2DU8mk835/3dEroRHh1zWrdGQL5xJAD2WHVid+eextqk
/ufPQRSWv590lsSHB6hZUm2zBUlF85+SbTjYs6QI8a15vzApdTYT1cI8+VnX075mL68WawM9xjle
SCjvmqw/3HAFMpcFkzdLYkebQcIR57De9/BS4DjSOgBQdUQjwIodoTSO3UQl0FIDkCI/7vepGePB
1dkeJ9MhTYr7Kx5um1Xw8Z7DehJtSvBJydnVNDg9hMiGRJ0nMqau9xKNaQrOoZ/l5KXkRpnH5eeT
QihsK4WI5t4LOQA2DZ08eOnFy4N0lGECssz3Dv6Tu81k5V3pg+m/flzOna+0LIGglvHiUm3okfok
oBIXOq50Ktpil9Rtn24sMDVQmk8UYDKb8WVfPFEBWcX6iOefKow9/WOYMHX26NWKe2WoaIkE1ELs
DvBq9Yd5z+cII2D610XYMzCdxSaACI/f4noDYaPM1ShEs1lurd9YEbp8KUWhRuEfNYrCy6o5HaHU
qwVHkCHIh2kaCXjY1uSl794/O4UfSu7KdXltpgWeWzdyKtp3vFWkht9iRtWO9jslquNQ1bhfwZeS
pAwUJ6Cuiy6tyJ2pxdOkSrlrtK5lP69LKKCFSyY9bto9ZVHGMvl1GiZNvRfFn2QwgAET0MRCCVbb
IwfrCgBinURLUM4IyrN/2PNt3khpVlltC8zTYjhr6EmkbUqVnR3fX093tt7bOX2qPADI3nfb41lg
byEBunUKLsHVjyaUyOPl1+dyUSRcE7B+hnVCWxrFXWQZ7W38iFA8KDjNDbOOShxF+64600aXeS5+
eopsojpy9aTZ+616uCaHft7LsLVHQLHRmWrJPuZU8xxBGY3qRYDlop6/BpXAzAqteNQrJ1RqaKgn
BYlQ05dYNtLzap6dQ/Y1cjSaf01q5L0hi+FeYBAeXgouovXtJYnUB92aHj7kPyz8NvnuNSXruPzW
T4yNHpt/1mMrD2RlcxaSvaHNSivfLvB7/eNeOxvxptI3+Wf4BYVvuo/4OAK+oT1QMikGR9BTZoFt
rPEhIosY3FAimplwahQiv0XJXeIKwinRCSfQjFaxexwdSUlfATCpguRmnOXMj+sNRHEdkkH5aqn4
zKcTSeaIAGJ3wnnTxiqHB9gWIGIElwqDGF8Se3Uy/PNcK/rDfhZAuYmjXRGHUagbzAs+q7gudO3O
iFBQH5ZgqYf+hZg8lPdzt/ISOyxcMSbX7RChbtlhA/Y5y8BqBGyEt6l3kdbx+65R0zdzaCynuhjH
ZD8sdWMeFmJdUbKpq70UnIglKRRxkN+n7QhGP5UXHYJeRz0hu2pEDAoeJEnyymiP+LCl5FMUL5vO
e1vp0QFaDhQaUhE3xtKVoaGUiaMi5siiodd06rNT6bbI7XzDrUqWuy8z0yjoCh0C2jxQ1XsApFRB
zFoL/250iw3u7vvz6dsgVgzS3Rs27v74TaDElx53AimKNFjgVHKTjBHpNJPK3y/2ZcVJvM5m2JIj
PMs+nVDe3w==
`protect end_protected
