-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
pPPgmg2bP10s9lVSKOkp9XhuiYaK0ygiNHctWT/pLp4Tsu5Re68ekMZWEsol2BkqoSUOG6TNbMl0
bboNO/IjrJFk1hLe2xpQpoihhNxzIWQBx1IRTHY3D1xQpUQQ1GFLac45Oyba/gqT0m/T4+NIaam5
WgVuTod+7T7nTa5i22ai0p+8QSLZ2NyMoc8pE9SQ67TilOKerCf9dWI0nXIk7XC33Xr/on1CG/0v
+DC4ViUdFEfY82THDQt8YTXY4I+G9OnbYo9ss2kVyBlSxuvV6u7UM+7h2s4eZJwMOo+lA5DKcGJO
1ykIuAH1eO0hdP9J2WmA+XpeyfZxsK4ZQDPebQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 3008)
`protect data_block
Mn/QLJxDklyW4wxR1dj0Y25+ZbBxdVbvTtI9ttVUXk5LaGKK7wnecjRrbYmICgYLnMHrz310ZlbU
womV1mZmb7yR1leg4Ux7f19QimsRPBM6LxabQAhbdNQXHf1Ou1oqbSiEp2jSV/Xg9/hghsuG6mxt
J4ZMr0SsUShcQgjS2mYaRo8YPN6ddOZAzA8KNpiGGbyP2MUPVA3y65SnA5a4Bq46OSL0vMUO41d6
VUbfEBQiIeXCTkpgyjYizRY3UFW1IEcJZkKpoPTcyvSALBhuexcXVJ8/x5A54qShW7InTh92yuZD
n+HjwCjh5TPvb4JcUsKz8WP8BQNyCYoPVs5ALibLeIzOkuG1OtqkBS+HDN1sCk0mQjfJYPjIuUln
xvODRHuGrfj34rmxHm0QXgzm1tiVNpfPDhi55vIOC8f5bQ7AORjxNMQpIPERWaefXvH0Ul56+GRH
Wwlrwe715DBjSTS4yMjeYG4UAHMm7+2MZAH1TF/s4BJsJ9ZuEmmB2eRSXOIQrSfpXKLsI3Dh/g5G
J7dxN5YnQ8mP/MUH4lpJPF8TAroEFwfRGDlCmUR1WpI0ZWsApZg5KL4b9a4tHJECtZv0T/7xr/mh
6evdyCyTPZm00biVQCKswDfp5I04R36N52Q0Xnn+lnDWHg13WwlYiBpO53l50bPTn3pctg02G3JH
wqEHF/ccuhxMGwD6fhixVq4yZRbqdo+ydtMAhbDZH/PMVjX5pM9TTJlgvhp1NuA3HgUCcIhljopu
OlqFHFKbtSiV5OgXrQNLxNs+pYvDoLZCW+pnSj1lKum1rfbHqq0EW8/PLp6Naot8A9x4ktFDkBLK
iiez5u4wBSEFKaY5s+VuKpjl6f7cufQyW+gIjLyePKo4MSb3rXjITM8fWUf6HJwxNI+ojTVhXHOJ
yFYovkwNF+dZ2u565r4ETXGoZPk4X91Z/GZFOkP7+tl687mE4epgsQeH0BTC7EmuhUVc5dG/uiv4
5cRtzsPVXIP9x9m9NIRhriG2PA+15QM49j8lw434MSJ4ggDddwKqdE1vH6j4He4hGfROE/PyXZzH
WzeHBaXWAya4o0je4X6sb9/yt9K2bOTPPrDqHfRSdwctwNUp65tBctlihdV2Qp/RwwMAxOiSvMva
esV2CkgYJFVu9S9YwRPx5/kc9cdZhSdhN7eTidrlQl5fSgt71Cz1cN2JMlz8L9jkH5BiBos2qCL1
nLMwAHgzZurPuZIApO5EXqPc7aRwjh1bGpFaqTA6w5SvFxKMBDGzFJNOdtnM8QuzL59WGMhN/dq6
+fKah7WTbVo+C6m1RHaa8snAZPAGWM1kTZq61atEjFmJInS9omAsoP4OFnA8/8zqkWKJbT5lgvJt
X8U3vFEyG2ynFPD8CZ5mpLdBE15Uk2ErLexefPCZfmW1r7L7npT9iUT2cEi7O7/rJmythRnmecPz
CXFYI9pe1FfXPdiSBqixU0RlhShjFiraDidc9Qd+BAmyDiN3cRx0+sRteJJM6My/Xoxr4bWxbasv
MPIWe3qqA3c8dtpclQvCh5547ohuSO4vnohkez7o6ZN9ij2QDSYiadKonGFEjLVB0tvFObfIACxX
pSMJuD3pgRgOoy5J4dPqm/hPVq96okK3JMDzCMMY0XJDYEkWj3sPmJVZPrrK3i99G8+sbFw946Sj
YFZwpIPd5fnh9j1d0jhSEwiWjxziGmrFb9B+h46ZVDFr4eguc0bP3SHc2xTFhPQg2pZ52E77oQ6t
3NgJiZ1rAAXdHEoSZnOwgAMYwnCFEQqR++GUz8DQ/xWv0Rp4mxuSHmJKcB3UZ3XO8z4im6ujfTH9
pv5YoiSutFVFov0HMWoBtGg42CdgRVOBH+jLkmxTh+uxG4/gNS+VpIRs9PNfgvpaZGktoLW7tlxb
pVoAQ07CzG49S9WCRf68RQbLRgUrj8c9Y6mf1oxNtealWqydHW5m9CGz6rpVUCq5MThKktw2ZFMo
vA7pbwGOQgi5fHRB1F+b7GCqJVGzFmn9dOQ2WmgNbVGOCOFeGMPRrpZxLfBzwjim5F/KcTVrTWeM
f+HOID2jzLQaUZUnG679AxAOOL/Hpd92drE3lmTHb30uY2RKskK9JqusxpzJyZGyP9zcdTMllP3D
4x5Wm3fxkFFbcXNHlmGYmZWR2uCmyrpbncfpu+eTjzEgUAqjFKJPhAS89Mk9Ga3SCqNVTcR1+FkS
s2xnRHMQtRs+jAAyp5lnOV2PkxPyfK/FApWnlH1GivupKtId8S0nt6Cz5k6o9XZsDFuCrsL5JvQC
w3TQ6RuIO2CIUgcwU9RjQmHWED8iwU9mjkWS1RT8d/TcoT00rHLvUvtFZOVLHmd1f21acJ6wu1/r
pxdLe57W4nqJ4nO7KQF/Bz+Jf5MK3vWrCIyGbi06nKY21t4m+eqESQfFbaVOYzYw5ZqfbLM7HWUt
FJghWueOENAu/GBYiT2Fp5BvLcTaiBO875QnbkvlBpQm9sdbbkHxTYLlDO0qawQR2sva5l8Bwg99
jRoKRcXZKW+nvC7Y4OcjVTDbGPlwci74mqTfmTfA0ZmuTRNYPBzafPiLgj5V2veogwx/hFCtCoh8
BQi8q4MyjynCakLN8Cj8hEo2dCP7+Yc4+nHoT4RToFZP7Cp03MMyKwWsGZFVOEeFUd76qH0YLnN0
oKXDdY0BejmGqwTXRynzfPKNeFjHfRHnz4ROtmsxTBD+1twYp8K9/5pdPBEIW1wqOKjCoFQZ40l5
7WjjnLY9oG55RUUBMZ9QqzGRj2fKK5sQLuzvSrEvTp5qaRu1DsUKcg4jfzDpy8UnixhJtkwDY2ER
kE8Azo38iaDyK9Hh4cmMsaxoFp/yPuJVMy0wx+EQPCveXBkATJOGWsrhbsemv9yi/WUMgaSJkK67
0PRJVofdtiUytjaghpGGiO18spXa8FPDk6dnHJ7hO28yGKHNyoYLf0h4oLDK8U7ySuMFoOJZznvC
TwVAB08Ozrn9bgxx9kAUsK/YtFCf+/MehWFoF6HLRziJZSKw5MOUZ5XTKwqF2hW2mr56EFD6UoZu
ZGqefqP2yAqd0N8BVjQqZogfJRhfwA/WqprYmAZ4YEAdiTT5FqKlDsWdUBR3X685a9H7K/o56eJ1
ux/LYvfSlLqqa8+0MLm5eDIzPK/JFyuKGHOHCTD8T28dCMJ/I+A0C4EMS1qH7A5U7r2fcZ2XNf0L
a2RKsvM6LrYjGVH1otfOiPrJGGB31ebxnp8BpF4xo1VMCL9Lo+/MhccxbjGo7ezF1kNWzXoaZNPQ
6rnKJcCy/R47UelxA3fznw5tz+uXprTQP2kWDB6EdebZZ/EXUNu9X9PfoJVVLwMf6ubyT2SMI11w
1ZZxjIfAMNg38ZYyGt8R3t6/C+f3i5vVGFjeBsWqoeqHPmEeCDDWG1AJmOki9ZTPFJ9gVYCOcFxj
J3GDuK4BC3dgE2v9a4Y/u5lY+7sB5T+/tmcrwkKmRpHuvqjWg1B0KS8yaML0a2mUqv+ne0S/jGpQ
mqSLCmX/OlWd9WumIa5R/HqAl8QoEm6R/pVIALfflDyxW+35IIb+V+kpkxJwXJErW5MsHRL33izE
YbvtpH4qcGErZgYHY5Js9CfHA1h2F0ZW944K/3vO0SJ0NLLSA0yWfHcJ57tly/ZucSyelOlrpUtF
DO0KxPFVLD1fElFMlfQAp7oh5+4+oHzooqziuFJaQZYWVZB/cjBJk8SeqOaGdlUHujiqPd1GiUsV
NuIK+Mq9UkNcjU3yQQtXgTkjB+kwdfFaLf7Vo9f4nhE/RWnPcADCwEPKMw3ptCgozwXQAWFFQD6b
AIjLQayyWKNKpjEfB1wYDNskceIPXXqNoNzppp3W4Ye99G0FRYpiklVntY6tOPWDwukD0RaaKhUg
d9h4l45tZtZgH8YdM4SmcPO8o3xya5RuhVQTJob1YqD6JJwNUlPpD+2mNf1rzgV5wCgoC0BR8MRA
v6/SBA9hwNZwyMNEeuKS8fpk+KnVaETM/Yk6CiiXH23CBelM3ORUZ5c+KO8=
`protect end_protected
