-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Jhn1LVzCb6+ejntjSsgDMFcoDNOp8kkMPjuvGgSZhaWCMv+wucncHH5RvD12rnrIMUCGgUfr7/7I
34DKyqOS8ach7/ax1/jU7gjnIsNUci4g5Py0iPGzWGeDX7ekKyDKWNCe3biNLTrdDmiMqk9HUx7N
vQKGLUim9Ox7c/6v80EAe3SWDZ/QMjqdUNK6YXXIJXI8ZqiL3WEht4Z56XWEVGInanxijjIzuYzX
9KgHcUVbED9xLdtqHksLEGn544bl5WTen4SCXGbMt81gCJwwlH//lTLcg/tpBlNq7/UlDYBGk9Dn
pk3u94oAT80z/0J+USok2NP2fQprX31mwcIw+g==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 2736)
`protect data_block
WRiZIKnCgEEpTLD/gJvQKcSTYjI9QiVltv99FukYqNv9VmQaiNvfKbSY4T7h9/7zyMA/xR1RKWWS
fuTgzR23glFt4mrGkg91wasVB90PAAggFG8dUzY15wmIJK5ioAZn8syYT0B8CezYEtfP+8+HnxJn
XVy5dexmQHTmej8a4h4Y7uBTEfepC1QkXzcx2NWRxRnZ9iEIwZkQv+Fgd2/ZDTnMm76oGgQP/cTs
4xjoz4+VOZh8SvTtHJQPeRJ4IKeY2nP77jcIsCT/W50gxk1tpZoAmoXyyEZj9Ls7k13vuV3V37ls
PoARyUqP0VEb4bJYTZhtB3xq8XAfHAp1pG80Jg4D0h5Bm+xc1Z5iGWYea2fJLxiDd522+GEiwHaO
Kjs08iQw7HdHbfnQlY2PhzBs6VHy3Pjc/017rtqFVxoGaJqBR/RCzVseVxZivJAab6jON2rGMSSQ
p6fwm132L0HAb/3Xqb/gubMGJS8K8eTYUukKzFwdWN4yisLV+u7MXzgvHQXuyJaHkTyMcjkt7A2/
FKBcydjgQ3anHlYtr/K80FlC2k5siGoKMDUOtKNA4rJOpZUNvkyJS+M0UuTGGisNRbb59+COGOsy
y1r4oOmC8jiszJJnFI+juT8xmx5qi+Xniu40Vq72VuAYyTqWbujBr8mKsv52VmApoWTnbR3+MKxL
bgoKHkIwULlg3RgS4PS1x6FKvam3p+3Nqu4048BeM68xaukH+ia1mCfdFwCwZX4W51YI4RczNTcd
koW8FfcwEp8QSBkJo9sSGJsDqAJSF7SliN3F3fgtfQHhoelx2hbWHO34L1L4Ib9XT8eNAoMLhLve
9GGCKZvzG/sodxu489LSiQgyZ4h1J2ED4YgsSLksM18SDBPn5n35aiTLKECDHMSq4AQdyjd5nGtl
YPk7+WSTs0cegUDbEGpigqsKPINhx+2iXj33HCPoHj/AuC04Lsz77diqa1+gQC3cGV81kmkgC+fN
lP9GD1zz9nK+HKYYv6auWb1B2N51Pflq9VuyBZQd2qCRZJ30ldhUN2fZyXLYgK1qzGEtNrKD8VAz
OfVYTIu2oYcbUYh+es+zcd87WNoRTqCajGrs+VpkzWMpcX5/RxvsW4I8oakQ4D6aL/Uh3S0NJafw
tqHjidfbnzyuYGn2w8UbISHHTDH5V/oYiydZEg01AEDIVvb6lSe++m32hTfPlGf+/sw+aOiZFmbH
Gy4XDrztZwh/modNkN9XpYLTx954QHxgk7U/1WEtyJY9KZ9xIKGw1wkxNp2EeErLAHcRS590SBII
RUKGgp/1Rq0dyAAjazV44oJ2oegzbmRNtHV9c9ZlyKlMtA/Y17PWywDXsvhlUBB7QT9VvVRCWbYh
k5bOJp/cG0qSUS/zFROuVeaGqqpKcF67+LABoNm9I6t4xptdvc6SSLu6z4iCBn9cDCBDEFQfywgK
MRNXdm066IpGv85ttjgBXuu8ORhDWeaT73Kns5F6PWbuWmaf6qOLDoDdnN9wtMqu6ygxlmwFrTZD
vAlOzv3CxhDuisUIiqTQIb9it5rbZLR50sANLnLAwb8t6wuEPtmPZqIfcOGksgzOfHezffFOrVRp
D0ak7bcHqZ7zpX+M5UzbE+n8aTbsNZQT6c1NSEx+EY+Pzz5JlYPbyxlgD1Aq5Jp4w2l18YRsdqCt
syv+A1hgv9GhZ6bA9zxtzqT82rbajoRVk40uPgk/FjcnCHVnSOw5rbXEbjHs8XQu5OpBLsVuHBg9
zt6PxciDWtu0Yj6v1RGkePMDiHLd3HBGU27A6s3TTjKfxtPg/IoUVhMcKyK/FbbnxUJ+3XNcsfGL
YsEVpx1ND9shEdRTzHJQ4lmoIf6TI5V2M0OrKN5KxKQ5SOJI8Kg37DYDWAhkJlC2+9I0TOeOUTju
hcZSumke4I3GWjewd1WrxpPf7K7Tvs5RcN7Asr6bj73FKhsWn2nJtTbGqw9lLQeoyGrcvm+NuhGh
6AJplSjSdNBOt3PpnFzZVHtUbA9ZCfnrwAZmDSQ6zy+IYI/Vm5ETokLH4FXoTJJ6YfqO5W6oEPw/
aUJXztVXfgW9jVcTGkY4Tnwcevi1I0NLzM92p3VSiSGPJ0h32xvdsI30dD0KJMrhYTNVFvNd1KRV
3baJIfjwHxgyjaFN/WdQMAq+XiK4EhC4N58qJwDJY32hb74Y0ZvlBBPn1UswJSt4OAHAfxAI+1ei
2O8mt4psKAY2MwGJSKy8CzvE9C8aGrWXHLdZnn94ubgejdEoLd1MjUa0OiGn+y4Y51M840GMzRSl
g65vSNG+gW5ZOt2hDlr0Pec/snWz0Yyr614ldFHHsiQFuAV+Re06jjEY67fYMc1EDz+pQsiXXEGC
nBdE0D3Xi+Qcs3pVwggWSvg0ni645TqxY53nxqiQXfP/Zl7offNbjR0bjvVlmyQHVZsHQIAPw5jt
Ha1J+zWzu2O22Vqaiv+wjOk+ry7JgLLOHcV9j3p4K1+pi3vhwJWWEnKbDGmqIq2OW+RhsWyNlnRA
mmtcX3r+9XJojZExUEG/F3Z68WhKtS03s2be2fOgfKr+NKSoCztStvO6ZtuBMaZTFvYnvsR0+717
rB3+XeAjYfr1xsz+j/84Vg7OclP2hsz1LRA7dMAX+20gN8eFCTQSgXiIcl924nmxrG4JoapFIcVH
+UB+ueUJfFTYeGNedRod0VWQSLrVykFKNZPbqnDmTtzrFKbLPMfVsl1ESVbbBAPWJMPsIX6T1QNS
+64Itwf4I18JqTfDX29rKzdH7yV3hKqGYaedVJxWCCZtwCN9xgiy+DIiYZ1IrS/A19Qv31+j3wo5
tsjPUfG5CZ1JSHH1Z48ToXW15shtmplFbsz+UI7zbvG5aYTcBxnJLUhul4gHrA7a/5WPIA6zI7zm
12NbAK8n4h7nTa5cZZhl8CDJU/S4E3jEy5vqwHNGVJtlzL3uDcKM0MkdP1FeOqw+vV3KbXDuTlws
AW8eFvhcagNcEucdN65UuYWYX9dab9AgLA9KTj/yr2PoCiQ4MxUYsly7hkkvI2NSGeVXU08PdecL
jjXnK3RYKHelyuVyzNj1P3mYOcGSOCsqQ/CwOz7WboH4ZrnlDzRlDzutJfPrpS9p9lL1tUWIv8Wf
mGSSIqen5bUtbZ5XkxEC02/vth/6R1vScesGey3utFq/SUBZpcJen8LVFhsePanKexB8sDsdcyHf
psp55lQ+mC6f5DdytYCC4iOLRsT6NAtrGbDPKp9lM+00Gg9/VWEnQKWD3LFdiOKSD+T477BoXqO3
QhUsLUXG8tYOz7Na2RiZmhAaJzgIwkFB6CdXEBBn+sNQQPrAZU364QX8n3kqhkf5JfAn53hZUB9/
QoobcQzWU/5Vz5h8FgGv+un35knFEnlIVS2izI81ZNrSvVSLjWvm8+/DLydCXhVvR/UlRJhonhFA
nHArvY8t8t55sk+HarE23iQ7nO3BIKsg6NUpf+slwz3JKPj/Ybn1V94qKVOC0Srd3b/ACBzDp5r/
WSpuLYVPGfCae/OJOtClQ1Q6VFhVFtynlqtuFxVXzKNwA0BGueweDXlQI5y4Zt36R4PLMZLQDHnJ
nTY//ZgdgdJMX47ZRQkZNhJy9NHEfMWaANWMfvBFsLu9B+iEUk4XgfprukTXvT56im7U6yJPK308
`protect end_protected
