��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$Rx�y�<��wA�*;�x���@�̦�W�X�fa�M-$u����n~�%���P�$��W��kYَ���P7�?UMfT��q�6�U��k�>����~�\N�(�����X�e���/6U|)�X2pF�]$h���d.���9E��WG��L�X"]�Ad����ľS���8od����e�GT?y	7�������ݵ�^��R�q^]�鍦�����s�ae���h��L��P_���ާ��YЭF���'\��68�b�[����w8�[X��V�F�0͘3����q諵�uW� �h�u\V�?@��_6G�_�*�G���B�絉�f������[�G��U&�����~�F��AׯK1�`c��[<��FY���4I� �#�G��x[X�=�Q1��`��R>(�w����R�O�?����7�,(�H\�#h(W�EH=�������yq��Ѿ��aF����:�U~m<|��.��0=�P/���4ǆ���T(���ORx�����h��)�hN���n<���e+�f�<��Q9e^�iS�d�h8|�O��$��@r���HQ���	rS����e89��;��X5�
�yd	3�Z�ɮȣ}}����pmMc�����}& ��IC���=���ey�9M�fi�)�w�9��d���5"j˰��� ���J�̘D	L��s~gpȦ�E�]�����Ʈ�iQ̡��o�F�Uk�q(�l���Ŀi�f�VyH����c>$? ��U=��>�[c)��-\��1����}lP&�*����B���_Eb��~�aKp�M��Z�Q�'�U �#�;b����s�`�W�Q��OΥn���q/���<����i 4Xp�Pcو���ڨV������S��w�tִ�@6�'p.qֲ]۱꽝
|�c�\� %�u�i���������~�<���{?Ǩ��(�h�"NB?����3����3�s	�V�뤰a1������f��ؔ���>v�a@JT�%|1`-�R�$Hz�S �&ex����9/�J�E�I��**/{�ȉB�l�<��,�l����bH|j+��Q�"�iz��K�9c������u�E�PP#��c�JɪT��L�i���ld��}&�$2mC�V�����:��0z]����͑��f���}����90��3?0�r�۫�2���cX.d��K��Bo2�^�'��,��U�t���S��1��M\[�q�r&oEȻѿc�P�(8f��:|v:���9��7�z�w^��ݫ�י�U��y@��W�Jowy�})�k�/}�	 ��Eq��y��9�
�g;r��J}_�㚜����Pe��"���x�����'V��fiT�(���DP���f/D+g󿅱���ew>r�-E�'�L�%�s�z���Cc�X����+0k��"5u�Q*u�2�P$���Vߢ�N?�Ǚ.(
3�$ȇ!υ):���=
����9E!]���G���h�ꪩ�"���1�%��/�����\אm��`	%�o�=(0�
+j��Z��M���Kg�C+g:R?RY�i���H육��l*�ߚ�tE�Q�"`�C�5Kt��F���1�W^]��wgUY���ta�/<c6�����i�މ���r�l�4~{��W<���j����#��°�<e�B�㥑�F�襤 @�')Q(8�X~�-w�q�d����:I�\>��>`0*����l}�<�<ֵ]^t6�s�ɽxV���mjh���w��z�P:�Ȱ_bMQ��2a�X�~=#��Kt�0�j.���3��@���+�'$�MJ*j�D/����I�-^�Z�]x�QO��~�w+y��a�gC&3?�D!���L*�n_�i.����_ڈi�j݋�L�^e���R�$�G�ѽ瓢A �]n��qJ�v�M�w�z��nĦL��$B��{��[lL@��z_���bZ���n���h-&`@�p@%M���}� co� �q,6�����u����+k�ՆZ�O�~��y�&e��]�9i���-�9o����@��s ���R4��y�k(�Pژ�b",�jj�(m8�sOЋ�wZ�}��IxIt�0�:�*�E�,X�pg����q�����Z��㯬w���.����#p0�U�m�O�p؀~�~C;����b|�~^	�7;��i���%�l7$�zN���u��Au��YrU�7h����%�shh�dx� 1rㇲ��U����v{��X�w�6�lA�e�b���#{z��	,�@pT������#�U*���d3�2�"O����&{�!P	����!�<�I	r|���P�[�v��ը�]�_�ڇ�XC�GPx�)��p.�h��i:ۇ|��������m���:�'�b��d�[���s�Q��c���<��p�?1�[DP���Au!��׎	�������&h�
pnξ�t��ڊ�>�UC��G��H��4��d�{=�3L����ZC�Z���_6J�K�s=:߉?��:*h�{��5/1����w(�/xV��=r�ɝɮ&�]T�rտz�n�͕r�Q��tn%o�-H�E�j���ւ!�g�T����>�1V�h��t}-#��fҡ*��1%,%�:����F�8Ơ��H-�Á�19|���������u��=s��+��|�B(ԞBR��gU��7!��"|�7k�+���2�H���~<[k"�Hܲ�qaf�L�c*;�`��u����ӂ�	B
�Ex{!a�\Jf�(T�&�<Sc�]���P/���T�z���]s��v,�7	;�4N��wW��6��n�1�y��L��ߍ�p�A������tDew2���*l$����������F�>�b]p��5����;���ܨ���/\�j]y�;o�i�!�k�q�5�TrqXo,� �7Uʦ]q��I�1���M�]�tze�^_��tvkHrL[޻��Y�����R��Jb��$��>�����HY<��i �r��k�#��S"$+��W�G��S���+*{[���#~�D�L " �<����/#^���f�ԍ���=$+\��p��G����8�ƿ�N�o�m@�;Q�U��)��0)�$��|�3�����H���;Q��
�%�&A�Ti�D�W���&�����W=lpyg~F��D����w7�����,��r�*&���W#�H�By��|s~�=D��)C�����EQհal�N���xCkV.UV�m��U
Z�l�����W�,6aٱE�ģ{c�A��?w���$D?��:ǃ�i/��� �λ���X�+VGX~<�K��#uULiٜL+h��N��w�H�_ �)�k��Yߪ���òΆ4N&��$?(l�������0�5��M���|Zr����{P	5����4����������W�4~��" �};��6��	��7��lP}�@.���z��N���k��i�/��5?~�^�/���7������˦A5��#�SK�L�1�&TS�������@/&�4V��)��s
H�(}rQ�S�+���͐�X�JF1uB�lȄ�p9���V���R�f��GX|om����	�c.ҌCT��ꬶ�7���.`"A���_h�w��U?&���ޒ�O��i�_��+�~�����ݢ9�n�x4F*N�\�H�'�b������(Nb8��	
��/x.�|����Ф��M��{��OQ�}�"��!��c�W(O�}\(���}�!_��t�c�4åL�
�o���Ye�4��]�R������ąqW-kk_�/v�Y��P�� �p�C�D�f>��H[S5ېX�WE�������%��m H�h��Է�{����Y������<��б+��^�U�����+ٽxB"+j�
�Z�Ql/��{��H��FʄK��v�����7x=I��r�ty�|ҏª�y'+���8.A����s�F꾡���j��7�QP��&�� P� �>�����A�ǳ�v��_T��W�iד��oFd0���չ�>�l_����x(��[_��%��}W����yi����uwD]oӉ����t�'�c=Ƚ�E��}���j��6���z��z�n��L��C�(^cj�mNN�.��U)b�#��j�:����C˝Y�06��w�d�8�^������尜�t��r��������:��w�
]j.L�,��7mx[A�ty�AJ*d�ދ��ޣ6uگt�ҕ; �[a{���Z&�\��@{�=����"�3_P���xH�,�@�T^��7ڪ�	����1V���Y��5���j˞�$�H�\ܜ��ֆ��s����5�%�=�����6�E����*LG�&��s�փ#L3VA�)#FQ
}�M��]Tg�&X���ӓƋ��v�LJզ�Ky�H6�	A��=���΋�lH<��0�aN��H3�@��/��%.��p��_{w�?���%kt7����B�W���^����w�l��E��y��sK�R���%�i�#�-8IoX��V������!��r��O�^���;�F���8�i"vV��L�(�W�)EX�f���0����\_ea� �1ndS<���^��MX�|`vZ@h�N�v�A�ÐT/Ulu�A"��K`W�7���Y,^Ҭ �>�� qd�Jy��y�.-OQ-���h,���� ��	GX	���נPg;��-bl6����yʏ�Z�KiӺS�$�������D/˦�W��a���ڀ_�O��^�5W�H��L��b�uB�ڟ��P�u�� �<�����s����Q+D!���=�"�䡂�_��{F����6S(U7P>�����x�E���j��Tjw�af���a�-@}�(r�n:��.��z�
�}�:O��q�;~u��S�T��k����gٮ�J�g�	+g8D0���m�d��B.�UM�vv�-x��wXגȷ@��z��M�[��sѬ`n�����4lc��2������+Ԝ��a=9��-��s��}��	��[���Ը��}���5���Ζ��\��*�B�u'��";Zj#`��3]�8ʇVw�EX��+��}��ۖ��`��Z$L�~sܚ���e�R˜!�]��BD/�/u��?G gK��ڰAn9��>呿���$��"���\.����-l ��eL���#���n�ز�Z��(�^=��O�[��:���1�u�RKJxw�Ed2���0`��׻��#J�a�!�M�Oሞ�P���
�^��}������E���Q ����z��wu[�0!��c՘���K�>y��2#� �خH~O<T�f��@�p����IN�{=�������"�@2��66	Iw�˞��&�X` ��OXy�?��h�ǻ��G|�6�J^f�މ?6�3[$�o��!��-�G��6,�ś��B��4S�4�
�d�%ځB�e�U�˩�un&�8O��gF������b�%���dQ���|�	*ˀ���(X�X�PB2@ms�Ӯ��E'fd���@�Av_^�E(ۛW%�S���/�}���ŀ�|�GgA?/����b��L
``
#��,X� �/�7m"%�3Z[�����*'���\T'��Z������!�zH�3
���Ĝ��8l|��{�_�a:�}����oX���S�}.phU�z�B��QKS&�i��&@A�v�M�h����z��W��b�S�a�P���ʔ���I�*�7KV<@\e�m=6N?L�bQ� ���_�:����8�GLHcJ��/´�N��M�ݕ�9̞:�Ga��?^? ڟ�9C*VV�4"�馈&hމv�����d\���&�k�y���:^���Grt�Y�?���0mR���(.�]}�P���iR� �g.������7�����U^�8����#7�ؘčn3�4�[A/���/����t3|Ҍ1�/!�e��?�OIFKv�b@�.���@\p��1Ay�}4W��/��r����SW��g���=�,�0�uM�e
��i#��u�-��Ey����a���Z��������u�L�%n��4�h�{�+xn�/��i<��S7�.
]��(o�uF����U��2u�����K,\y����Go�N
�D�ҋyG��i$� ��N���=�V]1&8���1VFX[ڳ=`-�G�]h`.�V��"��]�Gxd
p���i���tj��}���-�8Zp����0�]Ư��f��k=�� ^Rc�E-��_��&Ҡ���0j�xF��̕��{���u3Y�>�qvj`���e��U�����F��R\�&��Jٓ2/^(o��!�5-cZM&dhc�]��E��-�Vv5�ﯻs�}��UDЋ�r6a
�3Be���m｟D͠���i���J	0(���}u�<0E���TXL	.�p�ir�i���!8���U2 ���m-pݠ��y<�E�.���8�v��d��Y������)Y�y�������6�/�4"^�Tt�u}����h�ɸ{m�ei�J8Gv��*{Q蜱�^J�y����ǝ?��2r$����ެ۶�^����y[#!�ϙ�\����s�
��ǚ'��
QLKR�Q�}l^�M"E.F�ᑱc�X��҈���C������?�5�R���}!�!m�>��}����Ɛ�ݝ8:�/;��R�@+.�[8/�H��t�iz���������I�X�)ys�:dd�Д���{i%@+z�e�\����sn�v���Y��|��'���n�Զ�&�Ԡaǥ��Y:;��UG�&��jQ���s�n�4즞���}�_�
֎��3#|���VU�����iXy�2�;��M>ݑ�j�d��v����y�^����I �Άi�X�.�eLۤ�_��d �;�����>�c�$k>��F�[�%�$��^�����)*f�E�V�P#s�C
��z��u��Q�GD��	�1�6�	��`��f���ˍ��p�5����^���X`E���:Z+Ӎ�\V�46_��N���=Ld���{�wh6NH��3�Y ~�SJ��(8{���%������y��b�M�R$f'|ς�`Wܺ��y��r@����9�Ȣ),�MA�Ҁ�V��|:;�"Icr�]�7���Xk?(��_b�S��D��Һ�&��/��o4,�����ϗ�Yjǚ�o!��S��)JM��A!P�j$% �5 ��%3,�r��5rn{�߉A���3��M �Y�3�� �K|��Ȧ�4ced�G����UF~�oN���E��XHΥwN���m?$J_�OS����E��t���[K{�NH'����K�l�|Uo�������H|3Oؒ�c�gӥ6���j"��̏�ݷ�������,�3�Z�[G�6#E���i/���)����{�V�$�A���*;�`�LT���)����W3�T":u�ϐ`�C�͸5%v����͚Els�G�L�쎪�(�Z�Ìf9�U	�<��k��KiZ:�<n�I�Z�;�񘋦2ٖ����e�{A� �Q��d���xr�5x�����}�VM}�5��2<�,L<��qYe�'&w�;�-���'�W8�V�E��ᖆ��X��<?�n�	�M�eH�)���*��Z�Lp����ڧu�n�,����T=*�L�P&���:e�:�j^���Ɔ�Jrs���MQ��]���X�Oؿ�ɾ�-����kL�����8�25��/7J����?�u|f����ߥW���Q����p�ﾨ�/K˧��r�2XJ�к���U8V��etfA�K2��k��b���Ot �B�]-���oI�����"��4�����ߓ�>?�k���j7��ϋ��3�ҌIn�T9;�5Ç*+��&D�7qaM��k*��.��z5Hd&O
+�ôVȶI���#^9����j*b
q\=Ǉ�,��D�u&L �0n_��F��8	�ѝ�DgD�}�Q�p�	�8H���+a[�~%���[B���$0�%��K�.BɁ���Ӊ�u��^�� D��n��k���D?r)[�ݺ�k���2�$Wtʒ�9)Q��Y�3B4����Z��e���Bj!S��S��[�-ʞ8�	2�0���H{B�4�I�ݵxv<۫�@�CT��s\�ί�L�u���ľm4/޴�z{6<qig^6aބ�6h�su��ôܫa�wW,�i��E;TsF� ��I�}<C�a�IE��؜��_l�O��+���P���Q?�Ì&>N�]$a5���펡"]���A�,bOSl	�I�e�p��-���eR����&4�Ƽ�l{myb���p�J2���w%��kgDe}�x�Ž����d[F���W���i��P#Xc�Ͽ��JN��D�Yk$]B��,�7�c��.���:���p^�<��������T]]q��㖵B��+q1ب8[�A\���4�G�"�*H<PY�Ⱥ�I��~����uo��A`[�yvUA��������SD;����SöTq����Y�-�lO@��