��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$Rx�y�<��wA�*;�x���@�̦�W�X�fa�M-$u����n~�%���P�$��W��kYَ���P7�?UMfT��q�6�U��k�>����~�\N�(�����X�e���/6U|)�X2pF�]$h���d.���9E��WG��L�X"]�Ad����ľS���8od����e�GT?y	7�������ݵ�^��R�q^]�鍦�����s�ae���h��L��P_���ާ��YЭF���'\��68�b�[����w8�[X��V�F�0͘3����q諵�uW� �h�u\V�?@��_6G�_�*�G���B�絉�f������[�G��U&�����~�F��AׯK1�`c��[<��FY���4I� �#�G��x[X�=�Q1��`��R>(�w����R�O�?����7�,(�H\�#h(W�EH=�������yq��Ѿ��aF����:�U~m<|��.��0=�P/���4ǆ���T(����]�┎2����Y�����U؊�ȶ3h\��QK{�g_�_�$y�+���ln�l|�P��Z@z$�ϧ?_��i��牫g��z��Ø�S������	7�7N|�3"8yS5���A��gu4�EV���Z��s�+ȱ�X�++t�2�O�E�|,��?�:�%����[f�x���S����a���e�/�`퉙dDm�P}j�%�ٱ&7ٹD"Ed����=�V%J?P�z���:���.ٛ2�9�s����-4 MNăI�L�i�ۙ�X4������u�z�����x	g����UL\�;|=\)UU-5������0��9��D�K�:pdN�h_Q#;�{/m��/I�n(>_�"�s��V���k,�f��s{���ˊ�Ŀ�lv�Kn��$��,��eb���U��e�N���ϴVP���"����+�Hc[��$��I��j�9�ogC5��F`_��X��_�]]]O�Tn{��S�`^p�_��E��e����~����H�%�u
+a�
ˑ^�\�t��N��֪y�ǚw�ՙ�`X�3��=�֙d����1?�<�K3�:EXuz�+�
d�6�ẵf�ǹ�X% CM��h��R<"t�"��� ��1&�qʍ�i��?�Ё���64�%���~#����t�,Xn�4V�X2O���)�4�t9�o�p�ׁ���P,��h5y�b��^��u�3P�gd��M� ���m��D���
� ���:��̷�6Vט�W��/���	��W �M��AG*���)����L�h��"��2J��t�Ӝw��]��2�����Ɠ������Ң9�,���5�M[�m}��K���3�?�\���ŲV�n��Vh�Г���R/mD�7VQ-�W�v���N��!�_*�8�H�'��0�ǐY��դ2���<^˚��>�9�{ć�_˲�;��բAU>-����G�P����_�`�})Ύ����X�#�����E�#�\��3�o�qOhR�tb��*&�*���iGt�([��S�}w���r����K�+D�pb{w���m��Jc���w�������_�,ynu���A�g�����N�4�D6�1��8�{Z���}-.����*����K.B)-��%�3c����$6��o�駇,.�8�t/1g=6T�|:�Z?��Q~�j��F+X���*��L���
�PKܸ�K�&qs��tط�a��R���� 3���2�P��~�]xg�����]����} ����'Q >; ��#���3
;��Ws�l'>��)�披|�G�Y�y���u��͛q3�8;~"'����~��K����'�X��F)r�� ��}ǐ-��U���[�NO���+m]k?
6j�����{�y����&�0H��$��_~�VSu��̸�@�k��Ns�!�U�b�(��n�����H����C�^X_��ܬ�>Μ=_�m'����7�vކՅm�����-VǬ,v�4O��;�tOyY����j�C�o��+Co�|ذx���*ၻ���O=������l8/��S�}y)�[��r���}CwOۚ���=,�����b9��<R�Y
"o&��^�#�[z�3�s�h0?ͣ�WskV<����(-�#����[�j  ���4q1��.��e鯵�Sͧ`�zY�T�wc%�3Zܴ{B�L0�Q�ߗ�"�#I�+�G�c���~]���Ԉ	i}|H{w �BP�Ve�>J�(-/��W�#�.t��mP�f������sz���hG(�b��y�Rc�Ǡ(���:�sA���i��Z��*�*C �;w���
��IN�_��r2	��c�: ������xx�uK�^����x�-�ojM1�<�"2����lv�w�'��JX��8��e��b���asf�_܏3B#�J�Lb�#���|xķP���%�Z�X�0������>�hÉ�?����ǯ�ӓg|y�e��܉��t|�%?������Rz�ڏ�����(�W�@!�ߵ(>�����<�P~���c2�v��a�F�8mO'�VQu}K�ף�ԝ1$h��A��=k�PFWA�Lk���l\���ȼ�����8�r��%�@ �r���/ji�z��Å%�OkTΤc�X����DN�����3 5�o����_ 9G �~H���V�"ƫ$=�t��K�=��E-�*Ƴ�h���:G�W���u��'u�ϗ�n(R!m�sJe{�AOc�N��=�E�*Lk��$ʱ�;�݈b�,��Ȋ$���ϫ��H��N�|�QLO�=�~�)�O���BM����3'�ã���i2覨��7��*fR|����x}T$ ME��eQ�_�*�A�vV����e��>� ���R�#���� ��A�"`�4�h/�v��\�[N���!�#��ɘ\�i$B�^�3��շ�H���X��'�T��HgF뙝j(��)![+Y�w���"�u�8�Y���SM���X�#2ًY�������.��M���7C�B���'�<W�Ttn�ﶟ�f��3��R]���30�����׭���Z��=�@Nx�]�t��LeJM���X���\+ICH���<Q$��ϊ.	E���(��oXp����a���0${Ђt�:"r]�w]wa)M\�a��N"�hn��WOJ�+�x��mMK�证��C�h����%0��)��o�
]^>�[n��&�Ү(�mS� �:�x
-oa0�F����M:
���ۋ��d�/�I��W�����Mڷ��Ll�� 0��3�� �vj+���T:=��1D;�*���F�+Մz�M��3kq��L�
8��S�m��Ԥ�@T&2�BG��g�c��Qd��T�ii�ԟ�i�|Zf9Qe ��b ��aXZ8X�kW���>sd�kE�H@�@�ɑctqM�<�ߥk	���M�7���MT�R����G���G8�T
�(}�&	mG�r��v�\U�Y����,�������L<���({!��{�a0��r�!Ht]Z�X���3��Ƙ��g��Z�ܑᱭ�6���:��2�2�������-������A���S��1ez�6��簖��|By�@ͣ<ӖT��"<���,��g#?f:E���߮������c̬�0�&�����Ppt�q!�d,e� ��I��K-�ڗD>x���|)d���n��m�;I=?��A!+���I�R�r�Ξ��L�ND a�V*���ؓ\*,  ��3���=�`��5px�[��e8cW��x��寭�f�U|��ov�}��;7Fw�l��bm5� �8��@Ds>�z5q��x����T��	�
�8-ߜ�!����L�4I��/��y��ٶ���l��C�A4�-��F�&�cJ	,+VDTߩiZn���ԗ�u��RB"�\
���t��']���,�.��/ti�X�0���g�W�k|0S�#������n�c�H7.(��0�S�7�\r�D#��&�4b#o�yPC�?ag�z��KƄi�5rƔI�gg�����Mx�L�����т�MgN2��S���Q�V�됸Ez����XYWzQ�ԅ�WWB%	~əd��D~�lg�c����U�[cy8�_p��O{�(�ա��IE��-SvO��D�!c�sϤ$W��!&^Z�l���9�ws4(c�On_
!�xU��4u�J��z:3=�c�z�'�X2����Y*�
ϑ�Sx
�g�1�|�����!Ì�t�qءd��X��'���'�W�Z�PY��`�f-g�흲yi{�wt���R���Ѓ�;�����Wr�+�I�(�)�C�TKr��i�Ԛ��4�1�v�z�0т�8���ی>]VK�(x�\��3_�{U~>���K����������GW������ PV,�!JUVX{l-Y!Pt��P5avs�>��]Dd)�2������0EF�}Վ��[���U��+`/"��:#>��L����Y�C�I�a�Y�k�i�↣puy��g'�VMz�{ܓWKܓ\��@�	�����ʹ��X�>X�r��->(�bֈ D��Zka�_m����a�� ��U����H"q��`�N:�<~�E?=�ͼ#�Z��$orj��%;�(��C�_�k�A�c��."���!�{�#$��
�V�����r�8$w�?ڈ���F�����_�plj۫%��-C���W^i�=��uYqR�+h�<\7��7T6�4�K���,��?f��N��Zo5kh���ح"�U�]H��~]��@c��&q*K�,��]`�~{Htjѻ�MA�¸pp��������so���X�FS�,uϟ���˿��E���&�):G�L:� +��s���ŸA�6�oj0�6״;���cu(�q���u0� j�7?$�{FN=Y:��>���ʹ���m0H���,�33�$>��3�Ԟld�om�V@�.��}�yoY�ud,�J�	��ŌwjY�J������2W���
G�Iz4����S��^�d�ԉB���Z_|+b���9#�F�F����{f΅�e�*��������Ϋ�w��Zb�Z�[F��ѕk0mi����	�BT>D���tm ��<��,Zd�י�0��Acѱ�K�K+�6�ͯ
M�ا�v���2u�Մ%�g����l�QM�E���li2R�B�m�W�I������z6Ԯ>M��v[(�&ȥ�0���|����8�s�	'C�M/0�
��(�(敻b���Q�E,<T ���S?���d���1l߀l��?`�+泩��x�V���A.��/۠_�r�U6�w�����O���0h�����X���Y�N�����Rȫ���vG� �aӝ��$�-��`��">��!��'�ҳ̿Z�10�����x^O��A����;vz~I����`�K��(E-ު6-r���\�B��}-M~����c5M�a����y�w#�I��U��G��2'�����XdÔ�n�ԋe�]c��K���\��l��!Ҩ��M���?��g7\���t%�u�9�ڧ�PpG*�XpK��bx���Z�.~9ci[/23p��E��&�2"�Hj�o�p��l�gH�N���kl,I9N�B�z�.��L{gJ����UlI*��t뽇��;�ۣ�a���"F,�s<�A�s���5־�����΍cxWF,�i�d��:l㬻ҀsΜ֩JOv���/��]I�n���I���|��5��b<�w��&t���	���R��Y���~��1�o�h��-y{�ܺH?�پ<̱������dg��H��Pn9*��w�P���c~]�|BS�%굟��G��B^�����#2V���`0�M![ɢ+�v�g�����Lt4J�c��x��ݯ������aТ�&:;�y�LrF�
�vD��9(�7PX2���u�
�ڄYq�9�i�hE���1�`a����v�OrG�a�)7�}FK�βߚ���4^������B��:'Ы�����1�ᬿʾ���]�:]�d2t�ո7#��0����?��!%ꌧL�-v��$G"0�"�H��F)�-h�y��A½i�5�Ӊ׹� Ձl���Ir�{��^��;��^@`4�cRvj��Nx��$��ҨDe}�8�ނV����e��q$�gr��o�,sc'�B�o�yM��R��bF��T19���d_���O� ��T2�߲췐s-�OC!D���`o����+�[3iA1s���3���0_C|H��Y�p��B<ɕ�˿���n�2X@VF8ƲU�0b*3ޖ�c����.x�Ѷ��rs�h)����Y�<�*Y��E|д���826Y$	����~�Z��K�p�E�&A�� cl�Wp*�c�6�-�u��s��w��b��kc��.v}�޵���71��r����S?G�-]gz;���d�M�D�ԑw��`6��M��*���Jh%��A6�)N�|ݯ��ߗl�	&u�.��>�9F���A�*��6g������Z��P�
�i:�T6F#KIc1��]!NZҪhk]��)��Y�y����."x��cF��c�~�a�>1���&��oO
kz`x���`��}J�܂(���!��i}W����AL#rrR�r/hE��18��	mH̼-� )�@�K�O2�DU��Po�4�1.��>�{V[)�L�=��I`i��)�b�ۺĻ���JG�}�̎ٯ�(r�x�PK��ڀVWI��-���h���\�(s�q�@��$����A�Z:[)ȉϩ\:\+�(�b�-�xpEq�^�|4�g���F��m8� �d�>�^��t��b i�$g>���?h�d��[����$q�����1n���B����E��6'�����]�K��|�Q��E,f�إ
�7�C��~���P�)�1jG�)�Ҏ�S�U4�����y�Kv�4��3�b�8�}
e䈍���[L�P3�{o�
-o���ݺD���􁪺ĵ�d{�_�"�2/��n܂��,'�0q7�摄�	�``�(�W`]�S�}�;���Y<n���\G�Z�gkz�oO������n{�Q��ʄC��Y-xi��2g�dZl
�`�����HG���n]��:lG�����.yA�3^5s��#jO �"b� ���߶U��sy�g�iG-*ä.n������b)�c�ewD?�*.�,)]���æ�G�8�Ai-�CA1Q�W8��=5��JvD
o��>���P��&����,�CW��B;t�~X� �E�g/�9�1р�� S����9I Q�O]��o*8O��9y����f~� Oy���L��%����V�и�0�����)Cv"�=��"͔v̿�e��r���\�|��l^I��Ib(�YG8G�ߝ����%&~x<��E��[�����ٵ�*�i^U]�%Zn<�րD�&�@k�9M���b�*��^,D�&�q`/D��Ƈ���`vL����`*2#���щ׫Hk�}�Y���.��!�QmJ�9�2���t��͎���AY�/�4���l�Q.f�Uҝ�&e�=N6��&i~��/���Ux��Z���B�埜0U�W�Vp����7ά1u[?�N����zjcnh�P�tu�ҷ�������8���(�w:�����l)\G)(���C�(	�y��A������fQNm�|Al�����@�s����)C�qiDV���f_��y��y <[��g��F�X=���g�۩`#XgS�s��[j����?7|�;��i�.k`6�*Xn���o���z��">e�w�[t
�9Cٴ!C��2�k��r��u���Հ�|Mn�K�NS�r��jN�1 ��#�v#Pޟ9��/޴L����O��PuNK͞������Q9��Ih�O��%Ϋ�ܾ��4�h2>bb��/a�+��/�hxY�9����+hh
 � 8�P����+���l\Y"OJ�K:��}����5\4-��[�]tT�H`ߜ�����9'���em�7myi��IL�3����`F�Ͻ��'�N� ���^F��`c!�Q��� ��&�W�P��z��2Q�L�6�쏖�ˈȯ��9��9D�P���|����1z��P���TwQ_�/��SaϫM+z�c)�@�b�#��|��Sr���G��Vjl#�xZ����T��z @F�Ǌx��-{	z��hXzZЧ����r�I�5Ft��x��J� �Bǿ�v4��]Bf��w�4�]�W�\�<�]s�v=�̪�5����,^�S�/8��ѥ\U�)3v�����Q��-���:W�@w��)�o�����Z�L�X�f�H��N�*q4�#�x/���f�ȋ��[�I�5-�́n:;{!g=P@a�g�F��G&��f1eh��ϐ`}8��0pdnhŷ��M�Az��D͌�Xp�ͽ[�~e�ei o�o�f�ڃ�^8ZHҘ�J �Q5���2��D���zȉ���	)��tu�V	�i"P�	&*>�`�
�����57U�4�5*��PM��aw$e"?~z0�My�rg�P�|D����7,�$�t��J84�<1>��>a+op�^�AwOp܁��4O�}ژ��G%֍3���Z��(���j�'�e�h`�ɩ��\ma�]s�M{��y/�����z�~������� �(o2m�E1r���gZ��!�HD ��;����=��ݶ�6�C�a�ڧs�t��w�IXu�IO2��)Iiu�@u]D����lN��O���2@�� 0�D_s�"� �l�����A�/N�+�gW@ ��,g� ��|�%�+"�Qq_gH�=\�?�%��~�jz1I�w�B�[�m�]2"���TB�ѯ�p,rG��_��p�n�W�v�dt��5c||B�p�c�b�{[5r��7���M	�� }�U�����=��TߘI��� =A���ܖ�}�l:!N�:��S;X�a9Y�_S06~�'X7��}�`�Cw�.ʦh���tp�X�@4*��`�CE�U[n?�����f/35׍�GMBI�;���>��aj]S<���@R2؏�|0�,�U�]�iC��mS/(z���	�i}=�AZF�kB_ 6�X|%Y�(7�~�����/|����ʠ:��P������pܫ{U�Z]�7�A�J}���)��{�q9�Ӂ9|F&Ǚ
w�s)e*���x�xp�@�Ҙ��q�]�-���1��@�%)�)�4��"�X���d�0g�,z����^����n���n�}<�/��[uW� ����Y����Xq�o։���#�)�����3H^�*Ƚ����d�����\��H�� ��HI`�n�#a#Wt�>'`�\��#�[@�Yf�
�5��:c]��嘛+Ȫ�}��;���@�����R����D6�Q�JJ��k��f�%E�N���[;b�vb���[I�Zm��@������Y�eY}s�u���5Aky0�F���u�yqM�#Z�P�*kP�2=!��-uu}M�v�'j����H��SI��zd�{@�{�*?6����!��^�� �N� �0��O��� v���d�)�Z�?;"�1��g^�������O�L�1^�P� ;��Ӫ��g�2�o�B�fN��P�n���&Wkrz�f��9�g���$�W��D"��|��С��B���ɛ�D-&���T��9�<�t4ޣ����9�Q�v�&㚒*j�В9	����D�������<�I�
=�=��x����*Ysc����N��cAG��IIX(��ǲ<ׁ����3��%�<��$ϕ�#8���q�yD���F�%�R�߻n'�19�m�/}vk=�	�,��OƩ�n8�du/F�f��,��e@-0
�l��0��,���-���:�I�
1�@2`GȮO���5���C#M�s7t$f����+� �y	�Ȃl�н86���[�u|o���չLF�b�H�A����8�V��6�uua�I6҇�҉�N�����b
:
@�q�\��b1��eڇI���[�,��L͗���W��"��L��\��V���%\x3?����HNC�P/7�����H����)�<�����4�O���nR�7�[U����"�F�GD[��y�k�t]���|%�<����s�[^��>��P �(��r���^�®�S�������;01
�@A��)���x�q��Zq�)�p�d&AZzdq.���d�9�n���
g��yۀ�6���M��mxP3��ù`��!$ɑ�z�:��*�C�v���,��n�����&i�;O'�7bc��q�;��'�]���,�͛:77QL��`O�#N*w	�!��7-r3ĉ��-n^��;�_�JJ�ll�.�}_n��k�������t�X��rt1#�m�D�e���B���x�4<GPSrq��n��D���Hg��<��].�=N�&�x��;�-`%�Szc��I����|*�ρ�dX�U���:�@[�1q�1�9�zM�J��*���n^����ơ���r���t�����]"�u�X�TM���6��?x?��+��.���F�i��&�?��k3 �j�����i��\�#�:�pY�֕�aqu��Q��l