-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
dn77vvwx68S659+V4oQq7nY66ewPby93KtciTHnIAgLh3iNUd00w2fivyikrrSdcGkFoZNjGAK6M
73gi5HLbDz7i6sRD/R/hb84XFfZXIbIQdYIzLIUbaoMOj2CImTsppOoZ3wQxfvkckZkHUvZg8YbN
YJeIFsVDy7Ef6WXdL2+1iIxzTxThau4ojoGvSY9yaYVl6EKBXyaj8NhhMMhX0V2HWuDEqsCH0U4/
A+0/V4FH8M+OKEBScd4aw2mEGHZFLuEUMoaK4nAVqWGwEqp3UG1zSZuJo2zYplL6jQ8YXgLz8GMH
w1FrbKTDQwMi4sHz9/1cP1aQmV9NsLDgWKblAw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 10608)
`protect data_block
KlHYM4RcCiH3euOkwwUsRiYY/h1knl8KaaoE7JoZooh/RszA5djfIXmpG7Kd8J1gp3jiV0O7d3be
Ia64dsQZZfuyDqnWAPLQqzYwlsO0P2S5KI0NAsrVhy6QgNx7ZcBJYev4ds3Okx5m5yCUr9upfK7z
Rz33dT22eVi6ffAkAdC8PyrLigMm8SUBtSQbA0SKDDgHk0XLeP8qqyRYjYfxTnSNUh8iav2SIRFH
V67r4oHsnEPA3WZshd4ytiaYPudUd2DX94+4tvehyxaLJaLIP80SbCDpKZKczAQkIAXdr07JFQel
mYBVwDDSPn8f+MlarjVwQfIJllYKwJD2cd9eHu5FOKhrgxuGU4RubJd6jSwfi5Q74C1gImPMrUn1
cQ5aTv9LzAPHmDHFtWJppYo1TPAShd7rHVIy50EYrrB+HUe1VVWr3eep+Zu/maxzzRnicam///ix
haQG/bNGyimO3HDvU81lBCDKbF18dxckZEF45ikaQpvvg7W7FUY5WSyjuyAkJO6yptstIlcgxJkn
33fNchykW+1APV8rckfm4aMyWwePgdovqP8DQSs4lu6cfNZMId1iLjesv5Xs8ipyj9sSSw7GhBd9
cqobt0sutdQVbZ67UTT1mgJBzBu3CNARSMN7AhtqvZEYF28cvefZdZJGfzUUrYuVQE4WmHM+zMlj
57Gk5W7PN0fDUkMZ4x2K18DwmQT+io7567cS10LMUexmSSwB2LOWSoh7ETej7HLLXExKUtZUVPJQ
bhPJ3TvROQbvZ1uaZoF4j5qAx1GoMrRUSkJXfNMECNwKN862oicc0WtwT+QEnk7zyxTMGgy8L7+Q
56d9ufa0BbUB51Qg7Q7gka6eNAQRZqjI5WTjha1yUkW0ktaZ43fpvImZ3CkcxQSLjvshcLlImj4Z
HrfxZQD+FtDp0CvF0N5zaMPfAe3BmkM9OnL+UhssXMsd7jvEyHyA1bILzJ2NwbmUL3owZI7FFnLs
hihg3tyWv/F0emhToTykgr7s2z5pID+DjbKSYYsMLGrdYY/3OTg1ir7YLBQSjY7ghlOgiCBbaqnS
uggFs2ZwfErgaQYC5XHb1TJoIh3XJS0zeLsno/r0Coc4f3fM4bhALEhqv4h8yrnMI4j8MpjHkcXL
qxoWnJokfGLSr4h8WveyhfvKQYFFgQycbx1g84zQeXhvaYnoNtGqS7gU1jb5LYBZHjHTuz4pez6R
EFqdYtIso3y7ZQWvyk92W3vuBityU/MA0g2TMTsbsKjU5MuAsF3fZkmQRvW8ulECd0q+a4BEooLm
UIA6COd8ZmPx02l1qkDW7JrcBdOO/mnSKmo3uYTssuQOBz727+Rp9yMSqx9pxPN8zrfZs98vQV7F
NT7UH3+nkENiVy7oKB1CTMuxqJgM1B1MKZyHuCcCJbRoecuIWJRpbXbGOnd34TXXowjDQ6FTHw/X
Qp7tz+HuqBKCeYmKZn2wQd9ulIBOUuihqYOheEghRWjS7SYLv7uCEdbLX25U8mZBtk3+/2s1nBQW
Sz0LeZ2goe/9r7HwdFXAmtLOZ+B0xisv+0ESk/1sQolw9lEXhSTaHdEFBQNpRYNpPe6a1iSYeL+A
mfxC2nL2j6F4lXjbgYjfvwMaLHGTiFCzodntqQ2Evgru6+lxJCuws9oE2jOXmLO1MPM+6+LK09jk
08AgD7e/E4m6KoWKiXqJS706k4uwj+RPEUJI1MqyQHvqnY38s6oMN6mhfHj60pzMqH2ZLVhI4gyl
00VksnN379UbfhuO5CpP/0R8mt0IAoxBqYKAkvYKZ1MbY12cH03le4ioCffoGfvx86KeSsAJGBen
m42LHxg/tPdIuEt/7IayH8mVIDchBdAqzsk4ZK7TFpFQS44M43DSzqlKdaCP4xjo0iT/3gmbX7zz
wj6nVBJFW7TGqxisC0iwHDm/E8y1J+s8275ddftQ+I0l4aaY2Wu4+2nd1ZuKzifCblj4LmKXk8Nd
XUOz0GehUetlychsrLUHtJAqCEMghc9ltGOr6WwuwrCi0cikSOCAnJt7iepzqdrWAW5FCMApihGu
Dz5SLimVdXZUaZ9ckrYMk+2dOaVSQWbpnibY1vAZ0FItgcQaeeVZSrM2gVj5vtzTcZHwHjHCmZAi
nxkulVgfjt9kuvhhDgnD55aYcFrBkd/e5VC+Bs5pIgDMbcyePcjK+RWtESXD0tR/bbsUT3MyF7RK
RvMAXHeyOwamp6hwLRbND4Q0/nECpOPI7RpYxzYjKcHSR5waU4bRnxyn0dz402hHufRkpw5ZrLEf
teYXhboc/MbGLIwU/EqZvgArWdbSFG5klv92pg9GIGWh7Gk6p8vCwgTgAirnI57y9XpF6o88gO8E
lM/2wXhCYyKeKhWZZNmO4wQeMGFpQHCUOXSumkPAX9KBZyVQV+saRPVTfd01Z2QMUSgL/mKk1JoF
uvvjxI/FQyU45E8RYcLS/xVbJf/sVfoX0g3ddSSk13Po0bWkwom14TTb9LpdrZaJpBhWCYd+eHo3
SyOdp8EnhU2BzN4iiPZc01G9qBcb1fi3eodHInqJg/KhwK7cpH50l/uEh6lAGDnICYXuhlTxEMS5
KbeW6rHhnDx5SxsYu5e6TpOBRfQtM2k+qiOCs+/uov18KYzt/FEWa005tx8/O6zus4WZ5MvPyMk7
FHBb1oVj8UHc72YbqSTf6qL8965f3SZxYDjjGX2VTfeTWRw2cT8zzK9ENP1D8ctmIRlnzG5jyFi+
mAWXlmlfcF+M26tmAXQxbhEXq3Ddx9yZJunAPUrG6ZJVp/IJE2ie57DA3Z7Ld/iXa9JJjXw0Z6+T
rWHIpgEMjjZf8Ln4uzWJ0StC/MEIJQATcptS08s2It1xi8dljvx6g/9QwJHeySXzr/AYcjmb/qve
fq49wOuu5q+uoLf3yhWnzY75SNlRvD/gO2U7XpShDcXhVxG/TE2He7JV2TsnGLVBcGC1Hk4YfsJQ
gOTmnFvrBvgodzLC9fhWFSDyZ1w+oMMAbUQ4NXPpvVwUJK/56dYE3cTnIJ0Djzw1rvMZVcbNCJmN
QIEuz3ioS5WqWp5T6ESSCZJP/kYTt4M7uv1ebLhNlTWA7U3tF8iO1fctQLkiTSYCz7RytGOegDb7
XLOVQz4sCEu7Q82/uI9q6gbDBjdx6jMSFvcsST8POUcUp8wNK8CNVNHmF6MRBufHIeowcTsLxZr3
EPNYlBut0KqsSDiwqdecVatVAZQ7OeSWAzPWq6VdUsotCCgDgJ8i12IsaWyqMvaj7ECi8rHZwmTE
gP4f+YVB/bQRIX3Y20Hm0h20vg7+GuG0zFmOHqMqUJLQmYWKzSm7SwuFrbj99hA5INkwMHP4a0i1
eBC/pxXKBHuAmWl3U/5rq1x0Vq5AgkXlXEtIs+JcOgrhiRsE2dHJyc6s2Zv7bu9fbImLdrq5b8Wt
canIcJqig/ekxKf+Zou3GQzlKJlXDPJ7PdskcOpbPqPl7Nq4ohqNkoj2Uim5iuzcgWAbvv0zwYNt
laeqWQkO1juGAaOUB4Ec/VEBGsBFaeBg8Pi1e1XAEbXXJXkVHv2JHMfbDFJdA2JGVLVIPNy8Tc0I
IIsfHkab/rTY+YQmr34PQGVvc/hsjnW2gBQi2Ng8eFA2fYTtwwJoh8U1DNmrljLNvu8tRwanya2O
l3iP4vVEhc0Gkr5Lk9T1NSWYrP/ipihW9iPQUkqqo5h/TVSS8gd8SWAhupWSyzaSR2kBoSA3QxE3
keHT/XGFNOJUntsM5GrQ01POI/27OMxVtAxwr7wXuiRDUf0sSSVA0JscHJCsABe/bNepD1M8Xcn5
DtZExLHuCPrAppWX53/S1m9smJB/IPPzX1G2nfgEfc5xJKS7jIfVd4+VyrvLRgOB3hSxr/VisEi0
pO9qlxjsX4p07aBPUxKZVFA5QLpjVJlTKIG20kbG5lcCJCZJ+Y7C633HdQaEmbM+LtBUCEuAeZiv
5uTBE9tKMoC9lJrx/UGEgRpxQZW40SM+rQzXkOEC67yfBgYkLupMgmTcPEpeIWnqjJNRLGMBZ2Hw
m7sPtbN6oSSOJDNz2Ambx+0hpbp21W9OfMJNNjsGqNG2tPdnydjWogUlBYQSHILvVDXbIcNkqU8F
EImtBn9GqG+UcJT4FBSo13WqVbYptQkblrx8szMg0l9kA+RXWZ+HcgvrMZC+pNAaoLfuC2HlN8T8
T6AXAvl9+LGge7GgPMhQ7h10cxy+kB/P1AztyVYm75E4YYMqbAzLpVzjSSF1ORRxdgZJTq13OPSF
t4RRS5mqKsTrG3Wr3VsOV16Lg5qotWjA0rNDHcWOkoGLTHlrQJv9JZFZ1FaDWSBhd3qmFCmkuwSA
IIDwbHEZYTu1FiKQTRgxsmvMPXoy5hri2uJqpCBCasb5P7oO9NoyzOvuoB5/R4HYUTRL8KZ7ZZjP
m0leFn8riYTvJUtydEdlLfMAxtAzGB3fYOFEy7YoQKvBK2HW5Pz9SRp9VEe1UgcnGWTqi8DGR6gi
2iYTEe8jo8nGMxxMJvLf3BTJBggwaeRSJ98Beq8ZcNz2AMYx8dPd7yxAiKlLc6bh/MstskvrYLrg
ZayetFUcTjv94Tc5tTDp2EsNcTZFOyat1llvj2/COBJAeubmSp2UrPK8SSj0QGlPzRyZM98y0ogq
kHNRi7lRWqVkHzw0GvZiHbPHo+I101tLACjyC3lDlelj+yKHa3ZY70LTXuM+7+UTP9HwrB6DQ8vV
xAf3JlKmx6IvWmF4M3dnvNRWqTbQC68ONoCE7fm+X75mUTCn3CnY8sUX4EA4cBPIq5iIZjKTqh1h
QytV4WmDRnkESCPRrxwz+Df5nC9djnP9Z1RPvqGIuMBTtusQnIjw2Mx1s+qmst1aTwJ8sef/aCLo
9QL9ve9bllcLAPTaVrbuQFWl/8mQ64ZXELO/pMMBVtBwsjeviPQX49XHzRg8eKiIVtXLXoeBZqKN
vd4HVTrbYQmlQaWNdCKocvJbOT8hyoxq14aL974aVqhQr/XeR/yk2fbXiZDHv2uN6xHbznKrvbQH
VD52tuQg0RywebjHq4SEYVcULh1KpSACsISlHcSKH90z/TI9ByqaT5+4eC2kAyziV9OYPRwQ8Ly9
zsg6jt2WaZhEraNyTK1wRAw7438FPEqZiwLdksoCcwsngNuYVXjb908WvZWCmv1SuXtn7yxi82Ii
iek8VTOSmCh5a/bqFlI/aG7qtYOvYKuv7PGWHWpKXywx02MPGJR1sKo0rDwWVYrdZILNTH+1i5cU
o66GA4kS+vzXoRJt2jzVCh1nis14JrqKas1kys3pzHDNU090rzer0Oc3MTDzS7zuEBU3zEfmhRrq
urvv1ylqECbdgw2xInRdS14/Z+uhuAhSMsPSyuWLfrVPJ/eG9lfrnAiAZljs2s1QpAM2rd+Ilp9c
Ld7CjbIKwbBKtKlJmqT4N/Nb3YgJQObRGFhkSWERdXlVTvC25Q3mh6vKytoRchuudKvv+fd+GSgC
kwGMwUD3X44YNOF2ymT2GWvSrY8yfJODONyqu4EUZymCp7NSoxSLZAnjQop9yOKv2aYl8lF7PUbQ
aJWH1veaY/rqrAiV/brOIIT2PTJ493cilmN+Q1E/m8/X5NFwovxDBKymunXKkdbqbFUanhM7gJEX
aZJh6YFD7uAMZ/gI9Jv+YU4uZ/xDAxTJ015/g8a29adp6TiV/0w4m3f9Jm8jE/ODiPi1tZiCbyyE
ixdeqHwHAaTEcXFOK7R94C8Y9aKGy86d3KPCaRYD72xVg1HdRs2Zo6d1yG0yzkMe+rRrLd4Sgu7y
pCfL5qA3q27UmhI3//HDmpqxFjRU6S5cFxRrt2U1oA115qM9jymvS0YurN2Db+xGwgwM8l5ge1z0
W2IgyUIN0yt4eL7iJFOhBtvwNiZa02SI0Vfq+Tc5EoOqRbhgjrfOoIfEHR2GMu2ZKWMe6G8BxGtD
bhyLXDqOwmH3wYDFc5XVqOApq6vuA+Nd47nkMWb3Mo0efjlB1QRjephy7oadIGmy2urKlb6fSB0L
XMZ0F6azagUtT3FkDCrVlxCvpBg4q5ZDZcw3G2yz3UzA/bk5vOwDplxYMZgi2VagQwbGgzwYJ6CR
u2ghEzo2ySytBjAK7oBCdUOAArti8XSeBC3tSd2CoB9Oot2mACtJx9jGUc06eng/Te+/7ifj7U+p
JAiaPciuHo4ipOxVbGHCaqkwXcCvIxM9xedDCvluGpn7/pSEQtla6pZW/qhtWLf13eNvOGSnUAsp
Q9bdwKOkGysO7ooqTE+GQdPiM0KMIH//qkjCCeTVCSGgV/pgHyDhgyytr2GgNXSL9XWqwGLkaHqC
NdG4Ye69y7kwVOyRbb6XH+49ogGxo8Hs7K14Uz74EBRMWB6dRhsF5+kx0l8Jh3+24NGw3GRXuDoy
2PY6lLFQdVhzw67R6bRLAtvggw0P5whWaV2ZBPyPiIGKdQclwY55/4Kw9xlfTm9lHvk0FHyp8/Nr
NIhizPQ+bNSF4QsNPkBot8r1vQIGaZxzQU/pJxpTEFfc40BxUzV76J1YeLsr5ciZleiwTF+H4TfP
VyrCiM1D0TLII9SrVJpq4cd/61Mx8TcmesYey/ianKtXSZpl4JAMsqIkdCYAGcYzeryVzZxxqiWN
mqzSAvI0kzpEtySQc7aFNq7Hmey6ptk3cko1lv0LixSmYpVyyyzdZJr2X3I7E/MFlvUasXiKJJ4+
VAnO0I+jQo9BtFem9hoPfeyIfeCbG+UrIxYbVtS9wICdMsOPtu4VXQkXw6iEksyNhJwy0Lh1seWW
HC1AG6DkZFiiDKCwrZLNWpPVdkd5S2bvLmLkKj+iA99YBZ5+7tfecmbukG3/Fhb4jOKatcLI664e
iXeSUbuti9M6GCNBAlMPRhvP2ApkdbarW18n1HaeiAT9W26B4eIvPz8zYKn5OE62+/bGkZXNRoGS
xVkn28aadNK+jlatTK3jXd3yAavS93al8F00xZF0EjxRV9Cfx0p1c3QaJeCkqsPiVbUs5zZjg0YS
TXeQMaT0drYN1yJFdOOfrXpGho48e/PPVPaJdpkTgnETrblgXQCtmBH2TXTeU5avKsQTw5QSask5
7cFm0BEAEscOUtKejvjiIlfIiP/m7YXkiN0VD7dqsy6nAH6W+2xGaDVDiV70w/5FsMxzkMJR3JyE
rMLUCQSkI6KzDFT3W0yWzQlxRAtpD9yUKt1K3bAmaKkY5JmrVMFN0aDwNR4AN5b+bpxdiHgkDajn
FTt/nzAjGjGbo0pceGJLK0ZUQeyEqHi3tNEQMhTveMsbD40MVqsAERbizNmocxjgPewliFe57O6V
kpIXvDvxa0WuPrwH+cXaBBi8KoSezeVNneDs55bD1nGI+TWU+oGsB71qBckkE+v7OakYyM/+IdJp
OJdGfrNh0O848U/vhD1JwaWXiECZFC3AfjSA8hy5fMt46aIGl7m0wK8JNwI5kDekIlTBiyK573SO
p/R0vJwqjMS8nv4zHGqqdi919XK5nDADPh90vdU+df0J+T6Yaq1RqNAPKHktxiai07spEuUTdyc0
K+xBgGaAbPy28sxnKSS/7dXkmFG7GfcRR18fjwRck/c7rjksT8IwU+sYD94i9Dpep7/mB6hXGZ2K
d769QLzEO1XOsO5nEHRnBTRo6lWzqItJHTBVwcQlpjQSbG08OxbYyeoIGLamm2EXgUlQRhMZ43uP
59JJaXoTKD6BygGWMSq84gC17aGrcKU4JJZDznD/tdb0oB/feTZtOPC6wOYv35J5Apgm1fxbx0lr
o+514lAyX2k6AUg1P4LJl4C7m2spSuO2RpU6q7NpOVMTnI1lWNzEKHw02HIaQlU/KugZ5rbBSU/0
S4ue+LVxuVefjSERyaJMzq1sKvVm1FVLcicoWUhhZNLNmmDDdgkjXoOFkfQyaD5WvqcgfyaZH7xE
6BGhwpD3aIqzP1WUohZbial1YiTOiDFchx/SSjLawrSNzd+Z1wOTpxAzjr81Yqwp8elLnNYK4mAf
tz9JQiFOdoUj3oW0kpKgouqPxQk3wHLMLThuLiSCj+JcshvRgyOQcDhmUbWqn3alJoCvQ7RaJpBI
Nz35FinbXOl4XPU7cFN2557UW3OgLrD3Ob78S2oHpNpYf5lkAoK/xe/QCOUHgi4kXTb0W0X+Z9Q9
+FrUIZGDKfAF5eLvhBgYX02RRbmsNxr5JzcJnC5EK6v+wmPbVGCQINll4fq8EMod18gzZoRxXaCI
q/kePlEn9fH09iPXqhAweGfHPrt5cD7AHxyhfDTGMX7RW85833T7P05FO/Fv012k5nJktOfBxyUG
eiJOzrnVA7j6qtC3Dw6dHP+adVSc2xxsgS0oAR5MMYpEBVk/kbXFQLuAgthOxaA7I5bhlXxyi4Dn
5V4mb9BfeyhBZr3Xp0WJbig+27NrC7DX+724+cFSljKih0Xe9w7HlMIFV1Aa1PfJ+bdNjzAWJd3w
7huqHkgqpbtFlh83nu39pHsYosvlRdxg36F4tDQXNfCS4Ea39qV20lOqedNq+wmUVnLn9UfvWJSX
UjLz3xIJxCNTQWMtDeP5rN6bspVEUQwMEvtgpv+Mb/bZLNwTwbgAK89By/oefyfftH40vqM02uXA
mFQjMNfmmgfDFn4blUtLAtpzJSSS8Pa99rXGwMEDlrWinQ0X736/ttFFs3HMGCzFpROdBwVRpVIf
aoEZfiyULcKduhHymEwZqz75z3grj7DDqP6pN26EF0iZ0csaAAZct5B/5pA3+LoDpqCDfwveSwuQ
9i6K0h+HAszMZSWo6wyfyK0fugxL+dYScbbN+vIfKQRjpyHhgb/KFhmwErGB9EiHXFiquWhKHk1S
W3/hgOZ/IjcPodKJjGSYNHiENL64crBjb2OSrbb//AqkNGmisnsPka3VWC/34y090NaDy6/nMM8L
WqnRPxrPiGqHBOlzbyfq6eF8jKrJNB9OXCxTUCz4DTIq9qMa74ZIq8REzpyJ7oLFWGG5b938p8VP
hkts4xBA01mCgu68MXFxVtTWQnztm6Jj4v+i7Hna5oUnjVD8+xz7ej96jXzS2FLT16KMNd17QBa9
BnuG5hEwtWj6ExGVlapcm4UN2tbrYkuLKGxwXL1z11B19CE5oPCoLze5XvRbbYbwh5OFPUcFzwe/
HCgz7Y75gDF3EWQD7iMMMEdcXiSgcfOKY6KgbeJ/zopPQo9C8RuZHt+eAE9qxtnxLq9sYnRSoLxN
4SCiRfJJ5IbOGB9kpXj/CgRZQBX/nJ2ce5RlSHOOxGH0nPcdAa0IaiS6iMKTmro0aqQRf8F6KE42
AtfToSdSFV9co19QbcMaILWOST6lsw8diYIYpPzVibQGlONzyjxIxF5AUZuGFgtP91WfjQaphIL+
8JpRJcR+u+8HYVYW5omDZC58qTw2kqKptojDfCcNl/gScuyOdS/exys2FfCSleCg+VrGe66qt9it
0qVJ0Hy6ycUD3NV0om/mjkrm+hoxL21kQIToe4ZBsZ2zz8PWDe8ewfbEpY6/JUIa8K8r+dfRdEhp
wi82afhkPyrkdt41Y7/PQ24MwnDHAl88n6O7SpcmpBiV69PbtNxIzYSMKK6Nydm7f/hxYoGG3hy3
9ZMPf7/tEw50Ji8uXd46RgiOiQs+Rh8KzmBWn9Y7+++pqmmHryFhIpG3Ju9wTQwDUuuNq7sXC33G
AvLhOQszQ3NLK7ffIH304yPZTB4b5N8EKZAXhnS7ilIL1LTtCJHBSxbAWzCpE3/9HRCS4yVPZ4KM
IhxmitIxh5X3/DePtVra2WV8KMmv15cTEh8N8OkCQ4xnR7PNf2d6WqxmRcZaUI/wnhRs3TVejBri
utdjasEG58TRkJ93oxdMM5kDJVqxbUhH/+6Ns7jgX9iT+dTT4T5k6MCBzOIjuaT1FKVebNHs9AKK
YAXDAiztVrDFhqR8WviU6nSkiCrH9tIxz9DsIwZSPWyfLvJCeG0XXoK3Ei8YrqT1KANlBhdJuVrx
OpLHhB5BpG1zs/zeXgYfEUacAYW2DQuL3gYWtNmtXw3t6xOpxHsPdwEZKZbDZ5I/DdbViQK80L1L
lEUIe/1g9wDNDyFcU/Nh+XqR4XGX1/KhPYYe3nIXlmLKz62M7t+DFocJsE/uk/Zcz7Za6UPGrbuu
tKbRuzc3C6Gz88MGG28Ynh0XZCItZUqrJtX/q2i4dxp+YVpp0oRM9m8HHB/qZzsDPFghKZ6LsOpE
kUd3qzBhG5cDyS7aoJZ4kUg3pGKGAHSEDSGC5X4nY3hMMyJN9HEehS6Af7LPzhLAwHJgDuZ6bs55
/7v6X3sEYXhrC9NzYbz9RjZyHWmiyeoQHPI0AQLTQPUjOZlNNibRp++pwK5m/xUd2Qj4q7+ImEqP
1T1lgzpL+5DBQpL9aNi6loOdN9mVrzFG9oQb6IkxGQQkuFEm5EmoJiwiOgYTkvFbBGNipvmUu3xF
CKLy1mKNjDEuhjsOM6F8sleuGQZ0NbpbCdLlxkTNYv0c//TzGmq7yLwHD2t3LfcCT6n1Rle6oVCw
ri8FTcaYI7YVss3mhn9ObRJcnlG56lDj+ytujBVufNd+nu55JjadUwOSij5i/+pq/EOq60ajx2Ql
07GVE8l7Nor1pK/nENa1fFfmURwkU1Dyx4jsQx5/aDsdQJv0Eu+IHS6INqf3cTy8OJdq4ZdZFBij
wbNEcHZeadVsJYuspGQ52DLOopFLB5gz6vIFRuN47r6L42HyOxoQaELqe+OQcQVjVrHl4F1jWX/Q
VIXb8LksN/SRb3be79WhCVXNgd2U6eNDyykqIMEup1/gFcaZmidDRMWM05zMEF/6M5zEYKJl27BB
cUHuQfphHVEsDONLWF/oe5UhDvkGsyZcweEiFW6G+A5oTDtOf3yol6VKQwPVTCjJT4sksV9VPY1J
rR667twtD/xfak9NIuUG0n8OcQBR0Uhrruwi12JZFlWUuUH2lyFj6gzH0TYc2SY9/IHkpQfeshT8
Gc+/n/p4L1ofc+p314fVv7o7k2DpZcznEMSkx7/6at0apm8bX7UWIWn2kKzuvInFHXyA7rbh7Myz
CCTEceSd+9bpARUuAIPttlnUCCMT/O7yDAl2YmLrIhoAE+4sEzFD1NCWG6E3kBOVd5pAXratLmxa
GDldP0aB8RnUDnSarqnmlOpb2c0oqHAuogZekGSWs/TF8ie2YMrmwX8novnXasboDwtoZeL+k02a
TlrB9fZCr6WpHrL2mNQw7XDDJz1pV8inTAq5APSs5+5q429CFE3tMrIAIFqdUi5wph3D3hi9dh2+
/+Pm+L2cukrxv5lZITlGlRte5h9GcVxndZ2jhityLhZCH0wX/ZkMcW0sToP4698oLgLOttSR0ds0
ycu5hdVvgsOUDBT1kghzDILb9pzWY8hG7NE0nnDSNRnYekE55hZ//ASexxQYBWgCWiIXPoInLroT
hG9luePR52rdN2iyZKvPd7II4E+BMzzcdn2BKhydjFwB9nOXw60evctuPkHfOMRAIXoQcByvtsXO
Hy4XhDL8kaKeRntk18GhAfsQKl05dTyqqWVEyL0PK+l68YMc350F4zB0eU36zn3sD+NthbXTVtNu
X1yDQAkmPjth/07QdKGrJyVkfTBQL+EKWsmx71/MF2GuyERnhBADOn4/yfGpO+ufLPczTCwrpGLA
3n4R0+54qbkFZTGYt9j4ujpg+TXrEcDr/ZulEcNqHnpw6FM1LQpvepFAtDaVwfBiUzRlYFOt0hg1
uT1fnbszDwyKT25PLBcJLCuAXTSnlHlqMegVd/SXq053Rax70GTChea9cJP+rP+mGlbxXsKHy0z0
e/a7sEU6gv4PYvQTuit5T+7olsBeOEVwcznJL5z1vHfaVJkbnIjBwY7IMOruaNY0TgKYxzmWM4MP
DKDH4Yh2BJnEbo0zbqYHeeM4X5/rKHKOsFcbdXqFL4qg74xRrZ5PLEbwQ7DWBAXWgZEpAhPUmfLT
ONRjhT5c7rD8gh5e34QXKKPxI6mP+PCUjAqjlhD3yMgjUGR3BnxL1nvbLRXh01bqaQOJlFKoSTpw
hEZIC6H8k6I7eVMhrERr3gsoPfaj7rdQ/9tK7TfoGmJlhQmjDHx5dLUfbYZgBwMXJNhPpvtIcFnS
igeNRUiLqqShMVGoNfHcmb9M9GZaeqotGETysxllCF1mW700RijMfoYffQ+9KysJTDhuLua3w2tq
fkMuremdKKn+m7p8Ms06czMCJiri5xr4rxpKj0Cto7XLupgAvgpA9PD/CUhCx1K5GOi+hxjg5+B3
9GYmqPDJvf35GIEfUhCSKyEER/M3zuznPaw8GCQFA27O988rybY2J7cyiMKDH8HdtP3JmV8Jdwrr
47dVuHrwAhP9q4OEPLBYeYxMhwlcLlYVME7BI6dsU3HFWcsjP/DJ5L+g4oBnAiwzqcerwDyL5v8h
HgZcSPdSxfzd5nRulj2zhlEDlw7VeIVGn97nPskfm5aAGFs/8UzALtmUJqLgQjc6NeU/qzY/VgNq
b5h8u/V2PEr2eq+zt980/06Y2odhHbWgk3IPx6zqRDj9HYclP60FH+9c3Fs5bTqGKynXg880ojmf
krOJGgbn9tcnS/uX/DlhrbMeVl2aYpxUTtSp182fdC9FsuzVncDRMAEEGFP5idJhwkr7zeSufh5v
9iFHhFXpUYEgClznPXNA4E0pwT9oJCYHuRB5UcmOYQRNCr+s9QPXTIc1eZ3dTNmykz0AAs/tI9Oz
0cDuNmdaYG24lSyazlYyh6P/RlhiuSz6VCiE5+fe/jWiUs4sUYIkiA5GGE5l0H+6a11XA6iN8aEm
GFBmYBCa6s/8ikF+D4G+/bntGDIOUf9lZ0aGcn4IoPH6AdLQptSFeSeqF8ViOZ5WcPOUPDe2N3cj
XDl8abUjyXh9NBgM6NWSgeoRNlAnJJEpzF17JWnSo8DkXjdpLSGdXbKZwmVA57VFIK96j4OLFVmO
dwviRKoLPKswWur02PXZNcjnW/dSdT2/kPDbwAYKoDJAT/d88RtaDXtPudEDf4m9UfM8eFVtq9XC
vKggBbL9eq3E6uY/w4ZY4hf+IF9jJoh5q0Y+bPgfmnEFrG5Ce/nS8ary/m2FRe5d0YpUvMJUB1Xg
dBcSBX0UxAglWhHEbudBgHy2AbTjkeKhp/uqQgVBKCN9jrAb5iMhjVbAKSQttYdGyDGmSvkZyLh1
3PFTegYR7WS0Wvd+OxTcMfjTrkYGDTUT3GY/G2lpik0ko6IhwSwtQJFhzRoDRGtRVhgumrGWrCUc
+jNp0Du3SshXTpDmnT1MmthSn0ZvrsD7X+JNzLzK6Sef0CC8XOTiDKM9jHsIYc7MzVw/ToDcCa7g
eFlhMfLPckmluQGSJwRIC8kZUuwInJieE5sJsOSwVRlF4Jfh6TpPajT09Uc/puTxNeDtAtIuAW9U
zguF4ok1Z9S3eAGuzyUTjwiK2Cxhwzf0NIjDoMEvUYrKINuJ48HdGjFjOhQlPCOF6/yA/xevn99H
ax7hn18rhS+RdV+HtOGr7I46C8iIFvZx3Wwd55Z4uXfyALnswds1mSn7BWrg58/ABztV1GtEwW0L
Li+RTZZJuh6/v+1Y4tFCty9OKUceFxaQe8MbE74RrjtiJP1H0ZTfGtaJoAQhQnkVCwFW7EYounRs
7vXjdj7nW5/l3Hk51s6l6xek9JWKKrCx0lCJwlZINjh1MgLBKQ8yWzxfYMd9ORriUjDlH5u0nbci
H9CVk8JaFrqXxKef5KJDa7x5ZkRbXHFSl2Qc57sCRVDG3QlUwvyGrw8sTdqW4T0iJtvQ1oj79OMe
x25N7AXpTH9VeFouYtggZ8g/Z+HLax8xUSV7TVPId9Eq3XAByby9ngzeknDaqdZjy4xqUrrJW/A/
47W7Vog2e+SOtFkI9A80Fgr+t5QFj0+Y+0A0q7ty3GcLUfF7fHF0YWjkBN/XZUtMqt9qetQILqPk
MOF1g6KHVw7mgSQ7ldqG955oTowOEggTdOQTL0QEXBFqauk8obbIIHqmTmA8D4G2vEORjorP07Mx
+QGzklh0LfU8WwA3OziX11j3VYgerTphyNUdPnCdFfPxwtR6zbGF0dyEUkVYFEtQzBD2nKjIhHqb
rTo+U8tcAAO3g/B7HAVWDcVPrGIH/iLI/rumoXuBPpK65ko1Yd1xidWDbPzcJVJHJmXGF1aTVM90
3lwGNVib
`protect end_protected
