��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$Rx�y�<��wA�*;�x���@�̦�W�X�fa�M-$u����n~�%���P�$��W��kYَ���P7�?UMfT��q�6�U��k�>����~�\N�(�����X�e���/6U|)�X2pF�]$h���d.���9E��WG��L�X"]�Ad����ľS���8od����e�GT?y	7�������ݵ�^��R�q^]�鍦�����s�ae���h��L��P_���ާ��YЭF���'\��68�b�[����w8�[X��V�F�0͘3����q諵�uW� �h�u\V�?@��_6G�_�*�G���B�絉�f������[�G��U&�����~�F��AׯK1�`c��[<��FY���4I� �#�G��x[X�=�Q1��`��R>(�w����R�O�?����7�,(�H\�#h(W�EH=�������yq��Ѿ��aF����:�U~m<|��.��0=�P/���4ǆ���T(���M�������4dB�PAAڦ��RG�-9tP#����f���2�<�ļ{��4p��hy1&�OR��:���9��s��g��{nH}�I}���:����~��a������ %;Ҩ��9�;�ؑ|����g���s�/�}��q��AbC(�u8�y'������B�zO��$6��X�xt��o���{�-Y:�%����wU�^��W	�
*TAΤ=���o���;
q�s�	��8�Cj_!m��(%*�W@�ؑ��qH�F@m4@������{i��Mk���1�V�:yV�����Bx�R���~��|�M�O)}�ݶ�ϭ�L+�Ɖ�n?�r�M�6���� ���I�v,��1EY�7#[0�b`u��\������A�q$|���i)�H6¤�p N�,�a|6��W�{&$����4�-Z%���o��&���n�6�vfL�����<��G&QB���$������W�L��aߦ?4�\tk�o�?�Oz�|�Kn���{�T��h�$.d`�S H�v���&-�P��
�X�P�P�Ӂ��Rg�?��dM0�b�q��#B�]��Z��hډ��-��/�7�p�+� ���#Q�B`�P������I�l.�<�9��Խ�g��{�=6��9�6#���6Yl�<��J�*'�B&k���9L6����3����n8��큛��X_?s&gc�')�;m�>;����I��Ο�L�����-����/ ܝsn7��6�5�rT��̚Q3�]_�$qەĝ�k-���� ��Ǟ��Cqq����l&�z�J), w�L�m2%1a��ѻ,^���hdI�dv�_����EZ���l�Ğ ��\�ڴ�|���w}uN�M�}�xM���mF�[�|x�K�*{�Y��q�e�\�v�r�;^��:c���ZW��"���N/�����td�#����Wp�����]�2�4��~/,���=��yD��;�K�V�R=}�@-�C�&&�ە�
�'��
�v�"ި���^5lm���<O0R,����ܭx����h0#24Ώ:�D�o��Ԛ��6Dqe\|gG����m^m��☋|�BV�3���@л۫ �Li����ye؏��ZN�Av�QW8<��8O��cp�KV+PL�������˪������hJgM��Ο�fѶ�l<Cn:�^ܭ_�����b|�Ő���O�/��d���E������}� �j��V���
��qh�I �pƹƞ�2��n�L���s31}̩���O����1�2�	&��ݽ�Z��3���H��C��{3����Vͱp�slbbv�T\7��j�>K�sJ0�ђ�E"��5��լ�����S�O#iѠ�\��R'bٱ���B���$���~z8ۆ|��vHqVb�|�,L�����A唱K���$F�i�w< �4
eD+��o���q����xjP�^HdI��(�����1��� ��]˾��N�d���7D�Һ1:����pP�$�΢Պ ������_}M�j��׏�a~���h��#��s`�@yD�/P����+�YءC{�#���Gv�erP��gynh�@5��B�8�^�^#hZ-���(4��{���@���(�'��j�Wx}��ԚXB�����ر�z�"SF;⩫�]hZ@7�(����G�3P9����su��=V$�rN�Ñ}�9/E������u��݁�Ɓ���.�K���$=sx�iO�\U�jJ���Nh2�:�y���}M�Ai��WM�?ox'��*��jn�:$�3�Ĉޟ����2T���vE��Ƙt�Ų���Rb���r!>$}e�}-y��Mő���]��?�4�y?@`�%�ѮhFx�g�E��!^��GrѢP��q�ν��&�W4���a����Ih�	Y����m����끀�)�V�%tǮ�BpJ4��">��]ڻr�����).�(LگHU�H'� �O��x����U�S���!T�4׈}��6c�
��Jx�*�{���@� 9#uc�_V�_�&����U�_Q0y�ƒ�V>��\�a<l���� ;�B�!Kx����t�YAK�e�h�_��}%�`�� A��1�/7��6�S���]��ll7�ZE�aTG��N>�?�@Y��6�)���v��;��3����寓��
o%͉c���I�/r�$�*�s���n��&�4�;�if��&!ħ���"&�T�e-LbH�ϟVav&;x(����-����_y�@�+b#IB�B�����R`WH�#��?,8G 诱Uo6��23��#��?��w�l��R��Z�����h�ra����DI��*�i("њ���Ş�gJX�&'l��Bַ��/3{�]��I�O�<Ή�)���o#��(�J-FM|��X�|�*��	�ʢ�_@<�HѼ���ݝʖ+8E��/8\��l�:�A���2�?�K�C"�Ty<TTo�i�d<��>4��UＢ��N����	��b}>P���Yu����ض/���(�QN�
R��S��NK]�j��|y��0�4M�����'����sI��-B�뛹�xM�Ҟ�&���ǲ>�"U�yZ?�N��^���K���(u�s�D̓o�����#&Uz��F��3bB��C��������5��Z$	��d.�&`����3!� �^��ԡgL-�Z<�|�[8Ĺv�aO�a$4�6dd�\��.y������s�`k~�����3�E�<qI��^�:uSM��6�x-���M���ǹGB����+�����C�wɻZ	�0I��Η9:6�*(Ͼ7���X�4��"���[����(� T��JZ�Ly�-�u�4Șd� ���ʵ��e�eb�Fa#���F�l}9�,Wh�;�������L�gT�=�J��0��@veՒ��
R����q��{v27��=$�j��т��yu#XۚOR�o(Z+�0�I���\�R�vVH/y�
��|���O���
m�X>���
)^b}��*!8a�83�����)������1ez;z�8��j�0�)���(g��%�
+v)��gX��Y4q`3�U�'��e|�NT��,诋*�����n������
�^����E���,$�/ ��0�A��HdȆ��&�����g���%qu-�$D�C�lCF:B���n��T�'<o֒?��E���&���Ù�X,��tr���yO����֚P}���U^I!�Ԏ� Qv���
L�����h��wT}��[���͏��Y�x[%%i���'���q�������JE�)8S�O=�n��؂å�;fM�3w�U��q�����:�14�8��n7-m`��.xN��5:���C�1�*��~3�(��J�ɹE�k�!Tw�IC������R��#��y S ��<��m�`Δ t0}���	�cA�L+.mjYP� ��^=$��ٺBr��Fb+ɝ�yu���4 �!i�iao��q/�Y�`!3�����b0�=��T��~\����W�uO�.2�2 �/� 	9�z��Ԯ��H��/�\]T�S�4���e�08X� �f��>�u� �ɐ�����C3��g�'N,�'`v��'��t
rj޶������z�p_ߢ7���i�$��e'c�v7|��~h��,�)�-*ǥ>XЅ/����l!"��ɣv��/���W}1"pc$�$��B��	��0vtg7��)RM���4Z�v���@��m\��T�A�ϐ&��P��}t��%1j�>��x�?_�d1>Zs��(z'�\p�������ߋ�>|����7>���l���Yt<�>m�0�!��}��G�O�[�Y���A10�-����~e����m|Mqp�5Vl����������E��O��!9`���㒜 �oPD[��R�D���	��s�ޚ�E�L���Di�y�TR�
���� z6F��p����
�d�K�MM��y���7�ݺ%�/N7&`M�M����3��~�z�=騵����Y�i�t���ބ}���r�����m4Oe��էlR��T�*ђ�DY6*�ւo�A�x�kD��%ל�`�G�9��;ˮ�xY����f�VS�-N�y ��F��.�"�Z{� ���k���P%��
NR�3"*�w RCRV8�%4Ԅ�5����t����<�j�c6���d+��D��ת5�yv�]��!�iXx.�'X�=��ԇ,C��4��U=�+'�~�:���!�U�+Vse�j6N�	R�P�|W�S�rK���҅K�;(ߗ	�=U˒�Əq*�Wq�Dq��NǔR�#WϺc`��7p��^ۇ_j�0���hB
����c]�9�Do
�|H� �DM�e��x�>�����gb�
��/��@���:MM#����s��[��A0���<�M�F\�h�r=~"Y�Y�3�S��>ʣ��99}���������q���$O��JM_J��^>�w�>Fq7�W�A�b����g���hF�n{_�L{�����,4
��/�%�3ך��7���1g������ C�Qu2��<�J�q\��{��e�N��KEbj���Y��Y�~=~w�.<0{�~�
�5S��9p��[+�bM~��7�)G�l��q5�����ނ8lE���m��'��%rS_��=Y$Q�����7�Nө�^�v���g�ܖ�=�v�:tk�]�<~���Tz����q��`q��! ��Z�d��9`��Ny��>�������2/F��5���4w��'ܳgB��E���F�ފܞ̷>Ft'$���R4�UkK'(�����VK�䞴�~��У�Yt�V�6!�0���{���	��v��:��iTү>�I^����!)~E���h�(����6R�Ѳ�:
��V%�j������]Q[&~�d���>dV�ű��\2��pؠR7��~`A�;�OAb���9LܐE��;�9[�GD�A���^�{D��y���}�r��V���g)\.$���X$���9��*[2��!@���/��ҟ�����z���U���5v}7��4S#R���b1Ý�<֌�9�X��Js�=�W܎t�5k�<�8�U�R�tq��.��RxY��!�W?Л<���;,	Ŋ��u�S��/��8������f}�P�����;J����m��ԁ�MjYv�s�f�p�I��c�ߦ���8-�p�7�>��S2�ҫ��Vf��W &}j���bDd��8���2 �s��&�D>�|��db����M���/���ԝ�r�:���II%���Tf������غ*�4��8p���mЧ g@�#�]ԓ��A��jCR������Kʕ�Rc��M��7���"��(NOzQ�q��;�R�����:�$����X��)ل"�f%��0���|jO���l�RG�P�0u?��阯j�1r����V]��A�qY��rV�W;I^z($��ƒaFC�c6���HL��->��1�om~���yڣB���َR�G��WR�,�G(�O��=�R������㞭+a}���xK\.-��Bp[Ϡ�s@������z�HBX@��X��WM)��iUtږ��<���8���z�B���,R���\ZyZ��e�T�����v�v�!Hк��-jwL6�N}uk��Ew?�i�l2�#�"��j*O�7p�5�����̏��B��r�������v��0�I��ܝ�F$��mQF�֞�on'C�`�z�XP0C��Mp�%7����T\�s׵k�x�a%Ǡ=�u�t{K��W��/�6����k:���/���ަ�wZ���u�E#�����>�� S%