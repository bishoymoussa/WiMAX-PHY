-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
0Z3Rxgo2nM7JWX974LDtPdFN/tmXHYSCwchz4Oc1fWNdH9Sy1MLVH1LyPK87Jjf+wkGUSntK6Y5Q
e9mfAy4QPcAvptQjprGocztVdFIJ2eFua1BMLgEJJbMaWK8jQVoIhwoRq592MX8rMB85e9TtxK7H
W1jU2BFm1L50DDbXnx1Bi4vvJ1z/XvPxh2MqHSaN+4Ow1Hi0S0DfghmyMJhZB+fUhG27uossYqv/
hOvL7DCeB7npamuzajS4UuCHrbSRuvOJfrElXTUGc2WoZBNrkdMVhup/lKdbvG1HSysaa3mw8TmH
InJJ7PfgnRI2N5CD0FWbiRYgctDVtoSKv4ALUQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 10592)
`protect data_block
KASSJXW6lNs1gCF6GMJe+3THPBgqbWpwYNoMapz4vbXnmxENp3rONVJ4/g4P6Ki+l87qeYzupoqg
mS0XckblcOt0yTTbuv1V3p/1PmYoWKsV3qgjyB/IaxR9Aplcgy9lJabg/T9pj6m5aozd/smUFjjs
rd6ZkY58KQvHXbcSWBb6XJtGGpoR1LDb5naRuwYapTIgZ8hA0cayXHkFB+Aet7XUAQdsO6ml3RwR
U3g9sTEwRO8569rTSCBkUViXQJfbQgQlqyafTUASeKcSYxvQHvgaXi6tTCPW9P/fVEDNZqFREB1r
BXmuTV2dWqb6+gsikzpog3OjByXgS2Ea/DwZCecDPy1tcpV3JwL0KbOkxy/xtwgAE8stRb9C1t+D
iqeZ7uDXYKyiUEi+bzEWrRIVQn8EiWEnx4tl/lAFeemIX0CH4VwsZnm/q1I0IyGFkfBzcqBEAsUG
41nyOUziejmsK8wsUIa0IU3U2kyhbZo5tSa55u19YCsLhMe8S8Q9PjPVPAyQqdkiDRfJlI3nwV2j
OhzlPZieJ++C/dsZILAR/zVuYj1PJsqDXFVFutR9/IECKL2iYdmjkSUegcz8krH6M/CYaYVsDIFJ
ZrVx7dF/vrKSuMXREHpLn/oFlZLxUXBHagVyB7l5PwSovXnhYhBHZXCyHYTHCeRghHTbYaEyGIS9
QQHpZxUQqURHP7KRYunwdlicrP2TD02Un1Y59m7JwrDaeD2rfoWAu4ZD5UGlPoMKrUfRAfVO35RZ
IpUn8Mhe3f2KwUfa8YyjUDjWZmK4JVuaV5uFpidYtHIrRiHw7C/0R/ausRV/lUagEdG9x9zDjryf
5OfuA96GRwU10duDvv0LL/klr3iSVGchN/vunX4WBKgLI+UV9YASQa8MWIPxwE240zDKGQ1Khx2j
hRZ/yMsNgszjT34ORlOvsLoqkccElH/23hQvp1rQb5pEaiQmsB7I5h6b8egygTrjLZVW+IlhASQr
SObE/W02i9y0wy0x2CixlvvW29dCnV69W/o6xnGVpNHfd+AeZnb3DR2X3Bh8tEo5ibWr5CJvDcJw
NUaG6yA6s61/8thgctYwi52XE3Q1b4MQrEtKQoFxmRYiz0+pyXBWU0bfa5TRP3u1TiOLHTwLN8hO
VZkAj2MZ3d5ZNUuTosGKsIB4CjrXCjKX/9zUGE57aVlCuWfvnBzH7uwYrvQG+66I7JyqVApxyg7M
TF8ErIuWg/klxwlmcICD5nIyqrugOxI1f7xxQTLtVrb2lgKxBxZ9XrttAJMUTzNE1tWWV85Kgb5l
hP2b/qVUJVEagnhLznbic6vWMfYKspMY3HobWHp/JAGzO6nzZDna7aakDk8Bw823kS3i+XB8stZo
ndWxrmkRUJWAlzx0EOtHdIZS6R32FZuyYikvKxnb0wQbeaVVg+BqNJ7wU/U59SWP4luISZxXchpr
S9zIW6Kzjgwc60wIYiWQItY1iQdr2TPxm2UlgQr1uTwhUGaLZ2YYob36W5/pciy7QYE7L2aLkh5X
aBOOqla8FPV7o1i/AJEMcgWWDeUjaqRUbg8F3d12CU3FxhLOeBQaHf27NoNYk49Xu0in4JKCecBO
PsfP61JX+q5be+v8Z5zBPvu2aPYEwi4tXJRe+unmfqu1DYqSILPL2yfDzGXc2h/b5duJxSXAEemj
uLQRHSKMNmthicXB5VzHo8x294YBEaE82tzHQMlpRy7UiN39vzY12FJqqZyJYbtMXMMBMHT1NfaU
+tMjbyllX5jlJ0ctIGLQg1tCzJrMcxu24C3pbfrVdbkcVnjfnVroHvFE8zOZ/BQoJBCFlKkquw1x
ewTGAzS4x+hvoNNZKLP3TrvBSq2urTuZiz5wK7Al/qAxCN38FaTwpiKW29LzCU7PuvOezHtBkkGq
R4jX0Xz9+eNMLmjq4IqdylM2TGRpEu1AYLERkOqb0+VRVS7/HSv2g8VLs9t8oXn1XvrhSdKoeUwv
t913rYltSfavgI1yBZcb5pV+TScmtjZnqKxeVN5cIH8ipsqvEj702sraOhWfZCdRDE2fhQFXGpoN
DwbJA/S8U/zNUJr507Q3n3GPxy0U+85E52Y/9TGSFgwa+tXFRgaE+OdY+nYPQTj1XvNYuDGMAAut
7x+2sAVaB8tJZ1Ehu/ClBeC2cSwT32FqacxIErJgVdAE0SyejzSDvWhdPFPJs/UzGBV21w6VJHmf
FcNCIfvRB0TAautQkh7RDrFq2zV3b5nsIkWq4KFW8out3kvxTg/D9ySDGTc0jmL524EwkySLxWWx
wfge78U5sHYmkhtpCsmhFlHLh7FN0AgBnr13RNIX6aHIf9KKP1JLvVGRkaN+zbZl99Mf5XOzDWzu
zB7NdWg3QG1kgDyTW6LRjR7Nyf5xHR27HCrMlXnRBLuUPNi3Uq9DYrRQozKSx9H6mVGLPl4Hz5NJ
EBFreuO40hnJgG3mwP1GEaYNK2ASnBuzGzfh/A+tFzdX8Cx+GFNleJjQ+CSNLMoJPyZLNx6LtCYo
EflgCl/wjlxU8Ypo+CTHSZD6zYuv1gwbMSYmbJf67NtMUJKlVLypK8zT+B6x/uVmTxicbnvpWdt3
5hPQv4vWJlHkxHKQQXd4xmJvCe2hSltRDdn6VvzfpUDGefe8OK3JRIWkYrpZf4566vdC9DbEhU08
OQzMWwOieMha21RWOR+TibcCdY5SP2zl4QMS9gC4R7JrAuUIhCxi32OzfBXXLGHFALHDqcLNAffN
riw2tN7M10jttVJA9Hbh+NXBQK4vBvspVsk3W+jN5nRjiOWum7yV6w4kEL+maxgLsFFeIAMvovWZ
9HVhZPDt4R+lNIcDXljyzyPpqIgk/zn/k8nADyZeVjNGH0Zjdy/vx1nRqMIfn/Dkx44cOFN9R0vO
zlQeK9b6zA3H/sW0fyDWRSKr2MoH2D3W2K5y8+WqOn4o5sb+qyS6sYDs0xTiRW+oDe1pGy4d1ls1
SkXsHRXlZSiQqkyt+PSsJEcWrMfMNHPOnNyNKgiLA1qQzH7d+k3z2BAZ3vAG4o1Dz42/NrMJGrZl
SSGaD8CEldI4BR5hZc2UThBZ9jLvt00WG5Hax1PWN01v0H2Z8RxKqB/uk4xsM6SmOk1mNvUbYa61
PtTGxg2socLTuTm5ZRSbBUSO/C+UtaWGXdJFXDXjzkfDI1SvzJD0AooFCRxi+ry/0er20PXJviNs
XiWcSe5eXyuBtnJIFpbMt1iJOhVACufpXriI8Rqy6pznNT1gWiZVWZqb849r03OU2hH1UcJ/dmY3
QCnRz9GAiPcLAy2D6MBRE5DPb5Kwu65XcENZYg/XDcVjpapcs7gEs6UpnbM23/0u0j4xcWg/7BpL
Zp7lPbDsHFC9BrOguM8Du3L0FxCeSqxlOBganexaiDAUQx83mdw1JoHmzEmXjANOJkYUy4dRlYFM
AZMjwGPZaj5dpgQx2lQOpCSBUN9503WCfp3YF07oEpq8e1+nV0vAFHoUN5/jsAqMPcwHmMHBn0Ow
k+JcGewz69PmayxlYihlpVyFewkIxtQ4+UcOk+C3emCioWcFdNwAEn0KDh46Pm3bWIIkwzi1gE4d
g97pkRtgCctG7yatzf+WblzWb5LkS+e6VHktBfJB7cjFj9m/u2D6WhmNIaIcYE2cCv0GD4RDEVhW
BLLfrJJ72HIlUPZoj1S6urySgXimDodlTQDAJSjazCZD24Anf3SpiQDvjrzPxoGIg5BTQYeF46PF
GE/rBQFxxTUfgbSO13K7lWLmhWIxVP6Zw9v/D7mlhCDHjBNJflFF+1EPwb71SsGgPoDxj9PycZtD
LVqigd4334aXVt20UT0udj6BzgCUKhikRJaCAUeyyTIj9S0+riMftahYnOyCrowH/fvHLEwemEsS
30Kb5DRPtzvkOwrPQ+Aoa6P3mYdiOJqHBmFvd/0vESy9cSHUBy55IIXFjJcNPdtFjojfBAeC+Fa2
ZMf4FoWeK7FCtHjNsJtV3YlqNI+Jzxabx5ruTa86HccTcOZCxyDAulBjbs4oV6vJf7DdiB6ytSUO
vAFrS/+0YJQLR2z/T01PLk2l489oFfeT7eTJIelGxvf1WbbrBEMjnIAlQVLPL8a7oRGoW/cny/gu
5Gxw1Bof4qEvJi6+MuQG9LDJnM9PZpwvl0mugM3+kxAtvV4UEukh08RMkwnfxaNlGPYIWdcCwXvL
cdj8tyGO6oxY8pU5QgVy1+u5rSmA06jkjWva3qzodUN5SD9OBBPV5+RcomWA4KHHSbwdKAmf46yy
m90cl7pGYbGo6+Xn5zPeTGB0ZxW9fE2EwczrfI4BuK+cgnD+WLS3h/QI29hIdDlqotwUWXVSt/gq
lE8yGZqZehhVI20ngbTv6IGbEkxw4djA8QeGpqzT3oUeuuhCUYlkJIucaD4loDc0WzETyAfVEPqo
wchzpYNSmoPfURzBAY6tMbAmaSS+Hv/usyrJVxpiGppMV1Lqc7ju3hc9vTTmDLAzDptGOrLowE/U
6umOcqWKelPTMf4TYAVBm7YA1LPMLbftMAETPfVaEyyJ2scvRe3tYUerV+aiNKk0A9b468ctNi1B
ticw0TNqNtDTEEr2GKehRloHrxG6rF55BmRNH9+a//JT0KGkvf6MMjAka6Qf7pnaW+i6ZGO01gcy
hMY4UOMc5n0K18QqlC2q76mjysDEpnKnAqzJ/Ya1SlsNDFkbPoSWKPDW+Irp4S/6YfA1lF+wrbyf
+5A3Rsmx3uJ1df9RaUHHEamW3At2JJNRgw1NX8dC8j/OQSmcdbHOdCMj8TaP08LNTKy6mdG+Glst
BWWT7PEyheOoyH0FDsTxfC24Cv6vyLtkvAxh2fRA1vCRewsPZIP3XVsuESJh6ycAW5e0Eh7IF+U0
piZO1aMZlIZuSGU7PcuxI2erhcu9u97CcOkRTsg+Y5Z53DCynzCMScCWVA5mUagMz9Clw/xDMibV
shNTEkP+YnTe/th7O2w4Ki+B9qpil92DxPzzH9ZgiEEFH3DQR+EyAGttJsDOJfg8qwZ5HvMm2Nl2
3fYjNHlv8/atc13JBcDky1W3umYIoe4inh7cc+sdXf+dmXwkq5ypmgyVjpvKgfv7Xk2lD4PMsnf4
JUZBrSEfVm5YXz7VNydEaLACJA875JH6MFtWmu3PfupxOFdl6o/ENWYnsUp1hWumVYsgEZUefceD
9P1NUIUiF/LJt0/l6MKMKeBGAmXkgoXu7v8I+61KMlGxxdpHssa8VPzxYkZUxCVR8DgqxdoPi8cv
4lPNUCM+k6yoQu/R9k67oTtPddyN5muE54nTvn3IrYAnoUuxoNJOqr3EQLzK2TmxcobuVjkFTQUR
IgDOz+8ge5df1MF/0ly4Y0hZE/eqBrGfoUR6W9XDj/bNIZlNUbozg0TaC+P1LTJ84GQ5ySlWKR0f
AFgTZLf0l3xG5yYIAKvZEmdfSUyOSIpesc5tTmyr/P9eUEEflixoem4rbdBjNU6R00xZasSiHX0R
sHYtPbmI2z7jpXnXMePX543So4s9xlttI95y9QOQRqylViR4V7HGL6beAJsv5B45T1PtG6s8JHNB
IRqMUmgft3UONJHS4Z/Uq9KAawcVklDE1y47hyXRwFORDhxlCHx0/vIYVFe47F8bFrenUr4LYVSP
4osPSXB8VbCV5jLukl7wR57qjWJ57ITiBbCY4A9kDAbBW2cWFG1gu9x5mFovGvirIjSerFRnv4QD
GPs6/LEs1D2UEhZNxiEfs/iTD0wasthWZn8Ejy6cBt/o9AaR7W4gdZE4U4AaLdddX3DqhUQcqB8M
YJG0jc0rNhBnbk5F2riGSdHuQoVkQc7EL2sEqgMFw7VyNTu0h91p5kL2ArCLNPYNh1rTI4hta4tJ
dw3rPOx3iZNuba4tcRrbdO7ikwAdAq0MKKqOv4AwAuTBVazf7Qgtn5eh2Of8nq1rT4ULZVx02BGX
mNx36p0X9wvlelRPRwNeAnHrf2LftyLdyyL4LGZuPa2RpRrS7mVofE++3fXcezyec0+z6lp/CaPV
fkSPaI3L/ju+6AJ4LGe7O+4KGL+sW1tYYU5plMcKasaDxsSwhKc+jXCVAo/BcwMbftCzhw5pA3aa
pJS3S0wePEd2vtB73DZMHCXFTzOjtlVhF6LYrRYPxCxmLRy5Qn8G2xkuu7ulay/C1jwLLWecwagi
qf9P39Xy0Ad8rA2aN0odkAqAl6KbnPYw059NBYpfayzEwwMSFCuErzJh3KOQHbyGmOckh/NQ89jj
3PBpBEFhAlU5Isw1m5H7w4bQ1M6RnEHZ4B9Hvg/7c+mSeQELu+tDIMZ180Rpz2H4PHnAvirMpdON
PGexV7wWVR+VT2MZcEH7CcCO/e9fw92ApRKUGACaUh0Nmv9IPK6fKPNXVSaBHpS3R3jnLimdNbx1
Gm6YTC0KwZjoiJpd2cCfFfitroTK/RhZouSoeayZUk1kbICZWVNM+0xyIZpAYxQhpwfohD5ow3Qv
FgqWG6x9k4MA+Js/74DZl7slP6QMyehsKhTPIs+DrkNk2JQ2C5jQA1aD0S8KqEQB2BNUJID9IGHk
U9C2Vc1Ey2UJP+YHBZIIrqnWbUdX5FXdx/h1FxrqIf1RT7y4a2RSL1BH6KPbqhkEuwo2Oiv5sLu/
8BQLexpK/usA+GuIfPcbYO9QyTDn4KrzgP9nPSZHwS9AwS0E+yc7wE7rC1gQ+mnJ+ZlZesXBgNr3
GlJxh9h8sZznbk0Bgd/rxws9rOjNTv2tstq3o3r08Ups6VpHK/B28kWIVFQoCJYKUfdcGAtzUU8p
gj1x48GfQfvX82cpItSPhZKCbe4jVstncWXX19BTKhiiUkUz20h51IXyqr0DNiLuBKMGddHwCfZa
fZ2ifuWI3OxW1AowqyMwhy62vh0PwpmI/bjPVh4bepovGYo8DaZ0xHgBjY9KnWAga2jsReV5quXb
bPS25+d2IIYo47OwOnO0KHT+TK7D6zDLmSa7BT7ka4VEktD7Izv3DjKXghoT25w2iOeaKOUJqU7V
mCpYUmPAq8opmOGv9q7RdfbhG6+QwoKQPBgfdafEuH4Fn7wj9+JvB5Fv6CSbHBChxS/gjGe92sQ/
kmnrQHC0UFhdqMqYwZkhhWUlLUBbbXuIa7ixt8JkdY1RxeJvXIdmATDam7DQTiqtstVaY2HPOwiz
KrRrapeqAkL5770n2WMuC61o1yFV5Riz4hLdyIo5fLW9+FIcFKleQUKywpH+rDopDsTqFuTXW0N9
6VDq0Ug90slyUTXuUfw3VbtmbHQmmOCc7nkdalUzsI0LGfClEElxZFFS3qICURkOIBcZ0kZIP3HR
RWlzv4au7rPWe8Ovw88ibaxjUXZ5YqA7pcj0+neFlT8D7UBATzIf3FqSWnaz7VMlLuPCNvxRfJy7
1pb4Nki/6c3w9WZky1/X/Zuila/v+1wofdj4NRVsyDX9NoTmBMG9SQUMzDzuPH5rRXXQ59kwWVz0
xQPvrnGyHHSKQ7Z6QlvqsXKjKZwPcHLWCC2BoGGlC6J3tkTmF5qGn0xAM3zZUowsPZYzMLb7Ywz5
4x3OpQSD+w5H0ZrXc7PTwgKL8G/DqIYTxBDSEnB9h1DnZm4LO0xC3Q5S2kHULLUnsZC53dFJPiWq
LFZIvXYanrfTiuH2AmKTK3hoM3e4lAKhGjWmTn7NAyEQV9zh7Ug54nNG5pkuELIFhk0aLvPX/W63
jSGRYDYu8ZavLlpplOvkciYRbN6H2OB7UqXhJMnoo6+7/G9Tc2cAS4WJy6oU5Im7hpWvg80SLghE
9w2UXs+0fNpU9gF4jB40vQqrfntHqvDRrm+pei2XRy+KtSGh3yTce5tn1+pI1MQHxnNsP46FD9Bb
bWvhUXhlKg6snyj3yzn2hPtUlV2fER/ZduwhZVNuNeCfbVyf17+gmKcQ20rvUL73s2qWCyyB+BH/
Ie7OShVyA6s0U1rx/9U40+1Ce20DC5o/3Z3awxJnRsknhUaSZ1IgewoJ06FvB19ybUWhEPvblu/P
qgAYEKkaDwSokXwjFMPJ9ve62ICLNB+blQt6PxiRw1KX0Hd3UkLiH6tRYUf/4RSzEXxDks5ZLWrv
5Dmt46hnPc/4mzp/o4sHBoSktlqenxk2INy6TToj6O4akHr2LhmApUCKcFlJxbKYSVFSoZBAnP5q
ssx7AnDNyXT3sSv/9/Y9knyW006ObOM0OKbN0ixvpZPm8sHMOqjHd4PIDWPrtgokwPW17k08QPcO
yH58NstJufgWDuzEWtQKmAsjATvFJU0Fj7aU6CFoOxCP1YJSQu7Ue/ZxWm/BCGroT0yCoHvm6Iqr
4l/hWDNdGrCPvkQoBstkKUhhPycdYT7E5KDYvtnP8CzRswlkrjQo3dZ0y11opssHQlbxlv+EqBJu
4eivxy964mJh5MDm+PemFTEnpnKNRGN92mA7KdX6YLiDr1WXx0jQKLK0adeBdeSZ9I9rgxl707qo
U95LGOpjig/nt0a0hn+2OCKDpLyCDSP1W0QICSH4vpbcPaZJ1/jqoryqC4z6C2b7hWc+23U9PapD
dE2alHj7S2fLrX+0mgRa9Zre3mMrVd8A6VmvL7aKDxIXDSrqynkUX/fwbyxeZ97E+cwFp+rNtymq
gAH5GNeL9G0ivUC53VlBTHluVkiIOqIHy5WH9ZZpuL/mBbpBydhsQNExfGPi8RXhhtsTwiaIn5Xx
u/wkpPA5HLmT5/9dN2HjqvCfFZHs90Oevv0UOn9U98rr3vglbWFNNFrMHtkq/Ru/a0A2GNfbQJyp
4gdA4l3rzszyiX8j3O8D21qa5TAxQirdMvrRgRyCyR4+smdxeMPNMgKf4oBc0NpZduKshr2ohSFQ
09S+5l+4phENxYLEqXuj21/eXIa1ZI+dUhv15OY72E7YEIj0MWRPP8R1VJDfvaJhzIyzhmyvPtpV
1IF59jMZflB5UVBpZ14kEiB5Aj8dJTb/52Y0BBzH3FLj8QF0JlNP2hhK5To03Y22g6OMzlSzHkW6
5NAD0vog5n7poIdiOmRVaIgZnuq5N+jir5/zPDN2ugwtn2ECjUBYvmy7z9e+ez+4D1jL36xWbBx2
6vgGytjpQXLuuy0Wbyq28FzonhWehaiT15NrB37zKdwFMwk6MAc3GVrkNlMl9mQbgrB8F9OiaT74
mCBrR3Mp4AMdFcoFT1HitsgwcJ+NK7YWF5sUTDZlTWX84+FZCtnGyNbJigPm7nAXbGfL5ud2tahw
xZGkZTxwRQgXfGwjrJBdHNO9GQPJ24bbSiiyCd3cC3CpcxuMsKd+DAF39c/I5DvgnkjkpHT+qHXV
fzDwoFjJjUJtR4djhGP9pykJFOi/43fDxZLAKdNj+Y4lwlher3YgO5oBs/w0KzVkzC3C5BFBV0iC
mqscQDhZ0HfZEsUIC4GADVM+lYpkK73Tdyp9mohgsq/hN4jvh93SNTgMGMwlatnPZc9hZ1oTF1VX
P4o/rppVE+E8okgQXxZAroCifta4yilIg7qmt2Eim1YF6b+dniILedFEsQnl45yHoHhADJIWdB6N
CCkm6m/FQb4guxFSYU8h+fQhvlrPI1GjyD4P+pHr/X6+mFzVabND5l2y0Nq5dERo9Y6ihXnwo+A9
C78/T8B+sojQMXXjNaXA4UWhelBzXhK/knje4JQKrQW1bqdM/Cjcc1fdBOcGQ/N/KfKSAwWAOZfa
QTwId1FPKdU6St53az48ko2ZSXY4mgk4sc+nOPbwasjSPiARq+zqM07A70VUtEOuK0dnm+sxWsXV
ZMEK7tHMf8z06nZpGG9o1praTqP5vr37uVFCjSAQriqDk/k3ocj+xcs5/XIu8mJS0VKQK2UChyPr
YqegRxQhWCU5JzSXerMENc5gXo667LpPPFGNE2RbvDHNvYJ+aRnKxTv6S0N30LBsNHYQhjF55Vl8
LyRVo/V1IBUovNBDnJ3jagHyI52y1BB2vu5PSk3Z5wbbQ5AOLqB2rraCC4Qmi4qq7vgMH/iC1e4C
/ROgQ9EPIN4v3eSgonsGh6DyZn5NoNy5NXwmWO5Ry+CSV5hfTT4bdFoCzXza18xk9lW71qDLt1x4
si+/mLUzLpGrVj7Qya6gbndg0ZzAFKIpyFZZH0Ctg6s1HzvINOtOrgZiGX9IMjJIxSGFHVPliXj4
J3N/V0Fx1fIh7bivn7OaCD3GS8fWbBv8NC5at7hWkweGbxhj681O1vXDYk5sPAbqVMRmotIE8oVr
+uVtcSBq0VfUMob2Ve0Eb7VaWPtWR0HQl19+2yKDn2ILzxPYYJ2U5reDfnj/CDLoDveWmCnCIdFn
o2Mzf97wX0KgCmuAAKoXaXiII76dRANbqiWmLQvBLkxIt9SEs0Ckgf74AgjTnh+frsT3pel8g+yR
7Hg26ZgYQojSUA5wQSVxmPrxJccuIlYCAggCUj/NbQfsMurrL/bvwOmNiR1T6cCXQ70XdobpjfPw
ZiGAHBw9o6enwEE1TV+DyIH9HLwfsWmHHIxCLXFb6rW8j3NpMpsJ51gkYThzS/0P2OpTS6l+TiUm
ybKjRuuNTJ0HJ6s3ycMmHfba3kh+I0aX7gYZGd+0SIBiz74fWTe9omjJzPRVRTMV9gfXHAJ6y3Av
1ksNInOYsczu9rk7nCO8bwxMDHWXZuYvqWIgBijiEXMQ37soJ1hQduSHRf6UmhVGzLVzaV9s9Yte
bGjUffnPjclTjwwZfSg/5/Ymi7lGXnpsIy8DE/qflmWbj3Z0y1sNTA2J/Bvj5O6igq9wKSr9NWIZ
pvYorEDaxtoVqk9XIM/KmojC9vBA53JZbT5fPhsSNLE+YgZvPjqoq1atUvvGURcp3JnZ9PxrluJ2
AAMNLGWc5nJL5uycadwLwd5VKpcThD9rrXR+noY6gnsWtltKxOFopDpseRV7ACf88Yot64Tl48qE
q0Ss6bqORhhGvPcy2BuSsy8QLSoEYrRledORpaApIhDjxo7ggfRlT2OGsN3Lcfh6YDdS535h4ZK4
g9a/UTQGhBw4Y5uz1bJpsxtXXPnC4ihaAbAeyEz9OZfivPbDpo3PTTlLzqZZHXaofX5ZdTEsXyWw
7Vavr2kyI42KWTH+nzcuR4FjYS2UIPcU5aSWc0VGvjXEXt/7FR1/Xjp/fgdg3WBFo5lEJwRO73id
+ljKfapADzVC7OWzDZ2lbbG8jS2MRrYsRm8jO+k+K3IMtWQETJoslAS4ta56PtXyivd0Fe+kGKk3
jMXLxUVhP/FTP2E8mjspHTYPrLV1DOfZdZ46lJgr/vWLuj6byHyTbHmAH8WXtrXC+96WluatqkOz
gpxfGJ13w9gwORERNeJrOuDdWqg02JFmhqbbT9pE8vEr+YedJm81X1pEfxKJU1wDta9lo0uooQsY
oob9U62lmieiPDAYybOdXup6nafN3eonL1nfcPyN+UcrTmfQDGK+w14HQV6aFhffI5wymt7hapM9
phDpej6TEWKGUuxfVvzMPsXb1bO9jZpK52S1gRHbTPGleMjdw3jlKfHTN9WzVtu9o62Wq4bRhVJ+
uD7c87x8wMRAbRkr1y7qz+qlzyc7+Y2z8uyZ2E+35q2bPfM2XY10rZgFmcibjdoHffnM4ci/xeiP
ekfB2NVnKWRKPf9LA8FBPwvwg2N4NQLwoonqhFxN0ZldlS0gP551wip29r8/vM5XUp7Jkwi4cXn4
FvaJqsQk/Jng+8BHa14me0M9MGetTR6k7Kn/TR4yEDyZ/34+EbU9+IuPwQbzljiQvNSxex4Gx7TK
NkzCrNto4rJaalaFSXaxW3RyuAAH+dE3zRZ4bQETgc7Y0sM2oWdn2hvwJ+lLbAkoQEZSGpU/aDkM
0QL+eQSfrlG6WdUf13JzFV+JHqod+qg7oeqE62bqs/XkYu2Iio3PSB12ycLqZV8p34wXPCNOpK7P
1WRp4zGVtT/umq1VxntW4bc4cFVxKkMtUBTA0FrbGzR00r6uBevPcdjPRnC/eW1xdS3wP5SqyXz7
pjYuoku5JGEPFTsdNIFIFWNrRRuiLePMbWpTCHVf9LRMj9erq/YZvVLEbrn7HfhuiQ0P/uGBQwlf
hwExvQBxFMKNBeE+74YJgGcAfowaf0CRSI5lKJk9haQx6wXqZaD7k37i2HwKs1QdMTKuAcarFDr/
zkN/Ec4BZUbwadNqIGiVQFvz3gJ8gg5sjF1iyeNq/AF88nArTeztcmStqXv1Y5ouzEM78/Yaip1d
xl2Dx6+d/EZugkcc0Ya6/W0GbNoqEFk7gGS9SlbMxbEWUIqJskAjb2WXk3TmwH+orlH01K1Vv0wi
t2cZnMV8gyAKaJWXH+HMiC5g9kilQriS4Hlp1+DBcLkhzSCk/Zy7MJV57fuzoeGqbmHR/8xdpj1U
etHjHpwJASum3mC0inlnaCTtIDOwsisiZpDBhjHvfVD0lLrOFYKGlfDG0iiS8b1+vzSlI5FoUUMI
gt3DauFHvdnwYsse3LRFEeVmL0OisZ7ywRpiCqmeLDJ3d2MNJkcR6TyOz+Nj4cffrzuOUZaI+8IC
KFZu/8QUveyhWhUdOUv1TArshpibbKsj1t3wGb/MEygM9w+AXXuBMomZAgDX223+oRkoeGXJoDCG
ptCAENuc9Xwzaig5UX8e+9stAOQwKfAngz2AhXo3LgnhccB7WdG68zdqWoTggHek3ppPCljDy8FR
J2XReyJ8TqRJJO7sb0/rwZvEgM6z8DVAW4amuD5vNRfbeU7/tJHOyTxfYkuDzdE1GN8wqK/jHndw
kbN5q0wO4/ghhZlwT+xxJuuKG2EIbjs/sP9V0mpMQSJa4Zw8bZsdzGFRjo5HleZoeFBIKsl2E8bK
rBiK5rO/qLUnK/borPPGSOfLS/I5pFdFDlRNkzv4Vpy53dENdNaa1zo+9xfzyUtvztLGn540OzTm
W+f08h/dtgI0gaE8AdFxGsIh7BAc90hZMh9S/gkytIMjCihiwkToF1RJUEi72K2GtFQI6J75y5ji
8iDlqw/wxb44Y6AFnEnC5ZyV/T8BGfMzlRBdsZD3ZkMTBd4umCVmkeH9ki3YLN3s9GelHGh1zO8/
GW1JBRzenggrbcsGWC0ZsSKITazLjd2oVeGHJWCSg7MP8wrt2LFy/VBo86YHy0YjNZRezab9vT3j
smdigLJGDdfEyAtgr/Lax445FjkfnnG34iA2/WkaSvJwgptxmdoFOtQUzhJG553t/qXK7NEvm4+s
pXZYXKZ+7rv8rsE6ej+LZoVy4+QgaZmQHPbbeshsJ77mKtGe4YBGTKwX2lC10brbpohkUQuG1Ll0
sEDxU92vVnCCV9o/ZyS1ECO94BnFz97GOIyVugS3iqsdUshy0f+oeV00sgIyQRatpfs3PzOJMUCQ
aIhfG728hzelpMQw4Rak0aardZApZ+APIK9NcI5sv58gAPzJqZ35/2GXE4Qnughk02/BxDA9zBuX
xRdpzArIqo+sfQewYp5mxpDg/D5R0wyw6ut07JNPEB8zh1Nw5BJSQrthbEA57LlKP/4OkC74yQOi
gz54kpmWvNzNNrxSoZBwEYq9YFbhSdzNVkEArd3MVmPf3Shn7IkUCBBMBp+dFv5hdnyZleB6yFra
TQ67jgGC9kFDHUEf86L7dPWtBgjnG4WA4nsapwjtxguTlU7hgZ5h2r6CGkIdwNwGsxnoi6CWUY6s
65jpC0GRwA+zhsD8xVcBUSLQYylSNdvFF4hnCvJWw03gWFOimZ6J5AXH+tca7GklIjcTM8+yIS1L
4J63QMpaX+tHzCL5sZEDm6OTGQC01Ku6CLq/+r5QcF6mdHMQxY980hLK6FinVb+6+6hC+HGsnIq9
C/jIh7Cz4IyLG3+Qygq2WFjK/dp+Dy1u55lEly9lS+I4/L+IeUMAjTfbJHm46gX8BrOPCCgduB9l
PK88kNhuwYEiQuZzit8CkcTuZryRjyAubrPFHR7c2x73B0BeXLVPbirtbqhVJ9mfVOiG1D97Dnsr
Dblk42KRrKSgob/aQRyy8nPFosDulofdm0l6BzN48pcl04vDZrYJs/zuaDvwKKcFHCMdcfzVnECx
y10KfjjgjR1ctmx5xq96WW+c+QjXPWN59h4yIPa7QBxi9vtRlDaLuWAbo+v1z8hqs4WGMwhhOWj4
nONFDcMYK1Xv/l6G/73lZJf5yMVYDHLD/XR68/s32IbvSWWeRA3jC3nUzkdpHC8=
`protect end_protected
