-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
nsJMDM0wjERKYlHJkAlz2l451XZ7PATNEuy3ayKT6IZXM2NX46Pvm9BrlARuaNU3+0g2hoIPA6No
atG78kTUbNHEvbhakHkfqcndrXWJl5Srycmchx8vD/4Yej799ORKFSM7boiTy5XnOdnvSuIiLT+O
sau4z6SF/GiRGM4UNtqCIyZtQR6ZwKEbIbu6FX8BqWK/Gt560MNR6OIcbYHp2jR2JYcPBnN5kqXz
adyNnIGjjmLEV0ptKUTnYLuXWIlSMYbWQo/KeEFNLZ7I0WXAIM8UkdL4Az9C3JQ7ntqvNarjiBRf
iZocs4Xh7AHj/SAOVmZDWtcgvpZh1hkkPhjg/A==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 37584)
`protect data_block
EnZTao8CMXEYy43fTrYQHuZ1pwsCFmuKMYBYAp/Je36MrKzA+JYF0dNEwCQndesJb0V1MxvH1MA5
0qO5TrW84RWb3WosEI4TaIN+7iOPXkZjh8xDuigKf710HVCEIUNjYc8hYxi57Pee1bVrqAf5g5S6
QtvlJolZ3iy1WObVWHCFkD7aBsk33LLJy9oKM+ByJLyVSKcw9dhG9r8HoMrzgGS0FVnBOTpIqL12
0CJYo/0Qoy0kWahvpG5ksSbMxXvNRBa5e8AfYUvYlAxWCMUrlmq5XdTvHtAaKl8hfIr57ep4w6y7
VHwe8oYYEhPhvisehl00VSTrmd+EPPVW9CrcOzU0CZVvV2E0w1US8RHAugl66Tha94iKFWdDd3+n
aJzNl7f7g+xqSkqZlSGuP1NZTu5JfCJI3asMi65g4+5bLhsGOHf60YVDGTQ2qG8DLLdnrlapw/H1
8HP022eRpG6MRvhpPO0Z6J4g/tsHkLyTQOBVL3s1CSPwzIHNU/zBvYzbK58V1S2g0uYDd4iTMRA7
uW7D6ATFei6gxXPh4A+BWe3jImvlKukIxW1NOHaMvz2VHrqkiTPXE1OoIl8OfecFkxiNL8rC06bQ
R28hDYgp1PP/vFCKmFf/xauVOywbgjvZgvYLtturFaassQcXWpWs3ShzzhKvXAKgk0L+nHF29ehy
Xds4TrAAetINSdMtxiZhb0hHC1Z67OalbRkZXyK4AwhYslZf3Z3bjhGtpcljzi1kkpD8JbasEsSD
VIMSCNBug3sPS8lP2t4wNGhGOVErWVxTBXJ3eCScaQIHTqsHjVm2fESB7YUQSeZt+01H0Ye8GKCx
NeWUfnAFNbJ8nmmOs0mTDiMXkpTwonL74sILUkH5m1meFJyZ2QzraE7fkPNbOS8k7ICwQxyk2FKe
mRN0A96Mx6zYraPVSK9UTRCw4kijK2PkJoEm6C77eETvEJ2OQ+zDyYHxdim4nXDiP9jl40/m2h60
/uIfyj8YS8IzbS7B8oFzeRgVBJtqFbbmVfu1EqJ4UfV/rLo1iVHAudLitD0ngHkf+QZcC4/dB9sx
+bbpfkad1sDJJ0ItfZ5jclKEMbeFRJdf+XBpcTMK/8cFF+AEO0vPzQpb7VBCkJyJZMlU/8ssYjmI
RaStJEf31wwG5IL0ENyJz2EW146qbjnD0pJ8v9FQBTd/Jsr1Ei/r1pZMbJpsWIlAMwNVyCfOIrGY
XSlXz61kgEKWxClrciVRrUSvz8ocwVDx/gdG5qx2tJQYgYY279GeBMX48OZaqAbw8MIjCCnu5HaH
yy6VUxyXPYgCYZtAGRCb3nmQLRa8LZWot2Gjc+AYe2sEDQgZk4D9ygcBjXwFSfZWKkkwEX+O3lXd
xGXE9aiAUJ5PVSh9K5PRhaOKCVUv6kXw7skBuMDGpQHmOOdyn46ntHEZ8QNEPXGtPdcD34nglkf6
HNM4e+6B1NSKxR+CQCTfjsMlS+FXcGrDKg3JEM/WxoTc7MdQZ9SA0GUYLdegCyOBpTfrU1JQj+su
yhixP+v/6LtPPeliB3fErBd4g6bQNAkAD/O1kyJWc3D5nTtVC5puNZLferd2dJlp8I75t+iZwqfP
/YRUoyeMKOUW0r2ELkewwcKo640c0p05D75inH8aKOHMbhLck4HSUZTWc6YEDZuovBnaCdDE0Ybt
ZKpaEL/NKHAuLoRtbz7f+MkaWGzzSf+EG3sbZD2eM1bqOU/s3ShIkEpicoSF19Z27Mc/5ck6oX9V
jW2yyu171Vvf1cCF8sYmeWBXe8rCbuw1ahV73hAVS2AOSjQngu9hVSkmETh2yULm4gJ4z4+7EeGc
tgCof4e4OZ3xqIvZ4EvzyCpZzfL7wVgUVoeBC9cekmpsiZVA0v3OoSS8erkOIJPQoEmYSXT37vlT
7lzB6G1YSDEnK/17tQc2pGY6WVr36Bb4I5vlIPa70d8LzdKW/PIWLMV+RzsXcjPnegS3C8nw6G5Y
WWvdEATkx+k6vENAOjTThWkzxtsAT+m5fObMPpBh1BDwHAd9Z4g1zjUyQKzFJR25hzozlS6w4zPX
WbivdzuAispK3Naf0ygzKsLS1xO8ro6A0JapSGEMwbOGQo40bOgaW8OSFJqYXwOZl13kNp5pq1Vz
sqMDkl+n4fWqOmXkfW6SXSlxZNSMRMuf6dJQj7XMrD7p9azsnvdHxvmBgK83OiEkzS3xk3049RhL
XDvr9meaJh2mM4ZCtD1myojqAiGFDDpP29WaUPoJD21aANu/4/Fufkm+j7dCXzrLovfzEUzbvasU
n/CJq7Ep54PdmcCsL3H93DQ+zN2JTrP7DLOXLJ7JC1Pp71v337kRhRsX+7uBGKEKeDEbEGcjhd3u
rMJzVdFo0gz5fzc4aljpbMgGrHNg0W4zXawWb3R6bT9ZMYDYcx3+fMftLOjTo8WM0Bs6e7JsnPHH
K8XN6KC/RYiKd2tYRRiF7MAgMqMPCUeIJYuh3q02lKp2RAT+ri2ZtPa74muixKKgLpt2EVt4on1V
KaS0Vzzhg4O3YSfXhu8JA+TFaqz7E6EDOyaFZCobRf7Ao++GcKktdF2lZyC5/wLuzPTTP9dUCtzf
rks8llOlvd4pMONQ7qz3kJ79BNkERv8n/23kOwvcSh7phWI0r1TkDp1hs9j/7xJBt4O8ALKJjEku
HJX81zNuXMi5CNkpJ4PO7CtvmlDyzNCPZuVzQLL1ftkcUndtMJhHP1rEvcWW+/DNGLpI1o7zLafN
W9mWpEAXl5ijRQ19Cd5bUw2+BDrQslKtdxGUSCF7oqAGHivZP8Ek/zVZCSLvuHmRmS6LiCqMHb5n
D+jZ+RjM2ZKvIUNsp51l4R+Uhn6TcoKqEuPBOOZqnuQPWuSQKUWD8jjmdrnsjFMg7hheu7Ttd081
sn0qGnlUgGQZQJZR7IK5yZre+vG9L9t9usZk6+zAjH9qckDd0zaj8LPwxKGKQIISt8388jjLXDQr
oaX3XepO+wJ1JlAKRTxg6H7PSRjZpMw8v/BJKrUZFL0gelwjgEIT1fhTMukte6vd4j6rc9t7hI9R
ZCIKd9XhFBGru17JW27dhz4Kuf7lu4Ihd5SGO1ZMgF/CrF4XLos70cKkPHwxRwl7xXjlZnduKTcn
UQ17Gt5GzVN+URbbB6tbPpSKQkzm5rWyleKm9HtvfTGv6AKzlHP/hcFhCqIBtzyfNp8FBC5/k5fk
q3+ys6Bh7tKqWsB0KbXX04Zh5lM7jagublyjKw33Vz/+CJwupPa4udqN7oMxOGV6eU6qOY8suCKK
H3lBPAiP7rHIbr0OOIqo34SlXBVm8SYb95DvvLKi3fM716JFhC6Sx5P+2iJb9C2N4pg5doQ0L3To
6tCfkbp2t8fLo4Ub8LBKyVRcdsGp/ghE6DgLiUFors6V65VGFG7OAhNHHXs0qWpJ8+zsobLfjm5C
m+BAGd1PQKpyT+lhl/7nhDe1FV4ILkks9yUycQFud+XIsZIm7jpOgtfTX3TrNnDzUN4boiHKYPeJ
woXqTTpY2YC79VGkUjnMQ2H1R/eWmAEMWgdg/+22zGG083pd+CFX8Iq4+wzTuPBjrOhz3T+r0FFT
D4hD55pwnFMd2CdT0rKnVBqQP2vdr0+fLJsODt1DzxrZUPJ0rxAup+o0UPoiUnsHpDE23amuD328
65oMnMxkO9bQtJ5AVQzDf8vYBVzmR7/AumgaIZi/6jYsb5WXL7SyV82ah6+JW9FNnWKyAKIZGtIj
jZbVJvlebQl0jdNqGs/jOHZxoYp/tpLOHNA3D40fvlWNgSslY4GI11a9Z1JvG9ZTlLwGCRepsAHE
mLxJG/rgUEgETl+lfBtMxhMkFLrkqHejFXpeV2j8kJVOV2dSmhir3WK6GQjFao8qFf8rh6OTBEjr
fJJu5PP40Nkt8DBwseMDeKpEU22h0qhG2GyNocS/pbTymBiL+Xbo0GjVviOyYS1ogkQcpZQgi/VS
eKSlPZ3yn8Ibgvdc7RzT26kUsw6/DL0bCqIXvfLh4taMh0Hq5QljAFLEQOsr0mdq1buESpZEoHcv
Q1faWHU8Z/qd76Um13/QXkXpTd6xXnTGm4v0a2p/5lc8Z5QaM1QRb9K7rC43OU/iqQDrAe+0Rcwu
fCtODtyHMzRZUjduNUk9jxT6/usQ3DR7JVhPI+afVjAypRT8Yl8fxsyZV0KUbRiUVCN4uFBDjCw3
sysG5TiibVKUH2xyL7fX05jAKufj2/iBtx++b4fmigvewdnOvAsqqCFAZW6diXQqsWC09DQUwegi
wPWtogjJQmTehIjQkbU+F4lKkMhfh1Uj+aKGNKaPxIQ6jc8OZ2we10CuKt+xoTFrnzVtGqSKpxxl
t46mH04eyd5zyrAQHYDtgl8/q8WSOWjRe2wBPd6SmQVGkZw1wDI8tMOkkVUDYaK6pZI08yc8EPeH
WawNX20SsEuomNlSlTQrqgtxGpDk7/4Ato7Oz5mrW4iSspeca6NyK26eppvGvcf7t/eOEpVU1Rq+
kH2mA712UozSBJHNYs07T1QSRiMsWneZVco+PY+Xhlr2VpqGW0crWx4SSsmH7ynkEB/LI5GChLKN
GyT55d65qPgrIUXXmr7Co65iM6f0jSG6u8oxStbNSrHYbKTdBIF7AxWCjajtuFdX2MM+6Z2EFCEm
CKhWIfnyByNdBujU1VTT9hNPHBHQ/AK9TBY0pxg/at7y0mCnRfr6FsQZk5pBkXQdVE3PKQ3T3X1e
holyEpvVAgDJhen+VHbUKcd+1p4q2K+xiSZJJVhFI4L8D/aHnVp4u9XtBiQ7WrUpvuOa0Y/rXy3i
zb58V6FzPvGkq8pHYoxF+Q9x1Pt/HMddDQNNeb9JjDPfoBqaLL+lcH33kT+SBmFnygzjItzhh8BD
rbKuEoN9wXDaU6CuHK7pJkHKlLZe9AELdmpxZiiJCUqt9BeXcDuWAM8ueB8b6c+KKcjz3H8eLma6
hj+5AM/3MCCx7I06bQmltSBhJmiwbTDlXEOFCUzlr0VCzFW8VouhD/ju/o3wE1DFJ2E+VMbICkMT
bqo4rMp3KVHNjky95lefegoQl2aDOCi+IOjq62fgtg7sApW8JZ/c805oRHkz4YwiykfwaGraDLX7
bTo3sWyWAx/slghOK4dt8lQ0U9GmZiyORCmFMCQqk489Zj+9uy9jdNS6yO5x4T1Yf2L3L8yzTV4+
eu2AZ1sp4r+gpEAu8s/dY11j6+PObM/4cgX16q+Nrf6DY/HeiatX4PeQKGmlnj8kcjHfk7UqpdjY
ACU92LDrLatemy0BeLilven8ynkluoAgRGH0i9bPPoln1zPSizLbeQAMQ/vVU7adfFjEw6/g0rHq
raNbxpoUDgHdss3qte14xr5AKNRihgKSi2Hsb18/iyhbsa07SY39I+JtDLQDq5VhjIPazguvfGw2
BRKQYGdu9bXM/mM5flmSI+y2xFup/dxPJA6i4LXPXxqjA6dhhRflfqzNDC5uJDtdI2h7g0MyqHzb
uJLtBSBvn5wlVPOwAkCgH1r0JW5Q4CHh5xu8HLlrUnWN15JMTRo4vWp34kKeDrzQVRZiWvvS7Xb1
9S/2UdxNffJoFkvdA8OovqLy551Nu/zCTBLZ3qEFSGkgVeuWTnwpYxJy5vx+r8mD86Q1RBabVFhV
V2jx5+m8H8nQl/LEHiRz93fdrBc0o9fDtdTErXbh8VxZPZUvO+URgGW7R+jdJBnFqYVNq6dtAKXs
q5VB+iZklCQPV4JlZsfofawRPQHL/2SHDEPC6r4ul9DULyWlw9DjQMnYhj5zGmIgJDS9kjyzzxl3
tnTUkueaxC9C+cHG/vm3athkhVBnRMTzIWtSVujugU91FoS6pV9ac+4FPMc8FJ2WmKId9beVizdK
LolXyRL8+zccs3H0K9NQyNed6VYsNc0/36XiKCr0cfMzjEwEwmZ+DlD6PG9GWzWdRTtYBK0RAgmw
OxUYr4k7Kkre0oBxX3BbZeZI4Vjn5hC7XaFczR3mq09/t93yl0ACojCtZlxcuv33YwCh/XXJEXa7
LEbm+8mw02olUFnpW8G9Uc+zT4EcQp3MR3DnOyc0n0a91wNp6RU2GPokXt5KesoWFpNMsTMNFmHH
8x0+stiUCuLFtrzh7OWT/lVWKGABEhTSAQw9BS4snt/lrgVYSBbIGmncFIeEgL5iWQioi1S21/OD
6kQ1t3ECy32wJ3gWXNcLddW1ADW1NJWv12cuVurx0wJCYVICTL75q+dUni1vj3xhFLyfe/KbJgwE
eP1+Aseh81tayHuYamff+3NKAxG08e0gQdxj4verHQMrQQzP56Ja7/LD/GhXXuCSL1LqMj7EGp5H
zL57gD5a3V+aoj9taUbRN+aoEaMnePqqqOR1Tg5G0RFVnJOUZhx6J7+cW4xyz0jMFusD7bFziQQE
PS3KsK+XSsLZAO06tA33a5L2ZvTSH0XQJIitMg/Dn1d13W1tUmG8hu7HrH6ypBVfczqp+jmLw45H
aCe6VYahBEVp52cj8IGcj93BbKGPQou/nR1Jrh4qN0Zo0t88m1kmhcdlBDIHlZOVYlH92fkmIwWJ
hbR5jh6wBPlHO+1Ejw2xQ/2ZiFBi4PoJHyepyLaxNhWeL+XoVOmmakAXesAUq4AIIMSo1VOCtc3F
w7jQ6OYZ/0T+HONIIVIg5WmzsrpwE+W5LBH8pR0YF/blaixz36xxQuNezFBbXu8WZTjIWSn/SeuW
RgLEvw5Il/ADvp8W7v1hDzWu42w12nu9RgW1LxdI4Iol4GRDH/oxTY7nFXsxzVS46PJHgeBLRIWG
z07nfQmHc35p1cGplVddNc6Idk9nrdGt81qWAcfvWIJlLtjUoEU+DLC7yAWsEWEyOAXnSyux5aw+
3kCXRaCkzWiByANHWu0VNVgR/iGnI0eutejIPCwgg1HWYotQuylO8DdTbBy6Igh7Fffd4H7AGH/b
cIsN+G+DDR9RYpop7NckfxYWUVOesHodqJQnRnt2Odvyn+KTHGlgtbT4a5PbtHvUMG/ltWYavU4q
rWb0hTCSLHMaFljY5qWztKBMfCWEaZWVR2AY5Pe5lCXpIwo1Tip+yncN9qj+LvSSnRhRRQjypgh5
0Cai2YN0N4L0wL7LOJNwxA6XAbcpfs+naet3k7j3G5sEHUu03rWXkcPIbufAR+pTymfx4GvUu+kd
qZ46S5m+cfN4JzLiGutqzsvEl+a1jJQ1PU/FiIDTCRNrPqj0PnvAloaILy/y6vnfewfFLlTR3dO4
Ftnyq5yNB+ErxZwLvIhv+QbVHSqjvhbumfQNkH3FEweUyYIk6+X8keXe0kTAo2R3gEypfrbLzslk
Siv/MTKENFYL2vk1tpX2Zcj0DohyOR7gMM72bFsBKHtqwgp9bpGAMrrECtYbah/HlFRdP2yB34Am
NGWSYwBGgUBjVpViLWm055f3D5FcdYsFd8XfSaAShP5OyAdfdZ2X7yrJfclvxNhKWxAEVrbWlVot
zemASJk4r0zZ5qjGvDjvZg5wmogT4mcHtqFxa1LuP5nx1rnotsXAOmfYAjqYqGW3D+ZKd7uvcIMq
CxWelx2kmAVX5G7rfrvhQRhD0KBorbJhyXZiE1jOMkERvhBQv70+OCoVuSXFu6b38192dbiEPZQo
zP6ipkKWwWbf/xPEGiMuVvyeuw1o0hGSyjdt23UoTBO/3EqJomresfQ70fRte6alUwmykl4RE7B2
/eo4hMLAdAPDO4z2v3o4N4q046z8kTM3KPtPj47fjDY8KhhLBPF9osrp+bBFuGpfFSKKTamZTs64
P7DTyo+US4bmVdAkWwsz4kVDZGrFxO4sPS/6IEHGsuSm05fQX+u310DZewK/LIEV3sHLdYb4KLyW
ZkIQsmVsjA51NgSU9Hw1Y90e86j7n7UM58ZoVgrdsfVt3299CxPpMK4z0OiIW/gUS05HarExejBq
mECnG0Hj1/OoLM2SF8GIAwu6fw8wLqSY7mM2Z6qUNU/2wjYlpeWZS1M3RtaSSU7uPya/FmI9Um6r
cgYrRXqlT+cgxdUCFzZIOsmk5WaYeEWvhomOBCJbZod0HyGVYG8K364BStoU6TEqIOBuE6VtOLij
JUH9TttTIOGbhG5htI/zttGUGizU6//DJetyyo7GrqIpx7FgkOpy5lyrIoxEygypqKdqXw8vpem9
yQBi+PbXOutw9InuuNXatPF527IqjaK862n1aR7YekqBMp7ksQ4/WIBuX8GT884DVmNin21CHlqk
0Wk8gY0lW8nfNwMlsTKYUFGUIA616lCQDgGNGJGXgGQGCt3jGcZPZXr+lI+B4tyC5xafI3mS5Zs5
Sl/bkLBh8dI3tshscWBz4q508Eyp8AwLTQYOmhMnV7H2HkTz1b8lWROeoLQu4eX/mlM0vE3KNoXM
/TYUh2tTgUTotOgPVdvA5O2w567Ck/mxf/6a5KVYFXqrcPtFtUD4tmkB64ukubwhympD3/kqlBLX
72XArhJpYhDEsIpoBrZLIJH/z9Dvobf1YYcrQYThgiiQtw0uT0eRDIYJY8cFP+fhTSJtzO99YZ2W
4LFFNVQr2gwxSMdZGvBXJof5P60owNyGgzmv4vM7z45CWygCTWnDU+MwwWu3BDjxo8PVckai+fGb
AJuPErZITLh4oRvK7ms37eYIVPhYQNeBEuh3wRuDJN1ByySH5ZIarYhyFrRegcf3RHolTlnxM4oj
84Sr05EH+ehOzFimXYzVtcmyFX94un/caTW9AfVoh+hfD0HoOHggP+460yyAaXCjb+9q+pgYiFd7
7xbbjzsANqplYqFzug2pQTyMEZbYsDGJGQzyhb0yWWHdidmzKTmqWQro6az9CzOnAkX7MwtcrKH+
MyQ0ghBm6SixHAjaWe5N6cUtJY301pRbSBFDBQdC8KBGWMnXdfesLiSw6sBIfsK28ceHkIyhwX1E
tjk+WBPweG5l/N06NaWoTf0ZQWbk7HQ/of8fVVEt5K32WTbO0uh43R5k4T6LROtS3rOtzw9cw9kq
XwkYqYVfoHYuaqLA4g+8QdS/M/jpWET5cgQeY3EoUTlD/rr1PA17xOpy3/OWxMMMzQ/E4LX8VXsN
dTd+tw9qArDptNGb+L8fKTYsxhnIlwRqxlj4ql/959P9Az55+bKlO3YzlG0cJy9Zd5hOgif6jRJe
8o5J3rPLhi/62gd3zlOCZjZrQV9e2gBaTpsRXJVSvhpeuQth8VLF58AGKQfGZRadp5+ogMJOSJKv
iiyIvKUXUUlRAo6gynojAW32VBBVi5p5EyBGRF68pj00OziqEO4x4LAAq5MZS0fObkejqoQwaEVo
eKYpRnftIG6E/4bILZPetmQ03VarVYceLE/rglcXyaGJlyo/D1v9LO9dcgUg8PHrnSie9CDdrmrG
32w+MekrfsmvgBs1owT1V2p1NSQtYRRCmhlWtNqat/0PPxvWIfI4dWLIJ+s2I//Y9qtrmerX64lS
eFC3T7499qox0uL+XQjQGu4HJe49DtiZvjPOgW+Ct67v7xilRr+piAkKI1dBKcHMHt8a9vUD/4rL
S/JFoOihOlbV2isxiWhput1uU/UN7AWRyAIuGYtg/WE/y9mVWus0nC4B+M21oYwaQyKCglkVUL6V
ORLAYUgKWxuJl24SUZs4BkN2fEQDK0z5diIHjU6yCWOL3EmXXePHcWLtg1kddijK2ct+fcxKQi+8
VwA80MxfFpDW6neE3rzkKh2diORlffI1VFi5LtFsic7l7WWOuAeNAEUVP5LJbPK40gX0kOLU9Kqe
zra86/4lSPYvKKA2EaSVS71Ic+ab0gTQRsRAswTswNrFmQoFIq8/t01ZSvi3JC+PAp+BMNr4OYBh
nU3tH9hvTA/lDagoOs/EUHFF9tMOkhVtBN4nibTYllvaSBq+T6U3iudjbqZaLXB3tViSCLqGb6v7
A98P3TBAAeWRn54pkSRmQpc4xkEZVG8l9w2ahL8NqqsV6pgcMCVKMxgE5XNFmZDQgUxxzlputtcM
lxeHd7VyM9pc6tOYYhKduPNFhHfeR/UyEsGI93Fy3ZYF7vbPnLCMZkwUw1rN08rrsdMGZOdv2uos
v/gMV0dAAqVjOwL4WpxXzAjHxS6aTfH0SWCfWdeJxuyxf8BNqUEuHzDSVOqypU6maM6SBkIol2VU
EKXAbpFnr8v9+oh3UMaUiTE65J20vg8UeyjDqN1kYUssWqIeYvKlUbWTNMK6LaHQ5f6UofXE8fiQ
jdryuNH5HigrK8bYY30dAIVEXtKex3uNL+zG5EVtrYsZ4KdsFDluN+y/ljTm8hkO+Gp9IdH7fH4a
OnPG1CajyErgp1PD7mTDSTvFKXEXBheSP5qJigchZBovfEwXuQLipT+2yNDqiZrZ2kyCSrEKY0r0
z9NaEWrNA/Ri/Sg3XU1iqrrArdItjItwPwlnTLnEIVXhPeJS38L0QdE9c0hbscD46crmnWNOA9YV
JVOJh+DjbP5Zg9wp1hHIKSC4z+F5fQoFOxunUlAWfeVWSmlvsA/ZLiI72PeoL/ByBFE6GX/uLtK1
9VR05I6BELGhoxWu8J7Mr4E9aJwWI35h6NDtDzaHWD+OzEyUDlyPeUGyGG32ugFrIF6R6ibZko+b
hhmZNNbxtm/qSqU5EpeU5mVfweGbFslB441YfFoY7TblKXrDT1wNrEaLpV9fvqbywolgFOUAXa8q
kbrm2UzHlUg3P9jkVrb9HKYdJVYZ16TdBjFVgtMGgbZHIse6e7ve7/gLqdkf41sAyWGcwukr4yHd
APpNNqTnjY3oolF0A6NO4jxL6ZmQLO978ei189YlcwmFe7gF1ILn/fmktMepAXEHQCrvS1UKhVe5
xX8Mzll/w73jgbCzmCFIi/ufghykrm73cwYMKb1Qatn80IgegvzBdZH1ewBk6cPl2V06EVgZi1qN
wfDwG9XTzQxuUSYpd5VGNTIbxVXZZr+OuPHu7Y9NCFqyvLfqInLktw3xnTKZY1fLW+hmeDLhzs32
cM3sUTq2E8pVr8AJ7IevtktZW5IVAHQtoBt5oZxHHaoaEP1vqddEt+Vj2R38OElRGeejHZ+t3KNa
b3gQk1WscqDpR/qie9Qbk/S8RajMsXPW91s6Yd1/N4gQVJzfI9RtFGP9fN2N9K0mhqS7VfO1z69R
xuuw2cmQgZ1fiB5tDNFl9Hp4cXcc+KNRDX1MWnWSwn4UNAyiv+dq1U9Q0fE04CBE+SqL7cZxZrgE
uUQB/z2HpmUBuZuIivzjzjh3KV/g6DEjeUIlDgmjPaw4PtLpsPlUGGM9ChbkFgkCe8vddf1KuHfa
NO2Vazox4zIhTCsNGnzBqlo6emVO9rWIui/A8SRh3iNUrDYJrd3KDnNwkMv7T5uJrtRSQx5FJFkD
n8XySk5fl7JHryOkq4nnpcaUdk8KDzKGcpFDf4CeqLMDmBEWFNjzOxdD9SN0sn77Q2EviMlL55gf
ccrWM/HEM6HgDn99kNKWp4OWoBogRx5d11ZkN6GXPloxTa3uR9GN8MzF/VXapDy0fgCovcsmTqiW
OKz4TWml3mv/0E9ggCE+P/U/MRKTBXDG20FTnwN/Q/pfoD3/qVWbGV+uWLhD6NIbLJ5IFbePlLx+
wJlV3IqM8lcUSTO3dhstuC99ELqOek8nDCRcpZ5bl44TU3k7N5ear6tMfu/aZME1uqaa2CUpF0ND
b7qoozfuXmVDnd5vbyETu75fLjjIoq/NhIEJbEAMCTbKRHse9TIX0R3cawgCJlrio4KvFZnNhfpq
ouwMaoF3Xr3KcKzCzm8gOwOypNsAHj9l1oWo5z7N2AGgReQRAfOTP0PhcnOK7ywTzsgjSCYHYNXf
UiOO0boXH/tTX02y8A8VvcDJ5k2Gv6tMVCdRgPp+naUjoDiiPAAvvW0YzemF/sQ+LG/9izF85eDW
JBkErO7DtVu+nEDe8olfu01/Wj86n8LfxAo/YVBFI1aKexuzkCOrmait2Fe1CzalK8LbHfknt4nI
MNc/DuyN+MW9XK4LBQm/R6P0FR/xWEXS7H0Er8z11kf0Z3ldXP1qjr5tUkJYQJevrtjxpPc690sU
zZr8Q4pWW/UT9ZLh984hcfK4UIR51xCq3ONQOF98oQvyxXffy6HDWz8s6D0CDuTctKJDAmC6b4Jv
oS60d/EjlkrEOpaU/MzCCV135uJe1qMqnXo0g8G267hajXi9Y1IUIpoG/LmTROqGX8CK4vVuDI65
pzTFdxNYVpSx618/KZH59wjNerFKFse0OpncAMw/ChdC9z8e9vAIH8qGgiXs4x60Kg9MNU9XsGb3
hs0Q2Q5lCsGNe66l1NVRzm+7ZB/hb9Y++1uIDkbCtiynxroqBSQdmc1sDrlDybQ/p9qi405GbDoX
jLJkRV+OoH6n6wuHqV73vFelwgSoLTs1CvcaM0+GY7ObDWkBV1FjVfaWB/tl5WiXRDvJTgc4bfQC
0ef7sFZnsZkAZkv0ycp5fZ4pi0akS92M16Dn1toUKmy8ekY5IGTBM9oFOSlHoNs3AXSyIfwXDTyK
3U5LuHttTcddD6EIIqbpqV3Z7SWvzCqNuybDOaMgOVh3RUOlHREVuzPm05m1c3YqZknc/O7WhxC3
3QaPDBAGOEu5kLAfiIaF+3WGlESdUyIh7pIR1d4UHrlnqpnOe0cy22Dqlu59C+UOC0Vnt4AO2I1W
PNpUEDFwotWFcJdGHh6/VfHh6mmj0/lvwoaR4C/18FTlOedpDLgsv6O1zzsKj40MrYelyLa8L1lI
nF2FXflplMs4oRRNY9j6/Bzz/Wn/HStMtyGzgxB61zi7eRF54K8RLf+umNoWqye9witp7hn49mpZ
xYgpk9Z9HS6mlzDg6jpknT+ac+qhdao24/dPLxfleU0q2AxB8OXftpGyzfibsBc2wF2VHBLqR18j
yKghHHQ+d19vQYHPcCYm/EogRWA0Jm+lQQK/en5mrl8nRX/HZPuxDRSAh87xsXftMWwdrZHE8QW5
R7Ybny4EoAc12suTafBYCUUeZLPRyz04E/Vg6JT085zpsi9TTZ64ACrdTurgR3W38wEJLHqgv9c1
hn8g4QtXqEoEYl0pW3XsgzEKJ19PbMq1QggqjM3pOaEh/yQvRDlC8TIor2RqZTnZwSJQgYUCv6m6
dI1pMILVYFJH8y6D6NpDrvU++0xtVd+xnfJQUA7BKkWz8nr4W8NvNGEcdlt0Ba6USUmEOkalV95f
dDq4J7WtdGjq2t7Qqbqk62mCHlU2rzJ1kO87VLdXJgwG24AAMNHu1cPNz4QYq1E83pvQ++2hYs9x
nJXu0Vpa//sg6XrJ/9OvUGddc8s3XyqXMPZHB3cdSmXCbc22+mUfXe94nwDHL2khlb/22Ba/STeB
voA+SizOQeTOcK3ojKQKJKiXNqgg1NZ3XAVW28BP5U4HEk/EvCwhTYONbx5kBUphyC5CKS/6SiMz
2nEXMENSn0dshHVhjUu0RUOQO8XMgETqnHTFkPz/EdkW8AppeLoFJyPl0Zf1tGwPVfNc5Li5+dFn
afhEIxdSaYOHwyJYmgYQaaBAcL9Ww4tp4yiJtc7be+YroJMC7LCw8vuCRGEyrkAKdwqZrOo6+er8
w8eJg6IDD1pweXGQy1cPv9ztsZ79PXV4MugH2PPa6ZLiPsmBk90B4sO/b01Svsn80eWzIQR+DPVn
2KLLxjfHYLAiVwWoW+xOrU/TjXOk+0fGW+ih5+AdPAYnKP6V9eC83HObXHvsEs+2dxLH+ojTdqJg
Wr+fCxJMOpnLA7bE9IRooIPytCpAzgIXMEFAz4TKKFEbDmFvqFXZ1xI2MRDoyaqDw3KoNWSIQRcb
kvaUmk0UVcwExo8PoTR/wwctym7BsX6XOFGNyHLu/LToqtjj9U79Jps8oPUckH4PYEiXuLQvKk6/
Jr6S5efEJ/D2AFSiJS7kDlQWWBJVz9FLPNXwKIzuHEk515TAUhHbrjeVY3amZc/Kcf3irq0y0lq3
lDWeckBHwJ/fEslwl4WAoDcemrXZKQO46naj0Zgbg5gR+ID74nkuRPt7fdmn26a+SQzTRxZxzxS8
cHzM3nh6giYy15TNJyqx4WGZM2wHkxAh13MJFo2Bn7LnQ7A52gQfZ32fT/1bYpT6FVu5W9+IgOF9
OuxthWbcupAM6E9x8s0L6Q1eDrDz60lmeERNVkyegjkjmlaZ3eRWlxtTmUEixRx/9yCSyCyKt5/+
DOQ0N6slFpcnD1D+WU9lg7yF4OMe4wNGyLn4YcpofYnbiZHfGaEpsaX9gIozxk8/4160TttPo0iF
OJE0wZPlT0uzm4QBN3FAbQuvfxjhdpDw8hB1EjmC80Kxr1D0QS737TVQgv1kVAyTup7AL7SdY24e
pClM3P5wAD+EujJgk9ZJHlWposhnhmbSYb8BcBBbnWkVme7PyUvDweLoHuiw7CE3ROTrw5Ndmqow
N8OJ0GB2bD/xpip3kbRlf4yEq9f1Z+pw3Wk/U+pjKsE3iSo1CZk6/2Iis4Q+1/9jKjbecag5XIIC
Padpx+nhxD95e/H78GCzOHR/fXzmIqfHPNJfU9lRDMk/w7TBg84/ifTUJENYE+xEwhKqlM1cg1Yj
1pZW4bvmYOP9m6N7Qurc4yjcX5PWT/C07EIL7X8vA/a7GM1U00u0TN5JM+bO4n2Fxd0I87wX87Ey
orinUfEvm/w/SsO0VV0+wRkKKRdOMXeE9AZxh3pktcdwBL51m4jghh9uiMPhCbXy2KAWy4Hw5dUC
HyPiQG0gFIGzxC+NE5uvCeoO7lMebjl1qYKA3VmbNKWezp2epfllNPzzttzEu+VebNmFDPQFmsVv
tL1TGst/X3Cr4ISz3ZWf6YZTAHWw2iviZxaWLQg1qU6qgS7nTbCEAwI5TaEHz0rki9y/uwdUdYq9
x8fEKQ+xj5U+sJRz0NJpxqO0jUPFeyAi8ZOiJoS9s/slq3AGe+6Xb6KwH0rsJcMhz/rDz1vf8VU1
Otouw7bjGUf34XWF1pKL43NekoNQVzjK7okc9LigRdOFxvD70Kt8El6cacV9e4cSaLK3B4PDhuvX
4E4V2pDIYTnY2IvjVMsbnsZS2S0+0ZHPTzKnRewyViQuUseaMYBKf5pQIgXQUYmhMaN4dsqVjNXx
greoxsD7Vjtxrn7Ae+RQmb0Lex7IYLGo2btLJNpxIk6BoAlPONZUi+h3ru+Wt4+ggamvLLbeCH50
zslcmrFdcCYGirJJaDlMmAXw9Vn8ewoX174d581atxprXO/jklJKcVh/8ujdUEsfb7Fw5yk+uCN9
vSM3ia+8TfCDQeZPwF0SBnwNowUpNuLtAzRXg6ws6k8gpLF6RGEBj7MK5el3CA/xq/iioW5GGTH2
xWMjswwwXQcGbkFENxysVMfJhkiPsvDPHZo3LN4+E3D2tM6Z/Z79EwdnZ2pc2JAtpA5xNaRppgxX
DuWZgmRyR4K1yBV/e4BPhdP5UOkovuGUtXTAU6VTiW/I/0TEttAjyoqZ7lvBRwKOGXhc2QKB6l7C
4nY8lAy5Ku8ruYu7J+bMSVjMKRZEcvOEf+mynY/pV88wlX1A9DzhlwQHc4OAV0e2qSDkKUqb26bg
9/xw9LNDmOIaJVvpCDsJ+kdqvhDi9Z/l8iAi0wjtf+AZQ8+d6dxmlJXRyI+3xLF56inonNvl+KI+
j2DfhjT2Modl1lUki0zZ4WVNx72nMRi5FcL+NXthLdInB0QWigLgMYEBLvEdHGHwgxE1m1VdAyvG
cM1AbLsl4VN5sdvOG4oxALanY6qDRNnAO1BZfjwARb9JIVR9feLif31WJg39LhmfsOp/E1FJM/lr
nhDwSMBXle01TZnankI+Z6kpeha1wuGRyc6Hwsgu1Tq0Q3lFpEF7eEP7rS39361R1tTO5Ch9Z7lF
BuhOpvWAhJcZwDuyaU0M++HwXsqZaUspfQTwYXz1nKQ1jjP8+Fcf5psRZyVN/dYoUg4kJgHYRPJD
1cLEU4H/ZI4EmLoz5Lq1E++YfJaQaXMQYaZogxhqCafZn++m28VeRjVaS9QxVbzoaw+TQpEyYTd3
oX3hWga2VV0KZSVQly0PRU6gntMvoC9hBTP5eh499lfGqsOJJCbh0fdZoo5Tx99AStASpI4K+13I
YywhXOEUjCZsFUEU5vJeTnZtIDrghiyDeSmCpc1vuhhkgM/63XQd9HphuddyXuM2MJvYejxZc+ew
YxidbpdxMFqItIdfWk03dptqrbvgU92paoLSIEOTmHanYB2Rq51JmI2f0WydBOQ8nEY5QJF5askH
8IT6MhGNGl56gJmCr0mAQm94TpLRUzahQfdc1PA/kLpYl8xapQs/R5KQZAgCmEAMWGfhDtZstYkl
KJwAur6byOz0U3Nza2sYdCGn/QT+qHCQciqf8niWKMvwhlLz29lbdN5QmlS5imqP0jR/XtVNk9Km
dhxRFpLy4/BtCMoS9qqUuFpRqjIxwNXEP5XC+9ar9FuK0OcmDcHlvuOkG0qOEIBgVWd9lpktNYqE
dd2/QronXo06sllzN2K8/0r7oKMyJhmYkaW2CS5UZIcXQCdTUKM8P/dA+edLW/Mb52Eb6pbaBtfS
VRhVlwy4+944HEbXBFbsfdfcMoORwJ7WuvrqMNAFhJKmVDVB297RkgsQDx5dMaHE71vFmkpGBOgj
lX1656nFnQDdkYFzaxcRF+7y2ew717TBgQtYh4Uo69Cd2NZ/kohzUfUL2VbhjLThUD3orzuM84Z1
gYe/LO8EEdJAJxcJvrg/y9jGTussugI7X9U11HkVOzJv+PfuQvt0d0lwwTL0djiUOmUfksSZoHrD
YtG7mbarMyQIMCNpch1tnaVC/JK//pVpXYe4A6LeQE22JyyoZZpVKKfo99qaZvMIuHfZEDYITAjX
bb8K04VhKGx2kn4JOofUiaWXOFhyJSFlcT/Y6cZevbuAZBJDlDi9FbL7ez3W2NBoC5fZEU3UBEDr
2LPxj3UAq+TgByaV9JcfAuTVAFk8lB0PGwoGFLCl+yCWx0WwznnBpKgrKecjzyMFt1O/fBfwtYf4
JkjWAZTX9JNN8nTPKa4rP0IiUGncbrROVxwHwUB2spGswByHXuCANFyrmiGXH+Q57ALcAr0lgNDv
Wjimy0kBPCm+8oQ2iqb706DXjc6x4lwA3iK8jEvfMv9p6z7GQ29yp7xlxgzgSDszr/t3Gv9nM+/t
/ym/VbDI3LzwFU18kElzEjpQDL7sRdfJau+JmZjgobNVDpqUDRoukjd6nRafdqqkDOvr4SWAVwqJ
Ll9+74ycpL6Eg9WV3bQSXlslMSk0zA8TuILeddrLT5bVWiX5Y4KeKgWQ9DGhc/iGhueRc6E2vVnM
Fwyo7719wzX4RSwUx7UF3+UlRmkn3bNYAtQ2OIXsPhT24dsr6U0o0lopx5XGz88MVXSFm9g1Eoyz
aZ/MhPubtkUtuAHNwKpveIniJyswvXP6Q6ds6LTCUXP24ONU18sfyGmM/dfmjY/gxp1gse3/Q4p+
VbMJLatoZvaXIuS2D1Uy1KnZpC8T6W3bRo37QnS/hprtQaFRi0M+H5vL2qO+9Uk4zLuhYLX7MQdA
oHx06Nc1VOJCRIjzWuCL0YYPYjeqEuhvH9x2WCy23QLpTCq0N8jYbZbUDBd1TMJdKCRYc+fnAqzV
iNhsVONM5wxuuraSVOh1aig+7Et/mEOGGc6yaJX6jVWMuyt/ne3DA4UYPXe8qni3Tr0xrOBomDG/
aDO93N9iyhJPGNnJ/xboRN048UrBq7uDkIOsimJhzeyrtHSx8KZ8mR5Zj2V1THDaK2fxPiEJtUIS
kdF13DK5FYCdqbOtohuTxr6IfvHe4Xq/EysH1f7edn8wBO1KORkwoKWABrUKy3wUcV84/c6l6tHF
iN1Acs82sh7wT1JqHOz2sSx/UtDLK/bX+esZFbqIyDl+v4PqexH+zkiEPsMMwJzmYtDww4gmwI/l
o5ClNZooW1BKBKqBdDH0aw0xVetie5GKSPp/hBlAKJbOueKOGT2O+ResvIdYbxDhuLbi+zsbPvjT
P6Z6o2r8PrXV9HWeCevhFRHzodmEwL1rMTIpyBrLFTgQMaA6ZKNDfHB+VaVMowVDt+hRJnlVGeUZ
rl8xgFUwU61BK/tTz+gsQKLCYrWsrVfYl18IJH69Jy+ec7umSbJmeKEf1A5ltNqa3ODudxCsYGBg
RNe00GUlqU3zlIY/J0n8YX1kMwNk7oRJcGo0CkEMsxAKclyknoiYw96BUT2CdwsBaankhy0NB6tL
g0SHNAlS0EHMl9EznF8UgnxO7D3aC4ErhPCwFWuTre2x0Oi47FEtrCoQHNvntzJDeLdrGVgqE0Kv
Ar4LZsm6IF022Z6urF3MGN/q7ZEvGTd8UARPpCeO6ZFodMx9mNc8+JLBQLOF6GffaoNx/iXtB1Q/
L4umT4cnwHwmtSSASPQlW7PA3Z+EmiBivqosHL3uiApQrbTyGkxSWceNZjvOVMHiHuGW4Dn6NuSw
tLVTHlyiR5iVFJd4WRXlxj2/hjUG/zJmnhCRD8OtHAWIYoBEhuSEGF6QPd23cAHU1d915z/74Dz9
3Xm1RjotWw5VsfvZ2CKiOjohH7+AawIWu1W/znWn0AZQ3BVUqE0q2cDf6uvUtgra+mH36J/DxEaE
p97S3bJfMdRJxQAwXvJhyKt/lk5BgyvBw3qK32TWkM+aBYJYgsZN0slqyHqLsyI1iRKQAsndl987
9b3Uy8cVvtogfApRI7IBtPlA2BW73Uz+bnkQKy6zFmBCDiy3gQd6q68oSFyRlGt267mTmhYt5APC
XhoE62nXTXPFSD8mtZkA/BfcKEB4VndgXFt2+aNWQ2MY0Sby9GqXlOP5udIJNHxMsdCHRWCeSa7/
ai1+SiwhDBMFgNfM7HXb+s6iir6g496ZyQLAByRprRfros49EFVCo9gmtcrF3EykRYZKytLvhfBu
sXDEFjuXF4KpoZPVXeMuH9fyG5Sa9OgVhnn3asxHYlxsd8vn/xG365ZDytKwJvKRy0FkMucD3t+S
T8PpsDVmDzs293dYGHQox0YWvC4HBL6VYF+A0DHV2v2daL6UH5w/HsBAf4mzGEHY3W+qey25KfRX
EhaXuqkDZHPOgvaEw6KMSJFSyzxBshwbUOhudq9B9y0q8Dj8tZ5G97gbwmrRv4f295ZtGB3IVj6w
3LHgM8OtZqwz7p30bviBKzLal75u61yeOZdfhvr/3S4hVRoG+mNEQ464iiHlJIKkUjjljQjEns0T
yTiydPQv+k5eiBJuk5SfF7yz6JTLgd2VqH9kslaZYcNCDs9NWxifXgBfRGUOFwwlnZ1loXqV860B
IY+I6DU3+Kc8VfdnatikrZ8vMrJ5ju+RJcFwrwsZ3R+YQmd9AuvfX3JCn8KfOzNJtvmQRjAQPcqB
ip6EAUX2S+rZf/Rznl1aw+H7q5OaD7+wxhf6Zgh8UI5hn3n73hBLT7rx7sy3MzjYQRNvrauWhoEq
CGAt9/Q21T690ytvKMzFI08p8Eh6m07cBCjRZVy50vc43Sg/8r3bjqDlx5mTUVpGIE7is5C3WufM
l+wpN/gd+o7Qv8/wvjOnBY8Re4/0JwXlJOOsW8IOD38cVuJv84Yqs0bzS5mfird0WQj58zFFJGba
cwJ8dk6rcfdc98FbK0a50+tzQRhKqkBNpTA03UFusOm11H7ZfhkVrjb+2yU7BcIa7DrEd6M6Al/O
xJlbXfD8+2wGYd6ye+3okz7H8nPmXER5rv5G1UfTrRwBjne48gEJyqApQqMEvIybVtGRmZ7mVem2
eOxO/ioaYnXXuQ9ba54b2BsB1OBwna/oxYZmfgCRYTCO8GRVhgkD7g2amALKx8VHGHjiXwJW94kh
V00b0BODFX15pijei36QacP9H1wbMtxo3jLWYYuDrez0kxEAUPKPobsGg84VjM7H/t0EOuhpn6J2
dkHGemFejoDs6TEIbHaZAyqvRPfYE1t/Ws1lTPGRXWSlkPLCPQFgAoobL+nJ/ic+oXmmHtIhTMAA
yPbyRQxEijKb53tw8YKumYqlGkcGhZMeX8UuS6C/CFoXHAkiLaHAmETISstEAEOzp/Jb/87CErOI
qymdrlHvkh0aAm6/0CQOTQuSNB/GD5nsX10gqkAuKpLnBI7cC1yvBCtatygsuHF3F5mEeNiEjSco
8JMDx6P/bS5tnYTMNXdx3SHbu5Z5+b+PDiL12s1Zd4pqAoFxPuVdGTPVjUHOW7ycXC9CVX1D0+wt
fPFUSrmyO2x3YFhIDWfMjtXIFVBMI7c3vVzmxpCJnONcXGyj23LTrsEdLXtxBe2H75wx2zQ03DCM
rqsTYiFkr0DkBNjRMOkYY0z0j8m84c7NKJppJNirSDPItZAWqYFuvV3RvHE4DbQZw4Nz30QrLkWk
jESDVznUTHcnL78qBZcWgAmaIqigzT63jV1DMu2jUj8wtOkTtK3R6RqkCzJVBMiT4GhVESbntcEA
PFcyHpwkrfiqMwaZ4tx9+mm6rk2t17aYpCyZnHjWqonZJ0jRj9Hg4XVA/cGmwk9JWp20zOWC8WW8
nO3kBasl5hCzFx/HdVIgqMuJ1aWLdEKqJMR+PQCKlPo5zAMgUOCDRVEod4U4Unt6BR2t7y6E9MRp
E0diJ1p+nd2yR0vjHCUJVQdypA8G/uo+MKKP0lI4B+WbTIb7eQui6d9kPBMCMoMTEfuyt/kQPj4r
1UNzKHBj6Vb24Nok4Jn3teJuu5hf2lmqfMBLma3rwwWkvfe0hlah31sqIhnXHWiEqrfcoM1u4Kl8
d7BSSkyLJ0mxfHSvR7kl4rLWa7cJ/LdypPokjBqSu4yraEnxaMG8M5/vkGXPN7H1Tniok/1RxGIG
vZSUt0k/z1aKVRDjBCbrgjJchtsJYkNA69R9xCDloHjBc10IrUuxDVhNvdadD6cw97krIsvGG5Oq
w/UCFrctt3h9PNmc/poNA7IleVYRXwIpornQj9dtp5f5J6iUjQLFBsrMAvjDVkaVDw1tz8qZyclK
IjMaatPjnFyQH+5ZpvOTOsAH8ci2KU7BXOkH9WS55DsqawjGNFHkzQGyWBjiM7ZvHQ8c1vF2zUe9
IBTSdhE0Hrr6PXe0OIXQOxCQXaPtrg7cb3njvqF6m/UHHF7nB8a2ZnrH7viD8r+O4drC/hRRbHwe
/OAtr3rTgVkS2pJz+oajHCTOPjoKIevkW1I5eFVwb8iSVlqB02hvjhxYFXkvtFAF071saVYzCQmq
JcGIOj3qKfVUKNudySDfESB6IGO5WHCiL5e2UJqbMXRE3unmdtTp7S+ieH2r9IMh5z//pwVgiHNJ
Nbxm7LvD3/iIg90UzKIw61tCcNBVYP6jMSJ276zBv9dNjR5BxSn/JDwkWsPAx77Xl+HGSv/ysYWJ
g50LBgnrKf+b4alj7fLEC4lGU2eKPQwLag4CNZ8SZmS0UgyhHzxxbDk3A6bM14AHDr7pvDWi4hFB
9KR4j5vK9ehBmAFP1W+nadhAFOMAomZnAvMzsA0ASce1PYxnzpVNdm6C39mQKvzy3pbrV+/uLk8/
jkO0XPdd+w+DJamHedeOWe9vr3/ulvlP20BuSNWLMIyxPVbGMfNkO8vPDklKWgBfYg3KQWB5HU18
X18nAqtDj2XmRIDk3d8lFQR1me8T8Bcflu5HiNTmNicdwPeTlnTkMmy03l5vnoYIW0kvUAGER7QC
jkBnoc5yhrWCg8W87B29exMcnzFmiaJVaK0O5z5LNsLZe+3ATDhda73aQSBt3503iWrC3KTViLVU
/7sz7aHKaozNb79CzsGlxLY5ewDpQ580hw7GvXRHF6k1UjoFS6B/LFhaEQ6oHHjXWXoit74FgKSF
RSCVm4MHmQvkMjbtFBGyTjZEMzlLSC3c/FU94RPYZILU46HzFKS3xw75HSVQRQJFmPCI9+P6TJZY
qk8fKg1bWalZy+RaKpu0ksg23ohX7rDOaWj3ryMuACU4G42T23mo1+ABLIby2HZOoj/CgjksM2xI
X5RVoQIBHeeBRn6PIGpYITTJrC0PrTz7vXIXwtYfGydtAzOuowApZyX8qd+ZLr96+45oo9XFX/Ah
X7n3xRTIdkPDorGIMyin9Okb7O9pbhfoghFELakYC/JomHhZKDSk7w6lmHDkIyZyr1JLZM1ySr4N
rsfUQYTgPuY2Zo7sb3puEz5c1CHkIY254HCJtwHg5JxcAj82TUiFQxk6DIf110TJDD8UfM0uT/30
C4uEN1uVYjpcRLU+zgpJri2ycBAaEzI2uYBl+A5i2pzgO0TuT6PPPCpEAPMJIoVTyBGGP3mNcxLm
gzZzJonXL1dR48eEirsKZzYTpBqKF0QGiGRY+xeUv5dbMK+XSOIkJAinG8Xjns41w1cBUPVbp9j5
eM+Na952PKjdCdqdCIwwDeThJZSjdkAXDPEHv0tZyxDBacx9kXxHnV9XjkU6/BLEF4GqVELe4+jT
Jh15/JRLwdMChTgf3afaR0JWB7f+oSQyR5Z1HJQcKhXqZ2BWQoS04YSfDaf0GrerxSEc1P3LgkRd
aDClQdt3PyjWrwt/uMG0jE1ha0JIQ1O6PDMj8sSDCHAfVXUz4EHTySFtsrMptrvO2l/LGBYT7EY8
sXsG4wNvvGJGq5nEcKi/iogmSTc8eHkcEzxqLde3fhZqeus+/mfu333xSeX4zv80HzF5UCWnrNp4
4QMJuYZRH8tApEGjW0jmpD+ppCrN3ltqPe20w8Bp1qnONrn1lp9G9gZh+ZxpsInmBe42Kucin3Bl
NCm7yKm35tTc/aVZOJKsJfB/xHSfu/WgH7VuQDX0DQtGtycBtXWngnMo/41cOL7Qz7TygSawFtyT
jHrRieylOvi/0pCir6YbjSYcDLRFe/ep2EILAMH5/uhylKWV8vJSlMRLhdCSXodQk65HCaTg1Kb0
ZVmAnxqeNkLnurhStWKEbdMgUCCGQVcHBBS+VMzGSlM2jxSIjzsOw2vz13qlDQF4mgaPZLsmmPFQ
+u+PAEF7SJp5YF0O8llMztMyCSwtuLj/TBza+rMXJfE9aEaGeCGjZtriD5gi8TZz30hc9UXUStmw
1FzrJZs2DdOI3nLmnYTKHs11HgbzdSY5mRBBqIxRCekomTcmbH9N/ZzHco58xYMPr+52rZXqjvtn
c4kRYKY/thD5f+J8kdMDK4e3eUXzti2+OsrthB8o70NzpLSF2pSrzx62/aPdtO9ZCBpBqtIZxVXt
8TSjqSSxgCTUJn4mv+1y2TKmlrKc2/CzWBVSHO5XhoDnR8ubmoEE02pb3u6RfGcCITAhI/SokSYT
pczDyyfwLTX+bBJXHnFzbFc024baVlLPBmQZyZLQFPg/U3dHvWrUAm6bMFRRzA+RJWKaAoBFEMZS
q+AJXPkqednavCXT9Mnc/UBWrTp1QIRObGaR3rW9+xh0DDcCUtlzblUQUevKG+ro/soHkMouLB4l
74PJzKY26BuLWbRyv1Hqq57yulAx7Crl/1neALkDScjaTkwhWVeHuXJBL2nr7nk8M5H9q5oBgjju
fLuh40Q5pIRmG2B0Gan8yuqNejKDbI8+Vzleb95l+Y9DUQ+z5r6XuYEcRvNUr+pK0O+JP/agke5U
7Nq61KFDf7Msttbde9WTu56qy1uLez/iqdnQT+E7KDwZ+RbDI88bccjlFHUpDZcraPLCywwn0Y/a
zGre45SE28gOhITjFHUB8VMt9ZI2qPis9uhSDYB5THu+2AI87+crJ3D/Ai1SWE5vg2DGhvsA5Fni
bTHNz4zyuvticKctJ8pBHXvypVsfU456uDg9ckxyJgjBOeL3laDSezXpYWvb3exe5OB6iEsoy9IV
2VW8x/iYupz5PITV/tJQbrAM9TIFDB6PDLPxqMKEtLJ4iuIK/avu8fzBZbdBqF8vHQWpNc/n2cvZ
Ikcpne/Jfvy7QwKXolz1g8vV7rC63TbJJhqY/ym/50TiWiKjeyQ7iC/V0PMsoK7fZVQ24Y9WTx1Z
h9djq+iei3ugp4uqK8DnCauw+u9MFuG5nVDEppZsBp3D/qmcObLX5mudA5tApIOh741fZ+tqtzsA
3E34LyJJIbhfhibdQOLBNsQMrAKT4tE7IQOfvBqCDa4WiGKFmqPy3VNdVU9coYQObwXe0ml1PoAZ
jBE66OE6o83FLAYAl0A3LzRjonF8n+jTkz0+28X+T+SerCRfacE2G+AFf7o8JBJmamrJhvr8Y/4p
bozFawQ4G1tgQ2Wl7jHzWc/FAzavkX4sedvS6/88sZ4J64MKlVF5gp029SyJK3Hd9qHdGy5RUiKD
ddpnPnpOpagRLo+keJJKQosqmEoRwHzHwQWlA7Q05spDNydhBpbTXiPfS/PRUcnyIQoWOs1YCjTu
pA93dmh2mn7skm5uDlfohokknxL69bLiq/YGiaCt52ilOD9sNXJCHpCdz4FEkR3/30vxh3Ar0SY8
1Ehe6Bjkgo0kK5D/AuUU8q2t6RkhqZdWwPBD6LRVGqWXl8VgZY/0bZ/e5foZdgYUAqXwTSO36qqQ
Az0binrqs//tnfVydMLq330KqiPIxEAY34IIauCel6S69lG3SUFAEjcjYY0B1ztFWtJ7o6FDQNT8
cScoyuKQ1D/BPcMnUwJpgZ/jlufBPDeNYeVqOt/OBHEXYOIQ/5+Qtqlanu70daA4lVIC3LZZmTlB
6QWlBSKa3l9GAEBT2nqyG8dil2Yc9tzrLh3uZyUv4xFXJA9G2nTO253zeBAQPlxMQZF4OWw30eQa
kRKvO/y7HFgxljPD6jEWWc4QSzMLIsLhkHTQxPPFvK/J+Gx3AsI6Lpdn13G+1XDCfvrFofmxIelf
WrHqTrNqi1QLQoukUGZm8Ifg1o68jimvE7hBvr26kkfYF6vwEqXgaIjE4EOPJTGwdeYtak9ThxEv
YQxrSojFZZLVZ6NUdBxLG1N+gTIi25syeA/WexRaZDMu0W3gU+ALdB6AUyFY8RJdf9+ohsGwFjW1
RkygYXwyubZhx91C6lRR9bu7RCJqmd/3RgJEgnvwzlJUHOM1y8FDHPOF8m8uxGIXGpJTl7x93T79
IQ9cy9M/7GPDm4gpt0JxsvSMBXQWHaIlfbJ8ZGeiAg9GHHZdPVPky9IlLQVijPpDbb/FgE18r+FF
imYytPkx/FLxwN1sh0pQgPFyL9PCo9viAcVMpNE+hfr7QnzoYcLV1FUgQjNqKAJa4OaUNxqZeH75
lKwOhsiPsSSzY6tWM3YDWgGOuT86p31IoTHL/JJW1/zeKJEXru6m8zRIiqlIpenVDiJeNMwwEvgt
zJE1d9MBdzPvOlCGXXSmcDV+u6HTbssg39PVW8yHUEg4Kscr6DqZ6RL/gb5NHGOvoTYavxXf5LmI
/Sllwaxz1UXP8VvK8IA5zjbnUrbrMvY2uUXzTSFt4OSOYpEBQNCfP7NCMY62CPW9+nf0G9gWQQDa
92/BIzIpcbD/0P2J1YRrMWDAfe0yqKJ5WC4nbiqEF/Z1UqLuBWFcUC+6gbQorhRkTH7fLGC4Md6Y
4XtCaPiXSn3O1KFDulHCrl5O+ZmGwQHrnaGHl48loo4lmgbw5djZwimp3+s3yg3QlQ7ACR5LNeeV
acMxUoi87tx4YxDRfFdwbrVm0xlmpn3SoI4+4zm+hpI0msQeVwBKDpEn77q9EBjnxbWJnXnMdEmD
Tz71ZAdU/FrI22wQ6Lq2c741+tivytTZ0/nJifnHEZq/5egGdw80pAs5UkGziV3FZw+/Dz2p9jgE
e2vlDKCnRoiLfMRYCWKrcbbo5HDZ5bedVghfStD7hfugzW2m+im8hb/56Z1S4BRjzKGpdOUhfvno
/k1eNLL4rnCThCEE0SXGFF+3a+pcp9ikx7hRePncRHsr8ceH1f96AyjygYugixP4wfRsgEXywhEQ
X36hlCkThw7L3+1+Hq2NYtCcPG5QRimF9porMLKrHOekRJ8xps7EmVPCSIl7dkD8pU6PUjbI11Tj
adrZflvzDORvyB/Tb0tSoAsP8t0SBSjUvc7fexZ249r/h6PDc25cIjg7c30uTRynLUcFIo7rFwJO
H7qokXHjIpNhTv4dvBgy7CDrNoDLiTWps6BdkvSqFMO7ycjtAJ399FdEBCasZhrIV4T29Maf5yWn
01m/z+hv7Lb2+TUoqIUjVYH+SHHifqbHimb3fBjOJguPFpihR7VbFMwsoVUhhnw8RlXBz+6cFFij
Gsd/waFgcdbH0JKB3W1/ES45QVjo258burZhz2mnzmc2GZ2VwzdJqdSm+StfZstHxAurGVHTkmuF
Se9fIe5rkgHVNwZyNwPzDCh2jKU6H6VXkMr2mqr2zqj9b5zoq9/n6/8jMI7qauU8mP78+Z0Ry6GF
YVSqmo8sJ1ttfBUXwndlZ+xRIaUCCAlMlp44cd/0SsGdr+BKlM2NDHodk5exhHUJSCDy6uGFoiQw
ly1qk0QG4hYOHpNJ05ZMEAWsbC8I7BrQJi4Rqpf8XtcMCBsq+Jy7gjdOClFaxD4DUI/OgHU4ZIxy
8+ZzgBPn+0AIrZH0x6sCiC1/rY9BY/6eLv8bFzt96UnLSdJbUCf5034I20LD9bxmBFtuA6qbdYyM
+BdqMPyg5t6tvb750G9TnBYOn60MXWxaAZMhywixVj1+WecFDWHRWE7OrDNJ1jw1AKqGDDZi2VUy
s+vI17F6WIDIpJlduQCeaBrhck1yy99DuM2pqAL/yhvl4PGho9zpaPzlxs3LJhA9tELDfWSaFgsp
eI0zlAIVCiAPAh9pRQBA+IruGtLjcLve2XtPBJR77JVFmkn0aMoJ+m8czBAOKugVzX1sCW775MF2
ckJHOLBxgZR4IfXOdCZC/tA++mmuNbRV4RhQtGof2qSEmnZcN1CbjfKN5FyhXNBZtKobtubBcAPc
sygJT092X77dq/9TKh+d5319RqcOD9mD2yZ4u6dpK+jPOgOTNAxHRzpV6wWzrzLrgouzmpVxlrW8
wIBRVpdSJubtj4J7EkpulcWO2897qoHfz4CcpwoX+s7/gFncWmLQJgLMPtvQQde59E4nYfGkfCXi
Xv/n86EuDdSkDuX0rkDpJw/M1O1SMUsr+eYHKkpnwDbEw9yOh7reIAJ8A+nzt8Rh02cQkSObBIq6
TN+Ea1Hajw2D8YvOQCXxT/zmhYE9BTMk6PQKtI9x0z8BdejC15gBluHUFJ4l1IFw2rl5bUlmIL8m
gd9rGufEHww/pABrvwpgcQlSal28C4Oi4GvADHCJelOYAENlrHvLn078d4+fF29NgAOm3SK6JvvC
kGku9HXFJn9gFSV9bh1S+kyzJe7dKbdAAvf9XGtY0ugrBbZT9cWo+dzXCDHlTu27xr4aF8V/ULFc
2avVEUtvnB086ldRYKUEaj5ybovyzVulAzWBGOFnp2x0/wRpEoozCxhrzHWVcYIW9XSzqzCfHOe8
klhFi3hqoWLHaeZF4E18mUJgochQfAOkT57uLAdkeSq3ss29H4R2+6Wv9MBjkgEKY5awXkp7ga8V
y9lmIsVtuYb+G3qzlTVe4VWBbO0CUIm6WciW1ek0xVw9DMx5EFLEPcF8zU8GF7XJ8D4ew9FfQF/o
CqNCzY6QUggYDoE6E+CA+9k01EMhnwMfv93GZIXrLX2k7h0S1klpDAbWg7zFGr6AnahmfKL89FcZ
7G4XuMsgMVkSUthrWRI61E5wd1X7rXWHieko/4iorG2CxqwEWQYioPVzQBPNHh+hLs/7Fam/ONZB
KcPc0dH7mFzj/d9xkiD2dQn737ZdSmcP2ova32Az2mqa4uXDWWuTAdVFXnENHmlJo2kc/vsA2VHG
9oNxxXULEY35VLbZAbZXTw6VHtQpeSMsaSWzw6bRr1XZ+pa+9qZfkiQvgSkFZymP3hgA2t3KGHjq
2JH08zCz9c9xmvI8Q4zb371EDPZzAVzgWKzTuahFuD/Zj+cvhLWU+GkEm42zU002OMUCG5v2dLqp
cpAtRmISKgno/R2Slj5hmELulmAXpPc90FbtttyCRlx15/FtI0q4xW+HpZ/Rp3BEz+185grEFa8Z
ojkSQEKiqtu1B6QYa2jwZdBfcWPxUc34wWnRSODeAQmGD7IJn3KpCdFrWiXN8pDxJAwKJTY9rKbp
1FVaJk3zKGZRV36/f45Ddnf+nwiFCJNq9nVuw+4wOgL1Xz+l3IQMlKtl7AMxoCnxzOmmqj6C19uw
6zm+25kWvdJ83Q+o4jQkwTlU8NvlGWRwraLroHlbKEMzcI8pDmKfWq/3urQwbSMVmz8rPr60dmsq
FpfYTBQ88SkdHLlwEuQdOytjkzObEa3+q3obY8vz0ySMhiUpTmoCKxrp7zI+5sIpPdrEvkYDE1Xm
Y0qed2mjnR4ImOWWX/ZvWJNrAdNMTa+GH8gMnBoEuqKZDXRR93s9gC6MhmdTcJrh4Zptl2hL4+Rv
KS9Ckq10FKq70hXoG4b8ArW59xV+WtKbgEytzOAKaZuFcsdggYKz+mh8caHv7aBMSniFyn5y69yg
RhsDRyR16VbmQ2J3snaADqMjYoCuyNWU2zRgTrGFPNdQ0Dww3lSLUwtQVp+E53vT/j0tcnNMrkQ1
C0TPqQROFJganqztQxJzCrFJXtXBkvhxJzX2F7UT9rGJdrcNmEKm1Nk/pZlTwCP61UdAoO2LA5/3
GENn9Lf9jRgqlRmPwEiyF+vj3lK8JMtIe9hQ2qnJx2Ehli5tL6oCpHhiS9WCGi68afwUkngZrTxt
E3K/DNObo8vg1VyB6/BAGmWMHlz1A+7ksHgjh/D7l/d7tGxVcxCQYOsetJMVJlsDGOjfBeRtd0XD
xY8rLbkVEuocsW2JHyxO/kwwJPzZ9u4QIj710biAJzk3EQXQhD0O6xvfF9rm2SqDzuMsF56HkNRN
raNspWnvtD41BzyZKbDsIiwxeq43lLOEJ6UmMRGASRe144TJ+RsCNVZ/7a/JEBxxICQbrglGBoV7
jCD+nut3kYqAk3GXK05HbV5CIPHv5anIg70SuCx6IaSrhYkP4iMJP/rPO+i5zyuJKiEbOdUoXLdt
pa0W2+EVXwFcG324E014bji+OcnBptAfdgJvhbiSTxqd+33PPiCr2jO+plcDudf5KaVY65zYtqWw
gDhC8XczCyJJzNL5HJQtUB/l01vn0xoUHaf4eqV90bl6i9PMs2LPpIAgYeUkazm4UOpF3IwSQZSN
u1TPbhgcBiKiXIGoODsqyPjQFofYpE8JoB/LBkbQoPipM3koOQnUyKt/oAJq23DOe9Qy6RFV1Vtf
D+TO0o7kg+x1JMxJYk3DeD2HLVBUqJ1H8B1eGAbrvP6HnJkew9HsI9xL2cIpjp9mG/XepzZ6593t
GBl8DkIOGXxhbxEGOiYVWqTjw5vGgPbr6sNCkD+OPrXR7xn3KONuIZx6pgRYJF5sWNgzKoW9pjhu
uFpZf7kJWbq5/R8VFKL3UVH9+jA42LoLZvy/9hMCYVKCyh1T9vk3JNn1r5VtbhjthP5CBso2WSSN
OQnbcONuqPgbUF/8x8xlYU2xPhiRaOvLyKPtb70h0705RDMnani1hvdnC+gDtKxNvxYFbtrUcdHT
hOYBIzbMy3mVx2Lt/vR4JtQiU6E2RYpYXrPjAfJpzwRZHDLAjBTAsyRYbWZb0MaY1mp3RW4dXRLR
brnbF7Vaco3BBI7RR5SSUVb0/kwl98MVXPogxSDyNqPUFAhuR+l6+SuaasZhxJSMxAdEzsas+c09
HiqpdDs6g0bbKyQWIFAnJ/6G5QmshM1mOj3JFMBK9tSh4DBFET5JvdBlXb3JcZ+VLRjpoFyF3I/6
KyhKbR1XujKYdVWobA6cpIqQ3BEtba7LJKIk/6N4tJSu7Il9gqQcbvjuHDZYGryqpU/mEo5Zv/d8
qu6fcu4DIj94XEYyTTVDgflAklS//EcdAtrwBY7+syNI4vjzEzs7DSPOD1dyC9Dyio2R5PZanwva
7gJLHR8JevwVFHtk4iQrtshFGSlxQ+L4iU+pbVEnZJb3BGF+LFt7tCah87TBm6XUGTFM/uSThi1W
TEjNuCCb53xAoJ3hLJNhyxEXulm3gqh0nnxD8DjYtiYyMUwrLnVXGSp0A2LGhBXbmuNNkQy7feth
7F4i+Du/bCUZibehP0YhnPDAXL2ZXoU70qfxN55D125JDAURhemvzRZEou9Kx10VRhjpreAKKAUP
ONOzZrO+E73rMtjl4emwUQ8kHjB1qxdHOjVEKvXgqjcDC1ypJWQLgDQtOniM276dwXMHR2cUlmT/
COMNU/22I2IQpJDIa2ueB7HmUt21SB2eckqwu3BWXsll9CvYrMHccQvcEmNmERUjKHh335pMvMFJ
NZeQjR9lCGIUcM/85JRRNq6JblEZsZZTv97sYaMrDgketR1FZHdw849zsbJt3I1HGaIm8IAdjSgf
u6S5trbsMSRLgk0hTG6kBvLBB3tU6snIR+iD0z+iQ1uZPFOyjGYVviQ2sEs4Km8bCa0ilWSqYMRF
kN3/+Wo6tFRuT982tBAw8kfkNElXtYjSOBDMkxmnHWYyfe6rOP5GUSJPgh1++jLdilq0CeyjWexO
4n3aeqpqm018QATERICtITKRi9P5+uszEMUu3rNd0gZQ3rFs/P7sUUZg108ZhetBeZW9gO5gEsCT
RuD05G222xhoFGglEFxorFKplWPX2EjwkvCV7J8N3J06Mrv431RLy4OLu6DDELJff2+GKZ87k08R
BGphmc40LgCCWO7+jPwon/kwR/9sMSZXUGl6bidLrbINeL+XtOWw9m+EAIi0sBLT+byBF4CQrCr8
LTUX6stkQr7DxLqKjC3vcmlZpU5QfkE/7vL4cT1PQOq6eENIyNGRuCSr24L1ddXHWA7yD9bK/xa8
VZmh8P/FlKMjIU6k6mVeoPF14o9jFu7QKdgRN78W9AZzmTwAuSK0wiVb0r2QvWNOESCqYfqOg8HP
wQbfUmjs7671vT/yLYnhN5jAc1QIsRdfecJ+8GjkljOJEyetKybA5WSjR761HTYBk5vqK7xT8H8x
PZWN+RKJvNEBndHQxAvUuRDovV+E3Ha/Xe/MxVt7jyyrAK04Y9TUf1iTXXFrwD6IqqbL3lxUSueX
1KZiMKdXjyk0Y4cxHWp6gU9eb3YCtys0DR5baCA96bWxfYKoTPBkUHAW9F2xeimQKGlmX6PrcMkX
rAY9wk7wiDHXyW+yH0oHFRI95Vzz4egE7DUZhJwkJZPw9bY90zxjxYPA9l9ChqYbS8GIuPf0Curm
9HugC+aPKUkXtp8WOneQJrsv5QNY3dw9PfidO4s/BFinn+Jk16QMrAXv2fLyvAoWOOgvVgujOaWu
M6fW3EkqmVh6HI5Vqtu2FcmX+y0YZbzKKae6oZmhu9wwLIfwp/Fy8d0l5Kafd3XRPK2WX38MXt01
umCygpZOCioTm7llSAiVy63k9yI2HFl3A9vQIVq7nYCCY++jpctv1P62MyL1x5x/ZQ7rGv6AxpRV
tnKyIeJuwUtA8h8y4v6SjXp8fTWgc65UD+AqkhtVshAVGwX0L87wVKdT9+TdaisYlLN8D/OcUPbR
8ruv9AgeekxaaiOKvPhhaKPfhQzpKSWk4EBSLlwNt+C7baZxVVF/zB6xnfHS945e4ej+7YGpgm7A
MFgpW7FQdwrjeVFcHQEKvzaD2j+Pl7RAo57wO8A1+NZsRMtVEXGn/JsOSFIohnWz0f7boD5EEAZW
PxGA5dsIkKlpHoye4Tk2llYGS/T1pBNqGBP40VSpNIVuHqTbkCvLscvtPTnKLgFZRv7ELQZf/CdE
P+3VZjLaWyyF7OoH/uOwcgZRCo4ITxnbeSA0ImyBsq762F+1LTGZcFa6/oXoF77wwo/HneUR7Kg6
l95+cPXVv7U1uNZcGTgzWtS/U6Ju9k0PBdt4LVqMZqxp81nyvMO4n5gLTr1JzmrCQSNEJdgLk6lg
q5sRjBkICH+Syaa+7EbcdB8NtgllSeU4BcsYdhDQR7GmhtKN65wsq5hG8KCkL//y7ncwRGylnFPk
VU9VsHndeEnvozNm32cPHWkP9IoRVyjBiBk7n5dLD+M2C2rKkn2WglpBcc7DL4H513PB3jXqC2qA
Z4fC7JVlj3ykHiKuu6tINeTcv9PSMTrwTtIVTA0bRzzikidaOCVCOwUHpgOZZnUyapmVejN2SJbm
nJjqgsRXXdYnW00AarjwscMWOfpkKmh8pgFG9ck57q9JuM7AMnLy+B9Lq7J+1oRjeKJeTlIw9yFS
rboiRT/LW8T1Ks2768I+tMf0rv/ZCGjwFJdaDH+o10Ego3uSECfIbkfGHq6LEYyqi0uVYk4W1gAg
vCqNF3lj6JD7nLSF6Zrjva4PhSwzXhmQ1y0XvEMs8oDraQ2m81Wn2EsrKLTYt1OhQARFq+0+xq6a
e6ylVXqpnSjDoObT2A6P48PDjcFmJQOkRYv1R77QfnQSf1zBoY1JLgPI4BeyMDGWnMApJ1u2CmgD
HqGykSp14o3YqXRmxnAusssEtHXxsWuzxNJGXt0u10OYgBCJAQUv+LHqmDMDiEYMUxiA6v1BUMXM
qqOz2TqVZ3IWHQvTyL2rzlThdcTjnxxHDghs9pe5wtAkSunJGK6huN0b0z84Bu8qgro+6p7iwjOi
FiWG94Eg7+CN7abswO0maK1FikvviqLQVpcax6HLpelhMCeMP/PYJX4jNQr27iJDbolpusY5g6eh
+xtJRbdk2kf/PX1P6dA3a1Xa6aFNEhAkcZoGg7OFTLy7F4gCFo/RMpbHl4NBEoP8y73f+1WqhWbR
UASk9sAhwxWJPSZVZu1atzGtHCEt98XtgM4TvXT9yGN6VQz0LL8fNUvjPkqln/Qs2jjQu2AkUSmI
jPlzsns4QuXv11lZv80ODkt1bkN43RYGmC0kKy7V52C3WlZSUOlk0xX5teEJpt1vjJVTHCNeaQy2
J3XtH1WkBEgpZ5wuem24Jyjx59yGa4n4pbhSsZWNeFJCtxSQfddojrg4v362jSnJ0bZJUlemJVle
TUYlCfr54DAvdIJympn/yNq/h3qq0y68eSWNrDPcvbBEeKkkxDNpkyJ+k5IuQGpLcYs+H4MhDKRx
/ms93BgNOuBh3pvxd4s+yVMkscmOK8UCROxcM+gTIjqTB0Pvp5rYDxBHUEVJExr6CRr1ThAfzpYt
eTo1YuKWpVnvlH4bPUoqAlEkLBmOO2yTOLBxmlwtBos8nAd3qN56q90NgPHpAae2H4Ql5NQcPFbd
QT7ylKUTi3ymVgfB+Ilt/+GTlFx5/IhECCps16Ccg8bQM5mm6Ei1y16RRIGmuE+p8KG/y3N8V9v8
L0U2Wdaz1Ak0Icf0OBdqzK5z7Q5PeRnOz/TvbJR8mRBLEC2sLl8YliNqtUbdgWjrJtjAUQ6eFGLs
qTACoaK9JCfZ8wo4Z1w54hb2PfefDiVpGms7adCmrsBJlYEExAi5M0Lq+eXLrxFM4Px1YTl5w7Jw
IGCBJ0pzXCXFdMCzDHwlUzJfnIeW9XTUiPyC2e8ZvTr3GcOkwoyWoo9LTZzDSiui71sNh8xLrMn6
2jZTbxKl5aoT9r/ECjAPgTzFMjbZkAKOLbxPuKaZRb+NrP33dHAmoabvP9NzkFJWIBNHlMJaBAc6
gMcZd+UyFaZmTTvaBK1/C5FOnOI9FSgic90QdS4WG+K4DrAhMEWWvG/5yfbXUJG0UeE9DOmmrlRC
P4v0YsUWfDcXK78pVAJvALW8MILmxLHl5ZeNLI8lYbWD94AI1LzRoM6NLM8rFpCsQrStxV6NAUfD
L2eUE5eeJWVXyR8s3v3l1unHkQzrhLUagbyPb5nv7wyRsDshYB21qi9jQUfb8yN+m1XH4uXoNGk7
UyjdErhwoUA4snBibfSVqUrj8m+x1OScntJ3m0MxvaX0vKSgY7pTQ9L+jRvJRkstCuhVYs8aC9xl
t79qgAukqkTit8T82Hp8rf27KVh8tMpuSE23jRoILi1xfpbeF/ZFg7aUa3QlsP9+FLAN+klTjiD1
skQ/iCbT19KNo/0nYHxE4Yguk8U51R01fZfuMXiJTox82P0VFDVEj/K6XYXZBqfJ0MQbDL8iM6zV
9CzOpaJml9SOyjm4TiCL2S55apmn1TQ+ISDj21kxYn4AD1mcnx/OGHPiODK0wgUOWa6WV0Qi7TOv
YG9PjCr1jaTRg/w0MZQor1kfCYo1qkryTxeyQbsZf24kgsEdHTmNTNNOldss1jDlR2E/m8AflgzV
AsHufu6Lfj7gfqtq7Hr7L12rfdq23HM10rWYHestjz6cqUQZM0zykVo9eb6J0zfSQhXal/DxRkw7
f69/dTxfM6bjyDG3qYKYJCUaN3kneq7Dr4Mk3NDFTkNQxvNRYPUwZ30S503PkdUUWdeo+cwS6YQE
Xox7YqFBpnZ33On4miFe90oTBLPH/1PEROvzrjy0ncfufw4QsGviZfTQOUxn4fX9uXJipQazyls2
hOmxzGDbWCBsC/8E4jOelrv+UW4eHT5PcsLyqQTcQDcynyT394JKtw9j717Pq10H7pg72b5g7/BP
mSFrOhzTerOVUe5/kt3ekP2myvlLE1XzMrX7/rv7yzYdqXk8ZGv2cLfXEJMtkSztbyr0lcThT5QT
nWZZJYNJnrVaVkrqw4Rfvf9uDR6RRZxI26KHdfRfNnO372nhSLL/zcnHc2vxw5fB9NK4GPP3LiTw
2XIgvGr457YfrlD3v1zv+ESmNUrFjLgHnrno/99mWClZ4/2l9QDrTDj5kOf2I6g+VNXN3/zotfwy
9TcxDiYWYvyrfUvQ3zELUyiPu/Xg4KNa3ws8UrXDEuGHZ6rKJ0m6mx+W26o///AVwn1gvf+GYaA/
hPVgZRyA5mqNwTO8kvS/TLahWhzFYeNN+ovImkruJrqXAkIzD0SwEIjwHFNQgPCfSiS/a+FSgdKr
5muJirbJ2lEZADKk9v2om1DvoO9Kk2b20ybml6yvZLjhK8ywORE4l84ccf69ohJEXKL4DQwd+pWn
8RpQpRTljf7x726vuNTcXeVoJtDPAZjuhP9ISpTjh71FxmMEGWFRef290D5WvAoLO+nvaqbePONd
k4x0xBht9WCqjkQSHBfFv7/C+v9JqK4P6djUxNS5IZOsGPnQRLz6cUk6Xv0QNB9BWURE30Nqq8Kv
UODlCoWTw8e/aICiR97ZgQf9iZ2ZyiXqhbBi+1Ni/usWbedTQm2Q+sPTUEv+3sTAvPAEDR5ZWKhh
tP36bKh86D/38gi/zeTF0h1T3dMfgClQ0Dqmcebk/naQaCv0YI4oP/CeiogRDExOL/4LIDKxGyp2
ISpwds9iKFtVTLEinhEzGGhn6ONdu8sQ4cGtaufXux2Vm41L4bcC01Q8CLrxnExcbzunKQd4Dhhf
zIiZErRIra54NCK5wB9LfXKyroe3fvuP7ENVONYWMQHA5u37WfcDkP3at9IpR0HQCnIBgO6W8caq
us6ayNZF7z8FqNBy6KbAHjs0c6Co8x7P4Apk+mBWrCmxMAVXQU7OXpEGqkNRo2U4cHgbFJG+S46m
lVjmfLjP+TYiLTPtdritqtXQoN7z5XXPK9Hdmn3Sk/KWhlhwvVlglPvAGTi9DSPVZd7JHPw+hPjq
j1C3CFjxwPZ0Kpq18SPBwL1/NCW67YZsN58SNElCpzJoWVsX3hUqOZFYBs5ssqCH1wJdxImQoiQs
IztkxEiWvxxz9x8CHOHQcA7RsIvEMOC0fKkZ0l0I73kpyR3CpG7EsC4k0rxwSMdTOzTfJWc/EwlQ
mppuWTGPSkZ2pcucRG+IjcJYIIuCbkcSyPBEEZiF/jdQn03IukNAUKz+L/XBjr1kZZfYWLNgSEi+
QKZV5VAZC3i6AB4UGCDViV/PX9aaO4mjL89BNQI6ofUFk//iejtJm7yGjZIBntQ3xZ/cxmEwBO4U
NgCRv34tNs1BcSAdygYpfl+Ipr4ytLaeUV4sakqD8USBKFDW1voIixhEgtS827w6h86wqkk97cPN
Yor+Jc0rpSkKQXrC80XbYYP+GlddPfZvR/YZ/Ap9U3pPk+4xo8olFFOBuTBDtolCjqda6c3MvwWJ
L/niQffdyVwqFQ4nmeaR6ABqV+9NCI8meLFQPwDgvNqDwPp5H5dN85Mu61gizzFHyJiigmU88LIj
rXFf2NfPFW4UoCYYT1ZuKGLxVSrv26oaulSUbKr9s0kQNC6vJTo7FnldmKSPa7Ppkq3T8z7jVZlX
a1lxMjHgvN8yuy4cfRjYS3pWiSt6STXik0eK6P3H5kCHLNWJUEDVJHivUt74H6W43HZNOuuAYfgF
G306DkroNgeYxzvkIt02xqLaecKWbAW70sgoY6L/0ebtjJB2ILMOOYdAisOaUj30Frv2t/ZyAmTI
3CONy5eJfwuvkmqMhLvl3ueIDquKpxalNpyueKxaHqWpF2+hVB9kfXfyz39Pvpu0YUdiTTuuB4Ke
2S9N5KQqac2MikuW/IuepdCky0oUvD7uz8QYM/Ov5SfB9V6FlPUp6J0nl8OpT1nMBZCh4OhTtLxl
+Bzs2udXdJbevlVt4Im9fTq7ilgsoQdq55OV+MIphu4WNToaqHwlIdkM7f9E93ujLf9t/byXZSku
aL52zq+UWH0/wrxac/EpKDX3SSGqZlVW6DSaH6DmrcCozXNb2Ab151RwyPJ2gvtcY5VS0DUKNUBc
achTWfcj8c7TsgMfzsfSUY6HCszpj6d2XRP9+naECh1Zp1W54N0H+KuiLmcyKFa0XcDts5VugSUn
eM/5aEkZNRIBL/bG2QWp1XrlyE6DzNs8NTr5n9XuIgvOkTZckxrePNNoMEYnv6bSfRcTdZ9uMMfm
P7NRzwPIz0/HSm11pvVt6CyRrsVK8/FQR0Tylyci/vnj3pSE4f/ohS7RHc4muBSMkW7NFCr5RCcY
TI8mckalFcl02LtAdQ8H+7yVSiZxYLLHuyvoSlI3IqFfS+YN/oB2BzQuapNDgazwsM4Wuh3YtrZC
1fRNFGteVxVJI9gzNbP3Aj+wdCCRnkRmoXVsecWmqe5C+/RjTuv7LBaKcCXIgTVH3NrA2MZzc2Ms
fcvlGp0GF4lC7ItpSssx//xTwlHupZPkLArmoWUPNwCF9O0GHy+uB/S6G9xfjAjxRSayzqT8mbek
pupK0xRveBjCs6WluxC6OBaE8CzmAgn+ODob5uPTrZvJto6TBjOgbgbLwUisVehm+upYrqAiDyUK
HypRm8FnbuXzibm/zQnKDnMaWue1OgiIlb9lcWtuS3DUNbQ1lyOzOCbPNXR0e2MVDxHhT1mayrre
NH6n6Qajg6fMvbtUOIQaLSqzcSSJU2looDXgOW1AcrtoJ7KF9ElUBO8FCkEHJZZuyKkOZX6ViyaT
v8regZuY4h7cyvT/mA1ldXWUVYdKKyzkKcZLef9mxFYAfy95c58jmrxGnkQHJk7wBW516taHFqeH
l1eCiWRggJ95a452DWGQSRo++60v2hENiOg5QIHcNzLmJpmZ+AZO6YWLqZ3AcrQXHXrOp4Vxr/OA
uYoks/IhrNYbu2OatMV3A4RoCMjnfRFdENTxWrSXSXXVYI+jMrCFAggckdTS/Js0+H6w0ozWNymM
dJhwaFQ5i1nF+7WKE+jjM020GYiWDa9WRi1L9Wn+j65tdHbo0VSYDUuuaSP/GtVecQmuVrTDK4E1
0uRK7BGNQsNKXCgUXd6e8bXrxgX8kD7qMpS0Vkia2XOYhmbGnlbVDG9r6ZY9FeEJVsLqp9Rkf3LD
ousCWP4RcLsYaKzPWUr4PVRECK9fKEJMf8Cgt7yBHGHJd16VXsjeHeqySf9Wn0Eb9P6pYWqLBbPU
tpe4ZWZR70bqWGMnNZBrvYJpgGy3QKAtYyi+M+3VTzieCGg5PwTUH2phCtDCPs8d1/uQhlUxgIDy
vycxtLUCGr1p5hBc0dVPfpGsNZ6ME5mxPlTfDgCfKEfeZD7NLuZ3FTrrSq2RnGHBc4Cl3J6VhT85
WdG7xmTUcz+w0D4F+UTPt2gR/5RMHasSpDRg3vgfIbtLF+rZxAZ9dfJ7TVmXmdiH25qQGXV9u8uS
4FgvKUO3UBH/ocu7JM25NtlKbaGyOkGTBkMNOGZbb2C950QTFZ34WCAuiWDx5z40xf40PqXbPrP9
/ONgphqsznvnQluyxn+l48P0thmviZseN5DGCku4Szo5KtkSBhKUXR3zBn/o/j9jrrzQPSc5oAjs
E21w88wPCrWvwPi+R4IgSm6KT3VeISa6oi4N7K8bvAFU4xiUS2nTVKZaC23dhGwhDTh7bby8hlrf
5XADWj5fdPisnTjol1LVY6nwpxBVxRsODxlz1XeDmt6vj7NLmnR3u6FkpBAYIwIvKuqD1QOcQMDR
dDRDxl9nb/QvWOf8vUgIC/NkNZdeIHGjbLFNOnWKr/+zb/UEbiM+DMYCtcmBWtWNhha6LinxaW5n
N5WP0lxip/Bjm/lw/vNGYbrdOhUXivOMsWPCxZGFulByA1ZF1q2TVuFW5/Vd2lzF0nuP3ivkFKaB
OpkSaCI73HEEutFlba9Wm5IxdxgNFMppWMJ7hOB3v4QEu1Ny5hXvdxoL73TS88wgkjpr59aic341
kE50MJvlX6D30PrGNwB1Wst/TcHmOeUqYe8Ao4FL3hJtuurHL7rF2FKG6l3SwCI8dNlitY9sOKqI
arBDJqVN8J6Dectfr5zadGxY9UskDx2rkF46n4TQKYsunuOS69QN8GA56yDTh6yqUY48XdoEz+Qe
+40bI68DmH+IvNEEtz7761UFfdbZDoXGB/s9zudU6NhZvbc/9Ldli/0zLAWX1Kzyh8D/PkG7pCyq
dtwXytKrswXDf4f9UxcY/llFE+Gj24PdD6qjjU3gTT/zFc3OuCpbvu/SLYN86GqmWkNfnb+HWlrC
e+2EXnomtRy25xW2iSvYTKdzR+QPEErHqCPFF4TYth52j6l4/Zs7Exbc2tnAT3PMt5UDQEFIKxrs
LeHsY8i/XaZc259OwovyhQwiesMRl5J19vH8ySnLcKoQ7Qk1959IyVaUVJ7srIam1WEgnfSPmIvT
0w3UkMdKrIEaOXv8hrnzs1YM7G5E6R3kfJUMZHC90fC9ywZEJFgFIjC3wX7xiZYaq2IjJouCs+XR
rSGs3OK6k5hxyvFLTrtXoHkneg6Gqcxo8NSBOkkEM1uzOqbiDSyCwNvIM8T3bvsW+rdTtphr89o9
p+anuYsqEw6/tzE9hE2jU12vBgwYFEgDLNkbWA8sm2NlQnvgHZuDVfujI1otQVaqz2A8/tUGNnqS
4Gw4fECDZ/i3Ke+iHX9Co4vSbGzPRs7TWlnyJEotDWB4USwwwoV5O+NV2k+ZSBEb0rdGUb570Bij
Cfl4yrTDRLjS+crgRTfHq4WD3lvUN9oBZm22kILJLEAQcYcDtM/iEc8GQKAH3ZfxgDIumqyW42n3
gvaF3rJT/0wbm0DdpfuR44/6JOi+FgZOzv8rcmLYhkwp6MeiXLg6vahtQgfJyTSlqSNK45q4XfpC
aSOWhNh7vKWOz47T2cbmRIxFaQDaNqU+6+9UbYi7GNdH6kxwb4tlMpdCvUPvroDcBC1nphM58yww
yTL3omqmeomg43dBz5f1f8iE4HPofZ+8AhZrbbOQaQ/cjV0YOxAShmKduS4RMXqUkR+o3VQ6ctjz
ywfNdj79jiYVI0gF/O+HfRrlVHQZkudwyhZmMPJFAn1v+7YTt0RhbWHsT9b5I0x147s16ipbVnxC
AKTA6J6HV+lkyxEMDBQFamypJiP2sQ9bsl6bs0HrCfhE2SqvwEZZQs6dGsRAstJJkZBTaGWhyj4+
/AWJmMcNYXAIj1UlSJdf8LS5hfUlF8lvKjQkImBIiHOJ80/m2cmwR/dxNIsdiojTgKn4W21j6Js6
oVwLx3kciDdYc8ywjaO+aL/sPGw0azFtbPEknOGUdiuywqRtQRiLMyC91WAWgqdpVIp3QJaWDUGo
M24pPgQ/rz8c+QVtEN0ZkT9lwM3KxQMOMaUhncA3hy1ibsbI1oWoyfwb9p4/LHAxyfMMifgY0nrx
MDIUHeIWWxvYLMr9zTWLrnL3CIczOCHaPLy8pXlUT7NbEeanEtZtRfhj8vj8Y40AmfJ3pXgJ19P1
NF9QxJHHiH70FQtIZzhKtfhmwAYWGkUzp+huU5DqPmJ7stQ5PhMaa6N+1WzvzCfAEs+sD+BThq1W
yUhIHigyaTrOzKl5L4jQa9E2hSTaDpHASeMwTwWQuElUTO9R5H29cUnBDnfFb/7QZKu9DqTlvYzS
cIi+VT7df7PLfLcUOmAcRhtv9je+OKoQY4R/2xKzDnheyEpi2Eb97Xz5DftnuRY6KLoOUH+XxQpo
VAuEh91TXHFcRtYIoqBNXuaFAyOIxmijrVzYxaaB0yp2Rub0KYNN7I8WEnZbSkKc/gqXx17jhg2d
34ZbKOjLnEvFMEzziZQzpN2SqUCADavf1GcicaNUD0o0oonfL6EQLjHvK0i5WpvYYZIJY/P5QR2z
yHx7K0ErCbpEhlTWAN8rpIaGr/NPFMmGZDrX49+jFKTIk81emPGDU+ZPjYg50ZYt0i/wA2GbPKzO
1nsTeF2T+AoSHr4pZSl0STNnH39MSeKZq+PoxwZ7MxNs4hJUtth0TPztGgmn6gxEm1J8xr/BgcYH
XL6s7/Yvjo1A2jjiRuTIB3Eg0YmAhO+hWCXp5UdTcSxnGLwiqXSfNcM1iEH5Dn4v3uwQhIQUfrmq
A0D39frZPa0dA8g+05RkAp+8UOtsl4DICPc11mwA3nnUUL8SNT2EMRUkTenYBwHqRjHRIlEXHykc
ln+cWtuHsbCSZrQspggtQlckuL3dISOLJE8ob7rEaJXXMEt1VP6gyIRF0GuZ8Au4xORccO9c6W/d
OSKYAIggLYFDqI30+vmqoHNYm3MfPvQaAulLfinzxH5n3UmavwU11+KmZPaQfFnWG4nvBK5mI1eq
RF4olhCSusKLipGF+H+yqh64zVFKqC+0y6pTjdlhVVBkTioSaajLBtmxTqKdoDd3M4gj1M+4zBjT
tsfLuhjtpeMgBoyzOd+GcBKoGd/2ZbeqRpdcd8hP/mReWvmD7sfY32eDP/k5iWBktDxyufeIsxQm
6eDEVMSMORwVPc8vvGwCqnvlSgH7Gfygy7mMPvS2cvi23MZjYKSq1rknixLP2M9Jo/5bWvFIUrBy
RFFHpkVJ0RQTeMK8Lf1yyJNNbysnJZozBlXMqZxigb5wmHY1jtC1gXFI2WlRvedrfNjNZ3/UpP//
y44akoFcjw0Av1Q4zqn5fK8CBsNwgsKov+w+c9i5L2rkZe39HnuqOJPXYhgcvNLXuOn82vHsGmpP
9Kmjk2TwcItaxrQXxUTMkD1BscogLLzuVNf1ho2sOTJTDs1GPhZNBIxCxAqJK6ATHGlFD/l1UJ8C
mY5Rr+xuYac79Vs4DS7BqeqG0SJVto+g/sgHRZRN2OfKzuHfMMNNkZKZ1lJry0IGewqPE+sze0gw
2IRNbTrCKR5lyXy9G5xdNg3qeLDAv6I/4OmJw9n5+7x3o/0FLPzzQByka4MRBossoQnFXJAxpcQe
Cu2zbsk2J793+pM+CJnBtpm6vkvQajfpqDhlU4LrcCNAmjgfi7si7NmbhB87Yz7ofhNF601FO3tV
53xhkX59WLgZhPLcs+VqRzmCxZ3VMsLzfyG9KnvnzHLjgLZglMWlDcf+md65ELSsY9UN1j/60BxD
zDzSsbcg2FccmfUhBEqbG0NUpMoAU7crwKIQ17Ck1o6sRRCPOuIJrSc33GN10GOShtlBb0GiQ+El
uZtMvjXfbJbp5JojKlodpDvYRmk3g0iajq7aKMDI87aux8Ct1U0Xz1AMndYnTijXMYrD3Vx2QlRy
7S5jirzKw6egxsJ/Eixs/DPo4eoN/5qOF27fDzHkhL4HkyT9lvZqOcyYulDaD8JdxhRoamsek+IR
rfm6ReE0IO6V95GpXzMbW08cBaIC1Jb0bkTRYg5/NlBZIrZhkAorqISVwcH9k9dMQ1y8FHrYzEip
8/4yMTzgOIHynjbweq+qVOe3vlM6j1e9cPq/LlqZyFC93Bw2nbm7sFhhOAbb/CjhcVkP7RZywyaF
y9CnnZ91yiea5Gaky23Q7oPcv2CRbhT7DLAjzoEyyZZya99PV9Nuq/Mt/mJwF+kZKjQyKu0EMexh
YeWSmacQwSyiFofl2vlZIun3y9OH83uyfaBh8m+O4EMhnBOheVlNRvex/ol8Hk3/6QneCKOfGDOK
zzEMpY4/zxO0UKT/Zj8dUq41fHw2zu9bbh5kUk5oVfotX0EWhA6QmUMzc8qO13sWCp6wfvPBn8Wk
kONR3WY4ir+AB+9GEEdg65YJTNpLvk3pNqxJnWxU23qhRjdEveLZQhFGA2QL85YojMWWSD16bQfO
KJRBDU90kP4XtHzTY8NAcxPbJBAH8vxTZAf051RsvcDDvD5fTjQ89Tq3mcddi+/UFvqqRC8S9EOG
ynpRGLEcPZJDdd8pDvmb7SwOYH7QBSeNuJIhjuETBGO7tt/9yQVwoH1alIfmc0FdQUk/6DOXc8g5
tLY6c3ezjRA+KoCG2bFE4zdbq6cp+n2r++2z/PuzA9raFe99y8GlO+o0xeDLU2TDwNzkQUD/iRxc
a6VUg3EKZBPpD7/p+7JlPhtVlk4aUb651y/fpjqehF3tB/VlnoY6gdZHTxccxXjm7KRIWK9xFZ9z
sjO1ggGEu2YMAUtGi+nuUdIs7tmvHMiSo2TlLzub8nab5fwvW2vNCfgTeT6JbvBk6N3mA7HE7EKy
bQUVANlhsoyjHyMHrnNHygTI7SXS9wmW5hpTrCkzhJQwb3DiCQVXF07SGgZUUiQtN03lR9giLoTe
otwK59a6mZZ42i2DXTlQVJezccTTLoDtXw56B+/cWd/8VoNmYClJ/QaoJi1Xz761EpW0o6hayMfr
atSZ8sj5uiKICtjYcrkncX45EO5YWyBXsUUBhZuviIQlUpEcbWMdNja2rrWkY1X/K8MMsNoywKyX
klSqcbICQ6p4/uOWSYLtieO9CxJ9ATReCQEF5yPTDL1XYc3NNZEzLAIuOXyV+Vzrudw4mYIkjAQt
+ug+y2KzAcnqcWVILrh/AUUcWc1VshNiC+LnVzoj3rVfm52xMaD3z8uLWjnbkQUpc66nVq3uh6FU
WuZuOX+Th9mPtCVskqi3rY/r78GwlMyqCdRi2Sts1OTy+zL75TeXpdSV94FEhLvqxV/XR11ZVn4u
QviS16Bm1idefRUTyA6YkH3m8qVy2VlBymQpvZWOizGDQRRI+xlSzDPdrRjvZNP1juPizyYIHRSo
H7/CxAGyRad8GTgbNuj/wMW/5YKcAezG8RWLnhDvv2V3zI0iDorZLeEXZjWFqMNZ9RBRVyX+yDVI
bu8DtWY1D8Mq2NkJgI7rAmBppwIjOGSfnileF/wHn6fZ5ecKQtS6NWZJGR8iX3QjIDX7aQbl9PS5
yC1tEdPZvzFCixrwgkANoC8L6z0DR4gfFZO6UQ4E45Ivqs11BvUfmB+ZB5Pm/y5U6K9107++ZmF+
mR8xzXHXJF0+LudsYTWLjVvZZ/i4bTCjqNG7aqgb2aqmzL7GpWCqnq97GntjbOmn66yo7W+SOHXb
jRoDaQg181xc23B27B3lUG9eMh+PW2RHkwrcnKd6SfJDLui+b428MzKcv5fS6/KKx1Bw9mFDMr6q
88KkntYbn6vU4SEA3N8z0olT3JW15f5VyW7ZecouPLx0BlyrbUDIoAlydOySnv4/SwbVh+nX9Km/
h2IQlWP1IjzHZVjQek/zCuo3DidsYKss+vOxxWDMHNAENG9ohsfF/l/0kWurfH6jTOJ3xGf6xOI0
xv4hDEj+74NnQ8knOlXajApHb/ZkTCgBHq9fp174451iN3b4SdTe2ChgpzQBM4o256Boa9GLHPhU
lvMv0acgN0DOWz3xF4UnQe94xM5aMvStQwvF6oXLUSsKeRhyCf68UdEo/XuMOH5boP/GVOCY9UGr
Uc63tOlU+DI38lbyGIN3KoXIbfF/PqG4h1p6bwfUrxGI12q86ou6DN0k2gSBD/OAob2iOdqkxFYH
c0PeLkvKi1P2iSGHh488h8pCwQvoTaBrYMTCVHXDrcMCHpos9DCCc0CCDrwdZAs4+mN4XwQNi9j3
Iq+jqAX19brT7XAm4PTy5BEsPtB/TTTFq+tqNfoCJw93S1QCYr6OM0G5zxGTWyN4l4uBbgeR27sr
XPkpo0CDeVz3qKGObhQTjYvECvch+q+yzOhEQbQor/M/EWBNJsZsOhvcSFg5hoaFlt149iHPKXc3
J8hP5lrTcLe+KKKjpJi5nMw97Ocg8goNSNKOdIJVp38zccYbPcloI3hnECYKuKDGSCM5Hu2dwn04
6Nf9fVRXVDZ3B+0CEj72j0MnfrRPUYROzI+wwBrnHxz+8UdGmG3TNXStpFW3KgKNjz9Ic5zg+mFp
3AAJMvgByA5Y3MuIJ+nN5Jz67+UeL7RawCCpVByTzMUPCYohN3IU372pAG61NB+id/QoUJTFyMmU
nS5Ncl2tkw9OdPVwYFo8vjdrFGKxb4O0WFyCCKG9NScH2E5StCQ2oktLqUI5ZJ0DEh6BD9SQ+oSs
6H2uoD8rTAarx2IL/Q29bXZxDlPPIYZwe/9ZAOsPcO7CdmM/nE6WWeWbqzroucCw8HcZKPnmrExl
7KE6n4SPobqwGhApy/loLVSOChXftGsLDTeqmCi8D7KwzCN412dCwLOPScqJZ2VBWRxvhVFQjHNK
uic+HP8qLpoSCW3Fkf1O/J/n/4VLOK1vCT1e0M8sy4h5Ypq9t6BQo4yTiyLrMj2ck8tBvXOdGWuG
pS/piPqkXy7rnu/jHywdLAJSBG2npnfyRXNJCxvtsyC2VgpO/v+trbXtIYMaEwl9C9gdG4R3i+cF
CPG2QV/NEGBaZ9oaWfVLNkrnHfm0dQxjieQboPZnP7Kl7Os+zYPfKlBx+sHs3CTHR5lgHXNzfv0O
rpbBuPTYW2vB0FlPLqHdRSzKxXrot0Lx7T0f3trNr/LW44zQxXFt00y8Mq+RD9ZTQfc/Mu33/MHy
PkW5aVHfCd9Qg0+TIqdtQ6g26jyGDvZsp+FYZXvqWa+a8IWPz+qhG4Pk7IsS6GJAS3L4UUO+bcll
VE/JJnfVo2dbFK7cKrGcHsKKpVlwC9QXeHZ9Fa6z+f3wqw9YKdPBIvCNaNhhpV0+klRB+cNdvp23
XVbe9jxmb84byZ6luXs85OcBbPJX49TDjunjxI3R/zDq4pfmTZ7/o6RDuAtevSLlKOAR0wzEU/Kg
RYpBzsodmveqymskssZtxHC8kSKnVAiGNd6UwdcSVUIW+NOOuEmTm3AtQYEfGg9YqhaRvemccJAc
5ophc3QSie9r6+0/CsJlzkGDNk7mXSstZRY2aXsm7xFxaIwDOl5XdtCvKZOERM/RWWpv768qWoei
Jh8YOk6as+DTyRz6Q1s35Qg3M34KBDD+RvQUeXWPuwV6Y9AVxXPKcNkJf6iPvB0P5Ahn1LtN/0as
CnWXceJdBrPiT+t4FRJK1fJCBrFsoSneavvd0FexW07n4huhJEA75uS+j2r3Ef46Z3iXSmlEu7mu
HJP7mw/k78M+yEwsfF/BTxDeCNv2BRoecoQLtYmI+ppqYsPKgNnulLaLeVBTIIMzW6NZPNBd7ACd
5F4kkDUhO16eP3D9Kp2E7KlIo5/v17pFsJcAt/ZpvSxV7jTOTM7vew7UhTo50j62LHo6icx82EXK
tTW9ZKIIwhAjOkxMfpexgSPaDBYwS/5Y+WUuCgBNnW6XK6Q4bnt13Qihf0NRZjY7lEoUDEJS6nS8
WQwlLGspHetiTbZzmkmd4YSmSsZ6bpSpeWtJOkgVP8ktWA+NGX2WqMYbVrQt+Qs4YmRYs/vGpjAE
VpCDXUZrYKjmBWY1q/9F/NUpyUpqDo/P5BK8byaP6Kady76WdJx1aj/eDVUFCAipFL6ZSl87ldWp
Ds/KTO5dLAd4XHd94KGUzOOReJAdT6PqKn2SKVHkGq/cjGXUs5lpF1n7J+5sdWzOnkMZ2WCFZxRz
PsVJDKY6WsjZYdHgMP71Unhg+pubihzafkcDQOyMX0HWUKPgqWMUDPNksySBldr687ZT2+ig48vE
j5jT7R/t+NcGSHbbE01y+RN8TabJv5UmhLEOftTDVjUT3sYIC5TDJKw3xU4Fgxr65FCBV21hBU7S
0Y9PTaTcwV57ouwNuF2m+pHtcj/V1sVoptV3T2BChRfcwvwGUPT5NCrARtVGGZL8bA9m6Jdq8rmE
L0NeP0Rilceq8qVJ50abJYZvpkVMlrzCXEXIoUVW0SKZaVqhQ88Dt5iMdY0gjkJpGwCYpEzovN+j
ERAV+akaVb0E8oxMsNCbRKDBarPFjJqFpImGFNmRpwvgzRkUgGA6J5U5Z0q+qv57/H36gXpGVtRQ
fZoyz3PbYon3gIvhXDgaBeub4/Y4r9aby9oOHnr/N8/dJV2VlW60e6a7ib/Hw8cMQVrP7RYV2Li6
AozWv6RDgGl1ZeVd1vwR4MJTCO6bhfPbmyqG4EPpXE24YP+/IN83dmrmLCtOP9VKZSh83susLpqY
fhMbhkUh711iGkNUxM0L842m69FqCSKZ634GCLUL10Y3htdYb/mfCe/OQ7pkZpPIuCpzwgrBC7da
0QixSffR7nH7Jjet3fzoDzq9+odQEN0A1l34KwqrvdL5JIdJDebl+tEGB+Oiy31o7vcwbDqX0hR4
c8E955i5WDdpkLP+OGPhsCwzuQIGoR1W1Ip6kfds0jYGZfLv+rf/OsEoG3ouf4nK6N/4glTP/Zib
Elo/8NPeRlVAeZpskU/Fug5h+4yIOlWEjxUTgVMZzDM2mAVCA0CLCdhIthhPdGO9LRQLYWng8AVi
VBgYIcwdx66ZlumQI5Kpn+h/z29Autjl0SHI9NessZ+Mr14li86C02sFAKLGa8l6QeAsgQQTl5E5
mUDnfWmU6uFV1AsbTRtyTBPpFOMRwUm3Totwmv+HlEeMCcCNOBVD0jlHNC6FNdtQx+v+fX6zfIvz
4lFKFbqGhdY2XXnIFwUnrdL29m/qA6tIp+UL6U5tTIC2OxS5xeWTwFSWRLR0bxAt8bsQjWr5gcff
kA1DIDYor3ezf1Brpqu1a4MteGhkBrE52qAeAs4HrX9fbEhoZTpW4iWWlgWPaLtvjaTJXMLsBd/o
ShEZbznB3720mQoH3BeKFEmuFH7TkT/DBzU3iTnm898NZF8JZaQMhcIGPUXatAg+1p6PjR43buxp
eiGyAIBj0ICTlCc62yoW076bQ9jcQOuVRqJS10jIhT4D+cpYSdAvz1U93W8nk7j/OqPbA/kthvNy
y9BJGDpK3ntLAUNZB6NzmtwIKdAhrdppfPRrQ1zm9wlAJY+iw39nol686DYpaNQSa2VyZ1NaU0OK
2Ah4ofrJdLCJqVxzPzfnCNDhRSVfB9m33scGD471cWWmSjUu9d5aUoS41cP16HQcenrMcFK1P2s3
B53avQDFZ54DeZXkWgLn9JqzuybkPCIdRIW6zsIlD7mtByVXRHrkl3myrI9qaGx8G/vFTf19n0ur
dhH+PSnF9UxQSsGZVw1XtBqxx0PraUTvsAbskMWRafmcAc7G1PJWBMIc0hCVKft4HEucaTXkbQ4V
DAswuJ3p8NAguyU62PKXV4A0xSELI5cMqrsQa/BqOUfbVpaOgH+85FSHkxPv+6wCIZfED9MkfmOR
fJUF6t+W4lrITZmfpTVMUeEn+HhiU8aEcsk4ZKfL2y9rXMceglBCHOghpQ8fHPWof0nRkdrE7XgQ
e7mHxsm7hp1BmLhnoSqqhCuvzNe9Z+lKumUkCKLkMGeFNaCtzkdjkHmb+MLe8T9UCjUJMPT7VQrs
8CrqrS2snsoopQ4q+VjzCB/cKqucjDIh1jWCAs+TfD/LfFR1edQL3VWHy7g7qUiWxSUwROZbAaQI
So06FU6+apgobuCCIGBo3BZB9Vl2KW+6X2JZ/BKRlhlKJ4RddE+FAz+DLdkoV3hRv2iKL9ewzS6M
hKoUwCOKX7nrZsnB6KUtOaaUci1sDA64eip3dB/5otCiSOJaHnXjgm5yAaKvZq7qkaIOJ3DVZ05U
UBzwhgGJuBXYRj6XnKdeQ1Oak/g8yk5iLpjuSdkxh/UXUFkSSCnqJTSk4lXIFq1OxhnopenLo7Yl
8JQBZfN37xxelRsMM/CQ5Tgj5lqV/3Q0/FsSIk4lqSPOf0nPUAbwA/c6OxL9l/KEF3ZNP+yOVSjM
CAOjiBffTAD3nfySOwKvXSmr4uT/7da2SkPqIFiQ1Qu322BctFy1JQ/eY8dAdffodhedgReTNIdb
r6L3SS0s9S6fyAd9eqqBFgois123GAolVq/Enq3gMvT4/GN1IYiEEtSEl/ZoAWuh6ie3bbnmoNtL
4l6Vqo5tMV7lQpOo0diofC8kcdfVhqBP2P4vNHE31FEOuco4/LrfChWPDmtqLBbqrdgN4LUknSPP
2dN+cZ2X7T3frjVKAbu88Re03vc88IXJ8G6Ettv+MiOHvlfOPiOyIEdgKf547pqs5p5K2FTdkdBN
n30RVIafGrZCWD5d0HMsMJCA4MOQAmPEAzpVigMz/NgADnXo+PFpKBYBaiEqRiqGO1VNe2ZfBWeB
Junjz8ZUiK0sTzD9iwr9RDaPADYKzViRglHKYsdVMHXNKQ5X8uhDB+tuFrKuBKWuQcU1FCxn+uXY
GgC1ji3NjOxoC7e/2HezPT9XTev/t6y8Rp8XGPvmcVOZny6fu0bI8JO33pGp0SxtF1Pooq67w4Hw
MjDKl7rKl9fwiHWY7OTAbdStHTYil2Xh8lN4kKnaJzA9QmdHzTMo/6V5K07VHI1Gs9zfo1d2avCj
dp6Ekei2Tq97VYfaFOnLBfCOz8ylc5/JGeR62/+LRNwyVIOkX+T5q7kgLqEwicbE+Wv8RWuBort4
+fGVOQXIgdbwS5LsOc+pXzp5t1hZoTOQm+mwfS70iRcLMWhWF/y6ndTM0s8Szu7eOaMONNA4htA3
oIaYYkcIipNgZOR2zyoWw0Heo2ZNjZj4kBpDgjP0FwsNydYRLPOIzRyJNOibyrZrgkJvxXwbJBWo
xbNOLDnfRWVAur4nqx2YWRi/fPi5SxmMtLcBQLRdZySDS2gUM/51Ye21ogUe4HHmeqkPBuRYI5bP
32H6BpYj0KLl5qwCjYKvlmWhnHt9VQuo/0eeLdrBFyyV0fapiS5gQ4MmuAHGaRS6swaJ8IiMmvmI
0vqy5YVdHQ4r27KMDfgM04QKojTfWjl8zlVMKz02PwrTMl1Wfl4AbKzkUKnVipMoJ0rJIXORdFGN
xi0KjyjUBKjIahWI+6LFeOSR4sGjSp+MAeP1wRxS7CHp8l+63yeVbti0Tb/lbobRgXXQNJIgapFj
ZTHIIi379MFg0hoA/0Nwd+KIgwL6LbhZyWOEYIQo4wY+eOKH5cnRLBSliQy7kvu5Gnl3jmw2vsfG
Bp+uNBVs2gXg/KNR2mpTWG86JZwgsyG2SWB5ELRrt8NmxKkx8duHKqri4Y557GlZVfMJEJsQvNi/
N/L6XisFk6r/LT+Rgsv0MQT90VAzJd1mHMJssoG2zpNn2gPfc0j0CfmdLdCTsQGhUNgt6GGfRlrS
zik6736taR94LUPWCDbCtRNVuxAhvN8tAhuBK4kWiZlBBjytSKmKnUN1seCGGJIuepJOqgdPvd4s
T3qORlqcDTVu1GlEYFqb6ETdL8fnGq9zbLH98PfEYZFK5V7i4nKYm/LR+ktQU8sbK94/pQ8ovdB6
/1G0zxDDi6VV85G/gKDKQQb6TzYBreD7bXhMQ+CNOHiCL9VworALEx0BvWBbpU00XoVZO4vN10pz
NLMK22DlHMwmMuEPN8sIld81foCB3nt3EbhwSS5JxKm+a1neXI5fYNC78kaZ/F4DFO26BEJCUyhE
yNkTnRt3Z1qNWZrQmxDtnR3csPt0n46kPJChOyxRgf6IvGYBmBOSrlMEw6Yu2pR6pdIcwUtnkIeV
RvX9gKsyyfVPXB16R6h1WIU1901BJ678vQfG4YXS6fy91INSXd5AcCNVScBMGiNVtXGDuvFX+sKf
1J31zeHJ/fhRdJF0pUQyJZKjnAWQV6nTtsPs5vEDzY8E4xeZj1PVoTTdyYhzQrzsSgN0QS3Pnwx9
hdpYWGlAeRg6gR4XrHs7AJsAuQxt5ZGCZHA73TX50w/0wiLSE3MgBiIGiKfuJDB0k8mpdkopWK7i
kZGCtiobM4yuX53/N7heHrB9iRfev/rfz0OLYpzEAmrrPZVvbiGx7bENQKBE1zycvGlwzKeLIOv3
Wojjfme5cVD0l76ivyu2Q6RO2TxD
`protect end_protected
