-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
oOytExz693d7CuoiwDtWuhYyPqChrMeBNwgsIX3eR+OobK+gYdGnXbSg6l/HGFe4O9lhKqM9ezCM
A5QdTlJMbYnRUBChJXOhRURTCdJNbNM1wb/LJ8pWDI9pl0gqwGjcu3FATDubhDXSVhmdhfWVCuxb
fmiqwHABy/cKUVHq/ScUtTVRzrONPHB19oKyTMNrvoIduXBiBmoUcTlAqe4Goy2XhcDHP9M74lX0
2tiiFSoaRkbZjXviY0O7dMYMBlo71ABaq4mpFjFROxMPEnQ8pUI4Yn/SCYv8QFXriYpsXkJjsdze
GV6GJChPNEAcQQ/drx7jd5iuiWXfIWdZLWhzvA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6576)
`protect data_block
eMu2A7ATKs6ASKqsI0XXNKgec6F8b9FvQovtL46hZPSPc2BYYn6+D9bs/kJf54MSo3QgIa0TDMzT
jcTsE1HUMrc/4yaGM3MVNz7RGgdPsdYLOc22vZmVSxIuTjo/n2mrkprD5ofZ1Nd6PP3TbU+o2Fr3
PuyjEO7ViXdyR4D4zk8MuH1+SDJeHee9KruhnAr/RGxOfLysdZRmIbdNSH5tLUHtsjnJiSYvXh1v
6zFzTPK38ozeCxuBBz+IAMxSkH+pfVOgnUAtFxauJ42nuuZc7bjODn0q1ngfD5QOcFpXxltKRIBN
F/wAT9Gd1laf2NrSIXRrPgkzUkOh/9TgwDGDRhsbXj5VkRhcX1kb0IymGX4VuJRQJGz1z4t98bIM
uyy5SsVq8Mfa2R29KJE7AMFtYmWpVpeitqQtNUkxc04YnSlMRrxeSuJKdzauEoqlw6JZwgpx0SUL
ernK3N1wBdsL8cI7OSbFUl7Vh4tCKNBQ2N4Vn7SUvC9HyaW8ZbDzJPxHlwvtwFJEzDFSIuAIR8CV
frSL3S/PvQEUZnavkIGGfiQUorjOfGVQAIhZ0Y/1pv+6/ATcKElcCFZFW1kzXg5pVRjJmBE9sZuZ
KM5CmKbAj58sbMRq8VlwEFCT9erx/TXFy5gTwPd6WHmJqB6omxL/+/yAAzg79Hl47E8vwe87da63
DiwgyQUbMw794/qsS79hK8+uVt+kI5mRZqZVmXfhC3ElJ1k9y7UVOQjwhnhzvQZmKs4tssvrIt9L
mY0WBRZw6lfvUWXgj4OnBefxFmPq0qihXwPSTvA4ERZoF0z/9y3OeGySfePqF1Glyitu5bRQE9Gf
edXDtytfkU1RSvfBlopgOdrA56+15F9g44UG+0ZWXJCdSS0Vp07E2KBIaEM2v6PRzxQFjMDxBPcQ
usOBRhTupN+9AAEaQ1fRl2JnKk0pK2zKkNKS74K3OwvcxXxZgfCxIaC7WoNER/Cz2n9yDxI0W6yJ
6ml3xgYOEz6YsbyRO0uMbFUN9+DFVKArT4j4wt6NgBgcg0R1PZZURKvTLPY5BL97VOXR2KKBEKXE
vH1fud/KqI3+k5TKOr6CCXxCD5Xp7TgN06nLgfo30DFoF/GAzgwmUdjR5ilFZthB7Rjmxyaq/MAb
ooU5qaVEU9M3t32akM74hY6x9HqBLFy5Y+NPHfIypNpyAAstHeGMtroeRmbCBewjvcjC4ZBcfFMY
kPQLoOhxpYzerPe2Z+iQn2/yCHz9bNZMA9F1ft2HDbRq1s1HSyTUYy6goJmoS+HR+Ab3u0zYX1bY
Inu6Ao9STpSaz4RRCHdfEJ3wUp1OU0Sepb00yZUgwDIquiMIPWCdeLPKRtgwwBU3Bqqtfm4Zy2JS
QA4+NMpNnsr/p6iFsHNnsjYK2BIroH9Zk2H+4HU8EbnEcgU2ag60ghB/Hl8XsBD9pxVqUY3iFeD3
srtspXB4/FY5W4ubJm9oU8erMAcAQ76J541z2gBaGBqdKzjMzen7X1ZnVOwDgyCiNDAT2STO1OFW
xqVp5dPmUzusp+wd7xBfPv9+Ic9G3JQ7yh5hNbPklv0qqyyWfSsaAL9Vz6OrWX5mqeSGTRl57qYD
GGBckgTSWm7O+rnNvbDJE7FVZwtVtUFaAjoVH+A2b10PWaeQWaBVhvrwOmvvWIiUftv/4TY7s+TX
m9+WQGaboSt6ku+cPeZzvSKkm7P42LlPahCy1wcD7TXV4EVmAsF2X4c4y0DN6AvNBtwt7iWPGKjL
mn0ZHeKKGlPmhAgwTQzHe5Zfo/c1KWhXruX9WiEXMuCdSTHk4lMoRUP7yRbChPb7o6oR9ceT/zav
ihZERmticwrwhP+2Jp/jVR+3bN/6LBUvmQoSs/E9X4dUxb2ygYLqI40gquS53+wp6GT9CxOfwMO2
KF3xuSsK2pM0m7t47rBh6+l77Zf8a12PPEBWKxGO9/BNoT/clDt3nCkCLPMwd497rMRl7Vwhri5G
9BrLvY4WKBTj3eUakS2ifHcKqALv+X17CXaUAD5f42DNu7RTjaDMa1A2QGdlDDohBtJ7a4l+xkst
678beTXhWtkCT0OaMTw1FmIRcJtm9wjda/ALFHteQOGp0NwqdLkoTXAFezfwN6KarppFFD40kcbm
MAXX3BQbG5SRSBcn+MQUfUMf6SeeYtQAHm9APlapvB1DBBv+DX2deTeBKIBPHCJjU15+shp9lJHg
zTyBZZtl0guiMhZErs+uMYjMpLsLRZWOqphI0FJ2MPK81a3PSuj5Z47hBTiM4VX/dypel/qgYJn1
vXWjJ5UcN1OcxJvwxFAuL47Dqs2Nyh24+WrtVVexlYHoCDeYR74m3VZff48zjYPBmSOURgy/l7XT
N+ChItJrplZQgYnHdN8bD2mNfSCHDQwbsHlY25aKj72lPl00lqnNFXi4Q/9CfbXLwAmMR9FLuRYb
0nX6EpOOzLuVBrD8lU690Dp+BSqY9Gd3V1WXc1TKrLo+n4cQSJGwpOGxxBH6uOXQ0kQ+uuKKp90G
qy0lJj46BpeVYHPBjqvDk+bL0RclUqRjDexSVB83g+8s18C1392w6WasK6GQKMkKG5k3QA9Eda3m
KAZhHEgeQDblD26aNHIsIDZBMXQHr6ZJvbNxM13+8pQtBowT4YzvpkQV9pce7OqP358kyg4KTdLX
LXHpdMhGSnejSSuiJ7qSQsNC41U4kZYSB/qObUXwLi30xRZDEmAn+FR085Fma2osXlAaGck34Udg
baW50dFZoUcyMvHkrOXXpPP5zCWcYDaqZt9F3CtrBsLl6iDMUfeDmE/sC2zTrg4+qe9erJDU11nf
UgWgF4G2bpkL7ig6/QoktK5fpFiZxNxvbvB1//DDMpae4YypPt1WsiGsPC1EpdPPPHW5raQTVzB1
o0Jj3cT6G5OjJ4jJ9RgOfT5Q9wV2b406+RKaRPMi/zs7JWoEQ1D28T2Jos+iPNUbpGPPKaalghYv
hPOq1dKvTr82/CGJA2oSylZ32nNTt2XuTEaUaReSJS18o9OP9R9a/5qIFOPO70ncYd0Ayq6R4B/T
cVNemfyPkvvNUMR/e9NLeMjGm/V9LO18P1PNGHClCUJqwxZcZL/Rq0hZhUqQxxdWgcKIlMWhPJkH
JHEH0if7z9D5BTZ7DtK4e0AaqVnRIIWW1CTfIsKg8ZoHVQfAAR8xAgqKacH97Yk3XXOYG8HD5zGV
e8rPJjDkj8dbdi/4+7OvjL1+7ul5EtChW+/aoQYIhdH+JF0noO03EFkRbDdUHuBv0U15yFMFeXSX
cCfhIlLoGRZMySf3OAcMiQKbprSWiRKrZ98KDGKFU9ct7Pba89rkiNj2tx0rFKzUxDrAZlFQvGjz
Z1x/MFr4kvAgRGjwN7XIhnna3kwR4aF+EnPokPWFy4ENcUoVwAU1g6tEYzGbt23GP2NwnLZJYnOe
sG9vpCcdyMHirM7Mtu/MCIFb0A6mKiI9xRLOk0PV0Yd8FCzMx5lrqKPmYXpx5HF5CzAxBXea3uHY
em6CqMSp3HvUAFrAcsDI8FYHSdP/xUjhUV4FW2Htfapv7GarcoxJloZgkwwxNpXmFhiQzgh2S6l0
Fl6itsp3Vr2mQ5kFpe7Ie8RLELlo/pYL8xvp8uFF+M2ZGx62RwTOrEyVAxyFK2bXUoqgGjRsVz1L
U9/6mWHj3sanml2lgcsPkpRQMzow4F1CzYogDuEVKDYFX+ihLJt6hqiUjMMGtKtu1Kf04nLydifR
e+ZAbkf60Q/sMF90qACW+rx3CSIdFfjDNC8rjCSu8ct15am776XV893viZOE1OHTemDNewO1w37V
G9JQpfXnIsPs8RT8GVJQe10SLaJueYCuIz3KopVjq7nS/oflx6W5uk5oxpkmlLUoxLtfiPX7MaAy
ApzLg0WwhnvwoyVcycf47nXtQK7KxQaklTniyLUDQkI25owJobuDkwyUo9sZWFJ17XkY5+HJM9B3
uv6oUPx6IN/+he0Hkm50WnT+JJdazPJ2qqjam5xlt2NlfxA+egahWRXO8BacfIDJmh3sr38mSMh4
6JU2gAmj2M/4Nrnrl/Jb8BPyE6e06WznqW3PuL+BIfgDSOWonK8L2d4E9Quc5ngBu3y5swxjmAsc
5XhwkOrST6Y7zRGRVrdB7hHIShmGxw36YMa5jBqQh3ZKZuJpm787BMB1pk2EEm2kYRUfanARefuX
cL9NWd5lVBpPgZwyTDOr2sjLxoiq0gJnma5vj/u5UpmqogVym21hsDFEjlNKOUNbUR65fcccYqAZ
OACpQpFd+w0HXpUE3DvWDBiXFy/jHCzuCAqYavaRXbVe13rLCIofkIrYv7Y4cA1I6rIldCU7aNR0
tiPt+Sk5+P/KyUeYfKpDJ9b0ihFteS74tsRwuHap8+WMxyNC4+ITQfoMoSu1TrIA3vovDs7jvhjZ
o+TNrug2MA84WzCBQsVxz191UYZxPSAPjY57xifqJMy+Kgv8XprANmGWKpMZdw2lZxILjUlphYJn
RbCjQUQ4FKXgoslRpFMDuv7xMyl2+SCVshgWz6xXs6RU1EYopJBKfzFSNY6W2FzdMxU7B0EEJnJQ
nwF8EonzED7KtTU0B7G5587dXw6WRakoZwuJ76685UzHd8CFTdfC1JIej6XgqqlEQ22dtViZGxrv
PXQTY4+bP8z5rBpfQWJKvicAGmUjDTZ0uM3hj9FIwgF93Beulw6UuMb21bV61V+/LEuzYw08sX5t
lHYwCHAltMPofGyLIIAMDlEXm/FTjZZjW3E0VGfRudvQ+JwN9tEzhYDD2DpQqSNLunkDH/sYA0ZN
WgwZc/qfOSHBAnyu0z/LUtTCrWzCA1+ghatFKqsoVePw4ibReL/LNVnm0e+7uExABdiGuFz5OIgP
3ER0u8rb5lRWOGnFkIo2XSFMubJjNlSSBtZx+ciAkGKO/N70OcoPLKq7b4ZmsOUPRLxVKL5jH5UX
eGARh+MzB73eTqIVBAv4NRvgBPZdw+rspxcxTJXCkRb4jGSPfr7T696OBn32yvJUUmw6cXWZdkED
cDo1B18Ab64lqdDZ0NtTP1RtSdswO8d9NVTxiXDn/2XnMbkcMj9FUwJ+QnposwDdJn+IHXzGrK+n
My5MemjAQPqm+jTieuQYz5S+BHWQlokN7VnPr2r17Rp21hD7ki16H0PHdVN97/+nwOw0qU8+0G+L
SEhvCAD0aU2l4Dk+bbMshTt0lfwW50gG5JTBTYyVOeur+uLm2Q5TrSCUCiCBaLomKI6W3WE5Cz5J
mZiys0dX6GguknuPtdXogDAndsXwYvocEooTNfr+HjVJ3ykh0uQuWAEkdhSLuBAtmauGsNcvRwln
3jISjIt1rd6tPRmpx+Y5hzcLEhQhGQcfa/MeuCFa3IxikZ4rxsAmjheFbqwxSaBG+2WqweoBzq+M
rkIVurDuYn7qTjbmzy06DoIrf3k7Tem7WUCHirC5FFjZR5u21g3RhHdL4uIEA4Y8aRLNrGHAu/B9
qFONSFOcGwDVjR2CKgPV8EQVVF0fO6bRoU/DBk21wFsLPAJERq78E3UNP87njnoyA7Wh6kM5Lfhz
hK8WCP0M/k4/q4C7AJhhJfxST1mpoH7iOHFgo09qzlRCewSXwXA8vs9M5ytGmCSb+gxspFU4Lj64
Up4YW4J3lacCjPWkvg7IiqCb0wNCImOqu67i54BsT3HwZe6GC2yl+yRiAsnDLLT4YBJHqH/lp/t1
1uokck+an58rLAdZIFdUew37eGVgwv/ltF81cnb/6f6KSiqbiHkE7YJRaikcIT74yqWfri+UXHAC
ZaiD+HgFiAT5JujWDywJ+s2sL2oGxoAIPaDmxU3w8PJA5jRg5G83znTFMxnofSboeYgEng+Kin4b
j2/No4gWqiIxmbJq/niva2PnYxJV5KOAtkIEO5Kr8brQ9Guae+aSKY0NOwqk/dvGZUBMg8Ghy03q
gSQzAVUURc3/ZLy3ACmszkRLzcBZ7mKoxQJEuVCIujG9c0ZgbTM547se7sqT8OL2MEfPjOjaQwzu
ajN2CvLXYudIPAKVJEWqxADPFeMsR6akiU7iovJ6dM+iiNC8W7it9BEqGSG3RcnjpJVdxBzVg+9n
ZHCB4/QkavuZAcM40nCjVdeEInuqA9B5RLy5Ik/NL5NmdkldrwadjudIRohMm9+5UZUTfTfpcQSi
ygOlrkpu3lNdDBfsD4a6JyxmWLvicZ1etB7MGnVKbqJRclS286U8cjCs6QOvXjDzpWwX7Jb7XeAa
NmbUZg3bmxQMNifVyaWlKg/guJELoZK8jjZJbt37YfreFqy4Ila170uSQZgjS450ikW2uOPGs4xl
CRp4Yfolx2PRs7Zy8CcEsCOml2xlvS5kaD+eXxQv2wD43LiGgEofJRWjpPd69GosqOb2+a+Lrv6P
AhieQWJHLD3xaiE8B6P51ptG8/5K3cijX8TbYMcfJ1CkVo697OSkp0OPpem66b5XnlrXdr+oFGZj
PcPjET+E6pfIGRLnF/A7sPdi9PH0za+sCFVY+OxE8236W9klhTFCVhqzNx3HXZswCds3eqHtmtF4
R4S3mgalZruOIGaMGif+tuWyMrJcwjPzRtRs0tn6Gc9rief0TFKWlljtg3DCkVnAkS1/nUfQilWt
/kV1hYPO4jpBm/uz2Z/0L9xGtnkDbm+vnLfnXZ9q4+xbONFeC6pZkikM0dFU9Fem1+cofLJhGWNr
sLR2Uf5SIDOB7cBdgktHNf1BAPs9G6hQp00q1z6CahiBkyXJJInFAfVJNS3z2sp5nYz9eS8hbtz1
aoRaSlwOqm1Ad9HnbdCjIiSRzbm1VO0D/lOh3px/963G0KbgKgJ+ZbERIT7bNOHFiNnasnU6ztSB
P/hin6IHDhpjvfqCmRFkHQ7hHGi2YsWQ8PW//yUH/5tWpUQMrIwhkUt2KhWyA6flyF8aD5CHHb3T
Q3FGHRwyRZ2BpZJJjpPwAzqPKKBH4MgbccqzpyZfRBXUlyUusZQTXBZ3eM4LM1CVe+j1WZbrYsF0
f+t3ZT6dnsE8glpnCp/RelflEzicrXrYYmDgQUzIpRJHdNlb9aFZOdG4Yo63QOwuOKfovHc44y6C
CeGZPalm+d8MBwMQdU+EwYDiQPDahuRCoP5vFdXZA55EgM0RdOM5FVEkhxXPI0mhtjb6DWWk7o2d
MydrQLrdyQaQBWu9yUj4DTXQhurMi9SZx5gdSizjALzSSv6lDNpTSqLTiPosQl1dO/Izx/XmInh1
qI8K4lEnZ2EmFwCXXUGxxH0qc3Xp1Qnp0l1VyHfOABsAM+aOAFbqugJNDLo6ETAMfHcTe0i/TTAx
nSYag4hBKu9lW8nzngidTNaNhLin27ZNZKRLzPqO0mj8q+kNqAm78x5ibgp8pNdUVLf5lmWRD0dU
NCkuM/gs4WSIjRhwIHqmdOPOoWqb/k3d8QOre36X9Eu5s5CqrLyXY2dkLiUI+TGuYN6Mgc21+pzC
YI3i6QLvwMUL98pqNQRylfHfJ4euBq1UsUHNzgCWsySHEiK11K4W8Yh8mrODaQP6nGbVWPGe7JIj
+R6s9BhYirYpmZa/3HwJ96k4HjVWP5ApNG46ZlsPUyZ0pr6i0xeyixUjPQG7uO9KHB0fPOvkPxQp
xQka7wgAeKumGsYBHIgAExmak67FMhA+7kF1VrfNbiNf3b/R0c3c3ERPGLjeD5UGwe5cydx8SIUC
aiqHsXF8zqYqOAyFo6933glhvFj8eqhUzP0z3NCoa7jUVFj2hm0M+BoJMmlvXeCFUGvz5olMnf+L
KENXP/wUVUYMQsE8wbDjLVdwpEaeKk5/Wtm+TEkSqAtX5cM/8Hn/CYLGanzSsVVc7Nk5Ld/9A33H
oQZ/Swq/YOlRkTAx0xtyJQZzSsnpYCjhaJy4/uREHLgpM59egIROG1I7pThNXi1pZDfKyNgc0hgE
Xl5ySe0SzlTq/qSQlxuiTPlIeqYo09wlwnzzCMaUPObLGz7CxVzpOoG8VU99j6T6eHoiPmVV1gZm
tY9W3vEeqyUxrDq/KvVtA5uaW+nBURWPXOS7Qkor0SP6TRmKNNT0/QwNIKdECOsHoYa0fpI4V5ST
LPQlhmFx6q9ONzQ3OLZecOjMu4RRhEqHtFdM4kx4RmHIqHvRK0gTrU0Wat6KcxJ0Y7XZMODsBtcg
n0JCTay/pxoUql4xtioUovANaHsjOJrTAHuYI/KrLYbSY+c9c0r6goBKYvg+Lh3OaaYhCR0BJm8u
KFBPX+2DL4mCVtiUKfiq6UFXNkjBJGpWoy/RG6FTgEM56CjE4gh0u5YXPJiPymgYFfDQ+QvaHY31
ToY0BAONPeBNfNn8IkQoV3qZ3Zhjh9VViP8PBqwx0qUc1M+FSSh7TmthcZs6kKmPnMIyU56zMYNQ
b+pVWpequ8h9VSKo5mEdTsTY8UAlyiHCU969KdjrC6xSSL/A1x5YkiAG8VBhtSPFg7++PuhJXcwQ
uIKDgUfxk731FGpV2bykyCgk/PYwXq03+usK/EzrNpJaH8ZYs9VOaVGmP3jqaegRx6GW8UmA5XPm
SIw3lwun4xJmjohL53e9aljJGwvEIC1aR/OH4mpUHRSmRtqMJh8ZCgNQ+uWKadrmzehm38EmHIRU
DN3MI7MqCDzqa9k6C1YIbu6XhiEG6nVBtMwyESxQxMGhH0+wvqsouA45VMTCrzYdPLxRmSntWX7E
yrw/ckV005BgWYcOtfsch3Al0mojrLOoumGU5tXySvsU8ONnQVADMddG94bNLobvnBTWpBy+pGZw
tVClXqku250YaZVbcxeoWNayEifA
`protect end_protected
