-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Vmw/RhCPhH23iFMWe2tKynbGa36Ra1in8iTQ8N5n2GMR71XoG9dnjzr9o95EE3v6m8GvsrXWOLlG
ExOkzhtGKgEEIBz33sAwMcVfNN9/Qa7BDHCWIhdHJA2n5lJh5nxJpIBUWTiaIllTG7sgIJfyYNJ0
YF2ZylE4D02nTemXd4uELNRJT61Pbiw8/MduQom60tof57NIsW5/0VcuDSSEjANg4fEdiz9XLkWp
fp2UatcMxKF1sbljG+NS5z3ZiBD27A7kQNZQHqIrpL7EoU/yKgUU6UAmBzI3vRpVDn307+kp5MFd
e19PGTRA+84SbNdzpBRU4CgVuPRyOFrPSK6IOQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 9600)
`protect data_block
hXI7O/UbU7UwEhlzAjmkMqq9V5guwCFmq3jz7cF2kyi7VPk+m7DoAWZAeiWhQvDkgKEVQPn5ax/5
GmuJdnzxwqWIvoBkMa/zPLUxWhnC31KgZyE1dReuIAdW5dYGXERckI0rpjxaBoxg/Incwafyt/10
65x0q2hR0agSLZMkHCew+ST2NjutEc0lBKvJvfx3eQh5J00JxVmnLKuJvELyx7r631Ya5RTLR+gJ
4VxfqP4X/+Nhujg8tZf7vUV55nD9FeJXs/k91RnDNBfa6uQYGWEZxorgjn9TNLMteyp3PFXxBJa6
HcKbRrv98vQTiAIBrivOePIWM1ZQKVnJ+sz+fjzmGMNLLIPCQwERd6+yZSOwYLmYi9BwQegUCndU
BpHgP/k/cwQmGmHUjCvcGMMQBkNsIz/6418REiG2ScC8nZa4mE3JiGCgPdEyws2WXDCv2imeMFXl
dqKSfhW/so9CJSylbTrq0a7/cxm8KWdo6D2NdV4x5Qg8+rD9vd/yHi7KhMs3fpiTwmDWYYI/2uDf
FDuVzhxHfE/91xkJuvqIgeVudJrs+DwAHsNxSsNXUkSwVnAf/bBnRnOj0dyOwXOgw7C0wrdRGqhm
4qPrji3fffvigoMgH5zpTO1fbYaILtXb9ppagcGR20VLBWPAA8p/b1tCWFxbtSC1gdtrODEmB/uU
GyT2kYybpzzZAqilhd3UoLL11yUfILSl0kfi4lGXcr8rp4Buz2T2UApEZNvEvtaHZceLQCbPe1ZI
oAV03xr1OXW0qli+uDbMcXODow/M/sBoExoEJNLFzJmRLbzB1A95JVNF3c5qLBk7enrgF1MroFZG
j8JpIq3sVcO1nMblONFSZ6ai0jJF6OE2UkBlyHm9gQo2RooCoh6U9hTFLeVQMVOUBwTmKb842ZsI
NnNMmIxZ1zSnxqQYo6XvIifRUsob3jSbhq8jEfHYGDw+hGzNy7n3ZTaID5+i8pcrn3+gMeabbKmw
pdCSvv605mObY9N7PxCtow937EsZ9zlbFrr7rZD0jH8SmTOWwcpnbmT26sei5mcFdI3KAIQDaW1r
5fj5QL43Fr8vGgTDR3W52iRgPmwg2qu9EJT6IVtu5YOrAg75PWYGUoiv6sfOmKAqKnsJgaS23JlB
LAF8PIGARiaEAQgwi8sPV0xuxRS/U+7zmIp7Kn9vhpPutLC5kP8pOIWjKiQDU33lxrzLyxyQ3l+2
miTbYSH3W2yZzIRglZyKrKglonPnTGqj2W+Yk8dkpwv1ZuakJRDJREMAxjxLAulznxbTNAXJT2T0
7qaWAyV0QdVi8oX8FTfBrdPtErUfq3bS103s4AfixzLwaJCIW4O+6pya1/1kdfg7ErctqBh7YpPi
10f4rwZKU2DNtZvJOKK1lgBXVGgb/UoO6r/ZjvsH35KHfM37g9JW2BOCrFT3n8673Cgc2HDf2y19
2URs8yM41Z0hSYmAwF21XBjEK+JKH0nW28NVyAs2i8TFUfBDBB5til0Gi21cT8Pka/BZf3P4X0b5
1l3ywVmNyfqmlFmzMVmu5pERkr0qA00VFDNHTq/nuOX8+STklXIcjAy7TuTkCBmEx05SHWmH913p
/vV4b2VEhqfQnRYawQbPxVBsGh6xZQ2Go2p2FgVzo5LR6WhSHWfptrCjsBORhwVHvdNYkNtZoUyy
TfWXa8AZdtYR0U1UlWSlzoZ8RQaLOcy1hhV8PTNG4LCAEkpVtkgLq1GuBjRPoo6wsDlLFqgj+3pi
6cYcz6paxMPckWeF8lBcev2Sm3lOt2hlJur0TrP/WPHxAQquXzpGgZauli/9Vq4RHF6zEccVWSdo
AOuPbDK53ZxTHs/Ja0qYvFo/Mmyubig3GJstJal1XYA0jSKCUPTP1cwUbimLsbO21M3ho7bo0oxb
B6/6Sut5aeoNEVYjj0wjEn6hpTa1XhwJFhgAVoYmBhYPnFWxmr50ALTPTWIcoiaGrxqn8kGqnF0a
AFG2K5kNJAopDGZJOKdWVp/ZSkR1di5N9KHNgPCwQjIdD1WUrY9cZR7CdPh9w9agVD8m9c74TEjp
yw7MJuUOJPLO7a42VR0pf/b2gfZ5hoF2FOX6cJA1HYw5PrzvHNigyBBhyCgzuD3sgL22J+qQNqh6
EK7GHuHxzaL8ojeEef3ugM6iAHb8H7E3XhnPmU9s/XSkcuPROoODOXJV5zFa/+Jh0um/raWaUiu3
YwWyVk2aM45mbLVcDo3HzlB99CL3FoW5qAQHD72pwyZH4kai9gKT7p2ZI30WV8wiLw01OfADpFMr
gl7McSaeIxTgS7h77c0GHQK9OBs7tEvNGA7TyhRpdkZm5SLykPuU+NyqGWnRxmAOt55tQr1G5CB3
EcVP4C55WXRuhz2G7YFr0IYeNhti4wbGXcucQXymb0QiqlxMS8AgwXLAxZbGC46M99BwU5ETSa6R
hFgznlmWfkXf1w3mtjaaQgSvNSTG1fVfTh/c8UNFoij1atwU/GjhUVrjDipcxuexVqpmZtAD2h83
kfbKpO+v5cOrQG9j/YMvdAeYpprPWJ/+/k6WyYmKAncwwfkEJBfkv+YkamfJ95wCdUwTaMwmWjAR
IDh1wX7Byq7gqBUUArwktR54GWzF/DOW8PLvWWv+bLoek0Od1DxG9TLG5vwQ8l6FKmukXGHyZcz7
oxg87M8fRm/d++YOZEebrzdoyMkenn5sEEHPfmb2WZlGqEGwoPulsFIjRsxk5UFXWczKXcdGOYoT
Q9iXDsgXmqCap/gJh0+UsYlekbBG2CaicAuC0t8pWFO7ppDHPxp6ZyOKhs+wun9Kg6HOCEnpc7p3
i5z4JaEH+1+y+zBlcObKc24UdIHO/j0IgcPjMRBNmTo1KdaCA2hAiJwkKM9cwwxsiSmvf11nt1RO
MK5yMUpKwOGvhz2YtVcrX+u1AlyiYt5g4DM90Yj62685skDBzu9/WMSW0FkzlFoiPDGL/YsAk1qD
PxYe+GIky9u7H6+5WurzB0+vrZ4SGLoz9Tj3KHyWeoEpavHgKV2bJshv4QK/iF8xR3sCMpjpKGY5
Z69KrlLkJV2ciN8uuVG9o+MXmSt6ZsbQIY3L/msvC0cr3kBI/GwiyPuuTWoj4LYbPkoot5cTWkBs
3A1h1WudVjJxCwmeWmO/12iAC4Fp/XCSDhce0m0bDxX+YZw+xs63lg21m4SJ9fGd8QvBZF2kkGcK
rhW+nXkfuhNrRz8j9cGKizSibkIpHL703Q5bcUEr2nNY2KwWA66yciSfygxJoN6Jji9RQ2NBiaHH
sEiPP7vW3hbAtkaudKz0UKSipJO4PLsexQSZayZXvFN9glwAeB1Bnbnrul691VB9Xl/26ntO3ueN
CXdFjeyBcPwMqZrDLGWfMkrVAuXlpLSP87fGl92bjMOTiEcmY/UPjLFU+T/UV15i/fcISBBHPk9x
zqOc5VixS1+18I2SfSqB2GTERaVDBFRyiPI7lCqqk2YLsaJq/Ybi7LTaoryC7NFRXc5MsvaU/Rpc
EmYV9451g+E8Hw6513iYv+nkSEjKEqUpjlilQjJDty9s7YIKxGqaNjEiNMSRbjXUKPGtiUOFBlOE
Mk5M1QDJalwCJWOKefA9T+57GA/VImcHZlmptIP2NtYL4sieUsRWB84JAJNp9/fH6SdBxzqcVeZ2
TZegfySUFzi6a1WHATrUEl4li7yh+pch9dkeQd87L7AfoZG8POOuogHGHijk8pH727ZFCmCgbO2M
4Z0TNVpJONH1/lq2LxDViZNGK3jF4JfPvcRaxTS+1gIeam1wTiKreoWHRU8orz0T81Qw1edKVHG6
iU2OJKMFk1Es21TpdM/h/V+3/G4+Csn4iqHvcwEoXOJZ3FZ8h4zJmSmnglcQ4GQijJzZnpAUDc1L
lEWI7b6ML0sZTTBKrnMovKfo2zPCvEg1C44HCUVfNPQ8gEh5SR6rtOtWmfLwvJnVtmceyMGA+Inh
U1/9KBjBc3REQbU9m26i5hjW6wdUTjlh0gOaquqW8U2QdeoUbqm50g8mDhJg0eUHd/3i539KoTCi
MHCKqKeMmSzx1knuHR1axteodNAz8a3zXw0qQxsf1jB7gdbu7+l+/rZLrDVzeV82MsV7N5GkDD4V
9ilWFblKbrMfgCk+yMbo3NO581Nfz0JfHluDnENDrth1gkjNLFd3UoEVI/tccuIEZ9SbPJ7WrNPu
JYGgly+ajtJkTfLC9C+uzK70/SlyCSQuxgbfJ8FCy497X485LNdqdZGephNJPkqZghOfD8l1zUZz
tzld9rCHeZ6Il/k7TlZZILyF0SK/n5JVwG5WC1fDrLpMzzxF+xJUH412l0+dlWz4AZA8ybY07R6a
sNDin/6pLxNz/IgyE+kInTl9KJ9MrGRSobu/3EOeKMW1s6b+uVjTDzxQp5YoP4Hcz6mv+Gda9DFb
bzNlo0kXdYSZJBKo4OF8PMCE8rzElp8JBJho7N8mfyDdPFDFmVYETX3mJeNSUz3c+Lwvc0Nk0om8
/AcLF+dvrCKX+ZZSH370VssnQfB/ontyJ0rYR1wIi41fZ77KRzvSdZ70ZG8vc84rNlSQbZyqz2jE
SikZg88M12hcTmC0KrZnccRpGElpPmVD9nnOmMUbvB4bdv5QBUh3ChKgg6SnafQbJdDgHti2Lg0+
KnoaISs4giU9fkR4bOaT7mY1BiEHLQFjM9hTGKd9LPXPUccFKX/8+QpEyIrWxZAGLMcJbx2K6b4k
p61yeRawsTC5lvYP5fIzpw/2c/FwFN3+feKbKUT+AYtwdhrWg0JrM2rE5oTsBca7Ha+oj/FOaJJe
0D1wStdvE5cvtmsX42LsX2zS4v8P24+LnY5fZPtja6S6n/W53tRn11VcvZoeLZb56+IyvjInCfAM
KZW5P5kY6Ve4Jtbp1MvGz3H31yYDGc5NHreTupll4n+gzCR8Q/NWecSaMDi3pTFWXc5e40tB+Ah4
pPvfsB8ZHsGfhNzo5LSytXqpADwlxR60fruiqFLxRYuGoMK5GxF1vMVMBKmBNFRE/7QKeQlOGMCm
EcVjrTsW5zvowaWQrck3YEQF/TWhF2etfYcatGzg/vhQG41tna8pFWCnvDaPy8P2tD9YvQLBLD8X
wUHkLlyH8v0mvRl1aYo+RpCeGxW1i/RpoDak+6B+Y1SaO+xbzeNJiHK0CeiDzAV1rHrZdacviIpT
v6uCT37Zsbe5Z03WSHSAAsacrtG5EobsK8+wu0d2Kcdkokq/mldWgstBX4OPAh6x5XJTz1vDOYVq
EzY0N5yzc9jtPGqZsu/qrmVppzW5rqJWcWbs7mr+EpeTec0Xvu+AMYUkUTrqvpKM1eFlyEObk4vt
Nvujlgn9LkThC+03ZWYRzKz9w+ZGgLarcbxlmucXpmxUBpWP/128lHmxyqhE3/Hx7XbxpebR9VJt
RF8mmkhoU2+wgzRoNgw8zvVEHZTnt1DU0yoeNxGjT9bf68BAsG3tvAUHm4ImQybirC0Pi1jIlXY5
NmgeLKl0BUxqPc4WBiJlXWW+vAGGoa2T3cBkD3F4yvmtI1zldQQ0Dsvr6+dO8Bis1iixTrH+B153
6O8LO+Uh+hxZyyi3rSpKdz3JIimYLwNb2iZ/PBgvEbzNqrc2+E43e/zN89sv7jik+G+LUtWUK57b
08X+OMhnJODnqag0Q3BY4+gz5govDC8kOitMjDD/5FLlu1EcC5MUvIOEq4OTqAKySUGmp8TNOPyb
bsGkC7NwXR+LObCS3g0EXBXEExK6pNTUO/kpitNYPcozBdujVfKFu3vi6Gm0m6hSUAxPM8DSURjM
5luP4IIvUyUqcAaDu8T6qxq5Wsf+7gfO3k8Wb2L6ASy4AgY0Z9/NHB6WVp6l+QBEfQPxQjEq53zE
K5GSINf7mUPPAw6pNfvb/I4ao7kQg0cq55cLYNm1Cl1xorgqjPFjZx1zyKVxUwzi8HsWTnafiVfV
SCpdGaJeDQzDE93lkBjNurkgIrJflARmBN4Tqt9TO/Y57jh87FegUHeHflZKcSxErDyUPs5mcrFT
L2ECamAleThJTDswHfp91DglRC/TijW3egjMCRJq8AqEZOH4gmTyif/GAwSlHqAhkGFaPTwusVR2
tsUmLkL8yfQWxUP1s+svhCD1c6vbB0NQeA9JNhU9JDfzyQO9iWtuBNiFZwXLjhcthAMvxyYhbwkZ
WW69M4AlxzYkajtgU+Voc/TgTQts0enwCxry3Yz47Fm9z3wkusFhlaa6p7JomWzPyxYIxup1K129
yfKk9fHz4PY2ZNmreVMN8my57c1fNTex138EtYNREzTYoS5AkdnJFgP5U+oM/+IH3F6NkwIpoB2r
uLCRGKBFcDoOFkMFtD91+U75aFTOXvkt51iwyLp79OtXwE3g1Yu3DQwJ6eM46DhfpBiAPK//115L
NhUJDVUSAKPDhp65wXEQxtKNIPlbDv0vcFWxdRkvO9MH95K0qOJDUymBJzALSCDuk5Ad3hwiBSSt
78X94Xkd5PL6SFndgjH+1HvtKgRwrbjmx53428ZIb/QQpq+B9rEBYClCA0c6o15M3FDWMJ/fjfys
vqAxmbBOlb5hUhsvp6qmr5FKNn91xlhddoJj29s876RR0CfZpGRepsoMVk4xMNFpm8QD23l5iXsx
Dy6Oi+fPvDGhm29WIQrlVixDmM5UPiwd6vOZfukS2TA40RSv+bCaF0w14J46FFfMCvBIMgmjMkie
V2oMUde1vnAEwtuSMlFQy1aWhZH+J+vwSnOHuwjfIb+0p57Z70iO6zVDMbOqh2SAlFOx1ck6cVEz
Vo42XrssPScA2B1K2lC8CHO1BjtMwvlkQHl4uAEa2KjCIU76SXe31DbeABs8E6pPS8uJoSxRXtjI
aXDG/xmyYR9Ntxq5Y0C/b5ajLm73UyVTI9hXlT/l9f0F+4hJWkND2BxAdtiLYGep04yi4meXxE3N
6HU4OXbTCakmzdMaKJPao3uDWLMCTvvtddeVMhsmqqvo/3SwouwogWo/ioZSayKpckZdSzskRmeN
zk5hy93Y9skj1s2HBjzrDyvJIKoYprpwe0MMWxdiQzBc1E3vEUFn44o9Mc8ZTjYAbxCvBfknZwOB
O124xZbdfO0Zci2VTir1v4VtX+JpUiHNOG8J/MrHXS6PbXoVjekI9P6UlNw7e9LpDObgkbdorS2c
p65svzWP5qyoCWLTYsDOzhTho/uqwrsamqcRAhzEDprfOWGgxQvUdyUBgXDafqrGjuWIGcZxfWV0
15rzWfmkWQP3F9XTMZ6i7E2cqQl4i8b43x4xxdHsnDIliZ8N2vQpx2zpWVwMfn/UFqIC5Wu6ewoz
NCNFzqHSKpZWNvPn8hj9TGuLLPe2/KG3qspjS9do7trE7nDLxe1RhZBiowPGTZxieKnpidqdZhea
FTP93GWJZ4etPPK8mbNJSIo1f3cPjirRVTvXzsGymv3ePaIjOzr3mXgbVyGGNfM4waUaQ+DfZs9+
aVhUFhjw5cNeZ8Raz0xZVau67K8KwwLlNEBZ8pOprdtHiVPWrWJ9i3CfDi9S+y1WVupfmlIM9deQ
0FNK7GdH9WKBpW1F0NkS592CsIA5T6GYFeSNLhWZ+fmFRtd3bvXBD+IjegzgUK14jeumdDrIz/ce
x5OVScn67pcAV5IhJjc7XDolnO65Mu1E/iD6EvBWYuWwdpgzvvbm3dmxdIZMmJV/iOWYOyiy158u
2qzYLJiARxY3Bjuy8SNqbtsCb83wtuDZT+o+F3DgcYQ13+rrK5PJhns8I9mJuVBnVtYC4tzkZtmz
lTsjm7y/AxXv9OgE4XgJyOHLHV8AsNmIJmvXJ1Wqc3urTDdiXCNDAhaIIbl94Zl2y69nnJsikJ2t
QDHE4TeNGpUnrh4WMz7pm1mNL7ZGSfOS7Yj0TerVpojrhDjXLLJKVrsr1kpSPE8I2ocXYx+2cZ6r
9Tip4eDPrCFexj6jjUT6P0yIPoWQtJv2Qe/88fHbVXwrks9Ty+q6lAqf4ByQ4xV0Tuh391KNYb2Y
0qzZZuCBz+89mKceFrnWP69wwOqn7bMTvDX30QV07kj/BRu6+D0fW5a2NmMgdWEn5XAyPYCEJMNe
t8oyBvH+5Sm/t24qUxDNzRtNY9fQ+D4xRIzAKZCtjdubxK5S7Ng1ldcT9QBalltFJfqBrGw198Hf
LGxLMAh0UvyKaj7jBly4FJlj/DJO8C50QOHLQ2026U15TBZwgqocnSwUaKZcI6uBGQ7miW3XiDkh
k9wK3TLj3j3hfPRjImsrJcySjJ7Sw2C4zpZTthd29F/rWV4aQ2DlvG2j4mtSCKNofHtgH9P6H3ws
nXwINO7ay1wZ1gMb3BlLQJfDSMS3dORNWqh5jF7EYoy203Fhd+nSm8fMXjfhYUNN8fsm8g6Yy7Ep
LuZfeGrygIXwuWNmRHoETIMVm3ZjfEqaAg6q2E+QOb1M2fTipoTvmXt0IOuFPfhvPlnl2GBixxYa
uyNNFnOocTz3M+IHabWz+FNnlQlAmQofHPYqbTLgOhpRwDqu/n/xKc5Gkafymbtl5bP6ZEBscq4r
fYWgsSSjq0Mg3veVk5ex3gruP0IIAUwq+qO2rGDCObBVdXp1G7Qzeh8mMf/voukzsvm8nq+Aa8N6
oe1D6mY7au4cFgPpHOuXfxBiQSiPCQ708rppUiGIcf1axCIbpr9i9yy5r2xXQX5qOAjj7skMRdSA
o8tBhb9bo+9EysxAo8AVmd5F8V0J6n4vVwNqN8A+Ys1HYozHnY6QCujhPzPpewfZMUSPlGJ211db
L1lSW6/z29PA/aeWZwg20E2cS8dpT5ZSQ+Q0d1T/KbLGyCiCTZk93VK2AFq5DdY6OYPbt0VONjYy
27no8B1Qul24Np97Ax8ImXobh5gsuM0YVS5OSw1rYc1461tNY5Jq1g7rdNWIf7IozTx1rKA4gx4B
mtlygWCzf7A74xlmFpZu1AUi6ASz5WHjRZ/oieUB8pgzNLy9ixp9CIEieCl9nS0VLIuafjo4527h
0rvAMBIcbSDvpGpJieNsxtJxJOBQuBOq2fzRHx/LvTlffCYBJu6HP7GMp6bJFtCuUr8TkV8rfk2W
cmr4yOp0+Y0sqkocKv9oGM3oc/5VoVoV3fPo0fPmODvn1j96iBJBaXqt5lOPzsI8lbhH7zCpDy9e
hVxIj2FdyCJLFPbm74/IJ4pc/rnCdOJWGod5G5YX2V2zGKD2pbJncYNeXtBHtrhdLYOuopiXME5R
DXV/GAgSW+z4R3PQRB+i0xQeVle/3D1958W9QJLjY5xQgTuG0F4qUJRUDj7ge+kO5oubPfK377oY
RWiiuTQdyhVja89CfpGi9y+jJFS4GhmsdB+ooqXw6nkoB9aXceKvKdftySNt8Em2IkmAmM95/uua
k3hGCjca9KXq5QBwzthk8+tvXvWdLLiMmH89EoEmyTkYKcLTrDv6Kq802cR4EYcXXkxqCju8zrp5
jC/gCt7kkA58Y+KLTRLHixY4sP8ef4SmVDKRTh7XX13WF8Drl1xGFrsftSJYLSD+M+ErXwkoFAb9
cmhy2ic15/Dgmt+rkezCfJVykw2nuOdsLLimVaaLv0V6XffzlE/b184sRaWMxy/pxrEWRPczMFe1
tLYEO4zbaKqqL4Sj6HDvZXvG7OI1y9wwF2oLo9/xRsVpbvID+YopnaZlrDRd1jJ5AvzVzlPZBR97
hGe1rMmZRLhoX4y/KKydMWKzFMna9WiDs2rzP8C2e30aYsT7GMdRYZ/VlJKTahYpUutbb3Ftof62
r9xjOqeZbuevia7/TMT34Bw6Z/wwsWl/18u4/r9EWtGyzgZqZilH2K6djBsleogT5DJHXbxD3R2i
90thick5YKMmiEohlBFpgH9QDoO2jPjsgBUggGkUuxkhhGHI76IIR4qQmi/6FbZtHriAimRkaZ0x
Be31pIjC8D+Q1L+K7f/hXfzdqSykv7EndDBsldUinoapnPcMQjZfCDKNLWPdV3LT3ctH4fFWDqQp
vw80JpR4mCgktL9BS/tAizk4cJWpBg0uS+PIqRwpNwszPdZPx4p6TP7BB0oozXQTo3yf7Ntyf3RT
tjCREisp2iTWgurOlHD0BrwUcXO0XXOb5CafmuBiH4SuRBONIljMZrFbG7XKiHUwxvrI4RKVhriC
Fdrtys0oOWKzD8lxBnuOSe37ajukXDhG6xLlycguStfDjsDuoEBUeu9I4QWLivVjaHc/cGwqQEIN
T3G4Rs4DWAUmprUZd7OFPnqY+7fGrtbEBDORfobQWtCeyJQ7gKKJI5apTtauhC4pX8TInb8KFEbi
xL0m97E8uJJ5gYgr4yjCI4DdpN1iMygeQ5kiZgFgmguCaxzRlp1CxCI8Yx7yOJuNc9aWHe3Cv7Qw
C1iR+WHzhhwosLhBrh87G+saVM0x65xRnnvKLPAqGR0Kjhn22OJgz7NH72rCRodgRzNqPvQRT6AM
anZCpPawGbi5U2aQi1Z8Qto+Bp51CuVzTnJ4YfWieeCC2pPgJSrOpNjwWM8J6d+zehd/c0Ct67ac
yx/qRGH3TKgLdxt6xXXqTfC3P23mmRnLZa44Fx1iZLC05Pt7sRbMkdH2Jcv4I2Xmss0ocRWEM1R0
EQcgn1QvsqS5F7WAjdVqP21xMtXzQm5v0mpz3RQZK9fSzAOXS4RPK2JWLbjnOUWeh6TZrAEY7fTx
96doTDGnDXGDnCQxvkBcrhttISeqvi+192QOIUx7Za1yRo6p9nHMOckXEglkKa4LmPdbsOKXww2P
fzn3W4/lowliEsO6vvKRx5JSnZN3r1R+rMceFSacQbQOWCio9fR6nlQZoRis2YwcmDQNGgOJvnld
iPT2Maqr7l+VMXBpykMrqFgDEX5kpTAxAivZfPHssm1Ll4Y7/XYmpKWOxAGMZpwbYVUuSltN88ho
3yZ8UOMF/3XooxZvzfJFNSSOzE8+zGXvLutcagPcvEG5XbyX+w1TIPHZCUwwhXbsBfH51L0iMPoF
aa05TDQAl1Q0D/UWTopHMnqPR1Ykxey+LN98vgUBWc4pB0SvoTdtZywJftiMw4ML52tMe0x7sRpE
zopFjQn3dioNrsGDi2ITI6O5zrcp26yHhq//IYGj7neWWXlIjmJLXKeTjqTMvVl8fUoGAi6EtdpP
e2Fz9Mowyss7O217yJdMElaLv475Ov58gxB8nTZOv5eNK1bnDXqCCTJE1h3WTmmnU+M2jci/fGzJ
rL76Xp7QCgp7ttA5m+Uv+lF3YhCbKdp0LPukvSjcfVpZaclc7RJBkWcpZ2TMIiFGebvJVg2kMT//
m2eA6R6HnPYXWO5wd08I8sERAOqAwH88m7ovRRtO7wFHrcBC6vialTwbsqgNtMhi9b2QbBqZKOsH
GL2tdzI1ekGskTTk8J1/2aXYG4W7Ka/rXT784mpj3rCJHctuZBIldn67GShVQiZkozPI0Ig2wknW
EUH4sHdNiXM+8EVaHWHfJMINWtTCmADuNBqNNYpA61g1l1/VhHMJX5apCUY/a4tVqMa8ZzSrKMfS
pAHUhXHxRWgGTidm5qhs3pJwgR6xMGRLykDP0ZQyAzW03/HyFg6AEA7NSOSYIWGCImJhIxuM46OE
Bt03txlTscIxdv0qWhT8OncaO1jCBTopwMy/rg7UHzxBmO54jJfEzYXJjSXfyFdIsbfk7jTmN/ta
JKteIsCYFAcT6dX/gyem6//VaG8BV0uxHqGCRlwuV20IXFOaMDLj3dbR59ygPnUsaRaFv2S/0Sob
4fIB9GyTEpAeLKqA1ABXl2Ctayf/FHWDeLWyfjMbSNET1Wp9jCocplfKQL2F9KrG2IGP6muu96xH
8fuAqeqYybE3UhmuSM0IG5rEklBJv+Ln5tOZRgRqn5q344InDlIy1PJIWlheiaNpFmeuYzpgnxxf
5cKIzqwMFa3OLM62YXPXvp0K2nEvyXWo3+sZRk1wuAjxxQYnFVBa4ABydbJNGhavlNtJpYJfA4H7
wSfU0uveHpuoOvCHqH+g7ZN5jTqOo5MsmvB81RsUYwNKdpAylcslTxYwGG8hqphptAHPEZbKFxc2
4fSInrd5L60ePfCEcRYadWUJqgx13ObzTeocjHK+Mi5ZZ8tU9QZlchhmHPN2JPGuRha+UezqiTV6
AtxwyHBaZvqPGfj90eu4i20cFqk7VrwLhLlf1bZ6vUIXhBRtot2DS8DOSL/ngQs3BxEB44f3QzSO
U+k6bkY0TnlwPL6fg2b+yJunb+ZnBgbMWTFBf/OIrCQFLqd1liy99nMNk6qCiFwJr6Q1cDtw7vsk
/2Hzjc+x+TR4MFR5yNse9h0LlhsUpU/ESE9GlVRAh8sce/J09wNwkMOIBHNtJsvo5+fjfBQkWpe0
0eTUzNTDPMVNpfpOWpjhIUam8ib68BlEqLGorJ8oMPn9QVEtT5AdlUXU1966usQE3SGTFmYUtd8Z
U+4WVj0LjkUfsLSJQ0fuUIycFpyScckO4vFfKZCApwGX6TcdE403cVZXKPMeonyVF+IMzekdmwHJ
7dKEaKFZGLjurWeKw6Smllj4bxhtqVvbHiheko7VoeNuev7WSDl+vIIew3Ykwj4R3Cg69nUn+GUF
OslxP0/FTplU5Ucw7NXUyDu25kj79jBR+ZJz9P/26Ae9IDXgaMooN6puYrkipcoowlZM0SeHq6lA
kQTdcBw0k/VAtKr7AqIOIxQnR2TXnYZjzbzE/Hk3atuVdi7EXpfQsLSOPEK9hHFlCgr19BkZh4Eo
3WHtNsOiwP1KMcaZoohLo15yBfuW33yAavr+Hq1b1ZxwGA4mvhtKvru1hn5/ez35GHCNf6pUr7YH
KGFhwb2DkeyzqG5u0YZtXtiNDiJ0N8NR
`protect end_protected
