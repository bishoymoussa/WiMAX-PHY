-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
shiwr2MycvCXxgBx2r0e515eLMG+2XPOhalm5rcETQAGUx9qmpdlK0p9cPJUOdmqlYUsFeKWtQYx
EIj1bFFejhKQNaiPUJrDvJeuzgilWNJXxwMq93j0aQ4MBS1YPQJq51oUVy9rvxnwtt2UVKRmRwvU
tRSMEcncAvjJYDeltvrTurzHtu9PHIS3qnPhlDD9ODhsRddN4CUgvCIp4C6TnKqTOJua1juh2wMw
drh+RvD6HWFlm06JE/tAa+pO6f5VRMelOhP0H9qRFnyuM1nzOlOqMz7SiAXNmsz9VaVB+0u5Ew/C
wPJ3POvJ3Dxttk7ICpOzX4wzM2WPdDMQLPj50g==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 14528)
`protect data_block
mnE7+7bJ5uXqqnIy9IoX555LpJBAm4nr8frHycdFOHAYNRH1wk1nFQVXpTJv5WBWF2nSzSFS4aqh
ksWtvlPP1aI3lz6YqJdq44mtIAvFU0MQ2H+FKkqKz+oNN1hcbWAFTjAUtwCCBc2SU9T831tkV1Cq
Kzkx/XTXgwzcH65m997vQydKLvcCTUOOfys48xb8LUZ2v/sQmdTZed3BCc/UDUyAQ+/3D0B/N/Qq
tWRSs2iaXTDCIt8Fz6aqk1S7njscccafs1g/d5v0jAkubCL+MxGECgCNHryK+zilXdDay/4/CBR4
0QAFZSmR+bfyuFEvQ1QZ764vuEWQxj09ExIXApCMe/IsDUXUWtIRW6gImA9AVPXMmslMf9g6j5U/
THjyt/avyl+c4+dhqtCJ1LsKkj4Juf7YRq1y95WGaDp4d3EWaXWsnC1jmcLZKFjmE8bmfRmgl0Tr
ioFU2uguCWJPHzE62aDAYCyUI53hx+BdmhsrQnHMakpo6POFYh/P4Xs+jwCe8iLBIyP4rlcV3MUb
bZKrRL5vC+WUzf8e9FrGo2cchnMA5Y5T+WOZ1C5W/6fVQ1l8Cmnx5YzHaOn2btTX5Un418FGOJll
1s36WPF5j58kbEp5j08Ryiu5ROUOIGWSHC56GZJPzyfC687UeFZfgkKLOy4zBYb9jCEDIksIEyxO
EU7TvwGIkBEm2zPFhkKplpkRIWq2jBb8YgPeeIH1p9u5iYOXhHmwj+mFyXLcA2J7/BSd0ItySFMs
5P5o05QOgGVGAi8TM8eMJU1ihR6gE6WMmNXUnZ3sKcYJYieSkU7siJmQ4zAzvkIieiVlIiC2Tn9f
IZRBnG5TcqrH4IOYzl5SnFsWe+oTEPW734ycQTJdAdLd4kUPEh+nNchIfvT0OwdZIQaUcffuT7HK
p1r5tGnq7+E6N5DUwHHMaieKwskZ7/pDRZJ0ndPok9qtnp4QMxe2czxn0lmKMAVTNueHfxJxYsHW
c9ng6DnIyCOKgdlYyrFi3E+VDipw0EzNFu7Enqjh1IfN2rF4EDfch3dIw0nPWiSEAuNxMDLYSjIp
3icjoNT7xJL8uvXArhFHitcqWk1DYZ1Mbmvk9Zk6EX8nxmo8jM1dQrUJqCN++pd5E2VGqwW2/rQB
CyqjX9M+jUokWBG2PbMeopOhSv5LKA6ZKTV6zCFxnVVun2IRwbHt0QIrtGpgpIi8jMnfghtCfilC
0MX2E60HbX0+3x9osYkw/7pK7y+lc3EZ/NNTk3tpMQtztIvydAjOkDdEa03JGeYmbJdme9M5c/Dz
ehp1vvpCkjBZwWvXXn8ChQABPRYfh4vl9wKDk1YRubUpBqrrqO6pi1/5+1BCx4YXyKW+shFjmIdK
nb5lUO4+sSrJdVVYFWnOSppgfvZKEu9Ud4w+J3bnLqPbmda3aElDtH3UsTlCeZx2iMQNw273mABG
IyTBsdXDWn1CpfrI3vjCiRKTX+8lSFB/Ek46LVDdeYEdRvfjsVAxryHyQ+GqBiPcZWNlzPxSeweX
i3Rmg29N1Gn6yG2JXXnfpDUH9ETaSkdYWnmTD32SrunR61B3y9pyJiT7HqpWApitJ+fG/HTHs9jH
vBHHrWh0zrgNNHn7r9mrk2se2x3txFejnMBWY4QmKjX4U6JstztyLWLl63D6pOWUM8JNmhqG/xGB
JHiIjZAkbsIrN40jzAjPb8lDAjh2qrknV0k4xkzveCHijA7RoQI80dcUNS8X9UUKThFUNOcmVRqB
j9BoB9rpCWSJcXkQa14NLlA8KomYK8FNB5gbw5DDQ+YrUA0duZKR38Zga4/GsVOn/kOwVtcC/0cy
CSTc2j43HS5exRq+ng48o+cLbxXuZvIGZ4b10TSflVrCyOS9gF6Im31Alu3lUSjlYc3Dfa3qm+5O
xFzki90XgBOkF4KmKxPDnK5Ymt2VcECifIjzqWiPt9RSi9QPrY5kTwlHujUi/AzD/nTC5UB/meHJ
S9mG7yWR7rCBgV04LhtAUP5B7a7G7EMjWnerHy26OYCiyL7V1/TDLRmqXoRr0hhmaosvIaW5HgQd
5+ON9W1L5n6eebp7g6v1ZZnUqnHkpiX9VFsN+6NgokV5pxlhfvx2SHAlQ6r1453t/quev0pt4XLD
voIQAXH2zWMU3wPUDGV6mxKbF/3/w74ngtM5jh9sVKRNasUm92ZRd/FZcLBmOvS1cHS2LUA1aDVT
0/QRpKobIewur8HhJnQxaSrMr0jCrLneMpNbhalNPZ+PC+MPFY+NUh7JzK8fAgATbNmyseY5iev4
mPjJVkqRTpeiWv5U/GuRf+cNc99UiBEHAQJC5uOogpKVQyvBUEzYWJ+CN3DQCybBrQbBmr3s2uxf
4fMiP2u1zJwQf6wGPwwQLXgYrOaZhFhMvYH5WNj5oHbWfypY8mNdpaR3LiNs81AXSMUan89LdNNf
3Y7G/cCSUJYMzC5uBYb9r/cnXbTaWaShCRxGFddS4eHPq9BFTC5NeEnNya/31C1C208s1JSS0HAk
G0+8QlZ0F0G6gjkAQR8i7PWA5s6pyeBtDAil8+uMPPP6AXZZXTgvpeph7H/CQCyyVxP6DfalQhi4
4gSjlLvYxe7eq6PQXoNS3ZjlhivRLxNdrDJtX0Wt4ipJjBKS8y3aKXGFrN4UL1crtJzvvJsvX4RU
2qxpf3gr9XdxfEla91Q5RBI8KKwoogHMUw9xd1Rn5xKr6rvX7Ymx0hcB/LNiQ5uJLP8XD1Sb6rcj
drgc5y7cfiJnis1rHOo2WJ5u3Cz6U7J6b06Arbdt+62l8vRKVbnqZzQDp2UVySemKozOb6a/qLCY
nx8Isjz+MEwOsWKV7JNGB4scaK0ylinj/i151i2gbOfrXOn04Uj7T07QP9CG9hhoOeaWnpyMwZ8F
Pgfzp5eHhL1cj+cb5Uq4CmTowJZuTOQji2FsVzn2dZLNobzyCYoZmd1qoixwtPWjp+D9PxPNROmz
QZIE4uLzpN2BQ34j/p7L0Pky0fUlVaHoJZPMIqOEfn+NFh+IRVU4NdoQi8obz1nvU9KtoGRBDq16
n69NmkwWX6hRPFhReOBtNc2c+yJ2mA9Xb+EWEGaF0cTrexRaVaURFbnEgcZc6lXEkEokJVuNMEgS
19zvvjl5fSWGijkAIBYmtH7Uyom1Oq3FPIMZ+myddc7Dtwzen5DTUumRl29kyqmHquJ76ZIPMInf
csu7JMQ8R6SWDAUJegJX6AgsXt7aTCuPaD5APmHmRG7kilzix5vvtxmdfeERnnRM8N+N3RNllcPn
5baOE4XJag1s0SYMGoeKmsm/uv8WSnmMLgFd20RAZsSSQMxs89/F7agOCutvXM8QUj2X2ZPHJwX3
ii0XOiI/xzOq2uGq++1x3ZdYXV5g5KJAXsEgGY7BZfC1BPdpV675Ocyj9tpjEH6fhRpuQLTRzD7f
6CiHuB815m/byiplOqRaqHA4meH3IgTaK6Q25q7q99IJHXie5JP9vcoyvJ6ISzumy95uYigBuPt/
MjJznH/i52EWRncICQIqqRFZqq8KRXo4BFknDoFABWuQsFxHkE/LKiHfnzuDHCFB4l0h0PXAgkgo
Y0Nm/LfyYeCvzD8FwiJOV829OgekK33xDr2aKTud56riWuaTLBIi5eV3aL0ZGOu5P3UXt5ePbsIY
PCNaZT3GwfapkKET5jrBMsLgHpODwZ4B4va62uihfr0H/X+HFhUsmW2FSAcAaijMQ42/PHZRKHLP
C+5OK36S20ZuoAPIEzpxHmEdwT1ZzCkj91sjksr582w7mpY53OYDJdCtY7SwXqXVAEvX59MPciIN
rXwDvvx7kTjjFZJezdBjW98QAaW+aA0mR4WWu6+dLSbuvJzclaivzajcEe73ojmZK1vXcnZnVQPV
fLOQ7qcnuneV7oDPWS6sKwbth5e0M1O8+8SN7ZT8MktbsM2/Ij70P2V18bZ7FSV7rGbE3SP5NA9b
jSPkeLcjlNDyESX1zTydfrysom8U+KGp8FnS9pQe91JQXLmPyM6jr9mq+YjpfdR5pKMZefFrVMLZ
xdgPoxrds/yymTvTppwAsbS2+zfRNwjzpKkxgwVSuxj7kkxUYwChRl3XuBLh1Ze4Du79KPq9L2TP
i0Eocoj+WFbCB9WpbABrIDVJijLcNqo0UraDCo+C3qn0x69tRkECleCA/6W5PLmbHeUuj4tobaZi
fPujRPIV/pQ3puiU/T4uxEkvlNBXFS9nOERvKE+RnNabGFcjrJ5QB+ABchAIdsufo7fl8UbXjF0J
rgiceZiSZfBxDNJJ7zAD4ppZC4GBw9/PTJLrBU/TqhC3dMCGEiFesLedoy9sedHqFp7XDRG4ws4J
3Es315Ugp1ZMhVAJ0Tumlyc5gFG/wVOni2+ntZvnwAqJlQ3+29Htpbn4irIrpddTDsTSl2AKhgPR
9WZAgZk1oVb80ecqJeeKsMJD//EB3qy+vQZGvCrRa5Mwk329DO+wFGCpkoQkdZk0oDO2MH/1Ig9p
hnatyO1uibrR8bkW5tK9Qj/KVAdhvfEYwRTmmvEsCl+isxQgnn14zWI2KpsyLPPXcCq8D6brIaW/
XoS004eQPKpDRmeN14SMYid6IzntWu0yYs6cOEO+bl/ecCqBe4lfrzxm+lj4YxXEGKQkYT2Zrmvk
xg5qnP31dscYK6x958E/bue27bqd//jmPgtJWl+yqzrOm4e4TNqjsodmQDcC6EB3EpYquc0gUiHF
/mqah3flFBC3di+Tyh1eKLKGMV0i4n7FLmaryRhyIBTGg2QOZ3Cy1EA8i6ggIsR1KvSNwt5weB3U
FBstZmj/j6K/OYd4h4zGtAXk/rQMzWfDQjuynRq6Y8+CHBYtcTRCaZTXnPNIAoA4z/708i6YFFDR
9LkgLh9TvHWcLYbjJKAXJphZFfn/4MnrPKOPEIKDUHqHcg8Q3KnN/HKVAV35ebLSFJeeS/g0x3hz
epjmJbd7LkE99lZZ3sBbZFUV9ZrKWQKaVUR2znl4pa2OsipLrUsCL2mDtPb2vti+pqcoTxlqXNhO
GSfAtOPzqGWk0x4wdWOs9Vs4BNCcySdQSuVuOfwuKHgJUNKw8mdwGzWVh1tu6DwtmtUfOQlh/6IN
Bowagya5xcUhV0bSXcxVJwuisgtjVIrkQ4Z4Jw1+KIQXrK6kTu1jMJTNYqN27Gku/FNSUBBedV5f
L45PVmk2w8mDdGTArw0dN4wEBkscds3s7kHa3HbkMkt2QqvVi1Y9gSQpmWfTv++SD/LPqgCvZgVQ
mYJf5jxLfv7lOuv6+tvJ9D98kLKCHqRw4fR1SXLWEkVI19J+DLOceakkXp6WCTRYLmeovAv8e8RH
kaOz4inn68/9rhai9n0clKWDEJJZR9bo+j6Zs8zk01Ka2NZUu1wY3I3NGlwI2eMoPqBUQRQYEF5A
kOZ7FZ7wQyZokipRYdZp5lvoTXSe4DhrU8/4ohLLEDRS64xj6XyiIGAs46KDlhQqZeJeGWUfxkNG
PydYvFUgmvqNApemMeqDEE86ekKFDz/lnyAMsmxlH/8y8mqQfp/zRJtlJtYRZcJRFq7qqE5QDH33
FXn6AuaZuTTxLXlNWEU8zeXhcwTJNSKhatb6AupYvx8KYcgDm9pYFIxLNWHZ+Elz3Ojyw33MihcP
h8Xf8aT8TAzitk//qpGBoNaYpWjxqjG95aPSyViNVSjuTVIMnJ00MTUXtIUTLVLsSUkTLPnQty9X
T/lxxDWim8S1gjMElDG6KBKN8ttL5LrigDa8r5EAs/Ptbs2PuPnkwVDoizwu51SBXZZHqxfetjZj
tuXAy151ysFF2asg6tVRRpQdCQ113qPnl8qwfbWisZfk8qr0AX5DJsXuNcVY8YPV0H2BW1nDuesQ
8nP6VJlFsuj7Eulc2tCyuIuEWNQlkLNPkcYFPCRC3+fDusr2XcVznzIsPZpnHNWiLVrlcwhn7+2w
90uzMiz1z0QNOjTRJBjEFltnrXFfI2lOpO8wIqPYd0E81e3rCS1i7O0aawppBfI9/8lNVzzeIQ/d
pmrKtCH0Jps/tLI4iiWUrJfZ5bDgx/DJNhuA/CTqczsORfXYhlCq4ZOwVgtkZBAnCrckQtF6qvsR
jcdBtG4ph+0BPHrcy3oZ/HtHitf9BRXKY6EWp7tLknm0xDruTeq60lpqtTr/cuY4c1Csry6TGTyM
FEpGkZbhdFkPGciGBYBG5Etb39wfjNgU9sBNoH/bxh/mTLKlsklnuBPBKBaZr1w9dNkiC0WJD4Ei
dAlKK/n2LRAW94vvCyDLNJnk+Rj4+7ZKVqMTa8nwxaL/Bkfxdmi21KvNbz3x4V8IT+DXFKRiaMDO
k5g32KXI69EvN/TAZ8S/+HIVqXXwAdB8vNQR8by3VnobzDmmbmt6jcczqqhNff/H1y2wLAs2iUSx
f9ovcoJ7k3uftw16COEj0w/orFT15wloQMBC4OIFZio/VBfxcP+k3DKCdUPjOcCpEOuY1EiCFPiE
gkiT3axt5sJrgjus4UTbuzP77ae8T7H9Whcaf1Ppo7sdkMt+qVvO3ubEtvanCdPsQ2flnWiYZQ3M
q5YiozNl4fDm96sZvzcfnj9aLz+hnnEY/XTI5qeXKslQXbtdT/ve16f8HJh34cK8wi/76f/P6MSO
KvDd/21qhaeqC1Bwo3qsICkeeUgG7h6zgNIDo1T4L4xMVTYnUDC2EhIYwv66jPH1HuM2j5OM9PfM
isWLEtu5Hh3g47dLSepdkOavKKGZiYu5lOQOJ1w6Po6pCt5XfiJz60pXfKwE0nDx+XAkiVLifkNq
l/UrlD65oEGW5/K6fG7riSmtRWBHJJSBP8S2DIJ8/gdOIpHCowQtQV6LuXFZP7XJKGEDICVEFkEc
N5UusFKUKHqP5ym1XAjluqfIJJwO8xhRidGP+stJN6pLul+8UPLqj04DS6Fvlxm9cNdaiCBNHNLc
CKJu5t3tevbWmtUFDRMNbywAjxv0HNv/+jCCkXlzNSe97TJL/tf4SJOd4EKyP088LS9Mp1OATy7Q
hGlU8jYXsxgnXfdQ7eO+W0RRUoQiDBXvoKN4rl7b703SMBaAfD6ARqlf93QX5CdG5LQir6u+fD5S
3aX8RFrWzK3T6Ljo0vveJYxdkOqt9vB7N1r/HEhdlIp880Kw3+I7GrD2jnKVkjlNN6lVr39W9auB
ePgfL3zCq/lbow/MAi9pdFOe2dnDmEYS1bji8i3UJt2stJ1xXTjVR4QzHh0YDSbz26CR+yDGfLOb
mRTH6NBftR1Ki6M0/ZO1SSLBHbCQ25H60PWQtxIrw62EqPMTbeZc+6aPzUQh3mH0umh+M1rPnS61
pNuyuswXlAkK9iciImyvrag7rQybaZ5W5BGmCOe4623c+j/Zf14EBEgiitSnKHZCY9lFBVgG3byv
P3toNncHFhNY3AVPXAz3GL+40Ejefn/DYUVatM8ZA7T7bQjSSRmuE6FgtJyVedvVPl2SXUzR8Dt4
P0GD13N/W+dSHICscJ5uCrT8cHVoFk2UB+b9PLDcxRDZzHjhk2F00KZF/3NM+XmftHBvZs+k859I
fr5ZQEi6iVuIeZf3eX9pBMm6rShSbdjxu08YJMaAEjf6fKLdL6zye2936Gg3VAB4uRQGD6zWsQ0p
nwFktdzrFk1O5Z4uW079jIFmjvYFUYkx4HUaGUXItIs2h3AKqo8fLE4+rhpoA1ghQ3f3QA63R2xp
7GfOHL5UtFeS70Np+WsltFdsVlYcHGx0qR7Pp6XiOOCHW5c9K3LKHMWnXsaEIdSdSdanZ8hpyWZy
U8P4mM4x4rvmFgoU2yk7xaSDNjddB66qS9vTpR0FgFVyScCoFdOgxkRIWZpn8ucGG95nTDifv2Lz
Ef0gNB6aRXXIjJgADH+2sYV5P6O0u1U3FEQGa7pSYMmeu7V9kMPPFbTuen9x5emF5cLugjfpCqwd
4UwlyUe4YxwB3vkSP4M+0Iqj6f2URIBGXzTxp2MqTsWEetaNnTtf4FKHHQQMcRNhAKBoOa/1O/P9
N0sFRZIraZBsAxbTayseZUAWv1egc7pp+QJ2+Ypfq6sZv/6dfxHk1GKH3XXIj6iCiJtUkX/Cfmte
tKkCi3wj8Lp99sg7qrjBLtOJSLgVkRgSny5uhNHlFLaczbBBxAopTa4o3QOJSKeZN25+ZIe5Zr8X
RAGP0JcL+htiiz2jsBO9ObzbZO613sJlejYo9DRpIoj+xwwcHQ7g5GfchTEeIVjNpF3MC+ce9m82
NxyL0D/y7tSqNFYxx6QXXFfnSQSUIYmCSydMDhSM5m81a49S5WIwyWv13mS9D8BmlO/F/v1qTL7A
/4jMFx2+i4j8+QxQzuiFmpzv16xxFNzIWe5fuFR+kscg514qLSGxtFBKyuBoKgSG7ZyT1TDchxks
CEyzUb/xDJuzcCIsgoR9IowoTvfDiXFQz+IrXXPZo/zzV7PXnC8lXN3+nj/UFc5gApo4IDWwB9eC
mXGzfQ/aoZKKmST391nuM7DMkVC6BYmNQE0DEq/MDyY5t/AH/E+JLNQ/8op6RkKnqhlocLkPKQ1a
B+mD292FS7pgVFMPkhBODR93sFoctGgKlP3Uy8FNmfLD/rqMxTJQ9F7E1MV6pGKFQ7zivu9zyDh7
Mreu13YX/avZDLbk5hNo0xZb2G7SfadJvYdRr5UupqqmMeR1t86YEYp9+4DkVilBl/3SD4kIu7ya
O71fHjHxdNp+AGwdM8ZrDpizaCYa63vKD9HAdqom/Lh415zFDeWG5VVy7tXxBn9R5TsBn618Nz1r
mvkD64tNtS7OYpQeTSsLHBxVSVvdw4j+P8oSiCMzrdrfiH6+btmm52CqUzVh/wr6R8ytmEnPCsoe
hrY7njvt2k++ZbEbZqnj1DAY2vU8QrUWyJfy1Uy4XQsRpdk222Z7rSRnpRYlGGXSAZFWE558yw3+
x5Rpjne8hK7s0s4+J1QnJgXnJzwgrwEVdvW60ETs0OGcZr8YAYrnGRVlJ2QSRSq3OcKmZHSCZD7G
XyuncqsSoLwc5/8RW0FoW8/NUmBp6SIRfPm+3koPetA9lsTtGThqa4SEUHMJWv85Wc+par5fiDf1
JFhFhDGNV2l0f5PfiuDjI5sFuEHb3/l+qM8upKMs+vk9opaIoXuJpJzKDzq/tEKgAiPW9pjzimm8
nxY8hzNJGM9XBP0zl3HGJn6n/pDjKYJ4Jfe/9p7Y+heHw3AkkjmXJShYmi3YOekfCPydedPWEe+Z
0/Qds+E8sClP4dVmN44IYnF8JvUUrA3ieDQ280cN2X8gu+hG9YjBzPTHDdZS/c1V+5xUB/vrAH86
KzeRVH/yhpwS1SWRl+6f3nUdjk9bTYq5Zqinp7pDq+wePCQdTgdxAP56er5IbpB7TgCc5ptv0S7l
bppekrICAiKMRGBXM4mcxTbPESbAqARb9z0q0MPx6W/S0eokNjPOTSCR9iFD1plYlfsuyDI9YvEC
2sNAVRSMBgs9vveiJjx+5Ma0hDv/XVyyMNP6TSt1+Fq6Zy5FnCUlBb8FYOr4tEtJ11Imfvo5Thi8
RukobDI9IYQx2ZUFDqf0MvYS5GLymCue+BlfOLpAne1zQKqZ52tEfTG3MtJDjW3mchfICPdFedCE
fBp4+v4b4Z0ilLGCczKmFiJrLyvCMuj6vMPiuVY03mzu3OcbKefG2jpwPl+Ed5/YDIfPFnZqTaIY
Pjt34p4n+NwZpDF8POZRwmC7EkIh2uHzTUtpDWmzKU8OHR6OBtQ57oxGSAbFGRbbmgA0hCEPrdk2
ZcvrhDT/VuQ95x5EWhwn78CgnqwDaTJe2h2q2apsveZ/4QO8YUxmvdsNGKOov+VPosjvX9Ehwt+0
6kF9Ykr9XKk1BqsLlragnh2ILkkMuUwMDpV+HIJ734bN8lJ058TbjN/3Yc4bjoDR9Rr1cr5ZskP2
HPbJzx5P+zQpzWCzGuiu5Y/VoOLOmZE75GnRiZFWPQjLWCsXYoqBR/cwsrSksbscSd7VesH6JvvB
HdT4zZ6Z0NitWJde7CeJlR3a4lHGlVD61kwpObmXwutV0hbaFcR5+NPuhkoKXvPx9nuKTpIBidqN
k3gPazexr86Oe+IuYacKMiXZahopHoCy5mgdUKhfY30oEnVbaczFKOBsucKypyi6SEdJP2JuQrDa
PqKl6rSJVDanchlQHIOlgWE1krkCemAAKh744FemFWtA3tlMnqN28C1RLGSxaXiI0pMr463X0PMe
va2qXzNkQWtIRppi/Tz6wC8QK/dI09rTEak6yvcTqd/vdynkmiSVsTWHYXRYIO8nSuAPd+Wqsh+w
Qi7p5itkzKELYWRZQ8jSPF6LN4/Jy23nNS1bOwoaAhTHik6XAhiq4VgpLG2ij/oR1EylN1yHHla7
wB7Y/d/SXOtwdaaWiyTrQyequH3NkZI4e6AJA3465a32L1TZSrX64hYbpdRfnOETWX7dRETu822/
GH/Sx7w6G+CA51hl33J44yFOTlQVLDH3ND8MAcmhtaQmgUQpisLUcNnHwkRoJa1p64sB/FiPWUYk
j4yjq/m75Vd+GHoT3EUB/m2igqepNxUekPD7EkRJtOWP2FA3Lhh84hkJCbk2lAmKtK5GXkvz9S74
Xrs1KewymAN0ejnxfUjC7oruc8g1Qd9XkewG0bC387Va8scktZ1qhGov9Un94AXeNGkOaRyNtFtz
h93MDm3/MNDTG1F+vTc+EOy2MQKW8lxyCb4feRULp4z+gUqrLK6Y+kpX29o1wEY7Bxl4x0W7//j0
D48d+eMoD2zpYrK4zemZViZymfdhirH9E53v532soBNw42PQq21JBnyTWS8VEymkc1eeV0WKqbg6
e1Gb1I43SRTFX5fkX/ZSdYeLnf7rlaWQMmUoqclL61sq5MRTVBGFZITRBy4ka7qY34rRqZG2C7lP
5kkdokn4t3NPzi3lzrPkqXfOGGX27gc/Ecxu6Wgj1AVkZjHOi74nZ6bKDctcwqO3Jeykm/mSeORR
3SXrtghLbVTLrB3YrmVJ1EN85uLoKy3BsXSyTaWNiRZEY5IPg+RIyGrKJGOHwJ1+INI3/Ef7uye3
i7k+WteJTuelzrhjv/KxuKSzTsn40CCeSghLR9SkchileKAmqj08s8oudq0jCG1Pwz+ZqipTR+AZ
JUAZDJOvzubxR5oqidSVNMXrUCj4Iyk2KaKwmz/5/dLIWgv5Muhexm01g5qNrixeBOYOX4QLXuIi
SpeN9CBEznWTjdSVOJIJqDwJZIsbNMG1EpPTaRKJUYjBC6OBAyx1/a0rV7/1goOVk/H/jkB825zV
sKCefRmnxN9cPp1iHRi7d8HRtnW24LcDZrM4WqmB6PFl0GtO8YnrEtXtb+pm+MvZ+YTVbZzYhkYy
tdUsKoU/+fhVLdSjmjYiI5kbegxtY8n10zJMMU4QQvv/SwErlZyM4cTqX7bMWOvKZJRCR842nZsC
c+YibHCusnzeBTvgJfolLN6q4b4m410eYIDtijJ9YvqBmL2X+9uZyYt4hyrJbvsSt6/8x/z/2g/Q
CM7qdiIThcNw3qegB/UlYDJRoClPQ2oz7fdF7q9+CxTk2Z7Tkps4UOfGP2w+SQGyD0RCxNBJsQBI
7f6Bh95J3pdyrkoHCWTme6V5jObTSciXAymhTGPOfsNhjjgiHD9KTNFok4CNQxFu5dp+LDHALqWb
/B4tTqs+b01GdgBytSAUfez4gqkEj/sgnF22ClR+ixiGwVrXeBA3Pk+M9gSfG9xRoGWLLVJKvgB7
4Y0z9NuMsxbXixeq4E+swU8RbzUhcQTGTF0hjTr4Uw/weBFZlITyZlovsl9PpSVoleINqxQP+aHp
CsSiM4FDTK8PC5JPyM2paP71vYN6NzBVjK/tDPdNjeBC4I/NoMzYxQ2TAOWowBoe5db6yww0gOU2
Ppv26buz2h8wxQnd/Lz2CVKxMAldBdBRyW86A7vrCsLzfnAJbe0mgWRZeMIv6Q7kndY7y2LtpQwO
mD9lpokpW1sReDeZMNwxnXdCdYu2jyuNqPsulu1DpSShvdA/rZXvsO1+gSzZbe4BNupIjQgcJohr
GhA/BmOaoLtUvvnyvR3ZvrCSRg+Y9U1EoJdR5tBoN6OG8bYTMRK7EHaGZQ6hdw1Ph4LEbf8EQ+Vu
35kxZ/zFp2/7KQuFpuxeKSWU2e1F7aCFCBW1+ZFDZCO1EN0pNIbiSmr8IrEqkQ75c6X0TUMgFUcS
avBf8B4Nw2jjK9uupgVKwm+3NUVdXfric7t0EnuWRlONn2SOMKJvPmeGLA1kCBo6tiIn958L8Hz+
um+oKKqlLOToCi7MpLXs6deU5DVxJLS0XWGO+JNKIiEX/pm/q49j3XABnVlqWE1Aq0ZbmV0qu8jD
Vs7ZWPmb9ThNd3yxf9tp3CD7JPdwv1KurEVKbLV2x/pDjRT+qCecUoda/CuiZy3Ux0/SmPY8ev60
yZpNZEObaa4Pq/MemTdXSLSOk0VphUZtAQwYbftsCE1YE95clJ8LVXM7m2AQ6QaThetXgUW74TMm
bbhf8UPN+YI/qm1wmH5oGsSZX/jmmtIm9+iDmlO9x8zd0G9W/cUW7K+ZEnJGbBUT9Sli50Hv+n5E
FW24iZ3j+7+YX4f24cI17kd7m71yDsJsCdYVj8vB9ewYF8aEVmC48TK2bLEJ4/IS2iTQdghxEHLe
De/0ACbz9Ob0qA1fVFK0DfrzjLN8HCuJStYPQN33QJzpWsxMSNTvLT/FnPYIxISV9qmPbXzu7ddN
46pr6hg5ajpvlECNHR+N3Oe8WarYW+zr4ucS60h0x8eG7iFXPrbdi5AH8K9eVgQGtCFxuMIt18AM
MLkNpkoq8CyuMKaYJo+DMfhRFs/zFtx/YRPXJ1gfr3+T4FdTqAVwr7BjNF2hZ90srOTgZqBG/XOo
PXUZZTk9g1PHpJ1TSnFMU9/Y3AmpEUhl0IF4mfqLvQ5PSp6G4F8e8d1clYbOdLh9qP/NN9WlvHyw
ZlJZfEV66QDUDlIBovhgxf7tk1EWhnrHlZmjDNPall/nQJM7M0a0QeYQ5P/aTMhp1OYtH41VCHLr
4p5eTfxOi4/+SVH1HhrZv6a5Ftnef6syUliqvrI7FI4jSZgTi2MS6dYxL1T6A1sA0aOaS9c1ALf7
SB1PL6kJu7H5jl+MtG7Tq7lP9rP2g1B8kDOr26D8H2j0GnlJJ5z6dqPrZ2rN51uDu7icFerJKfpU
7LNpEGM5EdV0ZREFUY++dkSum/XkATIo3KbavRyMR1ykBgkhKQ+p+VTHNpIKShWj5mjKB4AaLKoI
DHjIB05QFCvWd5pMLVyT42KfNrvwHvgEJCa9AZKmrOt1bvHWCIaTtRFDf4CfqGWwB3MGY3uFt4Jl
mFRWPRler9I13eSMrxms50rssxFcoFONUQ061+CJE87g4tMI2r7XoHZnxBAE55fZz3FcZ2m0QlUc
ile8YKUAYFlbX1e9BcNVRoNyKY+IUF4Ub4NLhVhhp0lYPrlX7h/SEFu4I7jEHrbYSPup+RG9ZNag
Mb0lUFtqHj0BaXR3aFDl93C9LYnmiMrzF9X1ZGent06jr8f/SDdfERzazXvVEJ53zlkJlZF7QuEs
ubNDShFvWMCqGnSHsu+f0O8TcEqfxy5Cpmkq7SkoZPvOkZwLWepw85n86llfaWW0k/pn2ZOKXtfv
pYepGL5j5NsTdQe/Lb5IQWTfQJAl7eISfNu8SkfY+uHUrTac8cNuiGijN0lDsHg3VS6VCLX49A5h
c8hAYWix/V1TjgaWUUPeedOcr1dC5//rZL95MiXUAs95v48GRaEFuSS7B6aiFW7TW9aqTByb8YMR
DbEytNMzWX3cTO/bTBo9YfPgWVV0LTWUDYatBP87Hfxlv6dMxGBHnbeWsZgzEOYXBnXTb/LejenJ
JWz10LuNHWl4C7oOx02clZ0uXOm9e270u0fGT2aQomNsST6e7wmmkuLUSxQCEUkrL1NrShsGIL/d
iRI1+SE2WMTbW1qvstAMuQxkMBeTiWMsk1c/2dEfVW5Ce8KJFwMcHsxSMofyPWdV/LA/0n3kXs/w
Cv0TbdTmQOaNPdhg5ddCNpLSahaNhFBJnwWy9jhQbezccOG28048jjhCmktYfXk2NqiOu1aRq6qL
qQSTihGifPrW94LM6kc5+2g5BHiXW2fVNXrQpcd7HBdD5VWXkE2C1JkP/BygARMsr5jmCBqjzPak
kvqP5FedhCse+nPzK6YMUf89RiUO+j1Zuo7WHI/Mkv9SauFPIxIvaVV5eCeIwgNrnzBMeI5Ephu9
wMbSTtbQam97bqLcOnqQF8cmMBdd7oTumFvLHBDAoPyGWWUXZiYJtKb/vRDqPA9j0ZaWkVNm7hRg
y9xUAh1w3gJMXkrD6g+xFzgifkp0riF890lTn9/veEZ9MoB3lfmZL6kZJqUDpdjV+DJTo0MvZJV3
vsQ+RSIY5dtzP/4quSpSBRpkC5w+djPye+xAnWg2IpJH0Xt+KClLGHkVgsffX9viXXwfQUEO8f/k
FtqFNfilc/PRnaqbjtfz5lAlZGQgBNBqgIj7w+uOXp5Zvd/tUcMnhK3dtj/KfQkgHT+h6UeFMdGo
BRo4JtSDEZsdzCHLGSeP8IlCtJ3BaYqiHpu+Zkl7M4dnRmgXf+fVGeIZUExukskBc9vyTe+779/w
3V/RsMvHPdbczV4/YNpPaErqvXJOP4B/7PAzxVaYa2SrQDjKaZZmVrwbNtk8kGxQWxtasIQ11KyF
Ub7Bg60+aDsVRzNUyW42/eh3kGOChpZHomQWVv9lCMH1vGyaF/zLUjSciPyrHKF/I3M2pEF5N7sE
L2vIC5VsPvu5z2wFEoOJA4y+NbN0BIoKtzjOdILrNfXDppT/5HrWfVLqUg6FkgewSlj2D1twb4B1
D8gOynZezC/pUqQ2BcUowRVwseF2kRLtMhmEPK4ptTX9oH8TsSFYbD+8LXW9grA1BVsX1IlM4k6N
Nb10PmgjjO8d3AkQEeVNiG9kqQsBcq1JvwnKcXOPOvmk2nWZ+rQD5EaM01xjLF6+DxdDyHgNeVpI
Bgwbiguf8w9tKJmuT4PoPYlwpOuR0TYDX6oiVah9auWRSO6eTQyvfS+RbEU8LPCBkPNG1aMG60gJ
9O38kLzVDErxYYtEVqbXJQijFWK2QI081d/0GmuoGH5qu6tCr0y3+DWfiSl+IyPxCfK0ysY84LhB
mc0EAbKBbg6oe/vwNJYjYO8TtVf6gU4hU2vAScspuqSQ9y0r4NCeqX1xWTkw4yStAqVaWa6AcHCM
t8FPt2Dy3P90HrUDI390lgbdqZYS9kEwADw3rk0KxIfanKcJr+XFiAxtke2MPeR44C1xKF3JGcVV
EEmfv+vVzvsiOgurZO6ob8kP+hk1uPSD+KgzxkIpNQRnlQ9dMZnRZM3fX/GHUWt3GDqFxNtmungm
T1MkhGhFV6Rfcky2U28798SPGhwABfKI4n768mG2Qaj8U1TFkanxMCBhS28KYQ1Lv9GnFUF3OMkP
9b288ar9CRxwrAMqqAgV2iMLufb7CBxuAMzGGEfAbKD/yWvN5UleE4KBg1rH09n2qnHT8fVmi1z6
staAcdH6E1jhZ8Kn4E5OQHevcnUgPFJjENeeMnTxFBDea18KNNYbRV8wkBnllTKJPWqkPFeJiJNj
LFNWS4dfNWOCrOYampJWqkl+1OJL+YhkKsVAhBlkIolgbct4KxKmgJquyI6Gk4RL2sg9foFTDZH3
z9o918aqI7I04a/R8K0hJuxFJ4Ifc2ZdC5lFEdI2fmRDWCOHq+v+GUiLOOPGKP+bToHP1ADOrMbg
wPqDZRBipvFPpdba+LCo7qMcVXTLyLfRTNH/rD+yZeAk6Iua0whhf/Nk4t/mKXy7fLR8U9YTCAf9
KjmKq4j0ieFUlh9G4zwr5po7NhuddXoQ/0cOf+ntlxHS1XNLuJdvLYL2lh4JH932mkUXqE0QMOrs
y0aXfPPASTugut0Xo8D+3umD9iCZqA8SF44fMdhOlvmOcgqKCFLaF9BoXGHSMss7tO/m1MrEJKnt
rNzcM4rD4NaQmjN4kUbgPx1GOzfvI8sY0ZpEX67AXPHi+CA6uWTy7aIEV4T8eomvtPgq5VMZYTJ1
x7He+PewGcmWDWjTfcJYRPrWlvSrU5XQNt4XU+wKr8xROQ4VAw8JGe7W4a1OqNZQsf8y2Ua3occh
lMHi6apC+LD/NH1nL82C4IIDnyqWyS9JLhtRlAdYgHxDUlXu8+SxGeGtbEuw/nPco7MlhH6nQXyX
tgU2LiIl7jwlL6oZVbKEbMHXs7J02aE+ptm9K4UNXbxHx8P1goZCgTbSoAM73B9/n3Px2F4jtG2V
+Q84xhjYlN0+ffVPwUcv4eCc+lB2HtynEGmDJ99sa4lwx1WemJljHHwpG1K4HNFQksApkTH+VPOP
A6Q5KJIBYFbNdqHUfdUQfuYRyiobKcEMCjW5BNmfMFk70om8ZgsDOoaeswPwSBrA7C0dpz9ANIQf
YrBdqt5C2+8vHTZb2qrBRYiA/3CjEOLTkjS5HGIpqd0l/MGSJSTQA/NSjxI3hWLyWrB9thFGSiBL
WMgxOm/YCy7P6n6cq/RoviHvW082mqY+6T9NnzaYsuRDUnuj5eqXyaq3jCJG16VMcCDxAWKZx5Og
q8dDhkFJcooxKkh3Yjlr/6PTODUYxC86wfD+WpCm6NGmhT8QFFWgHtg1gRJwsGKDtaab+bzPNva4
ThEa5c9VhFeYf5O8+qA9tNOBVrLnYEWTqv4m8MfjhP5Xs6ugt0O00wdNoX3GuJHIilllZIF9Ffqt
HuUOPGjQ2mu3ELey8JBwlptKtf5SCXxO0k2gG5LApRhhgMwfkBK76wj2/jVG5VPHBBNqH5/SuUzn
e8FzJU7h20bnNN0UozzrfSObxfuaNiJiBnNrMKLe2BfuZfkv1g/QD895ql8AkWHc4sVgUkq7r7rP
jesqVwtnWJKuFHwpOYS0cxAZAVcBonfpzswM6rk1+WmO2viqL2HnBvKDc4UUZLRr1lYOLn0DHhEF
XyaGPSN3KA6zBMooox74zzrnbJK2zj4KPEp3CHAknYYiWbmuUa0ydVO97uZGzP05r8dv/1nsawgB
zpjNLvuKulu8aOukIYGzYx64Ikh7nADIwN9xqUL5eN6me6zSJCRNza+NWt9AT+9Biijth6uxbbqr
iP15Dn8gFTnR/1gZna4KWousdklVa715Bk+v5sEAZRKAtqCx0B6Ka+VdWY8b9TufOfXX/BPLWgmt
aZRPn11uW3RkjQCGJE9am/+FoSnX+YVtN/5A1S8e2ZZ3lH3rkyCwU3sMczxGZosNgXALQKY8WFkY
9hghaUf7Fn0Mff4yyJd4iGatSpmSrrzsDCm5igKThxW2tpBU/3nb9KEFAIoOUQoWmgFNNKysvMz6
h/8mx4uAFZKgXlALRF3aI7tJIA5KMSS+oUnaBP3R0DnuF5oTNjv1QT0kTW3zfmDoI8q0eRKx0SWT
piIKIHsFtt0uEGoDiW8SQRr/u8ucII7JYi4yYqyccy2ZczhzgzKpg9HBJwTo5mSmAeqM6pTL7Dwo
ac2oXCBF/ZDJDW0x6xBwYEkRhh1B/cs/PYnO0BOOhdWgr3zzRDyruQ2m4e+p7JuBLIxpx91JZiYT
eAHg0Dp6CQiBJbyx7ugzVSVB1TrZUUO1ssBSHEdNhUZ10RpWr+lwLlBnuHD23fTHq+Hyv5ttTvOZ
rEkv4n507i+bDNKyE2Nsja4H3W1qGALYOK9dQiCiUHCaPYhT5z5S87QiA6S2RJq3zK6A6/fxUgaI
X+tVVjT+2q1depJCF40+qTooUfD+RRjFN8/bjAzuVH0Ud9OV/rlDxd6DydX4pgzAb5jGvUJ0vwG7
IjWISULOWscBFdfkkS+TTZjhhtx4AxLr8t4jtxHskPLbbcz58CyUFrAdd/HnpSx0H6cAa9/Wg8b/
yApfd0VonaO8N/7m1bIGhD7TJA7xee2yrIJuMLkpgHEgeO3+uzQoTh+nB8WqmIzfEnaIsoQtp9Pe
uQUDbbhQXfM92AqUmmINmfrYxdZ4IwFHkjwjJssptI3teX9je7dV7Z8OXYtf1tkTJ6rTwz6Ri3LQ
4MoBUaKtblehA3k4VmvnTIMpwxi/DGfngVFt49TsH+elWQ0nkeI4xH2j8eHTZYp09oQykjcDZ6Pl
ei88WSPEosRvtutK2zQpPqywOnPfcvK7dxZ5W6P9guCoY3xqRUQ29QO31VKtLGq3/9l0pbaj+JB+
lVrUXi20PzdC4NqimV7Ktvk9aQv8E8IshNhqdtuguJ8bhF71fX5KD363+555eG3Wyf9fntYRt6b7
emE9BDUlxigz6YlC6YZH8kccjSNLT6FOSBW00PJu875OaHsGYkj7MkReft9sBtOHBTFddLpeC+I1
Y0Ag5u1vaYnOPstOo5RdwGQ5kvzGLC4sTM0SC0eVr7Exg9ZKTZuu0LqXIwf6QAZQxtnluuR6NK/B
rGvbkEtDow5CbNuV/aQ1qB6aNdwubcwVHg0vxSPBAtWGU9JnQAu0TPpTNlgWQ5vyaxX5K/TWHwRS
C0/YqMpgY4rVIMrZo//6pKb808H2lSJH30VixPVL4U7w+qo+tZJb8OM/oKVkpnEFDr9+evFEPiRT
EDPS96VoN4tiMdwvZiPCcSK03t4abQakCZx0B8qM8PHw9K3pnq5QNPXNEVrd/SOLRIKWfKdhswu4
FWdRQjsD4em3HTZbfwX1mVbtlZhO8o84wNuEvXWqd9Lavg/Xai4c26CuUXdLFn6O6lFZRmX+bx08
zq8n4UXJvbozTh3YIYu4XIFe3hpsqAe8dIo7lk0gLgisfVfxetqkN77RQ3OAxoUtGMLg4YwalQUv
HFEfdquFqDhU5bVuN1p3oAt+wgeus86SfjWHeQuIjxi13Pi82kTATMxNMZT4RF7cX6icT15/90d2
AwwjOGrymfixzZhsnXd2xn3aS4W+lsdGxlAXqN0qOOgW9DU3SVBuRBAU5QTJkTmNWpHY8HlRrV9X
hXlmowfpoLpqg/CNeXUKXQcVLGzLtveDFbTmu3Ea7GMc0ko0jfSkv3v0SxCK5mZEdiXqFB2tgAlj
Er2a8HuJ3o72M8KjV95RlqCLW+hQWmglC9cUVKwWSyprKzFyzBCgdFUDoGeJkruyzfENHco2SVsh
oZh90WVsiqJ+cOPp14GpFbil9LyAGbmMMxMl4zptLQL/jg1/ASVKgXHSVvUsoi9a2EFmAnSk2Uvd
QBT7v8UVf1dtmuEbhUgFdQuNaKiCtWOylBiHcweTvDcpPTzjlTtvm74lkawicEy+4gvE4hs5XXgV
oTvC1apRlGkTHRtldbeENCCfqhF2+5L5JHh4AO6JIMinzEhsNqt/nNZbfT9nFZg5xm+/sY2m1Ary
klvTBDETNa7Pbbuj8Z2Np0JB/aWiFjVjg3y6QLBkcnDZ4e46C7zhSdczfpGqgM8UndI=
`protect end_protected
