-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
xqbgKu2SlkDU7Fz7iF+F6B9PXT98f3yxPZOKgbcnBMu+Ezb4OXLLd5E9VMIE2wqQHYzMzZeR/i3Z
1VHhlTToRq85z30rJ9TpyTJGXIds7KByXR3bzchXEAR4cfTPoHu1ocv9G4mRwaO6WPjZdqaQUHNB
fp1F38l1tad0PLFIZnEnzgeERw/QEfNQTO+umvfyxnMyOnLCrLAoQDU6v7mI6JJYBxL2yioBJtPF
+P/PutqN2HUvPKIU0VVX955fBu0LGuZi8deeJnrHnWNpxSs3QJicu6Zx87y1XcMHi/G8Tktt+ieK
qH1YJjqHJgTt/EH6/76g+W85aK5rVSxiK+/N5Q==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 119056)
`protect data_block
/RPAtlKTCW++fD6ydaADjcNQ65JSLcYdtKjcPblGv0uZf8WohwUhMT/5hHpVdB7H/umU/e3jo8Uo
z8NtsCEpsVkng9e9QpTOo6Ol7L4omgD4esHa1pKKqAxoQZiqLynMxtOF5ijsbF63PSWYilyRKpND
hjf4k+7SsqMS/BKpsSOBfMhS+TPeTngG8lSivk0ob/oeumqA1LkX2SZl6nO8SBQ2KWO1uElfrWta
MTmKVqiMisgdbWYYXKb4FGtVeX5evQJQVeyrYoVdBo1q/XJab3f4dp+BrbUpnrWh0d8I4dH36Xo4
L/mV9qUC5X+lhaR+NFKdYW7WJQNdO2p8wax/uo0BsvFV9Yfh3xuHyuwI4uzRUZastCxXlt6TRxLZ
4b9PvlcKsE7Bl3U9o24LL31U7R7CtCuWvfa00UnVjdCXCSq2mCMK0hct1iMOCvZlMi+aRA4kS832
CZ1fSKTZQJWyDa3JrXbBqCiJVlV71KMCkV7T0PLxgJKV2Q15F868+oQ6vdZDeg0A/1Fx7SgupYLe
jiRnrnyhi8qGDoSpvu5rFm9SbPpVQ2QoJhK4E4/KvM5e2e3yW1Vs93VNawlIKPg3P0wxP8W+Zgi0
Bd01hL2nPczguGULw1SlP3J70vIO2l1EoX3wecmqXBDwak5uaxasaAXdDHPF/7bJ6f9TgnWCtg50
hHxcjVX0Kj49xOM+55XZxl4CjB5zjzmpVrNkzznMj6hMFEfm4WgAMxv0eG4o9Yz1VCWOEEIUw/Go
ak8eNE1JwLrVQomS4mjnxj7Vv15Yxo5w4Q3ODaJ0zLzaQdlM/UI7vtz6zAHx1P9Jutdaj55h7BqU
47necDKVPkF2YhZXDkwfOYb9XxcUg0A8wYn22HyouY3BXv6ZQsWGQKD5/CaSEBkodJiG8n720T+m
6POk3gMHfGpU+OPW1axnQZTSrWkTcsU3wXzefl4LM64EhtqsnPLl3w73tAqofYzCQXlZ97fGOhSd
VHPtCIguYi/S66yNDF4Nm1izXZItI3BDH00ZgRG5fZXHIEfadAwLMwiHAyXIsu24h/7jatxA8zww
hpbZzBE/rnk9O3Q6urCecwXTEHnyR/nDBMuFA/CjYoiybj/Vwe02hDu25sdsTqvXDbAvAI4tcgbv
b2UUhGSPOPJMDEZnOqihj+7GuauWVeOeuvNdEJRS6i6uw+L7mbDyaANdxmaLqyeLIfj5dwdxG+a2
6fPyXDfDAgn6zwQhcfpydigR+mdxhU75XCUWEI9b+w1LNoMGZbBxg5baoXGl8t/x14TRK8TK6MX8
1VPgQzM/IgDARYWiLzQEN0/UU60C88MZdFZHXa9d+XXIXYZZ5eE9fC63iy6wf4BKjCbnAiPl3cn4
T3y34XkKQvEf990gcTTA6xppbKesKdaTCkD+gCGwPT4QF5pc93yochui/keu4HMQW/IQhNNH5Le+
lmS4W2uRC8JSCgG5k6LDj4qH7b8okPVLlL/HdlCFE48g3gaTytWmkWIZ1mVImfnwFNfAuMG2SBAg
Ujs95cMdtJu5TXLeyq+V/+P961fdWc5644QNc/bnQVgLcEoM7/G6c4xOTPXUw6kMCKWqOaD/tE7A
YbDdUiDcPklwTG4eG0I+4GzkQW1wkvh9y5fAmJUuSI8P8xGc4/o32eCfEXLIak069qCbEZOrUmbq
cUPPyvhY9UB0sakhuXga12W/TpqIbZd5R4AgzuFJDhFHw5vG4SkGW1/KIy0TNPORDApiy68Dve8A
YTwq/G1mt8Pxve24Dl1CcznOjR1zYAmTfRCqmd6WGBSUAlk8mXsTW3RRhs6as6Fl4csf33ZUcL92
XBzDQn34259SImrOs3uupVhYxNRMaq2f4woEBipByhE/fkELRuYOzCz+nfjfd5F/bkWrCIkdFpw9
VSZIndDhuLy/Ng1uFZKXkGBpwL4Uunqub6QGplzD+TcuHKXhwrBmpkcLMZJXSk42OoKKTyvb4Scb
8HkKq8e0CS2Bh5Kmd5C7d6yr6z7tuVArZo2sZGHLGd1uPvryUHNlF9xPIkssaMlAcCPuxJlRKIP/
MqgywQ+xqs8NmNkjj53iqad4InEYdwrLfqDDvdjb1yTBcaI/gSc/sSuxjVwcZ3qhSVOkFMDre0Pk
KnkS0UNA2yDmjnuBubq2bs2murK2TzraVjYvnosgA8Eg4Nkdp4u4d6e7cJZKi8ksbSEvSh/tYMwA
elGwfBodRLqTHvNh7TUZ99WEOeB142nuj+jbBR6jiKRTygObWDuF+O7w2LkljWL+BLmDZPWbGzkI
K47QjEpxsc74gqlTBMVJi8HJQCQK2S9bZBjq78hIcvfKAQ5P60OSJGB7rCqnk9FZAV4X9iEZ07iE
ZYCm7nRv3UytM2yF3I1OMlHT3DJRD4XhHRlJIAcJul1GXaZg0g4qjMCJhYtGVRqpdskMvxPOHONQ
SBTuA4/EApoh8neW4308en/MgX20pVaOakZ5NGZG/ccQKv2pRLhT+Jw1OhseDVJIIQulYwiBqs3w
LJMKMH4hmW79ugqE/9Rc4YbYxD7Kpyga+4Ni7pt/W72OtAZuA2+OWPJthr4xP15HjlXGYkMnVWMz
J/0t4MDpXb9/2EjBsLl+sva+R8cTsDopdpfeTE2x56GDEs+VAdawQsccwMIvotpTuzMrrNbMKyJC
xhziAGOmbglvftHqrRSHP+XslCVXGMp1f9wBF9BUspsV76W1864odBLeTOfb2P9vbX/YimMk+70p
dsLpPTIkK5v35aMZApp/7FIttKSCIT//LlMN2bbaX9NjhU/hBZsRTLyG3ZrItuqWi2ETI6zZ0N2z
wcOptjJnDh2bQiOrN0nH29khebiFECwgrgrdvo45awuEppStHtv0qIMsGC/tolv4QA9N0IoTGkDR
XjOeodJAIkbtG7iOGrHMdwCuL8ybxg7VNVtMiY/hMC8gE8oFSwEnRemD6/9fIR8USqRkHt9m5Sey
5BiL8aJfgd6IbYfYXODjwrSWNx14BeHSAUbLHKZmbpm3sFG4HZfm2dIzJFKb228GQsB/f92OXmeO
wEoaC1BvRfnIIjNomzmzq1J42TZzolNTekDHSGsoQF7r2A75TRQek2pixWtQX839a9w7zluF82Sa
xz4AbHvuvWD0ur76qmr/UtqGOwNuz52SK0JVSDb2OX0wDw1sDptR1aT3ZdzF8i9xC2iTC2RIaP0s
grPXY/6JEkZL+HK1SCyIus0a7/puCBjDeKh4H6AGfLugvjS1aslvf5UiNHgVQIT1tKDt37z5P1+E
zw4NN2chKhsn5Y2RlsbictYmTySTdM297vLE8yDBLjk/WwpDa/pNlh101gFtT9kevGWg8yeCAP68
7SzctcBrkBXjq4cVq0o1mfroTTSlWYbcTE3Rr9yV5pSCJ6AYO8O/UTKj/scIl3XwN+PMNHTEeYIP
ZkKCqW8gUPjofY44YTaA2zo3omPFV019yV1hffE3KssptPHobeQTc1I3UFu6lHA4cLwiKRGMwZi7
OvMET/H140jDr9u9L8B0tSylMNU4uVpDUMUCgk3oQDqWAbfgmYbZ7Zt8tEAtEW00evKU8ZfT0S7A
o0cCS/aQmUDQA+7hvlNaaEnXN/X0XU56zqBsELcZgf5MNxJdT6NSBFN21Sa+jkQl4r0CaEAxRCFE
yon/Wp7mZLCF9Fqaq/i+X1xR21oRXWOIUPz9L2w3wjDFOjaPG0sZ2rrZCr3C4Gk3cHFte/3XSxvr
Pq+L+eqL2Ejwn2ElG0zdH528scH+24gr5/Itaz/aqSNCouf6yHDHemUNMF80ZP72SvW292dDsoNZ
cGkFY606jI1KZmCePQuvKlmvkXP9VjfCJpZmDIkPIgpEY/DNRBuuG676FpUMXaftDB11X2IH7O+L
CI3bSw/269efVJzSWblPuckbwdBxz5p480iAVexAxPTc5NfS4mLWV9uQc48V9ikaLQMZYL6UKHSp
xs0gN1YY5TTdz+EZsd0uBLg41N0sufBRPrkdKrNhpH9IxAFH66fQjPb5QhagEegGuiaWjAPjtbyC
Ol40f9EexWM3hivFTyCMwTtlnEd0Ypgs+1m20tFLJ1H8SD4cikMQK6mRoy9/5wOolQsUniwwP/E4
ZCNFO+q9kEvQiHTbAMwL+xWDZe9+1CRy3xUss2tON+kDBhoedZKmw5i4drx1RFNtC9AnmXqPGEoU
1/CAHYp5inNyo1cTZF6cdS9lBdGPRkjBXP/Elz3Lac0rSF2SVZlnDjk5+u5fXzW3lGjYnxwLJs9G
VqLljopqbO7hmz0eiEZh5/b4vFflcjdI0StXPglOFJ7sbN4vpxcjzb/Ih+8xbiCSFERXEMgAjxDs
56P7A3DlVTNbzZiDpOd97NuTsU8NrXeDP4pSiRgMY8ScUxtb/jNKfGsrKrPUcu5S7xEvNo4O2HBt
4CHJcw7o3Yxlzsab6PrkDOuefmOADLup7jXgeTxmZeNAZpI686SraBpanQgVp8rIwl3MKeL9X6PL
MnYxdCBVWHrbkMWGntuNTI9TRfUqR8m1MhgwYW1kBJHelUx/mXASBA2mo69T+aEfT2P75vdgJxQJ
NcbuWFdt9NIDJ4AZ8scs4M7MoMqnyt3p881pr06LKpK2amjxrYtzWe3zG+7CJXcjLzsDxT+mRKjr
SariZenmswGgHEHVwEAlqGaKUHnTqIbIQtWNH7NEpuliDiXJSHuy9hXSt2FfSHgZrJHtrx6+eBGD
clhZKovW2S8YpDUf49xXMOCRqUjr1/iE3u1YIFai0/+tcVMX1sO9UC9o4aOkBS+ZKdWbGczmnLfT
H8UrR5dYf/HkNrwtep5gS+W+tcIpEbh0JEiHuJlBT/u1c8UUcFqZ0Q4B1ZDi155rBqpZOopQTdPo
1HrrIrFPFlU2jitb7OF9QpTR2ntMZpd4QHz5hMRCQinyQ+Z7k3yjSKZ7YR059JU2KFMVWpbcGJF2
8LkQR6Dh8CIV5hSrEJoIEhKIlZZjM5gOPq42h9K/RXPt/vb2MjAECH9iIhxOP6XWtrGzdhkjZf36
Pkr/zUvXRF6CikeQPRQb+Uaqt+GAcZbVu8x32ONK3V4FRj0DS0nK/NE0O2dUeATR9OqjKK/pjP1W
Sk2pLdC2d5U3GMiy/UgeDSFAB4bcnk65HIn8PPD9gaYCKwH8ObyarL2/7dLlfgCDrV6d5LbouyCd
oFA/YKszXTxNqtv2WmmWIJMt+587a4eTVNXznhTyHJ1koFESRT0e04fS8PLTFHGILl598h0TeTc1
Lo/p6e4JPHsJX5Xuq1W04Tmbma5v5uItkr28J0CmOrjQAwaFaWr0kWjTnkI7NsIaPs3gWFGnun9W
HV6uUPxCyp+z5CQT2f3ueETATgl6OJ3dj2eCi3h+Y23RtPw1QEq9A8marMT1njsgFOSThoev8pL8
HVU87/rGjJeIoEJ7wu85R/ITk643ph2CzgQ1dJNUp6PDcfQrzUEHmHwlDhhAgeSPRl/2IbMikqgd
id/4KAzuESASf5OXgtpj35yT4UCA7NhUX7Y4sPKVLefWkq0tu1ruRDelWAZiuYw5B5p1i0PpRsD/
oa1fdem1Le600NyC+08kzrDN2QOCsYktKE0ka62uHGlkPinWft+XynIzuqVKOH9Vig6TI59I1F+y
jCeszBgffhhvG+BSPYben3gyqsZp1dgJjbhaytiFaFUGOOV9c2r/eoFnLjlUcI4v2W26v2N5q/cL
zoD5oecBYyu0G4RJAjOfk46gX3NfAB4kNeoR66FjUYfw+UvwtQPMaDCAE9bU1q0ieBAeT7JT/6dd
JExDX6qjowduv2/QGSRbKDTye0OIfzNxWvrfzgOfzRBVw7sWAd6jaq2uD9hsmsa1evhRRc+f8xry
6s5sRhaYQP5m1Mloo81h7zXAU9fI+kwlma83X+T0zScADE87PUZJ2BRoyMrQCtSVzQU/6lY/tvUx
GczlnqsQmgQXx3hzv8xA4ZNtqQF6s+ZCD/V4E2/p0PBdPGs0m4UUY1sF/BCQgtPy1lnNXE78Ik/4
Ss3V81RxigXM3pmytjJwAir5TfSjuHNrp9RBGV2IfR2sfFrzrCpUulx8FtkjwF5ZHBM2uXUsQquX
R55fWgnAq61kSYo+9eS2KEE9yCrMeBs0WKvP1Cgjo1TLxPEu44AoFr5ur9WXKLEFrCbr3aGA0tyC
q6U+BbrjoqjIHHkawYXM/+9j75G4dTsZ6X7U0H7OsLdUbFKF4fW3zQ7lA7kq0W3kXdtmKlimYHbN
03c6Yfr8j5qeBZAjDkTNX3iSnC46MLdxvv/UzRWec0g0eHXQn8TxbbgKmIQ5Gu7swsUM3j9t/3ql
S/SEs2PA7YmZmih/pKP7wzy01WNo1x0DemIP4L79IMKLur/YS/XctFU9MdGEBpgt3vdqIyza07JJ
v5LiLcbA/UTDrUmhwlqbw+0pksZsywr+/HRujqigjEnXmXhlRaVahYzV9Nj1130qcCAJCZCmTjhM
WuNoZq7yJOlTU3EO/u553k6ZAspgNScGXPGmZw5Ky8fX3B/ZIkp2QujfmZK1r1ocBj5WA0+V1uI8
4qMFJluIU64s9MeFUsl6A7FSyzoCc+ap12qF9Jq5txOOm956KrrREOQvj28rueUw+Y9v4SkNO59d
VVuRv1EaJ07Vdeo0xnpUKCNES3KZCytXSUBLQggHX8JPOxoiRYik2G3HYqOq7kBIxX+fdyeRULaG
cATszqDKowDv9SdV3Fri4cKJM/BAvMU6/Swh+nBEdu1QxdLiUragP+fuYBrRNrSIK07i0HRx43nL
6zaf8hb9+4kZxxLbnDRX2m+oKN4GJ5S/u7kqRGFX30ssL7wvug41s7DQv3tmonGe/NU3Mzjc2DAI
AVzvRqkMEJAx1UzabKFadghkypaQ0DZ17C7TsvQHI6Y2/SpwwXA3CdkGieQGyL/NtoYwhxr2XhHz
Arzr7R/XtEhdsTu9lPWuz9IcDOAkAkI9y1SihT2d8lqwApbnwKkAlnOh9mp6rqLGbg/qOqCGxm4k
HqE6R26sl9acCF8JMLrqRtncxDPEzD0hbtWEs/2ggmfVFvetnoPQV4GXsJDXfZPcu7T+YIG95ZJm
Pn2MtXdZxTwbBOL6MIjzTVtKojrAAbBVugzpaE0ywRLr4WcyItaPUFCxGBme/QJvcu+stdLLi6v8
k2da/QgC9xq6pBs24U9EPtwgoBdzTjuLGCwOaJjV6/D8nHaZMKkmE7PPZCG+uqaBUDviRZTKtuDa
lGbZ2Sx+Htv4xZ3JE0pBtaFPCwDpB7+1CnN59EgxdqZ5BpZTOrhoEWoYCacygomaaGyNqhwngkaB
+zpEBi8NtsoFntLznwf60/eu0IZWB2o2NkBwUrIczKLxO+0SoP7IUmqOHgy/yv9/WZbLPRpbiIOd
rMLZ1fkmkHd9IpKAviqh5yfSCfMCmptm+DzIktbnUOSZn1mzhjORX4Dyf2gap/RkFEK5dTVRaSqf
w3LCFKfFEatixcLMhm/5N2jj5tYh+IcpjrTBO4gDosvlJK1SnW3/2SjZ8rHEx51F4/xtsBi9ae4b
fMzj7STL/UZai4cpR8OWXjwUqa26JWEVGGmKl5g1mIeRzNKFPdRT9L+xw5PRXZuXxtTyi/Drx6gu
pVP4/SBuwzVX7YzVmdGYjSi/Cj3MSmMu54CVtvFHA+L5CjhQxfq+HmXTTxauQEwelDHm/FEK+YY+
En7HYAE+qZWdOLA/87lg7yIEMTj3aX93hSXL0/TZAJIPfPFSFnjgERGNeYbxdhsmB+bv54hLsdoi
Gs2hXRSmoj2YhSeWGgid32tlChuhhpJEmj82/Jop6IpRMbD68SwpZBLX+K5GNIQuOW1HfJfOxB9g
epoLeDUYldSWWJeqXT/u0blVKSgqyCSKBXtNuInzrH4B51ObU8bARCXqJdwV9IzinPjr2ashx/GD
O+YZRBX/qH1IdIjUqJRPqBUNTsQeXt1CwOzSri1zpHSwpfSxfxJqZNq1uRM/Zk7ros+Y8JZQr2+F
qGqBYTj0JuMJ2jc1TcbqXIwOTnBtxlaDmfGpwTkSl0oxzvXx44JEgOtmpUX3MoN4734ArYJLDt7T
N9sM44av3ZmCC3Ufud7QPVMYr/ODZrTDoRuM54ttsl2c+c20+jimtt2YDKac7IHxSKyJiK634abb
6DijNbnLlK3dxW6EglofuDzRz3Pp5NcpAOGU+roULjwp0Qne+kTlUUvAi4jzB64seixkF5Wx0/3A
WHbv8T7Ci33EgXXEHa8N8mqYYaAiPInUSn6WELVMX3e4aKTmiXjbd3i8vQUnlVWMqcDBCJJTPMym
I47h2hmM+G9FlfWF2qOT42kwJhgIgaomdO07W7ztBCKNcycWA933dXlbbXKWM8hgjHpkQA6ET8ad
TD1ZwC2eiR7W7taO8uihksx3AFx1Opl8UJoAKsgpI7KjWmQNu5xJ/emgEEjYaeltOYph5ADsWj0e
FCXpx5rMbGoHNeS4b73Q6bGjJG4acWtFIx9aYa3b6laRIW2ItWueSQWI/oPnndQ+Ra9lwLgAlPXn
EcC1cNRTHqWAbKGmWuqy7Z3CemAOtmDzzrZKrnTpPy9K2VpilbN+/+tpbc2S3rQv5yJy9JgcFnac
uPFPuvO6hCcmOh+W0RxKVpYifrkuhPbdl7Nxl7ypsRbQsggk/LzjG3IK0PTRg+AqDOI4cnpptZeI
79g9ooMqnyNyzBXkFnJSASOYi8b5FB8bHuHywhXboAWuXuQ/tbdCLEMdhZDtPPZCQxS2Sz41Pbkz
ZoL2TVOQXZYO7y9H/6Md6XfTVO3l2lyrkxhZfONa8AmyBbBiTcYbTeBjfnOHsgR6tsy5s7R2Bayv
ks2SfmTC0VceUhaxOvt3oavpxHGlE+E0Ec5nmiv328P79AT4F3O5jqrc0XzEAmfc9DcJ80a1netC
21JmUv8aiTgIOnlnEQpT2cMccNloV+37IV8yvwWMMTK0FHmWxxbGzDGzXKBSckr2YoSNST4si+cc
2ZbM8XOe3V6GSB8idWZ34PoTt2W6XoIPRn7MXXUr4NI8CpRVNlTA7eMwwasnqL9iFI4rFwQuvbP7
b680vGcI2VZ3Ld6qaWO8dORAWgkzmpFP9N3vZONJOs/5lIQ438IQ46lqe86mC8BP0YmShKNDTPiw
BJXp1kn5IsHg6RIX3tmZdQW9nhZiX8gn877SqdATOV+yfmB65lxAnXVAhXl5lB2TlvLXo18Rq0LM
wWhHTJygW8iACnUZet8UpQDjW7mLv1gPz9+02/w5VR9UpC0DFhjUPNyYVBXJjZ32V9wqjUS5Z9+1
0pIIRjJ0TxASrPOlxG/LUXF1L7HjmSf0Ue0zQXbxllMX3aGzY/QBFgsuKytPdnBa42lpnNaDTyBN
DKjn9nbaUUfsT6KctnVkvlGGvlEh0LMjAViUV1rB4QWqs/Xd75ds+E5EOFP6cp0UKIau6JIafRO8
hQcPtnxMneUsKTM0gCpCcOoxHJdqssDI58a1EbtKan4v0k9650YwFxthatzyVkwHQIrXBp9YnwFP
EWjcgKV3+/Ocrw8qclL8TXQHdkTVYNhEzY17hTJEo6toykHVimQ1wKnwyUKjb0bsW8nxT/8Zl9As
vBaWG6HD/dim2GD0d4wJjCTh00Hx13ICFzsG8zAY6zWokHHaOZvItlxyh1y1Irg0lDk2jc9MZS+1
4xyFFUaO/rQ8Gbsb3L7on1Oj9xDiHHDou6kHt5MKZzzU3jsVvCaOUAZE7aoYlTHirmKT2iBXDs04
IMExgmW8ECGbay1OPqqJ2XHu8kf9Z7XQJaq61bYoYR3fTz2XY0zpAMxrhbn3MnEQWMkuErmBGaex
0jtBEEAKkVOc0IhcHFfvr/QCPNCF0m1LnV1Mt5S0IbvEg0YXfSgiFyKGGgY7u7StQaGPde5bwMQM
A9nhtxCJ2Upn4K0Vs/jRdPsrdXL85sM4m/QfqAcS6If4iqbS8kAVQdSHIQItiIDWplTtqHoKGpaF
Rv3SwDxsrII96gdDpHejaJkEcksTNlmMvZcWTgokP1EeJBSVuSLZhykxmWhvsj5ZVKP7032U7JIx
H/Wcz/oK8HBrZRA2SWt7kTBGvyp6kSmxILVpkenDXfqIrgCAnzPFIvnUh2cfqeDKvSMIhM5DOTcg
Crg4d2Sgk7ZgtcVIXJahC6ZsKZI7VpHfQq0nnIPgN3enex4ghP3nlRUv8BFLp2A2ceom/1u9P129
iBfNuFjYWRwvPBjsq1V93DTOUPFRW22qnVQLdC+WJ/D9pyAeiQefOggwAYIw+755b9KB81Daou5C
BHDz5+FIyzRzhYfrjDgPGWntZO6s6SLWSpQ3GF7WBKiMHecKNOx1nP1nehRExFwSt2r/tsPzSWog
75k5JgkOjKu0s+yJpKfSxGM3Y2WVmK/jp8UohCzk0Vvrwat59QQTGOzuqPC3MLQT/aUMlK+TrNfD
VgTVGzR8KNS+NnNxnqrHD8cvqft14ZiHlra3cmerBlaO3tZF/lgdavqIgp7FgKtkeEB0vWTyHjtP
NGhEVXQCaj+AN/aujcM1IKYSXm/RbMgdSez160LuBRSVofU1HjsI4jmCSWsose3EG/JiiMv+gxT7
ogU+sPP4/7PHXQI/vxZJ0lsEaEE1Eimj7/NXlQffOarDvixRKzGgkkzH853gIBCfjVx/QmYyvnzt
CuaYHCVhvXF+iG1hpJ3oZDOhVxk+aWf8hO5RjEZ6Fbs40io1KLf3EmswDzwtXos+//6i9O6+l7k6
ZVysdnhzTNIL9BaP4OUhnV2oE8KwTi10xBoUcsz7pWF0MqtLd/Kj0jGYNXEOFzswJywZuy3pcg+h
WswPbtrfmYK76l44Huqdyt2RLbB092iqwcfMQiM8isP1ZYIyGtNP8XvFKYd1Tlp0BGZ7wnw4YDT/
O3+o162vIi+3VlEQ67mdXzl+7TJlJoaHLDNzpDsyuKwT06gkCUkO6dSQ2qHZV3ObwvMx1IN8Lx+R
LA5nZgEiekYQS+eAw5rFFfiRr8SQ+3Hw9ZQ3Nw22dxD+rmgT03Jo6/8WXSU9L4+0pEf8DPKwMmF1
5ChSiPA3TpDhQ3YPDtKxenO3QCJw6xcNcLmI8EukbDiCdN3GV+PDdijT1lbVOzAPZ7WjU0hUCt/+
K3aLIDU8lmGhsRbl5JcNHo+a1d8npekfcpRc6Tdtn6iFHcd7jJDvYrT1v4T6oJfi2cGVij1kE+k0
ikLjp6lRmDxx/TlTSOXrY0GLJuhTsfS5YenzAUVr2SN3hAgF4VNQOW89HZabqi3wG4xOcNxEl8Fb
/BbkLHeePiy18Y46jVyOAKrCIwrLB4GmWHe7uHUnlcz4f8P9SHP6RYIHStfA9XUqgreA0zSzX8Mh
VzPKMFoRpxyEU176ou022JAd+Q+tvWsuIOrLOjFJtWD8grA9S+SdbnVemaoBXUD3XCXvuxTTdw/X
tnbPvSOFJL1Hcus8srqgOap76iehq4pKJ8rCNDn6XeFVIueMU5lViLMpjt46RT1NzQvPQbG3Jr7E
2LKRsv9DcPx+cqhbiYUtrDGelbq8XD/iaWZ2UMrFpwAxrn4FjusNFNyCB6v1oUDCCWeLSsYj9vXk
aZRuTAOk4g6dvpHOv0NorKDgD8nWO5v62gtxjMbrKmq0q+hvu05uS0qerYUpHYPSs49SJuXht5RP
b51TtgzgXT4PSHVU5yFR66zpeV+fqCHSH9Bte6gyln2FL7AjN+Y/fgjlHhkTMPS5NAil76QZUN6c
m2zqSWZnbFDpmRcbe0WV8/c3hDnk6sqP8dSOg+cdALZh2sg0TO4gJDyt3/azEHYilYept4/4sb7f
8qjmZgBW5t+uywRNvLWRgSkyv2/is/KjMbEOMM5FyQtqHQQzv99WWIq5K4qGHojn7TbDt+aUZ0Ki
amsnXCerzQb0SGzpoI0sjTVstQPdzJ5DRxURsT9vH+Poryk+LweQA5onznsp+NsokrLlGXvysxq4
RD38aJaPqQ/GGDMjY7+DRbg98oRdbT78nd83WtF9TqEqRaWRgTwCBL9i0ZU87WvzByvtycj/ibWk
MuvwxkqcrNX47c8aEk9hONYayXP4tAYl0+OX3dsgrD289YVgkYbUVkpcEwnu8LpId5Crw5i3nUu1
HwciTXCTTO3azuUcdgN96MRyhcdcUyjkf70lVHhcSO2KNOqGZVf0HeXoyLABc/vSzFspUUWGVAFH
/ltSmjh9sYi05zedlTdtP57vzGKIgwoxTuPpWW3wOSUdEGd/n3cPoNqaBMHZ5caNcR6/28cY2EjA
K+u8f+lzEa1T8qeFD7Zm1G5mY0RHTjS4KGqIymaT/Y0qPcXcoxFSzVKjBzvwLRy7ZUEEC93Z7JKu
/4xYUtervySeQEvPuCfHN2ZDXWd1MBRFUJyn1IW5mi/+m0tLKuuFGrH6okVp+3IFR3b9xLGf2JQg
s9Y6v47vN5QfIElHbTp1Tk+WFdO6JXsl2/IWjgYxKEbk9BQd3wE1P75xqKLr4sI1Kraq/5zlrsO0
vF9Z4Uq5JuIXEiruJaKE8GJgs8DM2WKUuPgLhXHc7aRUh96NtX1UChPFs8Ek9wKPJY3t3TlXK63h
pRolOGgbeHS0lHetllrofzIy+zuTt1g6/E87ijEybReD4GE0HnuqeFGFrcEE/S/Z9zXLqFw8XcBh
xyxEqmdfE28epPqx+CBVR9IH/abvOwVlb88mU6P9bixDrqr4tMRNIsTQQOMtQzBv8mdjVFOmke2s
WWQsA5mpK+stSchkbvm/wICDlm5PDobFhDP26XWkChuiV89Cqp42z+e6mMZtaPVR6RsviRptUC/+
5wG9h6slMa4DWpx075Tt8gKHKQ81QG6uidG0BLTCC3ETBBy2mkD1KqEYGQMTEdi+Zxm0cT63Ttbo
N2NUDxnC7F7YbF/AxdkGMu+J5YacuNaXyW1yXmUI0lyvhORCs5BWIbQOgL2WRPHBAO06OmDuY8hm
fq0jQMbIqLkRsEsTwgw4L5etoY7GhJwqoJfhrOfpKSIrTEX0njFm7CZmn5T4YFuPsD66JduwT2yl
1q0UXlQ68x3rCi2phT/TM1C498lj5liTy9Cbev+S9diF/HqvxzugJ+XM880RCQyizgPQBQaigy2c
3ECUUimMRuOsbIIu+B1kbAMyGNZCSQ/etcS/IuClpPgDeeQfuSbt7COhkP1JLOwm8ppHgH2R7tQI
snLocL7afQgFvpLyUX3u0q26F3kCTT6rYBrnxjlNetCEnEBRzImhIiT1SD+lkbuC4m0fQ9qUj2Rd
MaA4T8GeE9y4Gt14QDzWn0+kE6JIg2CDzhkck75hY2DbauLpg6a3Nk2T+iPb8DsYmAupAeY0Y+4o
WdF2UnvVS/nrEuFXZC7VgJQYKog1FyvkiaccwYNzREmteEGFBVgpAW+IFXZRuFvhn0YKxO4pF/Di
tkuBlLDjpinthMXhQ2JP3MOx6BtQ0rXxCyvhmozcl2C0lU6ifD6LaeVOjW6aiARzuuvi/3QP44Ff
11Gc/7SMsEhrN2g8C3KnJ4asfTsdeReNSzVdi7017wNJYT/AUhMqynuUfO/cNiE1avnd4/RXIFnc
AwQuQlfOLOp2JYvk/49MgQLHovpbIqjzoJWfYkDWqaxqPhtKAWuFlF/aiTmx+Qv0cFnvLu0JGTyW
YqXlKP8xOoFZx0honBpDLNfEPbg3p6JXl5JAb+xKgNy/Z+hzu269Ynf/2mUAuqiC/lYRuSlv7HRL
tCI0FfyGuA8AIUg1KK6TSmm63tTd/TYjxTnWFN8ZBQGMLinxYLiW+L7TybpxegG5cO59f/WXWxp2
8+W7mnn95atdGNRWVr2cK6e7Qxd3sX0nZ7Nsxy8Hj6tABjOTQJcsFsP3r6pvfskj9VTVC6jzEEOs
gz+zoT5SaMaD3MREYNMGe0U6o0guBhbAc+3nENAezHSVqe/YRwdqXueOdNoapUnmo2ydHRHA268q
3E+U3poHWFCt+8NUchkjrOQgq0WsN6YFa4M4n4krL1xX1hLZZ1gGyAS4eSwGRBkkoBa687/G7eXw
s260kHLdWs6SVEy3FavWKHtJDZGfGCWE6HJ9xZ1TXTCDqC5l8AuP5xA9377tHVF2dZXQsGDJDjjI
07TPlev+ZMujNVnqNgc5o5jk/rYiVkBNozAdSBAQWxF5u1fxVxo0NutXZr8g42sts+p7saIEmLmR
xe5hYhO/ctMfUmPVd/NhAFGNW3xKhFcZcYrT4OoU+DtaCWqADIWd897N1MwBeFAEIVaqPmYibAiT
1X6Tb542X1b1bWOOsJdRaJSLlfP0UlHJbT0Om7cjaGPDuEzCgL4h1bKz6G8Dq0aALegZe4GcQlsO
drMp++juzfyjkF/7it0GxFoeEokmPyKIc/B3lrW0g6tg8DS0HMZrgn4tYq12RggICJDmLREusD1b
/NfTMiayUn0powWNTR1oEqVg6p3Hl7Nc+X71MvxqWS58X4OmLuFTZZ5K6wKnh8gFV89smtGLvCH0
2alNYO1bvJO7Qq2iLUHa4O9Fg5RbrYooGnZ3H7LcyJ6IeRgmUQvJDr6guNK3ZT/KROObLZ4uxt0V
MPXlyE+Q3Z2m1Q78mFJPVgOPHEztpEfPu+oFAE1egr6z7iicmVINRBhjkM8oX10gctanaIPPASJ1
AP5gV3VN3OU1RYRdQOYAE7v91QdJWLI1sfmuOqSX1WWYyyYydQmgTLRsQ1qGbMn3QRLsHbXzaBtX
CL/53Inn1HaojoBX6VzB0tmlO3NR4e0cu5mR7bTcNINppPcsHmw/BdtCEaxogWj/JG/UsGuyGnYL
9sHN1d7WT+D+MMCtupHYXzG4uNKQZTPTgTq4zEN6PfXYTQ39p+klizkawH0naTORVMsEberjAiEM
ZSN6NiSGkBdI5GhUv/ZqeCGCFN/SL9h4WME4uE2IAlzyl8kGSH0UDmcn3jaGNp88kSKXSSQLY72w
nXPoKNLkqTD8F3J96a4fEUv5l7rf1Zs/XGtXwMwReP8SBLv2sNjMYwDR4oIzXhZ/eyyknj36MATT
JGkQSg3wvLj4q2DAYtdtkWYx9s6YAxE6GyyCiOjecaQyYbCOHv4LFzlzsdc+tl06aHrraDMD+F2j
N2Zvcw6xPT3BBS3tu4JuX3HADh4hTI8nFJBgk3pAZPpL4xLvIWahSCkiORvOoOihbrf+h6xBkZ0/
oRxp7p40BexXsSmy47trNddJ1o0nHQzs5iu2u1dTWxAjbfOYDM6mATqXRXJXIZluKZAEJMfOT2YN
V0clZxd86izgwV/DHa+h6wTtIqgcaJJRy4tlpwCHDxN8nwGG28XivZxwH1i2hOMX3qGTVWX+zRyi
z5OyZXm/cv03GtQQYY1aOgeiCxhzaoDeLoTLmQXYJTb88QFrk6UMIkEFIvLVpLRZEutNMtiE1y2+
+z1493eo127sav2zyoeY3xl4cYjEthJHfHKZ5Czb9dV2cfKN33gqWUay1YFzKVv11LazY66yJywQ
ECFBBBIh1gh3F9n63nUV4P+EIqSEC3yO2TMiOTkv4P3A4kN20HiKMy9XtOxxtlvlFBPaO8v0m8pj
xz+ZlJ54jpoISP6Ox0kt0iZHKBa/rcL4iCGaaK7zd9qBD1T4VtqJyjOCnVMMJm3qodhA7O29yESm
uh5ABNF92maU+2VjtdgHvtAD/MSvCyg0Ldxf68w+hsJ5LzA8QgjOLC9D3ZRf1tK14/fwmyK6DhAU
/1ve2TtjZyv6n+4c+QwCfwUr0n0V7L1tZy6jUYSyky/NKEYXZ0LXxdvsh3kUlrbMXTLidDfqq0Uw
WqnbeTORuCm8Yifg6j3j4GzeUrTEzCRjipWmRqYpxeFezjNMqXKrVGA9I3o5/Q8OQ/PTAhXvwT2T
pNrh2o2tskvOmvYAsZu1QtHHNfQYuU7yRWpEmIZ9E0jSBqnAAX+qHNxeGJO+r54LXWVk8Q+xFloM
mRZ2W8swCdcV48amaftgpCMco5ri+LShd8oAX2Cp5im4EcevwMb7qSwKzSsid2ivBnTnJk6/1vri
IpM9nCb1YH0zggMjdfGhMLwqj2suo9qJYJnIIFlhwzTtlv4rzq6ZmdszjIs7iPFIl6cAUQNYCUxE
yGM0CeGCdYPHTYTRhpJGLFoL/YOCCAsKfHC3pDrv5K/60/Fr9QAn7SIeG31ZOkTv6htB3AQTtg6B
wZy9L2caKiJCyOC0TKPRg5JTXZBxGOVpnt6/MAyigVVDQIh5JumxukMFiz0PRlbMiiL0/3+KYv+q
G3cdk4cdwaPaHLx0FqRWPqNZ/qxrpwFhfovntHTAIFE4dzbqVzAB8U8nU0T3De8gxiCu1ONr4Djx
AsewlOCZrI+xd5ea+hLqRKRMXuRdyJhWFc+25Q1QGYO2g6FdqYCES9FOY4YAH1QfeDbUusVqL/l+
BgGz6XrEu6foIwwDL0CUqhEb1BOBVubs1YwGR8UFG5tmzbyZN6QCsKQukTHQiEYSjfNciU6nzi1I
qoBm0uv41qzZ8E08BJamn0pUKJsz0U1PB7K/lm82Sq+pyQTGactBmB8VBWbW37ICLFdkVVdaNe7a
ADuSi/zfDvF8pIbr/XK/faSLLoNgjgwblJtuKu7qdDMUaor7I6DT7QIZjdBnC9LIcdEeLwbt9bna
ACB6S2snnNoQ/NOhmBlPlfAxIIongnEddVkFgFz/UmBtFexnbZy68/b+xWMXaUF2eqSgabnbnHCV
+0CHRBtjDGKulC+jV5oxcHkCSrhlLsIB/PyKTGvqGfCv76B5av0u4m6UsHzgdpaL/770P2a3oH/C
OPXGV9aKrpWPTyfU8xzil4bdNEbHrMm+zUJc5wJ+eJiCEIEAAFHf3iQ+LSuq558l+leQ8tQrB1Zb
KfNgCHqhb8/iJ8hhUDhkTI9IOhgaZig0RRxUd7qc5DW8wIZbM1IheSDgW9IyEVau4pMJ2pmNdNI1
IoMe3X4aP1gCvDs5oe3o4njihz8zlZ1eAe4yM0j59bAsrtgk77hojDEYyhaKIjLqLwjJ+nckgYsm
NmScr27oXdFzpvYsxkJoI6S5yRs3ayc0QWJgtT/7RUOXZwi00gdv0pmgpUbaG9zjeoNAOFqgL1wL
H/Aeeal7Qd/4GD7gU8git2agBIwTKLzlrf/mazg1DUF60bSkJWlVecW9c89VXf3E2kFIKXG2lxAf
Lz5vYXOIRHq0UTWYH83fF4P0Sy/eaHjY7QNvz785IJpjgJ7vv94ipul3dRFbL+DGBBDMZaXSnIsE
Tqs6+Wh4L6p8vkumCeq8diNbLRnKO6q4zDVXJc+Nxkm2ryhPk3/pDNnWoTQe8e3eAUyV0sFLaGVW
HfhjSztwCy5E3fvAu2T/IbKb5zWKeSN0K6Tq9XnypUx3SwBb4Rhu03PxjTtPrTFFJaRxx8JKECPz
IswgMVm7dA3gVpXtMSxAYQC/OcqxkV7/OyxKi7R9eN3ogkJbC7Y0FGEViGB633cd5isWappqRTsb
Xs+Boxx7iWhzsRQc34xaEvyKK5+x18X8r0K6Vlru1hyJcHDIbpX6qxEcHwVdUnZhcZzc1ceQENmT
rQKX70G6HC0oXrBWkzpcUF5F958dTURtCBSlhDw6upk+dyAUhcqIOoUyUT77qR1BCSEhYRmG92Xy
PaINPChTTLp6KV1SIrhwSIEjaZE14crJ8f2x3JGMaTVPyBwhehex3iazLbBHBsaUkvwFz7dna3Mq
cppDCDfPjN/ss6Vx41frJqtFTtwRj9JrtT/jk4QycYieaPkZzq0gp8oMye1kApYeNiYUvWN5I5jW
Uh/VcqZYCQjrs8WjNJ7UIHuMrymQtQlOuP+WLk/4rHkwyoBMcvjY2OHjJxG3BUCrXOcYTwIBEu2E
7WmTjlLoZeDxdHgnDugL7smEQozzq/pV2Q6WnERWdy6kFOIKz+WjelZgKbaNKOfEHR0FsbqI5Xu8
dSC1pV3L80jOn3hd0BaGFqsxqV3z4BacOqqwaqT3jSE9w0gT/eVX6cqZuvPu3ZKdxwKZxzRe52NN
4mnIIYkiRsuhNPyFh1wrXhx703+VxGsQVumgXYpS3IwVytFPcYZt5vrmNvTTfuIM1L5VpywXSX0U
wT239IQHFhpcxBkeCV/32cZjzPWS7R3BaDkIoYxYFEqagv3AzpaS1ZkSwIW5KaXo02NyoivkTFSJ
6gR/9u4AoJ/MrqRmjoDlcX21UXG+P7BvvlB4hlJn7wSOIIf9hrm11idFhH+IQYdfDwtBAFFMzu6K
nw03l6OzjFCFr4mhGRhREPmGmHqa/sSEL3CjDd0w4jqJAvhKBLJOkSL0Z0pZidVRSB+Aej5lcD6Z
Xtl+MnfsIaBoyOq8X95xTdozL7gC+RcW91HxSGqMkeNuQ9ka7seayd1bpmpeJaUpUlENtTztqwzx
voA+TCSuZ7B6wgSpVOtAtJSj4rYaC935wqtIbH1LP/9QRPv67JETnfPWUBpTo9kinJESAPM7YLji
anUfJGiM90Vhaf5xLgcA7lbUzz24mx33PYG2aQ9Fv/sEUN7jOCmGv9qqJxHtpv/unfiVND49qX9C
d0+isx+p8NVcV3qTDveqCPUThnsuS9K/+95TgrAguWk38oj+RJw4SodnmyiRTyf1xtYFpv9tOYY6
E9JWx5COsYu4j1tRZDZ1X7wh4/DJerqam3NoezxpuFwAGMxuAubp3znMr3xKGJnH9nG5fTYJ1oPH
CKcmMaRBTWIfYahXo1BsbrSENXgOP61Zs6ZI+hBS5nhTZIiEeSctMi4mDTOz9bWJ5G21E+n4IIUS
cO7TqvRr7mTGD8SU7t8NAJ2t5ZA3fY+bPoF7OeGbd7QDpLrPj15Z+iZbIzCL9ey9D9ZOoBWw4y3f
yayl+gZnNSKUcRHSe0EIBEu+Erx4ILXEzqZzMopdLLdLMkpzcv4qQnO1Hw/kVY8r00WEpMV4YQs5
d6skuHcm+MyKn/QgOYBHAm5wls4ssMxvD21OwxBeQ1ifBnh59ntROU/ZL6Gsaq1CnY5+pLad6Cdl
inPJM/DoCEZFnoe3qOwG6H7b9XkLpq2H4ThPNeNnHcFxNfooXVSNQZ+HQHfEL3hhXPgUJcJiu6Hn
eAEOvuih2HgUbGDp8qNEeyM6KCO7iLuKm9vNUWYrLl5kMvweW6uyiOeAzKw0ppCt+OuZA5P4EuUM
76YWm8Nhp4UO8C+wvYIm409/Mf281NJU9is/ZVlmX6t77IkWWXxTiVH4uks7NjElfUFmS8YKtgkx
nMxhgQkFjRsiU8XKsNvYs6O3Nc7GBReqWl96cOxGr87in7UkO6SKFz6g8hsHkVBtHQcWmWdL9UaS
Y0TyZWOuGeOVSK5cV/iPYRbUHDa2x31YNHbKyauK8fIeHJeqSRfFZractZuJHF+mE9f9NoItjtTE
qZ4Yyh7rEOiKnMtLQhq4f53G3S10QiXgNYrvNUkU2Kuh5HJ5wafY7yW//ZqRUFih4txS6ZBoYX+9
UmwpUVBQSvxWWziuNqobqk8GwjnOR59pLSlas+3lmNKDVk+cJV1YhlVpY+2p+eAGrCJ+FPz4Erz9
CfTTAzSS4iqh/ONkpZnf18NBKCxRruW0bSSvKvY48A84MM1Fg/N6t97QeTePvsx4w1DIwa6PDGSI
vGZgqayhBdsrs71MNtqoFDJdFJiTlUuuNDfXiyZF7FjxPTE6m+rl9yOXooUXHf81/Td9/oOLPr/q
y6x6mWsBtCvkrpEJ5D6XXCDIY9I3Kov+FlJWOw0LSCh1+VCtNu7HOu4aojajl9IyMisX4lUTBrU/
nbzwOZoPEypAb4fAObEO37k+G+rosQQk0Kop8otRkZeaHECc4DKgyHbuC9hG2Y34NnSV2/hpvicK
qPIfwH3cxI3OTlD6VdYos3MIauDFcQlMSJI8PINkz+yIb5Cdlb1FvtWJbwbAgeIG8Asl5Nsii/om
ER9sWhrTIFMt5p9po9IdiZVvkOufIGVZDubflllXe0psR+a/hCTLbB92ryPeXkUnLfiO141KSmYV
fVSzEHzVIFT0ks8iZeFH/gwh7Lyr9o7hS/H9iWdxcp58TKtml20e1W5xaO7q5tSw54Xl2GqQlO89
P7RUyvX9DfVGo6ytAdLNMbL5hjwDilNPXEc9okQPMtADujuAEDupVeeK7hMI+wPkNM1qt1U2oy2K
iU2hZJ9WKHrPA9Maj34EPlYAbI60/3OzRQe/QWKFVH+Le5UchofKP9hWyUgkmMrhK7f3f6aFJtpF
9CV/TqIDKh+l5id5rNbZjEvpWD3ljHKx31yq8tYr+lfOIAlPYxjA1MQpDk288hv6FUQXvzw3Fna3
6JEqKDhscVy0xf9KA1KjUu3BY+FDfmVD+ofBosN0GCLFHRCg64mMu5m3krR4oWUIK3xwKm/7fpoX
p7PNo0EhxHvpH2ulqAk4sO2DZIbxSVjrRqDqaB9XBA6rAtb6vZZRgIEmmsp3UQVev016LPXNBtFl
dO3lmHwQQ2OKT7ufghF5brwYLG0ohejZKiuWmZZ3rhS7fdSpe+hcu4c/OBy+DG/slT5fdOs2G79K
o9MEATXF5jhwMSfDxLna+12QPvDefC8P1CFEfqrtKbC1Ca1KXc+kRX5CJWsF4lXS8UMpiD/HYS4h
i8YhMgiCj2Ve7jruy6t9Lh8/xADDQkscNNdvFP0Tn54dE+b5fDn8Dx0Lyb+gIDj+Iw4WCBKbplbN
DkVdIqHNB1z0ydy5iewVYyHJ0nITlu1CcggpAMKdTFUEV15te8v8amI+1IvUJp7YyZy/HZZkbuDg
Sr6Avw4beEYLJacxTlcHNPUSr13+75HpV/iEq+/a+y9JyCuVAGQAgieDgWD2z1OjRE3lQ0gggOP2
tC9JhFTHvyxGW0srPuuHhVjZLHa4ta/zUmujxbrl/GEJdg3Hw4qJcROCdODFxdL5Zaj6dXR/2Spj
Lghc/y78iA5vWk+kh6y4Zk8nUpIHEHLZdf5Fr3+XQORND19/co51EAn5k3Y3dSkx3Nq78z4d1RxG
VG2FaW8Go7I2znu/rdUhMjiEO9neqCMQlVUxeKRdOwfnyztWjsszLC+JJ2s2VO+0Bzm6xaCTQZxV
0aq4E5KHZg1f4DQFTWHKzgyp++TWkbXe50O6ph2qcv5Vw0BF/mVejQn71jT+GB1ER8EsLD/8PUpu
HHl6rvgbL+ZOZvgTdVs5wmtwMCxIfqEZJ4vW8AiemwjMLwraJa6m/YL5ZnwXD4jlrMNzOrt0iZim
y9xhRZnFYDXS0wuA3w4X1rgHwPpxl7iW6NDYBB9zpcLef80VFuq9PMhgPGIR6ZCX+AjVysU1QGql
bYRsfju0oao42EfP0nqmY9TF9ZY34F/bl3zKBLcTRdyRrncVIXxaAqta8iBbStPHBLFSVc+XDSLH
/bWoIK9Im425JhU2wrSJeIqT7hq0mRrRrq1TOynq9TouQAo3ATDrR3ww1Ic7RTxxTogrEwmE9r4S
XwVsMxxot+rTETIun2iQ8JAmBMDkUSyErPBNblHHTSwIr6QG6miT3LdLo21PI5FNaqtXCche9xgm
lJ8mF6ORfdeUfTxHp+kpNGFzvXKeWvuUwF1+qKl0C6BMT6BQE+EiU/OIiuDm12AGTZYHHB3kH0io
uNG41IyOZbHOx4tNhm6wiYQBWHTaBROdXD2wiPHwdwt8emo81rBov9zc4Qu9Fro0XNB7Yd7hs/96
sjXP2NH1tF9LnzdHaUpjsnDF976qRWDymnIQIWeQNQtSUo7tBAIx+GEgtJrhoIlfMWNLpwzrTsOY
MH6/2i80l9OySygZJeQzQ3t4CMMNVO+tB0BCPAY1r60dHjgNuYjGXQt39Dp3i0jRUXkE8rUdxqDO
q5+Toqp0fVVA1ImCcjsOsIOB71r1YsOHPjKJfqFV5m6xkvVEdTvUUGtq4nvQwOQfkqN3YKHNRPbQ
9FGFjGxzTWj0oPkv3uOobC2cQYg96u3n0kRwAqmLG8D9NCf5h08ly1pES/DoXGYNpJwUGbUohS3y
sc27+eSgM9TSM+IvCiOVvqFFxSJbV8hCuOrXxTHU+gmig4roV433gN3FuYIC870Z9wbp6RstvYM1
eVpAyVpN2QbeYT7yziBOL06ut/ZqdaXrlfy9IYdeORPsuOyEx3BHzm02580QQvkXp3p2w5oHMYDy
SBtASWHfEqyfAbWW+afzLP9RLe5yWSH5nPnCTKu2m8p0aVTGRmKB6kQ1xvO7MWi/xk48aCxOV+l7
lPPWEAiYKLXQ1wwtFa0OUNhkLrUgH6Zg1FDOLLnDT0aBi6cKx04FG9hriA8KyAs6puYFoJHn/ZvI
7GUDtVAnbDyCRw0vRZ5g1vYF6zSCM41RY4ixi7tMlOVkcYCUS3CrtwbLuvyxWAdeAdPFKmmRa0zP
SR3qm1qrb2idS57jyYEmu/cwDD0A8viUoZySlw15c3cs/QBVyhc8JlcM1r19KdMFt5Niu1xwTNN8
h6r33SmsRy40PXnLQyQtsU29FywaIPzS9UeXpqEag7A9j4P/CDwrGOws4vDRc9bbwvAr+Gh49tHR
quRlywWu4STCqE++sf+0ygflLwyZWMrEsgbQTZ0RdzMeu4V+pKA+qOEuWyLGhjhvvxTUWoTa8jcJ
DMxa1vG9ihRuQmjmJaT0V9Pu24vbi9kjoeZ1FFKY5pQQDVVJKYIIznUR0W341GbwgIM3NZrYCCzx
9GSWzfIorgGGPc2Qzdz2M+Zeaa2MVHGdiwdJrWy0bW5gpD1TZ5o3X2zouPitpKf09kMfjOLBopHW
Sg/HfJ3fUA9zVnyE08qY4rCFEk26DWs46/xgoPT+FqVqas77FYf3QndmwAuIBXcMbe8oZeKHCmeF
54JP9rx0FBHKxN4Yg4RXXEvhlIcq9Ib9FM+46J4JT4+ZN+L6wgZ0cwpLBrGGPBKnwXRwgR59jyLB
A4UKHVu/++z17rHUjKpXX1grUZyyUJMHKnOdu4j7kHPTtp8+Y8H7ovRv2xUmym+gPdQSw8FxUQts
m7yaU7+L0vZVZqi9qQazSSbiLUczAoUQBqzXy3RW7rEL8yqOFTYBRyaeBG9RV2KHh6pBo1YZHDoz
taawVRq6QmhPrDb19vI3Nfq18CYHgSmA4Hd01byIluhk4pYq4YfJEFZUWLdeGCM6p7GAhT9OMUey
t/U+wC6famm6NN6VWCcnCoN5mV+oTkj08GEgW9CYtuzXnFAG+YRj3qfHZ2Nsy38m6BbnwTJDQPt2
yxwAcUPl0og0tZkKR+ABbgwt1YDBqe2onX0n0w1s+ajPWjsH6OXIomR/Ofr+2+pC6hvFxvKsALhM
N1gtmYM2Mahwk3vhdbAn7jjJE53ZiAOqVUjZUye2Eg69Xt11E4OeU8ck5wSib67JWS+3XvxM6611
umYlNwtYEkksQh7WNKbvxlX6EkM2g2l61NcLwPy3TAtehhj6JcKrkVqaQFpYd2APN4MOR21Pu7Rj
BwGRvlQ+lI76YRfS9iHMhZTKKsBUY9in7VoKhkdeje0gXpd9WyoGGX551NQ9g4fYQqi+nJcqayKM
sGo4m8nRrQuFO5hwHecG1YGfnwll9WndDWKAdYOYd3UW85XvXPkam8tq3fRzL1e5mnROg3C3xJ04
QOBgxiamC3+GFLe8i+VFK/ziz96Ea6RN6DGwPWSk5zdidAzXZjsVN0I294HNW67vXk31JfzAaZsH
6amAG3KPnxScSl/YysFZHlWOM3DeNH4QQkiLSLlV8sn+aCBP5FF550U8BGoLFUFMxuXQ56jQdA1g
D7l4lziahQpUeHSzbs23dd+C0hrfxzGFpEGSqNPEQF09FlaR+0EEwn3p0RYd88icm9WA3iK8E6oQ
B/rbUowYGTdZuygKS6HZDvhLgvEyfQEZLyTGAONmUNo3oZ74o+FPpEqv7D5SbbXgrtvh6ObkYn8t
xcby/ILl64eXWjDtXeKA6Qt/9AWSo97l+c/lRv6cxjhjPKEMYA+XVFa20I2u17lYoEKDXLfVcQ1G
MRSSrLoJjucFWD5Zrr3B/Kxz4qEoYJwLVIKJ0oQsVPdGs2D4GZDwjGjt+b3Z3mbmq6OMa0/3E+zz
v8V/HHS4DmGlsF/hfXPMPsbGEN9s5fXre/nRm4lIRxKMiTtjsxjpyLePbZIE6odtbqZh0qZ6cgcy
2k3By+t5FwJlikvV7Hmjo3zcymiTzd6YNrT0onVxdp/Vm6BTiAB6Ly0XRW3qHKzcPwtlBeUaNITF
3uYdhro1MZEGL+bIx/Nniud6Gj9rtHlaGmeCg7gspR7kwXq/M9hfiiYmegIvib0pPm6zMs2wqh/x
cNmejOhAri6oBLdPWp2LoBm2YmqdC/Pl5966JURpEbdNGYTwHI+lk7WL0jIDLxUEG8MoSD6l+bGN
icOEU5sqEM+llY9zS7Sx4bsVrQqrac18GcwGG3piS9GV1nAP13mweP+WwzXeWzYDNnA22EJXNQ3P
ZnkAgJCoiybSxOgyOSgUGwMiViIZmQ4gQSZuugbg6C/v9ZxNJdnQKMSephMmUfgZVXOWK/qNmoiI
oDBZS9dtHFwtO0NGnvGgDqJTm0/4uwL+E1EssP5XCtTaynluRCLEHfJkGp4RJcP2ODOEl5/PfIKa
lrlmYx/1Xn1QnHhCLrntT0SGCNxA4kevx2BhY8kXx5RyGk5bCMI+mEeLcBssN6Nf0KwKpE3rBH7C
wjCuEl4pQrS2L/scBFpOjw/17uqNa0X9FIY6cUI3TlfgXfTVY8XSGfse4o0DMQG3HFtgeX2vXK45
F1DAdUcqj4xCZpaBL3ooOmgE6rkIuJ9jbtuAGVZArhryL1kRMlKZJLWQeWZt/5CmUWqvcdwLDeI9
tDkNMFuGzj/e8gzCjnwXWZW8aUdOhh7UNUAt8mH0AZfrpn31nA40NvKqyxkYm5kzISZgLWnSiFCQ
oWxQDKKxjjwFHLbqSf799iYmMiKTbofq6RcgIlGl/C142tX72pRncHHtL+veLgoHdkHp85ZrqsaP
eqk5nr4Yg8Sfl5g/s1KLXh0EDMmWojwdv/sCl9pKkdPEb1jFEFfVCLQvCpsMxmG9WaRSzMMLDi5j
uzknEL+/DKCWcwyVJasqAukps3j4QMDfLHilqO1L9K83xH2PWIpWdBQbpMgyPJKdTHawdiXogdQp
WKeGCp1bZ/RZAJqBHDZCORcU59nR865Pft40/SRs13G1+GPiDV4aoHMSlqKT3KneCpMyLtDIrjpS
YMoZUDfBV7ht9o/0tL574u+KGMrmAICHB0IJj1SjDOJFMftMIifUTStM/OpTblTDVhe8lKLqgMBj
aHw4zdEjVdP6e54sRiG+9kRx52hHzyaM5goEX6YcKY1STv/n+IpWwksoVrGmXeTyPflqq9/HuS1V
PYdaRWnp5QqkbORzTw8EWag2IO4fN+3WrVLE1keFcGZyuNiQI8JJ3MBVGMm46iJJBHPg4WrzzGFl
uVWmQZdyAIhASx5lVl7Xn4vV/A8JpwwBSjriF/+lsBbtt/KeCbef+aDuovoNjch9JPJgSlVSLCkv
he20sEQi0H+dah3pXd3NP6zTK42vlrwNkidhUDi3IGTsn9nLFhsOy58E7hTN6VkOqd4/Vyo83KmT
E5+1QtNVcPKcvAQJgZ+xaFMdsJWAtAXqlz2vO57/02ALVsbyfRna4jkNO8Va39DRaBa/qceqQg9a
/5ZCZNxX229xmzWj7xHB+kJzVDcQYE/w3/JOUfGOBqX9oyeaM38ClKCgRDVuew1G8buKzmpKE0T3
Uh7MNvmtwqQ2pLcbGWke4hDix7ddbcIov4uEb/nZ+9O8IkVlL3lxXPaQmietOkq9u4LgSv0H34Ob
BhZzY2omRxIMVE+XVZS1+9wvzo2CvZ0w5M8i8L5d3PBDFp2n5GJxjyYeXiPns15RjezxnIGmVFyz
5dQN4ft3fDcO1haPWX9TuD/ZslBAmVK0q2Qa8bxeqe9GGJ3weRNBNpjWJxN4ozGY650pSY9PUkZx
Q6yZMjpBU6Ef73usUgegbQAoj1UHyRZmGg4OZ1cgaXKbqlOiAiBPmeL0lbPdb+XrL7R5zkauMpWP
Fp31GFcTOEkLerfJGQL+Q+N3nI3nIHk6iIjUDJq19JRTHubznTPJhIShCDT91oInzCPw8RNY3bzp
DIKZ15zdHK+WZp5zBiXPqRGyXVRsWK429uM6sUGijWrmPZaUrXhZFPKGwNN4miMbotG0rL4+u/x6
PVLxedzu33yGCuu3HlBNV/2/2GtYt9hKLSx6aHpNyWYyeft/p14BjowMzHl3RufEIaWelYyD7yg2
9wY+pT5Y6rnMegyQEM9mDjKiXwORO6X3vLVW4rCi9o2oFXEDZ10K41yNGQzbErdBpbsz1nEZ8zi2
Muw/IyNATqUafzXK4knl7ZK1tW+DcPCPbpsRKlFA8gH+WnzjuWxs9gqOPpoFkciNxkSJulbWMJSd
PDaLlG5TWr3ERCM2IH0dj1YLi9M7SR9WhZzT4rHxqUgkmcWnUIDca5vv+5AUgl+ituSqK6OTDGOD
w2IPCTTv4TpNlAL3BauiLFydhfs7OfIiyR5wKIUTrTtL1ie3nlrUCvlYrD2H4wJWMIQ1H4r3f0nt
vvlDmjCk2BbmB7f/HKsmSMFv2sW8JKY1zOgxp68MOk8i2F2S+OdaXRwtKp2SvwXCZxgW78nYSFeU
7BRTyaPfo2U563YZ8sjQuK6ZhqbiUxi4Cg5uYcxDSLNNuc0Y9Nhsd3zsBG2tpzcndRPrDGnsZHe5
bywwpy0nzl9upWBQC6Nx17EeYNxw0rJNWpByFS6ft7uMBIHTPe2jfV32aTpzwPROfr/KQawemKty
sbc1Zeo8s1pvrmjP5pQ98aG38L03t+qi6XciMvIpXTfJ3OWz6ud7/8Vj2sBQ47H/LCuQIgo6wvFE
s7udPY93r8B3SELBZNhssBsQaBnbPyHduQlkczXLYHmCLH5aNpJwvpdMiAXyketSpUmiGzXJHMMd
BnViUchU8S+ZGcyVzRZP1aFmnkBrJwvdfrCQFn4znFgTeyukYnuwPPAIuREJfGJMCmBcpKvC75Kc
nFhleRE54tAVS8AxmNNCEb/mWXCy+PgZkCk7Nh5TkafdynMdtaPV2c92qfV1sAonYHUTgHsX6cU6
YWulHXfNBnIUss22aKWyZsBW8aNY4Crrq78uTQ+Og7xeOSA1GR0x1xO7GhZ3uv2C7rynUG+xdupd
Ws77vbjdg/IhKN2cpA4zx6X4PfIwzqLQnLGWbL1KAb/2Xj4gzFNZNRZ7SeIAt5fiNwf71MzQ318f
esJVmrtWjc4xdPrQl7oBb6pjSonnBH0etYysWyct1dc91/GKm+9nz9cd/zx3d4SDmXskqE8Q6vVq
7UkJTgBDmtjDORBgGZYDvUMVjBGooK7yo+g20Tis4jylFcCODLMRufBCWIpVRy+U/HzeD1Rv6hHZ
OYov2rARnUVVImePtGUGqgJGXjhUNtscQaEcdt92gG41zZavNEI2ax8ZGsXnmI3Ip86LvCV9pLST
VLjdoFtEyFRn9ZIviCuU0EamhVwNx9HXbvFijyQ8OFgNc224ncTOYe4GKCpc1dQEO0KblTdKGact
85vTUF2jppyJa1Rn/vicG8BLTb9WCz15ngrj4Wno/imp1uDkg6qZCOGC0UK7qMKn8H9U1IJL986H
XNI81GVswhzn2w320f+/0wtB2W99MBHSTI1DzDZ8lRzusgDZjKTsMzObIU1F2TFmPuofEyfdKm3q
YAw+dILjNJMvd7w8RUjKCT4mOKvKVUpoxzdkLMPss+WTmVlx7sB93FE6v9Rr+542o8JWh7xoYi0Y
XZKzk13cwRUNQ28t5whhKFUh7IxB6nQGVoyp37PnbzJ8fyTPM8/RZ2kpjrFFkPaZWQrH8uJQJoYl
D/dIz9nllksQUB4RdSfJw+hT57qsCVFzw18z3Lmq7JtUSSgSQtVoIMdVnvvf6WFBNwgOoFuBN+jz
bSNBAkOA+K+BZTumVqxs1MFHm4nNmzyFWH5dpuS0YvgPZHSuqcqMoeXHFDMIrFnACffDDYflLmKw
xwIrzR+D2dbdd+mkc8yPAHzkURcFRZhyBs3XF90UpaQpnFfoPAxmkixMx7gfFlUK1/DBXZeFzo05
FHqT0+Pi7UZuKP2c22DFw29BD5kaIEZG+tWZA/vOLp3PcW+BeM6Z+pF1Wb+eCTZCRF7zNDUF5Obk
6lqGOtcqTZHIBSUv5b0DsKhZLN2jKKYS43HDBEg0nr9+nJwvO8Y4xnH6prLXbbIt3TTGEt9LXT9c
/pJmYRv3n9ArgWCVhRMaMIX7Qug2cXvBCdhxOqmeHb8ELQXO6yDK0HpGK2WtDA9iEl82Y2xT/1GQ
cJz+Pk98sX9ldDoZY55ExT7t1jS7PGt5I74KoaLQWclN3kINhDyIk10HB3TCPYPfdSNpUZvIaXAq
uIII/M5HP4TLtc0dc8ar1E1zC3Yr35AvdZa7h+ItRs3/rkru8m9ARlgEdGwFmYkURYiDnXlMLUBc
b9tZJXWMeVmZLUragM7/INlM4O83wW13Er6LbX/KACVjQhxpOhlvC1MtuA99ptXou9g5jozhjxpP
EteO5Mv05obmud1KZHtQ/qgVAPqhmJKizZOhRJ/+pYvE417Y/8Chto2thoSmPgKYq9wuVtpoAIm6
vMkAdGpS8G5yi68rX0oDDoArcm1xv7sKvuDSSgBZ/u9iha10+5sf04t0rexOysqTu3srZGD3I5LU
rj8ofWbaviiXqWvt/h6qYdc0vS95+FTjs7xzZu9G9TiIsyRV+O8rLIVPxD9KI0Xxrr4G9QL8BJeI
6+/XJ0oIyo0mMCQQmwwlLS+iZdq9yCqDTS+M39dE4eeXNNgooZXq0FoWU7NfinX3X0x0oNCQv5+1
JfgaMW2+7B27w6zh8TS3iYccvxuy7fX2iqzhusaVb/33RSoqBKDSLJ6eIlHhap4Z35195z16CfTX
4f6D+RNvWNgUMzPZ4b0AluCLA6cuTNg4CWKBVl7UL+ad2R6SewlSR6bMToqAA4uSnBHWx0JiTa8a
yvWsLj1dImmqlj0aIL73rpGtwdI2fXoxtwYMQBJCepNXYzT3La40LGGuxWlYjphrUOvBgN8kozv6
oAAP0SkJInFTegFCm1anneFSTfORDba9t4TRaaVhh1w2Np2dcdw55pLeR0J+Yd3z+e5nczBJ2Orl
TRRxEFBS3OVsxG5URdL2c6ch9oA4Np0ytASfuF97w+NiHfioPoBkXDKpozqJJYtD7i8iHkwTH/k2
EyN9salvVvsbAATAV3nkpGnEMqCCUF6wig0cji5R2YUkGJX1iK8fhckRgh3Cyu3lANYaL4zxNqZX
ROyOb79l0R2lcfJqM0IHM30S8ju+UuAz9oGLnXvIZ219irSMI6i3NIOdC/EyPtrpouHAo4qNTdel
TsrXmYW/30+vSIjqGk3/feZpFAt+OM6USefQsduXZJZQiuKkYUmedLe9zHYgwZXO6siazXbZrcbS
xaCw8yj0dMy7DX+f2YbBKHoyeUfOcNgwwDd/xhKFqeFR06C2gh7M5JyZ/nEkZvqLxlZX/Eb4sKXX
Im6gVN3ioU7xVoJAg/zxPsv2D+JjNIdzaQKIqDRxBgVKeNrCuTSEPYJJ5HoGrLn0Y86Oa9GIHcL9
0ZOkZTuq3UAkNd0KRvm0nX1r8F5CfyJtc/4kdqqXaleoIVxPnlSlXCJrTwsHJ2Pxm5qcjwPCvqFX
5qVPYBhnsjqn2nvdCIUiU9BxerTbYQrlIav2j3r85qoZZIYYfCHTUbZKKkrocfTijEJM21H7fLwJ
k1nlMGgcG9AQDaf74vlaRnAM88nJ7hbsTvjhUcvHQxOTktNpV3vt+cOPX+lxYstg3kmNFBCqc6bL
SVFZ0Qh0DPA+1m/DxU7dfQ6LPTZKMOpoGXgtUF0GSUs/O//WDJm+sTF+gcBc0HFzmeWhqws/xhrI
dhS6ANRfGIJHioPMtsSvG86tOs8CORT1xxAp8ahjcrGRCwIqiS6M89z/vF0qCR40hG+/TCRyFr6I
ctyAnSM9lLqGu2OGKiP3JdAzoymxIU35Oh98wM0BNIRrc/3U6liBcoAQ7tiYGuN8JIQEBRV9X/PZ
DaH+HTx+YagND/e7V3tRnQyQrXgEsxLy6wyrRbhfuZ01cIEUkjXqLXPG55qBTvtnZlX2RrfeOfET
UOonhTGJM+IsVLvZ00fBp1sE3puHT9KLUHTikLNuKA98p6NwqIWqK+v7KEj6I2zwwq8hypvavwqh
rN95DgotnU8bYb/4qO3XNl6v1IsGSrPH5rlJ4yHfLQE1zJ326OVXK8gZX/LFRryQjHneAoVMV+rY
HyDLHPuJtjl6ermaaBgaomt8hHiQkFXjjo9S1axtZnTbNbBCHu7qEC0dMrzR+yCoCuRjUcrBzP6K
fkbZsDKWEALCtX3kxbIwkDGKNin4j1EuNUm2NPlMHQb05DDk7S69cCtLxIyD/TVXJEyRgboOyUjN
9kG719svjRcLAMBpb3b+kuXe7dcqWCQD5Q9IUneQqg9uP9NvVH6TheZmb1Cxn23WkpG698WBk44k
+MYVTc0wfxleI010c5tkwNFbe45TvQ1e9W8NvxXXJeuA2tnmCcF6muNp9lNX6OIWToU9Qupw+0yn
7TBLO/uXRflPAJEJoiIPaWzZHaQdfFDWV+3RStXhLzbXE57gFoylAyaUHHsuyiS6/AZW+FoFS7o/
Qynf1q7uJNdrAYhGPeB/r2OXoT6gNsNjjxwq377pyM4PVzrmeSFYJkYDPvaSHvIqSs2pznj7+ZQv
2AjlntDt98nZhUl9V0AoYNHLM6AdCnDIefZZyyCuFEL73ORriW6jNVk9sanqMZevSNHr2W4T64Dm
rRvoi7jj6HOvcA+nFICbOd1tEsCGF+tZVXZ8GUiTlKX/zIAoUTrp9hjW/DwJ6vNVgVZkVSzAyHXk
fNTKu1fpiQZm0kcYM/N7xQZUQQbeJFognjQs9KxOptjVujAu3FImDfmXL3l1eQKrcgfirgWG1TZH
2FmoZ3J9sgHQMhlRjHb+BjznPm7K8U5byoXv0ic1vBZHAwthkzQB8JxRz7jSvhHXyUnm5t1xtYVg
SeNKZCmNym/4VrCNNRMosbqZi9EwDsTZGk5ahDMdFFqHvdPPUSIj9qFtn8WlCcbsrMXYsT60hm1O
5gczAOw05sfl0YYt0TZ/eKPwxk+eM8oAVuzC6Xcepn69Heq6umPdVSOME+78QfUEhBTyG59lqyqB
xuG6gSt1zuxbV0zuGNKMfBX4Ulox6Y2ZIf36l9RclZU/Wt7IEHvhDO8TSEO4anl9oD7ixu/aoFkB
CiS77Mi+y78DW8pO9mHkeVUjC0+OlLeMCZww2cGFK7tUlxr+zbt7BOa1iy71JIbtIisR0DOcRk2z
5aCOQA6+ih7rULY1uEP1gQn2SiS7V8UdLS1ys5tXFSPr/NDGwsK7t4hWcFhiZanma0+PIJK1Nf7Y
DDo7GoP29GvQItKy/6XxsyBOBjX53hYy0Wj5w/QY4NqvlP0E9Hf5Rkio9+w9JwHAa68hRDR2rfXO
Tg0B5DtYi93LApRQkIyGcobbKBi4dEp3a1gbT3mncSr77+5eoLGp7crmVBc2+F3YvjQDfjlj4WcW
rbb5Mjp60vd6mU8iXA4U2Rys6IQCTYuYfGTA1mEfsWeY5rPXr7vkxX9KE/QNg4NYjztQiwSL5vlB
qNl5BGTBApiCR9bK/s++ODUyLKqC2quD0DJFIHuGm8nRrcScG/kxnfIxlYKxmXQZBlGCx2MmFAqF
zn3j8lsY8/YEB2Ii24uavYEUdVh8i7+bNebza/qQHOeLtC/vFzrvhOVZ1NXB5q8Ruojv1W82G4We
WlpbNkqMTYGAwl8dSj1EpHovw1BMGvzoQMv8RnIpkRGLe8WbOFZ9GyvvqF6fHqgLo3SnWwwYL6US
LwyZacmc+SL/BQ1B3juX4vD3Go8s8D1GbqvjXizLpm4qIPI6kd4tHDUyt7b/KdxLYBXLz6ckCH3Y
DmO2UIitN8nFaiPT/bP80Ah3Qn78YEGQ70/YQKT2LHWtIAyxNb7OUCOTxPJSeZQgRTmQZ7vg1P/1
TBkBK0GSSViXvpZ1nFQfQc9UVWeMA7rz5RDPiV2BvVfLuhaj4XFjRvG9SV8/aLfzdE+G/pc/a1b4
OEWgpJixjPuVfzMjE2a9/1FIiVVPMdJFZ8FNum7J5hz+FnPrSAqwjfteU4J+OqhMsXkHAQjs6SOd
FiGtkRXj+oHYj64CCf+XHLBKdYZTvhqdR7uxIv7P6j9l9y/tPVY8IrSTBO1VOqDCM6hsHs/cQ2xW
J9pk1CKO3nUEaO1RgJhjjEsvkzCGFYAsl5060Vl6CoxdpiSNZ1Zz7nQFmkJDgYBz1cKG+D73VmCf
9AIuyg+DO+LvYOzzcZemtzLdqHr5XxnnbgPNSloNelldihuyfryaQA0QtUlrRzL3H9uQhyal1zfP
pGZsLNmjvfvXKD6OkwCG3bR75dWtanKes2sIiBXgMMouLCBJ/8/9PAB+MNvWq7WJywRLZwEW6IYX
PiVBuyqCw+HbcJV3FAQhu8ePVfmhC0NdiLqqWhlqZddYGLz/2bsdkd9FMdneUJcAy2FE9SNtUunJ
g8BOxiS+zXOZN6giPPkxlRahUFR+vk1J2sERmO6KR6+BGWDTxG7OstBzKrj/js1G2692iJOeoXls
pLyXuObuT+zvFwbjeEjDEajahQleVHh5GrBI4DOpYwnVnlE8uZAeTJryl3mgDyOnBVdxyI9rH/UT
gzcwS7YU1q1u0r4LdynFGm54Okqd0QWwK3XVuVDSvk4jaRyf0mkGv38PfGb69N+u0lFfHO3bGuNu
/P+HozxBoNivyazt8iW/zglF5/mR2bLcwDf60SN/QJDyvYb4uYDhDoxV8kY6C6Opm7p4JXqokTih
2RcbLCwiIbAPHhjc0aEOBss0VkhMBMSuqVO1UJfhtU6Sg2IZBMNRVLkcB2/uYnNjdbAMcjsP/ipC
39gBHFBV7sv9A8yz5E1JsE1hiLzc5w87l1ADqP1J1e4ydqcmkBPJgxuqw9q0Rszp/IByvoapthAF
VHzRbh16AWQv/ZVED7U0Zb15WS70grnv/4BdxtGPHw+uMhbF6rkb3Gg22n+148BOtx+zz++yzZ4+
eRxSrXV+SDKHDvcy1TBh6Y1UobT+H8QuU5xU3eHPcnR0i1NlTZiWBnn7sAtfP0vk0GlrGowbmaQN
yhPedJUTwheVPwcdkVCm1+M/Tm3gmpFITaH5NRYDSIBhL1w/W3g8vdO1eZYe7CapoISml9/ZqNxl
k0faFhX2p/crrUqN6H/tMAh8L38K7yG2uCkMX35AvNyvGBc9oJfwhEW0Or46qzHHsSTwnkUHssAV
wxFTT4US6gAxKwRrPowU1QIpgh1JqIt+ruLHdzAaIhLhNpt+jszFfT6/6qkbgzpcbynAajuawBfX
OLlQT39dsJnykMPemQvZH8aJ3Qan3zn51POERa4BjZ5zol/5UtGvUW1W+obr3F2b9tkKwiWtOojM
1vKKDNz21+HiG9WKkpeFaQJPV3CurHMbqQTXjNUgyFuMhYaMC2nFagQ6C97MkkpyGtV33zWNjPxF
HpO/lFXMuTdfWUS4aEK7A0HYlDJwcu0DvDCB7j9zL/KysU9LV9hFFySfbk6HsYevZXJjofhNQt6e
VRUP34lfwoi5M/fDWeetaz6V84LSWmysKcTdJ1gEUxQBjNzHDA2YPHmES4A7ZZyrtXjaYb7AYKsN
9SY+4P5aQYUA5ipWrZnLppPyRe6UWbnguqERFPlr/gf6e/ZVNmT6zEQZxmMeydvtQ1hjzjmOAsHX
jhCW7osxppwW2legBpIy87XE7QnmQ0Jg83mxxPCkxwSlqi8zTV4fBiu9q5ZEbnrSSCc81UEUR9V5
o5vPDKawGZZbHp/0YhFZy/AwbP1Hl4ZOdg/f6Pj/+Gey6rWeWEnMYQ6+Eemk+az/Cd3lDC/1FwsY
WuG3tc6kfvmdjyjQOHNkxd/ToAEUdS5dvXYMZhGGegsICXx7iWMvHLm5T/6EY3E05Vylmnv1jPfA
l/4bC9m/39BvSCMAGW9eaUzUcI9DeiK+KidbZ0D+IUtscICmSA2kkKXFF+QaB3Sqmf8R5ZzIY+Rk
N/0bcy1VOBG2R7WKVnvOM/Qv1tllACLxFy2ri0wBzFHVnW37hpeBjtFA9Gjq2ZSGlAbnIhKhermz
VKFPaZsf70dj6sT49ViHt4Re6+A1G2fg0acLlWp4HDVxcB6FK3ZxeAa51euCEH2sSGjkuPF6CvmO
MZGmr1GN0e2rxMjG7cZyvcTJ2x4y2GaPoeFyUTNBs9Yi1dACu66igltL2GJyVOBak9r4gXZDGxNf
I0jR4puqaF8XfUaVyViyWVk6DlatNJUAV47xAKvTxRlshuKahR6GKzGMXGm3dhx96Ub6gHCUqKGB
KhOe/6r3JBTG+axDPhO9XpFCkVy641W6BrrPjsaE0FVrZBZjRln0gTKNM8xxUpQ3/u1hNGVfOw4f
U7VVlT86OVi7aEo+orqutdLLHTeoRcCn/RC70iQwFJu8hLE9Y7LApeNVAZBTrZLYQWnm+2sI900U
VRO2ZlFVC5CTykUyok/srTpn21i9Xx9qS4ts9GLdlajjJUJ+byAh7AFjtKeBS+iW2Fze3wky9sPa
uWS9lSypR9snph/1malEQ/dLgyL6bX2zI7GjB/2eMyR1LKMaMThMkkWZE2KZis5AhVaaPqayDusX
svgIHYC+seT3XznUCBe9zmOUoyJ/SFLgOdF483MfpwNwEJcQIfjMNFUzLn90mpbb7RJbeJHhmyNE
RBSQ3LW2PwM3UKew0awtcx8xlXdDxO4Z94ScdMQyjTc76/jYR81NemSHmgiTgkuFn5UMfNG1mCHy
Jf12vB2ks2TCKDwbzgJj6T6hv6T3DuqtNK8n96WGj4HvaXR/sB1qoWS3yOL+rBY1csamBVu18KkO
xAgLTCfEnCTlg90W1JmEk2PD7Qanx5GAT2I0xqxm7sPetushbXxqT9mkm1Kjz/rLHVkghLcpwMGc
xyqCGwpuzSKEXe9tav+GBhdMALwwce0TaLDujghjIHL0TZyUrppJOcG2xpZsStnziv254uIKrmX4
MlxN8sQnRAYThMX0d6pGrze68Re12ffVqHJEGcQ4/bWNqWuErVykfoXAeea3wcCnKRTkxMWdLlh6
wDjStPZAxRj5d5aVLwCZV5QGRRWEvUyaJ5CuckLVKCRLG8aX2sD6d9CUsErSB8eDi+LdZ36MwO65
zgVXNrfZLnRBrUgv39Hyk8Bmlop7wu9WsW/zVo246o6yiF72Qvs27tbppWMBlqsOj8lhvpbCZuL/
9jDpgGvnCKZ2HpkCjrz0p8wKX0Za3Y8xjwl1zb2FuO8zxoWERYiwh4kMNL4och8/ToJrYPHybwag
K9RADMBvFnYa7RmI/GYC/OunHl4ov5J8ePbQZ7TgKyK7a44Xv5jV+skRk7k2LbVYeI2ABLSIaIUT
mv+6pW3weHDZx1jnCcFB9HlZp4cicMISz0EkRmR6wFb0SGQJi45D0kw1bUQ1I+Tu3qLq96xtaFkS
nIlgXFZ0pw3JuBIZP8begyyc+D4K0JuLQnsw8LShMdyn0PObdFn5obkqhAHk7Qa474xBjoZMIepg
oF34neSBUk+UHYW5rE1AiDtQBj/42+u/PIWTOCBASaVulHWxSTJzRg6Z2jLYgyvyEGpJ1YKOb++9
XrPv3FLcn42e3UwLogqAA6q8O0JBbLZnCgn/+QrBMUfmQeREfFOY+Sq+xwLUnzDahethu4wQk5r7
cm3l4VsvJrmW1b0ujFlPzCR/d1nmyQO9Jnp2LvGeCy4PuXlHB1J1XShe3D3ukLjjHUDMNe5xh5Is
1RUviB+/a51xFr4m6odhqyMAqn+jXLO+Fdvz/EDWMdr3UlbyRNFvFBOJEIkErfi2p0tqnSiFxo+h
g1tDnIKvk0RWQCnQGrXOKk6Qe3r1nlgVsgeGFmSI6W9xKRK10uJBDE+t8W61T/sWjnSBFrmehCYN
Up2YSm17sTDLc+/UVD9a30FKIiX7Bjd6tt4d98BxhQpuO5/Zwg3rvHjwpPxUkLm4rzAId/yQS/Uz
ebHNDA3DC/w7MPLAkJcaY7mdmSYrsfv1spyqXBtPPpR0M1wQnWGXeTFgZOeo9EW7xxMW6B6+JAY9
XHKLXnezv3QppjkEe2/J9DV+Rye7rDrx5AE5ybvPHz/id4bWCBSeN0OR+gsykFqtSyBGy9/+p7cc
PGj9b1T++E/PjS4u8smJuyFXAg9JKrE4/0Z4c/JsKkgHgRZGLWKxrqWTUR4YXKLQIeEoVkKT3W3O
UjsC0BZqV9Q6daeBUZwDSzEAzFb+Sxkwvjs60C9oWBTCnKbqbfmi4Awk0qHGRHTx5Y2IBRYoijNS
NQ95JoaPvTVUrfx5K9zYkW8vQN9Y+0JysjMbQ27vX1wuZZsy8ObuOKzgCqb+SRcJ7vK08We+JT7G
Fq4cdNekvcpeD6O86+/siFL8I0unBxXEQzyyngUR9HWai7G+5A6OZSuUQDJ1ssP3HVl6kKiB4C+I
Xoudx8qSpCMh1n3gPrvM7hismHg4H5ft1jdYaOL84OwFWf7DWqlp2tvJgJ9wZjH96F+Lm60qnKRZ
MYGtb8tKjtL/qUaxogPemqIbel9v7A7f+Uc+HvM5EItGSl2fX+YJY5fb/CVi+ko0TN4X2pNlyRsk
q6nKjUVm/DVYHstSThlmAaQ16mJ4OajZrO1BIu/3j6tTyk/ISlUG2aRlO/Q/VpVERqFfireSnI+c
3fW5GZSM9YnkQIoWo5UilqmtFaSKsJSv6Yqadmc96RVbk6FBASyjFbvdfUCRf2EY0oQ7F3xEmvki
FvXz6KXozgxVaB1tDsszr0f+bMvIjWbDBMJFWRVFvWbvEvMVtcHyaBHIA8PCtQQp9zeoSTi2RMKx
g8DP+NtqB8je4NNzg9YnniNPFmwhhxS/ysm0HMd2yQJySN7RuAEL06K9luRF2I+JSEY2Q34O/i06
hM4eH2Z2ULHbOoasBu9yJBit3rYdDi8Q3QuekJEKLdCwErThcFxtVWe7DkPdhe2gFH9fxzzmCdXY
mv9usZ+vpp9gtwyt5jFZRsxBrM9bLzAZiql1nG8JT54C9XJHV5umFcka9yxYJ8Kv5ooO5v0srYqz
iYZuGCkbOqOYAznZ3jkMDzG05O5XoenvN0fBGypry8Yz8n+zBGAmBRrbSLzZWQ4lDJaI/d2QxWLi
NBN1CXhuSiV/neLvHoEMUlhnLHCCy8ls/tL5nOCJB0jCyKIMoPDt+Jav/oFAd59LlzMTAl4462NS
+LkeAkPxDzbTkFSNyBHNSCSFH447mFZe1B8rvpRVJI7DPlzVVEcrBbKjXUeIaQQ+IUsuol1asIcc
SY7/7Di6e4gkUElpW7Qp0afyKtGy6dFjA/LzHtLkTB72TTkkNue+butO8EPulnZUUpptjvihV9eP
uKQvLgafv7jQkZYzS/4j57A1EqWA05sPblwqBSUw54xb6j6cHQkyjhKAqdxuj861vr24RuC9Vhqm
GCKo1nGy2uf4LK5Ov4X5DZB8Jsc1n6LZjc2O1tQSVJvpwTGxSFyWyjuL9BjFaj5lPP4RN68JHjtZ
696oVhh0hPYN1NLtOqRRwsaBeX+bmVHd8zaKID1jsRI3L2Q3Q3BO9AtPJJLAIBokDzCijM34SRtt
em8JhL03rEGlmjSAktHz32pIJ8WibeeR9VGPGFIjMjp5Y9zVllIUncGn8mjdVU+xJ9M/dIR6yCB3
fzwq+uJOQWZJn9CtnWHJaomz6f90sdSxtGRXGeX0qISPVJ3away/ivOWbVg8+UfXt1+Oh09BRVaF
APR+Zp+bZyBUxrueZdYROiTgdBN44+XBjqlFDK/rRNCvcnQ7iOTu3mmGQyP8uvtu3hC7IM49sUuY
lnuZMO31sSkj+Vg+wwzh75yvgeoK7W7zgKFkSg3XkDVDLrPKklA4vZhEK9gVmBKO2YF322js7P7P
UJ85zw1iCPzrgIZO7a5vHz+nqE+27ThyZ9AZffxvwV+Q9/Fy7CwlMmcDaBKkHityNV1NvFq9PUnw
Osmw0dI6rBiAomU53nyZdRCmh3mVN0/wZN++bU8iTvVEdNBoGxwSPgV3jEEVUYO3Y+voLG79Xrqu
CnoGq7BlL437bkzkVbGO2SvrdR0YnIc0sC1oQyE9S1xacFKCRpO3QHpkV+NYYELxIgp+KMLTEsSW
xs6CR8RJlJi262SDj2kA/YVofq8QToZAGV/09cwDvk4XudTSbMcbdhx1KiVg/PgnSDbgbiQkkqlL
pVQgpt0OGi5/mLoPhYL+IvNyQJj30LL3QARq/RFce8uP9a+moeBF283TINqU54n2hWsaVU0YSN9L
v1fqtWQNUBn1ch+IlsB5u3PdKewYOhZapY6i6zYfddUBiGoWa0ealzhqMFsK+tr94nkkiVDZSKV5
9C1+oMrdLB09v7+hQ7n6qkDyCVA1SctFeJYAHt8zbIdjW4M3FeWCSQ3nJ83l1xOzp9PF857GZeqQ
4uuZAPBOZ1NoKGmYO/bGKiS3zJ8JntedAWp5GKLwqyQnLt1U9rD9Tt+8YBLngLUq7haTWKhyNMbi
DfX+FB7knVg7rC9kjBwdq4ltg7Ilp7ah+NB4c2b4lL2uxI68h4jYAHDkyIhgf4SsmVEJZZc5IMNd
jOLRQLq8yD73LOke5hG3JKNKYcytCBUBD/PCgwO3BVsBzttvzfibacNnYpV6mOGAg9LBhsac748u
OJclGqoOAKAQ9OI3UTJ8O6T9VpzQGiFNuzt/Zk1g1u06eCN2L/CImKTp1ySJEz8IeGA499qhhHMJ
zhBdoIh+4eaU7F9KgecegiHRjSmxhhcHwyVCZDT6VwOMFnJXzI9IwqKZaDtuE4sazsGvzYBzuj0e
BrMauY0MNkqrMxFCQ9POidiiDGwqN7tS/96931PF8FrZXxtBpHrU84dUgty55TDceezzmq+wFqav
SVpt5jPj+2LzDCk06BgrcjY8yncwz3kY4FtVz0xiZkWFvyVm10cY5gZupZ71+rCVDdWi0kg0+dvM
78aEdIrrwO73xl4HccpoX3nqdYRYN3Gh81Lxh3lDG6UUzWSGUm7qpi2ylTSx2zxaXWJNEYlkdlD9
aeQAMvicNRWAtIZt65yoe9nSUBNIrlRyCIZZgQCcdGYFgtAW7WjTIGqSDg3jvkS5cR5TD0tL9NiS
F2qo9Jf0I5xU3E/R8BBTr1jP47pWsXVwyZb9zzCNMy3vo22qA+jTMcvf/qT1DANv0X15pIiN1eLa
oMOiyy2jNEJMtHQTk8ZHX24eQSc6Y1mBiiHSgTAOUMfvTDLrFb+BUyHfCT0YPb1j39Qk78mmfyuq
1hBBrhIuBcayxpswgVlpPvJVProZNrMa6aEwvzV4Xn8s3oYfj+zL+pibpuoHssg5ZkS7OMPUif7X
NrzbnrvjmpXJn5Ge/WCtZVDwckD6o2MR3sUYpoJpimUmbb4xsNCDtIc0njcuRW3Cg5WXZ09M7/uy
dqqAnqkQAI/+GdA6i3yAYxmdkOaYrhIqU2N2gShohsAWSRGI3MsNqUtjkCUwKevy2sCYWlNyhBYi
zpNRVVpTh65kLHiPdBCIr2iVOs4XuKRFyhD1nWNlYC0LMQ1VKG02EZkugEIrtQ8dwjF5+revKDXH
A6az4MlvPfZUwbD5Ghc8B3pQxV/otDYgwIEawLzJGuigEKqLmP9//4mW5WCT2Bykv5ZA5dS7N/d5
4iB2LNSCqTV1+Luxp8PgivB7pe3evEq+gis7zJcrwWY85VQ8fzKZusHSgqfvx6OiJYq+KKf1uQDR
E3QS9zLFiOT1WZ10QbNfmkHR6wZzwbqKqCW83YSWsY0idby2O/QBZ2ZdFIVCbEu/ukAaZLx8ppQq
7ZZbee8Uqd7Adzf9CWPh0oIMF5a9jBalzx7vpQmJNLN2HlOmeok28TLHpYD0GI6z0eBxVzUZD5+3
xk5g/mB0mgNpeFvhJ0roj4npH78J63sdmDVJxxN0aHeKZeMFhC2pHuQwFjM/3XMjNxWUky5GxBVb
Rzbdx6uN/vrLDb+rO6rKjJ/c6kBhZfQekPfJoOnDENxBrtypKYLB4KtJdg769FOHJATbUmDnck85
Mc03tzdMOOoIfhyw4E3dM6K83eh2Jj39ktY9sKdUyk/3J2MAOqYrbv7hOVkX9jn33eYuAs/Vlyjb
1J4zEim1qMuuRX2WdP9BrkkKBrkettEsJh036Rh+CE1iLCmbGOhfaQMKa+ZeWVYwsJdp0VxjLK+e
vYUofNL2f7NCoPYbOmdMKyMq4SbBWvtBqFsa0OPnmTsuXriIdrdJmw++X8aGMChzDiDDhTlU+jSd
3TqwKsB1RBa6hVcWiF0pqDWLpgCM2T4wJzyqdWNNJcVsmVkvXRQ6w+pskdhHSE3UuVvc3tno8JQK
RebyYs6sR8jHCGavHBh3MjmkF5o5yt/1kHDBR1eO+dPg5o3I9eEmTtwQmM5xn18FJ9rWQxD0ay0s
NBXUYoBd2W68pKmby8E29pahdzWk06emvuc4PMoTo/zEupcgfaOkBCAY5wiDbRl7YfiC2Bv7uaZ4
ZJOwIfcVb9dL6g4YmOtO2MCUhwj8XvC8iPiq90fVCgeifLXppZYKe6x5DD69rgRAYL1NNvVn/c/w
bN6BWr0/roBFA4D55xhWYI4yo5tTXr168wS7ogLCoUkiecZ6/zLkOOv301ZSfZ0LJ8sa2uLupWbJ
xRsJZpl8UXL2v2crukWdwN4FVa3YyKB45NmTo/z4Ym31oyuUJiPQEyqxZrCAxFU98y5v/e7PHwpd
WfsB9VSh9EhL/5SKZQbdfvpDhKkuUlX33jT9me0lOq2kJvBL5RDvdqgL5O1AfA4q+uc0HCwuDokz
Mtm2LIjyGWhJdfgUocZTuoBVZOAsFuvDNfX4uFxWQK8loKF7ukpSssho0gJ69k2RBQYQRlEeKcq6
7i4+xLoXgNJjM7OdzdxKdGgikEI9X7WpL6Bht8jfQIcZEA+uZ7VRlyaYookrH8DV4kpj0d8VNgSX
VyX/opzEh2xw4dbCmjyRpFXAZblrSlSDlm93DrlRqkqq1IA9BgkkLOqjvtK+lG5Kz6w3YthXCzQq
3wyB670+Dyck0+rOLCeuTdpDlOaGVjJ82s4XjPo62ZbKwRAZxwf2zsoVkPk+6E+WnuBLosRXH41E
PLnN3R5BNQ58s3txhsf228KtexSFivcj2ufjpPH/Y3rx8oRNIbAMFxQzMFpM8KrLRoZQBbmv8WHf
/KE2I/wUhrBGxMskoNd2r/tXNrVgBZaXuzB2FeCjdLOoc7aD+ZbWXQuYDJC3NS8FS+O2kxGhiyCX
4xcGRLuEzA1hHnbHsYgusCIWQRq+dMu4GLCrhsdgNWlfJnIyz+dRX6qq9TTKBOcv7QbqfvICwYWv
2/gARptN3KXetKxvo7yZI71hgvwycRE9Q4rMizMrMJ/JqvwF63ftJ0wt/FsOPxc65XhZfh1fFCgJ
yQ0WeoRLWvDwZlRLzLaBQ+sncHXr5BomCl3cf3JJldpo8W4TB5mr6KV7cXv5VxsEfbZSt4+IFRzp
h1+9JdpP2aTkqPeTtBF0sJ/u6GH8KqpN+PfwBv7gdJXTHAN7fNzmeiLxfJ5qmCZvOU6gFXnHTeoW
UwjZCvDDdq1usNdgRoxHXRMcKxA7KuJRFpvLXVj519CYR6ftwmekbvV4ImyqkOhxFVyLZlOSJ/48
avud1wDnZI4gbG9NcmYBlw9tCpT/EQf3i4YRXm6I/qP+NlcqM2MK1MJWkc2hiZNFo8VuFOz/zGlJ
GWLXP/HfKUvsPtzXSd91uYiPYIV7gHHp3tGebvM7sPkEPthAm+mRL4iXM9x4YRurl9X8UadnYNUo
yQ0hw5rCqPcNNtFlgKwB7gGuU1SaA0ZmQKuR+jQCrRsoCbg5BtBTr4wCYdgHXCA3QMsxbIG5i0y+
bsQuZE3wFIYRtL/POz0qUYUhwfIzdX9IbsijyV0p//p0V3mFA7gC1vcV6LyJI5/WO83Nltn7ili8
PD5My2bLKvOrkXsHmPJnXcS/9Y7rTQZJmiXUsli802DGCMbZaK9y/YMmzep7ViEDOE8Dhj8eFnqy
f6ypUpmUxi7o8szxsc+w2eViZP3U/AJ+roQBOlGMCjkvgYbDAl52vKwPmS11QJWcWtR0E69oJ4tf
+dXAX58EFlcJCrYcTmvFeuYJsZPxcOBvfq3ok6UBHMTyZWQ/UaW5RcOQGNV2RoOhm/kS77rOZlun
bu2v9qNHvzSJGddYEicK3rbki0ALl9MfPVIVTaYlyP+A7eDgMXis7bnbcrhU4Z9SByngMhQt1ix0
+MeVCDkRKZM0lSxNwseDutnMcOLdaE95skUbAiGhKc9QzqYCfYeEvyKK9nxeLTUP/Qi2pMjEh7Do
MNuEZnmSkwjR8e5VL4UJLZ90fDeNuWEntQzRgQHQzqHNpADLwNY0wFwxTSrPmB7QecvYdKr1iM97
B0Ov+R7DBtJNLNEqZjjrZ5ioz6sk+GxSePr+oePmyImsp1FzgyG0d3RdFJt/NXcRc//iHJ21nM8/
tlg9aTnKRMLMiNn7JiRjH2S500xnLGamwYzcycNZf9AZWPF7ch6fwV89uaUlcy1Y/iyiOFuoF1sK
qd0sfsneG7Dst4M+Jsw/pQxEXObxPGh7DzT0qFVOGQSQmrtwv94hPT4iwOR1XNY0Ew6gz6Nb/0n6
Uo0WQCKi4gim5AsESIdI5aQsHjmrfgWhwEAm4lqG+lDp9v3hMJFxZPnRxDip5MrEVqE97/k6NdKd
rW0+qn/VQF2efO9VQBFjDcjNStZsxV0qFV93GZdpOAKN9j/ZHaqY1d12EigmNywTG19lH6Hp7DZy
/tv8bkdn2B53h9OZW1M+DI5R4lQ1743gCinJ2NA04kLDoIJWMdw+Sj0AGtlpmlwn6ZOhla98qKrQ
Vbv5k6QIhoZ+yIYzcgN/SCB089IFA3Vd9oYvlAT8IG/pPZ11V+ykJ9+dw2idlhhiKVADPbul2pMb
4Uj5CZOaZNHyAQgGhtS9DxmG408HzbhM634f0jps9somEbxhN4d/pk7nMJw9B4JtWv2UIXqUPIIY
ft/XXaqA/JRQFAs3xOmQlXeiR9ehz3Ww6AeP+s41q/PwH975CoEwC5q+BEzbg4caWavKfJM+Kitl
bIY6g8hnQC6znXeAa62s/cI875axxwxXXnmbOxEe08b/MXRIqwbcYMcNNYzLWvLt6HaqH9JhCLbY
khLznGqV3HCyl7mPLauSVTex+88wFSZezL9murLhwZj6MR757Hog/kwGaDt+os3InXmoK2fYVAiF
yRcpQcRM2p1rx2b+/VZEfmUJKmSyxpLTLw96ybX4/rmg2V0NYpBU5tZxZQnRNpYk68XfIw2NXFgr
JuS0k9a8tni+aOBCd7SJEXNesDJTjdXQfatAUGsgp7h9D227kaXmMX7c8megYslk6+yNu4cBlQRL
E31x4s5++ozkDEhChENeHo6r+vBAT7bwXMrsOLkgLdjAd9kD2LiCqKIxAyNr22GA+Maxkg9W+k8B
Oei1hXHBOQkKbR4Kyf5mDAihX9bnqF32UhTHItVUjooLGbzp+T5jGMaDD4qUYsB+MQ23ZAkvgBhb
bX6SdXub2cPVUivbNfqDAhxL3RRK5Cr7bCzAVlAMC4wVNfSsdEbwc3FYJp/cXVCW1U/Cg43Si4SW
eLTgfhoVbEekRk2NGeE9eREaI0ny0cinH41st9hZlO1o5NxE6Kf8/5mIShCK6cApGjoXhNsqzC1U
Sx+2gS21h0S6pI6HmYxYTgMa8vIM9zJEjbK+OeVve6+HiscAuXr2vtFLqFjFEvmOeRW/1WZHrbol
fpiO9okOqLvqQGhhAeeH5762r35RatXrv2wIW3yjD6G5K3dWk0qIE3+CtJg+DpcuwAQM/xSdEXTl
I7wkCBT4lAQ+Qlc8nMayDQAYk2CHFCeG1QiEuGWAlb6Ys1z/+VPVckL8YIv63480qiZKc6IsK7g/
8CWqIH8nwc1J7w0/Wr5fyAvjYJIBEt1AT17d/bJs+1MOYXEAsqgsTEjDdzQz/MDEJjz8VjvnHXjH
4kHxRxtUBVFvMMDd2UTryqCYkhZJuA4g0pAHmwJbcT1YGzapyAn++V+NMILOocJZCAZ9wDHZH/EL
lkngE3nhm/ELHfM/2+D3MsF2KNSvm00j9CXjxncTAznTDllixBzBMl4jokHkv4S5q860ZLAM9pa2
sEfDWSnsGKyAdMhfE7imGKDxGulhTG2pkQt3yaW2UYTzRN/GRPaZz3WnD62UlCPbnt5nqs1lvDED
WhBWmCHxk8cxIllc3Aeh8zgKM1WjKxPt/kSVZm1OV54NZXcrerJUcmXtYg5/kI5DG8JuOiV1BBd5
+oaMl1i25GE+wq+mbGRO/AbdSccA3TWhYvrfUcxeXo5YfY0krCTFHuTM647zdSPBE37h71VjoqTN
UPFgzu3WbR97MCjCh+XrTBT8jEDVhPLzCtr+vIgXkxqYSeBV4WBwhazWhgH9BM5bLmuVaX9mr8vE
DO41OcyW04n+3+ztOLw70Scmxoe39iphM23MWt3XF3BFXIVXEkyiAO8TixnIJuj1ehjTINQ51TdJ
WK5+ktBenX8u+YBqAp2KaEgIZdw8pdjAmMm9qduUif/aVhNetO2V9Tlg4SqzGXKdd5TJcsJeRUCF
qx8OduPfQNQ+ag0Zc+FHAMclcK4+MuDrNYKzHmLDy4yeqnHqHnDAIQYmBNh+ON/f6qUk6SwOt1f2
Xl4h4taGLZ7+yXEg/gAR+Q4glHS6N+eVlS+OCEUDfHxWdJW47DL6MOezHA60sMlJV0vuQvBqXMUq
HM28P9CsMd6VUExMhOmpwmoRP311srsYBEWPBe+jfGskMJ6qMkd1eqwne+/kG5jD3JR3MlxVA/JR
cQJlZW9eybjTa8r3N1fpg0V9wqpeEHfy9HwzAqyrhSgA/NNWzK9x1KfXf2wFios3d4317sXPdhrM
scXb0q9HaKGlp48us0IHO6T2ZPVQ4PFfQv/8E653tKP26mgfOIyC3Yrw/NMhaz8OQQk++hh2UTiM
ZYYPm+tVxX6rkpKaB5e/P6aMgjufcA1HfaJ0E7rNWDgVdLQuhz/zNXdrT05geH3nExO1Yv19uNN2
HWF05clU4CppXLk8WQNyX72drCHu/N5K1K9+1XGJ67pTK7ZJYuhr1salQqoa3ksYj0KuL1dmGiVK
B7Il71er53X6QA0jfxP68pHg1q5OOFhbF7iPyv5+iWAhRigpsY1YViHUDB3GNDNVtTJeddV/yH3X
wcBSLnoRNiOzAvZWZ/xi+h4ZrFifnZUpvbtbshS6S+sb34FlcaMRRmVvCTwq/fLJnFBfpqZDKeaZ
ykb6L33uhpoZJ272ys8XG4VWYSMC498Nh9Wg2jFSQ7BQCgFLyyLqG/I2wpRKHlNz5m8BVLLJCc/L
YD0akMa5Z4WPHctLrb0FLXpA4fN3TMW5ZxIiXEDgM35aClDMo4XJOFdce6e1NDbDpN5KIdry3iHh
CZ/3WcMERmDIMe5AtfSSGdEwLVuzjb3lGV64BzSKgLnllJFtK8OUScdTjTnRsGhIt4joI2amVlx/
Cg3bQNPB/Z8q7ID8ch9K2Q7J/PtRVYjyy0zX5CSOZZ9jdwkcqsSS5oD32s5PjDlrnHtVhT5Ewulq
ongx8pNSuQtCwTJ9w9xr4tU+cvEZG5KNyZ+JiCgWe+m6sBdsB5OGgPbe8aNg6GdU3mRX2Fp7wMdz
LIE3vIW/jZ5x+dy1o7DuqES6j/aEt32QBTmVmOoi/ogT9GieNMnrdZYtXCe2BG6Hi12YhHC67ouA
yGRgAIIbjRs130/ntp9F8NCx0xgLx9qdF3A3vbv03VfIP8hfTDfD6QjCj6f2N0MZ5LHlIYm6mMuQ
TpEMFFPWZtmxaLmA9KkJbhQCrO9CYhL5jAF25ONuY23tLC7ZSWmFHGgNwh+O6PU1HkCqylaqcINS
piSxh8rt5LCIuv2W26Qm8q0iDANqkxsTzGf1CzOx6BrMCB/v3dkIs4QluliW0y2yAHZG3Q5HwCHB
NHHqVIjImuVCh6WrSaniU8pKyBWiDvmzOIZPAHnSfQBW6nUGsdkn/gwq/JhM6PqrjRHcl4dN8stF
aX9gSzJfawjmP6AlaCCfXiI3nOPRSJMDKGj7sh4mbB/mO6Wem/JzJ58snSwL343LiPkHkTPuN9sq
BfzcZwMRVFCLg5cAx7ltqoYzcqkEM80GTO7yNsOmmZ4GFNrJwI/GOzSxQvVQ7B550XMQG6t+F7rH
cO8YU3KB6VV0YOtK1GVfKnLTmySFjMJD9ZLDqVc3EW9F6ko2dlHmy7r0nOnNUXCPlgno5e75h8o7
+cudZfPqqnLJzYrkUlfgjyeCsEg1hG1w1i+Ig4jE6uSXhLJ3bIm1pDuvIFaOAdQ6h8E/kW9wk46q
W7NsyMxDN1JRp3Lh6hHSkEep+dPwfTS+Ni7/8tUC5OJsQGJnGaETXqZ4mlXemaazw47H4Ui5dLn0
JnUtlBAG+5bTTsmkRhO6/h/YOGJ+fF6Z0mneTT03WEZWsPgRpT9UYPCBCNnpUgPhXKNoG9/XgVXH
9gfYwk51QpJdvCD7bnaZKDp+VPSS50SAOcMOrK4iiQfTz0y0rQoMvofv8jgSHXkhGAnvFT5KfBaK
uJPQM0M/QKodvjbHkgroXhkQh3OWat9ESiPf8IN/rb4dkANogjBW4/4vDFsXlIu8plJ7N6LY/F5a
3jV9Kx8tUqViZCL6/duRwtrMgF5NvVr2nthPkN0ncRZ2jtEIc504OUvboPlzYOVambVgaIIc7Lqf
l9FHrCPmm4P4tto5PXFSCDBwmTm0GiN4C+fB/nmQrYIsWzXQbA6VpDgnrOPFvS6H9RUIiEo1Fbmp
Z5QrTEyhJ2OfQLDTaOPYWa7GxHl6jwSkhsrYl4a5TurjtzUfHcIflyc1kvLFMr9/kw1Aqzyzw940
fSprVuYrdV35MkWrAWMASrt0od8mLBrIp2NMU8MvS24UDFDc5H5VkQS92q5mLzvTqaOP1TDf8/yP
Fhkxbq43bhkpFUYIn8a4RPYTdcn0ADV6cDOP70L/56tzPk/CO/X+e0YE+7Ub2WMyC8uTwG7DduIw
cA8T4xpoaDVZxRELh6AEHC/X5uFzWFubPxnj48wc5il/mCd2tUxI6+NJZLFN5RjGjvyJKZWd45fA
xBjX24E6kvz7/dAPC9z1S/BTJnnovnXu5nO/y+v27MQpdP9Kq0eyIuZkNW1fq4Oan15N6oJJ9xmU
frNjsjBzBrxliGy6Lt3KW2D1u57BAt+tyD+PSm08vvtoWy14uEqn3HPtgmYeyfdkppfebvzvwSqN
vu/sntxjBUHObApEJLyzgoWPFDy8EPSgLz3dhMeO/cVOzKF9KS3JrXUpCsRUU9hUDHSO6TLLg3nP
ADFzOjzrDEx0X4WD7zWlQwvFt/NR4+LAo67prDNB8UTNqhR/oEbnnOYZ/e8loJ2bJZbShabidqLI
2ErguoHemR1UGx9oodMUfwZgUjJkhdixoxP4I0fLNmXFmDrZ+Azk1Sxm3TEY1UW3SPV3eJ0Qv0SE
HXBtzjoYoiBlYXX8vpRjKOT7QsEdruRSAwgAuQVNm5rzcyXHKnfhoAKC/EKzRclCTxItZkQkvf9D
ZdDBaXxgtWi1svSaozHX88U+nKaYNOAODlF3uCOdP0Axaikv/xQ8snuJ4+E6BLGVAXBqEboIWs+r
H1oQpK27klm0ZbMFKY08au+2v9cKLdeyBzpIgJkt07uSiXyyUiGmdmXyBCsqwpLkFmLSf6HPKCv/
Av5lG/62Luir19h4lCsbf9g7PQrUI1w1mtjomE+FXL3XEKf1XSXxqsHx9+aQzlKWi1CzOFeyTESz
79mPBycVmUjfVf4m+wySjmFUBTQ2mG0cf/9zdEAP/zKIaFEnJ5icYNR+9QDK4znZeBrw38Q11c3x
NSgupop8NA0fXo7Phx+F+jD7Aq71eSINwzBR3trrbPtPWdf+7nRr7FA2o45bkmWyyVNkbGSFkUK/
3LYZTnqHvJKU0fer6tT1Hc25htiPZjAXWAL7CdK7ujPFyFit0k1LAUcmduwKhq7TSfpNF3IJj1Np
VzzGkF8BGpof5GHzsyThGpdLPWgTQkNWiZVzOGgwMlyoLEBYYEu10lQR9hL7sTLxQdhdAzfgLoHx
Jn8Cda3YO/riGrG6OY1nLD4eatg/CLZsnH9wzV50b57Vp7tFggwjuQ8zbsQ8D4Liezgsi/K3M9df
G+1oE2jmMjrJS8+7bws7waebqOXi4zbtyetwDHPbzBER9sUmcjaA202nOeTMzmWFOVY7IKOiOqRt
DuVnIgtX1a4lBittNeuhx15VcBy8vFKDC8Zkp09d3+zjntmmDx/UN1cC3mbGR5Ilnq6BW/L0KXn+
0u9l0tizf9x4OsYWuvxhPbSPNwi26+wRIgMCM5aLWbWfc4yBFZfxefdOgoNAZtENaJ+1t5CSvH51
MkM1nMyvZcMkL10vbRbBgObyg58R+R5fOpwlvfP7UiWOZ8m+oQ18WZs6lqnxGY6Vpy5IofnJjEUP
+IDfKxhLAVUIqFBnvJaJtczVas9t7TgFBOTh/ojdFB6kB27GqCUh+1INHHkYGiP3RtS+z6bVhWZz
h0E14ZwHY2De68UvPEKBBwe0R1GUG+HjQg0Ij6ItCpo+gPgOUS1JI/xPTViOatwgz5HQ/X+V0YV2
l7aLez0z7T50aQkgklwocfiQ1BveE5Qs7B/P/U9ld9KPwByryVXRKCcB2xcRGCJyf+sXg2IreZCf
uI6bjAsz0A74C9M7V7yGFGXAIP5qIqEEBfHjczz/q7MfmvSgHQubiM6rgS59R+0yeeJnDmI0BLCQ
rYpdON1Gwl12aB2L9q+QRAL6+dXCp23mGTei2Q2vDkF6FXiHEClYa7tCDeahuneLN5Ij0aeX5P3X
+NkYsQ7vb6xnyMjbZp3pzLIgUaqs525eVaLcRSi8skTDrmg/fyx/4Mb3kFMBIfm5GtD+85Gm9zoj
mVGW9wgNrsOfLbDLECI2gMX5uid564F0KP9bZMBDr5Z9t2OABSOH9rU5PFpeZlOZ06Cj9CuJJ3iY
NfEHhjP1fjJLvxBjYF0Zu5KWRKRkLglDav21OnlEvZinoEE2cNVOcI0EJIpqn/XsSlZXjS1X1RgM
e0MuYp0DxkOfg1Fh4nqUQTQvkJG6nKlEMUP4MR2+KtPKFlyh7WI8mE2I2nAkEpcTLPEJ96DM3VXj
ogqd9NamhUV7/LAjU5jF8WDwyauN9wX/1kt9zrMr5D/M9xNEQBYBARhmg+RPkFAsg8DWC2cmd518
bDpt6ep3YQ2eRFVdIjVR7kjjQoG4vWotV4A+TPWGqun6Jrfo3/0o+lYPO/TCLgxx69PHZ9BVBgIk
d61lda1nQNuvmPPD7MmYRwwO0vgDUf0R9O6YWpg1rr4LJ6H/fYqnU9r7yYa6ELqVS2663meY4eA0
+jb6VfPVnyrqtgBBtFHHoqQk8Ui8bbaNkJh+jQ/0l67Ty+P+xLf+Z0D5Lzhb/OwyDq5U9gitphTK
sCdoLE+VQ/sXj2vJPR7jtqPc9vRNnRweLVqqVrEXGQs2YH9XQi5dDrzdsCsYJCc/rosUW6/8KcQx
Lspw5COfNDQFBJs4vOHCpVehURn4xn+2zQOSnd1djl6qWQkYs37VPecS3CUY9gY8R33vSt76W9zB
Hh8XP3/wbKkaoWW8H5dYrrd/BMiTDPArKTjmT8KU0VVflnjnP4ruzD1VyLezUaHC0Cp1WcmdgMqW
BgH4ST72fH6rWT+MHElbeXVZ1wsXg/zHKd8+G+X/8NUUT4Zu6GR2L4KF6xBPp3qSDEoOSfEOeXs2
RrLniJuNMbROCI/g6sWb4KNmZuAn52kjsuq379pQG3omILjE4G2eh4Hp5EW5bXWaLMPlgbHAYHlH
9LP3yKZog6obWg8dWBXJmChCXi8AOd0VZWjFj7SeughFcWfHKKjZGOguj2h21NNbzed5woxeuDP4
dcpvtn1hwOIp8CekEqwV+3qMI+WT5BHgWXO4koR6VKRu3eDXhQOd1TvliFoB6Xex+jpv9r/oO0EV
NA5DkB4P6H1aOoPN0x8GMYul9noCLP7PwcT8JvUXvU8D6mCt9tFJGomY+3jExdmAS33BbPoG8TNw
oVrVanLl2wJOrxLKHgUXrpuy2dmOfmLAS/92ZE7H59ngPRg8KhKV4+S0K1fHIdra36kA3EpVFO3U
soGC/Pyab4UF5eCDWKP9+35GLOCyP4dtBQrAKJYsgwFBJoWffUTLHf8yY0GzNYRtoYdbKW3h6UDF
aTbA3tK/bZ0z/9pRqka9/ZZGPkU1bUBhyEuGkDi+3g1Vyx47jYtPhLJCnB+qX4n9dgydBFbu/gnD
LFrXIFUAEaS5V5nBMnQ3TarwRbE8oWxRKWYCq1gwKpk1U7EkH69Cuar5xQIOpNGqzBXp+IUXeIc6
MXbcv+WiWOZ9/ZsayYYnEqtnHKFEdtNWsJQgSui59+1UMrqqyTr79ivAcGdgicISvyAp8mg9AuHg
aPYJmhnzsv1DwRT8gecgzn776qmVZtSinhrPwu2lOxeyfQ7tMys5ktC8jxzgTMcOkhZKSQVOLBVw
x6uxHe8y7JXnyXi7nCTOgMQuWixRNPoXf+JXl1dohcK2C23SVIe9uIi3VqjwYk3ixfE4kNYr96WV
reDiwO3d5w2GY+nz8ErRQfXZxUJd0ZWPSKJJwjZEFG0wj0HZniRONiIOcjfl1Q22CQpMKmemqPzD
/dPxmjohiAJ9eR0uLouTPkD+WW/nexZI0YpKCoJs529pubDI7JRhtb2VAxvo6c2kxND/npTw3btR
XJmLdnaaR3kkSfUCSbM/ucn7aKt5atV6Vma1bI9RpNsMNlIl1GZal1jK51ICZlrCmke5R5U1VD62
v1qG9nzGd0DgQGh1YwCLMoQdlxiuhyXW3OKONNCO7sTBi9xbJ/ONnCuELOP4tkSXpAEZHeB9Znzh
zbkO5Y66DLHk+C0LE9kACIZEoJgyl7hodHcXD0tFyznhIjqOUTR6RA/wDVUCKJ0HQYhlhwi3FqOE
P4eMs70Mx/aZJ0UsNSjwzobK6oe3lp9wAvsNEqoKpAKZlz+NKoWr3oPH3wlvAoEaO2vsS1GWtb8I
hHT7doJ+TY5vmx6KBkQ1OA1/G4OmQ7/bbhkB7S6AE/ThKT6nCy4fdtILxdFp75HLMnq/NgHJY2xc
xEkgVA241pV93577jNmDqeg5fE42t6c6RxPBiUI5+7cD3yoNDDs9ry/+wjP8G86B5tSz5GcLwf5z
XcKxzLqmAGLn2O4TCcJrsGeGrB3Xft6vECel5bIGHjPlmCI+WLmxfueJIfheJ1o+knLl2SN/bq7q
YIifAi+ADNK6cudYmbMnk7ftUu+faNkRbiWASWZlAqMnS5XaQinF1PoKJYMkZ5FQNs/z5qXwE78z
QIpKAngaym3+2uxpdeATPIQXha5Q4u7zcBffo3RxDT1aGENEvGK3ct4n3LrFEPaQOdvUszyjSyk3
zeYK0/DthUbjSIYTAT/R/MSRp5xnGe97+m9hQ/y3+cTqIFXxmtUjLohH3gMuMKiy7+46dGnn3S1R
wLhr9FOQdCrU2F1ZiOQPMBwtX6NS4b1Z1HwSBMvr5tY6PXue3wpY/vjUZmPewRiLzdD+EC64Q/R1
gZdqP3fNHM33GAisgTO50BpVkiUKfBqi6KFuTFiQ4aA9Zu5u9ZOkWCk2iekb2UB9KkndrOSpxdrR
JBFnj4jGBhvv4BAXMixmEW89RXVvH6UL3Xp1FxSIDjtXlUS2unO5E/WObxf5/xhK8gyrjpWOvddH
9Off82C9Zyl2YPru0RSLGcgLNyX9tDHHIH7GntDqZhAPv9FkP9/4VjqJihBXSiP3x9Kv+a/lTlBR
psJ8xaqo+JUgw9FyAYZD/yldfUvPV4k1GoNNNaCEWUwzGojalxusb8wpa2w9FhxrG60NQCm3AA4B
Fsm1K40E7fcthI4odDO/fFKfb5ZOtmvmNvJn/RBEFdx6PzeDcuno9+M725xJae8Q8EVa8HIliFSi
YC/uUbN3zvojt701dt6sQJ7iPKWv3vSmLcanxnYAT+mCSX4v7vz8tCnvAVtLMJa1v+MoNmSeZY2X
s4KpUAsvXej0eE42e7BVLPD7JEa+V0UA8+X4sEL3TWymMlJqV1sdmytIH+3/yjjB1nyBhD9f6SKN
uKQbzBNehoAdYW2ppmqyXJTjQG29faKIrlSxrYQnMwnzfZWEOwOwLlHgZ5DlcZJRChHTAuYPtqZU
SrDh3y4piobSxgih0nPUumNjthcALr8Ge3uRhCp66U9ilhIxD1l7JXH8/UaVEulWuicSLqwrGUPv
i1r7gJe11dYlb3cnz67VwchSu/qtplCOCoT+aFv87LG305DCtj0AmgPYhw1RBPpXxBZTCvSCkSv+
asJoRhp0/y7jF/xAYdeH43RZPO6YsdpO/JeW6+9/a81NmQDqk+fZoAftagDDP13Pqi56O7qdKD3Z
9YFwrpYY8yQnAvIZ3rMRGmpHSBgOmNQmgyeFn3DXh4+C+NHBJ5xaeqM8mx9Ef4qggpBWH2E03IjA
EfaGSBtyVS9EiXIdYa0LuLv6Gd4mbWs2oVrGVjWzIl+GqiDbdERp7+IeQvreA/hPtBMJGMhca1/T
SQ+s2agS3t0hVW6R3RbFNq/QB7BF3ZV1+CTrg4qNGlcWsiXgTRwWTi0Bv2GnSqqxc81ByN5I6WJ6
zmbA8LqcQHmjJBhL3CvLtcLi9iBRfUY93ihntgS3QTMVBgXgn+kEh6pLp0sX9XHUwkJZxWdj0ZYg
YG5hDOFEFEd4HxwHv6XGHwe1Jdqiwnv9ju43B2oIHJcQdpzO8YEY7chLJff8729iEp/SrRPe3yVv
mo4ZlHxKIg2s1IUPWquCxTl3tNBMWqxs7AQzBFueYTxm2xmDpEEFXC5+AxDzEMzjvnEFr+d1mQY3
sBhHqjohwDpGYprPV2+agV55AB6i6xi70XfH8A+vo9R4l66BKiEv6vOrtnvHRA/NJr8UgHKBrw9B
CvUSCt5ymiWHwaGNaZGrNdB3MqLGP9vp/Slho6EfyyHiRErLeViNEgFQf9k5xlZWK/AKZeX6nvkg
YbfhDd9dH17YYo2RVAekOgyAnVxZlqFVWeql1muu+y5h1Tbr0pjFgREwkmhVNcuLMDEtKo+bw4If
78f2K1SQrgTZ6hvhfdSnEzuHKzavVJwT9gI+6naI+5HbMtvwSNOyyvvs/MUZ0s0leTzTcfhFsrwC
cg24yJbaz3Y695JsSBlXe3KrjwIzObz/qRfxG/BoQ5xNj2SaVsYNt52H0baObPWPvMU1UUMfbheJ
/K//DrJuAYSlX38HMpS853AjTGNhqBpuNQV3jHRsSoKl9PtK94si+aK9mfiGx05/+8no37N5jJnb
knEe9Il3+KhT5ozIJqwJ6PNFi2tmsab1lye/FrXxFRbmk684bO5tL1pOp3HjBghyMKP97dLjfTot
+yIqEJsbnP7TLQ6+K7Zi0/WuvCO8giVGaqHQVo+bofo7fKrRepVfeknOg7fC22YW27U131H/2OhK
9uZiQXmX5Bcbarsa1wsbNYrP1FNwEYDG0akC+wRwU8L6ZxkBsuKJeF2clgjYgHNtsglgUBB76Ztb
cTlP0hsC7Lh8Cv+rUQLZwPLNWVPNWLLg/8W/ZDmhPUXTJcTlbeF4drLoClLWVEzIdr1FvYhrxn1U
kMkll3wU+Kcw+2UVUrYAihrWEFRi0wnhkC8fAXBSNjqHXXZtL075oa7QvSMPW34tLTFJjtit307A
p77452Tg71Po5g+RWxrd0dhA1gRziyMzsfiIdOgSJYcTrNz9Cg2KJHSsiE5THdkEFNVoKs7sCP8W
8kMtycVg/4Q+cjs+2WEJ8uvCRmnPtBKR+CymmSuO7pSKmE9PiOzyg7wUVtGZ7usddkUCPHnuU+TB
ae6XLz07p+FN7/muFfMBJWXFj6xJKqFdVTfXdPp7NAejkdr8TZuydkqzfowmQr3ThAYNgqaHG8om
JP6+czB33Zaafgb2wFb0ZTdwR0NQ8eK0d4N0ILXmY1dcYWn94vl/YZL0HBJ13PVpJ6r0+0BQtwVr
FHH/0xr1EprKON8/H8FLKgjyg7GsiMPEOX0mCxPwoqEFgJjz12oIJBvSPXknW1T6iqrci49M+Nnw
H3LcmjjK7A29Xh9y4IY4e3z1UIrDVwRJM/Zt27YI1RGDghCIl7Fn636o+JBPFjJkdwObgkam6/Sy
xktoyYQtOp6ePCTR12JPYKTz/zB7tGV2sPQVvorSldRlY8sJoAJdXdZ5LH2QMEUx4CClhaUovtXm
xr2uyNhUIsnzKbMcu/ar/8iri6JFv5KbPj0Qe35Jz1exMaU5HxcHFoJmcRlL7Z7ytcqviAV4edoU
SJzFRSXDZObqUR2t2krMl2smTIWyQ1ELPDHPJidQVyM0lx1hebGOsyxmlPTnngqdoyOiY9sCMhnz
9C5Zl48tjLW0U6ADsxz/VsXjiMCUBJXxtHxbyVcOqulCC1wdA2CMqa+ALqqoF1NaNsTWRp3KkfWU
xPklPJ1r8UU2czZ2MQaJQIT6+5Pap9x3ZJQLwgOwo+rwkq5WMWiKYQTrA3ZJ33cJqrcjDp6e5UO5
Bvt/4lU/+Ms4mNEEELOiwwQnA/wn8flnaCBp4Dl11ci/IcEd8tRxsreFrwWIENb7rHL0abRMvzGR
LoPUsqx3yRKi5uSfjs8mezbm4WHXik7Lqebfs3GLTrb9zDTBDqBQeTU8Zkd/VcSxMejRGIno7oad
XOg4/MnGewY9mfzDMNId/WZMYK7lcepvB9iglrPd4/koCMKH+PD9TZJk3zHD9TWh/KIAGQ+aeKHY
Kazv4EYUvw0i0Qr6McFT5NygC6QyOa0UVqlgUgHCqD0sFYMy6O2k+p8HjrmEfBdxaYFCifV3p30M
3P+yD+2xfrnf9qXQiUXXGjuZ+r9O69r/5TXYZnRt8hg+ItlOdHCHoHwJNEtCfV6cNRWbiEvijm78
0WM7hKzFVfip+H24jbjGW7x7TyeivbZvGQzOkIn58hv1kWqR4rckDRVtenUH0L6pPNPAzczMmFQK
hwP3DbIUMJGaGUmqc7QzVuH5Oqrwvb2sayuqeU2ALp75WbUe95zfWHbxwdiwT3V/VF0qZzIE9oTD
vVqYTd104+GqHbuFi4hwvVwW3AjSaw2tEbo25avkucJb8tL8PvkjPhTF9Zoo5o1z9gNxPxSkyfVd
/IUiX8b9M7DXQYUnSUKKsFnQIPEnpBrkPneOHHmfrs5OjkthU0Tb0iWOWfbgANZ2hUtTeRLxGe+R
jq3nMSjf33W9xs1kbgljrfh6kts+pk4oS70LXPtENwjgNtWrZgzSjOveWjI5uf03tOrJcEf57G/F
8JTm//aYR1dAzxchnCD6d+c4c7lXkp+igarLu8KsHL4joGEi7GaEqAdBMB+QnNnCRUnqnTovsRiO
cZmEQvWa727OXF1GFnn4YSoaA/FaSOklyxuoAKRYJJdWXSBjXY8Z8ZstxY8pWB0EFW0AMGMo7Fbv
Ao19X4uP0El91XTcVAGZhlaVPYxTPyKncrGVkmlCt2fQIbssGa5AaWyzukWWUsWmLsWH3atFV+qQ
h6y5pAxQBHRzRjVD2XgeVRMcmcBmj3ay7PCUnvnnwgIUwi8Xwt9K94hinVxKSEqDlteGkAoRmb+D
hta/Ik1UhAJp4T2g5SUxlh+6luCp8lA7qAHs73x7dun1F6Nv3zdshd+zQhidWYhtWRnFcZA8eOX4
irsiYnEx4KCZ3xvBTAlVjNmeyx98GacCdB5sxH6wYf1ks4Nu0KUDHw90rHARz/dGvyutw7/mqYzW
d0W/cwFW6Pj6IZnHfoq2pQ6u3OLPqn68hnHDRZrT7xx8HDqID30RsY1hzonhIUMfQ402yHNe35rX
9lyqOF9qnj3CFX997YGW7aHP5veNtsO2ltlvBNLxmrnr3FBhm4KV0VeooljKlYHUh36w65StNP16
wwfC08yYSoZzPkUdVXt8nVzu0pdehCx99WkYDcYFXLqFXQPTSDomQPmq4V4P0CtcN+L7p33KCxyt
xJYMccpc3/9DnvETg5AwE7xCMUgfogxVVACIaZ7eY62wyFM+YS0VFouRLxnj44GhPPwdjtcuzu7P
Iu/6+4J6LjKGrUZ8o8OP8JjygaWqvubmIL99X7AbH4VQSRALk6YrgdOGjIgodSFLFnDPUmX/9MDr
qH+pJPDelG/yiw40+i+Ehzofxula5GKX2P2c9TuifdY2VshpllHSX1JoYJffh04ehcxVLO+NUaBj
/nwq7Zbl2gErcd/nPOlVg11JSeGNz/knXJA4DHTOKVcsQiFDt9c2XKI6udrQB8kYhvVE3TfD+dPJ
0vI70HZ6AbnvsdxR+GnGTXNE6BiIiO9A9hlz6835H3ZvMozkXySrYqA5wwtXaY8lf8RCk3J/XhRd
t6XZPzOdJYKexU4f39DWdxeq2QsAoBhKwuRDd++vuWpN6HYTQzD3f6Xg0YyWRev7lZ4WSeHf1w5q
bB1/pxgeeDLHspfgh5PrPiMYTd7lMmO3LQXaZwE4xlfsVZrDUHUlwhkcntcUY9B1ifjUzu4D1Pa9
Hw4Q/JlXHzxSE+K7jSoaCco626j6NOuRfI/7HOOxr286w+HcxB40Tppeb3WFuPYf51B0pvvhvbet
TyMCwFsOVy1mS6F61IpagY6zOKNstmivlAzdhtQEc7FFM63nxI9F2CGpfO61b4Duw3qBh2Hd4hqY
LMt04dRBkzolGGspPVJVM62yuaruWv0JQfqpLUn/F4o4rjDIKEDYnehwd2otEjnydU/zRZhwaW3D
+02r9GF/hh+IjdviD3auYjl7jquz9AkbSG0nacQNXt1O9XqaKdEUaujcGzPn8jJRHYwQ0BkGPJOx
nN6Hys9ihBI97X5TweLVd3P79wXgyj2twX4L1PfSu7PzR8sGv39GQsWJnJlgXUkPUomut4y2FMsS
h7rpMrd4ZE4J59qwlp5M58BN7T7IEn4uyhcqGJGJV8AtIM9jVcwPamHCXQZITYqGyJqMyIIKoT+Y
yJ5PnFGt+D6sEqlbTiZ7fZmoTjsT2PDuZa5xSh68s6WoPnKsZADrCkV9IG3Gve01WdDs5w4nMEEz
pS2mxWVnOawiJ4QnKetKlGeX7+biTgTt/J34lzByLwjY8AgMU+eN/iRRcSUWJ640F7KMa1Y0GhCk
TzLJgEpNfoyJ04/ccrnlC4nE28Kxzj4lmLNEytMt6VX25mgEtt5ws1SlPXJOzOHybfvt7YE4Y11B
+bbbL4gCOUO7QQt/TsGfCmGuxAPA0H5yl3r6+cPyvozRQ7ctxaypPcrekf8oF8mK+nK4Q2C2uORO
a5CIncY/4vaSBo9UAi0wbfoyhiLDwz97EVlLJKue2wKYOSeGL+58y13efqeEhG5qWnK7tf/8C5IZ
3NkT6PPTTy3acHsHiH7gyz8b2ZoP+1MbONrMRrVNhZSqx1NyFEAK9Zwts8ZF2VEgEtAZ6CN0aYxb
lUdAAd3fwWPGdsRkUyC9lycjdabk4WvoBYxjohHv4jokSh8FnGI22E3ada1qYpAgJAE9AwCWAeL2
RyEO7SUZoVT5W5NH16qgX27xxg8Cwig2RU03xDnRGUX3VPTeYJU+XMTuASRPvGRwZM8qdZ01Y0NJ
7uAKtSpYHjgu8gf76Gv5gwoCCGqqSbNHCVL8+6AKeRbC25iycs7XFcQ6NMPdPG6DN7nDckPxp5kI
nIT1bSqxkOkYAUXpEW2FbbwsSM1DdStDxp7NL+DCyLwL2S5691MS/0OMm+iNjaAsid17tNgent+B
tmlMCIOTVmNI3Vv3/m1Jt4/L9EP+k/L4u9PfZq3yLwbpw9d+5z5kklG52p22X4v5pxdXSXo0WhPc
dpJckdbRTdqH93Ud+l6WEL7Ev849OIoDwXxQm7+azzBoX8L1V2eUWKZwWiFr3WKjgrkS4zPCGyWW
m+WypAQGG9Hp7RkrHjdV0x6ph2FsMtIqjFbmknexFumcTJBBqLjxOTf0gEHR3BVLdBuACTn8piGR
+N/5vWCAzRktoH6MfuKlSzn7KGaixTxDtrlMM6Q4v7iH5IvyIt+0ve4SAuF3Twg/Xd+sqbgPOCyD
sz3mSAUFvWGye9217sOz/rHo9PsbFy7lVsDuFojw40bQOZ7EApi2LInwGbdWBvCTftmDgKJoHi4j
nlDEXoFH7YxAmIy2LnfYhjQVSwBMXk79N8Xi0uWDZ4vuluRO3WKzQzrafzlPVzDArpGZOJW2kyaa
Vhqc+/8iUvAUCYX51ZAGB0fKiV8aPzyaGCU1FwcGEjsz0+O/nD780wsfHAV+gSRKqQkz9PQYNKff
syH9B/9QtaobHxuPPHzkKSPXI4ULI6gE7bXkAjZYqvFf6QqhNh1xGDkHewVupt79oEKMZkrl8bTT
bl2tywGydNkMBbO1N48g68+3ioMvs4y7PNupWFpz2B7uT1uRcEhiRrjObPtPuUUT1Eiy2qTRxKja
5UiNx8VY4o8VDToDXEv3sYTNxrFHEb3erIXvs2FaoyInD+G+TxTqqjS25nTUPl7TvV9RB/+376+t
TDOZtx2is60sjIcMvWEmrJPP8pkod7VkSM7TWio/K8P8jxGGaWyfsx43TrDScdBaBVD4d9RxndCc
7yabpMvy4kP43SuCDVbpgkcwWXv7N36qOGKPQfM39V/UvmjIOLWlZE0CQVSXg7W0l3Pq3ZGc3fAa
TsQL0Q8rLBJ61U885FXlMiQ9KLt1+Vzhs6x/wCxURdZHas8gWp49X8HbHBty8s+J24VsZS2bpT7A
ac0qpCximzBLtIC1J2EFbWhwnq0Lx2caCOBUBnpRGP1e3mgvWoPY0scgOQQSIP+NM31rLmWLvMY9
tt030VgI0nElXccpjVwN5MXu5pTHtsIGNKwLxLS2UlmU6jGy3TLR3KK3y2xuiZY8gQgKfJKZR4q4
Qi3IDF6p2zdHWVx4Hjs7KXH8smgFoD8C4javUQTAp/lnNzp6Yn6egF7U2Lwd5NkaZt9F06Im+Srj
53Pdhq8/1osLm+txCGeThXYTgTEKxPAQpOiP/eDNiSBB3F+IG9x7sppBAeNDp5PmsDzw3wcFT+NB
jpYu1/mtav2ZCFBw7oZwlugFTQdpAIB6MCEl++SzWvz9tuD4lEJeAe+sGGijZTFxFYhLYreSBino
tdrB04vDS4TE4DO9ZIEqj8/s37Ou6gM94IwIu+AKiJ+xtyqewCOxDzewonqs9sd8MiKR85Cnfz87
67h11JCwFIvntpJ1kvTd81TCNVzIlfY2NbusYCuOih95Fz5sBnX6GrKLLxyYfma0szPmjMboBFvH
o3DlkMOkuT4wSUnH2eUhHVpJpToud1SI6PhywzEBOO/VvA6uoget8F7gvgUyPw/1a28YvJmPto3Q
TR2Pw33XBN+BvEtSS8dy8vGHeJblu+UsYofJZjZhM0/Xc0p0UfaI5fceoDm7Hxn5riHn1vrYuHPC
BKQVCT8Eh9MmICxs4mIavmdSldkeh14aJQ8IlIKn1j57s3GdXoc+DC3t33c+QcTX+I2j7w5sULNY
bT16ORVXnMLgbKwzDkvU/OkMEM6hJknTW8fAfxNnUm3Q8DANqsWVkQEidDAMqMx4uG2j9+t1jKNK
4bmK8tTqeNC7NGuxyBehxPIGg6cUCeWldrf+ZYm0TIINDKBpIMVjjzoKIVYcFGaPJ2kEDY2DQW6F
BJkXAojEZAj9wSrJhbOKH5qaCM77e5g3Uj+c5aLhKT5xg22AeUpiFVHvY1aLwGzc61z6oT4EaMLR
UtcVAm2FdSBR1RXrJz2avw23DWe6Y3+BO1g+c52JG5K5gFCQhP8IJBUC1wm/oZ0lXkAZBjr9WJPL
VDkEpVJnrpN1L/jrgKHtk0jMtOiyz3TG0S5ewIxuhoJDGu5nt6YYxdE1C16upmzmSA+FdUId3KY4
rg6NPnzvYaZGKJPWclETA6PIKavTJsgvgvslcqjE7Dt/fbUB62Ahi6WBgGrrFY+bVSx9/+oWda/k
4ARz3GULXccPFgscOsi6y8hvmin7zzIXOa2knlnfC8ahYiHzjSD4IsVUrBw8wCraQyJeQ1dREcEg
aX1O7mRb8OgF8oZwryMK7xKrIchJ+XtrCnTSBZuiVpXhkcIvqUZDGf7t2wRzN3Nd+taKs59/Srao
+gqjIqA5fKUIHhoU2Ug4GcBXUUxOzdCeiFOp9WRZU0w25R+QNsIifY82xCoUI1qj0hPTMYb0WgpX
tE3rDCa5qy5VK1J/UX8r44j09H68yy6GkIBK5JYgg/8d5m9FlsSIZ6+IISDI9eHdWPRINhSBmfmS
eld1HzANAD8zb3eh2D6XW9KWFXUosFpqEpEVWk3/16byXwc3CEbLxVWiZCibKKbP+ssFP2UE+q9v
GuAzCeYhKUxIKBfzYz7g4Qp1H2xizWvOaYFU0N3gaPG5TW6FyGEiDyN3ADoBrsa50ZOFI6E+BRaV
17yXCgQpgVC/THzwuu9+sxtsMJOgB5E+m+W9V4h/3uv1ZB0qUM6qJa1cwp5bHS+nM8sYqXCnoJlN
/EZFz8kWvIyKlkTVtGPiN9t/OrJdeZARWP0GRdIWJsydRUQIYlNAXZQOa5aggmJqJNUC+9hs+d4G
iUoBQCK3EElP2HJr8k1Ns94c23PE3siAB6M73RGByVKIAUVTM0OHohbpJFu7o0NQ6FRPYnAst6QB
FtRlJHM8jnFk27N/JT0r9tX3FkgOrhBaSEG5CIj2O1ztaC7BDtGbKHK58gPa1kjoRMBBEXWKpbXn
hRawt97/tfEm4BJwIMQg5yq+4Adl2LgaK+Hg0J5JHYi03lF2cn1TlXfTueY9ZcUdYouQToKPvLDS
LlHtxnfspdBIe+WIQPk/Hvqw3BLCooKtf3DyPWLtu94tp8MX/KOCiPKsAYCe0hpBbo4dHpn6IOcp
8lgqQFIl+XyWGx8uZrDcnjgeE5YJNZlOjLEff51WPBDbQTOct8/WeLv7YnWySB7TwugFxs4X9QHH
9s+BPUxMHQcUAvac5waBLtOTOgK71jwWnmEEnVFOlp85oarljURl3iMR1jJshak3RJ8nWMc6EIV3
ow12GYDC2RnrY7mWiCFYYcjcKtePyFgfTOuDP+QzFOmYpSD75Ui4MJdFY4dOrkGJ3UGX6nr27tyq
FvLoF0ZvjaPwGGg6q7ttYEbhv6SXiGUq3XlvfvVfFaiAeBMs15xfx0+uSfJUCW2ztFF0hE0YUm0k
TMI4i4egTTJV/WP7bY1XBolhSqA8Q7psIScYWN966LkyMWkBvSzAOZN+DwjE9Tz999uULPxeZJ8E
F7k//YODMSGCebNbUa//WwGEDbdjFfWuCrZJr+AC29GA1rPVepy35DcSjbdPiKZT9zS+g6KQcLK7
0uHv+nUkGyWm1ZJkJz20bPO0FQ7a/WLRyHEYyQ2dxlNnjIBwszlBqLRKkDDgbJxCVqLJvFQ3X8DX
EWofeXvqLLfcxhYEt6KvrzbcnyN/oVyuYnZk7Y3/YvIY09UqfXv7xEq5Bmk+mx3vuUPUEWcIAfOV
vTQ3Hg4JM/VSy2ldWZK2rsgFDyAQw8odrcfu0GOAvsFhr7OlvZdvIkikVgw0bwH1iCfeUk4oKenu
Z9LmvwnXLSR7pT9JhkIlJq0VvE1WjEyIppMXkle4hjkKaiSwJNJ8nFz3tWdQC6cg/AdSJZBFBk0V
5dm22gt8uhGS0Ube/DiOd166FECi5eM8IJhCUzjDkiZGZlX1nzdjK/vpWlrLSFp0d6R7+EPIvF3h
3Hn18f2xSvOwcsXBouORKcU8BBykp1DmERkhnom2Z83jXw8re7dBj4oMCBuS+NiXcJcX3eeGdrE2
XG4aCMbrsOGiTIafJqVrPrWeNP5cARXmCSt0jNenioVB5plDgXWJY5nYnEFUckLOy7yYaUpWQuC9
5kXOUbxLgGVvDxwNVuWP3EzbV5sDVGVPD3TNTdPHIsr056KAOuGGQ/dxuF1Mboq/hUInP5CbX5Af
Ej63WsHNB0C0PGGUBtjt3D+tZE9LIvPi/urQWFcJstBZ5eIcBIQ3I5A4wkV/XLovd5iiVKnp2ZIn
8gNA+pmL3kezNnZUdw/ExooWZYjJb2ZnbE+HSUX6RcvigrVw6VoitYkyvnNlXuMbZ8L9KrnHwKAE
VyAcpbyArWp6+In8tZSTGeZ/rM4OqI5cMZ2HquMraV4pcmbUeWoBWAJRqwEXYI6v2Te3AWTP0bp4
RwzymPuM9zTccfuCFtTeEPVbnORHqN3KYG4O7r8S4tUGoE+HwMTRD4HSo4mQYfCpGqi5/8RltUsn
BRvKq27y5EBllsmGkAbev8tIeXKRdUYwytCMz38ZCe7Dz8nXEsMlwM3DZMyMT50Ko6bJstp2/CeG
2tkrgR3AAW1LxrPU7dwoH8bXGDE1T+Kk/LPrSHABbVteIG4SH4BFIUrmNdCZ8vFYX8ZAlRXYdPjR
Cb7KdtIgMs1FuarL48QV3SDgbpF4GXezJ5SgmVio846Zu2KQVIVSMhdpz3aqokMxQ7nxPvPsRkNq
ouXq82sn/1Ppz/IEnRVT8q7ocuJcrCzKsgovQ4r+OGPf4sT4MgVG9GhurlGaQfuVmKE3/XlIXmBt
OdGimGNbuAoDY1BsjnOnN0GSrFYo9tWyWnZ+mE0qYeJBq4jjcHVrG6aoCl14vc1J0qic0xLqODhO
KMkIlsuQXFeRnCc913eYCenKnB04C842Q3WpIdMLyzZhC7nMJ+OHH/KqiSvuqUjcQzHRhKs+ilTY
eweHBRFzn4iX+3mZ4XNli7eUKe7xig8EChdk4KAiNkbp2zidUzuG9kMrJV6+8Q7sJYQj4omKVMhR
mVU57pewStltHXa6drHtLeV9nnsToc4z909WjKLBVr/W1drN7fmzyZFZjWT5B43SpsKFBykQI0j6
xz3CXT7K2W90wh7XjJLq0EiY81cqK/QfPRGxheIoqowRkkQe8KX71hZMu1r5C18TIeWNe/03uirJ
CmdZn8hjx4h5IeKMp+HLcluBU1RqhbNI0Im6EjxZVVd13aTc+Xr8F2yoRPrljDnIUpoyeUfocEnA
BNeYOb2P0rW0G4gljBJQsyjLDpOzZwFYYNb8Jvgi0a2mK4c/aaQWkwN6kSMY2MMo9OGiIebWF8ee
EVpdox8hnDxhGs/WWLN87X9v1li0ZHMz51cXn0ETh45vP7kc3cI2POc92gk+lHvcrNp7y+XM/Ncz
By9rbdCLPgv+ANu6b2ZUkyd3O26sh5rRjUYKi1ddNcLKHf7votfOmN+nsLUadsQt5+SkrD66eRwe
oqDYK5FVt7k3VkqsjbECb40hrht6M+JHJ6VaqtzbWgMLmSh/YmiQDnyu9tUOWpEX1B+05J74XNLw
aGgUD0VFNkstXXW7w2QfqdaVo/MVWtIj9vSXR2NEWjWo3DdpoOs4nNi4+qO/4bhpTGrDBQdBcgty
0f7AfWlTqLQLK79kEAqU9VL8nG/Vs1pgpSsIAawO0LBMda9Y/0nMnkIoX/4Oc3fkyqFpe5o4v59I
nMeP1DCzgSxyqv22nDAnsYCiW/QHm6KEdEeKMaxXZBqAw1XrMFNttAxqFuJQDSnSQZnAfaATHl+o
LcKsXjmQ6n3apUrCuAgv9U58LOLGdWnlxm1rMLv720x0shDHVzlQX3W2C0n21VfoS/syHPLayIHZ
J05nJ33IK0bHgi/STUW3Iw7vXfYDEtB/3W3rDCOrkJ2WeMGOqAitxhlI8Fs9ka/c2BnzWdFNaPab
iuiKyftMnvXeYobsjHM9Uidcdbh9eOh0AofuYnq4RpoGBhV9YifZ30t+qssF/Fgqxu6smPYPH+9m
niigIeUiuPwED5Ld/FTqjQZvD1Qi/pg9zzzNEODr4iuckX82KStqsdRAwtEix+l6dLUOJvYKymbm
l4CyPBm/7FKUNYO2h+U3/DwvqqWJ3AQKwYqq1GuP8G1wms3PXd8aCy1peJkU72eLOi+rAUZWZqVy
GI2+06Qpiby50I3HfJ9+AMH+xsFC3wCKp/38WyvHMogPtvuHvUklEOYNXA8yzN7niiSqrrAuBqov
qQ5nH7Ctmh6/DzOTPeAQVOewKM4p+PSJB7Vwugmhl6QV1tLgBqk/arJj6F7jgjuZTn0mWyrYTM5F
eY5gPoyB3qnkLMFRFlPmGY+yWS+/X1yHjuMO5cdZSM/Dgx3ZTknmrZrr67eEmFJT8B7N/YfqQ5Rw
nUDXXO3UM+4SdnFem9DHIzq1I6QKmzAeLFv/Gb1/vNi1AAmrabCULZ4U2b8lbD3FFSwhaRNCiE0N
wiBP/YsiZRMdTu6L2+RY/b0JXpvP5adWonXKzHmeYc6EYEefP+p2BHCnjOgRXkEtR0ykREHz3uVA
aTia+rdTjkSEpdy2sIGXBc/f/nRJNCFPmUKdKBjwNR6Y/LQeIAw5yi0YZCrWQDHLWhNguDOrCiko
4N/jlq1zeErI4XpfttyeUBzZjBonPyrH1+VVGHgCRoPuXuba54FhoXi/Q2vvn57SdR394dgHXruz
6Bs3HEVazIyUDr7ofgiIFf95ASlOfaeX4UHHjhuFx8IinrUD5LCz8orypCBWmDqg5oTbuinhuJOO
Ys6O1oi29OhhcjODzt7LoMMzGhrZWvUyXpBfcuGWbLXOpO0ZtU199at5zQ7sJYEktNcc9WJuHpKJ
rB9JnZ74YuMYpUfx6sPyN2RMjwnitahvchvDkvWe8KM5B3ICCJPLGRFwFgLgKSfZvnhEaejX3SEd
TKpNTRDzrvDlwgpjn2RlqFoSvgMzW3zMEPkk3aHCL6z0RbIpP/k4x3wRiHpGjkdLCJhbdn7fBJxA
38c6tF0rCuWn3TNDJrJ/iMlClUzCFZqY9O+nc/k2E2R4DoEf/PU/ceL73t6Oip5w2WqFCYcge4Qb
MZtu9XUerS8Z57/PLV7++og/CVovf/pWW5CxpGFj7y48E+CEFPtj54bhZLVffScJs+OgOMt35BUb
J5CsqxlNMkiGXA+dl2RjwgslEpnudOFw5JdrixAvEKJPxUVwynhYGIplMBkNDqL/YxH0UveZU4/f
l13Ao9ZfIXMBYSZHKoACBjABprPvYaiDDfsjBHoIO576QZmXC3fdYHoPgZo8oZz5IyFeE8gyFP8y
Ar2lcXwa2x+TrzEr9NW06N9IB9zvgH0ZlSCfnSN+xLi/3lYJazYLK/zcbKKU2Yo9oDnltEkhD0UK
4JdFVcAcTv0z30oOwTsXyhw+L6pJV8vQ90ETGThJjLHPVMR8YPsr3DooVVm2XU56lmIogW3lN3Iq
MJ4Jj5Fo0vBg8FPNsZtegEkhKUI6Q2WwHfcEi0l1B9P0zGM4D1oof+Jw/A/WIIbt7b1r7mZ2p8rv
6QqHfq69ff6Ei1vmYVUPBqXVKt6sGnQ6kKFanzc+WujsEbzymw6V2v/pHqZnX9HdFEbgXXiF4U2X
5oAdLyD65WLXO0rkj/T0a6uudWzKXybFElUVvPx9g5IR4LDQBVReu5YE5vZn6JNDCf/QJmrtQICu
QNFbTVcSzIoJXyaj/kpFamR81grcsPLZ5B/3tWt4VWJOKmEiMsH+hVFaNbZqOJSfRxdsYHfrDQzL
dPZA8cKzYIBJGGhFy4Zy6G21vB092yY3yOahqCxvNI6AhOCSU5i/bVW2iC9Vg74BbscRJFVyXHRU
XHKKx06IhgJxAJkF2phcIQMGklD9Zn/1xbE4qm1xEs8+nCQ3Z9N6kugFXzKafTM2Pkw//chpWy4x
5CpqLEpo46VQ/Uas4Lh9KS2mvTBgMpkiJ5Pt7KsmIX35K9KEJGdvOqgdseBXmXz5fKjuC0zaPKD5
ZH6sYlT0TG6Mq5+yRT8iZWWtmUsUpV7BCmbQP6Nih6w9u2N+7qLzJ5jZxXD2NVNAamZVUvGzxNeP
fGPme5iijYrvvW4/OfqmfKsg41S2PvAxUghBovWhHgoadhImGCN8WOmNDHqL01cGIlNabHu+/6Dc
9Sg7O8501iXP47cXwEdu/e+9qUm26N1n1ja0qGoLeb0GSJHQDdMTFHYkcuu+MzK6XhO4f1PjrLkJ
Bq9RTn2yf+G6tKji9qyrciJpcuV97msiNOzfJF2SBMqtoa/5VEgLlLQOQvFhRqLIzqaLwUZUFLw0
HFk+XOnTfPDM9Y+4kAEJgDAMAClIdZm0h8sVbWpTn4RI5ozPf4yVwvbyMvbLvhjgCHJCtnZIDSmi
DdyzYdCm9V5F6XwpdOG/cnbmiclCdRHnnPnSkXr09rOC+KaQLDYxNx6qwNmn/gF2NLVRTy6m4Hps
wMhR0XoW+AWNKaj8H7Nz5vUSsfOoEZO1YK2To6temGLj0DrONuv19N70PYli1eHeNO12nSTvhb0c
Db8rm2Tq+iKHhtLLhcHT891Es/GmRRcRjG1pl3RrTR2Er8x6XdvefCgMdMwWifilaxWa98MwdAwP
Il+rI2f84WeXqMb6qr4Oau3KhOw9NrWS6/spZJcsgXn9xWXmlSO5dKeGky/Gu+zsvadT6lvVNwLE
P3U1/UnuhZjqNhJuDMFdLF0CoqXbbR8v6e52P4FNHpRPJONT835uDOmLctPAimpXcn4+27U2ve3P
Mx7I6GF/WFTPpim3J7td7ieRgly7Ll+NBqD1u3OpmFb/h0Kpg77ZI1CXK7ewQVmD5K76a0//2CXk
r9+0B7w6UencLHkvkh0L3KPfDciOwHBWMPLgdEIELnf9QxNB4ALZzkRQA55GK+o8kKDx34kMiN0p
BMAwY/t3+wi4BXtuzNkHBhTY7DBOwvhac9wn8ojD1nIY/rzl20AoysupVSqiRjMErnfO/UlPzFuH
maItlSTmZgQztWirgbPWZlTnntO3XVq3SC4uvMmOarOzTnuxfx+0C1gaDQXl+3KDRYuqVgpWuUbz
M1ER7n/Txo/d6m6lo5QvCW3xt5trYmJe+N7jeChVmJ/opKxVcJTVK4gOKWXQJuwNRdJ7cpnnUOII
peA/G0g030VX7YBErU108CmLqJQ392dsC2ufArURuoNWwwYqLCTrqDeKhuYkjIeO7K8EKM3v8yzI
lIJLV6PDuaLbE/XM3cKcfbujNWR2dvDCLVnNi4OFmvsCTEZ2yYwCQu+Nv/T0sG3sCfNpcSCZ6zPP
FTMI0DNn4FsHv8l7kcvxaIMvj9BbT0StuhFgo9yoL7UPWfWIvl9BegZ9NIXjmkCmbmjw5INSax8V
RT3rxovVS5hNCk80L9V1t6th+S8Ejs5pKCv33nUQJtY5O7+bqXCNcjGihYZqxljdRjGL0LJju0I1
o63rE40jHJRNzbgviGLalDlRO4pMQd1MgkvAUY1V9H2oVGnbeVTU8LSJ4mBWwCxbK5b6LWPCyPeF
KUr+1v+Z9xni2AbHjO3h//HWKUEO4hb+WaUD49AfHCDirCSjuVsTTmowKRlfdnuBCH5tZiWldE9Q
MH9pPHew3JZqrTMLkyBL2zEpUE/t46A45XzqkXkrJr8LuN3K+25MmbA48Uv1e6awyomi4mrLDk5a
jbav4f+rIRWATcbiUcGKg0pc63xts/WSH+Ga/qw6GpfLqgAiWUw5q7QM190w1kHMFFYBZGC7+ntM
s3zT3Va/TcG9QLELLMGDnHC2u0K493YDjpA/JcbNTF82S0rMlo3A5ZylXzOSUdck0kqxtshMZxhQ
7ImBac+Q2ikbTT5Nr0a0UOYtem9MQANkT2TbWG4Fa5+grXYCbgLl4f8Bs/8HLvwVTzdiImHC8qkz
HxCOCAXbO//gWTnwW2Oj8xbTHirIviM5SwtHM7sF+yZww7j3QMuexJyRwov1Pk6pAUAomNZ99gc6
LBkWJlyRk6Oh0ROKDVeUKhfLOwfWer9Ju3SKjVthcKUmo/+dtcX3Osslz4Eip/qxv4IARRcaCCv0
GdfodO5rkpz3SWF9YROtgC+KGZ7nSp1RP4soG++d9wAWktK6xN5w6oeDJpRBZilMpKi4r1DbTxQo
0GkXgQ3IZho6zCRF5c4xCmSaRB3OV31EyWlomPHQOn3v0FqYF9DU/wSaZSPFfOXssXiyqQNXnEn+
0W6S0DQDBod/w9TX1zPwu9C1yf+sZ2M8U3/i0PIEWYfZUQ8V/OQzxSLY4l0rnZfXWRpqtEFjA76G
nDL7l7e31ILpJIYH6qdbY2SYO39kY7w6iDoow3EJCUuh6us7K7JosKiOdVtxhiYhQ2I8LUEOK/4Y
ei/6U404WMLQm9AAfM+ppS+wnAWVzu20j4oUOp2iuStt8wSl9H1cgYtIMLBnGrPy/FP/2dkxLTe+
unAAoyEmqNpTFPr22BkMMDM9CjETCPRYTyajgGD4C1w/jNMd3MQ2Aj6dcC+B+KdGPJiOOGbojAM5
CvYo2jr25+k1hVhSyEQybohU9Bk1fXAZ/fm2X5DG8QvTvomWiY0D/yUS/FcTOPCvTUKoNHrHpw7P
DQvgqzaMd4FYjrYTRW3R9+hZ17XNcibixjTmyJ16d5UkXVHHgQMk8Zzj7syBw2O7IJQ06gM4N6m/
BB6SrhZIngNY5DBg0RtlBzfMzTG9LBtqorjcM+Q7yOSytBG3mbEwr6Eu9IExI+BidFscXXnHbujk
5FeU5tOBwMDVuFZDtNFDKGIsIxlMUdgouJdipX4ngo8HlpdfTh7F9RNzGQjrckr2XYfWecG8vQmd
EqOvB6dZEsCoZsiqTGg4eaIlnH6OBoHfayeBd0lCkhfPAFhSEpnEWads7FpOfNvY1ScFdyScSYtT
aJdYumX6bFN+pGA4a8a/JCslrM8I7z8iOp6fZwfkMy/QTzqi9M7b8xFmqfKMqQYk5NEBQH6Aw4MQ
Tk/dyw4BpR6uMqPF1LH3SgY+tl7HcPdcZWhuEeuKDKnIdoDD4C0tMtAc8cYohd0YBTPEAUKueLYh
En6v9Swzm5baSVVhJBq6RA8ZQ3ORO7znUPUZqHu9Cyepw9/UOteT8NFnyuIIlrEuJEqTZJWV4epH
VlhVZ83IyIMuaJYOsSnaDFyqVuQW5GEEfMji8MCTzyDlVm1cFJ2klsi4mVDJCuZ2ITp/nn3cSqxO
sLHPVRIQrgEVHih/C/A98o95TJgkwifgGjEAES9nQw6Qk+VJXTxbUWyf3MHnCnDcAZiZoZ70oakz
Hug9FcRrCzares1u4mEkoOuu10jXOJdKx81YhKvnSCcqowK0uywwtLM1qdytzxsfqenflafKOUj7
erPVOj889jHhbTVfVMNGj8jMHS7A4gsJHKRTB6in2Tly6GZbzq01+Ptxg1D2tcd9+r7wBa/HeY42
JQdbiFYyYgf2wirez7EHCLttpZvM7CxTOj3vFUeDcbxK8rBP9ccAlEk/7OrP92tJvWweV5M9IY+c
Ca1DWoO6QMIks/U2YW5iUnK2WtFGzKBIUYyDXvp0o8tXwWUIMjHlSobuv2we75oma/5pQNSKiZGI
5JSqK+9mRH+YD/ojkY04D+ALb0F5NnMxA3C8KGZpdd4qIl4cYBtZkFw7MIIDJCcDUEl71JYbtZH8
vzQfAd7kNlQjP61LEpK4i0NOyADC+gGqlzdugT8swmmWw6M5yraEzx84R/X010+IrGTe5C4Rhn1D
tKhO//UHWtRT93EkCaw51VnvBcYjUWdUUZ6cGlWCVaQcMV0lrwDl44cgtLBhy2/O8tEZocsgIH9d
A8e6X0rkEJnHx8/TEoNrKKyt29ySDd0VCUqbLU2kcQACF+ol4dL98w+2FWraEq9ivpPX8HB175dm
aum4Jpk+ySO/vGrB37oyV1eWb9jbmUwVo0HFYQbhenzGC1TV3V25DOH5k10mBrwan6+/LGdSZtBy
QFhQSawQhUiChjPQ3YU7DEhRMzEl9qDtE4CRh75Q72Vh4ypFXkG/5DHqa9wK7YeyAwnUywp0P/TJ
+E0/hWgIbhcG9Z6yq/bf/xj2C/ZmOVi4VZJVH8zxok4y+L2pg6tgaYdLe6GkBKiwNlowqEXsLX9E
uu+/3pJUY47Rmln3Faq2959vAIe7ZS9h4ArIwlVYab+Ph9y+rGrRLOgCQQ+M9ZwC2oDbev7FuEU0
1CvD/Az4+btZmBcg2S5ghedt1JJJ8CVfEnucV2QFIe5acymfe54w4jlDFFswdPU6R4zXzZ4Acy5v
1s8EBPyuJQsaZfCeqkmjvefxT3H7KeN0Ao7gMXvskIbxLPjvfkEqX9+r3SeHi2CT/1ArWt1gUwEi
15utMhN9DU3dupKmgnEBr8nSyUgCZqopjROHyx0dsXMDaS1ChXVLfhA7xtJcpXyODAF6EESL66mg
BjbEs3BAp5nc3dI++02PwxLmeAq81cKZ2aymX3e50J0Zdxz5QCQeZScKshraHh3LowaZ4oCIqhcu
SquE3Pl5iBWehFYQTDao4ZgWSYrmlziNwrIVzAT054OwZXZ61hycIC4YKRanUozKWHPfP+0SYpXu
ZJOcrmqoRfHYquwBg13ocDlln4QKkxpbypuJyBYgOPJVwo5S0ZwHBBwHzELVflEtOTHOPSoKiZYk
BaY62hn01Q/xuBT03M5zWTltCf4hlwRGEKv9dyJvwi8LhhBrAPE31Nhrd5ls+Rl+o0eQPQg3cmhq
1fCjtBTzRw+DjwgViO3OmMM8qEJUdn9lxUMH3Fmq6PNE/rVFsD9MNVegxJU05fK2dyCJ6EIKNdJI
q5RS8qVPkhdvjGuuzqvNBGOhGlGp0dzjbKCofh6W5HHe1cTZBAB+bb90pAVWhu8bVV+f5gLHOuCl
FFsOceOgS5U8EKgSsNn18cds0WL0XS2H4XVp2XJTedeEwDl1pyVsTCaLEDSqWaHDEWhPGtteOL0/
+YKpcyj5mt+R+dOi4OUPc7scFOvuW4Nj58q+9+ZBO6OBVBTZx5V9WFHwhTPCQ2wAZwr23HIuS6vg
3rIayrap5VXido2zlM+X7MoCWquRSaO6X7i3nsKif4Udz6RNwlenZYjtEJurh35G9THkYKs50RLa
okVIQh88pc5/Kh+OAgSRgtz7L1eJyDxKUb2rOTHvhADM+9y2y5igpzKCDnJ73Ijl2S3cHVwJ9rQr
L+ZrXjUJ8RQpawb0Nt7UDiUuP2o3pFnwc8vLcWDMHMirJzw0rjkQVaicuRErgxr4HCw1bpN24KeO
7J6VugBaPUkoPvaEojG8+RB4/Z5X052JVprLjCnu4UZMzehR3GeiJBuy0YVgYM4DHOcIabcvgwh4
ILu7hYtlC7AE2nxnQ1HnLdo8BwL5Bj5BPMFV/Navqf949xIizB9SiL8vDLRa28nNGAhv/2L7C79T
7CVBLsqT7d8q1PNQbDxFbJY+XzUfm0s6wFGGue0z80cIOusAsCBLOx7AylxauKjR95iWstYAoevm
cpyLe7mwf2T+3dWZEUrKRvVjG5LleV+/Ni83C/JgzEkIZcJ+ukxg0yMEV5JfH2HjpKfauFaVXiKu
jdiokNeYsb0jUfX1GgcZFBPHueH54TvV3VOdh6s41DBU/cwmIRuul51+IIzJNV8230vBZBWuAtOq
6wOChCSfp0ZY8HOW5BIOcVWFMFmjT7jXEVCjwpRzaGxqYI4QDkBPGf6sy19gwptDNVi06B4zm/pw
qpuzfXigvIoLaDdY2KCEVUIvRWILj4xBUWyiGNq/514SxXhvl07675uRsxgzDu3XKCn0Whz7FhQ+
Pqqk4gPfZhZJ/YSd9J2GWIBZQnfKBHwOvkKNdQ5oBdgbJo4fMDANXGsrciCeYDMSQizebbYntk+O
MlsQqLEPENdcQ6rcM7/eXttQr3jEmIk6Qqe/8RLbJYOqI/l4bhkk0nhnr+UhZV2J0yWa37CY+qX3
Gj/SuXuRZFQ8OoPAkqX9Gy/Ln9kRDpjp5QWJgcDdsSjkW0Su6ygdd408x7o4CtmtKzSGNFHDf51M
6RcV3PHRbyPK+r7qrs5u+2wam0Y8dg1mPiCeCkJlJ5FSVCD7vHDCCeNBiABaemQ//kRW/ztkfC4W
F5Oz2JhQsbgnLC3oHRCSdUiAMTID81y/yet77Wyuo+tlkJ6f9jKn8Cn1dLgiFDgvwud9C4ahWhWh
Xa7/acxn6wHOOB8LRAwVIFEHc4J1Lne6pzgkXU05J4Xxqeygh3zQdgD+B8MiPpmLtSJ6xRuICLuG
R6ERENZEud6RMwLrnzYD4Iov2/zh5gDnHqfsJ6z3NtWYL5H2sf6ZeyhirxHutRg/1tH0HZeeEV54
9q9zdQrlisnRT4xvU/s+G3SA7M68poVezZ9NXFyengtz9xFWs0rJ90U1OxjYMc+mJ9Hg5kkILVuI
fsj0mfUOj9ZSbzHH3rHpmolb3M9MmfzdU7hasf2cZCrcFSgF9f/6v+VNTYn7xYkBwcXdZXQuLNoL
a3kv7RD9PAip18J1yS/GVJtXZfrtijapAL4EzTnb83K3dzPB+gKE/Q19NMkfHWW18/N9J+UKpemy
F0WgRp0YtUs+3hWx4LBDtZWyKfcTxk7wahkaXLbxR8OnTit2suxglY/fWjVmNZfATE0gqeByhHo4
gx9Eoyj9enCBDn0aBvWwsX7tIPQCMCSPTNwpBlt8ctRUuBg0ZVPTYt6b0iWEZKAunTcTVD49s60n
G8FFI/lCf6ax0Nba6EdtRiYpqBj/UCMMWAOqop3j0caIB9aWwAfZZPuC0GST2sCiUGWVvlWdfJUT
mCk2yQXLUN6l7YbgS34dAOIlGqZyHgqz1RXrZs8rpcKM4bsqa85TdcBORnldDX4jlEsnlzw402VW
i0KJ/JEj7uP8VEsC7ON7c6f8pwS/zDrGC66eXFOpzYh1OIwjc7qxhvqiyXRxVRXAiF9tzBcZQFU4
ETUnFbeQ4TFDodmETDUM8d/LLoxitzOhSjwrvlw1hUsZrovB52l6iGVttjoDBWygLZkiEIVyBeOD
v3XiVj5jH26LlLIZHNlLwVJm3UWD38Kipw/8qhpsnJXE32ZUBKlqqJ3iLGLqY9e9RaD4urjTTkqP
IpHBHYggldhjUxwnaRG+y51xZDgNBsKm4Du8KqM4relSL2aIixQKQ15NRSF28eDHnE/ZbBoc0xPO
Z3ZPVVxkDtVGpJEUHN85/W3jEtXUWReGZ6C3ZFfpyDXlnQlevZrOlJ/wxls60fbZ/HCqjAVz5sPf
mxfi0sw8kPPr1MAX6+6suvhD87qD1EgRwwQ0zZh1szKKwrJ3F7+1opTjeidrd6wM4xQQ6npqCcwX
9JouJ/Pa6z8wzchygu10ioX4jTDG+F8Jtf3+otAkzlJmTdh0BLGjJy19XpA98EmIYxavQqMkIBKr
ZA6CYSI85KUu+P7Fr94L10hZCMqzStmvdudv/douSlbqotuPWBsbgEHXREedNrVARJg6PF2UJDvz
PkM57kuhTvXpfKcAHerVHcAQ/PJgRRRftlMZ4j5VCAPkLF2oNZTOZFky8HyqxNEH0xCuLOORmM8r
ZfxANBE3BmniEVDI/hxVCsINwOhcUudXC6Rv0ijIuGCdcKKmU7+G6Dmkx+fOBeB3p9KEcI+HJkn3
Yi6Su0kMO+WmWCYeTCxQIF6utIhwDiIIWjOBisn4OtceYKHZuPnhhqaeTKp4Dh3ObJiouikeAAXD
6Po0fMphoGWZ5yR/FamCk9ptcI9uMuhTc8SdJa4rpzQtzJuHh09F5bqQST3I7jQmQX3UGaua3pu/
bd/VzGmEUiOBRr5UWsIyl2TP7f8OudKZuigFtvwTskAjUYAx+lEJYU0iCBF6wcuAXzCe43l3T+RU
RAJGNP2U8jzW0O6ZxbUzQNSdosEi9gH/eSDt+qbcIH4bqR51Z0dZ+NrA8oo78YHIINUSrVAL4Rvr
5ZQtpkp+ehE6RM1++2u1iXbgvSQCO/qGrY1MToWay1tN0Bwu5bBjsDyrGfiRQZtf7qTCeG+Q3o4L
gYDB0O6mlLP6wisB++Ol0fBOsMcQtYEY/YdmFnCz2ySBTnxIXYGyNdxY0Q42LMiQrJyx13UrbfkG
0I5dOhS7paBszsrgnzmWeheG8AC0ZBcHyosRXIt9FKLxRHEBZqseFNQPfh4BQu4T1tpFjN0nXVie
w+bIUVGy1KQlPcOYZFIQCAiRZbS7u/ggTI4Usjf4giiFc7hEljlNCNS17nwz+/j9lleqeWVOmrzE
mayB9ITB7fKc/iAKumHFUJ65zHitbnQaA8+2mbuM3G9wLTViicURqEaxgjxD4hn6qoz+BXQhJssL
yaKeOMqKJXrXYMhmWxUmHqb51kNOTCew2shwFPhTPDkKJF13ZRO2zvfTzS2ij+kf0wUJkNqw4dIR
ZSo1fS0PeiIT6sHL9uG/RVtMgO7ErQ7YzY0S8A+6lZ6v0XYKEWKyW5+ylSi0ms0M3JP4c/luVfZ/
38nycz9Mamg5W44jVF8YWBvuEJD6r2BrzObaecBH+gMu2xCcyJlXrWIGFJA/jXboTKy5Z3kykHTJ
KCGME5bQwmzcV6UqAr4pv04D05ZCWWTyIrbsiigTnWvyuQGGhpWrc/XvP0s6ihYsGhlGVBlMvXPs
khheqhEm9qNnDomnrFv2PbJMZEIRmZTqOKOXA3x2XKJlVejMgBElXbyWpHD3hTL8foc9G7ncZZ/G
2vcfCvRtr7IyCSTt2FAR0fMikJT6uz3BiA68ZvJaur8rQiO67DgTgoZSJpLcZICjj1tJa1R1rlgg
qK1eAS2rpQ6xm7FBaalU8mdSceVYiNbHSlGSKKjGrKlXAnbo6YV65OwLDNr5Q8HjsdVZbbwLFbWE
gu8d4+q9wJ9Ktw4WR9dM/sJ7qATi23sbUd0hn1ljur980Z5imbgre0Fnra3bbgac/vxBMDPfykh5
ws7gVdJBQ4aZzRAvFJ5oRcvqeTexdi3sUrrBcQxEp/HRHRRRcSLE/YtOjUQltf5F6xK230jbjfa3
8IcYz9+jqjSTRGoIaJVksi+XbZHPNBoOBuYjb4rt0Q7pPeUqxEHKpwS72uimAbBac02EApzPnKjT
Gh3LycINWBoG0LaFQqzMFCOuYoE39ZcIcj5sjty199eAnYECMyzfwhxiqNNDf16Opl0a+ityYwQU
uY7JuWqUXokltBx3PDnTZm6Mp8ga7AKpPt8EELrJyCAJ+CnCYu8b7Mju59hGm38AxdGNl42RPlhS
ex7EsqvlGXVKl7/NxxCZoPWPqp+rr4C+tiCOXPmo0GxIcvd8IfQgu3LmptXI9Q+0NX6zHZR4buyG
Q7Ng1scQqTqPR37gn9/K6vVQecm3Zc8t30bS2lg44XldiKuAxSB6wFUE8DvoqCL4ohxNYD6LMzqK
7xgadJzPHbv/5+cBOhyxJ/lUluLAGSzGNiFN0Vs8NgwpLvCFg6F7CHBq7l4TxtWYj26Bxvj45ylV
rTraRlfk4nyUvU/ASm/f0zH5QWLGJJIg9KVWYTx3vKTZdm8DSDuGImDLlY0EZbcNjjEklnqHRFv1
koFwHYu7taNBLBlqZtCyJLhitzDhmXU+m82oyH3bf+VsqhZXThKFqtrvpcqXgTKotXQNP8I62JmC
duo54OeRvk40KKsEKH3wS4QGGG5L2xuZXRWAa4HEPNvQW+ErG6q0l7tAFI+EIuLe/rj3+HkIe9Xq
p2Jq4adjVzNzrEh5wIbrbZ0lxzJrf93wIfQgWOVH2XNFlS6RwR9qKh54XgzhTEW7irrH3BbjbScd
sPUm+rM5gCnTrb7krG9ZP30fBhedtRXHXCSACQrOivE61WuCE00EZsmL7m410zv+LdXpf9s8JSIr
j8nb7JGirBq+0YUUC9Kc52nXrIdjzvl0jfzyxhZpzz3wCwOcU8PHeVz+txHQrENlaPVeNDd8IRGn
A5kxWX28QIE8cC+MRRyNES5DDJj9VEB+pTUkZBdsoLHCN/sS+vCjFqO+vYnrWbwSg+z82ePEHjWc
ol9bECM59iXzbvWZ9MlcVFU/OBoI3Qs4XgokiUCamByvIkLlFq4oTOelzIwi7StAuscS3ydG+sVB
bhNwsxTlA4jejYOQbvVQODINCvmBA5v3NR6Au5G34j2ipoEmlfTRXgVNdgOQAUzBVyy0vGptZtY7
BdkvEYpR4jlLQhmUcKwRXmbHnCn+gQRoG5Uy0B+QjAERStrz+8W+RqZ64+rVZO+LPmMsg1nBhH8a
pi6AudVfrrgtQP2gTEar1nQf8L4yRmLZCHRGurVJW7OC/ZAeZXmfqVFKZJ4kgsZ9d7UanR/7hnxS
jF2rVGPnfazLGOlJgdpm4G89b8T1/DlzjUxbAEs3bYzjFyGgv1k5sEgKIfU0+jT8QvFl8h906HPf
cI33r/mTlEpuiQU7WJdNti0mYQmiucKoeQPZtCHQMSKr4lOl3DZrm1maJbqmle2KDLlXYDabdrXQ
fzrUSnLwCmHat3g0RQvXXWxfA7C3FazVlQJUa640pGoWgp/y060ALHnUsLk8R+CvOxfjd7UuP+fH
Wfdf9MtM52WN3rIuVb1O8eWtRTKevdISewtu69gjDOnpD29HFJqGN3Ar6bsdrdX6p/VLhILM2hrw
bAPeWErlQeOXed4Ni/kC31yOC8r5jYxtGo9opYJeH0RK902E0B1ITT1j+Uzyz8WIS6pra4pM9PUX
0+CcH+3GivmZNo5pNRFS0WjX4zqwsbN2awvoz6CrTJVWTiClrrTX/3Un8VRbuaFXz9JSLl5gYMTG
Rms+YF6SRyq8c9+sbws7Gp5iQ1yCW+LCXuPMYg8m/mhxHLDZHugmptoJCXgQckxqz8U8+Fp6Fplr
vlgZINFQT/AGpQRVTlCFrTu+WBWp44L8TRCLDRa8xYd1s3+lWtPbPeCK8m3ghvkcQy1jtQuSmEmk
YXSmpNk1ZBCaJ5rY3rtKpTHU2iyY8F5zGG7nBYuIMODGL1IcGM+Bud01GZXNDWVY4OuiDOcCa8hY
DMjRaKliDUfQ8jnH1b6Smfw9Y8ZVX3+6p/LrnmsZRsolJiqaXDPnlQbJz62ZNthQUFZqOHRCXTZV
7wiOHofb9pRDDBQCVGTnAVuPvoulweDtI5byiRLduNuk+wy9d+mIM0pKJz0dP8G96V25HyFUYu+Q
N0CB/nZfpzuQiCztwnKdStBL7uNiUurmRt/mi5GtT2uE97hFTzWqROFse0jgUml8Zs0edINwJYg5
xQ4JVl5Ry/wDmhu3sKCj3/TWTHOGvfONTHI8NbfJr0TM+yb9v3sugEGtQ8y2c+9Bc7DaL7geK5TA
v6eUA0OBKzMXM6F1jzQG6EAcpVX1vReP4m7+oFTNGHzCY9WDLUwwoLol8wiefcCWmkcQsFLcGZ0V
xBAH0fx1GoBM9LQozbZBXs45qJo+MNjaBbtjxUNf7YxGpfldlw93SIeF2krlAsoV+YWWd3Wccb96
kWbU1H1MuoM7rfZxi3kslRyOL5Q++bdIOOVqheQkOn3/PtRh6N7OgBN9hgnm2g+aBrNkomftDC+0
hW4jWipA8PvvBk27KJU8Eyz/wCsOSGRdG76rGjg+bzoWPOQj4Kjqlvyna6mCdtUsPV5nxVkPtGOx
Ckz4mi1AaInwXLV4HZFHDUClaplc085ruKy8s3qQI3Yv5ZNU4KzzCffLt1s3a531K/SnNKgD8Wba
9Tud1ieJ+3LKN8q2y07zsn9bpIsuA6oep2eMCszVW3XfYiAMdd3Cjakh8wD5qhLPfEnjRikpqVO9
bHUHnvmHymKKdSLcirA6K5dW239Kll1qKsbMmewvI5mYwNKDjhKh+nFjkYvkOvM/zg9QJ6fgK/LB
SBUUgIMrzYiD4fVPlbIh99DLRtCP+u79hR9YbblKv9ZwyVkyqDEbhgJfeuDt2EWTY7Ce9FHOvR+g
FNrr01j70w0yffxZWnolR5VC9xCczswkAdDiFwTfeM1atFhuER6LFN2qZTS/GeK/KpBZVgRJp87O
FsAekcr2C5VKW628rAH1Ie2EJTWTxivR+XMiJkrkKVA6VBSfepnCIINkJsdQpcl0Fo3qq4HuxgxX
74jZfJJ2b3Bg5fbsaHsc2arpA+W+2G4NUwb+wqQRUWN7Y0B/dFfKUR67uY+CtiaqEFIUGyqw/hat
gWF/AtcI5FD/NM3YdXhMaRuAAOjUFrhogu7PhViorRO523HrGFSJcml81N5DRPmQHWHrn5s4EDjS
776ZxCppfGAN1XHoKnEZcQNLN+WMlZ/g1jTFa8tod09tAlIfMfvPH8LmCboLZ9VkBpjFAwLM654A
ExDugV+NuAK1WPAyZ3sSWUtjRLXy8mE6A+HgWeppTVJUfVDmoLMhvnMoHSBCmt0Bg+xIbgm1rI+Y
ZNxHtmNlbgUJmNErXd7DWmHAJxhDFNSUAe1aOwkGCLVUDR1WIw6TiXxk2htz20cNLaMwpK4rmQ9N
MeZNdtHDjMUEB/TyYRdIpFjQ7dW5fFdS5wU5muqnjWzDg/SqHwxc8nzNrq8a5cZGMu9mJ/HbIm1k
/8HAIQaOFe7tOG9v5C+Qg8fO4e4jH2zHTfTksK1U/R/DqMqpsnq8s1Q2LJc/CUYfJzsjMp8eso2b
MCTpxAbp9X5AVjtCH0V8Lfdvgw7ZJh+oumzEyRE2zi83Qh0xu0PxdSDv+RzoFfV51A5JL9JcZ+if
aCYQBEtOJa4RkkEaw8nikRXwDsHCelWq/P5wf5gcZzbnHjuM1BeM3RtOgTgD3a9SWBv4Tz/wUDwl
lIDE2+8SrXzuv9FDdCPvDKbuaOwmYhCNub2egXqnSTlMbVGYX3+W5vvotgSTLiQPWMKlA11zi6SF
sacJ+lqUSnAM0J+KX6F+dg91gDAxD5cHRLjc9854lSGqVoSPNlHoGJyrpEzmqp6alVX0yLO7GTc5
+ox9XuKP+zrZNdB6gYvXjpK82/WcwO1rBJy0479Nqdq7tFcSOeastlh2ABSPNKDr/uOYX/RdEC4f
b80EnEhk8Rsbxqt6YXmNPL/viCmWSOOcGbvs7sfLVZqUbwv8lCYZn2da4gOOJ4bRmcowl1Lo+Hds
c1ie1iQ7bbDRMmxA3DQx7W0p1nd9aBu54xfaA4KdKHJvqBfFp8gcl9jqLjWkhz5ci2fvVfhrG5Ft
+VLqFKdsWk8CUW9LBZcQpRiKlEBopp8d5kegjZQiRImgNiPF77xpRlBWuQMQLGYc/LmH1CDRiUCN
wGSG43TAUmfEdSbt5pnbNytajq38NbC+1JzqsQ+MzJhmJUfJAtdJXa4o2qCxaEJjJFCA3m15bQDv
Ys7rX8C8Mw2eol5rT0LYZuZQkAJF4zpC6nVpZ1LRi/0dOgRJg4cnG8V+A67lESLDOiulXUtzuhqj
S0eyL4S6fj7vMbqvGjlUFj3388bc85qygcPLXlfa8lveZrR2H5gvoPrqkvjEsLUZaQQI/jTdBgyg
3sjgAk8lu6zkZWRAWOD2CRq1FEC+uwAvt1NDUEXM0QBBDco4Uiu/qmd+yL9BgRy1P8DvJ7O1BD6F
dspp1jWEEvWneQPyxuJp2V6ufeV8ezOfrwYwzJq0ho1xzwwR2p7PQU0zzTMNQj4A8PIa15AJcfgU
wJX8kyuodG3YbRFEPnRIPLoGkGTV7iIUrGTSIcs/ibX8GV9JtmDQ+CivGi7czhWZRIMjJ1MBJ6kc
JgfW4ji3u/Y0GnH1s83OJyhvex5V2DR3IPxpJxWW3lt9+UjuXUtUbnZJZqk9pS9zoZqz0eLBAy6k
Lx1lFS425Fbvqbr7ellsDzE+9/yleWuzDFgaeV7JwHwYCI0PzIkSAOR83T9VZfiIYdvuT86EJmeJ
w4htBnFbG7qElBAYVsI9pxMiIp7uCJCTg6xPcDDyDpPXtM2AylSFEwbcBmRYVfjorhoM9xDsurqh
J+maNW3fgww9pGCwHFb+Bu69AUHbOJ1IbESK9hiyScBfIkYgyWpZlUXV41LrBdKlIRY0egdn303W
kxRYExbol17ObM6KDvoAJEP+nmNXPVqjgEemcaX+JHvifcP6/m+3+EAx2rhoYkN7rFS8nVuiMEfI
SHNOJ1wxnHoFab/bF8IsENUVb8EknIhBcxFdYXS4vG/qvzRvRV+H+Chs7rVSyEZZxkpOhAzPa3vQ
rgaieSmE7JbUIuwMptBqNC+oIEnEi8MyR/PTW90OmTuF/Idy9jkQ09S3+A93NTHqxk2UgL9PT+VL
P7gBHQ9vP4UrSeowrUvNWSKTcf7CunJIQgWphYW8hRtK98GuO3nsGbOZuDrRe4aegfSwNZwOYg2/
uNq+fSDwyBp6ZFj4uenKwyDyxAhwi7+XnycMP0JhOxF4+btK/F4uusDwwimjS5CWQBD6Ui1+CxDS
K9VdjNM1b+FtxWpnXnyHBb290Ucc32zqcRkd3dTZqt++V5uegPnJyZso7Q+CezvJxobGH1gYPNm3
ificEyVsEGZLlbeplv11ne9aP66XuECBJlNgNQZYBeUsMd5Pd1xXstmHKx8X1nP/lu0+QWtg018a
jpi1Oi3uLTGaXkx/26V1qLRN87nlzzeWrbTaRdWZOe9dsL+lQvx8PX+g5GhGwUNpGJoq7DoV1YFj
NtjNC+sZxPqOOnHLjty4scPZNTQ/TZySn4US0H7PoSs5lqaXqtiO2y9LZVTr72M3W07BkU/dNmgl
qesvRwzOMSUjqancXEc8N5y53yJs+3xbylsLH/NsbswlQ21D4dsOMglVSPGZHYQ2wixyHLE6aMH7
yVUTQDIUdNUDFsmnpIThI9uOV1yeHVtIhCTUzOX/VR1ILdJ1/i5vVT3cLu5FUKS1R9jy7IHSx4Y3
Rz2Qo3Dk2/D+jZ7baItMwT0YZOQ+tAtuZZOQVZyuG5pk3uYRFtqcsN3aWzBHW+svhtcEQnOPjShU
kHAs/WxK9GnMAbvG3+h9wXLuoIt2ZiydEd4hbQktK5JSqpRGjVzMfrBUP2t4Nu00def8MS1xTb/t
WA/X7WiRCjaABasAo9vcfW/qxk/Cz43Qw4jZzE49JZky2/4bdAHaSJCeZsQiKJZEHyQKNNQsYxJ0
aPOKMANY0byibGhMWx0+G60EXKL+kP4vm4mfGFBfy5WaAjaMZXL84AMjOux9ldtT99Go/Z+nnTOr
l2wZIaZBa9GXZ+Krkus/EMFHlzlIr//lqqj9iA0bn/111604bdpOhKk922jkEnEtukrAXhPkS91O
65nGQxuJgKSV1WlqyjJZsm0wzhGdAcccrLg3Ridn0F4jw/0OIEaPl3Ge0yLB1AthiAJYL6cqlfKv
DKh+s9kyw8cJq+jcN8HigrXfqQ13x5ch3I7RjmUxmREKX0dVe52B2JwpP27af8oJZR1pXF1KHiQA
uTaKTcggnrD8IoRLpPj1ZqafM5hRZU2zvtJ2E7gP8o55twVxAATIDHkIhGEj/6YnZXVVbtTfXfVE
H+CIBTTokUbiiHCZThlL4GSjqPzQzhc1xae1wPd6HmfIa21WFDdnQY92NLv1WChnIoqXVjIOloOP
fLnAvnMiexnqJqKz6fKtz/177f/D7EpbwFk9/aZFJcnt7LoF/awnOV5I6oP1nslnsLPBDPItJDt6
9iZya2UL0u/eMxxAI4q6GL7R/jpjVvb1LHAU0JE/vKLc+1dUsLjmhi+ftTjH+NWSfQvj+sW8Nh5S
Gjztklywu1MpoMoKALOkmkMRNEvVoUzq0JxR1oikibOTnvzXsER/vgFjOSDMhxIjJ/txe1mvZi8t
1rswbKj/or4Q/xB5BadEoc9AQ3qOLTUfveYaI9M4qYN2Z+o3Ozn3Roe/0UOJecIXECmXM6ie0RPF
nFl0W3nA/PYkTRvAm+QCLZ35wB3/KmrJVtjIo1fzejAWeWQDPvc6i2eA5mKaoO2yxV3rQnbMzpFA
2RsWVgYLUJSRfojzO5tzAZxwKOASmu/O+7T862U4jeBbHxpM3D4Ek+czoG44tWPGQ87Ul2yMbZLl
rNBO+at99awRpDB3VsAtLg2WN0Pk53oPr4jrapn4pSZD8CpNrcJ96OyfqWhsp3yYhA6O6kmzoItI
RKHjvnyfSlLzn8RKuh2VyG864LCPSW9WzVjFjbWKIA4tHIY0RLXDuuJnOZ7nJh/Mev91DfOXh9fg
sNd9/8rxS428mOy/JYdhU4jf13fhcGQVCbdADuYmFjzva+tJb231A2Cq2u7fWIpU+UHkdZ4LIjJ/
lRarcK4X4bZ33hI5tvehq1/yJHD1JJJf9XqVBh4s7lZzh2OlvROAIDA7Hwqn280v9NcjESLSnvm0
bbfHkN55ocByWEMF35bo/t6AwFGLIn18CoOAeRoSHp4mNEZ70HGQHXEK+ShrFvyoPkSMnQ5ipTuy
ch4qlonXOLKPzVNgy6TH5S1eMiYofcH8LGrNw2q57A33sHzjUuGeAGiIim83D7t2RMsPK3ZfqeB5
xF+iPWuJKLYdcDk00pwRRWPkseJINFZ3FPmw4yIRpK+Beg/kSPxYgU55lnZ0XoW+L6XbDFpKPZSI
06JjEo+QWjV4HKriZqtT16MLItqsgQXey0rRcKj/MVq1VeWN559Lc1iurImXTBRB0QwDY2F2s36F
SRNlgy8R3LzE2YdV3Ps4qTkv0ZKqfMTGSAmVMTXhGKm0AbUmQmDcZHSwMeKhYOnlDg4xzRbdsXJO
48GDhT+X8GI3I8Z7CyXbM4Smf6oYMWJiw+uezZxLaLrpYjnkndFQ/NFoLWXcINVgDSpb9S142iKC
uqi786BwbaZt4/mnUbLVFzW0eKvq/Nj/pLKADsdokgZ44gUj+XN9kI3aabfsloFk48yACfKQClsa
5vuEcaV2yqBozZSIjhKUCNdvlGvfAwQRYMQWeK+8A47fafOQkLeHm4llkYkDmfm+TiKfvbGfD8Wt
FAsvdE63cl19uezZIdN9Lcx5pM3Bho9/SO/L3LRbzlKjWaokpqMXdo+sIpysDI3XYJhUEuMHH1LR
/1kyzyL9xhm5cTbvriYEDnbpPes0ScyNdqP2zEP4X15MC54USEPn1hZE+JQrQWZsU2aNjSkPWKTS
HMa4nvUni6nMu+qKkunZlfoFSnp2Vx6IzNdE/DIdR1Gjdvu/YffSXcx3ljwkHG8SBmRbB2ml6655
7fe17RFT8WC6gORTVUwvT9YYSBauC4n6/XjcJAEuwiAVfNoIDSVpGIull6rT0UV+pMwy24X8wmrG
pIpSvblbN5U2JKEK+QEuviXOOHtixAAPtdDtquHZq0aFmb69xBmPDXQMwfksdUVjJMfZECW5l9xL
I3x2AQNu4O2QnZY7wdWx0SdkIh1nx7Gwfpx6j2ytfKieLC0fUS8oLRm68QUBftxM5AZQUY7jLKkU
tKeD10Rklb+WYJGJkpDZmNHGbXllHg8fBud40s+Ok1oSoqTN2QhTgb74n9ZKMj8se5iuZAE4C26P
4TDpDhtJnV62oZNI0Dvc9HHmHJkZU0zQ9XmGh+PZXKUHejSrFVfUDKmFhAoz9Xi8goFXXcpzO59P
oebA4lurEddxsY/RBQy2H4BrbHIyNS1rtW2FYHAJCn2RukFUmXV7+jl9ZBWB+OpH2DbNhQf93wPJ
eBeJ9SVHeRUBih0HO7J1MnxpTV2LobaSfZMPArzXoI0bKku9WfWtHnkgAAwxz41tY+7142WXsuNN
WAtgW2Dmkhoas7+Lt+l2rEtDxiEZIgaZNqsDUsleF9m/j7JgXzQq0bR0rTePLHvxWxrtHam9t10/
l3U6GPZq0Z6zCn5CcFCluM+JOmEJCAKrbBtzb823zEfdMenki3CQk3Da68AvKMZPtK77HBHTTa16
MJS84PKsZyEI366UGOlOw80lWtudKHrV1A8azCaSG9FKUN/WJwojtgd65YJ7buN6HhJVlQShd4Ns
mETIKrvF9TNXbaIaSJKZfqlg1i1nkc7Y4jWSCT9vu6uep+86w5Ls/1xk+3a+Wf8/GfKUwd9NKsqU
vSZdPN5BUg5FbKMkTsskzVTnIUOT5zXrnqOLqKxGhTXuDVUdrZKKN9FUGiWQ/RAOMcHymjcAqBDj
6ShK9I3/WY2Ih9ymMThDNhgfoVf3TsCrYYMskgtu8q8ZUxpmllf1J31DSHjMIV1p7+0qV38zBK6N
h35Bvyu272TSiQ8oO33stgvlBIZOt/Inz6ElQgj6C6oHH1nJoCN24+7EM7DtOzAiL7V4PMOdvsTw
feu56I1Ru2y36InyCZyceXLK2xq1kgRt7I+0nJINXpKx69Rhcev/NAe/kmhW2qLa6zgVFT95CGqe
9oUuGiQRgFJnrbiC+cdKNI/h8vW/uF3/P5nUmka5lFS/eDC1chl7gXcKN1o5pyqHv6eLBmRJbHL9
FZaoffgj07FrSeQJNb3r0JnPY8oAus0hm055aPfVpDj3l6hBur5xTbxF9BzZWggPDqYqwMgrkBLa
/cAp//Vnq+NGwwd+HyJnm6a6iNxW8YwTWRSQdO5isfiirVFB/09uoAjnmQN4O/6h9noeBpyLFb3u
BLvbW6L6IrwLMV+7mphae7cn9SDFjqx/6vwWLCJbpiMYacxU+MynT4Hv1tKDD7MJL0Bti6l/i+sT
qE/KsLteE48LUzyqMRRkxoiOuiWqU2rzf03r2U+cyiJCQ25MPrMULIIfjQcUMQcu/WtDqQadH8C4
d7gTrcXrjst5H7W/d6jpbPQS8tI8cnBQFdKO4ISuO5TnbclHufO097ebkrTPogIqGuVczE4oESqc
rPuLSql69nBqompe+hTpAojfVlOI3eSPBn3sEx4CZe3XhkgJHnpNiV9vC3AYeIKPYykh+t+5p9KW
/ywwMYjn6yw+CACz06iEQW6XdEBizYI6RKX+joCwCdH2o9DRZ3CsBgGtf6m3fjWFjNBCpOuELWks
JMLpraCLzo9YpVYJ+NGrllUZm2npCVvH8Ffx89+eZw0OMwEYag7bNj8VJnBkKfRnz5dmof947+9s
K8qRtSingaLExgkaihiGpbAs2T7GdKcczOaQfOLFQqmveFbnrxb0ygXuaQGZwKN984CpkLkTLuNc
bC7qjbeUk1J+bQGfYbnD2RdNzQDjcNc91AUjOGVZJXz82E9ZsQRGPHm2w0V2zhKBK6SHM4RlpJgx
LwAUUfSfJsHa5aa3UUvqaxnYJQa2510hlu/yKAqkjBID2jYNz6ssbFha5+5hcbxCmaTl/eH9BJ3X
8+n/9FYJZyjSoJ02heewdSkccBMBs1bkJ8BbQIIk43RvsW7Kw/5Z/4g223WDMZYJj5wXYpBlmPjD
eKPZ4HFm7zlmkYKITDyZpz8AfGYF0L5L5ExMH8gjMHmj7aS+59gnecvaJJ2Az5w5fwcR64muTvO/
cSxUFOxtSc8TB4glvXDV01Paq+uF79UZ8x3+/g3fqLv/qyVLkdek0NceeygsvEwWygPyCMkPDQaH
k6RspLCxX3oxFI/a5lI0FZVJKG3z/RrPJi8eRSOczZY88VZF0iVmwywxrQMMaHZtNy8SlsCHc/wt
epESThh/9Rs8yA/TiRAamdqeMvgA0xuJBzIDLeF/B5QxH+NI7ETMK4F/2E6AjOeanxBNC1VmshpN
NWvw2BdNqXojl7DSzHmJ9N/8d9Ri/HpDLvqwmdelWjSG3sl+I+wg1drGgqccFOCZuDeLJIYHCt9h
3gODBq7cpAY8b4m4rhMCovW/slqSnGXWgzoVUIxdTleEpM55DGyd2TT/sce/xUNJ9V80Z0jHVAD3
sK2HBbdOaJvtghUn/8biue3NpAS9AYsIxxCawZ1PGPMN6SXoUFA1fM15khFB+nMAAGUilaV/XTA0
ePwPls8Kt3hICvuq8Vs8+A+PCEJ873WEeIH+1A14X+fbyWLjieR8FB05vSdLS568DRyCzNFpOatq
Xld7WFLCYaM398LjtvjQjf/9RBDIoBMjXOALoS2q9w1CLNPVQCcF6HGQeqM9K26keHTI4oe/cJzW
XUUet55mIzIUAfovsVZeobGcys5it/xAo4eDkVTZEQCrp3o1A73aWuar5u3QbQbelc07gUrQyzPD
z8lJArEmN8CwcldbbCKCfD2PCEogAZpp5cv+YXzVkRj6Y69eMvaLPK7xb6hJWVvLylKOLO7m9S5i
aMQzFY9ClQLntg1pbsVKUVL9Nk6FmlBao6olH+dt9yeUnngzsMiLyUcPvlNvUQNFn/x1Zk3kEIjz
Iv3Xklr7Jet0l50waEibBq+a8NtZZze/Dm/ouNAx1B+8dvELFet8DHBet8i30Z5GqGu00w9y29hE
PXBBkvdpja4Tg01x/i91W5Ikzv82xtJvpSNFpEvfLHEEncHuChfRDJgfhKVLa5U8s3UF8e0JIMYG
JAj/pYWSdl1f0Zj8LPPcrpqz0LS2XGY/t6BqeP4IB0OjhQwvNv2sXCXimu/c7lk2tn+j7qNvq/p0
E3eI2enYgA+gztrzdQXEooCKEdpN9ZagSytlAOLmkKgZKG6ORO+OeS6kMjxVanKuOHSfGCNpLtBN
BmtQ8yMRmUh73ssS3ozmrKJcRuTMd+Sr+VK4lh7AeJ/KV3rzina95fmpVqVwJX/6hiEFGlHnfh0k
UG8ersLCDBWx/fm6Q6kOlRo/J/MpstEfb2BtL6BNLOXvFOlNR1lW863d02ysOo4XYLAjYdC61UkV
VftxoXiIekOSfL5YUBLcklFJo/H8ex97jW+Sm9dEF6XYj+3Zxu3yx20J0iqYyVJgVCgwiSGcA9K7
J2xadko3688oT9gjfTeToFdCoNTwqG/qjyDpgk03AdjBc5C95P01lXaoqwvikJTyBTTw46P+xy3v
mblHwpuFG9FrZWY9vhwJqWwLf82Rgy6YtJv6XEg58FQ+QcgwvBraTgVCN7EjTRg4cILokFKPJZhQ
jf0C20dqr9PjV0MivCqCmt/qhQOwBTWG+sXMqDL8s3NEg+aRh17sMVzf34w9hsHwlIYnWfr8fUSf
raKFHvly44C1jZyGsIqOZoFnqLM7K6Ydr8e0FScUdBz9/WVtAwaQFHQl8LYY6DmBRM22JsCjU8Vi
h6VZ8tvZNoLqpfVvxdsGKCeeMKuPBoh90glhY/2vwlkzz6OIyvUyiHrgorON7pvztwMSBh5z7zVc
D/q159e9qdhSkoioBLjtbLpvVD5eYRdDUWgSJ58Tm/MhrRddMI+33DfbTgnNHElxEN4TMfSjlEix
4etVFh75BZ8PwzREEKNIefanPyYclzFu3ouX6Nv5j5VtamEErqXv6RYB2grDzTl9F2gb4KGybuox
yo7vv2Z16QlViYu0xoBCGSp8eJYyI/xi61zFXJLH1AOhkF65j2szU+P2jj4F7CY7r1GR6oMH0Lca
zacU/JmFS1c18URvzzG1g3n/hJheXpwIVG6y02hk97Js5n5q6PL1Jk6KyNZafJC5GI31M3RbrKtA
PH47t1dnF0RFvfb2QWffExk9WmoE2aKOfPemAwJjx4GMYrLyDAP3G0cWWeEg1Du0mNtGFwdwrHLi
IO1I6JnekRA/YAP9v8nRTmU4VT+QPwaLqJvCl3er3Gq9i67Yyuo2YsUKzVDcLBqkyTp2k/odt2tW
XdurHijWeHK9sYGOkPMzxieIoG9kceQb64aIjpEKeIl3kba9Xn9Ne9pH4CdkB3EiuxV9o9o5oTz6
6MeAYGIJmsOgHJTiKgJpL1K/+WiwWgp818a1HANmR9uLWjgEFz0YCnEBFJcylqxHUkuuZVzE7rw+
Kv1F//N9nnYgceEWwA4M8RwTg8100zMg8VXjTtAjYXl7kc0MTer2jJLQSgeFdoI4zib6dBt1YDU6
hHaN05aP9RrMFWobDqr1Hocrp2lMOyrUlJuhRWsT0IedpeDLvQL4+VzbTiMtjk0dyfElFenQofSb
yFoy5dpzm6otx4UuEsUEAs5PcwH7td2Cqsy2BiQK4us0DnXUdY+v84I7wqzNrlxmQ0kfAbw32cOY
22CsWGWTkuWVpeIU5YVk5J06/nvNJjVyvQ3YYXt50D9A7jjaeDsuNZ3ZqdbRA+vHkpQEJyaXfEjp
xIsI9zSLZUIflVJc4dvMSNmcLnopWjqdpMqZVmM/I9yvdLeHjzWbPMEu/TxLNfxzwwasJSPSjn3M
rkadZPBiPeZOXLrw4Mfs0ivZ+P8LnIDyhZlCaf/CypgWrQcch4YwekColxoB3FMlai3CNe1f9No7
8JMRky1hGBIJlT+Wmzv8/noYRExYqDzwl4klyMu1+dA95LvDpEGbN9mclGzNeLB90qZxKEdVpF6R
JC8b9bIKuutHaKu/lIUAZHscKD/UJpxPLcYABnHuXS8tZYrqsSWjiEFpN6aWrysE5wA0GK6oJSUq
3gwqQ+uSp2fv/PicbnqzZi6PnUjNWj9BrEH1XbD6l2ratDlQ8mV5M0D3ockO4Q/7YInW5J1wsMxi
wJInDHLVJ8Rz5hz0ZwLgawMrZefPuoakG/BbOMghPgpA5DQvDgsV+LdcsF4wRA0Fs0S5ZjFAJRKk
RgFlby1Bq7lwbKP84+qJ2tBjIv0Zqz34crbGR5ldWaKhXtheRXII9+RI4YpHYUAkXlddSPujDgVI
7ClDBeehdohtaZ2tyZkw9cnJlZMzMwDJfn5vJlW4jP/MoDOhXHxF5mKoJ3022Svnf9G+uAHmaw1s
4Q8g3fn9cmdVEzekzE+zFs/P8XZMVoG7y44MxPpB5iSS6cOSHD3EE3Qa3pVI81cahBaoUhs9XqP4
5EqI/QgO/IDJQak1DHnuBm1UOnoxGUxsyke5k0MamuoIbMHZ5I3llgzo/0CKk+WpHKO+he/RQNMN
quDAqbBugdvQbt1kL8WGbqGN7yi0rM3TWL+IhjCpFs01xj7+7PItQjAgKI/vtdBaWgi2yt1Obrsc
hPV6o1t1Q1WKdSl1JQ/wWHTGtcPG3Vq+C4j8kbjnZtHOiZzhrFpdm6tU6BI0/qbtg48Vsu0zyA3i
huSRHsx3oJXFcMmnoZoxo8QePdghXISasSxiRyhDNOi+YmUOCcLJsKcYvfJaJwiRFufiyZIMQk9J
Z+J6jBlVcVF7OqE1QK8bsMlQDK+Idh9xMvxxMEQxtjpElOhLoV9wN9KkBQpTL6lrTYH5jfF+ojy7
F5as2XQ4ewCWMroAxJmfKFvTuUPH3RdVxkhmRu7TU/4qHdCoeacsSEmleedXHdrqFo9BuIbTl4s5
C6aNe9RTrfZ7qup5ADOgDOU6dAc/0nE1BqKjrCFGFOLNrxpZiqkUJBDHmpnMLKd7UWesYeJHe0m7
gyU5bJpSnE6h5TJmHZRoTsMH9Y/w96Mcu+lrtAs+vcauUSXWBTi6cDUJpHN7EyH9CukVhd9CW5Nd
lz1mjfkQJw8MMfjvIOUmlzALDNFxG1mYrMtcC+GCYDI4Tjn/2FtddQk/beA5YfA96V6mSnQOvJV/
gpBMUJ3RNrIyw/ceDsPSju5DapE+nY6Hh1wiK3xfvoUTGC2k+oeYeyFbJ++NY71yOQXNe8Zcqn8T
jFeixxS8nvPu0bLrHngRYfJ3e3RfH/PamkdWnp4Y6SJT7Wujo9iyrsoG03nnCbR86WrEDFErHIHP
ffBL6h/beOI/C/wO2rdB9ZJayPFpGfRQn00lW3VXpWwdvrz5ViVp0fJOYbZH3C5LUrwIKe8J4EDd
DhxgCeo/OP4/DOdtc9WK64lU2IkvoSI1DJophSyKwi52Ng0Fqr5OM+g2u0EHYv/zcEn+gK0Jq7WW
Bse0uYtLvQXbF5WnDPSuJfXbUJ+tLmsnibTIxZ0XwadWWuMk7yhbk8k/mKJpQMuiskdvK1AahgkC
8n95gCJjdm+uL0JiFiS9c40djWslvVjKaNzsRr53imv9CaebHH0/0DErwTUkSJjSoyub8r+oggP3
KsHnkQ1vvXU+G/JOXjrahyyCSGFG8N28v9r9Gi/LaTO25qJFLG4FlokIjwI9XIQOSl5rAeC9n+5T
1q0D3b6ztpkOmtpy2768xyioZWMGdHj/4Dm81RIYx+rqot+Sg6L76PXdgXsJwf+2tlE+wsSeHHi5
ASZicNV5XL8jX+zmSCkRYFaG7hPcR75npRL6AMSiDIup416jbCij5OX88bjhYbnKxTYjpTQfvrad
CQUIaphmhK+lsZHKVSq6Axg71v6LacHAks117hqtoztojSkZOP3U2g9u2NYyGcfqOzlibL0x1erq
+C+1QnVXbn53MFYWNBkbfm6XTOUSMSpRba/OyxbOiTxSyyhlh/vO0zmxVieuPzYgo50CNW2sWtWP
g1cVUBJbL/YoRDaQFbRTDTSHfLwKXT1iDCUIYgCdn3JEHSDwaj5J4rExdTThRayChsS4hBLAf8eT
OYC7Jof5MPDh4VoxM/n0Lw0xqY5Et+Mcw2hmlaNBpTRQyNx7qFVnKDvyKeLs9yl6/fW5vO37Fjmh
v4MQTcxO9sfBIz4TWawdJAlK8eiwCZNBigIWYKmRxC44KQXXAjRRMXG5mqPYR+p7J8VU0a1GhdZL
jEb2ML0NQQh7jR1UP98ZeWZKAqiKV061qYxKK7yJQlLLbs9mw6JCCTNK8jTAFeShxowzg+5gmD2v
tfsIsXlwIGqFHr7JuhbrcLV0nHtxID0w5WEci0fovX5Evkg1QOoYRtqOkrgRrtXi6LNwGtIBHCzT
vVtCqZ46E0Ydn1z4SS5tS2zFrwiSS3muStnlvOOHFSapTtd8B/acukkatpTq3Bh0mV9YVym2DxEW
i5lOd8C6QMMphpltxh0wI1uqmGCJXS5DFjuq0kirRH4nAc6hTg4FcEd6qU2TGT0nhPQoVNforTQA
2yD1IGsy9BnBadXpNGUnBtzIYwNtcVikKpXvOZ8qGqV//2l1nh7Q9jAp1yV223f8t00/23emzOAD
XyMuXiyxoMi+xyYeKDNB20dUr5ezeOHhXBgb1F7q9Ko9JBIDq57KE4Avpx/3qt/2o3b0Q4bV/hTl
FCMQs7SmC0k+P7m01uzT0ZpEPDnMOehccNOkhMTGlv2p0/1dXO/L5Zq8iTn/YHt75lZ4IA1HakJR
n9jbDUBcuYjMEiUQnkv6IiKLuNjvHpLAHOQl59uPi1eseyE2L8dKyKXxXzhP5x4+qK6widFqqh+g
kjlHqfQ+pMtgOpy7vUFRaadByWOpkEC92RIawwR6Ut1phD3fOxJBgImbRLAArs5MioC3RG6u2uR5
6Nrc4Ffda6+slMDEZOh3tLVY/trccUOWq2n3lCdFT/a+9PXt5WDWEk9N6wJ+m87yB0xhNDfW0YGI
+MBBOSzHT2staOH/OCFfx3Ci71a4zFomtM9gKw3jwCwEEdrsfcOmmOw3npbLM0FiqYRCkY7LLIOV
QWuubsI3Wl8dxQFQo1JFAyuRXe2yH3Yk+SQ0n4Dnu84W+Oo+x7/Z/JZhlFkBpy2y3JQ+A+RrxMoV
H2/CF6swXfJpm8Q/NzvpD9iPxkjZEsPSx72B59azU+afScvej6KObSOLQzjFpvicpnPwORWKqhDP
MbuqcJS/XMIebuuTeby64aV2mRHtr9UM/SPeQ+/x592NuLn/ttdrQX6fg23rf+19/pPIuQP0eu7l
4OfxQebzEoswjcVXfBxPIyDyDkiOFMHa/OIl6ljuCri2UHQcijm+DyHi6rr1e7rT9sY+LC/EaauL
+Yy8y0uS+BURB3Iz49xVMFriIjrSHbx5KkZePnFH+FwJGdqLZyxqoZpL1lt5LHESEuTa1Fnd6/Di
DI77wBuKDAN5Kp4aIPL6Ql1KibI40FMIW9SuYXMs6eCpZLp1z96g1fEP1PFVH5uqoIvXhLvLWNxB
sistNJ1N5H63ysYDhX593RWnmdqxFvV0snaVo+k73uMFXw6oXGJrc6dsZBEkiHuREvWGWC0geybO
xpv7aCNjG6rfmX7W2Ixiid8YGEVC1kVbzGBvdhf2yJjUEvdoBcLWwgRLEaTIu5QkscZuk6A5MGM6
7QLhRIkISQC5K0KyI62xyNlGLzMkcA/gkRH1sNWb8N6RxGMYEbR4e+mrQwlt6eTFeDIknBeiMpmQ
2g640xdKBT4y62VhNQTNvJU0LIWQQ/4SpzV2TBCUX4RKQtO8KrMD5pkcZ/Alsx9oV93QynaatbOx
zDrvHvsJfoftD+XRFPtRdFLLvMQbP1qAWVjBygGBwlDLPmJtl1k2x8FjB/CkOmZfwVrZemp8elKB
rFszNdMbfbwihyZjz67mW2q5son3IKPMoD/78J6Ds3BfRck6g/Llo3PW4YICRT5i2W6TKQEfoSJe
J8GOjNmrsNb6gBd1kbOSDsDP3u9jAT8CasISNG0/FujS4bqaOsTEnDU4gt0oH/q9gVyVXyQCnCa7
K+OdrgLwXOTKodJTykrSqGnJd6OzQtf2X9RjvzHO4jxXl2gUUlit69vrxV15yX9cmsCjvPhMkLtp
Wfodk5Gv/V7l35o06Vt7dgGTZnowvQLk7hcPaIy0Ua0BHX7GQu94zauYdnvkPDX+FBDfLWslyPLG
eJXhLk0paLX7nsryHBwHugZ8tyQyLRGMmwU+QH1PQkiiEN66NzGd2a+gJ3eARh0a36QN4RQYjrkF
C/BZNEGJpLWO17udv1vO7bFDB6ttzzUANcBKNNW9pqm0SD5h/1knQQygph/X5pBC2/mRGn0o1+bY
S0kZxH98THJbvnZCoNjN7LuloUB/yy/Q7AP34W9//NEmGPeN8gCWPoT/z5ElJKNFUF+NhOUYvRsX
+7pAvchpl0MC3WyWhwh7e/9PcMGhOL0UXqD1brgezZpZ9sxsj7Xcb4MUf895pdXXUpkcIAsWWimc
0mb9QgsjhhY0yT1c6gaZ7GTBeuO2wc+viKjNHC902ggKMKYgTvJNzeKa1DgwvUybieXKk5aCyf2a
oPWDdjKmE8FJJAbVldNiX82f2frwjRJq9eG6FloTybXnsE4m3H4EEtq+PT3ml4GI1fr1ZhQqx6TZ
D8Lgr++p4Q4G8wSGIOmA/EJrUszITVO4JSHEIv9k+hmSeJkccgWNVD3Znt3Ko+sy0+ynUqqWDnOD
5f4AR1eVqo60LRyDYC05dsLutlOtTzsRL6b6SOT0l8A9LW4C49Trhu1EuY4yL1lHCOM/3oT8nmwB
RWKI7LnVC9z455qDI6rHurUlKcwARNMi/TD+4rGATu8vfq27+CqC35jmbU3sKOY9csY1DBy4q+HJ
SwkkFPIILSG9egqb+YYV/xq3YJPUrcSvl4/4ISz/k+tGqhQANh1BX2FwyvUsZvmMymIyMRHm/Xe4
eJHcYFAmJuBDXrDNcEvQt50mi7Zinf35RVQNLUmFR13svjGPmjauAS2suoT5fEWpNmVWyWyik9Xo
+BcsLt+8Dr7BWC0qcO+q8T+4Uc339lMl9jWcq9xby6bIIms4SOrkWKadrnPAt6u6izt+Tu8h5ZoA
rKZChlv8UzAZ/9xtMM5ptT71iwllVWL725CNqFHxcDkeTy0bvHQHKKxkgrsD0ZyREUIn7ijizcLm
qzvg7JHZ4Nryzi6jI7AqG50Bv8rKU9VLecEDq6QDweTEdNp+VMmqhhuu0Vx3jB49L5pNr383Lbcj
6FD6jIJ3OES0QlQR5/DG9u3lz36FmTQzh0HOojCRYcTc7yQBi2PeP2FBbbV+Fh6QCuSnn3prSZt6
D3WCr6Yn98Pe23qK62RLRvhXxxeBO44IjgblOAGTOlWLH/MpDZr1vUvQZs6knp1TYPXySNNmLjgm
tfvPLH275pheEEvW626KkNx4Br26UlTWNaY/sefX/lQxre21R1JVRNJ1JZ5j0k+g8i+tbB2XuvQl
94Sg4ed3L0dYKYmevUWfyQNqEMY5yb+hCu/YRM8zSqdfK7b3otYhw1GCiOrMLmc9TfOh6Z91DafL
gvlYJttYFdIT5cw6mGgeFOwZLW7BOhUnQtyvhY0/S2rjd8F2saVbXxI/raFkxfzRlMKLTso/FjFz
qp/2KkR96YINWx/UZfm3DWt+bvmhOGax5wXyrEQFlurZ0wZ0jTAtitgGCrnsWXw9JcmYoVP3DPJ9
S/0PVUJAw2945+o3ZkqcB0M6Dq1VhYOlnvpvi71lYjI9gPy5yQHBoCPXfKZZEK/O2PrM6VoVt3IJ
8va+rABQwZe/slBv+c2ZnXY59USGaYP1RvwXiwSWq0LWgGQmzbNYH/17jb1Dxq1f4Dfa8zUEk6dB
3u0evP7JNu8cruhCd+WNRQmhFq8V93Lth3aHg+wrO8wapfeKkt+2CeVFZPTcM1y9Vb+nVfClht1T
buO5ABoaFs7KW+bWNmF12W1C95iq1rf0l0G/HpRun7Q0OlmfQTecmwN7Ea+rKVeIfxhVAW1Bia2n
r3z9e9T/3NgHGFaHCN/H4w7zKRekggG+GgSSTNAXKmKE+90g69iMncKYbluRdo2mFwb9lCKLTpAg
oeYUnbR8huUV7M4BALI6BFbFA4d45xfdlpOw/iJiyYm04iNsM5aLQUuahwHiEZ/ZNUBkDojIR8LV
wxJqS0wV4FBkcddPxCqLpR64ztthLJwFUn2DR4KLOtXC/K6Niy1l3SzI9H37WkgY31n4e7O8tiqy
EDlKa7N+DLeh+PmH/G6jsS3gyb9TbVqbFhb3HWdjodfS3n6qZ+NoEMjCdpRI+Nu3liCn24oiKGsv
M6Sv5KV2ylI0XD2OmWUVm+V6743r5FovRhvFV3z34+kd1TrkjScpN4WVQxyNjF1PiRufhy5bzSCv
FnZMHBNgpg4Ax5AU1clxSVYDd3ZKar14QPCG32HK79Xqbn3rZTreg5vXRpTgYH/a/eULckFRMXre
nIg3nu4cOvGzgAQfQzkqOeAYqPiGQmG6+/zdYqZbgszeSH3QNsxZLS9MgwotY0Yc0P6O2GgPZjoE
eMvV9J9+Vsp1yhbZvSCWdtDCDWQhwCH5dncbyZqi4tAnMty0Gmth/IaCYDxmq0Q17d4z3TZVhTLd
O5GaxdFeHpVOdXPxSgfZ90OhU2uJ5t0GaK5CIc/ZZsZzySSBlv6JrbsY1P+t34XpFu48T7D1X3NN
uvixJLn2NCzTXFQUWfddgU3yaAPBQpk23oryDxsuvm8tAy0i49z8rHzI2Gc4dTpYfWb4t/IQUPJu
9jJoE4+bphiGXb3CLCxgJkMhJHTetHQKmqlymlttLsioPt5ZgeygxBjl2Yx12eWdpDBnskSXdBAe
YPOyXG8pjOr/YGpH7FrN4XUMarptrnezp0DU0NPccsk0yV9N1yUWEgDSQ+pHIgk57lqvbRjqfsQG
KDafGjc/YrBYSiMdkpT0zfiR9dhg51EeVp6tcYqnbBVDrTko1Harpsn07IZYAkjvb/U5Tkl4ZlXI
9QRXT/SgRd/P+JGhldeCcikYV9D9C20wTGxvUiOzgG8gnBfNNCwFgHJMDjEXFTIDg5QHkfVbXxfE
3o3Q+oB7XndNiMNPcV5GJGwKKTJMYZ+S/ILlOD/1mi84qAbxGDk2LdI7q/yjpIcIAyaRqrCy2l/j
ilyz6+hriNCh7HMTv1xeg+lDH0GKsAGO0voiZqoUHlMGyWbVBa3oH7ib3z9WoVs0v7kFYRMWyIle
GqluPUN80f1K0gQeOU8B3Rc381ZsHPwrsLeq2G5cbx7s6fgqpao6rTDiRDp34DGiQWl5Ax/CBYZ8
0Xx4NXwqzuV++4XJvcdmpUg9o8NF0kTEF6zr29JoNfi/dDw3v+cOHa0hSKEoX+oQnzkYhRC5/qA8
iX8yCx3s98yeXRq1MgG6y26WlJ53spJO5s3b4NGi+yRfGOjkwhFcrAzpLunvxtcP9z4Fc3HtmMtB
nLIzve1N9eC7LP7n7Y1aZ0FGGNIw+VpNrebkhSA0J9gbBNNwSEbJ7cofbwCHrjRrbrc9pc0QrkMU
Y9TsTeQXr/xgrfrKKwgYm77jBjVHMuplYDp0bnMw0ga6y9gEHRZEZxXMT0UG5x++UN+7XUrgTZLe
8M8y0LU9oB83lIhWNezLpwPMb0aQKQU5pRgitOdh+XCl4DPljbgay61AW7lGWLgtdndew7KEMu0i
O/2vhK+ygPZbhQ25xJ3jvKbiciRWhjlhx1DJqV06ct0zFT06Semvmt1u/jL9rmyXQ3YG96iVbkz1
NBA0j80/UoLrUceBvXIMPpBtytU7khGlxN2+W9MuIZEteQqjguVhqa+dm7GYZx7alhHvZ7BWjYsO
+8ay5E3hYZn3qvFZLGMY2TJ9c9pdWTJimGd/cWyjEexgApopsKZm5d58tpexNM8KvoegCFS4fPdO
K3+XZpfzl5aijtS3j7rOLaclG+tchfs6vrSffIZx3CyPwbr65qpIvXBl7CtWkebSwoBfZ/q9Rsd6
u/KdacE+khnqD12On369Qu+HKdg4gyvG90gxEL4BDWLXCPKwcPYRXfgLgFaE4OYujQpMF+jT1ovH
SVMWFpllnDYVsKJVoMudDx+LE/Wn3guFfofnyTqXy82sVvSJbmJRklyhiWRSp1IFn37wDICzrxkm
bg4sRUxarJFcEcEJY3iX2P4TYjgxLdXC5GKxBzc8GyTPSGU3vmm5M++7tVOR1jU8KVqTRAw2/lW5
iFggDrLvcpr3g73+Hr3RsPB5gWK4Ihq8jau8Sc/dMyhN9x9Cmou1w99/hlSnrnEUGJ1sFc/gN7Rk
0BQPxhCkrosmcpHME4OP7RmWOzJn3WEvQMa9A34ZgefWK28FxzdWIUjT03UPpJRhEstTe/y68lif
Wj5ipsHU2oPXAVAofPAu6pOy3IrtvsmjmN3xnXceqFruaJz/GUXG3KoQsPCnEwn0qeukk34eDzmU
pfYs40MYGZFVyh+WAynNfYSrAOplueC09/PINo1/h8G8iQg1aS8dQdOihf0U9qmoKpGKCjmQCf39
l2XUYUEBKjo7zQZJqR3QTOur+x8k3mUJTZ9Q1mml+f9N2grMONq3EDMze+0tBdWS/ItZpRrl2lpN
QGakvxJ5e+46z94JoTnMtH+4DzRgCRrBI+69pxNWbMpncfs1erqGLL9TYm0Z1O1Z+HKxHQLd/YGg
yzxPA2fvqP2agnjeKgTpyo3syCpuQSdcakLaREQE6joAsoC8KiD/G/YMxDuQAzBJhn3Q5HVhaOKS
+W44iYmC+lcVIWB9RJi7Iw9/cmcqhVRO1c9934jwAH3Q/lhHKeO+0u2y232CfG2+EB4OLNKfWF/h
FRcxEMzY77uL8E84JmeItIM5k7Nx4dJKoB1e16zzGJswYaETbWmbgM32f9x8HecDqE3MeJHYlERA
rGgVV2cq2iSj+JAz+5dMXj3ZOnfGDV9S4PUILX3K6IsRdOn1xOyNfHCHHQidVd+meUqe0ttPusHG
N73NjRJ0yp9EGw5dAJ+0f/KzE+dDwzh8lhgoNt9/Y69wuVPiyP7UKshvJiSbmmiUF9duEb0KmRv4
ql/bV3AX4R2Uai6ZX6oXaoUelVqAymOiyttHFbWGGSW/wel2Pc1La9L9F9OO1I9a3PZwSH0dF3ux
099/+XhTrbLggo04POUzdw9iiwomgj8JgwnKlX1pdDLZTgQpUQvoTz1CoJnJ3Ot+bmNTNnnrtVq8
q1fV6nLI4/5xw4p6wx9ugBOt992+Bg9ZmF5t3fFCkO91Nt0CI0o6F6q3VG+XI5eykLDC+7+QWjFh
iUi/A+y1ksfyClqZSAz3HoKWfbdU9PteMLyfghfZAfRvPWtlYDp2o/gB89F3NCxWoDvA1eWw0TFq
gC5m2d2TX850taaX4La8p+j2aRj49h1vxUInJu4vOC+qkjZ2RUFWfkzxS7DwxLTsdv4RlVN6aokh
T5O7YgdTreAhnBD1YqP7SCEg0ajHwloBGJ7St5+O7+1Thch7iZdWP67rP75xQCXi+2jxhF/Rwdep
BO8OdnUsO+MN18drgYmGIeV4Zar4hcRBR3I709zcu7+BXsLsP3H01nHCU4Hg1XgC7tpNQTaeKx1b
fRU7HtdGqu6Nm/OMFwkaQNy8nxIQXNAB5twA0PGqL2s2gMeHXowCjRxz6w7K3GryLMUFUbZGF/gO
9tQErjw6tyBHD3QOFe8RgiwD1zlwwvltv6HxLGHQts0GJhhCyErBGGLrgP9/kyQ7kDd9/ND9ZGAR
nnXuLmekYolSUtU2o7g7rXVVM5ewCdmp7HpYXFTy3XkxDZQotaRmiKPp/YCNRym+CptwRB2Yf39Q
9kLKDmZTwVnffLuJAIUXgPiWE+pqKA3zRQl60kf7pZM/t7+ulRCOmp1CJ4tnUUYQlz5VHSI0WN13
RAMP4Ql5zzwZIQjum69oSVF7ah2UNMmEOfvAt7yJc9v22H5DlXQmAVU6sY/L7lzmzZhArBAuD2Cx
p+eiqfQrsURkOPE3P0zI9Ht6kRicOj7uvCiC9Ly7MKp6YnZctBUzXaSY7a55S3Pfm1jswmlffdMZ
oJ8Nq+EcDFfvUrN8CCLMi7jN++2h1SWyqxsTCPPNB1Z5FqitjPF8y35dEj4Py/IR5cnbHEyHEp0V
5Qe27FC4vr0oU1v1sgt+SKhvKb8nsrKWOJLZ2jar2h4bUM7JhQ9NLKWsMjdjetDy4X3L3QrfHFdu
mwFIfpKGtKmEhhZRGgNkgCWb46Bk60XA/SerI9lkvdKAzb77YR6U/xSZA3SPM35ZtXnDxJOpeU/g
+ytKdRyus4O+fYMVBqZfjXVELEsccIEGhOmHNNxQ6qjxlGDHICFEVDqrUkJ+jQRvd1j73q5Px3Iz
vuH3Ha5TrSTNaF4qcCEuQh/kFjI1Q59NxWwTjvCKcZP72BDmwYenyY6AYtFmS4T/itHHJBOqTu5Y
dX/QCjX/E3ZejSb+ATnSL78GxxF2X0IEFB7u6qgAz12CYXIIkFv3w5po2lgtSvlA2fVe3WE+1nJm
gB5u/SsVRxofl+THNI32vPxqFLkY0/bw0QzlwzNrYdZZHB4NTd6Y33yhoYXhUn6rA8iLCFmy8P7Y
Kd6hON+HYAB/zJ7/N4Jo9BvUjgcxEKDzciJVHL8c5jldqf38e2DvQnuK9Og8KpBw5IiFxrD4ExpF
z4gqk+q9bCEJGirDChefCk3yPDheYd1UjXnrN7OsOM1Wxf1RaewfGiKIEoTBBKoOTfgySJfqwDzx
qJEeICI6l45z13qmBEvD8a60He0z3UIVSpnLRSGpRe+lFsr3AE/2r0FHGp/JCDLZFmA173IruKRJ
5vdATYotJ1Uqsqyo4XjdVBiIMpjAKyt+3YUDkp/2ox6O3GgEBlzP6wSLV2zypXpZOCslBA7TIBpx
TfGBXAXY+aT6dJa4NwLIx/LFjeZK4pgR4NOQ+FwCQIjE5j1TULoTPpWMKmzPaTn6VYJMdJ+uaRrX
nJNvRh/HFJppibQ3Ys0YD4ECit/nRwmtVgzBj1ljji6pxfzAmxAvrFcL1Kqv74vkxEz/UuSbpLZi
oCDjXqx/qwh78+XDd2Rg8PmKwfE+D9PZxzWvbcNrTmEGdifNMslPYXu1cOlzNjzPvQGbQbqMm8fm
bG+GXoUCnX1z4XXLGooeIHZFmkaPQ7o4EyFqnoQrTXOWtbzSy4uhtludK1tJWbcoKt1qo4BnIPGz
dFnMTu9Ri75grpNrR/CUaqqLmJn+0cSzucf4rlvolqAo+MXOMy1uVxLvJ7+zzlYhhdaeNObAOlXR
QGb3/fk3nPoE5Dfwpd4lI/ypEKWrIuE4fe0cvOpBk4Xmm1131S2tQvL3RU2Om2zgrSbncCFXntZj
nkQqONEXm1zxQmRgKDCClT4mq9mOz/XtIoQ+LCmg/4Bt0F3uA0Ah7mQfdXpAKnviJe89uMGu8ZBz
1uyNWsCok866uhHv12ADUU4rqQIkF90ExfIaDFpIWgZA0rJh/ORwtuIpx+4i+8ssdMoAiY8oDGtT
Yn9O7Jfsx7o5zT4M8fFc/IiNH+tnfBpTgSLCdnMOHg+RowXSHAuMsP8OQ13AEio5WlDggbW727Cj
RkjjSdB+QaKMKbgVLuahWc/gJ/8b5j4orIDNxU9p3g8QKYWc7yTKwBb47TJGhkykfWlzQqLJ3E0L
dubMy/xUOCmWBgrUeWmnZDHrly2TcR5E6Mz+bNV+wI/9KDchNzz/X7HLl9kkv+QfUAWk/Pa2GxVK
8faQCoAEeXIFybgXNeiBTiVvWWwoFRyiHtG7E5C6Qfx0A7Fu6fOzkDbMZm41i51HLNpt+pE1kfQ6
L4gDa5gI23n7/ufCEXMWD+OfBBYjFfCTZ2Te1xTCd+JJVT9ODM6H1m3KIN6l+2BjWqdDi1jifvSg
NR4apMM85w4IgqqrbimTHrPJYS1djNwRv5JU4XbruyfmlStDXUD/ETHM1H5RWyrKbe2EqT5i9Igh
YNu6xLGziFAi+fn0iFuTF5Yajlj9gKJRE7bbMpAB6Yqf2MVW7+EiBmViox6nFSOuaOWoEoC/2HaE
NDB7sM7+DfaB6u/ZEEhPXKjly28oHmSQXaKqBmpbkXDHR2KGylAo2Dh394FSd2r0p35gvYIY1A79
PCURrIEE678gg7hs7YnK+LtqBzIJh4VdP2pbxHXiwOsyTfn++ELPYRyIP2g6RJls9tjOsbXTg+iG
nxql7Y3CLx7dpQrg8+nm5UohhHZJT3WSK1O5d0qQK+eaAxshlbMzlhW+A+KTntQCxER2pJC7FnRD
gMkEDTGe154UF3YMiYGZH9bhbYuiM7usmgxdjzCbDkYtzQ1bpteC+AUiQQ6ehAkVZHajBoXNLOM9
gCd35+5LYOFkJzd+YV1WyLzT2QPkibLb9Cr75PBE/w74J+OA91q3j2p6yTUbdnEcqSBx2JA5o4mB
3ACADxBftbwHyeKWEhaz+wtaYItXU6dwEaLXico1aTghiWE2UUV0I75Ns0UgW9HxmADLAzs9hQzr
JYwhWZ1rODFOv8MyPCt76+zIZBZYmVkXDnv3ZTKHGIFAwVqwb2IwWBxQ9bMU7gBz2sOtGh5O/pDL
6g3EEGIOMlgL8C9AtKyV1tufoPisM34OsscN1ALIvCatoOUIKlQ8UfzzG2OiGY6Cmy5KbZgPCfON
8eSB74VkcOlk/SvaT6+tT/sCQTMxv9bBHHlWzypGn6TfPqaCdUoHp4z7MBYigyvRnUG2kWXzUhF6
/oJoeNp3FVq0mnnZuXfTP0O8e0SyfacANq+VmrM87F4pohjY4SD8BsRub3qyZE7g5uBMbPXIaJ2M
D+h+NA44z/0T2XZkfY53wSuFLxJQ2GqE8Q9qby29u/iQ4+XwP6XMg0gjTUBUerD6HpaF6zWLUr0K
QNX9FEgPWpalBY3cYdm7x2/lNb27Mt6FgdQYJIh7eDc/OUuZze+5SQtTzuoHlXCVv0LZQpMEqj3p
dJj39hbaXw/+3cU/kpRTXpAaYpwDESTD3+t+xokTuzVUcJmZSBujq4S17UJvCuLNexM038sgQQQW
su5vL+/C5iF+udau8n9HjnFpxHuLVoKHF1EWsH2IQUJUmcNJLPpR2EcMrMBJD5WJ6KMG77EXhUo8
4TMxPlz3/lH04Fk80z3JvvihtDTHlPxR/Z21y8XJIyV0sQiYLAI5OtgnqOvxD04T52/pD3nv0IEG
YzyVwLwWr5qLucHeytu5ilJRnTir1j/Oyftv5AtDK++VKw7gQ+xIvMK+BGpjW+9iQSvIq20hniez
P33DaYOaK59u81A9lIcm2DjqlAUpY4yMKHK0FLKZmNq5mYYlDCP/y+EVGdQQmp1F9fq0HY72v279
a5B9VuQqHYNXCOnT/h2uFYTCkShcaPgFG2sqeAHINptOOC0hbtTlkP02Y1eAik2YSQnvnyTndKZo
ZQArILTRTq/VEWDrCbrQES4HFY6BcQ1gRtnoH6qH1wJIcKhzi2w7Ya1EY3zHBsKrBo+dI7emn7O2
IrCKUtNEjrHmB6jUL7ThhvSgcEbd+qlqzvrGbxaQCZSxeMWIriKMXRSHVdAr7wcN/ZoiagfUW86k
A86x0cPvmZyejsbjPTNKWUtXJbYh+COHr9uBhdU5riSp1STdMhiwVsLruwVTJAiX77lk0v5qJw4i
m23x3Ag+/dzjoetyATpAkq1IOVI3R6pSlqlbfAqqYsukcP9p7MLHiZtaJkzMzn34EdxMk/w6Javp
ZFji5O0WSd2ZXSMuLcx+m5R1ubetVEtxSxmryQL2whPt/mWY9fQ4qky5pLh+ZV08WUuVwzaEhrlA
fr6V1qbnRb8qm37xUC4jAOpOHDEPlAugx389j8IBSKrxpfcxKOBUwihAicgGeL2wg+SbYC1LAwgG
SBtdzHwuuvo5QKIhJx9go0eljOM/9MraQiwC7pgt/gvCyn6D7vSJMeBecdgX2BvO/HGwniLM1FI3
337KT7FQO3MP1PPs6UHWG/CYD1OYFXWdkUxKQNArdVc7tsFNwgS9ZjebjOJQICptYCS2drEd18t4
OdGjGgPtF1lckX5FzDmfKyQonDofSuXSINn+2Kj/l+YY2Nh9akmWzy22SSlpk07Cen8fiGUgmmBS
VB+8w9v73R6dpcbJKyguLpqcjCpfjgOcf78NVMwyV7lzXdnqmaGpugljFNMlbV7Lb+2Cq9ePLrXE
EdmwzE7DYRLYjEHsoxaTrwd+SzF8QUh/xm6nRGlqoJl/4wm3SFbBxK+hsvsqFC5VKpl9qJs1xCeB
oPMywpxJ7IFfehNsqYkBrj1ka6m0Uw6qmNe7ksLZp9sH8lMiR8aSB1XiPz8uO3OwXIOBRK4NFJqS
eZPmW3oZytCB/fI2/XRh0BZmWQLg3/FMfJtjenY7g1tFHdi9BLwXSHBjhONkbsdI+SwPvKk9Bagb
ILZM9EPKlhervZYnSddUA6XguOFopT8g7ZJFi8QA3oLFV5MO5fwbWZgZrbcN/BlyaSN+Uq7Ss3Yu
uH3zube6kfPzCJHByfvbyf0SfV/TUKkV1U+UwQCsXtfDXwA2tDVVDYXD2RnG66RJmzNigB8OQz85
8zeTSPo1q3UQsaNm6yoHUhc2W+gxGjD5iM9XBiMfk89Y1OyqlpYEhzEX2RzQcS2FE++ty0UraxIV
m+LXiPuD0ThGNFHKkulkgMDy+8/SI9HFWx2n0y7voPSrmp/jX/FC7W7Je/jM93VNQfvlVOTfUH6v
mXyLHhcylCCUlODQXrG3YHmv21ngVZ1a6ObE6znZ4B1192xKYNKTu8BfaCJYsWTWeijBO+pXr9RJ
hfz0IyyZjkM5NXFvBE3OUeYAk0RkAavCCQbOAwt7kpCwHqc6C2Ci0Uhy4UQ1IbOoPGrDc8A4clhZ
6cPQUYYzqyl96yxBOnJe8Jk3dyd/s4d60T70DMijqgtyOrDgXGAuH6L6dY+w7MCDO+9DPON3dntb
iissnC0KfVaAE69ByWW+GOsaK7KpesiWBxyiZBT06R7Spsna6ewRYADgR0IVhDX3YjpKK4ylbWsM
DLhNfl+FcJDATLlGjW+N3Cff2D5QURhjVv1NPZg54X5xER5oyv5Shp2GwDAofxWqZCBRT8WdMd4c
E8ZmTWdwPMR1z51JTj+vKJoX54MGBhrMjm3dxCXEH6161nT0e49BquJQuHz3bY8xh/ea7qVe3vrw
cLicKvk806YJ/iAMn0Z0uz62gDPaeNcxqZc0nHv0yGGXwNPK+7fYWJPVvo2V13KNGSs1Wl0NGMsy
kW0Nkikai3D9XKJhtSIEkhjFc7cSmOW8PN+lxQDk0PSF7UhhhLmw5mzzaPwtei4K4ASRMvtvIJeo
5tO1N5n0wkBrgh/zP6P67cV3MuHNladYVO43WTcNsuU+OPUMXV3Hh8Sn3CPOVhqnNonSBWbVqkJ1
TKRCgZOFtCmbqeXaE6sfWf1kt9Q+QglvkMpL+hlal5O4SdNSPKrJ1YzNXdh7FdBGaoPmslPAlGQp
MtDMmMLVsZUMyFgfUXxoDQNUPTVAHYh9W2As5/506+OJb+ShodnyQpV0EOZUzNN8dveawQT73ACf
1EklWMhTAAwTOA4UPPRBh0elJ5WKNV3gfrTAgw+3IeDHZxBTNB+yfjzbdX53Y3x76bRF8d7qcot2
+GhsCOREyDB8E/+bOpxNMKoVOe2XH0Wlq2YOStEmuD78FOGX6JkEGnb75yLmqN2cdgwaN5SVzIwt
YhMjAxziqNlqg6zLZfJ1TTNkf6gHG59VzFV6DJkyCtxQOfFc6r0GKaW8kkXllHuxrEq0DcPlQXLO
wD0z1MdLaE436RbZ7NhsmcvfpnSVfiUExLQBInfvYQNMf+CiJuMiBZtYC+e0WVEq+oo27bsFssf4
NF80AfAUIkrTzXsxIb7uiip6POd7iqfhCWIQcOa9fL4Q6SONsL+9/qawdDlWNa+8qLx7qRToIXzH
A6OteeATLB3pi7SREDYynG4nEkspLMDnjaIgWwig7covepsW0zTqz2xfY3etouG+qWdHdO86G6tl
Y/LG65BvNNeynQ59lQglPCaxGrS4GHw+QXBptcZ9v2p5sWbAuHV9iNuv+joaZGUCUYNGd2kMvKJM
xbUZVpJb/mXspxgBZoJDSVo5Fvimt5Zxj7RvJg18ZG3qHRH6z13eKcaUpCWmPKUUckZzobcW+OVk
d1tLjZ3ZnqHXiPkbXz2p8JIOikDo8aHXkCSw4/4vAxzqo9RTccg19M9tZFenRlstf31yDGg74i7X
gjW6ekmaJPJZsdssXyzyL5WJbd9gCdEQz+ukZUpOThVXv5oj1Nt3FtXgGot0fRakAZQqwk29S7rE
jmC28OJgL6LdMry+61kkzDqaIs29GXAnkvXY9afYUOaSu5QQxCKg7cv3TeI05mBPpQQXPAi8vlwA
RZxCGSB13+35zl6MdKf4txrnP3WvDW8HzVY06KxZuIDd3RXGajNlO6ZkIiFijcYteUDYcG2Ty6/h
Vp1adoOwEVXY6RUtCVFMmRA3cKt3+owGSYkl4YYykXEgpSxqwuJ6Ooc6mCbY1rNVv/WGR1NNLZ1f
KiQOXlUmmbDINeXPBAvzSsP8X1x8gFNZeNxHKOSeQrceMf6hlHzd65a5jl4D8VnffxauGHsVCRhL
p0+9U3o1C9TSwXMpOUbnJ+ZMNMBX9261OxRIF76d61kkthDqkq+IBi/q16FNRNyIbGLQuqxpWR7G
EtY//bMkZZn2oGrWkuW480mIZrYUgw4xf5yOToqBb0fGLpUw5BVmddftTLPOo2ZsPKk6hsP3DrWT
vj44cyMzPUtpFWpido/ddi0RcoO1GdjCaEjnz+vFT1mwEsPvRpZOnfvIftOswlnmHtFpwC2ugR5R
/yPrMZ2Qe3EKQzcsaRl4tlOH2ny0iMjUPS+OMI/BN8z/cnGv3Igt+3rgWpX6VRQAGrXCyzWasB5a
nNYhh/sgCLbO8pD1vlsXxDWx8Z3hoKvVvrcbfOl7xUkMmnXvTAIdquK1skkDCoLYtJf3nH0HgiH4
/gTjHhm2g5IExxlIvG4fNmz6IsLP2tEIg7BIksN8AVFjufWbaxLh0nC9Io6/6F3uViVGywmns21y
7nojwvyy9Q3DsIPmM8EfaxHag/em/CSptNWhtoZfUSg1LgWbdbYVt+xlLaRDf+y3E+haGpLtHtar
7iMxz1oGnbAe+Mt0h9MsSzt6qeaUdh0Ap1tmoha8zEnoyEjnhtZuYQNFM48Y/KpCwFyinCVqOJwe
ErqNvfZg7UxNkv4d5SbXyoQr/j2Wqcp/8rP+BpCvmpZ60Pwbm8XhHLhCdnEa6J7q+CQ3cn8GkTlC
oW0SaTS85X8v96cgNL5Kp6iZfJe9zEvXNn5UHOJhg00muuRT/y89iDVjhnT2C8lGIJJsL1i69bMN
MgFOSQ/TXTQWCZ6KyEto4yqt6QWdWMo4+xMV1C+k8Kkh/2ZVFFPZZd1RzlVUNQPfdSw/xUV4omnJ
Fg7h21PCA+/pQHHVvTU5oZKMNC0DgrWc3/aQz1pHo3WImAy+8ze/x/l62P/ZJsgm0yASodMuAPQK
GFEDlI3ttA2bgfF8a5sOO7DoiW44KuCdMQHT1VWCNGdRpml/goLY52aqURemOTP1nvC5eCk02fVg
4y18ZnrOJ/FI68Vik1yihmzkuvFjGaxhXn8oN0Qo1TCtOju+mCC/IaJd+xf2aEnkwwYZGWrsXCFm
thcgIhmKXuwgJVMofeyNRiDKkF9GBPVgQ0fXNR37FhpzXkLdbQITBfYsrBYX+tle+gsWFNS24ZIl
e6t5qHhHZsUhxNVXGcbd/6xBg9RQuswJPzmkumUEta0lP5hOnWxM9bIvOnEfRb1bJa8r5fSOiBgW
W2PHfJ/IhEGiVx0veovQMFEsG3NpElp/hBRrBF0LNQTNutqwN/QMumieQz3qghZIGO+MqCRoaOSa
Xwd1QRLuMn0n6XFKazLM6cYPO+IxHryv16JMogH8IvwgHJfLj2m8X1BSQPC5VdIKXx5al54KzvPI
rBCdlqXt+GBM3i83gFLvjTWMmm3thMrqt0OzvXBGuSz/hyW4GGImQCUARl+HLyZRRQHj07N7ysHH
2SqXwkwBmH51IWyECkHGZfEbs49BdQu2+d127n7xvUjmN1HBXMKlEMtJElwTk0O2WqaeNg8M8GNS
VpptfJQxXwWl5R2183OHVv9L9ioGNFnGycTNnGXRrzh2xsX5m3JcREoPmqvrF5zP2tbgUOO8XM/K
PDwkK/44sXW0ODs96Y0nSAm+m++VM+HpP1+TksZHteXPa1/2hDvJMIv17TIqxzXI9L/hW47Jtn75
UV6Tis9HjxdVmXVJZyXGi8HgrksqQ1cgMhhUCL5j2WYahyXhRNchaP4e2SwNQ4f5n6MOMgA2l+zG
N68AdFpGTUacIDLhj7mFLJJG1ZJe6H3voDml9A1KUFFBA1Qa+ll+mFhqEHMZI7ZhQRVq4gVfwR35
PFZVuEdZpl1jkZnMeO1HJwdaFdAuHDZV7W/Zop4c9+j3ky0qPeylsQx6oXqNr4dHhHVRBNL/QxwR
z+ciK6Jr7HzTAmTUya90SFXDTvsjLSo9GxFiufaK5IjD51wrNau/PnoiZRLDa0Vw2D0s/CxnPkPQ
gWfY7r4EMcV3kW+Tg1VOLE8QdwJcoOfklneU4oWe9mJmmXVPXUJay1H2pkyrfKbrGgKR/P74iw6M
rV82yXw8qyFsej5DlCYg06UKwSH+uSBprneWVUoH9rmjfrnAi47o6YbuaHFH2DlFQXgbPdA+4hiC
gYMCg4HGssttXZODy9xDFgI2KJkk2AYKsd/tc6fR3rHj9u8oI9LrRQKPkjQa0XSdlL0s/ZUpcHP8
NNx/KOqokBCdyO8PlXwNl4i+eaUgzrO6Mv2kjWOn3EGGYRupDTkfpWiv+2EppK7SfIl+Q8njALLn
FmqNjv4ScGfvRuXXp1ZH5SwyBe1lMb30AW2Z+xR1Y4U3+780sFm5OB4v5o9iJK1GcqfOAwSySDeS
/IBbV3NJYfRkHSOrsrXjBXFe07q2lbsi62TRYFRXmrEVrfBZ1RZeo2sACKkqjCReAa7e8WTNoRtm
SSs+Hmkurw8WmEGlMstdLI1qGoGOhFSpnQwOSgA3Fk3ziNzBPrcxIQiHSn9ZBVGb4Ig+8kGme5Z9
UKpgFEc0wXwTO2pcZ7JLMrwWgQL0ZOdYSrW1BeU8UX+m1AUZ10tBNTHpxx3XRvU00Xndoe44nWfP
MHXjjjYH6qocgMQvhA0W1rIIxO71o3GXuvisEI5WSMeVElKqOjrIIdIArFBJV6+LeqCFAhkOuryx
dkJdKeGJK25GiH0dKrGUJ+wB/PCuhD6S/AdJiQbrDlvJodTRDZMixP/oVKjY9030BxAZawF1JyNZ
Vowx05bzFj1Xvsu5nnEpjUjV263Q7tv8fAQCEU+3I2TZ2+IAhzARSUqfdwhv5oznHBQEXQmlhUqA
TVMTB0CCvLsfFnPgdMLk0etamynTICsrJKwDPFsXbkTz20UN7f/BULjPxaLFZzRMR21iWrR5Y1m8
2ndRAaPDYWwQ02dwMxJlqyzG5QSTnGMyyG2r0L3/PhCYDRuolu+24i5QFRK4M4hLZ+rpXdSgEsVP
HNtt7Dk5P5+j2g5F93iNSWsvIAiXEuIL4nOhqVgwXwTSSAaSAIjXuGPm9oJ7gwYhrTzoeh7UfVoo
i2OPX9UDIkCe6pSE1h9JUf2YkbZWEM6v4Am0KBJICyfM2QdvT5iY2WTUFOI73IOhDqFYuvDnivw/
PQ7kl4xgU9KTPPWqLti9APmeWP1JMyPH0GANE8dXwc0U3ieBHjdFRo6z8pMwyMzBC3evMvBB+w55
fTbvTt/bgUCIXL5kiDGMG6ICTVecu2jcBtydn/Uh5Ut+4mNgMskWLfXuPLRMYU3qLMJkpEgLfGud
j7LpuekXj/wCw/5pISczb2i4kh7eFLi+JIKgGQfS2VC+LuKSCzvDtgbaCkqYRx/WSDMZzL+Mplc4
Lc8TFbQkJ+a5oyzamwBxXMV9TH3w8kjKmXGSas2jUR/K0kEGZtJgqtP2+4WNhK9H8ZEUqnq2E4NJ
ijOkii9CT5Y4WteS0jExuq2N4PVUsdPL4hnO2p1o1sWufzOPs+BoLpcgK1kRae8PHpHc5izK1GA6
h/+6Wxvd7iKsdEc3NXGtIMhlaGskgH6iQ7CoASIFHJYchnymfL1WlB5ul7h8oInNGMFzXgOq6t7F
thrYCgsx6QbM3UkqLs7V5MfZniCTJ7AhJQg08AGNVn/mLu8cxMn30LBnZzHt3KnDPYg8huOmsQlW
XigrFIHa5xIIAtl9HBXLIFT3bk0eYiOiuAcNWWyZGG/sMT6LE3WZ4uCN/qcUZAeiXkl5gbdfyqjB
m0xEYpF8sjeSOHXk36PFi6hfdwYEGrEb63xCVnCIPJQnxrLQHQONk3aDMyhlR3X8P2nbLwUUtYBh
VKeo15GW052Wrd0GaIfztwt8tUEUdYIaowJ038Z13XNCZzAK2G0y4q2zILj1njJF53bgnBUPnEji
MczaGySKVKBsDjOM6QnWYQnhHmc447cx77bFNBmGuH40/N6hM/U2c51R7TzeWsd2ClFrAIGhvTAL
wdoIBfaxzfWDajyU+uVCs9DzP/mNMq52UjFEMwu17F+7i6ED8hdykQCPLpEo967IlPO9srgzuJ4L
mcLzea7NwSXWqhI89dq0hobwjR0eFZ18eZyzxxxohQTLq3zM1k3Fv7lQmI7QGaT2BogfVRXDJXJ5
vRuaiH1T96CfxETkXeiR64FDfiR2cEQKO1L5KOKsz0DVqJeWPq78iO4qfidHQefYlcK9o4Zy6rzR
/9WvoKY3coiSBizHvmT8kNAZrMI/ssxiZrfLcr2a8JteIhYAMJyMVlI2eMKZrIEbFnwZGGnN34uV
rgSgCfWMOC02u57nFwgTJAMgA2sXolww44aEUK4/km79JoVPAfgx5/UzzRtkA5Ix9hCbkGahlRBw
24y3v0FNRhOSmGsF4zq1A1vF5EHgLWoA2nypPBPYn+x8GGxUiSK9DX8nGx3aPGCecgzFCxxFQ+1p
UI3t0ce2YQaqtuZdnr0KTHsqpRUiwD3ONjoiahavDsVbAGHbZbGC6/9nlew/G17RFIB/BDIuF+sV
dQS//ts2kDd1g7XcDhAk6kjmcvXtzWqENC085vhe7d6jj7i+SgPrWMMhtOXYpDVdV4GCLer4oWwm
neOHZVQcLTqMWgMKaWQQsnD14EM9wqZIvHzOb7hn4CQ45dLkqzCP3ZrxUQs7nmkA73HvXt+Ud90U
Us7uWPMdwXf/mi7//oocgYYq9YtnbS1mJjN0adB9N06GFfz18VsAGE+l1VrSpNaWbPRoSdEBa2Qk
EnfcCNusTvkY3a/UIbyjLQY+qhv+RwQtSyr6vkaeEGVQVQaXGgCLX+PY6PamvVCOJCSCWWd16/7K
oEcaMjjflxOeyIz9KY+MWlcGoDruNUl/dSO6EFzR3TeVU/2V8p8a5F7FXOru0eLEUeaSfs/Qq0Mo
IUGIHdo41mfPvRlInMhN4cVzCTJzlhg8NH8heqh6dw7gggWx/bXS60gOM8RiYjlzG/hbxn8DQzy+
bg2aPaWk5GOncrLMXeDQYnGq9xEpbV7iURuGoOgsNnd63hG4sXFJLDsvVb/kk4ps9MInrWuwG5x6
/Nkt+2VnGaBT7DcHULExrN6seKCvGkBSnbQr8gW966rYZxIf0mNqX5UtF2ftWN9cayFShvotpp5P
mlLfykYaM6MSOMqGMz8fQRacCC+L5q6kiF5LGQaC6+kyo8SSrp/jTfGBxD+JFzqNmg38+cjVLwG5
DQe/0P6KF0jMMjfWBK4m7gs6nXU/J79njisbjvQkJazTYPHHPICKjWYkDAov/n/LGvZtSVzYKOfM
dc65vTB3Tiw7U9RbWgfzYdHR6hPqy06Ch5OyeF25WlYloSJaR7GYZOmzw3o5zmEXMFVpRXSgeaJn
m4d9J2ct8Quo7fiTwFR8bjfyRHnJo7HnAbdBIRVqd6rBhEkzTsLaFesG/CYeJLFte2biuRRINstj
slQBgV8rSZ8hXKDQIsfjZR2GxNnMVCxhzQB/ZEPkLPl0YqHznFskrmLV/edFBsmAbp6g2ySuw6R3
Mx7XjaQocMcFLHcDM7GKAkXBBct6KQrAe6XVo2sHBDWHchLncaOTK8hQSYSxO4gG4+jph80yJsWs
3T4i0g5P8HVyaEomB3kN9tYhB6oZyYXAJH8afDX5tJqz6YBIU3X5487BS30mqsE2yHPd8XNlK9gs
vqQVWuNCnRhhua4G7QIUONPGE+S02ooNHrXCdJH7maWBUBVNUzLZeONO8XlMMDhhMqBmId/j2bkj
1xTbxIAlzO8yDmD44rDfMSF13Xtuze55DV0Rwqk4bcC0papeLsAXI2pep75r/dUG433JUgqgSk5T
y8SwLgvRJzi9BBDataj0VuBVl0Ifl1ukIXOj+M2NMByUxaMgoSpvIdgxDxRHKj6o3FpxliNETjUB
UP3uUXKCgFOdQ2M2LLpUKGeCOCruIPamt4I4ADJUmh0LgJFOs67Ir14HwX5AmMItq2HyiYfdmQgq
vCl5yM4BRAurRNtgbLym+GBb/C1WzTG+Vg9g/sqslsLIfKTR0waL8iEYHqaXULt+NfN8RRK+ala8
EJ7UksHx7Bh5X30x+Joy9CYcW2HCBls4+I+E/GzkHvOB1IGUvP0Htr5c6s3pBI0n9CRpyR2D4mma
zEeul73r8LXfiF0G1LI/CmO36aPpiqZYpCV1Oas1r8Kume98m/hynn3+p8wPHKwlrXw+XDdyjqsA
BphMkoxGYbkf0at75JQVZXUvvz7cFiaPHgrkO8MIs7tlM37UhsuGfvtFqTPqygLrWubT6MD7NX/H
0Ok6GEqRwe4Qpv5EMTK8003OP3IgaDIr1Y5hlJhQiZUlb9vnX9MMiPs54YJu16SLZfMnhYMUkK5f
OBxYOrPVO3zawFciqpa52Wcwf+6vahei7IVQkI7Jfv835FJDTKS84c41zBoSExm2R70623hKstVy
UGZNCf8d7B3X8N/z9KpA52ORv8CPnG5hVmAGthsqrMWjlYWUlewGw5JWy9Ooir+1owgm+qqA1Ebw
ggIN+N0shrmIhCUNVVujWR+ENwPCM22chWx/J1IhBfCGJW4BYRzuSeuiHpAlNvL8OmUB+BMry1el
ACqVLpwP/TLxuiUy43krWkNZZ+ANTpnbtMMCqaUbOguyOS4Wi9H6tvzDlaWq+knX5FpgfEdB3vzD
6w2fV20PW0O5wB8l8QASpAU9YPyJUJfgJ7DJLKcEaVT0IfDklzvlbAhkmF+ZbZkjSBVZM/8LIn72
YrbAu0UqOdMcX99QFwhiY/ZGnOfBRvRW2lvjkQm0u4kmz4KOMOQJ11EYKA2NcXs/FFtYAtEi37CZ
NR7k3cDctEXoECLWDyQLYWGu/3synkCZ0vmXxqtbdmxKEQv4QI57bf6kLkxQVFaSnJDjUJjOSlrl
oM97p4uOLsmFnHIt1Dak0tj/fAhuKP2EI9XMcfMm4WSUEwt1HhF5yO7paQ+uIHUXrKnwi3ZNvTDo
hoFG+NFUrIZzsHCKxqNtn9hGdYhdiokWjzBJ9M0VpGhH4Vm0qGnUVzD1mFG1Ox4RE1q05iSMKOlR
kwatZoQ5f1IkGsFrAIzptsmGu8gHMGIjEQpzcbyAdRmVegI3J0ktT1uLHBDYVgHoFwwwBaOMmDY2
ulolqFATHn4SREf7yX1rF9chWQmEkr4sZnuF3vGEXjpU9sBqP2NGeaC1syof4I3zPnX0R0mgOQc2
9VZmcpn0++7uuc+F94rJE6b97asjGZffDUw8tSasTPIbDjvopy+znWHJWbk+ZFB2acLyEGZfSObY
vcSTlFfAjTutvcetm30o5GCLiXWdqbIn1k94TllMRDEivW96x//uW3DBNGTwRXTStTrN4rmSr5WR
vmCGPryuGS78+vqXQdvj5lfByolyZ0fM66vWyjs/WfliVYXLLYD0jlu0z71NQ/wvpTy+Aegflf0G
1AFon7lk60B/PX06pIkFMaJnx4KytMYqYcnD71tXvqq6FeJjVBW63OrOnVQG/l8ukdlq7Tn5+SwH
bYpkSeajqKv5LtIPq8JFhI8NJtP9GOJED7dJrebfpj9w4sk+0cERIKORk2LyOFQl5Kd3ogGYJew2
bP1UKEtMX7Xgfv/5IKTnieyahqCCt8z+T+K2iwfORkwyaOleg5GJ1S/Q3yUFRJLjVd4dCD8Po1vc
Uzg5vXeI5JwLaGjfA2YpBqUt4TuL2n9KF6VrzgAr0rSoYWe3idXVUqGP6S1ticAq/L2Qo0jEEsk/
+T5GYVbuhXTQ3zB9d5gWBFg9IdXI8xEuqUxpi90kcGns0OvLh97ulZihMghxq4oCOU8ctMg+h9xa
4dYJ0pREiUkr701/nAUxr5TxOml69eX5kraNBVvZE0rVWmHHBwb9aVCDvDSN9HviIxFtYOtKXwVb
vWWJuoCXZwt32ufXqPqO6ejVX1ke+bvWkYIv+8nipgAKxMAsCaLKifHnTbv2KsMUkm4Lq6cmzpMs
y4NMzg7CaP5S1IWNGsNHG/eS1Ds6lHNK+TssEKCiRDOL+Oz4dh0Hk3g1jKvBhbomYjfehowNUYVR
m6duHwZlb0bj9KuVpjCRFqXR/l3GHuMb1cjz4oTfx+GvR+86Y89SI7FVagFdp6nj1zlYj9JLw/GL
lU3IpOU3rxZr3bv5ZsBhowiIhzftoRtn4rgku+0Wv7vfGqev6pj8qeJL/OFnymujWw+gJ5hW5sjz
aM181dDv0UwsZx9WuqWEBtvATBQoI3uiQT5+rAtgmSHxDnxhMineH4QLdYLm4HRGaAw2ZjoHNQjF
dhxBS/CK1zoDfBMBhU9jOBNhZzvjUP4o4XKXfOPoXaa+dTD+k5PZ4bBSym68t3mxfU9MeedriXzV
JbKPcWoNQMPyvWtrCPeU4gBsfsKDW55c+x93SDSYN7f7Onn36/Oz5h20RCyStfIP3RkOyaeogcok
Ku2DehhC8N/zEy7Z7HuWxDSS4cTgcuzxOf/n92QbVKDuh99TKT3S2VdkFQryTtGDxOl1sfUQz6NI
CwhKjPLoVqceuKMkT8oTKBeChL4J/Qp/r+Sqgv5RCJL97b9C+Kn5kiYMxs5yufnWAR0djvU2sJzx
U8AYKYssftgHj5Rwioj14soeifbnI3dhwwOx4iwDDk9ttZow7EK+ZPbnvZWrqNVIMqCWpxMrd7ce
AV+bSqPv3Ys6yN4VtzxakkCftE41SYgkyvH8aosb3xhJmAoJ9nytamCUuU1H5wTgjMdouYpYMg4u
HEkhJYB2Q59PRp8JQ6WYfaWy2dOCbLnP41tDM0gtgIlgIlKfum5yHKJfFDOvZqpQB/W74bEVPMJk
IeUj72E8L1/Nhl6yj+qu4iW1NlbBH+aSH0eb4nbswNlkII6ZN3j9yUhesMLlAju6PSaRMeONChD+
2bycPNQ6vvB3wz3kBPLhSF67dcoX7v0D4mkAHp7f6syZNaTCkrtAEzThbGNi/8uafQzYB2ZhO7dd
uStE48rrkXAph0q9VvEQXTjX8aSV/FnGsbuXaH3+12Vt5cfs6bjs2YKsie8B8VzHj5SXFFmHm6sS
mc2tjtQ/zhEmLKNw1i+c8gG1gQnnb+AbtgwsMnLHvbzbSsB+Zah5hmroWHGNH9LVCvbpDlwwWySD
2a2eu/A+7ArdFPCRTBkWMDsQiMwfyEjpSRS3sqdJ2DJNlw9xYmgO0wsaYtCt6Qy2zVGIm02HOLfh
o5d68heLZuy9TEV+mJ8PH1qIzLTRK+zNYIJtG1Iu0o9jvrwyTUKG5Tz4s24TbuPkxkE1j84hvU7n
3oX7S/eRpU9R7FvUclvBxtn8cy685w/r4TRWgAmYwJ+MgssKWxtSkhwkR3vP3AnAo2tjPBy/iIcN
qEzVF1JLMjV9z5Qhd724sVG+R31M/gyIBYOmVcg9R92TkXKRoBYHESDB+X4/tsStEEpGSvSRZsXO
IevlwFbl53QN3aRPmRM5QVdVzUf/dI/B5GRI/B7Gt+pvX3pv6DIjZlOEZdIcx3tx+gGcAXIojNGw
d+LP4Mzb1o/i7ra3BO8N6BimTk3dRk9bSKwPu6p77afVkASKGeAY7AwG4Yr4X4/x6jppTduXfyr6
W8Ay/xQamyxhQLTVepTr0dyMTRIJqDhx+56LO7exGxlaS8dG6mPlmpMV9nwuevnXArGNBo1FLbRA
D0VxIvCDQkaJ2/psqBxNhuUlyD1zNHTts6US2uowuoofprU76Bb+qf3olAGzIBBLxbv1mCVkHbqO
bAPdHt/XEHXcLd2Q+L5FciaaDOkKfjcQsxhTR5IzAnUHzROMn3Axh/saNUPlG3gdIAdkSQPrSUPZ
Tg/szaenIZzXE1FXX5Sozg8ScBdQPrHjCX3zPuh8c9v5uz7aXGDRkCgZzwJzJGOEVGu0hR816c4z
Ibd+UVyFh38U8mFK1dtr1ZdcVdxUHUtF4pQHRrV7IM7zZzYp/tG5aoIseVwCjwyI/K6xfbLgeJDB
PIpXCaCzJvCqCY7TV0Y5cuhJWHw8U0siV9+9BIj5fI1+A/C4Cgmxb4vmEn+VmB8B2VOmnnhn8NQk
uIuKLKqfasN4+nSUTFdRF5EJeaVpGd+OT6aGPL9p2huxehzmMwJdJrrZs05Mok7n6zisSdd4pV82
MfsmZNYpM/0Qg70BvZyiYvwGDCiO42fDIkCxKNxz2cwl48p58/Ic8sa6J5c4VOelfwHhHbcppER/
432Xwb08/3g5A3ElhuEf5yAdD50oLy0pGMfGk15owtnRAkFaz3d2TFAz3KrcmrBwcjaOGbKzo15/
rk/u/8ttscCCZ+itEzl0LNlbWY99MLzrTp8rmG6jFYW8Puo1J6KQCRczbRwcUMbI/7O5BUSp3Dsl
dIfNmHI/XpxQX4/7kjfQgToSACwFfDWJXNHOCu+yU+8Tog8vvZxKXctqIXf6evzXMCf7LTs+V5XR
gmAM9iSeWW04YNqSP+qebnyihZYKoGPKxLdkTmj3e50tiJi/fr8tzx3Ni5XCxF5RIPEspigQF9ET
z24hvukmgipqPrF6d7wXvSngtahx28xIvnng4obfwL1I3aEEsdRRJtF99bZt3YJ9LEVjPmvn8Wne
/XeR6Dns8n7T3lHBLLkNowesItC8aL32NvCSEQ56nO7ccchsgU8XVWr6nZ0jIguQNxNsJnXYEZRQ
B6F8NfhvCoartIIon7Tq2u5YwngZGjRN/aXb6gfGRtK96hmgqEE6fFcqpbniLgaiXVtmqAvTDX4y
M7G/273DHGt05RK25S4xsiOx13tKUTBX9wetEZXpuJe0cKym4/UOX/NnseGrQY2ZnXiUnTGaI2cI
VLWeA1DLsIzKAB03qBTK5i3KqXaGGDDZ4i2lkmaWswKbJ3/rZ+WHAE/0JPvGsqeVsi0x043PnvfW
XPIXhm0HMuRAG5DoqMOiMUOqudd7dl4Mv84MrKgUlpsUqvaa3/D2fLqCFk+nhILgPYzSI+ZvbKYZ
u11ILlUwPhEXlm89uIGbbCnad76AF+Kem/Vy2b8jkB2MYyKJxTDUmVNlDugjd6z8agIgvz6xgWJc
TPOc6TuBOQxqKd5ZrdNaICoCG3DtxTBbT4VT4liG+ddUOE58UokD9WsiXlw/8uhx6PW3vLlxbabU
xWSkjB7BRQW776y68NzRY2qaHKGzP+1QtCsBh6FfGBNMFrVw3EHNdgujkFHGrYeyUkKzLl2hj7rc
qBG034Jm4T1XFGO4LzQzxrGeSM5uF6/eIIZYgZuTd6PQXThUM2nT72c5gCaAMxdFCG3ai5I6M8VX
zv2/TvBr3s6kOVaAGrGO3vGbLOjktwBsUGLa36xXtlzvxWFynqCXqF+0oEO8gxvg8Uc+VHuV7Wwy
USZ8vbP0GcKNj708r7SWTfRtDs4OTWqZt2pTHhdICEVFnfyfgtfaAFNkhllXb0i9iR5WIkutHXlu
Hq/wa08Fok+N4hYpei7fOM4xrpNvVJYWS/blOdnfcXV2RoReC+/Pv8wWc/bbtTm0aa/N2xroW3kd
imvaZAzY0A3N6q1kMaY9UYLdswCvio4sodS6JvtyMtfyhj+AzW06puIPnMTZhv6TgxhDtGR6DjVf
O14WUkNBy7crxhK17nfsr3p2jj2WKgZ/HIi+L/AzYXJTmYR/Jl3tCYa4LM9sdmig9naIAC85Tj9c
uEAH1Hi12yiu9H8deEXOeFN18j4MjaDZHZ2jo2HohqXMc7mwKliOjX03ogW0ao6M8dv67MMFNBkJ
wNeGvH52JkopihXVhledshjtXoFMTts//OdX8MArY9UGmI28pihtQky8xjfgJXmpQO/ZM3rP+Sw8
szWE2RPKFRZ0hWe0SNR8latpz+ThdgskMv5hHNEWYD0m3E7m7LFQUzF+t2QGfyKztR+xf0vWr/2m
sILBbVB1UlqaygTDcdUutGwevKm5sq65ddxG2+pFeET0z31bH48LBUIC0km4zdZWZlT0GpBKTrml
+zZvx0U0GFiGo5XlI/IXU8eD1eVjcSAMNe1CoWUrp2jh+WT3hzZTe9s5RGIlCth6LEFyk3TaCUL1
DxltybxfPiq9NmfXTNhT+Gw0j9Svy029XrvAcyd9k2fYmpCSMJmBu6ErT8ffeiGw5PvTvpxEvVPP
NC6WveUa/uTVRUD8A6BMKwh7F8s3FWHSXv+JwyB62dwgW6zpJhIg+zTZ52LG3boQjeDfDXQe6XOh
GizkpHfY7KVZMlVHxFsDdL2XFiduDleBrukEfJabgNweM3+D8yt48ghkq5TYmjcWSwt3EqK13FPa
vUjHcDGFxGpAF/1TtZ+Vwb2hjEtlfObdtE4hXAf+ZbaiOnCVqihyZB9d8aQwUCWyYt9Kh5mzuksD
bhp7auIc+WMiCnDB8yOLLNVN+ippgw18TV19Yk1JVWBs+wmiWDvllHy6FmoPhSQnk9Mw38lWdmL7
iblPcPfoIKCilrdTnNPTnTXVj9JJFtCF5IYF2SFZq5MIuFJ0pNOL9SLyWfqAk9iQ6Xrq02TceXgJ
JbZe4TLMNEROyoEcTHtLIpF1tWtMmRRTpIiFTNDviiBKDPY8TC2cjZDi+Qsbc45b+GIQdSVJ73nJ
wCJ/+A1bwcbX6JGViXfy+4pOJvqQ/F1oU+6T7P39i821u8kQRO6g/a+GaEOOnb24jVAqvokejhTX
oRaG5TCjFLhIPSFylysQ+EibLvo1Om9bY64/s2D4pujwusGu1ufDgxDA2POrznQIIvl1ZIpo4AKE
SMBtFZZGjAEELKu5mmuh1a/RRAHjuO8o1Ec17H0IPyVmzsdUyRybkPSlVdqFppn+fvVKx5rf9t6U
d5poWqbY1oD4hTdF2kGFISEJ+uGUd0Fa56yFLBtidl0oLhcE+kajenPJ4ak4pQF/eYKxlVb57d43
40CtAqKB7VfKsEdKnEUFuD4uPNFoWn1DHsRvUcOt90AprwZ1b3GR2+mWvl0uFm0FREiYfNLl6ZXQ
ptkNnOFmkA5eDUeP77uKviMaJt1LzTyI986Dd+JN6c7uP8u8RlgGe+FlMuxEzcuzYH86uNkF16II
P3wHSrjDMoDdXMuXuSGcwrKW667PH2mlsb0JhCwkcbSdx2XWsBE/0KkVv1t7MK/xI6Hmr1zzAaU5
8i3oDu4P6vkGhWPIFSYBOWUt9MIS+7y3NJ1trhieJoh0yRc/kUKDLkvfmNn4ZBvzauPLrOPv/tlu
EmK+P5FWDb6jqWoOB+im3lu5uEOOY4Q3SzdoBK1JRxmwVvToFRlntkLZpP37hQh6I01S1wZAz72/
owttNiuirQ8CQBpO1m6lMLVZiN3D5Y7CQJoCtaO7hIc9J6TYJmIdQtJ4GoFzJtdYAI5kj+j+f0P5
bhF6u04QLWUdY1+G+YqbjjHGLyMiCDBxdol2Q63jmaqEiZsUFloI1K2AFU1+NVbT+SepD8HR6mZA
g9XmBKX4phiO0SvCMX++kL9RTxZiYQGzYPib8e5rFEp64BzYS9INUZ4GlBIxPpehqXHAJ32WD/XF
57KgIRcaFmnjBRunYVsvbrNLY+CCZq6ruju96nT6SbOvlI4LQA+ER0fgIVK0WTZVKWQX4C/PcLSt
oD/9nZXc7KbmEFUuzTrVH9CA3eIMX62/CixLyop+weYTLY0TePgVAIA5s+fD9AnqlDWCB7WpveF9
L3sQ39XwKxYjjfowozj5jkXc1Laoj2mJd61u4XeOCB0vJOwISH3NLwZeiTAL0m4m4Wwt24neo6Qy
sodETV5Ug5ekz99xYg8smNOCBMRb4qo5dZ0Z3VEXB6RVaENvzGgYr3BuhfQYMVhveIAgykDWhP8T
MmMQT/Ok7nstUmAkKYHdSuXrXf4pQLXd8luBcvalr+WF+VtpmcoAtIWmQLLUfQR9wGqbfsKDNTCU
TJAdZYxztktERv1XuqeWZ/eGibPOYpRH6XNj/oCGjukOdHbPy3r23DQaYx+EzmIrdVV4oghK/F2J
a+m1J5gpPu/41WqO1+MhBgieyN2MCKu79K69Zy5urysCzhtsB9ad2pZTPANhmqMuYRtdx4155qMh
0M4pZssurmATvLjxcaoDQS8S7sFwD9hINA1vCBSHXIaVrm3PLrX3aEkPTKkbf7KLiGC6S9nNggAV
R6MjL1/I88uv1pKBoBlCm+I4PHsTkN1+y2cb3RkkqRff2vZ+k/qLvs2B4LCtAz3TQfXvvKHsIX6v
8LPAgqqK9Jg4jDuQtWtnJv+iEdsgR6B1aLjceA0ilCQSIR6N+w2ZshAHWPO5cXf0JqrMfP5Cd4eg
CLkCAAeRD7hjuNDCpEw7yK+xjpFs6yI3kzArWWpCq0SC689r6DDeKAMSvutRcGYfyIzfttBUp4u2
sBy4J5Ts6sm5BSPLFS8dIMpuTFRU5O4BLzLGQs639CN42IUgpLesXqpsDeqbN6aQZOYVAmdmuntb
4XMTLdBVObQIUuETdfXqf3aSx0mXAH4fev3McVrsLUZgN6AUgeJNTdgsbpNezMyEjGrjwMi03VNp
5ePcKS2ne5UchzNtBpyt1KrqkAVwDTIdYoTqnBl49tcGPqBBWLpx/OP/snc1w7wtoMewzfnQmPT8
xtaCOQu5lyc4lX95BdFApkrdQchjE4Z7q2IifxZMONl7bb4uI4I+5YzAUKwAJhwhjqK38ci2VUaQ
oOjdP1qnz2FoPZXwGv8pFONeZ95bpEGf7O4uD3de5ITZkRbQxr2kUruFAz4Je5rVef4JPV2MIH10
Y2ipA5wS1SA8iHZ7HP6lFZ8IHskkke+5kR0JCC5AxA2ZF6WjicCehCFepT0CysFyZUTicXK0rZBL
KIzMliYwWBEf4+gG8KwzVDk6c339CJSxwnjdmqz5qLfDo68QRVjl9AT3H6QcKsz2OJfLSUnBZyLv
L8ni5cMW1PBJhfRkNT4UwbVTd+K1hXLAT3GZQclzR4CdB9/WonfL3kkjZPyEreAhecDuKV6nsj6r
Wmm+VrjSVxBVWcP42Fgoq6L/OTNOyZUZcvvaWT3Z1wpHxVE/jkX1f5dXtENv+Hrv4D5oIKYl45Mj
8I9OHdIT7LqfgBgVTkqMwTW0XEGteSqlNKhtl78c3XmGNhdEDAq7Dy/WFtctZ2PdVSOZmyj/ekcn
1ujGhgUW8RgSBsm5g51qyckEpaXaYYkuSW5o8zC/nF3rhnqqtmVIfWQbMra0WpMyst34u+ZYj1Ak
/zSyP04PQCkwfoxzXt1D+j9QdaTmrX0iHesJeH4iSv0Zk+T8w0z19n51HtB1olN9SunQ9l6qCSVR
k5m+cDskDaheYZ1nJQPGPrLK43vesfEjVckFYUcGFgsNkdIjQeyXJwY2LvEU5vZDJB+zi8gzUb34
9Ps6D1pn/jyD5ndeTegePGVTA9wwIRoCCVL6dfpQ7+YpVbqL81M/9YsYtCKvgg+lMoX/G7aJRMMT
yEs8LoKl3WNf1JGzRLls0DISwUbU3wVfMO995A10u2+qN+l6LdaNtdkP9pPtKhAwvJ/HbGrZk/Bj
r8EUBZB8ivcDj5/4rV7SdYA7vGcas4BdyaGUQWuQM8gbWB5YKLWsLMNtW6xhQLgvNqeLeRzDnvy4
kYpCAanMz0sWmhRmehjfUsFgHmvSR7naPhc1oftzCUDYXS/kka8qejnq0hZBgG/TD5M3tdoFrqqc
XAW3Fyslj8BC6d3+HiWZ5JhlXvwiXJ+bVRANgqbAgDygrobTsygNrUMPt2U+xtXKjd/7JWCRyJtj
PIYM+P+W0Tw6f+S9qB0vl4phsaCUACPy11J6pZpBcxrlVPTj4LjR2wYx04MfBIuc5kjsaKerdo5b
kwDf2iI1gKHfBuQX5gbtC/m7ugmmf7SJCAfO8l0n3rowrxZ8rw4ZW1ySRS4/B8yuH0mzU865jeiC
YiRkgyMMHLH+38i+XAZKrwT0ekiczqnVbcwb7cCJCK2EVADbesGb+Jj5fwdlgY601kfIOAp7FJRS
syHctkL74zDy7aJY0GgaBhRFLifYzhLuTJwVe6bSRhMLt12/ATBRiIBkaKMUJ/91ctVuKPhfvEei
nO+QSi1qAbPGh4AfD3OuuAmzqhVMlnpuV1fmqZ5jwXF0vnhbeWyyr2Q4OhEYV2buoijmEc9aqJTp
+rFjKRDXXGhuNiksXBewpD4TfnkFYP2R6pWrDuMPnxYh2gP/zdHeHN5IvmgHv4voW/96VdAWxZB5
0Qyn7UGMkKxD7PQF4kNG1HYXcXYO/z3waFI96H2DoH6US09oZqNB+sQGMd8VpxmG3ZuK4+1Rk1hZ
BXtgkxfkGzqcqKtqDDpAaiNcV78pdJlhNf17+FLuok6ODG66/19KMqUkCazHEj70Vdm23MLrtDuc
xtxSnjPcl3MbZU+PwHJb+amw7V38WkVkS34bf2XD9RiRHBnZGrfzr+swd0JKF9MFxy1SStxK2+s+
ezOoyJcoOXA8BNAQA6yOtWylVFO/VSS06gG/NRabMYnPybss4+7GEdMdVY/xCKsuY65kMzTGN5z6
uxPqkmoAVNvCChT/jm/mT3sxKEWeXQ9Qn0so8NEfGCUjLO+lV32CGEchGnjQCxgd4amg7jS5z59l
vPLVSiZMhbyAeoMtcQYt1BWB16bXfCpB0zJ7M0rt9VOfnM/qzU6uVVKhbLvi0Nyo5tRCdqkmPTVJ
QBYztK9fo+Flm639EU0DLwLVtLT6iTi/WLk/PfhkrPZuH23h8dOzoCeRLezUyoya3SkHUip7bKcU
r5/+wc7Du3CUYcwomF90ZcBrSYwAq0TDSkyp5IfN1a5dmf1qWiu8VKAca0mBtnPtTQrPOwIVYb30
A5/tGSO9CI1olPAv3KHtT8Jhg26zLKGz4RvGv96lNelN1b5UR+PogsaB4yYgRJtaJtXXgCdxxUL0
VNksXzvl90uh8LHP2KVflYNEAy2kPapb1HxcQ4ILrfX8PxJGJlFGbiyAYxIpNtJbrvmDtWF0W0Qx
NgZLEjrYrWB4iuDolRYQpcq2Hd0NBO/IYgQjP8xJY/Y7vUplCmt5wivFj0WabhmrUKSvfy7UtOaH
J+VrE6PKMHJBBaL0hKW6RW4GUAO+5KDG8g8LfRZo+K/rHXG+PsrCQwlKPrkMEwXL/3FEkEX2pzCN
SaJOLLbJ6UnSJmZk2KIo0ee8ph5kI9tnZwB/Q+dA+IqMlE1iyHxz3ulCvh1jtGTIw2152fUb3xP6
/VPWs9Qyh2KN9/vwN+STIjqtUd+Mk8vuRzi2wakZR7UULnb+HrdyWg8iHpP+/q/lXKXPCfCma+S7
EPfGbVwy+nI6kGewhIAC0BS1dta2KOQT98KczDc6TGCvDakrX0i736BAslkThi68ChrrEZ0T2i2b
HQeJlBY79PbHmWccQGpWN0hcwniSqsbaBD2kPI2wR2+6YBokevE/qN8LQZhTPVSC2Lsg+ZIZE+JN
NuYqmxQ3Cm5FvxC4LWZfCSB+K96pvtGZHtjk9/9RYCdJvDdh0JmNY4sAXHAEeMxN2jlljang9XwW
2/KCtMy7wqsdC7wkY+ilE99r8A23Lsu88LyIew6spij772r73/7LAMESkyXoxTudwKCRJLNjucX7
z3aHprlS9sBhBScxrpOiy8IkzV9yUo1Fw+yBreQEeuvx+zHAPrlneUhoZ4PsiB96ElO99sh2IUWZ
mi8UD910Ra/vuIpIWdQgZFzujOoIMX35yaicftuwSXn+vUtw+e8jDVTar43jhqP3FXTtddyA7rqH
X6THLu4Ehl3YIjOYG+DCc6oceC2wgLjw8h62Q1TvT5imOGBgcGCRimpzgBDOMYlIMJLoW2zr208n
zoflgokP/lZSyTqSfX92TuO2IsnIIC492ywwHu8CGz/w6VOWoPJtUeKLTPR1vIWUsj2oRHGmp7aC
PfIYCKb2AZkHo4aBSUVoNQfRHJ9FuMneYD9GQMIDtTHOazdwwpdte1xYfOk3LH8Fa+kf9S+30Opo
gRpqcxaYSWrDyADrkqOxP0QyxjfDNiUL22HRclUJaBBA2yHrapM0pkUGcj6pkdFlVwFM8aV9k1hu
6bE0JOsV6q61MZ2WwPAqDQWY5SUVEvi+dREdvreAXhOlg/ZcxpV0dEVMLzOt1h4MiZm5twfJLo+C
yOrKwwLQ4YdIViyuYts5QzErNlan3AylPjh/pq/FnUUvCr847/G8RPFv7pgVhECQ21DowQ76wjf6
oHEhbrWnhp27m6IrbFnDAuxelPniE0jrmxvK3F3lC1gsioKd6OPHKeJIqJSOVN4sSB3VWRbFMDkC
uJZPd62r8c29CKSD2XKM9nXQRRyQ05ZWGCVu4ehnlBIimwqycz8sSoH8wW36XWAR5m7skwcVx+w+
xQZ4Gj3yMslevq3mlNLfBNPL8p/rjzuin/plq7jKh7ZLzwwCsZaA4ORDVs5OxzMIrWTjbCKrS+iY
Dmzb/lFmlD69iRNiR2hldK4+Ng1JjM1+V58ukRSaH8tEqenFDql8eXjdQu3rZWs5CLlPKbCGzE+M
5zCwZHIKD5CtvujfILh1U2LOiiewh7FS7k5IgwT0WPKg+isNmp94ZzlV5kIrz+GfIiJcHxDPsVwE
OFriA/1JbJfETC4QaSoWHTQ4MgEbBrCh2FIp/BZd4bNZrF3T7USXubd7IgmQVxN/Z+QuNloDcjAg
2PHRlgSLN83enk7Uu+LH/Ukr/Ft/41RHUcBu++1d7f2aVDz5rg/cosCzrK2ALnlcY2LdfKvxNpav
GzkSSqKcXs4qe2zjzPj7ebcyTH0iC9848xaeSy+q1brIoAViE46Jnn8HKB2V36sVh4CaeI7qnSdw
YnETo+7rIrGQk1IwrlqayBxVkKvTiZPwQGECZH6NLkTeaKvN3rsI5WPlbbRjQT7jJyu8Qgh/MVQE
ThRxloguhjR9NPwoZ42zXJ2ajfAvLxijE5U6rCMeZC2jD2hG8OSR1TcOCS4ZhPXdS97c/A05afv8
VI7jpY5fCcYhViwh9FrJy0CKjdB2lkkwFFMzyLfRZlJYRLiSizz+5+lG8jgXGxI5SeUAO/dAXcCY
DtML1uM4/4Jf63ZaFro4+hb1BKL4Lid5tH+1ukMmlVGpiVIzdtWJtrVHCXk9CYBg1YhZH7yVVyj+
XNRuTWeupNiXZNgL1HaerEnbVPm1FVDLpLi2FVScUr2YFgTIg233Wn82WI1CfwedMiNTodML1OU8
pKe2HK+7uTIf9F6TOEYCRk5ifUQzf44jfMv+SOTvdY97LuQhXsduSeqXJMAf4FgrBmfjTIUMRA93
4cv0R31lsY+58Ewenn3fxc+RwCtHeH1cntcDgj4EnDqhooiDY+v2+fXTcDrZxLNhl/yGpRlWtE1D
yJymW6CQqAvURJnz44gOBqAlz+2ZujTrM7M0nCQJnhHXswhqEEld03olzeqo9tB1139DMToovrmH
Yn1wPODrdJO9EPqSPMxUq7S+fYTs2CQUK7zLUvC5DhbKy7L1pgjoTiXiLbWml7vlsoYzKerwiaLW
Tlcu3Rqp56FNp2b+kYhkAODSu6GEBawUOkXiF11SOoPpzWGE/c8HMlNSZHHDkx6dh3H16qJiGg8G
FvC+Uo3OkEVaaxAXMnExdwkRNWjCm/g8R+dxQIaQtsLc9kGJrolyS1n2/jETjdngUErr0qGR2SZa
L8517JDHZBvHv5aEbjNZv6VaXFob1K7ye02A+qIwC49w6gKYOvt/6eQEpVpwMEYH1j8iHrUSL4yk
VMBGD5VOukWTyJgvG6CNQcVg0PYosTeR61D8jrjVylhPsnwhPIGKPohs1USTNN0z/9x1SZcUD9Td
B4+gFqp2Gm/YenATltdGT4eeXQAufNcNMFmLzqzVxV6XvSynM+9aPBTEl4kaeK6pUQqoRSzn8uMD
L4Jj1/LbNn6g4HwNobk6yd9nvyV4bvfqZVGjGrngB1ZSoUR5D5sbARGIR1Zjs5QTAd42QfhYitQQ
QZQcim4pEmUmU9uIsxaHTz37TG4CHyfMCJoXyyf/vTpWp9JyuBb3YGJ24NViUny7M9PIP/UXe/SN
Syt92fkc7GeAJsJGTmbbV+/0fPw9Ns9sIQi029MjQv2pJ/Kz5D/i959QVDMfeu2vkmAZBGrJJarp
EA7SSDdm5WJyx15gNH5jBRepqN7CHGFOSfC+p/LiJa3SXdr+YCiRn/RPGdWkm0D32ddi7VzVwRtR
CWo4+3t1Bn0UuR4B5Qo2BzY+BC4s9zb8ZD06yXRoHJm8By4uPPFySOcI5G5744LGNoQCdwDjIQYX
YjxaRePMtS1hTFHo4TsifIIOZ2nBrsL5hp6hbpFvrvjN3p69deJmXtPQqQonyZN0BgG38fJa664B
sUBhZwrxmIqfnpBevqYi6KTj8oPKTOJt2fHCQ2e1zazE5gxufWZaNVPbdiCSfKwJTb/GNwutDEzo
OYRbzJqWj3i0QnzGr8RVJGUfI5T9K7WgXTXnd76oqIMZRpNBudWsd+asTeSXen7NU8N6sEIbFvBx
Fuiy9UXLepkQd+bgOxW5/auptUI75EPlqTiczPYR32AiXRlpSafV1z+VqpeE2uOlLGFxavRk5hIX
MdIPnJZkDkxUy5A8tKjbi3RltcZOPiEkJgTwUn3wKIIkLlJUtuVANrZE9YQvke6N/rTF3pUGRcs6
f3N333Hyggk8g4kC3luo7tbSTS6DGqiZK37arTlqNSb2YocI0i76u2CKetB1bZimB9j4rFN2JHD4
PW8a4I+3vhzKg7lRSVf9z7ZFt9cjqKRSsoDrsK+UUNX4xpBe+FhPl3HScCu8XSYDQvKUmq6SWqM3
Q/MzSYCE0WHRNjV+YObysw/mruAptMb8H+C6MU4AvISm9cNOR4/WjlRosneowns7sZxDyAbrDXHL
vKD5bQ6EiL+nCR3UcC2KNAPRQh1wiNatt879KWKdQJHZknDRyzbPHV0L6hd5tNb580Q7Y8FHRoaq
ty4hTX9rSSKdtG1iAz8f7gjY0INth4WqysE3+bH2KKFSNm7RoFScyqC+O6HslPnMnkjx+EBzN15k
zxKANqs+Hu7mDz0n4HUEnBabe4yR7KFVhK5KhE4pdz8/dNIJ0msDAufD5IXg6ZBxrNVQ0PUS2uqO
dTxmf/bY63d+qX/fL9GDb6xK75UaaR35rKjLmUYf6f4CLrRMWfMnbnbTS3zfSlbmhhwAXc0UfKUd
bGo9g22wLqT2eWoKPrJktqTClMoDvDTU539gO3fgWOaVBiWzjDivsu62iI7W5lleTinI5unGbOnH
/TEsqTOa0oaRos76OO6UtHPx/qSpneRL+7CeTyMv51uDjbVJRKQc2RIVxhNfcUEzS84BVBsaV5l5
+F11BAqvedkfZds9up/3VQEVICe+kHXBThAE9akTE5kXZZNLgmQNNmPTNZW9NEiSUSczcZPedAsG
7HTbq1iGBXXPlN434i/cKda1wMgOywzZE4Z+8S4zKOW0lGdqBe3U3xONjXVLNOw8Ro600pyIdqF3
1qdmIryD4cGdKwCGAVfDsFRYPZKan7gKAqQ+2nuaZ+OI95TXqgNAnuz/QWRKgdCUPzFd4yx27ior
su70emUxhRohIGh/i/0d+16efI4nM+H2ttm40URQluCqtYtyQneJDEM8R5WrsYPT3+qfIqpQ/+bi
cQegYbCzH7leA7aZmnCi86LIhS+oPUEezV7KHkMgkUlYG1+hs2r+2V8yDzUQoMYtc/T0NYPcRy0N
RfowVQfCjyRepTU7sZgR5NTGusQ/HtfZiYO6Zf1sgifTuvdMr9OWOCLeXv9ycrfPJZfTPNWVzXak
GZsinUJp75LeOSIaoCoZmyjnTGD3BcYG//cFfBruJZu5spy0AFZg9mlF8cxRwvufqT6+CNvC7DaJ
OboyiEk37mL0OmFGrKH9rVmQnpr+nyYCMSKrl/jG3x4hWjZ36o3ceGhC0oedBWHUo/RgwK3qNj4p
Ir3yr+Qjuz1rPMd5a+nvP5ccE4R1ypzlzg2oUG22jjeHg5KqUfOqmEexbjjoVCOl2sfXMc9IeaEN
mAEqsAmjLKP+bj5g1Dfxt8KAwsNwEdr7t9EmiD4SDNXJatolO+fi5nt0sTi3BLaRKZBsfk3Z+vpD
NyAljYm94RuGE+kAeXTRAiO99rWauAmNfNS5Ryk5X+MvPjrF/PiL7a0YwuLu9ABN50zrPeO0T3EK
8LhyyZcMWnq+nP9Ml6q0G4eosrCtoyAiIacXOLqc78kmWv5HO15vxluAc0KzAqAHnP2/R0ZuzJ8V
6eUhAku/5JpQpHqcvPisgXXJjHexaNzb1stbKXHfnCaZMH7y0RYyLPO4laXVNzToCekomrJM33ed
RH8WCq+tR8fliAYwcU0kwk6j+D5Hmlf3CMx48jPmzIMcHJfyb7pehLnPv/WJXdEGfHSV8EFCL+S3
8KqLBJuu4KVpXDEj8Fmt5X1CUwHnvz+10pc6WJ9Rb9vwEDzHcxY5jGNlnGNi8R8ZcERHB+yFzR0k
j8EF6k8aXzRZWp/X9usgRRDSeB6oxEmS69bo5lwlsWU6oVyyFm+qngzIRmy/QPLwY7DLZy+vS7jx
Eo0S2DEQdIk+tXEYq6aKxKrlcyep2KMvi5TQXIcGgME7HODtzwSKQV0sSFsSqlFOp7bM5pD7n/os
ODIGFEAIlCcszi7K1X/guFHN9rY7wxyuOM5stJrpZfJQlhXP1vysqPIYqAX7EPkl109RyUAyIwQE
6Giov85xTyN6TiO4gn7fi+2fu5Hnfk1exexN6k1Np9U0dvAREjOXvUOaaEU0BZs4JR+kZgWctPoh
BJb9hEEfiOWkBpuhYAG7BZYja/Piy3INerBTkgikYZ/uTmFsE4o1HCQfXw8yXelzwOslMKzZXdo0
a4TES3z0RbqWw3G1b2lPZ4hEv1i8ytk5gUb/0mQU+NtvGfdmouw54uccaPAAjPaQuODZFqkjdXSu
jpqrgaXng+bXMNKY25zpBXmLO1NtoQyp7EH7EYdQGJwivKssRbGcWt0DYY+subQYT6ovDyl361X4
fji/QByUuAdIddX97zvy/qR8gavLECSWtLJ67wdJBgHbjaXPmv2qenua8clfAhhE6nML60HWT5v9
rrI+z5cRe5NfQeQDZTspBCRhHrKL2ZNRC+gjBRt+6LrA03ir+qQKkKqealVzIm6XfvVjAcB/EOAh
3kCDWNKrJQy4mnenxI8v6xpVXo3NY66vtkl19XKF8O1613Nh1Jgk4xsrmt/tweRwplq8AMU814z7
TZz36vKlV/jwLJ1p5VYDMZtaaX70sHMOIiChW23as4nscRk0epxz7KsESesAK2lRoRBwFOextmWR
On7IaDqC/w1PVhE798H50ZlQaR37g2xQGaWEhx7EZqJ50uil+Gk11Y0wLJazpyoBb1TcmfADlp4l
s2lER3/DlFlYhzMEr3o/Q30Vn2jodU4PQtJExD7ImNNQY3D0czZ/z5GfSD+j/UBAPznuTZC3+Vqw
KAkv/f5Gcoh6NGLZyx6xFL8TrQT3c04PhbId4Jmsi5wLT7zpRh1HIY19xGD4yJgS82gb9CjLe96O
OgXgu756bEHoh9Zf7vilJIT8pNJlQmzqrt7vjJJFmshFi8fZ9vmqFdU4MVT4e98kM4L3l+r7oXzv
EtBLzw1/9BwHDlMknuNkoH78tDgujYtN0hdl9UOzOvm4cfhlQxLwRwUaYY/IpQpObA9tcIcUi6Hh
N4+7//8EFqbMDU+g1LqTXn+SXHnPXZnhE+cc+E4m7hcU5uPkJSJPhp9vRgOrf8dQwlvfIC1zV834
KRZqn9fzoi3vZ0NL8WLoZkW0m3Jh9ELsITkOPQgcdpUR3suJiJTYazSX7JrwJUBUBNLxb3/4gY/s
7hz/7AbKRLyQrFgmxTP+xHiGn14l6XvMDYpPaSQrEuNfl+9vBbVdnyYIv7JquQynXo3elPMbtQoD
iXIHhVfmc0mNjYq5fqM3j0QK2MKtH6tKLmyTQP442inZhVCGJ2A+HCBRh5CTNUWAbCg7X7CtGSia
pre1IIcrM5ZQMfnbVJnZbHvKrROmJsWTRCfsrAJAr6Xsbao7MNRkgwUBtfm9tRfN3karNCY7LVOi
T/ZJiJuLkigvTEvj9AAb9plJM1ZQPitffp+FiEQwdFFuzJRvpf191BlhtYXRl8oUOBCjJWVyFu64
2I/PI6sSXtMVF4rARuIUDJFUjFSHFZWFIkwAUbroT2O2TWaXQZMt9A+dZNVYm9iyIiuzUzEjUVM1
UOxvzvyRPkue8Mkoa09qoGSGbR3Hl7WzhC/egbRk1V4UKSOyaLI6SYcWFUmtx2knwmVKwoKSlTV1
HAukU6s+KON4xcsrsPreEwAqm4knUPcMWJK6oZHw0uWahRfuvPOv+d0/6GtqLILtWi5nVLNCaITo
04FoKq5JHl6Ikmyyt5cmNxW1SbbyU9EDNZY2ONMIN8ZnFlimoB+Kbz/h+Na5Cf1vt30cdhF6e7j6
WiL61ppfwx5+I4im4vyypuqJ5wbRl61hnVAcnAF1FOw/znkGKK9AIgszcZUNko5OhbA9EJWOTXy4
5HLjPAZ8tjeeEN4TPaYEzuxOTkQ6yB43o7HHeI5XhX9AHWpRCwF85HwzY82TSCZDBua8KzXTpMEb
yV0RJeQD7bsmJQhv0Cf7fGBO4QxhbPojEIliTRMUcD9ZRn/ZsCdvgqrbN9iGXbnBwOhgVooEajHy
OJtAYCd4kqyR/Oj76ms0FHkKuyFEzobISobYMGUTnz4zvNPWRs/eUO3Rsz8JZ5AP7SWyH6DgH0xw
Nm8mBACaoM2eoyN+AuYlA24Ge9vHPTO922FnexK/Q07Kfk/Cqk7qmJK2Dxox5WyqD31+ivcgWp5M
lvp63eg30djg6BCsrSATXyqiPHKpOVoUvyRjzcq4mAY9bmQGj0lKYFluFNUhvN6QYdR7K/L0glwm
7e4fqjrGT58LZucBtHM7VVvvwqt+JqYAqVgVZtbu0m90TFfyMAAK+JceahlnYlevDmWAGAaOrJkk
dnq91efRYj/PZ7/Wb+1M6KGpkvVoBnx4swqX+8Nla0PjpyoJxHaXp/FvNXg+u7DlsQFL3RmWGjGx
VYvamNfZtVaChvR6eOsP1sJ7halw5cPq3EveGjI/DpBTCt0pPUJC5/wxOX+lJVC0hgCBV56pp8DD
cjPr6I3/5C9NBBXNlwY4JuA9VGD5ZVZ/eUswhTL+H3X0yJWo91+VXLGLuHtohB/3i6xEdr5qNkOX
Qm7sN9g8HKonZ5sGCcWK+D0ETU4N5mJTp1wss86GnPAqhuV8MlD10gHNxax4eoI6o3l59jfrOeb8
FfruEAMnzcalG8iinXcE+zC/emL8mJeiNWlZwtLcOku3M5jx/u2tMYag6hIXJRPeAeq0IYOkycF8
zUhD2adZHtto//lTlaTaOQhBYavoxgA/eamvKKRPX25qT4+ImR3tfWAPYEPmnLTi5XrBYK8WEYmM
kht5521OWaSMq1815D/CweeVYzob/fxH0b3ANdRw08hxBV144dj+rC1SUvj6Rh0SiDAuMTShPGEG
ng8MtcOs0mC3J334c/iR2MHKO3nFLuUDShEk6QLLz8YJqiT+hAAD7iaH+B4b2ji/7QicXhdQq84B
UH905lb0RYE1NZ2QUx9djNt9JLqVrD71K4cFqIyTbD4LceHPA9oG0ZUePLNRcrV3PulipftlVLGg
7H74A+apnnF7uBpUo9Ai+Kg8T/CVsefyS7XiHGZHsgbUtMMVOIkCcI53xuC8vUuliEM6nXzvZTGW
8mkU3CWl8/61naWjszNW069cwOG/6RU/H8d3CrYt+3s9odOc2JCO76q44Cq+H0FQBO64qXRx/RcQ
reB0JxF9A6ejrzQhhJarL7yGi03JD5BQwhb0kjlleC4ghqRzEfMBAT987QoOlvNSK7Xt7ETMVf7o
BwiwUoiN51u9vchb+rEC5aKHFbTsB2qpMmriMi+y3ztPeOiRW95IAzlMQUnixDsUoJk6OVftQdjE
QWU21f1Zo1mGk0ImEdJVmvAgHMDToImOA1CVn/ZjjU7+Q6lvQk/90aha2nmaw8WV6OJwx04mtS31
UnzpylT9elNaol6tvjJ0qvrVJWXpsGiYrDs7f+XR8JDgTZyeZlw3YLWsB+fWGiXPir9AdhDJF7f/
4OBjwfwrsJ3F02YHp1xMtDjsXVqCpCfZJMRH4mqHGTzBgJrI2YmT0cWysvhrQGXjtM5LCu5edG9i
TSIrNXyTAyyDggdGO6hd5VJuNbdKkFtwvPbBypYwOOufSjjbWgsPg46pn1D4wTN38NCSgskB2wMJ
w+iv8nhsiK6EgDWowSUB6Qmfqb9g633s9x0w+3AFR2WmBoWjRqKmep/FF06P7v+cSswA2WFKzHAM
OgyCbgxGloayiuCSFKolSmnviJhqL1wi9G8JEuhqRzXc+pgf+PgHvoVUj+OuGqxpLPBrgAnkGf3O
G4oEMCES6VNWGnO6Xn30mhQuYr2xGS4SMNwGw+0dCJ3mGSNWCcEQmc2lqZu+UH75okDJ2YBocHRJ
e+RtPjs2xUoJq5mefQ7QmhrUN91YHGmhyZ5j3ImGwobld7rjRDjIwk1Vewgf9q33pCYcq3u9uRkY
g9IaJQ5u/lFHAckMvnQ+1/sch0eR+Jyni5vTWbt3IPsKAGQ3dBBdW2EipfH6vI0yKAjDQLaMool4
5QcZFjh9D1IDSd3hCwv8qj/Kl+zO62JTLfmazcmPWorbt49/0aJsomQvPNUAbn/wfZvimyyBj0S+
mDl03Oqmf4XrE576KJPI4NXgLhlSKtYyZwq4XapiOWeL1AZT3UNMvoWq/0mlSD4rqRcfAZMgokNZ
NisEye4yYj7zPrQUe7vzMu517RLW6T8XsjgSetNeDnkiq6f2mCS09obi4PdrYWlkRosQeebpRjls
MKZ9zQY2j+9i29uPFlTS2UMCmavAXcg/wVb0RDfEQwxoa4geuCE9NKL3x+udYplvIX2fIYD32Wl5
ICXa5k6KC7/auMVFuGVRZUBbvw3vnStZUicqP1vhLoyCO5/I/5t78G3gX9iqPusY8Opx0WZToGow
vTVA+D/M70lgvrfCpbgv99A9ckMhu4BjazBqUBbvi6IyUy6HbM1mP47iWA3z2ncAD4rmS/K9kAbV
03dwHDOuhcqzJbpU7NwfPOBEvYVyQBJyunI+tjSltEvrWQBmvm91zHAzWnTu13LKRT4uf94lj/vQ
5i0dNTmzC4KNUImwKWpTGWDSuAtV2hnJe1bMaeCa61hnoado0arN/6KHlbsjAro5DJMDMc9EM18I
Fd+CpDKvhDYi1e3+Ukgo4oaXy5Z8AmsFidnRsTect2IWdcXQo46w2splKieqbW/o/WYEJX0GYw7O
NmpEkYIXmLLEDRvN00PBIS1ew6HMaI5M+DYr7uw0ShW695SBk1rFcPH7zuWPGPQ9SOs6JaoaMydY
CuLihH8SWN6ZsJj/39y3Perl9j7PhfjDNlsZlleTHrHy0AXOKe3MkiEjOy6t3v/YEWE7dcH46jbN
tFcrU4ZxYH/D7FU3rWABnjOzzxZ9XJ/qmYVwoJHt9vd1e37lLW9Y7+TqoJi1oxrzny1u9WhdVtUS
F5lyHN3V+uQgyMUl0VniX79fubSNOj8zCigFL/yFuejAosFhMwincif9fl4kqNzJTlXXqj0M/5YD
Be34gd9Upp3twuUUSQhwa62iBESn1jCJ7xagOqdS3pOE/KoAH3sT0d3OveZm4v4OeCpv6rIpfVJp
oDVfpxw5UpoBWHrvIYHbrod/DTbzZsGAjQHelpAM8CSnVJM+N913RogTIk8qev88rWKepG2zpgwS
5CEKx08cPy+oEJu1hUg4ul3SAtfRRTIczYV9XYVdcwrEHh0TUFbv2WLGAhQcds1udDyAY6NE5hkl
8qx+hDNrew5To578mtD8dRn7Suh8WYNhzGvT93ityi45eC2yrCv+snc05A0Zcjx7ANYMw9cupDk+
+FyllopkO7rh8pRHhRM3KaSrWbfSi2kcaaQ0PMwjSjxa+dySA5h4L/v6X3CzyT00Rwjls4W7xc77
VpUBvB4RPUBBMJRWmbLxno0ag5pAol0PTj12T77sunqzMLFbxdyqowboU+2IXeqwf3DmsdhaDesQ
oIHfCxTA+5HihAS9ynpCy0kl2LwaDNe7+j1x1o6H6iOgqo0J0Fb0Jr49BM9RXPi4XqCAt/H9Bg/u
AGDMcRkf8tfLmqjbkRurdDQK3n2ZwLCeH2Xqpvn6n039fB06DXf9ljm2xQwnutnDl/+rC4Ea+wnw
Mre3qPCrzGAUg83j4nrpg4aKkjTYL3SUNvQJ/b6iwAI8VJiZPeA6WpL+7pTqWNaVlyk/OyBQr7oW
kMNA5lqj0DLMnHabhpnzo/mV+0+erseQ1vARDp49Nfa/8q2gPAh12lawK/TyY9I1ezPUHQ8E4f19
ZRY+ZT7CW8Nqzwvu7dkaN9bZceLykNnkh0vMaAanf60JZmxtEdwcteZfVddZk52j+ywnPkzgo/po
4K/zg3Y6/sxMCUO7WOxozl/uh5eTJwG92KvJumbMJYyfZDKE5mpcl1QUyhmt9UTG/ZKH83v/HnlI
GjqcN8wzx7MLYJIUQZfFiT9ZnpZv69B0kx/pp/KJMPdiu/KgmjY1LMQZc6JmEbJk64j1A/da+whv
oGnkGQ/FQjWzQ3o9pbdiCVCm/47CxPMY9kk4qXGG06+Fk8xKXVft0XG9Qc8Vn/fLC/uCx5AzFHqJ
CQZ0qBtC+8Aiynn52UTutqOuh7JfBHT7MBFUSag+T+thJRBeIlql2Dt8rUXh+2Xpw3wl2CeIbTW+
YBi1ylAum0+VKW1idXDQpdNmrJ2FUYnjyGuwlXFhvc4dCUqrTOGDqbrZy3f7vLPgfsOiYXM4H/87
wYz8fQSm+JqQeG3HWHD7VXenCwrHVy1UDrbr/xsz+wbK9iwHzBBy4ErjUBt8Ez0ZrTNTSPi763Kl
8DsASSTzTTIZgz/b2xVrh8pQbWJ13z/VcSSrT/m97n+ICersoci5XHEFl1dmVwTOcuuwaSQ0jp1z
fHvEL4k7h6l0VPQ4EjNR/Sa+calEUjf4w+7j1S5zpT12wmKxNQXuKWrbN3+FPjHXrImk8Il4vldN
hw9c6+WWyPfnK2Rk1wPiRi6jKIZTjTQHQO5Vd6ASlYWMpW5KYvlDtQyv4b9WQS6YxGxBmTpCj916
6xSHFGxs4+RpcCmuZi9557O1Le9OC3rMaOme5Xs+NrJVHHWcOoKdjmK8bgqbzNRAFoB7auFyetSa
F2iCuxYOGrBhWNoTbzd8lYilEwBo5ssPSw4ElsDJOZ2/mjp3nW+uglvsI4ubzakUzMDxl/axMSfa
6xcjoGmb1+v69Y84qjsB8oGa/QMB2wSyhffHI7IjMFy8ZUWzKR9H0gDacGs1ilKNgjjcEVUs3iFL
IvCI/iW5Uj8hugvJyD2w+hVYoPNqlBhWye4i1MshBpDud6yj1dkR5ogKHi03mE4EBI14Es8PWR6z
Dj34jkAS7HmOIu6iQbyd6g66gPkdzWUGjcbsVfjXeFVLJ6yX4fZbLhwxUfJEPwg2zYT9X8l3Tjjq
CVhrcKUNqB5hAo0EV9b2PULKtd6JFwkQ26gOKBvZtYYahFRPXOjXmMTDwD8adBIn2QrJLhP+mJno
n8huxTKVGE2vVNDJxbetobcx8LS3C+VAG3gV8gT7vohRdkfMSzepk4AiCYIaktzsJQ9IVZYGcXPT
BG4tT4DL0AErAb97C1We+lu8TwgOCu0i4WZC8JxyjZydytXP9I1IowJHKyBqtgCThkM8nQYP3MBr
f5RkRTHxZ1KL0DcmUxA8uEf5RdNz8SiKURnD3C30zzLkCp52rtxladG1kRJDrTarEmdr6/SSnTEe
YgMR6uoAM3Wc4TykTpHtZ0u+tSVgiHndWAs1GCk0BmvrRcYyfp1SVg9nm7H2ZH+doYRP3NPyrYWj
aaxuhE682M5cElwgaWfpkfJBXpv1o2Z6n5jzN2uiklL6ams1F7F2KwtfWnWMmfyXn2F1iNaecfpz
Bb0oDrRd0BRoLUiyhIHHq2AeXtUF2WMZo8ul6Hj7TR56Ee3rxJ9n6EB/l83UFe65nLdEM+CLz/he
4+jMulz+4GNzNJh0puucKk1WhhFSL/yNqizzmGzrSEN8pmL5AyploKCcRtJuRPI0h2zi0i1gQYLu
Q2FvqOzx54vQu2dYUt/GOMDmpM19uG94tYmgxiblnfdGuwjzbag3SlVOVBbKJXiESEU7fXptgRdn
ayaD/TZmdIYO/Mfpd2w61rSuf/mc3ygYbdWariEIZtQhYT7CWZ2rGIdSmR0+pX4R0XEl6gkM+K67
hbgJcLJMC5dO36voBmfzHOflNcOTR76HQWLOmu+2smYeb52TNBvfg1uop0Ae3ZDhd4g2oapI86Eb
IOTkN2L5AtI1uZmoTNeNKRHjSALIWHqz6Tg2aktlE9n/G7l4DER1vSkRB3hDxpPEMmSC91guj89D
bqdxfy7G+YmbhlcRuQ5eJ4CjVyvc4R9W1dRvPm3azIOKBXRzGsaDhqAeSm5gvq3XQvIAp/Vb78Kd
r9U4U9luQhO+QerKg2GCUvN+ZXmVZT9bqLneJBvo8qEhFZlTa1aZLXbtLI9UW7FWEwlXP1s8uKFH
D/oGtA/0bOSXHKSIJqFYyoHN7AAI4QcqQGvqYKyNozyZSj4Tb4uKGZie8P0PkhFmdYBrdGLtX6KJ
5qVFQPDrPXQnideFC0qr+mxlXbSKDHo4u8cjCgLPYUuUfkYwcz+0x67uGOIlS7CtviQ2gmwart6s
sYIQfm29pesvNm9oxLuxRV3lJI0nc4gRsrLdh7OeUMiiruHgEKaJgAtt2FwZWhWUC8TOdokUN5gy
ehGyaO5Rg1mG9G+KZq7j3I5HHE3TliInDoWoAlu+Dz+SjuvhAoxy8aRpDj4RVGWXCjOiKcxY2Lia
vw7Nk4u1V5Rh18Pwb1j9s74ZopArGLJdUWvj3Vo+gQVdUqdxm2Db2KspVBTdru2lc+q2n3KSPu6E
crQOp0ukIpX9s1RpBR9MB/A/jFERxD9QoU5aOSwGc/VUS2HOm/lSi0QqlWA/SCIVu4eITDwv1vz1
yPOk/+xs7nDRcrMfI/Fx4cF10KUGGlrNg3b6AciQCsFrHPk4wuPadnSp8R7XtFEpgDdZ1KVnMhU2
PK2/5GRPlqxL4fGnposJ+yH3QmFTtRHF4IY6pIm1XbkjSUjHe2YgNx5zYAiKA36B5PJWqJ7O04do
EAzRVNlv97J3r7FAu67EgjeSBE/qiHkGLyX98dz7PKB7X0HLv2Lu8UyzuxAC3Wg9eFZm2VpObl9e
QgMnMmuwBU64ITDW2mxxwFEXGimrk9vRC4tWlnuuyrZMDr5YtIrEj5Dh1wQDhWdR24erOxIGKCYC
TRLVLRKOFHHI5s/+Dt7U4uqBQtmzrG9AMgV06QeF9TRQOzSc8lgLQ4WWTRGbFy2Sa8xtwp7WT0Sx
ny1fhRDKzbMEiDnG3M1Z8vHD5Xge3qxrSeTEznmM1lZTcSyR5U8CLzhupwnWE4PTyT7ZGd9ChQcA
hFZsWliHb3gDJ+zy8pDNcP68e/lwvqp9bbcyaEhZVSNhjmeiBD6NxVeBviNuQCbUKkMut3T6/JrC
q5iKpxnUv4sHeECk7MgtYCx0zB0DSXphrv+2FWhQRbKPQvcreRTvaCH17kySZeboIY2dTKzDifut
vlAcDwQX/WsO+FDLT3NAaVOClPSIuIjs+CB1w5qhb+/i2SrGkAd0K3uzMV+DvybUVi1q8nRouNWq
xGrZHwzMZVyfklDcGzgSPPg2KUryMFFdiAe23uesvBZJG/+Y+E2N1MAwyHzBZ/qrCU9j4voGsE/6
QU+QWsZLQ8h30N0aSkLqPaC2cg8n5sZ8DYWXtgeC6073MgJeVhBMDfK5/PVSpRavHLbw2fyWXTMr
zxNOiLRdA6UDyZb+aIhidq4yiBbdX2h2CpK611eR7KpTsU4zgGb2QZG501tDdy4shPvLHvGUepW9
t3Y5JsjdTESSZIcXf4D5+nJEQw7va3g+eRphHZiK4pMz3JscfT8s6p5nPPnvFz1xLgk7n9rccLTL
B3ltoVcZeJFs0arBt/ZDbc31M+D6kOgAMzR6pLiYByZCzWgRRNcPTi5DE2dEzlA0O/WaMZfmU6AF
bfxt86q/DXkjGxymVXn9vkK3hG9RRgwJ3Iqh3aiGQggTA17A9BCJIF0j5zoAsQrFObXONr0ky0nC
q8jyJK6m5V/kldBt4k8EKwbXiFAP08ulgB2sse5fd4+pTbJIiMzToiTTKevIHM1QDFYAjQQZb0Oi
MKtWDfOVRBOJUISnUGbuY/sfl6hZE3Xm7WnBrpk5rUXCToGKClCsnjgWKYth1erA9pO5Oz71nQ7V
wj3gWoO+AAao5QyG5OgvShhBnuL8pSE/Yo39gZ0/mBhcHnSS9YZGRy19ZVGehetOichOWYAY6gUH
DFcovXS625GqafhnueS5/jhNS+4Wey7HfYMQvUcQrn8UhXCa8hKCVcv+rClVA2wxS/AefSGKunGc
G0HYT6aQuuvON95m+I42oYDYAzl0jAB0dp9EPNLHkttIrhU7Pe3uRjoGcjt6dmH6dWJY1gRp4vjk
81UNKbbJqbwrm/l/FBT36XFSs3iyFULdRUNQxjmTGNfk4U0dfdPnppcpippYBF2QzMuO4gDG1fcC
60QWPmLg2C9nYQL3Haa8alu4l3ulDw39HejUpzIipULiGmTd3QsvoOkvrEgG6tyM2v3UK6sHOhnZ
GvmERfZDXx1kb40it3809+UOiglv+8f0PbwrMCDQuDYcg80JDtEsNLrrq+1xtVA/OpPhJpVP0rVY
DiJyjVCh2f8N36Umniy4OGXzhLpViwJGcYzjsrWIwFEFQ6b8GiQPMEY9CRTedvmezKH0qPa/+QHe
MHSKVDUf3Jk9gd7unVl9XWXQ+IxP7+r82gXNIfKsAZSNdtIBRUKTps0o6K+megiaNIg2e/mLk+6o
JY2OFBzHeYmfchgztwWRqFgs0TR7PTls7Fse3cVmNdgMyN9F+1jL/8rHxGmUI/1RnRDqCcJbuMdQ
uRdh4cbM7xiH/kPpyKs+ZMa6P04zlnoH2ra88K2zBvBVFR5+qQDQEmBT5q8VJEsLvsmgdtCVyWRB
6t96vlndVrIrQPRHKsFiEGesIbi6jiEVoSKd6j5NhmNNE6Klc+5nt6gc5yCv1VFZByZTf15ehCGY
i26nSZwqcc8RgMOIpOt6YSTTgZguznfSccDj3+xpFPd14xLMR5XrWN87gf9X2dPx2LnoolYCZO/s
KtM6xG5wiaBRY9mPX1E9FDqlEgSCb7ekJnbRF4kZCfQA0O3BGY2vwzzsjP9Zyy1/rxqnqj+dNgGP
sCti/T1OHrfgQugZQZ5uj/CN2IxN0oYzkOpqKHPDFyIim7GkoBhp/alZf46hEV05KfrIzoUQwzfY
AhogiEjh/1gkrbrwMZDo4sHxV94llampFKnPuor3HlL8r97cZ4dfm2r+hWQ2UkVS166uVgMXg9F9
B+J1YWjKthVLa81cPKg/EAXCKPTs3lHBbTBn2XO5ilXzhkSkX8nSZQJyyk3lVN3aREgJr9IN3KgV
LP55hAFBOydtBPwLrFl6xaJZDR3UaS95rSPrIDIWZwwVgQsfanWM7pbEJgS7rBdh9VKD0yygkSZo
CZlYIiw+9in4vdQYmx1oB3P5ziEOnJva7rIniJxKiNyTi8MfiF5oZ+MHdOjwydrwmjc+dWg91bJv
VemoubMxYha3iTZO4juOhGX2K6+g81CWPWx5JqYIBrtqyn7K4RUoKehJ5JV5veN5JupbRVsI8/Em
cwwlOZtIvJwdEKUd1f8Agr5LFOqGwBVitmNog53GVfxiyKgCrTgtewDkcNsHxbpHVV2gumVe3zdt
7P6MkeNmw3xNG/0eolzGv9qcBB7hBd33jhU+CJEl02J0z5pdxHH/Wez2dTUxJGC5i9NQl60MQQsW
ZJIMFQzxY9W5Q+h7UefrCfxMwOjk6ouZeZ7h/lt6+5ldg6sRN0BpIngiQM2s0L+3nANpy52WxPsH
zEbCDHQ8m/goF+5lAqcSh1Cb6rDZuUsLJbHK4quxgYuNi6RrqU3qZfV3kMD34HYTF9yMTIjFL7jC
npfphNFx1nJ9UcTXUK/1JhnfkXPZ9o9qA6d/iVQfKujpdsfoZJdYRm6QFdZZekRVo3Y6hoJGK/Zp
UuvVPs8GWg4N3SuGxRQH7bboMFmsnGltbPD+O0Hfjg6CJkZ8+9DGw3f63OWZM7lVQz/vgh2szu3l
S1YnI8uFrPU9XkHodKZHKlal2kaiIqTBqDBbegxwS44KqBNxKBgZglIOgA82waDqh7FezoNsEAZr
cyLh4kN0ccIFjighP85HX3k0wheHpC/aLtLg7d3Daqlbq5tpfFpKXlnfLzjEyhrAvUETWfSab/QF
2tqRyh2dvx+uKsWXxiRwUYl8K6cN0TIfJCAJQSfzKUFQTi9PfturfECG4K3Bb4PwnGKwk70A6zVg
g/HgEfXQ9/6+9HgkXvg5n1zUfGJxXdOglj3Q5xWcmeo/SwR/JeNESNROoeonsYIzFyqP6pEeaJKZ
Jyi7M7Kb+9ylhkUUHuveqidR0juDeBCsndA2rnO0p5Gzsd7SV30H1u4aCCNe/JyIJxTeIHl+qNk+
sZKwFsE9nuSEk+jb7ErbY3bPLwQu5m5zDQuZtDa+X6n3WcKgvawgti+jBXgJpl2fblLBX1opA48X
ezSxagzSR+F4KYblmyy1/dd14evr/y84Mjutxfmqw470IyKM0gPmPedDiIRAJh6dCvrPjCBSJ3I4
ae6TrivKNHABuOxIWkRPKSrj4F/Y1zA5ZUrOVSuOYDLP7aNeOrgkWmwLlsCsNWsd4b1+cdXgZ0y2
Gq23wli2LGe6MMsEPAi+QN13tKvY0uQ7GG1L0PbrHnirw2EmLViAiz1UKHra89vFqIlh0KDGoFNz
B3HH1SU4Obew9y6G5RPo0XZZNkrO99Er83JvbrtkOm6VNHDswPePgo4bBr/Qk+AK5nIxvRheeMYu
xFC58wBU82W/c0KMcWUq4S0QVxyDsoYDYLKaPOZLDRqsl0EPJeychv1T1PvOGktAu2kFVgW4U8km
RWDmhLuWDzrw2vTQ1z4f6nxRMawpRzr2NlbXq+IuzrMLrGYs0xuKjGTr/T0DRQW3pFIkPJODo2TA
mhyuINLQiiyzZtD/aLzY5tOgmVT5xOph/w1AWqBQyW84O/iPHU0t/sHwIFw7YzA2+GxTZRkCp6Vg
bH8w/IrdBpWV0oKiBV3jMydxt2xjWKun+tBpfNnWZezRsgsiIEVfTbMwFOF1nNq0BZ4+9yBb9s0W
/2G7QNxO0l1LRJxQMnwgz7ku5NQ8IylBAFNqez4pvDSovpcrEtOkPw/v9BTQ/WKWqqL+Ps4q6PFl
H0eKsNOtxP2iglPAdBiuYMdp/c+3E/x50kIxtNGbmKFFE6NTNeBlZE2WJF+sRDGARi+TGMe3kUTE
0S7soUtWygrPildRK7/9umtQzevPbcE+siB9eNb9lf3z42mjJEp/TMRsR8aKKiHk4V7ITRFJvgO0
5qzEdeVepdPURa35zKfzwZ23vjgwnTltF1I2RohxV8b+2JU+X/oSzYZTTfRz9uv3hx3Dx4GUZKEf
2p8Rx+yMjfbeDm/AfNi0UxPDvbhZg4SvytU6mmFX8EK450MKY+T7BZ6xDz1DuwDHSVMhuaGU0Ygx
HB1vYC/40tT/V8w8+3dQwcuZ5OnTHIZ+7yqJ7ACNVzT4G8LYQj2FBCmHbI7sQ8BHSFiuPhAR9IhQ
3Z6kJv8EHDPb6mayU4/BPZV3IcxIOZwDGUUopR6TDRn6TwQ1ViJiT6JflNCUsyF3ZcDRGQcaDIcc
zCXLKR+A8MXc38CHgySdngJ0dJDE+1zInNM4cBeLZjLyQ8N+iN2DFFRW1YqLoEg14Cq7d68fkZBL
n5JZD7VkrrxfDDTGWA3h7jDw4mahTlxNy2RiPJsx1GM9k1hoelPtawjKwiUQJtDIrweJXWDRDfuc
zAHMOsRI6G/jPIKyEBgpIcD97fc6dc5HTT/ixhuhZZFk37p12SIkQgjtum87B1axFflixkY9MEpA
nyOT84cXa95qLWvZDWEHUBkb5ISe/5wOViftBDTd2sW30sK9dTY6zXHhDDz48WcqVg06/Nz7FiUZ
4kJMjXnyKxxj6G1rVtSEsk/m7ZAqojlRTk79RqBZfSTlh7jrhXm7ZkM33UQEzLNmJleEhLKyrG8W
gMl8qw/CfdV2dtpSy40OeC+tCjV7B+P+8hEBCTnNTlDJR2HpgNsjBGc8gNyGZBPsNZfR4ya2ljZT
kTztBRXaX0p2d9pwPfhXBL0Z+PmzSYkUJAyg4KSEEzNeCVIOHW3Hm18l8YUbggWZaDJzUybl2wxR
WiQcWKNQVIBc9xkR8csiBaawZH2yXu/1rVw9HJZnV/5npn1ziK5PlMOGqQhQJQOmMLVUUSGuTZ+s
kzL1NS2+/JEuQzLw86ZS7z+z4KSE2ZtyYVIDLvgFmUL2380rFwLbMSaNhK16/a6nqvHnhIhh/Qu7
aa6QopilrqI90LoBmlelM+pg2xSGOGPyxV4Yvr7Li5o0wgPx/OMgwKewDPdr0/0DRY/EWQ3VoIlV
FzSTMH2gTAIRF7OeAGj7HYqBZuPENbWTThSpGbf49H/ZXVhtHjRFH6QSKH5JCPRbUZazszPis1ko
FzuMisrl9LEbpu75xU3ObZJnv0z8cvcaIrPMz798HfkzEeR40HlbRNqzeC4XyqeBDtNRQMObxY48
+Y8CqC8uwgftVlY3bN/xUShdSUtqWqnj7GXnq/1ss8XQC25Gxp3AvDenn54ZqYPOWuYMkvUtKU0V
AuoezzjIgqqBSqR6fni74izCx37jdxK2LDzihXZCry8zTg8uHI8XYucqroAPvXoJBjULuoPbEl/r
tijdt/hgwv0akd14frhLocj5V4go/0wL2PovilRDzkxTRgcgD5tulIPQENA9GBkKFBa8ZhhxDCi7
2hbPUJnl8D9fvdILEyXrZXRGnA+ly77V3o8WfmHfCLw+AxelyZgOsj7uAosbHrg4aQvK550fMYD6
75qtRQ7/7H5D0efZL5U2pG6/APjLp4VjRwlgaV71xi9g+lAPhAeWf0jFveGDdupL22lH4C5ggmO5
rC+Nz5/9J0s6LD43Tv9KpOpTAz1JNF4pPK+0gkgAo2wnLDRfLyqnp9O6zJvy3LPdciuTLUTh++/6
KUm4p1ioolMJrAwfsNPPMZhqeVw16LQppDksAILthMYscjs+IvJqbYrPcjVz5tyPde5OVb89vYdw
+he0pEFdZV74hVlpbwQ+BXiI3oZdiBK6dbc9IU1i4l0wUoty3c4dnbEH85uUHLUZAyOPFr6CgzaT
4/uWPThEy2Co9C/8h8Egoq/Lgmebzpdri49cxAk0DTgOqNKeLe9K/WH8iV6qMKdzxjPQ27UJ/qoC
zeKNFGb0dgYpcEObJVx5nrSXjQ8vQsugJVUCC5MuEsk24uWeQ+8BDUkP13MFuo8/VkzuQFlw6GqU
OtfDE39C11N2YQpYIbdd0SsdJYdPgmCAPqukukX6DuuWRDJpGC/5CT6/le3Pxd0x7f9DFA0ujGGt
28m5yBtAmWBMoc3q5CJEXFq3w6tYDDK0j1W4OOonQhwIG2YYpYzMchFp9wOrUrKv8UwSMhiPUs9c
VStN3HlmuXrnJ6CUtJm96rvZdwOVDHeSH0wH/EWU9h2XH7+yHnlS0d2kLPgYjlKIzMY6Svo8ONeX
bCZTEb8SG9PLEA3YIAKIact5iX5zIUXuxngO4zFxjBRKPK8r7qeC+w52mMlbJ2QSSey2UfKVMLck
jZY3DEmZFieci30dhepbj9/JM6DARK08aeUYHuZjsQ5eE2JQfF8vW59cX9GHeV6ml5qrQhnsNO5e
9huEsz/KEo8uO9Ubc/UusibLjy/JXGIs4PVi5ku6wrg8yiHEj93oTwALJkMb2q9qzaMlNLZKznca
eltGpvL5JR4nrS6WSrV5RW72GGY7dR3/hoCOMcSE/tTYQq986z//+V4IL4l+38fAD6MWK/QuZKms
VjeCwVOq2/vwPhfSWpvtW9Cc1X9KdPWJeHv/7qHg/7WUEHSGzKqaOc74At0xLZDQEgE7gmvgLhmr
oHHZEbQi3DFlR6VDIgceQYGHfPsGfO217a/LsH1jYPhHLLhjNykwzo8WIpdq1hamYc2EGsrRDjKa
al47O/EgEQiytX9PrsLFSWMVF/8ZUOe4QvM+eYemLqj/mNKztOjblOZg7Qdx146sT0F6MMmOqxkV
LFB8OAw19UYq2pcLaC44HX2BVpO+BGd0hf+QBovdDhRTL860tpvASLpz+lxsQaC1pPSRkwXp9/3b
OHCETjdvhHCzonSV0tSQIw8jN15CfNBHCA1dsPMyu6MALXYkBd1DAVSKCmrJe4tv7NBmztvEINiE
ZfdiKY1dr3NWh0v9nAAL39BgBY8BSqNEiyXMRBBk9+1QktEHf6PCmc7LTfUKmh66zdxUl2EbpOl8
96tRsuSozGJIOKax2mNjxbnTsSsQVrd6C3Fnyz5D1vvcUmvTi5MSKZ2pbgZqbo80CU/06TGJZwOH
YUV3UiVkFp4p9fiBctn7EhdnWtpIsE7Qw3/D5IhD1Pz9Y7WE/zIH1Y+N4eFpVDUyUlpGqRbM3J7N
PcKaEb0/O9oTcbObQpBqfnLUa/OAoLJtFiBo598AWcJuatkkmYkTHa5fZyODgS4VhmGgeSXLBpon
w2e2cNUCWRvDJKV3NTuIcmzCZCHhOUlLoVr8/lxrOk5s2lMdattB1ILZovxn7jhGOU8sW1nJWGSa
GzQ4ZnvZXsTXuWLaGKUWUyu6YNLYPzP4ljHNHUvmLtpy3vz61F0tmAEmDPUz5css8hzsCwi4Hwig
gEL9Nwnq6+ngdNsIYO31lEfhX5NYVeO1L0eUIvHz0JaaAzYDyTnNe262Y8H9H0zQ0DBJ2xyBHrJE
pTiyI4YzGuDHvrKVN/3dbLqJVqqE63MRPjTu6Bl4oa2bpHYZYkXsvT0RDC/JJxU1fsMniKTeViqn
tT6XYTT4AL/KqKZ8O6dGjVB480uvHY1XjcOKd4ADUv3tl5XL34//PyqJb7TCXVEDwwi/0faapppr
IByImmOA4wPnIamJpuVHzQC8ibZK8U4K/1qEkkijDEPday6XbGp4c2TuMl3bNL2vm3+hLb5MXHZm
zaauHdcFT2Pt8ES7O+B0ZQ+1Kly4ZORYGtln0Zd/oZkoNhq8CgQn21aimnlxvD3aDCIDJ+OFIW2q
msxAIMCvypOAPYWTmnZlpUHeNcYkQkbFY8CVjtj9ezk5UXfknymHvb1aEQ28HasZvtMiOudxwFv9
u7XpisZpTh43vP2572D7DKH7ITWE8RxiAeZd8oLVbZJjiKVpsLXPmnq8oyxeYyZwwdLJgmD/xzc2
sxMTqX7+M258X/uY8TZ5msurwX7E35lAnc+vwDa2g+eKulx5ZsFzXLLmuE8i3IHlKm7Hbd7iSHQl
+21lkzHxCe7OIB9VWD0LogDyew4RVaHSNoTv4rosghSPFRpmjLyvh1G3XUq7+gr9LNFGYwisPwcA
xdEgAg8csMoAah5if5oAz4SJozwGpZg+6RBw3VRtRjXe1CW7KO5gPj9rjjOP+JlwN3LulzRfmjGV
zR4L+0VsCyStLJbqVQsNY0kaY29Dz+tv2NgbPLS+vqUdeJpiHNreA/V60vqNogGLpa4onhybF2y+
4IZlE7ld5qAqBi52KMvhHOdw7Hrxil/pQf5msJyEzOoT/TfHJ7zS43cRaGiYlpZcGIi1oGE+kGkZ
Ot8Dm745fR2/dHKH5DOYTX4qyMni+dWcFd8yrZcVoW/0++0MFvbPoyBG2mXeQmKeIu24aQuOfc3W
G142eXaoJ/zXDzmQ+FCHrtjtdIEMOV9mleiD0coNCYLnszUKBKBstUbjkecMzcSNUqbXei66piRb
CpUDLe4PyFzb4FQUaB29cZEmQ3ij2j+4takhh23z1e+kaIWCZwbhJbOROyahO1/g3dVzeHnjyMln
OTy8H0w/zkVy4VEaNU2g7Pllb1HZ76enbG9NKnx3OONbPKdkLkAvwtVeqrkPIgdWpLIMKvnvuONz
1BCzbjxnIz5zJGOBRsWPqIRhw7S9s0VDFtz1v23SkrX3UwPxqw2JTOO9r7tRiL/ezWhBicaqtD9E
jhwMaroKsneBU+OJxRVbXbr3IZ/nbqVIH0S4atzNu1/3MlhWmry61tI7GDxe2NEqiU0FypjA5leM
5Gj+AfiNTqexJMHFfEdBTuAPfBBfwd2pAf0hFXwmbCzM/kHkypbSxFAuRrBuUnMaCdy89FrLLEnx
uQOS0uRTmCVZtN5T1Gr3HvTaJTRjob+ON4jjPUS7jpFYZhrNTfPjILhdhAQUbM1W3waM0eBVzKlb
XGpfboxUFLkRqKC+81j3HxmepI8IF21/lKWwDXt9ey6ix0KqiEz0Q9PcKJqCivGf0Xm5JxFzG+SY
WgyIqj8qP208JJ0XHhhhidQWgrios+BU57gf/6eBRA2xs+7WJVFty8t1mrGXdWQYIpgPxDBaSkeJ
02lzq6Zb1ALuEAZC3bYPmQMb3ANlp49jKKevlw0ta+bDd2s95Osc6BvZDB9hiJDHVCfKEUAZLjLy
VsF7nbKgctXfOUVsgeecBQVN2bU+/GQPaH0bemJnvPrxyS5m4Rhg3q2FL0Wk/lqCXldZX8nps301
7UDCMjUHcYv0CwZAA0fG4/WHD67wR+e5KVV0c6XLJY8EqsvEKWQg1EE8A0fNUYDGf5mw36G0Y9cg
e2hfDrtgqR4POblYHDQHlmlg+qsbnTnCPk23qLHgslgSo9vU09mkpFRh3Cnj6PTncw9/Bmqt7kyH
iBYaEN1L9nauGQr9TVujOsIvRGQFpt5HuPE+3EEgspQ8fd0tKL+8lGk5HypfyFrHQmV3c9weVpPf
zKjtUprUmePUoyU0FhU0eC2c1VJBkpolOfy5HmPljG64i2w1LFWM5AT7lNp/ltFW8F5B4h3SUlGy
uHWWlSSFshPYvvd2dHMXDs31w+Zc/kdKqmOe+AJC8ugHWy2whfgsDilZj6JUM/KJQYamIQ0UIxxw
Ru7ywGO804FXr2Yu9AAJFv3daeNCvygQ53eX7IMIsieRrtaLkMV1tYk0F/sNNbawq9APVuVU+dl/
Y9cvG8eUFqvxam+QvPHaovo5Ga//u18zUGtX76/VFULfmcEtmZhxdvowVJywN+PjdoPpgoKPe059
7I6FTe7Ot61eQIKwwNldFyLtBvc3Vf20iGxTUtwmMzZd+AgtCrVPhXMUQ4bobIqkOMarF39qeRoo
Un9LqbRPIXZijPdPkGBmrEr0a0uhNDvfuNPA89j+R7hudiNJjnbrKcaX9Xx/A96fwdzMYnZwADpL
ctfccPojzx01xWhDxTK/t03gfDUOKVICyV8YwLSpTYmHZ2HwZC0b04qMqqqUXF2MITaQiNLuA2QQ
9sPvAutezmbew2y0Q34nFPisYb196KL8xXngrs8uBjoPGbUUx5IvlDk3NFC6mCaOQZouCFD0EXUv
58EbagyLtxf322Uy6v5ZbcnDfO/5Fb38NvIpL9aY9RbJoBabANMpvLpcnd4MHfXywTgQALyqpLfi
Q/ItQPlUw8EjJUKibAlP+jlI0SiYxOmpQJfg2uv2af5LlN4yUEvanyFQePghWa2R3af+8oEyDKkF
R+yO4ba+a/9VTc1ivZxiGeM2NsEx8z4sJee2DOp1PkNqWhznjgQzxeWbL/5Oi/L3YTFLGQ9rq91M
52EeZnYYsR8x4p5suwjdgPcUSJN6SO4EjwY68DF00NESzlJAlMKZgXTtt+SrKdcfLBnqJzcp0EPR
oc2ETuiVUDRJ81whoz8wh+FZga1fCSGE80GitaO06y4pgA3fhAzW5Yuo6Vt/70ReBfysdh3HUGTy
yApIILqL2wMvO/F30FXJvgkduGX27Bw7EjmXwm3KLFMWajQljCKtvwC2g+JOQuhEDA711wSnRj45
LPk0nlySTkEmmsGkLDylqb7Q4qmHHckw+oSHGL1nhs6dHiyhw8wH0NsdLtXTj1EdyU0i2C/fEabC
mG3sOr7ZWgKhQUZpdYwwCqnbl037NkNjSXYOSvWXzYYy/CdQ40GdNGmKs4G4GNNvgfiILA3gTSEU
ul+WQz7AHPd+Fvd9Drd0YkikATRuER2t+lwK58cwagMw7yAmDAOY3lMWRKc1eEvAlx0MRev9S490
8Lp9MMOLDRL+flvahXzpgV/QRIRKOV8sY1UH3r4R9KCrA4Q6qVvcUPCK6PBN0xpWj20gCpcAtrbz
iDCrYA0VDzbbr2msDfjL3edH5JWs+E5GUuFqnJrc42BqD32zDSkqxC1IU5ctBekvS/2/qqZ33EOs
nOdPnvwnsjDa7Wfz/7EIggO27Sq/bdzMoamEWe33IrpmVf9SbhVj3hD6eLY/qnOuIa3iGrWHYvj6
srqOMYv3KhhLPGzGGHjJRdQVWLNt6cuvY56ORb+jLtFeNu/J4uwTrgoiWTVVzyt5lWjS8wb641+7
LMKoO6UD/7PA8bRlLO/S1lgut1gH8NhtO5gI6U9gWGdWQi2AuqEToo99VMfszA/iegM9eNjWuRM8
zrLFSa4xrWioZqPhr7CZwqzAKgPgCJSaRpk6ZacG5ItoWsch0OIwGPWpL4KS9aw+o1chLK/yT4Vh
N9UjsDsmZsBUQh2AudMNXhr0hs3VGsWvaTfjYS4/aFPhsprO39HO32i/fYOwD/ocDkYCp3tyo+HT
gw638XDGM0JpBF8XoqqMPzuNrFJAw0dEJZ3WnGANo9RUJunPIRYILKb5zqPFDXXfRJMDFQ/rY5l2
oUakR+yLiUM4m+8CP36Wa+Mm94FQdb+AtPQEp3xbF4twGyHkjB/IX2QYSLF1UV2Uiz9hTnIKimPR
LENXgHcs51Vhh4Rvm0TKMUE5GFhuHhkilIAsuaVK1d7icBuGN9gBIa6cKMvZpovKMuk7WKIUqFTe
/SSWxLtaEY96kCpJtF/ykmvMDwrEB0aN866zNl0IemfMzFWQ9IA+NobHIQ2+24i2iz7if3aa7rK9
fPKud+S+ksSiMU2HKN9zvLlqPHZLer30/eY2Oq70HKr/CtDrlDQbN7Tf6EzYJHuO2+KvkIEma2FA
dPI2R47r5I8sv/hRKRuAolixLpgZ6eHQy4WfTDq8uDugLpJKOyOOO8VxXW+wBNy+h3CLOBTiwFd6
kkYb38xRyMohZE5DKEIc8pc0s02LeZoVO9KGRKDFxMnliQTdbQx9Gi8Ay16ycVAJiIin1iuAY+Hj
NN+oo3NJ3UksA0EZJiJFhVVISZaThp6P7bm4QfXLWgpnZEDEPtyvtl2CDObPXDboviKPnRP+tKLy
zWxOPQ9HuTPb4rV6ygtKCoiG5+GbDCVU4ereVD0VO9gDOV63MiHyPJUvCEUUtlfXohn0Fl2hUjqc
+V1sq8f6ZO9DBIeLNsz51XjpCLb3CN9LRXZuZSsZIgbb/QAS4YmLg2iLSOd/6Yau55x31jGXol9M
lmxMbLFwkGSKVtzVnj5rIP8rEFHOpT0TDwP3SRY8Vua48oejBhLFhCfghLFAKzJ5z5zw6Igx9kz1
N8kqLhlmka7W2CBkiyUnzdUWOsvnVF/76TAqKcgQs6+y3on4zc7YT/pOd/u8NrzBW9sTNt0KWVRT
Kfq/DWYU4DHGiwFl+ctgTqYA6AO/XuBFNFHEEGVTRKo8viL7t6GxeCSVKOUBGALgH5wN+Iwlm7ye
0FGxqJ5aXfifCmLvvA6m2ePcVP36sAWMxGBNQUA/llmoX41xvT/9toCBpQQB9lV+jfh5mHth7g9h
PqhOoMlqTPqbH72dK+Ovbo1mXPQxkuSArNhDBoi2eUxGHNqp7vaDAsX6WrrkWqxFTSIm6O+NUS/H
UINGFuKZg9ItMghM9VCy7jW/2WgxJu36l6PsH+Ng6jYFx1vad78WFmgxKi1YHg+BgOgTmZjLKFsi
qfOzNju4uyjB6kJl8W/+yyAMmzPmJAr0iAFmHpNe1v2WBW6JmhDF9y4xJA789lXSKONEYZtJS23Q
m35P3uy8b1HDd5AOQz9UHMxBRaFBU/dUp0gKxRbiTUVOCjAT4niZAwSyzmXiYmX2yO1Vpasc6Xx1
p3tbLVDtRLlbCTH/CRPaf1n4BcN54VVT77GB9YcaFoRUFH9OtX7Zp1/y6X/Ew3wdhFvJbiSLQEyD
we7b6n9dlwsUQ8fOh0C18WrwPickFEUJDNdSAhqam5Ps9yulBuV/elVfNT7yWOkW7EQIgzqhVl7C
m8xIFmF/inOICjN7a8i+RK/BHPO3CfJ0cF7SuPkkhfH26fX+4sD1vjSfisiqAS/Xb+M6pRW8haiP
nrMvWkLvJk1rL8hh39xXuB8Y5TIPCztTRAJO5i3ps++BfdygJB7oAVlanNmiCK61IFF3O422rfZi
mLuS0igtnZZCwvhlXMc2s99KOYBdKyq/T1fle3HLyAd9roQhKRPov21fmFveoxkiukE/Vhoybbhc
TfW+N9E70Y6Uz6QCVEgDx7QPGzImBB/qylhXny0EPVBvgQXjNWCkNoTrlS7JxW4fFfxf6G0cVhu7
tLb8Fw4WCZnLvhOT7y6avWj4Xf8u34Bpkzr5MxQAB+bXiWco6a/GOZtIIto1qcve4NpySdQ/DkAH
R6NJIpZ5erxG4padB/t9xkmz7MeUY8kj3JcS9x/fxVVzQhTZpByyL65wUqMlW1/fNMYNLZn4DhCT
Ol/cLhmGTnx+hvv9MzXiNdOicCl51JOJVvvqFEErzPhaamnQbTyGYsZRQfa0DffeoND8b8Sjz9v3
Sxxv7eZFlQagOqoT7swwMmfhYkARXSe303HXfHEUaG+vH71Tryq8XpIgAkhua6uqbD/9IbBz09zs
A8TbJT2FS0XuptyL6cU2NtxeAc0GKE9yQLC519rcY6t6fKq6ELIyCAFuOMAt3QC2az5lG3SUplxU
UyDzHVBXkE9SjAZ/yPQ5e99IF4au81SLfKdcIn9LNWe0UHs2xMzWrAsCqDbV6BWWs5yZad3GOSp1
HdndF6VONY7CmrTii9I/+3pYYQ6vh7qifuFAY77/+hoCHb5g7n996NPgaTFM1FASvdjCBcm8IkRn
SD69phvf+eB6K/DtVa5zcSN5f85CptgoMG+hrMYPT4VDTW+hsIXm/wL3EwRm6EggnJNhjv0T0nfu
c3dw7gLf7UrpPPeozbeITGhv+CFArOWAAmkqDYihV1DnQtHQNxV/TALOhNovLbYUhqhrGTyN1DdN
jyHsdQpB38EFTme8enV/K2HjHj1uS41pzEwfRYKyGFIEpQwvyXS0dds4n4fNu1VU76+yMAMSKT1U
ug90oVMHg1SwF3n9lNc48LwjT5O2URBot5tDtAQAsLQoF0DoMfovLLVRSBbMFiF1zsELhgJ94yxS
d1pETzWJj1fn3HJRb8v9CsFL3Bh84negKLOKBX4jyn41L2E7B8rfwpT9KN6jw+cV9qsI3hlEYsMJ
wnwpWJr1PIyPLZkcTRwsghQ2mmxEsHoVoHZFyKSpcg169lElFOFL2MhZwrrT81DG9uprXctVP7QW
gxl0bhNcsyK7VT0d9pYiSRy875bs28R1EOBx19PKyOYjAsMB6YsGBBAYDr1FDzyIL68AZExIVfsy
0Wmt1dHYytXy8H1/L9H/PGa/nyRpJB6smonB+myprYpAeZ6Py4g/c78kLjC1sisRkqWbEhTIvw91
8/rmMDFYVg496xi0vSSBozKMTU9Jp2Sbjbb5nMmvzfsbvi8DhiMfU4qA63wfnmkRqOrj2+xXwGJi
EdWdvlKwgB58RuEaHw0TkQCur36cmLll4L6Fvf6PDCeN/03bs7awDD1305naF3+WwK/IisctJIIs
bZpAT06MLqqvE4WILcelh8c1+4+eBKxrHWCqcbQeybvcGI9VuOhgz5de1u4ft8qZxCdE4ex7bmxE
9lA665H3ODgHqUN4SjVFHSFhk6NBM10m/lEvD3n6Jl3WV7NWw1e1EXn8wVd+ASjDYKLJsLXNdCNJ
0HJoKAseVHzR2jcx8M9zXM9sA8KQvASmK0zXZ/BTUMss3rZ7DzYH5VJk6p2w4D/x8b1eugJ8JWUA
tsbtKlrT8oGYfJ+Y9lr3kVF2upEkvp2ttgfXZS8f4wjsbnVQ9UJlWnPHv/INGg5chNVOH8jwP2PF
NxDZK4RpLjsC6T6JORJ+4IOCzpnWeDfnQwV4HG+/cNH49Nu8gNh9KU4VAhPkQmQB49iP9twscLAU
GJHPbGTqQai+jZUxkJm4t9OR33HHZWD/XcuXMxGBaJQaA4yhpYw/6YBSpLds766x79SJuIawCgpG
8bjNAqLyrSC+0FsJQr5opNV1rjZnaiU/u/QvOLQsL8zRXpG1byqh6kWLxNhxUy7DHgTGpmJGU/Da
y1+XGnUiWJCLPVealcec73UhEy9T+NMmXHpDhSIP3OuBv9BG3x8Zrz7tbVc1jR7Qwk/isX30artJ
RwDvz5EMg5igWypO7LzPG+NUf+BZDcYaGxlT5CClKABmV+2u79AFW0OBsdPehRmBZEQtK/RA3KAp
FiN8NfCz9EvlN7vWjtD6/K1zd3u6rSQcKNGXokfd9B/piZ4N+/VPCLfYb/pABLMJVEJUU6jYx+Pz
xvVciShFFvCS0X00L3YAuiDIrghHPP33HGMfR/bphN8KoxpCylUWpkhMtL4KIU4Hx0/r9g+a9VFA
zwYxjJXvaQQLTpGm+8a4hhllizd23BBEYtIaSA/eIkj51SgJSSRNT6a2RleYmQ0NwjVAlAPV8yNU
6mOPiUywKMYxwHiyhwlbH9RLnRjXm3NBe94G0aIZhxzMZEIZywblyMwLwPUqiWczkgtjaVpeCuFS
vHEKcEf8TsUR3cjQRc9fj7f0Yo9yKUVTiACfo0nE/8uWaDbbNiTMbnuMaPl57fJpiQ6XYdfCcVke
CnaNNvw8HltN7E1DiFXm1l01ZWD6Wcf3EqWh/wy86jjtT5DZhkFmtJ8HC7wOFeah6IYA9HSFE1Y4
UCOEgyJJOwKtheBcE5r6C20gq71xQaz8pmlwKHMv9SsfzwOHXiMctj+N2KuUvlZltjV39vEd9lL8
yRn/R1KUSxxE/yoVaPMjEK5uZeZcRGxGDI99wWfk4BdLF/eRP/wv3B86Mx2o5HYg38XAVHDMTf5y
Z2aqbgGi3Vj2aicMjoRC8A01919S6mGokmsjv/uTq7mTRXZCOxA0FcSPIQgToBNzBRdpp0tYdoyu
0q2tOrMUwQm5F95vmA+tt15l6x1Ndretz69QeNtr6Y3IZ2LiUlg7NngViqNZ+xdtgTsAOOVvlIc/
y1uXPitLllplG/AHLZSZJAZ0m48IDOmnmKSkTz7uQbLaKu98Dc8PIDmNamrg+OtKkObe4XXGWEIl
ENt6Xg3X96SAI/B2TmFdKomjyh102fuxz9BEZuUGU+6ojiSkdwz3pgCznSQqpKMJe8YHQaeCDQzK
+mlZknwZoyxaryd6vPH1S1rOCvwlR1PD2+b/bHZ5C9r2KsO6+mXVUznj9131Eze4USO0LM4A04mv
sytTdoRYEdlsGwQYuo6nCrciONirBpSPCGxDBNIDTThcq95zJ+r8fBvXVSJzIHkRa86VI4dmBFvz
0pnxEavul9BTQaj+UyZHSt1Y+AJRxEf0KnrLSu4aa1JOSUituL0DSglLubpkSev+8mmBE1OjIKdd
qS94wTPkn51z8V5u6A01pP+zFcmF2cbKtgaEGJKYAgCd59T0a1DEFzZ4TMOqT6sjcZednwyjkcJX
smXxglQkrQnpKoq2X0nblvi6lCc/wirVgSFJWs+GOWYa7dQseUp4vlbo502Rqfgrt3F66j7la+iq
2yNGN5wWRGq/mMpdbCcMbdgHBWowJgwrhwi2VdXA6GpssrEVWBItzf1zuw1aHzRyedAwRSpJxtqJ
dQSmMWVvvA95EbFMbrvGtJlLGZG0agx67hPPF2Ds5v0sEmuy+adj7zsMgETcFsVNVmB7Y1Nba/pb
oON7Dt/oafbrQiBmmKJ0XLjO9oZI1bsvS2CXc1Rwv1oGc/+KtLCAEWcrjvdy+00/GCA8eCh+Lu/G
k4dI9FFUvo1nkUMd9l1HaKDulRE65JrttGAYPC231gh9GiEnn1PG5Ih6AWjlq9XGO4ftgWE+YlBJ
EXAhgbx2Lu7W3UT5OGOvp8rmK+LhaLaZ+uAtpH3KzCaS38j0SWPiSCeND6HfR8quqT32QLOvkHwe
lnfgAwrXhj/CJgLjmvbZZhgFiIP8huhOYFQAgJK+3S2JoVOonQ1nLfamdcq2BwqSINomvyboKpKz
BvnhLQ2NSVanfJd/6zGLsKbjvaWAttr34h4Oc2UM+A5PlgmIg60WVj7Yh+1YoMgAJ0MCrXvInKNR
eN09SWTidIrcx66DmUepK9zUcQSHJOa/Tr3apwdKuq42cboxCDMsrJE8OkDBoFL9bjrSON1suaTG
i/uI79/U8yWk66tyeiXiAO5mchIrkYGMPxOw+/7DVSz9isrgobQT7iRTsTmZ4f2QNImJQzKpsnOw
1Shf3xJCYRwJkM74yYIA6mZT6+QuMVIAgkrkSG+5xWRglW2rIaqXm6+g/DqaF6ownCh3Bs50lF2O
M8IObIFPADlu78kMJ80PnGAveZ/0c6OvqOrvn0uGZY4dbgTr4jNeJP5IFBXpZvrWmuBRlhio8QF5
ZaCGIfryVqahi9yvdfvMa6uMe0j1W7wRORJq0+nZ/tUiuZJaPr5KsdnKYLB+vQpnqsYbIDuJzaUT
riev9R6ZjpQBaYYMSurhcw5GIvEGvgf4Mu8CSrM8+y9MvKQTmlL4swFTFrHNpZqY1eFg5gaHs/N7
GUTIYBO+miUW7HSuhqXFD+qpXXrqR6jK/n6Yd6j7Vg+czwLJN+m0yn6BnV1z2xVT7RJYBkVStWXS
T3oLcLy97VjsxmVljUJ1rF7ZIH6iBDz0C5jGtJsxRQjbzJ9alyFdOQ5IzpSulJCiIoqt0AqPnutF
LWUinPAZReyWYXof+dEhRhl2vI4+J+YLncggLPC7DGTU9iVkaGVQf5KaLaYtzjCBC3k/rupU09eY
wZFYv9JtJtpg116BfCbHVI8eb+7BCQ5aoNFB5RowHAVWz/01nCpGDVfZxpQiRcNkxMxcSD8Aw5qf
nMz5/vVoR6pnCRmy0yuP+wsI2Q+Uk46Wy29ogxWb+VNN7Ghj9n3A8Q6WFw9iA7ZW4OH7wI77cx3+
LxuXxqooFZkTun1hII5S4gKheT/ddp8LZflyVtp6QTJhsqTXRoZZue8TGvd02MBo5LSzilLwQ10Q
fzPvRB5LcWSVbHHhbYLJvgJQsVSehoS9CoMutvfoWyxbiy9bjxIc7O6ubfYOSqnMcPnVH9cveqNi
v/pYtii8V9QCO/ao/yD7eTbw0Mojw1yLPqjwZPsC1BOepsawMO9BcVlavp/OmZBjUboIdbdJpL1N
Opn17GGRVsPvB1S3nWoyTq5NYtCFxQfhXgtBJCSlIOryZKt4gpLG39sneCE4BKxcXljQuQc0nxFf
RXj2QS1onMbp5Av7U5MNkyyyTvr54wDczeReZvbetfLkWx6ZNnkwOGZVKnHVrchLo5rOh8QILDNF
xE4eArWOGMQ7F30jcjLFCN+vhENFCqN5LhOazcE3evemdHQChOz4HVQh5xiZdnSzcS7VxTQ+Pagu
qUq+crflZYLn0VxTpKfNUfYc3wRLGTblwwV3GMy4U0WUS0xMwxlqte8dtnJBgqzWcU7Qf/YdkUT1
mMiCKBoq15MI5A0jPzmbcvvcgjHDuS6nmxmpQLZjJknxG66OsSW/q7L4IOg5RvhfFI+84myIEMrx
eTwPG1fnpbRRo3o5VSQA1ZUaqAi/iTjgY1xIeYndtnf90CFucUy73xDR6i3BHtDKktvz1BqtVZgy
AsHXP2KYDZONPuM1qIui8gjtzTz4lZQC2SdKvmaVAwLGxXcTYaY7pnGztqqv/XY6R8Y1swN8O+Og
8rdrOQ1iVQp9irlX3DM0YYIWuIcfNCsVd1CY2rHlO0g/32AYB1Ve+WC0/2U9+9JpBgiKuIq7xABR
iTDQ9F9DTne+v2oMTGV1IMz/ZWnXR8fduKJO/3zsRdUlmAbwewwD2vJ+ltJjMU9b2RTkIrvGMi+t
2GsnP+YOInsUBrLU5dlIL4esSrvSSA4GxAjrAlu/loH17H5T41YZFl4m5W3BUypcaA8f2D+Y+7QW
5bbdHY1AQfyeZ+tMBE/8Hd/wyhpNDyq6fvpvzhgZ2hBnNhoJVWn6c3vP5ieRzqkjLIKyCCdsr9SX
03Lxu2UulAOOt/fldYJIOnauGVhANJWeltqmh/KIOjiENBTEeeGAQSxuxiIMQiIvgIrZiSuVSVde
FIpn9P9YXYDdJwfK32JRyCijcy+hsx2CZfEll77ZUVEKvNR+Zb029q1oDuMpM86xpnfEBW45WIFh
tTuFLQCN5DmR21rqOgbqeINkWsAJ9UxGb8CAN061Jn3CnSlXmf+s+YQ9se7Vo9D/PHI0qRGdMrs2
joUxH8K3zAISyP7hRzBEZaBdG4sniiQ2LBARlEMzKqQ5DbmdCom4kwdNIz65bPtEswSCbPYayNNg
bCVxva5ZSX7Lq4QtzueTsSvJY1YDqSoNNM1YEhb8NpQdZFwALiUBklabbWJZofuVEJtonIERlH06
jaxKAg7sf1YC+1fDeMBOcsu558s8Q6i+VIChvuBNdDjffLc01lgWPdmI8HhivIXtMeqkiTpB71Zr
9SAh8zkw4RdvOH+OWgfkG2l8Yt1TbZwdYsYPdC1lenW/4KAinazDRgi9jBK4QYhOgATYUGMj1MES
PVpGJT5R2TpYNhvD7bh1IOR91JtUNijurDJEvJXJhu2vfhqXBOm9i19EGWEhpZSWfJxZKC5HKuuO
+QyBIGndJsdXHhUN4v0C8bacOPMsieeYJdDduaPBhBuVwXq74bx7N6S1Ez9oll3mvYFkuodEWird
2hkwhHtafBfRULp7THkxiY2BYezknpMPfSY2WcHqKJZcyB45bczO7iuT5HqozRpA4Qt3ijdD3ZR1
QDCUBnb6CNaqHPY93za0RVbx4EOyTuUqZI9xBwdNJceoctQA+MlsY190qVL/QzA5OcV480vv/Ga4
tjQYNirOMDBhzb3rc1t8TCP0LNo2nkrd00g5lh5IjTwhyqdc7+7VkGOm1k/Eh+afP2XsfWXHxhcX
gDTahYsLVBoeBeekkhAHZaK3YoFQP83WfaR1ivtEMPpGOyT2Gh7WvsO8gSNbGeIOuiG2CdqOMecB
/aY81zqij9r9gTOj7vmtEQntJ5ih1QQSlOr3TodM++iW1tiNcEXJhu7CmyLWwJONCMbTxfbFPb9d
nYKMhWN/bkgQwI1wxIcjolc0zeQpOMvVV9hmlUWITQZsaWuV3T/+SAUTc/a0PON1rPwfjXEYyj6c
081M6q0CrBsGHv6xOMnrGZH7VLji/Z9me034DNIIbn4NKPTpmv+pwQiLZ+K3gSeEi/BYP1SmEGOj
B480Vit159S5DDW2PPsmKy6yeVi3+RLSiycjUN1MvQD67R4w1U+uk8EjGeus3RH3LKAWhLflwHnt
1I8igkywfvvnpLS/sNkRVmF3e9rgw17IKpkNWCKPI4GL+UadNBeVz89wE2l2X00SCFPQ4HKkrOkE
Xi2L4cO91pxSK66cEGbfT3qoeud2SneteDfkNAY9fWe/WRGjGlgdAtf8aX5glN8XOpEfCAqLVWHR
tqEIT8ja38rc7+MXZZckEpGQXtcbWoy64dmCxPKwWHvJDRq7KdpgrCicHr16dp65wo0Yj8cSOBwA
d5eYsexjFs2cBsldEW1kw9n7djyaLe9gBd/dy5+a9QOyNqP3d3dwIuMHjMWY3z7ZmwhDjZG8P2Gf
2LoYhE1Z73CmfhZIIq22xI+isDOKOt0kD4drl/paDK7cA5t+k167bHaIIMChcaee938zEt1MH73+
Cf/zNn1yo842vRlc6AgAsOBSsTkuw8C4I2vKxhTNEgeGZAzR36d8AXYBL3vT6ZxXxciRhwvRxGDV
4GebBsQvPtqofoU37abhNCoFYWAfvU/Zm4+ikvAiU0bg9TF88Uc8RMMoLlwiGggcaPwOON98gQR8
zU/pj9raabjH0Br7Q7QP1eI90Nv6lvUO1Tk+AX6wYljPzS2VGvWfRAYGI8thvnLEaNICGFdlG9TH
sBIJL7L1FbDxqmQN4Er1vCCqNRdcIOWau98MsRk8aLuzeKuKovWVtj+sPOqrJ04mNXg3PrSoURTu
RTAWcuu9QzLoSWbUYP+U6s0sre3JHjoFUDgIpi4meqhbtjmvov4gjDz85+xAdGx18/g2A1AEBNoh
0nzT1Yl9ADTIAbdHAnx+CHi1GWjogJq2z3fsJsX4r8X+9JMkd47Qd/l2ZUFyCHhrNzKRxbWBBRTa
wD9WeZR1Ajplwp7+3VvEfdw07OooMEJ9oS9KUYX9E9hrqk/7wlX56Y9w5ohPtOCdSdnoY4kTYQBb
QWp/FcqTA2JUYSRMJlb3xi1mRIS/ADBtyVxJ2gLawrHkzQXnbSjSNac/EAeK8qwAVqvY6UTIrZxV
cqh+h3tnSSp5cZ265zT1wX6HXLBTo8TZ30dfXZID1urlvKKa3HKy4NNfVsiQJkTY79zRyWwBOCpB
P+3/p37LvCRq/qC6ITRE/V4nL3g5yxab6tDqG6PaxAjbPbJb0yvYc+bqc9Rx8fihwiwvxWSqMdsC
3L+Ts0BnFL2z91xuwHgg7HYnqnXpaPoWX+VtzU9D8YdMxFTnJES46fpQRssYhPgPto6wq68kmcZe
dwBtfOTpdw5vjQbC3+4iId4g1RM5DwXxm2SbOKQLmr8RJPxZ5Us2dEvdox7G79cymEUQWDtloDZp
L3sYFQ7AUb/J9VAqR+c+4A8XDtakhgDLsdLmLYC0tHiCeKMn+/BPA3HVEFHbgaZQ5zDZMn+lKXIn
BVfT/l9V4yY7qg/psLjoeNj6Wt9D8eDE1zYQovsoHQxQLQC0D9DdDFuaqZOSylcpAHd7Uu/7YmQ2
m5Lq4TgBSSxvAFhjoe4s5OKSc5ks9o6iiJLWu+d/l4zKH1+M3Nuj9PPC7vGLd54/qoGBl2KtINix
SDXzwu2LoeGwxrjVhr1lLle22RgWvvu5vGJEoEflkhCsZ/Cqoxre5LlGFTaE3MT9ipfI5k3JLOVw
qftSYIwuhwOCRsHtXp9LgyPjIeMb6mCDwRj4o2wa4CkZ+FuhKhIFpILmZ3MDpetuGEw3PWeVsR9S
oobPjTfS4hEkXnQiU/vdvtG880LpljYxn31N4tm5/1e1D8RWxGzYbkJfuLhlBwSubdpC4uGQ6XqT
CSsLiXOd1rGzj6u85LW/1b7NKkFIsjQm+k7M6NJgbenLcr811owRrWXI1IR3YS6HF2PBM1pQ+Drx
bgUiO/uGMN/PpJkdktc9/O5+dbdnqSqWnOeAGXdZRCEi+wTXc0EJiqSZCUWYPQhPu++DbU0xF0fo
TpOaQ429/KFCM+zRxkXFuZbyumNmtI6oRKgnQPo6j2c0VnwZyCno5ZminUUthqFO2somje3fvlgu
TZs1dgQZpiLQbgsjQrbvzUFHd5w//uxGTUGRIJen6AjLpka5dRLWSrv1tdjwDpfY/KwGEgDyopVE
nGwN9SRlYJjdCCQLpEr7vkMAUY/vl8D2cvFkYOUwnWkMPlcBBWS8y3Cf1A6iSCXxrM2SV8ZKGcy+
lEHm/G66dLaaZnwZmXatvWVCgVDGvBgaPCLBADJzyJYJHTqQGN4CsUHrSqFKnlaXjoa5PYZUjsCI
j9nen0oMcycZH8FgllfNt8iHwk5Ujysbfm5dm8M20Ly4ptNyrapmT91Zma5bTRd5sogxIJMzLoqM
C//mZt/RRY+cGu0IqTzpTGZ5EDbJpJPXVxfzJXVwh2+7ESEBdgZ+eE+cITo0JlPn8WtZFSHLwt+X
umfhkA/GhVcEg8WzlRqH0XtHP+sQrQwhvwQRY0FFWY9AW7VeIqn5TZguOM8KqiJauWpUv3jTcYgg
//B2cfkyl1IIKY813nA+PZvSMsykkOj8naHoOL19HiZqjiKf1nxie6BfYs6igyivKpXJHJlQWPPd
+p28u34cOSS6F0Z6CJvlI2oEY9d6iUQsuSi3S3vcOe2uf7A1VzHtNSVLcvdAPDOfh+OKZx4VSYqF
qRoBMbXISAnSCzKLRsxTXX2202xafD4X5wd7n/Kjm25UJTGeSd+CGK/50QnJUl0YuDM5tKY/yXt6
TmQnLXu8chtF0WVue7Jlv9Z6LsXRBp7M5FIqCLDQi+poA82O4o99xJAS1GdGPCMrrETlh8aPN8iB
1aVkeQ1KDE+ogcGKUifR55CFpddCXuyegY908zwRuxPu35z2IfMx6JfsZjus24A0J/RKsO1VCUVI
S98NmL2ttYK2c5SkHAOm/BLErFltSJizUVJFNdQZerR2mVrCRFALdDj2WGoZn+TB4mvcOf7fCEgF
K2HGwprvvgj6ShleQD3kufnzeapBixoEiqWT5bZvjEVyyS7dCg7Pz1qUo6BDZhN6qc4r4/5tX8qr
qHLcaBCPG4Li6YsBfO69jPXH3xwZQieTpn44cDEyTAsd+jK1J+TWIA==
`protect end_protected
