��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$Rx�y�<��wA�*;�x���@�̦�W�X�fa�M-$u����n~�%���P�$��W��kYَ���P7�?UMfT��q�6�U��k�>����~�\N�(�����X�e���/6U|)�X2pF�]$h���d.���9E�	�IN�f"�\��e�z�y�b�����Oo2�?�qˁ'�͜k-�K�P|����y:����3�l�d���bl��ˢ_�d���kx�rq�mh�MذM�`aS�.�DW�mS�9���Y��+�>��!��!�T�uOB���,��\L�7m�O��W���6����'���j)n_�I����2:��$�K�2�Sʫ��l ��!���{�l����.�j4�	��很�̢=�����N��s���s5���_�R�>����ТP .W;������	�"�מԫ�����]�#7@O+?�⡾�Ԫ���e�O�\A�	�ͼ���ƹ�d�	@�nQ˰��E؁Bf���|D_�%au�-�'���w�*%��"AM$w�*�!��os���͞X���'C����n����.���Xga���㔿�:����6g�4�7]Bt�4���4/f��A�8��L�Ӑc�T��)A�����ӖA���L���5U��v9�^�*��.�%�H�j�X��<&T��=M�+�>N��qo�*�6!7���,s♴��~p�A�/�����K�^���N�J%+m�2N`�F�$��-��;�:ETK��/������r6�V�J��B4P���؞FI��I]LI0p���5�1x^s��*\�vE2�}��7%����P�ck�c����j��[K�#�9�Ғ��C��t��p��9C���'��a�JF�Y���n&��C0��D�j��L�>s�|<,��@�oL��W��(ȗJE$�*�%|s1G=P�cL��9ȫ=p�h��("���D<^����>�Be�+g���ZV'xY�^�//8�o�� �L�H�=�e�Omf�r�	l|�iS��*�B[�p o��Z�tf;3��?(�b��6�U3߅xH�pÁc�Y-0��փ�$��mX�~�AD�+P$D�x&�Ph�˭�f[�^����o��L+јV�a����5U����X�t����TP�Si��U!vg�ɔ�V����)Of����o%V=���'�Y�8��Q���﮴��8�//��:C��Z�p!��� �i��\�g]��e܂'�w��OyÕn9���up�_�Qsn71�vT>Y�������գ�Q�uQY���|�E0���趟ͼ��M0��9�Bc��\h�_ ԯx�;4^�U��{��l��|����4xtc4o�=�M��F��ywT�]M3-J�*��!�N??I��_���S�E��\�z��	�Ȍ�� ���Fk����W| �z���`��5f�͚=0&��)B��!ԕ��?�� $�y]z��y�x���Sӿ-�̟��<&�t|ڈ�xJ/�m��>��2�L%�B3�~�?k,u>=�$2ۆ;7f�t�`ߠ����cU�&�ٚ3΃�3�,C�x��ϯ7TIɏ�?Q菨�L��[f*��M��l�`/P�)WI�"	@m(*6�����A|_Z9�W�Hn���1�DW�7�`4�5���qȋ-e�2�⹭�śi�b�$������| ����acSD�.9� ��gk�Ϻ��p��E�&�b,��-�6��'��щ^4�k�E��P��yS7F,��k�}D��u�x�s|$~��+��Wb��3���H)�0��H��U(����:=�@qR�<X�T�^?l�-å ���q�)��E�d��8��5~nz�H(p��:V����+joE=�n�s�Ĥ���$JY�
梍�!��](�wQ�?�L�K�_�\��ӗA�@ͨ��Ы�.�b+�ٻ9*m.~g�k�R�9\�y/�ZK��qT���ϲr�7[tA���C��[8�t��̡{ϟ�X[���x{ y��R�.���J&J̏��"(h�`����h��q��=p9�k2����J=�aBj"@a��w��m�|w��Z��7�d����_�3��\V���.��7���>�b <'�]�,��t�k�~����:��:!��+'������Su܈n��B3�1%�Mͮ妣ªQ�3�0h6��T���%\H�?��ސs�Y��'r�E'z|��qv��ᬯe��+RXU��PӔ���8P�ŭq�/ӣ��Y�߀2�eT�R����̚��]�`�ʳ�TK�>��.�q}�(����-k�X���1ҿ�NR��dȼ��2��p_Oo�_Fdk������L�el�6�߯.D[��աdB���NĐ	���m����$��ș(�LA��P+���!�IK�[��Ԥŕ�>*`�=���&]�,D��/Y��*f/�
{�s�|��t[9�E����Y�e��J �b��$<��%I�,m��J�4c���������
짺Z�{U�j3�X$٫�)Nά��e��*�iFE�/�8�\�{�qݘ=e����0BR��p��	��W��!}׿�K��d��Op�����B��w�����7��LX�ˍz��_t ����� �G7�ď+�:�uC ���{��V�~�{`t J�n�_��w�q;~e����n���SyY�h�	P�K��Y�""��:�����v�{���[S��i�q8�������`��X�uD�a��j5q*��J�A$4�����ے��C�{ى�wXFqOn����4�e#�B���HjdA����$�|��h��U�0*���1I��2d�;��)1�9�	���N��M�$�+�)�ǈEs>�Ra"~���*ik]���Jk��p ���0&����Զ�x}r�VG'��u�}���n�I)&@\�E/e��QTe�Q��R/:&�g]1�>��٢'%u&��M�'l9ņEZP��;xq�,u��{ �H��o7;����55=f�c�LH�r��Na��a;S��O�^�7I��W��X�轔" �p����8_�p�����)�����_���[i�B�\��]���f� ��l�2ߤ|ϔx�c�`˧C��y��f#.%��/L|��:��<��Ef�,��wr-���Vԝ�>YE��zӁULJ�U"e��YI���X�[�/�ӣi|q�[f'���]C�׺
���T����9M�F���JD�h ���s�<�%3%����G�t�d,M�y�&:�M�2���rB�Yk��vB��`|�ط&AS�W:{���G|�����NM��kH�WX��E�����ŕ�AZ�E���)n�a�4h��ի�O���}$!�OFu�"7���������P����%�X0��{PIutْp�j�߉:�X��P8���TAM�#��vve�U����F�lZ������Z�ʁ��ݾxp�8Yg�3�-�9n�3P�?-� ū9[v���	�i!�v�,(U� ���b` �M��q5�_�P������ e�0�VxX�����T�4�O�������j�E��_��ue�EX�A����ڶ){,oL�j�q�����x$A�<���w�`<��`����~_����>ޏ�mP�p��#��R��g1_�����(���� C�<L����S�M�	Y⽬L�ó�3����&G��jv�����mYn=�7��Z�j�[.if�l�[r=�����z=x����^���NdP/c�?��F	>�cO+����@��{ ��iZ�L����]8JƎ~�����s�Jr���EW�x9�G�cw6�J��Vn�-�߶z�\J,
�OwhG6}`t��ሊ6�z�ěL�+�u.�l��W+��/��y�#3�O������Y��?����J�z�&(��JA#V���/o#[٠4'C�C�����c͔�h8��q�\�8A:�hg_�[�#Iv��+Z�p��$��,�т���-�Ty8b�����m���5��=4#ZٹW�B ��V���}�50�*�;�w�~ O���#/� wa��4��o�572���b_b��59&Q�V<d��9ȳ�5��3��/���-���]y�kOta=H�'t-��p8�?�9SV�m$s_�Rܾ�?<�8��R��=�Q��O�������0�gI�h�T\�U$OVw��&�]���ސ����߻��  ?�o���6��|\'�/�j�����kv=�O��Wa�^G��_]Z����D�� E����n�c�Z�g����H�f�Y�g�pnT���R��hWZ65)Dp��JS$d2��c�R�l}&�+��8Cӌ�i���!�Dg�A�hBs
ɩ�H���bHS��"gy<̐���
�]+�p;��ٺɅ���Bg�L��i���L �].��S���LĔ�����tdK\��A�����#��F����	�"T	g����]W�BY�tx==��:C3����])��=�#��5���TD��_�/����]ɼ��7bj�	Ռ�z��̗�8n��x��Lo#��=>hRa�r|P5�¥(��e���Xz��4�5w5�E=ju����h�}j��]��A�ڜ=�G�_� ���|�2��E,����N�(˙��]9�X��X�/bg~[�{�-�z���x�8[q9Flfs��o�`��)�=����"Cd�S��T<?ʵڅ��H#8����)sK��� o��w� ~Ή8p�q]����v[�ksg,k""�0�VaRQ{`��-r{���9����GҤ��c� �gK��K ��ϲr{�FX2^i�\3ۤ;AwB��ӛ	i.\��N)рt��4��P���!U2�8�}�J5hyIxq��"��G��5�C���\&s�꒷D�I`�L�I�.��"�����{`�ym�
�� ��숨�.�c�u�x'�����
�I��ͽ�E��z�����)�@"i)�`^F;����-zI�{�QЈMv�I�IW)���bqUKJ�,�H:�����64CL��f��n��O"V�Ե(�0U@s�ҟ]Q�Ԛ��]���~v*��@J��ʀH�2�FJW)a6����]��#A�p鳯ɹ��Pa>�ʜ��!�L \b�96���o1�����ϑ�$��#�r���P��c��!�,�<���cpC�uND]���M,��.�%�))�(3�x+���?�d"ߘU�¶��XJD��O�ي>xS�͚0թ��Ӹk�����3O�s�0\#���jz�� -�M�Kp�X�~Zĉ�x�$�A��X���-u�ҁ6'q*M��՗�<�yd�b�Z���f���K
e@ㆽ��S(e�A���D1��h+�w��ٓ�4�n9��I�V�V���H�a���a�y?�>��8"\]�9�N�e���*�yَP��(Lۿ����";�����^o����kKv�Q5�u��
�JU��;��)K���
A!��{�Y{�]H\�֪�-'���Թ �2h�XH��_���-�0���!��5��r��k>�6�MiU���~����C�vBu:L�����g��u���N�ǹH���A	�A=�m�fċ�n.���L��p7�o��Ƞ�����^66�p����E��� l�������v�i �@,���0U�mk(]�$@][�WD�M$Eg�5J��:���ҋ3�ǌ��AQ����sY����u�p��_6uW��)��i�&�)NԒ�
���y2_�	��z�K�6�xl��w���M�1&������ (*��F�Q�Ա�	�J�Md@c��6GI��!��&�N��~'�����Y>�V�;͗Q�|���w�/3f`�iO����4 H�8�RA���@^�=g��^x �ET��ҳ�����rK������w��N눺�ȴ`b\Px��	�yBw�����N��	m⼗1O�*x�.������dqGK��(t7R����?����q�lb��q0n8l�j�V�� ���ɟS�<���/S��y����U=�2����||4m'���߱�B��c��~Þ��F��$9z!�o��y�3Z�2?_���4�ׄr8�`s�Ϳ�-FH��~�X��2�i����Y;�����F������_/X�7^WB� W��X��P�UD^݂�����F�m��`�� �b����Z��*9L���;0�������!����Tu�
7#�uٌ��a�+P�0�� �"�j0X�v�D~�z߄]2�P����'�꽒:�a��H�dfl7kL$���0!>������)q��j�)Y�%	�D��X�ƈ����q>`�Xj�"!�҃ `�9Pi*��x�㇅ߛ��� �v�O4��H�~!'mjM֛�}V���\� :�F3�|���� �j߷`�5ui*�B�=�{�Es�`{E)V������}�,rb��J�@e�4���~�8d'+���iq)>q+W�8�W�2sU���&�i�.}S�N�-bA�ޮ/SQ�؆W����6�[!;�qTqQ�d��[�s��}oB��v�C�� ۜo�|e�+��?�\Y������V:e�M�
rr�#�i_�,M^|l~��/i��d�8D��l��ï�X`�^{��W��q�WYo�Kݩp����#�X��0�Y����m��p)��{	l9�;2 ��*�ê�����7��F��cE[�mt!C8{R���� ������j/K�L ��`�*�z�O��W�����j[�������٠�4ўyAK�_�#L"X��_��c��
0潊���M�n�:p��6[�Zu2Q`b���dX�0�jl���[)�7tN��<�N���Zu��_���`��p�9bA��M�E�Ɋ�� �K�$PQ���Gr�I�" �"�V*�1Pg�s(���F��?�kk�;s1�
�)�]��u "<�@��V�T���V��HX�m9p��M��V���0Pз���l,n=����|�Ej�`�/x�{��n��v�^�����t��2��2^p�����L�"�n����-vW�y�H@ų>a1,g�0j��ۀ���`�2�J�Ј)<�������<!S
ⱛe��S�o�)Z��\�j�5S헼(;�B�R4qO���('!I��D�jM�N�P�]+T��'��C]�hMmY�����-�����b�z(��Ib��.H��G� 7T���*�|\����{��
X,$d}*�U�)��,a	t9�Q��n�Yo�S#Tb�X���	 ��9�X5�R ~��ܳ���V`y�N�ν)ղB��.F�Q�)����PA5w�W-\`GW�s"� ������-���L;�:�dU����Ub����=f`�����i�D��vDё�,١OJ�+V����}u�ܹk���q]��"sڡ�>�[GS"����?}F��"����Y��AKm���D��$K�r�k�-zw��p���$���}>� Z<�n�� �!��`:Fs���!�}%�Q80.0��\��� �fI��[�E��A$b<:�H^��d?ĉ�K���%|��C0C���j��y-+�	PO9�N�α��:�ad �;�"L��o��:n.T����M�����.��yh��^�|�2���|��p\
i����z�
�Z�'O�PI�� u����C8ƦX.+�1��l
�������`��(2��b҆µJ�Y����o@]��ڸ�C����'�+.
�Wf%�rf�[`�YGI�*�������L%E�ٔ���O(�N�*,p V��J5�v��rј������?�W�-t��pn��(M�����O��Ю_�1E,A3͹��D�z���*�m�)s�)>�6���5����ϱ����1�:`�?���E4r�9�̏@/�\�$��HCu��Z<������� ���SY�7��QrzylU��Ph��A�����D�j��A���u��.3i����Kc��qƳ(��d)St$�{��}�C���Y_���X��$��u�:ޥˉ�a��C=מ��G��Fd�H�Pw���.���m�a�&�9��Q���+���8�3��xٛ[�����z����3���>bP�;b?��`� #�C�'p��*Z;-�(L	r�G�/�c���<O K�7^�YԳP��E-�"~^��*e����4�H7$_�n}tNv'!������������)�UyS*�������tF�8��p ���dh:e���Z�q�,��ҳ6�z�ܛ�&� ��K�������P�����"�U��1���/_��Q�~shkh��g��	��QK�fE�d�q+�Fm&K���7�h�n6wpM�l�Eѣ-���*��i7�Ev�L�C�̔3����L�R�e։��n� =�xk ��:91��Лz��A���Ѷ�`3l&�h��(!:*����~\����;��?��%��J��IS�;HZ0s?�D�G)��iZt͈���Yh�����4c� ��9���*�*k�;)"X�TB��wyL�uC~���ؑ�FWE�K��㸔ƪ�΄�ĥ$J-W�DFó+���Hz]�H�WS⹄��jx6�a�{���}i��VA��>��sK�mUuX$F�7�N����=l�`y����O�")@,�z/w�O�#��:�)��Yj��g]�脾�.q�]&������^�����hpκ�y�1�9l�1�f��"b;�C-3��>$�S ��(.�O`WlS�n�j_rgF���y�O2eܸ�]9e�Rӑ��n������&��Zm�vl�Hi�8��)�r?WmY�����Z�3�)*`Q�ʤ�;f�Mإ��� �!{���N~[���=�k�^���t�ɾgXv����1��!Z�B��T��m��ɤ{N�|Ɲ���W�9�|���[b�+a�4���{=�]��ߧ�9
z�\�7Ę�U4���&J�C�[��PIBJ��Q8�Z���\]H�He빔B���D�j~��A����p��2LI��Uw��/���R���j[N<�9�l��Q����