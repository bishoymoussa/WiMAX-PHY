��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$Rx�y�<��wA�*;�x���@�̦�W�X�fa�M-$u����n~�%���P�$��W��kYَ���P7�?UMfT��q�6�U��k�>����~�\N�(�����X�e���/6U|)�X2pF�]$h���d.���9E�	�IN�f"�\��e�z�y�b�����Oo2�?�qˁ'�͜k-�K�P|����y:����3�l�d���bl��ˢ_�d���kx�rq�mh�MذM�`aS�.�DW�mS�9���Y��+�>��!��!�T�uOB���,��\L�7m�O��W���6����'���j)n_�I����2:��$�K�2�Sʫ��l ��!���{�l����.�j4�	��很�̢=�����N��s���s5���_�R�>����ТP .W;������	�"�מԫ�����]�#7@O+?�⡾�Ԫ���e�O�\A�	�ͼ���ƹ�d�	@�nQ˰��E؁Bf���|D_�%au�-�'���w�*%��"AM$w�*�!��os��X�{�lPǳ���ѫ;����K���V��@r�b�f�4I���Xg}���*����I?����c�,w	�1M6�e20LkE ���y@���j�2ɵ 2���3Q��WQm!�2.(4��z��g��R#9j���4:n���}��Xx��ZX�,��W.�sY����k����.�]r���0j���c��F������bPX�z�_3i�YN�; ��g�~6��Y��{`��A�Ueੂ�u��H�oVy���n��-7kޯ�-^�_��3<UmF>}"��Q��W���?�i5��Z3�E���,}����b��>��K�G�}~��d���U��l��1-B��2�.�H+I�Z�� �K�~�����7�iįщT0�g���nƀ�U�		�WU�b[Ɋ(��D���][���J#*�˪�>�0Ԁ!��0!�'�Pu���5���j�ێO8�&M�ob9����7NXJS5��g&Y���ְx����d�4:��i���d�Hwǖ���ݠ��Y��:!($�ц�H��� +�A:ܜ$�9o��MD�Uz|�����L�Tvu_�]��qo7�M�V�����V	J�����tg�Я���%�֘F4 z�Y��,����E������ֆ�w(�8�Õj��������i�h�����nq���%�\��n���lX��k<r�am��B���bTh�>-��{���[�7P����~�Q��H�)���"��/�g���$�q����6Mq%r���)�|���f�G��5O�=@Rݻ;k��x
Q�N=��.�g�Rn-�d���W�'�TԾk����)Ɲ���yM��$�	�C��LC*1��r�A[\�Z8�/��Û&����1J#v��~�4�������t9.7+��Z�]��6e#^��)�}9�`#z[��T�1���j�.����\{�����CI3�$��H�|3��[EL8{�'P�P��>ѓ9{�������x-�Dk�N�
F���e����7<5Y^�-:�Q��^pۏ�@1y �Ku��'"��� ���|jr�� M���^q���D��H�q�J��a��p����T�]ҲƐvXS�^,ڏH�P=�R�P��vr���JUn�OLJ��=F��@�b��eٶ��u��E��bQ#�` ֗��刓�u%%�h�����ד?�I�� z��?���z����A��ǍC/�����y�P�IнOȒ�Rx�S��I\"���19\jߎ`�	 ��U���)����(�;f��uJ�t���1*���r�`���5���y�Б�Ņc�č�H+iJ��D�Z�%����>���� VVg�,��1*�K%I�e>����N��WV2 �. 9үa0���]�X~I؁��(p��9�w��9���m�1�xxe��H�����SJ�g<A�.���YR���ss��Ў�cLS��d�jl� �¹�aYV{r��鎈��[�'K�s4�Z���,7�&�!��.��sM��S�s��\v���I���ֲ{Vi��"F�l?�Ed�^&�����iS�O�b�l�R'J���Ob	2X'"�:��>��I������ys�[
<��R9��H�q��Ľ�,57�E����?��6
�ZX�#�\j2���y��lq�˞2�@�f�۠׈?�	�Ǘ�F�9���_q�Q#.z���t��8���u<�mI���(�ЙY����2z���X��ł�_��nj��	� �1j}���uX6=}�qX�8}VL�o���eV7�N��f�K|�zM �'׿g�~�c��X���W�x!``��e����Qt����A{���W�x:�����PG�G�l̅�X���P��OF�;�@f���w?ǟiV8���o(f���1�!��Ӻǘ���c���:�]����m� Fl�V�5A��!˶�CoI�&����P�Z��X�9��b��B��H��Hs'�P�\� �(Et�^����k^FCJ�q���]��P��m�`c�%�X)Y�����]��zbcdIY�w�!���ɝM�e����}|yy�H�hoȇ@pT���҆e�W���g1���iw�ʾf���GHG��2��^���n��\�g���-�Γ�"C{��'�:���%�����n X�d�h��ӭ&)��MJ;Cw�7�{4������zTv�ޤeW�V0:԰�=�G
���h"�O7�ˆ�esԳ��i`v�9�^m���eq皅��m�
�HZ�rp�x�����H�n�H�[n�:���
V��,��DFEرt5��(�o7�K�;�R�>���u��&3r���PJ����-���{B����@4���=�,��U����0�`�9����̩a��i-��kji��7p���=���D����p��~���X�/���*Y���
}iI��>-V/('��B�WGtl5oc2,��n�|l8�������Y���D�{벰�~��F���<�SMԵ���[25uT���ܚ���"��6�w�p�;n2��s��V7RuyP�8R���5���]�O�-	x2�R�!ÜV��9uJ�ӗ�;=�M���*��
ħ����9� x6�z�dFg���]��r�����w��#�M�myK���G��ID`8[�?�Zg�pt��.V�)���$9��1օ����_�h��ů����叀3'�G}��[Yi�(���^�����Љ!}i
� �x�kuI��2ɾj������vO+n��Jn��@O��_U��N�Gz�d'���u�Z�H}�#M����U���(
/i(� �v�r��E�gv�YG�:2���Y=�EQ�	���lj�V�������xDC������:58�*+�;	�3F5%
YK��E\kpVG� d��;\�߉���Ħ���~e�`��ڕqx�2���1q�&��2Za���E��u�MGB��&��s��i�ZG���v1�.g �<"5ҙ��o���Y��yj3��A��x�+Ꮰ���/��褾�V�F:�l���@����*`��3�}
P��|Y#�!�8����Ҿ���2��)�zl�X���r�VpnB�8H@�$�>=��T�P �t��"ϵk%���Z�z[p���������ѥOb����R׷%#׃|J����������)ޫ��C��,����9��0��NP�P��>�Yl�+w�G;VFǋ��&���n/��U����!�}���p��4�U	��3��r�ܚT�\ڌ�z�&s�}dM_�m���܏����/`+,�3>��P����� �^]�:.�~�OUvN�{ƈ��7�9q-{T��\J�V$���P�	W�7W2�ns�g�]?`v�:7�p2��I:8ѱ����.M`�Jm@�]y���U�/��sRq
�h�x1�+s_�p
�"���J�oy(�wB�ǀ{��ϡc36�/
�a���k��ۓ4�. L��Um���1��G���,�k��Ҋ
r�՝��c����L�o�M�쿝pd�f���9 G�ݒ��M�QW]�I �V�*���('T�4�r����
�/S^N�/�9ݎ���Pg�+�2�'_�y�}"�!�Zq��;�Xs�|�����9B���>>o��� ���N|ӉZׇ���^l߂	��4�#��o5�R��R1o@�z�5��xs�\%8�>`9vm����с+O����E4W��u��J�ӕ�9?�M���ӳ�-����z��A+I����x����w�u1%�©�9	1����oWq�/��''�Q��~qj���
G�Q�k�orq��e>��9��\�%��(е�䋤/}�Sd#""�ӟ��
�VՅf���2�6�G�ŵތ��䜝V���X�I�˟��us�W*.Q�x0�i#�Ձ�DSA GW�@�qT�iV��g��L�V3?�a��r��1cč���H+�޻���WJ��}�f>�'�pXw���A~5a�c�Y�:"N4m,��l�'(m[��	'��HGb� L����Sւ<>՗�c�}KH�W�A�tM�(���?G�B��@�����"����qalSߺ���7^�i��\�e�,\�t��?^wN�4*�Yh��8t�İ-��9��[v���-"��od�
y�5���VGc|f�P1�_€�D�����ݰ��E�	:g1���Q�t�p%��sXuw�E�<�5�f���!���v�Uw�!<o����_'P{6u��8����f��LG��^O}�m�>�VgXq�xX2�[o���5t�{b��a��O�G��Xū%E����ng6�V�ͨ%[��|�b����t�ܓ�a��ܸ�\_�|�&/�!-PsZ�+�^	���'2qG�������x��*Ҭ?m���f�(�Gci�B�ښ�O��Lz+P��I���aY�a����޸����Ծϒ8GZ���)�%N�h׉H��#G���F�#,���C>.|���0F"H�������j��$$lB�X�6<�:�R[�f(��$��)h��\)-E�u|������Z'��b�Ϭ{��s����o|��i17�ay���u�!MT�8���A����vSz*�~غ��j�[b�{#�iy�"��Ha8o�ң�k��X�C���(\��h~�ff\xM�)��Q��~hC6�Ֆ4����kE\��ˌ�JT��_e����t��������T1wGؼN:�K�_3��(�L�G�gwMh����6��Uzi�T��w޵׸�<7l)�*��+�Xd�4R���R ��0�^F�����D�	�n�e�kG��9���I��j&�*@��է_j+\��MC�����0Tw�:Md�(��+�5,^��=,7�T�������m��Dt�{�2�0˝��ÒF5���1�H ��Fd;@��������8v8��A�9���w;���C�-Gܬ�Tjob�
A!�r�wl8�.8�����S�r������i<��4#�谙cz�Q���a3�a@n�B^����t.�K�9�D�l��AX������iIߊ���I�2�{ B{I��3E)|������������l@�WwĚ��m�e%L�w#�۴Sn�����|�ݏ�D#U��DtF��>rZ�
I��u��^�F	{0�������;@9�KA��P��Htނ�#�P���|H��`�u�_�y��@��]\ז�P&�Fa<��B#4`���R,�����ZJ�y'�m*����
�bV
'�Q|)��ۚ�N��i�h��0�~n�|Z��W��hM|��ɀ�C���^�BV4��I����IY��W\����q�ecE�UJ��9�.y�Z�8������u�Qy:\��M~��\��>����K�︄�0�b��_�� ��
Z�w���`a��(<>��y���x���4D����:��%x_�l�a�ͭ�.�?j��f�Լ�X�K=�O�����������D�0�ɟ�]ݧ�+D��;�t��M�MK]:9`��ս� �*L��z��!Q	]��	@��Y�EO�D�6N�B`_K?��\��z��v5Q�P�;����X����pg�߫���O̖!'##�cg�����gvL>!-l�i�Il��*n)��/{$g��b�f���P|�x6]��tR�������;�$�o�!��h�l�w[�����W~��YZ�܏_u�5+yM1�k�j�&�=�G�:��Ѫ(�B�^ܞg��d���1 ���ڂn�'�𔁎Sx���/�0z��'/kax������P1+����56$�
T��הCrܚ�i�v|�i!�+����0<�3%X�1���k�0�����hF�Zn��,(.��vq���Zf��et��*-���S��1sCTY��<�Grl� ٖ ؆�mf�F[�@�����U�Ŝ��%��և[�Y*`�m+$$T��d�`yD��T$��_�O!
�$e6^���L��{	�9��׃�p����R��/O2���+�9�}z3�*F4�.�/�|nΓ���o��̉cr�儓Q�XtW �e|�ړ��L�J©��U5�Y�9�J�t�/��㯴�<����k֫2�O��d�բ�Ʉ�n�.��<P�M��x�{eR{�#Ġ5]z��cf�����l!!
���X�k�[�f���{|Ǚ���Ҟai��0���I�1% W��܏��2x�Ӯ�I;�h,:y'�\S=�X��u8ٯ�8��<�m��I�'ed����k@~zj��u�N��5(.G6��S�1da�8��*���+ 0ݽϡ�ͻ��/��*z�9r��&�r��foρ6}�J�19b���
���ѻ�b��vf��T�C�e����՝!V7�kW�s�����pzMf=���VDCh�>=�M'(�|mF������_ &��J�/qc�P��e����c��c����H��?����f�*�����,����� w5_�I�_�{v֧u4�$_-"z&���8'.)>eh��|�����Qt��\��yV<��9��Z���#�A�r!�:?'�y^�H���wm���;.s֕y���'��*5��|3&PVI�.��բ����`���T8������0���� rZ�i�W��M|U�CZ�Y�<����/�Dt��^��	[��VZ���d|L��9)k��> 0;Ԥ�)��C'��Y)�,,vv2]=�i���	q�"��o?\/��n(��4><.�zUP2��+�W��Kg�{u�C0�3m��n�?�!LXDd:��H�Z���o��������ɥ�7�&�g��h=�7Jl��Z�CnQ@ԙ��E(�s9h?�����R���F��5������R�Y/J�w��pU}�#�����(z�i�Sw6ݠ6�R9�L�Z����/=��~BM�7����,�UIƤ7<{��6��\�
^>;A������f��ۺh��E}�i&��F���J'˦O�v���e�Or&�Q?E�5�`v`��4Aag���)��>*mH�(�ʁ�ؠgސߏ>�)�E���$+�{MKf������U�c@B,4J���m@Y��	x�4�ݯv����V�T�f}4����pf�K��k�����2�G����?)?�~���Ub	�V���@
�n�Nj��b�k_ub(��� ��-��kh]�^�r:o]OT�pň����(�X��}b�Jvl!W����Uk���׽�3a^���\v��g8�/k��