��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$Rx�y�<��wA�*;�x���@�̦�W�X�fa�M-$u����n~�%���P�$��W��kYَ���P7�?UMfT��q�6�U��k�>����~�\N�(�����X�e���/6U|)�X2pF�]$h���d.���9E��WG��L�X"]�Ad����ľS���8od����e�GT?y	7�������ݵ�^��R�q^]�鍦�����s�ae���h��L��P_���ާ��YЭF���'\��68�b�[����w8�[X��V�F�0͘3����q諵�uW� �h�u\V�?@��_6G�_�*�G���B�絉�f������[�G��U&�����~�F��AׯK1�`c��[<��FY���4I� �#�G��x[X�=�Q1��`��R>(�w����R�O�?����7�,(�H\�#h(W�EH=�������yq��Ѿ��aF����:�U~m<|��.��0=�P/���4ǆ���T(������v��lvh�凩����=(D���P���W��x=$QfB��ʮ��:]�&�.��H��bG��K�a%��m���)WʡC�m��n�*U��Szo����D��/E�ق��:Sm����9z3 ����\�1r'Ѝ?<��خ��`�����A���O�$X@r�1�(F
2+ i#d'����J�,qR�/�w�����
����1��v�B]�8Y& s|v5_3Ie��]�]�LQ���f!�hH��֐7�U���al���©���j�Jwk[>0@����d�M�>M��8��ԛ� )A���wE̶ҽXgȻ���Uyj(�� ,6�+}Qwٗ���y�ХH>��i]WY�DIe��_v��kP���`˸�w։C�����@j��8w��Jpi\d�0[���|�ᔽ$=h΋�B���$R����@��G��5�c�0��,L�6�@/�<��;7�j��Ԃ!va���'����꽞�f�w��u�Eq�s/��$B�����f���!C�H`��su�ሟ���}�f�́�5z����d���5�f��L�w����""��$����-��.ˣÓ�)�ұ��1��{ޯ���$���q�Kp��o�J�.�-Q�b�^^.Ş͗j�"mc����mh4&�'%�9 �)��ң�pԅsU�*51%��0�*�޼�� ���ef;�ph`ǨHC�����%�8]d�[Q��<��T�U�w�D;�߾����{���P��.�u��o'ok �
A�4�s��GE�$�#^^u�P,QS��<����[��|�Ex�n3�o�m� ��O�r)�>�?�E�B�P�<G��q M���Q2��Oi�o���]�v6�?��Hv�ީ�0�VjkwGR\���� 7V`pPq�鶿!ꤖM�N�g����2�d�)%�-M	��{��`KG2P�d���8H�#�n𾹥D~iu�E�R�e����Aq@���կ�Ӵ憐�ڱ����%L�W\O��8��S��iϱ!����	��C����C��ө=��T�����ˈ����Ѥ3��Я��N�820���������}�o�ܪ��ͳ%l�tx��U2_�qv�貐F�4T�T�`��;$�s���]�=HJn۹�˿���^��@���%ς�YPj.��Q�:��yw�km��wT����O��$��g��1��� 8#3*�D�>�@�z0;؊�Ag|��?��7{���{-�؃��q��n��g�@ �LH�����8^�]�Wh�G�� ��79^��M��_-w���S�4�R��nf����8X�����!��^��:��(����Y��ҙLY��jx��fU�~���k P/�D<ƽ}��G�/�V��_���(T{b(=pt�1��NHle��� �����Z�ч�=�4k�iǝ���yw���9�1�}oe'Skȃ۔t�����H8-��{Ŏc��'�ˤ��������&޸&�Mm�Grܨ�yI��g�8.��Ҩ�#�^ڇ��+$W'H�񈬎�Y�ԢnxI�ht9�a'xlY{�_�hK�V�]�$8�i�1�&T�GW \]i_f�� �w���c�k��P��:PR��{%��fP#lȏ�Qb�_c`�vݢX{l�ʺ#(�bV�/-
1�V�4�n�V��⊪�g���5�'w`�R,�a�r�g��r��t��Qؤ,����K��Ac�2/�k:MȗǴ����Qd����D6�&iWv>�?kѰ��9�y�>R��K�����/������}pE���*\�N-�}W���)Z���<��	q��
>��RNG#k�r��|{�������m��������;�E�	/�ɷ�
��%�.A0鍔>�ʃ^1i�0�-eo`���S�E�����wg�{n�������i���7�vo�\(W&�qG{��H�O��Q�jY+���8ի�"d��7�3B�*��b��Mǟ��P������G,2�
s�͙K�p/��?�����`1
 ����,L�Tܴ$cT�7r�=Q�D�o!�|��ޒ�V�u�!��dR�[�s�E�.D�kp����%/<?o06��8n�Cȁ��K8W��4�����C,3�>�;���v:z\C��<�����.��(�N�E��p�Q`����(s�e�'���w��Z *����!=�B�9��T�S�,ݸׇ�����mU#��&�ݐS�9��b���o��J���<���#�"�Da6Ȁk��Ƀ@��2ݡ+��c 
l_������`9�(|k=�k(̈P�vǎ����R,;��RDx_�Gw�a��T���˷�љbC�)�pe�MJ���ɿ�b������G�(ܮ��$�ܬ���oǒ�{�ڗQ��B�Sؑ)%�ȃ�ԗ�B�J��i��=�Q���~s�Yu��S:e�mI��8F���
0y��f�靰4/6��aӥ�cZ�n2%�\iX6o�ᆐ�q�,5~N�x�	t��Qߵw\ht$
��,�ɳƜ�V|� jV���~3��kq�˵+F������>��@�
�(���k)�{��q0��t?!�H�H��I�6�^�B���h# ���^C �,�,�����_FR��.e�c�ϛl��i]ֹ���s2���������D*wQ�|c)S��?�]<����N�hB�5�iqX_��T,�َby�o�Y��k�W���bekk�Q}��!���FӮ�Qb�p��Y�2HxAm�z�dt"%���x
E(����Zh#�>�P���N�x�<�{`�eU�����. ��&���-�����*ٯ��	�r��F�mڰR��/ki3���1N[��.�)+�q�*R^T�n��n���;�j�.��U�Y��O�%��39�G�q�Z_;�<����C�2���<"r��tRU(��͂n�ÕpsR��E:׊�ő��;߾���v#�����0��� >1�%/Q�8�x�C[:�c��q��(�c�Ԧ��7���q���6gh��QJ����X�N��ŕ`X���bTkЭ���[Z&��x���7(�N�x+��:gܺJ�\BmE��4�,���n��0��ed�s�w���H �h��7:9G`��{}��`훽Wt	��0c����fg��&�q�>O��ӚqdOSN�+;�\p��w?b�#�IFE�I�Z��&�L��J<��zd�鵜�Z#�V��t��Hu,�"��OKe�6�':�
�X?���.p��7`!���%�v!ӑ��"��(m`�+r�G���t�sG+oGe�(d�p��uV�KqW���8�xY-@\��A��ښo��_/�C�%�㚻��ߪ}a�	�{&�������>��<z��_�@����L<�C�h:��es
�3a�]�T�NƑ
�x��UV���"0����?�l�|���_�fV䯇;N�/�ԫ�0&.͂+�� n'��4"+��L�u�����b�ݜ�~��	��fd����<�m3�|.¥@��:��������w��p����+}=�I!��
7Y6��������_���s�ٱp�Ҟ��z�h ��D&g��d�����gP�4君�A��qv���ޅ�^K�0�L�����Yl�-����0KֹI�QKg6"|--��8
��w�ig�.2q����OCW#6����ʀ�!^�K5N�A=v3zP2;0/	�ha`���Z�uZQ$H�`'�z�Nԑϣ��hUYJ�@Zwt@�E�>���yN�-יFb��4{�w ��]�建�Ń���_?_%���.�y��v��Ss�.�W�̶�Ӣ5�ǆT'���^%��oA-ޖ��D��z��0Ra���v���3�Q)�	��6��ͦ�O��j����BI��\�gۓ24���4�2&C#�Iӡ:M�mD!�&�J��⼜}���� ��>g���,���눃���*˜�L<��ٓw/Ͷp����B��	R�1A��!�}�#o%F��Pr���4��$Ds�]���*J%�4��c$��2a���|��wln" ��9E�Aׄ�.｢����p������Z��JTn��I胥+���{~a<�D:K��򗂨IEl��z}�4��_������lQZ jX� �����sH�;�yK����p(>N�x�x;�R��Ia�>�7��WGe����� 4���@��v����%/�s��� ���(Ub�����eTx�t����ۣ^��`�H��M'+!�{D(��J��֎Pb7P2��`����#�������b��seܑ�C��4�F���H����HF�BT�*2:*�*���a�XP�?�U���#��9��bbޚPV��J��~$Y��`�h������zS�{tmL@�^i�$�S(���dҭ0]��'�.��M����]���ۉ�7d��2F�8%?k���*�����=��7c�;g�H��|u]�<�I��b]V��TM�I��g�u-7n����ac>T�%T��8���O���3w+Қ��[?���@w?��m���зG�0HW���]+e7*V#w�����?R�w�mQGS���'9��-
zo�Fr Qά�@!���2����5H��)�>�7&M�O�f�C@���I�J��M
���xyJG�����[���@�Hz��E��t�c��"A�	�q6��S��KqG�uZ��Oڽ�f��=�x³O����W�*Abڸ?˳��S���g}U��^�4'>/����:�g.�z�tf��	L�>Ԩ��S��N���
�=��,��5���U������}�wO��N�������F��/Z��U�o�P1�ΒL$��-�Gw�T���|c��v�LX��r���[�ۮϤ��4ĭX)�-���d|��2����~7SwIi�t�kID�:�v,��ksXԶ���&��;�^��Th�ytq8M-�cb���n+���#u���o
`'��i1,i��̇���8��*Ѓ�bL\:T��=8u-OD=���__�:�?�(��{>�Ϡ�:�]�[�R`�}9S�,�� 3m:��lWe&�&���ܢj��2%6�OR3�-�B`uñ%�;^e�@��1�v�v	ӣ�]�7t��~�#z�S�Ҭ6��+yR���D`�����ŴcԺ���OAJ��a���Bb��K�"�Z�5}]Q��l{@E�Z�����1b�w�.�
��1���S��{��&�	�\�h�7�ۏٔ��"|�����b���R����ǲ�ᙘ�l"�(�Y|ģ���sF�2���?sg�KY�������.ٯ��Q��be�]KHz�JF�Q�NXA���R���	Q�w�ʅ�:��Yw��ő�}�LT	s�����>��S�|вD��P G��8���U��n�=�Zj.-;J�K��PA&�tp@c��R�-���ȟ�����޹��N��?G�T�=��1t<'1aO'����c)|7�8� ����g��H���{xSAHU����x	�|�X2�������r���	���U�N����y5<^rjo��s5R9q� d�n��>}yA��b�����"�p��	1�qg�c�9N� h���b�Fb{裰����<O�� �s�ݭ��1xq�����s)_��u�|�����y��~m%���r����3���8��R$]!�9<\ίI��v1��y�����=8�956����oY��G*I��{�>���W4�sY� ��ۨ�6����q5,D�	`�CW&3�w"r_b̙a�*��=]w��쭥������ݱ"0F�5��ɚ����kTKFEǪpE\:��q���H-�X���	�G	Z��:TxR5n��ҽ?m�����NВ??s�u��1��*�8�?^�����]��0�qKeo�i�l�<A��*���|@2�YB�v�[5w�nfax��lyX�{}C���BUg��ٔ�Ȟ�S�Y"H�Ϧ�m��\	G���g�W�rf5�.����m"�A��D�88/e`9�T�t�zP�� P��m�Ue�)5�2����@$2	�E�b ��#����0TF��>�q���W�	�)��o<|��Et����ܣ�ɽ�UVNw�Jp`��N���/�dt�u�(�
�����bO�߅�F��nX�%�,$oE�(���*�K�p3��~��vx��S��*��n�+~���@�cݚ|��/���1Q:i��X�r,��r���M�	�=�릐�~\r@>}��J��6���Sa&[ig�G��:��/���4`-AOT�^�59�Zރ�5!�F��:���>�^fREEL)9��0j\qxa#�cE�Y[5n�Ǧ�^+y�"����H5ր�fU�T�a`t��c`/V+.�]{�L���%IQg�q;|6/`6��6�	������v��1���V#��{ui\��X"�?��R�q�Ǔ>��갿�u9s`���6�q�	��,!�8��M���"�/(:�e(�@��;e�m5��[$X$q�0�5��
�'�T��z���Mץt>ۙ��t�`Kj�㧷]�b1z�����<z�G:��d�˅��z4�I9_3�2��Ia-04,�p&R��m"h��/B���*`���Ʋb`�j�5��#�o��9��"PF�t��FL��0�	��H0�]@���^$&�"KF���)7�g�$	��7x�Dkur*B�(bYF�~w�L�"�|h��k�vn-F5�b�t�)���q�Yh�u�*�4d�-.����&_�8>S��8�k�� Û��E�Ǜ�,�E5��8�[D��}�|����'+�p���ks�Dq�Q`����"&\��pvu|_���U�Nkg���ƻ�VK�)7 st���բA)��Wm�X��{���c���޲�bβ��9������ƅe��,̻���_g"��]1�?d�x���~-����0�soh�k��>1�F�ӑM�ȳT׆�F��\9#��rf�b%�ۼm����#���p�U/�^�w��Û�4
�z��g�|�)�M��1�t�&ҧ��T��v��=Qx4��\c_��,�K��o�S-��;3g�Sۨ���?�[�nۧ���J^��~lj��q�D�Q�4o��6�3 (- 7q�ݩ3�z��6"��b���yKu�eX�^�鿌wӇA���Zju�V�?������	��6��� 	"i_w6���4;K��m5x��jBۑ?�] `�6ܲMZ~���`'���%��8`!2�7�����ܸ	4�t�Qo��FC^�;;�	��h���33b��������K��Gυ7�q���ixgO�{F9�j�<����P�NWv@,la��I���@��Ú�i�$�s�ig'?;���������Р�"L{Ds�
}M��=T֙�X�`�P-a��	6v�K�M7nF-3j�8+�/�Μ&�7�S��!�8�T� N�ul�?�vw>"� ���D�Ȧ媱��u_&37FH�Z�G.��t��95��3u��"@�[8�,A˭��0�4�iZ�4�u�3���o����:��IxG���o{�,�R������G��	�W0qL�Dr�WFT%�2�ԣ9 �+)�V�!��2��H
�(�TqD_P>�B)�O�3��%��_Q[�;�P���
�x��+)��!Et�AD�
��s�	�u� �sӮ����>����k>�{�*�����OTj0 �U�O�ۑ
�Ǫ�͙iy�g�|5�],��c�%5�˪� �j�|	�[�A�
�Y$Z\��z���T]�Y.�q3�����y�O�+j�$)#�`�2��!��Ld7�胶&-\���dJ�pT7?a[�Pc=K��OYj4˙�H��^��q�f��!�U�ZM�O-\���w���^�5�܉`H��A����l7��_{o��Ӹ+ܦO������
�����e��1�`��)�z`!�RW��hx��A��O��9���>�4Gu~ ���?QI�t���R����=��Б����G�Y�������Oɴ\+�(�ʍ����}	ݾ|��:�V!���z }wF����zް��ԙ�4������|���>�񛲃�8��*�A�Є�/��-ֶU�<�~4�<�H�Pld5��O�Ad��ȿ�-֓M�ۦ�י��I��7`!j
R:���1΢�8��xO_(B-/%V7S�V�p;�&$�ѱ��?Ϝj�y�\�um/1�����=���>�����s�W���Jjd��2�g