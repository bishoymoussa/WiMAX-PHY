��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$Rx�y�<��wA�*;�x���@�̦�W�X�fa�M-$u����n~�%���P�$��W��kYَ���P7�?UMfT��q�6�U��k�>����~�\N�(�����X�e���/6U|)�X2pF�]$h���d.���9E�	�IN�f"�\��e�z�y�b�����Oo2�?�qˁ'�͜k-�K�P|����y:����3�l�d���bl��ˢ_�d���kx�rq�mh�MذM�`aS�.�DW�mS�9���Y��+�>��!��!�T�uOB���,��\L�7m�O��W���6����'���j)n_�I����2:��$�K�2�Sʫ��l ��!���{�l����.�j4�	��很�̢=�����N��s���s5���_�R�>����ТP .W;������	�"�מԫ�����]�#7@O+?�⡾�Ԫ���e�O�\A�	�ͼ���ƹ�d�	@�nQ˰��E؁Bf���|D_�%au�-�'���w�*%��"AM$w�*4���J*!Ԟ(�3/9(�o�P�lq��e���v?_�j���-�����[c*+�o�g��Q Ai*�,?�Ko�G�ϳ�n`�%�)�#���ض 97}P�P�9�$��[�w�7�A5�cď<AMkѨ�P`�ϸ�!�l@%�bgT��;Xb��웭'ԯ��k�������6}��%����A%�$z燦�FQ�	�
����G&�6'*|�S0����P���`_!J�-�4L�ԡ�J�z�<��t�]����+��ZZ�}oN�A+��%������JDY~]X���������0���_d��:�f�p�p9����Z|�(_�8/�|�V}�����~��F��v�A?��{{N�m��ZI����iZ}Bc���� �R]��Ҏp��(�,)y�dL&���"ʱ��6�
��{���ռ�B53W��MG�R�&D˘jy�]>��b�T4򯮼$L��n ���I�-�"�z9���nK��?�e-�/lU���|�y�W6b�m	�Ɖ�y��1�]Ӆ���v�:v�[�y[�0fN�}��&��A^&i���kg�����4�H^�$�I�N49��Pm*�*�`�J/�q��+�K�Ow���>�h�ҩ�A~��6�>��c�/����kK�Ĵ��Z� �����g�S0Ɔ��+y�u��
��qJ�^?�k`tʷF���y���Ǜ�H{姵�u*tэ�RU�dp�4�}�<�`��-4��r�*e=!+0sP�f�ܺ
d8KD7�t�[B�?�����E.?L���
���>�� )�.eq/�V0�P�HO�V�-;Hv�؜���!?+RBL�Ϩ/�?�SС��IV������,Z�UeE�\��H|SD�
I�-rE]
;4��B�0B��0àQ��/�X�pb;��zJ{ql�㷾к��uT$��������Q��2���X�_I�j YN0�2X�|x@RކPmY	���J��A�
�W�߿��X�q���_���0�tI*#�q�:��V'(��W��R`��'$��͝'���\�2>ƥ4�F/#+����{U����~�5�[)��UTyLz#m�x��I|r�JƲBK�,�W,�:Ff`lh�˱�+�H%��7��������~�郆rs�j}�:�<����T��9O�� �)�ο��%�8�#ɩ6|�z��ﮣr�h��8��P�0����^_X� ӏ�:�
�JCFB÷\�2�/T��S_��G�M��5�$ ��O�R@w�W��9��|q*T�C�[$�/��.�7���^r�Rol�1"Y}�X��	�w[�K��N��,2}Ȍؙ�<ؐD$�3Ȏ7�1~��a��`8�5�r�3Mq��۸(y`�Z��lt��ȇk}�ט�H@�Ѫ�c2P�òrs̫p���qq��g,�&�(��h�6��-�����|�l�z�������{MyY����>�K���6�#���G��lC`R���Z�0��Ȝxc���d[���ѫf�$��U2lX���$��\c�(ǋ��5z��r׿�!B�J�?���o���^@��W�o�X�[F�xt�:Ek]��&�.����cB�Q&6���8 �Y�P`�n��wC�\D�� ��K����hP��OlZ�������i}3�"��Ǉ��i��d��(�5[p�A�H>�'}4�Z_(��K�rX�_�.�.!� &�3��
���C�U{G��b�|�g��A�].R�� I`wb]-~J��P�W�}u�*��#������k��?���/�$����u�3E��xM<���>Umq͝�7�rF�rE|�!�{��}�ꓗ�<N�N��wc���艈��ͳ4���v�Q��;f����s��^LVQn��y��5�P�3p,+@#�"���>�,��	���;T�̩r�e�a���,�E�����w S{�ۭ�î��_	G3�6��ܪ��+k����gO��p5�ʭ �mD��5��"�W�$�B� �&�	���sr%��;4�9$�)-_��rM����#k��D�~%�9�N�Kv��"Wp�.I�	���}��u���T�)ԛpE./��۴����Wkm!��2c�i��+C�O�|���ׂbtBiUE+��X�����e�1������\��@�oC1���
���MIQ!�,�޹!��HO2ko2��j��;�	9��`�rj����=�-e5+C3�A���W+(��ŗ�hQ�~��IW&$�z"��BW�ؑ�h�� ����4�B�ֹ�~��W��d���F|��/O��J�nI5z�%d���lC�60l�!���)̻ҕl��j��j<��7��)2 ���PX/��j#���eL���L'y&׶#^!6�)��a�F��-p3H��.�nB�2(RR�e"�/*����s�ǯ��Bs�ׂs���/ p4�y!e�f)]]���,��!�Z�ҢJqrʺw�����$�����?%�eaq0_%ě]�i�RbE�u���sg	���9�2ZH\�5�/��KZ#�?�-s��d���\�-��G]	}N��Э�pJ�.��LZ
tɜ��@G��F$Lc�<4��X���(�G��	�,���:7lr^E��ʶk�єEy�������H7n�ࢅ�\Ԥ�T^�C�2�m�i�(�������GH�%o���O���?͂�X �a#��9=ʄ[8(�8"Oll�z����G]bo,W:g�r�i��J#���FF(��eySQ��RM�1k�c�\��Q=\M#j��I�XBT��D��/^���\UK!\0-W[ ����f�p]g��2e�jx�n�GT����6Q��|åI89��3�c2k�f0�q�aeK=�
�|���~DT^�@�A!b��=SM�qd�2����N�E]��^/ I��$3�ۛ�m9���'Kp�%���+�����Hh�4w)��؃�ɲO�%�De�����^�͓��ȹ^rD�����sׂjͤGݼL�<�vr���!N}|����M[Dh+����~�����d�l��q+�X}h�A3y ��3i�$.�Y�w��5YL]�޼Q��b�m�=?&��p��+�W<|��l}�+m���p��0(���_(O��F������7��jDk:@Vb���V���ݭ�>K�Ѯ��"�`�Ռ��ג~��څ��'�c�4LL6G��f���Xl�xWHό��\l��xByэ�u a��H���;��ad��e����9OW ���3�fA[��|�4$��Ci��~�:n��N����z�9+�}'�:A	+:Nd�������L@m��x�^ykZZg5dS��z�����>�
ý5�M��-ɲ��L܈Q���.���y0t�:��c�O�w��X�����4���N9�Ĉ��N����fS��<fx_Mm���l��.W�o��m�mY��e`pU@�G�^sGv�!�=�^�)����I�emo��#�-�1�Z[��|01�cUP{L�4���=�) ;��Ka�wrk]���+�X��������G��Kb����˦��*�R��T�TT�)�86 ;������c�:nR�?x@ZD�>�C���_�������${l�O�Ss��ܠզ�8��횁���R=���-�\`P|�X�e7e�m)S��*W����r.u��w+f����`�ֿ��<�Rs�p3A�1��b􉫔�w�c벷ok��m���GK�SN��V��Q3��i�"��Hd���Iy�[*�~w���S"ɽa9W�&�u*s��Z8�Kce|y
�w��hU�?������O�ksN�J��!�B�-�ퟟ������u���۾q�W'�C$������`�I;��,�|��\�}���9��|�S��P�a�:�:�s�a�Gg�Z�R����I!l�����kb;{�'���ɘ�������lc�!�|����h�R��T��)\$��޳�����ȖY�`6��"�T�� ������PIՑ�I��g�)^%&is�lý�7�M���h�-35�:�p��)�^�뫦�Z-�W�F� �Ű,���Do��������k���a�l+,K���d���UL�9H�����8�����EG��Y 4��/��R������R+��	�.'q@>�sk��#�U=�υv�%��{*��a��L�f�~�m�(G4���y��@��򦿵V0��͂XTK�|��g�G#�?�<jᳵ"I��+�=-�v4�&[�Qzo�8�p��BZ�H��Hfh�C��v�KzG|�Ԩ�p�s���(���$WW���tg��3v�':P��P���/j�̑^���^�QHs���Or�Zn3p�Aׄ�FMژ�����H6P�ð�v����APQ6��B��p�@����"-�b-�U~o/P���4(F�7r�&�����3Q`�d�4��� o�PRXgA�8��^N�1��Q����'yBϐ�����[�FP�r�������&![d�a����ڟ�߯ U}O����Z!Ok8X���+9�*��S9[�7��w��G��L��ŗNL���f�6E�p�A<X�� 1���r'n\�����˕{���̙�<��ik��C �����P��j���L�K.���)F�����)�S��HY�N�������2VG^���7���\)*!�:)J[0�;�#R�i�W�9�z�N��i�4�/h�:���ѵ ��j�x)E�E�XD��,��4��W&F0�D���.g���ѻ�t��v����KF֝S\��}[^clٮ�^f�Z�G�t�ĳ˔�f
���A"6�3ݦ�֓�ɲ����,� P�'xR��¯g�`L~K�OdG/�W��YI�F7Ѐ����
;��%%�G0�%��C�N 1��rѓ����Fc[�Xy��s�?rLC�4`l*7Z@�<X�qu��Z�#����Gs���p�B�:f#VU?_L�ǈ��>P򍖴6�v��n�K�T���);���N#�j����D��%�z� b>���0���5y2���%�K�*�֐8���������yb�w.�����4�
%aR^��v�\0��:l>ei�i���Y&Up$��t�1�W�gZ'��>\3���K�5�_r��(A�7�c�џ�G�������d}H7A�abD��D�ܹr�e����0�@��f�Ih��Q�h?�_���ͨ�#Ƭ\?�ø���jSn˶�yL뒊ٮ�pcsp��>u	���U<��+yV�Ss_Νw�'>�R�4>�Đ���M�Iw]���T���`�(�we��{T���N�V�6l��\�o`֗A�Mæ��ǉ�_0�Y���|\1$3�d�1��K��.۔拚l��[���s�ܝ�G�1��K�5I�t#s�/�m;����y��[B�j�e�ƕ�%Ļ��>��zM|)���[G�[�:�*���\Y��0{0��Q��[k>b�5s�4�pnRU9@��>��8��׿�@����fC�B泱|��XI�E�;��Uq��:̩��ڮݳ�X�r:����ʌ��G:�����nHs�ŕ��./��>w�a�t��!�����Q��y���&þR��Χ*����=�">cvo1��@�����L�B}�!\j����zE��A��0��K��s��fĽ����؍�' �gX���J�6έ]/-�c���L!D���י�F<�4F�G�wH�m8?���"�0�⚹wYݨ�EC��.=��{����*���6&�D��"��b�9j�c���}wHbqL���
��^���6�0����X-U�~������ S<;�
��	��6:9׊�=����`)�HH��vh�A�'�G%�Q?Q�Ee�l���^/��ls����⺫B:/���D���e#�2�𭴋� S����	3�+�Ef&��l�z�ƭ|#�ΞC�& ��0:+/��#�%��)
Ҭ�y�W�6�nI�n��0�c�<��>�a��)�Qf�h�'�!�q��/�=��=���yl����ƞ����F_T$b�h����<j+��T� dm�3i��X{���~0���m3��֌��N�ϵ��l�������,c�v���rY ��R2�j�L��(���|킩Q��}�J"]
�J��|����e�\-�l%�7������-�6���!������9D���C��Р�Ih����Z�������hz�'!�yhS��j���Y`O=Ab�W2	�&�a�TR�0i[.�Y��������~��	hC�����Оhب�̕�;$S{~��ӯ����h������]��fd��A)F~�݄���k
��{@ӡj�#�"x�>��#����U�-�=-��/Ҏm�x�@��p!~��ڟ�T���/\ae��a��[8,�,6Ӿ"3�/SHS�Q|�_������W��S�P���`#&��X(���*T�ᄦ��r��8U� �g��W\�W�/�3�.�q��Z��Vm����B�%FO� ���ְ��/����l�?��9�#&@yW�貯�_]볤v��C"$n���2�j�ݴJ3%�u�Յ���Y�0��@�kS�)�ʪsg�<I��T#	�9J5�@�'֭H�}",n�b���EL�����i���"�b� /�C��SJ�g6,f�u��N�p2Mȴ��L:��/��i��e�����O	'ⷑ�v!�V��.;�х&o�w�ò������@j���+���܌��q�1����a��I�
���p�2����ßЎ9|(�Zz�4ҁ�C�����S{$�Ь�\�g�k�P�;`��-�^*��Qr���To�sJ�sk�
��G��E�P�-�^�}��*u >�� �O�,�d�}�jkE�C�!�>��xq���@,����e�H���t�a�O� geg��H�$$W4Rdqmv��Υ2F��-1N����4RΣ�ɼZr�M틊�]<����(����x b���K�:�2�qh<������@3�H�H�F#�\�}�Mv�¥8,���|���v)���$6{M�:De>�Сu�{���	~=�坻)q��9؆�T�!��cY�7��@�ѦP��uB�~���OH��z�|���|�Rd�����I_�6B��j1t����c�V��+ҫ&DDt��o?$}��<N�)�e�w��-fvQw�S��#�T�*��U���ck*�5�XL���G�?@�G��������N���WBq�/~���qP�RA����{
�{H:�B|�)�[��Y��نc�	,z�+1]ݦ�0W�Xk�；�Ҵ�L�_ǘ��;��5���)I�-�x
�4*�:>����05��$� C��nR� ����g�!
o}�`A��+@�hƥ���: Y#}a�����LT��[�T ���������qn�f��pK����}_N�+IP\[��}S�<�Z��Z�K-�Ȳ఍KG�fyӟ��h����rb5�ov9h�Oi��<�E����mr�0�H�Mf��g�m����5e�9�2�2�Lِ�<Q�1�����"Z��@m�B��Il�I���CM�MBs���7�H����T*�Y�d{�<q�� ���;)���"����P�2���yU��<��G���pDO���;M��M.����s��J����JE���2P�1� Ʊ����zz��4[�"5�ӊ3�a0���e�V�����PH���OGo�eQ%�LA|���d4��%�D�������Qӧ�[�"��F_�'�����	a�)f�Ҫ[}�le�$�v�#��	�Mx3��w�}�`J	Gd��$z������1����̸����t7Q�f�������Jrr��h��U�-SP�!�÷,I�xd�;���C*�r)
6��c0��(TؓZj��~���/���7���hV�a�~�bwcy��_��i�7��%��ϧ���˸�AeguS��G�(��OU�ysf����ί�C8t�����z��r�ظ���c��])�?z��ҡ3OLDӄ���ʍ��ȧ�"�k<9_���u��aEF�0:��F�T��}y<�Z��Z�0�0X��%�!ۚB��E�g �Q�! m�O�+�����:����gW$�jvx�7���q�A�j^vTy(K�jS�7��yr����ܐ()�/F@��߷�O���Ŭ1r
3�k�z��!�id�?9y�'�2}Z�|A�1%f��9���ƍ�EQX,�w�sθ�� ��M�S�R�����2�ю�4��t�d��n���C�r�L(��I�p�9f����T��J�?��p]⸏��Q���F&�;G���b������q�Į +�u��G����y}IW����Ѷr�3��?�I(�̢�ڻ�ֵG	?G#��Ғ�y��AO�D/uT�e|;�0"m'��Я<`�)��.��@��)H�3,6k��0� ӊ�� D���#Ɠ{ld>�C��"s�r�^�L$��] A̝t榗��M8"�;W�~�A+OZ`Sè���3�~[]���x�"��N�.�m��܂l�OM5�㔇v�[ D����Y��V޴o�ٯ�i��ǂ��4�t���C�"d�ZU�p=o=�N7�jl�,lq�wn��k���L;s׈�!��(�P�bD�Y��1�rQ�w����'���fX�x�L�����n]�{�Ѣ��7�0���9��C%���a��٧�ˠ�6w� ���݆�jQ[���5-�"�}��5j%U�5+�L�5�UE�����r<��:y�x�RN	kx5s�\70����)tvk?��b�g�8z���+<|�7�k��?s�Nj�M|CQ���01�=���U;ݝ�c���
\�Ќ��@���$?r��QٶF���31'���o����������M�<N@+e�]A9�y0gvH��ȅ���x%3��nq�a ���� �W�����^�=��/<�� �f�~<��N��z�4�ĝ ��OEѴi�԰���?�w��]d����߮u�Fdl*x9IM�Mx`	C��{�]�S��F�Q9���J-����ܳ�
�Ӛ�O��tbd�h���S���[��J��ո��q�i�M���@�Q��x޹+��b4����B`o�a�㐸�LvQ��)VV���Ms�"N̍(��
�:W���0�+�<V���T�˕
=>�A;���� ���e]O%�?_(J�D��z��3��)�3ˊ�ȷT�|�u��gm��ɮ���XZJv|����B�'t��e���. �5�V�g�3?�ˎ$M#(	{]�g��'8]r�˄���6�)K��у7}Zӭ�)�sJ��9�<Ҭ���A�'�j����8蘬�\�Y�E����3Lr�XqCh��|(?����0%�z\�|o���q�]*GK[�YU~�-��m����W�s���f����Ö(�r�Ȳ�h�u�����+dS3ZV��&�%p�]�B�ߋ8��.���_ �>l����?,��oV�����:U�Hhγ�&}-���MK�ⷚ�S��z8!g���}�^Y�o�f�Ҳ�{Y���w���T����K8�U j>�CZŤ'{�j2�f����<�_��K@�ʘVmb�,p"=	�7�i��bY���ǹl- E%��އ=�?V>��&�Y�靪��4����������1��'4.NW�3�g�C���=��s����|7�TMC���|	�r����������4��?ZV�U*:���g�ǎ���X`�w�e���̌'�f�Q�� e��|�8ˀ�N��O�Ii������S�uKV�G�(������E#�9���N�l���z�ΠЁ-�n��
<��>��5iJ�[�]{�y��B�{�W�C���7�� ��h�n�T�8���5����փbulc$���)3K.4����z�i�#݈��?XqeO`��� <��FQ����{n�_H��>���@d޻�]�a�]��+VJfߡ�=6��v��>Hn�Ҡ�+�UZ�B�_0��&!߳X�U�J�eΤ�ds(j����R�F���u��Oy�聯ĕ,؉�#7�mq7�[�)X��T���S'זV��f�Zc�Z���\ޒ���%m�ӐU�$Q�]}��s�Io�	����9�a�6�(�{j��^��n� 8�7��x�����@*�H���Nre_�n��;��uZ���sɯ@`�k�m�/@A<;,���e`l��g��J��wU��X��Φ't����.�ns�:�ae�9���.l�C�-��~��Ծ:8��&� ��(O�xf�!���I��%ρ<�R�/�{X��ndz�^>�g�~ڈ�x�HP�7�2��J�h���5����R�����6J�L���s�]F��p�9�
�w��?�����юs��}�-����Ue�dYf?�	�H<_	$f'򪉓k�XN���B��"�+�
�uךd2o%9Dg�n�R�Zp��n��!�����-�[�RM���7���Qz�_cz��RQ��<�'�x�ذc~Ig���j�:\�q� �������>ΌR�wE#��2�`g�T�����p�:�Mhpq�j�2�J���X֭=�_�>w�u��h����G\?�U�~&���߽Ki�M�{ZF�������g�����j%X�	��3�2�cg�uڳ�J���42nR����5Px&�S"�3L�\�,-�����4�ɣ��JZ��vw����t�E�TDEOo��bN��ǘ���hO���p2�W���DZ ónƍ��
H�<��f�\�eR���d*J�P[�0�~��ˣ|2nD���C�������^:�zׇ��t �����Ap?l�+W����]���Y~�U�\M�+UX�>�TnC��E�~��ST滿��e�Q�g>����2K{�e���i�Y8G���N:�����g E�x8Y���uE�b���i_���љ ��W59�\?�Nx�5ǌ*��qa'RV�rA�c���� �;��
��n�=C8��8�/��:Z2�*��^C54�;~ ��/�GHhv���ݾ���0v��W�VJ�A����������-�P���+SE�X�<6`a�
݊v'����~�{�-�wC�$��8[�D�9�P0t��T��9#�mj��'ȧ1��s=����'!n���$g�H(�0�	b >o �n�v�{�ZC����@j9�݂VL$3����K"�Q���&G���*����q��,�hjЛ�@P�E�0���D�c9��ĥ�D��Sz$���'U�	��h��Is�0~ś�4H����+���%*���\��9�O;!�yoЉYk�ůe��AT^/A<�jf0�#M`2�!a����X��0��<�D��I�v�9�8}F`Du0 ��Ҙ+�0�s�mWF,�y/��,��*5��f���'dC[�K{��c��?�~��L���g����jhL���b��jd��0��v<��<
D����Ob��@��6�5٪7��B+	��dR����{��iޏ�"�Â�iN�C����!���|��������f%��~N�eGh&#��W$�:ٚm,�%|X_f>�%�2>�M���X�x@��6��Gz��~��b��$�}S^o�����!'�s��b��3�<kD�W�����,��V�1����Z��hW��~W˅�=F�o �����Fj���|n��Z�W'Y֭�^��	V*@76K�g��+%�ZDK,Z�.��5�I����]�r3�ݍW�0 t!O(��|o/��G�(��.^och�������z��M7X)�/�7��2���ggޥ'�{܆/����qu����\掂���a�'Ly��p��z����P~a^�)����&�&�9��NӨ^���`2��}SlW@$��/e���P�!�+k�~���<������M�6�,����E#��� ���8��]3s�r��2#�SO2�<cw WV�y-��ޗ%�?����&2I�U�}]o����
�;�T�&�l�ET��y�ȞM�D;���`=��Ƕ�z�(�y ����"���{U� AE�۩�H�H�( f�<��w��q\������K5�l̓�|����/����T�ל��0��.�C��˷Z�Kp��J~����*�������l8�ر�yrU�#<�A��%��Jc߸�7/ʵE�nG�y^ߞ��fȒYJ�L��⌉��%���I��g�o��ܼ�K��bP'Fm�:�D	#s�6�E�\��S�
p���Hg�1�A��g(�Y�9�3 ��H
�ٗ4Ih��Ol��2Uy{<�+;;�K�)� ��d�
�e��5_Np�
�P��ei��U�nh��0�"K��R���Ac�rEQV���X��%�˫�6\@�+����mM��`GLyԠ��S��������D.J�di�Aew�����@�����|�U3"�p)/����,����}�y7�2`�W&F���F_�8��5�����SJ-�x𐪷<�|��{� � h�s�w��Z$�Mh/�k�]�t�R~�zOq��߭�����A>W�-��DAĚ����'�vĠ�MW�� ?��(��n��B+~��IN���,����S'�C�%�m-k���׬�b�Wˍ�hB� �KC��j�V@1��.�X����\&���!�]�c��T�	��x�e��Ct��\۬K�e�ɯ�p)�6�H: �[�Yi�`�\3� �x8�A��j�a'��a¡-�U�8�e�\XW,<��K�j��S�w��ĩp�W�s׵��Tw�[�9?��A����!�E~P�R94_Dm@GE�q}�wu����i�<�6�wv��&qO�H1�k�i�9�3�2$!�������3gBOKJ�w��� �b���Kc��୾GI!����=;ɫ��fK��0J�>��~l�T\a�֖۩2]@�hV�j��\��7y��>���&x^Փ�W%'u�]�	ߟ5�7W*e��������X �aW��k<5��$��1�_M` )Z�i*
��ʌf���h?0�	0e
�7��H=�n͋k�ϰ�9���ZB��l�j�<�[���| ���b�ɍ]_���U�p��H5*mI]�eAr%FH���
��	@��Ma�LR}|��Н-aG�*���5����m���_/K�Y��;x�`���A��������G�y+�mg�5+4�V���oь��� 1?�2<P[����U�&D_�x�x�B���*AJx�я/q��������Ѧ�,����_D��l��������c}��5�`:����1�<�IeDp��We��څ�m 2"!�8�ǫ8�-v�'#�,�EO7�t��9*�g�<bX}�*�|��H�����M�̎���@k������}�"{�6��4L,	�Ԫ�|.�!����!�<�1Tt~����~��������ET3"�=Ye|��c�j�Wgٙ*"��?�-V�fS�Ɋ�BbF	�}�Yb�x�	�
5�>hhLONr�"n��ca�!��CR%�(d�ۆ2$��c�Gg�\>'�Y�m|����@Z1�sM������h\��P�C2��^[��}ѲI"��vUI7Oɛ	W���5�>�����c[�3	?�ޤ�}�\�[z��z�
�l��㸙Tu�iJ����ܡ@�^m"qV�ȍhՀE��9����F�w-L�ɇ��]|�P�ճ?�m��][3�E.�)���[]� p��J����ζ]]m24^M�_3*Z ���o�6��xT ��F�"MY8��Jy�	|H����
�bE��"CD����{x&��f���'M�R� '�V�^��h2�A/��e�\��w�e\q��'��o�b�
�)Ę�l&��Ӎ���8��B.p%�u�񼗭1}O��Hb����VA�n�K<}OV��5'���=9$J��?�\��OoY�D�rYq���Th��xB=��%�!���q�S.O��_���m�	�6ayG�����\�pr�c�v����yNd�z�;3����]��c~��Z��gE����K!���ی�J����HE��C��S/Rb����՜}��*ģ�K2�cb_���䩤� 4�?�����)z��3�ui�E�["����+�O ��ҝme�6M
Ú�Nd^ԆZzMz����7��|�&�+L�t7[��|�oooz�/����s��ͻ���ͦX��vy�s3��4��1A����z�8�{у����e��޳C�i�U�<E
ӗ��.��D� l�+�r�����w�:U��I�����Q+F���ݱ-��J�N3�m��w4�s���pב��n[�"��\���r�>�-��U$*�0�$p��1�?b�,#��j����k��B(]W����̴�1��o��H��H}�7������>
_��2��fK��+[�	ް�Ͳ��[n�e#��i�M[����:t�D��w��VE�J	ڡovC��$���B�]�2g!mĬ�Rob�Lic���}æ�˴ y������8�9�}�V�Wș.������M�4��-8R��D��*�svS��eI[ ���H�.�NO�\��	����d�����<дO$�6^ W������b��`�j�;պ��w�50sO��a.���?|"FPK�a�����G0czCj�����Ha �e��K�SO�_B-���T�ҭ�,N�+�3�@jA\6S�J!�ë<��`X{]�%�h���/���lc���r�\K%U/��c�97���P�CM�&����I��ǉ��;���3O���ȍm�����sy�FT� �m�]E��_�~�/��@�`N�@�7F�GNU�k��w�c!A�Hh�Vf���ͺ�qJ���4�N�ޡ������~	:���M�ܫ+�*�X�ɾ���ƃ_��i4J|�Ɍ��*�	9\�7�]�&n��!�[�X��`F�w�G�R�% �W��~�-qG�~��[�����9�̴����.ݥ\F�D����l�Wԗ8���rE��_�I����nt��j��)�����S_��s��'�bVL���-���)Lc����s���jm|X�]73�W?���r f-�0	A�RJt�5�<�Y��)4՝��~� ���mL�'
d��Æ'Y�nzb
|ಇ���WL��)�ߵ�R7��+�Y0�P�w��;'گwI`�h�Lj=U��  �k�-�f�%C�6q���}
V�;t�>�k�@b~��c�W��X3��s��T�Gc>�ʘ`���k*���	&�{�#�+0P4��e�J��(�-����<o՝P�h���w'~� �k�tg7Z<T}�r"+��9Z��������Z��_��o��4!0��C*hs,ƓF���h�h���8Ĺ�d��e����z��p;I�yN��2蟰���S)�z���B��ά����͌�_��o{j�=�%�b���`�*�!�X$�,|����|m�{�
X�+)m����f_����N�0�z�j���2�x9���v�p� ���,������8���uyYk���!P�����4X��!�<;����m��S����� �q��0�:�E@��sKSS�أ����d�Mpd���LD�8�M�-�5S����/��eз���0XTl+;��.J��_~dH/�n���/;�﹵�I�w擆D`:����4����{�@��5	�ZL���y����%�\^��s��Q�mI�P�D5�����7�0#^c��Dr](1��%2�� �$���B��؈���:�ƶ�Zy����o�i���N�nt���9�JM��vɈ�t�p�4j���b�L����^S8v�U��q����8�6��_VR�ys�l'�/hZ���,����_y�EImz�ؖ��J������k����]�A0��	�CEYb�׵q�]Tf�n�Q'!Xămn��/�*	�-La��i�\y΂{�!%z���;�k]�������8/ə���m���2W�s)���yf�����\ �5b�æH��"�bݦ�b���k������ӫ�4ya��.��\�G�ݷ��q�rr	��p�'k`�e|� �U�sΘ�z�BHn�� dC��$���Қ� �̭e`��n9�$��n���q��BU$
��gO�&��Ἳfhݥ/���⍔��=J�4�삖^[B6����=燗�3��Ćb�>� �~�Ud��Y�av��¥��=�:b���8M @�
X��7���ٮ�Z�C�Яz�'��Ѹyأ���D>�ǹ]}��F�WI����̏��Z6�Do�љ���핂2�qu��Υ�b���7MY�z����z�����S��/[:�h����X%/�ש��z|�`Zv�x�	�|��� {�t�51k��t������I�+z�9Qѥ��NV/nS�3�&Q��ts�Ys�1��� �Ӱ�Ca�y��,��-��^��Q_�6��Yb�m�kT��&�et=��o6���șS���|�_�.���^��?��, �SsW٬n��Rx ۞������ �%A�f ��m��;M5��C��1�S�sRC$��tV��&�x�������w{�l&��P�*��.�����ݙ�k&B$Ea�O���v�/l	��f��Sn䗙�����ıe���7^��u���?Š�̤���
�:єEH��V?�즞֨����è����&l�R�P��:��v9����U��a��$�q��,j9L���G!���>�2y.��T��b��y��ZNS�SDOyaϏox~�X"���gp� ����ރW���T�ǝ{֞�"�Ġ�
_��������E%�gQ�{��=�g�������L���Slptk���#�8����g��揇�����X�U^y�ۻ�L7��<�8u[W@Wv�q��r�A�H�X��ݴi��b�$>6.����,��#�^�܃	l�g����<9 �-��*r������o�Vv�Kn�����~�j_}}f�U����ܸ���6��f�������r�5�{O'r�����
ߺ������HM�|f׎-�GnIR��.�Xě�5T�%L���<0�F���u�ms9�
���=�k�RX��1��3��dkǢ�i�[��Lk����3�|y��¾�G���;�'+5�E�۲8���ǵ��s[0���́a�h1�0h�~2��J�Qp�����x���`��踜����~�F�P;Y�dh�ɊE"���br>��;��d��*=ߣ���'NT)}�1��Oѭ�����N#~6�F����%�$�A½�-O.>�q�0�fY��2�	h�)�#fy��m�ǁ�(�e�s�!�'��Z4H�
4tr��vR����X>X!&~���9�F�= �ђ[s誷H����պ�J��(6Kײ��{*U�N�uRP�l�I�k�c;����?�كt.��}׫e�� Qa,L�O�>W�߲R2�G�,��e�LNX��[>�M<j��	Sc����i�=�{Z;8	TW������� 	��aX�'�Vd�8�4�����/�Q,�i7N;p���p�L� �|ozrg����Sb��`ߢ���6OB�Iq��pv֣O�b��v��հ^��G��I���tF�A��w4,v�]�_�L����W"vA.�:�ց䑷Xnw6�:OVa�^�]��D���h��*M�o����Ž�K���RefI��u��v��wO6�w/<ʩ��gI�Co)�a��nr�u���h�����f����2�;�͡���������~H���C�.�/�(88�ؠ�K����*�S�p�Q��=�ǧo��0N�Q�B;^Y�Bۥ�RP3^�����s��7�[6nA��定Pβ�*�	��t�YHh��ژg�C�~���;}ʈ�8�j�N�w<P��ka��N0�rCƛ��"g�>i��'2��/�̍9�B�6ߗ�$���v��A� 
)�G�q�Z-��p���'�A���~��+x�!���Ż}b�mj�N,͹�z���{E��e�N|2���?vo���?�0s��6�qd~���琵L���n6��@�Q�ޤ�9Đ��n�"z�lհV�Lk�f��r��0�'��4xJ��M�Ҟ�)/�����9�uZ	f���H\6�R�ʂ�K�����o$�,:��O[=P̸��ֶa~#u�Z��D��2(�`|��4���¸y�<���{�k`.�U��+��6�Wy�}�)kj��r"R�4���Tt�'h�h��L��pM ����7?��_E{;8�-j��<�ҠY�,�c>d����y�	��@
��ƴG.(U�����L�-R��s��i,��V���|γ�e�xXڑ3�eX!T� �")u��۠u��"s���i,�����tB� p���ν���6���:Я��"�>fA�id��Ů
��%��f�(���V�U��!K�t�S��g�T����0a�I�x���6 ������1���	��;��Ԅ�PVkM��I����p��#���hd}D��,2m����x.��:���Π��R*?��8e�� ���7j>G�����b�|1�e�ˢ�Z�y�4j����VF�JR>�u0a'��m��+k4���:������z�~��!��$�Gf�����ϭ؄6��]���<��`�>�z?3�&�|P�HS� g��'��M���{��I���?ݘ���r��ֵ�_�'���j��9��X�]$*1$v"�>�8T�}��ҽq)���8t������o��������<���#�- uL��!�h/��pF�Zp�'_�L����(��>�x�G�����C4��U�y UD�gBS��TW�Q����4$9�YŻ��C��y�m�x����̍��bQ��I`GY˒i �����.~�k��
@[72�	4_F<�)�i�N(<�] p̌��Kԙ��Ȳ0AM�C�mG��d��ǐy*�L�7�h`J����ME�W���u��U��>D���'C��e$G]�����ٍ*b���2�nN�"+W�d����j�Ά��q��>�;��R��
/{��^��KA��[2T�!��v$�ǿ�&k�~��GWN��Pu	�1���=>��N��	�f �2ā�2�+�:O۱�v���欴�CV�>�$W|�O�1�z���w/^N���c���
̹X��9�;�����qg�V��kG��w��mGF�\��bb<�I_�V*M���
e'#u�Ot?�T�SF���>Rm]���*z$^߻���H"mD��@�5� ��zeLA��u�Mgx&��@���ƾ�}>Ƅ�hc̏��^q�'��e��2���#����O��y��h��j'R�cݒ�㲺��m����� �\�Bǜ�-���G8T{����9���樌#���<32�~��3���GL�
�]�bO�
��hX���:.�����_H0�	f�!��,r/x�,+�y�F���U��1��I�_6����h�-O�����у:ʡ)*��0g�Ҡ`�`'�0�@�Ska�(��&l�q]�Ιi7�A,b�z�܃�2�|Grf�{M9�4�}َ�.Wֶ+��S��,i�cYU�8&KsR<�XB����#a�;�<�`=�տ�GI��ǣ�P� �F�����v�!Y�����k%̉�y��o��B�x�3dB�x bl���3��&�����s�rܱ�'�7����߈�=�Wn�> �����\������b�ޮ?�����������&%������)�,�2{5e�y�W�
eH����qG�d3I_ii�|@�����W[�Y�夺�!�́\�{�#��¦�������H5'�7�D5�Rq � U�;�Іrȧ�)��g$r���we����HRH�Ei-I��=��@�k�ǛR��7	.����w��/*�����:�©A?�[c�)�H�5ڇ�z\�푰�c�g���I�;Q�+�����G��4�M�Oڊޘ���$g�Lrudݟ�C��-'Ud�.�%d������K/�vL����*�ǅ۩'3e�=�%2H�|;�`Ni��K{�7�	Ӯi�� a��-��� ��GDn���h����_�����m�Ŋ�X��ܬ�V}��a[>�zu!0π��$��ዏ�\��,��������rh����"Ԯ6�@�*�bS:$��
H���sI�q�FeG H	�){ZV��^"ݞѷ_�}c�ר�4�Nr�h�_Ĝ1/���v��͡��V^���=<\Q>�Ҁ��a{�Gp�M!����I)�X���9��ln�ū���ic,y�2���?`dDބ�	���Пd0Hqr���:���yr���"C2��0�%�@z�G���e��Ads��g��.��{�v�^��>�ظ��@���-�ŵ��S�n"-��8������W�ǣ���x&�N ���M搜!�$GM,��W)V@�Z-�ϋ]81����$��b�{�(����G+>=E*<%��xߪq�Y����|d�٦��P���:�c���w&�}s��~��N"^���1��oF>{\�A([��cR�x_{2�F��0�߅c�2n�!$I��x��P!����u���|��^&�6-���ن!-r*�:����؂�nD�_�A޴�#�j$�ܽޫ����cW��8?,���7������Z-��
��;H���J���v��-dJ��9DG��ñ�@�N�7�PH���z�a�F����!Q�u�ĞE��*�nN�;B:���j�]�z9+1���8�W�S�w�fȡů)]8?T�5�QD�h!j�[c6�g�h�%��WjX�aw�Cnhh)�:� ��Ĵ�R��[v}t ͐s= lѩ��#����8L�$�v��X�w�~u�N����}B�Eq��')�b3��^j�.�y��(S��$�i�'�$�MQ�v��x`�/�˨�s>�:� W �Q�C�H�]7J�����
}J�����1�u��~�~���F�L��#"^8�B{ӘqqσW�3���m��ӡ ���P��@�LF���r���ϲ��^�����mK�g�/K�n��<�0����s� �H�o]���-�TҎ���/r�c�(ׁ^sn�]ߐ
��E�����h�u܋sq�*8G�t�x�q�0bWbG�'I��nP��ӧy�=��4���9�_�������)89H
Vqh��=�,��T,-L�H�)����0��CڣՊX�[�u$��88�L2 ���m�o�R��tH�Z�z�آW��_�%�ДcvO�4<1�L�=�qV�"��g-�d3%�\��)��qm����ր�xAo=M��zE4$�,7�z��~J��Z�h��o�v��|/���@�}�.|�n�b���0�>�;N�����T��6!1��"���ɤF���0O<�wJ��<�%�K(2Mz�1yXs�A�-Aݞv�9b_,Y����������g]��"���z⛈G��lJغ\��x��0��[a�nħQNmN�|�)'%B��2؅
E��\�!D�҂p�,�Y�w�}�ɱ	����'볩�ыث�[�n40Y�^n{��<d�6cNS)��܏%�<�$��":����D�2�W�{�q��pH�ζ�
]�6lu��XkIH(q�4~�ٔ���n�IY���s0�h:��K�|�Gw�fx�I�1j�RA�|�	�uUԓ�en��^��pU��!���7T��A�}\Q]��l���>h�t�~�r�nI���e���
�Sr{U�X�M�I���?"���t$�⛢�$���Bh/�������-��|��ݚ�Ѣ��P�zM
b'�y�Pa`����X��5$k� �����]�{9�A�"���e�^�W5��2���?���-�u�H�X�t�L���L<m�@1A~�Y�� �rAH��_���`�d@Zϖ'���+����n|�#���r	�F�0�DYb�_�~
)��4#��yg�&Khe�����bs]��&9�y亘�~���N��S*���w<�W/_�V��^":H+B�~�7�t�aف!47���M�KԵ��Y�X��,��&&�inu���k��)sM)۲�h�'M���)<��&
�9� �k�7<`��r�L�]�����	:�N��S�e,9蛪�5oZ.�K��U�:.b��6ē��+�o��|�8 �A����`�f����;Q��pQ]0�6��m|sN1hA��&(	 0�� ĳ��\Њ�h�i�٘���V+cu
�_� ��|㔗�����7?hɆsw��Kmk�����+��8ur>cݖ�ß@כ��|_��7������!�{ P��2��o>9�jʼԻ�H��ϐ�@�q����8_���8�5g&�&7�5y�;~���]��k�v�[�}ǤAy�5�n]��� sM.z��*�!(63z���=��-�߉���$��Ժr����#ϱ�1�_�7�cs�j�DL�iT�<`�+�iˡ_��|*3�!%�4U_]���8_�RT;,���t��
�4���DF��]��kų��Ջ��T7�Tg�r2_b�=���Y^���ٷ�RUh-���k������WΘ�x�U��y�׼��9}�ڿ�v��40���A,M���>L�t6<o>�mՀ g�q`��(�͸-cR<�H�
j6S�h������.����7%��!f�4��aK�"M*�c����}x%��2��c͸F���uO�0Kz��\ڎ|�>� ����H����X�$*䙚Ge"������pV4�φ����v�P�iC/��K����<��e*@�׀i%�j�s�ԅL�ٷ�#�@og!�v��pK߀��5��>߫n4!v`(��G�������.,!(]���D�H�Y�po��PF���������}�)o�j�0������/#�o٪0>�K�`?�ղV�g=,�=0��T�ϹeN���_Oz׵غ_+�=VV��~��I�Tq*M��1!{��J��u��L�P0���f1�)>���z-MV���V� Iق'����S!�D��C�x����P!�1W�]0a9�E�PP��$U�~��
����q�.�ZR��?��.�ѡ�B\�2��}��B�	h#����z0�����%�v�� ڽ(;�w?n�R�P�N��a��m��/�$i���L�k����{6q������P4Ĭ�;��/(�j	U�d�c���PQa:(��?J�A�i9�n�1E���o������r�.Cm3��>���Z����׾/v����4Ɣy�[�E�3)�[j�"Kr��m�%AYV�+�H���Ρ���u�b�?M�2)v>翐��%SH�!V�z�>Y�㍺G�:'Ԫ��d&�����֩�ryxi%�v���[�>�B�b�Z�	T.���&%p��@؅F��T�z5>�5��y(O,mӈ����`7N�(]��b�]�{�����L�=�v�r�9�bA�����_���gY�(GL�7�)�EY����1���x�I����h�����.d1��(!��c�4����?��Ǥ��w��1�!�R��r&�<M:��I�&JuE�~�
���?w&zt���P��V��6��Og�;m��5��Ώ%~� ���0)�����EJP,�a�+ɬ|~��F�;�ܤ�<�s�߼�o{�)dSThT�ÖmvZsoڪ̒�D�1���fb�qOe����� �3�E�hY�h8'���2�x�P>�"$���j6��٨��w/�P�ƴ���!�͚<Ѓ�g	~fVv@���(�9�/�:?B�"�{��P�e��l����UI�U��tH�7&�����HT�x����H  �Yx�c���+�K�/�ȸ;����}�"��mވ>��r�����$�S�0�o����`z�τ�1M�*p缲^]�&�`<vi��Z�.������
��c֥�����Y�^~���%��e��l��݈�K �	�e�_��Բc"�g���_�C���=O Bv�����sڍ��}�@P&#�/���n�zA��8l���֍�A"w. ~YdꊜmWH�C�w�
�I��c�-�':�%z��v1a��b9׳Q v�_)��v��6?~���e�s�_�O���9�Q';�Ge��^�c�h�D��	E�#�"�W���W-��I�Z'U$��f��~@u������yۭ<�\��.���]ṗ�<�ŚBb����5�?è��*�ԓu�Ǧ�c�W:�7	�TQ#��`����-[��l5��(#��M'��~w}����
}8��{�)�Ev@��a�=�Pn���7@�?�1KI/YsA�j�/Ȝ�qf��[[���(������\�ТX��(g:]��6�YؔA�9{=�*�n@�gR�WY�E�'��.�'կ��M�i�5}z�G��-tY1˺ɸ�7@չdZ�\��ғ�o��]�ㆂD����x���ңz�\l�yO��)Wz�(�+��/�q���w2_����쟞Ƅi�o���}�z��9�)d���-0\e��TZ �Ri�g�ȁ�M�l��;/�ds�
͑�h$B�:�U�8�˭�M̽�8}��s���5���j�?y��O�}��:��vӆS��\1�O����>I䣑X���S�R���bﴳ)}�p�U��~k(X�;�{6�k�l1C�}�*+�H}�U��<`B�F�y2���_��Ȼ��������J���n�5d���꼤L�;�ۑ�Z�m�}��=��7X�@#���a`��!�y���^���4����f�:՚S�{�-!�	�l�>$w�9�/� [�p�r���_�'ʜ?z	�J7o���q�g�w=�R!�=k �j>��������w����*����SG��Sj^�k)leϼ?��������1���b���&�M�E�P�|wbh1�����iCs$�������R�	D��3a<M�BZ��7�\ѩ�Ȩǭ���e8g�8�-�T�b�9V#I��e�l.ٞ��z���^yC���	�h܉͠�
���7��YF���9���x�pQ�q�׳cS���*��(~��+�H�.��a��03?�i�^�����၃o_-�a$~Y[�qC��k�E���qLݨ��@��_�p\[>u
�kD�`���dbȚ�(ώ|��iz����)2#�2+ZK8S�D�/T7ę�y��q�%}�\}�1���"!A�`C#���Ƽ[���T����Gs!�~W�-l^	��{��C���wjf��`��/�D� .1��A����M���`���-�Q�����#w߰�{�	b���e��귒�^�Z\�ʶ�[�����4!EݦҌí��nRH�-�_(�Dl'���!��뗀N�H�y�M��etE����t6�;���Ĭ�zP1=��H�CA�n- 4��W�����K���9*��`��	���%����reN�s�U�l�ٜ�����Pw��Em�1��C5R�y8A�� 8����aT��2�ml}�����	E�N,�w��y����=�ZfP�^�H�"nJ��&��s���5�=6=0�`%���S;�JF%m�֦���c��l�L0���M���R�oj��&QdU�6�P�����s��@��#��TZ_�?� ��r4�-��N��Z#�hT�5}Œٙ��vâ��L}Kg��J�̱�b
ݎ�P�rr5��JP+�M��fU:�Q�L�5I�e�˯r^�9^���6P�a�aX���ˉ�G=`,�qV�-I�@�}�7���u���FM7T�X�-���߱' �XVWwy&�b��*�Ƴ��'����0[N��Ϊ���^[�˔�9����}��H���P|���z�|ִ���
n�N5���Xy5	���#��nD�A��$U1ۏ�Q]��� �}P����U1-�E_[x��;�.]�!��XW��+>�#�Mo�S��� گ���P-u�L
g��0�)��ak9��ݦo�F ���f,�+X�������5%��fs^+��  Y��VT��4a����!Q�#�5��J��=)g�-,+��խ�Ѐ-�cu!�Pe��5�j⼕��"eAea �̮�a2J�׶p�K�.�\�ҮZ���8 w����(���S)���$A��n�*ʄ��W�/��NX������ �{�^ʇ)��$^)�Q=FD����,�[G���������B3����G`�F?'���Vy`٘Jؒ�OZy5L�Ơؐc��,�z(����B�S"�R0�Phd��y3 Re,*�F\�E3��\��7y�*Q��a�x)eV�n��F�G@["�fK�+w�2ސ
��H��R�kA
�\b�l.�h9S���*�ƁYiK����26_Wc�d������ml��TDB���ƙ��fEr����m�
�5��Qڤ���:s�c$�3�Pj(���!hJ�g��$�_��mw��Ց7��=1�r��:���!���0PV��O��%nDd[�Ȉ�e��J<bm'ef�U���C�Q^�Tߞ��uB�@���ẅ́p!ĳ��x�_->���&�7/���y�"U՟K�A��H	����N�@F�Mhg���fh�K���i�>=O�϶v��>�}�v,ߋ������"~:\��,7���ڌ�ڣ���m��xN�����c�L���WGQ�#�?���B`�ĝ�ۼA\0vi�aAhC��P�0�꬯z[S����'�<��D-����)+@�,�ek�2ŧk#SV[�c��p�h��X�����|v(��Q$��7�v]�Κ=t�g|�:#�ϕ�	�$^^��O�3��n����2uo8��n�bg��nq�� ������JQ/kV-D�v�Rdu�m��S��`Y�S��AN*�Q��imK{5 Au|d����!���9mc8�t�?�O�"�H7���x�G|��=�V�{�蒔SF�5f��Q_0��5��OI���ob&��lR��p�xni�%���!q�;�5҃��0��n���������o)AcZ?����2��O�L���님s�tyJ.����P��»0��P ��v&;�	j^�j��-%��o}p�_���Uv52�F�}��f��W�%9%�RC��)pV�����$ɱ���e�m��k���J&�8&����>��9(-�{oٶ�$���U+�;��X!��f���[�C:;+��Yk��]��g�3����vpjk�U�U��'v�1TͶ�c��X��6���&9�ވ
{����MuĔ�!KL9����K#�ħ�\�%�i
.=a~��
��P4���]�l�.!�"�2�Q���	 �N��\�&�c�m,�ɡ�X2��?�A	�iL%�CD��;cr5q��IC�&
�gn�Q���?U_�	� ��)�0J�Hku��̆=!᭞r /�M�6=ϞKu�K�ZS^o�YUcj��H�7Fj[��1�����m����-���Nݬ!T�d�4�1�>���O�ޗ��x��n�6���Du��~��0.�,���ټ{�5Ƽ��8�/#+��t�F?��3�����FLy\��|��RC� �Uw��3�u��0��t��U�[�-� �*>�1
>��S]�$�]y:6��:�.�^M.zT�{���&Rt�B��fܺ��
�I�p�j�cx,�~a���L @rU࣌��v��6և��^�5��"���+Y������r�}��Y���,��}�H��9Ѿ��ۡ�{(1H�ڧ�?���ƃ����l����Q+�fL������;�7�	�2�7ٗ�~S����n���I4��r�i\��k�鸊'b���Ѿ�ۓ
��%�%0��e�Tbጕ:��$�{������Ɯ��*��Qmy��s����_����]=MS����%��_&|y����9*h8�C`!�Ż�ssm��J���|]�t�o����P-K7��4�^�9�w�}�C��*h�i�vh�2x�D���}����>��,g��=�]3��)%s���+,������*���(�-���]^�ӛЪH�ϣ��WE�Y�G���>|k��#�Q ���W�H� rR},K��b�d��SI��Q�_���cR��V]! �� LV3����7]�M��J�`���<��D��jn<A��,�/e�V_�E{ HO�(���ӝ� c;�a�X�N��C�E凐J�]��Ȏ����=Xo�+oy����N�{+FK���:�(rs�F��*�mA���e�������X�iX�/t]t�F||{u~���;�ټ�_V*�L�{H�����g{B��5�ȇ�ݫ�D��g\���9�.�r�Y�C�C|���6��-�� �5'[���H�G_�I��.���a �[RZ���nj���KԚysO��O�r�+ ٢��o�`��YY	1v�N��m!ƽ�����l!��iS��`��"2ӤӜ�
꿷 R)N_��	���Q�~H��z��%ht&����{u
��?��A9�Y���䟮@��x�u�z֗:
�59�|��.��~���1�b�L_��w/ԏl�c�7���{Șv� ��>昧FK��{ʉwYm^���48J޾7"�[=��;���^�M�)�;	�ᩚ��aז����sU9����2cn��h.A{�1:�5��p��3�+G��%|���B���  �O�-{2Ф�ɥ�Ϸk�"���Sm����l��{��!�)1�L�s�&��|\s1���u��#�Ju�]w`�Tfd6��IM>}k8���S�Z�ӕ����;���ך���dtk����?�M��ns	�a&MK8�"�W��$���C��7K��jqz"� Rv��]��aO��UZ�UOO�j��C�kpaإ�Aj�^6��3��f��@���rYs�<��=S�KڧX���"�`^�3���J��n�U���vEd<�Sb��7��G؏�����<�IH[�&�,Z��5MEnd�o2��񥑭��������M����>�~\�)�����C�S��}�^;��!�d����O5�J�^����ƞ�j�aL=�V%�X��iz��y�$(4��d��ɐ�Ү@�SJn46?��&V����n��To��y�0�^5F�\��_;ӂI(`;�Y�����y��3 -�e�(��!6t�M�&]ZE�U��9�(�h���Ð��-�@���iBI.��5��#F�m���µ;� /o���	�I�a���d1R��Q�:P�"���)َ�E,#M��$HV?�~g�\�/� 瓟%�_��Cb�r_�����];�8�@�vt� �숶'�Q�T�
 ��P
H^;}D�Q!q6��*�<U�	�"�í�x�u�	{��Ŗ�Uw���zG�c�Y��SG��+-'�J;#RՈ�v6�>���k�ձ�%q$�L<h\8����~�I�3��<�l�qX�e���F/;�_��⸜�)����a�k�]#él��Y�.
@Pv�)�j�:h1�]%f`1��՛�#�����H�oc��%�_Z����4х���^+����]�2�_�"�b����z�2�-����K;�i�g�=�Ǳ��eXC5y|�o��\*z��ik��n-�#�<�;ECH9�;}��P>��Ƕ3 W�%�H7ӽ��k�^�0�璝g��W��T�GT���2�`T��-$��^����|Ӄ~��@���)�R�F5�>�p�R���zWw�pT��B�g��B�93���<����v�����#<r}�����?�Ɏ��r�7f�������b��,�DE��~C�U���G�����oYx�j��{Z�x��d�f�U*�:$��=�[���J���Uf�L:|m���)|�3��u��3�,i��],u,i!>\��XiT���v���iW��7������1��E�Ϟ���gaV��IT:4�׵��	��mWE�ך�)D�F�#�pՆ�Sϐ�qС^�Mv<�L�S�O�mH�T��S&'�A�`P2#�K�Q�6��g^��(>0��Q���e�_�TuU�c�@�и�r��#�4$�ves*�>���hN�d�ϣ�*]N�i��)#�ň�a]�Xl��k������df�ӳ{��lm��kMm�/_륅&�x�aΌ5�E���}����<y~���*� ��S1�w�s���5�$�f�)�{م.���++O�$B�6cP����5���s��Ԓ��'�"�;�2�*���%��H2�#޷�=�x;	�<%��u�;\�<�����HDҖP�>>In�K�āo`~��H�l4�d�jD������,��m7ߝ҅m{�����M2�(R���Ԯ��fmER����=0,�Lf#������� ���t���c���d{%��o�P��|-i��@��8ـ''K�-s<$�P���}P���X�z�~T�Ċ�B��.�W)6�Շ��=������2&t�0��|�o��,��٪�x/W9ʖW@��e��_���E\4��6�Jv�T�L7�{\ug���/�f�XC����!;{�>��)�����M��9I�pn��jƕ��l���EcEGj�t�Äs�SC���V��Ŭ����A"����WZv��wl\��H��~܃݃R 5!L\+�>�ķ���T)��z�2�@8��<�L&eA�"owN���9�h�1�=�=�v��L �!����uo�[e�ї��w[���*��Av���=b��f�:
k����,Q1/"u3[��[�b���"D��M�+�z��_�JC��"�d���Z�f��h�=q���N��o%�i֥Rb�����_�{�z��n�$�������RB�Y}5N,��z�=���҂yߔ�J+i��<2��A��*��ja-L�h��h�Ţ �v�m�`d'Ό}�x�sn`�2��������#���Z��h2�R�l_��<��^��7'��V�N������/=f�;��p��ͤ�����H�N���4hwQ��_��|"�L�}��֌��R�Y1|�"%�F�9iX�B.$����, �NH߇����M?�Ğf�g�R��l��VV�����E|-E.>��?�ѵ����ѷ00Z.�J�E�>�X}i��hpW�����X0Gu��7�8�7�H�ˎ�(����n(4Y5>Ī��b)�£�w����f)股#�9�(�8Xt�r�C��]��p����.�ݥs}�RB�w"E�p+(���;Y���B�����4�DU'��&%��क�����9��DW�m��:�j����q9��}�.@���v=[�w̺�ř��(��υm����0����=�V�ͣ!^DQ*��bj��=��
�jXv�22	d'@_�xZ��>'�V-�m�9��6���r�+�Gg�/�T#,|�#��{�6�?+\�+a_Vg�I�{��ݏ"��� ���g��qP�MH��.jj]G�v�-�3!oQE�lC���G�����\����ry�2��7㟁ꖆ$o�x���4_�ٶ�8�t�"�wl�bĔ�Q��P�/��G�~�s�o�D���x�ŕ����p2"
)�\��|X�L0FF��Q�'i���=^�;�<!��
���g���4�"Z��l��e�o�N>�p�S{9[/V��}����C�����b6��oj^M�g����Uf�ck��1N�0���YN�fY9���|�❖�^�1_�p�NX�$�����2���Y�ۈ::�9�)Z�0}�D��'ω���N���j���=<e�:e
�m���~,=��al�b��׺'���!��l��	�~K.�������Tj�����w�Y#��6A�r7J���h���#�I!ҹ$I��9�x�B.t��j�SC;��)QG�S��	O���T�:,�ڂ�!�4/�x�ZL��m���D>
�n�"��x����Y�}G��p�\�� �m�E>6,��a�N^gG��X�a��V�^���Ƣµ��A�\b��u�H��72�L���K7��Ӫ�C�4�/�J(��~��W�14�G�k��G'WV^�qgj�;�=P��+g	g�-�qQ�Qa%3`[�?z:�"iC֘�M��gZp��w���e5�c�<�W���b�.�|`�H���W:�%�O2�l-��W��!�P���
Qi��<X0�n9U��ȸ|���9'x�U�#���A��IdШ!��qh.��a�./�:*���w8o�l���Q-��A,��t%��0��~[�GT!�i"ݎ<Ņ���֖�-l<�=K�Fw��w�Jp�m���!�;�a��h7�!�� ��˼w��m0��J<����2g����Y����p�LA��y�䚢G[`�JҠ�����+����Ee�/��_6&�`�7O8|5�%�Q	c���$=�Jڕ��H/hd���I��#ݔ�<��ĭn�T�����^I�Rst́���)���k�/�'Ҽ�_�Ā��	H�V�9��R8�o3�fv|�NO�,���AA�K�!�C�<GL�k�ٳ�
4�F"'HMu :�G	�I?4B�J�.��(�S����ǯ^(w�[�i��Dߣ���~I.����[c~��S�����2�' �ըԤ�g�4OƢ@O��:v,v�9�b�Sß!٫o���^5\Pδ�k�����h�_"�@�K���p�[~i/��\���c�r:�����K��Z4��[�o�<�p�<9�3�3���ٻ�w�����~R�Hɐ��xIڔ�pLA vYUIc�Bp����r?#~#�ˮ�}�-ɜ��g������ȍ�&�]PGധ8�%FzqPU�}'U���..�1���!񞼽�#� ��IU�`�;�M�5�u�X�)#���2���w��y�YST��hm�~��9HtY�
}�b*����6�t+,�$t&/Z���S@)��K�t:����� N�OW��s�/�*�q��*<1���*uɘ(}�k*b/,1b�jR~�hs��^y��֥�,�ez�k<�m�%|�*:��Eg7��&�W�1I�hc��#%M���b	~��'�6��ꣃ�2q��ߛ�����IE�F�[b|�^)��|Aܡ�LK`�����5#j7��(��ב@�8?��Hh���(��ǂ$�����{�n����\��\Pc	-����	X9�U0ew��Cq���s�]���4�X�~�����і7��ڂ���?dP�������g�n��q2.���Bf���fؕB�=]���;��AS��zv���f�hzDܥ�~��3�5��K)��%l9���
������~#�|kg��T2�gl���֯� �������yrlj�Ģn�	ӎ��M�����>ɸK4�����r%����8�OK�3򜥺�r��`D��fE��$߳Ԁt�03�;t��>t����Wl�t��^�r>�� �5R��qrg�ʑ0ݔm��Y����`��a�0%iZ��\����M��m�N���]%j���,��__��M�ݓ6� ��P�&"iv�n��*ڹG ߣ7��J�W�찧���Vj�ͱ����Ӏ|��P����bh�b�͕�#����)����� ���$���vUk�,!�8��S�������ĢT��$��n��� ������|�$��������;�#K5T_ �oJ]�7���Wv��V��*��b:��Y�`�m2pR=y�=��c[���鯃Ͷ���͕ɇ�xB%�L�W����>M^H��\lʗ���o �
8BFE�m7�y:R�v	y����_�DT�!ds���+�7j8���ܓ\ձ�-��� ;�7L���J�)�Ԟ�Փ�`Tߞ���^T��2�kP�zٝ2�?]��v�W��
���Z���[b
Y�:_��1��Q�~�$UO+�Y; +��ᾁ�.�����;qd��pvV0x���{A5�)�q?�}�ȧ1%{�A�
ύ�xْ�k��k�ԣ� t9��<cC�h[���u�
�U���&;3j������|�yqm�htߖ�m�ʩ<��fyߔ�ӱ���1��.4KӲ�?�Y��:1��"�#��\NW�Ll`�>$��7	\�E��r	1����*�%;#��&�w�k8��h�.�=~f��B��7Q��"dHQ��@]� r��_qI3O�����M�:�X��'B���_K�&q�BN�O�e���j	SP%S����ww���vh<��u�N���E�;�}>ZZ��tH�OM�Ч!���t�w�ᩚ�|b�,ƃ:oh���6�e@�%\K��n��z��p���$�s�����]7�?m�=��KU��	���X��eœgٱ�h�3�O'��·��������љ�t�&)��Y ����6[��W�{<�
h��lq^ll�1|S�ـZ�;KHбs�X����b��\�`�ZCV�R����7���@x���JG­}���lX�u�aD���K�e���m���9{0�1�Of��M��=�j��{�$��f3)�4��i�ﰳu�kV�̵{ގn�I�_e���k�"�ͤ���������}������I2a�~�O-�=��(��nw��wּ���Zfl+�%����m������eI&3����෸�ۺ���>���b�Ħ�m��-3/K��y�ׅ'yӿ�|��.����s�[AI�hh�S������2�u32؜w؜x� U�5Q�����T�MkFk���7��q�����Cz��y�!��$)��/63��`�帥��F���@�(<�f$��*M纔{��l�#��*7��PN�<�0�?�2��n�Ugk�p?~E�E)�:����9�=cBL���y�9'��ҌmI�-�(rUJ�J3�����c՘p?�~2	������x�F�٨\/�o>G@o�g��U�g9�ZP����e�P+�3�4,��k��Ճ�^�� ٮ�<����rU�� ֘��k�W�7.rz�� o������6����»m�*������5�R�i˅5��<o�FipT40��v�͜n)p�"�o�����w��	�
�kܳ1��	��6{����ע�y��↱/�8F�il��Mx�;[d��l1%MM�4!��^BW3I�A�Rb���a�w�@��/����H����vT�w<9G�s�ޓ4u����4�}�����5�{��I:+��dI<XzQN��C[�1��u�IE��om�a��Y�sł�5�W�2��h9�b;�bVlq��N�7����v,B��-��7�T��}I�+�}lȽ���,�چy�����@#S�+y~�Ԣ8�$������g����ɼ���}�\�9�2S��Y���_��Qs��w���`i�e�N�������*^J
��_�t�ܿM�4������9df{7s�S}�:�Ă�q�F'<�[�%��zŸ�So���])� ��X�PGt7� ��#�����RV�Nꑯ�BxF�R�����o�s�-ca�s���**�i�����?��^�5���g�7�<��i���A��g{3X�e���ij��$J�1���T2J旘�7g�����O�'�~���������E�N��
�\����C�\��H37�[P�����O��hN?�u]�v�l9|6������^J�B���3��S�d/��>	�mM��2�4�FN���c���j?{��5�%�o9m��l~ӿ�3��k�������oyD�;�!!$�h��&"�Ճ���KkQf[�ꑁ�\��*���l�(9�4;Oa����F�YV��$@�rS��<����D4=��W�[��^j��R�km!����@�
���誮��s�N�%��p)E얋Є���h8�s�	����q��`���S2�m.�uݪ�~W����C�U��n8f
���YQ���J��?vy
��`�%�a�v�|�Q���PZ$t��l�*P��`�bN���_9^b��*��Z����*5�8�R/�^z�ǪoH|:�[mR��yH�������Oy 
����^H��/��{!�]X8��}��P��ӳ�{��aQ�(�`����M�T�0ǃ�M)��;�?��ja���E��63�OVOћҥ[�y��;��B��
 ���u�`��3�1v�̌���ݦg�y���JN'��5�t?��ɤ�&@{��O��l�{q��ʽ)�v��h�|��;�X�׋�8Ε��E���F"�l.�,����|�TyT��T�Xk�Z���{f�<�{�T%�p\����#N�.F���/<V�K�w�s>����5�\V3}���񱋬H����|۱�_�.��֯)/o��z��y��R��9x�����N�����{�cZ�y�,E �'.�� 0�F�V���͆*��#C�E��gd�)o���Ƥ�r���G5���n�B���jA��4�P��\(�!���4��!��Ҝ��sK����Y�J7��d<w��r�w���t��w�4���X
����p���"��q�x(��kѯ�M��#5ܷO���Ǫٖ�'����T�"�_�@7���nZZ�>���:+{��`��(�^�>��<;��b=���<�ϱby�:�G��&w�J�_C�'g��ǎ��BP�|�^��S$N��1�TԿەɅ��9�z�$�2�+4�����X$V��P��h��@2��u�dO������^�Td��_�}^&���i��Ho,����#I�{��ڽ6��������"(}��X�`8O`O��ݐς�4�>�^�������m�ΔA�x�?�n��%��u����D	�%�W�j(��nL�e�vƖÎ	�n��-v��VYoG}-�)Ԙ���]`P����=��УI"ud�FZ��]��[	Q���:Y�]����Òo`�a���'���Ȃg�2�RnJ�)0׷�?��l�!��k �3�Ҏ����Gl�pD�azڂ�"Pҧ���c} ����$׷�e��U�/��[Jf|Y��I,&}�W�*Ed��Pl�LE�`2/������M�C���ps��in���B� ��;p;%��������]�I�x%�jh2�����Y�1�z�#���9�:[~��}��a��~l-�	�o�)�W1_�iG�QF��W�h3�h*jb������H@�΅	��gu}#�ӠQ��,#l@
a���Yr�@�_u��l�OӚ5��4��l4�r�G+ک�5h��c5.�ձf���D�gJ�d�2�Hkߍ�V��ڴӏ�� ���m��|s �fFi����ᷪ=?�p�H�;(�����1��5M [�	E��.2�!$��8M�)��?�d���W���#r�a u��>�^��+�k#����|j�&X��<b;	$n@x!���M�,2�z)�,Z��p>�[im� ��	��V����a��_�T:бk���>�Ʈ���#�\c�K�u�����Xg�����mi�@xųcp	疿����Nek5$X+?�w�z��٣`�t�f�����ӟ׿"we4��}�B\���W��m���v�rP̕{z�%xf�иi6ؔ#������Q��ApE8������҉��UuD�e�.kԧ�Zm��Ӎl�>V=gYduo�)C��o�^܂)ua�v3��1�F�v���u!����x���w�cB�>�_�i��pn�A6�[ܺ�/�K�-�;�U �9�E/�@��_!��PµϞ��=��=v��íWTݲ��WG�c��������3�'Ƞ��)VaN�~<�[Y�C*�E�K��:�,��6B���D�lCǝ��NQP]o��<M�X?_ct+O�LY�8]D�61�ˤ�������-I�8�1@��$�ʋ���F��[}Ą݀���[g��w��Zw�����4�/-`����V���*Eq-��<{���wjM�BӴ�s̠��}a�f�:]3�������x<-�ju���w�'F��9A�y�,��P)Q��0b��@&�S��G�lo8�s�
�Ʋ�k\����`��T��N���B/{�=����0�#W��3e��ml2Z��k��#{�<���j�"=<�S�z�fA�������|fŷn�a�^�����c5�.��ZQ�Nt�X�<�i�}#j2O�;��.d������7�B���>{���!�@m��uXkҿ)�D>3��i�T����8����-{ם���[����M_��!#o����ߧk=�FBbu�M�Ou�z��Fte�����6�e��͸�A�9���\�y�.N w޿fم*�1&!}q�h�՝�}�H�n�"=��]�ʻ�z��~�zV3�)�n�U��6��{Z��:V�%B�ڱ�����A6�������Zx7��M���}�Q/oE���	�'eW[�=�i"��쌾,:�2>��Le�2H�Ի,*Ȓ�8^qwU�:�J�!��׉��/�����n�".N=5� ���npQ�|��<y�{��̕��C�K|-7������z���:�E�w�m*�:���4��&{��i�t���Ҝ!|z�ܿ˸-w)�?׵T����0�dN��p��
�qZ3�,����PVm)�9�ΛJ b9�:���PK"4jP�0ʷ��������s��l�ȼ|��Q �%�z�]�=����{54��[_ˢ`��K��#��ĳ 3���c�*�I\J�G{���O�pe�<!z�'�Q�Eg��N��_�*��W�Zq7Q'�i5�G�[r��b�:I\����/p�)�_�����d�[�B@>N��{9?@4�t��>G��e�"���ea~�����T=�u3����cyӪQ�����1e���?�ʫP1-�1�c��}3S��W��ox:�pe���cb�I��������)ț���_�|��7��z�|1v�g��2qi��z׎�Iwo�o�̶)�
�,ĩ&CW��W���6��
��
��t�Gk_%��6��
t�;ռ�O��ԉL�z������8�?�d�Ģ�emV퉭j��'NJr�W�w���-	�0��Y�|���Kc�fk��_���x(\p���hA�__�Q(�RD�h�"R�e�eL0�Hwx�2���+��L�
� Ƈ�[�SžͲb�E;��-�����Vϫ�,?�D�!���ˡrlQ�b�2 b���i~���!D����� q
��ɳ���� ,rl�Y�|.��[��	�1*XX����L��O�M��:��,�x�L���9��g��F�+��o�=;�b���=n�Nm�4&#�pbc^w;�a�r��K�;@�W:G�y�{L��
v�ȎL��� 3Fm-��ZR�U�"�]���o{P��ZZ��O��Ǝ�^u�e���3���^M��Fƺt`�)�T��cO��nׯ�ܒ�3m�Y'����Q뱺	N܍U�q��P�xνB]�-�8eX�V�B0E Ja��I`��Xi{ɛ�	^
�Em���A�&�눙��R�����es��rwRY^�<j��X����>%��]� �u��fh����F��R�l�����Cŵ���y7�5[��P��C�[-HT)M}�[?�I^���Z����1-!Dȸ���o���,DTnR|����u�3���̏��=˪
A��@'aYK+k%�#�#���s����q��9euX$�,f$6��.��.S�զ�o?)/.�}Y1�Eex�^�L�T�[n��=h��P�����k7E
/�M��>������x�A��-|��W\�y�����;A� �A�w����#�ף�#5Ϲ^>�.\�:J���9��iۭ��^�U���#�%1���>Vٿ��d�p�i�&5nmټ�c˶r/Ǚ$6I@d$���\��S��l��Wu���ZXl�fH��k,X��S&J�"�x���p�ҭ��4��k��}1���^�7o;�UE�u��.?4��"�Y�!��چ_�g��B�*/�(��Ч�_l�6���y���t�D���b8�P|�suP,yޓ":���a>j�c�=����.�W`-�����+�0�Dຸ�=�o-d�l�Ͷ����5w�8+�'�Ф��E6M���|3hpU)��c|��f��@`����,�aҵl}G?��n����LTroQ��`���	;���>��i���A�U���-Ȱ˫JI:s����{]A�yh,\j�&/���Ac�h�~��C�������%a� cZ�κ��d�����.@ L8�=D���8�N"���X["�0�ȃy���A*t@
uƄi�A�8�Z��˸�Z��7_+����A���_�Y��s90w<O^̈�^L�w�wn�4��E���z7 /;�9�ĉ�⌹���C�Pr�;��n���!.�i����� ��!�����J�YG9<��,��h�Jԋ൉ȱ��ZH"��Jk!�V<^B�t5�����u����?�C����*Zl~�����3��N�.�V�r�3Z߸e�Å-������gz�kQ�;��Qi��{%��즣��֚��Tߎ�G�Z��߽W��|S�ʞ3�j��1�@�vڣ@iE��0�M��M��?E\���e,�z-�?m?f����E�g�u�Y��9�ju6�Љm���z�})����E��>l���@l����!m`�s/)j��$�h��	�	$ࡧe�Z�	R�����3��f�%���@G<@y�����p$я63��w�^OS��Js�d㣔C���'���C�����|u_���ɘ��XƸ���v����U6OG���D/���~`�$eqtE�¦ �8j��8�[�F�L�`Z���W�5@#��&V/j��L��~�<�� �g>_�e&���o�b�ۚ l��l:p�bWȚ�!�q��՛��d�ᑜwf�f�oX���-q�i������rrH�Fn:c0����&/t�46���H����vT��Q�*�@�[��eNO[ޟ��w#)T�%��¯M���E0|��ݷkK������2].�p�1,�O}�:�B(Ȯv�=qrN�Ϡ(����S����7su2W��wM9ආ� |�#Bf��X�r�׎�J>��0 @�[c�V:���k�0�v��q��!`:#� ��"��Pu-�i,����='Տ']*�	�? �y�F=f<��I�´VԟՕ%��v���h+���(�N��r�������Ya%�q�/a-��X
3��DɉQ�3���I��F݁�v9��:ϣ�i
�qa`�x��LĤmf�pV>#�x���Z!���X��:� � _&�#�:ǟ�ֳ���{p���3�C~�(m�0M����P6��,��>�������֘��UqD���)�?N�n��{i��{iԽs��4�q�,@���(7Wl2�[�����7�0�>��kHs~1s��+����wzZ����qCp˲�%:%}*</��׍�*eq1�d�<=\��י�|~6@x�m�B�pyl�@1y2���~��ym��ԣk���\F[�L!�̣���iUg��cx*�c"������*���OX �z��S�.5ʏM�O����=v�9,���`wy��;��5��A���n<R��Y��6K}���$����IΓ������'���$��%��W���ECv�Uʖ&��O��5>��06Cf�GfV<���ɛ��"-��BR�����ǧ�zc�K��<>�⒫	�PH���z),�F��M�A���H�h6�(��*V�ZR�(�HnEE%��<�e������u�il��� "�S����׺���і�N~�E�'���d�כ������2��?�W� #�4}��|���
7�:j"f��.��s��> �p�|W�@�w� ��2��4���Z�B��?���,���J���_j�8&-B�����&*�U�hΞhF�X��+���}�Z5�k�E�=cw�4y.hX^_��s-�~BHT]��ʁ�a5�M7	UC��rp>�2�����<t\��bМ:�V'g�� ����Om�E�g]���N���	BSyE.U!�	�#��aq�w��h1�T����"�N���hE$c�ߕ��/��/�40��9%*�A�����#���pCn�ănͩ3����pC<�L����~��ː�u�T�Y9LM>�Ѩu��=g��������������{f2��y���f�P�V6��&�i��%�~�55h� �k:}�r��b}���$â�>ۏȳN��}��U�J�{ͮ;R�˖QTh�����B-�J2�������>ؚ�)&C��}��J���
���1b��>z��i�O�-�%����Qs��A!)@���oS��4!bD�U�L�Ӹ�L"�*�R����$�\He�����]�֙K�#�@����6�%�NVR�!���W�Ah����:x*D��ʛ�ϼ�X�8�ج�s�Tme<�r��Ź�>����#Tu���5��C7����Ѐ �O��֟�49�!��^�r%����bwޚ����e;69�^fQ��@���SX��P⤾�2Y�3ߍ�i�8Q%�p��!y���x\�E���|�0-ȅ�G)4R ��e�j����gs��!%HX��bS�!�.�$���Dg��~|�I`�CBb���8(ҕ �a����V���<���6\��Yrr�>�,�'��jNf�!5]����LrKQ�b����L쒆�����b����d�<g��k(�2�*y@�O���X3�D6�{YcY1�:y�V���Kx�����2�X��l��[BQ�w��gnf&���	@Z�8�olK�)��VKew�V���>LW�k���	bZ�b�~���e���{��5JA����F$����w���M�rv���>�NT��-.�fR�H��K��
��u�^�;��x6�>�j�D���w�`�� ����oymѬv�dq��b�_�
�xȸ�Q��}��a�#Vv��^j�Ɋ�W�)���ś�����@%���.��ܴ��Mxil>��r��߁�Q����Qd�W�@�u�<eo�*��M��`��S�	��}�ot���=�Y�ľ�o2m�_AǢCǷ\�,�>-�g��Xq廧g��G��M �I���cV^1�������(�!l�����'`,��,6�Y*���ys<j�G����13��*��S���FLc���ɡ �z�@M�j�������5E��S�)�I�n�V��+�EX���@�h;����֨�M��[�U��5 y}�7�ù=���.��d�����	䑢�:��{2W~��W���^�U���6'�:ӱ@zj�ơSL��t��.��B�y�?h�Y�z�V�l1r9��m}���<;6��s��jA�� S7n�}����a�/�\�l�jԛ�		�U3}��&��Y�;�W�x��'�T#CCͮQ.�[�X	wO�̪���' ͙R�x)z�w�/��J�}D	X�i�<e���c�9�r�-�Kb6YE���qK��8�5�g#�"��#�F@TE��[lH��J���h2�	���=\n�ⅭG��\��1M'�_�%�c�OZ�5e�L|�M��ơ��wn���Z�Ğ��t���V�bn[�`9 6�f@�an��Ԕ�3	.U_Ң	������'b(뻬�vNR�}:��_����k[:�h:j�a5q#8OW��GV������(�ѭ0�9�	��Nx�@�d��<K���`	S�>�.�Jo�o����r)d&�Y��bxf��{>��;�2��A��}��Z�M�&��4�o��Ǔ�6	aa�{j��h2Yc^���Q�?����.M�b:Ny���X�xj�K�I��O�c���-�i;��%��!�׈g]�b�d|�� @�L˄�><� ��tn*����C�?6���,�Կ���
�4��H��q��H>��M]�!R;�ٱ7Lh)��y�wW8��5�϶��7�
�!蟞3�	ѻ�)��&�C!@H4S��}��	F�G�>窢uz4X�	5�o{�a!�����˭��ݵ��p��,�'7�*��@,�}^��^�ʁ%j�=���фx������@�]I�ʨ��=��-{�Z��;�{�8��B�/ڿ��ʢ�`Cq"��`������Tŧ��T+v,퍒	��ʸz�s>���GDg����	Z��O��t���~��~O�/'���&T�������4�1��nF����ט�.���d��H����@}go����]s��׊%K�@{
�ˋM��,���1��w�7��E���l��ɕO���B��2���2x�0_1�\S�z]�z ��e�1�,�I�!`@P#X��5��[�+Űa�G�`��l���&���ي�[�M�0*�~h��;$�[����~Va���t�'z]�VQ�I� �r������&�o��=::�5�T(���7v���'^�hRƄ4D��
4�7f�p��������R�@�]�es�;�IJr`�[Hx�R�����?��ZQX�*�����X���gN��h���>����ʝG+4}����S�E��F��T�m%�[R/J����z�� �BW5��ѵ��M��r���|3�K`����RMvdi��ѩ��{�~�V7�];/�&E�!�x`��JԂp:��t�U�����J�,�V�'!�c
G3�KS���7Q!���x�+�s�W��o{��ZU��E�o����>����I�!U �Ɏ*�'l��
�H�Y��ب����^@��k>0i"��g�z�%��x���)?`o�֘x������?h����@��D�p+wI����ط<���6a����p����=M̴/��G_��M5چ�h��sE�SMJ��b�S	l����z�sxݮ "�	�DB�r0�K���Ʃâ%Ob��\���n�`3�����n(��hƮ�]>>�!AW�\�]B��ە?v���ض�5�FciS�OEQ�]ߦ0���O���#�~>�l������ V������ q��@'� ŧ���[+<9m:�BF��R�lz���23�N�%yjV�&��+Pt��� ����?�	���N�I����P3/��DK�ߋI��"gS�Op�: �ڰ��f��ӿ4���Zdv�b�2���i_�l��MH.[a賜���э!r>�~��m-*�.��&�')���OSG��v.EɡĽCg�x�%E��c�-��գ�� ��(�X��9c��-4��I�yR�1�A���I3 �9���Ʒ[��o_|�
=�~��ټ+��'�4����B�e?���s�0���	���Ĩ�X�8%c����Jq�h;����0�*�	X$_�d|�ɕ�옡ddk(����y�4+ﱚ�	�n����h`�Zw$��aK���zS��b7�V{�Z_�a4
���"�[���*\�"Տ")0�D X3���֛�n���LK��}H�u퇁��ͤ�Cԍ��P�t��_��gl�to��y��A�=	1�pynD��r�<3��b��R�(�f�b����W����^��)>&���E�
���32�.�T�C�JA&��(�#Y��E�d� ,x�2Ż�)�F�r��K�!	TJ5ng��,���c�T��@5�:��.����$�嬒����=[���T�[Q �P��dˎ�p��h�_�Q�2�{�f���e�Lh�z�>R�j�K�pM�:�dS,��I�r����C�-�bJZ���nχu{�hP�7uK���4�(0�@|*�8>6�rG6�� d��nz�=PDw�J<����X�����y�����h=��Y���Ʀ�I��de���%�ɢً\��s�����d|1���94nZڰ]��,b��L�ky��Plh�sW迪��,��6qDy�e��J��H�#�Ux�v�^I�^��8�auk���[w)�C�j:�Ow�H��_fB`y2��U]>f��}g����^ګ>�����L��F�ҚLv���e،��a��Kk�^��#b�GT��}��LH�c:m��``љ�IR悝ؠ}�*'�(��2��g�}v�([ߨY�ڃ�7�D������o�C$-�LzSj��6G��l@�=�I zu�$�TBږ@�.g(��d���,���+���PR�����D�Q7�o(��D޸8yoVN2��Oz��w��d��UǢ�>�*'u���[;}�`�p�a��8�x��S+�à�%�c�.��N�(���ag��a�Zt�����迕��D�!��L�����p�^�D~K�쮾P�� �z��Pi���u9в�?Byi�w���$0����:],���F(�l.�kr�_��U)LWZm^�jN%ټkW��v�G;	�I�%�I��ԝ�m3�ҦI�#E2)�h?y��f����;�c�Σؠ�Tf:���7J� ��.�J��k-\��v\�~���D��5N�`H��zl���3ع��Z\��+P����6�^�E�}qn���9I�8��UWX�1Ѥ�~�aX��}=�^��-�E������u�t?Ff���G�0������!�0VE�j(W�uO�e�}#�tJ:�ꭾ��

J@6P��RFCp���Y)�:BV�P��)���N�!k
-yB�ƞ�,�#mo^��������&]"����E��N�52*5>��b�4J:���d#&L�t@��Ta���:�`8J��&�.7����y�oɜ�9w���#^��V�=fD���*0��o/*�I�&�6�-���������
�[��Tk�C)�9�k�	����1ƽ��.�M�St�O=l�x]*άDw��'�b6�&%�t{9�/�m�$�ʁ�1���F���	Ϊv��1�#��w_�Z�g,�=���L����!CtA�F�yE=���=C�6ce�v������߄N���l�S�x�/N�L=";k���0� \��)��s���w�Vo��ښ/�LiԠBr�s>��9�6������ť�[�؊��67�\4}�._)�QG��,%#��w���֚�%/�^�g�˱�}�~���m��-A��`	GDuv�S��WD-�7ߕ&D\��N3�}l'��7@D�)"�G�^+;�#�ugj�1��N&O�5i8NL��l�"�t�NJ��2�=����b�Fd�Ǚ���*�t�,�����]j×y�e�W�1&���[]>��Ka� �;��fu�"��!����OY�W^B����#/sn��J���L[zw��v�yun����
zH�Ao�Y��߾��Q6]
Z[�ԧ#������|�pv�XVW���_E�x����/R5s4̱lčBwŴ��k��:j��2���G�>�W�@j%6�'&��َZ=y�rm��J����a�Lvȭ�����cK�N�ھ$#n�r'�l�,�(3cVv�	���?�,�������*x����r�R�)b����� %]S�%9}��+��d|1z$9�A�̪�W�AC���u>R���G�-�׷z9(���]#k�'J�8t�Wq��d�^	�c6�Gd, �\0�e�9�W���
�U+�6��h8@jG�ʦ��'��o�us��֤����)x�Be�K���ߏS��aKp���g�4+Qѳ��h:wq¡\W} K�^�n 7���G�\���=��;5q�R�k��8՚�?]ɯ�6����v���k�Ը>OGJ�&��D�X*�Bb:�`(b𺃣����A��o��_a��E-��G�_��p�Ȯ5`}�u��3�H�APZñ�3�d�#�P���h�y�q��VT�U�~%��h��l���/]ie{�5T7e��+�P,�%0:���S�|8}�A�`����7z�T��3��r��1�ҷ~��"�g`誇RL@my��"}��`�f��}�J�O�"3|}6�d�$+��+u��_�}s"H����xls�zm��x�id.*��h�����4�En_&�{�צ�QL��׻��-2���m�g���=$ߠ�;��i��K��;�cU@�	�5�H�����GL嵴W��[n>L�k�#Ȉ���ջ��Ƒ !b���W�"��a64�G�+:���l?]�w�z|8����(�:��OF��~�^JT*�����\�1T�L�1��a�E�P]p�����(@�t1���V����'�`�5�e�����46�t���� G��Pj���I�zL�t3u�ȝM�كu����x�+�o��4�;� �3����!�Pޜ�m�I��0E�;^w���7�#�jDA�/��� :֮.ܰ���Yes�*]@��-�(s�r=���R�i���m��D3hfO�a���<a 3S��p�8���u̍�������RX{��(�x�������:KѹE�-<�a^?J��ީ�^�4�b $5�����u�$幃�t� 1=��&���̩�Z%_�W撰��ƕܚ��1.Al���������28R+��|�L��o��|�����k���%��8<��h�g���*���|��������$�r�x��34��i2DVI��|ڒ�t�	&�ȏ$#���2��
���]�]~��$�u;r�Tu�����c~]A�ɚ�� x/���U`�*�H���e�2W|�:����il��F�h��%�橷�` ����t�;�'�{m���W�J7����K2{y�B�u��f���EΆ�ϭ�f��=7	�*J�]��ScI��&�;֐!Q�xO�IP�@/�5}u!,�f���ݵ'�7� ޱ1��H���<�DAI���hW�a��+x� I�gK[J�DA?grٌKo"�I�ȄdZd��t�'���Ck0���SL�/+�8��n�+�5�Z��T|f�a�"^��_�F�K����Ч��n޷�k��l�tgG�N�N���
�] �6��n�æ�'��덯�
82ȯ��5�)���|�=��Lt�l[���,ЮQ�{dcU���^�ݍ��w�%O�T�A�*[=��R w���Qd��U�C�$���#�~�l�Q�,d��LP�KIl�d�h+���$�\�n8�Wm_��W�yEtCv���:Q�_�ו���8K�}�Jj�6��p-T6�t��P�A�Ȝ�La�)c�|�y��s���� ����N�o4kP�] �r)_�"FӲ�$N0 �_�|���MT�9�q�[Ȥ�8����X���/7Ε�#-�pK��)Ȑ���8&���Ӛ*r=�W�:���s�m���"]�'�-��[������"�s)���[g�%h(���YY:��VB�_΍�g�� � �X��Z�ɾO+i�9~AN��j9oi�H��\����V���E	nM5��H�x`�.s�S0^DC�W�*~y�;焽����|��¦9@�7b�U ��U��Ecftt��\�)O�`�U-"���H�h�thX_��;�'O��|Pi�!Y�mz�L	/�L\C�C�N5��'���A���+ki�r�㞦�C\����x�6bQ�x��7��D|�j�	V�_�����ͮ�Hf���YQ7ٞ+5�Z��pQ,Y/s����F4,�$3�z�̤����Ir�K^��_S@I�G2��	=�D���5h.��Q�5k��s)Ҿf*��+�bS L�8-��{�����u��?K��z`?��f��������K�Ƅ�1/K�X�Iԓ5��c����C/�v��S*}�����%�]�R��>�qq�ބ�>:����'��b��N���,��zQx��v�G���BZ�D��3�	8��D#��rI��r��P�z�c�^�o򣨞��=Л$v{�/a)dS��&� IH��btաg|����Pp,p1���U��^������*��^" R]��ۿ��@!��xƥ�N5�2p4F����ve���#�z�ƍfլūE��Ҵ��it>�(b�a��Nt�
Q�h���#-�s+�:�x��,���Ɵ,�wBq��a'�N�E!C�̫p;�~���3al��AR�*y�}�]%�2���|�8u�I�9$YB��h.�	�@�k�}8>WDD��@��y�\�#I~���T�O'��C��Š����M�)�aNUI*��[�K����� M��I�⡎	�lY��wNdt*��*a#�96мͿ*
s���׺�p��>�|k�r��q_�,N���Eʩ�tL���*U�A�;�B8G~<��G3���ء���By�	��Wq�g����M��e`���1mx6<�·5j��>���C�L��Ay���,��đ��"������n�~��b� ��m����i�Z�8�y�����c�O�9Gp5c�(��J+E��f���I@2CIȖY?���׭����p���+4�퐍��Ddk���'�F|k�k�=�X�� �� ��i��"BO;5l��e*BZb��ZPi��f<q`Sٺ���!s���������������fo��@\;���>~���W�cW��TᕝW�F� ���)���0�d�30Ӡ-�|\|�^_�>5j������;�O*`g�C���R�^���*�?��`��y��$�@���R���M4�:(�{~LF��>�>ǉ>������u�H���s�ض�ס,�����;dv
�w«����v06[%_y��D��^ܥ��n]��'�i6j�y}��� ����m�EyrS���0��� �����]����[�h��|�֤'EE�H�J�+�<C.	�$����J�$*��.��+"�ek��j���w:9]����1N�-qgܵ�dd<�z1q�X���p!���V&�4�,��(>0�(����ñ��_L�4�z�;��e�o^��˼�O��� n�
�`�e,�/��l�
Б!��fp��:�6�}b�_��Ȇ,Ե������W��=����pr �T�u害*����ƒ?kэq�:Dki��eꁇeM���MN�s�ߪ5}�^�G�_4������9΂�5!>���tN��e��@��Iv�k�`�� Ɩ�4�J�7��4M�����n�<�g��&1���o .�|�R'�X����r�d�#Z��B�r��^�f��Z?r΃eG��}���3��U�nj�<�)7��\s�,��&8�%u�j�V�eO���l�!�M#&��Mg���n=D��u��@��Յ�+~�F�:�(�Z��r��ϨQ�"�ƶ[~"豑V��o� �3�E5$����g�rkfS݀:�ė�pF�����s�-���p�]�,�O�o���g����l�P:^�+}8csݡx����+@B|�G=`�zXᝪa|ؑV�j��Ok$��s�W�gO�pGU1�s�{w������,��-^j����[��W�]��ʿ�H����Oj&�,Ti����2Lt/ӄ����z�~�m>���t��Zϔ�3������`�U��'�<�c2�z�m���p#&��k�1�?2�S}�h�#�ڤ��|�A��h��A;�id^�[�p&�+F�.��Gɝ.�`-�|9�kᑍ���������^��I���,\�*FH�c��w�.��9�T��j�ɿ�x��5kV�4$?��v�<]�������G�������k��������Ĭ���V��Eix��܏�H7�8��ړ1-�ުTC� �Z��������p&���m8�&��}�1�ki���'ot�9�K�϶<���@��x����7�lɤz
��o��z�o[�,%KO5���l�m����D���!Z�C>���>{dM�Y���v=.�}0YY3�(O�?Y}f�ʯ6�s懥&�>R��i{_z�܏�4�~��reH?�ā:��l�o+��71cF�{D�q�yu���Q����`;uI-2⡵�����yY�w��䅳g�����~]�h�)�l�	��BP�)����B���읊w!{ab$�ǐ?2|�,���\`f�E* �6zbH����~����g�أI�Y��:�=gy��U7d��بJ����r������}�O�G��M%)g�Ȳ8`^>���-;x�Z�c�p�o�O���^��k�AF�Nby��@�ɺ�¹Z���+b��p�s�0h��K~#K�ٖ�h���*C�I؉D�)�{S�LȨH�����KX�v��-�����Z�%l�9�]����=vx�R:D,�!3aO�39�?�N0	���	s�ubZv�+�}�O���ǔ�;HZT�\�%���
���F�{0��3���+b��w	�V��Ggm����0��������P:IV�N����ca|��6'&]#:����Of@k�y\v.��k�#�́3U�Z'[븞&����H<��ƞû��Y@^�
(C�^�|s_�E�D��r�ZD-{�+�}�F����b`�/"�=^���(�	�C=��\v�x	!��M x��Q��I�_F�DȄ�JA�}����\���4C�ڋG��7/A�LW�0LoL`ي�w�9T�Lt�WS�=X7��l�$���������2�@9��g���ӣPw����e����QV��^@1>Rc)Y�ٳO"3�ʽ��o�d��dS{s?�3\�����T���D(�CM=��1�Zc�t`C��IX�)D"i�%t��y]�[��~���٠S���n�<�?i("t37��!���>`;eme:É٦����n��%� �{���1�!̷,��7<����״vB�Skb��l䄓��a-�8Z���ϰ���2L�x�ߤ��n�lt�T�1��~�1���L�D�am^�-�$j	[H^��\���_b����u���������%����4�E���Q����K��,���#q�����d���tPw�_�]$�*�>��pE��k{�8�F?��.��0n��v�� ��UF3���-ԁ�ٱ!rg&!{ǃ�?�4�vM 9�ܑ��P�Q�?��}�mP=G��5�k�ݴB+(��	>Yx�y�8�C�������i����d� �����Q�;��8!YFĂPӋ���x�h�c/�&I^��[���{�m+B�X��\&RvZ�rRM��5�b�gW��z�O|��m��5Kn4�y3e���{{��t��t�D��r��=Q+V���{��0��%���{�2��۞C�e�!;�=s�_X�S�BHx[���iѐg"���w��d�/�4��ڷ�#��`�c|���R1hK�X��Zv�3I�7�ڪ�������*Z������e����p��	#-��rQG��{*h���)��U��$�oJŔt��z�߽�����V��Y�������4��a6�k���h;�E����� Z�[�߁�+�R$^)���מ��箁��{��"J��Y��3*ra̓������3�Z�$g����
)fiZ�b�B�k?a� _�Q�-�iA{`e`��_Z[����J[0�R3�ť	�.AZ3>
��n@UX\Eʜ���
���4����&��b�7ؕ�z���a�YpF#�GP��x��Z�D�<B8��.=��<�c�Hn�$͒�h��P�׿I�P�(z���d����O��dYD{�z����`�t����ki'N7�a��/3d�"�~��Ƅ	ڏf3�M�A�d
щwrn6��֑YS��4ɺ�aڐP�~���+-c�U3��/����s>��)	�w�x������f"o]�|M��Ƿ��[�\�e��RW*�h�?&�s���N��l���qj#�`��dU���Q�8��)��C��-c�>Y�?�َ�6�����I��>�Қ%ȞE2>^C/��F���)7���nҒ��s/$�<�Zx�;�D�9$>z�xA���d��5%��P&eH��R�֡�8���
��Ж���Pt�ˈuz���-�m�;1��8����Ya#��PS �R���ʇ�l��.&�B�������M�4!�8�L�v�"��g�<����|��J������JJ_����"AGrC0�F������6k7�D��{��6éB�s�a������h�C�T���7ٔ�e��S!����\�OJ�s���v��\G;��
�ـ{]oXz%�����B�Œ��O�����WN�����j{GB	Z���g�Ic�6r=)�F>"�[hr�#1��=�����N��9$Y�������(ڵI�K�+M;鮭x����Q ֧�:� '$1�X;�j%A��^V�I�G�Z��ȁr��F�跉�7?,��N�$�N�
	�]��|�BJ9g%؈�sJ䡜��T�kѷbS�\N
�"��Z6��piW-b`�}�M���p��G2�˽���y(�Ϧw�������r�4V�6;�3��F���=��3�rFl�r�	 :\}�_����̻��wm3��R.Ə�� KJ�Ky���3�M�����q+�W���#���N'!�j���.'C�S��ęaJy;�h���"Ʌ��R���Y��s�|��@$G"�Nƴ�)�/�����5ՙ�@	��V��Y�)����m����0(�R\��2����R6o�� ��Sݷ�s����L۲�<�.�,����g���S�`�9R��A�K,���wd�Y���>�ܮ��}�[��¬!���O�΅��&�cr|%�e�BL�b�
{�xj)�_�φ����6����y>NĀ`�7�d���.��V�P�\�(j�;��=T_a�/h�N���R�C��LZ= "<y;F21N$�fZ��\~p�5_�F���Q��Jzظ��ރ�2^����
���(��'}�n�h���*��L2�B
��:��9��ڼ�/x��T�����W�C���g�c�eI�w�7��ӳ�~҃���ӗ��<< �����,Oʫ;�����R^ȣR��	pC,�[ �{����樉M�5^q���j#�ұ��'��[���T@�����p�b�� ����Vd�h=g�k��>���$%꜑�;�O�\�+��������P�A�i��&e���^Y%����wI7��\�\`L|	�{Bh���V+U ��)& ��9�4]2��D���y`��)���fvb6�i��ވ������o$�ɒ�Z��]'oˎ�T-��0�
�Cv�� ��@-d5�č6�Me*>`�s́ly5S`��T�/2l{Y绂���[:���[��8�<Ζ�\4������ë��a�R�NP��U`�> ���I���J�
��V�Y�g�b]y�a���i��ԉxKc��Xع,�5 8�)�;��:���v������M�����\�sGdI�tÀ��{�do��É4A���#E��?�?��Re�\i�	�|��yO��DT�=�Bُ���&����p$_���|�f.�ގ�$R�o[�ņ��B-d˻���r��M��Ud�g���CK��+��E%7!x7�N�G��Eň���{l�Tc��=��,�X��SK�VJ*�Ԧ�X��t7�zt�H�r�LcXQ䍫`#���	B�9G	����!�)k��l�2d�E����mm��1r����<K��+wd4�{c��p�J�h� ������]+[x�a�5�	vo��-a�[�]Q]gF>e	�Sv�����~��m�����aS�xs�S����*�����,Y�(���QV���_䋐�W��b������/�C���tݡ;"��Ѭs�ɶ��TL�-j�@a�0��7�U�	�+��oC����J�����
9��Pr�@.���b��x�LZ��T�O�"#�����ֹ�c��� T;����>���4f�U5����77�՜6���N�ktNN5�wL`K���n�">������G��|�1�b]�E�@�J����WHq��+]1�l�n$y�V�z����:~���2z�g�{�.3e� ��D�Y��S,���t�C�����oe���J��?�{,��v�|�ǫɱZ�`TS���z�YT↾pE��㏟�}�l�|�H�:�%�%��$�}��k<�����F�J�@[��ܧ��u��ᾚ�P2W�38���_��RQv�l�:x����M�\h��@��G���ሊ����y0�����'3^�$l�p�ОT��4em�j�zqW�Ҋ���A���o��H��eㆉ���TH�`�!6���pC��p8ksߧ�bl�~�	��}<�0N�y2�ʡtM#���c4f�ڃI�D��=ό�@l��%�v��Z�saػm>���X�Z����W�[Ew��ԕ#T:�d�MU��*������î,1�f��r��s3c�&?��s��Kߋ���N���9O;���ݸ ��B�!��{t�NފQ��b˜�R����c�[�R�)�b���o�Ll�ï�%���4x���bX��ic�Р܋=)F���Gd����p�����<X���{�7f��.KH���|��gE�~Y}����5=>O�3����N�(���Z�پqx��1��9)���Kx[�%�B�n��յ³hJP#нyFl�Cq�O����P�������a�{�f:Axq1���M_h����K�P�>���KHmUs�j����ͬ�;tw0�#�[IE�����)DA��36�R���=h:�S��F��W�+�����p��L�	�L�Mx��a����"�y�4�7�LY��!CˈgHb
5�R��	��e�q5�D�P>|�B�� U7�c�9�T2��-�쫈�
m�Ը�/|���??4b��S��l�T�0������[��, NBL���Woɲ�\�g��V�H���o�2�;OlkZ;��^��Ҭʵ��T��X`��&IIdXO0��&�n�Q�?Ҙ���3�-,��G�}�*f��e�h���/?��R
͡��[G���V�V��ep���bR�X�e>������� ��n���7�����L��z��K�X_���K���r/��_Pd���iM����oC)�'A�����X,swL�$��z� ��X!k���/�ls�[0��������H��m��A'�:g�
�e���9��Ԋʡ�Wr�^�Jx��?ĚD5�V��~t@8�#�(�]��ï�����W5�pE�q�+���4������]��8r������Ro~�o����6I>T# -�^.���eJT	Z���$�9oM󍶰��L�3��h(�]��F�R�2������ŋ�]�����M	˰*4!�k햞m¼�-����o|�A�٢!�}i��@`���n��䝠M�'Cv�����䆽�r����t.���ƪq�>�8<�Q���ǟ�����V�?I���X_��O�(�9�3fb����WRPC��LBA׺����:ғIbIC.՞���쨾@j��)n�.��91Jٽ3���L��鵙xC�� ��v�U�"s~�'�U�ׁa[��oq�ŗسW����Y���@yܝm��A���v�'a4��]R��.B�gH*��ET���P&28٠�'x[�U�C�黌}�_M@gG������$m�5Y����a�#[��'��t��-�p���d�}����^��y���T��қ��f9A�8?J�f�*���燚��+��y7��<��58*�k	92�c�֒6�O%�E�^<���|V?��@�b[d��`y�� m��:K7q����߯����4?*����Q����2�x+�b�h��������Id�˥�����~��ocF��X��L���w��P��\y��:Z� �kG�i��&�A������������\F�z(Q���F�ƺs'JKd���]��:Vi���|����1����_�l�N
|xj�32潲~s�%�/����~鰅���I@�[�4[[~��)�&�귺˧硳�x������2v�._�]�Ջ�2j��t��Ř�89'!M;��O0�a�M^��[��<�a�w��sV�e�^R}�ر���&��&�3�ɾy��);?��>�FO �N߶��#?�X�H�\�L"�@�1�����x��v)�j/�	!t�vu{@�C��(���x�ݮ1�~$���pL�.�	�'���O��y�Rl��C~}��㾜�����w��Cg�Y��+=�bh�����*�}��6!v׿������u�d*�=q����~{Sw�,w1��Z1ŕR	��〪��t( ����~�>�|�:�=�H�}��ff��ҷ�D�'��5���0aaE��j9��~�2Ҵ���P���״����*M��*��nu�|L�rr_
�hE�s�ٺ��b�S����k��f-,�g�y���jXg����E/`�ZR�&NF�P�$���O��8~�Y�T�_���7�ُ`�V��Y)�Z�F�t�������&(��	Y�X[௤A�K^v��5�~،4���la`0���M�Xudbc����z�ɍ���g��^�A��Z�M��
�	��!7\|L���4���	R��E���
GN��r~�5�<~w���m�_�������iX�BǇ�]?�@���'0(�����nt����!)Ue�)Szk,??�F���N�%S�_ƚ���4@��>B����#c3��i�(��>���U���=/�9\i?�5}c�'��?��p��؃���$��ao����\��ȶЭ��Ps�,�d�E��Ԑ�61�m���bH�`�r3�ʏ�!�i�d�^��.`C�[����� tz�u���>#��=ωar��s��͵���B��ٓ�ⵯ�"��^*��ˬ:Ņn������x�(БE�=F&�>
�C�x�`�b���&��
�2�I��Pu(��k�$(a`��.����� �S���x��_�pG-w��A�3;~�����k�a<��A2+ɝ�0�2�Y-��;j{���Y�?	.&x5C}��6�������w�50s*,^-g,��Y�{yc!U�Lۃ	[\�_��ga�Z�W�p�R�;`G��y����:H���S���"_�TZ� Q�fo��P�8G�|<W���0��jN�:�cH$�;���y&2�A��[ٚ>-��H���� 9f��B�`2��[�uz�钥���*��UOxq8T�c�Q�u�ٲ�S���B�Q��B��Cv'{ʴ]F�gi��ў�~�K~�[�?���m�L�G3ʹaMO�8�vq���GS�/.�u���i]N�'��_c��_�/�T���'�q�IJ�9�=�L]�����cL̽wȿS��$>�����ܽ�̶�'�$�Gy�򃁕�Xxߨei� Ć�zն�!���U�\Z݄�2I�4�^b�����D0�!��RU�4�"�C��8+̫��
����a�o.S`��Zb�������j����Y|�u1D�@�ޢ���?V������ǾU�ة��R��Z��e��>�V�>i"��'�^ݞ�GE����~���G���Z_	��)	2e2.��~q]hz:%f6H��x
��U���YQ�P]��zq�k���Զj�׳h<BX@+|�}�%�v������nj*�\�%�̫��o=�=�
	L�k/�m�h�Uj��vN�j$�gjɐ��r.#/~���H��p���0R{s[�04�j�1�>�ãؙ6l>�8�/��oh�������ƞ��O�K��r8ϕ�\�����ȏ��!-et�����8�� 5}�9���J٫b�l%�����K)^�/�ݯ���Sז�|���{ �v9��|ʧZ� �������6^�����Y&��e��Y�Q�Q�����}S~u�'��1��yQ���`�YϱK���^R����c�Z���*%���d��
�z)ʅ��f�����cbK�.�,
�]$;�k�.�$�V�W}m�r�\�"�K��K"s���������Z)gW�H+��f������
J��hV`9q��N�q�)g���(�I!+q�/����;ۓC���c<~71�� ���+}HC�G �ϰ���d熾��Y@�T%P�)��Na��[��ޮ]c��r<����7D/���|�[��P�K�z-8��.���g��J1xT渃Hgj 
�q�qu��M�a���7�� ����ԒyTp�B��4��r��nغLl�n�����z��Vm*�P!d���D���)f~�����r�1Rt��%��3ђ�<������O@*�m��ٱ�LF&�^9ū�<�Y�#�i0#�\����L� �j��qɦ��k~�&8#J*+ϸ{�+Q?�AGi>�Z7�L��H�JTz���Q��ɥ9��ȥ�(���-�w�)V=x	.�G�������;C��+0�	y�� �q:�}"�P�ͨd�F�]��$le��z&�x�I����ݢz���!�F��ntv5�Y�G�깒�{�S�-82(�<��T���G'�*Q���"��S���%��.�+���f��2�qrr+�{3�q�gj*Q���ts��o�e�4_��`3�6cO�#K,�l���)[�1<hE�J�u��QJ<}�P��� ��8i)�����Y�w&�	���F|(_�R6Ӧ�ex�n�1�%Y�hU�!Vd���-Š�K�2��<�=T�oΤR6��	23No�VzP��վ;(���5�I��tv���B2�<������$�	�+q�a��T��zS�2��wѓ�KߗN�w���@B�]گ�g�8	��]���U�*��j�'�����d�ON�M�C�d��x�u�3�	W}:�����6���5V�(�i�w�+��0 R�p���-oDK�y�2�D��Ƴ�j�9����B�zG��f됀;�Y�0@d��{�/�A����[��(Z �ݽ]
����i�B��D��+�*�I�=΋��Ql"��m�޸�A��k̢<�ntHN�y����-#����|]}�G�^>�5�m3��w��Y��~a�k�5Ҡ�*����
urjPލd��r�@��;ݣq�
��EE�%��j���#A�ݷ��	�Բ���U�7f��{���&߮"�Gs���Nu�8����Z��h��C��)n	=���ʛ�q�0W(-L�l������u%��Aa����ڄy���[g�u�!''��2�Wl���´o�BC��gEY���'��[�В'��s�̫�-�'����?>p��{�M<�k%�����B�	��܆�"w�p B>�� ��KD�X���%�U���D���	���+^Fo�&)�Q��̓�Ó�(�TVYs����xz�?3���������-uvF���Z��[_;�'��{Ǒ�y�^|،�W!o��\��f�4f
���طR����< }6�0����k
_�n�f��}Y?{
��,ɂ���h�\p{���$c� �H�!�F+u�.<�f{�+f��F�/�K$9�n2:�o>u���<t�+��/�X@B^r��d:_I0KU,��ӌͥ�n<dxÞn��n���*�_��H�IHW�'�	>�W�T�@kv���Ȯ��-C����W>A�
ङfQb%��p ����-�l}x��p��S�p�wً�u�2je��*\qBn��^�x��:P��6���P6K����W�o�OJ�̙%���k��<[�Q���W���S�.Z����؆�6���I��5ʺ�RJ6�Zu��I;̲{�Oy���>�d	ۺ��MI�9��#���ã����#ׄ�Z�'�h����c}��d�V7R�cT��-����0'�$��!nN�@^�E£N�¾�:صv�����x���k49~A� ��ct���VM4��_�ݝU���A���T9���X�k�
�q�(ԇ�챚R� �:-��2vBN���*���z3̫WC>�H��q�/�HM�oY�S(���~߿��Ly���{,���_����e� ��IJ�p��/�B�d�W��j���(m滴�ݐ��$���`e�R�b�H�.����&�0��s� F?�95�������T%~��F�GO�@0�f�#R�?����W��p39���#�:�d�:�5`���$e(�{c�NA���2*$({�~��`�W�����a�=��}Ш��@?�vk��%	?Ǝ��)�1!1vk����Vm� ;�^cu��LN����l��>�I��5�-��U�0�W�[S n<�Kbo�sv���:����s��;�ʷ�[�W3��!��A6��ݝ"��-����qO"K��D�5�o��s\DK���_nGt3�n�"S�����S��0�آ�Q	K�*�B��f�x�'���?Lk�e>ui��暥�DQ����Ȝ�%�J�ˀT__�6�m�� Xi��{��O�Ekq� ,��#K���RErF�=�0#N��yH���Ϝ x.�N앴���"ɬgrOs���O򾫴�r`e�9 ���/��ڼY�k�=�i
��7���=�I����"�W�]�9����+�P�%wo�/�6RVÕ����q���cfC[��ڲ���� Vֿ�s�v�DK�z_H�� |%�b�E,���#��d+<�.VY��V|��W3	��"��W�KZɁ�D�VB�F�#*�̒�+��.������^��|}���z�d#��bUы�����~�����
wXXG�9�"kP
�ѩ^?�X���!h5R`ADQ�%��h�f�c��������LU�,n�/8�U�+D��>��j�H�m�4� \KZ���yKS�I"�.��}�#��L���u?�m��P�ɯx�Oٕ�p���ǫ��oX"�C� �s��dB:��D|v�J�����H���OP��˙@&�����`��������:�y��z�ة�z��⌏S�����`�@Z�-�JÁ�@��W�������g�J����e�]��=�5'�}2�He��SpJ�vj��
e6=�"�>���D�X��{�2<#�4��o��ޮPCg٣�/}�)Y�,M��̒�D�*n3�5m��j3�Nݠ����'�76r�lɺ-��ANu�	oʖ���D��+��g8Ж�����2⹦�G����/�Xo�%�4w]�,*.�<N��/{�ԍ�Jb?!1���<���%9��k�M���lrN
J����T%�����LL����`�k�v�,�0�yspa��v�c��ʰBÚYv�&]�֦��9�֌���B��yH�[56^@j�z7}kZ�|�(у��� ����H�#�$N_S�����^*)bV�`�P$C�t7�M�y�w�����m�A�G^;���9}����j�!Vo��2ߜ�c�b���:��]� �I�iq� XDni�/�[�6V�5.�M�独��:�m]��=��xn����7i���o���K����I���7�v�L��$� k&H�)��d=K-˱Bcaך�V����븣��!�[�$��8�]B+��5���-�C�=����	�.�p�W�S.FBy�(	Bo��y�Ӏ��o�d2ßS&�rdt[�E2�Y	qM�����
[�����g�TG��mIf�m���r)��v����}�ٽ�N �Qw��3��V^�����F�6�k�S�aC�o��H��N[r���@����w���p9��	�:J���v��V����q���x��A����a�k�}iI���On�X�v�  �:�E(���b���2ƽ�{��H��v��B
�>(�Ņ7�J�'���Q��q�<��?+�Q>�m���O��Ļl
1���l&���k�� \��~��H��z��-��#F��RA��_2�6�n��vwq��.(�8p�I�m
�r��a���"���ēH�;�F1PO����z7՘Md:r��^B��Y�~���6Q��g*�>���Ǔ��6�U��M8@@R��,���t��դ��a��P��>�,�14��r@�=�>Xa�d~B�lcn�o̦=[)]���8�Z=R�֣>�Q�I����ם��^��e��a��A�Q��vĩ��!vl��K���-�ʰ����U�h�AwL4ΜüIg�ؑy �,Գ���`j+.��}�f�9A;g�����:��{�EZ����\�����8!���^y�$kOOd@�*,��O��i*f�}�6�g!i�u�7�
�xm��Lg��E��U��c׮������]�.���]cT:�n]C%���3��ꪱ�1�G�p��F�
�3����0�1�����n��8cd��\*l-uT�>O�&�E��םcz�_,A_����(ή(ƍ�q3���u�~�o�5��P��
ֱ��Z;�I'��s�vVe7�!���bs}�3i���fZ�Z�cd��dM���m/�`�|1�j�	~B{��B-�WZ��ru�������,s#$��^x���4�H9.���w��@�q�n���m��3$������"�e�WL�f��j����OO�M"&�C�W�sn1�D�%���03�!3�̏�^��l/��,t"�6&�OP�ƞ�g�@�Ti��>+� *w�ֲa�!5��� =�C�Ō��(f]����,���W̯��a�����4�1g�X?5��پ*�������;�a�C����ܜ7-5Gp=�چ��~�hCzK��iEZ>A5�J腢���ڙd{r���x�XN��d���R��R~�ݢa�J~��͞W��Y�V|�Ϯ�"�~(5�ڕ�d�:h��-W��$�A=N0�O>	�]�5�RDw����t��ދ;J����
��`S
��A��im�%�#(�9/U���aűM�#���9#t�`���0/�[rfg�f��woފ</��S�^G ��f�N�����`�/�y� �t�$���W�'_�K��H�R���)������*�S#3TI���Cכr"Ăc�:)���P����)��"�<=R���N��]�g���LL�eN��-zp��&�K%�lA!P�J:~�d�'�7����"
sʟ��I3y�
 ��6��g�²$o��x�J0F�sh�q�?���t��_V_�`Sl'�s���Ӄ���l(����߯(�f!�ݼ�|ϫ��m&x Ma�3��o&�����}�46�ej�j����zAU��Uz͈	�zJט�����P9x&��	���ш�I��Y��P��=ܽ��TsR�E�6H�ͽD�ʁ;U�E=�Z*旟	��=$�^d�G���2A�-';d��1�9������S�\f- "������]��
�7~�NÌRDi��Wu}��BR+-����V�ɨA쭍���yb��_�X���G��ۅ�R\�B9�7ic��A-S�	Z�`d�����Zt����`SKp���d�7��Rj���޸�k
�l ���3\�/CJ��\�:=�:l�L������^1 ��9�ph����
��<K�qW��Pqq��jv:2�z�RX��A[�*Ķ�"cɉ�x�GH����8���wj���ޱ���c � �4)h�9+���"-=u&X�4H��2�붺�ٺ��۴h'��(�nj�^�S��Sk��9��A�rs{~)���4�v�j� ٷ�^����1!&��n�|\Fԣ���,�ۂ�^wh��~X���#��c=��M�̬�7Og/FZB$���w�|��� �grR�Q*G��ib#�9� ����Ix��}i���ǅ��f����o�U�3��~j���ZL3g�I�W�%�2oU,qq�bǒ!@>Z��`8G��0��N��ҤEp�����z���N��v�h;ы��찝�N>�Tԣq
XT7!��*t\R��K�|�ܙ�3Ǟ��� W��!�u�a�2�K����\���*�`�&4%�=5���J��s�о���suH'�E���<�HS�ί\jP��wğz&"">2K���{i���%Ţ��U7��ȓI'l�(�6�m�A�����ZBR��C��\�����3\����k#ӡ�.�}^��c�jŌ:1�1�N>2��B���{ԝ$D����gD�Yݽ�>U��ړMZ`-|R��x\�@��ǟ�r��(iwk�7INBL��a�d��V4o�X�V �~6��,1�H(�8���ڲp&Th��ܩ*�J�R�f_�l�Bqy�:�EɁ�~��8(=��XT��f����q,��67�o�~/��8��f�75n�4W�����ܾ!Ʈ�^�y c��c{��;�)F<.������/��nso����!��iV�E��⾙-��,J��*>�@_##ߠ��w�۞��3��-WJ����
���Y�M*�!�&<7?P���W�G���ʝe�8�m�2�9o�d���?Ӹ�n�JCuh=��h�Pk�����㞒<d#=RǖFz�~�o�=���|�+�J�����dqt�$���B��k��v�&�;�z��=��B& .d
� :y5�'|g��#���Z�%�Hږ�)�fm�ER�	��c
���a=[joi�&rZ1Y�5-CJ���ܚ�\>a
�,e\�L�G�wT����#S|��
=��d]S(��y��"����Y1�u� �qx���X5���5�^�?���s�}g�(�H�ô����Y����%��/�i�M5�%���w���M�2kv�N�vE��Y9>��pb�_�΢W��$�8�6�ƒ��-u�X'��:!'~�V�ʼ�/p��	(z�A�2e8v
���'�6�tN���m��b0��a�4�\�����~�}��`��F��c
�v������6�+����ܭ�5;�����ؑ��3&�4O��aN��g�əL�*���4�?D�:2����^���'+��Z�E�N�?�����dم��bKm���V�|�c�f3�B��h��+Q�d��+���E4���g�Z!�� �X��IK�:'6�{��ß�<��������>$�r.�k�����b��� � �M�"#���m���K�X�Hw�Y#�	6bJ�O,�)`]�"�����n�sL�`�A
��}Q:)gC�V�C�U�Ϙy��-��y<���f5��j�b�q��:���DG�aph���0{���ዢen�Q���ʘ��[ �0�^����N�=��nϱ�岛���%�z�o��kvh/�����@h�<�M��]y�5`��r
Jyi+���e(��������G���zg�M��X&������iO�nt
�S��d-�Z��R�Ƙw���*]"��� �`.�c��F�@o�C7��T'e��ws�y�!���[�W��h'z*���2��L�����`�돞�ٖC�}֮T�4w�/=V���1�q��?��ml�ރ�SLˀ�!�<��'�N�ρ�`���C��R�6y�~lt�TQ�D�!�����X�<��7���C��>g��9!�I���~���X[����j���E�Gd(	�b�ح���m
7����;Rf��(����JAә2�0R�����<�ΧBKs>�	%��r��)��8ڞ{�����'D�rP�OAsz�@F��60Q�f&�J'/'5�4@?�[��Ctx�$n��YHmD�ݓ�� �e��qL=η�D�lg]o�?�-�<�΂E �k�[�W\�d���Bf`��v�U���"7M�:~�K�>uE�J���n�h�L�1��,A�:�"x�kx�g��6��A�$XLlݵC���bb�1�cd�b����H�u��i�u5��ͺIELDrKU����ϣf����FR1�(dl	8���f���ι��,�:��?���2��	(�@ C���v���T�/�����`�y�>�ʚ���r���`
�p�UCk�k������Ǉ�'�]b���T������-�n�[!n�dF?T��jYo8K	XV�ب1��E�;��^�n+���礠������� �%�4=���@�X	~� O̚�~�k.HI$DL���;�� �Ŋ�Y����<C�\��l�t��"����!_��'�<��ے���V����U'���Fģ{�����+�zs�|���G�Xt��;^���f<^f�!��̗_AA�~U��w��X�z�7���K����4m����@#��ح������p6&fs=K���4�N��]H0�.��G\��Cc����Gxy�}J�����+1�Rt�ѽ����x!ꉣ�(Edi�+���ޙ��!~��y�g�w����pr~1�lk��&`W����Dު2HT⍶��q{�6� ��`��tn�
��YqZ9�U�m�{����赋���
��-�+��E�C:�b%�K=!	���^�]�8�����J%݌��I�T�ӥ[�����Q��Z"`��{7rEo��f.�9�|{�0�����СI�Y#Z2{�Q�,��I�y�Z"&�E�j���bd������QF�����eJ�Yp��<��D�"m�+6(7�@dEA������h���u������p�nUA�&�Τ�M	��*|6�t)����1Yb�Ҙ���#����k��i�z%UzL_,�υLB��|��؟�y�*Obu���s��!�}��'��X�ӷj|b��hw����X��3X�A�Aҕ��S�ӵ2�4���PH�+�7�4���m�+��\��� ��"^�^�K���
;��g5E� �t:b�2e����ɠG� o���)T�R�t�4���# �-�	��]>>t�a���>��}k�is�=��b�l�-����)c%�9F����\N�!����X�I��(窔=���n�E1������i�֐x�9��[������ʀ�����u��B�2�Q��^Y$�j�4IC��[���)00�!.:��#��c�F�����/[�DSǸ�OoK���l�����0�RV`/�i�=�
��JՈ%X�>�Ȕ8��7 ��N�����˧p�=�M�v��1�V�J�(�fG��0���r�ʂQ�'�%a�E�L���iQ�;�Å��CG�f��^'>1" h^Mh/���u1�Ҫ^[�gr���=��N�b�yu�����ؗ57䷼��˿U��SZ����n�(і+��/��[�-���&3Oo�J�qxĚ�F����o��{мv��,A��A Z}�(�f�����2f�ʁ����*��䆧������ܽ��dl��1.P�� ,܎��Ҵ��̀�sj�?�N�q�<G���4����-=�%4}e�}8h�n3o�p��B���F���K�E�r/wJ`i�|����P��-.CG,�y}���Рy@�_O����)��BDkbϲBd
�BJӢ�k�"W����:����y���)
uw���BD��$.21�|_���F�Ϛ~8��~�0�s�8:m~���>_V\ڒ��:���R-�臕9zXg�`�Bj	P��.ڃ
�0��bF�H�6��ʠ�����V�l�.h˛�z�� s����!�؏��W-��ുs0�0f��O!"Z|,�t(�y�������M�3p��ý.�Yn��D!�=ӆ�Fp�\R �ZY1�c�P�`�II��z�[�x�)�#�o9�7��Ơ��1���u#`M���e½���ub$��?��Y�Js?�Y�s�==G��� R�(���XD<�E=Gf��������b��Y�kxbH��/J\*��b=_;�]�
:z(�t��Pf�-��*+�v�琗H��Zdr����AAI|�R�� ��: �a���fQ��MQc�_�f`k٦��1r�`�*[���~�:����~I�dcې����`Mک5�#nt�6q^�E���1^{*�C\Zcя���o�`�a@H�v���3n�>���%�<��jXw��5��,���w?Ԥ�EF"���Q��ܤĿ���|=>i`L6vU��1�V0abohn͊3�J����*$�b�! �4L�T� ]�bc�t�K �4*A�Y	*�M%��Ov��	�Vԭ�+����:��Yٵ.��M�$ծQ$�=�|����'�(��"���*�k0Q�Q�9i�nV���r�A�m�7�z{wW���0f�+��j�,�V;��h�9M�㺩��g.�?y<��7e�)*ъ���Xj*�e�kJ//%oW�p��%�
 �-g@��9���m�kN�0�P�Ě>IC�h�z�ɩ��O1�����ϋ~b+<"c�&Ub[�����1e��+:D���#xꀬ5�y��yN�����s�Xrq�$��8j9���̰n/�*�H�����%l'�/���.�K�XRF�	�����g
�5��":�>��#��ڴ��hf�阙���:R@&�9��s����߬�ԻL	Y$j�s�k��H����ݱS��{z�=���rv�H9}f��a����� e�Ĩɀ�����s+C�OV�!p"$��5������ޓ��7���>�@��7��H{�UA�b�X ��tpP޷���MiZm���+X��N�C�iQg�.�/=z�/�68�lg��U.D�u&1Nk꫸�����U�I��	�E�j���ǜ�p6	�(/��n(�l�z��P��(�׳Y���4o���V�(M�L�����xm%Ј_ϵۤ�[���zb@���!�S-�y�N��A*���s7���l�a�!��.wUJ22-?��n����v-���//��3���['��v�������'����KǏPt����x�'��8�������sy�-�(�a�ȃ�n�� 0��� ;�wh�I��hU���4"Vd�0��S^t *�m��P�FO�O@#j���{���9�Qп�Z���̤�+"+�Wm/�~��3�H:�=[���!V�f�߼�5 ��	(�_���:E�~n ���aB����{�Z��V�9zo����n�]�,2��qf*{�,����K���	�ѱq���$wS��`�۠���"N�r��q�!ޜp��h�X�L;;Z b7c��0%���\h�f�CXJ!W*A/�ş�W����G �2�yF9"��]��8o�\�c+�r�������Oc	fu�����.���]��������qn/+kw6}��YF؍���(ܳ:�m���`�N�PYm$������۪o
VJX?�=�I�yn*�}@~G]�B}N-9��p�A��t���� f�ټ�e�� �9Ǫ\���`J
`�̲��)znPz��50��d���B�M?��g�_tJG9�#f���`y�vU˰�Z� z)G!F'9�
}:��
v̟������nI+_N��j
�Oww�w�!I����f3"�c���K<Br,��W��2.!8�/��X(C�	��i
�l)ё.O<���b�+fM�L8�?��G�$���@ڪ�n�Z�k!Ҙ�tA)͓����?����K��$�Z[%�Dݴ:�!$�^���I�ֆ�^Y�2Ȓ�����$���i��I<rj� pWV�v�3�o�v�^����G�ؑܿ%�&���^��~�����z.�I���OgG?0����Ξ�,������j[uu�ѯ	G�ZyS�E<�$�����gB�����ˉ�����T/����A���{D@A�#}�o���^�vn�����^s�-׼��wߎ�sG��4�5&��w���F�����j�B���	F��;��y:�~p�~�y�J8�m�,�Jd*> �؀I� ����@9_.���T<(#�mGa x���SG�l�'S�
n�
�@�w�r'+z�3�+F	C	:� �$�2��L�+�z~E:���{ȅ}��KaR���������ę�6���|ܯ��y�O��b5,�>3M;1�L�60��q.T�c6��L�!l.n�rN ڱ������͔�(�k��yK�gU'LЦ`w��$uܶBU����Y��>��c�ABR�#/�Y�7��(�������q�]+2�~�h��yBi{���2��
"��ň4�1�N�E���c��k"�=����S����F$^U4��:d�u<�DG�X�<��>o���`��O�k�c�_MT��������@�2tE�GL�������"�h��.X�����zs7jQ���.aG��4�ߖ�Z��^��	y3�k�������{����-����qE��1��K�j����M�><nb�L�E�&d�N�1Y>�굟)�KF&��_@�Vf��"���0�{�� V�lhi^�T���-C|]�	�����wj_\�����H�|��ӈ����_?V)Gu��a�N�*V�(ԫ�.<e.�S���8#rw�F��,�2���o\�!d��O�]�^w\J&��N���J7U��1
(�������"����p��` �Y���	�Kd���=s�Fd5H2�k3����SÔr��,~����F�sX.0�Ƀ��̸c�i��g�M�Ȟ�y�ᘇ�v�볜������t� ��_M�u������$v�������&�H�Ӛ	c/Y�'_+��̩�[<E������(�����o����6��������T3s*OߞXcDĉ���wߦsZ^����<y��X�޵ML�%9
�c����B�4{Q�G��q㸃��1F��22 }Q&|F���БQq��eʏb��۴�Li��:�xza���L�p(ڞ@��Ig�A�q�Ԝ{����#H�T����az2Θ���U��L�@~��Ay@-\�ŋA����T����PU�lC��lzw!+��c�Z�Š���f/�e�͡?|�z����^n��ȯL�ɞ6b��&]Y�]#�N=>���<�Ʃ��J�������}@$�Zm/rJ�2��qD�t��4��{Ew���xq3>�����)��:�B餶�NXF%G���>�?L�P�ZX]������Y�W�$(4�8X�P \J�;��8�*������)��^��]�77�`P,����C4��Uά��Bk������Bm6P5���(V�z���J�AR-m8	��1�qu����q��z�o�-W��� �����������G���D�	���f��X)tR�����ŗ�g]�Q�L�w��dOy4B?�qJ�vw-�x�i՚w�@�)�y�!�-Q#�����/-eƛ�nn�$��/��OIk#������Z�+c�mD� d���Fu��Ue�Ǿ��pO4���\�ߜ��e��0�Z�C,���8�\$x�s�L3�!�U�B��2�E0�t&׷烿!vW_�ő�O`nnx}��`N�2H@����"�k���?4u�]�E�:��5��� ��|�1������W��!@�� � ��K,�a*F��v�p;F�~�w�%�gF�.w�@�Lk����f�l�(2D.1g7oi�J�5�M�`��p��O���qu���E�h%��(}��J��:�ˋc��73�i)�\�+`8��vC���D���Ū���~�*w~gfM�l��|��1��}[�)�������j�B�1�}����g����,4�������c�s�����dF0_0�|Sh8����.�T����G��Q,�WP���-{jL$���� ,�G���D݁Qz�T?��]Ey@�C��n��ކ,A��w��G��V�5B<H\F�����=bXi�j�	���>Q8���A��R���͌���b�q&�e��8u�#�k"0�Əz⋆e�s/SC���/��]]%� S��CQ�%W�\vȷ���Q�~Ti�#�D��@
�d!ew����+\� ��(�����G�����" *�
�
pT��Y�$- �|b�F�吂�9�ܦ?���t-�ʑ�S�p@h<�a+�R��u��x��n���C:���˭9�D����:��?��XII/A��4�x8�$4������R�k����D����d勪�jY	��vZˆ�Y������ E��V�,�#RmN�/����P��N�M�D�݆�Or�C�4����7�c�a�2�EX$/f�� D���k�*�5��0j�a�;e|ßI��F�Y�-3a�ō��Y���	������b�M9'���o�:�3+T���\C�Nq��Y��v�������Y�y�]^'���=�r�.8l3;�Ƨw0*�)�z�K��^%զ���l�.I^��}�`���������%'�ȭE.���Xx�";�>�
J���-�5.�*g�m���(��L�!�p8�wGc��W��]ݯV�g���W:���o����u>��~�����Ǖ�u��!�>�D��NTY��٩*T��+�XA�Ԝ�kŗ$��i��4]<��?j��[9f�<=Z��6 �A�C�����A]s�`���I��m��
��s K��p�ڏ��(M�0�ṙo�辭��#_�p٣ǲ/⁠�[���% >)�����}���"e����v�;1�yw�U���C��= ��6�6�Fbu����#���%�44"Lj���S(6�&d����w{_��������7�uJߌ�~�Fi�^/���X1�cM����l�k�R��0�42a��Z��>H�<�оd�������.l%�����d�G�s�YC�S�L��q�mjc���O�n��N7����g>�����(�{�J�>�|sF�]3Ɂch���=-ѿ�����G�1�)P�ÒhN/S�MX�gXy��FI�f�ݞC{������)�v��ĕ�q���,Y�&���&�]����(#N[�� ��7h�W�+�=��'�d����J���R��)�������R����+�C�c^�1{[�3+�늘�s�T ��A�RF����rt0� a*u2nHMg�� s�W ���1e�M��� 7(ƅz�r|5*�8C�J���KM��.��K�J��^�m�хp��ɍ�� ����~�c,��/H�=���O��#�����	�*c�ǹ���a�,�%5��/�eW�x��V�c�
�nhAe_� �-o��!{?�y�bd�q�f,�&��:S�v���&�C���h��3�f$H�Vn7x��_�~	��iaήQ �v�>����"�!��;lP�J�����r-P@��b;;o:s�R�7���Qlv:o=�ì��H��u�"��$��gP��n�7��a��� a������,���0	�Ob��4��z��Vm�$��T��V��^3�1pM�<dyg|��N���6��6�s�.&-)��2&��Q��Q�v�QY�i}gh9NW�󣧵L�6HӅ#�K���}�W'�񮎴M�U��j���+�qO%� ��13�.���X����+���3����o�������]���cȡ�M
a=�j�M��u���)�O�Cfe�Q8�A]Q�w�,.��\qY��$Us�Q�9:N$nJa�#��$���:���0��2ė�U-|�\�c���XJ�s�iT	�v�u#J�I�����C�f	֬��Qg7^�ê�P��ڱ�
܍"����3�zV�0�s�b��锨�+g�]�-��-ߗ��T��&��tз�\��.k�ޯ�M��-MYLp�?��i��e���~$�pb:lgՊ���b#P�#�*ؔ�
ֺ�W�S�#G��g��T��~��Y[��_��k��C,%Y2��a�y'w�Lp���ke���
�ԟ���e�Eۭv�Htn,�4�2�F;y�*�r�������O6'�T���7�e��J��L�˭��.q����nZ_�&ctѝ��֚/��-W/B&�� �K��d��\t�
q�*����$�f\��ww�j��={bPunH�/�\�V��� '"���e��}��c^!�=��>?��S �xo4ȱ>r�Y����O
��udҢ FX��}�Éa���5Dz�k��gՖ*�L�Ą'L�D�<_�����XW�޷)V���@c��)�ewk.�����V���4�;��!��̠��ۏb�V��oԲ��X֔��,eIV�[���Ya4��R1��#�_��=ႂg�X-r�<�����j��f���b1Ce�3m,m;�U�0�����*�γow�Mg�/~h��,���gmH��Q�q�~�Yzuhuwz���T`��X�����}A[~�4��?p`�}j �0�[j�O��d=����,BF�c��2ґ��ia���?�swd�
����"�QTּܴsc�e�'��H�c:��b\��ަ�'�x~a%2@��Έ�8�"�Ix��Li���0X�"N�Gt�qfh�3l�݆�5�A�h�a)|��1R"�=�g�V>q[}pF3+57����]k�W�U��0'�7\-�,,&e����K�@�����"�`��(�����7�\�1���uKŸ�h;�麷���$y�v��'5��-|n�0@��,�]ʷ	��y�6�ی������8>t����2�L��t�r���k�_�n�E��h��x�vM�8�Q6&"�eh_z�>���ur7d���+ùy�p6Hp0����ar���S��C6Y���������6T��g;۹�u½اD����<b���#6Ό�rVN�ԒI��pb¼j�Nƾ�1�^Al�Y��%��L��|+��<��d��|Iv�
�f* ��۟���p�T]���G���z����n���t�(�%'aU��si,�L����p=T����[a��#U�F��]�s�7��W�������c��^�+�1�t�h�}�%\��� �\�ŏ��=0\� C Á�cE�w��5"?�P${$�&`�o�!4g����ǆ���!�d]f8hh�۫Ȯ�=�(%l����p&��l��)����W����d�cj�(t�{}��<�B��n�Y�?�%��b�@!o��hn�H�Gb�N���d�D]�H�|�DN�_p� s'Tĸ$L�v�?�&vɭ��y-f������,�u%5�W�h������3/"���1g�7��h�L�2PߠhH<g�c���hPcY r�ޟ���X��QajǤ>HS���� �<¥�� �,ןɯ��W�r����cv��ׅ���8�����=�\+���Jy��y��m��l�Dp���W��Nz�;�:�\�м�,�w1���_s.8!�m	Z��nGh2�&�M{F����'�~-x�Uf�XL}RV�[���U�`��}�e��@3�[��nq�a����i��~�Y_�������0�Y╜&mTO'��q��2�s��\�f>�+q�;Ԥ�PTm�$���E�	����?��'���2VV�Dj�w��H~�(��a$���ܬ�V�?/�T=[<�����A���Z���	菠z�ϡ���� �cQ�q�k��%���i*�7�������:v�w���~#B����p��q���#�+�iCb�9�(C�!��z���Nσ��X�9����A6�*�C���.�u��9{�G�B�w�n:����_�����.�GgFU.m�P���w4�r��U_Rw���x����*5�(�Ƙ��f�n1��N��YfL�ǵ�8g�Νӿ4i
�7���
չE!�z��u�����b����ʿJ[҇��up�擅�[�$fA��K��.�{d�v\��H�����٭���n@�d7>[lN��P׼E�Po�jT�	��!���{|���2^L������=��g}��v���h���8��E9�;�v�@r�䓻�4���x�a�Ҳ�MH�$zaw"æm�E�h�6��e��יD���9� ���h��n��"�o�"��􅩹���`��������XAM3�Q��Eu�0�x&F���Qrd0��1F�q��3bJP�����R��:;��h�3[k�7�]aS�bE�����'y���Y@nV}�A5=z���_�H>vz�i�̆'��C�'��F.�e�R�-#}r�V�N�6��a�|L0�IdpA�_K�yl ����~:)��/*�(8����̠p��Gi܄s�\y��tVB�	6����H��(����2
��T+c����.I�X��'\ *�K)&ڀ��`7��ІĹ�zt�࢝%.��^�� z��ґ㱳�2&��wR��Y�'����ܦ��s�զj`8T���㭏4��&[}m�IQ�`/ ��j]�̸���'oӯ���ۘ:ah:�KM._ٗ
�%b
FU�Y�)l��[+�Z�t�K!�tc�5��e��B�{�rJ��hWo+����I�_e
Ħ�})�ȓ��k?t�N�}�5a-��ɻ�R�>�a��ɏ��3i�B��nv[LI3�h���E�tC���>e�
�N����oy}�e��{���ֵ\:���S������ �*��D!Qj��-��klk����u�"�%X�N�g��)��N�#c���HA�#Z"�Q����'H�G�X�/f����҇�eˁ׺6�6�e��D��PO�|���řEZP�ţ��Y@wH��Eq"���`b�i��icl@E?��5Ȅ!^2{l&���S�P���-y�<��b��_�d���]����,LCO����������\@!��p��'���t�X@O�.Jީ*s^�����c�<�-T�G#x#P��}��mh���onnv3��ˌs��`{�Y#��Y�R�Ca�J���v	
�\E�MwyU�6-��f���1%��s��?<8���:���#�.U�[�v�oR�7D��)��e� ���	ޔ2̯�D&���`�r%��C��H�}u[�7��OJ�g0�T
�v9�\�Rn�w�hr�]�²5ݐ��7J[�3H%�Қ�W.��:����7�g��^�#ڹ�O�<�~2�������{'���C`N�4B�á����`sF<ɱ��1+�ƻ��{�^1Q�� ��ic{�*z��5�8(�<i2r̉�h��{s"�����{vɌ's���`�����l�ԑcŋ%�g�&�GqwO#/
?�44Ǘ��M����5�GIyG�-�d�>�!D?逹�	o�Z�ʖ�#z\���1<a۱�\`�&��IX�x�0F0=id�[��9���=5>>�*ud�Z�ݵ�����]�%��~���*l��Ni}��)�/��W٥�4H�� ��O	Gy%��n�G��G>y^��l�L'ٔ������m�#�O��s��b��y%l�)}������"�S0��y�gT%K��f�^�=�?? ��y�E�����ϙ��h��@��%�)�ͪ��
J:���~����C�V��(�4�ɼ����BCX��TV=� ={[]w�����f�^JM
��\t�����G��M�v��N��L+6�ܲA����9�XvR�2ѷ���.���+�U�e]R q����|�~L��'E̸�-��Q��0��v�E�UT�XY�9N�3��UHDi��F��aۚ�PD�Q }���(b���'���!Q�-��}����@��Wמt$��Id�[�N~,~�3�:UwA�Fa�E>}γY"�y��|��t��
���/t��@���
��-�I����C�P]�,n�b��yY�8I���<��l��چaS�*�=�6c=��rFy����{"�Y��@{�O�8R �o�ؗ���ڴ��N0��c23��M:a�e�O�PE�;�Q��_�O��Aӓo�zd�j��?⤩v���-L��N��l]
��|O�)��,���v���2L?u2�Pm�R�bٱ_�T���O�F�K�M�	5�IaC��r׋a�Z9���6�JB�DxI:n�C�'��Q>u`��'�&STJ�)W��2�qe�غ�T�Q�g�=wi����]�.��7^�3��W�B`�&˱�F�0�C5-v�������߿�5�w3���پ�N��a���Κ�iW��F*�Í]�3��D�d{x�/y����ݾ���ܐ�!���&[kY��q]@���t��~����l��UD�P2��˂G�~�֛"y'��]� p��E�T�ygVH�V��,���j�^0�b_��Y�)�n��,�+�$M�ki��驭�	����ݿ6�k!)�,�v��E<�\��.*X�2'��5,ڱ�Ăt"2�$f�@�Z ?��o/��qd2��BB�/u��tm�/�ꓳ7�6��p5���Ί�aB�>�[
5zY��t�5�5�,��C�fȍ��t:Cv�B�o7�p(���*"YI�@����vnYď�Y��ww\
�*i'!����y�7�/�2�P�O^�R�+�����*���¡rXx����|^��n}��'DGd)D��M��M�-]|mh6آ�nvv����F�e�)��6���}��=W�˚���"�gޓ�@
�h�F6�c�F�;9[g��cʐ��
��B��٪\���=����v�B�:��Y��.����䝝��a �����̋�i�[����"NJB-Q��,ο�"���6�z9+�^��JY�D�O=���7��1ܫ��`�I�-gm[+"6�S�p<���Z ph���O�?��Q��3����g��Y`2bo0M�k�:��Ɂ^<9�!^��U������n1��N%hH��&s ��7�����((��-\:��+���~~�|%LM���^�z�'�Y�r2�V���]�f%�E�/��+�TG���8���3t�ho}r6�T`�Bi�/#g�=R�i$��;<�o8��G�N�4�iJ�R�8)�(RUS��m�v>�׹��0�$�x��(����~[
�x�Ԡ$��цC�;�$מ�b	���T�\��!S1��(\?bѻ�7�w2q_/���3��>��Iw�����H��S��g�= 2��L6���*� !y�/����bƢ,�ő0!"���0:�[����gp8L�i;���I�h��7e��u��Ϊ��)?K�۱�X�������1��j���5N<9.#��?� �����j�b�5�H��s�(dzjs0���O������u������!�w��ݝ�O��(�pC0�"�Re�h�#��蘦�<^#��u��)!k��U j:8���kы�b�huՠ��]3:�ȼ��и6��ju���*0��0�,�ī����3˄3:�w!w�&b��дC�Tė
���S�QRc'��Y	w�O�N��s9?�tZcE���?�M����P���vA3����A��g�D� �����ԏ�W=��M�#����zX���s�Ə����7��+a�跁�Lb�:���+..=9�F7S(o���w�I���ʟ�Rj�PmE��թcy[����Oc}���0%aagD�tE��J�)�hFT ��ZG���p�9�F�)+�S�^��j��(��Z�MP�)~01��6Ѿ�d5�D��0*w�XR�&Ltd)"������b�ރ��r���"]c�#h���:��� ��Qh�q�<7 ��+E��20X���ɬ�&U�N_���]$�r�M�� -��&1Ǧ�w=̴u���b(�qz6�@�{u �V3K�=�g��̕W�͎C'w ��lmո����&��E�+w��ʯ+���es��r��N��]J��p���́�C���h+�n��>媊h���E���e��������^ߙ�^��+#z�:���0|��uZQ&r�#;n������{��[�Ƙ��ia���������[.2�}��Oڒ����g��$ڮ��(�e�
����{^�]oxi�dF�T#�Y�5!P�dX�7�~�]u���_��;���w�]M�8�yފԭ{���"�Ď�Q)��7�@J�� >�Һ���uZ7k�)��3l��_X�ਗK�qP��`
����ITk 
Ob�y���&�"��C�+�n�7�p�0�l��7՘��,��� �u5�uB��y���F�5�L�im�d�+�c���rNG���L��&����m�q+�>��GX_�ؑ�K��aFȥ�ޣ�v����P��?��l�%��gԈF~ rx���V;&D�*3�<�i�dG�:+���pχ$3��Vr���>�֔���c}T05ش5�5�g���e�R��͠�jyb�oĒJ�|�TJje�Y�E��y����1��%�Jf�᠟��d�ho����X��ާQG�̲{8X$G�>�p;TtsO�C׹��9�ji�:�~���Z-���s�ujV!=�A^��S�*t�iZ��a�i��n[��ڄ> L����>��Ņ����cv��d܇�ǌ���'����IK̹v����$�C��:ECHwc������E����+P�H�p��a�9M�O�8u�N%��o÷4*�0�����0�<ZZ��glYIV��Cm���1!��1����J��YN�/繍����K�(�$���Hӗ�g_k����tM�9��f��9B"�Y��0t��Y��'�K���i���<p�R�>��j��g`�>��-m�g��O�:��(r�����U��1	����S����:���<| �/�{q;R�Ė0-��;Ϝ��P�q�m�B8ƫw����!�ި�I�bTJ<C��V�lү)�H�z<1�CQ�����H3���b�����j�
�Ҿ#e����~����]~�`M�� �ܫV#R��(�#1�F�en����ar8c�/�r)LזND����N]¼�3� ������.�$m0�����D8"���4t���(�Et��!j��!��)�����ݲ�Mb��3n���6qx���w��P�Y�.OS�����!z��Lv@\����rh�ue�y\l��F<֫�P ������vv��}�^,��[��A��7_����*B��>~��ZK�����0��y�h��� d'�X�Q7��n��w�Z'�C>)��k�H��/s���J�G��%DO`o�w��i��-��Jɕ/��v��?~/9�E��~��J*�x��95����}.���ix��i�v
Z�7"���c��#Ǭ�����:Z�X��'P�,b�2�����r)��61�#F*Gq��Y�8煞L���	�9⛓.3|���U�+.	c29�*���'	���6��ڞ�����bj��1��v�^ț�\ڞ��A ��Ld5�1����u�����oW϶Qܫ�,�ɍ��/��U�,��>��%]^g����Xۗ���-io�@�hr�_��a�:��[�]�84�v~�Z8�2-)c�ͪ���߅�TI�Hu�ţ�N](6���Gez�?���)�AԂ7$�/�z_���EVu����e����	zMp���B�1i�}|rE>HM¹���H���A0/R�&��^Y@%OV*%�#p�GB �U��	a�6�"@��D�`*&0�!���z<�{q��j�Ϣ��|A���)�����HMM�'����쳘�T�A���t��[��7Ϛ�;��Mmn@Iה�[�w�5n�N��C�%%���Y"/_u)v&�ސA[���-u����R�V��Z$�ʸ���r�j���:����f��5j�p�r ����r�����ަ�沧*eT�(uU�R0�Y�A���Ãȿ��ĩϲ�:8�?SE6�A�fq4�4��6fh�=~�F��.~�o!
u�K�d,Զ0����&D:��M�Hb=u?Y³^��J=D	L(�ޞ��UQ4���rc4�V)�-O��B���6v��l\�܀�g�,˲�/گ�Z�D:�XG{t�RI!<�Ib��K����� �����f�Ϛ��h���nD9�V��������s�q�s7�~�L���!Q�wnQ�7(�홶�}�}G�	z��n���n����8�	�@���s�"�h��-��߳c�V�#��a���B��e3��<�*���׀���)+5�f�1c���)���Z7�􊉯��h�B$0��c h[&�`��j�;�"���	 {�xI�'U���	�rߨ���5���ڤ`ŕ���$�~X薁�s[<�t��a酼�2��&�κ�[ƆZ���H���B�a�LW��̛��tԉgBI�A,tu��[�e�l'�P0��k�;qo9��:��0�P�����9s�P���䌎Y6���j�Q�>�i��)��@,��'"��tB�.�B�7J�s���d	�WV�>��¾���Dd�A|�n~)�:)���H����W1�n ��T���}�|�ԥ��v����F��?���<�|�;��ơ�jJ�ĩ''����@m�EX��8�Dz]HB�*��:ڬjWͺ��^#����=?�-:�d�U�a�d��Z��ό�p�f��3ܶ�	�!|�W�ir�o1�Mt��� ~�
 �Ҝ�������I�xGP/��E�>��&Ǯ��E�b���mieJ�<F���Sa�S��@�!R|����װ���<�U�R)��}hf TN�G��C�Xy�Phe�Z��ZB�^�S���o`JDs���Z��?��%�ăOS��I�z�@��i�>�
����^��>�.�G9N�:���.9Hu�"�k����Y� f:��`�3�e�����ѮO84�Y<��ȅ�;(4���ZR��E�!q�@/d�[q�����@R�`/K�x$,C�\�P�Hߨ�ĳ����/��r�i �W߶��LF��j�#�O_�gl&�38u�����+S9�]}/&�H=��u1�qC���$�/~-hć��!����3�o�S	�< ���,!��W��*� K=�r��@��7!��f�zZ�;+����&��"9�r7k/��}@�`ARG��(��Ig�|���/#��=	�Kn%P7d^��!�U����#���?^��|Wã+������x��d�0Sa���Q���u8G�D���s�e]Ųz��̺N��]4�F;4��RԴ�y��ޅ�b��������~��h���P��QD���F.�ທy�W���aE�?,~������8�F�JV��&is��Ї=�c�V����O�_����M�?`e:|	��>�D̃�3�ja;"�6A�9�\��	��V�����[lAtϒ�b7g��R�b^;u�κm�Z?dh��z��p}���%聄�(m�J�Pݡ3�]#2���G"m�Ti
r�W���P�d��-�vD��n���I�Czs�I�@@��.�A���
�<*c-.��h�خ�b}�e�2��H�YJF'#Z��S<n�|�yz���W��;i�����Pg�~[\��˝/��<+�[��3 ��g�?��|y���~p�8J�ԙ~jJ�;1P]a�R<,�*�k�s���DЧu �|�`�ꋽ�]na�	��uojSewK����1=�n����8�� �e�Zk�+���)q���6�s�� ۰J��ݵOP��l�U�񑐐�F-�@��1c5������%J���L(�W�޶�4s�9����O��<�]Χg����
�����^S<��i�̔�����ESX�6@�(�,L3�A�����
�ǳ�k�[+�78�~��n���r���zä=ۊ��w���a,�I���f��	���0QuH�|���m}r��������� ��x�p��'�IDbA��YO�K�\%���Us Y�)M�N� �Fg��q�,:V$F���d��[�ԟA�`�Q������%*�ܫ�eKY;4�[�')�X<.��QD6��?�q�Al�0c��c���&Y� 0�#8��/���S���
�#CR]´`�I�8�ܝ�C8`�	��d�@d�_��5YV�8�r^pZuS��?ylŝg��蔈7��Z�,�s71 ؜]��G�D���T�,�Z��$���-Ŗ�7�/���u���Z�:ȋd]Ãւ!�EUm��?���-ϐc�*W9�h�H*�'�Z P�N�&XS�S%�>}Y�VN�o�x]o*(8���3Y��|�H!�v��i߱�4Ȇx)L�f܀vxg��P��b���X��ɱ�,e����}�~�{t�tj�J�H��܇��k\l��F��[6}�^'�� _�� E�"���=!�����N�v{̑D����4?�� ��8�0,�x��R\<���J��8��ף���D@
[AX���J�`��gs�M��ϦW���m�����ٔ�U�Z������`׈؊��I���|TYM�#�Xr������p�!�o�r����?B΍P�h�w��5L�.ڟ��@���Kc ��ឺ��\��)u0���y�ݗ
�K[�?}�A=��ОP����KB����d�nu*&M�s�2qM��߭�ؗ|��R�ɸ9�~���:R�	_���1�ii��b}0�����-�N?�$4M�9�;�)fg�]%/3�2�i�m��P��LI6�g|����S]����bBB��t=�T����nuj =��-��n�3����[�F�"��k��j�M��A�|Iې�X =Vh<ء|�
�q�Ch��7�ў�R����N�^�=^?��4UCc�*m^d;��$|�H����C"��فQ��u���foJ��e��*��x���:��뿘��H�)e?����_ɭ;q�vQW�Hx*
�F����[ftI)�9|%S#1�ֽ�k:�1cͩ6��Y��ۡ�MN�����-i�u�?�qa��ح�9ng�	�XB}��n�Q�E�o+�]�M�����Ĺ8�*��M(�栢��A��\�ݽ�6�jn���(hl�� �k�d3�{�Z\�W#��4��&��B����f��}�r��+ZXz����3]H6hgM�rQ@��;�����m,�P��jr�ԗ�/W��b�b��XZ���~�	1W�"1�}�~Ż���@�#]כ��A>:�\j0��f��#$]��V!+ x�$q��ٛ\���N۵�Ap�.��l�k�2Ɲk���aL(�G�i�&gI��X�M�|���8�f���ca��Z�ѕx�r��A���/XZ��=�
eZr����t�MNb�ԥ���Ql@��S��B��"0�s~�Ƀ/�r�ݔ�r����*���=�]LKV=�(�������d�g�0C�!v<�E�9��$
�3�|ݭ~_?|\к��8|r�y�&1g��=� ҉��t�o�A��έ���I>�v��FQ��`xv� �55�"���*-ןo?�$�d�DR�m(��+NW����r�D%��W�I�'�U�$�����V��7Mo��]o{��WuJd@��{M��A������x+&�Y�꿙��t�\k��cT���RBD�LhT6��T��� ��P��is)ttے�k����0�'��1�2e��\x�t����`���{
��] �DŇ�r�"��:��I��L\�V̜Z�J���qu8Y�r�Ma���i�̐�w�6�O�i=2M��d��*�+%�Cvf �KB����7���9<�d�E�/:3}�I�m)���Wz���%@���rT9Lo|p>l��0^���3�?�����܅��>��?<W��u�N�ṣ%�j^.�,��Oo�B"���yP�ϛZc�x�Pz�뻈����C{�.��b��LT~	1Y��������"V������C���IW�g7�L��G�hnEt��b��X�-o��t"P�s_^��@�"�l��<�q��
B"WP&7ɏD.��������a��2}���w�X��:��ɳ��/^sk��@mj���Eg����HQ�I}�L�U��XÍӒU,rRGդ�o�ʟ�sN݀�e���R�c1��w�u�J������|Y���h�����=Sȓ�I�!��wh���?�ԓ��P����3�͢o�{��G[e>�$<,���U�X������0��$�Q��g��B������� �&��}�V%H6�l��gX�#���C�Sj��C�6��;�[��1���~=��l�>�� F5�����Ƚ�?�LL�P�+����1Z�'��kÞ8#r��'5�r�7^>]��'�����K��G���c郟Q0�hmlo�рp�a��ս�	(�l�qm�%���x��vZ�,��m ��'��"������������Oö�|����e�b�rD=O'CV���E���mѬ���X��?J��SE�U�� ������j+:�ny�i�������]v���cj��s!��������X#�����ņ�&`.� �����4ҏ*�̟PU��J*��:��h\���b�_k�	�K����	��� ,!v}��'��"lc:�t9����+ؚ�9��3�i:�<��Hr*R�c�O�Kݲ��,��r��Í䳳,it��XR�&��¸�2ѱ�% d�X�c� F�5\�z�1��Y��@q�#�4�@���ҿNe��A"�p:��\�'u�8��y�"}��Yp�:��:v��E�/;�TM��k`�^��T�pԬ�{0@���G�*?ŃR{���6r�|�!��E�;aY�+yl g�JϺn0�![�z���:���O�"لӪL�`5��GlQ!^����%���m�s�C�c[�TG��ҦeG�'�*I��s���1�\�)�e����bN��T]��N��y�ÉZ^gfb8Bfyk�]��$(�^��Ȫ��اJ߫��l��\3�у����Py�ܾ���Bvۧ��jIyk�訓Yə�����n�.{~��� +~�9����r��m�����n`�C��x̥�� ۉ�t�!�$�8��qN����k�nwLT�-�H��)}���k�=�aj=��;���z�ӫ���hJ���h�R����3�I2B:���P 3����Q�]��(�I~�|�6�ʅa"~�麂�F�D�$��Q�� ��{-B?f���N�AЭ�'��.9$�$��Qw�WB֟1���ǈ�
���= >A�-�v`��"p�>m���؞���jԚg8� ��3��J�AJv!	� Y)J��ȩ_�F��p�F)`�\�_�3�G��L7�t�,�^<�8.��B/]IEIQ�%v[$�5x�Į��|�{��I���u�i��2���sb�4��K����p�izcoP�/���VP>eO��ti���3E�bu!|��~;a�Sy�����01j����M��,CM�����d�����8e���oI&N �T�I�����%�>�DE��1G���f�G������������i;�������n�8D��(f���0������󨞯P�%�uy�
n�_�ݩ��'�7�۷�̔��̛3q�����,6DK5o�-.}( f�[��s�%	=���s}�A
^Lı�K�6��; ,R�J �is��m��A�����jDl���P��)AR�w�^�����g�ow�/��;��P��#�߅�:
>��_�!8��T{�d�����L���-�}��$s��]���^�c��m!0V���dw���y�L�i>��S��R�h3�Wt��hf�=����U��շ>J���W+f��,�|W���[S;��˄�Nޝ�c�;���ir��8�B��Q����nS�Y�ˌ4��ە���G^T�6Hx�3jM���&$����A�)É%|2���1��r������J8��zo�Z��!;L#(����_�R���y,� �i&���k���糥*�jj�{A�N}:yh�����	��Y��@	��G+�.�D��H�-G��X�~BNju�S]BX��y)	�*���_��੪ZD���x�a�H���GU�6U5q�O���AYB�v`��{9���|,���D�n|)���L �Ѳ���?��`�������ڐ���>��'Qcc��!���é�Ɲ�J�����rc�0����!����x�\�qƝ����q��i��|*bĥ�8�wC{�	�[B�s���g3Ͽ�	����[w;��A��x��u��EI. �r�pԃ�(�!�`�B��Rv4s[=��[Ʊ"�Ҭ�}����ݵ��y�9������٠d�Ӣ�E@��HO��p˕�o�N�˙E�g?bV�m�^Ey�����i2]W�%�R3֥SZ�П��D	�];ed\�Mմ���`���ZN&	~|�5	y���<�J�LW�)y3���/�I����Ե*��[�Y�e���Q�6Z��r8��W:+ �1��R�L N�c����R�7�]�_p�[*�gg�`��?��W��MYV��~)Ճ�Q+;@"���6�Ĳ]��y��J��)��2���Z���!��3xFFB��O_�q��z<4V�lY?��8���4"���3l��29{�6K��?���gRV��}R=�#���T��ˋ�Zѓ�X�J2:�V����K��Pk=K�(��<�d���F�M^#ڈ>���3���-��q��>�sd众�,ƚ�?@T��6ѼB��X� ���k�}Ǎ��H���&ƨV���9}ܣеbT�u��� �j+Q������VxVFn0f�E�����;������g�^є�kh�%;1��q�F�Ǟ�v?�*�E��`��!pS�#pƣ�h���`�Z-����M���6�ё���:�_�`~fr)b'I��{��0�����T�)�ںD|D�bQu������Y�쎠��U��u�l���x
l�8	�m6o�{�.��J5��8�^��Ue��:6m+�Gx��g�xA�NE�F�����ZOp�>h�:)`\Q�VƔ!���N:N0��MX���$wuJL�I���k��`��\q��mJZ�^����T�����b];��^��3G⥷P\Nj����$����GZ���&_���TD;��{V�{[�SR_�<Q�7`�--��E�a7V'�&Z���9e�����pq�i��؍��'�X�e���0�i����^�wnJz�@��"�>("�*L����n����������rU��0u������0��R8qX����@�
�5��m+��7*������Ǣ�}�͗>X|�]��_�|&�LKp��/��`�1��r%g^A�ɣK�����Y��嚐���}�]�?��B�-�	Y���ڣ/�xL���6abB��w�E���W_m	y�=���-f��蠂{Ȋ�h#�Lj���I���>�"�CA��3e��oQ�)j�\����d��5�}�&��-�G�2��ӌHv�ZU����؆6�����XXǍ��fD^1�a�����X<v��1�+�NK}�Z�8��Kk�Y�Zϙ7�{��Rg�l(l�Ҡg���~���>R�A����%7����h�"���5��Z�}���;�O�A-St���C�ܭ{����m�0���ڛ�hyL%K�$�	�C����B��);�o�������f�\x8�G"��oqO��g�* S����V=4HZ^O�XU��	G(>�<o���.�^˾w�8pw�,��sD{q�a�5������-�����3h�k`�=;IKm]�����ς�[aiJ�.#w��~��SNxb,!����g������-TvlI����j�J1`��4.�$�)uS� @�|�=R
|��.���xZ�$*0��
�	tH���F>��(ݛuj���Ͽ�ݸ�8+�Z�׼�t�@8b�!̯�,,�`�
d�i��x����P|&?z:8�[��f��~�_$��M64c۔�;G�odq	a��^#�g!������w
*�T^L�'_ɍct-�%@�~W{��
�R.�gΓ�)�M:_��EC*������Cϼ�2"d������C��ߐ�]�xu�ȌB��Gaxr��	hS�ĸ�����6�BF���c�7��?CY���#Y�s�}b�l<��L��ඣgmF>��ԾՎ�\��*益���r��ը����VF��~9��ѭwnZ/��[��ma/ת�C���;1�D��Ӂݦ��3<����aQi�+�uJ[l��ag�����q�錐<'�=�e��F��Ԛ�7����:�ڑ�� ��������D���k��]:�ؾ=z��_]���n�x㍅oGQ{�	��K؋�ˡ���i�.#�Z�����-	�1TIf �+�F<�)1�V|:�Y]��a6뚑��払.��Օ�� M`�s��\�%�v�[@8��9���Ϻʁ/-6s�S�R��8��3ps,� ��vV�.EM��HTȾ��l�s��;��D�d/,$v{�!�̧5��qL�$�U*!*.�4g��H\W���s׽m
bZrf�{RhA�Ϡ�fx�)6�b��j�l�VNg��u+��Z��H�-���O�ܘi�2r��'^�W����P֙����j�C��r5���&�a�|���k!�@Q���Ҭ�!�0��I���^��w����^�*O65b`���r��'4d���JLG����+�@�P�	�G��0�߀���f�|ӈ��HeUv=ݷg���G=�����G,�
F�G���et�u�ҽ&*�S��h�k��N*O�
Y�7QO���x(zHz�d� ����w(r�s�u֞9o�?S��4E���!�	ȋ���[��+om;;m��h	/;c���1��)�����(���s��dS��klL>��b2)�q@@>�v��f�o���_�E�䃮���ZQgdo�Z�kF"�� (�l/��l�*ΒfM|�P�tYdtHO{*0cGOKx�.�1�W~	XƼ����q�΄��N}�?�4��6��q����{C��b>ǧ��>�t'L�3Gs���\�#Ȁ�d��w\��)�*��%s7����N����,�,Py(�H�p9�O����%J�=�\$
M�p]�U֢�dQYM��{��CAӦS����r&W����!���z\ΐ5H'���l�w�ѐ���n}��N�Wk5Ԭۑ�������Tˠ?�����������*v��=x�G3��
F��!m���ͷb�b"*�;X<F �d��;���׬T#��K<�ز��S ��q�e�����N2�x[�CV��q�"�� �(�ޟ�����x�A���gF��i*��Q�
��ﾮi;fT��7�n���UϺ_騨�?��-�(V�7��w'�|�
Ȼ,�T�}����2l�zS����vW&��=��_��>݀�!�;��.���CS]�_;z��r�:Y5ػpn-����Ϧ���Q.C�>��� �Όݗ#�#�>\�2�	i�~d��3�0�fp�7:٧�/ۚ��3�V�bo\9���$��(H�����.Zd�-ۙ�z��A��J�Y�s"��V�D�^I��xV��M~@NN�jل�q��,��d��H�
�w�6��d\�
Y�zkqa�GN�*��-gh&�쑣��k�:�9�)P�'ă1�@��܂yOl�*Hs�����	�����*��p�˃P��f��0j5!�h36��?�,b�=�����c���+��w�0hH�����G������g+;��)*��è�&�Ȉ�0��'�R�f.�f���i�����{�eX_�ru�5�j�]�H��AxS�`c�Rb�?St�!�	���S�@�n��������p3h�+�v����Ԏ��;q�؆&dش����!5���E�l"_)k�k�.���Q��ǎp�uz��H�ƒ��d +�I`��9��l�K��
�JwY��z�{iF�]�ϯɺ��:!O_����Tw`s�VL#)�_�T@�n�ij�U�Ľfl-�΃ǳ�����Ϥ�7q��]�DX���5>Q�m4�Ho���`2ȅ������"\�S�+�0�)3k��D����n�XcX������*�㐛,s��j���ރ�����n�˼Q�C1X˕Є@M��Aȡ|Ç$˅�B��ci�@�wב�]�L��(��]�Ȫ�q�����oA1f����m�!�'�����[d�i���tS!���~B�_�u��Di_��LǏ^+$������JH�h�j�5�0��U���r�PՌ.n��J�
V^�q4�ۯ�Y�]�ͨ��&f�m!" �c������ޔW	$�Ӫ|�=N��m1��XF"�f�z��_��p�q��q_Y�,���)S��]eA�2L��F�j�B�.�A�E��wNw,�E���aG��X�HD�����|?�� �&�J|F�xK�oea>��j<Ú-�����O��Go}r�JM'y*�DX_�A��Oy�j�P7bB�WƵ��Ѣ3�1gL��ր8Y�����:�IT�P�a��ѩ=<s��3I�!v�=�=YQ��,.���*�d�Ŏ���&�Z�j�NA
!�.��O��٢�M�9Uc�q���y�;��g�xZ��'�!Y�ij=��47�F�tlM�=<����9���j��x@�� ͂ԥ�(x1+'�N~��X�1�Iu���0�j��>9�(c�fH�[_-�ӷ�p�Y�\��kp�b3� 9�ǃ�:�O���~-�\� �����-�=#+�M/ˬf�G�d���?+�n�}��M�:�(��h5�iI���ӵ&O�y������H�����5������	��D���H��W��Q�o�ʰ:���7����8���"I��
�:��<<��<i1�����yà���߉��w� }�N{��u$	Z��;>�*c�\N`GM�Ϻ ��>W�O��,��E��ړ٘Z�ɸ����f=c0-o)v��~�U�n�l����^��� �`�T,=�K�X�?�N%!�[-�>,ڀ/:W�ۛ���
�өs���Q(h�-�?�	t%��;���aV��%�x��󯕱Q �Y�~�
zL�2�9���ۄ�
/��*B����P�|���;}��.˙�-�����oe r�*��<,Tu�������z������:��)���r��zY)d��kw��ܜ��d'�A&3$mG�^E��u4��A�<@U	Uӓ�cqH_�Iw^>��rL}Q|�#�m�	mZ���{qYD"�@�'X�������6^b�rb�ݏ�����b�#��<:�&́}����݁NP�=�(6��y�0���XiL��T���
�"��x`6@NU�\C;.A�6ٱs�>n��������
2���e�0�ǅ/���)B�_�Ҩ�c�w���8⟿�6Ø�(�f[x	�[q��k1�t��� �b����c �oB�I���Pe�%G�$|^��`H�bh�v�E#7Dn�]�,授W����S�]A���?�m�#@-+" ��$�&��Kw���������ᢉU�D��RD�K�4W6#�4O�0����6���>1EҪ��3�*u���Ā�3�=��.��P����oL��e��̕����F��i����B<�
T�qGF>�fP^<�}0{~���ẔW~J�S<�>	��'F��d�>�Vt�+���)K�rD�b{>fe��M=JM�Ў���i3jF��8%�R�3��0l�_%��������a��s�	4��s��V�8s���Hܤj�ZOV;�B�Liyx:��$Aߝ�^�bW�V��א�>T�S�s�C��xÜ`>��l�*(`���}��5����
���^�ښYb>��iN?<I�����*���d$��^���c.��dndX4;�ǜI�jwo��=����6��2���0I5�$�Y�q,�h�|4w;�wϹ��O����j���h|c܍�Q�&�T&EU|���iF
�Z���!�F�#��ْFE��U�/��U3k:�#�n	����C2PJп��f���"��gqG#���[M�&�>U.��h��i�z�Ng�F;�Oc�ȫ��_��}�����p���]��+O��$��s�c��p��M�$^�2�R�x�p������I��>�`�98��8K�,A�@��z�f�R���Ԏ A�o!�^�*͂TV5鷠��:�=��z~XU��~ϥ������&�嚂\�{�Q3����	_�e�"#EC��Zv�S�� �C%;��L��Ԍx��j�Qzd��:���Y
��
�����/K!�%��)�%�({̈́��>߿I���gk�~�.8�;���EcfI!�-��a9�a�dQ�b�b�lh6���x�(i'���:	 �!WQ��<;�ZY���o�%D^���HƘ�G�~L�) �]L��Eb�6ql��e�ti�/2%�FX������K���@ud��F� 4�����co��jm��}7�M ����ZṲ�C?[N�,C���\Xo{�
��H�Ý'���n#�qH|(zl���muQ9�] �Ժ�К<;�.���f��o��Ἰ�>�J���؟����v�26%L,�W��</^�3��?����
|��Ω�vx����������o#Z�b�����$�ҩ_��|F���f{1�;-����������D�ŗ�5]��vf:w�,ہV�p����+k��s]�#4Sϋ�������ӎ��ܹoB�s�J�?R����~\�5�ć��ѫ�<�"�f=)h���8�?��!������=@� ���f3_����1���;�W�{a�̶���w=��#���T2f�j��6�����wE0���U�`�T�G�f���CO�����y�q�V�E�F��:�^��/& NO:��]�k��h�tl� q`�oe��ckj��?q�"�X�o��8
 ۝8O<�����	�\�i�`~e�f��Egb�~1��?�{���=YȅϚ:]����9�L��l��`�/Z�t�b�Y���U�\�M}r$�̖{c�dܟ�+�����o�7$w�����9{���-+����f���@7����Z�7�k��H��؊�t�,���Η/�>���a:�@��{��|
9��|
��ܑ���8t�3��:�P�".��>�5��� ��n+U������Tw���&s,��`M�`�Wi}�A.�@�4;B��H܂ؼ)y;Mi?}�P<���0�k�����2���8p��c v󺖾+����H�]tj���!ԗ=�AW��F4����f˭L�zC:Q��_��ݑʨ��B����4l��o�@��F��٦���bp�m���O�O܁$��,ϴ1��7��utw/�?^�N�R8k�7�m�Ư�+�7�6�ڱ�,�i�__@�����=�#�fS���P�Q�����&�F��'/�gP��o��<+�7n(3]~\4]�u���:�ԝV��,K�;l���F�K��,���S�[p����!�$�0V^�
�G���=�L�N�v���9T��PJTE���Z,���_�m�⫀;}K���S���]��2*c���xە�qy�ԅt�A4���e	$��F_#`.������2���������(;�^T#��IZ]LԍޭoL�|�e����n�,0��a@�^0VA|��DWj]��X؅��<_���mds�[E��/���hZ9��w�;�K6��fv�iR�6�Im?��5T�]���� �i��HV��8�s=��ڂ3v�j��M