-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
MTTfIAGS8bFgoR4CGwUlrGPvKgDY0TJ9/vuoLTEar2nuM7gBvMsNqiHTFO6oRbxGt1wEMGGqQ0mw
B8u07sF3RA/TFqpFQxhkOl3/CZdoMQywHCwWeZqfBokRh/o1OxmJlq9ntxoboR/rXenjb0EZuYHn
x7eyDZDC5FGGir2zmKnhM6mfjE4bMP0cOYSAu5/iW/l5ZC0gS/p4I00mgkBYTcHgARqY93yyAAlA
yyH8F+NXZTQe6Xfk9yelpdddz3jZxm2rPkHwDoGjNIXT5UNjgz1JRfiBXIn+8QOsRS484L2mzy+W
qTpWLCe87lPZMc0Ofu6UXLqAdfyLERd8bhhiIg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 50592)
`protect data_block
h++ruC3uf02zb+5TRlcBRaIp/RmbxWOWMMg5bD5TH/g9AVJKzjugoH8eLPoqJNOmvnIQvKema3Af
uy1RqHwV8EZEllGbPEOmbwlVw7fdaz3sf2mayyLE7UD2BDjgCgWKpG/6LOt3qUlnCMsci1YQoIHe
ofM0mHXGRS8Hvr1pz7xQkpdYAfVswVwRrNoIvw5zZri5wQzZbf2tuWJSCRmAtVthn8DHZ096YKzV
lf6TDBFG8RGQcq89h54beTESLWc3AeXZ/TM9qUQbygY/FHWdv2LzNQfiOlZGo6B0/I9eJ2C4AVjE
0I23pDDczHS2fw3hEQglQiWwmdwF4w1g7aMQYZViSrNwckvIHP1r0x07LsZpVtgXY4yFHV/1ywyO
o0bKmJCPWWmxeOXrBR3x/OOFDsGi1GErGTFUTJysYN8dkD4mE1EXwavg+riEnsLy8JWc6zxe8b+3
Mtw7jbH3INW2nsJEMPL0lbEV77oxwmP2iL73Ag+dGtFoQi1lNKcGNsNFBjbem50BI1bQz1iaddGO
hpqjr+kgWYLe5cEVwvTNveUUbIfgOjEuowcHwVj4Z96zPBMEbhqXC9O9fHe8Q+bwQVaswXoV2uqr
YQnLPcU4Tpe1bqE5vxGNj2pZ9uFTH+Zk2SFFvYcldaF8Y3TnGLvplpZfQAySmhR0SFHyxbbXEk8k
9eXP6Bwwlgw1padaJT5huUn5ru1hMr0sssr+u8m7e+ehVS+AbpFHD6+K4WDPsodT5NA4u0crVj7s
ahS2V/Eulhz9zHTOw75/kObDkqbs3SDlpdVMKzoUSY1ItWEHF1KWaGVPSG3FPbKyEOXIy9vHchRh
34QKetH1Me86c4et7xTTQBXTCDsA97HfZcorrQn9veZ0ZbgAXS0espMg7uouyTOhbmjTlTqS4aL4
sV5nTg/mO/OmsJ5dcgMZAsK7d5bnbjpI12TgeZip5IButYMB6qLQR2Uom7fpIjii5F0I+Kk0rW/6
/yoTaB5xD6c6WfI1Hb5KzpgiV4BzbCCJjFFt/AYzs4Lnba63/4XXhjCAOXssHMYnzedOHAbuLGmY
bzXp8bpFjJ14Xa68XOdvkJ1UlaqS7GmOiJ3RljZ5G04kBkQvwXBvA7RD3QBEJMk+KUNScmcvjz7v
qGfzRbr6/hZkwqAPi5wPtXGkbODqaPYo1gOPKfuJ9stppoI1UlhTlnu6QMSZaHooT7sANT3N+Ijc
dqODWpoOb2d/NXe36gsd0Y3JQHW1KaPiJHjNW71pi6/yfZ81JHj5kbnzort6th3QbIPzvm/u6Iws
gUaUuzCjxfGDiYLN3wlInUjIq2EmjtHFKduQQVlHDha2EtsyjZangL+qguIlw4+zUd/zKI+vHfTC
We/KZu4BgvJKDbWScUtOXTpXUx0EKcucZEuPmvcivUyPmSbY6Q9vb1+XfKg+utszRsnMb8MetsDO
zUT3CAx51F1pSEVRrQEnCUz500mnlt/MYIwlYr/a2qzP4qfpYBR5pTfoN5jAHbvh5F8pyH3ma3VO
OReOHJ8olcz3/UXovDyI4zi5wZ8AG+I7y+AeqIHEF06R0CejqBhYGEi/Sk5An/2KAM43oZtplKCf
FVJAarAVk9jQBvaEu2k1yM2gq7kuNhqU9dfolkavwwHXUHgbo6K6R9xBJuBarhbdnmkm2F3gLWes
gjGQ09ZilVoOa3G7swbqJCqADZLZgI6CNtjVTPiuVtmR8Qf2FZnv5wQ2J67HTkR9v2FlfLKQiJFp
8QaBhPqwOTQp0Lnit4QcMuAPma9/zU5D0l4PVao9GeP/2km50g8vs/iAWelfhY0JdfvVx87WIeZL
r98+dbM9dEhCRsc1BYc5uA4M5BtopuKZhvrklgahLu/Y4MTVtHdxrZI5S2/rYwcWSElw6m5Jng0Z
sbgsrtgF0oyPX+JFGgPKx4YNGxZfGzFGpWQfbuD61yFLBGmImP2dpeqZ/q+VGAzAOUNtMhw6D3+/
0OT5St2e3MBO4RkEqBPgEL40SzzBuTozk0Z36rvEgWt0hIMbytexLWbBOwI9XFRC+4/MsAKULrlW
mEuzigkbhQIK8Oq0HQuz5cGCWLSaFJd+bdEcnZky0Q0kErSu+VM63cYCV3Fbjgz5rhxqDgt5F4yE
voRJjTzXzyhciFKCJdWA2O1pWdlKckcJF3rOkwtg6A7MQo5sRTdfCKYmGbcpKjSUplWtsSW2aJkz
0p2SCWl+BUe2tfAC27TuDbvBNNBm/65H8/6rLFYgdMM1SZWjdpBVtDHrlw0asgoOnW3hKY8k+KlY
WQdaUAJRasssXIMY+QbsXsSzybEIJCPjQDHMxl3jGkK4aCFJugeOc0sy6M2/X0irZVPOFh5OddBj
L8X0Dz6Tiwb+b4wKPe9WDM1ywV93XP4KlnzcLfh4FKK4Q8/kbqLLMXZkofsO5D0nX70th7hHjGbe
zqAPfKE34badEMJUpCb/OFAl0HJe0gsc5tSrPAYPY2nXr4oZl/K4cKe4eDOx7OGefff1V4J9kjo6
gF4BUYVXH6l3ndeCus57eWtl0K1SIbrimTjwf3F5ifoOsY37rPJ9K3hiSBa0IkdiqxVagLg1hvo+
8i63KyvnUuek1Bzp9KHBKL5dR/yKNttpJRLUieNf6aK9Ua+hPgOvTeL0REmcug9Cvvf17MfvkZj/
up5qji98USPvdqKvbcQkZgEpCHoIUO3ALSXz4RMi/ZM4CPMbfCbRLspYzl2/55uPycjc0pB9zNK5
vpDzztJZ3igV8+wl/bfI5TEUjLXjJWUibUPq8iZ1ATAPQ8yiwCjaEFJXHTaUG9EBG7+qAMX2wJEz
nyrnLuG9Q4oxfcWhgvw23QiJ7rMfMMO7tJALrdpM4rWXuPe7seUZmfaY7yPeydUqDsjIJM/9Ehyh
liNxtJRJXN9U5pMas1payL196WjnSfI02MBR7bBoeJ40ynYArgl4u5x0PzBsBnMmtVHbiFsY32h7
yINw+rLYYmbQDbw0ro7Mkk90i47nhdy8DVWW4HdHqDpsjAAbZ/DuK2+YlOrq/HsCWgpA/08cRzlQ
Y4kB88kgQhpFzrl0jhtj3u56SAwBIc/p2i11xHXp8l6PcsqJa/R9/K5Z0EhQF1hqthnoPA/5lbV5
86OsL+eaZ69liSBKEzv39yDPmFFimYA/fT4jArvGPYn901IS/IPpU9xIv8vgon0Y7UdFPq1j99h9
wtCLkIpWEjtFErxYxS1OpStEPs7eOj2agehrfAqAh2xPA/ikFe7WLfpg2F+fiNJuCQ5LJMp9Lahc
I4vXk1u67TaIPiMfvj4UZaGQDknnl2Ojnjk89oIx+kGxYR42j5Gj8rOo6cFmtnJ+M/ukhqWBzmgN
UCxiuvRFAEa/tVMCcduxsrBpZ1GcOLlcfRczpDPf8F9znQyRfahu0zfWGYbv11fNsm5oCGHFA8on
Ttjesfk7EgWo+3yzrPzQJj9ytu7BwGlEkqKt9tFofI29rUloMTKYABtUsnuvx3Um1pM3TZP5o1oQ
iOYsxTtJXXqdTg70CqgQhZgM+sf8CYoiTyzbyxLQlSidZW6Z7ync3dFOzgLw1prpdINRO7mATU0f
AsrAxpk+tAocuJOs1EzzMWaGXeFOwwpnMw00t8EJQlHGX+sLJb+kpUpo78iamKaSkuzAwJLfqnEo
DPm/9gLrWE2G+yi0dF5HtXg62bXN/Id7dGxU3ly+Undlw+zYegsinieoybyJ+ABKWYuSTSAF9CFD
1MrMpuDb7unp+PSB28Vgam/f4knud9c9Foq258zQKQp2fWQiudfMMDSULRpkP+R0dnF+a1uACC0+
rCvFTz1M5EscQ/3WhNAQToWJJDw9JeNrSWL/9MnDpf+YQO3QpjGnlZGxWqt2Cxf+ZE7KBUIe0krr
4DfLrn1rLKiP2I8ksjphB8abDQnqdxGoAa1/FGYTB5roFd8Lmu6BfE/4MsYe6ncQ9MzRbFh6A/BE
r6L1+Vk1QMHCg5waskyRbXA6saDpvNXHuA/aJdhdynxuISpf1UChHH7IEPIoXGmStQewWhFTjk4s
kxxdM5l8NlLtFvzpcSJ420CEKFygLsxjpBkDB+MWR+YE8EgGEnxBIWMFJQIRMUaXeZpNi5hwHtmh
SasAe386YSf0kl7IN+P1bxpfyx0cHI6Za5dKVNfvKXQOqWrhLj74KgiobGgRJg/nmii1kneXoOVv
UMgSljQC8cWiLYg8oDjvRalAGTP/jmsHmZp9NvIFi8DosLwYKwBZrTGdUUtC1YIlTMdDjY9CSujH
zJ1dCffGn7ozA6fMVURJAjD+mkBnIi91GmMtTgMuZGbrOxy7Tb5kfknHK+5ihKbTgJSehAlsyp2f
xq8u5krCGPt6/JrbTYoc2KRn2XpZDYtlWefrkuYS+LMnRWMslupjlqlKTTCWjveQBIug4/DQkNdi
aT/MRwrwzqzrTtBgzHiTIoDWcPw+4ZZd1RIFK3oDd3HzbiqQUoozoXwb1rDl0XG33MPdv3ypEjhJ
5aWR5vCh63psJhP/FVFnNPRCYnk0EFVhDVDSFmC5zkv946+KgZiTH05IfoOFNMSH5xhw2u23oFHl
wtnwMPn/EujgJCINWgYaXkD/Z4d0OHnRgJf/5XFfpes8O2V7qQlR/aeGo86PFJ8Ef+HSmnOPHWov
d8Vo06Bq9v+BVvfSpCHwBsuOND9+SXpEH1IxdJFxFdFOght0wO53ZFR2ejMC2sKYsbsnYNkA4WSO
1MLd05v3V+Kg/C/WVupObQRZ+hiWl2h4jj/WAR1y3lXHaZv7irBSR8eqE49Liui7Mh6VqED437Fy
AQ3Xoiok/aJYuj4KZW0GmP6flrCV+jM3PDVHHZP/9eirrjQS0tgvcxpp/Eqd+u1H1Vyrk3hfhAiL
uAWRd31kVkXMRdyUhH6QyxNLAHkXgqfANNRbdYq+k4I6fdsqCGeyblFfTg8+ihtkGt08bXXIh7bI
jMoTeEMGhdFuyuB/WWae6sLvCicRAC0MWNm2u0KREbupvOq9TLdmnyNmEUI3CJ9JVKIO4DkdkO6/
yGRnsxCT+bL8RfYhuKND2SH3zrhCKtRtZNwn1O78DdaAwR8BwRAZGtI7iadd6fAHupCEKiwZ/TgS
pw1tqy203aHclBGOVonyKmt8N9jMaPUIk4sAtuLeAV5cglwXsJ/y07v8RrbPHeLjL8qJW8TqA5xP
AU5IfRq+knRQmkaw+u+iqvb/8yFuUIrF4HEiSz+/1MPC5kAtPJwBsJb4kSS6sB2yS6ZA2+BLtI9A
KpwC89UOKBxL97JP3z0SpKqWYnMainTNhrJMjTBzR3azs0Xd/7xmQ2EqqAydUZEa7UgH2KpZquRt
JPBNx0TKVdZdi6bC0PAqnYQFpvFD8xz5QtG0O7AQwUskQN137tb+f5ibCprXP/+pas7Smh0vzX9R
4jQwxM4qhPbzb1ES6fWI3nTbPmZ+P15Nh6GB6WN3KLsaTo2rQ6JdL1RVf+8kO4umrWmtrkNWc8O+
kxgoV8TWh4C7ONPRlTo8tSkU1Hcy6bM5e9AMTGsLTg6NN7q4+ItUgrMgeRXmfBFMuFj6AmRcIBa3
3EQ4aoJ7rRYohFl4qe4GFOx3o3A2Q7BGDuRoTPT+nIcrcNRnOJqiByLvFNXGbwULFRQh311hzgxb
esBX0Zc5p7EMCVPeFCnI0ELAImepBmTH5uopIvJIGrqE+E3nfgXRoULisk5O/xRrUbCB6Ul3QiRW
wmnEydVvUZIb6hcbSxsm6tGqW14RU0RDYkRvh2dZT9TayWAQwl9ecr3qFQ4ETQcEu2Kmqees/FGV
je0Y2EBbwRwXndB863LCBEL41TI2g4WVvazm01IgKYfX0+3ef2+xcLKnQu8Z6Y1GwRndMD1PDXl3
ket/K+0KeGT0MvroLGaW40+nmABhBdnrtrEiBQSQw9iNUh/gxMPPHy5NqZtBwGnuUSMURl2FwHhk
f+dd52P3NPq8Ka/x9lxUQJHM3ppzzONrN3AolAyO+oymsZHn66p42qmpXVKMxk3Pff3sJsqPH0p1
yHfU4ZCOD62jvfb40GtVWQK5pAcRlAK+ccjvTDZPsNIfYr5k7q9o9bAMFPwyMJqVT82EJqmgEebp
ZeMl8MGu3uVtqTuLQ8bfAvoUf3fTeE5/wJJQS7I1D38k/cyu44KA8Z0aijGZe934reH84/RhWV4o
DbHJV9QUpAvypsyCZ1RxVYfNSG6rW9BXgb4Yh5VFthca3Nr7NYKVEYsuNHCjLm0Zu9SbwvZF8hYe
wYcAbHCLNwIN+I0WDTmaMUvCzn2iMebiCa6njKwPMC30x6tOB0AWbPX3M493gIQV/CzbDhdO1sl2
vuFHy/BUBpegaPRI/THGx+qX9vpwkoDKa17Pb5Yd6MK2NtmJrsR7oVzk11ytsKxaaVJt9uVWHTjL
s2WvUal+ecQ0vQGaKG4b4dKd8ZOmxGK3IhmVKIS7mdCP0NFcwJGbmM9DHmpdWT3zBjLZLJTduAZK
c0wpT9N83C6VMdZrNyvJiR7zTbIIx43syZKNXOvKxMT3hEZANNOyIVnvV03Q9gsxIjwYi0Ne5BJH
So4Pt5xFW9QsWJpRoZV9pdpUp5vY37PgTIc2mWxWIanBEdViIoUCxDbocNFV31cESJV523J6TKCD
XPgdnuy6vcDcpwrsb+H75x/z1N5UtXvKiGMCUAJ2QQDG0mFcrwicRDh3w4HkSt3jH8wDUY/ZhM/l
9k+UNpZrDF6a71ObfbzItpr4OT8gapakJQEo0kdrQO1ZUCZAs+gD4+adu1hCiqYpXrMrr5KtRcGv
jBcDlPEMabMzZ2AGoloeWin4f/peu8XzYJRdioJROXaIXa6WceqT6Y66p2ye1LxlIsTVvpeh+3GC
Qdj5QX9RULzAE2ZJ+7owM8aXau2kA2uJd+EGUYEVI3q28X+FlesAVu1O+tv3V0WbJwnCFGgl0TF1
OLw1MSUlbV0ukEB03sdra1LrxHsmPOs1/fyi1WTpqwKqLI2jBQqhykAjWJni7dx87/MWpMLFoMQ3
KYz2HacOp9+iL7FICrezRwem+oiPzZ7fRnnOOvJPQ5l9IMpr4+rdloUFYfTP4QVaD2G0i3tLdtwg
SRmB9WCfMPeyhD6MdP2g62cTgwfuJk48BHFl5cF+xL/+AWFS78vAHA4XVqwszBlUbS5w1hSTRxub
iSA2EamQrzti+G37QUJbIu1NM6Adf+kNlMM6b6ayDh+jnCoA7VP2n1Y+6DTCLVWhi2y2Fh2Gh/kw
CDfPmVTj16O4cfSwajhyjEG4b54peBiN6VXV3SwO8BWW1fL05anBtqUFIueQCZ2QMLNONztf8mAw
qJ+6MJxcX5dvNSWRLeDdCCgfkqprMA0bpVfAyZWsGLW5LugOpnioJ91p73Uq4vYZVX7/9N/U57qI
PiaZJUBfQwTkOJxroLXtXh33TNDq/5qdSOXdXat/lMCDBVTVLOHZ4RE8TkmwmvPOZA3yVY/zwU8Y
REemjv/yrNffc/M5u4hv6i/V4S0Mn47B/bBg3rsWX3yYgM2tmjNnZ/qAppuRUJthDW52WeUGPvwS
PMZq0z827n1k585SqZJE/l2mf/m4zhPxe0rmcBr8lNyP6QJpxhCmtbtASKrSZP9m9VBNQdq0dmZA
KphyidiyW0VVPWp4zBOZiVNu+jXAA/kmChNh9retX/6W+587h8bZCh3mVjmY83PJpcBrOkxg4+bL
h0YzK+lUU4ArK/LoU5IsE6RJqFt6m7X7/n+myLN1d13KnP3GQQjqZCS10h93LOA4vaFuGpMxJzRI
BmPVeb88QxRpAjrWywGPOBZl2YIahEV9leJykXP6m7KDDjwuyENf1tXBWkdEztCg8zOojDVJf3wq
CI4H4CRK/qiatG96S/nITrKfI/iyIwKN4+SFPjdQC3b3avk/VCMqZIOCnhHqp8on9hfkbI8JuUFF
JwOpfzwQYpI/duvbO4DYtfr2XxnHJxQOXmEO4ZVqbu6H2sSZMvYbiVVOh4jWHxas8wFJXvlIAemW
rNcEg3S28SEWM4++W2AcLolrCEqkDBWbCChuO4xcrVZHNya6k5CW+kC9QSc0WdjJNf1LWct5cZ6W
snM4Lj5vY7SDMJ0rNRK0tgvMadH2KSIVi/WXnseMKWUaVZQ0ux5WF4sFVi3zOK2yVAMdwGfaqAAv
O8aLu9K0PopaMOouwcn9S+WrPY7b9D0foVwcH9QGLlHII6cTpvJBhKhXvERf/l2XFYppIY60XT4S
jdNedNHqAoeGYDWLLmpR2tS25eZD/d76b5ejhlxF7L2BahJgJujVFVXPbR5DHKsp+q/tk169np6H
aqrB3/hyLOC+7FJn9qX1H5hQvgzrwGtpBi9XbiKEMnbGONcuJUNkzasD6cgYOwdSCXXKeuJ7mijz
BuAJoMxBgDxF7ktsaCmFv5k/hdxHPCKkw/8bI3w44lG30yzxJu0qWz5BMG4aADNKhhrpOd4enzvK
NSAOM9vs8DKHulAJ2KwN9EWuttUGrGILYbFv5H6jolL1LrWo/J3m3AycpwmMNHdacFLHyBlywRc3
3lA1JaYV+do+QnKrGnGCWty4yNl71niRxQK6wyziPP2E68e02DmjfngLuYSfgiPpEPOQiQIgkSb4
y0Q3aMbBhnnqWpGm0DsgCLQlqjScyd6PRfzQ87/I141+K+hVMIDjBIfDB2d6FR651rTX/Ydpvnfn
yQmuJNAtGzEc/zte5DhxO576xOtw8tCRZF+NKHpsIASfUvHdrR5C5bqTH7S+FLnzqYFrvbEQm7OY
8sh5hOW0gDCMsxFenN7L/pAxsokIVvSYH6XF9Lh9RDyJ5p39P5yUz8af7wXAhZjT4+eS07oXDqdw
+JFNJls6Rktowgf5YKl9mT+DSACTKPYkduYxNunLd4pVBufRlesgpnJV9QipriSMBQu3QBi0MmaI
u70sI5xekFdnExoPVJj1zcO8xx+drhn7hbWtZ+eop4oNlwL5A1BJc2FCXlmH+zPjZvaUsNFAu+La
pO++h0HCIQXbZ/z3v1/THZOxKfKyuI7ERGR0MjRzsFywXvDMZA4BXBSSjeoSo5AYRx/mV46GsrRm
dENnYsQDX/LOjUEGxfPFV5vbA01umpIcpRXf4dxFdTRepeqsmEaTkURT/jYYb2gJbxA+nbZ/m7nZ
aVZBOjNPYpVwQ9BvFNX4fN3aUlra21pmnos2fJLhHCRfyX1GFQrAsKp8yZgvQlr7f9lPxUGZaRdn
m0Z9ziBU4OwbwoMDvZMIT8DmUh99pbAy3fEIKZnXSVywRY/LIJKD7PzdUVYgNr+GPmFQb5Mzqauu
afD0a70TZ0QAaQxzzRqsZF0H0u9Wa2FSYGAphnbfuH6uQ54MKM01fvPDvoHIZ7iRpq1KR8TLvWHM
BlXgP+S7v0oCq7X9wGNuZiL8O8is7q20XkA2sbww6yXbkxVybOvbAxTwKC6oi/JE+qdvwjoTiU3s
+/yEHiePZSBdLeIXEXfKFHns8qBNHEeco/1TeIQZr+R8p9sPrpLezYilB1ofVSEuLus2c8tf2PZR
B9c5na415Qz+iyud4KnIhzpWnFuCHgl5iztDUCb12VMEuxzSc4pOqQhIGTG+wh4JqlIRiqDvmI35
71FyNZedRk02kuh5Vmx++HsaCzoD97dsb2hGfuypUFedKNUxGzjB5oWQvLuQJoBB7duxl3PScMtR
bOlaBaNePmZX0pZADWfjakCfFTDdnErdGj8gDW+h98Re35yUhzYiLNNfhToR6igl7smq+hCzhdP2
c0XR8Ns3oC53dMDjritk9rr+Cnb0RFAJ0plpmwqJokoWvsRRtXOkJwHbPiHns/2Gzy2UB0h4I0fB
Oqv0QE4IEdKIlrFXrcmbdYEAa5kS4rIMsZkhP8QhVnh958AA5f6goqDGZSTZZBpCOECmd1Oo0lK0
35iKfvpNSjEPQUK9kbs6cVxpeTZb6QwnmE7IBL4pGtRwkUfXFxWF/JlN8YyA/9upENlPtD303Z+L
4MD38gmpvx8ZHksq2dvWLETD3HAvGmqLdTBTM2dGJUf/QO93dwwo+rDtQ0Gnb/O3uqVNpl9/m1pu
kMh7aKzGKhMW4KgD90Ji0STPMl3fsF8Vm8XfY+TWMWC4Lf1KWDIbdnj4AUhcQIZKG6iHPmzbRs43
JIar90XSMQVzlOF6szBeVg2gEXiTuq9058Lp1kg72Xp82U978/GBBmajJJDVjAdBHnptwg/7bQWi
sW80AiTR82f0Mm14nZRPWUG/sorjtAFga7s2lUfwkI4mQj2cnDGcRvP8PxqT0wxu2bAYkVl9J3x8
k/JKe2wRGm/Kr9WWK+B/Zz1N7EyF++oF9FsdhpswOHGoQGiSgiWPYojXCSwVjB3fF2F6ke+hN336
WRVfG2FfsIywNEvYqVTTO+zn4wozvhrVYBx5ldddkTJ1nqWX2NUYynL/x345z/dlDs+aCucikxoq
Ww4oqYUne1kk2V38ErbWZ+JU9u8SlWSvcLNqGzhtGxeVqkuHkmaffly8CaK052keuL7KjU/9tXJ5
mWhRseTlsLWsf7UZCHDmcJAZLICKxCmiI0qjD6WayTlEB1HFloWycMFZLlP2ppMmbJqYRDJMRzgL
eChlr6pzMTQ4cj6xkoD9pI/CAKuvxOCAXpbL5O91OU1v7RPIUK5d/PX8hY/5x9Jc7MYdHYYpIT1J
Feodrb6L6HIWZEJDyvjMCrWlRoKerAZxX89THuzPV+KoiMADSzpxw7w5o+68j/hZDvH9ITKoecPv
NO6ztYCdLsQtsWDZMonJvRxAEC4BARVENjnoi965tftq9yN42ZY5IYY5wynenak7Mdd8A87GgjAL
MSN9RTw4ZoIS95gq8jqvp0XSIUd2Hq290Y6Qf9y52zrTAhAGHjzzyKlVvQmj/DHrtuxF6c0K26cl
oJkNJa/MM/dO0tnHrnAOsAiP21SfzI3Izes/MG28UvVPXthtQQ9oYBsL++nJd9aw2bRmv8eAAPfZ
S4h8nzh4ySGn4IRwJAL6C6rh2VNpRoLNJDjDRiRRu+gKsx9Seg4qN2VG1JyRWLjGBujxRUQQPEbT
U9l6P4oFxLYo4GT9qq+OBd6Pgx1T9UZ6y1xzMMFZ09Ho9E/JE1M9QQ8yijQcd9NcUSG+5v0CIh/g
b5GlLZXMXBQDffA8LQhKAOS1YBUzqS4DIrgJXpKCXZQhJMKINFQuMAElfPK49pzUAyzyf5eZvI62
2fihUGx6/O/GN310J73AS0ye8mSpFNcs1BGcwSVPxmd0BijzCGQXFDPTYsQw6kAawkcYwKXtAHJ+
K1g4oX8vT8ilpbgW9TT1qPPHTqWtGdgeolEgoFARyg55xux1AzYxo14c3TEHTU1A6DBApSF+29i4
yQ34Dfukxr+AtTq70HyNho8MSMqL6JEILJWR/PE6xVKUEcNG7q/inqodLDM2dPmLBj1TL7Eox2xS
SXDjROCrFpWf4EZ2ctuAO9raaGwkWUgn5PHKO1PiGQ5k7VEPwb+94cGNjhxc6VvJ16RxbO4JWZxC
Ie8ILQt5T0VyWIbIAEfJHzKetyyVVUx+6nPfcKmr8iC0xjUGgQrpLZDhRTCaS2QIKM87JpBMu7Uy
Wf4xUikp6RdQYz3Ag2PmV5v3puY/vVHeZyBuIwADqKlHCueaZl8JoCk2bQV0BZeSpAD7ySFdKlba
+jDeJFnvlXxZBpfTpDaFCpcRygytd4Hp2JTcczuSEKLkAJUZmSUdZwEyrbY6itSjwXY7Fc1aASWN
bpgWJF8/wqQA3XFML/DoHHZD5nuujH2J6NMHyfrpx1kNHql/ssoeBp4xQVaJkjJfD1cgbLpSiqIs
Yd5R6pTQ+JJBn5eu3TVDoaVJHxHgsdTdRHgqgocW+TpGL72yD9Fb1JFIHL66NE6f8Nxo64Ffk6iL
yaQlTQq4PMKbQECYhjwW21wLwaRmQE31F0UjxPv39oxKT5jzSTPY8qjI65TSxcnNGHnfSv9bX6T+
1Pd8fvrorl4vVeRMROQ4w6WRyEpest4KD0pBRAR/hqOlOSXmp3SYQI9ksHFbOl77osvnz6I7YGrG
5n7XpG5K6JyM1MZgPtWwn3ENecsFEafdG71Yks99loN4IzxlNC6fw3U3b/4bgubZzORyDL5+o9mE
zwXWpLx61Pf6Va6ZFgs9bBQ9Np42jUIS3HcfA5I/c6xIRWaj94IPeARzvu1IpJU6e6zlAxd0oK+k
K79EeY4CusHftHmzbLHUa1sWh1aOCe6DHxuRXHBgry2pIsh098PzznS9o1Ll7x7DYiqq83AMYDS0
7My+TXHWLXb6Y/AATaEPkoRrln6GgAyOrJkvLUroBtH4W7AXnUlMBkk3uVSymGuexkeThHEKZMz6
Lhwxnq2VksmXpNDPesZWVQZJm2zglVRvAB55+NOXDud2M3aU4tb/A6PqdvgJVSrkxRHu11xmYGCh
e4dz+I8Q0/Ox4DuqAxFG/ExHCj5dVqcdypnsQu7mtcXZUn/NK7MLsX8mE3tMzKZBECOXGlE4ZlEy
ZjC5CZpU5XRhWhkCrYna9sEu0c4PHzRuTv8aY44TKIB9d65y8OkuWRgL+1HKFclROwBa1rxEnRHi
qdqqAAQCjYkRZU19R6YL3RonmOKLiOHOL+7kg02caF5XXALDIjZ67YdRIs2BR3Vh3vfW2Ob9jalp
7VKMffC4oO8xYZuiZPLxcDh1H30OGSvlgxGj7BUEwLAW52KdXYtvfUNETkbctQw2xNZ+TtRoGBq1
1UgNVS890I+y1cpNxj6ftZTZpXUFLAEDEBuIFqaaoKAkAA0zEN7VSEjeRFMkIxwxXtqxMw4TyGsp
S+m0IxKiy2GmMGa+lzvhB2hgRnnApQWv2oqzUMrPw6wUXfwsfK+AcdquiVDAbSfkOU3+kPW64Ie5
CnSHcNgAHIpmiiba+Q0+efiAwD2C//CPktkPxJSjCy06x/0xZ3c5DP1sRvJ8H1dSDueqSHw78NjI
PnRKzDPBguJcU143PligBGigD50e3ZcMiUttw+mxHKYLPHkKY1ZmLIPm7JKzA4PQIegRh//SOtse
lfq5yGWNLzlv18zoRxH6m7lIkoVQRCyF+BlgBFW/P9W7ZqMv0tyWCMcuyqLvCOAO5Dad4MSl7Aaw
p/JlcOGAEfqg7Q2o4JIfolpNlytWKpLGu2rJYj7HGgv6nLIIgqnv0e+CYMiJgSTGCSIpnzYuYYoI
u97qETBogiB8lc84iHRgzWvHGTrdaXPhbaFgJE89AdYnseg+joOKKNvXlJXoK4U8/oxU6F98zD1J
1M+gur+Kenic8myQAExR05oDaLOa0/doLeeTvkjb1qmuFnsPrdB8WjpehUhq30yZS3CZHH4VsblW
f1gPx1Obd9xrBYmIs418KloTYtOcqwlz1QTHORu9E7gm55hUYLkbrChhAXTKR7xrvX+1xOcxO4y5
ydlSWzZIxFdQMztwHfCuysGDQOyckJOHpcRExhD7pkgJFalfZrc+XUiEdj352Y6IAuJC/B6jGplv
DtA80qEY9A5MC0T1G2CnSvQXA5TtE0ysVpGhF9OhKfSFz5J6KShpx5DfHRiMpbYF6iHK1A3cR4ue
dJBA/wIhyhRzKpxd8YjmRbtGgYD8j7ulPmqHAAQk+W41EHBsmEE8wwZ6qhrtILDY/wpE0tdzNCGz
0zQbnnhfOrWUSJMS0rKt5nHEcxolfysVOEBDlS0lE+/VY3XgcIdXjQxnRzZ1bY4LtoDgh6pdoL3v
fpdGDiod7MuZgL8JeWrdCwqtrc3sRACJqlejBKIEBGUAVcHcBLpwPedrJpI9zRkapltrHEKE1F8j
aoSVg51TyMSyLFhJYPsWkYQi/wNJs8CGW8loNQFbZ01I+6uxAnMDoDHmfU5fSMbBgltm224eLRXr
jzx3gP82Pj3rSmDobH3g14KpVHaYKqQ6QHRNIr/XuCtXpzUhV6xCwtrmobZHw0x92z3k//VxJRmT
7tznaaPiqEeKBDwmCmd8v48fzc2MUTH42x7CDOeDHQDDZDh6G8/QVWy+60AYoUZErObeIy56Ceck
SUr4N332FGTFWH3K5NwszCQpyNZK/D6/KZMdHsfWisEuJmblFTmY8UUS0p4uQg9zVDeKVOETvAKs
Ymc/EObnDdxa73aK1mBG1eO29N3/ncXkcGKnmMxyCGkFg+EvQ9QL4Q9AwD9sksZbnxBz5honv1a8
efy1J18R9RVyapCPNXL8Q2/hGZwJbNHv5crXN2/zWAwYSThjzmL38Vx+YGlerVMkgX8OUjvinnSS
FjAiC4CjAb1XNQfLZhBOq8kcSPi3I218FpC9rKq4dUBWdfRxvEstxH1cpPHbl3k3oCYeL2HY0Z3S
V1wWfL9efLxFR6HDJnBquPHxuM9QwyaZtRgI2Uglt9BQ82WfUBUZ86X3Elokd4rfaBPeQT82HtAp
WuH/06BZSksjjbr2R2HTPx6bGN8nwTXBc6vCW2k2IM3iIdWpKE6pHD/zOF4MGoapjZUooq40IdsR
RtSrOfGOpmfVTxopFZxsK3qXZzg85lbx3l80m5gRkqsdSQZIBWJa9JQEzUXFkLjtoxhcp1IqssWX
ui3oSyekdSnQn11pCMXay7jwv1gYhNS8BeArWnF5aebACSccU1sHmDyOef+IN6L1fyPCXdo1HOXc
XFGHpJIq676Y/55lJkKPpEIUEap13yYRwj+ELRI2otkhADmPcn2cV+emu1XfBoDYg7okJawtPE2P
z7S9BgvooyExzf4twPmcP+fGgc2i7kB4/i98rmrX3VkIA1PFI9CpiQ3DWhEVOE5VQm/8OlV0W8+j
OFqvUuJFzPqJqZVeoe2t3QfWarrWWqFUgw3O/a8/kelxujy0+HjKdROiFh/PJB0VEzgBQnKUwBe/
VvI3yxC6yVNW9H5Y1F5cExVKI61tazcjc8KFTz0d2Px48QDRtFsmFmO7Xb2CrAsIpiz/kzS3JTlg
/9t+cRlAX2bpDDqOhQXK1sGYZWvZOWleMLd6fNjNwhqspjqfi0FLYViUJjQQ6+AGrB4AXVbD22kj
kap3ytsmNQDF+jLA2VbTpMIuconCR5EbV+4zHigZAUDYnQx9mwJIuePYTjhfz7RFRA4CxGaP+Izc
TUdrrhdEuZcvujVUtyEWVrVCMxpXZ45/zt5npGvEGaETa276T6EVEMbPycVNC4RDNnTZ+I2wfqjZ
QfZeWMsW0peymg3V1ErtJ/KYsLVootYQvPS4tuih6QOkfbcqrJsate95gyE8UXqp80Y2FYLORHuA
zG7IGS6TSTNLL/QuHm8EaiJvtc7GSjYk0pfhE8NB7mIwvVoZKtbaFwKc1DhFDsRsssIz0D/xm9EX
KN/pEZL6CTY5pqX8lnQzcq/dC8LPsDwFRx6OoO/fA7Lb84ymRcJTNQ5BRhMvLY2Xmnk79ElZmJJ3
31J4SlOvNYt578oHgJ877ews57XSemJAGHvnY2iJIhodol16j1+5+JlJRSLlfF6JrZwUyQMuwR4r
EE9csOGPZ12I+NApIwfjcvORCp93hS+PAmTX0YDGgVudeSrRZ4iE5oJ6pyVVqY7xOGDARaeIafcp
k4HDC5to7pHFCdZLwt7S+mYGZv3aLPIhribEBbfzBGBHAaPPxN07n/+23LWUvqdNIpaLtZm7PsK0
1JSI0W7xCcjDMTSSJ0mNFSnV1yCOPZdlBSO3J9qd0EefQGM2faaA8+fLroHEUOm9wtRfSU84OJm2
6jy7oZuQB/CN2TtCBljivG0+99SPrCkee4FVThoW6Dvp9+r8UYjZFbDXAVSEUxseepBhenWb63rA
4QoRmsKu8UbhlJeT9ulJ+PQ6yWePx3WVjuKhtQpBOl9D8zFyRLRdj8JP72ttpJH0X8uWLBtDBHUh
+V1rzG7lp+s7PvgybyXEjojMPKwmFnrPtavLZfb8eg3HCjlw5k/oy6uYLeCWwhCrVb1XWaF24Ukl
zjmym3ItMXstrUmMPtaQaReEIVqT1/d+//mekD4DrNYK7C7Muv6bH+oqiI4J6714x6ayWnIUPusU
4igNNS8o5jhF3FrjEk0vPOCPntN/jp+GKyZhcq/yzGK9fUyLqKr/9aniI/3JPR4RXgxMq56vw7ek
TfgMxz6dBpKa8A4Xkze8FHZk48xqBOwDdrs9ce4P787Z1qyQWDbtDA+hslKb3eD3DUF4aEn6kPSP
86mb1INYkYhjptc6Tg8gP8Vv8sxqM8nfsPx8jbD3aRkKM2LXPaLM8hljKa5mw56Ldp7yBemG9g0i
xyEnT39HQKR/3NHtUADKeLCj7pv7UlWgA8B36FYHVEy4ar8FBS8J5Zr9CxrUbQmzW5MhbDK/SOWg
Thbi//zb4J8YI7n8nzX9xMyont76TzHRgNKqM2HGMPgIRU5XWvkiZRQ/C2RKy1MjFp8uioEi6XkS
mQt3HMd+M1EgLsWU95lpU8sguibEUnbYcFk4sxQFIv1e4RAFqRVtgyJfwzi9gdFdvBTkNCV1zz3V
jvuGNxI1VLujyjTgbcoXzVqJmG5e0GLqx60P8G+Vu5cKDX323w62kZhdPQKmI8CadP+ct4PHLYv6
52i3w8ITP2dUPQlbW9P5nMV54c7YJBLDCSZsUKYHYkXpN6R9HFj51Y4U25gMNTD7M8E+nJ496JbE
kTn+nmM4Emo2dfr7pkOCtlHHH43SblHBdA1NKP8DGhHceE/29jNgoOuHCuEoL7cxigvBPwwJ93Tz
XMjXPmwuI9mA/Yb4wLF6nabB7DEGyfVKSwVPF870IX8392atVQKQYcIhRSfB2hVLmg6zGWS7TKaS
j8lNxZWxwS5ZViHdE5EgfGp2lMmfgLzIczJ+EXYaqmgzvHZS8T7CtAiGMUpzTV2RiczN65UGbRyC
6fLKjJ2McjtPUO/vl2EysGKSLDDXRNWiF8uCj+MenXr1UHiJGDQf4dPP8g2rMfG7nrpxdI7+w+hl
qmOQwAm2iowjUCVfeGkj+p0MhPts2F8wKpHt8PGmVmFGNEn3VG0ZraD6n8htByIzo/95EujeHvqk
8aFE5zh/lZYffE8+oouyurJ2df9+PnKBq/DOw+9d1sKQR06Hy7Fx3fVVIXn0urd3kr5ZOUm0UhOY
B7ytwWGMCBfxolwYQ0keI9X1je62HqbrY6btQ+t2liz+q2ymhxqBCyjEcJGabGu9pPdBjiVRrTXU
xfA6PuaYBwAFz2QgUPhfW7TEeL207Ng3HkRgnxYZ7EKt0jc/d/Wo8JrwPS3WMFltjQi00QWvFgQu
JyALyyiSvl8chRIWHtuID67LpydsEDFEq3FIMFZrAx4NcOdx/K2avrpfUpgaD0B+6lVjfQOlY7Ba
AcZRV1OxHhscBgcA7+oqM0q1ErGlOfnMpA+PQ6QmseVDYL0c1XlSfzmikoMOByLJKYs9zGSr6/lD
P5bt9Cl125blvRuzBq4/QdahJONKUEdaPO9kdMDN9pWEw7wCYIz0xga5rX857u4LreL2Vow6uthf
+jVu0R0HDKKqzaNQTvLbhErQcjeVPR1jXVWLFbCdaGp57vG9sAsbIbvwWGrBz3goBKDnpHAz53iJ
lwyhwKrS0ZfZDKADDNGRmihxN5lNdUMlwq+tSQyhS47Qok/gUrfz6YCtM39s9zvkzOAh2KAJom20
vFoYf34FodBWNSEwA0UsWqz8aedTsUwXFfFf15kLQNkPXRCofPLAaE5ZAj1glZsd1j075ehCnjzK
eEzAWEKkL8DRL1BvfPGfHUiJeLZIta/07DLCvfnni0IM01wmiUDiM9r1NfwyiOBusIB9BhH9/qMa
8pt4YrCAJgV/Pt6lFFbbTM1iMChTaLPCdVeNhgR3gidQzyTANILUZovf4HIl93DBCNjWK4bzY1x4
Enoyz3gE89xPqFoTmZ6riXL6XSNWB3mbXOjKoBY0B1Fnu4fJ7ecv25SYv2/qNJhCUieuyNNIVdTs
xCUe8ZikujpslXONXhC69/K7FuKZKygj0jDY7O4URdpBf4HCWf3lY+XsHYA5IvR+OW4yEG622YZd
zxIxB1+q1U4mvpGmZaRS+nMHz/BjKv0df2cqwJ/i4bYbhFK92Lz6bPQhcYXLjFXn/dCVy2TrUO3e
tQj0vYGZm25LKeMkYp8lTEb5Tp2eiRXHeAGeVpNfCHuMzr/P/8oDnZVMoUK+ghcFPCHgtYBoIPjd
schQpanfDAlyZaY5mMj/NhbOGewZt/gW+wKFLyn3dsZpZ6QplBOjX4P9Va75hVwf1gCErEBjtj8B
JYujLR/lGm1soHb0pw1Ca9sxY85gMgMp7QWWDW+Shs8QIoepI/Ev5J4TJd1JQTw61GY7b8rQpU3f
VunYXFzngoJuBXe9H87Y0xANqFy/kdMSlGJRZltCtX8ZV9h+ZtDuUMEEmEgMBDSACBG2QHgGR2Cl
o2gTPX+5oLh/f2TisjnC4MVa/P4knYRTvOcFouKDybR/a/7RDvcFzDwDQIVG6bDzkAgQ4JhjoBi6
qr56jb+y4LsCDFXomDZOp/q4szgWO7915Tl7/1m5fE0sdjfcmgCAZLnNHmOicTVMcSfTU/gswxer
gzd3wxplIiIBEUwyLk83Oa+XhOQGXSaT13CQY7B/YvNLZPxSEdkbbiE/tuQwo4Xsy3F43LVAhDt3
1vU2KW8lwbkNPauVcQIMZH8jwcMBxIL7lPeRbFx7SX5jbhbzFyP2jvtb9UgDYoJg0zCvS+V74F/M
Ei5V+mHbIsnqMf9es/Vey5iEcOPmbKWeHKkTtljmLDk0qJB9CNY8eIbm69AxaKh6mmbUa8ybTRUC
oTA7cG65C/SOn7KG6dK2y39at4MuaIn+LofpHoh5yr4LOrIemmht3l3QBSQP8VUpQEf6YzeIYqFa
LuLYeSNYCvwtgzdX8hVR8P3CD6tlzqYSHfTrfzszT7NglJMNf0GS9vjVSO/GnNsRBfEcUoWAmMJ0
9C2wWnZzOd9gfkKr8nJaGhhf567cvNxCmTqaCkhXgizDrudZVSHmtBUQkaHQj5r1QdCvemFVyAuK
MRQE6wJZMQWFzaDgaB14eUpTm4UIg4nc2pVufJDnFAfz1B98w4UYquxYIXt6yDBUKQG7q0jarHqs
6ZMGAv/de3j6kmFUJmwx23T0Y/8cw6pjm68op7b27kANMFiQnEt+F4QSshsKtE4xk95C3W9Y5mpP
k0NmjaMz4cpjj1hlQ4RhFtbeKLrfEj5/vjS5QVOm1CBCYaBq6290YLGriCzXIfmpRCVzQl0zg5d5
jF1qwQnjza6BsdFjcS28iobIHaHzPLfbhtCFZhfpKMuJ5c8xHjAALoFsKTmG6/5Q5Z4GH/ZzJJ9R
3btJ8B3YrsZfEyXMK3x/Wh2oJJDxeJjhMPPXPqbSsXG/FMRG1c/vIWmZdUsH8zaEE2MAGmBap3ps
2arRzdUWswNra7v2buZDGjTRZkxFCQoSkEbsV2MWbShdnbpdEDO7vLIY1zGvvDjeN9DbcJoSVszg
YamvYJch4ADR0AA2THnyyxekBaMxr7duQjSa0FrH5l0AQ2hqBMWqi9I4KsZ63ijfLmiuWM8DcAC5
UXrjoVyQYbLR2JjDPtCwxcu+f/YjvarUJx55xDgTMf9gprrzqgCLZD6nWHwH7QbsWD6huD7H43hU
FTkuQpSlSVyyUzAUxPo0bNw80u4kQwLGqMkq515tVo5+aezxX0hIucvdlZsd/HAE+0FhrCAuZZQ5
KjUh7FYxUPFMRC5C6d5HeuUh0k8BwYzRqOPCdb8FMS3mOs3h3+1d4zTC/FukKJUk9I+pOXmRajZi
yTwaFgna0EEyd42ODtoM4BWa5QR8+nZcyjmN/ZdSuNbF33A7xisKRWZt8iryZ8dJOYF3A7IwkNCh
Q8rt/CMLkWTp+bjZU1E+gmUYwimehHt8bOivR985X97MSNB/cRJ8XINxnRps4lnOI3lsS93rQ+zV
AjeKMXk2us66IWZbNMHHT3aJe1XU9K0x5j0TJ4xwMpzk4anqWMcS5xsQJ7Bq+RawbSSw9vsUCp8l
SnndehYp6rxnSqMj00Ot+nTEFEBQjRgk+AqYRLquMdHCzvKED+TpySTXz4WrJnbxIEi5YAP+xARk
w49pSNR/WYoExUx467ZrmUBmfi6CLQuT+8lSAk9mQU6yCUMYQzhEVVYFA3Rg1q5OFPO+q2z7Fayr
aE4F/UKamAKkl4OzceJpJwW2hGr/J6XLsbmzcbLug7LImWS+ZcZAc0BaFXnAlduLrZOgMWK5vrTj
cl0wR4mQ2oDyMqUNKL4yGngnkDoiJUe57QeTcBkmWF2jZfu14ndhfnkMdCQClPWUAqFPKtHLJBjN
nbH8vYMi53DUh0zUQXYSjS7yRi1QrBadd/aUxvC/btH6ze4TucrsuCJ2P3eTagyRDRrcc+JnK9Nt
iLMVb5WazoyVx9e1GQc81suAyWsCazMGPWfJhYTt7q5R9x59hXoL2sHA/RnZd5uclKjvaG3jRwmN
qdXV5orE5VxG6r2+QJbHlC844nL5nYL3UQ6D9O2Aq4ZTa2gLcp93o7U0ujR4Lii5/qbUX+txaYms
lao9iBXoysGrCCZM7wLJtzlNnQORh7y+r/iQdHQtHMVhq/GToqKXNAosQATL50fAtEC8KCL5Q8kg
PWiKPefRb8aP9XA9MWUCYiUSd+mRDRkZJkRqmyNXCZZlH8Hd65RqrutdSnUJcrf9fs+Srv2uGzv+
wEkaw9+L+HgZn2T+ANqXO1PxymDxYabcKW3JV8O4M+hfNhXh0m/lA1qc6a0nQ0RzWg3FPhqjZkR6
gtTA3vABLI+HJyeRb+7O6dpIAVsqZti0vxzZv6jrQukLyYvQo6k7M7QNt9VP9EF9DLH7Y3SKAEli
81lhFQtuQ75rPcLGz6ltXUoRoAEbFplAUCujaVpP5HjVvajA/G493WSPyq9qAfq//aGaRQHPrQ5I
QurIihYKdixB4mQ4GYBRKoxLc11x+u8hRXKntWlEUBG1l0tl/sczxHjs/X79BQnWPeyNYYFPK0Ww
QQPWOOsxnS87CqE2GNRvR0MqIolWx0zdkoVTB805TxSbhsGuzRZZd0CAeGKzYKNKZpJ+X/6ufSnP
WHWaHpLvuGId9xAYUlYxhAA2ww24Q40FhwyGXculNSD3dteuB23uSgs0zQbEtl71qRz5qvRSt0lW
Ai22rlHh+uqKVCPOmhrGySUSmtdGVv+nc22Dyno3Z7XFiNBo1NqByFVlxmC0KKabJVEcjgQI8H81
UWt2Om/JC8hEQevyQwnL9lMPnkq5YMx8L+zXAQTiKgrz522BSa5Wdf9Hi9Hi11kG/QOT0cUBFKde
GSwpnDrk+bFIubPeIFF1jxV+KUm4aGqByetMY6x5EgBmlXwcRoXXU6iDt2rrOqNz5z6/g8up84Il
DyzFg0/fd75jBYihfxo7Zwg8wKchd1X2avjgjkH7A0wW93T/O7Xc9Lpnxc91rufxsYJWSmtvVu2b
nYeawwtzTwApJUr2zI1E+6eirZbdgDafYBJOprY3JRPGk5xmJOgCuH3eX48L0IuFqGj1p8DNzUEP
UmnxIc3CG8Cvw+PeF7JPp3NXk5nDD3aICKSX9c2iMnNJCTb3MdXBMVoGVsj/86K530UPyCrxsiEX
ceJO6ek4mcnYcehgK7SjPkux3yN5H1cWaD+TUMB4ovzOHo8BD1RAXVGNuTD3EDVlLDR2kRx77SQR
4Kuz/hKNM6zfQ7XxsT+4nA4xqFCWh6OfiNzOujNPwaMErPfshgt1VHtzw0wZoJx03o3+NNSw8ING
pNlDQSJF/ioa2nGsRQTWE3oNvQUrKaLjWal9md9yelZFp8MdrIT47K52EV0tQ/1r7iikKt7zg7Ee
R9dLSO4gHi947GR4exE1pYla8j5aSDm5UwCaLsO3AH5E+SgV0B/ZU4vuyAhxSjRZMhWNLEXBXiGa
2gG0B8iBhslCq3L/tO1dNCnVtMmJugD+m7+3ITU2jIVKZBGFuVD9JSS1wQ57eSc31bVJcivlX1Qw
TqvdH7bHFMB2G9bVt2Cc9JCOcgGZLJynW6zfDN9T8XuRjriUYzLPwWsPmfKXZ9q8Igqn6/HnfP61
uadfYU0CzTPQmXIehSHmxF4XuxM8wpFzG6vpp4xKZ23OBkM83zBetWf5Gootny3WJc3g+2R9IefM
SuRL3UiMUg6MrckjifiWW9+3TnaOjV1V6KgoFZTq+If5bjifyI/LtjgnBWIB7Weu10O0ThrCS4PU
vUTAuclqf+I9KjCiJHjnvJlJLVOoYbr4L0zhJup+vDHOtTujfgepiGEH3ds7DnhpmD49DaZ5Ds4S
uQt+5GydX+vGM+Z0Ux5qux7bZ2vfdVOnXKbaai+bBDPQVK5yK68Yw2OiNJqtxBCMp3zfA1IkoSyp
bxHnvvGR5ndfJuDIWcEm1bSaPhHVyJLe/dvLNWmjipgkJKtix+1V1RlG4RQmHDLHZp+xBQEkpqaN
lhmqLWhZnTtWkBLKLCayoUn4KqrZNSL7r60hPX1HNlhiRQ5P7dOhvSARPyKOkvSeSzLkPkeeTVCY
o21P35yHnjxXYjijDNx4dBuh+p+80XCclMI1dPQWuI47OiPrW74JyCrqTTqDbVI9ux7JjiuomJVx
t841+XxxsUOeZcwDigewwRZggKuzuZ+pgyQHnlSlPG3XBUhBDedidZqZRAKkr+elWel1czqxRWJQ
vegGoeS2osu10b2OLj+S4Eql5VaaV/XBcJ3qFkqBXAEkRfwh3VfbxL2qDugQqICyxAer0iOaMahg
cJQ6mVz+LQbF2qzCPcyik06LjW/6qJl7ry8OuWxZdNbvDt2DxQFUe1fRFfSwpSVgolXEMuRAjSd7
5EMMwmaWzXKd6+pbnrKYFhF56hf+9uqo8IXSFYdXJQVK2oCmMUXY3VvbT67VVp6TlQzNd84Faoiw
SDAo80+vMSV8YSzo1t6P1E/g+3Fpu3Sc8fNnlhg36vtDMeQXJfu4ur/2tWlHRamzaqHkEhENzZca
3TmaU2tCnfUu4jk7HjGCvoAT8wY8Bt5EoecF9vpJlD9mLtR76k+2+k7go9rtO3pMTiD4TFEHrf8q
tG2u4/va4ruF3QPd3DwIWyLKtqZ92scviTsmdDFX2CAaJGMtCmDuXkjKUOTFQJyAJp7IPbhXglJq
JLU0VmHSyDAMLG9bpYYrX/LjrTxI3CoUDq56d5SGRfMbREZdCf5MppqNUCBMRob9T4s/QNshN9Cc
jaAXHw3IlyENy4IaIyXlmDZkKuOrlyAk+t2m0XQ1RsZ+0xNPgWsmKv6zeDJy9n+f1THQVjXL5AvU
dFGa0BW61he1Ts77oyg/WhLyzDvv7yxuIl+/UJVS2JtFiAP4COiRRNxI7zN5BV88I0ydXuY7XAX9
Sv0vDlJgJy6AFjvA62R1+FkkJhNgRu6AqRhaEZJFtyxDsdyPBhslvnoT6ozxyt+1j9jcKTGkjAt3
gIsNcGrPM1fMBCJngUxGJprJOBZHY4eypDDsSRpEBjnywbZhJwrmLeFIuFRV6t5j+9UpiaOlDZYl
Sz4fQxJzKWuUBkz06kBav6MWjSWSDwG6emNmrEvpj6EHalrX+pVzkRK33F1HQovJR7qXUTucR4cc
n9yc+T7oNwdBoOz+dMn501oveaGeROS4ZdUCvnBC8E0Hqj3Rjk3/PMLK/bIRWnAN6kkV6Hc/Y69T
CrXudjDRzISpzNrYGV9XPIP1bMw6uNXrD1Ur+B5Yj8TgiChJ+YdL69s65x+EPA3vMFKMzo23GpE5
WDxzwP4nXxSQfjB0pn6wQ7M93zlvZvuLqpSz8tcDZ2LVWKSIaH8ljE0xZ2uFyQ2fvd+0a9xSy379
LspYM+6votpikErv7APG5o50RQ2YpMHm8U55ipM5Xaxi5eDVA+kL6qVk8jNvqTl2G6LIomTWFXUp
b5R2/xP0CAgo4Gl/6S+IBDMv1VujpXaahPTfRT8FTcj4V4mPaYDGPuFHkvo5SARySVFtE4NcrWdB
p8pSShUubTfdWVNSqzfu/8pbIY33z2j6LgrMvHnHTZhJ1u3/BO9cdhH9wRMePfTUyRB5JByYeGGc
g6vGm2KAb32jP+Mt2/y51454sLOLJGlVhmd5/AdmI+A5TDO94jIgI9k0mk3q9tCe4Drlfz5Rlba/
a88zZGvHsJZ1f60t1WcCLvI95cfVMqbEneBtLuPsPMMuOdmZUNvoG5YfGvYIgfOUbSQm1uVSEV03
LajiYoHPRYJHOPlh+tTJkKX4s4BPYJDcF86Iypj2Re1W8mHidm9hpWh60CXjeQvI9WpDT45ogbTx
luE5omgNK9nx+js3WrB5Eojr6DVHxVcBSnKgzrZvrqFY/9OQ+U4pJV1yMTTYVHlimEwt6OMs7vKi
tzCy45r5IIj0Hx2VIX8s4aAnHW9Rwz2g+0byOrr7aiO6UJ93tXJzHvK8nHF02LMwZAfUjbzB7cQw
YVycjFFE0SQSh2JMIcwKzhD+qjk2wWluYVKe3uVA5Z+2K9EDy+N5biz8XJD3ezXGiQ2tHAuCbcKJ
EnhTAPxJn/VSSTLX52DP3qeaHs6/tYVl320VdkmJNxcmrDomns65EdeuEWFLvYrUm/7z+tZmR9iW
ZKjaHbOj76K7iXR37nDZXGQEDUhUwSKHwc7AT+PpUEXBIvZRuD3Zk83RWzwjnOplbeeWPnWiMwhX
X/jFqfhEV/tvjXiM8hSWktXDvvCxfLhoKDvOU1hiY66fcdr1HTSWjftDUn4yfDxQxltdk9Z3r0q/
ogXNTGkfPrdECiRZs1TSb8mrYcJgoPvA3byKk4KCr1/KLDyXfgLlT58q00KJlyDigAXZZP3MbpgT
DXJ9nJTTqKnsi9UgGznfq1xKNB5ALpo5spRmayTklk+aBY9nJYs8S9/RgIwW/IS1QDYK+QcaLHEf
LPvfBOsJZrVefGc3s5srYlFO6E0tDg2sWjcDtxyunH1BgKnDBhw+1U57z0S/qmdoiDryjD5S0SfU
R6Y/j5mF1LlooZjxgW2GtbjBen2+qjM8Wei/VxGR6KIFHWC7bCzkDvu8e39/giY/YLDQ1hk3grIz
fPnMxDo+f3Bg681QP+2Kb9zDa39xD0WLyjv4lcc0XF5uOTCWTjL9YqOfNFL0rPT+SGyUKJooBBIV
J7jaX4FuFcRknga36KEY5q8ieUkOX7eSXtTytxPfcSeRiDfr7+8wcZb7FScTiA3C2OaQBivU84d+
kM4fDg88hlviCIRHZ6hq84H/JoyjtlpDq0NONO/zfd9v1U5sciy1LIlPZMFbpYwdATn7q1gbF8df
AfthxFP8194XlC0QtZIDyqKbc3A5Bym2i7k56g337fB/sVwQd9YHm2GyLw8oKNeGqjeDATtwzTyn
ko1xCaKpslCVa8ZqnA5vtid0Yd/UmkvcJvcoWS4dnAKc0eTR4O91sONoIi9mpMFCt7KYj2LIttwE
TFni2SgxEGhD5FkrHSwRGCy8oplpBMaCYTFb6knYpoKYBbNcbx2Zcz6SD1kgvzBLjXzhTpkkRWek
DVshKvtjRqS84rXjcRt1icXVM1gPMbcKfnIMC69R2ITvN8QX7v4pQovLM141DPip7oioZS97OSQq
QgzaYWeogq6+o3qkcbOJ8LNZgItlHffl5oLAjCHOb7N4Hv78A4RfOuG7xbFYNmWkHPTgPiICM++1
SaXzgUn2IcTa4wDGxCpZAOyfLbXFX/085U4Y5KmriJyA6Rnke2kraF1edkFpL5Fpj24kFcNYJ8xL
+8DJ+/1ja3tl+XJXYM1BXI1Cmi+CxZ8tDv/hUJKXUY7OlIuIfo1R5h5+oCgh4Qb9hgUviwm+7nNa
cJgtw26E7EZ/EbhMliz2UiYkNq7xnAW+4hDViJGcQ09IPWdMrjkBeCAuvV1Ruj66oop3NKT+CXlx
0SeTDBjTW826QRmK5tj/y5rJW3q3GbJF6F31GSxfIlb+XFFy54I98YWf85yuKtDLK/p030Gy4X5M
k2M4jvm+1q2Q6dVMnf9vbwntSNiMdqLRJ+vwW2uT9DXte1JA7nfx4+eXILe/FxE047PHm7AhM4Zn
3cHy6PNpo2fW13HDBiy5ruiUeErB0YApv4DihAiQ+SgyXTj5RAZbUeBH/GHguVggeT2PFQ/XuF9R
8xvuWm6DW6BieZrDZHv1JhEF5ekM+S7M2YzmurK3mwQtUdBpSxtCLPzmhjdGMcuoYlFtoI/+PblW
qkiURCtBAibrEB1IzbIa+QTg16ea2AYtJIcKttNQMZLxcq0CAQVZjPYGY291M0VcNuZM3M40mX+j
PSUjpj3/pdmP5OXzK9CDp4c9cxGAc40VRcvgcZLJaIM/VkWlXn5Y9Tc9bLET/VdM8GXMqBXK+vai
9a01kUKA3nB17LXtAxyel7+8urNbrzD+FQdzuQgG5t035/urlN0JoJ6qb5QRMTac83anTDCvNPas
A1sglpwlHgg9eMBB9bsLj2McKCOwIWuUW6tQ1i58pK2uHVaWwdAOZsvK48vIHuPpdbg34Tkpm32L
bQp8w3cej1/rUav+WASrAI4ZbWjAs/NjPANbp/dsYWsGkC3483Rnf0pUo0KiQcdYTOGguRRrabNr
NJvl3gbZDREzQRVzBKYAj8Kk3hYYvd5/Z2TwFSzaatNLAUEl4dwWHRHkKB+eAPmhxAh0V8dOKukw
QtBCYhhnWjXhRMYshF7ya/zjoylzNCLJisUgKWDpJuAkp2oiJMDbpkS3YvfWaXM9tnt1JN1O7M7T
CW+m/FFHzoBQWMhPOPDUCdBsFM4mEM9vdidzhszEYSmWJZFuj0QI9dyM7DilJNan8Km7e5mUOxwS
gM1+xvBOMFIlbcTzECr9bbZGw5j+d/sDM71b4BvGeBO8TJTSlJ/GjfiXLpAnj8/2l1k1rXivROS5
D1OoDgO2bBOtJVXqYurG3pPGTixzGGPIpS0IifduIh/W1OhqAd6ya8mc+x+dmUiReI1M21ekcVBA
Mv4fotchHVkCSWg8szoaE0TtY04jl5j/cnQ5JSa0QH4WSGm+RkJ+bC5Fzub/KJDiX94/XfJtgkS4
MEUi82wyZcJw379erT8A/s/m+GgLG63Hn1KhyST4NIHnzKNRM1NzIYjWEIgob3mCts54OgXBf114
9ehZ5ELxc2veX8kHRvo13c7LunQJiWoswP40+lYttvvlLd1zQOm9YuUoD6Lt6rRnhEGWNW5PKbpP
F1mSvWh6SRqTZ62gKMupXdXPgsG8Ol3jxGjeGuiQJdx0m6PGdfBJL6lvVEG4DNRa0zeZ8Qb0aGwC
Vq+hDayLWTbjyOjA0kV+Kqs7WjKIGWm6Lp8lfdetVoNDLCQiSYCo+tlYvbTyNwHjLdl4MQdacrrE
xlWOhvPX91mcBuPVs68bDP+sCBUT9B1uoG6EeTU3RvpBGCr6X3zcyyqZ1x5QOwCcbH60syfdgxyu
hWYaPbVnqlNiSZTFUJVnPx0NRyYoZ3s/vXJUdi5pxoxYP8BfJcdRpUMX3TxEp1s7VFT8wHddgptf
FPExbNFk88iI0Xcocm3RE6wSJA27Cs+hWsQeuzR0U/5SgexDFEQbJh/0rZipqYb8EHpNBVaHsBn8
pXa0DfzacVzKkC0mIBpv2/uBeo6ZnkgYOVL27SsH8TwQ+6XrRE/RfaJWljwjRh3tpmFv3Q43np/d
qatnddKMwfhQBmBAtZvlFnQ4vqr/sx6SOI70XCitF8C8REVyWLX00MLvV5LBHlywK6p3Vw1E8srX
HGfAaoM1vL6cZgl/dYzLzievqXlrJJUkudCYH5Kt6bgIJsLoRXfVo9xrtKd1pHVmZO0yJdguSElm
cjVOKAbSilQPZC9zaV3003i6R2GpXCW2lXFQ9UBXeqfUwAIZSHeNOvFnTqN7TsWS/qvdepdZgBy+
G/wFd7TuE5uiwyVVeH1tZiTI04ys/nW5fqA9DEJ017a490xCllmPg/hrj+a7Rp2FoK3YLiSCoyEU
0zaZA2bUGFHkO6Tt50M27Nucd5GiGEML47aeuAMigdYLmyNIZeIwVOsWuYkzFvkzbhBOzMnrNm1L
2XYDtZNxEu2pPsXeHkktgPpWJNeesJjuRB1MiaCEXSCpHV9uJ9ZyTuFdQcbjUPzhELbtQxbz2Wfv
Gixr3jBNLOQcUNL33ZzMzhg9Giqfdf8B7d3OVgSfkzki2gW6SQ0NtwC2xq4W66/xp3qOV1LwCmnz
IUZ4i5wbFOPJcGDxZ0WY3kjbkEiTPdsm5RPnzxw+5EJ0fRC0viDumKRA3Mloldt4Pesyjq3Dtkru
DGk5oDq6JT1OeNXAl5mNZoE86c2lg7wETHVp5wYfjaKJ165siIEgkXPuG0alOgNhPFWENFBraDyF
Sn5WLnrJCjLeuDLxlBdWwTFVxQrwLF1SrS0Nnt4NwW72F7NLA30udRGdsbBaADEww44hJDkEs3Sk
0IzXgiXeMbhrV/dL+eb9A4+SNLHgvL4YAmeuEcWlhHAwsocmWj6RljE7DVC39GcPqhoTfZQUpzNw
VsGD6+jJ5gwnW4i3p1Cq+O3lr7asfqbZ1Sfwnb5kiuU5PTijHL1/NXqp7nNsy1Jn6RvBrVznHfRQ
6Usuvz/WhJE9hGOMDrQtkQ8pf5OaX/Wj1jxAE81WDyHXRKhgVIQXnX4IRd3dN6Uo+xtOMRCQT2ij
l8Eg9f970RldxlpUJrz5MYN3Y/1TNX/Gp+ypqe0tFBiL9gU3H0TMJIhmEd5mVQZXnwhDZeP7ONbW
3ac2C/C7W+ajmvC3wK+YTgmgq0W5bj2Fo11AEMkN8Zte6NRax+GXjU8FSZUdipmboEM8Zn0/cn0Y
rrZQ0lN+1DVjhzYCqARddviSqmyQUqFekwK5CRWc6d1cSZ1XNgNza+AqQM2SI15bupMfwYWoJVmk
WxipZuO/QMup5in5WUpQW5HP1hVlyRp+9EltnG4WJiBO8/h2bixgbjYL4aFpz8v3/WziNwECkjqJ
0ex64DVaxoJkUFqII+Btjm23oIEMzDdt3AQqn17BSiMF215c8qvYvqOvPb66MRME1cu0lR+q7x2a
K6l5XgRC3T858NRhBQrOeBTAjBS03aWF39sdUwJy/bfv8xswa0Quvf++plj5JAm4sLgz4h/Zs9cx
I0p5u74Q6ZzUQHIUvjJpI2Bly1d0OXqVCEMy8bj01Azem4VCX9kIhqdDy/+d3TOpGX8WQIiICi+M
4wAeIAXKq3YL+/4KDsdpThxG9G/c2yYDHJ3uFdH5Y0pMLlKaXIn48di5cGTNlN+GuCeA19GuuoLP
9ztsoLQVgnBDSZExlTCEjsw5CAYipY2SIT+Z8ctZjpyg3xiDSj4VXisW8T7JeJFY+Q9BYIm+4w9V
tPYrfnprG4/X3S8GUVlaq8bSMpyHe+PfPf51qVWmAxN/WSS2qpgDSSGS74mW5GZF8cLZ+8pdckqJ
c7IstwtC685sskvx3QjmLRAkpW5SwdOYmBv4sVPZlmt0PooBDeMZzro+Eizbzz6UE4DZRRLQLa8m
H7NdPtYYMJcEfvbi18Y+llepJXWwTwISRKUy3eQRY8I/nshKmW487JFS6ajRn943VnwrI7APDV9r
OIxY3jH+SZiQ36ZpZk+cJkbK9ept3oUrGFPBlT2LQhejeh/Kx6ociKv7hDNT5GHfEbKp1MAf06/2
R/XLkCt8LZb42avdb0sXfwJFm5/aWQXE8c9al71DzhTqA43ZzkbP69frXp0XhKMfm7tx4Bl6UDBT
KdvFz2NhRZn8j8yc9u9JYjFixosfYOrUQpghpQwKMKBkkRK9+tBOqrJNwmnz1X1a6U3jFYuVwWux
5Aha+bhgKU7LuQhB07I+O98BEvahPnCGoEMbX4NdzFMVKLyyl7AL3AqVowh8KQ3vl8OHjvvfVq9Q
jUfRzevPQSk6Z2+8LdWvm1Ih9llVMG3pl5zJnS182e42VthiQdOCBuOCzY+ouDn/v0GfWgYbmtyU
bhC2+IkrWgrIyYtEcB7xzOuQssEJrgn6jGH7TtWsT/EViijcp7vDmCZDNHGRfmAdOSWZT01N50Av
QCuuGhoAkxk/D8iq6HoL9KnYk9YR6BH1vMTAO4jutAodKuBuufRZmPdBwSKyC0z3Aksrb/5eCf+p
970jxn4VRCr/p5LIDnxYc5a30V1Cdbie/+b3876N1S3bzzhllf+MZq2CjEzkoOYbQzZiKasU8wqQ
2X6QiTHV8VU0IxAxNf6OvtJw3zIz9S25K2c8AVviDwl2tp6JNeYHFZ8ACaIks7FdPD3XGNoRqg2f
pAvUBbPxRDMoPu+TVpesGTbNrrrueZWqScxNbdXSB1a/q8gkpbsFPHDuPCBxkQNxTF9mY20Ksw6E
B5FDt2GRSoMXmA/mFd09PS0loe5yBzNngwSp5UOVDgEdpBreBz9iglitLCSa2j97Olw5avtfoM5g
bLJQTgYFWnxZEhJHwMzDWVGvBRO1Ct5cVjZ3dVv23o9/gt2zHuVmnDoEteOxjho/Ee/MDfwsJwhh
s7xrs0ff9iEjVoTYsWBlY0JHQhfC/P+3FC0Z/v2bJnlLhDf2dZY6JIXnH3M2ulQYGneE/bz4c9YU
oeye8U34JvF/chL+2R3IWjlEIK468iuAG+5ReSMuyxrzuBW6PKNIhebB2QFFvO/26FezNVVKpnIB
47YToSAoj9YmaQRyf6LmTo+LA3VBphsxH5wYXHbLeV8S5RBAEDahThjT/twKvgHhTYTV8k88J8L9
tSNPNwz+PySsFc+nbxMHZcJdEOfjG0h2c/g5gx2i1/C0NWGDeGdDeq2zchg8pLkKX/Vy3PFMy+yy
HqzRwZcj1dtLO9fxllbKOMuaiT9NOIlcLOv/iJ65lybh2wUEpi0YD/c1Z7sDvsH2vANsQwB86dWX
Y0YwdHTDQA+giZ9GR9Mgg8z86OwCpqiDK/6KmudbL+UgHhcOlRXxbLKYa3sJ42HjXs01/FbbJoBH
FClSjW0hdufL2NN3hI5ACvFsqS9hCeSLM7rCjiG4+ovE95TYgoHaChmbSfEAOsmCNzg/V+QAsXEy
zNI9l3rDzcBuk03+qwEq2IKZVixB9NdoJI+5CzyTq3rS3R0IfIYB4ZR8LwHod08w+/iEuxZcLbv1
0vcDImNXpW2x1buiwT+XjUO49Lxx59LY/vQ2zWzTWkuYbHxTwp71lqX9Ptt/ddU72iB5UjXO8cL0
vEx+55gyGUJfs3X5+d4rG1phNFbUkF36WJ4CzELFpbAtBDRFzDXvz+dLzTqZeZcj37QnVNvXIjg9
QRDNtJk1N7S+s1lTyfh+U2rM0NfAhnTOzA58/3Fc9l6ET7iLpIi5y4rQyP9oBWtmazCbBT+4Qikl
DfUJKkhEWU/Giw3cYZ7kQrPiOA5MDB4djgy/b8oKERV4ktIuvru7EYeII1GrGZMgzcVmvbbdk4lo
Bd4E/kAx4I/IowqmdsXRk72XnftsD8nxzL1V4WIk23Ulyg2Krm4LmJmBkImBDRYwQM5/aYjLyS27
vbSVfHa0+Rlfj9Ky0C+34P2cP8g6e9+WN7jG0lgrJTFEs5qsHdLQpZ3Q1dvk2ocAEr+tGL/IAurK
cUgwW4kAdw+0m3SjFoYK/dnp8pMmhIGA5xhFBoY07Z0DrNl+3WkweUjLpgB7ngKizgAYZTFTTFJP
e+pC8/CIFgT2LlGe3B7u8aFH94Z5BEGB1X6dJ0w7mmfAauB3e04ozvX90MA2vFU2LrYolK+nem+0
mmIq2wS/1IfCs5KJMuIGiej21QP72mo2eS0RR/CzBEsSjbHmzlbwyUKzj4qDIRWt+KB5jy0/y6Hf
TZInL6OdBHSIA2IasvRpi1YfSsbpm1l7+DlBuEeRp/bOMfGWuth8KyxiQuiZ9kxegmDN6+836CPD
1nPoquY330XetN+OpcDpJV2G3AlyHBU/k8ac307urF89fpAIJwZl0qNOVcc8TaXlzuhg9/yrft3v
wLXeVV/u1HVcHiEu6hn3ttvEf1XjeCIIzwt+f2AfIq8jdFeo9K0LeXWgIyAlTDpSKkH45t4v6qK2
Ce6S4NWsUcswglBSTK8aPUPfORhFZXi2YutL4EK6TRph7FMJlUnG1AvPOVJCvhBahyidKmoiEnfx
SCeudd+PrN1QOyM8/AJ10y94MWmQh6cGrJQ8C+3FM5V9FMiJHosXktwTZmnQcsfYqqzptoF1SHdM
foyDOzu4QMra1gU4QWjISmLcbnrD1J8s1oFAV9wRdT1d31QPJKlBbqxZoLb4j9cQvjH7D/nilY9+
ry3HsKsfXVmF0IbX90mGiO2ENbWJGUsWP/hJYJsxiECwRV4ogII8+Ht9YSHRYGPgjNeNyWuYImHX
YOkmYqq411D32VKyRUzJvmfpk0u6sZLvg+YVDc0fLXviXaPYoQlDJrOAkUI2FvHLswBrr6eG+cPF
THe+4sA2BlBgL9APNlweKQoG9IDzBj4CjywiK1oKmUU0lwaRFtdl0RZr/yQc0f16S04iK04ifNHF
nRoJ7E9ouSHQlpkZY/1scoO64rzDff+UG0MfiIVGco+m2VnOh3D8dBk+PhOhe1lWdW+lHHZIYIJK
vjNuHI5B4yeIgXtpfXaM/gkNho8lB/ic2L0p9qlL/KwSCzORypjCcsR/8Qe4Og1yVeU+tpKvqV8M
gZk6TD0tuaPYYlJ5K94KUscFBqp7YABTlI52cTmcA+01P9K+pv+8TNcpP+uo0fIgUjF/DEMuIxdY
iN8ftL9640vqaH+RWWMBsWnVf4YW9aMUteA8goMqEqjuY/PGB+sSRy9O6JEC+DqFkxOh6FsAsQH0
lEuwWBdCUexDiSCj9s1CMH/cq7+uGxmffxc7cXHzLTVJiwVIi8ZHlvQbpJ1wbRqRI7U8jBaxDaDI
WIsK91EfHoxnaX4tZkwke7+Si935r8og3aXXk51DOVtkKkxgc5lUqp/1l9N8Ny5XD0x+wKKw/shR
HOADiSoFcOvd+44fijkuCBBCyJb/W5oITxqft15B3djTxQE/LnKQm3ol77tpm87AZr0oSB9/iBWI
h9vFaHJ1cdDnUsqo84LWFIUUlLx/GrWE/MnqEZPgR0v/WEfhujmpCrOxgyZWHMcwzPqUTXhqnK3J
l+ByEvyEeuRbxeQEcCc23wrHPnMuOEHCFgUWurNotFWiILebZQ6rTVRLB0kbXge/amQsH6p9/1f8
wxvhIrzZ87vtocU1Hi5ZI5tCaTSwe7hzHPjOz6/X4Ls3v4agisySr4n1+5JPFfo5SLU3J5ohHF5+
Kd7s51qUT/NMI5Nm4YQJSOdhuDY0a3pmN6RoFTYFG8EXwlEn//0qh8N4FP1KA1cUke8lOl3qfAHg
tfgKmEWvF4eJByAqjAvhslG3vmXW4CU25LW2Z1M/UEq1Jnea2FTIh7kSWdDt49zBDquxnLV5JoXj
pKnwKT9qb+8wpRYd8qRo4FUDfg4zcUtNCR4doxJBmw9Yl/FJe30NXvlU3LSCtfzO+mibKFDuVaGk
5riIIItEJ/2NlgeNeKX4GokyeBCFd2dwjqTMnpPUVaon8CLEJHnjS13qpM3H8tZiYT6tUqrHq1YN
Cix7nXw9tUWfpm1tXjmZmFPxSZwYXThLbHhyhrOpfJ2R6SKACXV45dcNJY3Z/Rx0Owb2dRe0uJEo
wo12k/YAQgr8KXtY6Tb9BNtEMHwfpxjXdkB6dU0s9yLjTDt2K1Oj3kcHB4qHHjRZUB3++PxkKl12
ueL54Ac1vUox/Gnu234ZIeYaenBulKhfty6D+nM022ka7+lQh+ZRWKsXmIyeRT/1Td0B3vtb+u2S
Z1+ARcMrIqXbYNd2mRExvpKtP7LdPFTXrvyE+PiGqFMANHC3vVOu5qknGiUhJasODa+tKY5D4rAM
N+V+wjMD5lnMON04IKSWuDn3bZRvs4WEwzHP1+f+xavbici5DMk4odz2lbb6nVEbrTCeqy3UnK+A
jQY0gXo5DnnDWKh2oWQwf0fKuPmXX/kxh/OGdUrYyJM5wI0LxnbvJ2mSFu2yuv+E731Cj/TNyqzX
RCRt/1KSIemQxaUVfPgT5hcjWJGkCDqzak746H3cOM9E5xZDaVeAG3qRYpJssEbz8AH5PxCwvkmm
E6Bk+F/HMz/0qK9m7mT0iCNVcrcJrOvGdCl14haF5hEuM+EBO3yFWONY5hJYY8Ei/mQFOx62FxmD
zrPHUk9NaoJG+p6W/iOCpWXX/rVMT1+PWGhKYi3ynuvr0JR8T+NY2VQLN7rW9iL1bp9s2u/C8Ror
1D4efjIcDZK8VbkJmHtah501o5h9dHldWcEvtcaT5Zf3facBKo+WV/YG1e3YHxbBcCUwqgLcoZmL
HWoFBrac64zRlZ/KSjqdrSgk2U9k2eH+QtH0vNfX/qzFHrLJ4uHTCx6dApzdedNAEpRyYxCKTWco
Bh4NKK245fMuqWhG81AvmSvLY/rwj6/NPP0dbtKr/+UVqWNUtvdeD7jfiGl5sxxBRf5o0FbyqkKV
V/arZIcq2kIooI8jI5iAj9PWUDji7mOOKowoO6GBYqcKI3dDvWOVnt2c2JwWS5nNIsO6Mw91atBC
lmMpLLF8SUUJ/pvtHUvbdHMRa1vvCqa/kLaOewYYflXxId3w4DqsPF5fl+oAbam0rSKELovpnOKY
3WdY1oSmcztmLFNlZ4vPx8htynyRnivzD0hJGBb/0O3sXlJzmw28Ozk/PlcILT/ty4/rC45eop2D
J4QdI9zYl2bdDzdraShsU23wMZ4a0Z+N3hKgGp8FIqs686dXP4kedvSwEz7wimAd8X3n3KOlGcGr
TboeCeUEO2rqhJfSyYJlpoUNu6Bu5wsR957Gr9Nnx8K3rMSPY8ewzOeFOvm3p4TvnL4Q8VjOpcql
FfvMG111yBs29t9d2o/KhgCaJz9z+3b/pCwYtX+14G1315AXuR2fkQJwB89VsED6d4vhFeqxiqDs
YfkqZ6DAYxNyrDN9SsPzWpYfdBp8agS/FVd+di9jXtYy3l0AqzVu8Ixd+baOKSo1T2Xbby50gUXL
jjBv/T/TWSX2o+TpFFR5v8399TypcD+D+1YztRcJc/NgShsPC/Xta+yUbXlWpbSnuaW+rAbsdx7o
AWsCfHw4cvfJYxFNW0Kp8El87sREow844kCnMDvVMPo6XUIrNczkAcCR9QgF49QT1MEwjD6KVX+J
GP130WQXrRkWfG6KS9gacuxK6M6TT2APJbPRpZ+lzH2yuQdIiHAjSQfW4/Yer7xUcKkZGcSXD3b5
f1W1UHVH+s0874eZRaNeySR6NJ0FfT4txvdkJTIljoxawa3IiA2MSR+6m8BhbboWy9AJuvSniyDC
Sh4Cav5rVVWFkRSFvZ36fcc0NLbsJOAN68+wggl5VvQYPbfWe+0GHuLXb/jh+mesnAWEfCvt9a1p
f08Ec0mmFq0Njdi7Kugix6i+Q8JMTXKX8u5Tjn5K4sWpi5gEiUAlKI03Uk7xLDzD4SCfzUqCPBBf
08+U/5n7q16c7SQdsSxYlXrueXSO45/ZFMfyYCx/24WQyDlsBrBlELvJ46GLzuk6mm9OGmcGDxuq
Ygme9r4ThNDY6d2MoI25auQMhCXwrLfzg76CK2m5ZVwI4eopjeRK5rBmBaUsmOLY22NOrqkqgYDy
SxoROXsMJS0jPzh7jBuPRe7qnhnC2pPwqt1DsQ0JxFAs2YsdHNTlQ8BVN1QdDjJtgMr7h6wslA/L
HrpKpDa6WGMoisxxIdo22VR9WUpdDG3jLotCYkO9x4/rLEdx4asDWuXRWkcctXOLlnIsju+v2mfp
ozRwDOwtnP8/QJq+fOWg/JSSvr0Q6FGWohfHAwjVzmRRc+6XP5G3P/ZqoKpATDbZCzl0fiUosjvg
OLQyGDt33VbKDN++lWSS4hHU3Buv7xYloi8TugoQ0eOS2BWlcliqdmf/9nlHB+Fo4ubD38AaSV10
b8bGIt/SW0PmKwHxRW403/zWpQoICVHpeFxw0cdxG0/b8z0hEOAYtOwKna8cS2pWd6OUEuu/ekp+
FpyqhgdKaVdrAJ4nqMzDi/Xz9pYbnSfY+Jz/AQAK4mgakBE1RSD810dKuQnSt4EX9feyV0630Tch
VzEQqaDtINIfgdimydiFfVeOyGVQjjLK0OX5bVbjSUurvBWR+78NmzFlTOeeP4Mzuw7mxnF3G34+
BLRNYy5FZ+AEnygub1wvA9rdXXAl4sPmXreEJNFi2PmH3R5Lyafv549gW0T+pjW7GB+68oKD9SCo
4dHrzpo6TCWADmZc9D9D/qIRJoAWHOk7evMXM7+39BNyNNjwuDU6q467OuPZKGAjrMrqzXQn7tEo
+Hpu1yfYaPvUz3uhooThZu18hypjq2IpmNzUAOlriI0VF5FuwHfkWc8uiXzmREDauDd9kb9fBEqi
KDtC/L5wsS03HERvTdd1QfX79ZLUtFlBaDWU2/+oAt6N/wq0jB5umcjkotyZS58l6xPEZNYuUYt5
T15LUxt0/bNyGhmLQqHnFuSAqtOPFxCUy+2hGDBhJV1FJ5oENQaWKBLm52gAgcfP3vGo8at+esHU
po6IlPlPJQEBCpvqjKin9yOAnVWFZA88Dw8C5s6HByMYWLmm3sbPoeIJgXIeenO+pg7WPUKerKe3
nHUpP3cjGhimmqbBxnpzZcNp3W7OmoF4JhOfa1uLCJqL9GZ0PppaUgwrF1OZkL8kElkULH8tZAOw
7AvP3FvnKFwLomtihneF2W6rsavv4tsacjCFy0cam4rlpcI0+rImfHQ5ONXb2q+FCzXobTKm5hd7
WCoFdVGU0Y6gxExYglk0WBF+aYsOjiut76UgXBweEm+a+a7e11xjNntDwfH4mNP88gNC+wBxj25t
b0M4l+5APXIukvFp4jr2wZHvcrIWW0Wc+EgKkOAbad5bIWCDRDZsyvW6JUlxfC0vuXpkrF+y+XHO
sXPrVwLpAoi1g/4xp39mGQn2hPgGQR7uGro5wjX5cSPvu2t9WGqZdYyV7xXv0bH7uuGx1870kvZ9
tEpLiAvX6x8cjfRyAVMNXrHVyB26erFRJSllvo5dpWID3eYfh38F+anaaFbLaJgrnHij5NPxl2OZ
UzIcx/NMIwlmXDiYpAcgvZ6PNCy3Yjl6Ky5PNcIl3bBcd+i6fik71XiNQzXEK0xjGt8tQDxMqawI
LSu2Po4eoGOgq7Kjjbz8zo9IzmPqyhbP3xGfdn9S0Bppez3QugNqJchP3cTQ5Q9+rYCUIfrpVVIp
x4AjHsSzEh+HFz1UxnogWM53ngE6GYMF81rnUHmUWASV6+9oklxCSp5Hf/nNxXN34o0WGMHq+ROx
8V1F2/aexRu5GT3gRLsYHi9UULCmz5VA8kpnew8i06pR3rqBCS5rUJvAm0BuU2YmqdTqZAj+1VnZ
ZFf9ze57U6G5JPUq0MX1oG85dOtsr2lD33UEiQyGZVbx46iM0kpSscaumZwq11XLNGwNuzsRgUik
yK5IWewFpogMEBlJ8yWZfSM7gbVtxNesJoz574KwakcJsoCGXERv6pxyLo0nrbhSg3E/UOCUuTMZ
rzBXwS14O7HD2ikkCW9Jzz+zLEPh5RbT83HVNX/PL157FSxW8fDeX8zXw06lY47cGAuqcMzh7dDY
sRcTiL8TbTO9EgDkuH6iFFL1oz17yRzwlukGt8V5FU/SBYb+3jyUjUayxHXG1N4D5IZeXHKc/jgp
ia3LEDcucACiz7Z0b+wduT58Gp96u8SIJmV1+4pHClzAoV2gfTU3iFL9DLyuXubQDEWsZRqQEXvI
sxtoO/jnljMLMf0UaSe0q97KiIyDzWhL5cwTLATjrYSkP+8HuxqtXtVfg7SNgxmd4LaY4xg12cPw
gygJ1CHO7XPcbkKZMqdZKzW4OZ4qZIeD1kNqZf4iRBhQzTjVTz5sLEKxValn5/h8hqaerkzmVw1f
5C6FkMYyXbqv3cEUmAqPv2fjtpHqM8DwPwSZUOaQK2jPfz0qjpQh3NxixdyICwfLAWj4VbBA+Vhz
MmnjqVIZaFdDfs5l8zl0fBiMhO5MloIjU/vxA29BcQ9HBRhC55dGoty4Olig1mDz9YyeR8lhGKen
y/TxQU2VvcxW1+W8vV1H7I7n2oCiP85mv50iOB/OfeAqNkGYy64NbqqdGATwIEdses9VlrFI8RXI
RxwCqpEkkRGzQBpnwH0AJ9+K6XNwsq7MJc9RKcKXlYXrVAKR51dxJ6NKfVHPYnS6MMu9kW563kND
rKTGwHKDw3A7tAPlN8AU1CUXiZfaVtQrjRxaKZletpvqjIIBzwaK3DBJNS9NDgfsatyECpylDRSH
A2+Ty8jYDYEiZC29cSRMlhfRjVzDIAOC+XgkQsykonviNI0BQyqpWpgAq/08q0S2ltfi4TNZrJlK
eQdzqnaReMYccd/cBEzNw2bdl5mcxLs9q4l7kzE5c7CQzyD2d6AsibQMP/IDWEEkLCQog3H6rTTb
LOWgnQuPPSIZ6Wdy6bDB2tXygcqaZSImodYVIRyC0mcke/LUPlbtCKSa09Lrw82XHcPt2DSqJK/A
7y0SbdaN8y3P4bWLa/fkRzqH/GvGUo7yCDzjtnXJxrLLJWJFK+6g+erGkNNQH6IBHzkLvUYu4Rff
WjL7cGbHVgXglrxZGgWrdwBg7G5p+ad8bkOMr8DzNHRc65C5zZVV8MP3FeMDo5jqugopQ+ScXndh
IexN88tJL8mfosG8TmZhud/avU6FlVY+ehBTLOgjWwf+mkr6b0QrFJYySSUCeVR77NjDiiJ09Xsj
1GbjHzY/SwGC9VD5OEWhmWF7yz8zfKi3DRPE8PWvxXC4qURSLiGH6FR4Qk+Fj0/IdsXefHzLcN1O
lREIFLDni7AhVVqHKYX5cXXnkTecijG3V4cpqhS6pCQ330WtDpX1pYz9d/nK5w7Mo5sjxqo3ZMx0
M7+hWK2l3tA7f+jLtO30GSbo4/abYV1O4SNz93qRSr1FE1BSci+wL5z7Ijcdyk2AijtU/zKfDSTj
dZsb/174ePsaXlYzU5aUkgAIgset1j7T8g0x29yX9oXKmRO98iQvp6GtkuA26o6g+POzA7XoAKpK
OZ3e5Oe/1jfT38eg/MO0VYLbpsai47Ado9ftapuSD76dDjMweJX//8IY+LVBzBjFdaxPE/dVat6t
ZOcY9pbOuaaXGo3bAWhdK0A0o9SulFpY9tVvcnqRUGSZcZUlcXtcvFZoVQI6GnI0tW27faGhThbY
XBqwzysM9foCSw9mnPifqZw8PdDO6jnOEWsDY76h0GtxpfRA6o36MgbQZG05djsrvsicWbNnGLX2
FgJ/6poE6rLiTX6lxmVSolmbecsAZUHYSrGP7Gg6Y/TVqE52P9ZmyiHbs2uq3e7/7jMWAw3pFSIj
FEoOlj95HOFNSePSh62N2VfY6j7Q7S1YEwuocAtr21q/BoQMYlPlpGvTS+12STYv1fxbAJgwGCRe
JZxK0VtjqXGJSO318RospK4cdO8DzwQN2yn4nMcrxKl4k8jFy8qDBLqZFWCwIGifTu3gs6ZrrJUs
kiPaB3rGvREDk2I7xKwARocd8wMALuTj1Ahd+8t50CGJ+uQGe7YrIpJ89e3jhbtCJ43t1JaF+cl/
4GDU10iKJS4jEMDbUSVLEwoVPDN8xGES6cvlFYnbJsS9EJGJ2eIdVWhR9POkOmiGB+oZu1/oMdI6
MIGiaSrawsSo30M7ilkJb/3YYso+1kfokKGNstvFrXUUXiLeCMvvUWXVsghdoBiO57o8EwTjoZbF
n+N1Pu77t1IqfAMKGhMXrzVf2SbJzVzQliGMeDq12SvGlTcK3XJXKOjxCkLrbDUXfXGJZ8HSyu3f
XdLtCVf3u1GaZi3N1gakpxL19LeECQxnvpQhmZjeV4otvEtgQ5G72xIVgY5PUcm+6fVToG8A4Epz
T+r1sPI9vx3yM83mWL4Ot9br5jjn1LDoisra+xrx6EqNAB+Z78c0VyGIebpCcdNGfSzYyWFS72B1
EkwbNrd2YzeuKnKBTElk3iPiFmqO0JFivCnxpYxqMpo2MxwiEr3u6D1MTkJQkm+Vb6xL0M40/Bl0
IlWhIX5nLAmoOddGXgG4aUGp8mOSesFXmLSWojTQTkwYee7iMpy4LXOWUgHJth2EzjqX5L3Fh2+/
vYNFKyBxaARp+fGgv0NHlb2YH/2OHZk8OJ5iFXtxqQ06URdhggGAHrZy5WH6cO3xMOtJo9PNJzcC
Vmhbs4mQSs5iQYL6DkpiQHOzQVInDKfsIGKn7ryzBYNhwybWU1v/qKM+gKsC7Hvfcs59u41lhpBe
Bf+3iPGC6E9H0mw9Oe/nBePCKjLxN254lslyibhldfdTJ5i1CVTzJqv9ZAzFL9Oci/+rZwIL/y4L
+obRo3puhcJoojpIHUVxCuRWw2GZPny5zt4pAFALb9CMe0fa/57YPw+ZodULALXj1+8UWWFnsCuE
n3JrEODFDHC49aks139FKFg+fAiol5uIJQc3jWUWrWKNDvR50PXKF18PtE/cwQwNIUMwLDaE8cUl
mi6xq9XUB5POGOC6wuRU0CX/qRTrQHknpf8kyn4QwQF0GbET5OHULXywHv3OrIV4YPQoo96GSY+b
/vsJRLc6kRD3H3KVXemaE6U2CoOoVkfUqwRHUs08pbgp+zf8h6A0Ym64AKT19G/YVo+bobCTZkzq
U9Jmc3MOeizfFOU6qDvzf21WGhItIxOj9YBSuHtLxz1bWJkVrXztMlKhW9uOv/7amlzlvrgLTdvE
3BWg2DM+5PwVQnG+aGddsR0FeAqqWlkO9YZhBLPi+g9tl0t7sd0imhJYTTHwmMUfTI2ZC07lr6RK
hJzPZsuTDubR7jHgIqdN98woPED1DHuwmIgu44f2nr/9MAm1utR6xR6wGiKE9eCdTU8Kdx18JnKU
b+2wD0fSEvnlUwsP6Vi789sZvxAR1YV+Ht5cpVl8YyD1XdqOKao/PNw2a4mMK+m+eCI6Xzk12mLx
w5394baubuoT/YF9TqnkbpVjLvISisFuETzlLNPUNo4k7YvWMNtVidOHV0Exgq9pQ2lvUHqc4V4V
lVBDa6/Fmgt9lJH4Uthac2QPLZWeuCjEUUdUqTwGl2tylSYqA43tWeftGBHk3xLSIvJnWm86NboN
3gNHqwRTpB57M6vx+A8EFuoSF/rXP8XtOyJV3M9og8mObT3OGGUXuULZ1oBqGldSaAi4tLqEAs3t
pno2EFDsfP3sNGx6FePh1BfzwZOw5v9iSwY35x90+0iWKBCcQY0o3EcmdtaXYwwHMft+Fo0NwuFv
vrDreXZhql7hIHEhEDpzIvWTtq12mZ/HphgfikmeIY/9HUl4q07N2LgOB+fcrFvpnR3CXQmDva/7
318UwfBD5ldRS1fgYHwB5zxHzj0i7jqRuTmu90PdyXdieycn2EmTkYf2JfFKQ9KD95/CvJ8Szy+W
xcOr26x8pC4gSqEBOs0uhghKkpC8YJNq9hRzbeAFXYG3fvn/IOjShaq5LF+9KHF1Oxuq1EuJnGO+
8w43hMkxzyD89wwRy3Bvc7H8szr0wCBlEpXoRgX+O6l1zh4+PRPFeqhGyg4/9EPiFtD8kxvU1AWR
XJMq3d9Lz9bPT9A5VZ3IWSv5XOoXncx7Md4AhzP2OBc+NCDxge44rtcY2GQdYZRoKmtO89QOIl7T
DrwYD6RmQRM02Brvz5Qg9y50JhdbEt73YvY/B/uxKR4lloTZmhcm5rc2VQLJd7Yjhpad06OsYVHh
Ghb7Vl6CGaAdFHB3yxcNjldlrJoMC18Wqfa1DYStYMn6hah2eBwi+L3Bras+0Hsm+t2KibpqGpYc
xGwjHtn2LxOtwmbQeghByhJuNoy2TDNBgYk7dLpQdxhofqIU/maNuznw2VEh3QmXlfU1mjV7U+mY
NGbMP5xtmwEHJdQqQh2mAsc7OPdL1yVcg/JdwNizHU92fu3ADA+zDSqRvj57Hcb5AeciRXvLvTn8
ykZarSiDZcpb3ipKIHlptQB+h+oLIdXslkragSRbugt5E6S+JXXCNWcYi7nu3sNIiOocAfWWVx7i
XiYDXMTudaxQxvO+jMvBYYIVj1iuuBMFIWKJd8PI1LNrhEEraVR6Penw+2ACK6bKn0dnPFMxVBcf
q3Zfr7PrU3+vQjBSJR/ZUjowyZZ78EtoDHOlk8qqAIwX4aZzmloTr5xIX5wQ6yIQEdkYP5D5pn30
mvsBvygNW4tMobP7BVP9vTqpz1sWPEhI2t101E/A3hMzmIE2Ss54WOyQtzvNrjros+AcuG74KMlL
OwH4TVVKP/cQ4oZksHPXO/PiLZ0uywMZ88Prc/z6iz6yWcbVROqFACskG5gPFHQkZD/v0x9Aqp3S
IDkDSV5a7lmEKd3nvSMIpnYH1d6Q2gG59hRqmdeeolBrpYMy4CA5Atuz34CwLV0Yd0wV2oDCQC3l
ay0/4DcjE5UQrMzl1RMUQlNEMmsS1hKdbOFdAyNgnxxQRINNGDxfeVV14MpUn6HcS2226ZvNmoKc
Lj8Ya1csXrOy85I2K5C0dPmQ9i3/PXsb7rdejK2zIq2sL36JmcuxKXnQPhA5hYSxkNVYtMmNLznI
uCeD5cvlejmCVouxN+ntnYoO28RHj1U3vFQDXcBJIEnzl479uGrqUSic2MDKeRzTHwJ71qEKmfVf
ttbkbDxJ6jXi5xt5HnoOfhrimMLDCZPqw+ni0PmWMLeO7pCUQmKIUE6rAe+OZVyzun44dJ+0LczF
E1SqGt/qOrqxUJQID4X61/mo9ifYVr3nY4666jtXWXzQjvdSoZlYTzD0etYs4IA831PmNZUfQsTf
WB6PM6Jv/tb18IAUM+0WLCdG4wCtKV6ToE7ao0BcTsbYkROdJgxNNwgFPlYQMvwXEKFTVTWJhVsj
QEUHQpYY8idbvoqW2J8MNtkqlRDPwODfv0QLHFoJ6ZotFn2/yXeiut4Nkc9HJvY2uaaAKiy2Z/uu
G0Q0EbrOjkxshmdjxE2NQZ6QVW+QiEZa//s0KQPMCIAd6O31XNUtufvzqhz0BugfUqS48wAvzlU7
iok1C2m2i3QFUO4DRHekZF6Rap05a1Squ4w/E3ZI0Dc+v0kiN1sH4CVLohCNZjWFhwSBrEiXk6tF
Jmx1C9Vz2K3jmhl4vDfUqUqGwcgr1o5CkCuXS4yh3V2GPzRMLW8IrYmsmlg11UCwNglYvecoCpQp
9XPBim7hOMOo+kzNcPqse9ScbpgXH8Xxu9Pkpfk3VR4Xdz+6wNZnA8GpBVzcnAgbGoXiSW+mNKIE
KGNYpeSfL/4Vv4eQipnDch1hjtDf7317tR0riq42n6RVxVdQ7bmJ4MAngwMUyJnwwM45EPObuYNS
jLzqAtSUmJ7G9tK6c/9izMJ+wduBflcRzh6JyAvSg0WW/SzKHhwmVNmFTkVe1pES6UZUsW5m76KK
7e7lvYt0gBt1LJfBCEuSlb5djJ+M22TAWMP7bRZYi4hOS5hEVwJ9jd8j1q9xe3w3UhERyCgBW37h
qu2s8OeNGSec0z4tbzzISmW4OYgKTOo98uW/S5Fgq32F+KX2t7YxLdkYUxjypEdNrhICiXZJS3ZN
np5OGPLQrq21qlZPHPZmIpHoM0seoWFJrTBP2giXEdsBK+BuwliEKQVVJu5X/9hshdpfCP2RJ846
HujmuTmaEIkLZfAOoaRVBlncflGh88NRsTfgLicylVqzZwEhD9rLzhKq/5WJtYGX/0tjkitYCjZU
PHfY2+ms8Z/AcmXnuHBJn1q7tWaiGPViwvdMeJDTGgyhb02E2bLJOBX+7bxXJiXs2oBQBftFK7U0
31ldEX8o59JgkMl5bG4m81l4YccPC/kf4zYcETGV/AyQ78eUU6BL16nt8q5Vy1D460CbaSAo4l0q
pgxGbLG7cwy//jG9oxSLSdY9xEaYvytmx2geeiklt4MNkFcvMvsncI7+p2V6wQCPYQxvgpaScs0R
bbHZCd26BiCE15HKYj8p+0jyBE65Gxclz5mYxJA5aK59VsZAsYkO84ywhm9Jd+ykgDnfZpotUdCm
VdKVR07n7KnkdaSkFjPpy1bW7tslfxEwrVO3eAtSCvTmE9US7ca1BV5RiDyTNFWblCnoTg0gP1Qb
UMay46EjQ8W5IPK4qsoKS07lf+R8OM/i4ZzIdxVEoedQAfBWLAbnHu871iJSNHDRToJgOX/jhOp3
8hF09wwbAE4+ieeuMm7GkvBbf+Ntc41LMB9/0b0tjfd6S4EqyTEDVm6VpLWQ8cRiVP/5yz0gCpxY
Znm5bH4YNKXBYRdidD8hhDl+72OQAo/IsxMLRfaBMLg0Qo0H5op8Ofl4DW86bE+fwGIUNSGg06Y1
0mfhBaGEjfADwAGPwB4uPmeAzR9Nesqdk48GYJx1aUHi1Mi2LvH48L8wEo0qllc/dKvOlgRH26+s
dEgZEYcINPktZXpixSviaASPvCcStVPyEGtpFL/TBKGla1UOvqEaGDwAHhZE3qiqUw1k/qwBeGv4
VD0BbMx9TgD23l+QuJPUw3NSs84KetMYP/5xM71+v4BwTTiNcsFlMHGqS7GC2IDtDuRejWrkk7JO
AF0GJgH1V56qhLD/oyeI7lMCHby1n9d/MY3d60+qd8wdNqJ8z9rzF3ESb11M/rMlGrWzTHL9SJUM
z2NoIAOfN0sB5YRcff94G2FYux3EXMtM7+Xjcb3Ta/QWyemysWJ1xxW2F9rHyxWdv/UxRrB8BSMt
n1r0Y5+MsdEwFeOwn2O8LSVNoz+gjWmccOGzoMODiaIrh00XGMnDoK7EHbOn/34/bRSQpt3nUSbK
izq7X69T5vmDD7y4Fh9J6J67Q4Y/IQNoN0Oc9rzL0AaWAuDIsCreShHTrOArX0hX1C5CtSUvhZ3T
azJ4+XMoKPhJEHq4KsJUY37nwGLXyyj96Xi2SK9AeK0/GXqJhdZR7V39xwF9hk/noKKx9iJJYL8m
Uu6C0tYqXCB3VeAGV1i6yWwW81eFVqbb9nFF/pYTPQKt5DtoZciCU0ltesl5dpcCdvo54lELEveE
D6Xf5xXVQfCHGUsFoePuoWQtyo4KXx4WsUVqd+RCk2WOxBFht6uq3FAXRxb/gYV50D8qBSeJSBAU
OTbX62o0r7s0EjatdDxvklFETTY9tcQ79w7TM2BD5FbZ7HsOq4BeBrQ89zSnvT3Gc0sMD+9rcXpD
vxdZ4iihDmqvppJzjRHwSgsT3ljdTbpopzJauVWe7BdAxGkNxGaLzzE2uVmjPztLUU8eHxxbHMKR
vq0ux2+3ON+T3vQOWgf1F+eefGiNmqoWzG8Esjzr1gHO32ahRESX0BA5O0NSr9DGrv0hPLoDQ48z
wu/PtTf0XlVKpWpec8nbGFO4GiF8Ysj+2ZXHiY69xfotTmzKLmIrjqu+QeemuYynyZyVm+jR8kTI
qkBqnEgAxrYq/kexvPyo8t9gwClwu02GXKsRM7of1pypN6+DUdo1yECGJmsxBi0GSIU/YcKy/i7L
fVy30/0DNcWLkRHKsk+oruYCWFHnJ1Kb/ge5IVVUpWn8prsGgpq773LJxfPqmC8fylSWH+YWkhCe
p1kcFiNwsbu2N7IGPLQ7lmVzw6fb8zJu7STjpTzPkM5DnMBLdl7c8YSsfeFJjCv7erjt3yaCXQtz
JpiPYv0lhqQe9Mu6PF3Clot5b4yjJvFjx1haykV4D2wrqA9OM3xFxEqu48Kp+1q3Gj6gnDF0U0Td
VgzTvYu0EXyomZHngsLQpDgAtHk21w0v7GlxnkGYxmmgi8VaR+p1jzkoAqI0TQkBgthqY+rSOSD4
7Cs6ykYNjjy6pwG4qYu0CFLbqfU1kiCwS+NasQR2UxRLI5C48/S5ds5eVcv2rLKaGtwDC1sB2Irt
Jm4FuHYRiHFwh70TlkL2jyLVaS+5dooCHsFc2WUM4nD8F3OAdeoNdARlFTGI9YKkbz5MhnXj5p4X
Rcqw1jUft3i7YTNImLtcQYgRSI6zogzojowdcdHQoIDA7EiiniTWZdVygfYDf+DtCtecSx/1yRbM
sK9Gn2Dkdh2JZarD6yrLRUxPqwMbKuYdXlnE8gkItpFeZ59cs8JGddAE6NKVc8bugntedmd3zxWZ
wjCeBfRWMahDn0MzK7F86GtdIC20rXoo0qbBQCjWlo2oJ24wQd/DDvjHirTd4reuwjfPqzA9oWk2
JkZ4fHkMI7STjemnzHk6w5zjgObh0uC8HnUnNv1WtzfyKm6ycS0Ro9m1qIzhvXb0olAZyqon2hYS
ENW9ILn9hzVb5E0/DWnKm1EmDu1tED/GB/GA6GlJEZjNTl3bThhpqCaxFOXyc9pZ21VlycWObs+U
/Og+R+6DxyCNOh6wo+HNvxPPyTuvwYMS6z6WoNuPC5KmPb39ZbgPDxkJirRLDh63drffixiyUdbO
+X4AogO0DXRxMBTFaXKbUGp0pVk0Wpk/HK/46u3/Y6Fpsdm0L8e/dbhjf5LgFm3ya1YlJeMpd38m
HqY5e1TZN60XctBymb/rBpRrVzvAauOP23qHPSOqqZLgYn62AegCJ1+pxwt3Mg15IPsIiB6He6QJ
nlVtMgH/vu2nke1nkmHXXDG0DhCoS0E6xfa6Y+CADlVowMxQbEEh3ne6fkqaSLejYunaaXMk3Q1+
dypprGHhjygHmQTIJ2xqVaKfPlCdAt0BlEWI/HfZTWv9EKhOBmyEkpCQeSSYxXVeyxSfrS1D4In6
zuS9U2FY39t0QB+wQmIncu3aWLx9kAb4uQWrb2ASesVN9pxvElifCCOScR27iUrdHce2FSsIC9Zl
Fw/lIg2EarA+WdhUYUW1zjlPE0TUUKgn48fj4CHt9sUreiqmvECY9La84C7poReBiJ3Vq9NAdL00
gbx8NJgTC6M6Rq1b/A79Cw0hTKQvaAOMXl5NAqceKKpHlbWWthO85p4S2iFmFn5jOs52LF2EqnOa
ohDI02S2xPWWLVU5TMblOj7xjOZjtwTspURWD7lhW4RQ++qSmGZeV6txIG/t8NYltt+ps7XptRIp
YZA+tItGq8YCvCMG8y+vD4H4g6j94zlRJVpxknzE5AYE6cdhw/vp0JRYgswh2w0Ezih9fmNntyaw
oq1TlKC+1W4UQ+50Re2Ok02cjQXUPSjHBoNGQErW5IK02F0F9OKf2pVkLn0glTQbJFBi9tYfjqCU
1lW0s42P63B5v+Z64kirc/89cVXT+fOEAqJ28xBbrU7KUqmhDHXCnT9XahJdcrmr5WKdFeAW6yXX
idCWJDL08alGh8g09mjx6zqPhjYP/lGoyTzBLR4sKX88OibERIlxPMJg9DjXnowb5Ryt6X/EhVe8
/84dRmuI8yZeu6sUzr8D026XRs8Vk8TL7t+/oImtxzeVVpU7zMIm3+1vsAG/urZ2OXoWj+70MwT1
gG9Brb7a0X4ChZGLCTXvJAJjokZV5X1vAqRyn+bId6cgv/KbAok39bdOnjiuEtGfmnyWYl5rBpmw
gg2rt6I+2wLiEJqGzn0VapE7ryD+EbIB1FzqStSUhBhFM/gzgQoqQKpMI6uUv6BmL/m/Prl4UjZ8
xMWGHBFUOzEDAdTUuW7LMKwqcL7eBh4ZBLVrJYzPWmSsXRYGJ/M7zJKz/TOoYTVWADKNK4TQRr8t
zsTirjtHACp/PE0zuoyMVmSp0Fw6TQz+XozokRHCHK+3eLpuFDLHe01u3tQKJPx2SlhH6yHl9wKk
HiRUI6iQHd2fA0aCNQd2QL6NTLb/wYDl9w9ZsBg2sm9C/ETPfx71DdoVEugdFnuXS6FgQh05bAX8
Wq0y+0ioTJoFLO6PGlodgO8r3h6SdufC0eDammOinrDabqCIvOvk3IChYC2YR8b9rXr/tzSMtbOw
3FmYTz/QYlXKQqZdJIhBBCvd3sOj67l2J6o2p8oLVW1JZz6qI6jZvZmttkrZQ3MxQ9cV6V98thnA
vT13V+eMEHUQ8vxmIvElpYCOCSZCspmn0RSnCQ67sGK74x4WAaRLqc8E1Cow1l4JsyGohMQqFT+Q
rySzD8k/wB2dqXo3beQkhDATH18MprXpd+QF0VTWu6/G7xq15Yt02bWGeiIUdw5PL8RcMEg+zA8Q
js5vqNyozbsrUXOWqrg2v/EidiY5My98vFeQJlm4tHGVcMKVFH9J0OZefS4Jl5EoQr9Sdnr7FTg7
XmSYn7i/R1leUvZ5V+QPYEMNWmh6t1XPT1gL5+0Akrent4Ct2DX+nf7g2AleVfjJClXoEIAmQZgz
nB1bIdrE027B14cH2I5iAEE4soq39Jiq/0BiWzK52MwWiO5TBvJhddK4uCGTwD6ruqdBIeg4PMl8
fMi7QtQgLIbBxOw5gPZUcwrsN22NOQ6855DAJe1hTjk/tMxXe2l6MI5FYkEoyld1EYlkZDktlHnb
asdgTF4YAd+WGq/QZY8f4d0oL0EW9/ROfRqzSfvVYLwU8dmvY+m34RbaX3G76f/1Y0YPc7HZ5UYM
mn+Qc7/yAFpg0N8xoJjjtqI2Bju5rgfx6OyT0RDDBAA7C+HGufsd6m7ZmmAxhE0XyNO7Pyb7GkRL
fH3QdB6nOK0TY6hYOwrmD+7EqyjJ+KOFBxfbd+K0JgPhvFBbHQXPyvj2MFYYGd8z+tV+dnqlLQwt
4FXrNv1dKVSx5pdmHw/A4GG1RGjN7pR7ck0pOkI4vl0fTCVV2eP+miuxEGoY81ANQL+wP90ZVIv4
XbVCtjFX3JQ+0mI/9ZUff+oU3Q0E/7PJmX4mn1sqGaGb6YQgjH9kZlyR4iku73B8kvR2z2nDiYFo
OL1P9+ym9hXmmsMn2UedLHT3kyPRkPrH34uxqWDWVXNFBjPakfe/6hyRzb/JqMJwTJu8Nvavh1D3
5KDa44ZiBjn2l3xrKDqVvIWz3oj+jx6MK9GNLyaLhYyEzZqxIPEro80xx+ogG+jo+B1AfoB8gdX9
cwE2l3UTmDXijBCAJ2CMKxAVaiDzBlO/p4V+QTH7VyoaHkjGY8KRiYDIulIj94Fd1YbphbFV1FkO
PeYPXXGnc3YUa8oDXpnboDU3wra7B3whZULrcH+QmjyvwJQ8lfQG8Un0jVqxm08xXaVgbOxnJk10
C+CAkJx/35iSl52rcMQeaD/tL6VkE/eKaAK6MFaDIledlpx0jLK96oCHJ6G84FeyNgl3RC7mpWL9
EDtvtrIKRomgUHL1lIlbK/wVX8tmwSGcrVXnYf1dGsLcwwmnvenMlISGApB2IrabwTqrToUr022T
HdPxct53CxeksgHHD9RYykY/a5hhg4arSDzbUzoxeBZfDACMXkRilJpQT3YzpphFrB07gPCZsNX/
AyUOiIIYDzQs7zlxEM09e/bdbeMxULQy4wmLADysglCir3oYFQyEMeuj6voThn/W/5LSWDNtE8fv
LZGvXai+bb8ggc3Z5UmGc9LxfUKtPdHNVLSpL7lLqvKhvLl0+zzUWoCdrW26GnZzTh5+3FgHQIgW
Kewhd1NwfysviSH7cytiwyP5n8lYdBnb12NVqqrz5CoRzY9LElI8wtUjz2aT7OrKlDrrJEuvfhWL
Tqq1qxM1Vpa3qUHCni1mZ41wStbVrV7fsFWXhXApw12oi7d3iM7VJClWCs5W1pHK6SQ2Lr4/pK57
czsD2Az2nShDJ5kegIWhGGFufoZHwbOBy0Nnn2+1hseKsGzCehoyO/3t5iamQa7a9v61ATppo5+1
lunlBVaHbZ7QKJUhbr+ftiZX3OTQinLGLUwiQv57hv8ExWjoNWyMrxuJ2Ac51DxPKgPHNmBrdB8n
J5RjHQicTigVC5CgS/Kn5CsIOo0MPTH2cuo2z4NtwWn/wmFtEEVMKa1H4zxC4ognpTTGg4XktAZ6
0B5WTUYTbFXvNyo4FMvypppY/n6OWJZlYI7J9CcFNFofU2iQpebCtGR17mcJDvWiBHCC4uGHoowy
vQ19NqILm88aArKHHpKB/3kSVDDsaxrWjc/o6y2/7NBZtNXLjlk3UjNZIv64cvK/JQ4inkaifsjJ
FMZht3Cl8t5oRR7wQUfEnShbarj8Vm2HD8c3eey0hk0Sak7y21gW/F8yDaKFuVpcTE+ivtt0KT7S
5gxJspnh7S2qppJdURdfKCkB5dxqJCS8IW7+Ydr+mMNYTjfZD63JR7t6kUVMx4KKKDnNYfPP/Ifc
FQOtPq0Tlms/YgQQH/qyGk+t5XKnzzX7+dBnfd8Swq7ttDrFDUat2+XdhJaLX+Dbco1v7g1+bZn6
kmFVV1k+UA+DM5IyYH4TgGVhO8Wcd5YApmmPBQWQ4vPeGN+PpTOhqVt/le8Kh4wXsLs75cWnERcP
/GuZj4mBFzZfReG9EHNr3Gtxa4H8+Ls/agcDWqQpWhIo+GWyYMqAMM5h5Z6u1MajNpnKOxSQ8+6Z
YgsaEZaleSzutZW8A+8gg0kXPON60G9n8mQAb9lX9YVBX7T3AdoyM11ozt4YZISiUhRASBpyJlVI
9vj0bLt8YOCW4gUn0ktZtfKJp9sXMCwnape6ecBSkqGnrcV3g0XjvTcaAac4UFKBueguWgy7VA/6
vLnlccY4bHY+z7rVjYN/Iv/hYxNgSZsTl6QRzlIa/nqMGFPtGPGSt/0zHTu/16QoYJtpyVbPHm4o
flxrXWpX+a1KekzywszYJfaW6IQD3y48PFyIm3TFhP9jGk2mZDbCY/wzgnuHnfumDLVbPFQgyIFG
/jr2WsftkADx8/CdVd9z1k/xf5Oh0UXrKcvBQS6VcqQwKjnAOBCbLxKkxZpXqPE6nw2slugpbhe3
lrx0cE0XyOuvk2E1Ir0I/j28kb/gWPQax9fRa43XMntpUIXkBM739zSuQ0fQi5VUXtC6eOPMl8F5
Z+K8gMjKBJ7ebIzXa+3Qt724JoB06aSOxjzwlLF8JmM4RedN/h5cX4S8R/zn0iU3AFVGpETFSgxC
dNOmjxG7pkFHuVcYjrp/27Qc9lXvJ+fbwMVjCs3F6QOsNmrRJERaqWyeCK4yFM1cnHZavjoauCbn
0Msd2Efs1mgngivCe4glHN07IYnSVYrV9d5kuHUAcmTrDINLrNH4indAqd+meggmoFwLyWdFyLFm
umb/6hDCeND3+M5gj19IS8O1iee948onUn5U2wqLyRcVIiO9Hs5LjuGHlYXRI2iuHsn2GUAbEDvS
G7YsQu9LTbBVJNtxehEaMNU9BVgppczpfIyoKfnrrzBVyliROtboMNrvkrMqcgWDjxuKZO1qOpAL
8CzFQLeJ3+pAagbAWBkjTWcwhCRwi3LUMCKqSd5vbLStzOkGVaSDZV56e+T/Q17Z7e3Z0ADDMfNE
GFvZjBGvY9YYlxOZP/dD7U0NQQhp7NwIo7ZUaoHTFoLZfVEkl3otoftlWCnAlxq1QB7UB10ZB03U
GUyZJHGkJNY8JkhtfTvUvqLR1Em6XICravdReDKF/OoATgi14ozgKLwE5SnB8vvKmVyi/PIVUP3y
FlAzc6OIL5MFlJudUA6WR3INeqYeDm5H8UXE8P+NP7GRnipE9z/UlZUBf3OT+6nsnzu+638D3vu1
Ya+rl4DFKn3udrTn4qN+zrvS5ZjwKqKQs3vJ1Ku8jlDCCFF4+hIJE6V55P2nHf3qHHOPLMJJxfjR
wQ5emz58j5WHtDAdv1F7M64V2b8w0Nb4Zok0OFvU8YmxfMW+/dFxAg6FDspiAZQ3nrvG0koLRfvz
MIw0chR6PI7/blQ3KvsV9tJ3Bla4e1L/MNJm6GR4sIj7r73RXW2AxuC6+iswlg3pWOAuzOTkJuvu
rNiGjslvMvcqYQ0uVyhhTafbvlcuXVYtpfIlqf0KgiInlONk4YMO6njZAkLgeDGV5biNED740wq7
UU3falTOMKJdROdQ4xemQdoMf5x0ffFVbRog6Um1ohXiKhkDuLuusUgvHLjIp0FO/O3rrT/vxNZ4
114p2Xy2o4cb6Yklx8RmKGTywWNzR8dcLByJp84eIrf0jR9Ew18fVe/z7622d0krfKCqcHj/od53
yAdHbZZT+25khlMZKZx4F6+8GLfPvWW2wARPOmaLxNpHSwWHZK0fBf7gikHZEZ58sLhaWg6cFRYT
Ojwbfp8ELSAgE9AxRt5Q/sdzIN9ZhzfKS6enMCNKnQ5FAF7WjjmRtax/46SIzbqXO+slcMPf1BGZ
bOV1ITDmpWZ5Wi9Rc+UjB9Ngl8r2AEOJR53kwrfHePIqPkY1Po4uoOR670nbxBrZWPWtlSTnMp7I
3SmAQTzURihsyhFlA/BV53FAbVzCunGgvA4G2xe2qyy1vLmr0x87IW5wgkxKWSdDM/H1AYUs698J
wVFGdgWRbXNx+ZkiDea9y3Xerx0I2dT8pUy90Fqgpmd5DeYTNcv4dHUSRV4W2bK4uSkSEKs48NDL
1TQWgM43pevRxncs7Zco3ixkoiUgEwELBTg2k7VB4vF8PFkRWLOJUFnbzhOeAS7RLE6XtxM3TpVw
zqT3+e81fiSP9pwgFwypWteYaz/r4r69ydri1pwSPxzI0wdoMZ0CDjZZ/0kTT1JDH16h1IEoYy6Y
uVpgYVP1B2quEOdTb+FOf8LRswocY/NADlWfQIufPvNcDkz+CaFRfeOgKPoPXXmD1VuZpxBWtX6v
rkn/ZlTEcxHdYavkdK/p5PQaZhZg0CV4tI1ihGosePFBNwQpl2j8vm9NQa5OTSa6kMEqhq3W7ZIc
AXuHzBLw4S5aPQ+p4NiFuGA5ubFfMnmmyuVQaDJcS2yFVKR3cLyqfWYquO0BT1scEs8Cng6hr7zK
89ITN4RfLzK0Cd9kde9umUY13V1zPpr8WnPrpzx2qUCTMzniIg+dFQlt0LDuN8jF/UBPUpsvVYc6
CMdcSOFJhtnx5BY5/aJdWAQWMFIkgWhcqGjINaWYQ+egt4vMWhmIrriGLFGL6cmCGUwKurp6DjJc
nh+3o2hy6rKf5YRlWG2yQnhPFwqb+vFPWbwD2n0IZ4EbcCmmJaPVOBm3AZ9o+bPWPuDLZH513s/I
Dd1EB5reS2zR9ldVqEub01eQykyZ1w5GMfrbGjqy7ijJAc5RSbgZLSEMZABSJi7WSeKKpnx6fwUl
w286N089T/OGEenotT9ZTSJeguivY20nZxz+9kMsu6Azw2PUcIMpVg2DcIAJ+5YTff0ggyKTvKl6
d8kwm8YRn4vzgnC7Fxy56wL2dZMVuCpeCG7BaP9dONCqlyYL4G+NDNIt72xB4jmQ0Z8fnkUGzUHw
IckYAZSZ2UNhedkekODYbtyp97nMy7qQbrNurKBtcmKejLhLOv5qH4XiY+p0jvhiZQgcIdVoDW23
hdb/zRWuFg9t/PihKug79ZeMDcrD4uK15cR6ZKnTTzMul0v3WlwksCkcjiLfzKvRV0gmjuVy91vl
vMZfLocC1PHE7TVRE0cgGNlzk4FqRK0Ky4VYP2COwa4QOhgqNgqaas++YJT1A9lyAQmkXu7BmY1M
gp+gTpnEWUCb+YCFKoK/OvCUnQleyzVeKveumpdk2WxX+leF5oqLX7LFBKe1VZ4dxVXUwvG9G4t/
dL1QFOGOmFwia6Uu/tpx1xzhqKQZB5sk9AvXSlWh+eQpN6GKPviPyivPG928IMypj4a/x4Dh2ysp
iPTmMNjvn/asHRr+LA1mL0zCqqZ0ZlNxxTcQ09wZiugjBp7syPO9wU7IvNzrGHCzgF5fQOji2qew
yUxQ00h7UXS8w7H0OVaFL80DyCiYaIXSSrmPU0l03ytbUmm3VWLmTT0ZdsduOGCTRrJNy58E4mNr
Xj06IjC+AY0j/9ASUQL+jscL1/OQmiRFQbYVDKQQAmWdZRTLoOgqRFlq0cJXsUlT+hf7hMuQRsbj
Cu0PeV5uljYMrZJ2vCPIVx633SyKAlBeMapwGp/8+2jisnn8UB/TCbYqp3zUTstPysz87fAhyU4S
92XKqq9YpTMcTlw4f+qBgDfGBmtiJ0L+18N943wv5StmmxtMIdpHeyVyj+BmRbF0zLhG2YAXvFZq
oX92S/qkW/FQ6T15dRJMuQmUSqccLt9V62k7pcm9kD7c56Bf201mOaQVSVy7d2ui2fSCWIjS7tW8
LIJkjBQQM2Gsc3sTfJWrpgMUPHQpUOEn76jGsCV8OYdA9MxXLFBAcXsvstGmhhi6OMjSSeWxMQ3q
uBliumU9ZMtPe6YZ7LvVBDg4AS3qH7BHYTx40Knv90FERfTSvcCxejr18iNUOA6oKX3QdltrVT/f
2M2Z1YJD+HHqoJTOfK4BoRQokINR6vd65dVNuucKtUEU1AVbD5xiAMCYg3P0Sb5BkTwNdSesdbfD
wP286hsfHjegPYn1QiXUFw7VF0HQRi9b+NPIGyZ+73doAMmrCtjB74Qc/TV95dlXBAbaqy0zw+uC
q2cDEnOBHIcbjicbNGGpUn2alO1B72+AOHdsb7itpdkXI5dLWHzDkfohT25VxAtPcbg8eQD8Z0vD
2VZ6bV9cVec+Urp46yuMAY4UNdJ031+07u76cWDupiJwg70wza9D7WgoaSPSI35nUjiQQ1y5J8/p
ioAiBDZXwg3pr4igboZCXtUZa0RMUFBExGjS0ScOxA6SLqg0OVoaU14YkcXPgIbuLIPFtxvyCkL0
sUAU16Uz12qMQ2WA20EzHNz6rRO9+k8ZFo4sLxHNkMNOdSbnEXf2qXbPyClxM3VuCL8WgdENWpk9
qP3Op5jWsQ1+m0cl2kSPIe5lPb6tO3jWCA2TewSEpP1HHq19lQ+FjePWDne7IOTQ6Sap2GYdZJwz
ell+KOktgaprP6VW5OvrB/es4wTWVj6O43JHdy65DZ+2hIu6YUVBZNcBiCfcnas234Ui5a7LHESW
S5CLkiiJHa6znB74gGgH7htw/othGzqj4VgeABEF5plaoD5UuWULIlWDnzGQMKRexl/G1l8v6ey1
rP7IE4yFerL9gX3oOeixnVEH6sYjvyMFzjDl6rt8vq+TCbad45AF1Pv6D9vrb6kw6yb166uHLlTg
oZ8T+H7Lz5nKBChVdFJUUniKLkaoGlS6cN65TsXY+4IebZnenPqrWWGNlxz7DNFuCY75pgrIhrcE
o1HPsxK3tjAXr6UXG6Nfr8fNMA9yUngr961aVBxx2QLjK8NKHcxcrnMDSDFNxIhmYcKGIc6D4Fnf
hMW/u8YalT9dZyItk0G8u3fgdj36wRHcE8Sd7U4d2fD98ZLvy4QedKkUKS5PhAn5g5zGMIduHMsF
+DEigL59tZuwOS4TqRh4YJRCHXuP2QVUncMr6lu4E4ZnxgpRM/Msdl1tZaymbruks3FjGF+jRXku
+kQ7RobC3B8U+tKOUO0dBLbRiea7sJNJijXCVHbyE0cKEHHXJ/Dih0DAYIy4+iZjFlHeI0dJ8kC3
WOKXOCeE+IBHHJV5k2qDoYjjoCoKiOr+W2DrvPoHoYH+mscpF7H7uyvFQ5IfVC3UvuTkPPDReNV9
fjSKws46t3U/NvAfPKaaDxPUVQ52CeNVewJy7pM9jwneaaLTji2DDd709SlsNozDEqWzotKH6yba
JkCjGSFpfXO4/26rpFRSXZ3iHxsFwrOCm0RAqx8wWKs6GpqFvPT/IEn69kUyo8DJHbRic9IOrdCG
1anruHLZgdyHYGEbd/ByyjxQ5ZeSCTRI7hoE/fkT74g9hScJiOYI6l68LVmFUKrYU9alkHsAQwGh
oUVjS3LUfoooLnQwa9ckq+fUmsHboZDLG2RRv7OoJJv4e5ZRREpCsU25fRx78XLjEPmF+U57r+04
79U2cmMiZ+sj8kyjfZvuhs7BMkFHp3YrfrWd6r4iakoTcFaDNTEmZpObvjRspbxj5dDuQzkIaHVy
sF6lA/GBDxVWFU8TxpjRLHKu5D1QHyii6GTetqzfOXNfqJjzVmAcUd4JeFlqVxmOCeVrZvjYb2Ur
/PwHzlq3MYD06chJLFqUKA0UU80hEv4BqRnx4e30FBCm+IF/fis9ogMiAjQVrDF/SA2LAHl2jWft
gDjCGUihqdQ2LGvwpAIp49r06i8Gy+AoEJa6kz8v77e2xaLOuv76mCV6+XykIKW842nmbXCAasX9
RZpwhEQIzFd7w/1KT8SGmDOlQNJK4R1dCb2UUiwdz9hKwD1sSUxBwWHWsQe7k9f5NajHPztiRiPA
X6RzHfWpzISuCBjXFkRGDomgSnp1tt4sdMm/koAFFRrhJWX7UaonevzfcjFiNOyTohIxezJp2uJB
Pd5RefscDGkQW0j1bo9Q9LHADo5jTt7Uek5PLVJIrJzn2m7tIgpgqGugC3UHnb0FmRlxJaYrrgok
8fCR2KxiJ7u7zpIpAoaRvWjBsjbV4fGUH2xBIyxeNq01wEVkVhIZ4MaeEiu6RkcGA64wFoomQ7RK
4sg647psDOs+POf92vxnVKRUz9iXhSPS50WEqPrabsyIGMFxtBFvXpGZfdooixvn88qEh672D4aS
vCvBxyjoGHZXuKMrnU5JS/IDp5AN5kWFJOz7yeJlP3hRM/kaBKj/wYWHx8vULKxaCKz0SkRmsOk3
EdNx8CPYpz6ApNq5gjkQaYVqq6Udz3NYwdL7pnH4y4xDHyvAu7addQPXPMoyn3wrfo3TQCKNFFQ1
f5qkN0HiZBFL4hXrrBcgSPOCRgBSigf+m+4vvFiOGiOHXQdo2x9s8Pv5zVeRtC6YjOW8BXuUKn9f
tjoIhVOpiXwCqfTkiO9Ml3iqay/PgNEJ/3QkhVuMXqNb6bvX/arFWOJFarfsd/9QoQzewmVEt+RS
pvuhYvXn/mus4e/u8zlsla1sRYt265T3STnw1/wSPVVHHNqqiZ7rFjLCvOnSZhQMqh7ZE8R+Js9j
pHdaMnkfKu6cf35hUg3u/q2hI8LG7cw7PgJLTw9xfxuKGCrrKrSbJnLhmlKQp5cWnTdVfX3rVr9p
mFJtJ0pEmZrPICxZ/Ju0fIKF/nQju+u8JLmL1+nAyIkmqHH6F+aK9jMJm/MwwjIZ4i1QiMfheAlc
fhzFHh1SEsZeupeFT5D0mQiOND/AHrhzqN8xzPkYJerTM/rPJHlOFWthSqLjTKJ2d/b86FZZ/Aj3
Aa5YKO38wZCK2PTseeyQxV0Uj6p275aQm9BbJMHEnX7wDmKshoMF1KOD8YER88vBoTViE/l0hBnD
JZTQvgAircUKNtmiVikN+tvKL3g+xPCHHk39hiCqzllFYrclP52c+l9e5fX76+vwtRRROceKbiuD
6D7ped3jZId7w6FHkYJ5T3TqUf9kHUHC91GWAriLmw83565AaoLYQciMT4MuvD3dbJJO5sbB8l0R
8lHQ1bLE9V8WU0yx2gpE5xYS4tWZ4853FUkbygjFyI/CnVskr2LCWRQkDCXNQULJKSIuiKlyVRKd
iS+cKuoNNI9scWyeaZno5K+uN7pwltvLc80kunDXVMQhOsaZnnysns6TikuOp9Q08bBuz3xW2b+k
+Tqixu7y4gDt9D788qb76J8P5Y9gMlwXEnOm+c9LsHN8AzPrZq66D4sep0CeBjDNPpzo/4Bbn2mV
m4Q2cfjBRjYoYJb8xfLppThQpK8UD+zDh+TvD6XilZIYyclsK+lcoPY0qjkKJbc27re/UZhR4n9A
Vcfi6jjUNGRcvMTMUR8a/Xngd1Q4UpDMwqn/02bKo/+ioSKeJeYva06i2zKh7LbObQPr653QaWpR
V6RlGIWddu16vY9+D/GJN9dTqTc0nEOgF/dsX73MdEKdJFNxZCgAv6JUL9YFrywreOdha1HB1UXw
t8sdrqhoZZyx/4xvI6t0RWcd179diukKhRA7quTwAohS8ZcOx2mV2y3PGhJ4ax7FYZ5lk94dayXg
2xD2dS3xKz/IZ//gM9nYofKE99twF9XVvjWelG+gWG8qrJHiOchJZUJ9zlCnnoOzaSIgu8gevIbe
EoMN9ySmRTQ2OUdNmzSl1waayqkVOe52tieaEGUydFs0uk+i+vBu+4zidZtrfUuEHWIjqJiPJITr
tp0d27eIJ6/n9kJWrQ2j9OUtwniktefqOGD2lft1v9Z3hXITbi4D98m1w857zV7bv3Dz3OYTxLqM
6dQwUtIODDiCNSpPeIFV1yrz+roiu4yqGXXSCsb9lpQ8ufTZlzkQ+StaR4fe889WgPtCAZzdpfQ/
R9U62Jkr57NChPTKmQnt4G6Umqd49xDVdljlJM2KC72DxWA3F7wXRZYOSXX88ofbU8gM0zPlhI8J
RXVaJAQ8EiTjR1SZiQQEcLdA709l1Xgk/P4uxzj3tHIZYflXABTA/IehN2aAmi3mJxuVxuXEViq/
a2CE+7R1GLW13s0P6EK1BlvyjZ6hpLt7xk2Jm1wQE+hlwUXlFakqUQRol911sBQARDX7y/+RSTGS
Ix2m0KK4HW1w3z3wjIst8RvIoij3TNgb9QS24dzzx8IOH5VgIrFll6z4a2f9AR0hJukZoaubc7PT
3f7YJ0ILMb2mkqEefxecPew452D1G1QWrg3sN0VWX12lCkbQ4t0enoExVaez4DVXB7gFQZwlzBih
2Rnc+p7IstNH18isMv5wyAzodipakLPWOxa4NqA/X7pXxd8jxB1KvfCMyV2s0qfAvOz/7uN0tKuS
3Xr6nENNcviaRs2UCk1etvw5NLzZGqp8edKw2WpLS9k4Z6rOEtH23IOYwIO1wHzqSB+MJ21zEZRN
JqoGK3/WJK//+zGAWRbM8hWRPVrMUBUREyvU3d2k0Viq2JbMQxkUzdQ69g3KtY9Y7C9oQUjVyLxh
8qXRnVBlK1e3aU6pcw9jaecWAf5sTk3hDS3qGd6WPPoy1p6GO8HglpKnmOAL8NX3EdRVD6QLf7ca
Pl1nAR4AHv+W+qEllV7aa4jwbje7MoWO7ovY0+uQF+xo9nZv0N7hILwQMD57ccfUgGEUqhIhwzox
5xLTfzLAjgtcgyh/eouLBOQHS1E/suPMdjo/aX0oO5DHo4WkuJbCNUrmxgcGKbtB574BAKhvdc/L
ucpIjmflopKnhXMlbXTULMSqPzrHbywG+XMYoH1bP7NKjDhOly7JM0DvXwkDfWC5ce9Y2AnQk9+2
V56k2JI9b7wsAY3waCAJcvCIPZYar0mPCxdT+8UH2A3Auup+3KUzFlwV0QcZJW80qSv1wOTUuewn
Tz1UzlCCNtCuPy3l0SmU2D0KEjNNTKvWONvT/6OcTI3ytOS6bdBvLBT+Jq/NlW3bRRq615S2Epol
YYYh6n0vLgQ9+MDSh4TsjXkOyPb3wG1WoEQwpxIcMo3qRMT99q/gfV5xYMK2BAXkCcM8+YofNkmW
qSQAWOkCJfLKZVr59DzM7Nv6LI2oktRY9lU8lFXwqgQQqi1MxOZ7+xm/rnNCmMwgHbgkn4Ttc4HX
WJp5ghWsGa1lxKlmjVG25TqgBOlMWlIIig93D8yl5NJ0AlY84fS1xcPTMOAJAmnqKwbmFxz1SJd6
teYh0VO/lyfhUYLCQiv3JKuLQXIn7QB2xUSreByXMjmbUHY2CecLaQS+YxLF9Mhch9Ldqg3EGgyk
vnZ0vKv0cA2B3LZWOgM0oYnou1jFZCtoooOHq4soTDV3Qqj9Fh7ClneupyN7AjgqrdNqPrRWsAKd
9th1o5L3DMpPDS+8JKqHTDq6xZawj/ioC9frHIzv9rgOZ2envGePdkSiLk4GbbsKB8paCkV41txS
7BGc/LpmUdADg+HyrOh/tffv6PxUz+CGbiVhxX6RdyLEsoM5KZa6JtEWj1DAKMKQIoMvuGI6awnm
lyOGvkryWP+nu6pO/2sBVh+gMlpCJBuyrwCB611f9WcKrZx5OUk/ttF7Vx5feQ0vyTjzdd9IDGdx
pnY+7Obk5cq4QAvarwgc8Xg1pEar5C03gzMpw+hQYdBWggSRzwFnaD+ifcdrZkdTK1lWIFfu08WA
Lw6jMcs1fT1B4knWseKW7fr2olSeOzesuohsnBrdcH558M5Mxn25JguUAEZX+AzIWuj8Yo4zgR9D
OlqzHDm6V+O/vXc7MfObPQXeuxDy8ei9j7JTyqg0ap4um+GTz4Yij9JKHMaUXfNMQlh4+sLf82sZ
Flonlbny4nj0q0QLrRQg4mqxA77HJI2MqzXWcAVHS6KxVluaVpk9h4iOAfLbbZvmVRZBzH9TPT5T
KTUvGY29AICf324SVdBdyGk4wuQvvKP/ZCYRB0NfzIbB4X9RNQHZ3SsVFeNT/Xr4VtrEHIsAA84h
jUu4E6sehRPEhjwGepAaVdLbpjUWbCFY0OH7aaoKuzJrd6wmJKSsJxRv7OtY+48zCWy5tRQzOBAX
fehQpdubiBLrz6yq0ISGGVgfYl2Qt1eOJy3HjjMIuZPWEMZeoPtiex78N2ZZw90xF+e3hh5ELYcO
4/S2yfINkO5E8Pw3AnrBll9U5BXLLglmyeMm3HaN5iXSATgUUCcpXhL8D9vCHqBsqNPcoveTxyob
VfOYf+u+R0Hlef8iydCA+0SK9Sebf/k7DGspETnXA5dZCXTma2AT7YOGhaaYMVM7fgehlkWTIRQe
o2zwn5+ZTN1baVuc5JpuKpAtCSyY6PLvNCa4Oiwp0e0GHt3QIqZeAU7Odds5glNv7gK10+VZ5XD+
aPDJi5zWG4U370SUKxl1c5slychuAmq7+NR/O+SburdUi3TAersM49JV6r2KmRcJHqM/f2YZ9OLa
U3kHZOcVgLjus/KlrhoBrGQkjNfdt5uUzSJzLK2zVtPFj8+68TUsF1lTF+2Legw2HDBxGw8TtVKo
h2d+8DMQPUgy7nd3v0t7dZNc2yh+kFrxBEX/FXtTh8qyG9uqA5GTjivM2aQhscrSNzcdig44cOCg
Eu93+8+BEP9LUqkV9SenIpTEund6ykR4rRr/tAOAoO/TI702D28WXRTRWEENDK5/mIn/cl57e9PX
y9mFJewF4DTOpU1D7ZgDEATNO3hpc3ca7Q/K41oUo5HL/gf72qrTSdGSCA+Z/qCwXHX+3OuynXKO
bUN8LS3Bsj2MrkI9DtjwjLvTixqB3mjPGdJcVINHRao6viHpteXU6d86FnwAFUxeDszNUjrJnDJc
/WAiFYfy68K4nOZw3DHH5J9r0+0TyzLBnYnvpG7gKUlKwA/1g3d0hnJTIKs5Qvaes4m1m/07vAse
CrIyrgtcX1D5jYgmp4B5JaKtCe3kOADTE7Q6iy1HWT9TAc9zZVdYol4qdQ/nzQY7fxzlDhRMe+nk
p6MllLXUhloQ8h/ka9tqbw2eknsD9bqyMINl8Mztm/gZk+n8ZULcj4H1M1YPLREYIfGn5scO25SN
RIUitQSNgMLJukSw6jwkq3f8UyIkwTD4FcF8itcLGTw9qaZZtkJg2rYHzGHzbU6YtNYP3K469j6J
JpOKYU0iLoDnZsgWj25VZJYq5h1xb21mTweb70XnKuIemtUGNBGiMDROuVxPDN9+z3dq7xq1fiTQ
WE4DGND+cv5s7v2geqfnAG9RwSdUEukA3UDswE1SIZ7MGbTb2kEb99wu/shWrfaWHwNpQx13utYC
mvI/VsUXLPrrrtZMNtZoDATfKyUZZF34jHXcsivktzPwLbCERSoiVUWKz1FfYEGdyYWEE6Ju1Ijx
pXvDYoe7YNCpn1HVJoi/gAealnaegj+kyW1QHbidOuLqo9LwM//mxjdE8pqRzkRIiHY0ZaamHaY8
q83+VypsBpSpxjc1wvID6Wd6gofw0GrROcc4Qk+3mHXy4iQxz9SC+a2wSNpR6lGYQ267dEezd4qu
cj1xno03C225uwS6Novs5AsAjIh9yXXSBhV+qMiKNauiw6T1T6Zkp/OALThVsgTLzXD4EqH2Vccq
ZDfsQHvB8+zrfV2FY6guDBuBuZYeF0gELIGFkH6qHOAu51WFWN49tKfCoVqaDNjvUtjUWtP2C18+
tionO9ZwBK6dUSMhWcsdlLkPaWZHZ6LGuhKn99vGYEJHMCqy1ortdGaZPjfOvHvHg2UPUAHvWgPw
LsVAKLf/PL6vaBt0RPQhCcF3kwup1b4U6lq5glO3jJOoaFngo7tszT/FbLJACAp1MjZHc4d+x8oG
yRN7rJjBuJmqGit8yLKlih3zlRNVgPsB0pfYybTl98FRujdYhJkTzK4zQJF06r5/uQJM8ee3Pd3/
KUpFqjydf4+huRoDTS+67smtOQUXvBifkqRhc2pejrWqhObsXhjFptJZlH4m4HRwQyRei1xEaUHK
wOXkNmpTiwlbjsWviHFcp9s4hOdktuAy9o7CWemYFuUIrQ/q+zhvVV/DQ61BOXuRYzxGn//NjAHP
TdQkdqbVch5JbRgvmCTcpMVWowbEk8urzIjPTPWu+1KcEEUkxaMbOGkjp6TqQtz6vCw1e9fUQ0hA
ciOe1iyHGpOwa59RyWvS/Uddx3wRK242jXi1JIQBBnZkQycef8NIDkcJY2XvXetH3kBuL1ni6pv6
/HcZcCV1MGwxY/fHZs9sEzyunZEQ3SY8NZkveuGNL4hSrx4lt8oV+/GTXPAtnwzRPEl45pmtEui8
9GppyTYPYK+h9KpH6/yMkFhYN2OE8/0osWZy7uunzdyzvNCo7v2YvZLGx3D/mzxoBqHIt14HfdXS
l51z8RkQUoJ2b+NbEl7lEydyr7gYp5+LGDyTPoWZsTdxjv8dv+u+X4EWmu681jAdO8SEFZjgvkRY
blvTTiWPezP8QxjkgiJzAhV7bNmw8sIMBRai62ppQD3soV6A9oRhKF1Sd0jMLy6hYPP2VvMhPDVe
Wt0JNYLlpitGW1x9aUevgvWHMKldP9mhgwtIPAaEkI1gj3chsy4AepsIO9Z90Qg3b/Ta2JBoGk/f
ZQOlvk6mfk5TZWoftDVmiLsRW9L4ba3UymKv4ZPNfMG17dCHkNCHKlO6cH/fTB1wLul0bggYGdC6
IR2XG2JxRhp6f6X1i6V/DpPb/GUnRzNYui54vcsBpDgIZ/NbGBsVFugeqP5inBpfSddEh1Fwbj+X
0dB9+91/ddFz12BqIchLrAohUETkqkzJA7z+/cCN40TYEqT/A0oi5DUBgfS02XHI1e5wi+CIhR7V
HqBWepcTDf73COYwIzrkxmHsXplLbhZK2LHGiM6y/NT+qWjTgROc/Il0w7H8rmE8JqT4Nag92i2L
wT7dNbXaMLBswyRTXkg7cllO0YeNLyYqJZeoiDzvxZYM5sMA5Fb39vyFsUXkLxIGb60C43f0/xgr
ReLXnZQw0ZvZYsfmUEbSW0iUPxXuZf8I7OYo+kgG9WTZf7HGRiwh7h+JcxGQ2GpS95Ie6obq24Pw
XT5XOVH+EMAUv84RHCAGuU4NioF9FwWNllsUFy1QhWIM+DH6uDrhqk20paRBAloPjtVn2TwZuC67
5tBRWqjBrVMMuyqFgdaYUk5pOU5fxD7RGfNMFW5gTv2OUG3gtzJ5lIcmXis+A3gCynf2SuJ74+8s
KFHvaMkVBl5ul+7gZLlOiqj69VNlqP4oCiZRfJfe3Y6KsUScu9OvXfcxOrMRt6CVMF/DViUu8PV2
H/G6DaWpaFNuZ0FDHRj7zhae/z1WGRkn5EYr16E1T0Hvfgq9NL3wjCpqacOFPAPlRj1Vz6B4zCuz
j63vGwu+UxWggP+R7lc77ynZ1N6cHTZ86DuIyoooipTCLb5D2+1yeoQKOj8h5vctBsjE48nxUQFx
/4eO4hQXb7xK8xZswhxMjA79qvk0ylj1cult7TiwyV8POj5qbwcbLYRFpk5DNDpKmtYcPHb5vxAZ
LbUAyZfiQOy2gelHD3m/W/W2J6EdzO12IkqDOK4OoDWzpwqFE/Rlxs0vmWsf/Ql8p5jB/+CA3ra7
plzb0+VNR2av2KDVIIWtP4Ed2d/blu/trgcxbTp4YIzvcq6ZAlccnxOJ4UsGQ18booq0frG3aC/I
49uHQkGhibpjQwYfK5uTJXE1HRLP6zX4uBz4cQBK0FegsHo+tdSUb8nA1SxRmn5ESB4IqobDqSyY
nn1ccFbyCSrm6cSmL/vJoB0CB+k/Z8/ju/g5F636zFnQnU8z31EfdidAKAKTqhAe5402pKAYuJVb
aRwOKDk34yYoBrO2nKd72/6r2JRvkpKFTFGEZBjfeUuDjraFpRP2hGzYr56ppK0i/xcV3Nt7Ha4s
lyCHrYcqqi74FG1Yz6jy+QSnPnKzICpJGLX81TVc//7bZM098eda7Ispre77LHcMBWuixVjrK6du
MsO0dULwjW+AM8eItoEdCjquoRaa0OIk7VNYN9uuAbD9rpgDSjXY/uijo5RQhf4tJbzpftKTgLBd
VloA/D/wmsjVXA8I6TIL4jdc4EOCqCH+6g4LDrfMX/3N2iulkuBqzMvH4YDgeG8mEr5yCVx+Nt6i
VGcKxbottdDfpXW4dmWB3pR1YHmUO8wbZY7ruN4wkyLKAvKZNh2H+ElHAD7XqmRsS/rGYw4ZlJlN
aUgwOULLKGkWLO8DYCRshMJrVYP9H1NqYkWrx8g4V9Xbga7thlssZzTB923MTqMKoZVGipcTb6VS
+P6T3Mcs+7qF2T/uRdpbdyOcRXASltSh0pIghK68wXk5niH3J7ld4WaKa3Jodge/1ktlW94t35XI
YCBmxth7XawrU31xWuoXHkbY6BjR4iYg4986JA22a+N00LQMXHpzCja5xHMovSi1c79g9pPKtL0q
v0SvwSwsSS3yBUxxisoNQ0jEO4s/pciXNRr8AkZRfuIafbwrwH6B6W99MePwIegEoDn4/M+0D9Lj
xBKLeEst/bUF+utzFOZCDFM3BPrceMn9dwf73P/rQRxMKSBuk+8TRcni1pI55QnRdT1oWgfJRoCT
svZ9t5tO+conxB0lrFSnXYO5OIIjKemBqFxRE2YFrk+0l+YZhPMOcrhfVHMZgjLA0f79lQoWv/sM
FlOGbKaesRgf++EmYF2+wEocd2NMGqhT7BJmV5YXwoNPHsAuCT6DFLsQI63wnsCLimCKi6NahC9E
0i3BWULtGk6nRZCur4HuSKRZ1trjW86DumOnzIFblHLefKFWHk25rRONzEaoU7bnVJAeYSaMoQ8b
SpVt0yfQKzZHU3NuWYUIbzTI2KdBjIhGx+GtQlf/cPOYRNotoVSvf4sJBGckLaSkvj+SJrVEiifs
yToCYSWISMb4AP7QIucQN4kozO4svJks1QxgvzPndvZZkzQPYb9QSNPwAaAm+NqYXC7EQu93Vp1W
aGXo7QfMuVVcfm+1v80JXDXDleysjoIRQizXZQcZmCDyXrZVaLA6oMEAOEYwQ81eJmDRtKhIklLS
0fVo+PqlhMGm1uYPXmJUMANyZyC/FAaSm+1gbP9XWcvr/ekY8dWA5QRl+0VD8aXCtjDbtqy730PJ
dRj9RpDsgT+PVH9KH4sVaamgaQgKsIBiIRw+nmWdwcKhNRJhtUASx50FveDT1buOPcpUbZHVjeMs
GwAldAK9J0otNCChuTSQNupaA7HzZjlA71kR9+23h/R3QU0rIempR25Zmoea2PBQRa1kr62kCkNP
rd1yzR3ck3/5fEB1Ir8Z2aEbRhbXvXAAZ57H8QEHyN0sX2cNmQQ4TzAFSNWdC9vPw8a45mzO7jNR
iV7L9cWtRyM0gJMYutZhxiJL0MweVTgObVfD88laP1zrhZPogf1c2UVki1sZHhEOorHACm9qctg/
1cJrv4k6TAAJFEZSWZTXPqm4A8PY6ypkFD3w3Bjx8VbpX7S4Hr8o9Fk1D2Fuqb8AI+ycAfAlyVcs
1VqxYLO2ilzqCcCZW9B7vgF+WWf+YAxWOGeaciImmB6/yryAUGFCK1Y54Gt8LtaUpiUiDZ+vyrIF
eO3kXMEsRg0jUI/a3hsNtbahDGQLKpclzY9QWRlHVb9CctvYX3H0CeFVl0ZJ8dffm41EXaubhcCY
nDnBzN+pZGBffOx2Y9DT6daEloFpFO1Cb6lCzAd1qfUVQvX5ljpJPn6Uklksikc05C5Nc0rhUT6f
x/YAnT4THpO/L3WjdCO9p0kw5HHwFTBkkl8y21pZtZhZz3gOb4w/8lsDRPQ2ePaHdbR00j8Qmpeg
cXh3E0895BGL8Y9qggE/W6QX4whd5E7EShzyvPIY4tPzaufa5UxZb/pAxcxMw31r5nYgsNI/siqk
tiHIigFIVFkg6W1lxG2GZ6WLYH4zhBqF2uMT98u3tQI5BqytaG7EWJvVsPekzsGcIbt7jREa+Kwf
npWutfHE9G1VpC8mgr0K7DBy56zZfaoV9JT0kt2Qi0XkTE59YO+Cph9+B6iSdmW70Yu0eX1bUSKR
UuFS6aN605+/OrGBNXTBxlEAbnmAj712TOajXwZmVf7DEMwmf/kS7R0raAu3zMhloYydjwbXsyj9
Zru8/vwHNQBwYthFNYHCWGlppCOE6bjqHZARIx0S7b8GTjQSvqoI1nswfmY47N/weh6kVYwbqWI3
Z6UQkGVCkJyrYZg/UM8DXK3J2Uvf80pOdYr9YItoD9EsmePlvewI5WRHzRFhmINp7mLaW+QrE7qu
I+5kwlxSSbp40/U7ycATonlKUww3W8WT9S2FBXqHCsQwXaojDtuyz5aXT+5UrBdBvrJZTOVy80K2
7MwmO0OtSRfCCft8ANM+MiM660jXvuTzg9/OV8wpHF9VVnMd5YF6h7RlPiJiwc+PVd8OMihseG9q
Wu5QzCXCLbo9R/8SyI9/OtepEbvd6KclW1QErh3lV+oTF58N+gY/CyCKdUWEDQ2Eg2f+7ENnJyRn
BDcHN6khKwR1NLujS3IZU9DWdx/teaz926jEataVlSvePQppBiN9rn7umHMW7keD8Mmzsnj3b3Z6
jrdfObUbMYuJT4Aq2F8qutJIK3PW0vQoWVPH56awyVQci/Ydn+h97jeblWQe1SKSi5Fp+73bg71T
Mo4hBruOOOufFtYDbbP4SyHTR0YSoGMbz9MhU/Zqn7JkfG6T7CHte/AHYqlnBkN6J0ceHhIH78To
zdnRLuMKmdzdyiZOJNSCkfLKh3ertwFxhTUz4f9GSCJi7kvDk+S/65cffTucX8EbA4GQ3aXykKaJ
KsR3wKxH2K1EB5t5JXiSs8DVUqXLqDdZChb5J35Pyfn9iVHwOqpxPnjsIfG3C2F0IDNEG7rviU0p
sn6Wfg+D+24WSJ0r+bV59aZjZQW20DUX71U4RT0AlJ0JRZxxLTSFfxIrNvyACKwNvabAdHvSY12g
7amgxjyuvmesmmCaJ/XFbomlShSrwqMQE6tmxaDHdVPCXu6ZXYJ0qaTShthXOp4quh/M+VPx1Z5H
eh2BtwX0iT2t0FURlJVEOYsaSMFHQ/Qhw6uL+QnKoyV25tKpTnKXjOIuEjCmn88m532T1jcuoN6Q
zhhRwBWF1DrIn5IMZNBMRVMBJoE0TgxJq848GoFQIgli6IeyYCkh0HUIIq4wIJOOpvfmVtogqDQG
1aWeOzhgL3lZgq9cSztux5xhVZ9iDFgx4tgibH6s7MXo3zqPc4priOv/QblD8igIeIRam1pVg8Vv
jUTcAidR2tkXK9VgBGV3/u025tm4eCNfha9aVALtpjlekhO2mNEKlY1yJ/nHXHxXLTbJWWAyUsV8
CeRWBIywvnpsHu20Es0KN8p7C3XOH0YIODyasHy7EmOmzyrUwIf5SiauKlA6msePz4wJqWSaNta2
TSqJgkqArzw4jXn8vq6SWE8Ea14Gh38JZq6+XUSsyr5XgPd+cX+JT9acbyyf2K6s6EACXa2U5Wkr
cMUVWdW60tAvpoMUIZ5dqHdoRvf7GyFD2mQSekjONujHDx7yi8B9x8rBGK9UR5Nq7+kX8HS5Q4pv
gTRi2YX8kX0Qtec0sFjsDXRJxdH47+Gh9wndTVKD0GNxwsXHS9qwPlyEtqVKIWWxqJUFLLzXIln4
x4adLKc69pK1NNkoH/BQdhnWZ1nyv0ZnK0+i56+pBOzm
`protect end_protected
