-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
KRTErBJCD/LTcO4N+5x00VmWmaBWCF+eqiDAR9khBPbAuN3KL4HWBiOF54wKQU4lt0XIxGQ28pQ+
AxhAe5zGquekEZlWB75GY2Jizv4VmE/H0qsz8nWrO9cAOizOV+WsZ8jBaLySmy4cZiXb8hUaBYmX
vs0Vu1d7zcUcZZf8wkR5OATnXSfVMH42poX6Sa1E2Ss/oCCBwFNA8hNKHlH0uXOIvizt4Oih3OvN
bYP7B1vKNtHzph7ENQiar6moya/yCC5sYFoqATW/5gPRLeeqWn9ekjeSnsiZctG5ND2eJAL1TnWI
aMKhX+9XZFrG6aN4zB6EkM3jqmj7mKwwADayHw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 8848)
`protect data_block
/eVD33TafeUA1/YNAYNHVp9kEOwuucHwA+PoHFO5LhyHNPSYAS49RewW/ms5+Ig/rkdTyEUd9zZ/
gCtlcPKNaE+dufJe2O7w69epGuGSihDOb3OtdoCk53EaS3asrMGpr62isbj+OQYq9hoECPOJJ9IS
/jD3RlwnRLIwITeKczlCMc9K9nyeCxwrZnzma+5AL7vQmNZ137Y0el1FOSNPbqG2BRgerRIgMAkt
+0+5LYNBOgd+lAj2SmWncDetxNCJweYT6WqEMRUmn3UOq3PMLZ0KNXMLrSmjict7zN3SIyHS7fdq
3r5/yf5xpVr8P2n9yRjFJvjV6SqFnxiFXnDDLJaC2htFExKno2n6gKMQ/EcKDiDGia9IgbnbQhcp
rCCquoF+mkSSoFpRG6eeklXQNElYBKghKKbDUxG3e+Mv8TCMKFeYdKuuUC5NSestHTEXAw+nZULg
7gYS0nZHh3V5UC7HQzrFTlP/vPmwbXFcqHO3E+bdQhhko+wj8xtsuANfgBMIvuPnVHgInwxgWKkK
s6usUKDw1ktreMdD7oTuaT6PwNKjYwxoHfBtbqDbYreY6L5CzIFV/AMeKeHvqqa5gRYPNuSNu5Xo
USo2+2Ubw6/9dFMvEuYj1h3kzQLpstxt3QLInyHP0gXlawO1BgzKbTjZ0yUL+yQyatAeL1OOwTP8
JzFkA7iGEjP0HjWl6evcg3Gmt7OQ1oOnSN6pA+qHjzo4roAbiliQNhiv72gU5MN46M0IQZK+CAk4
3QIV4N2PvzzoPH4uAiHR2jb39E779p4Mc7exwAe5ewz3pKvbFv5hNscqVMZeYfEzTcq3wGeT/dVB
c1BN1xmz6EO/KvnxmtJV8G5cemp9PvHD6Vaxqg82+YK2Lvr1kWGfp3k6t3iWijPhOGRBCoEpg28B
v+ZiZ0ZduoJWAa0dnFLOSR45arZppTxnZqAHigk9gcPiilJWLZfCAvDNS/4sP1AAETGW0nCUHOZT
A0N3tMpsAzUrHSP0bnoO/a/hP4WreCDuucLuZQtFzrdPOi5m3wVkitXLX3/A+5EFrcnxblsKos9P
Fmln/Vt66vOiYP5zBE/DlVkXaPIHF9g46iNrbRDMSRwtfpwtnmuiNKv+bs1YFZXW8ceRWP0+6z5p
0ZtQ1Sp46UBHRKzJ1E3be+xf9/nGr74lnFMcrbmrFKR/NHZNAyrUY3x7ibzZE9x0JCsbKQ+urT+t
uCAL1j7/ZX/AgLSqydIgWSunqN6WGghihVo7Z/UN2xBxuL51t4Ek8sRnFcRp7dSGeEJ/hLIhTUUb
/8nx5DoVxOW+bTzMgDwGLzcBetNU3Nu3Gd8nbYwPbXZNKMBWs8tVZxRJffxzaKD4lXHcsME1xF9i
Yc6ehb9WmroMCS/vYebBlRWrgo83mtp35MFhTW0ci7Uj7N7DGqqUPtC6Eox/MHDf5ekw13mdqD3E
1WKJRxaj9W5wUDmrmh6SuGEq0xVMNqapybaFK75+8qJ7qafoL2Td+Z5lYcK2I8Nl+p8bk5gsSKxA
DZbb7OdpEcw5/AWWWaDrbZT51jaMQwTLttMPgPKbt1leInu3FYOawAWKgu3v+eIUcK/hi42Rpkja
KjEiDXokYvK4li61os10fGkRs+XO/8FUzqoRefq1hniK2ILnHRhVbtl1jc8cGJQ5KDI2Pc5ArqzF
au8tvfA3B1Y8GL0ekbR882GZ3t2d9KZV0338ew4ZZ3itacvw9sysOg/uhF/xy8sdZFgguZZEIYA8
vzLikp0kPRu+LOpkJ97raDmRrWW8hGpynzNS9UBK8LRYkAXWLbERRr/BMvW6IYdCnDV4SxqZ8lbp
52SSL+blYPSczBbggKoSTciePR6TvquIkGRk/2xmJY7Y1nBhDjC4ozAnkmz9wSmdKmyTsJ61P+cp
3dCIiU3UVqRuJ5748ZqdXjPaZgPoHTz+hLqcMCCx9bIOouac5oN+LdjEelxPpxFVpJd/1GsP3kMQ
E1M/ls3vr4AoOh6t22/YJZkh35x/SVJiNBJbBrOeYQYQA/SBUOq3f1sMAfe1J1dp1xfbFJxZ85PJ
kPVPKaDMOnrj+0tSrz3Y9ki73pRW1uVi4yhOwNKDMKNjg1vis8uT1czcISBMolo21syl0ShV9EYx
ncSqtDlPgC3VQaA/dyabwEyRqB5Acvz/8kU6zasCnQHrxuP8hua12MfMTSEyyg6YQioLdtbVxm8z
do5uSwLyybOqFqn+FSIXcUxAgsJL/RCu9g9BgckcFSsXGHVmgRbuijUhJK6M7/tRhsUF1DB84suG
t1BnKe/6sODGdxRmtoqe20qq+XSqRAxscfnmFS7FYY77DfqGZbk1fQ31iKbeX55jBReClHrmrZ9x
ef7/7cmntCz2+xha9T3VCXQsDu72D03qm072Iy67jGyxYwJjziczVTv480LE0cuhR9B+hZflt2uM
j6UtZOrPnUffcfrMqFuishhNEs8AxH+7vr26OX7lbFjBQo+RS11Tw/KYNi8jIsYzOte+frWZZgC5
8BD/CaVIIvN+veba+d/kDy+j9yg7lChgvVzKrrQd7Vg51xSJLQ0JOWnJcOZMkb8iT7MVsbGk5nTz
ymNCkvwwjM3ozkRPsPylvHHkVq33bo/qX8Sqk2+pxnRqlNpjwCuJ6DoG/D1H4+H+4Jr+NakNZq1P
WEra1gXS7pcpE8iMe1jFnf827CFQaCvLT74+bV+wZjMaPqJLr/SBa3m5bmhIkN5x16I3R+iW9Nya
Aq+WKFnpk4CcnYVsKzEQ+VL5o0f5XdrTUj3x+Ac5N3/ItqZ1fhUoJAhViJWXPFPGeqeP2P59Vn1F
mV18hvvWJDYk0qAw22njmFiK2A6l2saz37fXZvZNDz/1p4pPf+J1oBYhCPKTLYdACP1vQf52/kG0
4cL5eAbYFeQMvJfufP8cqcBe6lVAGjqTCBmDwT9j1aXKs6fii46qq5zekDJd6tzZN3Cni5scwR8j
yAwkTDHlT7dpv9OL4tyzq2Ml/hesGfplJ9Cb3m8mGTzms7CK+3Zdb4mSHKG/eo4Hv4Pw7yiwRbDB
TCqwAh6ILQ7JIZ5ey1SbIoh8EtPwmShDQNoS73GKkAApa9yV6vM+zS11EI5vNBJtGR4Krdg2JtIR
VEc1HoIhU1sW/o70nFdGJZmZnYKT2fNF2JkHwTeSAfmaVyqNTQ0W2HQUC41grs3H4QeKTpxxHiuO
TJFNir4VFzqYysj/4J1fxZOe0YsDS9b0i0T8alFN/vd2jHhENVLaUtifU9MdpI9thRCmQoIt5azu
X1YJY1NzAgBjwqSBqS1larar3nUypjKOXk2y5KftOvhPJ18evuc2guSmmzsuAwiwUH4dxtDqE1xL
iqU82nOwv8x/kvAmPVlBN80Xys+pv6foJJSSeVWsIJXN7cR0oWSCUXm4xnoVD1ppSKdyKoG6YEER
moa0ud13OpdzXKyxsuQmrHF0EzjH4igXSWNhYR/VWgI7o5PCjWOs3aR34X9DyhIjZNDNXv9wb9Nz
iLi7qrZ+UzxfYYsPk3enfEO3SnlyY90wyaZo1LILFA2ZUlr2jM/ngGglqoVfrS6tUURIWi1XEMEG
bvGe0821Ulin/VkpKb10X2rSLqS3r8KxojmRmVjivkWzryJj8jtnQL2Oo08KYDrsbzsuaBEDP3CE
AFxFjlOopFEHP4ozznRcbr/kTYpfj7TpHdxCsCECwDfO2SRVAG950yllMJsn3Sd04NXdarhyiK9k
HVpfnIU4w6UAFJJtvViaRp+Kg7GQZbP5E5UHr9bkss3MkS7/FVLdnmfXlU40sg4nPXXf1rB6/Q8n
5kBLVowJ8HcRXzXxep9b2cCTIxuQgQ1KZExfoJdOqavFCOIVGJLAR4yMklNGnOYAau5xXvPw8eIe
/Bzy1h7990IOzqgqB2n17BSU60G7AgyDYpN40vVjBinWB5idzPPppTYPq8PDa7OQy1H9RFVWclNJ
btSUQkPLoivnUNgqAKgolh8LgYVpOyV81z3uIo8D+yE4rM9iVX5IOtjjGmoyzkWsRyyZ8ecTGbGi
t2kUE1h9Pi6UwXujvSAuxLZ5acR69RWFoZ1jbKVrzt2woE/GeMlJHFRXlbs3nvtppCybaIj7pnWe
+3Jf+v9Uxi+1KKPTAKntjhXvzMqvsKbbNPybBSs8eKwNKtEIfuvNs2TmcMRpNP6F4BjcfcmSomMD
dAgvO3ekZGPru6dhAtozsbnQ1ZdnegzdWCX96sD9p9qOVifrBJ8B+DgsAWtAJua0roxWIOivpr+W
xnlZ/BXT93LdyK7K/1+JS9yzyJW0SPKA3T0uFp2FPam9WDhTh92n2HkL0idSMHQVtbeDJ2jf/F7N
nbLiYfaRg8r2xQ+LTz3eLgI/3lK/VJLiByM/spfX2K3+Xi7+TWEEx228NTrkyYnmKyLgAuOCc35a
ooAYohHRaKF0kDuXaLnJZ300w3EfEAQc6xqemU29bxIjpo0HC/owi4vjcfX4auahYe9GKOuihDry
etEEmUC8TJdYse/+NhQ/gainur0z/wHDkYksxcZLu6QYRKLius74J4aZWnstZdQqEL08ehnIWgKc
jBO6VRrCqgaXQmRCzeil7vDBrTd4QQ2dHNrMdVRdC183+qiIB//5oyxT95Mxkw10CUMOkKBR5XBY
hka6Oz9TMk5YlqwNh6STRE9fl+OEGFe43xDCOh3u2jXvn9t/9zVFr7NP0wssWMPYMP4bUTQNY8OB
TrIXb5+tDvqJJ5g0UjyZjqm7nNssU3wG4C+JU+LMJ7XHsQ3ls85uddMtZdQVUx0sTv6qimMkhdE0
2svlZT+aJQm2sDTRJvwKv0HK7CFWbjUNOWcb8SZTV6jtAtRwDBnVFPFfygUqW+JPF35gmRZ0ObJM
AAIOKuHY9oWbfXQO2dQgaPlGb8bkb97aLCZDzT52/wPl8AXvlOHR95S7vWBk80xZDijHbJxzGmk+
Ykh3LypyPHlGXrkl03igB1dWfvISjL1ev6k1KrxLUoceDDFbyl3wLXQSMXfthyv/c4jczf+wK5ul
MbM2tXTyPFJ2orRQ2u49qsAyGeGHrtwWJ6EDB+tq4whgVl5IiO8uEp7ifNpdpmygmxqWoPE2/yeM
juJcwDkV+riDREVMSsv6HX4qTg/VQxq24yhMAXsoXQFzmdSSqMtC/o6gIL2WAl6W06+oB0ukpnv7
pFg0petbJM/dQZj1/xTo6k5hdZ4Qyy017wZjMsaclr+YyDDZnBt1DOUNTAjyZBxiASwrQfTvcaoi
NVnCHrVP4pp7GRrr36Lj5EJYxilQqwKP8u4wLbQ0TR6zQ0C/HxcGFxl/141Icbm4ajaW1e1z27OU
AbL+sjims7vsgAnSMwgtwvSAO01wNUJm1k/5yYn2HP0DMG3r0T8WPHKPYFb9up8vsVjiFVDRFSx5
K0zucVuJkfvJgEBr9pawJ8lCC1V1Caq58exdOYsZr8xrNalC2izKHUZbUxKvWjgacfnHPbN1Jt/4
ckpCCl4lgUV14K6rWYCxGC9zT72K6nxuP8qNC+Zxc6u3Y5ka3kBiqwIPl44+D98hzcGtrvR4bBxQ
r13mv3pS9huwhOl8EzLM/wec3GvMgECgrbtO/EvOZvPWfU0E2N0yvO4AtliNDIx4hzuThLD23GkQ
6vQIWJlx8NPaCm/h+Ibtk1B0tRy7tNArkqo0mdpjkvdEzKji+46oZra03k2wbWeYFYD9Pn2HAHyD
cKc42bPrlab9G/BHUf0DkFjN+t2mkw+L49k4PKpWA73gX6bz0aF/CZCeWGxJvXVD9/zMnqFt6l1w
S3Uu8LZVSMbWShIx5ka4AbWSvHwjj9YKjEA8p1v+B2Tj0esk4bvN6Jc9XKd1Pf0npzna/eyRlikH
mNZsoMegFxVTo3n7NjCdf+dJJKycl4zFC3gpXPGuSvG289/WEdY8XgniEtIu+12aoDyg/qibAFjg
Dpvg250sHdurxe73BZKmahkttTYnMETfEuMgzPvCk03DPAlqDmDu5Gh3cl6JizX6hqCKNF2MalLN
BkCtOcZIJxCGlnsHdbKDbKSTIEGAIKoTSwiZSjm81f4FuCHxB4Jx5jJgJAMr7JCL/KxOvmxBGz86
7nbwXkd3w8q+6Fi/xn+YKwfVInumsZD+lqcHTHrsCi0TopVT1FerLqn0/jd1HdtKtI1ORUXx1se8
lm6ATvG1s3i72Ck7VVKNGubhaTqVJBjMqZ3I63NQgYyjLN4vTzx29+93lITHAvd8hFCifw31PZZ2
vZhKGnK6s5KS4PBcZAfYRbzLdzbFsDWb+Jhc190dL5hqmbHuvd/wrERu16o7IAOTk7c4Vyrh221H
pSWU32IO3U7uMWNmXYtVPdKfhxvmUcylZOk5YbzeLGrO5MUZS/UMCgpcxCHbJSK1P6dHce+na0/w
XBHZ7txM4i4YCq1brtNr8S7Wu9xrMabpQ7dbM3Ikdb3OX+1D1fUQl72aW1v6AsBEUcimigEXZqrW
8umfmcWVWVskCs1rj5/IviPKotGGmZq3nBVqHDhPodkbTS0SutP5vJO8+YSEtiGcmkxUebwwKsbM
lv6GsRnA3P8Qoder5y/gIXyU5yywMre3zRfimHDOYEAj+2S/6xxnc/qXulQ+BSj9E5slK8vkKKGM
Q64JRErRQe9MHvzbEFtY9EPTWtyLC4OlDT/TnI5m7hGn2sA9Vtc7StN6/Bc5Kmdko7oGCaiJaq5/
6HC7JTR67///0/dhAc7TloIDezUxw2WE71tkL6/kowu+9FOiyfsixJNAg77uI6Ep0jHNm+ALni+a
qkERKj1pQSNtVMEXLDJcULk/8E1cnPiEpYi6Fn9jqXkWVxzKR2zxv8ioeCj7lmf3hmcd7vXCMQzb
CY1dURevIafFUDFJI1eP++dk0AEy2aALi6/ghv10kObFQy5RedukvSxtfAwOZaM/1Yy3cS7rJT+r
vX9CVDXW5pMfYyOlUbao8yg1vZZg3lZXC160lDNoiS+CTdaJxPm86+KSce+geWjmAhWJqgP4KJBI
N9CORPVlcfHO2xgLwk2AOAPOfRIq48iBB6pKzTpkX5zJtXHYtieHx46tZUJf5E1E6zXmVkYOZuLx
rQL1yOpTqRyUf0r16kIthKkIqCWnuK7GTigEkgOCyCytO4/l8ETf91yuCxPs/cASETQM9BlBR6RU
MgCFNTgmxBlP9SW8EdGKcznIAWK+ezYKQ/pCyNE6TPSSDK2E99KqxQIH6Fn4c924uOCAfd76IKqp
QykeXdg8qt3avcqfDpnSKg0Di+eapmm7XgkaSYSti2DbmRcLAO9oQEiV/VuTgZmWVo1Whgc/dld+
g4QaiOOdCOSnSzYlWb+uajzRqEDOer+y4HhQELG3zskpLuI5ed+gp+MWVoIVkVyHSW4OrRz8jMZc
x2jdHBOGeUh3g7dQP+GZy4Q63GB52DgnfjztO+GFZY8fnfnykxOqLwsKGmfm1Fitc3u6UaYbYGBO
JZRnXQEUjLJulooFAL7oTlgpueVY3pquuTCtFeRjLvvoNp9AVeTMo20m2toG4l8KJRWiPbIHJTj4
lEe+Z4DDQ884XC9ng5u1JaYQQUIKe4YP9ZrX/zbVa1se1o8z4X5eRBoMav0i7H9mBwIKa1S8CfbA
LqwN4hdYp2XDJ7E8/sap+/LSxJIkJKYQf8Z+t84ZYrIAWjHAvKnaRQy5JldCmDsdEgmFUNkrxJ9B
HxCwKD9PHJ9PiRgD/AXuh78xIQYhR5Le7i9gorFice5aoRvKEYbZEbSciNEowQyT42LniPjLnXMW
H0hccJc7sUO4E6YN2uOsyG0n6905pdWOy42P30TA+RXdqP1oG4o2dkq9fDB+yYKlJab+OkKmvNxo
Snbs292HHecyW/13LA4URZo5ZcuMkzKjPtyrgs5ZaMKfhzYiEDIkIHisGxN+4PjtgiNZUMH0c5nb
/9NLSNej+xEENrGm3lTOrhLNIJLk1iZcCPEx5pqE3uzbJdEp6qS5f2E6wVCZnfyqI9ndYDGj7WLL
GB9l12jE0R7iwgDJYkhw+7PXTGUryWCamiTxXPkh/L9b+rDxh/P5KfOrACOlssb4lOhkHtfVi+5K
Itv+IwEjQwDQSiNL8mgW2OSwZFLdx0YY+Bkl/A6ynIpY6VDPfvCVqZ0DJK0TOer7oTPLg28015uB
l46Cnnb8GwYSPH8wla9hYL3lXtyE2GLP7qR3d3at9PJ70fp9sCZHsNCKB6MYXfJLBt2QmDA9by5Z
B5jaSgeVt+aB8dxL3NUNz8ol5iv7/4P148KDG/QPG9JvlBLJ3Cl8tMzxuYaYrP14GkPLsPLcpj2Z
F/LRACG43hP/LVm+Puf3NCGLgI0E2ehRy6Qq09lR/XcykMzKZUA6GCswCk7XeOmRivq94UxOS4eA
YtNk0dLOFH5V26YvcZNm0q7h6RTbqGUzOLnsipVCW2HsRS5OTeZoSS5f2YWNOchPODb7BorR8u+m
Ec6oCY8Kt331FDIJ/gAtGmWYPoL17yslQTlheXaoaangymx313Yr4cnFO2eTKfTcuSkHFZ9lv8Qg
SBMa1Fx5NxEk2dbFzIgIqoQ1nanH4Stm2coLkZ6fgaxjSZdnzfnFgmRMxRHuDXLIZpVr5D9ogYpb
fI8dZfIRawWQNJ386QaIqTjdTyN6e2NyxBD3KI5wEa/9O5a/8WnFfWUV41G2r9IaY9YrXWBlAK+K
VbdEdCrH6m3f0dYIqnGOo0MXqWWf6NKOXS9cpHnaR27UWOgByaCbkegaCThJWzTOY+T3cXOASMFG
i+onKre9r4pF0HeWt7d5GVcKMsP/UCdbJlF4Yc94m1X1BMPbXYliG7j7l563rLiLchhbSlGhNge8
Rgwwe3EOCOPOgBkMWJ36B8T6MXV5acQkpPFhvYPtq3wByxTygMqa45QdSZlSwVnqgDrJiBXAO02n
/UBdqiIusMIldWkzDD78F6McVqFcw4IXd0goi7KVuLXFi1W8mp0M1E09NuJ9KKaFBD7ThHdWUzg3
1CSyBQcIARuWbpkmcsvNCU868SP1nREbCYhS3CZa80C8YAPquzQg7yKQ8lMoloIQyj8wHgu1Zncl
6VD4tKH+GEI1EPDRuxnOpowbFm/WJ/5kOFrEt1n5QuEH1BTnfVrlo1GdTFxIt5/e+uArTbyR3hPg
Z8W9Cs/U3aQrjkJlUwPLm2Y6500IfG57PzowSr1kR7j04Vv/TKh+f665yZ72/+Bz5ftT3ArjVwnz
hZA/LNzVSCZrtJtE/XxXDqfTvf6Gej4K9Tp0T+Jw/2490hpoPJKR14HPfXxe977RTi2jPXUCKCyK
armV19Wlw6hq7X/tINyiTzeARZjQti6woJzYcbpCs6F9sl4Ek2aYsHRmjN5Vs0sfVNFFnib51GkK
p24D1BPd9rP0vxIU2KS8wnlmYQ63Rl9A9jI8SEkuj1Vs3tKuc1h/NqPKUuTGcJ58vU/XcMOX116L
2J/yLNZx602yIgWT25iQyDTI2V7LFjEYDtymgQU00REiRA4O3uLXVxWIHxPdiBZH14KUBdkqXMw7
ox1KHBg98NGCCpKsKFreE00jCvzIFqVTCTDgGJpPNpO+oGF1E6vuQpWsCERjviFR+mPgZG2en7Yn
mUq0jAnf6Se5+AEyuvpX5l8UsGFqqSOG6ABVRCYUXJZ+bAYZWvzjPNgiwl2VHrJjQZPwXhz1+raf
xDUqSOZnA2OeL3vtGiZDV2W9bLA88yfZxy+gqnTmRWALj3TCDClUmR1Qy8rlCSM/sNC8XxfOJGTQ
ow3S3RdeJBU0ZzL4wLoss8X3qHt3O5I90enTOctggTfP8bDhonio+hC9IqQdfKjKoS8PnIXAaUi2
BvW6aQmH6OEO1GgAud+vtbVUlXE/jrNKKEFClTigjvSUlQXhrvdJuorY/NeEGNsnLnmkZ5Y7GgJq
4ps9oZwdROwJTE8rSoj1NkTzKR+XtlSpTiBUCP3BQ+7QPi++xI3IC8tpTl89jUI2AyUQynYlrIbn
CJ84WbpwTgqEIi1/oySu4eCvYbB31lt4/KN63M3vRDtuHMUNtB/5yZ0ny8tSYKFqcdKg7m5FkOXL
orBLvWVS7IUysw0yeX10GQg6q6h7cOSz5hDAnMi5ahOYR/IJaIHiIl7IAsKln1ES3A2mJiNwOBdL
x4Glc9/s7A9h6itCFttZh5lkytNuW1z5KOGaZXwkaAwYRwLAfDiKDTFpdociZzePC54Asvp38cRo
FruNeIbS8O5qPzttC4vSocFEkWXyNLfa6p7gFXL8gz2hUiQFSZRHLku2OgNTpjP2cHFBVx48wC+Q
fk1HIDYWKAnPfL5nxJEcTx09escxbaaA8zneoe867JbQUPC3VlkOu2ISCd+rLXvru95JM4dRCbGJ
GUIdc1Xdm0ggo16Tj73A01p4sxx9FJlsc11lGMYKFAq0G+8jLBUK8/XKnF7FpFqeFdh/a0h5j4sv
3bW8a2PUhY1ma3C2A7VXUyrDBkagOWIgHn3ALAVD/Wh6SkLML4/I55kYAHpE03WgYcsepemwpqIt
gbx40w9eYQ5EcIZRssggDiUrm2d/3/+5NTMCdPEY5YYHKCKsZ+fvEglSuCko8lva0qSCmEkL0UGc
iBLtbOpgrzce5qGKvyasqhz09LUYx1+ejVmXy98xNRc7tCnuD70wKbObgIR4lRg+a/o9uaIl0xTo
ve4tSW+3HNRHdJnFlFRJkNIVqYNjZWEUjlozHAZApriu7EgOdxbtwcJ6idcVZVnlPL1UsXriWqYF
feU795TUfz76nOBRiwASAYarndVG+8755J87TS6WbNx4RIdrv7f3yv9kuGmfkh9fpa3rNK9Xsj0u
Haxu833RsH0+LuxdotawvhJhqW8niKp39nxrHq5k5W0l4O8KDfako8Ne2iE2WDf3zfuuB98BCY/f
8zDvzTS0yjU1jP5/K4mbdipdt4HxGILWhd/mNFTLEVBLNfJZKgwWBQYpy1yE7I+HDfDPm0932HmG
g40uGhjmylpIpEZt5QnsMyvnaT0MbNhEQXpHfJg3YbJuLipMyXdgWyRqtLCOxYrfMJlbVGXsZaVh
+9jIH+0ezoFwv2og2zqE/lDxE8j3jMNByOtrR7K2+2gmxpA6twSqLf9MHBVdpEstX3EURgBz8yTO
K1/bvbN4mG6M3B0YJe/QYbTPLbVg13ElvLqORNfIevseslrPNW9NNznutVljMIWoCbpK8DXOFuJu
+P1/VVqhTouIapTwmDW2t6aaXY13miuzt269J1ZzWJTglwjkFybTWlvTIdixs+w84Xf8liuXOjA8
VIWfpxd6t/KhO99OJwKjwT8bUXUgo6D4p2sK5lzGyJpnlXOquNf6xcLpoFZ+RmQzZuQPnBCZL1/b
rZH00i0uqpZy51oRQQnajyWPNBwBDR8mGuQh4JgKM0TytwT5dx8/z9CNPxF6qolxDn488vrzbyse
/jiZlEyE15TzsXR3VzawXG8On6vtL/PTA1mPJ6cODZpfo5o6nmBbiM+uqnuOrJGjUNqngt983BeR
QmnlvbnyGX595qKt/3ZwzKxLHGIqG+R+2WYUdC5/WaBFWHpCUKPK9+4Cj423W42fNscSm99nkCUN
GrtxTi88eLOGuDZMbbMcSf6oEpAMKOO3LUzH1KQhX37co1CwhHhDc8Ayp55p9wIQLh6dplXUeNsB
zRnWb3IF/qBLTEPraQI5J0deo4KzyzR2GINX55e+FsC89iu4+gWAuy3K/PHdw27nyzi9MqSlFP2F
28n7XQSyEL0TWVmW4TKn+Dm488LLqBC7my1SKFqEOpCv1DYQX87fYaxWPI5bghwwXD75PsXySHZo
sqcMIJWK6lMg+6onvw==
`protect end_protected
