��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$Rx�y�<��wA�*;�x���@�̦�W�X�fa�M-$u����n~�%���P�$��W��kYَ���P7�?UMfT��q�6�U��k�>����~�\N�(�����X�e���/6U|)�X2pF�]$h���d.���9E�	�IN�f"�\��e�z�y�b�����Oo2�?�qˁ'�͜k-�K�P|����y:����3�l�d���bl��ˢ_�d���kx�rq�mh�MذM�`aS�.�DW�mS�9���Y��+�>��!��!�T�uOB���,��\L�7m�O��W���6����'���j)n_�I����2:��$�K�2�Sʫ��l ��!���{�l����.�j4�	��很�̢=�����N��s���s5���_�R�>����ТP .W;������	�"�מԫ�����]�#7@O+?�⡾�Ԫ���e�O�\A�	�ͼ���ƹ�d�	@�nQ˰��E؁Bf���|D_�%au�-�'���w�*%��"AM$w�*Q�#��q���!��<�	+"F���E���C�)Jb�5�n�l�9XM�;~��[:��dl3K[]���qk
.%��T�.�Jz�f�T�R{Vuu�H35�ǩg��|�at�
��W`�"�$��=�{X
���|�����0��}4d	�?�5�L���ʹ�����p
ν�������ݭi�U_a�f}�B"�>��:S�A>�:iŐ�N_����Xuk���eA=��ϋ�k*�qw}�<�Q�E��?cgmʚ��XMm&� ǶҴ�YY���nEM�+U6��n���tp�*_,+W��Ax:l�w$��O��?H�lC�r~���Α�
��u�$`�@!	�L�����ɽ�\ehvh�+���.��+{�#p�m�c�j%�����hg�� p��x4,`J��h��N�1�.C�t=5#+(�3(��QI}(�k+R��qO��nTZ�E�����M��$�hE/ ӳj���R�K@k!��>
O$��w��d����_7.70�'^�y��*i�4p?�
@&���`��N�.�8��MԢ�~�D'�)�[�+�`�v���T�Q���3�q��$ْ�1e�׼�Ԉ{RRF붸���:0&�,(1�]6^�V�tx��^ѡ7)4�bCdJI�ݍ���Z�I�v�������#|�KL�c�^��w\S�E�b�'��wG�Q�� ��E�U.'cX��Mi���ah�H�����!�����;:��:�5l�H���ז���x�ˎD���e\7�+(kR`� �l�`����^���!}�i1^y�=d� /J��8��>��+qch��A2�����Q��q�|Wྐྵ�����5p�����P��ܨ��?�3p�'g��Mq��>�`�h��fDٔZ�lw�������o�*BAzX5'��^?C ��؛�vOS�`�<�J� \�J km�,�;B��������<7�����R���U�SO]�?,� �#�[��"'+�jÕ�_�L����Hn�c�n�zL�.'`�э��X��\}/���@{v!�a:�S-OYJ=&N䚀�{(u��#�Q���r�	7 ~�>�y�Y�G��C̈(�,v��Q����\�R�����y�%Z�����^���.�ѻ�L��^���O�lhs�֓�M���(�w�D�~��
U���)V9*�}���ߟ������/����̤��>�^�*���)F�R����L8�Qe�·��l����+��.ua��ǝS����͉ﳨ��"E1�j�~��7F ���x��dt�v�%���Ȉ�����ΞԊ�G7$B�a���JW=���J|_���-we���{<����V[��T�T��@��K�c�%`+�6D��JC��=`�x[X�,�%T�^�[�IH�r"�1�?��.�ݬ��Տ�a\�͐��p��O�UP�ۮwI�|����OU��%~��l�g�]#$�>�<#Pl\̗\?ג5G�P�~��U�Y�Wrо�3n�G��VB�I�iw:p��k�����;ۊF�H��+)�0E����ݧE#�0\;��a� �	�#ooD>���Æ�̫����?T����"q��â�>��O���f7'�AJ9CK�8Spar�4�p�D�"�������d�
�Sj*����S��>��"Z	`�gP�key�o��e��܎�Vo���I��'o�10FZ�E/�ǝ��K��7�@OF�Q��_�%$D]S�y�~P�w�Ս�Us�)-�a�o6}r�o���J�y	:Ѭ4ڙM]
�����X+kN��%�A����Źu�"�c�u���ͦYY�V]cJ�ɴ�uu�e��0�-.� ��5ʦ�����w�p�(E��X��/W�W��O�	d���mѻ�Ǡ�a0�e�b�Vp��	�A��N�[�#�F�+h7+�}AMt���;9H����ڷ,9�# }M��ܛ2����-$�٥��Z�Nϭm5R�3����Z#+�+����֑ݔ�]��/���g飳̷ΐ��]u�+�Mc]��o��!���݁�j�c��4�B��X��>6�aj8�"�f36ӗ5�G�8 �c0��9��~
��D����SYB pID�������:���Z�Њxg�9Pa������/08��"������=�����J��=a�v!<\�b\!������@�g3HRۡ��`���SHA�S�y%������L�=(�_���0mtR.y0���R%����m�p�E�,
\kC=�b&�&YJ*��@I}�E����ok��ݕ��K�7�φ ��.k��T�Rc:٩�V6*h�,|��NT�y	�^.�TebD)��a�o�٧/��,�
F;��90n=��:��k���˱pӼ��ubI�\[�^��E��&-c��I��.؉��P�~ۧ3.�lN�Ԡ�\h�^�9� �nh{*��X\n(=��l�ȹ��Q��J:�R2�u_e�#r.�0�9��~$�9(����{*e��B�6��!�q�ej�L�u�1UN?�1ԑA ^��i�g��jc=�
R�m7��N���m9�C1ƒFz��/��)<�-�Ǯ�j����%��(����;PP�����E��O���<ǈzE.��+/p�9Mq�W�^-�o&�d. 
�-�\U���ѭm��e�K��L�.ݙ�w�tQ��B�D�T@�L�RG���lh7�H����<�՟���bN`�l��ѱ�����垕�x<�1�S� �҃��jd���
PL�G;��$:�����|� �/UP�H0YW��6����� �"��N��ٔ?»�w��)P$ب�g�U��B� ��9� f�Y����U�(�#���j��/�蕍�0�By��a�Qv<^��(��+)"�_"�4�ҕ� 1���s��q8�,�{�}AS����i�L�6�a�5�8Wɸ�����jQ�m���eS�N���ed ��j*�-&fz*Y��C������՞�<Z��V+�|~�Kc=zh�S�v�����z%E�S��D+E���K�.�[}К�BQF���s��WZ����@�P4���*x�������{4�Z�9��� H'�a0��I�[���1 :#�M��$���I��ۛ�+G�����(@�I��_�	N%�(W�8o�����\�"{��փ^A�m�C>���8�92��n����XX��Ы�ctx�N.و��I!����Yר����7��kE�9���3J�|��H�(��"�3�K�l�X�&������S�<�Q���J�p/|���̵W��L�:���iC�,�on�x��
�����U���^�F2'��r��a�����j�k�t2�+�.)����.80S��K�^���hJ�;ɸJ�e!o�.n�响-���5���FH 
 ��rP'b�L�t4V��Q�c��yq�c��&1#�
U�Gvo��xί������>�f�-��ezs����'��7��1ۍn�@��H흐� 9oq ��T3�X��V5�7Ƕ�Bm+o�s���qjJ툼�Li[�"���c����O0��&j1" ƺ/�֜lh}cd��-�.�5��^�Б5�j�Vs�Ӧ����9�%���<�<˽nk��}����a8����<�/ ���H���|m�bNyh܎�f��\�P�D��z�з=5�Bڟ�J�j%�=^��}��e.�q����і�YU�����8�9x5���Z�B�q���s,1�E��?`��0��`�#�s�"2c�|�ځNw�+r/@C��}�gN���
���6�x�~�҃���p�X����F!H(M���ORu��Q���ǒPHZ�LbE�3	���gw��|N
��(�U���n�(���� N�)��y\�����`�h/�ջ�#�'ݬ�c*HO��ï���pL[�1���1�-vհڝ��@3СyD�dOZ�z�Y��w�g��4�|���
r���1B�aDV1�el�m��u���o@�Z @6S�aTe�QAɺp Z+�.���B���U"��mE�=�
�;5}��53%GtP�;��J�6��vIo˕�*	�A_�c�Z���+�l���)��*��G�c-��z��[z ��\වC����WtT Yك |�'��H1�mT���0�	p[&��J�j'�����ي�99�����.D�0�P
�̦�B�M�;�iI"u.S�_��8{NuȮ�qt�
~X�0t�Zक़yW��6�3�4ޱ����%���:wwfA�Z�%j�٨u�
���U���s���.,��T`k˘�O�_��7Ǹ\��@$�!�A�+��M�:3�k+�\g������kO��Y#r�P8/��#�2���UQL1$+ڲ�k����I-B�_���gh�����]�/�B�(�w�;���8ۅD�z�����Xo����j�ۓ�^�&Ok�%qVޜ�߄2/j�≥��߈
b��w���q&�-U�p��,���('.7v��N�'��/�d�m�����^Y�S���f���1 �9�K�L��s��D*8t(�93��ZU]��/�&?����x>�����h	Q	#V	>	fC�9��ύ��s�� �Fج���%n�ќ1����t�^��k�8���Abε���\��-\���Y���H�n:��T
PBIŶYw�$��t�>\�����	Yش�8}8���@��B沷����;��-
f����=� �fx�(g��=�J@��K�b�	פ��deniӍ[ȹ ��jO�+Uhk{��;��,��q��L��Ի/P�|����ʪ�%.j��"�}h Ūz�|���}p����dH��=@��N�Y��7SPM�F�B�̝}ɠ�W�|�	;�࢞\�!���ך����t_����)O�2�\������N?���J�,�⫾M�< e�K��ݹ���u��7#�]�s�����Y,�&֑RE*OE�`�{����J����iK"�`=��V��s;@�%D�� 73��!�2�m&р���'aS� ��4� )flcb�:�SL~��0���w�S��{?��OS���ZS�j��O!A�\�����Y̛y)���X�����o���R\</
���48Ѡ�)�30f6��Cs0~1f�������27j��!$0�sl���|5��3�Ż��Wy���8��a/mz�l�M�y���gx�X4�kC3�ƈH�	���w(U���c����u,���Q��բ'z3�ֱ�`��ᡩ�(mk��{��������Xlo�'?{��߾[|�Q�X!�5�3�����g9�f��Ō�f�]��y���JZj���6���DD�p�]�������);_<F9�Bi?q�0*�]���B5�u������*�k���\"'g���]���c!���s�Y��1���#�$�X�op��`�nq{Kh�X���=d�Q%	�-U�,�����rJ*['k.��F��đʚK�Gm���WL�ӝzq�TCT��W|%��H��PڣmΚ�_�v�4���>G[�N�Q�Mq�<R#��7H�전�T�
jpf�I���Z�? ��U:��m�T��Zc(Vɨ�{���rK1ح����v����5�Kee���V���kI������� �&�ɛ��uG�N���١j�=�5Ī[3���<'fӴ����r��\[Q�ZFǔȁ�;�D�sB�T�&Y����4��Z��T����_W
˞���'�pSZ!Ӑ*|T�-{_H��V����U/�Z��mt@��+�kpڌ�b	R��V	d{Ɠ�?�p�r3:%<U���1�iHǇC|4�a�3��2�2�B�=�Մ)H ��"%L_�؜<�M-����Y7��:̂�w+u� k��U�}w��d������`����\l�ZM������vX�EXӡ���`�r�j{*h��6ے�?����_ȎFƬ�}�uB�����������pie]2W(E�'�rxBH�j��d������������&���j����+DY�[,9\��og0WԠ��ۺ�s��F����i+�u�ɔ�6U���m.����
��+ޡc4�	���AG�+�U_i�נ5X����V�)�fI����.b�Q��vDB�7�M�J�S��:S�U~��z
�h~�t&ޔ��A������1ͅ"+�YR��
��*	h������j�6����+�f�(��ZK�5od�Ț�O��:D;�-�:�n}��FS�.�zQk9A����R�H�T��N뼸"����M7f?8�mj7>Zκm1��BV���0,w�;+5���V��Ss�i�yX�u0�
��J_��D��Kc���-Lb���ɣ�b���r:�.�����4���,N��I���so⾹�yҏYm��?]�K@�\��+�#��^��z�8=,R����m�w}�V6\�k ��ܨ�_lm�ƈ���}��b1�������������U�æv.���N|@}�x�pQ?[)�P��Ճ	����4��Q�޵�R�����e�d�lN��$��3��7r*����f�`��q�jGA���Ĕ�J@��i���!�w1>��ar,)�`��"�q�E��%d�Nv�*e�BA�^=��ؓ~L�`w����7`�c��#x���s��iU3�u��=H^���{�C��:b�k!M*n�u{<��j�5���$~$#U�����Z��ta�Z��cf��Ds�0�ӴH-1ϛW�HK���Ƥ���+� E�/���;C�4�=�����L;5�ǀ�.��D+�N��&�u�^i�_��h��f�>�P��Lܖ����B�M|ˠ;A�H��`��m_�%@�˗��>�arD��0!�<��X�&��9Qgl ه ���}��噓^�im�'���S�u�l���6�V2A��S�B��:FN����¾t.�����(����ѶoM��|�:M}|9��h�O<�kw�Y1`���i�u�6�]Sg6,��K����.'���e1at��V��}߯U>j���Fd����FԈ�4%����
_������r*���%l������>!��c��o]��K>�j�ܐ!�0mm�,��WN��C�ƺ$g��ńW���Y�y��k���F�{�:���!���ܸ�(�t��[?��������U�x�"E��1_4��2����S%`8X\�ʧ����|9�/���=M�Q�؍�k��!a������O���w�3˟��� 5�Y&����e����)�%�l� h������O>O���0����J��B�CB� ����z��4@�u�A��Ma�F�j��R/��=z Q�/B�(m�&HJI�y|*o��u<����f����LBA�"��k�@�Z'��v��m�<����*�J�J��ғً)��m�i��q�'�#�T@�Ǎ������_i6mQOj@y�]Y'ψ�)�(����+�&A�@N3��q�ߚ{E�Ϯ�rt/�Z�Jjm��3�L!GR�2[fC��@��A�;�GA=�� ��ɓ�z���\"5��M*�M�ȭ�(L�.�y�����`� K¡��pzw�;�j)��+o�VH\�}�M<;���%p��x�p����u�4��t�j��Q:1s�Lw�2{�δ0�:G�J{ܕ���Sգ���q��<�"�|�g�;�N� �jhS{���A�X�G��S�頺���in��q{q�o`bW��k�6�uD�&������Uk�#!�3������xQ�$3
\�C٭���#-1DJ�An ���<�ͼB9��`@GC [2��+�t��-��U#c�#���bOKJ0�s�lޮۃ�[D��fW�{\���s����<ؗ�Ւo<����g�	e0/�Q2�\ӷ2�ŉwdn���"�v�{�9M�]�䊨���0M��>�����toI�&��U�E#wB�3p1W�u+ ��.t��pw� xr�o"a×�^�79�d�Ř�ɴ�� �����9�{�itNU�� 7�C���#�Â��bt��_JS��x`Ϸ_<�/�f���J���69�����=d�4�g�fe`o�F�A@<���	���տ�As��4�,�k�i��P�|*��N�
s��9��b�L|u\����}�#�A��G�Z:�a��y<U��ͽ�WL%���y}�U_Jm�>II��Xve p�ی(�Ӻ�Tf�.�U�lj�����-TD�$��"�6�֞�o���E��3�7�n��Ca'x�KR�~�9�zԊ��O$�ΘW��5:�c��l�cJX���J��N�Ŏ,�Gȑܩ �I��Vީ�C��@�_�⭣�����Px�'6�5#}W\�_�a��3�:g�d��2��d-��0z^Q������������l�:��!Ē�� ����L����yo	� �e����_���'�1�N�$չ��ӡ���46J�%��N�ڪi^�y��Q�̢}Ŕ���W@2���/Mx�
��+���VyY���Cy����Z��$�8�}�eCP�uTB}�n�h������B�F0@Hy=�#x�s�x;���;¬C�T�Q������1��������Tm����d$��VنwO�B0O��<�6���H��+Zv}��*�[d��
��y�b�`�2Q��}���K2Tlff��+������*��%wv�(��F�u��)�>Z�ǀ`��]��+3�"�=��;W��#�n +O�M7*�O���,���3]�&��7�\Y�dW�D��)Q�����:��S�n�Ѐ�7�Q�}��q��M\L�yZ���1�@x�+�4�}֙ ���?RU*��G��Ip��Py�Ym^�ޘ0���A��$��#8��g)_��p�b��W���u��܍U�7ԁ*��)��P�_y�Aa\�zY�����N�q�W2�i��������r��R�ѻ�n/v���b0%��';k���9��S����<5�����N�ηԜ�z~��E�b�i��h����.�>�4����3ҫ��yq>��dT�ڧZX�%rG~���V��Bq0�Eq�Ρ�ga�A�3�d:�X����` ��b����Am�������Fn�{\]�ʊ䴠���݋��E�#��U��1BGMh�e���tzP��{����I̢r�g�$����I_M�j+��]K�� ���&�^�����\I���QJi�?e�>�x�8��&<�Sem�8�{�?�^�kD�	�py0i��1E�5%=�+L�����,kn�ȼ!@E�؅�Ea��.y��rn;��p�
[	(� �NC��Fz��6��Ea�N|�5��QoQ�>ր�_�;Z=DK����yo5^^7�uX�ћH$���5v �doK!�sa�6���ٔ�8�#��]�/��&t�L���2#1"'��p��d�-����s�i�zP���ؿ�YQ{nM%@����y���6'*x��!#wq���������
�-Q6{(���ڲ�h�,�$4�H�1�_3�Ld�����AB�Kl�Պ������23���Z�'�/��̒Db@*�&5s>�Z�:�77��!�!n�R����b�}~5�i�}�fZ?RxW�ĵ�*J�Ր�v����=��an��`�5��8:'�qo��݇��n�\�Nn��8��L/?q$����z ji>veŭʓؒ����ڭ>~�ۓƳ��r�\x�H�m�6�1���x�NTW�i)�Z���F��� ��x�'�$������
S��e�4S/��U��9��G���Wzl"�*��N*��|�j�������[��.��h�Q�}@^�B��d`6zI�(�m�g���26(����/��f������g�/��"|��������� l�bY�L��^yw]U��G��ӆ	kÕ�)�B=� �'���W����܄�yl�)zP�ڊt
M9�*���_���L�$}*PF��c�1�$�*��\�a} 抚1��O��������kͼ�(�8���N@Pf�k�D33��0}u`�X>�5��Y�֡�-��lO���"�1&B`;ߨ�]����#�j�S��$٫�_�����b�S,�G�/���#��as�"��O�۵����ۗ4WqA���P���vU�B����^xIÈ��Q��NT����T%�I@��If��:z�@m/(��W�W�M�U"
:��qÝ ,��s��f�7b������5�
MԌ\�k=����	��>ۜ�6�7]	e
s��?;����	�c�K�O�eY��Uy�$T&�t��R�}7�fR�`�9�{< ���hC��)H
�(D�>C!5�8g^�D��k*>�53]C�P���*�^'���?E:�ޓ5_���G eQ�	�'/�3@�v���\�Z�XGvZX���{�N�h}&��l)ҧ_#Q���~�J�!B9�� ql��Sz��6�{�^^�?��&�e��+p�� ��&�(~��~�y��{���"��`��Ku���'��f�_N1�w)�����l1�-�}pNȆ��~��a ��ӝ�NlӼ�y��e�G;Y_)�׌9��>��r{5�ȪՇXӽs@|n�q���65X��G9&iq#Eɡ]�h!�(A�ZG���AF��.&q��a_�<cv�g��Aƛ�tN����kja��vZ{���UJ��|��I�����>��/47,hy1���0v�%�J�3T�i*��?Pͤ@��&��TW[!�'�ޔI�������ͅ���7��4���눠1l�L���#߬�m�4���uH��������"2>4y�g,7�ب���ޣ(]���Pwy7��RO�=�.�W�o�Vk̦������:����+tٷ�c\o�c��o۷ص��q�
��=�q�^trO��b �.uh����?�?���,%�1L �k�{�CV�g���|c����b۝4$�c ���E�g�H2ˇ�&ĶRԦ"��ڤa�����E�<]7�
��D�=�*-�W�S��F���g�@��B��|�i�.������~eMNgU�k��CT)�<7����h�%���0Âzq6<��f�h�ᇤ�����5N�) &z�Y�艱.���BIE�J��x�<��H�ht�:�VҤsd�5]�P��f�Hqo�`M��L`@��Q93�<'�{��� �tX)���Q�)D�f���ݿ�]���!բ,�Uy�c����Ǹ�J���]0tq���JK����Y���J(aU�A�Tq5ٹ�I���;�~ (H0w�$�bg�CGF�@:���nb�*����.k3'[�$�P��s�B�̾���]���B���݄˺H	�i��P_���#iq���Y �X���̰��[���SӰ�kW�z�[��/�_����x�)�D8p�S jk�V�&F�VPQi���O�lǌ5�O8 󳂦72��8Ħ�Le�|�ډ�#H�����K)s��4ckvaE�iհHu�����?�	��j�����T�֤�*�-���)�oޙn_+P����~�7��� ��&Ǒc� �ݞ�7�IO�6ԿVn;�'�zh�Q��3c)�k�J$*���o'.>�Nª�Y�sS��8[��֯���\�ځv%kuά�1~ÂUjJ� �
�Un`��<��=L˛]c��D*+I�p���6��{�/��4�hsB��� ���.�	�����_7r�4w?L �^2$v���ӓL�t�wNz;ql|��ޤ�5�	�x{�g�
�Y����j�h��4p��b�87:S#)؈��)D(�nF���}��:�(t�_B"S0����V_& �@{�0 ���t)ȹ���5&���y�a�o���+��"�k�	�Av�1���F���[{��4yk�<��ǫ!&�zz�#q��*T#X`�ܴ�]I\_Ƶ�Y�2�����\��) �9�W��m�L/u����N�-R�P�Q�6fȠ�=r�;G�2T����c3���(�r�!���|X&�ۜ
�q*����p]�T�;��Lh���v-xZ1���F����d'���$��]�E�+�?F�����fU֚�ܤ(.���,:3������'��`�;���m��.��9$�_n7��\"�P.:�`�.�A
��{E`�Vr�uK,} ��>�w�ݬ�W��<���N��7�A��Ѕx�7��Vyi����cH%?�8�ӎ
�Ms� ��!�Z�y|6�ڏ��{b�m���D�?{p̢�Z��Y��U�pH��u`�HEP8�����;G��G+������8m��deE��K�� 7�UOl��p���/ՏƱ��믹xb"��NP1���Ԝ����v�}z��5���r�����܉=��㖻�8�	��ᫍ}��{YS/��� ��6����H��C2�����o�J��ɳ�Ѱ�LtZ�:Ȼ<Q� ��	�?��HUB9�z�Ň�HN�Z�k|}�xZ�A2�	O���:�ѐ�χ�~ �:8���`yA\[=�#?io]_�?�6�����`�o�3����[���Nt�?�\kG$��&�2n���<?]=�����m�m��N��eL��md@�����n+bwֳF�
#�ٌ�����@*��?�����o��z���t6feN���]%l��O"B2U��5�i��� �E�k&&{E���`����!�������>�H%L�^�D��bwi�m���R�Cm�Hn�)z!oV�_#��7 ��A�Mm�C�$�{\e�L �<�I]�:K�\�ҽܝ��B�@�omCwP�z���H�ϝ��P���'�������U������h�g�[OT	�%����S9����e��_�4�>;�q���mY��*���4��k�=P�ɍf*�!���.U�3"��+,0�[%�:�L�r�J���^����V�9����Z�R^�8�8)�"�rV	��.�_���=Ƨ��M���cZ��Ĩ*}���c���>j�_����ߪ�҃ũ ŐR�F��G�	 2F��n~���Z���'�_!��SVI����jջ�2���u����l���\!:Ga@؇�U��l���Գu=~9e��4�
��Cr����&t(���E��/D{D�C/U}�=�$�����~���Y��<�1�׆�n��sN�/�T��餵�˞�9�E��В���!�x�}.X��1���!87Pd���C ��+s��Eb1�5��.������Q�=������,�E�ޛ~�0��h'���vt�2������P%��#1�N�.M�}���9n�&@E���|��|�b�c��ۖ�����w�����呜����tTo来h�u�	d�Sg9IMp��"���Rqa�[�Ux䟿i�dO ���\\��B�R�\Mj��p��rjR����l]�24m��N���(KO�C>�!$��]�jY��'��������=FI��+E,�*A�U؈�_��;��(^O(�L
N��`VA�"�M��`�?FװĹ�D��	#@�R�������G�$�7� �L�a,`X<���::�=_U��m_K]���Q<N%�]g~nMv�\S� �{ku��w0c�y�U9���8�ݢzLv��>_�H��8���z�����`���C��!_�G�m�Q����g��2��u�nTө�Bw�ge�}�����OO=ѩDѺz���k�m�2l�1�Q�N~4��(� X|+�(�m3_7��I�LP��:a��\��fy�	w�R�).lB��l�T���.�w8�v��9�Ejf_���>E����!�t	�M?���A�I����JU�L	K�')(�[�tu3�Y�b�F�
�+�k��a;��Ge�}�$����!4w?œAT�/���d�E�/�;h@���\�aR��MٸO��C��a9	�>ta/-�<7�w�+ث,o��)�d�/kg�<�S��^���T/S�R�$�ɚc�~�,���.�#}�q:�0���ȅr�{T!c;��щ����˴��� D&j�'~`�^��P498�C�d�G<�V4��Hh�OoG��"Q�XE�%��'4w��o{Ax/�}�+\�����b}��}��̶c.��^���:U���O��Z��$wiJ�px���j_�ɏ��E�5����,�I%u�Y�(��*�kX��?�%7�^���&����' ݾ�ўO�!7�5��6��[��'��"Δnv�k{�9V��O��id��I[G�@���LZ�$��gG$nl͈D�C��9l���@�4�Zj{����o��z
��%�;I�m�--2]�_k���T��_�+�T+�����W?M���jc��V�E���Ԃ$�jG[��Ck������|:�b�`�9�#8��v��}�I��~p\�	�B�d2�����G~?����.�q_�3O
a�evA�aw��1���xD�da�>f��j�M�Q(d(�6�I
=ׯ���Ƨ{Z/T��At0\�1��7���5���sӢ^^���K�g-���h�U��(�Ŧc�"�:"�
u?�r�' �	t�	e(�CW0��/�E6�ý% �\�w�|�K���	�Yrԓ梼C�%�@�k���΅�?!2��/`P�m���y��r��S������-�@5��\YF�z�u�'��%8g~rX���a�eE� o�cf�����E����b�Bt�HA��B��Z�n4����_5/=�d��{�Wt�X3=|�L LJ�s��Z�,?�N."=�Q8	���MB��ؤ���KX�"�1�M;U�-K�Mp��^��Z�p�ja�Ĺ�*L�~�\�L"a6�	Z5dQ.��V�6��`�",�����p���R�l�B�@(%X�����l�U��(��k�O�
�ouSve��Z��I/�%?+�W˂]�O
F��r�=���G��@W:�=n���9ػ�x��5	`��'b��(O<�؋���>I�NF��k�-�z��d�Jmq�/�[�	��U�Pa�&��cZ�t�Wn��Er"C����)F�,vл}��2��Y��3��bX�,��m;�T��,{�s�j��M���ڨ���IG�R|�y��W	G���}��C���:�i�ϋ���i�'X�J�����L$`�q9i����lV���M���"ߨ�z��a�}��.B��Q�wF��]j0�L��A����/Y�Š	p���Zu.��7�4�v2�j�pƮT��o飓���ߢ�{��ݗot����п,��_�k���L����Bq�y�Vzҫ�����l��3����ո���ߠ_��-�[>��=�����^:���S�I�6�X�CW}/B�!���y#!4�>�o9�K�Q����lh+��n�t�'la~r�G�x�9���B '���,w��{ѕ����B��ZFm��������Qu0:-��,��[D���D��E�O��fDIՃ�Eyv�p'��c���2��s޳a�2�L�͂(��m="d�݈X���c�������6�'O��J%ޛ!-��V�	M>Ygɕv�pz/�=�!�����j� �/M��Wʅ��d�����6^��m��;1�O��Lv��A���I%fkZ[��:�b��}5l�#�@'����A+��H;$πK��&!�0�;�pF�[+$Z���vk�s�ß&��y�Q̸)J������Q��:S��̸�9��w�!�?��0�Z�S��`�x���Y˰ޥi�Pi������^v}�EFjӲ�\���@/��Y)��l����F���a���8��&���I��!ހ����^�!��D�p$����a>������%��P���}�x��)l�l$�暀��P�Tj��Mq2mqv��vN*���6	]��-b��hL�sݥ��V���`���cϜ��a�z��P$��_��bj��Js�T4�B�Ζ!Ci�
(�~�+����q��
�}mx�k�.�G�{kŧF�Eadt��G�=theSB"X������x�Y���qL3kuɂ�	��l�2�,�΅h D-��'�sy�Ia>ޫģ���Bڣ�)�՛&�Эuj�:���v��8ק�3Pۃ��'�����*򷩁	o����>��9]�ۇ�x��1��(N�I&��')���`�]T����%�4{��t"�V�!�x� EU����-=�-�E�ˣ(�[���S���N�{c�i���-���~0q�<��<b�{�^V_�Ӕ��cN�����x��_�RX����ě[�R�H힥�Mh{§`��K�/�(�e�̃�>R����li�DW�+I!>�X�zz Ð�����q�����E~e�	�L�P�.뀱+,�9�{�h}�������mhY���f�N8�)c9SFj˴f�_>^	��iM�:c��#v�mxX���%��]�p9,7��R���&����2=�Эy\`"q���a�VO��]R��5���?֪��ߗ�3,�L(�q�ʼ��ia��]bs`Z�EY��p�J��#K���1��0�L�T�ڮs�����I�U9L̇�K`bs.�.=>���_��H_~��J�xe�$V��p<tu#W��S&;iQm yl�~}��������{xJ�^gb�=G�J�������DnMJq��y�r�Ԉ紑�O؍�h\��r�bSd'�sXۄ�5e�%,��<��o�������N#d�(y�������Ϙ�	D��g��Z���0ġ5UO|7���9U�.�c�M�,��E�����������'��)��3e���]�G�gռ�Q�{�n0���)I&���ˢ*�G��uϭ_]hyC�1���IA��#h�1Pud>���-�`yL�^�-@+����thn�z���&'Q�������+�%�3����ֿ�.$�fD x������Ȋ��j
��2
8��K#G�s�i�Q��dݫ�X���#]𼠦�c.B�J���;����Mg�ۣ�愦�@ĀY�92w��U��mӼ;FS��Y�xZ6�1	�V9��`D��RՇ�em5�����:��u���F]ؠ���gQ��3!����^���a:@�A�Q��%��N��bg��?K�`����N�b)
��+�*��)�dڸ�+
ce��Z���m��Â��^��ÙuB}F�(gi�F�+�(�(|f�y��郎Gq+9�D�`w�l�	saD�����L�������=)'�F����7�,w�Q����K��iF���t;hA���W�c�^}�$}��f�8��P�A(�2"C� wF�m�%>��AK=!H �ϼ�.��f��%h1r ��``HT�+<���K�ݨg��Iݺ[�1�H���Ů/Jk�Uģ���ܨ}i�0,Mj�Xkp����<�����¢�%L�Pֹ�Z�yQ�MB�4�yFh����lUG��dQ�2�%'��h��Q7�/'��`[�䩓�ۘ�`�R�c�B���=f-���k����Ae�����vCYɧ�s��<1j�i
�<ekR�q 7]�$�S����W�q�Y�`�R{����V=�6�OW�ަi��=��[h[���^(�6��JB?�J���-�~��OGAg�F
�8%Үn,o =�[l�۳/�E|�>��L�с��+d�?�K`�E<�gx��2�zv'W�Ʈ@�A�e+�Z��s��BBp���}:!:'d�eIvXR��R�#/�� 4��Jl��zS��������9,�H��YX	������$8�_9��b����2K6���&xSˡ�����؂3�a::��X����d:��k{ք/H�b�@(�� ��a���
����=��'�']mH9�r���g=q����V���+b%��E�4��������p�i�9�4��2�x�M�z5 1�Wg��)����p���џB��_��۪�Y�T�4�c��ȝ��F��?��v�\�;���N���X�0�MMŖ�<�D���z����k���:�_���9|+�LP��*z�Q(��ťw�^9�W��T�`�DCU�ƀעyA��b�>$����.��+�w�-*��s� s��[_��g�|v���ha����������G�7]I;_[ΛaģV����V���Ո�X�X[17��dw!��K�8}��K,YRlU�5�99���F�~�[�=��W���W��5b�a�0�s|�	U5
A�^3+�7�8E�_�;RE\�E6�3��Ls1&���Q�q~���RV�[h�s̓!���nT#֒T�ٲ��ΩN^��,beܡ�������v���tS�#�7��^�FD�A��o�%V#���>�����3uu�9�"��WǑ����&�g����\e,�|R�t��BQ��l��B=c���Z�w=4�����}xb���ҵɥ���N�j�=��f�GF*Z[S��zI��zlH�(�]}�&��;챦�Ǧ�|	�3�6/�2�) ����׺�|@-�7>@wx٨��!JH��L'��K`}��iԏq3�ZC�����Dw�At���U��(�
`��$qɛC��mQ��zC��n��Y {O�O\���;����ѫ0��H262�論���һ�~���M����j!}��	4�R����D���H8'�+��< �M����jM�D�'���L���J��P��Mp6L�D�}�U����y�B���W��t#<8Q�Z�j���]��J���f}K�??q�K:o/߾sۢA��G.����~&�����%�]�8,:�"�̆�t|��z�g���|kS��nסV�b�4ܗ6E��ӻ3Pz��b���>n��<�Td��J������ݨ/�'�`U�jvX�C�3��Q#`>h]N&����,Ev>��L2Q��<���Z��Ѝxk�{s*'m���1Yx
9�F�X�^��o3��x՛v D�Ix��ǅ�{˺�nu3;����z,��(*�޵���k1�X�[H�L��J�K�4 d�c�H%��g��R��(mb1���#b��cq����4t�$�*eu�v8�%�~%��o�]�/�&���7��\as;i��ω�kW����>�&+$��g�ٜ ����P}%I�}K���7��Kyѷ���T�'H^�l �t������@��z��+���Cx)�C��%m��'V-O��
���i�zt3��Ő�ẗ́L>M��Ū��ݼL��� ���W=��?D坱�`n��-i~�M���\���͑��4�EYED2�JJ��@VR���8t#7%7�f"'G�EpLۜ��cq�av���0@�&'���6�)��/T8a+����n<2L���/M�]}�����]������ET)n]�lbs{ߗS�V��@ .�X���d���[�#��~i:�ҏ�ޓJ`ka^�W|� �!L?mlx����%bL��`� ������ฑ�^	�T�~�uZ�mZ�>߈ޕ��}�[�8����E�$C��r�(��,�JS!���- #���k\��{gh?�B��2�fL��V�;^.��1�j-=�����E��6�yL��1'�s�%����(zQ4����P�e;��5a2a �!��Z�|��[Fn\^�<�A�]��ϖJs�y��_p�	jy2��cF#���a�8����ν��8���;-J�'�y��ϗ!N����)��-Ri�L~�qS���������0*R`=]�U2��!0U2��XM$���A����¹#`�VYܳɍu��:-��~�����%)n���1D�0]V�MCo��KN2�v8�zQg��5o�	_n���cu�������hBr[�xI��^��އI������1&������&���=7�P�����Y�6K�]g��懦p���"�P�d�D>*��D%��8�`�ʤ�9�Q�O�8jpk��I2R(q�tA������p߆�(�)(~��&��̎$n�JV`� ���}�C'g&7�أ�	V� �K�W'�����:q�Z��p	�Z����d_��',�4[��_�ߥ��y�5t�dJQ ����鮹;b#��g� ��9B͏WFY�<~���*!��o�*I�����Yy�"fO�cNw/2�|�{��&�e)���5�d�]�X�Q�7����i����[�k�E��JC!(*�� O��d|{��c��~�}�}W��K�[��c0 M���D_��3�V���4%H���7<��*���>ل�j@[F��������x����_ڏv�E�E#�U�y-�����C6��W����&5�G2����׼K��"�t�9��V3��f��m\>�͍��=3[������ͩ����}���+K3�
k���V�t�tJtݔLĜR�g�T�\��`��1����E������i�-�S��@��7���1Z'W���?{��Y��,��@V��ӄD)��t��ڴD�q�e������c�悆��fpt�&�2�P�1Ej�/�(h}SS/O5'��[�S
П	VE�<ϵB�L��7���k������$H�=��+U¤���BD'��;���x[4�x6�u��<7���N�y���,��QǏN)_����Q��`Uy�	h���S���(�l��t�y���I�l>ֆ�z�q�#r�T��f�~�<v�A]��o]���� %�z.�-c�~b�jP��}CO���mZ��(��(*S�6	�2~o���w���BB���y���K�cg��O����?�����Y���� � ���ߩ P+��+�N����x�]�r���@׾G��i?=[�	�u�?�sA|�~˒�K�� \.ֵ8Q΄{�zW���/���=+��9��=�ޙ9L"��:9�Քd��e2�%`es�3�t꼍X�g� t��BoȎ(R�<(�ш���D6�E*ߢmbyאϑ��.4�`Ǿ�y�5��9�bi�p��[�h�%2��)��I�p`N���4�������YY�L$wTu,�h���eA���L�R����N�EM�ڣ�+�ád�����^�����np���-��%��)�=���e?�����;N+�[�g�pMz���F.I��%!�,���R%��f�O=Ə�U��̟�&_?�M��P@��αѹҞ=����b�0���=�����"Tu?��:o�x��Qy�����j�"����X�{��7�^e�y�͎\x��I4������k��R!�Y�~��5�<j����`��`1-(���Q��
��>���z|l����g�Ŗ�����j��_�xA�Y�� �费���/q*Eh��ih/�RU5h��i/N���Xb��ޤzX� ��DO~x�:V����"�������̗qA�#�:�������|�:v!q�b$��|;ʁ<#�K"���|�e�䪖c�Q�b>��'�"��-t2��2P`X-ׯ#�H0>�������8�٬����wz7i\,���;��'�5��(��*��S�̾R�u��;�
Vc~�{�!>����'��H�<[���r�|�����)t\������D)1����Q�P�[xHr,�__;=r�e���{�c��~��_m"�!���j��J1�뿋��M�N�V�����7FH�M�����/�]��]�G�����vE�Q�`<8ރn���cH�>�	ؽ�.u��tOu�����'�-�@�N�]���h��c�n.��^�جBF��GA ��Ź��V�� ��:�w�/��ף.NlZ����u�{E
�6|���6�7O�>�4���
C��9>��a��^���
�+	�S�(8%
��4��W�"��s*w����rV� ��yp-�]�R��~7��9//4�ҿ���=C����}����	�P�_��Ww �<��:���a�Wۇ�mb��T���QMޗ���)q4��Ӭòy�.�����LQ���*H�(�ʓ��Y�(�Z.�E��`d�Zy���2�m�:�����g��l�l�H���l�Al��v�5���N�D@�Xk"�6z���M�'�ּ��Ӆ��,}\�M(C�V�qm�]3+J�ޙ��a@�����<y�e�!�KJP�+����Gf�A[��/��"S"i�E���o3t(r�� s貕���r�%���Y�	y߾IR�4�����������x#1M����I>���w���y�D����j�\��������ki�D�wvvs��#U>�r[ R��ݢ�O��HN���OS�b�0B5��Z9H�C�0��󖧅����w᝴���(v�l)�2b�o��=yw�v�kr?j��c�Q�󒔥�U�R�);yϹ9h�8�>ھ��n+v��Fp�A�>p�t��x����s.�*��UY%�zl�w��48��ͺ��.��&R�G\�g*C��K�zҺ^%� O��%a�:�#�X�s��<��N�N�;�EK��r+��O��x(�C���� ���BqS�G�ֶD�Ž��6X���;�T��H� աm�q��]C����A(Sc6az_9��tEoq���tR|�	�f��2`�ȔC�힟%�idaU��f����	f�v"�#0)ߧ?�T�44��?�6����=/;�@>���o0�h�݋�r���n[t�Y#��E�l
+�	�o^BTL��~#=CM�  �ה}���s4���OM�#���x�ۦt�7\<�dB�l$���֚�:�VK�n�S$A��">f,�L��_�3�[k�uO���h�'<��w);�}C��^9���=O`ۂ���� ��Ö�-NT��u�e�YzZJ���L��r�)y�'.lC��� u�n7�!���g�V,���#��wҙ�8�j�3'fz��ꂋ�k�3�i�������Yl������#���"�/��Kj����z�]��_Y%U�=��[[]����3��]_Ӵ��]'��}H��G���qK2�3G �����ҧ�'�P������c��(ּ#�<��|�|�e�w�68��=��/	��������Q����z�)޾�eA�B�_��
���vܹ�ID��1F� R:r�f�Dċ��d�n"��_	�{F���_W�b��L��Px���i��g�R~��	Bp��O( ˣ9�Q�9�����X��h-�ϐ��F�bT��� ,�����ΕԚ���r�T�:���3�_+�4g�M93E�ǗC��pD-���E�m�A�mM�q����������t�N=�p����L�=O�h@�A��{FM?,���xˍ_�Gס����h<��B�I�lUxu���C{��z��ѐބu�j(��V���Y��~����m��:Z�:�`��]���ұ��4�rxÏ�T2nl1�����Lu=�H�zC�c��1�֐<�¢���&`S�ܠ�p��@U�yq������#�zd�Kø�����v��AK��IǛAùg_y������M�����?/��?ɰ�2
�v%�?��σ�4Eߏ8��ϵK}�Z&��b�*sHn����ףP)� 1aܭ(��g��,V=�4KX�:���m�����&3���aT�fPv�mh�R��U�=��E��@mʭ�Q���:�4(8���i�XADׅAި��\V�jB��[���DA7��ecT7hN|ug[�C���l����.KL
p����k�mc�G�8�,�5����,����NA+��k=��k4A�) ���?R.���W��҇�}����� s6I��(��o���V~�58�@�!}��}'P�'N���2,6�q�)�e�jY-���N������rA�]��M$tH�]���0ܶ3�-~�I�L�k��S`�O�f:Q�Մ|#��#釽��$(��?E��2-ƴf́�L���YܕhS�}Ǣ,�Z����~w��,������9���@;����܃�v̭�+������cI��^UHn�P����1�FM�2k�i��/�b��8��<N.$�T	`��Z!��Rj�í6x�D���.tK�l���Wv��I����B8��?BTUI�[��a��-��Y���MZ	��X�>���&� ?Xl���:\S냌���]��Y���:iVͦ���,i����i�^v��S
Wް� ���ɧT��f��Wյ���5[1/���C=�B�ٟ��_~���ieVF���H��s�T �{(��K����s��Os��x'��Z���i�vߟs 	�؁�y��K��ҳ�[�݃ � F�o���{�Dh�`wO�{��En%�z1�CU=2�#�W�s� *,�h�b+r��_��~�&�D7�{��tb�^�S�ے�2K(�m\��v�i��a���TК�9�{���&��A�$X}1���&���r|��};��Dd�ɋ=��dQBM��Az`I��=����IW��յb�\�}������
ڠ�P�S���<��)�M�1��y5qP�?8��+?0E��;���/ 㔪���L<eT�㡵��x w�3'�L��C(D̚�f��'�7ױ����X����PT���.=����7���t�V�k~g�� �x��!�t��2ޓ��p*i����^Q^v'�5R�V�)8���,L�Jp5�廷�ܾB��F����6�H�p��;��Ȱ�[�ч��Z�=�I�9�����'O�ոt8Շ�s��V��c�q��)4bAK� '.&y$�W�e��ug�c3����݄���J aVjO9�|Τ���P��w��R�����O���M���v���%�����^��(�2{��Ƌ��L���IN�KSӋrZ�P�]��8ar�������{\��Qs�]�.��J�|��;��x������s�b�wc��1�I#E�~�bw¡�8/"�,E�g%�2����n��=��v����_�m�c�Y�A��#��s�R��S��[�14@h�ݑ����A]Ŵ�zC�=�@L$W诔��b��y��J�����ӪtZ�/�.�'������F3��Yi����ɽ��!�?�fm��	(�g��e��s��UVȠ��D3��^R����2!_�Yi�}�݈�6�U)\5?u��Ǔ�wD#���t�5�t�%����S-��_�L�ZP	j�n,���F�4��p�}[�'�-�H9�׬��QAE�B�a����X������7�Z+gyd۠�M�0r��� �o�Tr�S������!Cf�40|��YXQ�|_G*҆�$�Z�R��`���Y4�p�v������9���)��E�Q�5zY�3��=�%�U�HD��u�6a��wy�)����>AݠK��!�I�7����YuH�L�=Y�^�b2��'t!ڵ<c�&�]��R֘bd�8�q©�i0�Q����ɺu�l�/�)/o�L� �C~�Fq�+�+u>�	�y�c^��m�`t����3���H�n�!�^d?sj� �%k+8ۣ���t����8�I�Ss�u�%vU-�?�7<�E<4���f|,�ak����F�[g��M��ǲ�&*�J��D�xR�)��VQo��OV�NF߻�;[��?��Aɣ��!x�A�~�j��v�V��ٺ�#j��$�<`�WJJB�nP��^1�hWͨ���-�;}�nB2�A$-�2�<]
UM!`U������#���ʴ;�#O�,�7$���{����Ԫ����I�K��~s�!7ÿ�:DX;�3��I��_+Ͽ���QH�yG�rO�"$���!`��ZmE��G3K�Gr�����U�o��Ǟc�hzz��|�Rɋ
~�˺yN)�TKx�
���c��ӧ� {<�F��;ҙ����k�FR���i�`탓p�'~��m����,�9�1)3)�t�׃NO}����I��/�s�W������NAWK��D��`��3R�,Z�ͣA@a����@m��=ڵY}z��J�+*����<ڎy����<�(����>���B&dv[>�?~~���oB���SW��H{�߭-K-�6��:E$�c�)�H*B��ӯmp��IK({rh9;���<��O��6q��XF&ֽ�4�r>ԉu��C}+C++R�s|]f�2;(��qv�[ѳ�+��wS�^�E��=�
')_��8�7epwx�Lyo}ru���z2�o11w�鞩xl�QS��k�WO�8n>9���0��k�O�[�{���[f�:��,U����R��o���rtXe�^��ĮQ/����� ���}�B��;�A��	O����u����WT�/C
 ���0�H�8*,�I �^R1&~��k�a��U^ޛE����CA��qx)aG.̮1PZUc��G��Μ�⿥|��w��:^�RD�zK}j�1�GW�x:䨢�$��#~����)Iv{5S=xW�u�}c���!	����z�"��c�ƙ�������ԟ�G�����$�P� nH���g�x&o y�g&����Շ�)z8�IQ��+o�3��D>�mh���ܵ���E�CJ�Y�FQ�$(��s.�5�OF��^z_��D���i���J�r+`
L�s�����"/wV�	��� ����H�b��'�b�/WK!�\��7	M!7���Nn�ט��1�a�|GhD�X w�}L-��J����BRd��׳�p?�0��n֑Ț�7�]�o��[�r[��2�qL�&A��x>"��L��E��[�v��>���
�1`�g�o�̑���j{�ąT�ɖ��Ȉz��Cz�|m�4��!��\�*�c;�ݹ�l�!�������ֱ�8�L�y�S×��P
{�{n�kګЬ��JOQ�Ų�%��;�fij1��$M����gOrH��Ϊ��>�z�Y��zu���Rx�/(0tͯ.�Go��|�#��I�p��rfw��0B��kSɐAD�/o�zS�|���K^S��濒S�1��m����=���J�������A����j8�_��5>E9;���v;�ї��A�.�r[��Z>�V���eo���_�m"��ߍ��y�
���z� �r%��㔛� �z�:n�ST�^�3�FG��y\>�J.���8�\���9��pL��=���!�nw�63�t�v{Y9	��%Z`�m�<�=,t�����M�1���p(�M2��@���f{gQ��!���)-??�N{�VՔ��x��ޑ�=W�����{(������U���k!��l��A7`U�ȐN&��I�t�p%o�%��EtѼή�^�Jz~>6Ԏ�{�P�9@r�y��4�"�/�lr>ǌ	�l��Rq��Y��<Sí-h���e�<���O��8���>�����sK�C���)n�T#��~�I{�.���6��
���w�%u�ЧJE��f�u]�F1;Y�=�|ʇ�U�!�*�
�Dg��3Φ��*`{,]��7�^�XB�*]�'��>zpO!0��j�����a��8b
��<\<zX�G/�F�3�/>2��@�����Y�{Δ��{6V{�[���ͅ�E����yYu x�x����/��&��V����/3�x��B�7o�F�r}
�l�%x���ɭ1��:�/�� �^mA1��ͽnq*Cf9�x:9|+��qX4�_HՇ;�4��u\�+�p�����#m+٣�Y�宀Ѹ��Z�Ę����8�h��WY��|�4��U�e��M���S�o#� ��z�Mb�S�!��vY�"���o��C̜[X ~��t�[�����c�,m_uā���C/.�̄�N�><��A��v"��Σ���r���`�q7u0����K�+�$�5R�T-�X�����l�*eݓ*�N�h��Њ��M|�/u�=��/�ٖ]Bվ��'�.`�&:�!jW� �6�7;������� ��]�.o{j�p�����p4�>�6�E�I����0��I�]l!~1�Ö�\57�H��� 6-���&K�k���-�SP^Q�i���N����\�K���o�&������f;����p�X�
P�!�ݦ�ג�� N>N���9:S�+� 6.��J��r���Js��A�]�
߮7	�w`!Z��8�'{����/��(wenL��5�q��(�����z �Dg���5c+�/�v����1�C~K��gԺ�9�n咠 �J�&�h�ݱ�H���V��ـ� 䔀,�,G k=�}ŭ�>����T�h=mV2G&������,v��*��)B�]�eU�pNR ��^Z����Ù���\A�v��H	��~��9��EC?�Z�i?#	��h�jU�����f�t�Y^�26�e)W]0�#!��X����9�5��虏�>@t�\X��xe��&��8r�p�Œr�R���T��~,;	��C��z�N�o�K^�3s��8[�kGn�{�F5�����>l9-���~*=Ļ,c�{�8�!+��'�`¸�=>���%D s}</�G��a<��Plq�l�bf�B+/�V�/�?�S�qq[��r�����O6��э:Se�sFX
����%h9�E��)s3�?J�,�W���7�Q,g�"(���J��9y�v7�L {,1��G�����/�]5Q��l���X�=��]���$�M��ם�G����@\2)Ϻ$��N�~��Rt,�(��rrx8��	���}��=�shu��m}�Vg��s%Nʱi-��S5j�@ýelkv�k�^�!<{n�����1�z�-f�O���*�eʺ��n#|�ju.l���6�j�!RC���7uw�����o������!l���
�G%Q��ð�.�;}3��OCKc�(Q5�#�p�+���-�@w������a<}�	}�@�k�++�d�A|M�W�C�j)��ñ��Y���e��~C"�E��|y�9�]_o�0i�����H�(b0p ��W�N�d��B83|QH 5֫�(�-*�k!�� ���W�H����Ue����.Y�Vf� � j�x��[�\���׏�����^~���n!�6E�ױz[h��+�Yۥ����j��Uo��q�����=V?�t`�{^�k>��`�A��:��T/�֌#,�1|kw�a�=&���Y��h �o���C{ ���3xZ�2S��|�K����|�4�A1�.��4"�~ϵ�����sĦ��z]"%��Ȓ�
!l\��bɗ�+VS֕#/c
��W܍��K�����O(�_���՘c}y9@���4b@��/��0~@�lE(��ᵄ�Uz��a��-�Q��б����<royĒ5_��2bSL1�[�m��sm��|4�*�Pؤ��W��j>Qx���c���^�Fu�
�~<�g'��x��}\���@�`�u�$ԙ��S�u�����[�Ȫ��f�Bn�+����O���S�I���߯�0�@�Ha𬉵���7l�v�hi_M H'� �^�cUP��#v	�N�t�u樆l܈��4:\��a1���߿���vk:�ju��?u�6�6���U�SWc�xXR�M�jz%�Y
�S+ӥ�f&cx�B_�p��fw`B�ְ��`�qP���d �S��ߟ�\ou��)��jTT�٫��=2�[�Y��
E�e��Z%8��C��;��MG;%F�i�	��������*뚾-�Dp(K;g$�wY���%��X�'�B[��3���Cxb�~c\��I:]������1V�H�L=]���m"��Xq�~��)�4'�	���sA�$�[�Ǳ�p�O�^(�����̞���*w)FΊ�G� ���2���z���z�ԅg�%�Kd�\������dL��������(�0]j���f��u/�t��MS���:4�`MQ�)ЂB�	M��0$U#���M��loO85��s�|3v�R F�-5�h5����M�����F�d�D�}	L�7H�u���'��49;�5�E(�6�����˗�*���qŔ�*��)�^��Z�O�z*�J%�Aɑ���2��2У�kW�Z���T��oN�����C��0��D2�-Y�7��]$8f��敲�
1c����!c�������A@�0��N�c�b�&mpx��	!�T> h���Y�psfo6��3��ya�b�p��|ڍ��+J�ThH��;�(��+:�M��!x�1��đYCK/�Ȓ���fee�qH�dmF%��F�c�i���s�q&�e�Y<���r�QӜ��n嘓��
>�d��;LP�(U��Y˥�UP���	���K� [�!��(��v�l�$Gko"��20h���
�u�xS��qw�R��=++�Q����̊�s�ygR��W-x:|�2ҿ_z-�����ˡ9�{�4�>�Δ���&˜+��U��,�G���J���}����(�p��ɹ���˪��2����?r�f\=��!��U.ر���b�1��t����񘴻S�{�l�Z�bS6h�л��I-��t	*c|�v�)�X(P�W�f�ΞK���Ғ0.�����y�?�y�0ZS|i~���Yj��7��1�ہY�g��yo��}�O �no�n���*%g��FI�~�fOOl�XrD�j��4�-�0�A\�Y��"Ӫ���P����B�xe��[k(����G���KCOxY$�A�?ЁE�C�������;���_����!I�^�C}3�M�Ӽ(�D:��W�KQ�h�웨7�(�� �`�
JHԌ#�+��h}����u*&	�kc�����<%�4y�����,bL�:Sl`�@X㠙5]E}8s��9!J{��6Ɉ$؉Zykr���r���)��֓�5S�"����[ԛu��kߛ��%-�M�*�rm��-n�a]�t,E�u��ڊ����Zĳ��ZO�q��=����eS>4\��&�p 5'rO�%\{S�S"��;�Sv��$4èU	��%�;䩗o:�&�7;�J���s=:|���=	%q$��C~���όuۤ��^�~ߑ����6�B�.ow���8OT��Mc�7�d���U�S\ ��!؏c܌P�������n	�����s��f7�2?��Ԥ5EB��X��C�!wܭ��
~�u1&�)M�IO���� A^%d	�}��)Ơ=A�B՛q*��>p�M�j�KF�i���h�e��ʊ���oV��B���Ȍ��=v�س�/�[�1�������? ���G�Cy�җ�S*������NU��A�F������M������Kr��v�'�d>�!�9�i���<��i@:4�b��'����b���������-���xHշz��V�ᐳ�(�Ƿ�����q8&�m��+H�s�<E�f&x![i�c\z����C��f��Df��7��>���\�Rc㽷�D����(�-�a�pusW|n�_
���y��P	���v��H/_�C�_~s6'�-b���Zc�V-٨�t'�)9ŭ���=L�����)s���,��֛<*)7�<L����������T`��*�/c]����}V. ��wC't5�\�dTd #̐���Ut��8�Æed�e�P��Y|��'$���;�0�?�?�������|*�W��v���+�L��h����� �z��$����xNj�[��C�{��j:=���ݖ~X�F�t��u^�2Xv�
Ok���]4PL��d
9MAT����ʑM�u�Bt:�Y9���L/�����!;�:V!c�U��X�g����K�7�6�΀�z8
��w`�Ը6e��"~�Z8}�ѭ�+��n��0>s�(k�opYA��
=�u��́#���q[��-��G.v_���q<f���*���cn�ۛ���F�����C��e�D3K�2�mY:`�	5��tGx"D�ֆi�'��FE�W>����2�1��D�vj`J�]ۆR�x�[9[B�;V�!Q{S*�\���Z]Sf=���o�����G�vL}�]�Hwk[gȅN�bwH�eN�B��m!�&�I �Ի����3�4���Z�iPŻ�����\����v*�jJ�ǟ}�?S ��x�ꮓ�"L�{ECL�o�!|�9���P�9w���o@!���prR��}�`���e�ǒ�����V/V�V�v<�*Sݴ���u$�(��܋���a�'�_�ig�l���\�cϒ�������|e��X�S�zP�o]��C� ���G��̐�r�O�꽚eD5���֨/����&rf{3�O�Ih���M��Rυ��@ �%�H�jo���:w�l��~5��_�rU�)�r~����������(v���R��݁K�	Ȯ�2
��#GU�7{��'��2�tv����{�F,>�Y���w��1��1%�[�欶��d��?e �N�	�֦ �9��t8��o��[n,a~ƙ�e��~�@5!����%�Eʎ:CH�V�&�ZY<&O��Ү��Ta�a���8���Eb^�]7vҘ��0t��R�&j؎��G�~��9��$���r�gC��bU���k���*���Q���A�s("$r�wf���g*g�=2tw,��e�/[tOTIS�-,
�	5�8�|��Sd�^*���H��S1L$�7��U�Lv�>{���N�M���J�Lr��8����uu/,F��yt� �����#SDU�ܐ�"���Y'P-F�ke�Io�"����(p%��omE9w��$39y2��_r��_0j�~�XnPa��uc2>7�X!�a2_��پc6f}l�Y�����7Iw[�>,4=X����S݌�����R����D�ߓ�#2���*}�������^Dץ�_[y�G0sI�{RɯsR��$N^���Kz�(ڎ߭�U���D��[�˸��B���wRygF�eu��H�i��u����ī���S�V�F����.�[�7I��熍V�`:�1@��qh���󕄭�����}����+E��'�|�'��Z�����<�Yg9=*
Ϟ�����[H=Kw?4�7��7�R�ע#��FY@�ç-�~����	+�5C>��;�����c��V������V��1�кWj����Q���t���Y�tʢo��8O|iɈi�85&��ǃ���M�)���y+(��o��ɔլ�����ێA)џE�>b��yb[џ?��D�Rk�k�HY�ǩɪ��>� �#U��]��,�����(�
�w�$R�`L-���0��3Հz �r�7HjH�
�q�0��4��R8Xp�u������Ӄ�Hz�L"����ŜGE��;�����ib %q\���%�nGV5s�����oo�o��Ŀ0/�@0iY}O�	-j_�"2�Q_����I?%ݏ[\
Z����LnoY�~G�(��g�:$Bk]J\�)[�"�y��dυexI��=�Y%�=vL�HU�����[��J��,��c��ł����A�Z���$��L"������	�\� L'Y��^Q�hT�Z�^��� ��oM�����@��'8+��$E�e&F�����^{DV�@�D"�B=InW��چs�2��B� y8p���Wfe5���:�����Nc��`�Uڮ�U�L%"_[�ڬ@.0�G�p�&�4����j�C��� ���P#"�_l~��h��QTӄ<u���J�_R�s���~t�mQ"��q�ȟ޻�g9��Au�0��"�-�I���0��kP�9�~� �+�׳���[� ���ŀ}HS����$@���"�@���\d�N3f��~ó�7X�t����>R{���3�޺*�T/zO�)������8���-���żY���P���i���,>���WUh�8L�0V��˜*
�.�.y!r�LE'z��� fR�(+T���M���]zE�儬�Õ2�\����Rl[�bn����"��</JM�{���Y��:'�0�w�^����b�|������y��dM�1��<Ho���
΂���i�o�®7Q��N%����ڬ���O����nࣟ&8���[V��ry���y��툋LK�Q>$zl�%ŅJ��su)-��K�+d�,;gڧ�ߞ{.�yw'D��М����a0:xʉ��.�$���0]�g��C34��U�o�
��ᒨzfmW�u�`)|�%P�d��^0���^��Lo�%��t�䘸�����(-C		.k��sk-�2�D��h���f���������u�u�UƿՄ�t�:�����m:�E� ��D{7W�磈��c��Q����|l��]���1,�7�K��oA����	M��fr>��$��#=�5u_H�ˆ4�gQPχ� �E#
F�j}+��#�����-dO�`WhO�'
��-�N����|Ӄg�J�#:��^"��1*Н�bu�3ܜN���0�$T�%���5��� '�s���1A[��������N�K��U�2� �iW��
	yJ��tx�b�L(���m�"z�T���cPX�dy�O��ۿ�BC}x�C�4�F(Y"��ehH��Z�~�*u�>@�\��E�FS�#��.�ܕ�s���������֢��`g�� �Rb 1�
f�v ?>��~���� �!P6�ϔ��M�#t���������"j�k|�(�^��r�S���M3�G�6/�9�?�zKv�6wVS3^���q�~�g����r�;wK�^~H�D�U6�������(Ԕ�Yv�.�b6T{����&"\��!?bΒ��`�R��;e0��b�--�������+�|���#�/J汋h(V�=u����!�	�Q�}jLv.t�|ǲ"䮈��SS0qî����zi~Lm�+Z�ɤ�W�4�,7g�0��[+(T�*�Vi��M��w���@K��L���;�l+u�>�i�r���e[1�L���~a�9�|x3'و�v��&$B���X+�	Gt�6�A?��VR�&9*��E���pt�#au�?0��1���l�"s(�5��*���wT���M�4�RE�p;��h�X�u���s �-E���s��9)W�#̂~�M��B�^�.���ѻ�O���K#$m��+c�e�K��}�j���S��V��v�R��@7"p�p�Ff �(�g�e�N3��y�AG�!k�[�XX�0�Q��sD�� oT��~�|Jl�2��{�wp���0�d+�҈�ڭ�A�vU�F~�Y\�T��-�u�-kj����ns+qAZ@�e�������'��}�S�_�30z�|�R�e�}���6��}B{I�ԅ@Q�Mb��3�i�tu�R�w,��z�+ivB^dak�@�y'���Ǽ��(7� �v51�#^BR{>5´� ��p�2�V`!`�(C�ᤓξn��2U��P���#R��S��V1��V�����"���0)��q|��4�ΦuhH��ZqgS;+�U[���U����(U��_�|2D,��W��'_"������;��2���LSd���Ԯ��-�{�j����n��NC\^��q��D4��œد֘�xio5�T0ע�\�h,r���B�߲���AWo���� -����={�f���P9���"/";O��t�oVsϩ��# ���+n�D�䩑f$t#&=�����W�/�`r4�+ ��:R�.'�$N��M��Z�<�����
Pק�xc�^JˆCx���/|@Cҹ-�[�'5�nP�!��u�u���R��E(t*ב6c|Dd�d{+�в�N�-&�5ǵ]�j���"����ʰ2Oh�N���cٳ��(�Y4�Y9�l�oĂd;��_�ʀɗ�C&����A�a�*��8M� �Ц���F�\1M���Rə�mk̬��9���[���e��/D�RU�݆����)��������[*��%1-���Y-V}n�ɣ|er�?���A0/v7��ߘ�JjG"��z3!�[7zP�x-��q�r���M0��u�\�#����?-��F�ݔ-#.�O*Η�68�,N��s��}!�|���E������Mh�[%��g/�*`�qlS�8u��6F(�����v�����)�,q4m�d)�+�����F��ħr�����^M39/x���xѷ���A��Mٳ�G�w��ة"oU��F������R<^�r�'�b\ĞL.���,*��ʫ�,����::��.� �E֍.(�(TP��7��K1j����4�Q�ԧW��Kz�.e������(e*�tB�{Y��F��`�ZrUQ&DH�{!WϞ�=�}��SWR�K��e���Ro䅝�L��P�����L���^U!�NbL��-�O#�k�IF��¸���i� ��}�ܤ�Y妬�&�M�Ge"�qxr�<�ƨ}���j�w�$P�Z`�	�,��K����<kA��Vj��d��D�ş��+J`��G��`$#�&�Պ!�n�ܕ?��n��eo�`U �-��Jvӆeh�-c�׫ͳ�[�t����]K�(>�@�A���]vb��z^�%36��c�=,�,���&	~�W�5/9��JW���8~Z^+�[V��j�%�B�/���QDm����~WU�i�̜q,���o>*���^���P�9��E����r���m�����5:�AVW��dt=�Ae�>W�l�*��+iã Ax��xh�^���?�\%?2�R.u_zhǞ��y���D�?�{D�/_�����C���J|�>}/�t����ϒnܪ��b9#m*aE���K��%����R\��(���-ߺ2>?�6��}e�qw]Cm]>X����ѭ���5�2��?�'�2��_1 ���䯂fһ������W�d��U�a\i�%r�OTl]�i����ZM� ��Zb�Z@r�MBj���R}@�++�c�����
;(�\-�?j�0F���L��x�0�.^�>�a���3�q\j�t��!��(Q%	�OΣ����}������v�caEjO%���Q�����QJ,Q��6B���ħ� h�r�a^�d��t���2v���� +�ŽHCTi��g�X���p�����d��O0Ot�6��f6�F�J`���r�ĺu�	��V�A��4Z{�7\3ܤ�7�&�O�$�:�M�$�؛r_ר�>�o/&���P?J��ω֗Į>Fņ�Ք6�PI+�J>HJ��$�z�ք����=|�!l�Ԝ�0����j�`���7������þ굗pfS�B��y\�F��������SA�lEdK�I��(!S�����QQ��&�Y��t������c3_��R���A���������������Ϸ�[��E���_��]Rp8�����SҜ6��C��tT"�ٻ{����B'�))��_������z���b(��ݛ۔2^�PJ�S|�zk��_�9��i��~�M��[�\G����z�w[@%a����a>�N"�0���<�jJ��f���F��t��jL�R���<_7	t�~��-�y+HI�5h"�P|��Ls���!m~��=���,���4�*c󿢉�`��j9I�^��&Jҙ9tF��TB��'�>RB5����|�H]c�NxV�̓�s{@X����2���qҕ�>�RPҩ�f%}�sv@�2u0���9&V�\��0)�o���Bq�JO�k�<ҤW���l-��)[�h�^����KY﹦��X6��3�90n���/t�\��$�wnd�<El��z=V��	����������Y<W�F�HvAP��T��ݤ�����5J��f�➇>0$ܘ�V3��z#�f���'�;�:���7`؎�Oʹs80R�Q�`"BQ�Hw�bp���^�@��@'���U3�y{���0��`b2
��@e�4��U!�^�Q�71��E�&[Lo�<�׬�Cr[r{���y�rVL-��'y�߯%y#�&HVx�[n�c[�u?a�~F�dA4�M0�4��-�Y�	Ώ�:nA=��M� ~M��R4�_��r�~�F��>WXڐ?�I�ܗ��Rהz��k�	�F���v�;sK ��	{)�#ң���M�����@g�
p�L̶	�?��)���-�,�����͒�1�M�����s�� o[E	�qھ��r�	U��?C���'i���54/��w���9N�%�4���䦹M��V�f7]�Dc��]�R|��#4�'����O�}W��1y=s(�O��^2�I���ϓ��]���X̷��I�n	u'�@qM�@w��~�m�US��=���6?���i([;�-����h�H`����o( gp�*ŁGR7-���|��G�f8��ƣʗ�Rpl��]FG��)��L�Hjb�N-̑������z�#����j�˖`#�f�(+�hsF���ı]������W��4!��K��ø��:��V��m�l�)�A��&�v���o�	��?�ȳ4��6��E��2�¶���N 8A������sS7C���Ysi�9D�Z�����7�²�4�4���H�{�[�ډ�D	_��6�JNƊ���\��]�ZX��\7����[[b������3��-�N�]�ߧ��56p��mКP�Čs��miP�)�$����\z� ]��zߓܭ^)����Lc���JM��(����Ԩ%��!˛aZ�}�r��q�:�����	(��YW�*,� ��	(�x�Ox| :�5������n&f�Vb�7�J�h��k/{N�%T0Y�u����a3Ÿ��#Z�<�A��+:�IC�J{ϵ4���Y�N!QI�׻�wcc��6��{u2�\t�"�5��Yv2��p��}P����$��6ф"�'�Pp�3�%�l7~ٻ����-����G��)�e�1��f�����p$^&�c���ׂ��#��!�������=KW����F�g�{!��g���`}�4C�DD�^oq��'Z���x��CؤH{�ʌOʕ����N�+2�Q���'L��q�YQ��w"�(f*�t�(�I���r���t�X��&
c!4�9�C�a�"�K�#�G�a6�6ŸP�r�)l���h�7oVN�\O��\�\�vpW)��LFƗ���/��z��F�zq�R�0p}7j����l�+,[.p`Q�@����h��mo�>b���{�S������[c�'UP|���V�&{|�>�a�������sA��uL��e� )��ڑE��=�1<vkq��Z`mjǧ���.�Ʈ7���#G����zD���>���w)g����a���f�q����I)��{ޠ���}?"h�����i��I�u�;*]���&�;�i�IA�
���ئ�������
��{��}޿:���p�WѿD�EpQ<�+���V�S]kK��9Թ�m�����t60磦C[CY"��@nn�e�������}K��!��Q�GpA�4�u[���g����wͩc�"
;�f��delޔ�]��i�����4���³%�gZ���uB���&��dzB�ʙUj4澮_�����H���������}(��`p�nq�@�L��h�V�N�72,#�y5�%P�{�خ� �	xQw�c�(��T^u�F���!=���DS����usTL���	��]��'��1�������cE��a-g�.�ՙ՞_<ǟ��$ޤ�/v�/+�1tW
؝cu5�@�FJ���r��h�r������{mMg:h�� t�ekR�^�����ŝ/��1�^9b�4��.�D�lF���C�Y�@�Gt�����(z��J8i����h�˵�)(̒P`FlX�MҲ�.�6wA��0�^qE߬{�]!|��.)�
6@;B���?.��]�?��|f����w4�Ƀ��/�`��հ�@n�Âf�b�L��E�ǊH{w釺��zGH��Mq�/�mk�h/߯�#0��6��w
�=���*F�gG{6�Mkk�!-DGJ"9)Sddϼ��ZMƯhg,�����!I���5O��0�+fZ�q��ݩ$t�
_��}��-�e��Z��u<7�:/�����	�e�����h2[@�ٚq��)�(.LM��ۚͧT�,�բ�Z	ǿp���(A���-�Ei�H��=;����ݥ������ȸ�1W�ba�J� �x���VT���������q�7[�5��H�j�N��?�9�!��2��n���.K����k]�חٝ��/��ލ��%����wŰ�B�j��0.��\1L�&�b�{[1�^
����Y=d�O���w�
jD�l9n>��kzϋ8��B^KU��
z��R���x�XZ��ME��E&`�fĘ`����#���Q��St��6Yfѡ��:�9z��X��(�Ǽ������b�� �7�X��g%���eq��k`Ι<���Y�P�,�۶�O�А��kU���hP�}{e�O�6�0\{�LVL�fV��bp_�Jp���S��Lx� ��a_�"��Gz�w�9]��Rf:�Y���v4J`:�~W��.�^�#��	H�j�`TH�*ʣ��e����5^p��7U�}Hcd��+8^�n�˸/�S�S��Y����'t��1k� �=�PP�W�|֎��&qM16Ύ*����H]R�4���RO�r��ħ[��w�і�A�Tl��;���C��b04�t;K��l�Y`�I��{"v������-��6��j�YG��(���/8����
�{4WH�r�A��2eR�(��c0>u(p�F(�c���a+0�����Ԫ����-t� �O�%�G�":�Cm�,<	���O�O=�:Ra��`����(I/��b�Q[z��^��K�^���=^�ː���iA����sP]��XG���~6%E�ח�sV��UC��!�o�@�3������}V-��t��N������©Ǩ �L6��e���1 <T��P��	��8�r��>�ӆm���y���䱰;lW���,mô:[�>��-�ךXe����2����Ar��=֡��p�	�>Ԁg:YR<Q�G��+�zùA΁X��6v4u�*�/K�5�K�cx����xd�^Zh��c�膝}�O�q�A[��z�㲵L3����F�3H��	@C`z�4�ʃ�l0����XI�����ۯ�\P4آ�i����Qb�f�L�Vbt��A�[��9]���u�̥դl*����A��^>��$�Pg @���>F��1�HD�yu��v���� ?�ŽўL���V=��F�5����V��p6<NiO�;~_����+���,�Bd2�m-��,v%V I�s���:��j0FT��P�_�@��G���B��a*
������PnV>|!IH�c_r~e�V�T��Ĳbw� yh�����9"�)�a���}��ڳ���S����ٍ���nQ$�AstͲG�o��@
,Q�î�� ���3��}�y-_^Z��h7S
�\�;)r�"�����6�i�,�A��5Ӿ�FR�}����l*LQ�G|A'��a��b�N���E��~��С�;����*�~�#��Dܣ��X���3y�o��=f;�'�~��6�|�Z�-l<�Xbr��s�ב5Z`v�R`Q���-�.&p� t�p�t;.�PY���#�me��?w���54+ԣe�~{*�䡭�c#/���C=�$��e�̞3��`�RlP�5cT=B�3�'bi��;*=�L�:���u�[�s�E9�Fg��0��ðpCm�� �ru͏�!��M��H KmXT���Y/�)O�K�k�Lf�{��7L�nB>&1��eq��j����%ؗ�*��"'������|!�T��r�����Fb���n\���|�?-���!zf�A��F����zL��+}�έ�1�7<(yڨX.��2F���wʜxﯠ�G���FYyI<-<�#v?.sK����P��$kS�A���Z��w�R��:�ن.�� ���9��,rĮ���J.��.� ���}���q�Q2�?�vۡI���V�g1X�����Aj�9q�iS&�L� �xe�5& ��:I(�9�8QfWT��@w�������A�|f ~ϊ?�S Q)&�uf����^Û����eܛ+\��k+G\{Um������}�`��m�4u����@q��V
�|Ill�
\�2f��G/12E�-z*o$����<`V�( 
�s�o��.�=�9�5z ��"���A-lJju�����SkL���B�	s@��z�UϤ��S95G� W���o|��m#�'pGh\%B�o��=���r�nK�Fe2�"0��`n����
����]�lv������wү��u���������:Ә���I&�j��@���2�����kX���,�zr*tdep�-���c�co�eo�L��ƁM��,_�3��������s�Dw��rE��M��"#��>wZc����t�[]���5�F��r*ې�����(Z�j�lN$��Nn �[�$�!�f�}j��>ē��}:ԵQH%���c���7�j���7�L?���\��TL�a?E	4-��_!m*�I�Y����@PB��{����ga��t^��\$�M,�	J���7@���C���I3��b�U����P"jgm�*�ǽI-2T�Kv�	
p��&����@�s���@*��s5A*K/��,�y;��j�@v��k�ma$����X�;k�l��������d��d�7�JPV��#�I��V޹vJuPQ��uư��K�������a��4j�lS�["1�Х?�C��)5�#K�03@�Ɋ��$R��R��~���<Jt��� �$��W;v9��ά�]��K�}@0��[���>|��!���W-�]i��ƾ��o�jH�$>�PP���DSDV���������P}F��pߨ*��?������N)�������L�CߌCo+��Îg���L����m>��}�-�&-y�
�X��s�����r{�U��ᥑ�F�T�e�H�H� ���ԝ��6QES�3�����y��d���B_cm��-�NH�*)n���x����4j�z���歼c���R�U�j=���_�fe8�0����L�����B٪����Mș�m(Ԟ��H&Y3�I"�ʠ�(��l���}�������ٴ�b���CB<��2���<�M�����i �1U�"P�Ƀ��BĻ�m��q:�-̍��ɺ�d�c�
�ȵ}ʪ����+0+��j���(ge��>�Q���O:�h��J�=a�]YS���l�rC�y�@8�ŵ;���yH5'��
i�{.M���Ԣ�q>,
���l��$�E�%�;��I�:$��Xo�D�DC�PB���j��x}	��q�u���T�ܒ��#�[��I�L3LuP�Y Y��£����� �e o�5�<0!8���N���[�`0�?���K�*K���"���t'���8��Hm���[V�����7��U`ݫV""X�v.�S��_�8P���opV��l��6 c��kqկ:Π��˚��02������L���;]M %���˪� �SN�(���t���s�t�dY�>��Ï1!
�!�z�����޾�7{��2U�V��=�G���>6	R����G%P}\��d`uj����ܟS  ��uF�����4�P�!K�cˌ���\nV�V�d�.9x��Q�̍�P7%�\�<��|e��]�yl����l�QM��3P���I��ў�!9���V(��jf8�
O���2����
�?!��?(�^!��D ���ш����\{���?��4�f����s4>����>A1�Ӷ�@��Hr����֋���}�a�Ah��Eb�=�S�⚶��ԙ̚���1}B�BPw�I��4u�>�����bd0i�O�}�z��ͰD��:
�آ���ݸvj?����p��;��(Lk]�V��)�df!D�+"̛�U]i:�0u��;;1�n`�Z������	R%hS\��'�1!TU��d�e�LI�1E����f_.��^?��; ������g�m�Y0��a>���#-����"v���(�o�1	��`�&3�5��(�>�_ �̋�(��G � ���Nr!?�oM��Ǩ�Z*���c��t�H*c�x�������_�½#�����OotHx�zf*���z���B���"�xJ�Q�c�C���j�K��!,)oWC�x(��T���C�v�0{R9�Y*W�	������z�l��W��p,nl���Z���f�nv��]zvc15Ȁh����r��R����M��3qU�'�� �aiq���1�B�:�؇;(��S$=�2�j7���#c�y߀�T�c3�t=���c���H��.oZ�P����B�gj�B	t�����ű��rh�! #Ԯy*.�
�j���������yE�ppbC��o��:�v�۬���!����Q��0W�O*����3F��Zs�O�JP>��:E������+�PKB�e���~�WX붤D�#�ш���?�jV�{%|��8y�� 
r"�%��P6c��z�z��e���v`=@�vSY'����Rp���8�83�$�ecƍæ��!li�o�����T=d���v���'��Bgdo�f�u�g�*�v�Κ���FY��|| �>�L�;�!j�%�Ϧ���)�!k|ށ���⽂̳2�P���O�Ƽz��fp�E��gj;��� [ ��H˱LF��>�)�dg�����y�����|�?ѐ(u��ų /#��]�Cg��$���j����� �-�%���E�"���`yvY`�a,Aj��G� ��)'�l�k�8�ȣ���w���j��i��A;�^ZK(����ka��
Z��ڸ��CT{�4A����5;ʎ���%�ě�d�������G�1���c$����xm7�i����$��K�O�^����.��<�2j�;E �A!*]%���]�rJ���������k�����´,B��hAe<���Q]2�8����$�`$�)4���D�K�4W%J ��M�:�h�kR�0�Z�a3�r�����p��{;�����&���(�A����=�Q��M��9��@Uz�b��ޤÕ�� f&�3,{�T"H����'���e/L���Ş?ʔk�Cj�&	.�jD�L�P���ͪ��s�`�qWN�3���������L�|�]y�S�����1!p��7�v�S�1�cѐч4@����[��D�A���e����O��
�OKnB�Ħ!��'L+Y�9ܤ�t��q��g�^�;�2��G����Q�es��[B��U����T��*.֎#Me�)�V�8���Aq��Я��L!�I���ǙB%xL1 B��%�{�L^?(ʭ�� �h�K��_F���K�X�]k]�l�S��[�Y�1d����v��+�Fu�HU���UZO��&�U��aA���E� Q�sI�&��P48�ү>���	EJe8�""�(@5�jp����C���~�[k�2t�zJ�%�w3S;��Z�n<"3P�)xrԚ����d�5%��"cTm����Q�<̿RȟB�L�����|��D)����N
6 �"�J�C+�Q��C���V���v�I^R�hV/�2��@fMi��fn�d�pG�y�\0ӈ�h�!�ǩ�:My~���՗���t=�5ڋ��Q�?#�w�хhNc����2]��,�ҕ\h��)1��!'�y@M�9���� :���c-����\���,�p���۰f��e߿��Ly]t�BRK]R�X���#�Ã��-����y��4q�6���?�.g����WXx6'�~���Zv�mv�����뒦�o��Bkz�`
.Я3ƹ3N�<� �`L�9 ��cS��ƣ��oa �n%�,���'v�L���Gey�����D���b�G>o@2I�`���W�$��a`�ND�O�KHw��	FW/�c�	���;�vR���#�}����'a�Nz	�xW��׾�q1�Nn#Pa��\�G{X�� �\�U�ڧ./m��v[ٶ"޾Ƚ��{ރ_�ΙV�q��O�A���r���5�Ew6Wu��$��p0�Wjډ�0��yߋ��X�u-�G��%�J����M�D�j�Q�4D�5�`X��3]@Uօ��V
��t�l�M�{�V�t$n	��J�OWU�^*ܷ��j���h�%��pFV�>����!{���`w�N?7NI57��pr�M���N|�u�OФ������S:ߺ�)�V��y��:Ly���yJ��mw��@Qc��1���f[�@)3�n��S����ee�C��흿F�uikZ�%F�o��I�Z����ۢit;��!���[ؐ�2��4����ͤӻ����v$��K�zqˁ�����4^o������$�n�� �Ht������S�{urĪ�tW!��]����;�5zvM8�r�N�j�v�%�7c�!`鈉
Dά��;C
��&e6�C�_[*���R��]�1�eC
�lB�c�Δ�k
��:����L�l�f�<o�)���r!U	@�"�*��v���W䊌��l��:@��X�bU}�do3���a�����$��/E�X*��CD�<�U����3~�/+�L�:��{k�kZ�9�������s�{N�CH2[��2P"�(4����2�֚%J��Z��� ԛ��g�#[�J��q�����ex-���q�	L���{�|�/0�����o���vON�!ş��B�OO��q�x8EưZ��*M�4��F��U��.B�Qߟ���R���L76CA&��7��C��}-7�	�a�/,y�tq���$���g��e�|�O�����u�/�O�(xQ'._�I�D�������;s|l�p��)�:�fv�2������s��C�*(I�ʦ|ߓ����hc���cK��u������uA��� 'B�τ�\P�A��h��5��aӼ�֪��S<�i{'7�jf��2�yi>Hb?u�)��7���$:���=��G�6��h�M"�A��o��sL%�2��~==��/���6�����F�|,*�|	�4�����a��U��\,�W3�""jI~�z�6��أ^]#X.ȕ��_��E�$�7)�U�&v��&Gġ���������EC~	<�mfj/(^7ꄮ�"�I8�j/�IF*�>�����E�fD�|�1͘&Ua\�w����c�at6w�LK:-U��K�@��X}�� ��D�߇�Q�E4z�П���:y.R��R�~������l�H���_:�y��	��9H�c珤iWר�׍H�@#�p�*lo�e���7�J�ɋ
�B�N��a3^��zx�׈������ygg�a�9%n�:~�\Ŕ0��z�
e-�����ʞ�.��U�}*El�����Q{�2K�4���g�R4��< ��t���w�.�ē�E;���|�]�.Ѡrtp��h+�-t�(��.-�{�!r1n�I)Y�5�nꈛ|WҒ��ۢ�[uX��z[�����j�/���tP��Am�TT��O7���A���q����x�a��	�+'��X-�@�M��J�ω�TZ�l��G�P��S��!L/d�W��b���m>�f��E߹���谳��yj�DA�g��K=������{8�����^�`E�#3��w��h��r!Ȏ�����w'������o���Eg5O�m�0�m6�W5li(5�dB?z0��f�? X%����H���R-�'���.`�w��1H4��Jb(ښ��,|�u_�,K� ����s:)3Z����jܵ�3ƈ�u�Nb�����QL�W���ȸ˩������@�"
R��s|����>;�k��>}�d|��̙j�T�?�4���'�ɕ����V�� �ބY2�Ѽ*�BN�fN�t=W�\�����-����1뙲Eɯ����>8��Nt�iϲOg��w债�y���s'�B:�CQ�+S�Ҷ��9�?������É�W��)Bw�7�����4��miox:-\^|���/��i.HWh�ƞ���X�/���Q>Pn��"qC<��.�IpF��zts��5@��S���� U{��ﹶ)o%(�Zvk��ӊ��ˊ�&S޼��u�
>[�,��L�>2����!`�4�����2�څwA�WMnSZ��H���Bi!$dH�����>�#�b�T/�sp��o��G����8{y��Q�Y���%4�R����>`v�=y���/z� ����?�#2T�&P��ٸ�g��������u|2��M�}�D���#�C�ݥ��"<:(�쑺Ȫ�E�~U�I�/�屈1Q@̞���!V�IyGU�_)+�����Ի��j{E��뼑�H_��d5����8��q��iG7��H#$D�ܮ̆����S`�	���X_̎��r�gr%UEU�7����u��Dľ���xۦ�-����S��g';�>�c��r��!ʄ�nɢ�Z&�6B�A�q�9�#~�I:��ea�-�i���[�,������{_�m��3fѝ�mv�\OޱeӓcD۶~n��eK��Vr�ɲ{q�0�⥆+
���M es�[�b�u�s�vw�a�C��6R/�L'g��-�c:�Y��nz�C�ؖ�Mq��g)v��:���\(Ȕ:)�݁�Xx`J����)
����V}3�R�����E|JLV]ȹ��`],�eg:QݾDy�+ߔ�x,��W�M.�k� Lȁ����`{�qK,^f�^E,!o�:��q�7��u�����sF��.K|Y���8j�� �>2D��HX�o�Hw[Z�Y	�}/�7V
5��lW��щ��u=��Mz`�ޠ��y��{vh�5��CԊ䬕�pɼ�@`�gC"R8��{p �r�>`~!M�M�(�MFl¡�l%R����8h�\AL|=�+3����>���ǿt�u~-{��kˈrc
�	��LJE�s�fvk8m2�P}gvG���/���1��Jן�b�5�>�M��X�t��F-F���}ڶ��0�*��ߑ�  &�}���j\\(�5D!d'�Yu��F��0�8�R`��V��W)4.�E�~s�(x���N%D�T��W��3� ��)e���ٸ�n��w�Ν7��zz.��Yʅ�[�ש|5����E0Pۄ����@��1A��f�|8+��س8�����얐�f�C�Vdީ7�dp�z�A�<��kP�пF�`� ]��-"�!z�tC��r>٢�����J���(H�;�%��Rl6t��FK�)�5��?I�xk��QE:1��&�Q�4�(x�LKjU����(�'rI��Wu�a<��vH��3Ĩ����i�b (;�qN3X��'���W��С������o�ؔ���d=����K��:5^xy����!�U�3{+Cd���s�3��(O�C��� �?(�s��z����"'���4۩W?5&Y�_3|�GJ�Bv'+!���M\�ꗨ�N38W�x{rN�d�7_e��G2�v2l
�aE��\)�$�F�;���Z�;7�E���r��(U�C��z�W�΀��'�:����(w4�lv����p|-w͈�	v!% �����v�9�����(��p��H��~����2�x��[M�^l[�q:�G���R�U�;"H���������U?ve퍝,Y0sL��DΉ`&$E���A���l��@����A�l��D��Sׁ,���I>7t����ˋ[C���*�Xy��X�/������L�ڽB�̧�X�5L���J����O�؛�4 r�g���=M�B}\�ѐ�?/?c��s�N	�^��u�Ø�N!�bf	��
�@��Λy�4<�w���2v�cG�,:]���tퟢ�[�� Ժ�2�f� �
Xhcg�M`a	?k��s��it�os�t��x#-�|���x��~�`����0z*�
%,N���5�@�,� \�t�Ki�dX��&��U�EP��¿����nc3��:��d3�}�Tٕ0��bGF5��K��J(%�[,ݟx<���wǙ�
�5N��	�K,�^J�Md1�{�hj0�R�~�?-r��L��E��۬��xU<�S�W���w:o!Z�=���؛�H���T�sSSs�B�1Y�@
PT%���lv>sLrJ2$�nW!kZGܧ}R��<B!`8N��^FP��ɉ��Z&Ʋ��?��u�
ަA���mŘr�ZIXe锲[b�#�RG֣U�cz��V��&Y]4��P9U6n�czI��B,R&�%�Y�|.�$�%��9����W����C���{W�h5���a�,7LnC/��`)|hHhD*ٱ���4��
��-8T=�;���j�+/zoV1Ös���!��}It �<~R�d�v�M ����z��PB�Å�؞�^k|��ܔ!JC���;5zpv��Ιic;�('^�F�>|�>��ٻ[�J����}�Ԧ��0.g��>X5W��	���ꊽ!9��*ы�r���`��TzNh��~����B:� ������6�>����/E(�%J3ۀ���լcut�\�i}l�{`;݂rl�:�������^��\:7$I�m�f�$�F�D������(8��C�k.�Z_̯%�©���������!�j�v����mt}�J&��ym�k����?�F��W��R�?zqfE8M�i �\�Gε���SEW�_��'A)�I��P{��ˠ,�t��w˵y���p����.~�� xiKS��U�S�O�>�1�D|�J�p�"k�n�fx�(���u8��r���
���f=0�����&���].��I_�x���2����@�8�����+��n!��W�e�?��-�fxow\��ԯ�oa煦M.�;�"����9� G�h�@3Є��7G��L�@�_e�Y���z����h,��ѿ���p����;)��*}aH��k��y����$tr�p%�EF#��ɡ�{�)�}ۣpQY�"
�#����.`�����Y�x>�ˮ�a%�Y�Hq���N"C(��SF�Ŧ%A�tŠ���\�]6�'��o�ؘ`H��H��+*��'d�t:{�h��!5��F�]8��:��
�XD�l};5���x7}�-��/B#�<���{�7e �"N��aJҋ���ث�sRC���N�C��H��k���u�[m@S_�c�{M�=���s�
�ѯ�i}b]�a$iH��x��a��h�lL��b(�.��=���m��D�Q��Ak�m!���
ShX^��+�A������R�3Q���6+Ǩ�_�BD_��-?��xW?��D�xx F�61�B=ȝj�J���ZL<l�DT�J�E��du����[m��E���^x)����)"�����V�p��?p�j��%:��Ƞ��zܕb+���A����\�1q�����t���ݽ;�����$���yD�3��T�u��s�?�3r��e���l���(Qw\:�9�&���I=D��k`���nfS�(��.�)V|#i�"��b��+TsǑ(t1JU����g��h���gk����F�L�q�7v�C���0
P�%�h�͍7�7\�}��E7��$]eCJ ���K
Q�l�Ǔ�TIb*H��ɀ���9�������/�����t[S$��A�W)-���:���%��\���Z��{���W�K���&:�ࡦ�E�
5u=�/y����8-&~hk��0��=nv�Tt�|BW��
f��K*B2�\�,_>��1�B��kb�;�{G�2�'�@zڢ��^���A^�7I4���LZ������B�:���եD��*���CA.�Ƒ��8/���,�L��#a�[(�1�<�wpF��~Q��d���{�'�͏�d���vQ-8�@S=��o��*E�5��&�6R��>7^���ːT#���8���W^��^��\��Z�����DQN��C�[2�G]�����o�A�J�+���w�_��.2�Ȗ��b~�B�Kp/L~���"3����ԜE}|ø��.+ƃ� �e �P8�� {F�Ѵd�J��x�vkɠ$��T��34:�xwZ�^������F�=S��^��J����	o�
󂅈�/�4����Im؀�&�_c	�v�J'���y����W�+:l�7�	A{�#o�ttH�:9L�^����r�V��Cڸj�BI�;rWL�K)	U�g�TK�$��6�%��������ΓE_��ٕ����bNU�*٬]F��`	����g[ߦ[�Gt�i�m/x�q-�#�d{��S9@���]���!k��a�G��v�Ο����h�r�9k�yc`X,͓�<�5������D�	��Q	��Ktw���ţ��y]�d]Jm{9AU���#�7)Z�!�P��3��w�7�=&�����J?�5��[���nt%�_��S^l�yEO�����b]8=�Bc�߿v�;%�QG�2Ķ���-6��!l��V���G)2�%!H�"i�-��r�C{ ���	���7���4�76K8����f����MA�r82�Z\ �f���"��'�:�U4�������e�s!�L���V���Y��G��h�=�˶X	U�����[]�%���6^��E4H���ޟ�0'0UY�>�;�0ݶ㘹~���٭Ք���Jh2RL50.B3KyHf%X�����}æ�f�u���'�|C�<�vx��ɑzni� ssUA��^By2�hdF�w���y���@�ک�(|A��w҇�����ٛ�B����@c��y�|T����D����	��L�$�i�����>:n'>��M���T����f�� \R��J���-���ۡ����1����QT6jKC}G�%(�(5��@�B�.���\�m"P����A��r$HN���Ł��ۆ��o�^�5d�8U4����N\�X�tsl���T<CC�G��}���G�W��@(��ߜ�RVT�?�)���|�pf��H��R��3��K$2�VZ��q�&O݆�X�����tVLir�q˳fh�SimI>z"����"�f4Nk��t�k/�O���/�ʙ��Á.3��qξ��:fZ��ܝk@�YL�M�VV���/ �����G�ԧ=M�~�"d���C*L��%�j�[?����!t�/������{�Ч����W,,^�
o�{:��?K�eʎ�����ƞv��ǒ-b�X�)����1�tqR����a��O�H��~w���d�͵��A��1!S��<j��!�z\ש��.����A7=�9z�.o����Oǧ�Ը���/.`���*M�8S�PY.��\��`ۨ&����Ds�"_�X�Ƶҳ~�Gbd�����
_щ$�%�X]J&�*
���f�����q�B.��19��H��J\v��w�pk�π���w�Y5�ͺ~���4ӣCB��b�Z/�5���|���:,�M3+#�Ĭ��`���]���dx`D�q-x�$K�l�,IaA������%{����?ڿ����[��G�����o���i��M'N�ë�#���Z!�3�3o�fzl���2$���3�',gn��9n���~szM�/�����Г��Q��h����y_�(�B�M�^k�9&�G5.�İ[s<��(�	���Nac�1c�����c �~�<Sg�k���H&��Z!8t3�`c���������"����H��CL���:��yW�����F ��9��t9�7̽�X�t #=�e!{8��#!�FXq��nu��͡�<_�Z�d]��E��K�p~k]}��m��w�5�mr>�����$��PH�D"��-�l�z{��+��V�;���D�OC �d@�o�bF1�s����d���9h����[b!5�BB�w���e�p��L�� �2$�#W�Y���_��9D��K�҃%<Ƿҧ���Z��Ay(���t"Eؕ��B������I��EY�)s��ޜ��<�.J�Х#3�N��<�Λ:p4F�!����P�gm��g��X���_/Ԃ��]��T`�|����������[���E��6�P��S�2��@�1���:�=n�Xu�!����xz�����L��OLd��<Qu�yXi���
AH�zL�b��Ԇ��x5��c��+,��=�{O��9�8{��<Kh�ŋ�W��*�ր���{��B�t�#�G	'A_���G��'�Z�)3cs���>�2W�`�?��$������B"hE�����2{�7���Xp�f�g)�Da�S�C�ʖ�R���ٍ��$a��2��h�7�5�,�L�~Um�p�i�$"f�b<{�g����8K��r?Pх|�5km�e
Ԁ���]����}E�k��1��0�!�������n��A�¤ְMm�cڙ\aJ��!�D_�=;g19.W\�E����d+ɺO%�%��ơ����]�9�n^W`4R,/1�ׯ Nk�B���u��+�zW�i~�LM9L�N�s�5B���a[A����M�l��˞݋f��{t�r��Q��e`��.�oc��'y7)���_v4�N�?^�R��y@�8�m3g����
:)���+�%'��b��)���T��%�3{U/\3%������QQȺ*&7|�&�	%0�V�R��:�X}�-g�d�@#��?j�S� U.���Oe�lp!�!#�JJ�}�sϷ?E,C���*2�?q@��<��8O
�#��pk�F�
��mT�x�����zҁ��̑�Ĳ6�g!�u���x {%��*�f�D7H��)~NJ�ѹ5y��K�@D�|�(f��s�Rr����T���j,���ڻ�f����~嘷j~G�hO��>T�i��eկWc������n�8��<�U�j膷�_�Mड��������'h/�ǒ��uN��F�>���� ������HAU)��t���P4�!��Y��U5̹"�ҎD�X��唚U��Ĳ����5,�˨��l�*}�
꞊l(?n�b�G�p��~Nώrn�J�J�4��X�M�܇�15�ar�a�����~*�)9E�"�6���å�ZS_���`��O�a�m��g<-��s� .�o&�*\������Y>M<G�kʏAi������P�����m_qSZ}�۳�%*���1��O}rq�x�n=��2|���'��mS�{,�����4$��qs���v"�:�T�H�W�L����N�<(�$��)B��*�ٱ�QT)	f(�M�`�ʢQ2D��Я׵gk�u�=���p���1�A�����O���l٩�v2�'�/��������v߈�,C�D/�j�����:��_˃����wA)�y��<#.͘^����d�<�~�T��j!�H��=S}����R������T�ԇ�G�r0�Y:�DK�s+_�z���Dҫ�=�;J|gVЪ2���g~I	.Nd�p-a<x-WqhдǢ��`�;'|�h��њU��&PZHA�z�m����c	x�'��jؾ�]��/ũ-Bd�hŻ�?���#������&88�����m��D��h�r��	?;w)�l\v���v�v����94�q��L��3�aU���>$qo�~��&�2������ECc�{.��̽[�/6E����'��,9��t~J[z��x�,�/C5������l��J���lh�BS��Lj��uO��3����IO�Q����j��Ow����4���K�s���+����+X���z��G�v�z�6	
<�5�2*ʟȤ����x0��d�E��`��K����""R	��f�ʉy��㼊�#O"��ݗ����\c��A5���K	�!J�9v��o:���e�G�կ�?y�␈�m�[����+>F���32�{Y�[�Bl�^��$�X�?�˺��[n�[	i�=���Ss�s�g�q���������>�J^0�4���,㏥�B�>z�p12x]W@�)�D�hDp�uiO����+w�Ͱ��ά�4Ǌ)�x�e�Ocd�c�bm���N��ȇ��9_����5]�R�[!-`1�@?~ϱ��OT�`0��#��Ivp�v:��_�F=�u���=� @lY�ׂ��]Tg���?���E��T�N��o�0�N��W���Üp�1G����m8Fʼ��O��36�I�؇�P��Eß%.2
�@T�+�,@��eU�O� ����?t[��͟^`a��f�&ڙ�2���~k�4�_��3�23#���Q
��=��Hk7�^�zN�K�H�V\�X/_��s��������M�r�5蔂�d��"�(}��#�0n�T�2���M�Nء��X��c,�\�'���i0@T.z�:p��	
`O�t#�PP�3D��/�
pi��������n���2���3�Z�×zπJ��?��4�F�dY��E���"0)�+�Z�+�J���I��âT{����k	V/�ݫ�{"��?:�B�5�QQ�j�*b���XlP&b{8[S�h��q8�m"4�����Ew���j� �������Q��"WYS]�]�@o��"�$���}:Iƚ@��wh^�#3�s�������t�b��t��T���#��޷��&���r\۝���Rf#/E��x2n�9g��bK�7Fr�� �� �yJ�ul>xk��j�{�?*J.T������#��_�Ȟ��	y���c���V|���	(�0�j�FH^SD!��Sɧ�p�2y��(*K=UmK�-{������Č%̫5���.D��2� �u�N�C��h�h'�K���^9�z�k$E�u6q��w��!g
ε�9o�
PE̽�7�Ж�;���Ȫa�˔��Gi��&gG/��0X�,ϩ{���. )d
[<@�ݡhA:	Z:��zc`5���+���C�L��mj�X��Nz�ȼg���������2��t�ibi�����l�)Y�������h��Z�jk�7}�X����vǫ�Л���e���w��mFP>����^'.׳>U�G�y�����X� ;�s�4ƛЫ�'pƪ���*?��CL
�FF��{'�?�W�����A!�?"r��z�߬� �w�q-<�>yaKw���;�A�G>��h�~��A>j���I�J��������o�0UŹ�0�R�HlA�1�W�Bw��3m]t�I��'+ -��q���i����1ܢ�AP+A����yN�{�â:�q�.�=-����ON����5Av�e��ʩ��1D�)a7S�Y$�*Zf�_����[� f���q(6A͝�".��f*�M��q4)����͝�����e����2�NKi�Q��[�<Qﭽ�d�Mt)�Z��H��ʿ�DR:�x�糎*&1'H�X�牠P���]ʸ>Iw8D�3����,9���åVלj1��P���T!b~,Ni<�X��82�3�d �A���t���!�N�3� ����2L��_��}�tR�ʜ�(��u`�c������D��^wߙ[��[Q|���2��^���T�X.m��\����p�B������k$�d�~�FC-�?=BC#��ŏX�����P/�� ��,��6 ^�*%X���٧�b��(���i\��\���'^߰ǧ=����sfB�.6�b3�dY�F5��ߪ(iiX�P9���fR�L@ֳ�{`�����K���w�8HCZ�휸�%,V� �a�����P��%�@�ut4���/s��D�.3KX��"��D7��ɔ�����=����Յ���&��*~���
���{�w�]�m$&�1��8I�!�E�V>QՊÆ���ˡ�}cK��+��(�ώ�o���ƻ���������tK�c[O�V���`fgP ߠ�4�kS�p"=;��A9q����^�jF8��O"����;EG̮&�����5�ﮔ���`E�ae<��r�����t���j\����l�d �*�2��9la!���o��2�%T��h&�,�x�҆����޿IEaP�1����@�9O�8�7�2;O�P���w��a&>��s�����-#iP���6�N_�ĬQ��u�;,������ޕN}��R�?�&S�Q@E!U%#/2%F>��E�K$�������f?<&|�I��r]��%KCü��ťJ9�Γxo2��k��Q'�:�Ӷ)28�y�C���o�4�}���|�5�~<Σ1CV �0�<[V:��<�	ͣ�?v��;j�9rCV�s�q_�HCAL7pk�7��C�_Ĉ/��Ԭn�xK��6Ҍ�1����6�?7->��b��p����8��='\)���U��4����ͨvZ�͔#�һp 9��S�tU�߫�&H\�U���{�C81@ͱa�ڍ�TK��kwr7b>k��ePl�V|^����)n�ɚ��`9ɬ�*^��Ā��1Jp���'9*��]��a����L̘(M��È-c���8����e}?�76K�Ҹ�'��}�R��3%x�ɰ�R�� �����i	��3���<
ϫD�p2�����/�ʏ	<K�g�?QW��@Y�v�6��u��A�Ϧ��q����p�t"$&�po�aĜ� yV���&��Y�����*���p��������è�#e��,��!2�C��\�R�*$!����D�S9�4e�Dn�4�h�S'�/�V�d˂�*�jj*�-�\�
����FNMD���Ύ6��z�7x	$����E:$W�/�m���b%�Kߡ_�H���i>��M��i9�ݬc�v��h!�N'��D5�`�$��R(zʱ���_��mؔ+�$Α�ZF�����n�}x�ظ]����I��S~��&>#c�
2]��mk�t��7����2l@�S���U�N0deyc兆���M�?y�t*�$x8��@Y�hP���+X�&��Q�ÞI6/�1�,�{}�@o�w��K0Z�=���ut�8�ʪ����]��+ߎ�ν�f�C����~^�N�~�>\����������w��4��#�^u����������(e�p&J�I6F�΄��α�R�ig2�@��N��:1��Ř�#_��bd�:�&���`!w�.Q|A������)#�.
^�y��{�rI�:�Rmɽej��=�U�ߠ��]��P���(=�D{O;L�����rZ��ǝ��_ξ�Z�$��*�<�Tko1 �e~�)�'��aU�Ii���&<�H�����*�<����~�~j�e�rͨF�w��N0ԁj�!AH�X2�?xIM�9�!T����J�
(�<hs�A�x¾�F5s�
���ux�ޜ2{es���斮��ꌆ��Pz��� e�aZr�pK����n��]��:�[�P�ߙa�X,z�vQL���_���\�β}DX���ߴ�E
B_�����~^��e�h�)[Z�c缌ߌ�1��q�llՒv^����g�����9���֤Շ4ϩ�4���"����=#b���Q��b&r���p�����a2��0�&�Ďa�����ڔ_o{����j!̘�.ʩT�.�&���F%���kM2��-�d� v������u|�m�?r?>����}"s�(a�g��wS�i)P]մ��J'��Udp'�����Yu�Ý��ЬH$�s��o�h���t��E���f=&�ڹ�� ���]8��6$��"K`Z۱�Hf��幟�".�<�Es򩗬Cլ�Z��C ��3P��y�󷱫d��c�f�a����WW��@�ϰs+'��0\^zc���"�D�#[�Fc�=�zI9q7�»]*2KpZ�����γ��r�_�`�� ���K+h{�Y�5��q�:O�zb7TҔE�)�_�!�[�p��{�@w�:2�~��9��{��(��!�g΁��q�6���� ��Ĵ�D/т�4�N�,ۃ�iE%�J��/��kb�??�p��{���)a��~�����7c�!�o ��+�M\Oi�����Vݜ���jܪ�#к�ͻ��s�	AZ_�HH�9+G���js�K�Ϧ���`�.�(=��4�N&,�kw��]s��\�)�\���A��뗑/g���"MI���En�xZ�mN_��?�D��$�>���y���k��$��دD��4a����+�lӳ�r���$P���~�c^�ƴO��	X�H,&�SE6G�7�6�(�� M�V��,M���.������^��-�g0�03�Nɨ6�ߟ���ޘ��͸+lߨOY��a����綼��/j~)�~�܈"8���l�{�n(CDeO������cw s,����1��ɛ�s[Mbq�"'����gc
�DK$��$�:UF�2_����R�͒����Q�������6����P9��P3	�)���]�'4g!n��7��F3�u~x�- �ˢo�P�ݯ_��Pf�㪡�>���BJg�^���������:�R��.��j�Ff[~���� �C���{�Y����F��#_��dN�.�S���6���әU��q��&(�gB�/Ϸ����焏L��A w�Ed�m`�_8�-Z�Zz~V�����w�-���j����`%a�tD�:��.�P0�&3�;'"=
1��؃x�`KN��yn4��2����&)HW�<?q ]5�`��񿑞�q?v�3�B�P��v֞�w3kn�HLQ0/_���~K%�F�j��\P�=Jy��g(�7f�}l?v�oM/���0{�Z4!'z�?�V�r[~��ZS�$QO�'62g#���]zBQ��6]
��&���@���V���3$DY�t9Ù��͊�{��Ͼ�ǅ���f����{"�j*e�nݓ<8�ŨQ:�N릙���d��zg��wG��;�UƐډE��G�YJ����F#gT�G�o��2��.R&��`\��+u�[u�yT-�Z�r>k����oY#"���E�5�%3A����J���l������B<^buJ�v[ֲ���.w��x�BF��,m8k�T_�sB�pq�|!���U�K�dP�~�5�]��R�ֆU���\z��l
`��獦_�?���
��4�#^�]��bûnX��;_6Ӣ����z���I0 ˼�5���RƆ@�q�ʦ������1Ϳ[yo����~��7�b`�o��tl}��3��7P��X��npVF��^8�p��7}�K�,+-{���Tiqa�l�{v
AY<ҹ��i���Xn"�nÀ@ue��Av���;��ћ�;H�>����K���> j�4anኧ�3�����OnW�Ƽ��/V�84gȾ՜�T[�4�\Hy�A����>.�K�HL
~�l���Ą�6PW�_t���N�����8=��6���N�M�n�?#�a��)'{�hˇ����.�`�
���u鈅��vJȐ����T��*����ḟ�i�����p�%W}��1�����{K}{���Ք-*�h.�)���K>�Z����e�{�~w��w}Gg��>>6��u�t+��H��(��.������ ��̔:H�3՘
4���g��/b ܸK{���I��
���p\�ϫ=S^��������]�`�rJ�8�
YS'\GQ�Aj^8�"�d:,|�6��a�[�̣�;��_cs�?΅�C�����0� .�_R�����3��G�s��G�b״��	nݐ��1RjÝbɸ&�D�޲	�$�4{���m��� �0�_�� �5Fd����6x?;�$6�3���Z9?��;�Ʃ��C�e�/R&��F���n���6�AZ�U��/���"���_�f��f�2����'��T@BW��4��0е�+s�k+�&��Zb&[p�;xS7�@�+"���	��A������n��ؗ	蛧�����}�`�AcCz�"�:��U�(���h�==
���}��PU��W߀ցBbz]VfSA;!ιY�V�S�g�l����(��!�6��
�Nȁ�L��S&Snb$��d�hoT�O;�yf�7�Q�!$����SJ6���	�� m}�gЗ���	H0
��x�kɪ:$��[�L��n�r��O5H��3#V��g|�5$mZ�|�Ͱ�e?VOz�K�Q�ׄ��2�������_k{I��.��䓠�H �~#��m�`#��u��k� UT��i�֐ƻ13j�a�P4����}�$n��C5���,������R�l7��v>h������1eu�	��9wjWb��.ܤk�5\��<���$� R�Q^�!��~����{z��!g���Q��m�K��@����Y��rj�f�k気sv�cV%ɸ���fZ�d]�
<x�W����se�F)D�n����u�;l;P���nk�:8���F�v�4>a �wGGyYDh�� t���2>0�#�j�0�y�������FK~��Ns�j�e���:�8�JW�07������л����N�F���7�O�̈�|�0c��d����1N�/�O�/`
��Nw��X��c3_�\blh�[���YC<�׹�u�YM��;�m��Q��p<�b���3Osm3�T�\���_Q�Z	F��n*��v�3�L��V�0�-�a���mx�Qё�Ga�d�Vmʨ�J	}�Z���v�g���E$	<�?�EW�y>�E�G��iג&v���f��`8X�c���B~ $�R�F�ށ���ޚS���m{���E����������è�a���\��Fy�`����R�#f/�.�hmɶlVؘ`�(�)N9`���gf{�������?�t�WJR��*���Z��[+
���wƈ��Vv	�I�w�p3��$��u(h�͆��.WK ip2;G~��	1��;�1ID�Q�^6��bg�)��FJ��ʡe�(�>�?P_,$�!e�1�r�nw�ڹ��,:��;��;���<9�,|C��2r�!���yw��8.��t�H#�$EXYyKB$>BofF�5���k4�2d���C��8��"n�ٷ]�ˈ⒠f���v����~�u扑sZ8Xf����u8����{-�~���3���ڪ,������"�f�%�V3�1	[X���va��n�k���q�W���M�3�O����8�8��L@�%�(�I�ŗ���O"�Ѵ;J�OO��Y����Y��|���`��䱈��y�����t�Q��� ޵�� ������1z0�G6�{�O`m\�c��` Vh������d�WI4n����&<XG��ޢpY����8?�l��o�x� ��
Tq�w^��L�nZ�È	�%Dȟ?/m
:(�n�S�U�-!��S8��ݻ��a]�J������I4����6/�S�QN�1��C��7����(�Sі���{�b�)���a���5��>��z��(,V</������y�g/'6P�Rc��>��NӝZ&�ZF3*��\�Wz!��1��2�E_^�%��z�c%t����k"YNu�+�|1���0�8:bU�ΪY&]ܜҳ��!-b���hszMљia)@�ߡP�i�)g�D������O%�P����)p��÷��8(�e� ������pX
�HmE��l7�����^��[�~ �7��E�����,�ծ�wTGǤ�K9�4�"�k��.H
��Y��T�$��-��)Jj��y�AE��� ��O�CL��!�M���k�����P��,�����	'+ɒ5��{8`���,�G��Q�д+ܫ�q�JWH��h�����r|�=VWA�X2��ۯT�$jZ~�,�$X�Z<�`1˲��8�4�MF��0$e���~�Ujm��:5��4)��R�v�����O'���(M�=���i~�2k[��"�����~��t�R�;Ql�*H]㰍�CG�֕6�a(:AA�h77�>��[�@}���V�Z���΃E�{�Z���R����d�����yF��SHMURF��BCjj����X�g�L�'DB�8�U��̎�*�$L-3�|�:^�/�x~�&y���،����Ur{e�w<�sY'_�g����A<�G�	%|hS���<�}���.���'$%���U�KDO5���@�=�Y�|Ub��@�7ۧ��չ�n@�=J�$�+���f(�}j��Y�*���}I^wH�����/Q�K	��=�O0���g_�%�g���נ:wD�+��,'�M+ .���ZD4c���z}PO�Ȳ���3�ȿ���mň������q���A��v�gOQd]�<�#^��TA��Dk�ʲ���G�,5x���H���%�?i�?��Mǰ�x���_��}��r��-xnP*{	".��2o�j9��9�����6E<�K'<�ui=��jDu�+���ٹZ�c�Mo_~�1J���U��Ĩ]�H�� JL���.����!�B��^@[������H���u�K��6>�1�B�,v1N���3:�x]YAu��i��?�_�R�y��x�̢�n ��#e��}�c	)��B9l
"x��q���\Fz��˲�͌5"���r�_&�	���Ʊ�7m���eه�W��Ṯ+�;��{m���I4;2טy�!_ ^�u�&E�lx�r˺<�JoN/��5��v�='\eƿ��ؗ�+_=�8uޱݢ;�-�4��jц[{1����s�yC�����ƫ�u.���&�^jH�Y�O)����{EzՄ��x�Pw�q�߫�	o"	������=ZtV�(����P���^�y ;Z���~.���b16���a!�PP~\���~�F�\�Ԋ�CC21�8dш���8�Q�A�f��y֮ۍm�;���P��	E���A?�3�Uћ���d��\u(v�U����,\��|'�ɱ��"�AG��Ǭ������`�
������T[Ja˹>7.�'���O��<����.��4�u-o�Y/�d�ACד���n�}�t+���TgD�d��:gt��������]���G &�_�Μ�nq�/��ihJ�.� �N��I��'�s�cfX�݊X�'g�d�a��,��17��ݠ��3|w���Xh�M����:G�h�m�I/���H��Q��\��XkHM�I4�����ȇ���˞ ������x���\��Ɏ7-�aVf�r��[��t���I
����iW�����i���O��� 5���a���G����cpJI�7e��XB$����jUC�dCi:��H7%GY�e���b�ha(v(���1i"��0�*=7�z��d��,�������0��m�hI�\o��H�,����Mq�8�#��3�xT�ӆ��N�2�H5d ����s�jEC�eL!R���HJ]LT5Ʌ�l��g2@��֎Ԛ��>��ت��� �s�D��5(s︽��Y(?|c�ŚN����O�/�ț9%}�­T�hhf]aR݉���P�Z��B:��Ȱ��&7/� �7�2�q��+�
Ԧ�Q�
��q ���h�����qTr6�Y���S����:b��l�a�(���D�eў7��4-"�i�&y�ݜ�Y�a����b[~{<�N$�h�/�fq��Ҡ�*�f�[w���A\���R>����[4b�i�v�I(%Xb�w') %�A�0��~�}�ꈹ�:����M�v�55�Y���h_%"`{��MH��d�ҍ�ؽ�e��ؕ��h)yc�z�s�3�3��EȑbRU�ApIU����{udս^UR<��B��k/�Z�ߘ�I�9k���� cA�u?�a-��j��d�@s|k�E��+�cncF��d��C�.^f��$�b��V%u�.'�HS��e�`E	��� Lkr����uz5R7����v�}\@
��%����]���_)dj|&����p�*K��9"y�(�Y�*ڐ�P��R��P�����d�>�mG8VBc��{Fr��e9ɌҌ7���W�x�t��u$��]IA�1�q�(�=�Կ���8E7���%�MpkB�f���q=���@>��1���T.����Ur%P�2�5�"��i���p��O]Ep�׌Nx��ʪB3>)@Gޖ���qxw)+��3��׮�7U�pτ�]��g�_������%냋����^��i�JQ֚��e�&K�;�+�g%���z�빱���.���PҋK����1��.��
\�z(�ӜE����� ���$q[b.t+���^���ym���=��z�5z�7/��+v��mT6'+�\�d��K��΁n]4�T��4A.�E
țx��8n>Ǯ�L��.z��^R��V�Uo^H#����J�w/�7`��ro�sָ���Dv��Y��ޢ�0�ȟ�MC�If�0��E����ކJ��}��5i����m�
�X�X"%��|�n���Mr�}���*UE�Y_�53���6{_H��*���_w|��k<.%U�<�N\W�]PO��+w� �g��>MU�]xht4/�G��L��.�{�l;h��?�:=���d�澍N���E'9˘�қ�8��7�e\7i\��#��褝�^_n�g�����oj���4<���I��^��|(Y0!�~�U�sfӀ�(��ND�G��VY!�� �l�C=p��%tA��'�� ����r'�f)����S���1BU��:�`$�b������9��-�3�s�6��7��F'�eO|D���$t�V��~:�}��R7��i*k'�BMB���hR�S�fO��*����24p�O�����bd"�[7Zz�§�4�M�S~���'��@�m�׷l�`��P�h�u���*�cz_o����v=+k�?�����dbd�k1�Eo���a����ԟs��m��X�<
w��?�[��X��{r~o^�����[�" $u�S���P�S8[x�6��%���9s��JF �I��T�
��mp�l�u���������3���%��o�
%U��.ȩN�_�*�������E���x�KD�oTD��or�4��U�K����zhZw7��Yl_��"4L �cV����_��yw�~�y�/"ݺ/��@=��)�n$�3{�z��!���~�t��Gj��D4�µ���"u��=�&����<�Ck^���&�ƫ�͗�O�7X�Q�0���{ӥ�>�:�fu�͋�R��o�V`�ת��m'��W�kƟnR�آ��������|�G�`Y\�1��(v��\}��T�@�N(`�a4>�ȝ���ڱw6G�*�����]�>�u߉�/��̩5��t�x}B��U��W��+�IqNSg	.W��l�Z
Ṇ���W2�m��'A uU���F�`E��qm����6w���/Բ�飚x��{K˂i��̭�wf-V�9��G6풍n$��f^�'߰?A��ޚgs"��w�^A���m��}n+$Ԥ�Þ�ߡ�|�ٽ(_(�6Dܰ��w��>��p����i���G�u��=��,���X͢�`�ET]�J�53�\v�b9{�)��-7����hwT<�����Nq�I.�C0�8�>���P�T���'�I(�)���)`ɲ��,x�VĦ��ď5��|��ͪ�Zh=�ع4��䖤�i~S�+���@��܎N�*B I�aL�L�9x5����z��� яȑNGY��Gӫ�iN`^͛��b��F���W�փ�q�d�r���r{��`f;��>Jz�t���5�4�[�_8����u��P�VO�Q;�+�x�w+��H�C̭�1��A*E�ܤ�qE�V��eqIG��I|Q�I�bL�_�ϒ�J W����ҞN��y:��9TA:F3�����TD�lE[��O��W�;�~����P���]7�z��d���j�K�8e���Ť���^�p��ʭRL&�L5����ڇ 
|]��n���>N�����?��7��S��rQ}���j�r�����'՟d�v���i�,k�/B�p׹����wJ	�=Jo��1)*1(PA��M�H�H�.F�a3$8������7A�QdM����܍>�:I�2Ï�����)M�'��db�VK�|y�0 -be�d����@N�MuK�p,��7+ҝ܊D�n-�&#�{A� Վ@�;"�V|^8�K|̊�g��=$����@�b>�	�H���6�]�a�d�89;��^7.���<d1w�[������v�X���̺"�l��z+RX_�G��N=on^-�ln�|��-���n����*�_���n��N|�������g�Q��-6����r�xC�_� ��3*��LT��S�,�8�N9��c=5QlV��e�aRN�e��Z��iuF|�G:������O�Sϵ�~R�1���l�(n��a��U�͕��/�B���%��{�f˛�������M�q��������7>���I��#-stRf�9"��^��o�(+��)���ܐ����o�l'ޗؤϮK/h�ڗ�sK�Pn�z	����(1��Z4���G{�KrE�Ӈ:b6��|5u��E�_X͇�dg�ŝ6¤�s���U�7���k:J�Vܻ���qj���5y��7B��-�HU'Ue�?����<���nL��F-�u	F^ڈ�пI�I�~���N_ۀc
4�V���O�~MhgPjۃu{�Ovb�`�<���d�50$5rHm�͙V����"�*�S"T����)�Vd�ܔ�^��׺����b�E���s�Dj����*x���3¡a�ʓ�ҵ��q��.��-q�4�_�����h��qpC�ֻf1�s�����7��%�S<:�X9ŭ�ۥ,<
�U���PE ��>>�V�(��NF;(���WfW�Z
;d�
�ɴ�uƫ!����ғ����Ԗϯe�A���;���'�߂��x����-̞��ʠ��o��8�-~p(0�)�tz��)]�׊�Sk�԰d脖�P� �K>�O.|���,J�F`�)Q���ՋWj�K.)b�k�!;�7�`6 Vc���8��BN�(*Eo���5�� ,�����=v{5i�	�Y&'�S��)��_F���;\����d�^��9�p�MM�',0�F{�h�{Y��'.�y~zΓ�����(7o_�A�Lx��ʓ�ۭ+)�v%ab-��j�N�R���f
�v	�]�*�'\�o� h1�$`$�`&�ÆK�z8���T+!�� ��됕�|�!`p*=����6���+l���ۇ�����Q�׸�yE��!1]�0N�U����
�ݑW-r���!��0:�)�6��g�)B�T�!$�PX0�����%�9�\:�E�g�;�X����n�" ���zȋ�q�&�|���Ze�6h[�^�+���#��V��1�郣-��[L\m"Kr������� <��j��L�+m٫>.���0/��3�2=U����Um���t����,�Do-��j駑aF�E���� z�E������&${�!��%ޙܕwf�z�Z�~@�P^���$욠� �R����|�e�aȐ%��0�k�1;���~��'d▭������|�i�X�ƕ�<�f��҅�le�'r�j�uo
a��v{l��������b/^������<��?)����,�:pɈ;g3�#��h�xF-�0�7z한��W�o"��py�ʹ��E��Q2�O��_�6m.�	D#B_��З�䠟k�k�����^q�O�������@��+��t�V�*0�
�i/4E�t!a�~ZO3�J����&]]3�	����#0}6��Nrs�8��[ִKV�\𿴹J<z�]�:�r�qr��� ��XƖ����)����.�!��Fo���Wa�!�D�W�s-��&���xR�6X�Ti�X@���D�w��,,Ο��u��e#G�!� �u0���݋�(�PNp��7D������_o�7f�]�^N�˩��"{akR��j:����Sm��2*L񽅡���q%��)V��)N��(]le�G-�ȁ�,^����eP
X���@�^���w`̮�7�p��E���J�0[���Ñ7!�/�>�Cc�W��Ih�L�e���Bs�T��U���߉K��o�pw�]LV���h!���X��c ����V�D���ͥ<��G���`��x��tav�T�^�^�t�е��ZJw�NP��=iZxqt�#E+�zrynt��_R�)�j0x����)}�Wa�ù3.
N�c���S�A� <8���������_I��v��~AK�Fc0zD>�`'n�jt _"-�ʿMH�9��z�����;�.�l\Tc@��$g{4wR-�h��yv�b�}G��3'2�r͚TNO�o��⼜�O6��`5�1]I���̻�|Ηk �#��Qq��@ JC�6��>��t�n]&ߒHw���Zm;�|t�C�"o�y�S��أs���"�%Ug��&�7�b�m����θ�M�:"�O�3E��aq7��k�,9����jl�Û�����JX����Y�����_|7���҉^��۵U����c,JFj��(s�vԾ�8t?����y^�-n&õ����g�5�7rGg��q�&5�w�i�ㅩM2@/��S}8P ���׷�(���o�@_"�d3NtR��n	����Ǽ��w�o�UT��cS������@�i�=���.T7~��'�������l����m+NB�ϙ����
��G=��(j#��އEэ���=[�'�ͼ�wՃ9�P��
�g¥q�?�(˶sX�?�P��p/�a�}�Y;lG��tB�`��:���隥!�J�f�,�������͟�K[f�SZ7Vv '��.���O���~�w�� �4�K�c:Qq���<r�S�K��3ȍt�Թ���?����9cC(��H!���0��R��o����)�ڟN�;R&$�3+�gf��QJ�(Y��/��"���ٶ�b�]���#)51^8���,�W"�RHY�=�;��QD��`�q#|�?�5�1��/)�/֔�Ap�4���<x�"���6��p�@��:%p�7�5���#��	��W�����d��M2B�g�>�c	xM������حms	եioX7 "S4��*l�fB��(Ow���X����X�
/
x,�$�#�����Ǔ�i���y�����e"�mQ/hIx��3�,z���ؾx�i�Eᱚ)�>�3tWɓ���V�V��e�5_QČÝ��HY��S�>g�7����Hn��g.#NAE�|�ٱ, IPG�d}ؐs/頂O*���{�!���UU�-���ɓ��8�#G�	�aSB�/]ꃒ�\x\��iT��:n���W�9Y�B�i�d2Q/�8�:�үA��jT��͍��3�i���9�����u�y�!Qd}��t��k;N��ҍ�����JgG��z��Q�*�d��%���ϖ-�O��C)��5E�Y�SE��a\Tc[��+&MC&x�M<oD���L	�����?8^�3�cE]��3�u+N�̓�s��'�<!�Z���e�Jڕ�^����Q��$>��O6��.|�ІzQޞbO5�K���Z6�;���8�ɀ��o�$�)�"(p�.-^l�5��usb@4�ŏ�� �u�P�3������x��� �f :�S�]�[�p6*ή%aX(�-Y����
�\Q�aJ7	�^U�X����a��<�w�D>�i >�H��4�h/jE~�����o���1��/��o3�([B�_��D}
3�{y+{a�sx����c��x�~e��.-��	z8��;v�e��$E����E6��4�Mx�7t���7kdu�^�;�Y;��H��i���Ƈ��/�9 ��ɨ^�:!�1�E�8������ێ4��M�������lj�x5i�)�K�r���;���O��O���,���(�Q�R�j��ȋ*<��eg�
��j��	C��~F	{��b*�Ԧ����b�d���<G�s5.>?��!Oܠ�Pм����Z"� �W#8�	7�%��_!�7��G�f݆L�8��^K�O������6\C�	#D�}���}�oA����	�uK�3eߡ�4�n�k��r��`�GS٧�� �Z#��(�g{��߃�}8��	�,�2�px�x*Y屌�@ :<"{�"��V"��@j�h�X��a�oYn�/ͫ��1���Wf{qӾ�K���|ӕ[(�4M"�'q�E�\���/�Ѷ�{�(���� >	��9��ku�J��:�"����]Z#nEk!�e�:u�7)�5h �G`���� J�摩$ y�aL\�q��zzܺ~���,����X5�hR�}\<����ّOU3�TuU�C��E=V!��#I�9�fK�vD_S$�D��5�tV	����a���a��?L�𢼏�ZN�yd�`�Rx$���-�Pp���vPJ!�u��ƥa�4�kf>�"\���/�Շ4�?�p55����-��H�3N>K�9��\UT�FPڧ����}/a��m~Į��iӅc�C����Ʃ�	;��WcO	�y�Y��Z�u�r	�+vg0�[,Y5��Ѷer_'|U0��ז����+M�Ċ;mS��\�H���ܨ�s9�Ժ��/��$ W�~w�.8/��P��2����j���ݠ��Y����6��P�-�3 H��w��z���Xgߋn�I�VY�� �g�kn.@�q`���2,
fi�"����e�B�D��xj�7�|v_�����<U���M��V ��,␳t���G/S���i��j�Ø4t̫�����`���K�r�u~�Y�_o�Ij�I�\z�Q�@�Hn*���x"$����F��d�%l=�w���*Tfˍ�<����
�2|07��0�;�Hܵ*嗽��ca栛|�GQ�@"�l�!m.4o�:||��l����T�o�Ͳ�@rbw	���>�v���D{+z�������x_�3o�#B_�Q��r�Y�ւky���uBŜ�E��p�*�%zfZln�R��)>K6O,a�kl��sVN�0���S��X�5HG��Y7�K;�P� kZ�民����aOu���Sg��ޣG����Ӟ۽TK*�׻�%:ի��M�~�g��z��x���F ����@Ll���k�H���^��M0|��Z,yuT�U\��jK�� ����	F��"n&r���_w.R]��NY�gpn&j'�O�R��f�#w�<)һ��-��\lPe���)4|�[��2�V�/�+:r�	:�����l��5�>pk���f(smʧ	���/�軡�[To)ai:��ώ.��bZ�#���/C�H�8��o~M����d8���b:�η�����d��
����,�~�W+&Rח�3���a�f�>\�o��@��Ƥ�B"b?;�:�����_��L���GW�H��:Ewv��*Z�1�>�[:s@����ٌR�/�ܔ6׍�y$�y(�A[�}ם�=,ŀ��d�a,ح�_@1���0��~���]�-@��-���}$�8�zw&��&�:����B3�:@�����w:j���H2Wr2u�*q0MMĲ4
��*,�.�.��[�ǛjY�a�@ʱ����M�>�a�Y�;�n]g���̙π��#PhU�eN#l��#e�*n#���`����6O�m�FA�u��Gӛ�[��b��'���P�����'�.�6 �����wt�;$����4�Po �F�|2���H�R��n�\�1��]j�tA�Bmb�mxU��^��f�F��Z{ɩj�m'C�+H%�d0�W`�47f����n����M{�x�d=�
M�byz�( ��]�q��3<IHJ��A�ɝZ�wѪ��K*��~w%�BW��&�{6;F4�1�������.����<.���JF���X��OR���p͡�`4#pa�1�2ē�+�B�5�j��0=�LL�gkY'#�Kj�b$5�,�I�l��-��28hϾ.�A"(_���6�N�R���A��*O=��K��]Ղ��s������R�����TZ�}�D�����w���AI��O�?#n>�!�0 ��X��_�~�?M{Т5mY�KwMqi��#�Y��ߏ6�J�W���W�\�B^G�bq +��妞�k��QΥ�2{叺������=mq?����:M�B*xt!HG�ʰ�� m{���x���~,ҸC��P��q�~����B6��r�i�뀾s1�y�섌J�P���@�xa��a����lC�����\ݧ(q��8)�!]r�,��pV�UÔ�sK�������tdk莘���������P��RyT�L��gS��N?��\"���h�4�G3��,�I���=�ɗN�[hTrOU�.��1}[ �Q�Mj�(�|���*	�x�v����Ov@����x�X�G���GZ5č3�a�?�|R�r�M�Gx�5�ʸ�J �C'��1�0�yr�Zd�O��C�n�4�0�*x~n�ok`��U�b����zK͸x�l8;�bb������_$���ph��f���z�[uct6�=���	�q�f;]�:�+
�QKQ��V��m��!1`=��TE�^h��M�E�	ȫw��0l�ɏ|�Ȣ��|�9tf7�Tt��+LG�{?���1Ğ�qv<��?�]X�FO�VY�؎x��
�Z�%���d]T�&�w���̉d���^�#��ռ��>0 W�J�L����W#�ڵ���|��N����ƴ�i�.�"������c��r>�xʑ��C^�m��tr9_j9�Q���ٕ*�q&\o���:b��gF�p�*�܅�Ǉ��p�鱰�[4(���&d�2Yh�@ŭ�@��A�>m�[8#n�����v�X[�f��:hG A�Yn�\ʯ�? ��a7�1��l��n����ȱ�'�`?��c0������5n�(z|&MK6�T�ڀe�c�_��x�
��_q��'�HglX�&\^S�a�;H�ehVfF�S=�|��+S�U�q�{/1��/�Yx��r��O��b�u���xr�J�O��RH��o��iM�3'��(f@�&1uE4��A��^�sr&�."o"���݀lW}W�~�@��pLwE����Ə�p�!�=��5����8����pt)���]\W�!ɐO���'/�e�di�F��_&�aXQ�k�տm��>&�"����3�N\n,�s���~�r9%A�Ѷ�UdY]��G���B �N�0f���O?��2f�5Z�L��"�n�t>\N$H��Zp�bGyKZ*��6���&�8.$��'��5ވ�Y�1� ]'Z��x�(��=Q%����a��%=O�p
A���9���9+�.������]�����&���'6E�4�5 0ƞ&_���f+Y1}���Gӽ��#}������W��T�,��*u%醅�*�~,�pCP�!��PS#��J�Q|�$P�F5��WH�m�x��g�?����a4���^Z7,�~�?�WW-��~d]Hk�?>�M�?S6�k!�Q�4�)�!��3hˇ�G���j)�hCujŅ{�e�>��4�h[�۹"��;4�o�+#M������u@U �%CJ�V��(�$����[�aʄ��D&�3�����¹����0�6!�?�ta �6�P�X�$��;������n�09sI����³r^�|��3�+�MH�n��/؄��Rf����Y'<��=�>u��WNnH�	.�Kʶ|%*�k�᱌���!�(���s��\DN��F�Lt/����"�(�ʑ��aE_�=x�{���h���ꌚ��C��ϛ���z�r5��o�kF���m��[�騷��f��}WѲ�053^ϡmY��]����l7h��׿O�ޚ�b%$�e��j�C󿟑k�H� ����PXR�1L���*TrIn����Q�2�RQ�S�Y4����@B�@8����[�?���Welj��s^	��W��a�ᾝ�(�ߜ���;Ja�!0 9�ς1:>w߈?:���`�!Ӷ#r����h�aJɾ(K ���y��;�-�S��ޏ+�\`)E$j}n��u]�FQĹy!�����x	v>�>&6�o�E�sϽf>���YUD����h�8#.����ij�rBP���I	��!%#��;7�[l!AE)��J��'�$��
�M��h��S�<�����:���A�񲙼f�#�XW�q�=��iڊ]�"�c��3&�3=��m�a�W�8;��b����*w(�E��Dt��h����M�3Ik������c�#���e<�ʩ���X�g�̩l�?�K(�f�p���Lb����B�� (v�;O�����R
j�N�5��P45Ԕ|8/���ޖT�G�;���o_��S�ݖ��2�l2���K}���Y�����~H���gy��n��i"�]�S�g0&(T��i�¬U�lV"~0�_�=�*�r�w&�8�c1�����FIK�/���\]�x=�;�+N����aV��g߄#q���,�2�
A*�3�*��s��q��]��[V���{!>���s1�_�LC+��km1�o4�oO����!%��n�����������Sb�чZ ��&�BP}��)�|����^��?0���JXf	K�iQ����4�[����b�)Q�s�(�v��d!}@ǎ��Jo{��"=�9T󔔜����g�`Olr��v�Io�bp1<�q�T��P���3���ME������Hv��+4�k����C���D�OT���ڦ[������(p}fC6�������\�9JI��[�m���O��({A�{k�N�b�����}�Sj��34�OE����d��;�G�[�w���~�_��Yx�����ֹ�`������g���N������*�4W`��� &���ƞ�D��@�5k�IP��'.��bQ7��1b�Hź�G_3i*V��s��S��ʕ�����HQ �t�,�q^���鬄 ]9��BX���΄�� sJ@�'�o�ٴ��b�;aw7����>���ߘ�k���`"CP�SG��rO�� �[ꓽ�A�!��^�>�����~1`�_��J��A��.9u�Q�;YZ\���s� R!���*�'X~-Ӵ�w�����=��J֞�0:na��/��C�ׅG��`���%v���y
ɛ^uH��c�ɔF�&Á��W��w`k\^)��8��u�$އR{����jz	�o��[8�����^��C�n�(0j��X0J�诈I�&�HC-K�Ȕ,όM;;X>1vC���:�mu�Y'$z�Yd�m�3{O-'*�I5�w�@�=xZ��[|�j���n��%�����$�p������a�t�)<��G9����pY&\�����cqcg�zA���a�:�n=ԞW)#1��X�P�	�p���Y�����M�&�0������s#��Α}GI���7�è[��DY܏3���1h�'j�!c4�
�"�����r��Z��� �\M�Xc`����R�����}]V��¤X���$� ?���0�c/iYV�>|v����O�CO�����6�o�fg{O9�u���%	zc�C�9j<�H#�����uj�?K�J��vl�7������8SNd:���hg�2���sYwy�6��mCG�J��5T��-�ё���٬���E�7ⱹ��
�˂G�hhq���C�e�c����E�<�b|γ�N�z����#ǂ��P�K�ޝ�B��ٴ�rGy�A�b!i�4��<�L
�mGq���_��� =�V_�})�f�=�/��)Jt	��������T}t�fC�`�jǶ�G�$38���_�`55爽�+ &����2Jhy؆�?�Ȇ���UG�����ԃ^M4��`���Vc�8���	����
7���,2�g�A���B/������$�� �h��Ax����� ����I�2��\��H��Î����[a����]��r�)(~�5܍裕�N�`!]/B��_ȯ8��KZ94A^�B?JЎ:A�tzH�B�(�� �ݥ0����t&�<�WB� aY#	� L	D�{.Eg"ܠ>�a<���*��R"�`p}��B �g��B� <F�i}�+c�5t��/hQ���Yδi��EnΓI��e�YX�V�2�
����|P�`%D��I3�Y\��wJ5�]�qJ�Ք��·����ۗ�ʈ�9o�����m�(��@�	҈��_Il1Psƴ���U
a�����+喹����t�`�:�r��T�(�ځ�L,z�K�٬���x�hDYA����T��Q)f{�қYМޙ��&@�a��t�(ŝ4���W`x��-�ɤ�Uܴh��t�uS3U˳=�,�j@s|��c'Tz�&�F�L����%�La�a�b�	�.�ZN�.��Ʒ�eI�%	DQS�x1h _iLi�V�1ؿ�r�y�-Λ��yiiʞ���xHO��0���%(+��#��F��v�a1�;B�yڞ�>�	���,	�r@�g�&�eg�X�S���ߎ0L���n���q%5�K�q:��˦�O��-1-?��!��ݴ�j2I(v��gA������k��t4Ś�$�<��0�Q|t.�1R��`��[V7���cf�<s�h��4��1��d4�ϻ��k=ޔ�k��7�_�NW��#�Ɏ���F�n��ʭ�8�����c�Y\��*@*��2h7�PY�	�|g�~[J �~�4�[��d����H�ULD7�U�Y�~�nl��Da)���L=z�Od�c"&�k�ʵ���h^*W�\b�)�%B�h�'?�I���=z���@�ć�LکE�ס	�ǵ���a���ѥ@_�Z~K$J3�@J"�v?L~��:Ϭ>��A�9N�D>i\-�d�_8
������ 5q��^;�X��BϤ�J >����е�R%��!_��:�W'L��r�pKf�\�3�l������b��:�P��a�T�c�2�a�~<�oXJ%��2V����U�k�Ep8���)�yB�	o���]��Gn�J&?��/E����ҁ���;���r�x�Z���Eh�P�i9�$����9�PГr��=x�Z�@��}�5�U�Y��)%�3�~$Isi�dޖ=(8x���B�g��L��������<�yIX'�O�Z��s��CV�(��*gP�ǐl�@��y�kJ����Ӎ��ܚjr�A�� p��6��Ĕ���K��,x*�k���s`� ZJJD}��{M�~Q�c�����R�@�A���C�_|�<�5=�A��x�q�«�H�ں��(7����s&�k�;S�@Ez�1�����
O_`-�0|��ֱ�
��QX�k�-�@g����Z6q���K��"JK3Ajh��N(Fd%B�%O���j9�[ۥ�ߋߴ�ٞK���}XY!��
H�45|T���^�g���!���uzX�B��7�";P6�P�z�	�{�t���l��P�|��G��w��pw8[���̞Eu��3�իv
�EN������
OFVi�)��"W�im�E��ek_��}���(��Pa�#V��;th���#�Y�1ЙʉYm�2j�aC��\����j�ʫ<��������f
w�V�p�0wڗ�RWﹶ�����N���Z�9�����ƍ|���K~P6"wf5>DU��^[�ۼ4��Rg�Є�&���$/�4���D��j~����bz��ixM��L�{�s�$�ϯb�LP
���ǣ$D�b|�������b�/.H$��*��¬ة۞�Ġ�y�2t��'tQOi�.^1��(��BH}��g'�:XE}ؤ����q�7gH������/���n�s����$���Cp��\9���n����
ؓ���k$F�Ӧ�N�~��@i��c�}�d��<�l[?�s�!A���	���Å?27�7<�X�k�N�C[��� ���q@��&J��1�-�$�~����K��w!z;Qk�X�.����А;�D��=[��?"��8:���!z��fi�E7=�#���KCd�R�-����0���iN6*�����E�r�+䝥����B;z_=��΢��y�JD��h��6�ҩ#�?_�y������RF+_6��7��.[��[[�U��ʰn����I�\h�&Y�k8���0�f杜��4o��o�Q��ǫ��T�f���e7�n�k�͔}�ȷ����Ԡ���R�Hޛ�s1M0c#�q9�Vg�ۯ�Pf=�[A�!	���E�`7����p�� 25���]c���J3[��,��tl�qg�������wj�'�w4��c���5�cޯ_,cǆ�'��t)Nc]�MA�}K�W9+�E\R���v.�yË�	Y��|V�V�񬢈]�	��!R@�Ě��Pwf�B�I�;��N�E��?HP��`�2�{���	��c�����KS]Zk��Z1u�\(%�xU.ޕ+�?��5�40�h��xo�k�Ŕ�O��u��(��KSb�W���?q/~bS]�)�<�U
���i� h�5��o��H���
,,_��F��v�s�S
1�I,-nM�&�8C�����K��Y�C��tK�T�2��L*ڬ���1�T�I�eS�O�s(�VS/����>	�Z8���`59���;2�?�Hs�ӹ��x���q�\�1/�[F���~�@����Y-%-�zRoz�W�?o�%!= �C:�6p�	�v����yٜ����v�@$�$5��,�2�7���L�૮�p����y2��E54���U,E��p\�&�Xc���w���#V$�Xb%' �;l�d�I<���[rx�Èzo�}E�8�r/�Gꖃ/��*1]����E��-�E�B����6_L������:��2EW!9����U&��]m��=���o"��^�,�W� �I�ps�0o;�ך��0t���������k�����y��dF)<h�
��P�H���X�i�T�n�'�/�7)N>���
��D��>�����lo)&>�v�y���«CG�����y�	^q ǝ{$��r5:2*�/%���l����C�$=�?	��3j}��g�1�0��'�.���f�c�T��P���o��`bC�?���<R���3!D(�ƐQn��^�`F��k���#�?�̽kQGʌw�Q�z���ru��֟��J�@5^z��S�y�7,9��`�Q^Bƭ�y������U"\��X��tX\��L�B;":��Kp����-�8B/��On]HI�L\W��uO�]��m*0fJB.�K-���/4�[�u��VQ�2�N;�C���_�[~����S��f��O�g���Q^ፇP)UBz͈?����	ۖn�4��:�v@o���jĪ�z-
ˉ�9�����
����g����S�&��zs�����0k�>���af[`ІbA�=̝��SҺ*��CI�=̪\7��H��I׬�l�Q��E�5|`��1��\H�{��|\��|΋e�𐭳ܦ��� O�	��ߞ}�)�����|�T�yN5H(��#�^Q��T	<����#[��B�KӰ�eh�S�����&��f�c�2D��n�f<�r�� �n3kŅ��n�-
�z���)c�-�P���|yd��NڑVQ�>���h�8�vcy=����|�BăRa상.!��`�#��9�	�2�l0˽*s��V9���ky�@�,qV�8�A���+0�D�M ��s�>K@H�d��z_
Dt#%BWPl��Ȓ�U�~���Y5&US>&���	[z�*� ��_����)���d{f	��*_������d+��7+4��Ki�ݧ�E���]�L���'�0d�C�Q_|�bQ��he���}�;�-[7�n��ˀ٠��q�����'���)3
5�l�-��tAW����T� �-֙,��.EtwE0�U'>awP����=�+4���%��Sq��q���Ef���&�)l�_��[��V?p�!~֥�?��h{�6��o��)�7����g����?�#f�1�|��ɘ�d��\�.��TdG"D	[^s��E����r"�����};i��o�[�'�"#�4cW�'`��<؝��"t���xU�;2;�A��R�&��3�UKmh���ZY jyٹGR��q�<p�>g}TĀZ�����|�W���ʠ�W�_���t#��^�ĜS�	<�e�gM.�E�7���'3̡dsF�?�l����2��� �Lÿ�y�ofX�X�i�$�3�P��nd���t���Ů�@4����7�w�_��"d^�@V�Xz/H�k[")�k��c�c�z[���N��Bw�-��=galUg��f{,Z�$}�\�*���/R�	�c|U}Aa����W���,�^E<dfC�W3(/�Sy0���b�Sqc�W�F�N��
����d�x^l��d�p�E[QT�wgc��Q�4��z��A���$)3�~̃F0aaR8�!ޭu����kIps�9��}��}��nʆOC�fӊ�O�]�mX�Իxw�>�����������U@�[��!�`��QGQӶ�us�]R�l���@�k��@��dK��B�g8Z{"�?�޿e���*���V�Ѯ-"iO�.��Tݏ�� Ri��nR��������#
��J�,c�̵3�Y�gK�5���uFUw�� ���>C���h:-f��\?��C�K��Ċ4 �8�d$W�z#W��ۉo��VZz��f�U��x3��\E`���~o��9|���p�rX:Y�G��?��K7�@�	�Ӂ��'}2�a�w�C��9�8t��쑞x_O�t��
���hA���)d����EI����&�L��X�"
����R|
�?���nr	)�P��}�sV�B�����A�E޷@��tw��a1�$����u����l��OR�`&V�q�����ۅ�A��đ(�ɔ�Z�LHJsh��`��(�D�w�C]_:�S:P���1#:�^$�,��h����,�j��d�qy�%���c���A�>
����<^��
b3<�G��ڏ=S�B����E��-�중�5���G#�Xo����v��f��R>�pU�E��%Ǆ�+�LMa H�(�ݷ�kS#՚�!��#����nI AH�$���C&o�M�*��&n�S؝0�Ku�o��CC��Ҕ���"Q\��b�cG�=�^����܀B�μ�q�f�u���:=�'���W�q �$���f��C�%XC�a���'���G }RL��w��q��Q"!V�D�QnS��b��y��HFe%�ʊ ��cU���_���f̊u����IIl�r����]ՆT�us��n�/�0�X�����vr�\ê��!�m��aV
�w��3���?���ǯ��;1�ڕ}Θ�d^_�\ju"�\F$$�&?��.��&!V��#�1G+���>HR�����	�����V^Dϕ�lVi�����=�B%���9U�����~�F�;�����'��-֙�J�!�8��'�Fό��Oz�"c�Yo@����ᅫ�������Dn=^jXl���g�`!l���A�=����m��[Jj����y�}�z�I�̤nS�K��G �����=y�1�U�	���&�wQŬPֹ~$�]د�ߢܘ+����p���#��?���|�W]m��?�b<�H,��.?{~Z���0�4:�����:��)UM���5�:��a��d�rn�����*e [J��V�n��� O���]��ՖX\K�\\����@o'�`���&�b�[s���շ[��2v@X̴�N����T|����?��d<���t�,�3��,���|�FT���O��q/�'�e��e@�e3P�j���$�$�	���$�y\ �����Z��"Q��5xw/�Ȇ<�d�=�;��5g��"�7?�\\�������T	�Ǉ�H<uowp�7�U*7;!���faH:bG��G�N*�<ʊu���N#���,����Q�̯��D�zYENo�t��t�pH|>H/�0 ����ȁ�X��π�EƩ#n}� ��Qѻ~z�Z����t������`�27>>FX��B_S �q�{k�y���?ڻ�"+�X'�f�`(��xA���b��/��sxC�tu�� �w\K�3X�v7I��������mkk�g��v�Wb���������nB?�J-�AV��2����U�u?$jtL쁌��H���d�M.]28:Ð�o�v�! �/�
�0E�׆�[-ؠ��
��Li�[xZN;S��>�*�%w�Lޒ��V��FHٺ���+�1E�}u,O�5�%�8�x���Ʌ�vQ�0>�G�`~P�3&�˹��k0�����9���<]W0��z�-~��䆴�vƶ�S��#��Q������u�����@��L��@�o3����C_�Xy
���w/��_Í�jT���<�R�q���E�H���_�?�.ּ
ߔ�wK� �j�qT��=g�54[}�O��(ȋ���3.��]Bqr����`nA��;,��9�d5�OƳKA�YV�����f���_��PT5Ԙڔ�'=Q��l*rZ7���W�"���o�i>!�
���aG�R�v/�k��_�G����x�H�A�X�����x{�����:�e�����w!�ů���������mA�+X��V:�%�j
�0�ݲ���C��3%ɗu4w��\7��ˤ�S��.��R���[ʡN�縉��2���F�����j����<�_��ñW��&�8�%Ҽ��PKq��:E���Ā�%N�2��l+�����"1���Ry8�΢���ײ�P�{���l�f8!'q�#�{;���Bi����\`�E����6���G��#g���8%�yqZDɋ�I�S�`��_s|>r�����w=��ߐ��m�PR�O��2m�A��.�(�j\���we3	�?Ι7Va�Ä�d 1�x�i���"%�D��Z�%�lٽDD���dSK�#M��q ��S^�9�e0�ˢ!ի�/�>����i��I#c�#2'�Z�3�y����t����I.ؼ-$1�{�pMV��������1�X�j�E�����Gu����-�
��#�r:-�R�՞�3N���[�G&c����hzC�a�N����Z��q���]#dT�Ō����@DǄ�,�/4.����	�5��g�dW�zσOl�?gH�+��Ц��_�L�S�I�w
-�NQ8����t���Nw�X�/��(��_g'/���`祀@�;:˓o"�W��o˜;�ٕ���LE,ʺ����_��hb�\���.������J.��Э�p~x4��m_m�$8V걐�asuQ�{EoZ�~*��\�3@,�z?�<�&\�S J�>mQ�~�;�9��@�~��,6V�����S��dz�G�߽,U��e~8������ZH���ܬ�y�Pa8_�p"r(�`��(�3��R�U��4Qm�;�\�]�G�&���И< W�]��_Ь�`a�m,W2@� �
��]���'0
4����Լ)��	ԗ��D�7�RN��p���3����,3� ��)��Gė4��@�W��=���A�&�Fg^�b	��Y���tZǴ�zL	��ݐfh?̓9 �硻�-h%Mu��ͬGI�-S��ut`��T���ʞ䫞5'.ש�LC�
{>��l}��1�8��{�v�~6�s}53P�G�������$X�����S�
���O:n�� �������� ��X��jV���n�Ɛ�mh4�`�ܮ�{�^� �a�����_I8$&R�9��Xo�QR��j�7ɽR�����hG��{PvX��|ب�`��j���<`�$�3�q2\�}IٞX����E\q���2�+�I\T�F�#I
�����j ��ҝ�D���',4B==߹?O�_&�2��*�e*&�B`�1S�1xY�f�MxR�vP����:oo��x� �&�L�e(�ʺ�'{C�0�4���m��!��\l�˧�G)�7Q��è�CW��7a�i?ۂQJ�����h�6���&)��풳l��6Ŵ܀2��a ��^�t�|�u9Qk(E�\ v�T������C��ׇN��Kn|��Eο��� ���'�P^h'bkّLl	�Ͳ��*�r#f��������l�[�ȊZ���.5(�����o�T4HI��	dp�W���� �u� �DDs����Kōa��J��:L��-�k�&�������J�ߝ��FiYG��|I0�3�5;�%�촌��x�y���c����ZD9^���i���'��i��H˗��=),�yͩ�n�<[bj9����j\|Cԝ���@KJ@:7G=�V^:�Û��F	��A<���D�[������ǯ�L�:�䳢�������'C�0 #�/ "e��E2ф�f/3�|�� H�?3�B��dY�J A��#������46��I86���j|�^������^��N�u�$�n���_�SK��MݙY/xɘ�L��ڐky\������O�4�B���S�C�jx:x��=���>��� t�����|9��~���޶ڌ�P�l7�#���G������ 2���Ź���K����t�-3�F�M~	F�l��5Ӫ��s_A^y��77���!o8y3Z���%��{���`Wov54M�o��h��@,933=���9Z�sz�����(g`9ʺ�nA|�J>ؤ���\|z�����Z�Xn���{���e<�S�k���}ѿ%5����I�9SGM�N$A�*��\)Ι�D�T���4��@I��bȐ ��ِ�lV�Ѵ �\�t�j�8Ch����iH�"2���A	��?��EB���+�|&�%��NbxR�!~�5"�tQ�;@��O#r׭D��+��n�@�L�����N�N�ʁ��K���s�	 �Q��gW��$خMz��D�;����/�uFΏA�Xz�fq�[ >UP���I*~*s�E���RkQ��rqƸ�y�Y�>[�%U:����ˌe�1�7?�U/��^�+
̥���&�qH��� G�����ϼF%��c�U_�ϼY/l�q6j��py!�t8�x�����۝�T���������5.1�w��tΟx)Fy?/[?Ё6����a���	�h[- ��ݮ�+���LY5$�� jv�Sc�_��۵��1o)>���P�ļ�$,��x�+4l�Tz��Aj�=ɣ�L7�ʳ��M�ğ��:#��v���[�N�0��mKY��ro��tG�e��\Ž���p",�nj6up�$y�²d�H�����_��4�GhuNB;D?�^J���֫	��@s�0^iP7H#c�jHD1�l``%%�2Q6��tQ��8U;
��!V��3Q�a���eU}s6W�+��?��f±����[�8Cs^]"rH <��O��U�#���$p=9Xd��PÒh�	F=��mL��n�����>�an%�ڼMG�WL!!���7�q_c�i���N�؆�׽�pb�ݓ���x�������y!-���Ҟ�BԝM�?Z���-T���<-��kc��ם����~`2�n�M�V���4�Xz>���V�f�s���D�K��|z˻i�:#�}~��LS��u��L��.�A��C֩�cA��%5�h{��q^�
��@�"Rp>�N>��D��]J���!:��E��T�b�.�ù����e����`V��׽����u�iQ|m,=9aԌb�S��PX~�`&Ծ$^���?���s�8'Y���(i����$�#@��A�k�K�2��>1�������T�k �-F\4���
�b 	�Jd	.�Q�؃\D.��ο�-�@����*HbI��ƾ�1�T�ͨEf�(�� ?5�*^.�iUʣ��a^��� xl�^$��|W��dܕԾ�y	A��H���F!���fݱ���Cn-7ߞ�Ά���� n�vO&�fBi�Xm�e �O��!�B��Y(�Dd��-���b�!C!���߰Gh�ߡ~���c��ڹK9��&y@R��"H9�>g�{�u�7t�V�#,�=?;&˃Ɣ,c�V�l�}͖]�R5�{�S�U�n?��CI�u��ߨ��ۯS�26�Y�Hm#R�-����cƈ�¾�l敢�*�~������v�1���"��o�=��E����:[Y�9�� ��ùG�������{�`����(b�g�c/����J5�Bh�5y��Z-�'� K��R��^��E���2���g�O��S���@?�`�d���X�5�yޖ�.�Hti��mW�M�^Ք�TB��VA��/�o��!�-���Rf(�)����� ~��U��.\��@h���,y&���h��ku@~E��h��ϡS��{���B���yI����Z���l�a^�F�,��z�Y���t��w�Լ��V���X)�t����M'5�6p�����,{�*��eԗ�k�O?yr$e&ت��O+=yMctΥXp̿�2wTT�o�&-n����|6���2"�����׮d\ܯצ��W$.Z'�Nl�&�
%���K�i��irv��=���]J��g��c��㶅��'Gqx��0YB.|��j����u�<�m�PF0`U>�	/%b$�R��V�Eٺb���R�*q޾���X=�ſ;�� p��U���De7�"�膼H��~*T�I]�e9S����itU�61���5�����^��Πj£�bU����B��Um��F�^[�f�9�.z3&#Q�&����0rbp��Z3w���%W0&,�	h:��|8����r���X�=��<��|WW�9H��6r���@Ʒb�0��A��KEdB'�
8���Gj�N�Ng�R����p����B�߁���)7<��<W�ן��ް'x�;1ָ�Au����e�f��i\�>��X0n���R._�j���#�T�z�i:-
��{��r�0Π����F���ۡ�W��&6|���:�d�ϣ~�H,�Ss�)�pՅ)im�'�C�K�r�c�
Ɠ�E���+�L���k�El�Q���zK�l�U����!#�O�&�g�����/8>��"۱zR��e�:{l0:� ݀i�o?s����ځt�a���:��{�%�lxw��k\�0��@�@vj��������Fć���gz~��C�e��T8�S�_v�v4�BEE��������vW��G��T'w&�9H�8Q���za�����G�פ%72�[~H��]�nǫ��������)�d���w�7	m=W\�I9�B��J���,�}t �ą];}Q������	�Oǻ@l8��JZ��TB2ܝ���%7s���]a�a�"��'�o� ��U�D�-��G`�V����D���&���Dn����xò����5k�:ۖ
���Q�����F=�׾W\�0���Y8�-7�M����i�-����(�YgKHAC�(,d�B�n���+aU�|J#�����"c��"���A�p�'2�g��P�G*��L��xO�&LHi��}m���:.	�0߆ ��0���4�C�RR$��Ҥ���C�#�O��/�?Zvv�s��!�i�F��-�RT��ݍtc��)S�C!�ob��<e��p��~<�Kf�d�tsH���@<���+C�_����xE�P�FAZb���Z�3�Ȏ����/���U�uw��<$���1�����@��n&�g�@��Up�ˀ��'��*Vc���`�{"{��6ba<&Zx��B�?/��Wc�����N5��T�*�Cj���>�g�k"*��O�J��� }:^�*l���<�>���왃�T#��R��M���Tk�"������(p�\�`�j�!S�T .����E���i0����V�a	=冪ZQ�����ru���̓�I��t�(�N~��-/D��S$��@�d��I������"�Lζû��r���%,��=$�r�O!�Li���#R(��lX+'��Z�v.�ډA}�����G�\J�~�-F�����h,X�x���	��:�?:8~ٻ�\p	���¬��6B���F��R���Tt�74�rf*��.���©ZYGii�y��dExr�i�{:�|A�y��>�A�n�w@~$ؗ��p��osxa��C���������3�%�¥xT���L�x:�Uv�q��U�ۈ�@�x�U/O�MgV��"���X�ᖓ�����+C��pQ���((ƍ���8�Z��[�|�=�t�'���.#��P��:����;��_�G�0����@���d�|�&:�'&��}��k��['O�ϗ�����ʕX��J�L���2��Ϡ��o�tD���E�yd�͈�m/^7�j}�@��t<��	X��m6��?6D��Ԕ喦�ɩ4����9��
^���׬��֢_H]�t�xf�_��Z�Cu�z]���X�y
 K6��n��,&1>�#+��8��H���T��gAY�G�w=�����|���B-$$�h�kr���
��?8RU[�u���ᕯmd��T��z-`	�6�Y2;�|��#K�R�]�����8�*��V��]�l�rr'e��Z g��юk�I��/�6R伆ZD���W�JX�4PF�j��awp�@S�3�<�k��6��;w����-V��-��]=ɸ�G
Նn`��<Q��{җ�u���r�NS�Ds�����>���x�uJ�������p���2�����Z�婾H�ԃz���g� �]^�@w4��zQ���x`��b����`������{gd��.B)���?�f��a߱�g�pѾ��zojj�^��0>� �p] I���z���02�.�[a����]I��0{��Yࠣ\���8bnP�Hqǿ�#-%�6���1��0���Vx<~H��C�Q�AeZd����F����;B/4� ��ir@P��E��d���D�p�C���v�A r���4��j3�,^�&T3�z#�At��-R�v��'(1�-(��s����J?�_3.�f�X�h��N{D����s��]	��s�U�
��s#���/'a8���p��B�����G�̺#���PF���L��z�4A;.dA��m��P�Q�u����;���������]=;ͅ9)�Q�79��W���֑!��H{ѤW��uc�b�u'�s�`���AFħξ�Ɓw�bq��>J���!��	�8��h�3$�<2V��8l/y>��R�(S��]t�MlsS���1�16��$ݲ�:h V��)7I.�9�燓�H*_�z�T�߸v5?�z�H�c�t(��>���VV����$���O�S,۲�i4P^6+���	e���k`�k�=�����Iy!�8����f"�QP'Q�}Uwӟ2�O��*�W�+ߣ�E eH��K��R_;��ӱq��s;D#u�]���I�����?y�<'�l���
^�&0�4���[�ЦA|���z����n��0"�����w������Ô��B O	��ۅ���C�t�X���7	����oӥ�L.�*��!�`{��h�R�CCdγ��v�����>�t�o��fܣ`LL�;%Y;s��.�k7�@#�`e�`r��l7J%зҒ�Mx�������Y�\� ��fms�"3�IS.�Ҁ��@ҭ$k�m��6��_ ��jk��&��@춌�n��aj���`q&W�����xnz��h�w{��7���V"��������z5b���Ʃ�Ѷ���!�O��;��(�30,�\����	�a�����cQ��������Mi-�^�/�\���>�H��0��c���dp���� R��8�u��Tͤ#{ڞ`�f>I�v�̅���В���J���!��y�`�|�f��7^�3�9��\���&��{�_����A��9B��0��3�G�ʊ '���Rh	��D����}������r[��<4+�g�&��(0��;���<댕E�{im��j��z���w�$u�M��/��pun>�x�_��?v0d}������N�8��|�k�ݏ�9<�٫�������Y=[p˕�ܗ�%��/��e^�e��N��l�L6z�7L�6WV��
cƅ����	�F(��(��;��8T�lH&���W��ӡ/_Kݚ�>v�J��`��Lk�x��a�*K@b#�h�(�=e�̍|y���gf�C������\��	�&+�.e�A���W��,*��L��Fa�Y\@�����&Kk,�c��!|>=�kE�/�nY��ꅥy���p��P�NȤѷ3W���6��RG�7D��	.�f�H_#���13lzCk�|��C@4[~�خ�����Q���Z&옡�����Q:!�@@>�K���M�d�#�z=&���L�JQ�NgYn;��S��@>�G�A�3�l�uO���T�+��w�jfۇ�!L�5>��Y�eb�`9�8)�!�!Zi�EM�"�mI[?[ZP^sφ����I����4V�Fa\�We/��$�t�������;7�i�&��J��"�a�5(�������e���G��sVd��2β�:<�-�Qgm�N)�?���$�oªU�����}�^���~�N���J����"�QU.�zJ�U-��5�WJRՆn���dAv��G���6s����u�ϩH}��,*Ұ�ç�;���\b#��������Wݭ���:���������4���%ec�f��-�$���\z���3�VE9��O�����\�,3푽3u	��ם_��'r�ad�>3��T����"�x��������(�+�vF�w�h������[���,|���u�X,������|F?�uqH�����Ԯ��7j�vep!�v�Yft#�5����Tq�fe���b�zcJ��
L� ���%7�� ���uID��O�\I$(r�b����;�aCk	�x:�x|��>�؂~4�)L���O!nH1��˰ؘ��c��a��O8��31PE���V�mn�҈b�B"���D�V�57�i�ކ���i)�<�!�5�5A����2b]x��� ���"�?�xt��:��2�Q/��7{����&f��[�B���!o��}��-Z�xǧ@;�V ��8~W���k�[�n3}X�t[�A��=-0\���##ֵK̠���p�y��p��֤�J�!���#Z�v�)&���&K8�x"��	��4�(,��A��_Qt�Ox$&m�.v�K #�h��^���8G~�@i����X~ލ
�ˊaC�Aq��u7M��JwG��*�T/���ޟu��v�Ę�`�;Àl�&�>��}�ǧ�����6�����"O6�/Z���A�I��V��w����N������vq�IMJ)X8��$����8ސr� �&�o��Uܞ{=徚d����������̻������X�[��'�NrpL�C.���z)L�p�q�H���o>C�Qe� ��1#'����P܈���g�[R�>��`��b�,�1K+��:����ȫ���Vh$��A&�
�n�x�6��U=�_���9�f���k�$6�\MU)9G�N������z�7�E�N
�*T��^�T�dG�N�&�7��%��Q@�ک3�gN̂��\9͆.|� Ř���/�Cz��>�j-yZ�U��q�D�Q���(!9},���F�X	���Z5�Z��Et�,�K�:'"8_]6z��TE,�.D��Gku����u���8lr��V�4����B���p�W�OV�i3)��n~��\Z��ʴ)fj���&��<��/�u���S;@�s���P��7��4�rr��K;�`��;\Xx��{	�X� !��}t�ɔE�+��Эi���q���vV�C��+���M<��Lв�x�=���4�k�?��)e��eВ�WŸ�d �����ņ
u�o<:�`V3��������" /{�'y2���f�YZ���|O�x]�"�E�^ˀ�f^CӤ�^jE&A���;rl��@���y���<�%��@t���)��4��E�uܔ'�]�^���U�&�1����������Ud�S���nC쿽�[�XÙ>��)P� �ݒ���&e���U���9e>V��/c��m8�"�Q��dE2�ǚ|�b��!�?5=Q1�8*����K�8���y���}H\��kPS������^O�C�!�-or�)z�1��ŗ��U��F_+%�����������2��ԇQ̽&��O�3�!�F�(��y��}������M��Fiv(
��H���^ܯ�*�&��FMy�hno��'R}�-�rw+-���u�T!�p�k�M������/P���&L=�W�E;��x���1��k=��m�ț�-} &/e�U�{�Yy���3���)�Z�3`�fa���|��̀��9���C���@7�QI�&����SL$lj����w�jA�K�+*~l^��b�}��hB\d �K�4�-�����J�rG�Ɣ��B�h���D�=CGaJ6��1N4K�_3WL�M���a��oy�c��7Yo�2+�l�!�E�0"L氒3�q�8�}�>?�Cs�A��IyͲ"⚲��f���Nީ�l�C�'�0D���������Q�6G�?��L�T.��8�GK�Ǡ���h���iR�l���n��fS�Bx���(&6d��V��.�IU��V��%깽�U�Щ?�`\�_�Add��>���i������j�1>�J'�z2��g@����:��R���$;G��:���`_`�"�&ɔ��ȘXҼZ�93�~Y��g��xL�i4�l�Ņ-+'�Q�E���B#+�Ɓ/�V?� 7�k�T��n	�b$�c	�-F��*$y%L��W.��)��V
X��cju�i>A ,�o	������.�b��L�;�*�5�`�4\��eM�얱8��)�&�+�����ߜ2��i�"�6����Q�P/�L�mr�Uln��M�6�yT���[��3:zP"��!4����$��6��6��Z�j��ƥb���Z.���i|��G�N_��j��[��}��D�6�KX�S�2
���3.If	r���y���8�L���AF32iV�3t���i��௖ӫ�;r8��rc�3ړOq�ԝ_��^�C��=%� �jS��I_w�$J��"�>fv-���%:�P'��J����U�.p�O���ik��Ҷ�Ţs��WA1�k�e�"0a����b�qq/ǲXP^�)��x�h�Ƿ���z�OȒQ�R�9/����y &��MtP�&;�$u��}3��;�n?h4�_��KRD[��R!��IJK����3E���e��$�9�+�!M�[��B��J��8W��d��Ā��k��oj�|Uj���ݡ���׈�j(�"��I}��R�pP�G��&9���a��u8z���t��h�[vp��XWD�>$�/���-V�=�H)���l�f!أ�O[!dG�^t@���,r�Y��[��>�� �2 .�!|�*tqh��K˪�B@�k){�F�����en�B�5+�A������l�`�*LUdS��۞��^%�4%,&�z$"����"Z#�d�ֺ[E͞��0�B(��uj|�iD峒��#�P�谼���S'n�Ŷ���.��E�!��v��
��� ��ל���F���]�ĥdf�L�~b���N�����+@�7Mɲ�����?�x`�Ml�<*L������O�C�XX�Q�6o����%G�ni��Ey�,��Yr�"��0�_(4k)jo1��}z+1�$¼���h)@㗉�&(�LK
P�	,�5qt�h�������x���	>χ�!f���2�D���*�Nj,��0���)�TcXU�3�I&"����a���v�H�_ ��m����/�i�:pa ��H�C/a$pCQJ�=u~$2R������\3�[�(ϓ�1��_�2ӣ���+`�$��O��U,�.\���w�f�a���J�
Sfi�B�p\u�y�������ݐ���z:�zT�2 ��?P|ո��!���I9(SF����
]V}#�h��,T�����Kj�' �L�r�W8LA�ݫ,~��[�@���0��*e@�!�B
��Lmۚ%7L�&������t�yz1��C���5[�;C��_��au��A@���מ�ѯ*�ͼs��L�u|�_�f�cKc�w�~�m�C��ω���ޡ3�:�����n�M>��0�����<�ħB��ʏ��OE��4�09��L����rk3Y��Y\P��,�j���<�ǉ��W�_��WK��I`#�!ZC0�V� �2�r�?̲p�=>�g��%Z�'9Tnu_�;# �WO�2=�`ws���mU������Tޑ��
Cb,e8��P\jn�/B{�M'1
x>�*#��Ӊ���}�����	�͟�y�h��\H���d)t��c�'k��9�g���Z����pO����^ɳ&��#;��Kk����,���m+V"�1�w��U����X������m%�sL\�@�>�t�ԍ��}�H��(5j��|�5=h&ľUճ��G���D�9��~a�E�}*�����G���m����.�A�3����m��[���lsk��[�4��
G�P���TG(�f	�;���T��؎���tT[��Zi�+���3��s	}�Hz|ˬ�����>�f��ǝ��[��\4���:6��nY�N5	��d���:����<���,\)���CO.c��_#�T�4��S�Zu��&dPb�9�vi0[�Հ �ͱR�G+���/o�/��,ٞ�V����&�!9�����&5B+��lE{>H��Խ�K��D�}n�~V�O�.�8<x[[�h�5u�6� ����j�_s���[���,-yD�y�ө)�1l��α�����.nx\/ ���`Z�5���]+}�e���|�/N��ū�v�o���=_[�xRH����tĚ�	nn�s'C!��PJ���$�Ȇܟ�nf����(�֓USt�)k��iPMK��|i� V�$P�,5_�Q@:�S��W< ��'���"��>��x��P߿33K���ip�˿,[fw���A!���,���T<�.:;�b���C`ߕ�K�Я��[�Ru������Sj����t��� ���.5�S���3��]��sUN�֝K�D7�-���-�gr� *Sj�ݿ��Ds�:,~�z'9p1�R�Mx(���!#Z�A�D�Y;!�=�� i�	�W�X���m"	`����J��ږ�>��{��]�qWw�*�1�Q:�o��R/8ˁ�p�fj��
M�-C;�M.�.$����IG�Ae� 5R�Ie�4���*"�,8mM�x���"0������X�e�l;��:%6�������.�Dz��R5�Ru�Ls��e.�>+�e靭6쥈�h�,ڷ�!�{�6r	���?��d��#�dE���_���%�+�4nxy�a������"zG9�-�ܗ`�97<�ܥo_`���o�87����￙z���Mf�WSC͙���[y\����I?�}��Uc���/�� �#��!2�"6��m1�@�V���=㓊�ؠ�q�p=Xֽ/v\JB�|��O>����мoX�7�DގC\O���K�[֥y'������vc ���o��M�6	�d&�W[L �X%�hj�]��,�q����>:��fnb��3KG���	%Ի�n>�Wث�J�l~��2G1W���Z�*qr+��/���nƵ�kS
B��K�j���П*�[�E�b���o~DԃL���>GUi���Rјp�?0���I0�,M��vhv�Zi@��/mpӶ�,J.�c*����R7�F^Ez2Gn�����^���1l� ��U�3n8W�-J�׍TL�`��}�|�Z��'��m�[�q�|��v<cD���hMsRf�v��
��ͷWB6�L�2�k� ���q=��X{���N�E�����?L����C��(g�
��G3d��n. 	(tXj����g��%wgB��y� j;����B�y�I�I'�>_&M=�������j>�85ꔿ&}�RB��T��(��el�3�D$���6��

گ<�rnM����t)8�/?{���#�_�c<3���'��B�!��u��aRx�:�2 �9ly�L���!���*��^��l݈�4C�������4� "�R�p ��5� ��+���c�w:f�+@�0�`��E��=�F���a�ȹ��?V��j���-޲��rЩe�*8e�c��?�MwC�A���+�n��O���kȗ�
g	�g@d�r&֝=KV%ѭT%}����Ҳ&�B���@Q�.Ҍ��������jw%{�C� �~�
bMZ1�x���t�얞3�Żq*��F���,b}���6���d��\���� f�N\J��~1���NV��.Z��:��\� -[�i 2�i	Ys����g��>)$*|����B	-��b��b�����L��iGį�8�lj��R̾�[��Ud0/�I���R]ׇ�?vh����1�ƫsY�Ǻ�':�	H�'�O��WM��{�ʿrs%����Y%��H��CM3W��?�.�W�M:=x��B2Q4�)�0�Z�HY*ԶWr������~^�z���&�W�`�4o%�  ԊT�%�կ��������۲oA����h<\�θ�<1uw��k���g�JŁ:��2�R���F$��k�f�7���ⰸKP1ѱ��B����)?�*Z<�o։�&��ؗf���F�vk]tS\�u<J���/B�rjCU��~59�.'�6�@���>i�m��mڽ����L�@����6h|r�65i�d��X>1�1e?J�1z��[3�dC���r�?s�]��UOH�����e9������J1�&�H�_\&{��ͬ�@���2�'�}��/���V�IfԠo[|=ՠ~lKtsnT�F�"����bL��2�70�{�����A5u������t��_9�b���Uf�ю �~��Uv���r���R�����_ˮjM����M�"Z@H��+�ގ�P-n�?��q�/{��l��2����ɣ�-T�\'����!֓F�Ox[�,���g�H�#]񛏈������	1ixy-��R�7(Ű��-���@��k�M�	P�&�G8��.��ҙj���Za�0�G^���su�ʺ��LV�n6^�v^��G[=\�tȯ
u[1����y��"���0�:&�#�P�//Z�%�0.�ݵWtr���kO��*ID����01{֓Ɛ��J��S�%v������g���h1䮃��G0!$�&0m8��`���|1�1���O��z���-S���:���H;6:Y�Z�����Յ=��9M_f��b!Ω�� 2�h'�/\ͽk9�P�S����r��	�A�S 2��<\�k��S���nL�y��z�}��a�l��*�|�5�.�[3�����!Zj%�2EUl�0R��6��Cg~�@��NO}��6+��%��N�����N�����i���!���y
"m�ґ���^+Ϲ�<9�W2�"V-�8�7\����O4��)� NS�NM�X���֟:�@#�-D;��$GSY�lv��6���ꊠ�p1J����Kqy���U�(.�R�k3$8�OC�`A�����T��ˍj��mf#x��v�ڂ�)=m<�h�1��Y�^�Y*g]�,�]R��ݼG?A�i�yv��6l�W?)���	��X����N�Pw_�4Ti4��ȕM�'��Mތ*?{&a��4�����Y�Ƙ�wC, T�N+��Qkbu�?QԶB�'[�.k��B���s�vo͖�n>}�Y,��mLG�����#���j�&x���tΟ�*����,/�͛A�'�	��9�eTί�s�OI��/"�/2D���i��/��;<�fL�y]T�v[~�% Y�F�p�$V�T����laΰ�.V��� Nd�
��o�$oG�n+@��0%�_pԕ(Q�SGa[�!���4�{����Q�Ue彦}( h_2Ch�n���v�T=P^z4��o�$g�PuQ:`=������_<�(m�x�xڱ�}O�,����.�o�#�Xd]��8���RVt8�V���ƃ�ʳ/<��N�.Tq\s�F���M�efZ+w��:\��ENm�R\��E����HP�I/_ ����<n��&�%ӢO2N����ZT��R�vK"se�*jm<66�F�<�@��}�[��k͐��o����{e�jg�1��9b��*��i�
������w��˸�М�������W}2%"��D�X��0=����~>�Q�7���ښ��I���/Z���M���℠�K|����J?�9Z���9A\��Z[B���l�pK5�U1��hi��W|ϒ	Bs��x��+����/�� c(��W�YʐA[:��u�A9ߨӇ*L"0�k6N�13�
�ܵ-[U�L�6!~h��@z@���ɺ�?�Y�"���P����O�&�L��_&�謲�M�9u�4?T�����F=�sP�颵*%�۰g�������"�Q0@Uu������l�R�Z��|�*�te����
N�$33<�IG��i��e���W��11W÷L�
N(�~#"X��#v��5=��_9]T.8���/r|b����r\�y�ݐB�	)�������Y32�X`6�� Ͳ݀�+��Hi��3�V�ە�n=��sBg���n ��u��{YCE��hh��{���m��\�����T���hfѫ���^
��CN
 �Fe�-����6��\�bPk�A��B�[��z`.���7Ye9�[�+��ѳ�w4fƲ���C�S-��5��{ill�SA>Nb���]�Δٞ�`��(ذ���*�����N[f۝�j��n߲#-U�+�I��zܠ"�W��rT/ I����'�� u��ִ@�2y\(����^��V쨓H'���/Ŧs�Dlz�P,F���%���\���2�4��m�a���P�%?�+��j����J��ռ�R���oΓ�3N���{�R=�~�`EG�Z$��G���%:$����r J��X�1����E ���?e�������P:���$ݺ�H?:� ͊#�ғ�ܻ�MNZ���k@�|���z�ى���'��~��tڅ@�B�,�8��f��q�<�̺��ϋ<�|�[�󢡙o�~Q$:R��{F��>#�s�#C�n�B���ΣɿJS����S80i��YJ��$-�f�E�+���|h�Q�()���U�	Vɪ�0^��U�,[��I i&��X���Nq��}�జ]��
���à��y( ��h�A��q�L�=5����t��*���m�7��ʹ�������i��s�$"e�|Y�:[����R�3�
�\����P��
K`������:έ��:��5׸��ͿAmaz�k��ӊ�f�F����#j�{�ѡJ�@˔��b��&(�4r]�e����d%h���]L�Ǹxj7��!� ����%��h�j����%�g�F�.�[��;�VBv�e���"��+~��-;��:��T�ϖc$�d���ѦJVL�'��T��Z�KΒ3�(`��2E���N�HS�_�� rV�ϥ6f�=�� W<b�f`�_�X�ɠ��h�E8�I�����5sk�a��[�t����1�3ջb8�L|� C}�l�}X��
d!��k��*�鳨�0}pdÞ�Ji"l�a]�O�:olI�ǔ�M,��#��PA��Œ�|E�<���삽uA��" ���{��|��ʹ�ʜ��m��)��#܂<ߧG�/
���i\��:�G��&B�`��2a	�1��2�-ڌ�&�OQ~�wψX�dG�u-�{��23%�5	�ZKP[,��}K���oX��r�W���d YYgR��|p���MSVU�-G?��p��ߝ�����rޗ�m�����bh����Kf +T�ϟ�B���~�z�qy%�}����ZP��@�(�N�C��y���cp��8c�?�l��W��m�)
��Q�d0J^Ҩ�2�A1>�Xjt)��?�N4 l%w����mn�`���ܕ��F�`P����:K�B��;��GP�`�ZF#��:)���ƅTW���M�)%�^0�2�ƀEI�����K�l���]*蘌�޼�ay���~1L�uE��,- ��e�|�ј�ߡ&O� Rsh��T��)����h6`�{����x5=S���p�na���� ��K��.��@l���r�$w��b��"����Z4Cװ�⏃^�����Fj�b�y�F�h��ϥB<Ƒ�Wya�����|O��G���1m:Ụk@���f	����|pc!��T%y�U,���~�E��$�k
=q��A���/�I�)R$q-z�_�:~����:�7�� ���V3��<}F��O�!�cq� "��O;NB���Kr�[���7[�x �03�U�9$i�)��'��c-��3��q[9 ����	�TY��H�~��w1.fߥC$��U��W%��Mi�Q���z^�TG�,Z	�;�
�~��M�}?��(�D%�|^.k�LX�����S�I�qb��T�I*G�����7�o|����|�%1-�;w�:u���߻��v�f���p�6zhv{15 0��=�#�k��Rv��y47<M��޽�;CśK[NF���� c��:nH.k"�Nԡ������6�x"О�e���u�7�BF�I����τ���ع����Ji���2��X����n��0�<�6��5���(��MM����)���@3�Ԡ�r"9��U�������	?�$o�Է�v$�B�J����z������W�M�����g�W�a��I}\M�	~O�����a6�� �܁����/���BHdO�n�5��I�a�Mb�V���Q�3'ʲO����(ar�\ I�g3�m�BJ��2i
s,���; S�����4�\j�)JF�����c�9���=��v��.��a�����R!�J��[\����n�!�����n̴@ �-�3б�ki���������)H�La�>�~�"wG�V��y�p$�H\i �E�#ؾ�楁�!���Y��T�E�j�`v�{(a�av���:�ꍙ�ۚІ�JL��|�8��m	H ̒�W<I����NL���9�V8��Ob��`����WDS�F9P���֯.�$����tU	����<�`t�dJ=&�z�7k�墐CJgh����Ey&!\��/�h�':4�����ִ�J���O��B�VQ��O��5�RGM]���,��ү�<r� 4)2:����ST��|h 55��| ���Aï�S֯$v>)=eŘ�֚�oЕ�*���b��o�PN�$擜\�C[EaGx�f5��g�PF�\/,��,x�Sg|~�dھI	���/~�W7uv�!�l<��{_y8c�@��ͮ����pZX*��ԕY��(�������U����]t�k�I.��[�M����0����H�s� ����� aR�n��9ly8��Ls����"0�����lF�I?�[��H�S����,A��j��� Y}@1��.�7�Z~�dWd'��|��[�c\o:An��M�
�v��n=Q7����j����Q�xZ����1����`~���j>D"f{��*��)�>��$�Q�_
{=�;�~!���Â���~��r�{j��Dܜ�롺�b�5���3k��/ lp�,�:�(`ǭ��S}��;	v\4�Fs3c*  �is�mH��Wy�@�W*OY����!��Y� ����IWS;�23��h&�=%���"���_b����_V�̀��g����LVv3:而��q�r�'��חv^���c��ЊkZ�q%�	2OWU�����&�]*���V��;����)m��t�x�:�&�㺙����C��su��J�鸮��U(C��[�5?x6M>n��Bβ�[L�
ZBLP�G�>o4� ]z�./� ��`��Y��4q��r�(չ4���3�XQ&������x�������n{J��� �MM�{gt���քoE�J���(K�,� Ű� ����y��@�����;�͌2�|�?����qܻ��A����s������	�g�;��[�2*�-:1�@|:����t�!�����6�th������0N^�+���S�:��ɜʴ���	�8��|�V�LGa/)S%㖶8JzF���	�l �gB��o��6}X���M.�쩬ԗ����,g��������,�+��@t��gW¾�
|1�����6�i5���N�yV��P,��6�Q��i�x+pz�L=u��
`���s'���<蜇�~q,5�%�FwG1�'Ն�y�3:
!2V,d�^�Z�&�f:�C�_X�Zu�{a����D�<i7_ ����F��0�,�R���>URL~�R����N:��J�ɠQD^�x
�J	a@Hf��ՠ� �ѿ} �aAk88}:U�\�!����ɳ��,1^�1��c�`�|�D0K{�C^a;o�iHe7�=���(�]+�7l��}�/�¹��Q4������&���"� (����Od9A]U@[�P�w
曫Ya��&�q�{��'Yds"g��jN�ϤE��.���أ�� �҅�&{U'rɗ�<^k�i}�,�+�F��F���z~KIvU@�y�r2&>�x���|�gʈ�R��)G�I��X����~i��<6�(�N�V���޷c�4h��XJk��C�� �G�\�:UZ�`�+�����B�-`������l�S�-��1�\��8��,�E�����(�{�F#���*8&�*�L�&�V)%�
!1&��E�̏��U&�P�����ݰ���}#�[!ͫ`��y�2�����M�u!�:[�1���:M։�4���@����%�шQ=�c�δ�큔��z;��R�9�����r!l���>N7���g���"y�sv'!\��[���s�:���pT=_U��z�;N��Z��aDD�{֯J���TF@�,��]%�^N�]������Z�Mf�X*����S/#���ia��b�߮�+|o��8w�z&��T��<�yv[��v�o"���m��URZ��&����j�x �7ss�l^�6~�jtH3���b�߅ߠ�Y�t�fJ�=�ʉ��EuG�u���R-n�)	�qԣ,���K���䈶"��`�	< o�C3ڹC�� U��Wb���5e.N������X��Z��O6`rFVF����7ً�� �!��cFG�)�S�ʬ#�a���V�&��X��.���鵁@M##�AL.�%t�`Z���x��猂��@mP��zH|^�u��P8���.!D�
a�V8 E�>hlY���R�;,��H;&+R(ҏ!�)nۑ][�c�!���5v�����sf���1,�gI0?��8�J���&9��B�o���x�7�����C Xd������v�����B�%Z?�����Y�Z t����M;)g��G�!�0���JsJͨڎ����(�rT�Gʒ���B� ��P߰�r� ���6V���T>���k��#HL�Ѿ�j���8���,K'�,����~�5X/|-]��b1!J���W�+��d���G��s,��i��\�A83#��~El`�A>���sB��1ā>)���x *�DƑ�����7��\�z���}Aω`0kpw0:L	�4Ѐ�e"���)܂6�3�4ٞ�ߒ�`�K#��,�ρ��Zg�l��I����6d$X?����ā���+��T�
���9nc�Ii.v��Z�uC�&V�g��f������
����ްg3D/���q�l	V�v�?�ި4&�����!�-�Vǅy�K��張�H/�oշȦ��kU_�
�Q��׳��D�Zi,���}6� ���Y�р#H):�KA����]��Zw{V���? �+9U�k�:���'R��� ��W���!�p78_eE�0ז�U�'H*���9�Q.��R ��]j�_�@	��K�k��o�ƞ��k�q�VBL�xU����n�)_�V��H��%���oN*��K���:Z��nH����%��QW��dC0Jj��8þ7&.�F_�h�'�F���Qѩ<�� D�U�~�D����
(�0\�g@���9��D.U9��7U{���p���],}e;xCo���-��4�NtF؅���)����t���ܓ��Y s��G|w�]���q�0n	N���S߮�^
9�>�8����� �x����Jlh��\�T��Fރ �s7P�6��M�w@� v�F��������?SgҴ��1̶u�SK�O7�j���I�(|������[���~��P�͵��9=�U3��Ć�Z;b������ŵM�6�8�⫥����i��X���[��e�E�j�Ww49��� �y<�YEt�����j:�J��YשT��GgIC]kN��"����b ���~�(Q�[��g��\�,�{b(v��k
��
����W��'nTnN0p�y�駇���O��S.r{�w9�K����ɶp�f��%����4���VFWk�A]S��|Sp.��u��w0/����8��V�%���ʱ�tb����`\V�zSfG�x���9���v�d;�9�+�����dS���D:���[}��(����%�ck��g���҃D�Y����N��N��a������uvmD�ɕ�}�8b�#��R� ߛD�!�<r޲Un�92�%��\Z0��!l�\�<^�C�I��|㮧/�|���(�8�9ťD�jb��]����U|��w0e��l�(�>c�V�7�)�d��va7�������u�
��Sb1<c��	�t���ۧ8�aA�5e����etD��+��@��{��)�;�z��-&�v��LV��DZ4AW>ys��/Ux������|���:؀�{Lq�#+;�YSA�Y����9)9Dc7އ�4���qrOnZ���ٛMc%Xeb�D�G������5��)�����B}9���֗�S�����Xh�Au�P����%ֶXP�#�?�S�sGdu�$q?}M\]��0&݀s�2p{̇R؄z����Hi e��͒����+�3��W�z�շX����3���[۟���Ŗ�V{\m�o>W�Ƚ�p�R<�cOϻ���#���� �j��H25��ҥ��pU�2՗ݷ�G>8 �0�Wb�����3F�`���9`�T�������,Zw�&� i�kL�A���m��!�(ж_A���쎏�eO�����_%d���T���-�>3Q��Yb�����^���pDs�R���Ƚ��)����l��dk� ��O�G��9�')���y����������g����"|	
r��.�~s������WKp����&���
�m[ �8��.�V��io�Ҕ�^�!亭=?<J����%�A��p�9��L�/��bn�.�=\i>�Y�^a��?�aД<E�A���x�9u�7E�����=T\T�=݌ |C
1�
՜���]ٳ�z���˄�����!�#��/�6�3����-O�:�n�/���[f�(��Pi�Cm�9����v��}�e�1���5����o}��>q��B%q����q���
s�UA]���n�XV�T�i��}�۽��{h�$j|��`ʒ����by�/!��Z>��*�º ��Gc��A���UL5�Y���]��VJ���͌�+G�n�"rкMfd����%9C2��YY�5WW*�gu��^K��K(�ǒZ�<��2�L:���\�VTܸ�c��#x>��acXm���^��	bex	���N�穠#�b>Id��P���UNЎ���p^#�h��:��z&aֶ������m5z��
�p;�=��j�&��;��]T�Q�R֋j�����gC�dA�!8I����m l��G��i˙q!D:��j^M��!��6X�ʰ��T�O?|�����b(&2���ʻ8�b>@X��2�:U�� �x[R}�ʉ��/	���(�ka���$4�i�+W�}Q.���m����k75�9{-����EWѫ"��&{�����|�=���"{�����DET!a��\ơ ����e�|!�=}2\&��F;;�g�t����op��;���-�K�B��裰Ų�<�mg���w��|� Xd����}�����u�޳�_��n�%-���̇��C�=AΙ��^����� 5o���C�Ҏ��E�����A�k��κXn$��k<B<w;~�x�Y�B�����>Q[bn�<S|��`�3�д���i}�CL��t��Sq��3VΜe/]Ѱ��O[��|wƸ	<�\��+&�T ���ػ�Y�1��� g��E��j�.�ȥ������2�����yb�`el��t �X�"�,�ve�'�߆� �ұZ6���`eCG'ꃉ\��#�� �[�Zm��j���g*��S�G�'��b4��%���#9wгF�������n������F�4~�2�#��%��(�z�>����,|�*+���yڹ��=�%:Y�u��sAG�#I�Y���_�:�I6畽�R��j�>��س�-l�+M;\YLm�� �C�R�=m��Dק~P����CL9?t�'����Ý���5�2�儇�d�����_sc��B�?�Vn7]�5"�����&<qS|���G��B�aquCYkG��(��X�-Fƥ�����u��5�菠 �c��ō���)�[����x�S ������߬����H+���\y��5)��ō�[���nC��1�N���e�;�fE�r����_pa��1�!�z����F�S��O�n��Q�9=x)����n�Kp\7T��\�R���Z���)N1Igv�l`e�ܮRX8�2l� �����<�,
��2��I�<B_C�Na�<�9���4\�;o����buWY=��tM�>�1�;љ��;x�� U[��R�ҍ�9M�У�׫��:]���4��-2��� �����k���h����藪^�H����KH�]	CeO�!�`�� ���T�xd;y�K$��U��M�/D�P`���
#��l�m#�����VfSZ�/�R���'��,���� ��Iߥ������)D��\>�
-O,�e�ST�M]��q�%u�pf�ܹ]�%dX:��ҟ�|U�l�݀U\��oM�~|�]�Z5B�Ǳ%e�:yZ�:�I�k�S���])Z�L����Ȫ��^�.J!b���m�+3ĩ�x8Z��n� W���r���J#���	����N��#�1�͙"��2�MzFG#`�rz|�1V�K��c��#[�����:�DYZ�#P�Ĕ"dD^I	�O���J��C�L��(�}��Rq
�Jp��V���x�綗�X�,u�!`��?���z^1 u�ȩ%�vyj�������-*6��O\V0�I�[��� ��:G`7��d�����~�Yx>͖w�<V֗y��6����M>�&Z%��eM�K1[C�H�h(H'L�un�Far�������,�f%m션���8'�e@����2�a
� ;�!{��U��_�Vt�n6X�����b�t����TP���v�-�lċ��A��ArA~J�iv.g�h�p~0�����?>�
����9���s�?]r\���{�,���0�5���+�<�-si�\���S�a��S��s1ASf��?��D�I�qVh�X���\����'�ȳb��U���oiT\��=Tg�%�Aa/=�[�/"&qPH�-�����g�*��p���im��9���kO����#����7 �r�1c��5�dȮ2h�ǋ�ۆ��/v��p��^����\�/�׬2�Xɑ7TI�x���#Z�r��aC�Z5��kW��Xؠ�2�����h�Z ���B�
_~��5{���y��^��eׇ�_���0;|P���ݗ+,	w�(Ὼ�$窼�G�oܝ����������r�!�)d�����K�.�hP�^J���>~�ܤ7 �nT��7X��1�i��F��J��0B�G�2Fd�_`"㤌�CJ��~��<Ly���aI�I�?��)�K�ꚪ�[���t��a6���0rh-���<t�u�� _�V��  �x[e�]n�	d!�F���V���d�H�g&�I/Ԟ(<��.�z��>]�?t�'�?=���a�&��<������F�#�≱�\��FV�tD/��*��3#��C��N���d�1iBf<wq ^�[�\�t��I��Q��r�71�T%M-/	U�e��[Z䆶�w.����A���9t��+�U�ؗ�y������9%�4����j> q���k�iA���2����` ����X�g9n��9�;�u�mt��s���B�D7��M�����V�̛�Ά|�	Yo��<p�_��n#�֨/ 7X�t�j�^X��e�j��R�i�;`�1�V׽z>�	�)�H{U���!L��_~���ڄd���u��8<�M��	�:LFy�� O����d��t1NZED�)Bv�#�蓤�DGH�-@�H�@�T�l(EG�Z�4s6ջɏ�|��B����@Zs���7�n��S�=�ݘ��S��iN꿏����b����	-x����n�ɩc�~S���[dYO��v��L����rX�x[Ӊ�����D���ps���YR�8\Xz?�~�p�S6N$"�@�2�N�Z�?��%4�'t"�f#>ͱB�萟%l�"�w���O�I[	���}�*k�kD0ʗ����D�7��*��N�	�e�|v�]�P�~�]�B!|v��aI�/�
�T��������I�h���7�.���e/ÿl6IV��}{ލ^��U�KUY�y''������wd�2��
м�/$��pײ�>*��3�^7���ؚG�$Ryri��2q��=�R��X��U��t���3���d��OAw��򧰥�c���?�H0�!��tr9nh۲+� k��҂JG5-M|e���z9N��t��.mL�?�l���T����Q�l�;��>��q
�.i�#��kl��[Qey㦴���M���{bD��l`���&iĲ'�7����_�����]�KK+��sP�f��@������{��ӕP�iV�(�|��@eј��Ff���3��nĚ�a~�kJs���4��B^z�صA�5���|���\�LR���6���ǪѠ�(Ͻ�ؿF6f�NR��\�~����|M�g�i�u��r\�z;�5&�����²��|O�-�nU`$P�����=w0戠y*>Yӝ���!��n5�H���Y������r��h�:?iY���5���
Z6�y8ŒQ꧸Q1.銲�vgM�-�#��]�E���6n`N�՛>�UHb�*�?�LP����u�P`I���XM k��Dd�J��\���ڔ�j�+��n``�J�V,��G�Yb�F/"�Q@P�4� ��6�k�?Ȫ���4�]e6+�J6�'-(�'Հ
��/�"����Z���v0�er��������k����Hj�,���m@ ;]O%���1�~�󮵐��Z�M�(�gG'�E�-�,�p}c����T�^.�`�|lŔ��<�e�79p���Ī�|�9�ں/��)��}���{B� ��ˬ������}�aa
%��\�l{Ԭ��y�G���_
(`��5����:��zf��^��P�EzPZ�;�?�F�غ(_��vQ����7�[�*򕊲�q���B��e_"k�.h�P�)���Y�_L&�V��}�e��+G3�b���/�P��A���F����G�>�P�8�u��V�����4q����ھQ��wLj�-��&A�Ks���V.��v���^�U��V2�ex!Y�U*/vXoE1-����Ó������&G�Ri4;���D�*G��>^o&��n��ו�h<�]Ν�5ˎ���rr���&��{�ck~4E��,�9�j�r`�8�v�c��H��
�D�%l��'r�T}xA������Ѫ4���*�o:������F��)`"Z|4�#sWAm�#��5*{N�>�۬�LB@����L��$i��u����a�K1��8S@��,YDV7�5_�����|�#��u续w����.z��d�E�ae�=+FЎ�GX�>�uE�8�P0|cEQ�ذ4]B/el�ޤ����9�����6�q3�6�Jm�,��)�`2m�'�n�lK��&����u���{J)��x��X�Ke�j�ޢ�v�1USK	�'�I��ޘ뎩�Zs$��.r�-�+���P�����k�;��go��#�ܪr��cD��4�OQ�}mX�0���PגKߠ	@a��se^BL�]�-�Cl�]Y���\$}N��N���ٌ)@�[ϖG�_�{<�o����*�삇�vX�h�?]�;��~����\�68�a�����?�s��r8��;}�  �dR'kߤA/J��a�	���F�)�������.�񩓔Gb�5����ؘ4,�v���l�$����5~��|��ۤR[��6ɰ�j��|��s>D��Ȋ�3:���}ͣ�N�Pv�֗��5���أn�����oY������2d�T�)h7��o�#2�&����6o^�=��1W����dD/�� �4���	�rݦ�SN�mBS��<��
}[Cj���m��X�8�����.0fd�����/7�Q4?�Lȡ^�l�-����3��vjOE`��]����|��$�%3�����7���(��� ��b\�G[�l�b}�T��Bd�����	�,�&�����65�����D�&͌-l�9_ ,�A��6eP�5f���I\�M��d���PaoH|e�I,�L���&����_�yg��<���67����T�$F�M/�@��A��3zͲ��N����ޜ���ixE�*�$�1�%<qzy�8a��da��)�4��R!A�������t��v��k9�c#r�T��3�2.���ZS8V+Pdm`���Zf�_N�ϗǆIu*Ắ��ߠ�"�H�(0��rذRiO_�z���w1\��}�T�β��t��ʵ���jn,J*��E��,�5��u�ԁ�7����涆>�߁'g�j���GZ3J�ĳl��a�Q��X޻����A����m	�q�S�Xu�ޒgj,��A%r�"V+*D�7+��p�>*5��a�y*s���$��N޵Zw��;[��8��.���qٻf��\��o���G.�|:��V�O�k�@���Y����ێt�V� ߲�7�L��/~7�R2,��y1��;����F�XTS|X�{�P*=
yi�(���yWn���M��9�Z/F�jXeȡw]�^N�=��Y�.�Q����;���c���CG���|}����E)��3���