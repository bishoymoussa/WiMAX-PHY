-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
ZhZEhocKr0rhGoNQPaLaD7rXEaJ0f4QN4+75vSXfLi24xbG8T5dPpuVZYm4zlGeBW+YLVMNa6yNp
Rj8OcfkgV6WFMvMWpjq0zq5N8PfICEGCZ7Tk4KoakfPXDKN4ctr4svwiyqWqUSeYu3TdG9UmvcS2
tqtB0aKbqZQKBCGNenMwGyLDUtAUecan5ZbRg6EO5oOHfXRf0xpLby0FNVm04BjmIT7GUcrl+Am/
P412H6qwnRaVhZpJXat5YCvz0LkSBQsrGKkJ7WxiFAjngNEhrqrYJrkScLhXPA2oMZ50RRC7vMOh
pgy4+EPyXOByxtXyF2TBjknNyghfxZ8xFdMi0A==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 119056)
`protect data_block
Ud3uLlCZgsRx/8Lqn7L2TvW9hwsNXJ+Gky1PUL5W+OU/sIm+M1Y/OJK9xKRgarMdYZUt6Jxyda6G
Y2P5oGBsOz5GTnl9bWDmIvcAdGL5yJmzIPOthfkmm2FFZglQOI3vBepLDfYzY0SofTEp2azepLXb
AouwKTO3NZXnoocPhPIjUOTbdTZVZOfe6+TqhUtzhDI7/IWbcll9aG7KHT2s2OLkm08RPgiXyExM
szv750Bj5LiD2mbuaNWHUNUAozc5Fg+mi5bj25+NCbUSTB0k5gaQq1DkZu80RU9bJELgwzb9F3cD
mNA7P1+a1Tl6gZ2bajJxvb+5OCnjObiL8A6kFY24Wt1koZ4Fltk0EnU/CQzG6lWJoDal7FOn39Ky
dqHE+Epli61qf7oG/6odue96WZThtR1BZXOS4uDvrZigRTBDdyaKdfgcc21t7Rlc5DW0IihKwwgu
VXrqASnMqXRpTabKTLWXJEYKVndeVrXUnYY9fD1EZwwQkdAzyaFtSs1IJ2yMb8ylpXt7bmhKiDNW
g0vutxbYWyIfPsw7uIWQppYR0wvRqXrBUL1AJShJR7pNaeE//+209V5FJns5WdoZCbV2OKonKJVw
mvVYB/p6B3Jm34VnS9sj8OVwmXcsMqt1y3w+x16ZY5TuIxP+0EXEpLfj/yLG5lkvI6BdfoaVxYci
PFXwd+t68Lc93rkmyYRBTcqENMuWw1jwUtfTOiCtHe0Pd3Vjpr0jIYb0LM3SQnnxJvbfNtLTqKdl
+pJnfarha9GNcIHLd6pk1CJ34t2QfsnuJsyhTvb6JQunUQ04zDf4bROQEKUMjkBbg3lsHKSOFeDp
UMaZ0AeixoL4quTyQ72OJnnuIsXQWsOQsmFFfm1Ylxu8J+9rKGRM2fcoiEmt7ejjdvuGCzj0u2Gy
lcceLJAwbtg/XJWqS/kVllJ+raW0w/vv170PCDkJpeTM0+nYPmun0UBA1X5ClevcpL5CTgUewUXP
6KJlPvB3GwQJ0QWnWRw7Awpwq4wUbmq//HBwCoTvVAzdrzO+byS6IF9qNFejdsRjVQWhbzbRbaCw
14MnICEUyZbFGLTFs4g7q16dOD03m4rG1ln01r3FaLlct8ol8lXyKUGhGuiCVZVCkP93/K5gd3KD
qMpiHvnxIkcSWRLONZSKpI6L8/mUCdykNLtgJc9UK3ADDDyD2o1yViqiVf5fn3HY1AeIjKtnyXW9
WHx2+aGrP44vz+pl/4WJwwAuaxegza+QYNAvE2w09q1nk1jAW5PVrtW7MFu/9IKrXj2ZvImexGo/
IUGZHug3NTU+fytOb13EN2pYsUA0C19Mj2OmoK4o021tBz8dUnb7PHgIO/FqaEQGMCequCY/R2Kx
MlDI0ajarkIzibiKIc1uPPJUcZYLNz2sIAMivr6MdxrhuyO6xDbgO8v3Mz3qOXSyQH1oba3/K6Ss
CbjAAJizaaGOC5CIUZVzdk1/cyQCdoBTal6+7qJM6GbkGIHx9aPjfBIHLOIqCam/ZQmnHxiqfA72
Wy3wKsAp4upZF3PoE7bxv50dj8LfEo/Hi2aFUyNV3HBbKFMiki5RIBERtDTCf6Thw4OifGSwKplM
ViFh0hDd6az8DbMNJuCJwRCRQQtXUlgR7Ya4OKnrCRoX932uxUWLBIjwIJZVShKxk1+aFlJm2/Fw
WDLJ7MraGX+sgFNBwxBvlBo+oTu5NbxObYBO5AByPfnFrj7ZpgijVZ3Ou/bO0mcSJttCSZkMkvZG
hO0WePbqGgf2ysBqiWga2H4s63uayFbsrzcFqD1LExujnezKRZF9Hnmfg/ANHO4qsNsNPGhlX+Hn
VOVs68/W1GoGIYc2c4ZppSWg17N6h1W7r/CgnMTDBWkypm4m9uxhAMfWFQD+SszOhO5tJTUs1tPT
YOHk6kHCaFX3vgCOydd0khwWJyKgHyTI7zRR5h1WU2bS12UJQIgIygwLpJvGT3HhKFle0gPZrBG4
1yB1TFE5uPTofJLjnwQaCIjZTJ37kjE5A8XW6ovhBEoBHL+I27LzOY92sAWKeqs9y8fZsJ0wjaRt
szqwX8JhlXVcVr+KssSi2B7Lc3rjyqjO8qcy/gjG/H9ITdwLSxHxAcrPl0wEG7IRFOsM733sVn7t
PU9lo2uglBuqEHCh9rlw8R+QznGMBwd5reAX3E5cFr3WGzmlC7e7pAs9nMz0xGEo3JLe1rGVUMva
VeX2eFBPk7qGu8X07c43j+8Ehm3b3j+1GjEMJrwJupnUE0kSWq2Cu6W7PUW2zPLlUvCh3Wm9Q2tw
wqtMYtJA3hAgeQLaqUK2Vi5ZMlAs0LmP/Gt/t614uJeaNAMnvf9uFanfxFPU4AZ6ThvRhH46mOwt
PHrsGyer1b/iNuytORYVI5HG0Dt5uRytVQWngjNQV1eFklpjVlmUjy86Z5CCH7YGsGskNxdfGZDG
FIOkeJTFNVyMn3ymVhXiq1p09l81tagsFv7+PfvO9cs289ywKlEkClF3Yhe5qU6VR30oJuwVpSnz
hQRBkrU7lvKTNfz5ncc6UPzjw68tTqamQTr0XtogwaumWyrGhZ1+PG+hl6W8HGzCNBxt5OlJQ0xw
e9BNHZtNPph0+GxZPVnRDdJ6SwT5TP9tO45NEvBWW9R/KLA/0/CT/alATYZJWYdfhyXuC96VB3WL
WF8jx4RRFnpYO9bgfNsA4Yew5efH8DodGOMzvmwfuzpXqyT83LPrbKQH0H0ZhDJMmaiKcRyoM2FY
2FFVy/uqXWrm8eMPPZc7hV3wJGgBee/gc5DNqxhxKZQFUusRdcPi0jMCh9nRj6Fb7amGC5lWd1Fh
w7F7VM3IPcQM4wymAkIm/EX7xdXlMtLlXKzYXqPdk/VC7bj8aIDJwI6xjsoJSGf5PS7vX0iiuERS
DovWWgD+qe3oaVRb/3kC8JI/h+BvFQVMDpCFG6w7tHfvc9MryCUqfyj+tcJIYVzndFIjlNIYZAbh
yC28+A4Y/d+2vlQlzY+gTxQ7ObZMzx6b1pSjXxJzT+ssLb8EK7G1+bMrlhjkv3z3zak5cgy3lOeZ
wV9yoJi6SyCir8C3KAI0u8kQGh2IkLKF/xRuiHVFkNXar1WWOtIUzX1kjg+dQcAl8v06Tq+ZmEY5
1FgrndJO4jCvjKYKrk+QPPMROB4Rw7xsWaboZM4o/xSuVdimARNAGMJjpcMxJJx8sj2H+o6n6K5M
WttgZJOV0/mZ/Qv93ce178K2PfWbK3mqbQHC+nOz0PEqaiekHJxRrlMHg+Gq85XSgaJAZlvma/cB
NMqx90GjQH+eKyE2gl6Ha/v2HkdS4HCjqM7iykkmg1ms8Ol9en7uwiCOUZHlgWEzE73ViTAKcNqN
1DfNNBbcP3V89MDV43iWTQOXbCQdFEzHnnAS+eANSXbjypLN/Tdu74CVeOxEvoJgEpISIpd4rHx9
E0yT356NoSLRpSCstn/OU+g17gu3ic0E/HYZyJuihKLxN0PHS9JHTB0yuOExXM3oPra01fL1zvNO
xlscw/M6VEneRgGMOOpjs9tedSM/E3YnVCc28BInBPgWSbVtppNTYWcim5gp3Ty/vvM3gYF92ofN
I36iCuM985S2y7PW+iv701ZcBNXR7WIo/Xt0uVVArKagcIDASeAV6ntGK5XpYVBdIMlGF0YsVMPF
xHOLxRZlQuShM7OViLDTXMh72YyO5SWvaxouEomsnnoEtM3vygYTcwrJyIBliyGWF6ImVzQwnyMX
buXVBVifttp5s4tahDVya0dIAr2BbY9UpYV7+nlC5MnnazH9iqOgsmsuOiVrnNC7+o5ZP4wUdvBz
PmBYM4KVsLiMr2t4LuobujnCmzh0fK6oOMEVnHEIoUC6OfygjBLFHNhhqnkfAig6IbpKb6WRGzjy
fcuioToWA7acoYsU6KUTZtI2SuDOmsMuXv0b3ZUvrwfMqAIS5FvsUnhV+MjGVml3UHNAuvKte14c
9nD0FDupG0XdAKRW63qGhOxKKUOqV84u/HVvil1OEXhwwyX3g0bhg5eRw6iWZB6K9zWImv9z2l4t
ZJ6iKs1xJRJuEwx3tVG2Sgtu/Pv4Z8h/A1o5FBdpwTQXD584Tot7NLVifdIMucSKz1DEuiGhj/s6
ujif5wzoK1MlLJSdSUuCZ5cRHUPKjYiU1CESXaAH1/v9NF0oj4cos3m40/Va9STJm+KuaTgOunf3
9Fcn56AkeqJ9E7i/Tv7DheHBCULAjSXcRGrNTp+4a/gYbBhB7HqqXQAZFn/jVJZ0ueYdhFAGSbUi
DAHnqZj2LacRXCrjzoMnXBaejZ0vVFxc3cYiOiNq5zagmyFBZQEvakJs45m4AjPi7JxhMbRIOfXH
1CxBtzy7JUa63npBqsdOWrpHUMfSlTuOKGQ9gPXQq+HohCN6JzQ+dp3ahhGwxRHdTpUvGz4rzj7g
sShd+0GE0ULyGFvAZDfXm+UbnpFn3g3VMyhc/x4tPWZuqbXX+e/PYbZ/cGw/5+ujx2G1navxDaYq
jGySK0e/fq0m2JC6jGtpWnmU8QHlHHqZgi7Vzt+CCyGYcGSkEYtinSFlJ2MxAh7X9i0OH3iKTSBR
oV7p09S1/RqSmP6eBjn9HmZ+DbwQup+oh9pgVNAPnQvlnQUVQKq5CK5KH44KYNhT0m4Q61MZ3Pd5
8Veoc1tyL4qmzAeTXf1b6B1dGoRmKWwBV+TGLUMucWtX90vvZTadvDJdAYaZGL1EtIEOsscMcCG2
8u8gg0shCwa9689iT+Y5zrY/6PxvMG9dQrYea5AXCgkzvc2JLpb7LnEvZe4/z2TiveIlzMYsHhOq
/Nog56oX3HpJF6opy8jYM7Rni/AHSlL/yyTRtdPMhNXt84hciZu2ShVcj66Jly7yLgl4A8wZNu6h
c4AUzSK3FA1juGcKWVXmHwEij54eOtRcdgbYXCaprfw03DCYeqt5uKhocgZbKLtGp9oQu7VGXNKo
bYPZtAvVcT4oBInFYjfeQ5djPqnCO3kRCTyN0T4tv9usAVN8MXbFAQ+qHlg8S36b7GD2Ir5M1dm8
/IVF/9sLOdwO19K54PrFReVVsK/jigtCwISVEQimU9N4650IYUSaRI2tBPihxmgxdH4btv4BvBWL
DXt2GFWW8Z1cymEVb9VR4lQvZw6fjY1vltEwMujWsQCrtQzIkGtlPCWxH/5EjjhoAlBvRyvzwPSJ
sQGAdw26VBjTkogj6VqUrEiyCMCiK1mlDjTsB+kqUQg8a4qntOffIQktTGRVZ+waxVBPtsmeogY2
Et6lSoEYA/SWo4S9slzx/moxMeNdRFEMtpu6ZbXpRQWEcCfqORXx73OtICvjkObOuCZo40iLRBgv
PKNh0eUCd7EGLUQxO45YXCSEmre77402S+dtEcIOYnL3iUgJy8KchPs2sv9M4O1nPE8kPLsBh8ry
0q3cZQ0ucrnm3NFLmYDNrSaBp+ZKZXDVa0Ex9WBlWWPcQhgvgAl6Pxxe2R8Nln4tg1FxchLxQM6y
MgCWtXjQDfXySyTgSw32hz+00g7J4eSeYI4VFwj7uIT5plexKxKUfptocPJzVyOIgppRbttksUNG
x881uDvu0tTT/2oxHexyAPLc9d3BrHuRcByaG3cEMZ5GnpR/lmsAi6j1DM4yOek55q6zAY7Rx5pR
lQzqO1MoyWuW3Uuz8VRl3x55bR/pWR9vFTsjkNnQM7q7KLDPF9Grejmvf3pW7r4x4+e1ORDTXsb0
MIk69LYrV36kY05hvhnxjvyDG/gpvjRvZiRLKQUQ8cq0Yz5fQIYM3DDino4d8Ndex81EGHZ5Rdga
WmGf4ejfnzi8TwWGl3Jt23+DKg/fGcT44mmHigjZMphR6nWMgJinHMJF5SaPBAgroGe0bBn4ODiu
uw3BNXbnFoGan4eN1tFYCyx9RPJ76nkjjBk4SVe6v8IuLtesrCyfiYdUI95glUfnCBQERBzrrWbm
lzLrijQz/6cCt4VCbpJ2YgJxO5s+lql9BrNbtw5dlA8wlG3JkkGCWyr0v3lNZemQcKQpWMFkMNd0
TWDUbT06t5oq6bzKBXPsYQX/irDkin4B06yUUYPERZUio/fmuDddg01yY6olenBflE2Kn5ChSgNl
OESHh4is/zpevP0MVcIaN45SHvKZ3aZccHxH0ERs2OHutNs3VkOINVNBYvvHtYWMkth1z9llBnIb
muYqCM0H2p9GcIS5se1NDcqZ/BiGT2maar9TKFfcX7DA28ROwl5tQCps5oDFE5FK/eX6XXCGHdoR
xrowdkwoxSKjkZC8ul7w/3sZprmFQyOjmIvlO5qcTb+dsKOcAOroCx/PrRh7JHtn6IWk/UqDlwTY
IPM+HMe1numDmXO/wDXI4zeLk2fyde2yc8OqHeVBTcFOelkGjNuVUPTwWTk1PwHx19CzwFVdO0qr
XVWr4Xv24Z1fAqTwHxCGiiNDjZg903pUBOsNp2kl9JdUZLlVcuKPJXWbsGxceD8lvQFZNngF6Tic
6i5eGBBenNbtmKpi0QDXYTPjN6SBFvs2VlgyGzHS8ajLwoIUaYZ9JB2N40392cu6YN9xRx/17Ksw
SM3lf7nTe2MBmOikRQ3DjRdA8PssjJskeqeJ0lk2le4x2C51l+FhpHX/iJr1Lsv9llzwERqJVn8y
VeOUXs5Hd/txLspzscZaMD5xtN2gaoux94Kdgg1PeMhYXso+H7+C4IFSdH4rRZ8phFukxiDMRcma
KKLAoiXYnSG5/vwanAXtCmW8Aw0pizUl0KdA4XS31yN7vXwK0rLsslVoSUycEZbtQYeJj1JXAx6f
jo0NdDI0ixgCJZgqubmc2S9/xu6002b9C54vRXf6cj1m6T/FM9tEeW+ts7AxR3YgC5YZwdddViaq
+DmEWXUFVYBKUP9iU3t4vpcoY0ggfRhwFMf1dyKtzxDE9Y6zcNy2/R/or9963ho8ZgPnSaS0TO3A
g2BuMKKK1YvcMT8cTb9YRNx0iLfzf0ZwSnHAN6lV/YaeDWgUhTN6YceMCvf/DnODoBM2I0Sem73h
6mFDX0oTkX+0y4YFGWClqaQppupI1ZXPhPLcccZDF0N9cRNESChH35astqzbunKHreeV6O7Oww9C
vRYjgSGfg8nBUriLP4o6sQBw3634f6bzAMriGxFIwKSjRWknH+jpHkUp3gMSrBvnIt4LG6wqlKKu
gMPD1yQcxVHnW+PwmKlSGDQ37LwU9qmP7s26OKT7XhB88y6StCCWGen5B+WH3yNK74RBkMk1AcZs
UOqQNjQ0JYf5f8Dhm30C+9Sc6X55RKsQyKrrQgNioTdk4oS1zaFVPWeq0Ty9MVKCiwDxL3QGLIup
vPBqcAphwdLpclsd+SYJVmQh51SXJWUL9nz4ZxOGyo9KaTvnlu7XGsLlTyM33eMWeC+Aasttbx0O
xSsXwNYqKSI3jE/VXFTI5eWluW4CYB3DAk7nqv/bzSam4/H28usyuyJk5MReInv4xdPcrrEd8lmQ
9Zlh1myLN7Qv4LGfstkq4o05vZOCebnmeWjkydhdNS+cEI67L0qM/XvYOCA+dbUU46zye6wZFXvW
E8hS6i2dABUkefdVGeC1vKEkv5Ibq2KYXtdO55VFpTL5ysCiqMPvFW2QnS2EQU0+4bC7+9EsWqKe
snhD4YlgWTqPcg3lQcdE5VlVpW9Hje/+fKKXH49dkbqIl3LggqhKvSANfXNP4zFbSsnRhpVJzBwu
SqGhJuCI8K0dwqehXTB4dcK3iqk1DU1oMher1d+ea/HDbY4iNrQAtWskRETR906eJwXFiIo0ll6x
qURozl3pATJQNr9CsDpMfqiQt/YEYh94hLN77An6FTl0WXZWxgKxWMk9xz5AA8qlAWO9P1ppDF3E
aIpV/a+13TSPIWIfScK9HUaQ4mw/Wu8yEdpcRVFc8kVSQQv0Nck1x25kmisSmS5O7lRSmTUTcIph
HbiPftEqGzgrVWU08YQMEd5b/QJQ0Ohghrr7VS3Cn+A6rBLfOsNlFbVAFVIwxQZXJXsug/D60ABA
9+0R5HJEk8T+yY+iFIeuBmCliDPC3Jkqd8vcXrujqXZeY3eJhuNhTTpCvwHJ1T2Kf6epT/O9jE0U
rXF3xAfkiuNCE46YDU9HX7sNMs7nCMjrRqgNTZkiv//f8bERPNjC12gQ4Q9uY8A/HCtnzptFkVlW
3QNgsjAq1YXnImgqS1kuQNkCsxXoNBHJm/U/9AYVrDnP6tuvpUUdmyKViLscpqsoulMEYF/iIm1V
CYG06rUKnM9lxGkX3au2q2crOzRQe9D+xEoDlUPAg4V+hg5TC4UIswX73talA1bFZNohZMP06vjL
XTyO6SCFSdF1MsgQXEenafJwqH/qpvA8qzu+FyKDONeDxbLFro2VdoFQuq/MgH4Ic0nx3gD3M6f2
+AJqfopoTRzv1aVVdVtXcwvLY7Q1B3KqXFfop6rMQOe1Dc1n8qQc70j/k8JVbSFUaRgIt/Y315B0
rFM3nqMpgiEx7ixvHqhwCi6GfKcJArx7G8HQ3Q2rIQr6SMLyHm5/e1WyIfNKMwlTS8L3M/WwWEMY
rOViL/nPTR2HrO/8KnDGJxEOfh1yUIjxY+o3sN6mDNuw0vPaKsmTH9eVKH+IWmFLjK27gHRI90pX
y5WQ24KDU8GXxECu/oElyp83tpt5W/J4Ptdth7PrcXnMS4U4niwVQJ1L87zDN2hnKrCWZpiMyuOS
EiFZhewxkYP/+4zT9ftsYa9cSOwVIjE3nzT695UC+61Lv/t6dHVwbGDvC+A0Q45VXPfGx+pHjJ7e
tazZiTYBJ1VGJvhQk2XD6TIz+xztsRGxb7qPVoraCehPHkq1N6mbRGgKlcXbiBHuAtqEMBbTZJsE
efqguDIBa40SGutTnTU08kghnu6ToXBn2QJr2ydyVas5Pg666pKlAde4NWizhkWIsDlfMmx+q6k5
ebR7ni/aFdl7Y78kY7wc6de0OnutWmL7MRi5TOhveouD0+Y30xAl4pceORogaHKPDiGO1nlaVmXO
+L/ILkmtTqIm07emH6z2sbbxyKfy+Tme7iNjt1m6kptXk9SYAruL74cE2rAISq5VVqOyEZ32uBMT
mI6OGIovwBcICee/tPEduUvK0TngzYFftNs80zZCBHnAmjRWmoZgr5Z6F9p/SSHkDveAol3PHeqy
aneyoM4qFInqa69UMeaozLejmc634h3GcnIJtNm3qz9RUAB3zqiJpGQ7ubz3lQzoix11iSiOFDT3
c00Ey2xiflO1//p0iFB1ENu0IiagaQS6b/8qP4MCM9k6NZDDlmTx5G3NRNm7EvlqwcypCT/8yy1U
5ZlwWmCFE8S+nGdvL9Tx/mmHFGPgo6aO2vdhowicho46Le4lncQixRYGRqJavzsBpowFFQvHS1VX
CGoiAgRwxO+pR5edeB30Iz+PRKqlBNTFCc9TCn/6qpYrBQY0LaloBMz+zRU08CSk5Y77MRagyOKF
Vi9MZxvwNojGeBQJibhbjgMtkXZDjapWASIZetoj7b+u/vFKeh/mnfjLC1ikqClHX4H/L4DCiIGz
lEzFqoinswBj4JPvdHPIkC8qb/Nhx5Qc82aBWOPBFnkuTFsDzoVNLddLnCiZ2UBT4ztIwEQgXmSt
xrfPhsms51QRIWNmIAc6H4V4fbp+f+dU5R3Fl3R4XGpi3chZk+PwizK7WiBOQVB3eaxrrGMwIRaa
zxi8BP13rpqSV9O5R/r4A1ef8EdFr8YsFmVd2HV1RBVRk8aK0ucUVNvUHXV0DCcWz6urCNDt7eHx
C3ealRS1f/+IWiegdgSQV/C7q1nl1vkJqSgfwdoMx+R02/hfK4FdqIm4Og7gPLQD7I7CIE+Twcf4
737NXJQSJYGiEph6eNFWJnHS3/L5A0AIv41wayypnhITrxAFNgkFMgYUTSwR/wNpNTmcDzX3ZUHo
70PvkLUNRwDHsbrMIFEbXtLxUl6Y0uCmbdeC6m5AeclNKBO2ZHVUHvACPLBANxi5XOq/39JXLsRV
CrU73PtAJq/owqfA1NQl5g1h0jtE3AjC0jMRxzAULfyCwxE2pn0PAS2WnJj8H7zfR8GbDwLkMjvj
mKMt42/Pmz1xp0ilfIrYmYB/RO05buxwUac4hLbjNukc5K5CbES7m7WXmgJpBqBf+QU4G60HNkHt
OIUUgUvaFqnyOpn3tK1Ab2RcvmRr/iDsXkf4fIRyVNZ3GeIhqWqETuvUtfo74d52C1kRo2FbU9kT
XXnArf/lDLROVNrkFBGe3ESNesmdKUzX+iU/ScfnP+tJ32QmxhkiB3CqXkHUS2fY5jH58W9I5u0R
5FENFfrpefh5P09qAUGgdnoUrJGwHc41asAfFagUZkhGg+jX4We4n1wd+gPZrvgWbtVWUH1CW7s7
4r8eO9EeqCcnoAM6gbFtq36UFjDeLu/iOhKW2dST73yHDYoALb0+ZxpYnnJtEDmUXDPAIlVSZZB6
ltTr7La2xN486KuB/RjM1nriI0S54CmQtwZheJqB+Wudc+so2iaKzocOz34sIJ394xhUKNuG5OK+
l9up5Ohl5xjaClXAj/GUQaS8EP5W99S3uat3t9pJr/UhTHFNHYDHpCpPQ75jffW9LWBgI7Q3+nWs
2ED7V+nNERL4/pEno8uTxcj+dgm162cBb3uq6E/Z7G+J94lNSQFfnqMPZMLzJ/Hp0L9pKY4tAASQ
FuFCtfKWOJ63nb/PRZ7hSQTcSEZBRt841mM0Q/iS3YvvsRtvABu4pCIqu6uNNjPejyJPPw7RxDqp
iqH/AG4xBkozeUbJ6V9gyOZHX0iWP7JQOXUGW0YW1PWysh04PswSlOBoXDLBnapWQ9HDlQtGrf2s
zihv1ybseTyVfQivdawARa0t8IJto/xI0j83Ba5lDH8ifsXp54+rGmhgOf4MS//sU9eWGdULXVwC
ZVDf7raBZ0pUdnNO/H2YZnVrvV0CvnCOIZO2BHHETe1/RImMsqcLcRdx5QcPCPJvUHSckc0rcxlI
Sf3C8OFoWQOtuaLOLycSqZZNP/mnZj84gDzybjoyRhwPDvveTb5TKicxijHaqt/auuliGxi+h//x
75HMTRPclYpkaNGTVrINaoQ/aHvR29YrgaJoJUOBfNNPcXi3DcCg7T9vh2Z/11G3WavvJk/WRXSw
DogH9gaM9DHqBVsYG/+I+OmvBTbTLuY0YMnit96Le9vOdKu09KY/o7zy3I2iP7X+sYnziMWe+2sX
T5IqSV2C/iHnvgB/yZ1Ho9CLItyAtnj0tdrCjw9IahvZeFpvYpvVWYDzDEsa2+BPLg+QbT1CML68
HzgADi6NcRHD2HNxL8ozhoTBbyPRByR4tE2nSxSHZbEwPKH4FEDh39t7V8t+7wuACu1k0CKWNKiL
lhjdyBtfyPgIwO9bIgxoSf+pZYIS4/aCDH1WC/SZPpUR5FW7hUH/A/0OR9UpgJ9p3WzKuJDcHKJn
r5bjoY+ef+cJA1CqIKc1FihH78+uc7XTtW3Bt6HeqQPtiC5pQwVsEQb+xLVr9aVpzqB90JxZnq9F
eLNr/OpwahmjerjVlDbGB4j9Rbasuw0aMoZ8TVrKGDLbSFeWf0V/U5YoYoNjnezGpxppvcH2C+X+
qdqfsQOEaT2TQWTS+3ZamuEhOTPp7ZvbrIE1mZg+c8Hc+ghDZ/jfo3R2ZAIH63IVvXK1Uk6IxH72
iLwHNhWqn1L9Wh3ZUoi5F7igVVIRmH8vqK/uVeWdw0YyTClAHznDefEVXDWlYpK5zdmG4FJVKXu5
YDwGt5NVmYcj39bhU7vRHdJH2jdmUh4ebgXKnTpyqCYW41p71H98WPeTZn9/LuPl2fjK8sLRMBtK
n4bimV1awL/OJXPwAILnQUK47ipJbREjiSbnTAJNCyryL3OxPzkAokYEs9Y03RdsnpnT2/2hpDzl
bPNUdNrBxrV7ceDryecKNvbMt0WD8140wkvijGLmj7/BkxqzNxOm+hvWIkedz0UJlzXZtfZM0t5t
d7gqAKnk0ICczDZrA0aSdnXsf6iVIcyRvGULodILOBDhEqQkDP4c34tMMnc9fPbZf8Zk1C7zLxWV
fuOS+mbCz98BSCV66DPiOaMXE6iU0OpIz80scMAXkeuxX3wouTeBgpmRhldawpAVk6hNqRYJs2Ur
TRQ+DwjWJmxcb8KyqGfHqnZ+qyI3Ave7oCB0zed93sf619dipK0ALKinYRgCKsZimigV4acdHnx8
WJxrlOjSZHOf3PhiucY4w7eqwua+0M2yfCqdFIGQH5AwbRqfvk9W4ZB9wjVXANlhTcKCQwtSj5P2
Eg9QgC4tHar14iCsaVAgQ1LQ/+753OGFvNs3y6jikzWnIZ4e+TA49GvF23XmLPqxrLz3qTeRp8we
RyiatGqv98+gaezAy6006HKCx3PUh/x8aaLugRU5PWCS1D4fxu/vGPVT+oPi/QiKwysh3OkRoNRq
OZ3C9XxIZmS7yL65cLPTtzQwtL2X4Q0L8jK9A1rDNzMue672oPjIlLdCwDnqhpwXZ+Vaoca1EVbU
Ne4NySNT90CVLqyUSd01RVMOC2/54bGDdApQCwHmL5OeN4PDLIFOMBe0ipIuXydt5qQ7tYIgmnCG
I0bhUfjp93EPxqdlpVwp7FoaCHx3rrHjAch7IWVKlyUU/Z6YDvtaBaOYigpDCXqbXhhadAn3GQiO
lV7PVqQFRqHpbeG3vPojvrFudg4uAHL8rUUonZEL3qKFOI5dHmIa83gvEUJN01wOR2FICbv8ygdE
X2azrj9vaOZuVR28ajYlrzSXIaZpAINlIeire1ptJq7h6N6DTo8J6WYgqrLWjKSqVKAl8YCNB2b6
I4gq274eE6NS52QBQdFrLe2I3mVE7e16H9Go65wbE7CjECFgLDrtExazu6syjfmJ268qwOJ66oYg
KVnuKLSvfkaoHxaOnZUgWaIqki1mz3XMIWAjYW9uOHTKHVFX3AP/gqGrrnBdAUITY+c0qDjSMCWU
HSHo372QP6YBbMmFwBOVcT/gwi+/klpzsEKVzrQOpguNOVczVwMSjPwORDq3DWgJXf/+hMxFQ7v1
9uYXQcvKwWkcbbq25PJPu2nM61OOpL4NHd8yFXODz69Jho6xt82k4IQCSzMbcLRq0XSxeGQlpaZs
oWPsid5H+csZ2MDfYGcQcnDCxtn+/gOfsUayYw9ppjt0gVG/qQFCf42nht/pIQr6b/JgiLiLRTvo
LKKgZXxTKPhyjAm2euoYSWvXjt4Cz0C5EU7Nbd/i1P9MkY4RTLp4DddcVvWbM2iTsP6f3gQfZu9a
TZpKeiLCgZJg3J7agSlyRJZFJ33M9WXzTFpf4k5648K9KpPEpbrNYuDNiacHO1ZjvlRAq+waReUR
//MJoTWe4q2Nm5ETN3+swc2ect6eTWii7S+R6A8zNHJBpTqq0225yk1e7jAIiNmP5pDyUOBAuz0H
CRgR6eOC90G+TscOYfdaunRu4A2JiZ9EPb1A9txvXqgywhwHP5N3JGOqv2BfkpKjBUDxz+SW+itF
YGYPbC7tULggso7XO8cw0ltVQWP4WfL2XJNSQ6pyFdQow7fUUdjWisP2eyG4MgaM0ahFQ0f/5/0c
faVldNKynGe/FuyK3OVXqCg7xGZWzgsBbkpNUk6ldV/RAlXqE+bNMKK8RkM/vrfVmOi3KNG2TqE2
APsooshg2l3EpVFYy5wPUnGOPNod702UVSAK2zoQD5YrIsUUxvi1H7DQVAIhEomf9KExjnBYQUxm
pr4DjxtIoPuMXTrX9g2kMdB23kAQ2IeVoxdZz6qstnnG51KDiFA1wpTsFqwOW9K5jwhPl6rZlEzO
ikJa4h+kI9WjO31LCLMF63Jv/KjJlXwoZYBT2EsZ4hqWdfPwNnACOV1IC/l8Gt1bwqNz1LrMoqVU
IifavYA3gp0JdEVrlpgFG+3BBQ/ckoS+WO6gOf4HJVJl9ZQqPM2aYXPMQlBaQ49lOnGHxhbUv3Xt
1cU+Lxf0klfIndL+Q1juVIwAPLup6f2/5vbQGUsJ00OvjvHszsNyVr4fgtPPj1WduEfpY9zqLt3V
UEGoJ5/oB7Fev9uFsgDXWUacS0MolOThLGILHyloB39ghDki7X6ptNi1WxIuKYvZcexrlWaSMkSK
U1RliSUy4+T2O5okIm4q0KVmn8z+UpIzI3zrGqzKcVrFIhKFOuXE22z2Fc+NbIe394thxkBLDXER
7Eu+zHb78A744P+vLIwIbtSh/hP4CGbXh2oEGh1K3iW36fFWX0ugTWBL8CPpIgxHyLAWYyrmrAd5
gUcUOcEOlUrwPmIZnTowo6JtEAhAQO7EdOR6B/zIRigVB89/AG94HrVHVXQk8we/24jymPLbkOWd
nIQSKTcCf0udm2rWhrSZzVpMctkSjg+LpYr3Vj2YmjZCBhU16qOtGa5Pi1dvqA9oIYQTvfQDDQA6
uJ6DTgiWq4JML5mIsZAcsWhXujMEJV9fFImbG+xVMMlpVslrEOqdX/8R2Oj30ZHmNYtGlTS1mX6j
OOGmvWZNLH9oEZs960XXE5a8Zdy16cIUXaR3Tf8nAI8hAhfjDvA/WEXg+xltK9dmg8BccELHBZ+j
v2qxZHrdd/mt8PzEtH4RyZEK1Jp7cMCjOOx/EPNq4Kz1GSqOk142eNFI7axmMbH/a0XfqclPHko6
gHC+vXCoZBZPwuBD5jqrDnC9hGL8kq3sRKdTch6DoDtuHwewD9KmJQLoze91taQDvSRFNjcpx3W6
UpsfJZ4bd37LU0WggB3jSBPm42JptfG8no5jSsTZgGyfMdDvUsxipWUEztMEXlWHPgWNFjFbiJq5
8x74ygcFh0vBK/BQhbcybjcKZ5RmHvuwS9FhsTR6LN5k2MJ69DtKyFdMCn+qiDfOGtd46bJbIxBh
It01c8gZu9eMrhzWEmPTp3b5ZY8hfN4f2rXpNPfqsBHh8rrJFHkaswAcDXaGjDFDgjIkEX1af394
BorRxXtwdyhahC20IbhfCCUmFD458kayDaDVEvAt6qv0PnlqSmuwomv5tPYIiKXor4UQZIc/24s+
RN4EWXMoDI4l2MC8Vs0BAet8BL7yF4r6szBgO7PhGgWlIGBBKAwY5qyQ899s27yWwK3MQG95ZKhe
rtBQLrRBn2UD2i10mfZK5tR0jACPYne+uUL609+8UqecSQdQcS6rIgn3PjR/bQKPSBSCksQGY4vc
/WpzhJzt7VvgqH47iYLnb7BqKexjnIq9NkSGpBF0vrDQgCNtiFzVmco4MVeHohM8yBdyPF3CNe+7
2ABVqrTjr2UPVRCcYx3cXZxoE/t2DGmvVtRlt3KXFr3wG+hm0aaldXxcZoY04ri8VPzYxSYh9CmD
cfMJUArX+gj8wkGMT0bhW128WgCqndmhu2/Dt8BPRQVQj0euA5wLLaAjcDgfF4i1SDqBLsmzYpzj
mX2nFnBA5mt6Vkwl03vrC0X3k11gFPi71o6Lb4TvWORoPh2rcdanZDY43+uGgNPrEXpr6aCA9MZS
D4taQLL1rVcBgymWghVKxkHi4YigmtRxJA+F4sVOsEj9wf6kXt5nQuiuXt7abPslH6flz050Vtke
88Z6FqkAujlX+8fpCZyA8HNIXXVjP3rRrrGgt54Wod4pjAHAflVZw8Zz46Q5NYgHikYqC2/ExeIe
ft0NG7xE6UUW/fkSfJLpIvHlokLBdqpGNn4X4mgIKGlvME7Hv8XNLOG39ka5U6pOad7JEaNHF3ep
9mRJxcoIhgvN0Ssl8RUEZouhMEIcwMAMdROztT/m/MucTNFKIB7cYa4UOGQkiVVOwID5OpuaEmAO
FQsyh6jGwoPMUDcPHB+vnGRx4+Aq4m2oHfinreM45bS8SqYduh+AbHahZzgtu+UMKs227uwMtuYm
lD5Z2UTjH1P8t+nxUofciTCInWfyWjRdUn4wN0wYfr6cq3Nr9qcDDL68uKVG4xEB4z2j+b9HlYJC
N74X8O8QFt0TAgoiwA5mSYfav1IrMy+gcly3gBXW5+fc8CSko4qwU1ZIGUz1qFD2Wy3b0OUfk5WU
cCBS2o61sDJSQiO/XpQ2oD10PgQPpqUzqBIIj9Edef7UXzasZR3uzrid+NQPdXY/BAjnOPf2/Im1
SGD2FBBCeV6yy10fpJoONRmjovLMJnk+w4TDPxi1bsNG6g0CDTGVU3c2J2KBFjCFqkzX4qyhrKzX
BU5esodtYDCz4YD/6JlkA2FpueyU4zzheDH7bE3CkbQBIsQW/07pBjFa9q/LgAwuoMujePeytE79
Tf9g0Dd33N59EvQbKx/ji1r/qwdEp06IA3rPo08CeWGvEXIhxKhpoO11T83S9vD1zSMZzVsVlvfQ
1BS2ngXXSRDHWgPhvc4gok5iXvG9jSTkt7AU5TA4e8ndVzwmtHSQ/JAT1OF6p+PNzpo/iMaB01HR
jU/KS4s/BTfBk7EPDYMdjsebiY0Kd3mlpTfLtFwJDCK7SC41d40g8kW9i+QCuf3bBBRZa+Zse9Cm
GmxD6vQ1HEOr5H6DMUPhNK05gEMrAfkdwiRhUI9B7WbprrSGzGZK1XzArihbgj97OVXXSMpIFOD4
56SVFSo3t03pcUDS2G7pzWx5w47WRu3j1uDJSxODAqAoAJX73503SbNvU16tjN/yvbjdDmxC1Kha
Xs9Yqyp5lExtifKvuieMuM3XpBiN7CBdRcmU+MJNv1g7QTdgncVRaZSRrtR/qTbE9vukDRwvyiMs
Fv55NE1Lv+01SOxOstICp+BmBE9pDMmKzAvJ0/4yNxQVuZjV5zu5lhIMs0M89gzDs5UslbOSWCHx
Phs+wfVinuZwf8FPqZmGZzzDhfhxOKRXitprVeeh5raB2T6C5JP/Cvvubd+a/tV346jIOvwzouoW
K+Q9amNgD7bhEKQh83CxaXZIJOXij85vteHZ062D2Lm+95VDaMHNG3VIFtY7vVT4pbOkr2YJ5/es
UQ7AbmKmjwvK5NnOsxBM1lWlH/QPIbn7Py7PROcGsooinJ50qQ/5neQ6Wo9xCsjrMjo+33XAUnNa
kpScHkBQ0JNko5iOQAe486mKfL/IURj3L5ZOBzJxhStLueW/OeqzvrL33V20wE+/mktwSskXiQY0
Wa6zwcHqMWmi8NX2VmxUMBqgA4C34j6wIvfmlLSLWZAIwGqlSjkXhDd0Kwh7YCQ8sryXQjoyqYON
av7mFCwdBr352qfCUnyRdvHvxzMyPQeza2uYFvfb3qS5jdBRTm+WkBYRVcSSLtKgv1b9RUtoyrQu
zUrOqxnRORx0+iDxx7aHts1mw865y38My16BQtTfVI4VR0MHBRuSI9+5FLHEe6T1VU+HOau8UAli
94hSVg3qj+rIL44LwQvt7OzQqFLEaXC4F1aA8Du3XPdvUmYjSiqVDg+vUmX4tnVkoe0bzoxLH/+o
eZKvf5Z2CxFxEX8B0lyfCEvtmtC9Vp24CQouJalbS6poxTF2HqMxuRUrvXrvjp5Hc49njlZz0nDI
J7/mZJwIzdZtmg9LgbPyGN/DYo6eJncwjKOyK5oMZrE2tuLmzaoyBq6nl0zPuZjKAoR7HDvnImEj
EtoErDGTyrZUTDN8OUxDozJSBXsy8iCmAABwjzt+L3NUk0iUseFw/KM3WDss+7aL3KoZ3AclzrF9
WvA3JTE2tceC33fE8KO6wiWyA8BYOQlXdsgM+gA2bth5bTN9YuNeodKpcv2pN4MHbxMkVt0y83fh
ClrZjjnwnVPpgJkPwmOPIwQqi6p4Nmlxzk1jB+lBJJ/lN1oB+qA4QwPf3fkaqk6MvbeooMgzNJhb
JR0Lh9E+GQekBL0zq55s6zzzPDfaSLeE8Ydkz3MpyhI+LLWJt0lGD+yzFRLtweWO79i/AlhnhwUh
iJ/T+QfSo8fdn22O4+NYflexQOvti2Lp3l+KFMViJzIPqzGpx0qRLIsD9AEcqdPSG+9RubFTHJSN
wdh3ZD30z19aCnt/BiY2KqT0OtWQqWGpYTAZ9H7q0+peP8t7U8EhdlP9eNPlsRi+ipoXfC2d6+MW
AHJWROkXHBvoBuuwpYm+g1JLEvyq6xuscY4LW5sim9LsmkfB6do4Gyb4bKwAYwm04zu4HCU35Og/
C6A2+7nDE8cxrjahala4qM4ALMYhum2Vqdk0DeRdinJ+M7b5HvR9CPLtY0gh+95PIpLbmJuLdnNr
a2QEhVCVjgTPsUotn0N5FX10fpA5LLoL8+ky9FP1/4QXyuTcuQhFkZuJLzomuulzhUgOV6ZRmzp3
bCawvhGyOGJVZVLxg+l4KCImsnrY6rbQYV2t8+VQzy3igVc/EXkwedFy80dxS1jso2wqgYFVu0dX
xMUq/hAPrFxRsaCp00MipNTAcOPvXcLvLJyn1iIdKlPKWP1//11r4l8M6P9DI4ndCkGJ1blPJUqN
z3Z3flWlNOOPEmIZQOacu6MR4cktqiVZJOaaKp89/qThNNK6HJKruZEfYmEzGaWFoz1a6zlGv43e
l+BrXx5ca6Rzxyot1wIwWcX6mXSnxDByg7mqQwYqdceqArpc+yRjQaG7JSOyL94N+UrK8Klyw60E
ZbqMPiu5/Bt14PmQZK5Y1oa3Woj8a9aBHI0PVmbaDkCnptSFBjvfnAIhzF+J/5OxQl+hjfbC+pPK
ZkSgLOv2VMIed8ThfLrJPhF1jY93v3bnejJATlw2F+//JtKoA8BEHHtLW2rfPe11PC4btq3aynm7
KkBwPxBjEf07R5Pd0S+vjlkXYYyckeFuWTSznN4xXgJnGrWOMumPVWmpusIp7c3KlFWt7W44cj/d
d//uCZ2JUP6GD+aYEJlUAgPebmTvYHuhmQaJHI9ZDzNwMVrJBi/9JVo1Nd+gKS6hoomHx/L7wqsc
AkHGYqUPiNKcdSJI3WunGDKKRod/P9uKypzanfQuzNt1kDZbvqBV4DGzAmCXOqqAaTLwVbKrNch+
rNddSTipMKJ7MalqyzHKyo5ThJKOvJIrp7tinyUfi6rRmmsX30KOHOxQgznUBhYSr2JcC6/DPoRV
4ZTWXXJL8Wr7mAk/iM+nGvk0PGspfFLA4r3YzttdEjFmrojhgNFGVYCpy6RYRdU575DiUhAAIbHT
0wwu7rsyXisK/95ndFrqsYpsgHQWbYFKnCyUZPXXKLPsJRmQWw722gfqE9FWkXmDOc0IjNDgrcwJ
5rlBoqEHvaLNPQ/oHlAIYLtIxCddlIWOoofFWoZBQxaYpaPiUpW0kS0iwX1Yy2LiL0nKyCN3tbsw
CGHNQgXM01mdILSNRPO7aq1hiPyxnaMSoAopSrRqz+fqpwuzDYB8WrVn79vFDarP85os7P1U+lF0
+z6chLEfTCPfnthpW5YicI2RBymthCKnC6fiPUJJUNJic0yo4f+A+IPr/IvPob0kzYWacivyuPFG
AlUIUw0meyhkOzSA7RT2cXWIz6ycMpWYaN3aE6R2HMFcDhlwjofMedikrPu7FKswNVZy0M+cJJit
7bUhqnbhjs7yDRB+AwkXA3g1Sx81pvt4UTSYPjDMpjbPQ/bZWWpChRf1UpVrJsEc3PxK0N9egRnR
lP/Cou5/y75PEF4JYcSGU2ymW2XW/2jzp5N8KWXNDKsFyMOdyzKc0twEobsX4IaiW7EkC43o7GUm
1gBml7Qp8Xuz731HMeBXGwMsq+I6NkVZGozTYLNjx4/v0AJs605gCq1Gyg3yvut78xzyDtWdPVTA
YMU+YrK9kRsoBenutH+3m47dIb0JCVeRelumHa1l8zxQcLhqCxYYtXrbAATda8vIb3JOxr0pzRCM
y2sdQvdux5qr/2TxevCU0bXVSNMDwZpb9eCXlnW66d/qXwg95m2YIQOvW9gsTocRLzvXpd83iI+L
0ur+sgcW8LjdSoWz1zf4fXfY/H8WvdOSXEgUKza755zujdFBdv6wxkKNJKU05DfFD4w/JmxVSF+p
eMg7iOPEA2VnrslR8hGoiMQu13tiUNzVfdkKNeXMtyw3bwfF1IFaZTJXU+2pIFW4zqSeQPmt8pEB
A8LzVunktovVku7+t/pkcyNeMIEdqb+WNTB3CpPFQE+3gqwavVr1eXrhEGrA35XH3GYRuSMSY8t0
f4WOQLuaCZELMJSxiBSvKwsalOPLZuxreTHzBiRVrJKcRi1t5NJQXMeAEeDFhGxY6UX1rbV7pQ+X
1AM+Mp5t4X3Img3TNbFJXKhXvJKoJ+/sKUVj5f5GKB7AQee923Y5w0UtW6/SOXYNbzU9exOqfAoi
hEC61Fzjtym13gRmje2irW+w3Ur+rQB/4qNYdetuY6HdtIxNIYw5Vk3YoybvQId5WcoL9pl2svQ9
33KXpCmDIYYDtM2eHWVxu0Fg6c7OHWD32uY3eAURxS9c1xbPhXTPzZuKrD2GjvE/2mvrRHPRpWJN
be/0gn/UjmPkPxrGgyFJkYlkLPwqapj03grJsGHyd8fxSdTGKv2/RrhHmjwVpDGEt40X8fuSp3Hy
0BmEFzDZ+9Y3Q1PWhRW1z0NS3O60qIimixGv3SDYz14u7yeL0PZpz3CapK7M8MFdtorXsOWpEJqB
LUGLqnLCQUznSfH/C9X3eKMuw2eIxl2+NVqTn6MN0s/zPXVYX0ShPQ3uKIvFWj+ZHFXc7OiB+Q0d
FJZUqlgl/o6R5Fs64kV2f7bIze0WeE5HmITITq2pNevZw9Mm3d5XJUqPhs+rdmgO58QEOPe7DB7b
M9w8DAHbMtQtstEl0vskg2nwLW0Uc2Y3SjvxpIarejlnFbIsBU1r0I8k6NXVKspVOWMl/NtS8s9+
5JhFa9GjXSoAwu4q3RpGe4X6NkUeHlh0t4I4WhNZ3OWAMyuxHmS2qURKepbXDTfzD8WLU1Ya2hX3
3ifbpUQ+2yHU3b3ODePk3oGW8LW2o7w85b9COOsDqGE0ZbziYkDccNitnbQ/5RDp/0tTLZ8e9CrI
iqoSaVvfnTsHZVLFWAHIVS9UmzcjL8+pkPiu3pGTcIe2ogBqPZD1viwpvc6am6Pi5W0yImKq0EdM
pWyx/UdxpqZ1uqonsEu+rWCGpuer/cdcWTpEdbc0iLByoWW1CGjCf+4osX06IWGyofwqh+Y9XWSv
JRVwj3dWnVAMGc9F8mWGw5MpHmfT/LZ/fNl2oNt4L+I6TphFmVCegWHM1+Ya/2PKll1xmiZq5ckR
Qm9/5PEwpN6QyN+ZcftFnlJGW7EZmZIbpCF2yjzbDvNs1zRteXVhrK34bjUu2Iw2CyG5v/YCXHIc
vfUYCwSXcKiGM/Tg7jmnD2v2IxMcKhebgrzk3nplQIp9mkpCmMt2hB9+diYmg3xzh55lSmx4LTIm
Rbk6fYxYxwQ+r4D+3fYZISNxi49FXBuS05gpr8mJRVqvq+8boHVt5gMETfX1a6ql8xuJAMzDk5gi
Z3SUQQkRupq3Hr4AA2lmg5Bf+45izo1curWGBYEbcwcdElfoitnMJTAAuBmvkifwPwd8r4knvaDh
/lSq2a8Nuz91W8+p097Su2ZPPhSAfwWHhBry9BzyK4+HQFSAc3bVUgmwIewqAM2PhK5ZM0dkKU9p
ooYWW5mfnWqUyN984Zc++ZuCmpYsJ0jBbvnwZAM2bO7130eoM9HoPJxRX4xFdfnTrFqy32GSDrbq
b+bIUrVLhgYX0kLnU7uPV6HAn+QkteJGG9Ki2O3AZBE+4oKLfLslQGs4riXDA7WVSnYey5Doy5B3
1lV+opQHR6zeA266FwVIpm3RrTy2ZYQhSfq+0VF8CoTqTx9SBQ98ZN4IC5C9p1fmAkTL+83YKsi/
m/3xrcSwHEIawd31HL0y9j+DaRR8Lm3wPnsoCI3KRg55Tsp4eS3oMi8Uz/AWkkvputAI9lH9Tptc
OnMvV7RNsgobtE01MGfY6Rzd8bRU4fIqeI68IHUMKIFUoyoDBqtZf/wXBSQBYXnoXaMNLuBSqYVG
c0r0zn+ro0o1Eq5bRCsf5i1aFVvPXBMqgdxm8JPLwHRc9xd5+x9sTHXjIP2So5H18Zy87Y1abuTZ
zf3ItcjCy+YPSWJkqa8kBCNEkAlcF4FDf+FCqsgCV6PRdXTqod8vNdSzICV4AsigRbNsYmeCxkHF
s8aTpiRQOnKX+KYRZLLokclhYb6mEGrR0EA4/LS3uIPQubDcIZHIA38M5dRaEF+CfO9XXsdHyEYQ
FTBdNdqr3swlupGGzyaIkd+TL75s6hX9P/WSiUzOx2PXum8fUJt6UqH9mcoe1A7LTPaZJ6Wi6gtP
x4Ike1JxkysTdsZ1McBqay0DS2OL7DbC61pPg/Umfs63YFszcvoINac/GHiNwf1uytEKb1hS088D
rHBKFnQ9I2al1x+3UpSHw3RBXTfNwomvEpV3ThqI9H8Fu85NC1+7dbeIyoYOJwTUkeZWV6CetcXA
HeEjWryUeh9+iLq+Oxuzo+gjdf/dRLJK2heAkjYKO02ScZlz6UGKADPjN52zf6xvrzr4RoUQxtQu
kxoEfr+0z8NZnK9lw+VY76XZgn7Gdjp2xvKuGl9Df3ffleuDdH3TbWQguFk7YbppspwD+4HehvT4
S6rExmx26WHnuTWwTqYRbBeCgDVwfZADcv8oTpw5jZdGFg2ODp9xv9wFf7+u0yktgGTvZ+fLQK1v
Unyje6LflCYztzSkNCDV/EprT4KaZAWrJNuC/py3JF1JPGnBRE+fMlnfiWS9dospLvB3gBwP32NN
dFHectnCasCHwlUwmzpdWrP5Rdea5o65b/6dxgqIHHRNWeaxzrVZzKvIeliRBGor154nKeaUVmdZ
Ug+z9fqJAG7UVQs/8cnOIghPuJUTcD1HNcjl7j2KYsDmSJshPEgCrVAgFJyS7QBp7MQwIfrFSfap
R05neZTlqqLbEZkjgMxpudXKfvOZBR/1EAe1FYdk7oRXyCkhfpphlfkyzoTgwSkCHrNaLSWoNa5t
w+B282fnkWFsLixTE70U0EDJUVHYNG7UNdGWfv6ervFrimlgg5sNDsYD+b7P69XOJNtIqEEwpLT9
2DtT8qMlyk9IxNGAV9c5YPKEpQzJBfabJcSBnjhPpykfKr98ixVV/DLlD0wdONrqRBVvYOI5Yj3p
hepevz2Yi/HfVV1dlxAK/YUXjwtO5qcNiYnuF01A5SdGzK65pX8bc3BOKdcK6gCPPfgQcbvFh7cR
XI+rn5BEuy6SQazpBMI3h3XlPUVB7YfUGQQ6eO3z4LJfe4iEgYVA4mDIspJOkJKxnx0w+9sBgP9l
NInCiq6YP6x8Yt4GlsPfh6py6oXIQl8eAEZ0fUerYBvhS4Wvq+PUB6YKykcXTljemM3NC1lJh6aX
vTAIUrS4HNWLMForYD3dDf2mZz89HcsFMBib8skqoRGHaH2JyMMtHTP+RdqGp5T2n9mt7gRJBav6
xKCCWtURqOtKr2E/uzSkKOdaQw6wZIaX8tgrckgIpZ8gobM73BJ4AKvTwYlRBbQGqdkeuHMzS1a5
hCc4KVKfvlDmgcRnFTyc4hsqub0YQB28p8Z3ywnFnSfrBgcTPxA8jeqB8da8xR/XRLqAfsNdHA/r
PPKGB6bReTpYMHy3wj6N6TECoXKLeXJSvilzuMEC6O2FuPd9m8saIJR04oxF9X/vjQJwBA07djNb
TseMU+bVlmlabAzpg6TUtwqFsQSVR2poiU/hWORVqYQjoe3KX/aCOKqrxP1bFrsWNCvwOJUJfoZs
drtSe9TucXtMwSqqyXrVT4kPbjmgzKb/WDOGzUmum/V19RLSxtIBAqh6N73PdLx2Cv0d8y3k5R+g
F846MvUZ0J65sco1OoEv3sG5aFM/UIR3scOO7BAM/ty/hckAy06B/3MmSnbJiS8ZAIi14vTcndp7
fSo+O9pktwKSP+XZQ82R/Wogkm3+DWbUC+DSLVWXmCcLd8gW5Cy1hVOXGym1+i11CeQm8Wbi+jSx
E+/S631b0CaKUfboJjmHGMG7ybp1Yk/Wp6djEZefue0SBzi4c/xlMCmTJP0t+lIrOqDfpX7+N8WH
wqP1eNFftn+1izAXvfzbVn3sFcYMKibR0w3S8S8v+CRjVrFHnJRN4q8tjODOiRGVhI4XJ99kaoza
RW1B3sXHKPOP6KcTM5yiDGUmOoG6CMZhrqfM2ftllqwwL+qAZXuqYiC69msHkd82a6mA/2VJ2jxy
1tJGWl7vfPf/mgYHYU5d60hwYvm+y9aH29RJYfoEeJlnDkiQ+orM5UOgtNCuG0eilMqTaJsdYjJd
ix6LBhsAKpCwNphSfdaMlX7MEAvzIK0JcS6s/GzwZs2RAlzBMasn8eJong7cid9GxWXwWBt2XsDQ
zu7OjEmm9Alggom4oKiwGQhGAtO41ZRXdys4dxPpSWB0ekVswpupoBseLAP/xbFtPTeMaJTk/JPN
R+t8ffAyFhc2k9alpckiPj8y65EHDMw5+2sV12TbDqNnZXS+fpwYvbn+ZAXiznUrw1ypXp/DIrio
acD8qz2C0GMe8LO5Iy//ARr80T0pwm8XBAIMsA/PeoA5Un3/HXZXg9bFuxVVEKH+z//fz5TuYzU9
kg+V459dRvaR4QTgBpEkabdQIVphi3Sb9KIQiTmquzSswWccckwL1qsrOupKMFugVE7S3rMnk9gK
6zQd8vWp4eXX3HGQTPWsqd1PReF4LYJhmYR8ZhLXfApwknrVGE8f0Iiptsjb3PGy1/JXv0usTTpe
dY9Mbg255U3t3ynxk2nBKrSEfG5oZcrOuqvZAXmiw8ZCG2YOxs/PIz5JmMs1hO/Oosqefln1kKIE
KYnhscIibPkmwiFug9/4yixkIT+UTKTjFzBQt+J/uHGBmf7iMcQOoPa4zd1VqbKNXxf9FbK8QID9
mColjOSHVESaKGDxX/lOVqVB26QU9khFD9gcCEJECaDAbInJF6X16P5N7IXgTahdkL+rBIkGQB+F
0s8YYWE1Mfa9D0iJ+UJki8l4UfYEcJGCw6nf8vCgfGaZkVOmyI2AWGaaGil0+nD29zDkMAGRGWdl
F5g9jFJGdCTd59gVyzafcYqkCpl/WVfW5OfSYxvbRDpH71yXWzR8uWolnIsKg770UGhaT74qSpeu
9ODZFdDkhQDXwHCbJg12DyF/c1M0U21/2egRIZODIuwZxJ4KOri2aqOMQ8Fup8SnjanfIVzeSZ9n
Nd1GTnqMMShgec4jwehvGFAsb/jtlOESrHFwaeNTjBnqO6HcK8TlvVdoGu3HrCwmhm+hP0ss/WFr
SfY3qaG61glbGrQFEw+nA3O+GAlKa1kKmDIpBd9iJO/1LZWjOq91R22TGWG8ta575mhiBSn5i+M7
NE8jOndgkr9HFcnaaZOMd9GoH6ydLC8M0DewsHaY6uXvMmUD/7/HeZL389O5XjDDkL6CSgdFeAc+
hEiO+M/5Fbgnhykf/Wwn7s1NYXvz5Q3HWhrmEz9pRWn3pW1p1Kdbhz1j3nDdz8cPzsrAYexx2zGL
tsy6wQTZPnXl4re5eMDG6Qj5y0WVZzbUUSYhl3UuAS7zbzLTd+yMGNZPzMuGe7p9EKcONSzx9QUH
kNnSKLE290sVbj5jFCr5k6IGUPHuOQn86JqdE43iqxso0kXKzF0kr62f7hGmRzTUvttftCkCRAYJ
nMiWhgzIhNHKhlGy70IIqoXzKM9kQm73acUW7DC77BYey6z6ioeCL+JdrldMAPHCClXEv0bb+Nlr
xxjfH5yLnHm6NTvijBKlMH++MoBpG6525IXhAL7eEYaAgXJDzR9KVlHr0+MQh7vHMa1iT/BAUD5r
CwdSdYUITsrjCjoQ16s53Z9JwwImYQfX3mio8LDGhdv8380cB+p8EnjcT1ar0HmSB7NEeSZQU/oU
CEyYgFaHG+esPJXeLfTbrvtzNGC7Cc3fgbhib3if9MHz1bXts+czjXAZErAy7D/d96KzEK/z6Ly2
kSLd6M0K2oYuxj/JVtPUsf/pN5HafK6RN5I7GxlNuYMssa8nDa1AElkYc5qTzYWr+aH1pbbjm3ma
tl4/0At/si7u1bq5GJGYn2/AtAUGt9mRFpkGXbWfseRZuTOrkfKfd3Rh4fWkEpkBjWhtVtka5jD3
4BXX+5sSPY4zLjXxtzT3Yrf1RkNRLBStkqaiX22mCvuPJM8FKLCLyjsCSQY6nu5ZG0PnhoMpzNKW
l+enfM7DC0yjhJw2vvnbNMgFffDnrR19HA5J9X1oNTIFDBOEZjs0LK63s0kUF2FYejTiUB0LbUer
JeRycrmTQiHVKuSORkHQOtvM/maZbUXzqY/LaoyZs5j+utGYlkpojqCr6qqxZSDSPnQqlwkZlun4
4lzgyV/kYirB6DeF+P0yE/dyD2cUWeP/dddDns1oicrEgBmlYvLZowYZ+ulwIErGudyvqRuu1QSM
EFO7aM3TfXKe3524bcGvK/9hi/KOqt4rGq6dGqBOvhQpmm8426gpwZ4iQsql1q/4LkEbwMMwPAmq
H8P0sZvtQbRt4xC2AKJbovseCAyVt2IO+KEcHUKZ2HxFEXMJ+4VzRHsaMEZCmbQs7PFW1mPvOBBc
6Pq6iYB+BdG2igePZASKWCFrPRJnPPOB4riKAI6LHzSsvLx2yTRMMEWLDNqOgb5v1PANTH7bMphN
k+LrpVGertb/MCopmNQzn9gPDF5Gd5HwfzHJLEeeFyKQTcj30eU24MLtzSX1Dqjfgx+HP4PIrPKy
HWOnXjvf4ePmd5fKxTMj4mxWeQ+ATotmqMiQBkyGqthmctmBE9nBvw7jZsWZJr1DZoQDP3OrZHp8
3uoJiCeXG4+9bXMCoKYStoRu1lv0lZUeBKk1xUql2AxLU+/CUVG31//JttU4RnT0NkaPf82IeyeX
MeQSHZqBQ5m81bVIaiGyocqPcqiO5KjtdEEN5ehdxzXjHdaqyVGg6Qrg8vrpflyTPNPTJtsrTlkc
eQCm2LZJdG7xz+rebUy/ayse1UXrXCvZl55/EWXBZsHEM8mUhvYnaPfq8vOOTXK/+Gklw41MaG02
+KNhGRYJl1TJ4jd+ki/FDq4HPRpPPHxia1ILucMPX9Egt1Wc1bzgUnRoMekDQwlkxcGl497RAtjI
8/jHTeaMjtIKMYHlVucE8SJdr4n/X1LQmnqiNqEjgEhnVgdWMYj+PVgH4V7TFmA1boRMv9ul5IDE
lmlchry8CWDnJ65viTWUpU+LJY/Cglz208wqQvOtrUkfyEIMTz6Fj3wAVjQFwt3weDqHBtlVdHGt
hv1vv7EFH7va+ynlpMJ9DouA/tjXCcvX373QbRswKGEvH1i+ofu6tDHC3jHhRVjelELChncbrXnR
J7cXYRwJ/tQzPoVIe6TlNXmSTgATE1uMNaQCUM7nXZXWlfEojXXAJ3gt1pvPpXTBFGxtJc6pF5XK
lj6NUN0Jy60U1Fkp4aT2v9MNUUHH6EakyfbFKG44IhK7JN99jes45Jy+wCvNKCut5gfwpgx4seW4
zKwFwLlKxGOsuaOl0mbGSvPUN3jR1O9Gw2ENpOKQxeI4RHCji4I+RS3l+udZvKQg6a1O/mum7hS3
/pRUsybNcVpIqH84ARjNc33DL14PdrOLGBjnQyUwzZup1MB5W5zf9w6RS977RdMz8BTq3xdYXrwm
tQ4H0Vxhi4Gt8gTxY4f61mckolirSRPKeHoICljCeF7EfgAZaIRp4LKStYquqCXmRZ0Ofx+7ReFy
FiitwoPVQtOT6S6QTDxgME5QiAhnyND2svPF9KYma20ChbFB84jpbKRnPAcr+/2zO8kG85B9+bq9
76W2aiS2imOUfQljfhaRMA/gO5GlFYaBtXSs4pgu5+U2kt4NLeJcdokjPHWwlQxDtuinyKDcD+UF
NWBg2eLSn+RTsUVkYh3Cqv1CmBFd/VWqYMdW4hNJDZ3hhwRLKkTfyFH1ywuooUue4yEjiWAONGlo
ox5GQoiElq+YSI75WMj2CL5NY16OjcUVa5NgmtbvGyyILGJjuBIHkZiomABiwx2wYFHWI2/qrUWR
GzNWywXKB/T0Hlp7NYOrLFIheuM0vp+7FjSPcp4jdilFqvknu5vjv8ROz4QX796mlbxkAzrb/qs1
aP333q7fbQGzWECWJoIV0sq+55qhTkzcuCASNzgCC3xo/i3pptoZXNnZYMWGTFmy36cLiRx6EbGl
vZ6/YaovbFijXlosAAlrrPcd6MXnLxezhPj+NI4vZBC+xXzZRe5s27SwKL9hYxyfaiBAXTE4kAG0
x51Bqx5noNzrUQ33HYLwArcx/eglqd+W9hP9kO0dRRZdOAvHeQAgVCatI24dW9kEodgY5FqeJElo
kw5HXvb+JqUQGgEp8O0k8vd4XkzdnV5mPkfHrJvKGlIvmb5aez0q0J2F8L1gBxj/bVpvjX9DwhXA
5chZAdezKUe+UyIlVJ4hI4+c6RjcJcygumQvuKcFOk1DZXbnTKDrekWK9JTPtnC9al2w2DVQn2ok
asbWSImqtHT+mHvWs5WMm96V93TUQg4e2ekgwffd+LkPoAm02rQYm2AzU9M3AkTkWif7F2/SJGBO
TpFbdYycZDWm/zNMWFNKa0tatVLzvLCyaN/hJmTiJWC+4+i1YoH9OIoALfzfxF3w6L/VmLU80iZV
EKjPANr4zAzq9AgRkd8s7kSDxbmqKggJbtg1iBXiuHVeQdegHs4yezazFZMZAEI5WATq56MaROMY
qfZ5rn46m8sSQcBh0DIxTlgesGNM6XZFJ/vIt98AJm0KYRtC1Q+A9EVA7Ai4aPcKxyaBFKapJyMW
8s7ua8ggTXCFwsXSpbKEECTSzmUxxpS4SsggGLCvcpVhMj5Hjskj4g1t1ndptT5oGXVBXupEKxh9
CYl4sPvNSRrlkOKHbSDF/w9GFdnvVi9FrNZ7vMEOIxhdA1ROiMEkRRFp9GHYBZJewRQ1RzVGIcMf
XMPR3icLITCtEZZWReQUyeApVpO20aacUeLV1AceFHMiKKFMLgqYkndNkHH84Ey8pwtgY4kZ907L
mp0I+KZJx1v3r9wUCxAtPuurODa9hHa2Zs8Oht9b3AD/j6vPFqsFH/9keEaW95boMeISnaRqumka
HLv+lynS/IDUeLOdhequF3bxbbwyVgUsAgAT17eeXj053ZymUtrPwYVQkpoiAkeBezpVu5XZHVFG
5UzRienavaXUyKfnJYkfLxaW6BdCgNDRcicATpOW49pJ2NwUcH0e/quGfLVJjypAEuWFCrM4SExW
Uycby70nOw0bEFW1knDQXe4PZJ8s1ZzJ3wyXP/IIMFUzozvpf/k5trD+pp3AqfT8K2sUPjEgWx0N
G/LJByKJxQyKmq7cG/KZkYJludPc62g+1f0s3GMf9m8mTRdRKLoXVIAF4g0yoJagB6g/l7DCfjVY
N9X50X5C5X1wPj6uM30J7HGT4WpslZGAMTP+gGCzyEBTXTfET0517TUqpOoTBwJUHKNA2+G4OTMl
Erg651bKTv56Lk7JaIf+X5cZPg280VXH4+KjcfY/vLHYRX6QpCkNs+xHWTOX+3yWZIN5kYzDSGJq
BhfSghFY9cWCxa87WZaUfAFzq7EQ7wuiH2T/75MVprersiY0hKJTsnyY+gN05NHzwNGtKM8Bmdhs
a0PMgP+AXzSCTEkYvAuaFCG+wn5me7VTc5+HgWU7VRcrHJtdupSItcoRHFZn2oJvWEXnYD53Bdc3
91OV8wIJPkpOygbJZtbaRDQiHvG2RYAOL5JJvDz89neLutHowyKrHz8Wz4inQw0suzLNUWXL/qkO
BODAEPffoWwni4rPgII7f/M57pT80mk30CYd9r6ni7gr7fcVShC+azY9ckLuDroEnk1pngDwJ3NA
F6lQRI3lgcy1EsTGm+zV8z51008t07FsFGs6fisJeCGYcJCkJY1It6J9VfFymUELc83a2TqsSSTN
Qx7/nM+pgymtWiJ9Iatc+kxVek6bMdrLyL1+kgchtm+6fjdIZHCkxVsqhlx/3Q8YZAEJ24w+Ducd
Hzk4BYWe1qqnVVVX4z17BGQ7FtVneyxvXFCb7LuTdHXhs5D8igxFYPSdyVz663ijnL+ztYX64bxC
g2Dcm4U1RS3H3ITiwAuktbxU8U28FGqBDi6EPD4P4d3MG/w8jRzhN5L7xAMKtphkRXFN6TqVtEFE
+8vpeCDz2mJykFcUrAvUn+p2eL4wUF3HstCoHhBxWzLZXRyR3EGu2AFt2otU+sWEPjEzPIkwZywg
+J47NL7lXQoj9xq08+IeSenanvcdh6t68tB1G5/q4Hk5CjKMZF7RkXYuFicX8K9kaIg9qQlICO2H
ui8tTblO90X7/5EaM3IoQDIcvZMNWVyknANl5bcdUyAD2hJ8budo624N+ABESfzbdZ04ATswDy0o
8CLWXp9x+0XXlXm0bY+vEBiO+a+xPdrV2pI5dq7oGTgDiaUdUOyPi+JkHjfi1S705WV3Nixswciv
BWB9R9Qq2VcsC+v+MOO9qgAJobidAWqpF6Xx7z3yrUNq6AZUXhlZGse9G4nHDkGMnzE6XG+caQSk
sItW0adge34uxWvzBvT2Z0DdXtATPns7BUHPyJ3m8HHXuNrkKLeckI4lZItnpLqEycXBEd5DlLhV
dR07x+WcJSzY2+cOEHwqob9ojWPJFgUfLT1j7MX++8JVS2YbO6B1th35ZJQ1/zhjd6cLkSWucrPp
SjLvqtazmofUDN2/IUQ2sq+JkMrarKqO0qvkB2vVe4oZA3QjIdZyykn8IRxWLgC76PKu+CIjgq4J
wyG7bEQlgS/CXmW7F/PlK+OiWm2lCUJQWv0jZ8b0RQw/aRlGSN28/Gihd4jeiDkqz8FYsPbEFZJE
4aTVQsq/mmE94ilw+kghXduEDUzrqX/ADOaVutyDSopHJaCT4XzZhtGtNoPqae94OLbs8ofPajaU
cRBp/IC7xRNou4+eslH96zGFoO5pby5WfAoxiGQPp82xBLb3tnV+m1IvyT4Bmo0Y6yeB+/x4dwll
r2ywACPKHGni4PhHobpSwnkU+CbXgzLCsVdyDYaVP90mhE9NvLlY5GVqJr+ZwY0R0yp0P7U5NMIx
BFfrwtjQFbaCT4AV+OSU5u6D+LHrtOD2PV0M0dOF86hF2v00glonCyXYqL6UjQ7q7DAEvPw/jCE4
i+wnRD900962Q8PP/Zu6d8MbM6PbHw7Ztp5RDzWyi4kb39X+Fl3KKVccRot4RnEp8sIyWl67Qf8K
euoRQbR9hAhC9ye18m+LT9Pb7ZyswW9xDy8BwphptS9IyFdSZ+Bf+gW7Yiv/1fGmQjgEHVGflnt5
FqLWUv7Y0kGkQ5mHvSfi9C+CAxfEjjdb4y5owGvY53KC9oOQXweJqdBkjxUhCJjgkKiMjQQfWzgi
Hr9H9o6bHhVFwr35l5yNzXRQGjFQJIDT1X8+b98TxIIDwCEt1c9Fx+9ZZiv/V3B8YlAbi/fM23Sz
Onu/CZlnT1h52pcqUk+I8SnUzggA6KmArYE5HYZFJQctWsdhAqCotlh7wjQl34F4d9cTImkboMO2
s8jBj+EuNjgWubC+/TTNclrtuSp83ven05c2Z1aqH1amrje/OzYwsgIXSjYwso+oNOZm7TQ4sK2Y
QsCH0iRxuaPbB1kFwsoy49a4UrkZMitfgpKgqpFSBKRyMmnkcYBIssX5oHJMz32aOObQrAVK01V1
2qqT2jfKpIkMPeMCu0PBQlJuH78PBgY9ZfqjmeNzdwdCdTxoVPPiDtxLJAqscsbo0UbWsv/wnWdn
e/m0NRcMJ6cX5q0XLVxx88dGjYsBBc3hlfSRTk3WG47RwNBFy28kRw4lcMBEiZqPcPcvY9rbKRRY
5hBrV3YQxqz8qb5L8yZ9gyDGCx8cKrQygqBsPwVGxF29xVt8dR1QT0gPxX2AzIQ1YYyJF4QdDqau
fnhOVN4PQDUbW14+UwCAMkLD+x6zcmaJM19I75xjA6Yo1oC0FgqgAVRc5+Qsrq5iLiJU0cbqtGnG
n5AwM62WollB7q9xKty9goa4StSxSkBH6mHaVqxgDbMy3LpBVpW1ydnlRqi0C4WFltFZzdmZy3xQ
QJe89n4DDhCv0W28VSMq38EZeQPjShTdnPmFDVD/kLhx46mUwlFRJDqJHHVMNwBaOLbfBmsaxdbn
kd9JM54dunv9TH7rK7RKd1Y/GliUTZTjfpu816YU9X95WQ0qlDTZTl7QCB5m1BnRPiNAw+H+guVo
R3ZxB3iPQXmT2K0Dju5ce4kHRFq5AFuiL0dxkM30nEL/ofgykoJEag4bUOQEvXPiLaGRxgDr6F/D
DQF+y+Vqr1Jf+2UNdb/MLde2BFnNeCucq7SkB+SkQMN5qMey7sYSUpE0I0+i/6pGaMB6sx1rAym0
/64FGV1oh3YLAqOKVEyFaa9FapKdqqxgD1cdEJnXZS4sqbxtt39G0oauaxEiVQz4wn3ipe0UYlaD
DmXzK3a08rNJ5fiNUtA5iB7zMkm+3FBjrU5LeHWOpqIybGKNGRtAVDZRd9YoaFSBpWsXxY4tz+bu
J271JGLmNYW8xuzI09u2+Riqx/NiV5iQQdcA6atLrT6ahQXzpFC6uIiuPP066QJ7N6oKrbeJ8zhw
js3E8hakh5yVPZ/MZaLNMrGkr35aQgr+vOQGH9zPlHmO+cLmBSgpkxWp8AVPorigaOT9az7yRDif
yuknliybYAHmyuMp33Oa6JcTwsvoZ7fjAulfPSEoyrUsh/6wPesyi3IzndMv4kBs83+lLyIz8anL
iq0DcmgOZSZEg4BV4rRJycodv3BEMpnKKtFYoTzOnUAHFatX/cyMOmTn+FO0XBWbTy64SnPjAa2L
2pNDHpJ6O/621xauZdjSTl1QqWv7cPNkUEjqLwyoanUyG83/KCo5ZdR2dgsVNQC2Bs9lQEIsJUEV
qfSPkJb6q4/kmBLV+fJR9zVbuxh61EYPWRO0pDdJOFhfViwMfCkzzQub0rMqEOdZdb5I6I5MbKnN
fPXYbM3bQ7jwaggtf134H2x7mz7bxCh8RKrMqfvoLTpmfSy2O5UgEq3zTTq9b6bbCeTitV8mciVj
LzYUT4Mq286AzziUgzN6sngBxnNsaYBXEm0Od8vF69uHp7pesRqFPjWzqQqJ85a3oMS9XEZhR3/4
n6xTkFsYU5cZFji7kr/zRSKxMrdiO0sH1OuAgyS4dgUOf8UPVyj3Di60sIfoRyt2O8Lksb9Zzw8p
W6PqvHuXV1GajxZgA7jFshcfBm0kwgNHPttOx0/Sk4C802yHAsh1bKx4k9i+X5G3MvsWNF9rUv2v
vkQxWqg0ZXWpKQ9rD12jjtCA3h/9WaptqhA7n4TszoxnrEZIchwOgbSHYPtewjOKxbcJELSOy5tP
Qbh7hbxyHhimW0ljbIssm9USuhrXiRw7O3dMYF8Ac/HCn/C7b66xjxRzSjxdyq0P6JHDkkAL2LDb
FsqzL6BaN4XDJuPtF7MTc9aQq2LmXiOm1LWHVKSvuhxzlYiU5ub2++NbvKH+XNKLzgys3V7DUmTM
bmLoggcGlt2qYJclUmTNMNg9tovh4bv2DNbLMKOQwf+RamUWNgAyXEt0N+pRdHjGrvCNDJ11E8Ly
lPda0yjqVVr78mfHsOaSlG+Jcwo+x6z2ynFtDp24Ux+q+ETtjWV5dy8UkBt1AMBojsvV5QYt845B
sa1uxUsO6Zm3xBaLB+RacmN0XPVyZP71KWQDBkcaQYpdL8hbGcvN6Xd9RjBkqen3PcuHpt0KAXJY
rM7HnB9+qxfNgvJjUU0X2IfHfrcXP1oMf6CqZXoDNUtwu7cCf4pOCCAkgJ/v5HOvdVdYSgowxa3U
gAFaWxjFdhQwc1JN+HkaGE267VvzbNwZ/plEEfngRLEtUZmOKgZosNNbDa+yW/VcWPPAGOihWXXj
GWvcMmsrfQuz4SBC7w/8bKGVxUP/SdTAYulSgfOmn87QrFl5iPI8OTjXr5NmKifTRcQgsLa6qUSc
HDhYdukhF0GiCS2NxVoIrOECoWlV0nfXN+VSV0cxyOEVQqTkmuyyvjXWyegj7o5Cp5Yj7Kn9kDM6
2ynwnuYztR9rGNYj/62C3N2cNBOPcL2r958grdXpnNfbbWeyk4de7U7rO7srSdVzZjiyjgJubuT8
lc95NEoJ+W/pPqCeLQOX7fAd89SzX8W3OhrFswNwV2sDUWlluALeU7FsqVaU/LYkBTPmLeS1z/Xe
RqTfWuptKJ2+qjRjcDAX2/66nkk3tC46KmJUGhNQLxArflw047jNvNkuUO2wKJuUwbuoe9ZahJOI
DQKylNxMZoenRGZbHEIYUpWHMtvJVn9AOmGW4NNaIXNgAiwftgCHrnnaHfv9hfQ9bILBmbVE0E/d
eU8gKCWiwxm15sRezMOKf2y7IlJHBPe3SZRUEyNVR3nT9KlmNkHqtClrA7YaRoDs0j4vutzi4+ti
va8TfdIznpupF6Bdbh+6Le+hRwWCzdhbMNbXcgtHlwrKxoKIoeOrDBpRS1pja5/6jcz+HZjvoD8I
rVmVkKtIVy/8s2a2WYS+vqs49N2D0NRoqTMjll43qnMAJVaXRLbH+JW7j8WjdkJbBh8FE8httLGp
pghoaMguib/xGrFPpvSjSBmRoMb6Oukt4MFvA3CgTLyycRt+CJ+JHKqfYHShl0/z/NQrne5FJ1hu
xvqbUf6gDQyh+M58BdvM8MIVro8eenyEubdyjse0247/B3/9dX3BBz/YqtXGgHm1CXHNeBdlFxAm
3COqfcZXaiiVWwh/KbMYy0eA0wUtiQEw7b1rYB4sQbpRvrg4lIEtr1uAUNMFd43wE2pdWltAEu4l
PP1FI2U+9fBGs2Suh6700bNEIGzpPm+UU5IzJnQCFwlobxh9FiN5rqX10OLaeF8G8paVSnS0gA/E
1LvAzV5QEpQloXac6W8daRp3bMsVUDVkMcl11fnFz9/iz1NiTQUuhIdiyz1uM4hWmmIR1JZsaQOo
LHBXb2US+3a4o5gvz43nvvX7wm6ndkyMaRQiVu6mF7t3/9tzFYI8mS1yynd/8XHcfRRamSko9wGO
74x85Dg5FGNou/tw3HLN4f2Gwbm248sziY4h/e3W8HZL3HHlKATPNXTjZBWACwrSFUsp+XiAVXBD
YyBMiAmSLfeSoEQbWo2CLFgVhEV9224b3OGUj9AFPx9ohdb0ZwH7YvbmS+eRg5lcdLilKGdoSZgb
VF5Fo9N4pbzvF611rTYH8TV0dj9K57RPHBVRkIcMT5Y341SatOu7hGRARQpI+8bZshuPnsa+1HIU
gRT1S6Yz4JivRkn2ui4ImjbMso+WHwCcWgiKfF458DB3CKlkKeeYoO0ttiGHN0DXButjJLOa+MEf
VvZSYJ2gHj0UF91W6RQzyJIbW/qLKiRBeHIJmkdqt0rmKkQMvQxXUgvdON0ry5PvRFSNGa1HtRvN
pmGVkLJhUWt8VDLB6QjjpXxIf11A/a718vbTAlQstRjvqdKn+2Fa/aMo4kvzmHtTE777HlSh9j03
aexuHeCY5csK0zBdKTBIGftMflHQKr+T/7Ux4ndKNzrDm26wl+aBabGxrZWSb40AajMLio0TA+VX
idkfRlnmd8V3QDbjz9BTIY0YHwgw/kToUbHqU3ZoLO7bcwQq8UfmuvY0QiLQXyScNd5th2aI7PSh
Y06Z4awixfM0AKWaeoloV7sn7Al14QJcRO2YvyA2xx4CApbDugqlo2Ihw+yZZYtSdQXNIosPYBxJ
xGXVb+7bBHhn1qHSkCIHrPFjgVltOM/BIunO6XlnFy0IzdyzfpqEWIwhRlvUZ3mpNqS1iNtZJiBz
/QCQGN+YS939JQxf18G+1Nuf8ZzNhA4GV+PIiOkQmflGXyhmx+YntAiZVGJWBqertxavIpojnPk2
6ZMOqOALI207dEIXftnLlQsT4PFKdhMxLlhY8c7dDHzAYYxOyUiXyC0Iqcvqwe6Mw/jeNr9MfVIH
X20HwA8b83eLPMJKrweBpd37VE9c8bpG//4VIbRc9/l8ehEbXlNS750s9DuK9IUDy9td0yYfxfaO
vc1b2wGWVX8hQ5LGU27W7Dj0VmmLmHdbLcoOykoFPrplZcHro/MP/yTuH0wDi5H2UdGM2ub4VNfZ
oC3L0pFklrdWVFn/WAAz3tyzs8X6t+AUpuu/zfulWjSxl1ZQQ+WQzLm3uuB4pylIp+hueEwoOkJ5
IIgTHcxomtG7p2xvqxZUrIzLW0Sdc8h5ud4MqNHCyA+Os/8wi1oDLKaL6g62IJC1qA2nkVbHsjjI
oeXFjytUG8M9q80s7762E0R5OCqKB4kvKLU+fMFjizZ5197Ysn4kXmbC7IcHWUv6K7+2M9nhioCC
mV5eMM2DFUtO+KnS+IIGGHA+yQ3mzjEMBJW2lpJWOl0nTlcRaEuxCd+txbt0IIr6JoMojAcc5x05
j627nMDSrbBGx7Wj74uCVxKWr0FZNbnLw2FyprXdo5sYrp6wz8kXXw0cQg/RrlxNWGDdmwVzHaTr
MluG8nEUmL7+vin/RmdY2H8xO6WcDYVFIKM7K/fBkpmorfZUBcksxV4SLsanQshVsXMLFuNqn3m8
N1OVJY+DhIDHDjZXN+R0eIVyouy9voSYbXFDYRRtdR7fiRQB7wcEt0uyv7sXju2t/s65NmZeI5ky
LhrnSJuPmz1fkSxglexFvhQlc5n+FGaumMWIFtyJufcLKpYm/wv9//GRDN6ZHxcbhPv3XI0ZyTsF
J/AHrSaLraJf6kDadJEZNV3cuPucGBbAJ8Gu397g1XLNprI95zvo/lytF4B7odNPqb46dZ+zgT43
t2t5/omW70WxTc/bufTNKf2+NNicOmG5zzv8ubUfWIxnit9Fz5FUR9CKlfXHEWXD7aambrYfeflR
fxNQKOJTBWctx09bWHz5+Hiws4J3FHZGzn5VUmk5lbqWeWpcEBJxWDGOpEhl5MmGNDqVIqeAchSY
dSY4JpTCucy5MaD76+U7prcmpN7LCyp7hEOCosXK5eDbJHpR6cTqWdsb9ypL3QeKa7JqKIz/++UA
j0ecyG870sEQ31qnDRu1opjJ6d0j+LO5+A3hne6b7t01k200fDhI8MrCg861hCILjBbnFJ6KaboR
bAJ9HFStH/Xw03GAcGQsljHe4lZUZXxAmN8RNSSaDxuPrILsyOmc0z25WNYSxQavKABqArQs7Sn+
FJswQnNi45L9m39OrOJK28x6SlAeUwboHULfOt1qazI9oJr3WWsaLwtEP43t6OLMbTITBhLQkM8P
HOxSerrC+IrRFA/PjALJ6cKfBe2bz+OPHGSpt4r8hzieBSLGHYSsqRiMO4fePoqw4g+QUXuhukuI
tsfI1pdXuXNuEc4H8hQBhhbS8kYwk5uftYE3xUTn48addXHfY4x2JoB/r9pSoJBT1nx4MHYT2w5z
9Wx+NlQ1ftR0Te/uzaHJd8LLDj+dOokkz+xIJ8Q5s1x1Jvn18J8ICZL7MSIgLiSIfGyotnTj9DU2
Hxcd3AGnIYRtCv1BJCQwj4ii9iyq7Yz3l94Rwpq6G/XffTsqeR6K2EhHfGCXuYgw89PTkpIoCua4
q5VeRK61fTwOqt3W7+Z5XRKPvSRwGHiISJy6S5lDP+8Kbp0PjcCLwuUtpBPrH2oVsXXjnlPomGL4
LQg2HUyp/97mVqpEHAjE5vHn908FcnUDyVJY6f3qfcCr2ID4A7+49JN6PK3U4VqHN/WX7Hone9UK
Rgl+9fAHYoCnt8OjAmz05NJI4uXehIinkJyeo5dr94xf/1hVoJHjQuPutAMSpgd50wetYYx8YyXo
VsHit4DcuTmcPysDdsHC0iANFO0YYfK4KPWIr9INwxQDDZX83+BpUwTv38zgNcdKFAxVbjE+tq4a
UBPgcWELd/dyhXC7porvdxz1mCi6kDUFD+ug7jmkpW8nf3LpS9zvP21SLBa2bXXy009FgEPS+YQH
zVio9OYfP2xMAh859Lvux7gpZEofMPxOy7k5ZU/Qu/Tk469swJGE5xPv/CcLtLXQ0JRClTo4pDai
Z4b7xujWUOSqBGckyjUze9jM8njXF8l4CeFEp7kCIkU0DyK7Dy0nBOFGxP/rMIYEFpGA2zmD2/l9
tbyibjka+DEiRwp/541lPlaS8pfxhjcoJfv4R0T7ZW7x/w3BTmlt4+B/jS4KxenIqrZ3Gxv36WPm
Xt1OxjCjGQkKGOFLHmA1SQ3SLlHBh66dPnLjmehj3AEYr1NvvLssKtdVzH36MVZEbQpS5HGkSlJe
YMM8F2d0qFNrq1JJB7VuuTJXxWBHD0PR/bpPsWJkqrGEBz1+utEeuctmP5Sb5guiNYPS/TOTxZF+
rIDG0EMtch6uFmMryalGt+H5hidOFEvmtViBhxR1jtyzsbrV+jNx3vlBQYRhBiCM/BfY95ScNqFc
NI8poHLX0sLlpoIVJlnIXQqYtN912FojAqpdDs5FpBzOf5bh6JhKqEOIkmLkghvdtvsN2sZCBut5
lI9b2UCAn/LLCSFQEyArXf7zDi8EVMC8AgyAOI4AKYuDnQIJ3v9tY8oHjzfRru8TtcAERFO91Z76
iMNYVJL2+FIu5EorH+5FJEsp2r3rR9opHwdC7JfGe92fo3FVbCLTrpUFFo1DdToY+vzD0gKPpvsU
ZcNHJEs6Dcl6lhPaiCQSJEsuBC4bgGCrc46NUAZBEL65/T80OwOQtC28CVI+fV8aTfgfm0qdlqyG
Nk3ajhOG+QBKK85gbhqozuKEMTIqVZVg3PIc51ni5V10pqy3IbZIjMs7v3aMUDVh1Ao64OzNd26C
dC9l8Z1ZR2/KsjhSZWaPzWh63yB/HcIOV7KV0Xj1Hfzx0Yk7F15tvDItkkHisUF0eAbQA7b0/Bry
sXSHNJBnl97SYqEooR/fURnFBh2r2/BAAnz3CMVGCEzmpo96HaIvzKAQQqLsEU+vN77oj9qmGfZy
ZUyqjzfGTbcxH9QhTrmdZJ+SOlXeC6FFJ/5nglp6v8gbaWGcm2WOPkYal3sZdEtd1BLmM2IsJLPr
+uxgdlPjM37T2gCR//rYNAVrPigzj7kDBH1vsjad0hnoYRa6ne2s5O3MvVpvafaEakMbadeyYZBN
KVXje3BdPHfVILO25YKjya1tvIn/m+yMJgQZlq1FElirjriWWOM1tSsvpEexNRsvy4X+Mk9HL7rS
79edc9JoZesjnPyU+bM5PfS0sFd5wQPYbnu+3H1+VPd5GKfaanAad/YLUBn2moIK5SCN/EB9Bx29
NvBJAmF7nzU4hGLAQH3aQhlOu4QRi3z0h2dIKPBL9w5eeiQNWsTcCV/ogVG4g7vBTHJbitS3dg8k
nMofBgIGOO85e9dcyO5JfF5QZBtChoLmRbUI11+8kW0swa2QckiRsebp/6zS/VWMac4v0CjQRvE/
qDlEq3Pd7CCHAgIn/TUvgrfHFzIkLVqgArdfSbPHjF3zQRmEwsEhHz/ItzrTEEkooKkXp8fc9C+M
tGTS6u8yG4ZK+Mg/4Vyka/3RwrTkac5mHgcZZIjJPpkn662XEqe68nUrXug3QWUGSJqrE2I5YkNf
q3ico962dCtZ046SfgbLrOhzsH+DjEZitv2H+mhb3oyIPnIYwMtWxQD99F8n66PIMIjsek+Lr7B7
Ee7A5JMiu/IwuCBkZmTD76CmMoWSbO2CofTyEwE5dV7y20ElwIIAOmULMJzyk8LqBHjjU45DmRkX
qOT6+xOtGQMrI1yy1EAmi3Sr464gUYpcc+YBjzeQ03RGIFxFtTeBGIVnLWtplbm24/cZO4xDHhHF
b7UcLj09VLZQCOlLN4bD8CMxEtyazk5UrrFXCnw6hO0dnOQqMpU2BMpNaSCngnEKGtQC3zmLH6Ux
+uL8401duLFOE49vEatYqbXuzb3/yl7ENir1lfkfH3Q4k+57QI3jqerHqPoBDFzl5YzDpVQd2QA7
v5KA55kpOZ+DgzWlg411kndSBq6p2UtG9vvppbTR+s/BsxFDO44el6ur+sXMAEoAYSqCVMZPPg0q
osnGQ59Jnc9NCVCSzYZ8LEkQ7fLmW4Ujqtw60SNHK/7aG1/4eGyE4ALRbqWAKuQkRbmVICjweVtm
kMvVY8ekwc+hlgbsFHzNa2l/JgaMyrAo0Dv7LAGuEf+gohT5U79Y1hukUqTb8T7y2wQODjBeY1Fc
nUo7qG4ZaBKnNQ3plG+NQETnKikofWFYKOk6vmGA/8NfaOJ02qssyzF82BotZ7PPgRoYsO6ie8/5
NZMLm64km4oF9VhhkGA0UxJy3SAwt9gW+l/eiHhvWCpExpShwYKdzW1hp1iaR06hhMZL/Ij+SDiD
Sn14E4LudIsJa0c0PJ4aPBRMyi/yGfWAgUaYPZlb6yz2mpYYu36Fhel9HNBzSHUFOmY/pVV6LCOR
QpSjKfLAP15BdctMxahUxXTGDdDegIsUx+SjVWwu4vqaC2HvxPXyYCknK4WS2PCryGj0rbUUo+x1
2pkYafzTpOd9azCsN1L3hW/AVJUWGnsDAORFmKnW0caN/Cpi0xaSyGYNiOQaUYEcf33Ni3lYxqfl
HD+uIpZOMJLMecAbzMDGEuV9/rGwkOVS4PSZ1TYr1EPtY6f334Kw4Ittr/FlXIkCXHIJcW+t18JN
hatZBXMiirWUN1Pqv2F8ruFwLG3CjpPb6mdu9LBHwRLIN/qHT45sjxRY444CpOykpHC7XnyIyKAT
6rDBTTu0MSv5bvATSFxi2b0D9L8pLERCBLzfsl+ufTw+7P5iyEVE/BGGEjNTSdAFiLYSoSe1IdIJ
mv1Mi1vAnnjU9ozjzkXYrGrzu7qY73HAyAsiqrtuj6+aEXs5VagtdP/+nw6lerizuzjSYLzsIYKu
9hCyVidMsvYXcTKYsLZbVeop3X8Q5kWSIzO0ppjkjXyhmRiXVWclZ4bA2zqaEphxp0K/sTVOI9dS
FAKAhpwomHTHf2VvuSnQhLkIMxPh0xbnX2Xj2ub6Xj0TKbT9wcHz6VD4AED24ylw6DLZc2v/biKu
F2Nwa/17Rnyup4NBG2ofv3bH0wdMuThcft5t6Qyn54rW2lBmcxdhvu0BVT2d+H0G4tFu19YXivvn
r9XxF1P6A19x2tmaq3PA2dFz5QLHVXiLIy4I00WA2Hio9xy0SZaYvMxoz31HHQ20Y4ysT8wct20L
o2T52Wypm8yPCCwhpNkIt+UvyjrmKLyRAT8oKMdwiccmDGOdglh+R7cD4AIMHOoQVgvEiiHFmXE6
WeM8kFMoFG6ZMTeSIcAD7L/VwDxyZf8DHht71kQ4YrqGFVh6LFFRDzwLOIoErpmJYg+pBLfqY9lH
b1hVcvo9kDt//4Zj8hRDekaUn//PLDnetuZo7ek/L/jzDYrw8fGPM9oO9E1TaKyNDzQ4tKGjn9y0
Djoz95LQg/KTTlPCMAbIqPIwSlzSIRHOIHwtTVwPvSibqH/F9fDj3l4sWDtRvEEdmIsv5qfDeT3t
ceWSSmZGp2RTEu7kABHy7O8vnYgTN94DAgQeRnfmySV8LxeLTH6t2z1gsLFBeo1EAFO0w9lAObN2
x2hc//+VAb8GxxW4dsz5J8DJLpiOR/R6I4l0cQki0Svbfa78sQAfXrRmjSnYNYPWJvLdGs7UGL/O
B4BnUDpTvEFtN90VYYkq/Qh9DoqGZ4bAlyW/HkYuWdEO/5Ez5N/duoNY/n7f1EV1sE6fOhFqU9Mi
aepUjvjLCzGicjs25dMg5+e4O1+Hd21YAtLCxBTQMxj9Py607tV/WGEAEqj5A7v18xKebbqHPnKh
MkRcdi1GviyDuTVJj9AvksJth9sB8LQgAK9pw85yzT+kE0It1Yllguz0ToRL4iEHgbPx/W5AN2FU
vhwKwJRC0qbk2EnvsscdB99m6Ap/WwtlrSMZr3rdAKOsT6bBL901mDF8VwIUb30MC7W/EXRnbmfk
/N55yrEkUIL0aD4jCcmdd5zY8pgduV/VNy4XumlUQxyIqNoZSmPCkKFmogYXQn2hna2cOZ2HGsMR
1Ql6ScVxv/pIh5byIFC+kQ8/ayiPLyazHD8TyvFt9xSbYfBOkqkjjnZ/U67uyJzHM3Qks9oYLqT/
kgLVoedyOsBTNZtxaRCZhcmglTQ26GnTbHMvagt/YWyEOpzu/yHcU3T04n1il+0cKBLYOZhgYN1W
RV4rGHBSIkafuxYSFeBoQ0tMUJDYwezusjtRrC6P3Gmz0Ru2Si/DQTbaLUHvR6ImAgMBzCDJFuSY
yQp5jtQp+uZCCNOBn8LbsnCWe+1L7DqSoR7U0t1I7JCkwvbSM4xn18IfKosl18WncEE5UtGzFiy3
x2Yksqe6LSZB6cYMKrdcMMfUHbOveVPSsxmqgGZf0jCIxB5DbkKOM3C2XkV0anbkrpo1mrU3kDdO
LQbNekl8qrSZdAxCtBa6LoiJSwUgTtdDWnM6/c5rTu3vJ06TPoTEqbkUrLu7ztXSZAnh+cOI0h30
tS5p4ukAljxKmFMGN93c5FpSZ8SBfff49JZrhwnlFaqWMjWblsnqMU9Wr9ISqOXJGBMcJKEHTB3t
j9RbYxPxidTtV4qaNf3iQ1oq7moeVD0ytDvqW5wSMKKaMblLUq30HN1Da/4Wa2OcxvPmn2c13hGe
+tW8Z+hQooVViRd/KvjirxN7+bOyv6wjV/vG8gQkMjBEgNK6qogBWFvyFZO2p/haebGUvBCBw4fP
2nCyaY6VtPF9SaqjX58N5kQ0MNKBwgXWPz7s1gdCjFgbMiKcIQ+jPQSuzoth86y5Y2iG+Jk2ECOF
b0wz+m3N/HXVPGrwFrCufRiUUjX2bm1tuCIx7zYI5V/gsyhUFDA26SxYZUQXk7uAY+vYuUAMI5sF
axvN7Scd4gzppAbeCTMuqggIjD3/c0NjAmle0HsXkf4cAXn3e83zYJTHDgFNZ5MEv9Bc9Ks7RcTe
zoB2G6JmEnDV0pNY53ShfP+N56KBjHatpdlTAWRuFYVkpwENitVBYz+sxgxLbqxvKI4nNsUVOoW2
bCd1ya/+IhfedkU37kSZKfKlrebr2FgkBY29eKpQPbeiQQNohfifz1l99WNtcD6VucBpdEhMlTo0
p7G5YpPxwxXalP3Cl8Zg7onhXCDLH4wGdUxM/78zuZcGiQRsGZF5NGBKmQbCGj/SL6eW0h0nF7iL
C6FlPwP0jyScdfoDC9g0ZJTyVc/8X7KeSkKj4eKLXLs4gmU9MfeTXWtLiJeEUIe8ehTv3VJwy/qH
ZPVOLKrXrOeGAptEC02ymNDLX76nSHk2cd+rCyvrjymC+g78L86liyQwbogk5viRyDFYeiUpWN+Q
jpDgfb6MtwIQJ2Ks+/pkCdKCj8BsHoRSiGpkNv3TvJOTpZ0fcHi+aNFmkxNKDIHjwv/cYXzB4T7r
GRpXudQMKc6qTLa1tjHLcf02qO11oVg8NHdFajTcbzqMqzAp+HpuA/vxKVzXaBRhZCL79iPrcq5+
r434Xwj1sMn4Ut5bRrE7w33CAvtxk8IDOsjkfa/zZPymGq43q5EbvUFPD4gY9dYEeggJiveYqDkN
3DGoWodrs86pxUdjuu8fz29EteIGjuLqQLQVh028EQxoO+QNqO89ROEKEOHyRU9AjyO+YTja0GOi
9+GUOlLRE36zV8od3zbruTXhpkoooM+iPozNwYZwF/opHtU/hESqWi5ztEd/5++t0gCynn95PNsM
NuYw1FthedVMlVl0XxXBdDf2Kz6ibYCJG1ZHm/5qqKTrfmthvudGbYAxWFWEAIxwEYvOUZkwosl8
m87a5ZLk/VBANLTHERTvVHgT7bzHyLv+LEkTrTQOIbmSU7hF9NnKWT/Yq1t23GfbpTBKeUZ+hBqu
b14frgRQIb/7hvH0PT9lDbmnN3VSfnItfWzVAfCv7cS7NkCB+9kLLhmfuByX882MEXLBAajygTmD
S6twlOxLR01OnaHfjW/r8b65KO2v/xmsJ39xaf3DlwfCHOV/NPhQ5yADcTFxcodzjIsHLG0UN9FG
iBGvjnBcIQ0tPA8LUCrmedcWTBIpucgnn9CYnrN3C8LaIpMrBsrw2QQ+czRL8us9VOEe3RalXEe4
XmbhfRxfQ5qOZTLOj539GgDCTHl0aqnIfFOXPQePED5j11KTU2NinWRqds+1Z6H0gUg0mK+a75og
0Agtmiy9x/atV4qrtyq9h2qMYDcWNjkj6NM289e4FFhD1vW9cOsMRHf9T/5xl1Yi77RGGE13o1f1
Ss0hHadp5tAhc4pJD0RRfXU6NyxJ7j6MYvJAtqrTAVPBkF6ScPN11/jAVKV47ox7yjUE2sAE40FS
0VM2RQPRo+ja4QSqKFFD7L0G64q5vScO/7afHFcRWJilUfe1TUR33zAEXRboCsmfSPnEE/sAQqaK
hY06/QNzIoRDQJC+NPxAIYywqTBJUp1bQvtqID+o6oXkyqBKg1J8ucMvdM0EgGOvOVSICUmJs9rl
7Ld7Bv7N4xraMKiKsKILebidsJdI6Lt3NYuxkkPNFL7WY1Gn++ISjVtTMUftLBMOkK4zWoNU8IZX
RBc5DqVApLuigzB2u9TZhnmkkqJDIae3nWXvZGMj73YUTyUeURqkf3P+FcoACqhlZKMpjoQwNTJ7
1oMERb/d2GZqehhxCexlY0zMODmqLky6Rc4QY4M4jN2mlViW+chpWBDkOkcCW2QuPaD4yLf1mIGl
6tQItiUQ7RLPlDLIIm4glXau8lEIulmoMYviMulqvmMIq40KuwhcxL/lYQNtoxWgyL+R8mcH8zvO
2LJ69X5ZI6afejNXadqTWxT2aHOBTLWBq/deTWhU5TBAu+veDtTc4SkG2DyllGvEymeuqDBPX7Ii
8HpO98EPtV2EgVGfP3feOQ8oPLQRv1JLYr2S4k6p61KtMlQNrXoupoNVwxmW7Obz06QlDS//S9TG
mWCm2aUhzLiduiiMdGftiAHhRDLOitgX+V9frM+xHQWrHBD8eOW3f9h7hv9kplMep5FTnZuLiBKd
cA+ShyrAXCsDFM4nGOgHPWW6zBkuJvxyfYYT3u+T0azbqK+fYZBWxD9uMPOskuA9aSg8qtT4eEoq
j50koCxD7c6e5YQa8qMQG765BGYQ7AH+SxZUHDKYg+PpFzi3+lrq2WIyblbPbck2IRv2DnaD42lF
WkNmjlsEISmAYvorBkAqD1CkKcPaGYX8xr0O+2RrcL/2Bb0aTi7co+EnRkMk5rWWWnVxRXt+jerF
LaxmUGjs746ws1ZmD51ek0OKSbeJbqcIKSYGEQwuUn3zaESfeiUR8PdOQcdBTMUejNOS4dGQ/O+j
pB49yWQtEQyqCXHZPdu8mVOhUynHNuQVyFQBjwwqDQEDTXjxu6Jyk2GRvjI5sneazLAvgMhvBh3C
vqku09kt9Yv3sBJ+ETTf3fwYygZtjyX55jAsUZ03B3KOBnwvPQFmaxad73MU0XMz7qbh0uMwj4dG
uySlVcalDCMDgjbU+8J33FhZHgu9deGwxitlinMzEH/BZ63581pUlYmIyRZp5wCf3weHL6eR0aU2
yR+x924z1MBd+0NmSeTLG/EiT1t/As9ByyIGekqSyb5n2/DIPVy+HxkirnHUncbWH0iAkigbdC8Z
QButthxv8SUH9ZFjGFO5msXYc1DQVwDyAlYPOnC0xcqoEWcNg37nTNXbaV42LwCeR4S+8O9KKgCY
D5kKCQdPsUojDDEU9VIYFU7Is7l0Gy0oe2v/YHX1iagRevIl69PCIka9jdfCGPISJFCf8Ueq0mQd
kMFh7owokes0+IIcE2zKLdQBEIyc74R1jgMc6fBBtxBYFjeNNTGEKm4pj/MgSdchqhgg4OD+l3m3
ZxbIPdRuRetGPiZvxeLRe1xLI+d6Nb1l9QJjBhAu+Yx01s1HIpcNR33azVTyUk3VXSyG/5xKhv77
j5VdnicSUOg40MpvDC8awmauStiIJEel4OkFzuNnB9kKekHndyGKC0lbfvOOmIsN2C/m0kcT51lL
eo7wKGW4oxBAhZ/UWtp6wkYMfVOmMJDudU6cTZ74cmixEEU+rHLirdBQfWVqzKdwHTFZ7f33O4i8
VTdmm9TEm0/S7/zt9FwkGVS1OTCp/x01oVXDT2wZ3t9Z9+SUOnWUgoxa+I5190bGpYpqON5s0DQR
fIEwyuRI9IcwBwh+G+IPZVWj8TgwtQqwTqynKXVwsqQ5Oofcz8VuF5lLsaXIxFjJNkGEAGY45tI8
NZknq10GctXPwE70DFI+jIf6XZiwX1bWuvZk5uZtyyN2MJa46ECDO1U/ZpLcXvwT16qZiT4rNGxh
GOYhyjMszM0JVnVFlYz03wWtL7llFmSvGw7Hxl7b9htpUXkmYYJBaErM2L4iRtn2vlZXL34TaGyh
xBWWaKNMS98Bhc8+ZDYYwikOHwNZfvslyqHEHnXQeSTjHv+KYmZ3yz1BMiJxmn/bNAsOXt61mo06
uQjw79chP5SkG4deZS8+6drzNiQveSvcVMPS/FvlZuL1oToE0mvFqqI/NpuSry2ZQTiWUnjAEZNl
5+X3WrHQO1hjXyx0w0Wm36qkK/IUw8DZtQCLCcXy3S8pxckWVruNGifo90t2YKxAd8RjQC/bpkS0
qOxfhB7ExNoN3BcQxbJSVTLA+oLvvHS9IHwqZBGjc5xaav3CiqdqVAOtBKI3F4hQ4eqUFkzmh33U
UOw9N/PWBF02E6yPkBS9oYShXPQh7pCf859lIxXVnrqg5Dh3yBivZw3VJ88Ran9aBSXO+cqSOxgW
98vgzjyyOCfBdu8YGE+bp4p2u8jXNOCcW0idZ60YgFulwukyyK8dv1/J1J9Y8L6Y5k5M2rI/btkA
+Ir/WRihknHw5SS2Q7S7iE3fQqIqyB1mm1VFjUvV0WGJegQKWgJrdQGC8OfXDiJVWOTLzwtPBRNl
od1bvCiwa2gPg++QRA+rpPN/RvLvw6gJPUfTqIr9kZGn8ePfk6a5s4DWTw39uxdaV0ljB5XRy6pM
m5wbL8O2OaF8hBme1AnvAfR/KG9tm8ozi8r1B1/x2cTC/P6l6f5DTKAIsACWr94FnbQhKtag+x0r
03XXlyitDOndWsF4Jx97CjU87sJ7fStXTsr7vFDrXyiyGWO5lyPyKtXUKHDvmevTklAewLDWoZUV
wSygZHEDkgMYiSP5dqLm3FPkyZ4ZltUJvRfG0EOUn677+++ZH4ZY7rz/ILOljzHcxlGtcuhauLVK
h157NOXHfuzyKl2kfa3jbNL9HQxz6C4+QeVi0xNXRBuNP9U18BTQ8bSdNLQMs+JOWKwkS1J6hoy+
px2NiTWcqDeeDYFut79+LEklQVH7FoZlsSW0i/1gBVNXI9nhlmxv/NaGUEguLGsDhsJboUyi2zUD
MCfmm8NWOffO9JPA0WbLr6HvL4lKxyrttrdFMa0+c6L2PEeS/VW7FhY8yXIMPPcu0k74kAiSBkWO
2qois4EKMB7RGXk0l9P709iRiZ/zdIoGRbBckIXB+20yA29dH9AhP2Ie5uwVmTnoDTyg194o1d60
GNyMJpM7+UmMtuqt/dYThZoiR0ZiOd7AzVsc2Mds0yoGgJyircLhsOEDl5a9bFs4NvY8dYSOIcPp
CdKimH2h71U7+xBMH6VrlG2E7CHH3ArbYsoJvUF6U4sV0JbjHCmR1JyXrMfjxnzchMNwnR/1t3Oe
q+dF/y+jDO1wYRX0sDN3Frw0gIKbfXIfDLZCmWBOrnH1GoCHkUh6ENbq4MPTS1VLoeKJqIVR3yLg
gBOzzXwXAin4AQBv+gig7MgiZBglCrjdwQVsVXhflU+ECtyV/s6kPwHT7eSZBjgHvpn5RbYtavew
bI1gFFOISMmPgLQ3FvXdKe+l/k2/n93aSeg/vPuYShqU6sGzgWxmvHWlUxevEnx8ZX/k7pZtvwVu
GbTIPJJtjuPasg0lIEig2Pk2Yn508nX4zsOMnwOsINTi5WxmFyr9p+2Nlu8DPhnjVQUdK9Rnimww
LHxzHzt82eGgbX75cgsWOB+vzryWhPVqZDAQ9KI68pdx6lcz0GJzmNFcvwklA8xDgTmWfUxzlhYs
kaArP5b6gHXXLZDpQyNz3Cuunr4/X52PVU5Kk277OSoLfMujXZ6ZD5C70caW3THoGLBbQaegMnlF
NiO+K3tjy7EDvoAF2OeGCbwx1fJ5ihnwXby6zhe9thDOIenymYdi09HXIYxM3DyvOA/vGWPLGmVO
RJJnIxU1ij+XQ8WFStppdhBe3lkXXs866LzodFvN2UfoGQeW97F9Ilrb30XiwAZj2v3tSbOIVITW
mkW5Gh35On5gqKtLmaZsdDyI7Yt5/TrDkf+aG9zBkgPgxIbQEQosBsXveF1ziAH+AZP2jTnb/NV7
vP0WMFGSs+BXfRmtlspOeBI8bGHj/jAdmfWf5sc0sqUfUI8vh7HXi7CRHGoMWQmISPUo7Yc0vfmC
ymnZPLzlGd3WFDbj2moQzp5G76g742U0ptpzE3JboA3nLHfU9D6EiLnfZKhsmMriewykvyn4js26
9WMf2uNkNVDCWfFxTb15tx+jTugjBijlKZq4FUmxlJr0JsHK+Bb/UJP7QAmcPY6K1R/ft+bWF9ZZ
Zm5BpfAv0l3kw+aLSjbI8DKEpatLuzZX9svNKBrip1v1EyO1rTxSpNNhePm6zVyKD2PtuS0+ccU+
FlJFobbMhihZfOamXOlmhnrYcNI9jkZgcriAPtBoFG2x7dfhCMzV3oDuvYSSyqWuEAn/wOr//7ND
yxtbpDKoH/UAHY0EGtXuA8iIcQACmF22RV7+xnaOfQzJ4eSMDjBVFRoiz1bvMZz9xwKZdypIzMdW
+ExdBdNivx5eaHUL+Z7j/E5zt7mpVESVCRlV3APgjgKjpGgL7T7ZcChG3zYSTkp27M1E7G3f7a+k
Scil7GH4LbpWf56OUjD5LVs1fsTUow/xzPXLYHSGIy85YPHg3taVKs1V8+ObwutrpPWdcmEw90tG
NSfNk8+z8UixghGvrmBXDO5/rb9Td5IGAYR4hzNYI76/brkjHS//5m5MslOOFCKcGV/xO6rjTa7V
gzxXcxJzP6FJKpH5R8bCyxLub/uB+qq0+STAPJj8GaM/NSep5CR0Fof4/jbHTUOhWJ9OqRsRiw3f
gVQ/70SIfJhgw8WPAKKkrpBesaw0BUSe3YYNekMO7uiPdsIegTUC+RAdlX/xSI5iUm2RzGnXDaJp
3sNS/sflyviPYGYVsy09VD3Ri+kiI148wr5avSf5s+nSE3Qw+96DvG7wxOzYh14xCdwZEOVYo2Pn
+2Ia8wUUEhkaWVBwlDicHv4BcIEIvZNVVbSiOAlEAf1rcLazc9rkst+vNAGynDa1QcsFbcF6+RWG
Fb0ZDcdNITNOBG3yOxQTkVax9b35Dkz+xyN6LA/P3qhIJY9oNsrXqSJebpP5GuQAx8M+5focNMVv
GtSIDq93nKfwloHHn16mh1fGzifzSLNFwlETLqGzAUMJLFv2g6VV3Iqmt+7imHINzsLHIG1kmUnv
F67gnHVy1QitEYjVJLMvER9NpsgQ788coQT8XkEe0kaMwtzQbPz+nRFOEv3oze5XMqYQTPeDlBNk
l7JmwkM6zgF8Q2LbiVnzapHWCNY72yAfcSKzA1GmHcryNcSsL5U1ke78fFN/0coVV1WSvI0pDjZc
ifWZOu71TSguvZC3iLFBYdBpdkv+bdLTAsvLYc0j674HLlsV4zYaTi8hzu2/HdLVF4qnGtMfxn8B
f2XyG+EAeS2svMgWIXJyyo0yoDvOc2Gv0DTReu4vuD0U0u0DfNy20lqWCBxnfuLfJtcmWT5fo3fk
x0VMAi0/mtxT3/8S13CvwDAwGj4LPU+V7j8NeTEDDpFJfeMGT8lgGpuUW2pxgzXXBbNgkVy2Rfrc
ibQqqVlM1U0bmYiL5/PZgEZKTCfZ9hONnzB5zy8W/VvHHskE1Dv6JrXnuC839oGwqbNqNLYBaHYr
TkwCyQw1rSyO8d9DSNJixC6X6WnJgdMQqPB0l/lfMknGrlB1Ie7IjUN8275fsBETot/mLsmMfvXr
h5wRbbqrdXgEu0N7ak4AePYjUo6jaFUMoWwlg0lzUfp+P2rd4c3XbFho0oISgEZHiqu3Y/4IwfwL
/jTB/Qu7BDrqwbvMG8CiGl+UkgTHRslr2cbbyq0r2qUmZr5CgDRQDmqqiwavFsFaXOTEyoFgBYnC
r6PA/Zq4Iu69OFEom63Q2ucQOCUMGTryO/YwnF+iCfZkhSl9SDs170yNDG6iU7V6HI4SsjZlQo7X
y57vc+QMSoCeI/earBZWVWT4x/OFZb5Zk988dJb4XRNmVjVVxPtFHrb/JcyDcWHXnVCqd7VqkEXa
Dvr8z4gt/4A7pJse+fESINCubdUnrXLkD4rtxRL7lodSZ90eIJTPt8uldPe+f89tU2DUjQ1JEdgU
coaQqlOLj0i5nQkpaYIb47zLcAik6hU9ZXRQizHeUXnJEefU8iw9Oxm/Q3O1X5RyrAmV4PVTzPoW
PfW5n9V72CU7ccFkqphEBdRw5oI0GPa8Pe6+zIhdKUskSyGDK9sfgClE2eE+wDnJJqNTu1M7dDjv
qbhuDkE3y5+izZw7R2ObqPi6UQykxQbayvWUhVDJNeksCBa8nFDkvie9zWEcw6rZTwJ/0XDsGTiB
JuwkcQUYEwzl1JOhZI9bApgccJIpXMQc575TuSoC40yOKoVJSk0gFm6uCgufKS8xklyqVZ1MBREg
Gh7cj6Pmxc4E32ftOS2lvKLUeOV+nFds8sKaJVLsjSymXKCeiG+y+VTx05TuRqeVDFekXKj4QSAP
7zmXGKkHtZvkrANrRbtAoVQ4uZlC/xwEbHYe+ZMkQkBK14Xc45LRsstMXZxHiHzpPATdPC4Jxh2a
VjLy4MO9stYHwa6/unE4gT94m7F8Pi6przEfzAqGgRpGnYh6d8kp/zbOPg4J0Ts5PFbvf1kEa9pw
8E1/Wme2ZVB+dRfoU+g9OjV64EeYqBD1J+y6mWVfS5slw+eSy9KCf4ecrJz8tCFnaEwb8Rw/jJTe
J1sZTqyu0gFqrh03eZDup4yb1r+A9+XMzXGol8wgvZpevCHSxernfFZGcuc2eKawAG4hyXHjP/6J
SV9YK1gH2/+27ZrXQ2AzmL/vJSxnG8mByAv9t29P+avfMamqPFbSo+qttnVD3KaI7x8jUm8alhiI
mWDh+IberXo1qHyCDdE2LrE4kFRkbEIokFmvgIxbeO/rWihJcX7zMhrT1NmueD556jwX2Du7HGlg
9b0HTKSCl/2v8Vviuq1SSFFFIPTygy7LUtj6bMhOhJblGwx3xTHrBUzRa7WhEs38U5d5guOJkv6H
q7QTj2Kqd38qbYtRdD+vo9Dd2LygfRlKzO/niiLpYvqTx45uTB7wivNTKsxS1RuEE2jRbziuI8IR
qwvSZI0scsSM3KzKUxcXAybuL6GRzf4TelxddEyerXWkLflgh2Wx+SGkuqpem2O/Yj2sFZ7qqK0T
hZdRzlHKKkKLWuL4ZUx7Vf1G9mOUv5HO9ZbBrjin3NcYxsKROfketYF9MNvR3hk2YOtFa97ewDPw
m7n8PxvTtKxMQMnwr/Ql43nV5oC0AkRyR1/M4AjjuXrldCg+Arr9keVzfjNQvSYVDghX6K3ZwSBK
YzqAi+fTyEN56BLbbIkU8T+flIx3ZMH0ePVYfivyZHuis8E7cHyEPinX8ux5Or7dqmJ12pr2JQ1e
28rc4jejooRK2bDFAhoVv8syZt8cnuLarA+pLi5yEV8MWpUCeSpL+fdj0x4f0Zl9sqk9saNeLcK1
IdiJn6nbgHkWMTWAJ32RCyep3Y9ruJY+yQAB7Df8eYsVcNIjxdW/MBS4YgQ0Xbg8cHYq2dBTuWXM
M/qh4YAZE5QqA8CqtQguzUuDe9DKQrUei27ZKt9d9l0PCeBZEIVBbWt3uZ1GOeEmuYPHmbGtjxOd
nDCfN42saiJjnRJoU2aDeIROr19xLqhSEYSqwL+cJ9KozJv/WoslUZ4zJ1XcNSnrC0s+Xs7+ch2a
aKDYXtRau54JhMyWPS2RZixaUXwEdejlMS4OXX0OcWzHXy1G65hh4/Wt8FFoxySCTKF6Mn9cj0ff
2Sc7V/X7Qn00czdkttzdJZfn04wXhhqCUE9UC9xXanba0o1fF5SE1xDJaU5CECq+RMfFwO0WXTnN
dPNMCEKWuqHe3bE+iD4Mathx8X8chBpQyrsWL/2xrp+0Eqe1tMxwGm4do+S7NT8RCG9njaXawh0Y
Yo7WRWEiOVyP96rdhDg7T6iXHeHdRMGNOWdlXJsoe2fb+cLdLf1i2CsicKgmjSDJRZIuTmIwQtwf
FV9VOLjUUQbMwqOX/lDNBNdK9Dk0w9D+jXAEKGBKlrIazUYllx1fIHNcfKTBTdJxyOkxH0eY+M03
TBKScqQQL72QHZe65+QIdTR6sHVj5YAoPkNadrPiwjW67tuAd29ozHV46nISC6297xHv3kxjGgMy
Fz/DTzbld1sYKlF6N+rboY4F1L23ZLM+OxNmj3A7KRVR4zvlXWmJDeq1rJWNxFDBsCcEPVMrB1gy
ZtTGadnZihTv6UdEQyfWomRHE85tqu+f/aK9Y75LqEgnMDoVrUH+2ppUgQcZUqkCTSyL28jSWQnK
K2D33x4ssq0ax/2TaGsS0G4twIdugybVkWN+kbdIwGTIyDKvmxQ5z9iOKVv8NWWr/H+6m311Me3r
6t+38HFulwL9Yx7oFQdhlTHdMcfpcfD829YfqtllJ7+cKFiKbtk3w88xi+ykz6Y0YK3nrlXgKP74
tR1iwkHSK7+nxwkLw+SB5t+yda4lhusp96ye4s/tudM4IeX260aL5k605q132GiioASGP9qSSMOf
stGg2Yc3x2HsKuM5BkcsMJx0+Lwl2SPt7q30CBt5hZr1uwIzA18Z21xbq2j2wxmOvKSVeucpoqh8
e2hhC8pqXUyUyXHAtZcUz5alwaXW92zLgk6nrpSpoVeNq/ST48l61qP+EvtWlI13U3Ni/QuOrwZ7
2LSBO6uo6lKPCkpExV0mwYzXQcyiOPosKSVpRDxEo43QV0/ET6xt4YNExlWge+ghoY42VKZ10b18
jPqfee34GW/z/n+BE7PfyNyCrDWq9AssuHN0J2AeY274774HmnNUtdfBJsL0ukmLusRWbo1QxUBY
vIT+J06foKgT9wAuEhpQYARCeZdP4wE2IN1cEtRFxouch0WkXQg9Jz6j5OocNoMLdynPzJbHsZi8
J/DzylD7YFvN6EruNdEy4R9BsEPFBMFJe/WSqeuQPBdHMQqG8RbzaADV/wYpfu2h7y3HSgpDtN1/
xz24MNAskE2bF817nvNFI8f30FsAqbfYh2eRQ5KZ7UWhqkn8CInO3ELWnqtynrUZZQpAu8mk+At+
aFNsdOz/TgtpKJGrkqvieu8ZS04RTu1BbkkzWLchSg0BrqRzl0awIASTbiGIzcuuAHQLw9flzL/k
VgOGpUCuGM1mmKEcQ4v4vimERStIvhrGrYKwtv9mg/5aP/qjhkgOaTrXhfoUdbnerZPvuRbgAxYk
ya0U7aaU3Kh/LQY+VLa3BCSb+p41PnLGXRdAunUIPqFX8mLseduCyD/wN1rG2/tQMCPQCtOaSb++
GCF8n5UyKF1j++E7IhSt6pY+AjqenD8jToQjOkC2KDbuKZnWQLurgZeYQI92IGbGFbd0+ztcGIdF
BO3o7XidQLYPPeFUaWhapjYO9UzDkLrlPGnV01pEpZ24AilwBt1J8ynj5CQ0MQ7jkGb8rq9IMEmz
Wb1L+uh9HOoGtkZQJveCTX5JOtCR4dpWQsTb0P0U7cDTcBQKXon8sTC+9rguk3am93xuyvsI4Mcq
Tgi66zJpWUvTnFysSYbhbJWY+VTroTJtl/KBjExjsMGqvuHHW/EIAAxzhMDPMtlFCcqmgRCoVv6n
3DFqC/VjkRrZsp6oCEUH6i1SMHUC8nkxA8yBZEdFXEamu61FsmKLEsK1kJ408SDeuGdcnDbt+Ff8
KgAmWqCuMQRQN9MlkVecxn+SyhQ3Z0V0uZplSGiTDO43UfYRrjZ2oU864NnZ5jSgKp53bQw2bVL0
6L/1fHWnakjCCrn4fr0w6RxWkA3LMlq/8e3h1hzabALayUtxphYfjJrnvF/9iI3VcbL3Z+KKGLtR
vegobeVr3anq0k163gJfKWtNp4vMH3GwBda+cwGLyxOWGTtyfor1HDKcPAqxuUmlkm7Q69TS2Muu
QvcwgjA8mquRGV8HX/3ZLOep0ABQ3w7bwbG33+6ekm+x1Ui656PNqjYmKYC5ZJCfICyMpic5iLr/
AwpgSUNoFgJI9QargiuAXlsPQfEEFQyPQS8V6xTRPtenEvQEWb45uwnY4J6zZrC9p5wXle4HhDmW
gPZCK/cR8b5EzDQUL9vpWOfOFVzrtn1QOfTtrbNMwRw0x3dFkZ7DE0y/93V7zw2Qg3uj+cXUVgQ5
w5/BGiAx1PjAArcI6xXtHFbi9loHvnga8Hx6etns9DBtI/v/17lQCqlpGiu7sGywpReUpc3xZ1Zl
2Shm41Im91hHFH7aZsH5Q2bm1oeVYN6B6PoO8AWiGY10Fo4BtLVSWaVWOGQ9VVVkHAMQmcBtKJOt
ZgqGnoIzUkhNFBILiXhhetrJuCBJORyyQZdqfFjd1SwMVE0pW8Hv4P77ZSTHKlskJx16g7cbS8qq
rlvLxjQe++liWnK2yjpdshg31wMS79fC6S3s94HSE4f/8y+vXjTAubfY1IaITWjR1+knsq43zF4l
eXb+S+r6oO++c5tknc2a6vVAi37JzdAqvCSmIhpAR7z5W+GipPfiEeBsao8e2vFGVEiZAP1BZ7ug
Of3PW+d1BCVY2hy6Z5trgdUwhS4HPGFH8UTrigOWejdoD85/ZtPRWAajMOrLMiii5pk/qIbYuWqR
Gx2x6Lmhpij678rOQcOnSEa6w241e8XFztCPCQCAWCdzxUhGtOiG4PLM+pJv1BJSKLu3EvyXGfOX
Pc0pDcgHNbSYo9gRdtqzicaAO0GXLAGUSbnuSmFz29gqpXaPjqA2jikOo1YNJXPpwNe43OfAhH/H
Z3qkOeuMEASCPe0eWJaYidlR1VI39RtxVvSW22kIOF49y0am9OMhMQF3CuYClvUj7jYM/iXAv36o
VfEfOo0wGtKk/G6bSQxbqYjrsQDmkjEot9/1CCX8LmgnI86X+G97V7nU8Kl1HMm/S2tJ8YMzCVH6
Kn/MbHkCgIzq1sESPqXPlCGOeN9qRbjTR2wpe6ogVaMMLTr4yPRAoAJyzpTcodFbBRPctNPqSyX6
p8OorTnNZCfFyRSwNoOp6XtuQLO/30XCgzcv9baoOpMMuwMSne4caYh2FdIvUpRrY+rpKgWW7g9h
OBK/uxKo5ipilqT9U5STf5zalt7BGwW+XrOQtpbHrR5WN+JxAqeO5OFoO98KnN3P7M/gQ/YfbcHY
sZVyeSpW3FCOOvKpo6AzEBcBngi57RFdpD7PzmrDo8msnW74LCAhSGnAFq1/6g6n7uQmKZtU47F5
HSkcR82DIUwkUMn4bL02Whc2E0rErRIFXjG3TbVa6NNo3T/MxWT3F6yPRBpjWotJKijuN5Laj5ga
ndj+jWw9e/zU6+RerEddXLc7kvGaV/3ZuwfplQGGJbZqQP924B2zSTMnT7YDjYcAxTh+/4PdqVTv
jsD66yZFEasB5fwMNl/6Qc7rKaosEgddpNSyudlod8RpIxTRGSblVN57wAyA89Kce/vTdKfHTwqn
Cl2dMt3MfomaeOiIG5UxmJbIMmbFkTRgx1QhtjR9cRCB1j3HRJ8RLSrEs5W5grfydKCV9Dap3cVv
7dK4D7SU2/2xDQ3QnJhWTbqr+bZrNgPOevGbo2L7J7ybHIdhDh21qON2pMkAzMnheTWtr1qXNEvh
mRj1O1Snye0P10TAU1K8gDL1OCGPj1U/Wa6XC/Js2GRI9w/r3D3kmOhtJ5y+eiMIPp1oRDRLCElG
WQavJ7tZXmGh0PnJPycdWidZbS+RcbwiWx01kfH7hikXxqwsdDSeKiUYBNPnnyHURMZhB8LMT4Fd
Qg87TzlYKA6XpRBU1iJJo+RKkiZ/KwaV2H17pR36t/uuEml2gEuN/8yOyNqPjuEJTAQl9ss6gIdX
6+2ZwMTWyu9q3N4d6QM3RsB/LDiKIF97Qt1j8pn2ZuQw0Bio5Gdknyk8wVflLa/0BRuparSJa21V
Agm+4JpgKzjW6McnzmdAuocTfEUDB0XXa9+DhO2FY7Md3Vu8TxwmXL+C+MGFgRcekOi/4UDzACDL
mjmai/euBYERbxBuacqQQOe00NOMbeM47kcIvYqneBHkN2enPb4S7UAzEkpyrMq2jB1vze6oExHP
lENNblYRDzo+3C2e0fXQGfHh1VBd9NJdKbM+n2Ku3/WJ2b7PIL6Ckz9ljqe5Yht62JsHQ9lt85rd
3xfNusMZKahI8Q+P3wD36TIDTYD9dTZkGCwQzxHm4UXEzg97eX8DIWKUm/GZRr+4nYTMrf3/sEU9
m1yBIkDS121RLzfeDC0Sp5qZ4C8FRngiekN1BnN/6FFu8RbBDG+43kdFF8cR7WUS5Bp0p1R2/JnT
KcYxNBEPxcUyZpqNqK4n1zlbd+18FRqxVeA4EcSQMi8oWbXGOCnOFG6hITPUthOJ4zqH7vfcUpPP
cbm322+Unb6L9RGTBjBM7vK/pj/TJMWoQakGGCat9CVaDlXLdFmV7qk5jibw5q70SZUIxjBhdu/X
eXfonarQkAExHIbt+xcFRUbv2gbPnGeYMbkP2Wxi7ACyfstAbSKtdLlczNVSVD5wC3GxmMh2q1qm
zl77TjHZfFyAFfOSB17BRKmGidXfovrzaeAZoGukwY8v3Luvxl6AhYRQxoFGYkXJa4bHQg+b+pRx
gBlXRgSMNO3BM/E3XS4LsgHvTFO8paVyCkidKCheVnbrGI789bVZ0b2kuZFS2OagZfsaa7W38nqS
EJ8OBQOiSrUaeIsUqJopE04rWvpeaGUolt+VVAnz+G5XJMI7arjBy9EO/fJgxZ7Lub7zTjLwGG+W
bsGzhtUKSpVvd84nh+W6EhsmWhIDVZ24soa/dV+xydtCgMWkCPT8K1DXOo2JBHPoMidYf7R6U8Vs
pLyHS0T3RJk6d/gZ75pE7Pfp00pM+vFlJfp7b2RSde5qn2RfAhCz1KtYeoLDRIgsJy54FwykW+Ad
ULd9C3BTTGLE6gJeBaQjMFQVnPY08aQDv7q6erRADLGdutuDZM9yvpjp4lxm/ApqX8AXSbKBEnth
MNUPJmxNxBoqKGBcRxu7OcEzAPHxm7HHK+eoVjIOzCj0Bb76m6OHp6YWZFuNENIxBeMY9VEl6/OU
XCQ5a2obyog1HasY5+l+VmcJa6jzClbSMBIv7RWWp1lOpt7a173CS9ht87tHlOjyPv1GxDonR9FN
h2sawBOU038SFf13qIjxCAx8uoBsTDoUajs34ORKIPGWA1x+HCyqaPFg9GzpsP44Rzg5uPofcU9L
SBbBndv3R/DMnBKCtIdzOVwRQm5zVKwydZNT09zosJEiOqF6rxtURd2MXq/C8m6AffQPPSRAYDhJ
+FUBMU9wby58L51hp9j/HHCweEezgtQVrnGbesp9lLgYxXsBAxO/C6CbOAKFvB/YV65bAU7oekRY
0FxJP4tYAeb5KV9y6nLdAJQ/DQlRqst36koprM33eiB0Dajqyf3J1jeJ3+9iPfptbLDIhzDwRzzo
WqeOqMcjOmRTmWEyDOB57e+pd4ayXnoqAv8hCVvuPMWDpc4F8WUTJ7ujMoo5bP8u7ajjGp4zp62a
ugYRUW3e7kWAUIdjNrTsnWduDcWszcFydyIpt5JWeozLufZ7eQXigh1KXWQmRWAGQMNm5Rvc9chl
6Sr6JFWXni+7EOF61x7rWVXSqHZSr6COcs3a8WLJazefk2B4H+uo0J64yX/WbtJ+Mq+GAzrTXXI6
7tdKJavk2+630PC65dK008mwjlJGpWK/RK4fH51/CVWXShfKGhVEgTsrZM/c4RU7JYG2pC5QmE/3
bR45M0bR6NnMUoGJINvvdYdCpxuCgfSxSehDtOAArjHIFCTJE6XeLriDehmwMJZMELuLW0k1wMJY
ZjV+L0Ro3HOiuvimfAhd5Gu1AbqqWAGuwcGISoBaX3QhPG8IKt3xT/HmlDZBh9nrc8dFp9UuNH6K
neqWWwdVi0X+XMvkExMEm6tLNbqGi32GirCnJdgeSTima7KrTGUrp8opKtTPZksBOrT/pNK5uXAI
RTUp9uN/uw7+Sw+138+ikoFzwAykrlgCTYQ4Tok2OzgmF2YLVqGmWT4A06MsMsKHXmzl3AAhNFBt
3Ta0DLgmXaIPHMghq6ovyvYsr2yKYWIim7U+5UhUAYJSk7l7LtQMmqJB3QOkhCyiWM0KqQ0zFFEE
nhndsPxiypawE7m+qLb5WuAK75TNB+QRbcvh+da2RR1lNWCbxslxF7yEKgS7dvi2Y9+2jLu9nRWX
X+jMwNGGZ0WdheHGJi2eNLwqXvS121FHq3oqxSRBDgMT+qkUjbYQmRIMdEJ7t+l635ymm4sQGfHH
JHDLFcK7fq/Lyw5gsK7Mcp4TFD6JCq3nOr0PnuN8Cz9pdMiyh7E/fu4MOvRZVu+KLrqRKjoDrNve
EG8jz0TiuOMcGHaF/v1N5k8/ma6Wt7dG6E9YVZWX1pqfG42wQ0TdwVl+bC8VticoAhRugzTXtiva
36UPGXkYz8iZfM+s9EHyDvRgyp3i0F2baDBDXWkD1wPBtzoNssU9Sl6T0mDnRvo/2DKJbRv9I91L
KYQ8yEahqLJq3BxjkjrsC2MoheoT0Rk6QARBhiHgDcjDaRXNP+WtoJ3AcP4+srjbN78etcCWlhOA
SEq3/J2hfMIIuMxFsTjI1R+4leWSGQ1gvwR53ZABolBasf1zf8nB3DexK/9lCOJQOZk+EVGNHCVg
xEoZvzvJqvMBghJCOoy1IAcpa68o8iwEkEuwpeEk5FVsdj6e3Z/3W+B7UUHP26xVaIZjZDWyv3iL
DOegil8qqrnDr2kzZP9LhSod5UKflN1/8/8BZDhfoBX+Fkl1D4JnDx6sS6OA0JH9c2Htj5K8/BQC
dRcI/zN8rRN/DFAuEEayiE4CxKy7fkdcwRpXfw8VvO5r6eCwvRS4g9+uKbOY4tlGs3WnoQGD7Xfl
PqtQ3i632hTXVxz8TDykIDPE6sO6CZb6kbyMBL8HukPFf1ao/TE25A6TeISYPaoaav4hP4AgjA2n
1uM2VC4xNRDiV1Jyh6oh0brNhDdOcvT0gHlIlQHVi4GKXMiWjtR6t9osbURxSbYq8/KjV9hgi7i6
zSlQBqO2Uzyz7r5ChVL7Y6vRt+Xaur95tMlP67rKruICfRpHiSJRQHbF097KCU4MkrStSVgOQI/m
1nftrblIVZPOTbMvEW1qZEV8w07XEi5YdlXn4srzae7xpnRViVxNIteJVHkGUaqYfVh6H6lMYldO
nxo0WHfc7zqEE776hdUTDmLrltDWNBM0BGDhIBnhaCCKw49PYgNTShx2A+5/67QmCdJKKGVipwaD
oFOBEP5geyCwskFGuio4LoRYlE2o/bsszenDIWHUm28Gb2QcgZvdw9TKJvpuc3L1eUxapEl6gp5Z
7xNSTnqtBtLrpNV3kec8G34PTWPUUYWwEqQ4hOoMSobiYlV72FNNTEJo1AQ7qLgediRp44XVxUxG
VWYqTRlH9uIGW6w1d7H4aRH+03PcAQXgDUhEO1GywqEzKspQpKefhKoGHWd8r7m9+4nozXTOso5+
AlvOYZzRQQBzL6fT6ILShCVaQZrZ11M3CTQfOmj6+wPmQKyYm8FePFx3RRx+RtdijMDOvgeoZpSs
rTkvc4AWLkILatqG2cW/4/oD+6aNOjO774feji+PUhWrV8ttgYDC33o/McLfR9EaUJurefkiDkWe
Ky3i88M/qocguKNjRVs9HPiCZYXiGXMSBeoHZTt2lYGqTGvU17Jjnt97tx6TgE4rcVBV5qnjs58C
dnTNacPQb5DBVPtvxwMufYTL6e1JkZvorz9Axm5n2H28J+vC/XCsyI8qD2eA0Ca9mVRcrrGv0Dz1
t0T9a1wFbyUi7BpSdiBmLoC1Ja1jG+hsr7L/z4tNC5f0YEJ9KvgB8t69xba1R3aBO/OG3emEetCq
m+5uJgo1u36/y5coGEhgpqVAQjNwjePSRA3e+9DnjvH6VVY5hznWQjg6O8WOTD1Nd0IsTS+YLcmW
1KcUF/3zDPvBusMtBT9r7RhDY0piGLO7NuLtc1UdNrAp9Jgf+QfzYFg3dBIH5+7+ab+hdZ1yhntT
ds320BSQx6J6v8hkCY/Two9P1BVDx7B08rPAW69YYY+E9VVkBX3Efd9vDfvGZwYyGtPeYDzDRA1E
HdeRjjRtMjfsrcJHT506RLteLpuLpCfmmwGEzOqTQvbMVrhItLAS5MrkHlEPQK3gqvRRTwnxFLgo
MNkN0Z3hDL9C5wX9s2yRlB7Jq8HxYX5CXK9Ot4CSGB+vonMiPY7wBi9BF+8jFk2uE/FYuf8mUCBj
ZgJxfoJ6+Qh58y6Wq3p7XmjHIxzY6SMi2N+9r9Pd76Isbc1mNi7f3bTAQQdnyZs947lYz3N6WwYq
WwbBBc/XFuW/7k8BnseHEVBDK+inSCYFS6e9Qad3XoISK2ayBfE6ZO6appmGBqB0K/W/3oEifgMK
4YiFphjXpJ2s9lVL+boQWBFszt6OL2tCxdpYs0LCHMjjxudgH9P+I09H0LiTgQ/fTuBraWrkkbEt
5QCPQqNPyDdm7Ud7JNguErH+LigXjv+qV1LA2W5gWmd+Yp/Rh76MDFbNWSRU9ey+IIByA4GSegkh
JXFE2lfu5UKDNshRiC6mLX0115eklg6C7/+a3dZTS/dV/qsa8/Bb7KP8QhIA/1l6aKo0B5Xnjk88
IVdkRm9Cn1w+dcgLb0WbBD9ZNla5WnBtgyzjP45LeNj0qpv5I24IXewAl8pScrBjMu3zVzvtnYTr
0/RUauROnhy6qJm0biesXySxQ/SNcIySALqAitYvzi2viG6t7vysDRLt0wiiMz+Vkr12WzWTcFR1
+d+49qViPEwVXzT+fN48tavKcfQcwp2kmJlq4tNfEbkXwdimJoE6OMrMMAdB/m8jMwOb1aRnE6wz
4ygRJIs0bXww5PeloNFu5nxeITshmn13RUg4b9f31pFywjrDC1fKp8/K86AqFKDCnpuIfm8/LBwg
RtQkMP5yqrQ5kKNUk3CiazE1lHi8FkR1RfjlQjZ3lHCPKlnjlxg2/7qlR6ZBJDm1K3YZ8QxywNYH
rKCBgHsU0xEFV3gHnF7AzC5YLo9QsABttcDBxprHqnxZaholBzTW0ssKr9SqymfD33yyoq8OftRl
EpG2dhL7UUWthdmwSxpMt2ktFsWLJQuhP6r/Ccmp/nA8GBGe6/L7eccnOPZJNVWjaT9tRrMc1A0X
Cp74l6/AFLIlE0F5DvLiASq1ly3BD3bYue850d932w3TGL6POgqx0hLL+EKOp+tZ0oXh3ki9Aqaw
GaVeASM/99gqNTdrnLITifUq2S/alm8bWFdzcY1VxbaHFA6oPaG6sOM0qnPmtV6grTmMTuXhRViJ
U8ijzbkzXB1LFEj/D8yZVuPFfoTKykTV9IWw/edFQpjekQZvK9M9ukAKPT6S5D+FkPPkb4HVWC99
DbHg/CpOJFE172zm3AyRIDFP8bVGjO9XqsQ21/dx+Nr6lEVP/fLMpXdpvynssOofdtk28YgyndMv
iP0+huFkoRqMeiYnlIE9SDhEafenUciRiKyedQs7UGTVlC6RXScATk7/ZN69eV7SESV9cI4qbPWp
mLDWtQl5FJaklSON/9fK6sEV5avZAQCxvdluXc18TBQa1rdEBjrQMpDw5gQVd0zuAWklXCyWIsGJ
dPWZAQJMKOoWXO4DuZlfe56v6HqQEbMNnJuSKKBbt2l+9BbYyoL6VEtEohpBL8/bTu4mmCqMHbXV
Upwsz0dtHyNRH6dJubsAKFS+fsfGHLNVp6KOjiJqpRY/WBmTQ+n4zPxb43C6DTtrYX4s8vZGQVQ2
KoXZdRTiYjVFedsUMSxiBTFaBxG3oV8k5mECU39+MgyXTwMN1MD2HCoV7+ZFO7eoUOk7clIXpSJb
IIB+wnVxfuGRQNY/BHf4leuCAiIgdSi11Vmrj8lLa5SPBb5msAQ9tM4DK0HblKsJjd9yR7WRF5P9
qflffXvvaKTFDmp4NUKxMYSMVUnw7EfCUr0pMYs1bM1BlGpk3A+JyhWE/z8KHjagf8gn7J4lQ07y
0ahfUzhrYNT7hr5F5VhLPZoGTlrXxG5jad6A5tbsvNtBTzPEPJxuiT4JhGrDIGZxBN4xH6rxHAVK
EMmJimkfrudWSUt9Aud8A8erCj+2D7YmLGUjpFMMHp12EhLTtMhfClUv4mfvAyjzf9rfOKoi76gm
k74vJ365p8Lx0BCN09A+PhvUgjshdT198YILG06iw+qbRdjEJRYXop8C+KygPaCSwLIxDu+nJzmy
6eoXK0TD8xhPgBGOQ4QrfBiefnfB9Uzh55rs9vPQGE7EJO9AqCu6+sEHXgUPePwvNmd1rtFiS4E7
JC7e3KHvM4YJdLVwZ7Alym/p0bzL9rEg0C7m0wjLjNmcVUOR/drZWF5sMGAumw5VbRXTqQX8sVxf
LuvSu9Rb50nQoqyPGHPBCS2pHitKIUQ5FP8JiyZp7nFLZZBqc+2iVfUMIb+xQ49WLhoOsbBEYs17
xqATBj0ttOo7oLD2fYD03hQC0NCkdI/cEctxiSWFgY0j/WC/K0I6qWn4XbywtVXHeWbWXPI6+23H
/gT26P86PPifnKMY4mKfptIjklwiZFBNHE2xcSaLPKQt3oZaf8QcmAMlQDUMEuF7SKw4GBTIk/O0
YnI9s/bNw/wzUfFnboss85zSYelzVVyYCV4+n14ZSrw1bSzvgPc3Zus8jwZ0Sz+Go1fVGhN+jIle
E5+MEjbw9LhX0SNtUwPzQix3DhxT5lH7obzIsAMRc6xYahwPYeTvFbk4AiEW1dkD+sdti8aipHHp
8zfPVJ73dCKV7qn8ursvna5x1K1aIjJVgUQf211N7vB8VallkK8dbP+byUtY1Z7b8B/kv0awmHmM
gjzXciXagraDJIG0t80gPD0XQi+Irr6mJfRl2AqKx+CgNbSUa5B/N4uNyvaCBuCeo0Hd8wzLUVj+
/1t2oxZy0c9ONsqsV1PKItRcdZ7ZEjD7MmBKIoHLQn94HjLwrq1pU3dItY4OGX+n7NufgPmWj++W
MNxCZlgyaTvDRWgrGBhgR+Y3GymXpC8VZep854ZhXzXMftQZ5mhACT+y3IJ9DehBiZP3n42rZJ/Y
Y5IHo0LPaqAFLfVTlynom8samc6qhnYX3BXPqXTeQOOYaYSCRGv+7v76PDant4ZfKbxWxSDSZD//
kfrztb7/kEoZHmheE8nqXAUy+jrtZtIxvYxqJc9YScr4DNoDHE5wtfJx7mMuF5k9TGpDURyVmrh1
+Iguz01280qdmrxSNjRJhDCJjvBd6fqX3hnogARirxy03TqqD4zhgMP98Y9rx9LXI099xYnrb4Mn
tlmoO6EDpNEL1asAsoNLk9N/gAGJ8TrPcukrPBcF+0wtUuhqkP6tI23E7kOYumwwNEpqmnIZ37OM
5o7ZBQx7P0QsSKRNknGqlqcZtZzsBx0nMVHEOWFpEoH1cJDqDN6PyJS1KTFDn7Lj09n4Fs3VpFE9
WRm1h6vwygP8y+2viRyrJTFIrWvwKekdroMUuiD49sIf0T5hTVvaF75IU8Toqko/6yW11R2uw4fu
GbYDB2fKfGL+9eVwr6ZPI2noi4/wD4pD2myt3yWH7gzUG9WXZl4QkPR1ihzLNJ0QQkV+kgFe3G50
/bhE6wkKrcuXxhp198fPkLpg9WAknko3ZxssAXDEJJWwb09cSI7Vaj4JzkODZOaWVYkmLPNaTifU
wylwrrVVKYz5El/rYKMVVrIGObye+uSZMo4LepgQQxhoCZUV6h5EgynnOCVmkNeEnKeMY+SnZk5H
QCgIYJYd5MtrQl6CgTh069e6gFWRfs4OFV4wvMenGPePEydnEB/bUl2tmH0up16cQQfiBgfd5mLq
agRXNilH+eV4SI+zacSzQ1oTHH1FbCORkKpI/uZOuY+jlu7/qcbf5xF3kNZTkWnm6Sd29G5pZxtR
yUpNw8pkp7feVHphc7V1RpEPNjtLbPmeLpB8hWGGJMsn6F7WjCUCwq+S+Av0x79mHMnxp6vkzxvz
pML64jKNZnBAlVbDavW/qetikFb1Hgg/m61tnh2Q3m4T2kTqPY5gisTdL4kFEBfbqzK+ZtQwUts+
+G0R1EMAUuwIY0TqAyV1tXljctJsM6ltgYorZFKANX1zRCpOFn3h/5S9H38zRpdnvGcjG7A2o8UX
o7YSLinAKoA3gXzOann/0ZeJcmxNmsHe8tPfrvPQ9V2ajKOSXZZGdW38WmNq/EQwE1Z4Vd4D3x8T
Z0RwZ7YM4wiHn1ECu39QC0xJad1vp1ANqxXgABFXK/jlUKKoibHnfOLEPXQneT9do8F3mv6TXVR3
6wEEbIiHTcSl3gjVbWRyG/2o2Yn1u8CC2HPGT8Gb6rkKTmOeXYV4OBJw3dLt5SwFlXENq67y5l/j
Ohrnh0v2prD2gNfbh0cE8klooF8iACFCON3rRg3jPeg1yeH1MFajYDirvBo8K+lFUyEuz2rZTvxY
JZtTezJjREWB405TXCPsObw40u96Fb8HHUKWsNTrailuQLH4q04gqlU3yMFp/+tizT+NsDej0HS7
M7uZbHhVKUguRicyhZ0yWaYpNFV4vSF0H21t8iv0LzRz9g6+0YXqF1PV0TgZC/FstjxFEdMMeYW1
emkLkB+kxINFyjlelpZls2MstEz5X3jGpk0gSmPZLBR1YxpiCcAg98kbW5Dg0Sg0YESaDN8VOpA6
UqbpT0ZuyCmbWBY3lnzfhHoW/JdPXeqh3qd8a/tsSkFpPFTM3iQYylHTVQPBFMvPHrjRPDmqcX8p
sMbo22TxhY2cNqJpRcEhdShYGHVneugxQU/h3dOGWxXg93mmN47LlETa5vGFiREWVgBq7/gDTbum
IpP9/LX+4EEwYlb1olGHeH3Y3tFZCbfgTS5yXTLB+Gj+S3Q8SUao/7QJ6Jb0egmgIORg3JskXUb9
NOYBALEjMu26cIo+2WUo6JhYwnxYhKeNJwnL4W7pgeZZeaH3bii42XlREyrDAgkSsEWnO2voYJgv
vpojXiGddAtgWnmQpdXam/JMsMN/7WZYkO0TFBOyJz/QURh+FqY4f+LTTX6k2PencDMIQi2kgp4G
VpPgOJB4cqJ1MELsvhiT7vpLp3gZ/jKZzoWYkiQLz9x0FtXbOEE/aYvM8LtOPq9L98jN+VYtjfuA
hx5jXM9P5vsH7pz8OIzJYpLMoD7emRz6IT8BDgMzyQqYg3Px3kpo6j9APtQVoc2m9nA3+JI+6G8z
kd6E9VMQQGmpYofaLOFAhFCQ7PoelS30Z0p27f36cGDOzlIjGY1Cy18a4oq+tTKTpatmL7KAFpVk
OwHdq2pDF7njAfhXkmV/MnS5tqMJ4rHAHR5K8ArOCewugGX7zu3kyRtgE1SfEm+vq5HUUaLwDd0p
L8P1nehOTBMrvYoaIWadhfmsSpZZwBD4Vtp99QswchOVFQIUM+0N4d2gIC+AKPXIqK5a5GQdT52x
Mvgrf5Na2OrGIslLSap7E5qE+A4YDeSppPyoUY7mYnvRk7SMlAmoQfmXaxDAY32vWF7UK/p3c+RR
adP+7q6TL1znEGLEm2sR2+U1W9VFz3wuHj7i6RmIJPGpMdMfJHHHPViQ1y9HpuW/+d4Z2fj9S2NO
yBd8gcBKldMR0PlPiIyEHgMA+I5q2NErRxUvnAs0GwFaPak0T6XvHoQajpag3c6++xyMxWMLj4U6
b4kTktQev3F4u53K7Im+gmDn+MSCguysdNjeL602riytFuyrqQxb+W7xkBmy6dEA9EDavBppMJow
jDacLuj9T37iiJJHf7L58/4G4cMV9I3h65JWzbu48GkHslNTT/LINAKXrjvnpCdart4E5FsrEsii
yheUcVpEkhtdU083Bz+gifpM2RaReukWNe75AqWbtieb4EMHDdJfduh1f1SZzgXZCpT4yMae4snF
VxwHmKN7bkvy01wX9f/wsXwDNustOmjHM2UaxYjckrC834tQGmt2kbaAg+zLmaUkceVOFAaJkLLE
FwboXNWO6f1jZMq3pQuu//EVbR1D1D7vB5hOlSEEZSRNTHFM6ikXzDcGvXzv9HzfPcnCg8B5x8oK
2YDObLA9iomLp/UjvayoQ2YSqbOGm8hDng0RzwUXSqH+6Va5hNs7BvU5A/UK4WX/IuILg+Yc4vul
A8HehEb/Lr0+voFaxqKAz6RngTyuWdtRhNlyMi+pqYMvGgWzmWdpOSBEuNCUX1/cjyKJEOOGjD0Z
Tm8jJ9IQTH9GIJyMYDNnAU86vbMXPFaAryNJa3qLZYivY4X7A/aHyoTF/bWTjLDY5bLd/8ShMPo2
CV9X4R+EjyGzenKRH5aKEHTNdfwgefYUt4Rrrlc1cOsOFeN/IgLeC2DmI57uxVJMDJ+ZuznR/uzT
nqqR+/90pCbY1x8f+Qi3AK4DAokBfFgfGHxghApmbtn+C/2Wly+K1so8DgrQ8wUHTTOsUX0s6H/b
ep7dMyh4MiJMMxIqXl3+mJygNF7NwEHqFYI+ryPDFaH3RqVrxWCTLLnxgRnEQBijACUvnKlU0maM
9uquwGUmKrhqrx9o8NS3YbRLJ5dmxMqf1/pzLGRG3dRXgdQmgazJockcvaSNaN7dsWVx1tAJxGVW
r5wDk6LLSiXihueYrIXs8zurb1fjkcbQ4T7ZumYUHLjOzMxly8KNIt+NLiO0cBuNPKRh8qQSKJYM
UuzWOrKvfPISgroVBsFyRoKbnbafOFDNMjZ6I4rT8ZibcIKcQccQShU+2b1KP/AOCfomhQ3rNHTl
QLnM6daSjlSxFg5mTAxaNvbHF3leUqkg07Yb2y6oJTIdRa/PfbBJOWZ/ARQPE6XpAObzXWpM9Yah
TflzAaK4W4R3uFlfwZTIjzKQ3vI4XzBuOzM1ET1agQ+4Fe4pK9BWV+WiIWAlfkFbY9mcOhacsfmE
iR30HJ1iZX8zlJ7YFVFBk4mYg7RbBJJHe+Gi0+AIUOHaIoWXScyl2h+PSIBeO02zxj53C0FLIG0h
23arDUf/ajsQLigq91zyJ4ZqreP39KqXUVu0Jk5u1g1e7zph0XQP7U6cWBmaGImTlQ+/ED4jullj
G2PhZjvluNTRhYtq/I+/lCf0UQgTgQWQ7vECAfvkURkUj9Myj5PGS0gOW8O+0udp5uX/ek875TZU
J19BNUufPDLMM39+QKvxwKez4Nvok/Op1JaQWkZrGPOZKcRuWAOXK+x+7k+1BNb2aqgI32G8fAQR
ToUQUPfaE5JFCIgU6LqsvxkRL4iUh0rsmSURI/6rpxgPY5eJr7c3Pg/cGynfDVkdz3bEY0VV2OK5
lq6+jcZgPUua0CuoeI1PX+v97/MDMljUuycKRXCR6gOUBjMNSe1PzxY6UYX/uEypXpv5gDvYUHfJ
OO/u8PSMFmzEoKD65ysewTuCY+yksIhQr/iXVh3fbX92lq0wvTZOPvJ7QsAc7cHSck4Nurttgw36
wbgCOIfRo9W0heveO/s8TCKU0bYVJGvYTmybsRazG+DAVnMuZ4PbTMB3ekHZzlvFjNoVFrJF1k/2
qtj6N+D6pkw6uofXC4XpOP1kEt9b4qKl6li4YomA2dnSCQxZvC6slmV82aWf1pjXYWfPqsJhgN/D
CiFC41I5fV6TvOJc83KxtACKWy0ZeXhGG2aob4DrdP0rKywjfUqZznyNqACcCcKvRL171RqSHt0U
QcUh55oWs4AsOwAnuFn0riXJfATfRRa0dch27ngLulTP//UVvdhxMQerHtddtSeZ6VVlVa7Hl+V/
bddZao8o8REZUzXFIFiinSbN3mYKWFaIMXIqwQxxk44m+e0dvN9QGeyGpya556hUr4QW7JwX4z4r
zhkU6X9DoRhn9mgg2dZt3XBeSZ+vyi+zNcTIajaZwZI8LHZ0tIlmil1m9HxfFU5wSS2vu6xHj3w7
e3OKEWwN9Vu3P98HNSZ2Wi6+ctOz8/v6bMIwHbtGsu8ok4pM5DaXiATzmD/poJ7AHsEzFL7rzTrO
jG80pMZWJ9Z8R5Gww9DK2vd9QllXr4hXH/iz2xmfBrJP+/afVS8PNFagFEGXhHh6qE6ht6PjxH9N
wVngCUiZRAojXb2KgteTsjCYp60EGaXkd6oV61w7h6AHL65G3/aakag0DIrSfxOf89szgYV1S+IB
2ZYuQISj7dQGLcv17zcNPvlkaUpJNDUuaJs/pJ6M37xmB65Yx7kYLZYswfZi2wtfwjedUxLByZqZ
fmbUS/EdBALZzNQ79OFTr9zUwn9f7fKmfo4wPTqd/SBb8ZnSNduiq+L87oCjqSvlE6QdJBNbp+t2
A96H1FS20o3aKp/oAhME0gzvgSMX/NXWnLz9UmwTVbTw+pAHSYcVQqi4aAaBrp01KurNxLR6o3C1
G5Q406AUMrvJqMkiHwfZ/Z9E/DlmqSz1HoUFAQC5j8HIBNNx6zLK6hYiF4zrmEQJiXhU42taiO9t
ZKFskKNwa5AHgiWZQxQsbHhjNoa/X9F7Mlc4VqTQBJTliwG37wDkyJ96MdlxUuIjzP3oiWK7OX4d
4sWD4YZoolM9K0YdSoPvoYOAMmFajmWVC7N/3WqkXhXzPbhhdcwVZTClEB4BWlOPeRkN8Z+rKF90
Q0TtHyng7POiFgrnrlR+435VP2wC/Z06LgJilbmgxVsjdCt5GQhdYefDQSAxAEDSGgNQHPOuvo9Q
9k27CcOJ0QKdXa4bQ4C9okJ2Ctv+YNUTqgGgRSz7rbCTiRt4TXS/eigT2JJ9zwGpoKIyJAYyZ/ZA
yXR2xQ4oOni3tmOoSgfUAS5dVJ5knsWDaCA7YeVHbDQPEOadTy4t76NwbXteJrNoF1YZhQpuEM+p
/Evn1mj1GKW88xrAdK4Lk3/SARf485o0lFWr+a2D8whwkIHAOTiu+ttbKdyyYuLzs8qtme/3tDG2
ImONOqdL8MqH2ayJVoguma3gdjFY1jIuNSBAbjqQKkEki5Eq/GHIXqVnGO1IbkpjBr38R5EY793u
4v0/W2QM2CaJmOu+bUQvAWV+hZUYIhCZYC0K+fZx0/Y9u/EJIeAm2bIXIsrNO08f6i2ImID6K4CC
ymjzmZSx8Ns2oNvqm1yrvlH3Qi28GESieFGhoLjRVTMNSCpbn5HHlFHQbmo20GoiNzl7qyzoQ0Ju
3BvPFL3qXzASrYHqeLE5EC+GQFdl26k+PLyGmSQSPsIM6CtqQ5zL+X/zTrfybVmmslKbRTmz4X7G
nNfnAUXPz/i09yfuZiiHOpoYWHYD2erh2FrJuwzmLLyqIVKuya3cOPpDUE+nBZOlkGHj3cRyCgkK
cKEAjFdbRox2M61+KyOB4hrY7fX/FQSLAuafaRHKlgivkhHwNzHNYLeMmTf/vVQOxfa0jXfZAbQU
ZMfGWsFPYkGk1s91ByFnbbh1IOwFdfu4O8Km9r1WfG9EoB2vtx0WAZWBxQe8ZzAtx7qwVCNhJGWM
DJz+i35N+ZXkl8oqTBR9F/rO/e+0T+/JbkJWmIa/nLJZNJ9Qha5YB9t7Zc3a+MRjq8s4oRzsxPBp
i+tPyW7zUTZeM0J6u+1WxPJ/Ua2diO17J6n0g6cH5F5bW41MuauA4/hlhF4IkHw1zlM/naNkYeyd
dC/QGTxq9wECRLzSW1JHPZOZ6XURM8GaBpiPXJn0LCMyUZgYb3KPPqygDCM1EaRGKFTJdOTtNAMB
qOUtaWJ2vBQx0NKHAzefXIViXfz30Lq/aJmzyhwdrwv7qjGDOFTewpnMTNtjDNBUKYufJvL9d6OL
+Pt5aE2EXdMsxCRtK89zSFSrFlMK92BNGj7tlw03WjzjTsPAYPoQGXz28xWQK6XnmKkwOg1kDRl1
lUrS5V2j5q2aewp/5/snNInUpoVDE8YfGA6GZjDuw/BWAtNW1vFr+1X+HSJUngL/y97/OPFlOEFh
rQeVsvA08Ng7RclHWbZMUj9ew4BPtjIMqnpg3R7ydnnPI0GOjhax+rIqn7XS4A4blgqrGI6EdC9B
S8EXYKflbin8h/P9QhE4eLNV8A01zuAqLFTYRQEaFSQPIUyMcCDcbAufmot1YCQsy6ntlpdUfBnA
ywMk6ytnCD1EInyDRr00XpyW3Um05bOrn7wtq8l5WuD7gtAw9zmrKumBkdpUusfEE92QYQz6RJmE
LhYNbdq2mZ2/yzRM5cdko/Ti3IAyevaX2AZfAbi2pMaGFcbkWugmUGOpCh8j/NJugQ6r45pYEQ0y
w0EfF7TU0Ip/4SALBsZqUmUCq8UexJt/cvzZI2GNnRBEm/yA5hnEEVFVa6/9R7QXo9cwAHW6FFlk
RJIwSMAxZ4mxmQf0BLPIHVgCNDO0KK3tXQo79aZ2k16ozpd9iVOVvWb2dL3Ye33ilf0OfPvye1gH
c4Rx9lc+D2OI9m4Wv1DC3HZFKyJUxPIIg0cr9K28F/dJ516oBjGyAaBGd/X1U52kAKzQ5ql4XFiA
bLjk2J0pY1vBU0EEbOpL8JsFI5Gu5rCT1vfesZ0REzyLDdbkFk1T/nHlbzPE52462MsCMYpL4T4/
pFkpvPzfl7wCcNhImuF2ktKuaLntpHTDqjweK/GkvqE97pdnaQsZwteuUopiNXo5JkvON+HovTGr
9FOY4jiGYsDn7SeZJavy308OJxc2+j0PJduYUhhKnP/Qdf6wkuxeukVR0R8hs5DQ96u8qPePCtxI
+rkTpy6p+OxMXtjcJ7P6V1ZNx0fji6pFBcNAsYWlAxCgxzXj6g8peQrQRtf3mhnkDXACljDxmyUp
EbtuMUy73l5gAMnzcrDWpRnH4xmAbuBIIIIwTquomJdhWrVRLkNOpiVOkT+kHXt1BVAdH4ToWSLA
U4KUlIEptF2erYkRLJvABF1y/NLBhH4g11Uc8x8knG8OlxAAJK+v2xlEEeDK7LW/BouhUGA73+Pb
zzzFzHy54C+Oo8vYdpFNlrb0YuZf5fn/9RiJDHOCSlshjdPuk3GqCyb4rlpX6xVffLecRDQeZIKq
X886kDq6xOhXSLxUpmtlL9AVynJcfN3Csa5NncC5aWdxWUqRUBee8WewEjiyMb9VYLX2ldAW3dsW
VQSOBX7gFwAbIn7dL3aIUoqV/uxodvQqPq9fXZrPcoT8udEs0qAS6hQrbpnZLIKAF/7Zgs3GDaOY
09bdmVnO7Mp1lvFFQf0rr7RRqOGmqrygfFOhbfYNSnah16x9b1x+a86myx65t8icSPSax127M03N
ZGpTY6Dyv73oGINdbM9p94RNixnZtlx8lQQQZMd71WdsA87PBYBI+aNi2IM2linAhJc4ip071unK
CESbZ/JQNxxxFAKmhz6d32C95CM6DWq24iM1O4gotSIy3S8dVa+nFWakuCgkNsoGb8tnmLrqlN+h
AUhP1c9RO6zAe5knu3F+mL090DdAsgM2HnT1BCLKrDQWqmMBETZYImOx6hJ/0qogj6N+bYdgx+VX
fT3ip2TzBxu2XuceVI2xOxOGyA4URh9PoueT4y5BS+IhRR8Xd4FIrRF5yBFI8dzCaJQsJW8TEQ9Z
PufKSbkiNSJW/l8io4Ps21sqWqyKsy9O9D9FZWQ97E6gATFCx7rf13SfX7zzfSjSDUenqATdwgW7
E7+aicWnL/y4HOYyKiGQdeNzSGjjz+fx4d5iqsf72Yz/PwLyDOtGyPnZW8KAsLTIK/7HBMtQ9g0C
JLHnNfP0Gr9Gu0usIIAXaO+ed6DtzlERWUGXJP19H+kmcK/8cUOJ0O0DWxC+k4HVMDuIhio4LbLU
LZ+uemJKVuN9GfXlK18j64MrjZ6WmZG6+DN3shpuEaZ9+sQYkIRuU4Cqn1LJxHpgu1zd6YvD7uk2
DdZYaIscYzBgi8Vbo4iA6HKEew2QYIVY5suM9hFgdkZIfge3Yl4nd1JvE2JnC73UcxZKW1T7d9eO
rWwqyJyRueAQOccz8HIOywDOI0//sGNUuO0x2tdoVBrN2KKd2to9cy92lcyD7Xd6NH9rNj1yvsjT
y0qmyJsdkHLXKFiabvDoXnuRZI35GJEXmb+RgO1F//LzunROAyVinAr5lduSn5yT30sikBfKHV5f
N0V54qIRmSa+dL1KndLP2ovMtYZT7PKbH7XxacXeZoxo8NHqZBvyAkbvaMCwKGyMOzIFMWBr+FBy
pEqfrbe2fTuPWcNU+22wyvN0Bl0j7H2SeFXBpAe97xLnJjh9tlU4GUYrOMX6zVD+3NIWBM2Adqd/
ANqyJeEnm/hO+82Ljis5yIQyETfIPJoCzto4rVgWNwmUpMbgYDlnMICyjc0M+y8lpJcIlUc4FHNi
O3n7va+vOg4BkvZyZ0qwROoSmfB/m8QwtWLpdhNROE1z5DwuoqsN7uEBmEaSxaHPEIIwIAv3ZwtO
6FSWLhqFV7jFW6fPfXF5Y/drPva3GALzueEfa5m/W/BYSgCEVJmpndoARImsnoAn1HeddfO+jSMC
NrX1EzHVSqgWNIS1V/OkYAbiq5UDK24dajAq1QYnNGILMi17HP71RzgqqZ6tsO7jvFCveSY/n8CE
VTTx4c02GLCfjK4XSUShDAgrleVfPlFLqslBTZfBfkwOQcZ3ljzLTzs3uqlOk/3/An80juS9ytnE
YbmafBhx15mnRbyRLdAxo0pPjinUOKRDg2iRAAZzIGhX3ytJ4k+FiyGEj+2GrYq0IFGELtlwt0LH
sOhtikxe2ruGtcr7be3FxVLcBtYgSA73PD66ami78ZTicSCYPHvXeSjb06KcsIaAiYo+7SUAAauB
pwUAgztLaVuyNjEY0RauWL/tMwMbbSJDFF8Cv+5WZwSV1x7XY9AzCdauWP9Kz5DnPZ2yjyBZJWuU
ApbWqbFn7PwdXLiPTjDAbKaH2kxg9sEAQCjynslnacfvo/ayEY6Ugu3fiWiUI5MrTxSYRn3smSAJ
2SrYD6TGbz6GrNnwfS/HUKlYONCz24Ss4au+60JG7SCltDtjy4IeVIrfcoPmETEzkdoguJ06sLVT
bDziewapekUrflYqE/xoM9UumS212wstEWQJUDcKyhIkPe9rc9OlSlT4UWtq+1Dh6woFd/iIvwHI
rrSKkANdcYSisMIGuMkqE0jimQeOGkE0HXtomZmCbmiIOnl24li5L6YXoSV++GH6CQeTTADOjBPA
RVIR4pCenpnKENpH4WfAkRVJ6hhZPtHu0l3Hk1sikHtVKhHv9R98PgirG7kYZHT5zc4m8BR2kWTd
/ptSaS31T40t0FZdbYKSC5A2hmg3dYqVbjwOv2x3cQK7oG1qjkAAEX5CwcueF0EL/uqIHR0zigvJ
lOrXQENJ0R1dsP0jZNW5RDTSGCOy/tKMolGOjqt3yAuQvgVcKjZ+oLgMgWEKza2sNYw6ndyVEDaG
8HZ33+0CvQR1oopxkWGnkWMrFMvEV2gP/d+7rBBp3PfWQZQHDNqEEzuxctUM2hKbGfFq7JjVgtSV
7XUob2Eo/dQiAhiR2PUFf0uaHGVINpZwtZcaHpjU9IN/5zn0d/tWYtpFS2IkYGYWTbhYfbcCJ7Sf
rgvj5vRl2MYwaQ/OPMVq0Xn2bjGm3whbv+Sbp2KWX3AS3jQl5JsEW/8PyhP3Ksq8J3JbOUyz+qLQ
UUnbSHbOyJq3DvJfel6RfGZQFlnu9yT95sTtgURV1RzvDwsV/lcT2gFwW1ggyvgLdh9xG1v3DD4N
gZyElfC7pYy3MB8R5bgaP9Fvu98n4qAncJ0Okj4yE0PrMqIQfQ2O6rwkcTLhDm3oNtWE9wEl5Ofp
3eDMhXNY4nuT0AXGZLQ5VcI71AFQ2giykk1LWwKjRwjB/EQV71U217s3CiZ81qq5OztwJVCGRrC+
bhOyU5L4jyOnOnpbqeyL5WpC+s3b/EvRpjSQ3mWUhn+O2zupZyG0J02Hej95kStnqaK1P3IWoRKY
YeUftZ7ZELljsMJ0wkrAhgpSWNXrDbCIgcwqxUVx3lfXuwaNkGTY8y3KHcH4R/W4Gaif7d0R9nbx
4dEU+rsri9mtkFwoCaMSOSSfrtd69hfm1ccHM0wAIjKyvTrNoBz93wkPO1uN4Fd8bcH9FpbiiNkA
SH06lIhpm46OoB3usYOvsP1aqoXIOmGGgobG7m0LrYD6CCU9lBZ/j8zErGYQLhtWqBRZOulPlDY2
fzFxaUtYkIUp18h/2KaKP809XDqmQ2BHwaDed8+gUPwwmghf65bvoxf8m1oiVn8SiLQqcApWNbrt
8iARLRY31sK2ucb5OlBsEeV7kgaofctW4IaGJlsbagchqWn+Bb6zDq417+ghzu5AUmaGuFTE0A2U
0Z3E1ONd6hQoWm8YDjtd1QWtlU6b1JBUv9DOUFtKSksSMIubbYdJRW2V2HjwZsRm4CR/QmQB8S8s
/1MMCBFkbd/CdI8VEIoPuae6n9SMjtIla58hBvly/MWXZGiUTbhX/ZKHXj3JakQxMjmqT+ge3cfh
sWveMBoUHKboq4b+q5hObO9ok7X2him+MOzIZpCV3q0eayPaPygwlG5Goo8PNjjoLitye/5zKEhf
jdJBjtTD7KUg8MdckfjjzmF8InfmPhxng3n4X8TChupuail8nPbx0f/q9FWmdpwraauI+LQfQ4aK
Fl8iNDnJvl1mQ996resFkgu85tbnE9XOI5f3TuyXAKG/4QNpyYn9LnwRkxct8Y+9cXBB9CPZ/rZT
N35RxpEncV39xNhji9tDRMM4+flRHizai1t+JCQ/YCEX4TznYnf5LaaIFYUVAoptQRl0UtTflRy/
V1b1Gem/yPdWJmW1so23q6L6liw7fQKxFAAtMKqiu4TBA5duYPJhzdFPATszhtcBHvge+EIsvHoq
2rmfDcc+rYlOuH4xAt9PcoeR4RnraKS+556fU5fKQoijWHGmLsMcmFXQc7tZi37V7fYd4a3qXLr+
V0pm/PIGiJ22HdesS8jEQuOHfZ9ab6OO9Bp4zqcQ2tf8KFRnBUooBYWzIjm5v6IuhGZCyJWOITvn
0AHs6y1pQeJHYWUj5bBaKr8n9SqcDg6+OzJZ4hQrinwftRoA8T+KFMlCWSp7O6wxTjUYALd/WIXx
KObiGWd7dPtRmcfshDkmmAMdXgg5dMQFRXHyhurwOUdc5vmpg1xpWvcctG8vGpyJHMzM9tibhXR7
WAWb3yfCD3TkIrUr8vzaNh4naX2rxisDuYNJMQxQIujX0eYWloJcAADXVsvXf/0nK9lFtcCNSmYI
6i0suHmBAYpzvTEWi4FaPCLG3z/Td6ESICHnZs5gFMk2fbwRdwlhF4JkQChY2c9M5OM5DydrT0qp
wCOY1uq758Z4fZV2WM660Oa0aNGsFbWd6kM+NEKUTLWx3S9g5lT3jC8xqLgy2PE1HQg0hyiAOYAW
j/9qOefd3cHdJqwDr1BjfClg1MU4mBUi3bDwsL74Haqd62qSaoCufZWcqxJIGD+p6a9P55Phq9D5
dNH+7/pqiK6zo3gDiHLVLZJW4GhPt6jMYZYfD0/aLK7PbZfbt8kBc8/67FmQSYol85vXoSlUvQJM
oSli7nNNMzQwoTu0txNrIel04kDxCZJMaYuokM/WASAS0eFhZ0+rpy0M+8+r9PumySTbiGGQiZTt
RYYSZFkwXqTyJ2X8oB6HUg0qM7D/SGAIAcus73m3lLkgOU36r45yndWNMSgKPGw68uPbQGepuWDs
LJFya3rtBgmRSMIYWYya1rSfgRBDS5MoGegyzNtBcD3fiAClCDlEYlmsCzNCfSKes1EzhvOU6y/t
zWGE5OvgHa7j98B+9Z8JY7T+lTE05+wGMhbCcZ7LmTBZf9U+4RZG9/BWuLCKvr/n3JtkU7UFLWmg
9/9bQWM0iIufW+0iHfO+wbTCFUhACAb57YwMrSlVexzoaPfpOvP5GaEhfgavoVG4rciUPDVGuDJw
dWUau1Kt3BR65nbRt7qGBna8o4yF3tRpOhqA+P8eLdI1ca/Ycu097Pf0ETiQj55CN6p571UuVU0Q
UYt86SCvuyRYFlxPH4NUQXhDqOGwXJQZyne2Jhkhr+unBs7skdanRU8rEdBY0ldaAgMvNzhWw66c
aKehFByQ1Gxzg85PmOUV+bcgKy5kKrUs/qswQhIRv+YeqcEMyuT8qz1mpBe2fRjqvolMHwmdj52n
BRYF6ULieEvx+W6vPaaUns4AXSPMh7DGYVtlQ74MHA/v8OJSB/zsd+q16pk3anApJorSTU67f4m7
giT4Ef2CKgYxtVaGcPlZgAT9bFDV1xiKHDM5HHmWsnrM0DMICH/c31zoGCuxEVEnkyP1ZoJwpJW1
NjpcfIB3065sTStBCkzCgoUudDbk7Bi8M4C6y8mxAaS62ILB4wqwoENpZ+i2ioOdFKFpat2+5cKC
OMEiarN2EA6/Seam83WIe+GfVTBCszc3VILmJ1rjxTTn12pMukCBcmuG+h3r9qxZ2GcEjrR6rvlV
jFLh3bUSR9EeobAefg/mVfpg9PUlx3jT5hm+lklHNoH88Yl5HC7ELDM1f+yUJxvjvcTSd62SbaUn
DqcoXjCkXZhcOshiuuBq0muWrEM5Bv/yjyw+sf7t0Qesoi93xh66mBs/+z6/m7lmlmIEdkndGyZh
l5Y403CTr+SEHvjRAmNNMr+TrptDttq2xF78UdaY6JU7NMR1BYJSaE1EvHRBb8GzBcXOf8JeKiyR
syzIRd+D4Qy0S+YRT9m0wand0vCflulvrmH7p8PTigAOgFrmJqM2/rXuBmYkZc3fceqmQBxVJuRs
24iv0JbG06adHGyAOEXEb/Xee5ylVZFsG850/hxvMf4EfsPV1B6BNSxbnyJcjlfGCZRQ505X3oso
TYnrcD9M8KW3SkHTQNXferTUVX81+MEtUK7ryXwqBYo0Dp9VtZ1iCst60RBDpHjg1nKK0Frm0qjE
brlKdcnMzzCoIM2uWzQZoHUtFdJPB8w5hGbxRyvLAJjI61cUlPbrREcJNnTz/oS50pP9+n4xJt5+
ltd2jLPnKSiKXwk7udA3VrH5WhHC7Kc3ko3bjOmgEPnGWoJZQGuuPCW4XQThrkow32+pRI14RWp0
3VNR8YWbBZeHeHVFZm0BoYbVa59NRpHOjxg70ba0Zb5VGK5xHbpp8kjUkBuDqG5GexCkPPHu5rdA
v6eLfl6nTXIkUKP0K7VE1OwIrZG8b0M5EJV+3qkw0jc8bcy994AA+C9milQSV51UJkbIxD0ZWPey
VXgKUd5T6eMF8d7xQTxmSs9pFmI3aqdhrP9vDTbmlxHRxviWTuitl/HE0K2Ns6C3t4geXkhNaS4w
KPjcGeR7uqONdv80c9wGIfaTHhxQIRomh5R9DduzD0Zo8WAMifFQ+cX4zpjHWOodqWq6cu2qKsJO
cy7absyC9T++e8mzBxfbw+m/ViGiUMQiytr+B34iIlNIFpcIU1Ml8H+hCzYsnoJ2Yc9aBdzUe9m2
4dzqf3IDTutvVkF/oU4vMPE15c0//KFd4Q7ZzG/W9PLMz6/RjEcBTraOraRGv9vye6uuvFEQOQnZ
y0Vd61yv/ggHx2uGaiBpfUrFLj270jM+t6hOjCQJtpWvEBu06qLKu/Qh/976JU0JJu/dA2Pd+hEQ
DmnlIWzkmVn28aiiCl49yo7jyEWcHUpwAvcbz8d+WIEqKD9aeXUvj6YFeaitxkGj8wBa7heabqps
kqlP3u2ppdmdcsFPDI7azg1EiBRphTbJIXVyxgbBqDjmV/0So7cWsRKA1EhV+iaWrpB+W14DefA5
kkH3wMk3KHehHcMALsPYK2UvznayiS/yv72aLYAlqohPPaDF00BGawjwn/8iDzO/JGlHesZ6P8Pp
ynBrhQd5z1kQuneeuVf8U0e2wLh1Hc5D7BDCcvsKtSvAiWV2VznAHI5bajo1eT1xMwwAKNVU1Vl9
FmE5NU5A02ROVWJpbNOxlfNEtdOKTOslnwf3eSeTPes+qnMBaCY6l83mo9qPiPXDONUjR35q9JZ8
Hk+zq5KCP6T0fl8Puqr4KYBqMRAE1AjXpETLYMXsX76AyTyMDGYjO/MegP4JH1TSrdVaGY8vV5NI
xzeA7EydF7rqqY9dI9eEnZjpcQio80iE0jmNMiNm8fIFd6unVEwm9Jiyd1h2rT6dKG+Hd89f6yjP
a5zNh8j6Uqq1XGa6ssjSLEGCbicXWw4tKKJ/Abmh1oWReh3yHUa9M2pJQPSpTtUH3CFeVshUX5rn
c8VjNQBtBWcWG1yi7/28ixjp5BahuXrBoqIjl+fXOC6hSdT1WZE8++FvSo3/pIaWy9vw7p960FUR
awEBBi27Y2yC49T2sH3+15s9Y28eYmQ54nkk+u99CM9jYEBrhQkiFMiEJOTAaMiBg27gZwIBsD9Z
V7CmDLHljdGxQga0ds10OfMgQMCNF9CqDAN2RYMOM6ox/SN+frtzdM2g7SsRjh26YlIPUCwW402s
qHlRkpLi/lCtdUO/ScXjStWJevvv+f703qqa/qbtp80m8lrR6YpLL2MlWT2at1w9lvfxSEgKVyTO
akDDOgBcD0qanfB+mVISDW2E/pyiloRz8bCggj2zAHxOgo5cxyh5yH7q4oxK3LTeHdYQX/HOhEez
jIlTwWab6vH1N99aHt/6eWIFeVwBx37EzXm3/wE9BOSXUlOUoJw43CQLx5tAm2RKE6lyqccCKR8w
i66aZZYXcfAbKjiGik4sHNwlbmuA9xUlU1VaG7ewcnvg/kX/lSTWH+Y1VsGJ9u7Y8GQTk1ZbsdT0
R151oiKxT4Ufd3wL+nke1B025R1w+bgGZNgYCA9LZ0MFRtrl5bVZ4fLf0s6ckPBeCX+4OeG0G25o
QxnmzcUGNSpMXLNhzFlQIOaGYEAEACuRUO50br+yzDZ5U7OyBTdc051PnaWLcU5FqB20Q1xuqHnT
U8DqUK/+xFhbVhpP7B/2Oc772C4qKYvlSzQlbKBdWTWW3eW/gM7XJjZ57UFY2T3YJW4BjSFxu861
KzTDt3fg6vz7woPK3gSC1pBorU6mp5Al1ELEibVaSk1++h6+shhF9L0UoLLhwONIdXmEN3TqJVxN
/7UCgkaIT6QZSMa/0dPi70rDIS+ekhhIm5NQy/dTxXiPjTbdZIRVxsyy/oBZWR7A0x1CioymVMDo
zfOw4BwT0J6Y9bz9vybLbA3Ht1MBTNkclQX4r+js/X4NIwSH4Q8WKcbxtSrwDuhojoxQ7AN+n99a
NBHDm5mQriXwX7b60rmYEwnOkSpb5YJYkjM/rQgNEb7DG2KA+ejVbKVQe050aseaC5k2rrJtENs+
KWPVtwJq7H1S42rNuwBuhaqdUkgNNKGXxze5NrqrU2n4GWyvmKbKhG4/84tFBXq96Q38EyMmb655
CXK2cudYne3ny51NaOqmamMbhfeDeQR4p2Zzvgy3F09N45HifXFm3OpXc27XLdNScihFoVbaEyJU
62IeRG+kIvDNsA/xTUqcOj/QxaIDJ5okgpMNCQBNC8aFe/04G//WrdKhm6v7lscC545hEWgvUiMW
7TY+FhkggUJuIWxcAq6swgj1DII+H3OseRvVA8xgEUyYyImjan8fGRouJO2RfuFFIZzd2zYwBC3K
Ey0j9rk/W462xpKWqNyU3idWMOCIzze/HUWxU9sDT5+hkkNnWNvJ7xqOPIe+ELW6T8hPBDKevF4c
G4EDwYsGE72qHZjjquSuSyhPjhdjOlFSra9v9bd7M+IOrMQ45w5tjqGcODvadGy4Dm/e8MQWV7Px
Nxjx6GCNuS4KxyzG5g9l4Os1S4in2h03aUK+BUFJ5R9nVDUDQjKIH5bg2OFhBpVmNh1mkHZrcU04
LeCKfc7cnWwzTIC47T9GECfsElRjPhyvwCPvrTLQ3BmKhdXxJiwTqZlWDQ5Z1Wzbv9wPkeAvTdrz
rgHpmzmW4FubAFpprk7kZ0OUBrAKstPZ5AbAt4480Kz4QSSz1rh/NfyEE9A37OacEyO66CS05+AH
nMcD1GqUD1YL2enaXy6P6TqQnnbMJo4eHlssRBhY+p5RoIR1jYE3yTv9tO+eD0dn2p6lFsdgFSUO
yQ6Q1w424pCnFwcHJYYl+2l6CMGN1Oa2x22n9pyyhQu2HAu09lClYtvH+IRwgPRVw6wRrtw+Dq2y
UoGMWGXQfrtTzM6f/8cAt6Y0ulQJ9uUCwpqxv8rm4rm8DDlgu5EnktoP8dV2foSxd93MY6Xn9LvC
57MCPfd3mwB4wxK/s7nJEMOitPkKR3Q037IqYa7NdJk5sMLVW7HozTbh48usLMu3PE5LRhDE6kmA
5Mu5zJqneOJqhG0yDSzyhRjZsFoxIfH3Gm8uWDQjGqFOcFt69dGPshbJ+PqLmp+yPg9vCvZp5kjH
+/Xe/WZ1UjEwzRzVx/GtQ+3VAANz6UutzjAKC9SC1JUW20JzHWAUFhAbLOhdpDvhjNhbIzNxINBC
t8u+SdkeVDto+ihVWB1mVsVQtGFlRTsJaKjYHJauQf/o0uJj6V3r9h1cC2VCSdcpCAWf5pHfb6sr
hSq/+6BuPwPu3zl9NocDtXJ2bvra0gylxgM4gdQRAsYOttmwOYLIeMNPwpVdi80MT1EZ5ub67HuB
tD8azle7GfGCPSNQqUbpuCE6NjT35CApAH0hCJWSY8DtKzxcufmpX8OlmDdgmWjR4/VLzKQtydqw
aN93vmTs0wj9NI5o4o6PPkUHHi0jGUAGE4jkffjAzktqK/OOUkRh6mUhHOuLtaIb9IARAS4sm4r4
T14V5EZGNzqO8rTSrCqYEbXTlzmvavg7vsKtkSKxByE1AXR9bYYjkks78M+qJ6fXfte6nps5JyRq
o74WZ1IGQhv5WTSn0L1FdMHx2sawKcZ8pmPzcwMT776JnSkk+imBPtWMCB09WCLErH7a8+RtetW6
nz3tsUc6+N5rmRefezn+y2iFEX6hXoLhuBTn61pkMmP6f2JqJ1nspNz9IQ4BCvJxVX8ALvKHPk8v
Gps4RKzCgT4iu+ABveVxx2G8Q2Thmpp/ZKP+8Ho6lQ9rYs7ZMCXN16fgIqjHuXO6gGQy5nwBtZuk
esxYOIXBFT2xqeH+qwTG0/a4Puq67FnG2tl5rg7MFrSAs5Aa9XWAa5EcNEum+nAC7J/Oz8bKaI+4
MajIvCB+nIl9zj5Lv/f+sRnTZ37PQuVSKSiAsIyxMseoAW6RLL/wkVHCkg+HjEAtAPkgcjCZU4Aq
Sn+rM8kwl4POTuAfumgARE3jZjf7TZ/6hvPPO1qd81zqwDqQBlphtvFOV95W+DDqcSkAy06O964i
irBEHCqCAUL5Iw/qvD2IRlEP3DHIamYEcK+MZEGiIMSjsti8nYaoIm8Zchd7JAjLfgXqnqMztQo1
wuJKypb7AFR31aNkCox/WqJ0njIGwiH13cLT9tTO+65PV2+55Wb4YGQlevfkIlnHBqeV6WX1J1my
txdMvjA8i9FCtbB5l6wBVtbSVHi5NpVlVpe6kHWrPVfMcSLCaK8Dd7OjIS71tmk2C+0MfFN9rOS4
dd+SdFb8wtEoSrcm6ikUexTtooGiP7G/Qna6dUBk5xGQg5c8BVTuAoKV8FLjU5VPvrC1+huRtyQp
FO6f0+R2TyweZB2nR0vBLbniferarjBNKH7MQgr83mgtRIbJ/5b9tvIb896rA973knd4bEY+igF3
kGL347+0/5Kjt8AzlbPxDsRof2ma90oy4UiYFNc+AFPBwjseSsXaP2xbDNI9MHIjjD6B8TJH9DGl
OSu3PHJq69QJ70E6SNIyUoXvx+tI0Rhg3tSTlsQ2h3+iVbWwEsoAizfCBo5rSN/tdP2kUU6Bam0t
DZxG5Jwaw6dnG3bjhqmL7TAg8S7eSBGzuxdBo2RkhjAMz0j9it6kUjLdGROHPpMDnWzPPQsltohs
D6AsbuRQum9T+yiNiuKEjcRlrl4UH70HPRGAQHDdQ8b3UHhj4pGkV0DIqLeYSXjD+JYwjSnFjnLZ
Km6RMvpnCWQ52L4qASOtb3AqFfues6qzK4TIPXSSTI0mpTIJOxTfZSYeS7zxLuiuPFVFKjXSeBvP
dQY9q8GrBWsp8KnvXt+9H19solOmL2Gd424oMb8hFJaclK8wdU+AC6qwJigh8WpKEvI5LE31WAds
wD5ytDUoAHdH2EUc4TABm4FgHg+a/5x2t8H6+dW1r1abQUxLRxf/6e29imzkbMSXjL29KaT2WGjF
8z8uruz2NLmHftvkHbXnlElXQ4y2++KQVnT1IBtmWl1AKqK05zrzk0giwB+Mpj4owkDtTI1fKcEs
PXflvT2ZDSpUsAMI0Yv4aDUeTKwts2Wx6bswXBH7gj0KiWUzx5f+2mSwJwoMpVEBhmmI8xtFlMol
NJxB95RbpdyZuGgfMSTSw625s95iouy7yBjmZNEl9JuZldTUp4pekfIN1BT+xVN0vJgClv1zmoja
/5AIL5rHBhSW5S3xBfaRRa5Zh6XRPfXyJN2F/vngX5jsJqFQIEvmiABQ7EipjgXBNqa5EETuEIis
eitnrn6XvpgexPTJTLPVtpAKFmb3Cki+dUI93K4K6mNNeRHWA7rZCyRraz0xYAjlBfXRwYzsVq+d
xOzG4iDC63RWX6uCJ5jlSxXQE+2zlIK5bzCizTxl//TpJAd2Bn6jM8s0SgQ5/vqVgOcnH4OandJ2
QD2v+jgMhQiL3HMtb0AwXRMXj6GmFgJXXG174iZWGMD0R994BN2P5ILm6ZgllgQmfbrXoQf8o1An
NZl03WsDAmCNcS1Ez7GfYesFydL0uK/ZB7aaalJxCDnE7boMfTEFGoDsKh8Tf4SRIWh2AK7yHwbC
o/9NKm27bjUefF/rMtquowjp3a795g+KQgKxx+25pG+k7xu/q+um6OfuLImzfCz7HWKCRayVJOzC
h1I/T1NAUzq/JN/zLOM5gvkBKgP93Q7Tiivi+b1uh72KXBv2VWOoCJviy3nC79hipt3Vho/IyK7b
u/Y7zcqp+f2A9G3xaBQseWK70yEMxF+sKPKup32cxbXpOqDt2ezFcZWqiWTDoHvpGCezskkDkiI2
TzOMTBndpIB0/gqAPB2yoESseUdG1k6iw7KlQFlNLEbS4ut/FYbamq6LaXUY3HtDq4Re1Eud8Jc9
cphSStK3oUjXawxS5vyiJhe7ZVyK3ZY7xKZW68vwWPE8Du752SNQy8YXkDuOIjqzODfR6ZgnJKJP
y5tEDXga2AVPIFlIGs73f7iHr5TqllPVZfqGjFE5clb1dqwmbHLczo295xwwO5yLRUaKwuV4EnTN
XMULyWLvNJ/gIUBaZwhpMsMazMrW+5Z9NG4OSb63JlbcCqShQPB+wPZnwpVcPcc80V6q4MhxH9WS
yGR2Crup+5/vQjinmmAeZKv0d6WwcaHGLwtKx7FNhAPcq/aoassWFBHe2ntr1No8bSabfTh1yl5u
P0MbUxyr0xjXrvGJAn9V9GDGPNrHSrFCu80B4PzH0NVMp+/xIPFRu9dGRdOd85CbaNuH68hQ4Jnp
a+qGArBR8KwBjYkY/7NapRmK1b5b3iwj3ISQfZbFS6g44axouo9ebXPODrAkfXzqn4jsRvQvqzQq
b8FEPVvEA9uvrav7js7g/sm69ctH6npXSet0lFwMxEbHqyJk0nAaRz5UMpsR73OFazgesGPj8JdR
B7w4e3S4bLQn78cgfOxRwRcoLarNp71WM4L8wSD0dlHtXwCPrQ74XDzJmfB3M6qXy14uC6HO1YSH
NZDlzDQSzzW4Rk7fIgfpBwgoPpAO2U1xJj8HCNLt9RPQfhkRJ+xK6Z2NyS3PLeQ8bQJhuOqMTRJE
JInkF0lWAajAuP1ccANCV3z7fNKtf+pnJY30LgcRIUM9j1MMaQEl16TR+xWQ1F+0CxlveVjt8L2i
o/Bd7xm3tcU7jwgNtUFVx5dk37+I7yUYWIM5QdjtkmU9viKa9vluffgBR+Rfihwhi5KVEnkKMsfa
DTwLr6QZu2HpVDDp4O90IIegOi3IH2BJxWBVo0TiVezXUzeTRpJi7XwuIRw69o/5ar55dHLX/FSq
9wM465MtxzJZD2pt3l86dc/rtIo0DRWwDfltQvw1+FhO+vh4/DOuAY4YkedZrxfLBYMFrE0TDHrN
7l5l4jVLphVNpRIq/R3wa9jEgDnZiRSFxmBpty/8SG1IvGDoH1S5bleopzaBqDXPjh32VOrjhaJ6
jX1Ga0aWA8KKjiLfxUXgnqZBCFa+PJkrjxJVh++fbKW8WJv3N/5E9CnCB/L79YmjN6FmIPOsjb8v
XOc1QndO7BXc7hkKCDpJzXblhw7epTonDsf2XBSbNC4sFBv4m6pm2jsuihtdX+CaRwm7eG/LDacv
broPyiEEvI4phOy0AqxGRZb0VlDZcGEBRHat+Icn+69Qe9D9tD8bv3oY3qAgyDbo773UfK9hPbTg
H8XBYqT/o2nPRohw1iggM+SaoNVbYYYMdqMwUGn5oVrS7lLTQ0+jE+QL8iSUIv+cXWZ+jgM0OfpU
TKVgnGh1s5bdb8XjHChN6uP+oOF8jwxPGoTyXH4LVDfODH1Pbt1W29XrcG8bhurHcgTQafJlsDkD
kF9ddJ5yqqosd1V+1zuvwpAiwWuQnF8I0SNJATTvt7L27pa8UU+HFBVHvnYv+qL1ArRG3j5X5l+P
auG7CxYhHJ+gXBLLp6+rk7OCqI+/9ElmXJPgVx18pexqszAKuRFgAMwCkEofMqESGocF5Nyb3tVL
c9TcVd2jSMfN7PHETQbpLf8UgpscJBSPEELwNFpXxR6a6PhWfriaHaISje9j+AiOlOTDDWwuBe0x
zL2HOhyMK0dR6ROPu2HmgZecvSAaVutdyJmN5d4MZtK4ZrIJhGwt0RC8BTD8set0rm4Lsgzt5TYj
tqXuplCu9zUEMtOqiNSsyqNaP3K2AVKETLQa1+je1nFslLAWW+VzQO+1lMQxcDYe3sLyOvDVJDpi
CgtYT1dEm5H1neA6bTE9WPZeKxvkJNqlmFl/QWjWg/wZaKNfJ7lGEfVXRicW19rC5fj3lvWc+LAw
dCGFtIjKS+JT4v5rMBw8scjt5/JDEKQ5Xve90jU6yrMzrJtJHi2xb4PQ1YGpjn6HvUMtDaHsqgOg
+X3zDnttLwS9ZFUkZ3flLiiE9LapMPdmFLKUGrPRpIIqznfwFWVReMG8e/G7QinB9dgxS+UHwX7l
1xVyN8dageRxFSZYQ7ZpHpFJdS3bk1vIU37InpOtu2B7HKVTw2chINBDZVsQQ0t7Dr5Yo6cIYNGV
3Wx6EQm0aAdpkkQOR3ByKClTT/TYh4RVqVg83cJGFsyrmwnKTwF/7jlncxq7dDremXhkH8OPvoSu
aWmrdtF8M2LwHCcoDTxQVMgbHtwavrTUmkP9jalFV/RYjaidazm0or4jA17u9+XQHw+1ZrQ1wHM9
N0mtk+EFMEXMb1x+8uKQMKPLSlh5yfXsBcl7y1thp2//BPXLqEhCTFqt2JVWXYQlOCEGYNRIdKAa
p2evvhVulir83hPOzjQH/W7nsDDOFWwYboObVJ4askq3qBqzfFgF7y51WftxWFIyADrrT7UZZuvC
kQvAoZQoPMchq8dmAkqW6NMsM76QbgaYICQxXgWLfe5XwlVNbcnBpCN8o+2cd77i/tWECCvEmazs
iikns2stDB5xGrIFuq+oeDGXM8CYlgfMnDEmAj3ZO/hZG29ZC+NJzjlbG9fxwwuFhqFCaNEyTiWw
H8gl9q/9MiLQpr5b6LHiF2rQ20Fx534Lcu3kRblAmgzZriaanxAOTKuCg/oQAXAhQLXIOh+Qqu96
RYTVWS7gLVXefwaKl5yntoKEOEli7I0LMpEf98lVWKlDorVedK5CQ47ripOgmwBpv4wFxTu8rho3
rp8cujeqYrpXdLnijn8SxsVafwHjvjACXgFPgVVn0voCs2rNESgfCwAZhJLN11WYzAOn2uRj3d9A
vbpczgKoMWH1V+d18X1aITA6nozZ+PETMCozDfml/9Nu8VohyzMagwJB4lm98KNX1eQPxcbhQKqb
N1fXWzE/0hZMoe+grCj38h22hwvbU98k+W3HAI34nxcnOSDfN+NL3p/h+ycQ8c0fKz+/WgmtR95+
1y47DgkT1QmlTV6RBr9gfG+/OfLQNIG6KKWhw+sEnqhMUJcxL1cLrj7Y6i6Z+UdDjMEWjfGjBR35
/oTpiwK80P6ULYIXItN8lbTgIwvZEzZ4O8LPkgUxlPbu6YS4wfTjNsoK/jT2ldA3SgaAwcMPKHdL
cj1R/fLVYR9W7+0lWXE57gWFuwrnryxUgmVNEHdACg8VpYegzYva58Dfs7KZ0nmA3yQezoBHdrfA
Y3+zE/iMUVbLT1IrziNDw8YT3mkAtxhlqIKt0QTI25C18gCpnPp3nJw1E+c7wQBb2IUF5bYe2Gyb
Eel+UEcAu1p6eGK1oIz5uAY18qx/23luZATJQDUIlJF6p1YY3G2ghgi9Nqr+K7F3cb1eU151lNgK
2hezDEiawi1fLilv1wL3zm1wbAXR8PPENNBVLEgY1trVmddJocAac01IW5+25JXAjWzP1WPX6rqt
G97LPR76WPczLatBjBD1/0EqRifVJxUNCh54Dx+eeS3gWRGX6UvAZZSPBq+47b/VvjshNMCpU08N
E/aQ3C7pcq8ScO1NY6Jq+TUHRQ07/Q5GgpOTLTIBCzlvP65DNfOlYG9+EPg2xJ+o9e103H+hoF2l
5fnD41lp92Ic1uaBfU/8kmy3vjBO/uN33sx/rQQdY9aso6yLJigoeZTTOuOLYFa7BvHS0KneybUX
EYfpEX7vQIgTykXmNnfcJh3v79AkyI7F1126AjeCWCgm8iigt0B2UyrAHzv7+UcvOwFMU8N8OFJx
5+qMa5fBaUOHzWVHSAwTA6xoFY5jL5wAFvzJMt0gibOHFLiFsN81pNpjdQ/TZqgr3Y4iJ1avIuAM
0pc4EX4Kvlp9kngCA2HXujMNImrBb1yZoMX3VsRdPYvqpuqBlJ1edljhSCn9ALOhBzntGcaA6k7G
KRR+6eUmxjow0rpVclyxtoi8872YCrWATJlZyymcv1F0jqdYOxlrXPBaFB1v0bpDEOXVibprTQfx
/GZsLFXcShTjSHU97BRx0uTUuh81ir6+4mK9HQgS8FEYRVF/Fp4b/TezRHvfIND1odf9zZAKolS1
isTAZtwy+14DhEl9wkzaZjg0+22/9R1V27PXot8ZhAANKUjbSmz0hei+CGUWyCJK5o8vsjUyoRPr
eAFcIml5YPyGDR81qOeDMkBXaDGHGcTFCaf3RpM2tBKm5drFFWEMn+wxp0t5IvB805vzuwWUSGtu
JrSYQTSr/s+VP0N/1sZQHYG2EutZhnET6STNkDsrUU5NAPbGeZLgqxMFjAX1O3ypItUhP1Md2mkR
PO45X737rxwRaFjf2J71zo31smKyUd+48ddDtIxJkkX2AvYNtp9kqmylWJb/VPSEeFMTLU4GW0mC
S8Dv8ggA0j5LF4qqs1xHYPhcpcQyYPdHLsUpWipq4GTTfUDjPOBFqtylMxNfHolgu5dmz5D6bxHt
s97le4Pgz8KyVplb1JbVF7cYcGx7ORAedHF9y9iYQlqJZZ8hLYrIuoJLrh6+zsMQZcDml23jR3+t
Q32HNxxVy2IbIlrV5vuQmOTSssEf65oKsDmf/Hj+zfWknPA3wastn2p5hgLpX2AWfm0wVdYke6ha
9N5tSTiw/Ud0F1wxLWvo1JAyIkCKO8/7RseIQ3afrk0sD0+SiM/wUX++NZUrxFCfNjAuZYQ8s7QA
bDCEIE6e9fMXrtOqWIDp03y9eEmypVNRqU4SIPXOUYwnIGYm6XSsJp7QQdegDnPKRDlBB0v0CMXf
um+UpN1h2vr2t4xI9ikbqbfILn8+J2dVZcZHrzYJy/i1A1l44feYVqjELJY36gmL9msDyUV7bDaj
WNazuU2tFiWi3ORWUpcBf+sWhcSrcKYLHyI0sCsp0/vYBdLw/nUNdYxRI/Li8AMrdNr6+Ja1m1gW
leZtuUaI+Ozwuvsl5kQrI7VbdHku13v7HKPQuYbckDvCWGXxxjweZWzKX5Y1SvAKq1PsFn65gTyB
4xYrOYk5iusP/N8ixn5RwfRNkixahS+FvXhDp8w000XJRfVvKrEf/in4ST45aPSJA9EVuCFoJ+lk
17EQCXBU85rTYYjkQP0S4ZLdgHblaZpoWJf1OhYbir7oNSqgPLaKwtnEycEji6tODlYKiB62OaVt
8Pa9Y7ed1FhqXTZ384BmwIFM6qkB8vqk066J4TfbCWh+YK0bca9hgPFgfSrUDMte23RpeDZ2XQmS
Jq+OVonyE9f8R64ef4AF5Q+CgNinTPfVAaV7uf4cesbu1pEPsYYGT5+tFMYMOw9WeO/P5ZacXFFR
cLB+CSxjtdbwHoT0F1xWdv9uhWKt/l/LJRmLmBZbRL3W+w8bT9VM2cXR4wQsheGlMTtIEXg9UST5
xdv/Wpcrlg7CtuOV/A8BIcaClySso5sOvqqBNHt8bc0t4yZhLmlBnglywvAHWhoDXSaV0ugK0KXK
JPRMv/lUWI3SRCxQaxpeH8F5onD2pA/DjCAqg/XXx1tvmwGubz7LuU6nlH916rcXdWn8YIiOoxlm
aQrmhqKiQf/T06MGu8oWkalE+ix1CPdUHDokxdPDnRh+jUQ92ojk/fM3XHslI2vboiPpjy+kKxuV
Ttns0EpiEr/ll+9I+lBSgS7a0lu2j9UOvO7GIz5nLMqzLhVzjiZj3UPzovFu3pn+zSx4jg01vcJl
4mKr4LLRvA9o9DXB9q4Hx1bFi4F7aRqWU9T3hg2rft43Kpcxlma/7LL4S3Lz3pLlugujKcfTOs3A
7v6myGS1k/u0CxZT6sZas8hOOMCMUXgOlvpkg4a0IwB1F7pYMFqWT6DHVtcEiLkEVLHN8TwavTKn
6ziiT0X//MNSKfctFyl0Z5NMwamt5mVC9oV8Og+52iBk1OgYN2cb8CeT83JhS+Uud8igiuctqRiz
PkcgX7CAGeqzhA2pqwUlnRih8+IixRBvv4B0MQnAUZq9toFp+y9ewYMrCeAbx8wMl9AeO/P2Mqqa
0NoQrvNCzsCC4DEFsoGevn01TN0N3br3sVKOy6+qXGLn6XtDqRC67cKSSRP9eCmNGxFoS+NKDQfo
pQ9QCsfDq0tE+LSxDLAAe/9tQ0F5bvfG3UK76XeKKT3uWPanRlp+UT5lKXWHpgSxFQNKfIjVmrdI
LEGFSyI/RRp/32YD9Elw7mdGRBxpEzl5Aac2wUWvcL9PSKdehIsX5LXomPylgPL79ztXqdfB06Tq
FO2YibbiXGli5xGEYsNH8Fdn0uDZy4j1RN31kPtk9ZttZBh56Lgn+RF6U7AAVd3CrP7nRaFcaRYq
MjhvGpMfquTR2k5covGBVP1/5J0ht/ExwnCZV93PtB0W+XQFntDcIxbEu791MmvHibZG6yJTygdK
xeB1CYIbINIJgKguwKVCPu/vomAQe7FRrDoS/zNpqs5TO5iu1t/64oVFY7AWHbxPUO3xCC1HgPi0
zPyxEgYr4Q6F9woekfW+REHVluwRZiOSqhYO3Ew9PkK3bwjrahqvRItzTT9bJWwM8qQE+lFmSbV+
CRjX8mqVGN7p35qdcspPR+hIaRTIVlbGrgo7Mmr6CjI7bjmSwf/6Zw23AWzpBpJf1FZNW9yyi12G
iOyYHmctvmJvoyS4YZ8/YoJvZo7nn6fit7SdhEnWizlXM/Miszv8g0VDzZ3EJhUk+/7cBQRhxmUY
V/rqkPvSkDeIcFXZP1l7yWp6Dd+jNiStRNDIbkQ1uAB9xEYRlQ9tM+fzRm0LYyeP5eyREtNYmgQv
AqzjZXedUX4uLqdrc+1zrYKwzFjcXnyIeopODLoG86GA8JVUuEVGmnn89Yq6TvcQXyR9Lf/Kd5w1
qlOpX6n+mvGYA9h/EGIExr93FIP/rP7etZK7PjXfPqPOahvapxvx05aMOYO9LrTDlTm0xyk9mEIH
0srJ5rFFjWrJ7Vp0L8CQrGHFPB3gzQGg9J/57zu0gJF2q8UZhC1cAcuDZKOnzlgbWTku3pH7tmh0
adY/TPL58atBwkzlXvvyw2IcG++Ex7pWhzuCNCFf848g+4fs9lC3oOv4jaLqvLONjPf/Tx6fx91a
gUwdA0IwCxYpoOFSIpGFWTIYQrD9nuMu6PwmlKBurULATf4cFcfSt/f4gVzpJMDii/9wQsX/Eui2
QBllmBX94R/NvKJMG8BO14Gk5aLeGV9kM5+s2hxgvk3KtFhP/az3Ce6lcB2SATzzFFHJya0cRzbp
3xCLGkDmKDlR5FWiwP7pfQHb7h1CsgBcR6Im0MzbGdXC2T2FHwm0U1P81af2O/HU64O7jcPcDtdi
fMK9mMlS1P1iWrZdvICygexs6vcYOcGKkRv4Z4FBkvQIoFmPlsHCFtTdkn9GhVSlnuWBgjUQY4Iz
SaMEGeNKeCpaXn0+Hp+5QfWhSjn8gOJZUXvT6OI0svclpQ1HENtYrR1C1xr1o2Yskh359pP5Zl/X
LmVF+U+H92CkQsdX09bZKuNDw7j6eEmRue/eT04fpmXA6i6A9NSnGb7a2JgSRmdGt+JK/SeNNGIY
rgw0WsHedaKZxrzM2g6JrHNQuiql6dNoFmMvPD08WXxMCztZyg5Q0D2c2q9CpFBaT+tr4weu20J/
WdpkS4JTHbTaMvooIwbaEh22ZtVg3zuYSxmgrICuQ32d25KOamKZ2nBKDF6DPpn2rNyEQCbpMkFs
Nvh3EgTMPDBPUlbifwcXmCrSl3mW4FQXMqdpbLNdfbXMULt3pyWOoeMPLDeW3PI4s1Pxt3yyd+B7
3oBK82P4eDt43OxoVNPOeo7Vh6S37ugRDLYOL375GX8Dd3k2yrd74nKuhwaHHHr5g9IvAv/TTE5C
GG1d+nJ7zsTjib8/M76VM5x2q1vQO9gVKoy/cS3Pyz1TZhgmZWgUTDh/aTZuQyOBS4w60YwYmX8u
WmJnNaEIESijcynLvF0QAsS4wCS9V39CVmU4p022b7Bp6n9I9nVUYbmAHmME17alKd9XgpKGp+4X
lJaFQlgId7ScS5xV7EiF9xyaYz2rfGOaftCt3lvCFJGyPH2oBaTRFbAy+vyXO4obOTUlKvLpm8X9
q3IWjs06fYNaRVL/qj7vB3w9GVBkM7FRoP9Gq0j+M5ZwUhF1/QpCPFfOmoe7wk7tzjiQocqqtwOK
RHRQQiALV0pHfpwbphsx2o/iCZcYGDZXFWJmTgDUxipsbPBXTF2c/t4Y+B+anfVdn1LDydtu8kD1
V7Qj4cKHyQ0khgm4sdy+Fh5atApcsFIqLmGOGZEE7O7YSNi5MIh9eYmclNZda4vWxi/+VoJN7YvU
ZzhsGiVqbx1bvfNBz296LkH6l+wUX3aVhAzFOFSeq+nAhWRI0fq0ETS4yB3hrKd4wnTZf7l3sIuV
Iuztsy5Kx0pFslCRsziUa/82DPhT9XsGE3KQA1wvmm45hMnFxMhFHe9G82XQd9Yha4VwU63k2R+4
uaveTYhcjb8qmn7c7qFuv/HlalqpHlXt8QOb2AujRU4WUUlxgTg9D+uIbhsJFauN4X/fHeYXjs5j
FH0jSnxgwTOhBHdrW4kZreRg8rMmzjtt6ardLESPM36VpPs8RXqK0D1ZC0R6llhEnGhGCcEvwaT+
xDAQE6j9lFX73aFR7ydp0FvnRD1hGpV5xYfqaHT8f/aepp91rd5LqcUs7q9fc4EEtqpnxfznkowL
1ZszDprURBb9gfd9K/W7OVl9z+gksdH3h4ZsE8rrbNAl0y7EvZ5KDoMSjyE8nlj0fR6RPjDHMfEk
Mn+qr5FuUwh3+Y7Xjt3FQGnzQLdnQOjDHQNbr53Gy/eIn45nGASzt+18nJqAQ8fLSPYUHo1fzex5
qisbSk/BPILkQaaUx1Iletp1BGMntETWgs3NQUh9Ui9ILD++TWeLREk9O/bkE3tH+6wiYqAXuUTC
S8zArAxzFA4x5QtIMqDEoT+0NGJf1jmuQzdLxIOfgMLRrdR0ns3+1s64m1WoqyIJOewsx8LhEAfK
9XAAnW4of+UpMd0u/kp/rxhXiWDxHICwEsVNh2oz3OLQ5HjfInvob5TIjOpIfbjnJUKXjBZiHJ1g
1rjxC6No0EKBRoTzH51TpEEaRTpnBbbp5WeT0BwboNHPJCx6AvQ08fK3PRTNSMm7jqlrMAiA1nbI
a+TxhrqrKICoFmrO9S/uO8XkYDxkNSkIedN08oTq3C1HpfnQPUgPQM7RTlSihmL3qDBN+Ym1YlxU
NovYslzdqTxx0uQauzkYBDkQzEPL4diCMpV7wnB0LcszVkCBWz3AXOsEx9UhzGWTgeM/BC+IG4e/
MfSK35Yd+/3ro3Sak/nOwPNrgpCIgd0HUR4EImLsmZoWRyeJh760bTVEd1ltP0Nm2UBeQ+C0Mgzh
iI5n+jlJIi+adGZtjQUQxNjXJAOZThufn/uFxcUi0j9MGNQQqD7NUuWBrWGxXStzIO5JVl5uwjlo
QMjvA8unQILrvsIuoSRr18BodtSbWU5y6jbGiiPU5R7jbZs52R6KHwNXiJB43cMf9B0jJwlB5aC+
EHqiyQir2xscbUkIwXttJCc7vKi+7v9xmuiQlyGOXz481aixo1UT8dJ68RHZNfQM3pJVhy3x9SqL
9ODgYIhtplN6W0jBOrqbEPWEtcYbK8psJdKYqSAgbCSEFKHKeZ8GwZ+kCK4bQH0kxaQ9eUj/CITD
yCVy2c/cc7olOvD8ruN8HFilHMs+IMkWwpC7grhJMbaaAtxepf/x9KrYLqhNru4JPW0nc7H1tcld
QjSmde1p9ee4BJu1kMwoyablwb4/KSv399hJ7ZdeVOAPPP9uNJEbD9Db7W/nNb3RlS/WZCIVVgXG
6FGJTDroJS7NgjmfkXDxa+shRZH5ogpIZCo4pLnOjdz8O72q4ddnwtDZDGU2Z6KXbGHgq/S8e9Z7
Cc1ILH8xH8TPma3XyI5+MiznvNPouv9ySmdq0RPF1+vjcXwPJS78ZPlmCM61haKe456m7rsjZeqW
//cj78W1+pBXmmJaJwVKpEvNj8YHvKnKMG11hOONyYSldAATxk87KwiP5toIlWJw4Db9SILjiZX4
CzByoaliYo92jcN3Rrez6BLIMp1uCgDD3psurmG+X320XJkPwZygQEY05991cb4I2wKsYa/43ae3
D23PwMSOi5lM+i29OxnjNrgf77vTmeOZ03NenBr0nUXIjMO7zJQdDB4tfLq0hz3FvcChM5OjXLMV
b+OLMvpBi+hjKStnQ5qZVX2HvlW5RAggU+csKMjubwSqWl2GO0XcOzWSwrzmzej0soTqDJoeDqkC
zNOmUltAT0chPMNWKZDYqPlhGELiXxhrYlh5yiADsjayLfdAmjW28pX0JmeFb9mxW1Xh4HNjLUoo
XW20NsjnL1moSSHRv2JnA5iEqVJRPfFwuMlOjmQQemM4OJiprapKlma7QwkXAu5NXLh1Rt4BGC/B
chY53hCuAxWRQ/3EO/G+0ccrNnjHGBkvD+oQEAQQzp7vNqysQmnueQbCsudMzk93S2GORuHMz3Af
wvCXxkWlnedbH8B/LJKgk8amcCcnSDb4yq7KHrsdX032yrW1HULCXr49WkkhMHxH7/rMoOmzAzW8
IXukdp7oMge9ASZ+ElF+2KlGwmkKhU4c1FfmqD7fw/GL7ih4xkqwnNeTBHMEcCgjsOdvzBStvI3J
Xq5pno/NgDfXnBNEs2N/n+JbbGExKaAJjGup8LkAzIEWzIEZjbFS9ERWIVvmVzNkAOUYPq7OHeFc
Q+zDx0IbA4wBHb+8T8kjWloPNJ9hf8HVp4GED/mU50xbsIssJL9FieY1BUckPNdMhQZC+p+yggAN
uVGjFMU57Brytinx+mQ+VRW69cC1+pvVtjmK2pkcb9UK9t+jTeqFGTVDPdkeT/sdRUldfSxQRXaN
vlzi0ItlwX4vuGysA75ZzG3cvcoTETBGpAMDa6egdU1rYqcDBX6UsJgP6OCAkL85jvYZvtiKCEag
Khy6Nzh/MiGvCw0oKgAheypccV/tQ3X7MRLUDQNulCPiu2Iq0OIrY1nSUq5ao5QSK4vd7XcVgH0A
oOm23r93if+6p7DRflsckaRAIss0JW7nVdNdJMD13c0mbBlO8DAcxFDSCytb80yRhE/l4WuVGEWT
AvmWQblwrWwbFaz/rkLW+okLirbhEWjQFLKIC9KeXem2GJ2WZkjrDQWrMr8JoBNL4H3n2/c8So/4
hOjFIwKxdVbvYDhRE4jKlncwFaVz2mSgzHocCwncUMVQw0OitwzHSH+lCU4YEroLgOGnrSDEQDSu
sn3um2C14FfpLxnpKYq1ZgggbjMh0ZmqO5VHHTEI6J/zk5WeSm8j9DUxs7bpItedAruNjConnaO3
xld6JBpR/rvCYpCawvd6H0uhEaoQ3NsFvLKqN5rzaBbhZOHYDdfYKDMRXyllX8k9iPrEsCT6+4/D
n/1LgR2bb6bm8myQPKKXTzEO6jFTCjhRO17LWHQFfzEGiw6tAV67w1OMhREDr9HwjM3h5qvUB/Ap
t7pFuTyPVdd1xfkBcf0GrRM0/hAGpxBdbBwQ2ID7OglAwYknfcMPfTaD+Z2ZZ9/pmlclRlPe5Git
YUoflQ3n/J/7CD+JZHx+/4tlbByPP7acZ4ZwQLPC3aOz99xth04PtRWo0tGXA2dtRq1TaFfE08ug
jKCMJx3ENc7tfWjqA3a0Cnzd7wPnwTpF2R0E2jw6664H6QJJmXLDQUGx0Z7e1OZLcak7JPqcuWzQ
YsuyazBpHeVI+iWaK3I3ZkQvKR2hFTxTLTmIS9rNbE6R/HXJAG1n1813bU2nbX1RAv1WME6dDX5O
Pn6EDRe3jR5kFBRG75qXoJ3wi8i5Jl+kjTCIPV2La52+1WfiEF2CLeYkPIv2KBzZ+lmSUEr3HaEe
DhHeVBAVxuEkryi3f+wrsGCmwOwDGTuff1op66pD3uFBaZ7imBUtYqJDsXUU3MbxE2K5q9FUkEsE
zONkTMZXSwgIUYt2tdVpcCd8GZc5OscVCo2vIECGNRcD9PGCOy1M2CmC0kUeE0dMlt7bWkkaO2Mx
eqjoGFiVAPs/kNOBm7+w28nw00bB57UlRDAItzpZ7XZWBMWFPGA2o7nk3/FfiXT42ZAf75h2Qe1F
dlZhQDqRCV0HKXkpvdPND0Swx322LUM/CVWjhfhSQ1yBJhB7T4h20lcWGBBK1GONmYHfkA6lB2xL
onmwp65pN1UZtVsgYCDunnn1VluUgxxKwds8TSbIpPSRl5a0AAQj7wU6K68lwUvqTkx34YQdfvNV
0odvIOS/gkBvXv7ORbx0c59dbM0mSVdSMxqEA3P6ESwiEnCpKQDn2K0MYpP90ho/jhAUBs9i6LWX
qAgDJvfTHcJA/VHW52vx170PigaXkjROa/AneXV+KjDve6bRqI3mhfuriP716ccLbLm7YdWu2AZv
7352R+xPLdlMH7tO8slTPEpED4oRLMQqMEqVFJHPC8ZTmJJs+yXilkN5hZ+4nRd0qgJi8zPAiMAR
dFkM7Im3SLt8ICOt8/lqPoh4RzKZfTNUkcFXVwiq/86AHniTqiJeVsbiC9x+lw3EPUFZPJ7fLdmg
fTM30bFZagvETRt3yBwncm+alXbgMyNpiIYhQO3ePWZwKF6BwLMWLgb+ROAL+pTA1yVLXnMre4in
HYCybBYOr20BPAGWIdKjgQqTtur+RjQ+rDwf7wKrdyQL4WjeaWVS36m39tKkf4NsYR+s6mzzLPa1
/UPJWDfZfY3eFBJaITSzMHzUKCEs3i57IcVOJ1CXpPg+70Xk5FUr+JTJ5lIphpMas9OjPwD2mBny
Zfwp7biAl6mVT6BbDgoapqYMbE7ebsQoJjmxARwlILjMAORlA5p68b/yQxW+bEfRMfFM++ySXNiu
5PWk52ZErkmrEdzj0NWyWJsAt0Vx28WgLsfOV+fV3EVvZHoVvorQEFplxaF+DX8x5/qTnRIh9oej
G4eRuDQUUh0LYuAEva59R/RVn6rlZzlC71XB82l8A+E8HR2uJb50yBk37z6gbYAeGgQV9cWKtPz5
TVNzCDz91kmvquroX4NseNq9Zp228KTN+JI0BgKOhW6i/ybDgwEv4gDDnn04RF9sMjtjinywAaaT
kqjIyGHEYEk4tK8gZlHyr1+Gbm+HB32qjgL/g/n/08rsahoG+r/GDWGFKJwawLoOj12a2lHU8dbT
lOy+pvCaapREc2BUATk7KIW83qbm46Z/F/ItD62dLuYCBrev59XbmGrsn7b7bkog/BX8tQ8MjgTm
Z7QuEBui8Gpo27ycuBUKiioIAkma0B/KS9e273NavU3SSrw5V9JwdCrPYkzy2l8AQMI7CK8+bq22
7BtqhKhBwF62WDI0sdWHGKc8Su9hwZikJDj2w15lXG3GSZnMOnSaOc9oFPzm14FRJBYsKUbsT6ja
S5ZKPrLQfFP4k5x4uavyRQNnGY65bHYuWF0OTBTSQVJtHzkHmTFjzQHM7RjRSAO9pnGnAfdsqFiL
GJ4F4ER05ppNYUM47WtvbteeBmBnHkk92ZLHxA/ITh/cRD1Ktyjg1sovnXed3F2eluiPmtKJbKBp
FIDWr9/GLixSxvODMKnmK28VwEJ2C3pXAHHT4RSCNdpKkhx0iH/3glHJ9AvH7qJXFFmfwL/r/TEL
HrW7VbAXW40STKr0vP1+/bvbw+ckvRmgP3wBG09gKtlazCPafZhuPTZ+Ud1nuVBYSi2NRxOwALCH
r6h3R8j1MgeUb7j+5j1iVBk8DsUIOyZGak5ZLw3JK2AUTfg/8Ox/5MQTjo777z+te8fqTRLJdj9l
wXJvuUxu2Jg1lrpmdGux0ZiYeFsXqtHU47q1QJyePVD6uftvCMxL9quBz/M+1z6fC7pDpfE1k1Xg
ulA+1vex5ujlnXoAVTD0SatBnh3WjDZsf0REOpbe6Sa4m9hHjXxqInJD8RkcoqbutSyjtZckRZeO
AlUuwJWLQ3FK7EL0icCEc50i1MIjQeyDCsXFiExA3yLmSEYf1rQflC87sMAdgvGt/D7zMjkSh6fC
rvUZik1WcZO4Hl2zY68vxNY9JGoc5LwXTUu4x2BXHIOvCX5ZfFwXNyfPkEZr/F/K30ntGr+c1ZM1
LYQl5GLsKnxjP+MbSKND/f3bizlsLzgwlIJ+u72Fawipt/yIMbPb0NMnrhxakWXaG/X7CSt8Eb+V
99qxPYFoNjXLAFLYNaaep3Q/DCKKF+sXHis8nDf+RCE0Ccg1IcupSgYR6FwPixT4k2x83TcEj6CB
JrEo7QYFpaoF6iocDTi7VfmDYBsaBrSxtGBynRKoj0bpv3mHTQqbUcyPj6v1V6y7jXDjPYxRDzGs
G4eshSZ7D9x3/o87vsGa2SI1bdjUrmRIDzWnc2aXKFEcqZk10PmRnaWhIBO6LI8IpaKV580oyrr6
PGXt+7rpCaVVGPVCCTkp7+1aRnL4MrIh/Eqmum8mLOjCzMjOXLb3P8QnQGZnq9Zy4oYSuPfBwf5B
5xZKgm0nEmJdLKzjQTzF9UzSd6sv5deNBrh9QfjpjtoYjVvFu8WPOkzTrLof2/ls7XtE9YYdI5ig
DKZXVCae31CllQzU+pbGk7xJ6giam2qXnkUyUyTX/XTNp30YPjbyDy/5H8NHpDZ2KrR2HGZYDgUt
PYCOu0FTgqd/SzpPRSFGRdctrWGf78/zeEIiUfxMq4goVtDUBxosLm2t/Ns/PG0520Bry3xlxGzb
2eUwk38A+wbTpqgc52Tg/rQ9zdGkzQcpo466xis6cXcic+1+d9238s7HRr1+zxoVzZ2UDUzEEGCx
Y8oH4kIANoHNt1bDtoVBRRq2HExF6tpQEfZ41UvQnFtGbcvRRBOWlq00mCmefCwxP/I+Lg1DKPKB
Ro360MuVch9F9rXotCYGNCr9dJVNiD8zVdnjZ9tMDVALp5HPyz6KjXvOU8B7ogx8yOq99QBtTuRk
jU+QGkZiGsTsTtHo/eP2ZbsS39uqZwgkgIR/mkUodqD6CfSbQf4dizDsQ1vp9OwgIoG/stYiVP5x
N8iwdJ/TleP3EASxv364gdVFcf5lX5NQRwJy1GaDbSKOsRuTuM5NrNHaslv41H3NZYT/Dh/Rnc6V
M5Rw46x8bPpNuFTJDsNQFtr5E9OuuwaxHasZzfmRukD1uewZph7c7TC100dc2a9bcBJn4NuY5X1f
nrLQSw51MoTx3sWXCkAtiuYnyS3UapL9ZzqmPTtz7vyiPDI+1ZivkZ4yIratyMyzADRS6fy4QVzw
eiqoR2qaIHsK5qfyQkPuer7wq7TxKTxbGGp1EdRcdH14NA/HFlvVIRT0G4/NZ3AgEy159rKWyN6X
92SR4NGdPZS6Um/9275vZiHfHWivFpzfM4nPD7T1RL4YP2Y8qDBBD9mCyr95811Npha0JH1IemGN
8Ln3CT2ihKza7wmagUHxLSD6HaMZsMcr/CisYEcOqBd1RSyiL/vQPC93w8qtqE5V3il6EIaxeJdn
1Ds4MAxDVySyE0jpXBvJP/U7vyzQo1RmhKN4A39T3tIEZALpWGfD8STTqhkm++Eid3Bntnhzkzyk
/n1BJdNBLmFXywoSimQVtQJQi9fsh64H9yZQjbhCEwHiHdgzH+dh5lJ93/MnxxGD8eo9zboCQ+tV
KJClVSfEeblTVozygu1QBfysg06pOLkkNOyjY9HRaPxCy1Ff0mikdFZDiHO/cs6hFzuT760nHoxP
mhArjHS/2rEQ3th6/B9CVthivf16lW/7GMvH9jE/xXcJu3tAtDWwIWhVcOOEOLG7OOJzU9ZlxAvv
5ET3jv9v4xP9fk5dXFOsWJMtOu4imwvG6qwnVcogTRGN8EqoINE2ZazO1UFHxfzhgv54a0t7Tp6+
9aWmmsAublXSSfMEA4GuSdrcBuRFzy5Ct8OFSY+9fgWF3l9QXYD3hUkIvEuppnYM/PIhAK2YWbjf
8RBQzYCNZd+XFHhZ/tipg+y7j/hP0WEL0mnVmbchK6BpoG5RfILLY6H6O/TPwN/jvGBMGEh0G/Pz
3E6zeWrlSr5lKyQT98kSda/3AGZG31Kr12rqN64Cxu/5F0qdYOWixDQjiGr4cGQh39b2FpbxcRYw
rLbD6/1hjoIhXP54LDDS72M5EPLMXozXOlqDLqlPOHeCFfNnje72peeKn9a+MSYUNIdGShEZ+36C
9Sw+kbIYGZ3+1ql9HGnttI7x1aWvYCXAZAXWcrlZSyKzoZExeLWQCyuf0YvTGJToxlqFTuXQLzZR
ChxL68DppSw3ELnzJg+2AbTTg+bfXjqAjwFOE+YUgfe6xFoxWfVNpL3gEQaeAMlSsd5zE+Yx2wrv
YG4uqAF+6a4wklhH+vEQDVzoz4YlKjV4lwzMPmCCzsWkN/KClsgeaWrV/l2kXtY3wldQV+Pk0Q05
ptOX9WGQVPjXyXZfPFzJmGCeU1iH6Mmb+hHme7V1VSWFrZ8e5OY0AKOfKdEiiGjLh3Q/Cgv0Fasf
BPUyY1kzp0FJgYXQqberqBUNW/LR2dHTH09SKrTFl1t3IlmCNJBhqmEDSa0j+THUXziJFonzQPgq
bznqlQ3wecvwwKWknqFFfpyr8YqJCrM4FIV9P/YLzc4frfE2/OxKOhwgDbawGY0BjSCzmH/NNaKu
PcIzGJ00L7wYjFUl/Oak6GNcYnjAM1H0biUGPe1N7VOHgDiKj7Q4HFml13jFmh5eNHhQaEo1Ax+s
bNUIRx37byQjF6uRwaHEMKUj7x/0B14mMfhctJV4CA03fXIdAX/FKdzE5QclmQ/PJh8tYiw9CA5q
isnaXA+7FgV8rgizHlaaXzUPs931GYUfZUp/j/amwQ3iLPWs4WQu2VN6AoLhhDmYKCWYvoahvm2P
txExzH2Mtgn5jCW8sJZdjk3D7j7XhmoO1Q0ZeLVXoDe8oDUJAima8jd4dckHhjrYXwui0hjOhbDK
wG3rMEjwIDQUU7acLzGSnUwzwuV99LeiPD5ahyQOWn+HnpJ9sCdCvWGn5kTF6ZA5NgxxQegscwTD
50+KujBoon403Pio0THlnl/DsQAGoSqa6Fu/EF7vn0WKDNugCUWuEmvz+5BKf2HQLKpOhKaTHow8
7+XJswHoI53ajbdQE2IlmrmrVmFCFyfgPFb17Ink5EU3FwX/diU+5ZEoKJAhJ8k8FWdOYoA1PIlu
s9OzwI6uyKwSD4paaZzPw7c+aBduMbQZRcocud/8uDuIcMqMxCirwcqwuq2MHkHkD8ImOCzw1Rvn
JUpqCLdp0yMTxnpGByO9oT3SBtakksJlZs45sG55ptfCE03SNysjJ4EaTwHxpXyI5AXaAiJM0Lj5
lV/7rMBRQpJl42IkOG44gjnfMWImxhil3uQmbK+BZYjfHW1a//iig+1DU0JFBq9Lfr9fjdfhpDV2
Cp+OgkjR7oF25v3H5sPxJ8o7Dvfyq8tX3/rFRCdMfhmpD25xMo3MTyp3WoxePXVOSpHDLaWldwJX
RrLYMixQNMyDqa7yqaQLYlDs7HrIP/uINjZNtGZUjXlE0CjiIA0o+rx5jwfLgFxXK0hs+7gLmkfz
kszXNL/taeWn8yOqzS3yM3ndbcu55OnrUHpOlLIqgLLMhwlDVR0hM2DjmOqJQGHPJAc51KrVtclH
GIv/E2fFYguFtU9xuF9i09NaRBvYDVuyziBDwa2b4Dn14R9qhyh8UF9dDlo/SiYAyxRScejioqAI
x98Omx8ApyVhRua62Thc4xcWGRNiVQf1r7zqP+p9LGDCLmzRYJTp7JCXaAfR1woLxLwmacU0wD68
pscwv7h0g2YqsmXGebcNrEHnG6MxhZ2Wxag0QdrE+wSj6WbLgWDZplG3tnR6vfi/Y7c/l3u38GfA
Cx6dQpUkZGeNUoBEYya1og/WCQNArZxjFxZqY4br65/f1TGW7lb9hVyv1DosWMWyfKUvDVMlgjbf
eKBzrpbamtr8USG7DgWVc0BUDUcBCztb5nlUThOQgXQhjqDkjkPn2MI3hs0XKRCKJCKE3Ju7Fa5b
mkYqtau3EPliEot3Vgi8CQp84bluTMS2a2aUJ5N/W+H3FHgiS9JPEqFhj7MfquvIHo8OaqGQpRWW
uUfT94/dAWGPUi3gOBQeDc59ujRw+MdQSbNYmWXo8sFhCckmn6Z2zYgFZ9u8hRR6RIYcxEg/w+CY
1F4oj4eQWrBzqNS40mNoVOawXREVwkRluT3tSPKtdJkQxSI9WRH2KUJrZC8G9bDrkZDBxsA/4Mdc
9NnawdZ0jTU6pF34erujUM7/+X0QmUkQIwqEqQ/lMVT35bErcKqg7VgrRTuFDkqeRkceGh1MlaCU
IY//iUKn3MvWU1By3VDmsFrARGLCh1ZJGiJovEqw2fXsxhD4pWCzE9oWfi3ZYf59u7x9iKGIFPW0
M4mJKeBf+AAh2aZkxDBYDlcbWLSW7dFWLZBlQaS5HzZbMWrohWW4UXMkTEMIutb1K4c1KvByqN9i
3VfV6iCyRczQRJ7/ujgHkglFAAPP4eduCqO0h5vb17lC1j5Oh/gmvYOjssxkWtjgWjHiKrlYiqx3
i+GqKubAAc95pTAScsUWkwWd1YXchvxQ2vxtSjGde7yxAc/Gh7iCZK53uo7eLXE+0/7k8V5EVSw1
mRFEv9Dx0+IB8/KUOQQEr87EdkAHjRZyOq5qDrhvJ7g/k5YiSr4Ar7HZvgJ8/sYEwFqFvdzQG4zw
WCzqzqRNtxUk1SVoMJnXDoHrne4nGjOUeXdbTW8h0+8rZfwkxZ7ymgqDiA9VXSIeWGdXudsPlfBt
qounMC3jpcOnapjjDAHx1bnUDn37R1FD2pflHB6ug6eY/MEBeOX0oUgZrXTAtHDoYR9y/ep4INRj
IS+mzbzZqW7FjcNw42Yk+C4fd+CjmbPce2IaBD+fYkuUtaJh7eIbHSVCULt/MswdKwlUrB2+1JFw
64ThVADkNSy8fbn5Fm8HY3kJSwOeD64s9h5flLcOH48TZvryTfQ9JGkGUFEakRsg4kWZHyePNb7Z
DyTh1j15e3pHa6vbnEqGFkSUXKGTp9IY9V7XZWAHy37MH6gnbtaqmqaNXM2kZH+R8DIWaEPfIzow
JNLvzGT32jFyIq0hD8jGDPQea/tiPo+RNFoywKzgpSLEey4Yb7PP2ScnJnyxpA6kdseUnsgWWgCF
gKMRCKDCUzNIXY2JL96nhhRaj4C2A6YSySkLAQiZ6W/eOlRJ1i4n3cVX729TltnMqajVR4cE/ly0
J19CBMwjAzOoam9YMjJu2xR15xYk1pXBcADNYAmDUClrzmnP7ldMboetuXnlUaUOqHf/XeRjYkHA
IF/WUassOZarP7khL7rp4A7fm15+gvev662frmCk6n9A2U2vQ3yUhbr0kGhnSsmnHdtY77chFER1
pZ6NO8rW4Ni5ylfDiwckGnS7k6MdwwhnRu+vrJtp2Eho/ZYJ8iLw8bcLzGqHquf4JGS5jhRf0Bx0
1aMKBdynJzPGErXYZn6tYS9if8zykkxpWRW6JDltWgLEgmOKKpOmTWSHy5rn3J7f5MQanQF8oz5n
9UxdPZpQKrkO7ktSQcnjXueD02rfAo46oLuuSv2fiat9Sh2sjJrQP/SH5D+57YIi3+usLcVXPIj9
n1GcVTo4//SyKlQSTngczOfKSZJ47h37iq3pAsKFEjuwJFaVK/aREaUZQnamx34dSTr4VTemhT9W
1ttxIgb2YWkqTUTxfbOoaQbP79J1JTZqrWoJVyNpM2tsVF0/Y7a+JJyqU+ViiX0FM4/m+97NpTsX
+7wuwmAaAZ0nWzD3kPdn06mABp8TCRi/O6os58HJkaIpjlMulxIANak/Z7mhPq9hz8Wj4zvuPcba
IfncgCZd9f9xWYLdvSiFSXQgB+QRnuClHO3o9SQiDtaTAx+O526vORW8FSUgvK5a3Kpe0z7BYiZk
pZlFe7Kkfaul9l3LORs/SVdi0zAehKzTz3OM86wnutaVVHFqfmioJR2DTthYlCqDPiq3kateSJkr
c9HT7DQ2XgyZ/9DX2l+ynjJMskbwX3Ep1Rr4XyTEYibYde5zFhwu9n8E/haz2Bj0BGa7RF01sr7y
Dg3GmYEbyKTZ+p4GlDM9tm7QojTnX2pwXY8BxZJm21yFXJDnCD0Pai2XjKH7hGT/zZReLmehWUuB
R00AdK8IqhXhHiOKrsTN1eOFmIxWTdg8fOCYf1c0f4uVuQFJXfMVzTlTVNMZSujBij7qjigiqVYg
Ab73wJ6dwVwputCf1wbMnMouRjQGlYRfYgGmcjlTVBILxyhl+sAo2miuBWKQhmC8+XCmBtEOrL8Q
qQ7R5H1wHPJuuvfV1t/Mf0PN65M1yMTDK10qDSmAeQdn/cDsLNBSKNGQdskiJlddcu8ImiIl8Fv7
YD9OiL50jdravYoLdXl9+yr4z1yYkyVNrMId0UDfmmkTzKBYqt0G4ig+01nGPYzph9aqwtgZUTmn
gfSPM0BaQ1uH3rR+8/BBGBzg3cm2YdcB0oMdgHcspsl5mF3Gq22yMc6HdI0STCMurI0tyR3DXlwP
rJHMZfKgohr+Q9L+SgVmCdLXMBZXv4kcMEjsIbzjETmEgmThqps/6u8SkfuDm6+RgQ13dsjIDWsm
S1vvFNzhVmyYaX3lKxFxjp9DnxPiEsmDJBQ4z7rVJvQfjy4q8Z83OojgSuqaLCJaTsTxbdSA70b3
IfNOq57xQHEbsEYBmDq3nzSTGIrdnKZrerY7mDz7PR8SXt4KhKrYoMYy+vlj9Wh7fn9qU21UBXLy
gwPoZsaifBgnWbRso/uvLKlumvWcd/Rc9hvNA9oqSHb3YT7sDgnFcccmEfyAmlB7MND/72R7armM
aRaPojxgeJJJfqhFzWWB5UfO3pMWIDu3kB+FyNE8c3ekwD0VcmXofS/W4J82G9jrlCR99SivBrpJ
EEnFvQR6oYNt+UyFbVj5xcRtXiVqgdW1cAm8Evho6n0PneiUZCHAtE7mFouAQEvdmwWp82it4Byi
t772MFkEsytP0KE/E2N8kCP/4R+G40e8rkEcF5sT7jRjvu0Udh98YyGLiDiueF+pbi3gH3cVNKUx
acZ0K1OKEFklgBJJj//IFyjMJ3gQddRPHYrwMSvIeM1oJG+6hYzlSH38brj0lw9zKqucNSpO4gEw
gxTVVzrY/zC6h5/vUd/Fq4NWVYmehL3YwzxLqTlnqxHxoy+fI3AG72+ga7qUsamsTxwbuR/IYRuB
Ltfjqi9+9KwvdkjGBVx850icT5ct4N674vz+7gldrBJ5MHFF7XrwuFhf1DkfFgmvIFf/Ur+aMhj2
IBCaMIGqx2UU5SOSbmdu3BSZhTY8iXVysr5q2vw+NvzkLun+CGAIvzrGW2D9d6vKF++KQFlbFccY
BOhdPkYnPsCZSJQ3ynauWbTiY2EksUHRAk982wVUyoVdaaoSqwUsj0QrWoV2ElVmPmea/1wkwXNn
Mko4RcxmCslKuhx8apIxUsuGPwljrYEJIz3Mu+eIR1kzDNtplTDdTl9vX7QNh+/Y/f7ueKdtRITx
O/sdTvvtVPSELHbKLsZKHWC65h1ttr4XXxWJvSg6+U8UkM39Ggrnri0MX74WSW3xi8EaUh20MJc7
dtmGmru9F3xHWw5C+fj5NNIFBVMPbLQ7t4NCpaxs4E8ijhHPCITOAPkGRIWMbF/kQLn2H71+lgSD
QKlKwp0gWzmmWLm9kgOqv+azohl4veUl6h7bpnLboRPrKOXna+VtKHiur4saSrPathvuWQB61znn
DuXFVKzhELgEWD49fAB5JEQ0lWlnCf96fzB2hmtWa1++HZ24sH7BiM6eYLjdIRq0P/WXe2f9rzRS
l2xV29O9cl8xWH9MYukWWJqKzXJIylSWTQKWNvFB4CytKiVjCv9CBRXaFVHdpJ5vhaLzPGF6C1kH
0XGcIFxnh9/PXLuGWWyGvZXX7Yf5xzcbTXGUpN4BmFk47a5YWFCZh2ARkV4I/FGe89YDCLbnPbfh
N8OLCuk7uWKSHEgJDmnpTo+vCAsK20SeO58FNyCkipDCwIaK0j6Qe4zXTab3CafYKuESqPFUmR3c
zcqjFU84AbGCdPIKofFUkMtjkquSKta+rqnYsyy/I0XDWvJY0qddn5ITK0y/kFjUi3qbAGbumWdk
6d2IYeVRyuCRde3ciIyujexWytxvO1VO2cSSTXwv91gjG5Yn5Ua17SQe6RXqgC4zO5g2lOZLcFln
pvf2FYLF9UZUbt50GB84SuZ1dmziAJHujAtsMMLl5AaQInr+rTlMhlxXtKNx/i54s9CWDza6cn5/
q7GjrlSCtSSBccB0XlaMWQBugsvO814TKoH6rms3b1eNnXDpNEF6Sl7p1jo5Tuj8PH2T9GNSssrR
UAyDW2x18Vo3D3jqv+OD/rca/W9yQ17we1o2/D+G1rY9wxMbT/fzgIfzm8DWjWLWgyC3NbKXflz0
YHj8f/q7eBsu+qBRDSWdnrCq970yFN7bJPQMc2R4i5VM3i9WBXIsHdKN8MYDSpgmRksFv+cSpWCY
JAPvJ+hl50Et6QhEJ3JHYjIgGfvGpG9edRgv//wMxsJTHAA0T1jlwVthrfTlQZcELLBFtaszRxlQ
oINC3PYzWgFdvtKIzUTUdAY2zgoOY4TwMwiRWBmkkMzhQpUgJ+Tbqm2sEFvX39xOSQmAhDsYe2hC
Lh5uDixyVtqb5gppshF1VY5YGLWrC1Ge0hA0sYuSCOUU/GiXxmxX3Zz8N3XuTU1IpP2UA6nBvBXQ
FjNNHuSebjviCejN33K0Lah/VYdN0+GXgCFtcqi7E4fDyXbGgx0GfH7bPwk9OqlLNhPfVP+v9CIF
cwHzUlkG03IQrpecmXIsCBGDpsmBYmvplZ1MfXHRMnjyte2fZVud5PFqGSTbrqKmVbTh1oSmGCOO
B58F3TXfu3qefOm7KlRtFMXYZWQ7UlEyJQsnLmf5m0HrXHqp/Pyz2xQR7PwjGfxtkktiSqsejm6M
W73QAdRKt3+Q9OBVPCBorBuw8jzvwE5d5dxcjm7Fbzu6hIyYinHl3YV5KDH1us7KMNCiKv5lKPJ9
QoedgQpFP+Cl5xnyGsty8GF0f/kuMZfgLjxQMrjc89dI7b0IFNhq+jAliytjdLyzYZYVBbdiP+zt
Ow/zKZ9ovCvJe2LiYJaExGLP/JcnnG6rJkPpkRWb5Syd98s4/xJNLiZ+RAiEbB/3LT01JzuynC92
0ydMSljM7gDMQfRB/Iwc8XcoV3hdsCcZZrqllJm4IrxtUvldWxEyUg7PEzU8ko3dpzJ1dx9gjh1b
/2HK6MqKflWJcW/rH0iJ8A78UkF2Jovc5ziuXc0QtBOOX5DYumVXg8dflzxWaoFC4GQZtIhNN3BW
J4EDtN8/x6ROwysn3z9LjZxYaEuUbHxxmNLAKpNzcOzyJ8Wc4oIiehruSZfkr6ystSMKwSJdpQZ2
+uyMZXUijNfWj0T11WBQM34MpjA19zYKavEyPnZX3Dd9L8EX5WyXMiBJ9fL4Eb5gDd86LFho56Sj
dUNcw+GCVvF/PjbO/zBXlhD4C4E0s0MQzC8EFOOzafSR3x6DuHkizKYPN4m01bemdCHkSW/JjI+g
xyZ/3AiBKlzer2Xz2H9nqpSK6Gvzs1hlsIi1ufsHwWhnG6Cf+6fTrllzev3jKNmiIbA1/+LlSkGp
4ebG4GnfRK6ST7gzW2P2Rut9xgX+c9xP5cDNyUyfmqroc5g9cHi3kXWdk6xIou416W7Sf69mzR6b
I0c1yVE9xLXHaz961RHMkB59PdWA6xbMNG0Macj6o9ykPGMELc+NUIVMsWxBj55700o5SQS8JjyL
MCNXj7IF21+vECpVREfmv9O6qt0aF6xYvskpKnoBuD21hPou/W/y+WMATDtmuAYfmTIONH3QDLVy
Dla6EwmCZv5Q0vLvMyOj9+7Mp1dRKQTS2ezucKhBEun8oiBcVHnDSKwD+UjJHZg8dJmkB6BWXoEL
+fMwN9lLe1uLir9nrY265WMkffQgcaxRabPoEenMAyJr6rVA0vfecivfZwl6eR5jMAOFjiEqCYWe
vszAQEIh8xWsLTOf/oyh10IzDBlti/ADUQi+c0Q5cy/WbzDBKqCIdQbV+u07RQbaaZEetjKWyCFy
pK8g9z31kSNKiFk8HPzGZZllY9ZgHtUZuKKe3iHHZIh2oAzzgmFEcZqV8CuuUBhi7Ir70V+i+cLU
Kt9s3CmTSLAaXtwbwkbo2U/NjSdliRr4BQ7DxIXuVcBTg2uJw9xmYdL8rNEsVMUrkwkvn4ziOh/h
wdecUW6ECAqYfGoDAzMG4Kjju0JtPYwPlXDmbZ9IYoIZFTclDx6OMvYuBkbs68R5mPiWn0jYap2c
C5kWqiDGMTFuQnuq065JiE6keqLre8E5u3bMT9IGyJADaImX/Ilx3ANXQhstSxH2L03pl+LWW2yD
QQT2QS7SNOl0snLugFga14DlXSLGTM2NPoCOhzeccdXShpDyKeviMca2rOGTaohPsK/fTPRr8pWd
w/qycRYXFBLMNV3qqYFCIgJHkepPqkNzzw0E6WD8HQw3Y8Po9/Z2E65ZGbZuN2wQJxVnJ+F0QIKh
gHF5HaSFvZXWdL1NLHW3LeGjEeucjOBnPZq1ENosT7v3BTG+IiIN5Pv86096SxfCeTkjtPBsUEyL
8MnlF3TzGe1vPzi2GT7GnAzqvNpm+aO4tnpBiGeYAuGbhT6vZjAgVEH6VTYVdcviBBBuXM+erkHW
gULDN8BRK/mcdGTuL1qMqIufKKzxNWhVj/K3CFj8J72C8L22UVzD0ZOSQXD8J+OsSK0GaHwZi+DO
DxQ1LMJj2rMn4BUjrrXZ8yXkTL8MaZ2n+SHxVhqpQPPLurDnYKtJ64xIb2JPiS1Um8EtrKT+z3Ev
5vSMPkWHg99wsNCkphvvXCHnN0VKssYLQ42Ow31/u7JsqC1BWakdbIDjxEXw17W9OTRdw53mdnD9
wi/C9thcV8zlWEylHibKHOyl1hGADsoAXk2iRhEUs6nEaq82YhCvOvTbU6d2j7yQE7XiZxL/pvYH
NWF0GPA+JNuEo1zJnULwiFsD3AGAeLKqa+j1He7s0M76OPoqycX0D8M5mhagzmZw+bgnckIa6HU7
6r8Peym2ilnd+YN4UPJ12gp5WQFcu5yJ+GGM+mbE9Tfe4eQ8GxYLzPaaerYuboRJ2TMQtyEhsYx5
FwjO6d4OV7KVsl8x0Ru0dRUHbJgacXhVbsvpJSO/AmF2mP0JH79XPoUr8vGOwiNt1D4Nxr2SXm42
9JTMv7GJf1mBiomb/LD5UrwSVK4fkz6C1c58Aw2FCk0F2VAyTvEfdNgT4zElkpD4vSUIXGFH8t7G
omxESERIfN+EMqccCKdzXYYMy6GCP/JpMt1Zcze7WyIWKCnqVAZ0J/EnJcAqYEsUpUwIwUIViNuw
ZgzchP/+RyzTybYi1qREoLOPfyl7FvY5QnqtwtYXbDMHs16BSINQyNwxMwPazvpQLAEGI8veq0xr
yspVxmtxe/K3BYEV+y2MTTpfBXfUmQPAS/mqCBnBB9K6BJaw5/gDwumm88/BW6T1MllvKCDF0U83
ZFss4HX0HryDwswNQG6urJk82dMXKvjUqrjlMADvA5dRDyklQFXy9wu8OBUZyRJaZpWHALVYAv+t
g36KJWSOhdsyXy+XThdq8/uLE2A636a/CXqi/dHJQsqO3LUHC8mRaQ6m5dSUxjWFzfKwDkMawVcm
5VrU0/Ac3YQ8h/A8Hu/m1iOhaAxhy9EulUhZvMvdvBBkRKzblhZyOfqfcszLNM99grqEigCtQ3R/
fNFVLTF7hhC/OJYYHUxDaj7iK2D2/uV39evKUeORlj2ja9NT7O7ymFagcFqkMh9f36gt762EpjFZ
9V+NzksjOAsJYO10Ee0GgzrwO0sXg/Anq14lXA8FUY/2kHAE2nyduZkcFGqafPxKx3DZjTwVdwKe
ln1JgFbYOlxy95+YT/4oHUNDgEdrYq67pORlUxGjIXneFO2xW49V+5eeWsUEjuZE+ZVc9geCCnBp
8u7p4Dll6GW6ZEQHMg0YjDSJ4ouGggWMsDhPlTXGsyAsfCXoGNFJNomtXJ5064Fi52eiOUU4OfHt
AMEy7Eh5bhYYQNSX8TfyU+pj51qW4+gnY5p/fhXYskZuRsLKJhJZSSSXDGAhxwLfZC99K9JsNXNC
WPpgbDnmFlizkngQCW9wnZRqqYPU6CwWeuQthvdMqxAezLfpySk7ijmQhYgk9drJZeZ1tzr1vDPO
SyoYseysX935ew/18Ru3M5+5t0vWH0N225AezZt6hHBsVZI1E4TmFwe9kGNKPypLyR6mWhExuhcR
hA316fOhZVhnQsfrioWQvdDk6R/RYXSscYl2ae88yejDw+POltgXV774IGmVK1m5Hd5rHuMA2adR
tWnhPGnbah7WngldysYrH1hW4duz/ZUfxCm073KoLjmdMqdENkJQgKa9uQZtxTTxbQQxqA61U2Ng
PNSHBF7ObqVtTZYiHGUpacj+D66E3SIoVkvEn/jIKYPMiKLah9TbC7OFos5CpvCgP3OWwhbrLjLy
LuK+n9/nF3d6dptB1S25g/bLVLxfX7iy07EYLYuTER9Rg3fDG69TYFIGx246bW85CYgv275jemRy
CP0vrPd6PKVj/mFSEXgwd88jTBmEKHeTpddHznWAUSYXjbpgpHuihbkLqz/HVN8aMu7j7z/l/bqF
KhYbD9f72D0I3NwflVDFcz4zMEsEtY/ObTO/aN1ZU+mt2BLL7wMNRuGrtDPYRAreo9tH1qvO2c20
zkWfQ02lxwFI7bgn6okPRnR4UqmIBIZWbP6a+2rHLhelzlCc6M73ZYrouLm586CO2O0tNLlGJgXi
ssRmwrQ1qMYh1wn0vkN9ihX2a8RIhDHLnKr/iRl7FVLQynnKiVb7KZXEiC/HgZH2LLkdwaZ1FBKv
W8bRsq4DsgTwoyozR2AR1ab4YvV31nbdJKzmjrfQPGsC8dEzHCjKH1D99qVtst6bemxmuPiTOKPM
AFBj5aCPfOfy6cpyWdilfbxekd7mJScX3Bi+lqyMdKGsBNHOcQk9Y7SQ52G3qKvn4XRuc+xGVL/5
DoBaY6qqvuStOa7nd5I7/C6FIPqg+uRmuVFo2DcIYUD3EW+FKFeB7wJdpgpeWCaURrt8x+sMxjmh
s3yJK4O8Ryd45y2RoNbYFKmzxsr7fjKARLkYV5qtu0lns3Q1/kQazDH0jMdPzODJ+AYyiAuZm/9A
0gbgxZDoNvsF8TYTOn1BlwXT2GVQx4Gy0u94+60MWq4tAwjf0No56ObvItXLaQy6/I6Rl+2jGqQf
7gzz1ByXve5BMdOc48bjBlsnzizl0Fx2AQZxGIPmZ+miLQavp8ATBXKelnxUyySRfrYdnbTSmCz0
C3kOpXIoI1wX6K6++87J55ZLN7w6WxzKbQAiKRDuZHlNZsUyo3GuzxdTL1nAj9wPyi/RNeuzLQ0p
mdxnxujrNmx9BeubxoumNI9qH/I/M54S0t7dUOg3bTrpjje0RwoFrcH2emUohVxqFqZ0K5NlteGb
qh5b6XUrSMzzm8ygWrERyzbOSz3bC+1lX27zh9/RYZ5ieMgeQxk9plDS9XHcrcMDBszFp3jMwuE0
2oWTqsBWUu7aBP4EmM9Ynx29pUJiOU4v6PkDuYis2i5Mdw7lBIwbRvkev0V1ggFE+X8h1AZU2NML
VeQA27QUI2eihY5oJI/YtEhXDvNSGO7OpcUM7NHazDs/Jn9uq5vm/JQHwE8tjT2qilVftfqKQJIk
Ltq+LLM2+VbbkKpdNYLtKT81XGcZG0guTQ83c0OkTEYT4r6RxS/XOljY69U9doLBklex5sE7CuoR
7CFnIvvpuvyRkS0vD/6FJtaSa+0/XPBMEsJJ48pwpeMZmSoXEt1q6dH/wwZo4eCBKYNUChn1cOrT
hBwpFXp5Ikt4zZFZ++ZrrTH8SwYc+BtNFRd737q77GV+vS+mv2D6Zhx+pBJxhbxZUrxGpO6Ojn/v
6IUswUfEnW8K2gjBx+DuDZ58iiu2qUzelfKVlSpaftKk870M5OTdpKUvapvFMzC/v2JFtdNsxSBG
ifbKgd1tTblQb8ijHCcHH9bAlEfF2FQbrk1R7fgSENTi8rCia/PuuFhXwcV9i5XjepPhfgYOYnGp
0soxeK5g4xgvMob5hThiyQq0xrnSHZPQ1Wjj2CPZJYZTnMKQQ8y3DM3z4QojKVjRgfzS60n3/8KS
QrKKkKJgWd/sCfYl7dV1dIqiFfgG+dgEMuN2vMoyVrQKqJ/QCuKRtHQqJTaqZr27TcAUIuW2wWKk
m4hr17HH33U/OFLL2vZ7fV+pH2qDKsLkkO2h+k7P4zrEAEFhycSmapeUQs1+pDz5SOmg8rczapc/
nykgIE8NeINYc6ibjClcfhrxd/gdTb3fG2qRddVSYnkayzG6SSdv5lg/4lM1hQ599Dgi9qSKTPLB
ZSuadto/7rNNDFtetScH5S/HeYcofS6ya1/r6/XyW0lNUwCk9M4i/Kcep49Y3FGqMSmnL+Q+7dKM
7oi/RAboRmHabxRzq7UO5bGUg6wzyUcs97S0ILUIRDmX+cRrT9NHiIxK6fQ4liVsMMx0wm6RjMvm
sBiythQgk/+6l3WPV8GZf+NKsalSDFNH0IjpLFQSISPJ4yiZA3vtQW2pBc7+13u9A7H/vnQ8Rgzx
thai+Js/z2jFhZUc2iGqZtVk7uYJELbGBUycN9PfzETIbYKAuMUBvnuJn9Avpg/2eY6bK4peQrjK
nPU1SmBDv8o4wn+H3Fvsr6hwfCFd+boRoy73nnOn9ayK8ROOoyNW8cPpKvZ8EAdjqz0zj9V7urS2
2DtU3lHLCpgTxYFSYvO+ftv0Vrbr899PxHKHFLspavWEAZGokvlnzxXHpM0gmHeY4gB5CBh/BuSw
Ry2Dfb6izeIGswntG9qvK8rk9SegCkhDuszXjJwdxtUH9cuya7dCKhmLQ3mzDmUSGsFh6fJV9ThM
/m8La+8iLuq/bkWwgR5unuXEV4C5D3scUGFaHd6nDmacsstGGaVrkFbwgh+E6oSDxBqf3z8I6RkC
FtCv6tpJ4DnU0Ui4obiK2fgeeWFblM+CqSTFNAysMXJNwScAfXfSMKEoBWF2pjnvjjd/mkTgj0Gq
1K3aLOF6ips+zA0Kt9brNjhO4quXxkExSfQ562RQgxDBOgDQukzTdTOlyStpVIFlgYnQbmYO91uF
kYbCRTx2h1b2K+ReKmVYbzbmMBGgJl3W1rzMIRW0ObZLFnIjXOwhGW8hR55/tcokJoutE5yrNkM1
ToEdOzBaCl3dWtJbJcwOswaV3v9uSyqkhXSvq5Os/elgsd0ThdhdXX6Gu50msOUgiUx75wy99YH+
/v7fClP0Nzq0zStPVXrF0lFQ7LGmmkNEHoYhAbCG59J2q9X89sA4/j4IBVy1pXQzlovQ71vLMP2+
m3kQxGXriozCEymXRUQH6Q+Ib8n+LArg/qqQTlbKI8Bej4EJ4xcXa8LcXpxtprPa0+dgIKShP5Mf
HN212ExbJTwrHqj90orcW2ggK/MTEbHmIDhCSK4S7hC4c1DQUoEfi5O7vNn4nEF9rK/JXrFednrY
hRjCTBc/ZaioMflttLoxmZ3m0uYyE1pUG26iPaRsC/8LLWQamcU1W4Z7CCdbxMRKJ0ODyVIOTtR/
//r68o3qK/F0OATmcJfxP24Hd0AukWcxjLu7gweHdyz3NM2Bzpd0w8CZEUnmVBoIzFOB6oxswihJ
vplnl2YncklevnGvsVRhRbA/7I0HQNfthCL9f3zmz8ri/c4UjZUDrEZkHbu3IA10m0c/bSBYYKaL
nBnjzHUimUHgCQPzebbMzmD06ThTsomPLIX2LBofx+3wqEHhoSwL6PBLj3qVXsVj5eASoGQtwWz0
l1rurOxo+s3qty1+p0mIqwA2qpKf57sFHdArdam2daDjc3RVo9J6KpG7UN2/Uk500u5kL80p4N+u
bLLc2VqZRu0mjvVE1eR+P9ZOme6jMxj04hKq0jNkvA/YjBbTrO0RMj63jdn+OeT+xx2G4+RZnP0H
aMHFUHaey1P8alTl/u4mRA82L03v7dB6fJZVXq+ahDYCWSuoVWm6dZc7PJcwxwk/8jREy/w068Hq
8eefeqcw249mNGUpHgnH3C7BprM62kER9SikS+K+NYWLS4SrbOwG+//28x/svLHgDbO8uZZHVLsh
qWAfoJk707Hhiyj+FzRY5B7KLbQLIsoXpBnUMQcmPHBXWO6dERwXZIFlsJlJ5grsUND3Rdu2PWJX
4xvURy62slPLBLsoNkk+4ukiCTbslfuPh5Lit5bizwPxc9kZVh8QyK6k+TAPjwcPLybGGI/ZHl3F
jR3oCJQ99DduVbc1Lw3q3+7DG5MoepAzfZQU3IQq4pmIrcPhpjCO06GGRDCvlb8cjsdoq5KAVUVu
4j6I8QAzwLqr03+f8P/jiWBMrdt7HUAG0nGc304PFKTQo3TYL7K3K+h9Fi2/ERsqqBH747NEwxSa
D3DPYpYvBOmFc72zCM5HcrslAiOMD50aSeEBPtSGtj/EoL0VaLCuY7DOaxFCsNB7LqdUyNWvSBmS
6JXoVE1V4KwcnnfIgBEy6Px63XJeHihmLjbQhbJkF2NMmFvKArDVv+QLLYo/O0hZo6R26asiLBPF
QqUuAeVefg1mWAs1hUSdtEQP1EWjDJTHxEZ2Vt6eTLQBtIhz2I+WxkPUwTpd1Mm9117ArqJ9qs/A
5t+JZQZGnZA6DoupKQ0j0YMjiVwIMog+C7rbEfv5b/OlEQlHeq7S3I+blXhCjuFHbXwQ8ZEqHiwp
Iw4uKjZkmxIXK+B7exH0Z9kVc8TGBdvhhcyDE/ZczzKnb9tIxN37brha9+fhlLNMmeUasJxzeOsL
RAobkLZInBlN1qs5t6ZulRXHfvDyCsp/+v/NaRO1Gdk7Yr/qyt+X0R0hCBcK0TioXJNHJoItBpR7
j96C2T+AwvoHyYFZzSYz1WROA5QAp3tbbgpKbBFTLsro89olMnMu0Av76VqjewD1yI5dGYAUC8Nd
VjyFchAJ4I9JTKNPAFtPaJPrcX8OsbwE+IXpQKfBa59dpPtRdxrRzXjDyjpvoIsOqBBiXC5BHGbk
TQ40sWnzAmiUa4lQ061UQfIGqjCqAa0Tmt96S8y1sX9pcUHyXzU1bJ+XncO/tPY/ua5Op+hipQKE
WmSkfbsi9lF+bHfPLi2kDn8NMIcqAv9iz8zmFm7n7P2TLJZy1x4YVrmy0O06T6PhI7jaE1Pa8epe
SY8Leaf909TJHDckRt6xvKTUfjHfJNo3YEH1C9KUh3cauUBfyZHfF4gE0eDYewjIIRuwTcTqY1sB
/xWTVjOHgl+o1dfFfmGYPN1SeOGhZJQ/lFCxbvoiz4XAF4KDxgZZV7cTfsIelx27JERtjFZMSirs
JPooKBwxd+JYDtIfRR8nNGlyivjQcayDLLO90nREOLSH7AjqZufH6tAbuXo8KcfUYbQHgasOLrkP
zRPfwZ83CmlQJ9u0OzCSs86bwPO8DcbiCcTgLchfbHDKP1QEe2aYrKm7TyEp5oqfGRNweNNrd5AU
Bs3Yc9aEVZEwDyPF08uwY6D19XG+59uRNXovmROISooG+C84bnsjmoEVFOtwtdhX8XECCiMoVNFZ
q6t8puRMSTXGh4z6x7kuct0LIWrC6W90GL8wMMv0UKdtej9x/oeNXt+cRr1GXvI5du4V9Kvl0RP6
9GzmwVPxQGxm14e2p6mXdZtFP8AxppsV+JdbbxJ/2enTur0PUaToFp+beiDYcQZiqHRZqhioXWfM
S0aZ66qaKOFIxVJiOAAO65NyOjRxL5mjaUuPgFkD1Lv11kvSP6e1kGrlUDTOtdVDiEjIzl8iEz1p
gN2ZZukD5QpS18qDCxMf8SxB6pOR+XrPtDesVFUQbnrPj7aijdkDX+uUq6ch2tiSNUepm7qnGXTi
vtzFPy4gG7VwdwdqrEKJQ0DM1xqQIzs/TG4z+b08/+b4WbnDSZVak7g1ACKIP0+t0622kpWQgN2b
moiGvBuJ53KnzuutyubuCIIk/q2hNYmQd86CsNtxIzBK0l4mAqnyxxgxxd8dnWnue17tdD2CjUch
rhd7CPYAb+zVIYo9MKAC7+IKBYagKZr3FNeUXn3b0XO9+bKSJijq4XNAnsvDuIFJk3QTkYXT3WDL
xmX4BRLs37OfMlV6uFvGwARaOx3nRrEaW6tsrr7tD6w8WtJ545S5FM/nW6ouUN1kyVwrtrZJUQQn
DnQlFuDYidmUJjr4sEEN5eaqTaBFQl1VhURD/diigz1ZA8GGNmWpenqfrRuHz5X7I9OP5M/DAEgi
IMDh0/3VIIzaFm+DyI1/X8s0GLaac/4Wy0v+kw8XZoFmDVVpZf/ao+VztWr/2O7nIiv1yy3jNHYv
1thFRm6iagNRt6DmyrWCyYHJld1ylO8G9Tbjs3wDUR/glR0ploRKqZxzQJzKi+HA7aNLOS71DDr3
EmCmWg0Du7I1efxrDPD/WMb5b6G7J1/oRILt+6+Uq5Lk2jFWfImwR98VOt0zdFzcV7mFtGXjsZNU
3ETbJ+gBdAfoXGgEDfpZg4I3YPBggJIGzK3BrmiYeZsjRcqE0M/ObU2E29usv8HrA7CpHwEkDxgP
k/lNcLKQOf4S0GwsBFdf6KmrYtL4p40KqNAOQ+a2teVHRCG/0FFzZ2plEAmn33qJTXM0t0B9hm1F
VCfXZBC0dRZ2SBPcG2X59PULE/akc7sPczoDe1tep51o1sRxvlghojYhZ1CnnXO95t/scSBhUNCR
r7e4JSIdsPxoPV05zpw4ESLTP7DdX//rF1nvxGQaIbWt/79IDxoM+E+2M9QWkf/ZxnehkXJ4o1E5
W9BJXhH5wn3Lxbsd8ctnP+SMV5qxPQVExziYPO618yavPLeJ96w4whKA3qq+a7pquan/b0/4poNN
ZDiEfdbLqdbJAhXVrjeUqHOakMZCmQwjBEqFyVid1G8Zy1/yeo23cIh+yNF0zmtFASkLpTdq+NxE
r+cuLIEV0XlSEuo7UjvrpA9iuJtJnuWdDjtAK05P4Bqg/GmiDCQmxv5wWuV5DJ6xUSfY8L5LMevb
+4ysCg4SqDaxRpwbXH4axzm9SxjggO7bi6380NHz3qFv/Bl9TL1PxJGMELqJ4EFGHOdyTUL6rJLY
mwg+HPD/z+khj1Hs+fwYEbc82qayylXc8/hFJgrWqD05Hbz89zpUqq5auU8z1f+IdUjjmsBSSFuV
NC2nKAVpTaq96uIahoQR4vGNWczVU0LW1gEPQBihVjnWw2WJwtkTNGzXJZcJHsxyj7Gwruu8ZvsN
qG6Bo1IyvNCclwHufqGwY2T3flpHMZgZkCw9YcLfcSkLsPUzSBT6P9VJNM1CnGdtwvk94PFrBh5j
zvLZe/Qe6PBSANbRM3Mnu2zSCzsI0m3s71GbpCLVosfelwteefdcn6W+8WIS7gMTVDvW81NwDbYw
szRJ2O6YK2vYXiYNyqP2OvSMa0WI8krW/33KcA/7lIf7BjdAaylAuMT7PgxxgGH00cFs+oEtUwe9
PcjEP/68s6ldOECWqd9kk/5aC6npwmk4XJ24Le7IjXgSD+d8cUw+LqFmX8jFkxShg7GQhQMl96G3
Jn6W/9KeQv6ckDIJlGxz/LMS6yFFn6pRGVZDb3blFSaGzpL98OfG4QD+uGfuWyazzwjWj9Hz8wI+
Bzwbfca669OAxccYfJQsUsyt11mrRg3gGSU6LeRLSlJU1nKApzHLTCHS219DZAjO+msakixJD2hd
w+X0l84vbLYOwRgXIqf+y7lsBQJB3KGxYJGGyQ5s+DIoW2immKCkEtLKRpoOBZ6zQK8HntZOq6ZM
wzrlOREjhIjDSJ4R8C3WLiCjxCTzhLy44RKKMswrgNIr8Ey9eP4tZtc1e3b50wOhC/DaM0tEvBMD
a9Ma1F3pzkEkNKCvLvHXzSqCX0FNe3nfWosiOxhdQ2JuF+Dbx5YN7sa+YyM4IRrQXyXktgFArozT
sY0dwi8Ob2xz/0jR82Lp1yhqePUvYLaq+TZMuS/y5+SDxVCYkW6jjEbjKJaUeSng1LIYJXOfRYND
54VtJRv8lofYwvbcue7ge+vsEk1E1253sapTyjYaBqFgazFDz7vGH1XKuL+AoQ8sSwAlpmxE4pcH
ISDUFvKiXKPuJ0Qwpg2mvI0Jc8lv3pkHe9JWEUh2jI5zb9l2LoFOQzxMkuaGxWLC9E/tC1VDH48k
Q0iEevTkDKkLPAHsrCGG5eafiACK/qae1ZiJst4wMvdT6HCGerzMaFXNo64Ls57tvtZdToJqmLrO
oLiCh0nU5C3fP7HuLRawIkFAQgdhQgObOFIMRfOuvKZcP/OFzr1tRNOwFQg97D+yYrEDHSB6SAaK
woBRQ5ROFUI7zKiL3HpFnOi/Cohdfl5Vurd3SdswEQy4IKj5f+Ca8EOd+FiEMeU1Xi24ZiB+Zmv6
QiZOg+muZhvhVn21c4KMoOXfDs7GTOzvEI45QBNDu7chjMDVocO2oaSIRH3n/jBYdi2RTmf372ZJ
7T4rzmmXNUmqZRGuRhsa8YhD+A5cr8ihRilMmFAIO8YOmtlc2x5JVTonjA/kGCHfk96zGN90BpqV
+LGfKt5I9FNKz5y/Sv5NgoB5vJlM9znPCcetvZlw59MBl6FVfp6vWLpLkx7YcoGOOiDOYJTYBPpY
hLuBQHSgVItWTdFWSE8zBTyAomC4dzJuet24oj1GUCttpQ/4kewQzITutNEzFW2XOK64dWNFjLK3
HI3u6c+Lq9rBW57URlYdt7b/yUmBSIESVZIkfJO3P04wIHCmuFIJC/UJSJzFYmZ1/Ddd7jfNI+X/
b5mJaRaDVQS4OTef7weCHn0i2ilG5A9srdur85x/A/OATiygRblDxEZAXyE0220y6P0hK8jyGrgs
FIebO9LelKeedw7yN9v5kYbz+myF+a/B6ttT+LIGWChTAJmnyH6jDoxeRXRTTSJ3iRdrzCr3dXSj
UXXNDqITe397bShSZEQt4tAp5Nlsb/51fb+LBfCMBrFkCYhcKm1D/PH4UZH36dlonX9qmL71GeQo
HMdYhvVSVTXWOYQdRvWnpWiyrc+x0smPP8cMOrpgKKpjGETseB5VAXFvqc1cWGt792IshwmuZ622
VFWDSUfxh9W+nGiSNcssD5JUT7L0XBgYbmLB9i70MNt1SpzEkTVUUfzMEmCmmEHXM9kcYngp5ATP
aAXtdk6GgB5bM50Ni8bvLPDyOlXtyntj6uoarWCOvN4WO/LC0GaFjzvsdkgLPTRzxrmbaTvbBUZO
E5lcgZxoP8AkY4XsBTmrGP3imb7hn5qcRX71AJHxoRlxJZPiJjRQMb5TB0M5Hl50hc36U+/ZCh3o
QnHs7/8KU/GY1QTpLpyfxhiw0J1mWsvuGg/XrKKKdXAH06SVAjEfuD/suigM9rBrEmgOQeCULalD
I7/g6669EO8CodDqyKQ0juu4W2wDSRcK5PEZTrMd4lhVTWcaexqb0esVhuXe+1X4BWv2MrAe3Fst
tsDhydV23c61H/9Bmx2NxNwOiCE1ehj/5HIY6KR+CuC7teVwHs97VSzxbadrONMCnzgO/Kzzm3sb
7tz8cTicyxYQtndDAHmi+hg95MsZMgAOHkd0BicEuGcY8URX4ASLVwp7DMZ82n9PHTGHHQ0HK2xn
6BMUiVduefUmlN0y/mBY4AwztUKrJz9XkhgT+2kRbPGwBP0F5d9VNZvGH3h81FXMdFILOn5YqUlJ
TfYDD4d8RNuJb4VgizrWyQ89UPmes657tKNdCnLky8hkqN4Jiy+ZxI6xFzjkkKMTar8T+Do1gH4X
oq/V+5S/Lnxq52uO0+O6Ob1+fOyxjrZBC0kqFpi9R1EcpL/bdorIzYUsc3d5orZYglPI9utT4L3s
3QuRvXxHNHcdfCnjgW/yZlUGPdXr68G/Dnj7vr0KMqN8DWlubGXdezq+qh7jnDSf6T+eGdsr0K46
6ifywCyzjJuvNLbjyIxlhu/jvJd3gUK3LjcjcKBbNkeMWpaBV4m/3SyKWiXBnJPL03+NiqB+hP8m
0DDrAt+Xc20xVUmvi9ukW4AW/VFkFBN09uEXe4nKbGS162R3IDIjJAtqsEZqqBTVXDjSE613nOMJ
0UtfHuvJoow6EqSf3VLHq0zvWtgcvrb/sUwUxkml+iJgEjlZHa2ENrDeA/TFthLrS8bX4Juv6rFA
5UJBsmY0QCfikXW3+tnsJ/w3uosV0gMLH7P5OLULvGxIQsqW8bGIvX4TffuvRxAWEVweaqdIdQkx
VqRXr5QrvjYIwPM+zoeo5Rsvq2zJ6GvjB5Vee0gErXIJLqG1G2cPxnFYj7IeEQUOPbojWYOCBLLo
zPK4X8L/JDl0UEwl3cC2HZE+XbIkqkLCO68wWkLMAlWFmfklvVlVEvvWXEmkNLpidtmzefjK6oB7
qxwBxnT7l7lvMOmxSTqqqXXVzCCG/qA/8ZfcToAKhnpEXb7M1PuvRWEn1ffzeLe7StW/48s/A1zZ
yGTr3uDcAld9l4ZjKSh7TtYL+Z/HLqhLk1mgQiG+7m2sTOw94CAfNvvE2dePlb3OCiU6ltn0tNMV
9nU86+0jlXp3nByjPSKwdX6g1vHJtpd0NfcAZx1HjJYTb4939ZTfrl84Yu99AkL+QVbaE1/ViT2W
cyZMWVv1yNqq7fEAU4ERSoCLLbo1lJhDjfQOS/M8X/96BZ3Xioderp03B3HGQ6QlxU5J4lqY7RXU
bti8F6qD8Tnj7PjNsFNh5hfUZPDVVEGy3hXTASJ4LwUd9AfeNpgjSo7WS1UQERuetZGkV5J4MTl6
bwEB4oZURLXCgirg6op9gyPx4EqmBT0vvuBMH3Vem28pAeds7HGt6ptO6aEDSt+gTYEjkqByeRZO
TrOlzibseAiSmRdkVvECrbBx1ja0MyCEpQ7EaJLzc98V9lwX0UEsdohXBZvJ0R7QgaOHoFyXsWJ6
zOFBQhQnMSQOXvbul/3tmAZ0qunPOpaCczNkBflxCb2bXOcRNKw7XG3xv0/5Lpy4BrtmTVXWPRAS
e5PCgBMGCc0eLl02QIbGPJ21PVfAZwZ5ZHFQma7UAfH0qMdEmt1DLU8DiFPlpfwvFQ5ue0v90YIA
dDaWiIe+ywy2ue2WvNs+TO0D2NLZj2JuaUq9wamfVyVL89VkGo8udaScQKsVsYy2thOfjUK1LgD3
LUgl2jnStfAR2vzsbyvLbM4B1BmTXPXlJ5tXwC0Z2skP3I04ag4UFDsINsThblNo9xRPz1dABk7m
1zHpyps73hFIAI2Ioc3XwcXNV7u7+uN4C5CW4pmsHr6yUIMV4dZ1DtOJV6+uHayn5cQmMOjIi2Z/
0YzT/oeBMgDYAApq9Rn84dz/iiv4NGdMS1UXNIS7WCHqy9OO1/+gXIIMzK+ptN/DbrRg1/XYKIFS
dfN0nST5fgKisIvDRA7Tl5RLUCy3cSvcTPgYLHPH+/VYoKZTrVTlMvXYIateol5XFbUknJXXA4qA
3VgARhJ9kAuDeykpR3WL8wkZezVcjrT8zXENpUkepZW+VMY1EyfC6pv7Xi78rnhdXv8GEKiIOXqw
bDk2inE/Ehy6EvKRFXABpqhsCwxciOe8dNpWbn2SuvO3kajOBwo6mPi2w697pys1Yi6hzfncl2O1
lI+A0YL5X4t2TaH18ESy0L7URJzDc3T2qDHmzdL/TriJkBxL3cyGEcTJiJSuXExIkPfQ9Fw/2GoS
wmUeLytRn9zUzhy0TQRbouKRnTYWoS+IqkYAD0YCcWEJTlvJddsDwoVNdHoFFD8d751zcyzJYgqw
sV3x4pyLazM7uto/T7GksEXhRYCYu9iMrtGCnjvafPB1q9QVmIuqGX9TZPzwYuALtorLfb2WpNwq
wmPXUF2/OGG1tG7/sBaNd/3PrBs9029xB3WMQlhcACdJROYy1T2BVOP4e1/sE2KZrSUyVkERK05+
m6jZkedOT8ThVI2L9uNiPVXtOrt4k65VikVtMR1LoRfdN8CuE1iIOVuRBIoOAaiL9k+B0vzv+Atv
OfAJ4tS/5lrcHR7wZL0LwYZhLcieV+2hfxB2kQ7RNReaYrGZdla5tL5a1essb73Wb+/v+cgo4Kax
v/thhy9fe8hD9M69RXWxOU+Kpb7pwCusqMwWh8Ojw+My+SnP9U61AifRI9aLZPrCnk/pTAGqpxpT
L2BGuLLUSgh6UbK1GQsq2dcKPCCa8as98z62vCeXuXbhTpTAMbN3TzqLB3Xt9vvbHpIGZ/TJ8xEE
wn9WiiD7vVGqCLfTaI6qTzTPmUswmFSgWWsb+vYXZkd8b4cftvznw/zz6Z749Q0KLhMezUhPFxJW
pmMkh9cJhpzmfQJ6X8ow/mM+19/J+rN9XsHrhbI7hOVONv9OwvrWxxHy4YicifFuxE5OfLIzsFP5
s9TrtLRftr4rAQwOBlayizLGBSiBt8ZHZH3jO8e96sQaQjElnuRpX7YZOJumMXcfiZeXHlSAJX5Z
PSXGIYBWkj6ZN+agMqZbmCiqaZl4Hfj0FMzydGdQI2xOafDwYDPQqGJlbLNS3Djrfjs7tCqX/8Yd
L2y0DPAQd+fp3KsBhCXmd5Q2guEFVrN2E4/y+cVWEZ8t8zfpM8FMsCRpuGu7NEoqYh2egrWpLnT5
59XHFhdBfHaXe6ZPw3vakqIaZPugcN93BTiQvj30GGF1N0fxfASO+MMmhSryboJjucubfvBDhw5m
GHuk/XzuQ1GdiKlx2P+hu4p7b3eOisBwbcCpCPRs7Ial/7aolPJLcT51WU5sDqz4gje4ULxIzByA
irG9ZtJNFcfau7e9LwYt5HXBOV4PAm6pRNjeJE488k4TfUFlaWTxe8ebm0vA0g2FHHozhiWn1EYq
70ubKnCfjXI7qbHka4SUvvLwMIMk6RQx1xGHCSRHpq8HYlddf4iWbp7kJrLW6zKPZxk1A2wPqBjF
aeOl6kCrkLaBp38M52gSg4Ln+FJl6rGo+augOMaGjWsnMsEJS0+jdsMsZF6kfSmqlxmWLqEAHJND
rCe2yLd66vqbKos+E3s44iyAYASNm+y8d+8KJzl8W4cVYr5JcjoGjOOCueK+z8OnxubbL5Rcgaln
WnBiBYej9tJmBHgKNifQiTd8/RzejWMztFTMVzXVuck5nLrVJUuUvXUlO6NUHU+v/nG0y7HQ4a4G
hePeBbdT9i3tdMO4vmg0CxVJovybPbfnxZVUF4Hn+qVuPdTdgo0/y8FcWNENs0BWKNspfXnzgxir
bb6mL+2ftjwQhLh1q4PBppZzdBJC30ZSc08snNrNGSRKXhdTxeW6nwZdLtfT/u5vM70Ms6XGIu2e
HAlNIhsEsanhx35WcYJFcpnyKIcOuw2NYTg5AKuSj9GZ4sC/p0uZ+p17CRC+uzfLIoU4wXiioA54
LJDHE5nkj2Zr/J7KTIZaX8bR8mSdJweoVcrD+UMqXhHD/wNFAvnnOF6/qg6Ni6DsC6yWoECxIafz
pfq12cpnVpDZS70TX8N1l+QJsA4BQCz0ACmm/rFDvZIRhAQbMscCHIgKIKkt43e2QzhUhlCkXJJB
bYEhE888izOEjLjclEW2LBGVVmz9yORxeNcm9uJj6k+8MMcEO8Bv7noiT9YGid1JNRhNoRiB420t
IzVhHXs/LbspCxGw89PmgdpHHW3zU09PAdsGqsj70hwKre8KT+fWmgj6tEPCWwL4oQJ2LnSoDiXp
qg9n5ShGYOWlQIRsUVdeRJQGNr/gwSyeY37Ku260P5Mpek5B4dBKGoNUcWpzxl5BfcW2kPx1PGfU
wISuzXFW6ivh7HVIldZI4v+TrksGu68bQ5YVBPhkXrwpUZKRPTw5LBzRwtTPptLVhZddj9/TvFv4
xavEeaqZ7fc+KNUb94LvT04CLxa9dbWLn1bn4g+hNQqrJOx4v2EtHNbuuqB0IycDAZf8zRzeUdME
nw+m7IAkfumllcSynziCVZJ58Sjc/8NU+UrtlUW3dTnBLgOTxIuJdKT7vOZU+0mvylfrQNtSTGIT
ZU9kNutDqXod451z4eRY6R1qO7IROfDSlosnleWE1MetQvqJ/TCfmLdLED+nbiL41kyDqF8ZxCm9
kak+dVlNxvcu0gAdWKxzPoO9V+ktni22xvXhHSBipKii3QDAMLy81kxg3pwuYm95aC8WNX5UC+H1
kiDM4G/ZFdDIjJDeJBqbpjwa9ghscAcXrYbV9kVjI1lp77A00bHnDfl3IP6cmP3hdnxuGiM4GXD9
GSiTeCLLyQivLnDjvaSY2LkB1dAILyJ1efSyYOcZ3LSEVMfhyT03etqqsEL8Akw3qq75Zs/dfsn+
2cDtdZHIzgfgtCvcWsLxpsw1HQiTLYI3zTLi8V8TKdqFIho1df7l1jFplTns8gajmts1rHWOr0NX
rDAn7ogDznf/nkf53HFDvQXfehaOawamgvar3KvhBMh+H7yKCiHWrjpNSY+KIYTr7EidESdMJJwE
U8CJp1Zmyl/KigYXm+9zNeZraTr+hrlAA6M4NIJJLFLGd+shrUdh3SS5T2IfagLIUtbPknGoUKtG
xQXAW2pKgR8scYWCQG74gnCHZwRj48favkxTbcg4cGFuLyrHfLytO6MJAsapbn0B0LWk2NQXszYE
Hoa6gwNIygnOM0TmW5Wk2o9Xir1yIr+2ruhxC4o69rAKkxm/B/goB2+yahR9jhfVCubmTF4TZk/n
YOQV3riSDAfNUlLJ95YLVIYDehKlSkIA4vHPTmjEz27TToMIt9wkrAKdfjUiApJiYWrnzmGfudRe
QA254L9DIzH1RqmoepnQiGFCZ5F3m9OYsVyRKGowbH+5ipReliZsWtSrQXih2tngehzt3me9rqWi
fAmG4Hy0PMi2YdPzGJTb6LMocQ4T32k52Vr9/0jrrWSdJWmJXR16gLo9KtPBdLm6ra4TvCCpKseJ
J4516k0PE/RIWevPt+rUx8DcJWf6xAY+4aLS59cxNMqHFR8bN7hHmVNVFsFYc9qaRTLb7GunZC+B
ImpOwUGMK5XctAdaY1y7PxCOt0eL1kegFbPG9lWyyuIfQnbOoFffgGj3Qq/UF8Pi1Rhm9i4p/aBe
o+wg2DL0uYA+bzpKdFEwbtM3BcCIif27kshApXSRi6xsyhSB5x0vZOjFAa50v1DGlDHF2LKp9Qv1
/OtA40NGwzNj1OSM18Ou84zVr3MTWkPleutQXXaHqsfID3w9ZJMx2RRszZtqvVK/GSJERm6bh2ta
0E07wyorrl7aaZ7ND7GlIEU8OOlCiif5qsoqJFYNkafxBxwH6fJtkcoiq5F/OhoIHpfWFqnEMes+
UhW3rVJpxmaDDkDU/s3Bgpnz4kQLxiocLyblKT9VP8qHg8Xdq3SSFhAJsa+1b6HHM2Af1mzhhop/
brXfajrB1DgIoZG0EwkILp3xX2D221YT7ujYp6HwlzGK6WdLaTobyTdE1i+a4yScJgTs+9EUAKpU
QQBppKQmJxTtTQnz4BxbLT5qbgC6TDb6OaNWDro+CMdEL3MS7AxK6/QzlyYljsmVUcg2d+dyXpUB
GaCzhRmTnpuxDgyLITTAHR/k9nprbBdgqLdoObMluI/XQg0CTgoTfdsTE8bTzmj/Pkyg+a+4bzVW
N5bJw+BYu0jUgt+qCioql17kcB9Hs56Ik+Tpek9zMdYFfF6daZurd12v9orlOuEGk4vk7R0/ZUZ8
YwgOp78qhXSFi31Ot4nq1UUe8xZ6eeQd/eMNO1HFNBSHZuhVB++Tqb7eMB1gS+j15sgKqUz52YnU
Gtn0P45WsjnJfDavJjM11nBfmgvklZxxudf4E4JQmqnVPO0Eh4OrK9bw97H/CuEsX7yYhBXvbtJq
I5oKQz7gKBI4lEIDlorxpC4muxN9fuRRlZZwwdjfcbvIil5yu68Uppxo3GTxFYy9ivrSkTXNR3Su
VhtREF01Y8u+x6HBZgInwwuauwzPjUxiedwB3DzU+o1MNdmWNWjdR+vkcXiK+9BKfLmQTIREjYvp
1IrhUBpJ5WzUmJA7QT1lAgPN8HhQlutL/V3Wth/NA1kKgY/CObuXRjYvdwm9LU/kWTX9Us01WTKI
nPqukDH77X4wyzPtmv4bBnCO+93nSZ7KUc1plnP3PJDEwPTO+RlUxExPU3cEg6129fxKZ8Vu7JeE
muQnact1PDeMo9fn7SfKgaHmSi2YhoMSiTSwF4+3WLi+hjVsxzmUv1rruP+Q9izd6jYOWat3rs5g
AsWvNLSaK+VDINm4wh2+MBuogpXUueDtOhNb/qWwE8N3rxFA0BGBKN8adMviHHK6kdX2AdLccwsJ
IPJw2dJ3d7XQmhk+XiL4SXPRTT1y4kHjDblhh+LanthN8cNjRMHpYZcsAAG5XXo9CLeMi3hCCMVt
R4MXN03zLndTQ0HAtha/5dYxyBSlNN5adi7L29FwDbAydx8NIIcsn0JNjVaBUYZf8upE+hvMZvqC
C6TyRZVc9oWVBpAO6d4DwQuUfaeRzwRU6Pc/pYFoM0V2gGNy/iitcknPbsnG7RrSUjjyUb9WTOGz
UWa2fLZzInnySTCKmmUCCJffK7Ypfz/xq3ovxMU4/5EzxHwQH5fXhYhS5EOz/6MR6kLoIXFpBeT4
cmtyZ1yThnu9tR1ozUEFd5iyhNYaCKjeVcDiGl+EU15SJcjn9pJI6GIoztJho5AF69yPUdJPHOLL
1Dv9ZUrTxlSeifirhkh8fh/C1PQr3Ef7s02u+m3YNcBR9/dYqRxi4S04k7ML/NQiMHHxckFbs6Y4
BdyIIJ9clBjaZERAvdPA9JKUHu6lusduW9QBYhmZ1m9WH70hXjl47D6y9cg63+DMoOOF8XDE/NOv
kcwbMcGJ+722Osdof1Q2fzqVp/1CK4JBei5JAlL96MYIMhzCc6m/yc1dywmK25Hv5Lek8SrRYhZC
XVmNyVioBgHoGAAbsntNPON6cJomlmWoPfhwEiU273IsAU1oLgEzTjfboOpdh+Vzzg1ersDYyWHr
+NRmKspaAPwIF71AHG1pXsJTqZ9byDSelMtH4RK3bmjeo8UG1A2grhgY3oya+LzNok+LENDch0RT
hbXFAEnqozb1c1haOCXniSe7nmHGVWTY/X8dn9M0JFT/yWKSqIVQcZwS1j5Rp1hoItCVRlcwmWNC
CaaJC+BTaYysoxyugNmVcOoLlad8F4OYRi0t50F2HNltEIPClt/jfAZSeECq1aSydVWfltZ49xJ4
t9lClDbsiKcrMRWcj+Tjs4tT9GmlVaegftzK4ZbxsLfNJORdr0+loPqzldtEYjyiStdqibLl1nQD
Lv9BL6OyY4BXkdzde+A9XjrhjvKMT1y0e7h54j35MLWGWrPOCvKIjDKQBkqe1RFONVOTaMj0VN/f
NZXdHaMpYjhKM/1/Pgvy0sSNjdQZnRoJaH9mkYmsu8yeg5Owpc9WbkaN5YEtVsEUUzruPAyNpW2n
4EJMx4c58poE45LCeGPHtAcSTk19SmA1nFo0KL3695+ee4ULoGiEZjvOrhqV42Gh3QDNERAgCbZK
z6vwuGNEQoDPo/MHReoZqJ6ZPbiwDZ80ZU1CO58z9HCUctQpoS3bGwTeh+xRbrGBNAAIh54P2V3w
6oyPHsT95htar1AtcghHTj82cgldUAdWkaQD6sE8FjNpYVjAwncKoOF6RDDBEBOn3irw+BOxpbZi
DznTiQ4FvpjbFGZtagDXjlb8N0dxLIJSBAirBs+y0891XApDo88GD2QPuTK0xTFKbuHOls9esWly
SVjZrAkqhGjl3nEbSgcIrbAUE2cnyCLVwXREeZp9P/g2bXGKV8oGaRQ0Nc0uZGlGCVO1ZITZxJXN
LSzPb6Z/KRX7ShOa08sck0WHHOuCABQdRkeVjFdYjPdpJ14+NtyvialnIAH2d7Dz/+xWFY9i6+xA
vtJLHe+hAUVm3XX0Vg39AnV0e9k+XchNKAcxOYT9nyfXRpAL3Z7zDp0FWpGXuZmmMlx49wzq3VzF
fycI1tNNqE9j1diNlIO2/GGOdNjXTPHMJDAdmHpxcwV76jjbW6fuhMKEdlQHs0h/BCoVexZNGuM3
F8RGx/lWPJtL5IsFH+ZSh+s1+Oh/IuWpWusMm41j8f8eujEaX+vVs0MCcl0GNhMGSktQPpCjQ7Ov
wLwcw0JDFpdXoUrK7aaxWQ7gfhEp56h5gematz3lQAD4pfCNlh9XYos5/HG/uVebuI+0LdFak8FA
6BYcoPaUmR1Fb3rGIMV+hVFtXFt0jnaLKyM9rSxBCDZLVxkXyCD66wDg8MVIeWnMmtbhK869EW4k
9J76pdQiS5JYJtgJsk5+P7j1Pci+4O7YUIE6tOEdG63ZQ3oTGOqBdzqSNrBOF1OXzc/d4kvbqxg8
/hx1+7eXQyEB8rAKnhbdzN5uF+rcfxB5kqcFSUiaSjzI9tf9iudfOCmCnzXpoLqVx5TOfiXjOk1T
O+0Zziug+xHxSjKVnJOzKg34kF0TR9ovhhfry0g9myssbnRT7CZ/DJBUvRH9/oPF8pasFuiHkrA+
efUo7CRO23Tr1+Iic15A4sHWLZZ1WaOHguPq7s6GmTcR+mNgd5Js21/bRKRmtriV3w85G65AmvGi
+xirzwsNGaEQJP1zrj+JsDziUjCzyy00h57rmT4fY1RbCcWLM01Va+PbsHPRo+jWHgDxk3JWxNVM
nCEFh39xL5Ner8jM5QuFI271hMzwxGEaia0NXXM+TIU9o7qMCP4WgPVkCIVb3DS3zlE7a0jrbk5J
rzrmQMdjXhkhZNPEJMVBZpqBkZIofiWhH93shOaTdvGCGN1Z48VZ7JjwZv5iCeI/BzZ9xtl6hyLc
ZNxTmXwcRmSfYGY3PP2JHVUqyJG9HD+SLfHQllLxPW7gnlE7DlMO683YqFvIr8LJB4AX5SAsanXM
c2FmbR2RVG0V4dH0d5rJKwQ+CklC/82d0vPvyUWZBF8vj0EJwuIpjrv8s3RvhgPyn2SAI2040b5V
Urds4/CzntQWw6+vUSv/YC9Hy3rS4KMDT1ohH75R51/bUId/Hz2sE/yTF8ZUC1pENPtbEYQNPst7
BChUoNDLIIFVpXdzE3vhdrlCoMs4DNSvlUVUU9Qc40ebEsKJDhtyf0OO/ioDqrDtCaD2aHq5wzma
hhMusQeHcgFrSsBALf+HuWsUOduAd2yGB1CYyt3QGzdkkm3/Snphoa8PxOjaWFnJujtNmqm22djN
6ibubBqer0an50i0lB1pqdX5Ws8hNZAJ5Vood7CK7R8lGCkcr16e119gmJJWjRmYgn/M6QE++Bsb
BYNuj/Z9O4Y7bcaSrD1Q4+7X9UaV7HTzRM47RcQGLKTZimxwsXfw/YoMTE9/58AIrhXbclIQ7Sxp
Z/igx6ox6XVVUNeGHXiThfuNZx/1GYuRdGSDWzDfKlaeAe3gYCvWcxH0sMobsBqna6YUFw7ZJfJ7
IFE5C5ubGcY8BbnUvtx1oICmjYuN2Jp3aYMDvL4Nx/qgYbU9fy0Wd5605P2nBAxevq5RLkVnGgxk
3nVW3AkDpNTM7lC3ToW2enyfdsMc4HrNHmDkadBsDR9oOHw49oqWvj47nFgFtcfRfAcdTkd1DUon
6jHsTT+QQPQF4lX7JjxiWykb9diJcnW2fUk7L1A03K7OFOxPdml1+QN8idcMVL3seKDeGXbFobYH
4Ts3SdkeIp3vpoSBKYs0P9a34MyhvQ8YAWePa1m97PT+mzusR8e4UY4iiXRKQop2urlFMeXCUaH1
5HU0myZ4o7Xt6zc6RP4N6ZSkdU0FYQIOZwuteCGBZbuKwj6L/Qcm7+uMZMfh3MrQgxLYdInQNW5A
0H2Hx7BVXEqFxC/QUx8Onv8EwOsK2InOYvaarkICS9rrxSFrBNl+3FtElk/+1uxKBeNpDsyaWxHZ
ByNwqyQB9mpzJ7Dn650CJAsJ3yDSEhwPPiNQgT5VhBhBGVhMtluXf6s/rsdTxD64mQMZOUWh5ijC
nddMuPvCm6kQTWLU1A72iKsugxhwDNVpwboMtO9woxyccuvHRzoQdXhRK5xhE9sUf5QXYb8tM79S
PLFYPiLZPjvVq5MX+cZZcZfcz/8yFBsfRbZLgM7VMslsYOUW+NdhDUsLbeyEFuvmsGgLbKwX3pNX
J2KWQhYIybosiKMJdGacfXe4lpui/3jr5v3xi6E1r38SNN6mhRaIbr2cxo31W1uiATwYUdl79w1+
wl75cr/yKNtWpaVGrx4zAKq3gA6Sne3tdhVGhOCl37QCwhbrXRavWcAHep9KgQX+xf4kQxp82GCy
z2FXsEHBuioTtp+8OTXuDjvypJL+hSIg5gz7ZSU3sbxsEoNhY6ncFFtr4Wg6CD7WRCC6ffys3s4z
JS7XQfZpwVB7LE/Wi2Mh7DF0sXnzPB9ibeOYuze/x2V8wJdTw6BUEGalU+g8Vic7bwkBz0frXcTt
kULkIKWuHLYH7evrUXCJ4MKnekVwW6EkfcksYAj7D8qr+u+4hVPANhkXHB1DbyAqPcCp07KKl4v1
qodoblTadXbugbm3nBEexWTzxJ1av7+S2GcCsTQ8KBoEhIC0/f/Fua8xMS6V+3TEtobEnISWyYvB
Skd1OYhsosrs0Wl3pSMkrG/OsyTfk8zfp7DNAl4roh0L2vUqJOcYNfkn6lWuTrlLdlAhAMoPsVOq
6y/pVC1w1APfyBxNekbkjcUnLDibXArhVdUYhOUjoFhJ3z6O0MBHHc5CxF7P9XnJNehCWUppX8Qs
IG8t8qp3V+T/rA5BnAZj722cuujWwV+/xtxg5eIRJPzumMRURiOGMvg+cKXaip+WLMjUfV1bGXrA
Y3xee1Ooe5ThQrwN+4ekGMueqinSGD+HSHXb4LrvJ5BCSoTgN8deaUZI/QDBbQP04vvyXf3gEAze
NCoLKjEB6eo3vdkju1FjPMk0KCOS6Ti0tgRcpiOjJbSzS2sxGFg48P5HenZspPwoDikxfIexJKYA
OaJ/4fQCikr8/WK0HLwSRHuwjL37MpUfh6MlrOTN9MuAbNLqQzhU3D39bcTDP5efgu24OcA01s8V
8g66FpqbWonRB8XtwbYPSjGtDvt2BAymeEAkWPavX5kkmLK7h2lTR07kOGvVhVZkYja9i4Q70gKf
FVJOQLQaPCtFnNlpEsIcxsC66bO8IdZ7Iv7nbENkgft1zyh/3asrOPWrARKe/PzWA3v17ePClD6J
s7LdL5eaGZSFd3Ybus1RLwlGBOTqtf4eJV6wc9BfRJsObRieAQikbEWnZAQ59kiuRjiv9f8Y+54b
mhrZVOUz5Y9onj/fgtIiWwrSZUtIGc0qp0LzSB7ka+rm7TmHaDVHzUhXurGVQ8MleqpVxsujmhsu
OUfRJTSC35lfHc+xCA9+IP+y0q2rzwBXFCt+EHqcIZrxIMzbdgB+JESGvKUKOt05weJoERkocHd6
2MCjpiOIW35T8N00o3l3fVFlC15yHnfN3Ll6TpV540ya8F9afaiXQJAQztX5gifwZfUIWgpyX1O9
eW+h4WiHrrZcpWC0aKjy8osm90u/vuvGTR2QQ4LER6ZuPXB7xlsJMhI3l156KGOQ7twFv4gRaMqV
mvIc9vS/T3PraXI/zv2GuARGyFYrgVz6gGNVIHmNMfTgdthjQ28BkcwncWmhipVcS9ZOknrri1qe
dTSt/+a32KMO3hrgB40uV39iz7C1vnGeimbisubqE8beSRCXvhO3jNHVEazHxY70fVF/w35kzi7d
pfIOXF8uYt455de2nKQFz2tU8C6rW2cXLGih0/wmSmknWU5MivBBcFevpTwnFPshKOt66VecqQvo
Qxv4/4JDEQwsAOyFkbvGpt6XyFX1NgtiUdbVFuh37EtWp8OxxmK16F++swXmQd9cTEM2s0YuQ7Xd
LQgdgp2A1Q807+d6SpPwDOz/YOAPwf0EPO0MRGCeCNCygVqb3vRV0LcSCNwOWj0b8M31kjxG1mql
WV8pMtcwshJUqMZt6Wm5PYrBOz88+iB/R9r7DFcdDFfLXt0X37wT7g1+Cdrn6Kcld2tfKFZBgmif
NRIWNL+PzBYaalQyn8NbPv94OEqEXQuqJcDz+WI81TXt8RPbsuikJx8ThhjAtSpncxIG0APdpPyW
gmzzrA1sH/IfPNgO20aHPbjqtTQqTFzbeczb7BWDd07cgUK795/DoXjbVFK2aGw26ni84HRb05z8
dJrsPJRzgFUwhJ7rshhUYAfNEzp5Gg+bPb4uT/P3iOqL+xB6KxscpOH22H3XvdhSx/QVmDSDKe6m
Jmx0znz2x4KWt03sSpJ9IiiejRdkWHDWnDecK7GBtcI7Aj7TDl+t5xxpbr178duW64U2NjnoeG+C
JHah4ephN8S546Rl94NYiFhALVrSkJBjZX7h+cn7YtJwQZ/+EVQaG26PMDG7Cfs9hWHZQ5BtzELz
cXO0ZG/mpcTufal6X/XaBMPHQINF1kgdIIAQumZQcob+xmtEfyEpBRyTxrcP1PNZ1VlCpm51F7EA
SYrXofFr5El9spgxnG/n+7J+6vw1x9mw5ckzC8L0Tg/Mt+rSnXNpXDVIrwBftp0PKN8cgEV5/Rfq
VhidVPvgAPJOccUCP4tKSvJj/zA2UnkdRy4mLbldsYjMDiCcGLdAAb6mPDoWLdyIUCMce52qdMAD
pL9/RO3H/M3NbFb/LaLsnz7j2vf8lt5KKF0uk5TGWNClLOR6J4MjZIFF19SjxAuDj84L4ma+Crgq
azTOOJL86ZmPfpbH1ACSPaedZcdVzUILawwkHG8qLypsyhb+1OkNypNCgrlLJ9qGubP6KFLig93I
DUxeCnsXWZ78zn7ld+lFlAAbn6b1JKdtCb+IKV3nTdjvW3S6IN2fnNJzDcAyk7/rdzpe8jkvSNGX
0YrYtqXq6ldwUd/bUlhGtjCrzs9Tp6+4X0uwCzay+gkG68Uci5+414IQqAgFcrTDMGcbFCwCquQo
Om4h7iT8rd0EFSAPR9UUKEqTq8W8vb/Txwc8huJ6O7rWC8h/LQ2bj6VqCJI4PqpsJNn9ZrZ+kEI/
IMekxWo9xon8MeFEDUBX6Bh/xzdr1phnwQn0MBW+sQI5lkOYLYWKj+X5iVKU1Y/hGURyYVIi+8Mz
wSyuHf79j424yjLDS4N3IuOfzMlnnAfbiLTAn+9P9JTcUdWadBvDNMKQKnQGcrtWTaaO1WCjSz1G
E4wq0qrp6aHF1wrfrGAhWmmQyUFvzAQQyQs6A3Rzefv3TbmsA7ig3aAikcP6O5jPlCs3XLIx5uoF
06EGWPV2u8xdRydRmFqx7fNm7hFmUoIOa/4W0JhAEUR4xRaxv2fekoKYHl/wRFaZokM5ReJOV+a7
+uE3hX/a+DYX0hHmXEf3zJSSuD1e8RelVL0DFfxBsu4YkMC5gwTSPJorRfTcPNbBhkThpX2BgWpM
AdiWnYOrMPD+Ltr2bJ5OrsJBzidtiFU+mYxW3swQccRxvuDz95CCv3n0ONK6EuWmQ87Zs2tekMeO
j/fMz4GKWh26G9v6w65DxrRz6KBc9kOyjxnWoGhFNBFvkN3blOKrF+TGhbjU6T+gglTqRTfwyjZC
KlFIBHoPynrYRJHPag4i0WWBE022ahWIfiHWU0Whl644WvLV3t7pFHoJLD57WJZMUVtbJT4F0ypK
MTyNtu2qoz/310YhDjswL1Gv6jbggj3kGcqRuFOTbEQqs4gX+nUY5Iks0BvKMCGnv4XvOe4lEGul
+cBdFl9QbCynpD5II0XlZENVF/LdyXHjhEIMa0xJljhgC8CTcUgZBiIARe9VPZMZnhOExraPPFpX
m3Y0TqjDil330vwo3rEl/JOoVmxuizXBQJWNg4z0itw2xGPenV7M5XU+A6SwrARqZIvSXLb6p2ak
mq6spGcSby4FcppZNw8aCW2HBoM2TMZaDf43rtrxkiOm26vx/EICfL9p1lht1F/dWrHyy1Yb4eev
fw5Y39KKYG5jUDOBJNg5ITDG6ojed0g0sffSJNsCFA7x9R1X6WnF5r6FwAI3/T3QvwkgHBuyd+6k
DyFq9yycKTgy298DjIFPeuBLa8QFCX3NHH1lixJDSw6QfS/64rLb/8B0VYP/Yal6B6+SXVLyeglj
H7+0bC55DfYGf8GASRI39Em+5C/jPJZiw9nsOCHl8BFYtSM54qDH4fcIxwIvroxNTGRp1K+Zs/yr
GJJWJElAYFWtdilXQvjNBqg8PdMCQ+hJtu3O0sUPo0MG2zfN8ULbmfhb/krf8YCsfI2oQstBtJwG
xyD1dKIoqVMCFk1F5+b/yTwXZT7Q8xnoM+9u3G6xrUleErssBVcNNMzUFj6Nh9o+w6gCrkSIQuWQ
R44NatAo9VjVNBsYO3j6w6yYEg0f5sDccV4EJ/4+jtkpCEJ0CYUEFbp7iLQBEFUMr5Od0bzBZQwL
qlxSHkA4U9sWxAx2sqxBf0wlwS/CG1GD7nfjza7ClQjnKxmaqTt/4i4wvYToUTwUAMAsH9J2C/Xo
4d4Xqs+3zwPEi0GP2qKY3cQ0BC5wKCD+ybOqYFA69NRaHQPL/hJFbswhAHN8JcRRCdPruC8EhegR
16L4YdsU994GzavmRGsZxPfgTERH8ANG33qJ6ChfPNAIZ5XZwc8Rng2uimRZwjSLEapQUiVqwYdw
5xQtc4IuwZPsmYMRVKrv7gYGyHNWGewXkXRiZE9Rq8xe6GMOnEkp531OpS5nAKhdDogwes+2b6WL
LcPBrZq2ACD6G3f72GM0rMdfxembUsF2pZsFm7/fEWvQpRWaLLYCg26Ge8Zu3eFSY1Tsk+PdxALR
m5ADkuGGXwmxdFvUDjGwqeU2EbDe/6Z0D9F8GvhsbRgfLAsBi0hhpea/7V3TG5bv4Jmp5K4utkA2
WUsM07KuIXeFyI4hXUocVu4FvQZatqxSoM7RfO18K/z7TnZT0EOdsdsh/1TRhUI/ohdpdqEceUFX
0iTNGiSnVs0YIIFvPNBDWym+hv4DGcf5g2RY52lfdMTVkK30sYGbOBnn6lsCwsNi8IcD/c77AZpu
CUV/yDIc3x1rGtOv513fcmllLAdlbnZyLixRRnkiIqftiXhZmt7bdygLkv1Uo0HO46fOQ2uAKeUu
DkEquVqwyTPgWeNFv8W8+OEHAQMialSzyXzTUGgv48rh8NprfxkMmzA/lauu3+MPUmhtpzyc4hoM
Cu0cSK3KK8U8soYmGb4unXx1oCCjBv9pedzdD8UHSPHolUWH3eeLTz0t+nzpgYeD2yTjwjUkDqK0
BV1E3Wzy5Piy5rnxZSCQ+q2CYKjBhpvh/APWOn6l21zKcklgB5h9a6o9+sPj7FFr+lhJrEtCxlg2
thP6fwDZ1rtyR6BdAkg+4sgTQex4lokBWD7h8N3PUi12iePX5ZGme+C2v7GYwL/hd8AS2I0pCjvo
C4EXzaZmAJ/s5i1cG4RyyWCc9Ia6IA+Q7qHwxsMLrqNVaB+EC2SXBdTBSH4Ma0/lP87l6r2I6IBl
KYR6ISuJR74oG7RI4N+w9sKT1EwQKJQQ+jux5fqFgWf+Y8ty/1ZCrWlWy47/DyEItfhhpZPofw5a
X8avkbJBLagWXOf39x7dow6El0ub/HlPmxeVB/aNTtdRU8on9LY0HAGRVlOYfeqyuWUsY+hDSwFe
lUKt/Lg0VF134aK6WphBFTX0GsQOkxWR/nvCGcsBbbm7/pwaN+osKp3nOdHXylMSh3x49jRZxurj
gLS+b/nGrxBZYlW6BDeYK2EKhgFIS9jfhrGtJrCmQbs74c9NSy0EqOqilAtNSp3MvtpNghW8pvS4
qJVrm9wKmHKL+3QPcfp5sbdtg+4uv34XCidHRtu99Z4/IOLgv7vbMiMgG7Y7LRcLedWhrdm18gWq
L52dODSqmj+CWBhvLSBvO2MQUMtzxoSMy0HQ3gy1XaMmZOVfR0cK6ZMJ408zl97j71zvWcON126r
/DLuy69CeCiVCB7muMY8T1rFWWAdGmjB23ltMV5MmChtDZ8TcciotMc7g+c1ChFQFR3m7jq8Sd94
XqI+w3Xsolf2I9hF6YYEBlv2bum6byYX4S7Q5UqNytACl4EEOvCsTmAWmZtgmr9PfDmhIiHAgPPu
ME39ENSwZfBJyg0bBI2KzZ9LvXHF1/cUqDJrZBoHZVMlmPZzhtFi14Jbv4fa4J/2jSgc8qOdrAOt
N/g3XaWDt7XspO8iUnU2+iUaZmBLCB43jf3aafZCIOEP0zjA6+59CURZiy/GCQ2tSydWfiraC3OB
2ebYp6i64LSyiSgaXwenPkUjj1xZelRXzg//ecXAFUcnhnk1Uqj+VsBsWCSlcnVW7mcufyMqrrLh
jG2X4wYbQl4UmMaSlwG5EljlbZpiKVf6eZGUw3akB4xbo2VpL55EcyX6lbb/tLRsyNMugpIIP2vP
EuMyxxdGLs9M5wcsi7iCet6Aj1lUEZjcuyT6Ll0NKmamVsE/joiXUeZaE5mHuWMbI2SgkR9OU/7I
UgSXqtrFtSYQg3SM0shWzWAPakuX0BRR3pEe49VYRI3oY3fkqtRPMPpWcbRbvKNJvS7n9tCShn08
1Qd0ZlB4p1/LQ10pKU4zqSyLSEZkVL2dVM16ggMOUB9XqMj/xK/iPfLGIC6f2/DvlinnaNCnoVzv
vngR3qxwwqV3BrVVC/zgP5AqWtFFI1uX71CUbsiL38vyABfvLJaPIuModqTGf6yC/pC1Wk1IOMoh
QosMXSs/VD0P3hOjoKa45JhM07ZH4+7ISSQmUp25K32pNRS7nuUgFlchpZGeJdh4qwVcJBMYd+rI
HLTMWSc68PAuksoe20n9aPUEB/p8QhgaFisZbjMLAOhs65Q4ipxb+fYmoD7BXKEfdL/H5VHU8R8Z
2fd1LprAfrjVJZpf9IOWI6/viwSa96k0zWu1//WD4I2owgIp+7Ktlks7zLah2J9d6AC04aB2x7Mw
clbDoKTtE+DgqAwXF/x+kF/CcaMVmomkDU4QsSRdxgBPUzIkvmOtqlp7A/oUnIINHCHFSu5d5dNN
qtiH1/wTOVbEnxOU44JiBXliDWau8f4JnoX3FoVGLodtIJP65g+6OafjtRkb4+NWginAnB/S5WLB
0bK8AcQyNjIiZ2MNwuLakiYR+dJIJPPFI3tH/r4gtQpsxedUSZN+QQERPwrlR8ImhnUfRKgbx3c9
+GjNdVjCPqC1tuVFmLCaW+vdF4a3ift3Baxxa+jrrI8G1/uNzDhwNcNgGT/4uPNh+JvbkW0yDHdf
WOKEK3qzQEihdt1akuYmMl2KNSsU6cTJ+iiJO/I/Ak+cxhJEnAfJfsBH2fPGO1D4aEDTZ4pYTxGj
0arD2oBNxrdBw0hUMOD1l7TVl5KWvdrZRsKqXyeOmGc1xnpxkdixHQO4K/goZpeSSxHGs75f+4+W
p0uwiIchnxhEvla6UixkC2oc45n0c6PoEu6TIirxGjScNNPy6X4WXdI7yuWLBnF6/nD4NVUPMrFq
DcsBZiG5+2rIjYjGhw2TqEG2bdLR58MnKJuv1gE7HAa2PliBB6YZG218qZhsA8sDaWw82t2A/Dxk
lKhWR9JmoyFczMNVhnqo8yhevvMWdrnCKjTvW+uwN3ix9+CkwX5X3yS9QvdIM+e/hhfidYQEXpAN
ctizks9OML3Z8h2zLvhL4z4jc25Mvmtuh1aR5V3JhRdDbOxSVHFDjWjlSUgVD94wcTUwQ2xhBY2j
XFZSc96Gg5fK92Cf9PeVc7JjikS1VonzId9c9bd2DzxGjacVM4e4+OHsbCn4+27cxjfsfkP/eJhn
VLL2iLOhvfjJ3IPbVefsblzfMUG6jM2zbRaxHykWgsYV6LgApZK1r+G8aE1y6k5q2UzY922jQnG/
qN6TMWNSVgGaxlfGDzQOfrgSoCoKCoTR9Do5q+YRqHBFMT61xbJPpahWLet+HrApExlO/72/FLsJ
YhIvbhMgDIvHIR0WfabWIEd3k9KKtYYiXF+0ODQaMJ34HdsvBJePoD8NrUASwsEuNUcL35LyOYmO
jl+Oorh3+4McKAicSbveGC3iwhy91MX04CUWV18y9Edaq828SY8hdwAb+3FWucZY8EKFgtVEyQ2u
Fi5J9Go/SpdzJksPnmhxI206hA/KHsU+8utu/mCOch2NCJMiP8IJFd21XNEJ9YQfqKxaQEA1Hw6c
jN1THBASwXsPgKoVnimM5Z1TogG4PCVYaUDiqoHFiioeZ4T40/4hXdJaVp4+RT7/TWbFgQ/Ri6Bl
LAYZ0NSb9d9CtybO9P+MOrjxQ9bnaoib2Yfoc6X42ZC0HSvaKKRVewGvvg0BAzhUGe9gYz9Ti+Bb
e0pOA+6vJHnxDrN3FEQTlMv64zCtCW+u0tDny6OkIl7eOuXtNscOJiKniC4pJS5fivtO3TtztUfU
0CegaQnfUtejbU6ivwLRK8elBfVFfDJlppm80BuZZB878Ctiw24NypIqa/7rXh1WyaMqvCvHAdDC
d2L7pqEyA/I3Mv1k/9R46WoqyTiezcVp8xoJSxeWk9adNx/mRT3VMp3l9aR92l7tcYg96e0zkcif
Ijq/g6Jsxi4YFD4k5E8obgpA1Q8g9no+LDhMgZeI1voU6PO0Z5N5YbztN7WSyouUKmxas4bohkEe
V9qW4j/Td+cxbhvFpgJ806KrvEkb+FVTOeKEtGqHdUinEh4KuVWIBKCHxlJs6ZMMpPH3lG3d8DZV
YeaN9VFevc/gH4Ua03rgEXoPGoZhHmDifLNoXryIgUT3Jh0SA7gbWRu+8ubRYPugfxNGku/mmsPj
+Vd8dkxdKwWBpdNeSboJdr5ycslqml/S2Jor5p4//LQ5DfKGBKBaHVd/H3YB8Z3K5ngYAw6ZekRW
mFNUBzytqEJ2apKrU7F/HmaJDg3hLouhPBev1M8Zc0zfs7/aszjj1CiJxJ/lQCULu3N4BPa82YBh
JgNdrAy8sctxG+GLLXNuTs4EGzlFuL66PxjJnbwLKZPBRv9TlxSYSEk+90tDDgnDfytwCNh3YTUs
creh4qb4QOTX+6KA9Qxs8Q1gqnY9lL2EexyJiONV7hICai3RJP2lHO1Yonar7gNpbpr3wZxfn3hP
04MZKxNZ2eRr5o+R1bf3riWYNvJ8WzVjN9XcjJ1632nVsA6lIE6Pogg9YSASPivAn6D8enc5t0y2
fnAuaQkYl8iH9+ywpRF1NLbijtIdJOm2+Q907oderyW/Hs6nN6EG5Cap5TWX8BltxED9qThT+lGq
0E/xtBVaeVJuvtUKnFSr+IR7PL6raJQ0RBOBdxGAzVMZAxVeF7MD9HWqgeNChh+gfWYEUY73qY59
65SPlRtx0P5pZAEm9OBLN200iNyMDmATh4vwu0N5eo4pWJeAjuDyPTAGs4iegJl5kHKltVx1OBUJ
/50JeFjZrWVNyFk/UhWD3WqHDnn1QaGCb68hJASLb77ehT7RPR26DF1biTGv/Z1PW9pudmiwgjJl
3QNgPDotRP2kTodHN+etF61INDS/Unfn6hU/oq+7Ctn/eroU8x3FqI5W9gBqmrB0JO2YcWHhr77I
h0tUfO+Cic+GpQ52dzKsJ+OF7+3FY4tdpMj7fbFKuzXa6Fc+cj20xJL9/VALymc9arxNTOLhq5sV
0YnZTVbUexrEDmajfxIdZfSgBiZqMY9Y7egcwoePECCV9qnaPsMo2/3xGo7SjC/b7UsyqMIaLkU4
UawN53Jg4RhmieCyDx5EfJtW2sIyN+ReG2MtePumtJukp25pWSrQdu6YYxbDxk6NUAp6ldpQVMS3
LLWv0e+2C6GxVQVpyajDQza5EV7PvDMMnMV3HlMINM2nm2vbbTKMdpqkpaAZfs7KdP8iRUoOgBPF
kTmy43fn1XlGV+GJZiGU8qjStuIQX7WwGRDgyeFSyHG71kyY6/cvoPxZH6Wzab6VdPRMqcNFzfXA
JLP6X6LVKQz6ndKHzg3XDA4l51mdfI2JfCV4/jbft1CrrB9t7HgCGNaUJL88oTaFOHVt1F63N6JR
pqu/X3eweUaD0ukNK3zuaBh62kE860z6/zVaOL4jNKnaSKR59t1BVsJIW9oUB0lIw1k5HF2M76rg
+3qp5+lQuxweR3Y5PW47/mtjWpeIvEs1w1AVh36wwke/mABat778O++FClFRu3Aam2gHsIF2Y3RG
1I+aQeb0kj4cTQi5VlTzku0xkt7j9/2xCwxRm1bI8r+/wb8qA2idVnElbZ8hA7surTWyjIsssIFL
evYvAsChvbNDLkuvw+Jnah3udQV8OXT6GOr9s08VP/MuxmPJGVUlJxkd5D32Jr7BLP7c+KEK797H
7G4/pAGF4p7mOAUeB47V2/dlYlrZ2GETq+eo8UxHJfcFRGsc1ujo2R0kbOFHuKvOJ+vG51gk/uX3
oYGrxajDQIUm4xv4wUzoYLfku+XmTrc1oxPWPYjjX8wo0UthJ/uddcNly4t6bGDDm9Oy22KGCmK0
vWN3S24nXbqymYuFZmd/Eu3jGoEnmvztm2/mQTdu9szbmjaAGN8DRKnEYNivpVDEpX7ARSnHzceN
oomb21h483ifH9/rM/bmZDlbC1vbqtZgUeAzvOs3j8tdpvCjQFGWVBUbDBGvDyILkghKWDJTPkgB
4ULd7sb3FU0BK3o1gmGJnvYklfurg3CHjtjyzS795pp9a1YGf2tLFz2UoexzCguPTDeF8t2Qkhru
9JPi9uzTr9nbo49QMs3hHN+DWprjBHV+DGHzsyXw0QbH4WzTTR36iFwbUfM6nC7GrzOxGRBnHNXT
5+p5G7KvwmxNX355q5YhMpr81vVdqf9bJb4SHkSiBvysPPuO/n290EnlRqvluYeJXFGvsOFzM981
8QbyUaB7Hpi3776Hj5USmu11yYDrSBWwUKkjmPHdLUy5so0w4ttQ8bjuZvfPgKaCNA8Q+u+mg/Lb
8ULY89gdLTFyxBqmqUwHUI4BDoQnRWMvYgl/tdMY2OpYas1hFfGAr66hLc5PLdLpnAPZMmaYYnSn
2uYY9KNFQg9khkJH/paKaQllynLmngd5lr4JxwF0RCBFsT9KrNqS8LtQOelo00BSwhjV+TBeJKNF
LRJwn/y+5RVb0UZQP8uGmtCxpHWL4MtkfMWtYE/wBCFElH1jlGZYBG779u+Kniz7140D9ArRkmBF
kaRc5rq+ICTKTJSQNR+ma8VYl/o5rE55RC4mQCybYBsprJs+W1xsLg4tefowpsWZTrir/HzHhGh/
boZ/eKHmIXbessagKmcSt6J9NWKzJblZbBE7Mh8M2OpMzdn+q8dXZ47OLp/y8c3EZrdBSxgSVRIL
utgLqf8QZgnhyqycx/utKKPapfjNQf2YPhcvsQIVHvTcbuTzm9Y1dRXyGF3/SLiP+Ix6zBKTXe5g
+7YZ0YkMx5iYrFHvK80/gHIsqMQxRQ+BYgbdJh8PDCl8OdTFo+5DbCwyCFOq+/v6dgTgLpY6gviI
ot6bk5s50B+oU0ZFheiR9uFEj0lt2vPC5YM7Jz/a9ECUlWU2eOJMvPWmO36uqUEblKA3Atj29w18
bq5W8QGGE0uuCYPvIoMwMEjnDJ1U/Paz91GXHyQOyGM5pmqOqhuc/Xa6jkF2zgqMEmtc9oLwrvEB
sdeKfD7j8SOoFdBz9BXdc74uFwEVawIpYcPeoJFVK2BLrFgAnMqQ8SoYvDd17HIU7PNDdYVsdDb9
ErA1bV28I7/AEAjQp9LVeJARkAeaZw3IA9BQZiTRnaFuhHYBptCdIkRTbdv+ZqnG3HfTT9/emkbL
zcMCkwqAggAAWBSwVPCpuC83sX/0ub4EciSVou7ZjeZ2/N8A8BLLL1D9Og11hqluTUCKnvY6RZyu
VRaBRyDwmw7TP1EyQ5d378226d5C60pU7NoYn7U9wtNrnnBd69O5/xvpHT20Cv8jEIRU2hiCW1Ul
hH/HAIMc51dtuRD0G9Il2MDSm4lOrPZVyZje7+WZeAK/3ot77A2t4PhcJ4y/WRP+hHtUmqLmtVFY
1kkMm6XwwPqJwVDq3/BHF2L6XLuARWxPkvYhfKJ2ixlrgBfCt62+8/QxF4czPY9BNTKaOwncTauG
iOIyPlh3Y7zLedADGWvjq6TK+r1nVU71BJ/kXOp7hQOqYPT4bkQCzjD/MoVvJznkpnsTVxSnVoxe
3HJnRwCTf1sP22ZAwlW5QH0n5n3SArxhczjL14Bdeyo2RGwHWdx/xIHgefss9OKIbIDzsWOknfwl
Ll7SzpbGZhZiJeQ/MlwoDKW4b7EQfT7h9aLXeZsFX0r5Roj1o8+X4D3V7H5RSF9vfRiPFV76oA8U
05rJOlfk1RFEqj+hq6GJQiqlSBbz+zuuBwiVHdUG+QTAwHcz6M4ChPHUKWKvAlS5pyBR0edmrJmv
i+Z33UrJNaY4kzOzE3YxP8LBo3AAsF2vZP/g3NWKUgT9YW8gtnL4e9nMEImaTNxx77Vu2mJqdEsN
oIN6/ozsEp8zEmhMHy054aFaLtjoTyu+9dpqJe2hsLk6wCVSUW2VOEBDmV/oHWBZjZs5watMvxnN
JOLwmKYyXU3NwVGX/B+RAl03QoLampNkOuJFWK36vdVzg9f2y575YXPwiSSX8oB7HWS3CjawJdMY
vGsiZneXswL8i7KBsIO5lM3xH9q7b27e2zKZ0fltZXkK9MLqtguwF83OunuVHTi9UdDJU7yfyJwa
CwRYZgcq0NFTORppYyIr7SaPprq6xNGi3BMofxLt202ZXHjJ3bSbFFiuCJgwfEw30NdivR5wwUgz
ASLIKwiJ6F5ttngRdJD3Cp4TIU1p3s4+kd46a0yAoSdWPM3ZtcYLUUtTXbQ45kxyH8BJC58lQ84y
LLK6gV+AWn0UkJ+5XihpEUxq5GmQdVmZmWrBKRkxJjSj0F2yl0r/8U3IaOq9yUPv1UI0pysYOKq1
ZoRxfzTkIdQGJiDOeIW242NstGPFbRVG3ORKjzuQFljlh2KPB6KRzqkPREdco88y/y8+WheNKKNP
apHGU603tBEiAzR/UR8nCCNetMkIXCW2ea1PLgndkfqIm+L6gvVZ2JR7j7sgEz/iVC8FqThGV2K+
v21a6GoBmeIihTUJqG82gJtQuhJELnFs2ImZazkoS0FD3iPQQxARPWluoOFdEH4I3Q7p5/u9wNmU
2VaDQWn1WUWDL/x3i5ZPFuFFKgFfoJYL7tIy3CtDFrj2gqFqP/y8nRDUqk2qavGIH2z8t9oHwXLC
wkOB6SALDBdx3fxWDeLhSP+0vnCp/DnoX4z98HQwEeQ/aOeCBTWgRb9mkDt8IJkslC95xdwBrw8z
8+pTrLEPwzhHqmwsr63QbV5eJc5qk2+K2YO1riN0vfv3SdEUjTkdl5UMCf98wS4JNlOb26wk0dvt
mLhRNlIZCz0ucYjYGKSrEjJVcrYiAVZUFWfCik7yVyJ28IW9KeNfGK3nAPlecyZDEP8JtwH3mPEO
84o/0PdTFXQQ8GEUjawYukrNN+namzRceJLUojA+RRUP41oOp2kkEnqCp31FDFRIg5796WcQCbW4
YrYapoAqpYKlfEptFA36vzke+7OsCszBst2LCSETgOgeIx+GNRsZX3jkOU0OTIZ0MUC88BdtChlB
RvQLJLXzPb1T5JhDZPn1IvSrbNhhwMvLPVFUFPgoUZ+/JrCDsTgQNt6qLUceMpJx361th9eST3Da
/ko2RIMjG+BuPeuYjo5ZqbfyU8nMxp/28ygyAuTHqIdcw7FFREOXDZbpvOuManH/1WyPG0slMRSA
nnhGNA+o7Bdb7G+TKqU1H3DLiBxoLzmb742iWHRsnZ1TksMHCX9EvP5s95lAHQqiBF7/8NX/6R+q
CYlwvec2mk0tyeF/lye34k93cps74YOEbpaOic3g3gSfgFYqA/7SvaVsxCF9BAxkn7Vb3hodPrln
j5KDY8FZLgYDbPoPZAz0K1uNxxHa0WS0+GPM/ILqzqgb7LEcNsLp1OoFbr/JW1KRV4JmeLPg/38o
my0UDRI2zdwk0/P0FN0UVhskHf8i+GgwdxmXcqVxRka2OmggtKcjAeijeBAvXLN8LWbT99KjKXqc
cNGMBVEFUOaIiijqzhmiPi8INGf/ByKKkL97emabNP+FWm1xdzhp5mR2PNy9atOHnNKbRVUfU1gE
W6A7xEivItRhN65mQQh6Qp2FsxestpDIdIslveEWjW26phjkNUD8tiDttUsvq2QhMEWSJYJsR7th
k6lE3cfRK19ijkKi5kRsuyRehF1SIiXQtfYYAYc/ZQqM8QUzMNNBrORYpJCD6yzGHdJYuKhoXwEK
eJ3S4bH5Al+yYRaCC63Hs61EPmj7WJSoFZZM2eUYWFEFQiZuHwm+dXeXYyIdAe4vuMOOBxTfMTfy
qE9hFm4C4Q22Q4Mryl3wz00FikPQ5BzxWdgabIWASqwImQ6KyeArY5Ge77deJQDzVItl+qN+GAlW
IXEhxYsvuyz4PEwIo+WWUsFkz6DdmsRNtITSfGKNZ/IOK91ur/cgzm3Z4cpjVeMt5rRjkLo8bkCD
fUlX4wW7GKoyWlWpNna4tdHdRlw4u8Nm9qRrwjQdrT2SC+iau3GEkiCKtJ3VeAavj7yX9JsJ5ynk
87keVdItBSckrOpZlyQoOgzFphtxTLOL7aZ5j65FDUpW3CEA2GScjs22LtxcUiiDCB1aOgp/MZ+4
tNocWo0mdRFKwXo3yEf8KoygfHjGpVFvRDsgm2GEFoW54/zcQhRuyP3XFEOZrD/sdfTscb21TPFf
oMZxNlVb18c8d6pUycNL5V4PUVAwycBLrYU5UK0yTw7SxqiHh+b2FsiQzR1nWGQV8t5vVnxgUMxQ
ancG3fXNJ8QbsozgXtSHN12+i6ZgQD1vlQwdMMOyIdDwCxETH86fAsdUzv6H4P1GCrQiVtKPlkDU
MUG+E+DYGDaRwAGMSt/X9KDi09gqrwersTBFkIUobNHorbRnwS//ilGhrySfEEyL6LfHzbDfoWBz
6V4YspRFESeC+UK9ebfG42jE0CEy4rHWRprSbIuos+qCnAn+Glbve+mNk4fCWhTDZ1cZV9SYiQl3
ca98OHSWJFtzz4DOJ8om1v2pth2hrB0c805wWETDCG/MJwfxy9VaTpFdN1wouX/BYgGA5o6NJKsu
dSARgXPnD3RcvmgjcGk4nVQCJeZ23fD1l5HCr6PQX66KaD3uWHsnX4YZR0+RIVOioAW4qD+db96I
But6S8ORpm/djL77ofM+3b69pnMclSThz5tpraK+nhn/wMOYnXEtPoShqqq+zUYV9hitdmpVRT7H
0tq9u1kuQPetc8wIKce995kT3Vfcpk5sn6jMa6XMlbXxhDdS/D2H4Uziz5OIPzZ/2YsCXcAGAxZh
uJ25e5onGlauOF/R5Jz+SSvXMFcZDC/150kcS+GhV+oYYu3GF13N/+iZQyErzTqGHGXR7Kukb2P6
5wLs/nM23CgmmOCORLNG77RIIR8/NeEICR7188kkqzpKch/QJV2lHoQYvKRThd5QZ3H1iQ0N8VSN
CDpDCeQ1x2PUGDoWAlAx3IOLfhD7Askmxr+Q/QikNOCOvmwIM6CQsmcTogsjyJ4SPPCrrZ8HYnoR
44YFzTU6370wvEgnNfKCpmzaRFlPU6gw7kyyju4+tda1sDoGFd4G5gN10ScOCZcjk+83VQn0q1YN
PsVqYWBEZ9AjQUzWeVVQWif1IFO8Z+v1u02Tdar2aqis+eL2XDt73nSng1l7rfDxR2gKpbQPQ/it
7lB6RYvOo0hQaRK7yPbsuS/gbNat5/ZuDocBX5s/aWFOuStxOvmJ1AMJS1VNvlTa8aiY35IcCJeo
wUXGGCxwQ5/jmS+4JIRMlAPmpWqC/B7lMoz1dJZrpOkgnKv0KUY3LS9gXDN553hEKCZvoL/4MjcO
wHVN56NhcgPp9EjNQ8AA8V/OCH2Hnic7wIeV3SMlIkrImqG+uH2+ps+W/+0QRDh3VMAiwcmLzKBk
zhGvL1rIxNSLpXe1sI5wdDRu8VKGgfXZb3Ldf0FmokHYha9hA3Qlz4K8rJN1InIans5Ix6JmkJR0
McMsoEHWF1UpRNkeUaRBCw7pJ5Kylqrv0fRXNf+x4kgBleCenNBSdMBBpfv4cDJWAxIsOKLW90tO
SiykitUp8oYfqfwMpd2ZLOFZ7eLtVF7Ygn6SeioY7IQc4j56xRB2VQp1NaHXmwGC71K68IDEPeSt
LVIwmTY/RKtDHiO9/72ptVeXyPlzJoiBwPlRZFJt47RLzT2dKjPw6T5J5XucbBzdz+jeFcLIVKb1
yoF97Xlz3DZdlPDbKmit1gEdLYbZVQNzIvDIDQjiwGFxIzZu5gVSdJizKDGtivfs0zPdZctxBXBh
8mEKuhyphkwUFMZq8NuLMbhZns2NFbO75s6pBjGtiBwR1s9zunDTfz/HYM7VqCVwhZSOlqipMN5y
vNuhQgh0xvr7AeFBQW5KZDBJvEeHgpzcxRr7xaTwws8NutqNYnxn4+eAuB9crg5BohUBsQiIuG1P
bEjrWYYYldrG61F/8TYQxILRqjUn5UiyGWphkp1KcwQaJHAyxO0oQy/2nqlOqCMUDXfz/7MMiR/F
n6sl2x5vUuZsIsiZt5Tfx/KYf1VkPSpN1OwDe3V7JYH6l/Cbt3PhgNdRK3D82fHq9XiP8RxaFLOJ
n9f/nXHVa9HvoBZB+KUON9Z22X+qRXHhw56KgehPIz0PxZZzmAWoflG17wkZ+ZVmjwHatfLPfciV
zZ5no5HMmOV0FPRpREZp+E3b+k+c+Jv0yg2dtgdKZdO/TNPvBfgiW80u/FI3kR7T7olEwIeHJ/AS
t5gyDQ/9OKr5xmBeDylcD+5flUENiVMLVnf/sHKC2fk+2kve5XbKAypvWNqwjLUAmXY68/yG0Ao7
SpxUPlSkE8utfR8NBmpKXnyxidIymBnw/y+sLyZqo9ocrAT/tH/XZlLsPl0wopNQjK301qb1dTO1
5VuCnRQgQoTNap4Ok/WkQWpTTnpKmU5phRKEJevA4gaSKNSqn1a3eGHLZHXVmS2cFVssAlZIBh2X
0F6QyYqF90oVBF+I9kzg8cggjfyrSqQWccBZZf7vKR7hXzpCyHkNiJRBi7+1ZlyhU5NUTAHPf4Wk
HdStSfXcThgUsGMEhSKcrxYwY5yLpKnQu2BjFpJWpLiBqMks9yZ2f5DezmUMsxnwX0v4HOt3LLos
vEpZ9Zc+YoGmrcPbLhdp0qIcUTJi3yUUdF2zAeVHDWa1Of+GvCr42qeOKEkm8S/PeFKyLB0wg54G
xLRQOtCias0citN6p1jpJ2Mz54qCIKQJg1Hi+nH/4KCc9MdrIXcKUIVVRTTXwoy5gQOUxZTfO+IN
unTwm+iMSomUKCkt/gwV2oI5LUpPwGsgBFOeVULfSpA43JxV+aRKtUaxXbGAvyfCOtn9sr2grhQz
WJcfewAdsx88uiqPY9YkBJeZ0T5gGdl+4S8WwjDXLlFtx/1zjLoQeBbtw6OZCXFhs0xJEiclN3No
WyuGChQ+y2GsI20Nvu7bwrVoovnVZPynPl7EeBMI+Q06F6U7wlsmlnbEUoIc6hxNLkPVWkg3p3Yu
3odppXkOgC+crlHiNS4ZMGUl8PSBnlbjMTob9GoS72X/rd/0aunr058TVbT4I4JG+vwUCd4XQ5Gp
7zJs3d+vrdueUTmjN1OvzHHBaKzc0ELckAM9Fuvv4q17u3iX81m1X9WWs7MGpxJMNe6YJpf/9B5g
6Ya5vjl3VH326lqvXqweCVsyUKcZzq+cYbSP5oRmUYZkhsLj++Om2ODHPXJn4/JNkyzYLKB/Beb9
lQD566I+ZK2yMhHVP+EdB58HD5TugUh/3BRt0GwmEKio3KJSN1yil/ZSH/GrT3Jl/adGtAA2Pzbd
m7g5CsCrCUJDl+PMvKF0qx3pYxmKquWLlAO8HxNhjqj81usRQReXgtCQ2Ghwv3v7rVOQCCDYshry
zpmZybDV1BiE/ELSXdAbQgEv2NatCv/FcvW9CJ3fzBLBFXGtqSz5MAcjpB+m2S7joyDGs32Q27hy
DcYj4v370qOoZpZZwGQGeRNzyI4cByB5inhvhvCm36E+62lZDuyk4aJ2Q7hBJXBlpPYIo90Ip+RI
J8ammo6MjTVC16B6YFywgPgYGeKmajHDzKVNfheJMNVc0qr/YCD+KOwpaS6E8jIy0T+wCbL69mld
+ua2Ux8lGmc/8aOf/D83g+BnIWBkK2zkyW2Xf6JMPYXe/ndZ0QVYmo4MQkXevQ40nbrzpICaivo5
YS0jA7bOMX0SbmQ4K4fqdPhipXwoZN3wklXUbmIgY/ArWWezoP95z/2lp5dl8ciQ2zHPNZWjCx1L
vgb7BLtcoUiDDVTTdD/xUx7uLzY5rtaVqAP148Pv4UHoe5W9n8qaVGNQs1MCnc0VEyr0+wyNj4nM
qwaQIYruY9fzoOrm8hLBIc0x622fqUa7NRSaRIBAvCnyqYJSA5Vue60I4WxgDEwSk5Jwn8WoVUFI
o6ATu4teufBY6l7JSGqOa7yw6FmbQ8XJohi95GjQlaqg2tEoLMSw7m02VPxkGAXNyGnZPSKQzxi1
KiLvFIzvEz6nlkhvmyNeiV31lrCYBz9vM3RbTdmzJDWsFkQEFzWuJHBuJSdvOKbsgAn21Q9Ot+83
5mqx9RzFP68SKF4o7RX+yJYtSuQtpNUvE+Rg7+ZESTWD6wQeifq9RqSWCaXmtiPjMQEOyAFpQxdF
26kJGMkMLOIrwUhPYrayn9HdTvRowpM42DIU+XI/NI1nL1GWMFMH3K0MAxo80FPLFswxZUNuQ59k
29t3e3ltPMwaHdx/h1SXCz2DmejUjsplbQo67mQ5qvPK3wwkYU/RtdzfhgEm8Pd8O5v8Bc5PCgG5
P/NROULrZZteYguy5NKjhyLCl/chXjXoq8PRoJadSVnvKbbMEn93j2wENmm08btkcKUPIPUD0yfm
7xUamEVxH6RWjIgvHI8z0TNdjlUuCtaWBEJW8pDahJ+DS10K/VevA+f8HNluz5U6gne6G/AvHUOB
QrulQ06Mgef7LBRouE6IDV6NUo7g1qV5gHgHRjUZQtetp4u/NMhBQ5i84bLbP+IotgOyXM8NLj1M
5W+61LixkHBMKbOhedL7czVM6WaAHRwktL867nFlxx2OarySeL+FwcLAjknINtMYc/5KllBZOxDh
TU9wrrUDCyAvQggMkEPzYr/ubkwptbvzQWzkhtEgrPfiDYhV4A5wIOIJnVQCh3HAw6TD089GqAme
Pkrd4y8uUvCaW/0hF+WaPkoREzVA5JQD5wW9lkV6w9blZQ5B2PRA+U9OcVWtRCDIoOvNJBeNHGNE
yerRwNwb53WDtqWedD+xlZ7vIqvpgU2qgHvCwjgzoAd3OMj24JWPu2H/FlNnVbnYC4eeVLuk77uH
1VeiGdu+7pjEgnp8PYRpZ1NsrrhtvlMT+WKqJ21oJa2H0kQ6HBzpf/ng0FjgB4vG3PSQha6a9Kqk
0Y9Mgf2LInZWuk6EyJo3VDkUaT/Bie1qknR/lsA0SaQ7Z1VjLCIS2nuH9mMvKxHobjZw3ohnsiej
435YpBTB0tH7xktje2s0DhiaURpOhQKGNUqiCzCR0tsWjm0iekDm2qkK6D20wjJnsJbbyKjhxql7
dlWbEOe+O9qBbkdN1YOsWI3yuC/y3YIWD2iYXH8nwhb/h/y+SICwr5W5kqLeiSNpqwGx6s7rVSCY
SInbLIJqpgWsrraA1eZbHtSytvf4WkNi1BUxxbXXiq/5eKcSCvi8rXxdI/INV0ikmfAQgSE2QW7x
h4bPT4DhprJYkATmDW0GJLsqBFkzL1aMZhdAZb9sxUhNfblgpyN9ZxL1m9zD01Q4r6U4g2GbT/wI
Ka6q7OvLjxQoQuPWjr0Ht8dCOiKTBcka6MxURzJoRO10tkVsPVa/o2gd7V3qdxmDdSH3yyVm3k6h
vVgS39PLQMb5UIsxq7GBC+3veYMapxLwkPt0UJflGjbr8W4A9RXhRQ9URlKb5HT8EXoEo4JDxIj0
aXfoTTQHdWMFQUq7A7xU8rW14+Z1pNzSZa14+792sVfqpevIMBy57ZVcQrUkeA5XHLdmBqcJ5gUq
ww1KwH7RwNshHYoGr9ltExzYXGIT5+xqmAUoiO1ricRfzmKdxhek5R0CCylb4MyQoMDWkWhAVb9r
m5ddpwpKWm9yE60EPOmFu+fqZDMlnuQ0ZpGIhOT2TvtwMXIOd2cbhyr73r6lLwGrIwYTNJvU/Pau
lbsUflCSDWzslEd9tH1L53//FIMLn1CqnK17YMoRy8BLyYRnNmJLet2ObZLUsMTz3SO3cqBz4Nfl
RpQgQ2GhXCmr3XPccO/4nEjBnPtfTLNEA8keM/KtvqElNxHNG6Q0oMjviToTns62iD/BrTorK13+
yOoopJCfNk9ox4pzq2Sdb/vQJNFiJsoTI6j/IIccs3sBpsVmier5Q0owK4SIVvrtXelEOzUCiiwf
QSUTAnyknihZEytdcvd7mCqS0zfbn+FzqYRgeaa1C3IcUmqqUzzCP99aawDXOO+v4mCBjBFUygID
2aMAgIEDg7EyBjdeCNxCdWb4HRSl4GTYDGRpk1DqDkmPpIHWIvnkDhKeVhpAkl5ylG826Oie8VcP
P9g8lkEBtC5678hEKnx4RhHybtrKQbEAQ/AHlXZD7pZ7geImWupCT7GAfmBvIvXBQ92hhzY3xyaZ
nMcx4GL5MkauymDdhzCkHUBfaPULPcR0YzmR6USd8MMzlLePLsG399vlKsVtJGZbWOiwAb3sAWWh
B9JZpE9bekPyvNPS4R5NRI/THoh7jHHXrNBDAxiGnwH2ESz9M8F8MePKWoG4ADcLgaycZjIhkJEf
IHOiBvGNO63wqen7lkcChtUtQfV65p3YV/8aasfaV4QGpa1zmWZxtktkTFdgVRPEcwxdmYWgsnnt
HHPsZUdxlqnr5EbuECaWLgVUiE5EaGzyz8by/mwOnH67I0CRgqrDtmNhYRzqR+XnU42doicfwu9W
eTXPbXVo+V7bHWQ+/QijRbJDfoYXKcC0EScH9Uj/qdRn6FH2aZ8YI8WgFmEs61HsoWSGWQW/DOaa
tpovObuAfJavEllo4/h0/UqWYTKy5ASL7WeO6SmfP/JzA9P35WwOJ91wFHA/pqUsrDlRmZnPpv0a
r7zxf3baIDD2nuMDrHuF6IInNa5u2Qb3hyWXYmUnSFvDCAAlbvs53HTNuLtsyJj9PFn6fV3odpWb
VUBSB3yKDvsYQK+o8sStkNl4x0Kzn7tLQxkLnyk8IQsdcO+OVYfCPrfyRFa0BYxXkA+NubFywM3V
D6D7zCmGIw89smYEYuLDWAsIVras18hIf0lDfVFUVJKMl42KUUTAaKMeRp831YVCnLeSjBaTIJmA
z0KKpdxA4/S8SA67/M03IET9H3Uc4yHCNWMA3LSh/4OEBtRGHP6zjpbMPOQzxBXgnnWIOy8lEGuR
VjOJj3TkvNbAwruDcoDB6wcO5N7KUf/FOXt6EfPS3j7u0SLrcaAqyMAZNNxSKQQOef+eqzwsIhB4
TxWqcqu0s48H82poz8HG05b9wJX0yqsllKJcVLfCR7lRBFHlNyKy+uer5K6lOfLBJYk5TAMnk01v
ppWnU2Moc0C54neQpIkODgugZwuhUiF0Ji9Q+dhqeVVANwu2KPRZKFJxQNy02/xe3HFVfHRMWuw5
j3UeR83bN7euvJswc3qpjlN6AsiTFGDxp4AbpQj5UBDvv9TkUFQ1z6SpJiTl0nbMCOEea3dc1TtF
uJ3zXwIva7QXmm1Xtij8iOOXBfslQ+zHHrqje5dWitpArsYoj3jxC+C0Jq8qDSRc3zTVeAYbh1JH
N5slzO6pNTiE2mGvwe2NLSqf5Ixp/4FfU97f7z+Pt90g4JjeVLe6U6zOZJpF0AOGPLksmdEBbWGf
8GkNpYAFrzeE79vcIFUXbJ+jMR2swuNqkkoRmDVAWjRcyqv/vGv/EBcDQlmZIdJpRUVMMo+AISku
nv2L6Pjt2yn9DeO/FDzM+ltudcuKj4LfGW6ODObqfXcwTp9Kx1W7x6W+wUS886WrCHNKA+UmiPCo
d7JhuKrRqyxwXzEhK8UU6RkRofns2Nq9YsuyDgAULMX/is73j6x/ZRk0EWRPCRIyRWFxduMU7QQt
YMS6qJ8a+DR9NH1JMNgMkG0oubTr9j4UQiJcQ4qBWjgLGOHT6vegjLYmcLMVVGq2lF+wKSGTXCFs
1C2Ok56icZH0EXPi3PZltViMdDI6Y34l8Cz/9ZyxVAdj6xjliRuI/kH+tU76Fg2W1m2avyibuxKG
gNo9oD478aa7RVFzjPXqH7u7uMLaf7hXfKLDu9CaxWnq9jOglGVf4l1n1+Ue7ottfHE4ovKCpTH7
8+gyzeAGrbWhfiYO+O+Mdn57EnMTnVumr1s+R6r2nGGvDOuA4t683b/LHbWtYuDyWY22Rjfr5t32
dyybhK4jw72G/FNONpCSL3UD2PwyIfk5O2J9WbeaTwJ5N7UjiRKxrt127fb0m/UifG18/XEq9x11
VPWfJoXsLG2Sbc+5xAeydYqWjU7z7HCN7ro0gM9oH4NAkn5Tp3XJMMwKNBah/iDaXRWJ38ldtwBR
hJYvllzPyu+6UarFZMF9wIOy9ftv4Kf93z8Wv1Mzit/jr2hOufO7iNL29oqbG+o02M2G3jfmMx5/
Pjx97STwIbirAEvU5EbA/XwcATXUt83OBkpRCBstXqYQlPaHlpDIuM6x6su0laAR+kJRoUWP5bzc
s2ZIGZ410bqzlT8RRSYuZbHouxsuJFEZMb1Mhmf89kSoSkDUBrIDrIE93vTnTPiljGMbdXXtizcN
tsrZVz3wa/jokWUa2EsO9Bm6CEI5ssn4cEsthHvjpe6NyhOrVDusns9hdhchJgPGELTPFlYC4Fe6
Ay9rn6IB+0+MMDeIFES+yKuv7OXlBySGN78xCT+tdCBHHTZ8dNZQDSOZLffEVF0gdmP92u0RPwqR
HFyJBtomOCf2Eusn4uRvv5IWN5SpRHOsHrLFC7UTNNQnNOJunPXSB78wFPQh24kT+JID292h8FOi
ieXHtXVlDMV4WM7wpToeBd4HrliKjZQsSfaczu6mQo0sbOqBGy0q74vMGCC2XYiCn3BedgljoEA0
V3krBtLlXjWV4Yw3M7wrnkOgUWzMuuaHu5bB1x63oPcR5s42NC9XRDFuvVKaxMHeA8wihFSciYl0
UaqOQebyOGZrA/kBDAVWKuIQYMgoWbd/jCx4GdfvGO7aa8wbsjY/pqBtoxkTZOE6KrOSGNdGCn71
K7lmxlfqST1KIpeqkiJaNWqyGQ/CnALtZzjnTxcE3pWreOnhV+RZLv6QpNwdSYGR3fTYS+u/lPk0
r4P+I/P7bbvNup0G9Kg06t3NSIlrC5y6f46kN9J4skgB2J/FCp7QAhcKQqX/UZRDlpJIvkdctix9
h/WrFHG0hoYquLUyCvkpOOJPxIvRcX4OvtT76HpzEBHhkp1toQpLzHvY8imAg7G5bcArAEkxIt+d
BWS2WF/RMJ/e84kiTfVyQjIrWGwSlmGT1AJ6CC7LChu/vSs+ErKt1P9pB7plPx2e+zNoG3Hmzvu7
WUTyY4+RkoFCFL6ZcedRk9DNP2sBB5FVyLn6QY92GxTQweg1mFTqYFx2MyJKsExlAqV0xec1scb6
4aERRr4iaJ354pFYkldMmH5WmpivJQUF3OypAbEZXe87H1xzp5ygvVcB9zvX6tiY7hapoNwDqFTp
cv6qFyNsSQO5RfM+opH88W0+Tw5MtG0XFYHHnkmvwFBHyhwUDNB5ZhUxRZ4qwUucfxz1PlxMQb5w
jHP72UQHKOvGZmJ/pvQ+n0MMVdGuAlfcZzeTlLaht10i5+M6SmN/knvysYsdEnh8P9l9DvZylBs+
poliAGgDb0vtalQwlKRVYT3MfPwBuLGoiUFDB60g5I/UHuWKdt38PpjQpW7bngbQYhv1G0vvKOy1
YERlHv4kOzvLWbtOmhi3LVYeqfqMIXyj7KyCcAPGwdTgEVuI5W7NbaocJd+wSsLM5439X++bSnFA
pY5jOp25jF95rVI250BiZp7ps82AHaOxmV6lzmGh6W5WGJp4uw/Jx+aksINn8O6x+GmnYAi+kEMM
b1y5EtFzU2Wzz6ElsW/G+c9En5fXoseQNc+sZH1oXMJJg7BfMFA2VxkurFw1HZT+YKIi4x8igli/
CXk2ohEgZwu2cCZBfQ5JZmg5oN+REk4n3DeJOweTmcQ6dZ7JO543rIRhC5SfdY78Re5r3mhWiMdh
SGP0ONo9LMNzQx48GvKOv00LWHSwUd4T/03euYjICt0UMbtHnpan+ZTfOfJSkrKLg1MP+LwRWT5C
W469ubdDu+toNgvaQhMCRqlyJRU3XDbiwE7Ii7HZw567g/DPjkMG2a/u/MgGm1XvGjpxjwwNkqlK
khUu28P/uYmlhht+K34cKpexAXd56kowNfgAn29EiXUOb62B1zKhGc+Ph2WQ4ZgMje8de6K5nexH
yO551Grk1tmLa5B/byyTqZ7PGaS0YnZ5sL8+1WE0CgY1Fc3bgQFhbjiGb2QG48eJMgpU5qfSNl5S
qA1pvqFie4+wmaSG87bolc4RcVgiIBjIMEN01dnmjwvgtxvq9D+FT7BmoFI0iMVlwaWoTlq4ETr4
ST/5MEAmwBIFT3bBiyRbJNxtK3QHst+io1q6AGdkdYm7ucpwpVjXDb2uk6LyppbE1dIEbmt2qzDf
oTaAaf83AenqV51gFoS8J/JtJfhbg25Z0RQJWWJ6AEcg/ovfaAaFdF6p1NC7ZLJAw4aLr+pGKCM1
WcsST9MrsTXNA2pLGSc7XOwnOgQAndn3FGA8LlOEzj/Ci5Hk33XpRbc4eiFinjykBSZ3lnfwDbfm
o0GNmEOtu01rfVp/M+waQ9AW3Mo0Qs8XVOzEC3z7hvux09b33IMBEaHOE3nMD5FqL1T+4V5+xbAC
N0hjIvSF395w3g4nLQtSgQbBRM9V4tACEGIMi66e9vsD26kuh7R8ybjWg4Wxf5aBcrmZeTbDCPcR
mAZyhQdgGpNLXBDyvIccZr6kV9dKbnCXV1LzHY0eP9zLMEtraWaDMCrcr8BIeWEPF3xZ7+2Jl4ZE
CVfI9KpfF9jCLni5f9KVWTobFh6x8qXAIH/7vTvt+CfFH94PpUrcAJqPom4RaCIV7XO+zvzNX0p4
HFY9DNVyiEGtEhEyF3IYol8oAoc8PWVr9JtLpHf6HFt2HMiGdIj+VQC7hjDdMAxk+DHLvX5gRqVu
Vxa7VHFHNZ/BRrKhbnLRM19CB2i15F0EEeh6lyGcN8iTiFrQk3tLOqWIPNqjnHXfwHbKr+QwFPVM
wg2lOantnpbM7qgGvU/ItWVMvkBC6Q1aq2G7cqlw5zn2i9zZMdE7Lvc55d4XzeIvyneB0Vr2QimA
OqtqJp+pPUblpq3hN9aZE+SbZju26nSqfdQVX5HXTUKDA/UelihA5PEbgeWq+/0Kf2O7IKjpWVJR
LS0H/2WthYbIqq25ufCyjpa55Y2lH9UDKJCsxlfaIJX66oPgHP27xpJVZEcqR54W5nWBCA5xaQJi
WtMHk35LR/7CQg/enaaTUFUvim/38aDKv79+f3mmbGJwUS1S1Hh33c175UQQG8DRzjO3y0MaCMDh
4u0uERpLgk2G6D9Ju8iPo0utmcw4AvNwdlGHX5UGj3y8OYTOW/inseu5Qdo4rx4xRXxlyP5oNuyu
LbPhWnIp/IulAR+pHTh5kfpPxEkixL+JnMSqQQSTkWdeXiR3wZwnzAcCp8Vc12ib7SpWtabdRq7Z
0f1olr6RK5E/0I5tVNbZ11TBWppevys3dbr1J1c31slUoYEeybulcpbZ+ps37x2yMIzzfMAh1Twt
yH3foPJpxWfAKcM7dTqw0DttDAXXRhGiWzRnYruzPDdrVoQb45GxLljYLH/wRETI1LB3MgP8yXth
nONXWgSy2w1yg7Ko2wbkMwrEXufU8IYSkGV9+bTTd00iyrKAPLWXBINXTRTkwt3TpiEO4o462sA8
Y/sEJR3W067pFCiVU1Ib5FIQNmfOTkdxcGRFd4VjJm//qU0fugbALgvhd8ptgLXiS2Yohj5543Bt
xrGR/YSb7QLVq478ideMGqKoggjoL8jWtTX29uDDGp1RveeVr2LEZgfTxtchZjzoBdfxKOTxf4kL
LBDxyRM6ClP+kQvPJ2ge/YEZpkZSglJINaAg/uQgNEufk41oAZbC1MECWpDF8dhJgmbkrO+OfOuN
/cs8/4HWCRrd2gHroDZUIPlLkofkSVfaC3JnBfTomCqrf7MofYZQoKsEmwJYH/po8ELiSKXUsfDK
ztxGfYzZfFJe579xrH3oCtf8WNa5duzMSvIBZMccB31C3AsC8vpd4n2UHaxFbDeLD4Qez4ksPcOY
u7jzYWC828imkos+uFvpxLgseuov3SYSJuIEyRcQpugeo53vXLG/Kwu4cnRVXo2O53Zp8OmHSHn7
pphBaFtJigjfIfIgNr8kuGpJs21LMOxczod7xFOyg9aPRYT8CQ3aGlHvV2GZQ6bToz4NHkT6Xxtg
OpSn49Ctt5RWKksHIrocLt/fhTRik2EF/L6NcfXIx5ArAjpo7cfhwUFH18Tfkk/drspLFvJMpC7w
7AWKCGJnFHaXsHvFA2O9avIZw5T38Gpba5GEYwVI/x6hwgWLk+H9I3gL/5QifwRAik9A7brc0xov
xy7c48FhZ3tyR8SmDoDWw/3Hj+lBNV3bE1nDWrvjNQQRD5UiSdemT4G0lGb+OCH9Voovi/ZbiJyY
YCFSqzmO367lWo2gQBmLnLUck/apv7ius2R4Q1WSVvWMAjKQYucNH6ikTOsmF3tXBjEG36BgeTel
ZOOt4GGMtZjSKmE0BLFAXPVaE6Sx40solf0jFrbOOB4XvYGTu7pYHxq/cx5fgyIziHisXjZcl0AN
R28L0g/tyVBgEtSyeEM1QJ9ga/eM+5pVjHbNIK2uFcFTrt4L3a0LWwhyYb4F6jQ/ekkT9zRgdhyg
bsLPPQDL4C+DsAQaQe+ZqJ5pWwoO/ucnHwB6o07GYV0dB+43Poz3pRskTTO4wsEipaWs7+GmdpBI
+Aj6XqnGGrlngxOe4zdmgUBUpwgBVmIv7mFthZfbDMjU49+WKtGLUdmYHh/VYVHTcMznmLaPVBL1
MjSArrHDEWYq1hQ1l4pDZipsOIcVonkbrKFMVhf1BlmlcDM+pFu5cUuBCh0xJoQFka2fWRORlGzc
tgs/EIedchzQXUwWiRTvQKFkgtXCz4joH1XEEZLYxArlCFJ7Vud5v77dj6lce+OEZujo2z0xAAPu
YqynRlUAfB3WirII1ljJs+HGgNLBGs4MCs6Q5iqa0Ib6E4jA5PTsRePg0jiev3PXVYf3IyOdXYo4
57YvQh7lQREko/z+IXZZRGzQVIEVO0S1fAYKzg0wzVcVJoxIsQ/W6HhIXNAMCu18IPO9670c88qn
5b9dfzc9UP4+HIz7k7NvLb4oKx9+u8e9GjiFnP/rXWMtPlMpD2B9c/VyeYfRdBEjZehFmDb63xnR
fGXNSh+5TjgE8G4Z06JemiWx1kwjiQyRjAfIxneje0AU+SGaBjibXNeN8Uv1I7AIx3HxqhgKY3sl
Bz9yudcUTiM94nEBqzQmaNyQt/+bI286Vl3eTR9d+jmvFAXgbISrul82+vn9P8qBdDCQ/rk3zNsb
TklwBrJod+oGFbuaaoGrD1LtdSeMMIMPgLWv47VhJgs/wKcxoKrDb0aoPVTjGWUF/dv5fP41sGxR
pTnMcRCK8XivWFk/VL5H9XpUoiA765dCuLsRdNMKbJVdearLZ19wcmpdVlHzv5V+6G66n4xfD0Hg
J4c4UkPOgvABc1WSpoQeTrWqiZ8tMuBdtTATixzbS7iOoweGXBWxaTHlWw3MHMjAKSEpbrwpXxh1
P3j+1e4s0SPMDaTuS+S88cvKm0y7S3pSpIIYhaWmqWWmOW3L2+39GlFjjlutzJjC7+cjkh01emmU
IsVv5OjJTdM1Zaiw+Lx8KuYZzMZ9RWr2JssSIFolfBszICV2p2rgtjaucV1R2uXODPL1UWlvSoGK
x5ovI1anxrEMNUk01qvApIf58iwf1Nvkkwdv67nbD6ujFXi59ujsyHT3MOS6hgFExTSoeH7oVEM7
8jxAgAAog+SYMVkC3VRZyMVrGlIqve3WdIJ+SEJnQoLOVIpu5Cim/GgxccSuE7HcqJtd6gP4FS00
iMlQYmSElNK8BtxLOJXfveLH+qTG5U7p9FEqTUkpZMF+Up0nsajw/zTOgb+M6cDFgigpVgl1EfB/
SBcUs8vx3lqPtWufIvYvV7O+tZtcP78TO7SYZPhU/1Kef6K8SMMbuz1ZyqxG5Bq/UhEy0MWDdPgs
kNxmANGLmd1NgE5LyzCs5OannbPqjF9eTPYMhACaYxqpPvmHWBzGEzBaijQ2cNJ78R3v4d4TY64U
EsjPMF6zxGu0tR8mYC2t65wj0G2zwqbpvkIvjYELwNsxQU46iQPA/MRxsivgtLC4YpDLankeEFCY
DLvH5VqLnAxL0gkCmG+DbxSbDcEoOFv9bHhrVXZzyddQpnYbbGDMWNWNSOIXiWdqtn44BytfZeJp
iKSZUoaX2dWcD0+NkZYJPM0sbZzFy0PATx1HRe3tp/Xip8K2l8BA4S077Re0DM90o5SJmcTQTfw7
WbdQYWLP/iW8IOYGkYc69ksM0oOTECGId5LvxxEcbLyJ384NztZ0UbvJF0//UAxI8PNs4/1+U6KP
lzm0gojTkaVWS8CDwsJByJU6f0nFefMaGgBn8KRaRWoQdV6JV52eieF4LKVCkhnhePlJlTuRjTwL
0gh4j8YS0y4tTy0Bzq5GBxK5azYC95Uc+/IhB38Btyriixgo8+lfdO6wSDKJtjNpy6XNVSfl6Um4
r+wcIip/jubaeo0GsIBy1EWFd/qJmBvJ+qcX0jolhR/d8e7HSkpbjS/VMFzHdozlMF6Q4t/KuPKQ
AtymwTYcYMQc2NIgvc43EBTzZ3ONVP8V3hhk2vHUBRmoGEyntiLmevadPQHmH8FXGCoiDzgtMsp+
8UJydhB4YIllPEZbg03g2kf/3rDg9YsAsBPFtpj8De4wRL1eZ/bpG2XRn2lhzr1OFFqhEiV3nZ5k
VVHqhdtaNjagLBb0RLc0ZKWzq7FwOqtePSo77Wem0+cakhYejJUKV/4T1VcXTmy0mcULX7bDegoh
4rrMfPap/w/GmQAeKYGf/ckvd/Rd8NQityGsISN29cNirhDhSuajCYPIPXkWekDeIy/WtNILX4eP
c7R4ep2Kp9vQw4uAXdjcXdfmntu+1YgOuKU438TL0uCNTGztL+gw/xcIaiK5zKmq+zDKMMBBjDML
cRQsEjuscXxqGigghh0z5hgZjYm7ITJ4+TqUTWDlvTlaH46Y+mFg3X/JzazmiMJzgYJzM6ryKYxW
gDEH9/2c+SF6qAfZkQ8YO1Gqs0K2M6VcY0xM3sWxTAapQE91/aO8noVvIhSrFWVE9zWS45rxo+FA
6C6AUhaSLFkDihjuvvjGN+MmPcI9lGitfjmNnPhFtja4nQ7Tq9+CGYIVgCttz5bvlLCgXcZjzdXj
y7reu4ag20l0KZl9b7Me7c24jVRFThHgGyXavWnecHXgdTOK4xRYeLVwmr4Wi7FckcZ7lGvMSpqZ
X+JotegmSNQsyxtmlRxv1Rl5uAuciyAg7fap9KeV3oUOPPAvoSksDmy+wtI5Hu1/BOP9rhW6qKMu
QEtAjwHSCRZnr052uO2fg3KnuceNJuWcEQs7I3fqEzEsjOwsyZjilsaSLEmHd8fufAKH7WUGZzD5
dQ6AnGFB0VzM2w315nSyM9oZzd4x+HqgPLFdWxu0s+yNYusdbTfYiAHw3qrqUs0FDjfQdfMBrdcF
UfO3QOBftpKNZSqiEKOF+dTActaZpD+EJYj6WrbynIH07csIgLTrNgeoa1HyK0O70GpcBQuqLScI
mtEIwGPsiCUcabOEu8tpGk51KmUK2MWwToi3KZdEKlJKsn0QXitfM6hcHskAhfeNLrg3p/4umbPE
3vmIYIjh3i9zuBbkF1SGIc8/dZwK3uz+ZHuZ5XwMyJYblNPJV0nY5TT7aB3toKX/XDpB6d9QTTUV
PHsb8BU1yDz0HB4GBAs2SusaW1AH0YT01sDux1FFFuRnbZF1dEMyio8cVrYUNQFMPN8gHgKUwKI7
7KkCoKC0ov8+Ye7Niul6AX+cUEHyr63AplErLUrwNEgQurW9jnSnLw==
`protect end_protected
