��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$Rx�y�<��wA�*;�x���@�̦�W�X�fa�M-$u����n~�%���P�$��W��kYَ���P7�?UMfT��q�6�U��k�>����~�\N�(�����X�e���/6U|)�X2pF�]$h���d.���9E�	�IN�f"�\��e�z�y�b�����Oo2�?�qˁ'�͜k-�K�P|����y:����3�l�d���bl��ˢ_�d���kx�rq�mh�MذM�`aS�.�DW�mS�9���Y��+�>��!��!�T�uOB���,��\L�7m�O��W���6����'���j)n_�I����2:��$�K�2�Sʫ��l ��!���{�l����.�j4�	��很�̢=�����N��s���s5���_�R�>����ТP .W;������	�"�מԫ�����]�#7@O+?�⡾�Ԫ���e�O�\A�	�ͼ���ƹ�d�	@�nQ˰��E؁Bf���|D_�%au�-�'���w�*%��"AM$w�*��d����l��\�Y��e+qFɚ�ϰc�{Fa�:�}���ln��)�������u*���P��0���({�!�.
O�0���ˏ�2"`+�Wse���*������>z�opX�b��v:��m<��ci�����4��ٸ��Q�8�F���:��.}
N��}�:��6��=kw��K]0S��2 ����W&)D@�+#��(��i���~ȷ�0�c��s5/;:}׷�@o���C"����w1�W�����V�M�M�u�������|~;�c�8�D���,/��e�l��� ��4��NO�*�]ڍ�52VhxmB�wEx��?E̦ֈBA�|3�~
"c5�\�Gs�r����ຉ7�_Ϻ�}�F���e�P�Q�Tح�";y;�!�4�����ﲿ��)�-�#qwW�9_�L2���1h��ur���bsĵ�2y�����8�,_K"*A���tr��.��z��Us-�i��-��z���;�w��iwҡx?2pg�<:��¶��L@yr�c�=��C��	B��u���F�f$�uV4�6NЉ�)c��ԋ�t�8�gLLT�$�o�p�_�K
3���	�^��+��X>[Ż��x�pT�"aS�!�f�j�`�O�0�Kɠ,��8����1�s���D��ߧЩ��;a�>�?*nP��%sѲ��^��8�ڶ���~������^�/�;@�)T)��8>��U=�qOp�i��sF�a\
d���@��dDL^�(G1�������n�h AI�;��~�t5:��!W�A�~C�G�X�M)�׳h恉WZ�x	�E}��n���J�-_@��?�f���
]���qG~��l���ЫC��U;�B�qE��C��^���B��'x�J�l�F�5Ao��l⦰��f�.Vߤ�@T_q��Ǝ�����Ρ�f�{��N~��O�0m�Ib�Ʊ�g:����g_X�`9'�-E<����s��橫.�}e|�EЁf�<����|E~�EWL�]3>�l��bV�jA	�a\��l����P��M���X�5ęO)�}����i�t�uQif�k�	��$�p�� �_�:�b33�d�m$P�*������{AHj뛈��r���"�������W�
��f�-}��9,��G�u_�Vc	�h��?��!�v����>�VM\j����TI߫�K�e�Yz�&����(�r�I�)�(B$�k��}waC�"�z��zc����'�=�$���.�&�=��= ���~{�C��W���i'%�5(�r^�M�����k1�b+E����[Y^B�)d��6$0��� }�,���z�_N9�.�x�<����m����������9�J�
3�k���;:F}a��9�6��>f���<̉����\��Ǵ��]��F�PP�`��xU5��Pd@z��͚L�-'��2�2L�'�@!�����a=��H�\�]�C෴�὆�L�O�(�	�d@�UƱֻ`GŁ]
莇�d?��pVrceş]2���g�@�?j�J�?F��D����#k�pl�zࣄ;	Fh[��H�>��t�T�n��dz�܃�e`m��Tb�-#Q�)%Əب¿1�8�D��H�Y��M.{����x]�k�vĀx~���柭8Gp�`�U��}]�ʟ~�6g�߼/��}&xҥ�L�݊��=N�M��9�H~:�-�
��5O�eO��.7�V! �Ȉߥ���KM�]�����M��Y�}�_�V�޽�C�1�ć��U�(�E��Cbg��Zd2�-�sO�+���p�G?�$[w{�"?�}3d��fZ��.�R�[3��*��?�{��!�tJ��ҵԙ+O��:�{�"͇]�QN�#1tWC(8j+�-<�NL��u����s�<r�!6`�Gy@ mi"f��)R7-����G>���NUufڿ�p��$N�U�3���9gP��~OFQ�l�I���(L��!���OY�T���L� /'A~��f��U�j_������]�U�q��s�@�Z�tFod�Vs��_��U���L�l�@0{�<�����L8���k���f�9k���?�{<#��C��9g����Bb-@���$¹��41\LN%�bv5����V6]�@e���0钄�2�t=���Jfy���D�t�O���p�U�u����w�<y�R�,�=��1�<�ύ��g���*�[�J{|�K�{X�E���	x���B���>a�ׁ�d�ǳ�i�xi��L}U��A0#�º_9u5�^�^�eJ�\��Ze�i@(tLŤ���խ��͕�o�\t|eݯȽ3���]�ѽ�<gEW��C+m��/�4�̱���Cw8��A��E��8���=��J�6t��e3K���t�e
�0Sil!�O��i�$�BB�-�ǧ�X�f�i�iv�׹?��eO�:W��j�f��X@��k���Ѱ�����K<�E��&��`;���|q* �1�丆[>K��_xΒ2�Շ�:v��<�ϣ�K�峋@�핚h���Ù��L���|������X�?o.��)Wp���|�'�M6�ga�Ls5͓�2@�x�/�6W��˩"t�g��{�<����c%�V�&Ƭ�S<�7@#�O�"�qB�F-��C앥c�=M-)_\�˒ڌnY��$)�K �?gм@���q4�R<.���0��J�/#�o�nk[	@��¼8�6��O�����=�x��g��=b��W!�s�B����.i��AE�p���BO4��ckD�R�uZ�(��=Q)�x����w�m�-aol/�v�Y�ԋ�%nۣV���dq8	P���6��;��8�t���!w�s���ٟh-�R���v�:%�?z>q��<�SӲ�,�S]�����yi�{��G���͸���?�QJ͓�aYh8��y��RN��i)���F47.R�d8��|t�"�J�88<,��ߧq%*����z��Z��퓁��YOG�p,X�����	��E�z짦E���q��G�{r���n{V_�Q�'1�M������1��f�i$RH:&ӻk9�s{o���(z�XS!%Q�"�:��>R�