��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$Rx�y�<��wA�*;�x���@�̦�W�X�fa�M-$u����n~�%���P�$��W��kYَ���P7�?UMfT��q�6�U��k�>����~�\N�(�����X�e���/6U|)�X2pF�]$h���d.���9E�	�IN�f"�\��e�z�y�b�����Oo2�?�qˁ'�͜k-�K�P|����y:����3�l�d���bl��ˢ_�d���kx�rq�mh�MذM�`aS�.�DW�mS�9���Y��+�>��!��!�T�uOB���,��\L�7m�O��W���6����'���j)n_�I����2:��$�K�2�Sʫ��l ��!���{�l����.�j4�	��很�̢=�����N��s���s5���_�R�>����ТP .W;������	�"�מԫ�����]�#7@O+?�⡾�Ԫ���e�O�\A�	�ͼ���ƹ�d�	@�nQ˰��E؁Bf���|D_�%au�-�'���w�*%��"AM$w�*`^��u;�^��4�kX��V��� dK ��r1P��
�B�Ӿ�'{w\���Q./b"�1%�d��"�=;z_|-��ʐ�3��u��<\�CXثj:�DL�S��yei7���Ș�>�*!V�j�#���^A�I�Ȑ�i��^�:f���W?ɑ<׫���b��O�
kV��D�ʪ����P:%��b�rjā�;��Y�����)s�&�|����ՠ����~@�;hIc�½UV�A�g/�ԷoF�*,>Ӿذ��^Y*����
�Ǧ�?�X��D�,���Ts��z�a���P�.���M��	tE��6�4tT��;�n��9���1薑�� m��\�5��kbA�����^!����I�.��|��^���n���
#@3G��#��d�C���\_�\-�՟'8@�Iel��a�b�y�w'�/��ύ:ѴV�d�Q��r�b��6��;�h,�H��\m���(��+)O]]�0��ցfVH,�$�\ O��z�2�VG�5���}�G�����;�=<��e��׈�D��nG�xȒ'�h��e���>��Ŝ�ݗ�6�ؔ�rL��(�ևBVFi�Do����N���r�=Ƥ��u��b�W�wX�*��t��4b;L:e!Ã��������E^��N����E��Ѵ������(ۜ�IVe�*EB�7ߒ��j�̍Oe��*��.��7�@�g�t�*��Ҿd�ZP�$�C}ڇ��!߭}�
~5u�«:�V�s��v;5�1r�%�f��d�b���m��-��#r����Y�04A�ɿy��d{D���ZK�z���jK�J�����r�� ܰ�AkC��cnQrY4ӆ��N�3�BJ�Շi�Sq����y�mbh�`�fӼ�y�J��~��8(`G4M<��4Nl�أ
�s�Uɥ��5��X!@��W��e+)}�So,3h�Iqݧ�5a�Hcq��n��cMX����K�|��~�1Y��WQ������k�	L	<ܝI���j�#�V���� �
9��5eL")Ðp��r^�Ҝ���΍�^��E'� ��w#����dy��V��9��]�l�׍��'�+pԷ�%�V'\� ���$�f`�ha���Voh�'���l��9�}�B�q��+z��*k�� 3B_F_/�wBu���&�:sbV���e�o�Q[��ߵ�w�o�C��'|����-g}8v<E��K6�GA`�d*hCO�]}i��p�
[�0��J�J$o�l�@m+��W/�� ���|ő�89�qn �y�b���
�]ϝo���(�6��n�����7;V�U���H/�^����(Y9���g��h�^�E7��ѿ�4�k�n�R����`?yn�!d��l�ʤi�]�=�����dR�U=�e�
�Z�^�D��/M�6����"�
�1�#�y����$��}��'v���X/#�X��/���_C*�*R�:��).��rPx�N�e3ՍEq��;L���d��j���QHݱ��9e����TUjT���$�͍^ �� l��vTZ t���yq�BuE<Z5���
>�clo��P�s]�-*\r?�j����i\Y|Z�)j�t�����71xk#L�����Qe+��bO8��C���<�إ���t��
��F0�o�3�A�=�S����#B.`��sd	�����Yl��CA|�0`���/)�j`r�����ť��.I��㞻�y�����S��t'�Q-�b3�t���#��H�ڌ�4I���
PU��讞Z|�	7$��a�lSSL����xNk����r�� $|Z���@�ZHK���P7���/����N�S/�����p�ݤ7�u�X�uI���df��Mh6C�2N�v��i���@?�^1i��\�};�ᎈ淍~�⡀��
KoE�m݌7������yv�Ia�L�X+�s�G⮠��55��MQ�8��á#�2R���lt��n�0���GݐGM��	> ӇP���]����t^k_�����imz�����h�m��b���E�K�V��o)��6�ӡ����&��7�8�w{|�F�j;F�<�Cx�å-x0�f;G�i��k�DIՠ�(P?d�x����_�����Q�" R��P���������ip$
�O��2��n��4/!��@em������J�y��̎!TM֓0e��/}��ADYK����>KQE����fؼ�b���B�0e{�y�+�<R�B�6��:5z-�N��ưr�eC�8��i�mݘ>)�=��g$�����:���4���X9���*���b�F���Hw����V��q����}q�NJ��ldh�>zf�[^a�kT��DA����6jS�}IP\���H�y�>�"��%/��C|�C/��-�E���&Q��T�U�nP&��N����ʴ�ʵt��Tt����tenQ�w{��pr��G�H�%�-��	X�;�x}�մ���ߺ�T�����d�H
�5�N&vaI�T�9ӾY�9:��hT� '�vVL��+�!�ڒK8N'��=<;����E�i[�'\�ܑ��7#���Bgobh���̏@	��#�K#��p��2w��ų����Ҿ���#~��'-p��q�w�v�493�&U,7Ya���&�&/�e(���}s�NpЅiQϨ�p���n?�K��"��ɲI�3 ����:�d۾A�~���.`AV�灋j̢��_0�����f8��:c��z�6S>Jy��K|D0�����Zj#�D�|�-�s���DH�ٵ�W�s��J}�v� �g%V��k��x? �E�xX
�����4�p4�O𧋖ɉ����,6��w��	4 ��1�ધ?�Xxs�[gs�(�l)�DIT��8:2"��>�ױs�P=$��]��6��Sz�6��!�z}%�1b�ڣ@�rW����Ec���\�a����"P�(���vY<i�
�y�ΨżҜN��y=K)���\Ƭ�.��(0E&{^:��Q״��:68<++��W+�_#�ON-����:H��<?zGN�6�(w��r$�ڭ�� x��*�	:�;�l)��=�	�m(��v"�����S@��&�H��cE��^?��rKd@}�-x��,��B���_�Kп����{��A�����xƎ	A���:D�2����@O���m�}ؾ��YHz��2j1hP�ƿ%ԣ��j���Y]U>������<�R��-�1p#�"��bS���)nN8;�!N�Ye:�e���D�f���,�ccv���s�&�.�H�D�p���M׉�S���*/���-2$���3����Oٜ`S!�n~���9��A��9�j���G�R	W}�%��b�
��YIrg���|F%�.�{>^�i��%!6���܅ɭ@L?~I�5�0�b�G��PIܻK����B���77�1Dw�Ov 	5�6R혧����gB��4�%�j��r��0?���)���d>c�%Q>q�@��	�`#"�ѻ�I��[�!� ����u�����'�_V�M���y��)uR��=/�<�C������&�ex�Q�����Q��G2=F٧y�����4�~2BV��ɞ�����"�� �9��ԝ�\}L�^N^��Y�':f����#YO�g���:�#UpC�T:��- Pɴf�^a��s3�y /l�J�D:��?��.�+K�A�Ư �rd �������0�O��~����~.Kt�$s��wss����b���@��$v=�B��o���g�*cz�fD2V{kQg�@]���`�}�V�	-ީ�����b�����N�o�n}i1�W�3mX�$��R��Vݐ�����bF�1!Μ~�[��5��Wn����Nu�����8��"�A�L����]��3ԋ�r�l���Ga-djI0�����.�����"�4��N�â��S��`��#0b����574f��f����
ׇ>Ь��p�N'��i޺�J�-H3��s!Ơ�ə���ŉ���o|������mW)�笳�������y@.��:�y�(�52LL��}E��"Zx��}\�P�Uy~��tw�m�C�R�U�� @h_�}�Wl��D�p~Z �&��ȴH�M�H/m�D� ���?m�J���?ʲ?���"xV�B�|���o�c찾��?���
j�(�I�2"�z�QU����/����&�m��(��0���R�*��9��>��
%�KRW�sA��W=\Q��QƔY��W
e0P�߷�����њ�����&^����/- L�.EZ�Pd!��K2��m톆@9�S�{��d#�u�+��"�"J$x|��e�S�]Ⱦ�&�����_�N�E|;s�)�:ߊ!hd�<0g1E�W��F9���<����(�$����N�CZ8�50���+��߉��~��򮜍^��7Y�ߵ!#�Kj�t	~���`�H$A �lw�?��;�]�����p�C���h/�Xx��`�x������Ј��n��5��r���
������{�	�:"'���'�\,v9����lHϡN��f��=$��CӾ:��Xw��{q̇��_��#ZC/�n���!�E��
m>N�y�j����Ԕ۟�Ut+_.���|0Ѳ�h?��?�!����ʓkrS�u.�؈yb�$Y53T��T��3��ASz�E(P+,��)1Pe�2�Z��O"(0!�p3���0��_E��tK{6��)!3C^�Њ?�����c��q��>��ԿD�����׿L�G�a�2���v�і�d�v��ϊ��&C#t�g���n�uř�M�e��PkY�G%E���%I�e|p���Wǋ�NVm�,��#�a�1V$t���A��|�I}BeHe���b���,N�g�j(>s3I���àZ��Ϭ��LSIۏr��C[��715 �0{]FB���l�&M���&�CyPPJ9�|��bOrhp1ֳ6G��4C>ku,�娟#��[�/@;U��}h�E"nHo�Q�v� |�K6>�S��n��y^6��;�R�y;������T���T%#�:�I��h
�-��2���4�g��d�2U[��9�}6Hc���k�����v4���k9W~��P��Ϣ�#&��7�rHIz⥆��"@����%s�1�b�T���,��~����P~K�����#����}ИY�v���@S4�I�i��	p;h�n�o��5�f���61��q+m�=I�^�J�Ǥ�c��ؠe�'2�-�	p�/��]7 �ΰ�Q2X.��$��z	Ae��! ��U�R�?NAЊ���Dr�Ҽz\v5������ \VyK=�ۇ�xÙ����<G���rGmΪ�h
� ���o������n���"����)+c��Cp>)����!��B#v�6�I�$H��۔:��粽�@�A~k9�@g��y��'�&�GQ���h������d�O+5((���  �����L�W�J�����ȋ��[B��&�;%&�X����x����n������vt���m��˔㞸��J��j�h'���~ Н��cg�틶_M�F�w3���M���W��!����)�VپJ̶EIJ'��6S�OG�DR�l���ľj�
�X�1}�u����N��b��A~�_�W�r� ���ܓ�B�����zOƌ��uY�t?C��U!񂇓���4#���,��Ӫ���*슂�̦)��~��M��>�n�f����@W�{;�Y%�i�����w��q�sxR����H�����˔�� 5��L�-��5	���5ֈz�� ���/��h�����Ѫ�/���u�E���x�"�g;n
}ւ��܀]
B_�rd�Č�n9�S{B�G��(���x _�Yg�3;ʱw�&2�M�[��ߤR�cpȀrw������Ӿu�*�*�����8Z�G �a��st֗igeO���4X����T1�V�����P�ޱ��^�71)�����-�[�P[��t�*98��v��ī��vͷLPw�-�Capy����v��"�
��t'mǣx�s�hF�@��c��9��5%����I��r�+�:�_�e-��HSڔ��$�Ůy�m�7=d�i|=�7J���{ke����vG?_	]c�?�ėկ�a�#x�h,�ۋ�f�;�X�B�E��1&-K.9���ڕ���K}Y�q6f�q���lz��P)�G 7�?v�l^��R��_"��8�I��� ����v���YI�b�sp�4`|'��0Xe�C�|���6��m���r:^ȅ�Pn�1��v\% �s>zF�r_�����0��|�M��tX��urt�>5�>"�`����q\�X�"ǟ�����D��5(�k��=�{��w����e����oh������0v�;	�8��������73�Q�%a��E_�A�p�Q�kvJ�u��u����p>-W�j�.h5�66��C�v|:2�T"3�8��|�$�cY$�N�4�Ґ��ek;�L<%�J���B��<�c%E:.�?٤�5���3�Cfث{�@ye7�X�I�N����X *�
���
�ؙTW���=c5Yf�Q�<'/��Ϧ�&P+�YYGE%�:�~�ܳә�b��o鼄�ݥ��"�"�=���z���]4��tʛ[%�JȤ����dҠv��lc��a"YS����>���j���Gn�W�Lp�G�P�n􀘀���ƩˋKF�lOZ'��疽���7_�=���Ƣg
�/�>8c{�%*DF���	yM8F/H6;[��t��s���L��&Q���Z\^i�J98����4Cٮ���B4�ڥ�	�
��O6�{��Z�S�p�!�-�|h9k�f4�j��4*��^amN���lJ����������	�3�++TO��*��<\)��?�Y�b�(�!g,%4@��WJг�Sn�j-�M2"�O���q2�/$����aF����"'.��̼K�r���[��V��<��!�m�Z�S�k[q�;�5���ޚQD��z���[m��e^�bz��o�F_Z!zEX�������;9�6���L&?/���r��yA��Nu%����y��ZN�&0� �Ǖ��[<x�4�S�eRř��=�G �[|�ƍ���������?	XT�	�f�W��{K����5��'q�lK�PN9,=�S�L
�F�r2�=%�>�A�}%�%��m�C�d��p���v�w����N�r�2�'��D1 �{ە�:��hbx�j~VB)�j� Ȱ��r�l�f��u;��:u�"�5��:�U��D�L!�&`1�����e/�P$L[8nm.!�u��^�!��>���E�o��@����̟B�r��l�$~Im1%����c|<'�����k0Q]�)�g�!����a����H�S߻���A�1o�GN��S*�Du|�!�_0�B4�d�y��]1����.h���W�׊'��IFA\�pPN�_L^���# �����2�n����V�Yv^f~F�t���-��K�%^aH���O	��$����zP�u>��I� �Z��i@�����
���Z�C��}f��n?�%Vz��4�|��@��E�1����¡9o�����dƈ�Sh�@�q���Dً\�zd
¬A�m����[=�䈻���I5!��V��P�ߤ�Pg�(a1K���΂Y�X�2#f"��` �+Y6a����E�N�*&}���X�dv�m��������l���2�������ę���|�U�p�W�2�A໬�3ע��˩��Ř5���ܵs6>�N�c�/.w��D����!�k$
��0ӟs���#Zht�I��O�	�j�q�֤>Bęn���{n�d�*G7#`R�T�7�X�%���x�FDӦ?4�ʐx<����ؕ2��Rɽ�
��d�tm�e��`h�݋8ط��V\�e1-`����5~o=���0�V��!y����� ԅ۳�ؼ$���r�p�O�]u����~�C�d��Gɫ 9]�
y7�eXM��ӌ�����N}����g��`c���V뭑P3[����_�Q���EHƅ0'Q�����1V���OH��Q�N��b�-��4��C���`��ח���)u����.����8�:y<��;�"�G4�&F��ߴg�q:��� b.]�EAm�a�������6������ۡ��՜S$Pgc	�R"ߜ1�Wn��zux4��Ղ�a�������Jퟧ^ت;����9۬H	V�Q�b����{� V��~�Ye�G~��Je�FnU�=q��4a��r-Iֽ��2kXl�Qr�`�����x����M KC
�����@n~�t�b9�׮���e��?�G?�p���#r�
��l���jN�s�{�&��?F3\�A]��f��$���Q����~�a��i����Kj~{ �9f� @�U}BTT�b�Ax^�i�4�D��L�E��Q�M� ~]V���
�0do��i�qw��K Ƿ'O��{W�U�n�M@���6�E�G����V��:��+�D�Yӣ�a������,��-��v������U�y���6`�T:+�ۅ����NW����FU|�h����|
̝Bbg� ��H����G8w��H�R�gPP�>�F33I-��9£��;�2�r:>���!Z޴�����a��s���8c����0ř�x_�}Pk�b�C
�����
EPX)
mj(��#W�)�ZFi���p_���.rf��V��+�pz���ak���]es�VsK��mb�������fC �|���BP,�u��9�	�����YU��*���Y~���c:�
3E�[$t������U�8J��s���Y��rlt��ǌ̧�o�4V+T���T������I-],f!�<�P�99d8�4��Ѱr��jX+��Z���kw��ԃ�������r�1;���83�]N�p��)�^���'2wO �� �aj�+�)��R�3�����#�Cq�Y�����B�[��
��Y���C��4�|�;���9[Tuo].�&n�� 70-Ɛ���;<����=ď&�rΣɋ�saJ|}|�59���3�G��P#)�����r!��g괦�̬Ҁc,�q�(�s��a�~yZ^^��j��v��|�l�
����*���Lc��_t���%���^jky0�Z�s#���*�`���P�4 �Wc47�EBEL׸}hщT7��͌k�G�*�T�UѢ-�c�@	�R6�K�����/�HJ�]�4)*{Ɩ�^�ɇh���[�b,w���/gzO�����'�c�jtU&	/qg���==r���}�Ck���;�a�s�d nW����ěsDc䞹�$	]��c-=MK G\�:۷����7�����o ��$���L`�ݍ= 
��/]�d8H��|��Ϛk2��*c��pV�E:n���#*p<�H3u�_����[�E���ah���R�ayD����۾-ݒ?̄7��S��թ�ø
G\���a@�Z!���M{�֤L�6^�p�hs�8-��b3�?|!r���#���"�~�	t|����}���~���'h�^�pdU�K��8�r��mxe����kʙ�P�O���r�$X�3�!�Z{�ѱ�ޏ��"�<�DE�:�)�{s�~K������t�q�P�W'��Uh�V���Ѵ��*f�fyW�E|�h��QzB��9r�A>P擂Q�+e�����b9��X\R=�t�K�\!?��~헵\
�����W�@"��K��)0�7�/8�i�Td�W�u��hu[��O��X� �-U�I�W�+T`a��΍����x�n�]8�r�7	,������*(����^M�f�4��
�������[��7�a��߾���V���xzGZ���5� �)�z���ɬ��is�Ǡ�e�%`���A	�w��!�Lx3��)2�'�����;E�$iX�)=�i2�R	�ғ1�>Z/��������>�!@[y��u�;5��|�tU�ܗQ'%`�m-��ёV�M�6ԟ�Q&]��w��n��/ �ځ7u����#,$bxթ�'�N���e"\m��h]��? �(�0l_�)F�nQ�`tQLMة)�^8�����p�߫�&o@�0�Ys����}��7���h�E+ϩ�}R$�5�pa�8*��['d���sMc��
S�Q�.ps�
�����U�)���>��\������>�ۙo#�������)!��^3��#��yX3�g��>ei�^����T�>i4�[VyQKy%;��
�&�Yh#�z?�d�a�|Bx�w]�D���<p~
\��k�%Fn�����*�~<�A���=�{ i�ԡ.�3l*����pDu�O��QT�U�x�08��f5�]�s�O���m>�M��
��I8���ط�n�Y�%a���
��T1�)?NG� � �[k:ʳZ0~�ԥ��c����1��ٗ���H���v�lNa^��6��J�\|Yp%�%FO��>zݥ7�����s7c'ԕ�eU�Bܨ����7/��Ñ_����p;-_@�L��&����ꑖZU��TI�at9P���V�aoArBRd�������7Yl[L����7W��S��c��?�@�{R���+��� ��2k7�Co�����=1S-a,��Z,5�=-?#^ۼ����8���}������[4��x��O8��b��Q�O��_ʫ���vq���L��	Y-HM̍9�0�I�XEM-.�#�)�����[}~8B�_�!�B^m~�!h�r7�/�ܝ>T 'M^��I�M!_~�#�׏�|k��c'���!�a�S��|�DCAxnZf- U����H�4��j�yПɆ�p%�9G|��t,A`���Nh`:�1�����D�����Ⲕ_9�����^�V�������d$�N۟T����,/_&�k&�q]��c4�^����r��=A��9���g��������7�d�c|C��M4ن��C�0��xۛ��䖺�L�m��7��1J���4��g(&'�ǒ�!ռ�D��o�B���NL^(o� [���U�?اP���qy8��6��]m��K���d�>�o����/]ȴ<��} ����)=��+=�9�l��J���	U X��y?^��̭��]�>�ݝ h�!1	����;��?F����QwoJkz��h���ܸj�����OU��;���xa�U�)RU~�o8�x\4�Ɗ�$:��7z�qn߸�(G�\��q������
��ǩЊ��6��o7)���!�������a*�?3һ��b���]a/��p��J*�nZ>�r��`�@��Z�B������Hgf�~����J��٪-P�8i[����F&@c�5���������k�ߠ�^�����9�<���b/�4�=sv��R�yo�~�P���4H�\�nG/�|�c;��.ggƏ���zY:Hߤ|��S���Q\��\��2g��TiX��?͔"l*����[�9
u���U�޽��a�QX9��܎me��x�j!��6�{�$����_C��dP��������JEVnn'�<��ad��s�z��B�ቓ�H��m�j�Tk��4���F/�k^_�Z�c[���0TG���+��fb�]�%��!K���K�����kb����a���5Q�����+� 
��4	�O� �J�R3y�v�q����Lk��XyR��`dF����뾼�]�MHH	�SA�e�̎Q$T�=�0��d����m�4�/� 1͒%o�����A�����e-�6%W��?�y�Fo7�4^��F7oL ׬�6���s^p��
��o��8�["��u��|���G�y�:n��2��1������h&�	�@�L٭ؚV�F�P`��E0TQ*���nԡ�=�Q�͸~;�&��Bf�=�����-����]�� �M^O��})!l�D٦�yF�����>�}��O��c��a	�þ��@��Լ˒��R�3NG
o(��w�UrW+�;J�-��vn�#lZN~$�q��yG�W߷�sb/Yi/-��lvI=�& ��d�/ǝ���&�O��H8�W�ܝ��7Ϩe�����^	��Z9��՗���7�:���(e�wT���x��{9���~�
�yU�+���d�6<��6�������<�����ӓ q>�c{S�d�-r�`KIg	cX�L�v��%@Hv��&��0$��Ɯ��A�2�G��҆0<���KAř/�z+%���|dZ�����u"Z*��'Q n���K֭�BA�GQ4*�ᴛ;�;���K�>��(;��D7���bƤ|8�@p;��6���$���l��$�2sN%�"d��r����gY~̞ǟ�M�l%6"w��n��̈́�`^�I��{ӵ�z�i?@%jd�Cz���Ko֑ȕ��d��Gz�2:�C�6}��5�7�^�̩���a�����������Jh�܂"#��/��c+�����!�Q#��Tû�"���
���u����br;.#ws�~�C������������k�S/�)b���!$D�;xfϪ$ܨp��0�i+�f��m%��B�i�&��V'ʲ����Qվ{���\iK�]·Q���E�@���dcadg�{U�ɞE��_��O�0�����F9Gd4�pux3B�2kx �:�;�u�������-��I]������SO�9���
�c*鏑�D���2o�ބ�Q����Cxfׯi�,��A�m�q��aP׎ςSA�V̈́�~T��|�/��g�U4�\�D_��鴔�r�
[b�cr�u�I-E3��<w���GG��i}�^
&ʂ��<IZ9�D88�g�� �1-T2���* lJ�.^�����R�nF�0b��W����4�M<��n��L�w�w�&#[�Q����<I��^A�  �&�Ǿ�l}� |��<W��5%�ܱ
���J�v垥�Θ5]o�3W_(a\���W��\]O�R��,WӦ:�%^.�P�f�t*EZ"%�+��r�ޏ�y�Ķi�$@Z���w\�{��03��!�,]6���#d�.��C��/���&�5INo���)T9��������睑�]cM,��#A2/�g� +0| p%���.tў��$�曍C�@x�ܐ@�2o߀� ���pb<G,���C@
j$�;3D���n9I�N���wCU(>N�ㄛvKl�س��/G�A{�e�ۘ�ބ�7�� �u���� Rr�E����/L�.I� w��	}��F�4�<�B:��[���`M�j���mȉ�K)������Ucˬ7m>�H��n���4��+�N�ES�ې�>�Y^h��a�-x�w<�Ea{�����/��M�gAE���ɘ��j9";!��sӈ����� D$$eL��-흨u�r�b���z�瘬~QGI�S��!݋Kb���Z3�W�����8z8��J��9e2�*{���G�+�3ڎ�t1�Z?��֜U��E8�-���H�bW�Գ���ӏ}����{��E��B���5='�e���i7སB1Ffg]*ۣ�>�PdX?K��|F�e{��MыQ
\�y�d�S��=�EI�4��{[��ˢ�����OmAHqv@[�}%�ue����z�dŢ�+m�#��o�)a*�V�r�S	���όd4�T|����a��hՋ|_]�w�&:�C�����y���W܊�_�M ��{��.�w~�V`��S.&uw���5����u���� ���df\E���D5Y<��mC4_vإ"�%�pd�2�kO�~m�fG�����݁[z���-ط��hr|�
4^���3�����y�P^�[��)ۺ��s�t�A@T̺ 9�y�x16�r�|p=�ĭ�̤t`pg}����ei@��#��;�b��x��ͭ� :���n���06i�be����ri�:�g��[N*�bn��ZmX�����(�Z�e�8:P�x�j����Sֵ�x��� .F���܆��S�}3�$�7�]�EU�(���9�^�;��Y�Τ$���صo�%.[�������Y3�hޘem��J�N�9��y����"���o�N�>Hj�d����*T��Z#�0؋���+K��!i�������1O��U�fn��k
����&�K!,����.�~G.pU����?�R=:��/8�c&?t�I^��. ��Mդ5����iM��Au:�_E�u�H��(� ��<r��h�a�0�Ǒ�/5�S��~;��8��8a=�]N��PZtF
y|]B�n^H�:%�~���'+2M#�S�ׄu�}
9���-��@����&y�P�կ����F��Ш�E5�������qT�f��@aPE��Q�$ +_�h-�b�&̲�ɽ���T�i\pqw����p�M��q�qCc=eJN-`E�u�h�?�"jPԼ�/H�iH8*���
�0�A�������G8	�/�^��H�OK��<�Z¶D�٧S,�ؿY�?��\�e���<��c#��Q�R6�g�3,7c��#����� �E���z�I
3�_�ɍ ��+��n����qL0��؋c0;#ץ:B�B���Gn�;�ȟ���A)�f�%����á����������-L�z����������Q�8��WW�w�BX��~������qf"��Gyt�(!�2#��z*`��z��ۆ��g�U�Y�,ȝ�)�[N�(����)���X� !ͼ'�*��fN����x��Jhڏ��&��Q87e5���4Z�9t�!�����a�On��9�b�4���:�Ґ��7d$a��;��cc�12]�;�h��o�n{)��C}l���NA�/݇7P���̝�R�I�	4���I�ɍT����;rBwr�!�Q_ث�x�'��vW����eJ��q����!��PY<�Y�\�wSH����do�_;��%�yTk�����D��Zxm`k��}���-/6�b�*2�ޮ�oc|J2F� i>:D��3�����e��xP�e�0�4#���4�x��j&�K��c�������Y!�;�ɐ���u��˥���Kp�ƣ�;��t��I�t�^�<�t���.��B����,��b�����J�g�8gn]ʫט�x��S�Vte���(`�U�Ӆ���� 5^*�ػ�l��HYƩ��L��ɜ�8�	#hʙĽcjk�c��]�F׻dj]!~��?���a���էFխO�����O��%e��o�W�o�4QjNf,��5�=�|���0�W�� � ��O}�L.#��B�`@ͱzW��QҎ���iS�øp�c�c�+�#v| NLi�p#�����Ϳ��d~*��_����X�BT�t��YGF?!E$�ZX��d�$�qz�l�;<����"�p�Q3U���:�;v���f��_� M1��r�����Y�Jʄn�^��(�Ш(b�����_Z�"�<,I����.J��(>Z��3}lL~��������hx�ns�,<�Xp� 	iQ {��\��>�s=;�8%�J�bV�P7?�-���5��t��>����U��Ρٵ�e��`C�Ѽ���0� tl���Ŗ`����4��֘���*v���f=�j�:��ζ��軅�,����Ԥ��ӓ�xc[����{�ݢ{���(
�?a%9(1v
Q$L4}�<3�P����4��mr����wU�6>�����n�K(5_��<�@��i�B��h	�NC'��aѱ��1��)~ܳrE����|H�Ov�G����z�υ�-�Ϲ	-����P�X�5�G�]�6����U�-��$^C���Zh�k�H�L�}��4�t�����A;�vcd���؇{�A%������ȓ��z��_�a�]���վ�����L�&�)����ߔq�3bbI�xO�����af�Y,��D���A�%�w��c7�.f�l�^㉭N4|G�e��fRLR�[�@@��/��Nx���ʼ3D-�_bK��"�(�@�Їd�����+(4��
�TF3���v���zD�m��1$p���k���=���c� 9C�'`�:��{�X�q���	s��W�L�n�_�T��-�]�:w���`�K���>���0\d�/S��y��_�Y�<�?(��v�,-\��U��-�M<�~!#�~����l�K}�EE��;���o!�F�y�#����r;`cRz��t�J5�M���*�灴z�D��L�$�Wx��(b�v�D���%"Xil�@���!ٝ�Q��N7�P��-vr����K)�4�ZZ�n�>.��t�р3W�D��A�<723����r�t+`bm�!�\��<��-���G���S�����ʛ��ڐ�:y��7f�Q�8����bY3x�=��*� ��c)[qRc���t3n�e*�9Ĉ����-QLt7��Z���6`�X��IM)�?�S����2b0ܹ�#�l�FD�1߅�����;��Dٮ��e��I��+��:~_ ^f���SAt��[��!{��f�4K�B���\"4��H����h0i\��I��=��m���j`����=3 ���}}9A%�믲j�fQ�i=\Hu����38�LN��Y�Z���A�`4)Y��SUH���䪷ʾ9������?K����7w�L]���b(�K��6�@�$��Y�׺�1�"��2;�/u�ȫ�����ԖY7�8�r��J�1�i�F�r�h;;��5�Y�B>S�"y��60�U*N߱fF��N�D}�.R��d`�|�rP���%v�fb VNM���\�f�������s���g K)޷"�K�.�u}������{��f��&f��yz��+�O�m�M���g&�:W�5
�R�k�A�1knk�'|=G\ʱ�C*a':�������MY��};�X���!<�J�1⨢^qp����1ڭ2My��R,h��i�����˓$��t��B ����.��G�}��0�8#�.:�EU���*��F�9w-ҕ��n���Z��\��Uh��K��3ǔj��e}�˪y��uO ̓� ��-��X�3Q�d�/��>���YJ�s��� ���Q��w��K&���ӝ�},���z�^sV$����埇}Ի�w�d�;_�|+C�	�c�ԋ��!��Y�ݘ��k\���wMc6hT�"�����)-�G@���W���YXBm>-':4�L��EQ[8E��N�7
ތR���Q��:��e*��旭��K�̓,N϶��cIք[ܿ�~=��M�|""��=�)B�oj�/4]��CJIq�y��h�����D�
�Aw�Q�\C��f��#�lvo�8�V� �R�E�����s\�ӥ���ܼ�i
�e�����H����,^��2�pM�E��S˿�N&qHQq��4�U<c+x4�gBS/�a0�������RyS���4��#�J�>��c�� �q=ג���_Ƹu��k}9Ҟa����b,$��A�J �;o���c
ۮ����a���C
� &/4��pLWbw�;/v�uI���h�=�c42���oO�N�䱛��\�*�i�+�2�a�5cj�<k��;�����`��Ie�I��l��w5����B$�4F�C����w~��%�ܳ8$��~�[�k(���k�̌��|[;ܬL(nt�W���x���z�:��Z_��1[V�����]���'&�M:3�]o%���2�\�ž�z|��3K(�ђ���i-86Vй��N(���'0��1o��h�O
;��Q�Qv��ƛ�
�`}�v�caUU0DВ�%����������T�½����o��3a�B
�*�����w������D�-������Ҏ�R�DP�<\uG�Ÿ�&��ݪ�����P=��	�Ql�:)�Kep5��M��S�'�ʀ���RC��� �A����;"�����"����0d���B�I�=a� iQ��D������ߊ� �����|;eg}7�grP�C��'�7����=��G�][�d���t���9��Q�&��/pZ�_$U���9�˨& 6r��\^[�s�g��	�4��~8W�����,��/��#ζ���9���m�|/��5(���,-n�S3�1_����|��0/m����yI�x�K��[e S��s:���M�*��M�ͽ�AR<š􁹀�˕�N}�ˡo�W���J���LW�Y�n\7��k�K�*����bL�Q.}�@�,m��Ni�**�A۪g��s�<gM����DO�����+P	L�������s�pJAoIN�2���~H���wN�3DjAlVM�^,^��i����/ >��N�,��_�7�G�����w���F/�U{��E��&+�����r��*았+�j���KZ�ڛM�vئR��99�Evr�7�`��߬Y ^]���렛�Ѫ8��2x�Z���?	w^���=�I(6��Ft�N U~q���ڀ��s����k�o�-a����Ʃ����:a�S4gE��6�-�ǲ
���m��)5K���h����_���C�/�	T�I��]W�Z뀔��?!���^�J�N�r�d����7pѫ7l�\�*+��d�-f7��QULf�(��|8�R�>6�����ЃZ'=��vd��^`kaB�i��%���c���7�\��?�Z`vu!���h�M�c�}�c-��I$o�U�nV�
�z�`�h�^��fa��,X�xM���6!Ml
���MeA�,���Oc|k�u�c���C!N��Z��AH�@	O�r�����*�
S����y-~������ (��Q��N��%,<z�ݭ!H�˪]�����Z���7䃎�>�g�:����Bv2�&��]��M+N4��Bi�]~d}>��H9N��S�۬��7���B(4!ItZ�gZ��� "p�q�}����b�ծ~��Ly�=�
3�M��HN�ܭM�S|j�O#�^E��:E������yKV���K�]S�0�ɥh��_<<b��u���r���^=rܭ��:��e���8r.�y3p�cH�8��:齪��@�O4��Zn}�)�7���Woy�r��(��&�K���샤(����d�����n\�2�V�\`����B�2�g�l��:-�A��<���8�l,T�/θ����.}
�R� >J̩�zg�py�-��]wZL715c[K�]S'�\Hf8��#�6����K��6�^Ay���k��qN �y2�=S�G����f�	����J���`,��qHF5��O�>�?Y=I�<�a���	�;�/>�a��V��빶� ��<����!��8+�
�J.d�㢾gt�"�AD����Ճ�Kx%Xߨ�����s�����7��7�aB���"�P3��h��v�tI�o �Y�}':��?�x�e	����;uA���
Q�Л��+�S~؁B�^���z7��P< |��8���@��6u��d�R���|���"��Q�Lk]؛w��!Sx�"�z��4`��v�ܤJ��5�\��ui�����DC�B�LhL�E������Oy�[engf����[(�5'6T�O��M�M%CY�)A9_���$D�}��oK�X��M���$��Q[:����V�Y��p�+OU�
#D�;����cFs�k��Q��2`T���Z�vAF��	0L��Ie614�;\�/��	Ō�=@�Z��T����� 2dvO�n9y�W�쮞�?�K�$B��#�\�^�4������PT��Ԭ����i���om�@y���j���`�p�s�uᴫ�~�]��������� �~�q�b�tb��qn�N��f�reo��f���@�)��qn����」��R�cw�\ݺ��by
�?���5�q�ƌ��,��A�8����SA�O�������<꽜���I^��̏�7*����a�x��/7�?����%H_�t��*^ki���#���ˣ��|��*Mɚ�_����4Կ{�iպ�*P)��l����OC+�s&�������u�7��S8�U��$c��V|�,��ײ�IW>Xf�iS��o�fr�juj;��5؀^�d=ƶ��?P{�<���}j��
fZ$����M�iN9�����ML�vlc&��~�� ��������|�N��׹�����d��|X2���K2��m�r��7n�3`��U*�@���"�BN�>�;F���'}� Z�@h����`r���������
�z�ܧD�@�^�!@�|k�\��FKGr�ܿ�sA�$-.h�X�CҖ ^m�i��F�Kr�T�x	�L.���ߪ�H�lC��|(��.M�������K�򿏢�JR4qh`��=��W�����W1��>�|�B�C�=R<��jl�zt��e�w�w�-���e��T�\�n�=�C`zFbȨ`��F����,�L�1��И� ����;�|��<�l-ʚ����DUl�f[$�26���"�i
��~�
�-��@�A�p��w,o�h��f;) v�ѕ����%��d~>l��8*$=�@�?Xh(Ix.�x�N^�C���&+�t���3.:�!E�+ߡ��,hw�fg�~�)��#�_h ϖƛ\dH_�Y���+��C�B7�IP�$����.��}i�T�e�ڜ�qb����C�a�Ijt�g8ފ3��o�e����5�|���� $�.��+F����Y7z�Ί�ndH �G:�o�T�����LF;�J�C��B@�C���<��'x����r�T[zq[{*�6��Gg�ozi�G�F)�9t1�ۮ���C�i#\Y�.9W$�
	P}	�qO�@�#�l��2�e�W
����5�:K�6�n��_�	�y��u�BBZE�]Zsv]�+m�����j@g�Q+kb�\鰝0Cm��
>o,�B���ۊL<M��^��ޮ�*��&],�4���`��G�ᔗ���. �I4��ܚ�s��Έ������G �sQ��O�|�.]�|1H���E���p5#��}^>R?@bP����$�OO�����1V��}�V���Q&?�I���Y�<��3R�J ��.a[h���u�`5OK���({���[h�B�n;�:q#xX��U�l *H�F����p�'�n� � 4%�L��r�(����e��dHm���U+��J��e~�-�1fq�W����II$Q��W$D�[P!Q�WV(��=��F��a�	�l�Cnj����F����}�?��*�f%������L��4��g6���I���P���ْ%F��	��c3B�j���JY+�$5;'p��L3N�ݾ�Ř�S�72��g
��|f�C�ĩ�o'l�w�0�P)25䗼(�����^ e�i��.�=Ft�U���.�?���aAM��SP�������Y�4	�������1�}�C��\�K7w觉��}xp�7_	$�<�&�S� ��)Q�9(^�Ө/H�d��=�g���sJ������-�[ʅ��Qg���Y,��b�f���01��0,_�
@7E���Lj�f),^�d��ZL���-�S��q�R� p�x0}��Z�"�\�������bw��	�SkH��a>��"�nyo��I�W�a�'z�(�E������*B�Y k4{�nD�%�@_9no�w���S��@E^֏��p[Q�g��,�^���$aىvD�H�/:Ie�w�
&��xo��j͢����#Bo���&���6�B} ����a�O�(	�Gq+�R%�	V��9~�j���W���n�
�а��WC�f=;I����˛���a�8��~�}�6sb3r
��e�.�bɲU6a�y�D���p*^V�T����r� �f��ŖfK�x B,[�-���6�p����Ze�Ðl�Xj�׀ԫ�L4��æ<+!��|�D&F�*D:[�]��#�ؐ l�<5��K�T	�����\�Z�ce�'�(��`B��[�R��'�_�`��e`�xs��ٝ��@Z4<Y/�j۝&�t�U��&���c�V$Y�l��,��ܹ1������QB��8X|d��L�d�ʬ,�_�u�2���羃�5�*��I�
���q�i��\7��k�'���%ٮ ���7>Pp��Rѓ��/b۪�2���� 7�sK˩��<��������Ł�;�0���ڕ:����kl�p��3<�V�ڳ�j@�F�'�ɐ����?~��X��z���=,�u��^����"��ZI������u��lvs�~ �TKp����H�U�˰�4��a�,#�)�`�4}$���D^{CĆ-	
������)L��o��V���_��{����gop���Ș]��;���k
��}�T�N�8�sԹK��@�,GpLaE{M���m�)_�� <��Rk �V-�{0���c_��pZd��<�.p@��������\�lT���`C�'����mx3��V���Wh�<a_��8�qQ�P�*���7���м��M�DX?�4���Lw�PS��+{b��hD^
˖�6��]��A�y��XO��;�H]�~�;�Z/�-��ρq�R4Ҷ4�3#���ԃ��@F��0;�䂷�;�Z����`�Y=�ؐ��#l�~�a��5��>V�T��7~���;!5>���5�#��TJD`���]|=�Q,Dm�Xk"g��-�F�[�~b�2�*k쀨�l�6�ϰ�^�����)#��'�^��� �Q�����Bm��[gѾ���>>���g�X����))h^/�_� �V4���V���W	/��<\����Zk"<	zd{��J���jC�=�c�)v��g&X�%b��d��~�5>���5$o�D��5&�TH6Uʛ+�!��5*���h���tJr�ܯ_�B��E7j�^���pcX�m���kF�aV�աyYU�v|*�Bb�ߣ�Uf����yk�Ҥ�r���=��������%��	gm��)���۶BtM��m�j�kd씞|�t��ր�(�cq���T��Ζ�Io~.�9b~r��F5��?nL�KUoMl�'W��_����<��T��?��6Z~/3*�4t��\/n��'CW��t�C�:�/l(͆��#�oW��;�z�W>��DN���	H%�o����ɋZ���䟒�L�!(�q6[��;�-pX�Eo^��sʌ����]%\�t�K��F��h�k�u�L�[CtEk�E>5��}�0/ݾ��b��Rd���Rd���Qe0'�]�P'-l�p,8���f�,R�01s#A�G
mE������wk1�
ఃX�`��\W�1����nz�t
H�ܢ�8>䎽yܡ���@:��B4n%럫nCz_�����[�2�e���=��Jl���ϖ$Πz�3��-���lE7��6/ZF�3��	��՞�-�e��π^I�9X���V� TG�
>A�Ioj�O����J� �8muL��J�K���G�(�dN;�=>T��MNݴho�nsi�e�ک��y��6(z8ŷh������v>�d)k���:1,75�A?���\�[�i��2Zg�V$�#}���[���m�!��Ep���_6����_��?�~�)'����/�z<-c^Ua�����F;\A��U��v�n�=�a?Pe��s��Р�B�]�s��-s��s؄��%��e�qhUڹ=��s�q��s,/���m�������4��)��r�#s]ꀞ	�8q���ͨ4N�:I�����@ꛔ�Lb�K�OD�P��Yb�Z�$"0H>�:`YCs�D:���R���x��S=��alZ����B�#&����Ñ����O���zֹ⪲9�@ ��^ ���
N��o�S�Ԫv�QgL��ut�;��tb��}5�<)	��޴`�*�$�tj�1�W�P䑡YӦs��"6�.J���R���Zn.7N^�%�L�Bmq4���1���l5;8��q'��a�Z������b/�F�ۥ�$m������MR��]$feC=6"�{��D�G^-��_k�}�$��P\!܇��w��)2�giJ�P��q�*(�]+��X>����!`�z�0@�ua��{��mP�D1�R�bW]�H�]�󎛶A��F��G���R�-�b'��C�_ܢP�VR'�ls�tX
�-�$������]�)�XE�ꤦArb���T�b�xS���ШY7==ռlG��*Ƨp��[�[�c�Jt��T� ܉:�zsq:�ܖ�R��?���T́y!c��UqZ{�D�gp�Jko�cZ�C5�rr��ϧ����C������ɕ�Ǽ�]V1�����i���<���1eGfT���+�����fŭVcE,���/ޥ�L��V}cĢ�P�� SB��j�a�2��ar��dV�.�?�>���~:r8='~Ɔ�U�N�[�.��	|�>�!�Y���D-e	HU��%q�ˋ �*��K~eAu$/fo��g9:w��/Ix��+��[�u+XY��h\���l*��J=�א{�B�W� q��%Ɏ��$* �ω�����qDf�b<��Z��/�o�xM�ur�%�HY�Pb��L�jR�	��E-?��E���e%��Y���Ncj�$s�C"�RپA���#���2���-��ѩ�zՔ��ףO�>3�o���Ы<���#k����ҙeH�������B�׵u����S�Lsf��4���-����j ^��:q�ܭ�@WoN�e�v�����O"����8{���LVm��Bo����	���r{���X��Q���$��I�8�|.?d��Px���|�LD&��і=y����0c�\�ِW�Yط����0��bw=ϙL�|�Ce�IcE� ߯ؽ���с�+/V4)@��$�_�E��i����&�k�f}[��e�r1v�{�Ҷ% �h��E�ńeٍ���D�����2�{
�B��l��s�c�(�x�*.Lv4�a��:f��!m`#�f;��lp�3 �
&Q~��z�$�����Y��:s ZF%��`$6���e�!;Dn����(�>���k���(����+BU��Wc�����|*�Hԛ��p�(b��y6����܄�!Tޅ�V���/�Ff2Zv�����.�i�T��Q�L_�|Ǭ?b'��#\�{1]&��C��q\�9���j4�f���4r��&J���pR#�紀��f�(e�@CB�T+�v�~$K�Ǫ#a�2S,DV��r�����D����"�ɱt��x1e�u���WX�z4����ZYđ ]W.�cY��wZ=�_Fj3\�w���^+�҇^d|�Ce���o��p�l����J&�2��fN9u/[Ҝ�Z�K�Z溉�耨_ؘ~���4���Ӎ&{��RA����_{f[��˿�G�N՟v��l,Q^�(�� �p�D��}�35|����z��nq _�����,����=f>�2Y6��染

��� �y��O����>���F���[�.K�5��*��c�2��N�I+��|�9e��c=٬���r����sXW���l��Z��R%IE� ��(��	�d� ϥ�Ba}��]c�r�nW3�W&\(T�:�zL�K����Y熒0�JǓ{�X	���|�K�5$�ɳ��%��$h�b
���s�S�k�Q�܏Ә�:�=j���.',S�k�3uMH�^��Y�2�Ňg%`a��I"C¶Z�<�`&�.TU*h"��U�o��l��u)'1P��I�>�����P��`�	�ʜ��J�OBu_l@����9��1L�2^-1�P[�����~N�U9I�,
sJk�OA��%���Bf ��b<vW�8�J�R*�}�ԤY�h�I�<��f(p�|� u�1���t��̅�[�+I�o"8��N�gV?Dq`��v�\f��rާ1���Fj&�s�����s�~XIm�A>Ps�^��<S�s\��x�	U�(mz
!n�bk�Ev,
s�Z�@�n0�7sן�yŕ��%���k[ۊ��w]���G�%ц���W2v�Q�&-���Z.F;�����)�}�yX���9+ߜ��ϕ=uAýẐ£�� �
�� �M�^�Q ��#��>�{)�nC�Z="����,�;#/v���v�T��w��,�d��V�,�|R�z�C�,ky�W��l��
V|��E���ʊ�|s�fP�lZ�ߓ7���'Z�T��,����3w��M�?$b��r�
qi���D���ȫ4��:��؆�����~����nZ��4\@]�����?%搣V�Nfb�bͅ�R�>��iN8���r���p�?+�]�X� S��h"������?r�V�?r�91x��<�{M� e|�[�zQ�U$��8*����e�b;��������!#u�؇�jc�H�n?<��i��ÿq_�:����'���o�}����b��_�y�5��mS���SZ�a�ߊuy��՜���V�����u���e��i�S�[!�S]n�缆�sOm�YL�qZ�:��du���(N�N�s����3��D���V�-yu�jR!�6�/0��c}wN	ع%�L������2p�,�l	�~jԯX�u�"�\VL?��?�	}q5�ʨ3������H(���W�bE�d���?��*�WW݉��U: C#w��i��U�1�\`8��+,KiF�l�hԶ�%�.}#` 6�́�jfl8�`���%�O��ϟñkg��!�%��K�{3��G�+��.��X~9Џ��ѧp���jgyu�{!)�:S�;��\����;-#$��R�M�$-��8	X���	$�m
�'����ӝ2[}=Y���ը���+����|�s%MtmS9mn3�T/Fp�/ϼ��� ����)F)%_�!fVﶂ�IT����GRu�p^TXe�Kb�
�>�F�,��<8ü���46�إ�*�`*��]~P�Ch�0b��,���g��'}�#Y�q�y����IA�gG%4���-��jg\�������{(^Āewɶ9�����M8��A�ԗggAO(��RT�??��-E7]-G�@�G�xh!G��'0��pJƽ��ѡ�^��J���6Kǣ����4R+��9Q�@�&;&��|��M���/�M<�0�(��*r�RZ�p#�lk^ΔX�Dԩ�o������p�@��y(V^`l��)�b�it�B�I�j���'ǾE)���M������nW~PU#�W>j���<�Z����Wb�z����#�'%�&=���-�����oo<���>�o����l���1�LH���-P�\j�#�C�H�h��0���7g�pS'���w8�dJ[����IvÀU�i���@�kj.�����#+΁afb�=�Z���5��
��L̡uUlV�:�]Qa��F�Ԥ�QO&�5!�e���B)ua��٘�yoe�-x�r?M�B"!<��y��<�c;�
a����\"��Ѷ$ω��pi S����s�Ǘpjd6�Y2ޑȍ�g�I� Yxނ�:aM�ܨ���Â�w�h�y��X��tZ�J����ڙ�,��.�6g�ƌE_��CR�B����`�(���+���Y��1��kt@�@��@�Sk��Uj��ݰ��U�KN��b>PM�$�7���5�y�g<�|�J]Q�>�ix��Q^��}���*�u�p��WҲ�]U48�?�hb�UHu�24���σ���a��4{�]�r�8_1{��T�� 	:βͧ����4�|X>!���H�%�t�E��oΣ�L��>7�W�s�=�=B���|$a��U6���D��W7F�W�����y�y
��_NV��E�[�zw7]���t�pP���Ɩ?�g�t�8�6�I �rn�Rكnv8K�$M���10��g���Ÿ��Q���e��j'������&-"v���ῐ���ʿ�=�o�^��J�f�=� z|�x��f!��6���\E�ΎL.�	"�Uϡ�4=�UXi������O�E���"��{��������@_,�B��r7��;�&Xo������H�m�ۘ�x��"&xP�C���m��ƫ���g��A( �Mƫ��F�*�������U��V�<��,\�:c�8W;�f/{�^���n��W����V�mݘ���������L���kЌ� �bH���2';�$Y�B�Yii�w,�.7�ٷ�..i���l���S�\��Т��H��/3���|˓�}ߩ�FG����ț��#1T��zFVE��ofC�7���u���������s�^��*�aa��9��Y
����Ӥ��6�n8��}��4�=�Q����n@��<�WUmV��ӂ{���W)��ݑ�^�S�A`Hz��p����pS��$�c�-w+Я�u�Ƕ�����T��n�G�W���ߺ��v%�[{!C���1����qc6�� u�k�����N�r�xRD��$�
��/�_��<��{�sw�c�.�,�k�D_��P����$���F-/r)V�Φ�DW���ɰu~Aĥ�A�I?�b��JM�\�@��W]�QcT)<��B$c lb׋�p�kBPb)��#z+�NR"�a:�M����^�c+�V+oاT�#Jx�O 7��������sl�1�((0N��;)�g!w���k͝�wb�e�={����
��"�Ɗ���I�$�));�#����s�!�Y.�2��.V��^(��᫴k:�"���J��	S����~�(����ߙ�%�zj߯膇6��oT.к�)��KL�PX|�+_�a*O)s�?�-%����]m�In/����A�� ���:t�\��Y��䲐.FH�};����;���%��i�m�h�Cϕ�����x������0�X���!,��Z�2�\�ZAٖ �qMz��5@�uĂ�D(�T|7$;3�Y.���:��@�7P�mg	@�M��O8�㳄6��ޭ(8pN:n�9�MQ�S:W���P�U����%z-��j�W2�=9e��忥��"=��.Z�I�b\�TfI�&�@C^�`���b>�*R���}�\��J?O7DS�
ޞ����G���)����Q@�SU��n^Pq���{�̙s<�gR��F�_�F�UL�8����)*At�܊]�lf�-뻺�l�{F���U��#���j�E�LA�G����\Z�N�g]�|}�8E��b!����
���XA�D�v��Nl4���?[%��VU�4���Ǣ��;D���1���>�U����S�y��|'��w#]m71Wԏ�G-r�}�����@����+�_���gzJݹ��K���#r:����ҡ�R5)v7>m�c�g_#6��ve��6㭲�S`����&v/�2g��yq35	!���=_b�7����g-Z�p�<�jQ#㔵3b
x��Kr3>A>����_J|��|H���O�>��?�ݻt�H�}�5�a�zQZ�U~E7���֕��mdЉ�e��`D�"��a5������ R9�]���v�ȥ(�Y~���D �Ԏ���ϳ����>7����7~�� U�����f�����g�Q�p�=c'�=���;v��U�G��äނ��~F4�O��:,�j��������^�7DE}d�SMb$�S?�i<�7��N��cS`���?j��~TWf Z���2�,�R�k$O+6�E������%�|��a���x�Y~�KJ���;� a$BN����D�d�M�M��yу��Q ������a���:�O������ΰ(;P0�,���v�v�	)y,o���~gY�$�ړh�5�ޚ�9�(b�5jh��\��8�j���6}���Ľ}y&;C�c[���o�����ڀ(iv0�)|Z�CYH��O��o�3ɬ��E��mv��iՌGG���kן���|N�c�Sr��$Q�co�9����ɽ��7_F��K���dy����Z�+ ���v�@�,���\�D��@��G�����l���wL�Ÿ-��q>gw#ʕ�f��On��m�6�bݖG}���Np�p��@����.Ɛ�IpF�.�C��2�I)EdL)Otq��%B��|"��Myx'���[[튪��  տ� D��j,u5�+���k�!���d���EP������`nG��(�C�)cP�6��in�mسֱ��T�_H�r�� �T:5:�WP���ղ�(��Ԥ�u%��R#������c�D�5J퇗[@���}F1�߾7�[U��m������&Gk�wK�^�Y���m�X��t��$e�<:�ͣ&��3ڤ��i�Ǩ�[�V*���3j��(�h������$,@w�RP���.[qvAxݨ:�%9zqaL�-�^p3m��������m�& hvʄ�,Pt�5;vF�ck��LSl�l��`�O�C����n4:u˼�h�Ȁ�}�u�͂Y�>D#I��q<N��D��o����p�,�H������[��W%򌙚!{qY�M)���T�]+�鱉s��ƀ�p��嗚S,�����őI����V:B����v/������ĵ��"���Ƥ�������!��g ����MX��0�G�3V2��4&��<l�'�s.#�AS0�4�]���8o(��U8��ϳz���}|m;���I~��u���d�Qr�2���3�L�X����cG�[91(_��(H�x���*������\$�Ϲ��DVDG+,�V��c�߭��C�,@%
�@��d�9�jJ�Qf1>Ό��Zӷ3&��b����yz���e�0�t���M{�m���Ϟ�oTA���4<Hǹƞ��֍��E�I�֙�|""�<_&�w��d�JG\�K�s혱.�8|׃Ih;��-��_]�� Ԩ�Ama�\�����-<��4dj$p��-H���3ʢ�#k�`�hw(�,���{��,��Z2����-_N��:tͣL����`rށtى����R��i��9:>$'�;��y�L�V��!��9}TL���Z�b@,{V�1�Y���R���o1_��]t���Rnޣ'����#7�D�ܧ~4�q df�zٹ�����E}���zez�T3l+Ip_3�H�w�wgr�C�t�k? �	z7����;/�p����)�1urHG����ƩIh+c̊��L���a[�E>vwq�2���'�9;��#�qs��ۣ�^י�o�c$�_7��_G�wX���m�zܹ�f{���H@�[\�b�X��r�*�YA���f:ݱ<?F5�(����nK)�r�lX�B}���I�MB��a�@p�JN���I���h$�޸)��:e�+ϳ�����~9�6f��5�i�L�vz?��>m�[ʋB�(����p�TG��C�7og�������cH@_�p�Y��iY'��)S�jx��Jφ�������p������� `����%���:LISݸ�e���g\k�̯�cA~b� b5����͈$Ob�� F~ܿi9^G?�H>��su�3]�J��។onj��m�5&E_e��Z�`h.�O�J���b:�d��	��mE# ���]�aU�����/n�u�쬄AI��lgq�!�Yb�g��7��̤��������q�w��Liq�ݘ�0ֿ�_k�]᠈�tT�K���92Z��d0�Xa�xq9.� '5��7�<�ErjI0����s�Ӓ*�u"<XΘP�k&hY w�F#�O�@�w�aB�X6n��'z
:��:T���m'w.�5=�N�S�iסq���\`b׆!Gi7gI���"ސk[��i�B���U).Z�6>���d�m�'��"��x�e>��w�n�x�JT!j]�+�3�Ux���RV�;�)]�H�G~�J�Q�e#6UHK"VٳѾh�1���J�=��n��D� FM����e�]#��SM�
�>5������^z�7x)����M�����0!�sc(�p�1��l\� �u����	֐�����?4żT���"<EX[��n�g�^5�띛Z�`7i,M�3�;���yq=q�
uO���iu<@�lc���0���Ut��DEa���AE��&,À�u�ʕ2�0�g5P��_��]ا[M��j]be1A29�����m�@��DQ|bl@�]�~�y��<sЛ�߫ښ��*mdu����)��!�_5͈5��d��w��~�M�r��2�T�A"y 76ݤ�LWQ�= �K����`/������
-�I�i*2i���' ;�~���V�5kހf�����;<�/�qn�+J=�\����*�
J;"�9�m)B���ǌ��-�De�R�{^�\q�/�e!�K¯���kՍ��HPGW{R�_��2w��]o�QFo�O��y�~����֕h��W�a.Y�̠�A����߭!~�1��V�޻g���h���\������ �	ׂ�T��7����g�\Q]Vsa&Wk���0 '������%,'&�>��r�_0�u,Y����˨$��f���UeC�5�4�� �~aF�H��HEo��&�*AuEC[�E��Q��$�c�g��0���LC�4C]���9�!'�����ܞ3�O'����~x���l��wݷn,��ݸ�EY�A]�"���
o�7ǥ�g
�iԈUL�Eh ܲu#��