��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$Rx�y�<��wA�*;�x���@�̦�W�X�fa�M-$u����n~�%���P�$��W��kYَ���P7�?UMfT��q�6�U��k�>����~�\N�(�����X�e���/6U|)�X2pF�]$h���d.���9E��WG��L�X"]�Ad����ľS���8od����e�GT?y	7�������ݵ�^��R�q^]�鍦�����s�ae���h��L��P_���ާ��YЭF���'\��68�b�[����w8�[X��V�F�0͘3����q諵�uW� �h�u\V�?@��_6G�_�*�G���B�絉�f������[�G��U&�����~�F��AׯK1�`c��[<��FY���4I� �#�G��x[X�=�Q1��`��R>(�w����R�O�?����7�,(�H\�#h(W�EH=�������yq��Ѿ��aF����:�U~m<|��.��0=�P/���4ǆ���T(���=�ըTW���fU-_��k<8Q�����{�b���������.Vb��+wG�����!ln���2-�䪕>�в[u���n�7rVr�C���.�$�K*� g���Z�z�
�	xXZ��K�Pn���ɼ�nx����!'5O�N�t�A�G���B�һ:�e�|x
KQ�p]���y���&}�	�Lc�MK>d�>FD�5dKZ?.%K1P��!P����w?*��/�/rg�Q��	c����&� /�&W�r�I˲��@�Q��2�Z��sI�DBo�f�X�a�4�(Ъ8'{���8!��+XC��M����+����m��HD�	(�錕�B���kF<6=V�
�J���BI�ԮwA�,;�Qf3��6�w^�!Qw�I��Rg�bu=��st�a�G�+�aq�a;E]�[Lx�
j�O�E6dߟU�����s���[��_V�}sy�*�&�<QE�?�S����r�}�kIM�����!�eF��A��'�R��c�(7`k(�.[�����Ov=[���^G�\/.���g�L;��y��,�/o(s:urGָ��8W��սq�1��H�"·�p�U��j
 o��'���}�`4'j�WU��8q���m,�O�����D���A��y4�.W �����/Ly.�'��:v��S2�@�:�u=�9���uޝL2�7hz�%O�6A��	f�sB�`|u����C�%� �'�!�L���c��Xv�m��[v8�JnlH��q�}VQ��㣧�.�k���W�F}�z�{��'.�ۜ��L�^�H�uw���i����O���8k�|V�3�K�^�u�b�K�{�'�{����!���nF�9�yg��u��'?�y���lHr���|g(\a��*���N��Y����s[���mQ��RɄf�o��S��薿cȠHsTW�b�8�h�.��|~�u��(���U;ռel[�NM"ɶ%{G�qV��Z�9Bf�HW
��p
�d�B�y
4Z�*x���/Bh���]UW��;���\�5F��S0L�C�s����OxҢxi
]=��w���~U���P��h�Sf'�芇�,�<u�d$t|L��&�^Q�#5��'���{yV��-|�W3��z��}�7{�ԑ!�-�|�\�z�L4V�È�[bR��K��$�/��V7�O�EP8�a9W�*^9g}�\��(K������N�
�L�U�x�u�X%�r��x��i	�-P�(P5�4�7�-O?��r���SXW��9z�};�ny����C�S�
;Z|��~e�Ŀ�'�(��E�j1S�_�u�-(}?R��agv�PH}5i,��%��4�^�fZ����Qص���\�+T�Y,�z<e�{�����Q�h���-�W)�RV����܆\����!�+�$1�<y�Yc� �'����ӵk׏�����2����F���㘯����m$�s�u�� V�93��7��B�Q�~H�x�)0h��x�wn	��%�۞&cYS��t�NA�P2��8�b����k�y����^`�w��k�!(�<m%��ٱ��p�O�s*<�/���CƤ����f�,{��ү�L_�tm�S��N��=-*�X�m|F�!J�{O 8���r��m�z�/\{8�o���(L��y����Fs��4 ����9w8�C�l���/��ԽQ�n�ޢ��Z�ē���$�@�ѓ6�L�#�t���\��
K�2,�[�1�G$�M�cڙ�Z��" �lNh 3�P���uۤ�X�?�_D����8T���k��I�z�./�I�A�Zp�h�E�����m�P��tz@K�P\9��=E��K9z���Q�B��
;�_�0�%���x�����ӣ�;���W=�!/tD6T�C���G�H��+}�@�h��xX�q2��#��P.Nn";L�e����l3�La6�([/�!����*K$��wE�f�l(�p�y^�ǺH �Š1E ��a��=J� ���痁���YF
�R�	�Z��m_��S7VA4�����k���i�	pR�����y�c���X�n����*_̎����Q��\ߢtbh�Cց��-]�s#t�F�3OwM�̄_N��l~�F��go�Z�\#���@��o�h1�[��6P��/���Q���n� �N��H(|� u_�p�-gqޗeC�Fi�9.x>��Cz~ K�^��9�r�)��㶜���~]m�M���D��������Q;9Ր��Y�v�i�u<T@l�C��A9r'��W�b�uA��Ȁ�㧱��\�N�!��G������6�v��X�~җ�� ����u�*�%U��b��h��g�?���L���JYt��x���"T6(cy��!ͮ<�*��N)6�q�)F#���o��\cp�9�,�SDp�>��-�B��I�d������5�n�b�$�V�8Y�Mp���+����� ����<�2���\q����F�v�nJ��=%��[���O,�h1��u����ȋ.��\q�&����mHZw���ږ��NuM���Nw/��>�'��m䮫p�Wf�0-/0���8_2�MH��H�<a��$%�K�6� �NtV�f$
���B�>8��>Pq����z�6�<��kƚ�~�i��lʄ����]��X�Es'

cg�6��
��&�@z�jk�>�R�?�����rh�^����XZ`�������p��\�:���)P�s��8��>�!���s8w`�����xg1���|<�`����F�Ss��J�;�:�^�������/��;��ӵf�����eŮ�L�����C���fg/ϡ�8h ����4��$�&.Z58Fd��u`յmw%�$���CR�H@F>㛘;�_��讀��
?�`�gW�w���M��"`�r���81i�YY��c�wEDϢ�lJk,����ޤ��Ƣ&"$�)_ ���.�{�Xz����O��" D(��e���]��(��o�ߟ��puh�]D����DAD�����4~\ �K�g�955YLnH�TM��=�`x2���d?۳�/�qA��ȼ����	�1��s�S��8�a�[� �P���Q9
��\�Gt۴%�Y�
�%�� O�˼�Gl'�GRp+y��en�N�G ���T
��8������]�M��| ��J;Q�ܫ�|�X���D�§aQt��G�&�&�}j8v_XX����#�oڂ��k���QYY��5:�o��6����,r��σ*�`��~�����b-�d�1�󗌪����<��]�ˤ�W.Vͮ�ea�L�ݐ� 6�ξ�W�;ã1@Y���m�Z��r��N�9��@�WHW�z�"��L ���C�淍��T���Ѝ���'��d6}6�0bC�oȃ�7<������Xl��֘K7N1�1��&�Z0(��8ہ5G}���q߆�o&��J���_ܣ?�JpE����D�>k���P��dXN-\�)s,��*��Jz�J&�3�!w�>�P,`�pe�nh
R��*�*��
�ABhz0��j�f/2n�M�-l��&C��v�'�ӏO�6v���+(����������d$Sm��8[��Z��j�|��� .��K�6��\j;�,S7I���Õ;uc;��w�x��<�~�9�����/gR�bU�Frǀ)6��B�P�³.?�KH`.ɈXGD�).�ݐ/F.�c9|���&|��n�4��I<WY-�XR� ��v�|���%'Us��U '��.�ьDĆU��t��T��j��?d��%Sh�K��8��bb�����|�`��Ͳ�'F���`IG*A'	iҎvy�م��}�������d��'w�rڱ�f�Mi�͋��o�%'��ًuL�س��.}���y����'c���s��Y.����M�k��*`,��{��Y6��n֬���/�%X����������0�{]ќ���P��)��u-�_I}�\���ِ&bLv^۾����=�����!�V:X8��}}���a��:�"ѥ�����{�V��U��mg4��;���&CT�!��M�S8� RN�$f iƤ�8�N,�Z9 ��`�,����gc����ZԊDt�~��1|��}�]√��Y���L�,e��{��$΋(hf:}q�&�]_�50���g} ��+���*����#i�N*\=�e�a��v}h���pi����]�����[3Kq[��N����u��S&ּ+�/YQ9���z� �i �ýq	 �v�s��r&���b��?d�������Ύ�``�H(�݊�a�'���WG�[�G�j��!/��x;� rUA�[���J8 ��;=]���]�}?��b�GA�>�� �@�Š^Ό}^�!�y�� �k���[V/fߠim���q�q�@ҝ8��3���4>�a�mj�]3���:dzjDYt:3+�@� E,�W��U���+�SlC;�۞"ję�L�T���W�F�>�}L�꒸ݗ� #q�m7%���Jr �u���?�N��`F���-M�U��,͡0ޓ�`��ss�"H�"޹�`V�g��J�cC�;�H8��gYi�y���8}����T{D����ꨎ��zi�_���H��IB�B
�{����: '��(M,LlV?t8h~6��G6ªѪm`�v4��W���^H����wU�Z*Ч��3����ż�!��O�$��m��EY������n]G"~$���u`FO� }�m���������d�����Y�.I��[ٖ��Dn�����,7v)m�%��J��	�~lG�f���8��l�S��ߧKDY	3���'�Vټx�I�я�Tq7���`ո�:^ ݊��䎥?�8�C��52��`���ē������eMEv� �����r^���g#reg����Wp|/��$D*M͋%�i>)�h9���0��$T��jÆ������� �L�g�y��[�	��h���+�aܓ@�%5�t!�y�v^Aw;�w�0�e�N�/�} q@g�ݝ�M�!�.�i����:�L�q]���*�Dtc�&&���[9NQ=�zi����%x��>��q=Y� ��ȯ�e:��s����k�m�뇠�w>W!ݞ�=��S8��.���6�㮿�Ř��}��QM�E�)+�=��������j��Dn�J�[��H]�ҁ���h��A�l�i���S���t��|p(6�0�T�/�#���1^ya����X �$��<�+��k��]����`����ڒ7L�E�JX��8��5�RU��r�B�w~�y��d���wÚN!/�$��z՝�~�^}@��cM��W�كh���U�`�QĽ�~���ncF�����*����帒�������w'�%����$˦��l�:\�o�%�p�+�̲]�ρ"P� ��п]f�p����&�k��D�����+sgz�9_��(5�y펯�eKS�u�o����k���eYqI�u��]蜎"���i�9��NҀ�`��#�bnŧ�ZF!M�wZ�'�K0��+x��K�2����晢��ˇ-��5� ���������F�zN{���-��pr��� |��M�E�3���ro
�Ӷ��a�l��7�/)P`��+"��s�?�������o�[^�wV�ȿ�]6��r��k��@�q���B��y��I~6��Ҏy�=��^��F+�����(��c��.��z�!s����GO��R���ގ�e�ø�պMwoǄb��rbJdB_�`�Jz�!m$K{q�Uq��gz�#�r#y0��LZ���4�\T�7|9�԰�E�����^��ִb,�E�l �w�����<"�+��^+�J�M�[@v�� u��UM��d�}�M�w�`�]��l��|<5S�CW6��I�&ۉ$帨;b���%///�gysF8Am��V;����v)��� ���We�{L,q����ٺl��td:T�x̖�`u0�ҭYp�%4��d����]4���hԇųw��f/�|57���,�R�^W�ȍ�ם7��f���s��[�\D��
 o/���y��7)o�щ����g}y�	Н��b��g�*�|���@�y�D!��︂���܊o015�R�<�2��
�i1���yN�N����@��^���Y�&F4<W���z��z��ӳ](0���ð�ֵ���U��*���%%0B�dVnH�>����^���).(6``	r�E���
�&�S�]F<���oB0�('pOX�c�*^�eqܳ1as��N/��������+5�<��X�""z�s�JI�i*���a D	�y�Eߐy�����ګ��R̀<�v|��T���ȴ�ʇƭ ��vZ9�^��c�,��B��Њ������`�28*$�%�[bQ��DA+��S@�����*�[�r�r�����0�RgT���6�>�&fh""��
�-�	�_�����c3Ua7e=�D�4� ���"Cឆ�Q�a"��ݦ�S@��,s�|^\�R����I� ��d���Wa���TV����DF�K�:0�,��#�X[���sF��ї�;�hi�����C���ǣGqp~�xH�=m(��r��akczQ��k�\C�8UH�ER���}у_�X�D{���<�q�}�^@���vD����[���<iܑCj���"�F���d�c'��{9�4���su�[i�\���#�A}v9�S�.�fcy�2��~��mxC����������X5�m=T����!�?�?�ӏٌ*@TXw=��E�	L2ó�r&R��IJYp�����2b����w����r4�c����?�yIX�خ G�Z[)���[w̩�{����h��>���l��D��x�"��d����0�ƋAtG1̹Ł�^0�X�ES����B*�r"	#W8\c���Q^��'��}�v#��$LTiiJ�2UU�à��%g\?9���t9W�U �g�<�m�)�`O�BQ�ڐ�o�%�@6�n�E
��,�-���`�o����<Λ)!l �ԕ�3�V��̗�WLS0B��`�bk2Rj!2�h�E�8\��Z1�B%^�յ��"�ƌ��5j%���Xyr�fo�N��9�����p��1k��+h�k��	�����>6��{r�E3�Kj惎k�w��&U��˓ͱ5������B��xo
-1u)�V���M���Ć̜�ea�s��C���=������n1әL�#��x���bY�pš�bu8�婱Tp�M����V �j������ �������W�H6y�T���-����4�=0�c�݊���Z1���I���Fꇊ�cj�p\���t�>1���.ʨuL6p���g.����0����}�����ws�+)�2���Q��p��C,�m�n���n��18/D�A"��b����'�൰�͌2p۫d�g�w�W9���e��E�r�I�PD���${�晜�R�����r��tĜڐ^;��\���\��N�a�BUH�����ˊ�� vg��w��Ѽfw�����M���|'���-	�y�@kJ�A�[�^ܾ����3������S��C2����e���$�(�D&�Z�X�㧧������T��lx�/��)��ui�VY��V�bl��<�:)�j��*#t�Z���z-����_�ԙ�ޅŖ#p���AW����t*V��Tχ���4�o�ٸ�W����Y�j'�y'!�]�M��I�,}K��ϟ�����IVԽ��g��HC�������I�'��S���-

ɜCC��Sa�L.&��vP�fJ����!J{ϱ�l-,2���)�-��)���yJT�k�}j~�<6Z'|��-E�g���A=�����˾��@C�e�Tk��r��o3�H�g� ��4������E]&��Fͭ��V@�	�`��1bƮ)_"L('��h�/�r��5���9?D�3��|�qF��9����[W�눉@C����?�s5�q9���8���aґ��fX����/�2��%[�|'fؙ�D���Z���?O�=�(�Z���7���N�RJs��p��`x�-f�rۧ�����Ȼ�Đǉ���^YoK$�hT`�|3��6��+����-���=@��%@��쉢vǍ��������e�?�1+���ī�/�Tv���a'��T��7�� �a�YJ�������(z�k�}'�T�Dmq�)�#:/Z `�@�����݇N�]���2�I�F)H=]��T�$�n��7�J�Ɋv\(�~f�C񐬖�I�4�q�+���Y���:,*��Nӌ#�u����?�d l��QRM�g�'��݂Z��M��{"�a�o��B�J���K6ISA �8��^��������[����(�8���"Za$&�vf�
�����3R��I�&Ha��:_ث�N��1��.{msn�L��[)��t�L��2Г��Pf
)�����s�"�J�1���ػ��2�ށ��(�70W��~"����R0K9��FE4���w�d<��������b���%L�/���+.���T�ET�T
+a�U|W��C�~�q�� ��n��F�F��+f�_���M1��m~S��D�L�zf� ew�|O��� ��d��|�lκA�ji�3��h��f�1m܀H��s���>|��bFK�.3�x�}dt���B�K������'@���N!_����}Ħ�'(/���������)�T����<g=�=𣯡�r~jҡ�%l.l�K�8g�\�*�������T��ا�[�BT'$��6��`�aH7}�T=��W�[#�jiцM�0�>��',
�g>�K��	�o��b�3'ZI���;	FA����-��g���=F��p���H�R�+B]���Ȋ0���LF��	ҶU67���G+��lڕ��u��2��M�)� �!߀4)���^=��}����/�=�j�vz]������Wȷ`�\��9��!�j��hٕů*՚��F�)l�Ks���%{iN���t�����o.~�� ���n�J����J��A�������	��2�]���v� /4�����}"�Z
���(�����jB��#v���o�Y!� �Ѣ�Nf˶ ]���B��ڼ/Z�0�集�8����-�vx���ϛ,��P��.��!�X��/<�Y�sVj�X[Lw�&���H0�A
�,���Y���4!�)�vm#$�	��^*�B� 1���&�6i>m5�����%< U;�l��[J�nVp����n�bi�RϚT�jy��6.W�m�iɕo�F+��ƯX���h�NgT5��=p��,p!���Ѭc��2�
d�#���hI�(�x?M�y��P��q`n5�� �
��_�=��lW�w=�ҫ�M0�n�C����>�`w{��1���È���k�͡#�|HcI���BYQQ��Mb�e�d4\�HG�pa�-V<)���p]�����]8�86gFY1���V 1�{���Y�1Kj��T�!��6T���b� }0Zh�KM?YL$��Q�
e	�.�u1fb�Q!q���߰Ե��"����mP�+�)��F����V��Y7L�O�ۘq��N=&6���+~����S�rlt�=�L��8��Q�B'����A��{�{�AO����Ǌ&Ě��=7�u�,Gͫ�6M ����cu7�_}�U��%�GA�碼��?��ɴ�-�����H1*=2����E��BOY�e"���� L��M�
(���^�	�ύBu��H0q�w�oIB�G�1�i�Q��E�b��yz���Q���؏��G�(_4	��Mk`M�Y��s�l�Ɵ+Cи��4!N�n�^4�V�7y�T�.&<�PF�F�oY�uՑƂq6<���#�"v�zC�ٌC�tV�	/��z�Pr۠u���?0A<Z��U�,h���@��z�F"Ä����2�<<�S��9����o��I\����u8@�&��k?kU�P.�C|2	��7�������5�j!��p�.M�z9���~��o�#j�<��M�Ҝ�Lz�&�B�y�Kܧ�vac��C��!��9��9$[2���bH+j��V���l��̉�x�/�|������i �p�6�����~�f���Q��dǎMN�t7���HT�(C���RP1.�=�`�ËHl��aL���|���~==X����97�L��1��X�ŗM�q�;��4!�#5�@�^�����ua�-W2�>Z]����'leI,+W'u`���}�,J�r�;';^tXae�ѭ8�%�#�Fs��I�I�J�y�0�a��"a�SS��\�$)���c�N|>6K�VO�u>?dD$��B����U�15���|ϩ��S�D�3W�+�����
a���d��!!�ף�5������cND5IP��JG�&���R��m�lJK�{��jk�uӴIY)��3u��7�'�)��("Q���/q����4���MҊ�qRbl=>=�[�c%��%��Q�٦M��X"�8��ͱ�_�
~ۘ��(���"H�5�.J��X�II���c^w.��4r��mxy����C*��	��"iW�{ޝ�Q�_^��&�:|�l�f�*w{��	ڴ8/��U����z[Tcy�G3�2DL��46�0���7�2anD�^RA�T�؍Z%�yuR��j�B��X�#(�J_�!*Q�f �����!�t�Is�}��Ϳ�2q�D������S<m1Ĳ��d�2�lv���j"T��svsD�	(3���<��X�w�,��u�+��Xۺe'�#S�&��n��JIµ����j���o�\��Qa����I�B*��ކ�K"W���̬d �RL1�!}�w ��XH�Dn�C�Z�W9��i�Ԥ,���Č	i�r��,hp�(@�8 .�t�p{��=/�vn��޸�*�5d��7\_�p��O��X���t��
~W�3[>h����t%�Z�2�PC�ж�Y4�_�2��wv舎b!�+e��M��g'О�[Ϗ��KD0	DE&��,��䧆2��I1d��U'2/��B��o�Y#���i�d�N��0u��F	,Mސ�ng7���r��Ŀ�x���<_w������O�ʑb��$r�5c����t=���$����;%�qb�A���f�
�sU�rr�I`�V�$<�D@1bb� |����q�����vk3��T}~R&�Ų�'�E�����9qֲ�{���w9���q[��E��߭��J9�5(9�V���\=XC	rI�2Yv��L�x�9�4�֧][�#u���i����d����߯�;y��N�9NB\ǳ'��1�������1c��7ڋ��μ3|���ڧj�4;��k+O�HS`���F�(��Q|��~������=�K'��IOyW0d!}���{�É�)�<�	k>�x�#��:�Tb�O}��;����<������#�HX8�ex!/��H�7H��:��agy?���r������_v��KI��j:4:(��l��+|N��fr�=N;j"Kx8Kf�� ���y(1���&j'��3�9�>��{� � W���'U�8f���_
�]�>��i���$����<Z���5-��0Z��ޢ��]~����c=
F����ʇ {����Tq4]$E��+��3�[S3<����2�Z�J�¡RV��[��w��3E�2#�mD�<��}6�S�X
��9�[8�z������Hh4`�����R'Ҝ~0��-�=�{v9�=d0=pP�t#�̵!��kka��o��&��Y����ӷ�3��eP��pL��LݧUS�5��Ճ�k�Bmz�8��ҳc,R��RT��P�B!E�����������1oa�s ��˭�1�[��y�NJMJ��Y�;y��[Z�[��$�v�Y��`5�'Lb O=��e��`7��@r𛭺��L�<-u'`��H/d͓��!�w4PLOg��U�R��Ur" ��5��K��54��eAeԇ}�5��)��FA���T_��{=��G��.�P&��Zŕ&�6,���[�5I)3�1�EpP��<�y,���o)�a&4�l+��`�Qp�$}�������������8}��M.K�fe<������(��0��$G|+@�}{%�N ���H1�%����!����f�S��mC�N���+��n���	��6�.:�ݴ��n��M_�("S��G6�ZP�9��?�*�٤3����N�K�l��8	-ɔ{��]4�X���A����:��L��(y�8'����
;[��z�%�0�[I���+/�T�Pe=�ID�&��`D�����3�!�4���'��2�i�A�u�;ވ�l��y7+����Yf��jl��>��c�M� �_��.���@ڜ���ܚ��67�<cw|�u�Ͱ�	�5Ǖ��L�0Q�e�����^��+��|�qw-Z����+��a��ޢ-�g���@Όc!��+LJm�kܺЪ�lV��z�{�Jc�xWp!~�?�u������dE�������n�s�R��6�:OZ���K���:���L`��^���D�>�b�br@��T#�']�r�����r�c���G��-mX���❅�t`T۩_�CX�F�F!�)��z���*���*��p�P�E�֏!I�:��;��c��En�4�bxUj>F��ୋd3=��Bx\!矒�"��I�.n�g�z?�T�/�l"�d�]l�r���9&�̂Z���X�`��9kg�M����{D�~Ǝ��u��!���}do*>��0)�W`1�W�x<�'�B��S+�@|�j?�MgfC�kKԖd�M��d�������t�K�Ba�̦��;qO��^.�f!}=�T�a�M���D�c�-�t+�wh� ����s�����\�;4C<l�
�w�2$m���,��W� %�c����\�
Le�~9Z�]����sذO�CI��T�v+�b儛���7nƵT�������x;�X��f~�e�o��~�.,M�g����C �i>p�n�Ѕg�4���eX]�d�,'����2����=uy�W�
��B3���N �Nf����X��i��c#��u����&Χ�l��%�3V�7J	Yi�cP\����1=4fG<�JMg����::��{�{8��S�,W�R4��^���� �����~uz9Q}���+�FG.'��\E-Ք�_����7'��BF�Z'?D��#�4���f��3���ڷ:�Xj���3�!��� :,	)����h,�x��-��1�'8^�]��P^�$+Q�.\���]Ћ��$��Tʩ���:�5&4��)ў�ڝQa*#� YX�
��K�6��H���H�Tb���Ԓ��5�Q/��u��3�A��ع,kP*�b��̾����ܩ�4��m)B¦�ϡY{zIE��Q�2iiu���K�z�8<d�E3z�I(9��<�HzP���
���w�s?S�rO#��U/{�Wy���E����W���wQz���ͬ\1��b�̸Ĭ�M�����ĸ%1�q��4�-f,,&��o�r���1�D���25��帘vPw\&�6��l}�u�%�u�Wf�@��FӅ���_��m�k�.����C$C)��j*Q�rʁ���c�cbaM�/c�.�LR׸�s%�눏;�6�VZ0�Y��i��pڨ#��.�e���E5#^!ɋ�$d[%�D��e�I�+0_gn�UX)�Iz\�Up*�sK,�_f�Z��2H=5L�d��[��	��Ȗ�
�a�O�q&)�B�^����Q���B�Y_�AF�ل��t�QK����Q&A��V���W�J{=�퉒���5�-�El֩����񉕙vv���(�����e������(��lnV�.W�E����;4�I� 2�����L�u���2]p��d��Y���z�3���ie=Vp ������hUG�L[_�J���S�t���}!��[�}�����l��l������r����:q�E�u[�៨�d3�>1�ʱG�=� ��p&�y�o�jE�I���G9������u�FN/�\�/p���5{�G��l�ˊU�y����)	:�q`m���/&�����X�������&+�΃;�	4�X� ����
�B�Y��˖x}U�S#I��
D�����'��TU@4qf���j��LB���~9Ҥ�P�%�=D7�������I�K��=ފ�����JW����w�>��.����Ƭ.�5�������ʬ	%a!L� 
����:u� ;H��a��1a$�Ϭ!�9�����zv�أ�k2m�r�F~	�
��V �`��`���;L�09սOMCL���y-D��1_��<�|F"���V�0]�[���;`~%����i��h�^�!u�P;RH��j]/܎nhi�hK��7;E�������C�7�,�e�i������D�]�g��d�p��3�rJV�s�ԏ۳��Ua�o!^0�����F)�[H��!��>��5��l���GR�����V��b�*��vT:�]��PR��.��)848/�fc1�.��E=m�T�Mb�-�� �#i�O��������,t��$����� �Ǯ�x��zW�/��䷒>B�F���d/�����z�B+�/��V�̈�_�s�y���cc����RU���xu��ܓ.w�8���㦾�Aݬ�F��]%��

4��i`��|����liS1��� ��}j�����V��̿�ܕ%LF.�O7F1a�����)�E�.��$+W���E���Yr_�вEIE�B83�R�`pdcڈ���]U��/�q�#��#��/d뭌p��q�׿ۗʡcYm-B�C��6��+*
������8	'�k�u1	����j#�Lq�dK;��;8L;ï�֗k�0IIJ1�o��A��<��� K`1/�����p��������Dn�%�A���Ub�5���}u�-�/&�������V�a
fI�_�t�R���Y���~p,�/E�����@bZETc��[�+c��i,=%�=��9URW�L�'���&v~/ӈ���iX_Iv�k����?�t	<��T��~+�	�6���t;�!E���zD��Jl������p揦S>R���m�O���[cL��
���E�=+�D�=L��ֲO������}�бE�.�� �)��K��9q��]cƢ���Bv1��uȏ��\i#�짾,@K�)���R��\�>�R�^�gxp"`�/��c�8h����
w�g�7O��P��p{�\%�/��h�i�pQ��O@6�	�Ï�{��SS%~�t���H#IJ��$@=�̈́��w9���ià~�̄C=K�O{b
�ܔ$��X�����R�/(^���=�+��d�8�6��^:[oPq�?��1��?�c�kT~E�0-��֌R��F��ݑ�}����ߒ�d���V��|;�����8?Z�Ŀ�o��
�l��&�^�7��f�a=+���d��ME���}�?@���T�K���S
����ֲkz�A�`����ٚQ�nF�J�䮕A�T�K0v�����.���|I��rP��\��Wg
���+�d�9�z��X�W�=��B���;�;O��d����ˏϰm��/G����<���U�")4/�1�w��A���M5�G��Ͱ8/R ���$j�J� /S񔥑��Y �����U����ѧ���s2�O��$��iI�ĿcM�@S(���*��Ϛ1���i�!zk�@�ޞ<�����k�kϼH%�1Q�\��S��W��BXZrL.
-�p4�ȭ���hFk��b+ӳI��ӅM�}4Y,��їKk\V��>A�u��0�ᇐ���d���; !YE���/�.k�nOA]��ނ=�<i ���1�j ����7���|�P~*�*�����z��Ō���&fۢ��]�r�s@�^A �Mj�z:�,Q.�a���T�̵C�xؒ�RX����W�΢��]���-H�������������:"�󟀘��Q~�Y<mU��2�Dk$�m���N�R�z��|��'y�S[��i2cy���2we��:�9:/���7��m�lw���̣��XKӏ�� z��&�l3�_Yˆ7���{Uw/��n��0G�*R��>�z�t�q�]pؙR�!�f��wbfZ�B�8T1yD��k��x.�sOVQs�KA��ɌG�|n����K�������B��]���,	�&~�Gx܀���hf��A���1R��͈ �]�F;�K�=�T��$�q'�d�e���	+��L�(�"}�:��cf>�Lv��Rx��%,uC�2�/�u�و�P��'IC �34��q���4��?�H�\��ģ��$I<{oB��>��|VXj`���0�w_=�Մ��yI1�c���fF�Y����/�O˵��;+&���o�}j�A��=��z���]�>�~4K-�M 0�r�VдSN���P�r�Q.�������c�d:��v1 �;�/�M"�ȕ�t�?���|������=�
'eX��b�ג�0_xT��}=�
��������9愕U
�P�/��}ff���51�C!<�U��b���i�;��Q������e/m���0�cQ�<^^!�nb��4%�I�T�/��>�|2\,Q�_��O9X����r/ǆ���Z�/� 2|�>�� ����39�8��a�^��Ș�Ր��f�B��CCʴw��1�;0�.G�$'���Ɔ���o0O-��z��/"�a���E�*��]��e*
��L$-{!��A�ie�����?;���]��^j�Ub���G��d��`��#L~�J�wj�Sq.ڡ�Y�OD-<F���5�p�6�s��>�/���/7̘=$�m���m�M�o_Aw��4�G����^Y�Fn�_���GH��g�*7��&�JQ��/C����# �H+�꒑t���*�m*�i�(��Pi���h��q��IŰЖIH��Z�}�0�By���z[sN���X�< 3�9*����ʤ=�����92఩��܌T:��r��+P��]���`�2
FC6}1[w_�A��#�;�%:_�ȏɴ;��� R9�ͱ�k��d~z~�&=��������c�4a�{�@�$��I���qc
��/A�@�9ݕ�C�X�2��Iv?ʥF��Ci���].�H���:[�¾���#���7V��P�H[�d��3"�o��h������jʊ���I�����{��T�����JK���O������pn��#
s�}���Î���l����4��E`x��-������N��ѿ�n�*(I,C>w�:ZT�������ʉQSX���)�x�êM;�_�6i�Y�D7�~�����28+�D��=k�2��U�nv���}:~���|h�H�i���5��g_ѵH�-Y����?XsT����v�a��o�\GŒ;���e|��9~a�F�ʛ��7��J�����?6D*MG���i�I�E�j���E��=��k U��{����㒧,F4C� ]%gj�JQ��nyKz�	��4�N&����S���)�g�{�j��!�:'�~\�U���m�"�1C���E�f����^V�^Y������bVh����^�'Y3����ϋd��.���-5b9�)�؏a�X�xO�p��俿PEHZ�pb0W�5�&'幾d4�/� ���Ę�PF3��7�.������*y�~�{�ކ�E���t��&
I|ү�pz��mf�"���A��q9�XzD���[J7}$t�.ިi��ْ�y��Y�2�v�-b��U��烐����Lռ���]��>�z�Y��jճ�ڧ|ȶ�?���t��Y�1Ӑe~�������px�Z��<I�`1��$f����B�0b���L�׾@}�# �֯��d�V���u�0�e����u �l2�y�\�M��e��i����&M��L������6r����E3N7r*<�VJ��#kI���j�P��Z�1�G.�O����_v��K���γ0�A��^��j��f��oi�B�v#�����2��0@D�I&Q�iW��96Ë1���j["C2ϩ��K\#�.��"�������|I(�%7�� �hƷ7��h���]�~XmH1��B��V(�}e�%r�����\���r�X�#Vn"�����A�Y�e�o��}��_�v�vs��#���PW���@��d���޴rʌ�'�lE"�	���S��ZM����|�?��xl
#s6c	��ȠT�N1�@�r|p�6�l�f^{i���I�8�T��&4C�S+���M�j(�3� �@֊�����Hq���W��S]����ݣ,L@\��	לb�[�:)��Ax�.ǹ�A����U������������f�&S�{�����K�����Q` �TL���`���@~������~�������,}S�U?'������?�> |T���Y
D�3g����������W�(9m��Sm��G'r��l� �<5�'�%���~��x`�F�m�Z�dJ�b��v�F�"_֯��#z��-��\҈g)'�w?}��3����I�����dy�Tm�I�]�3sĶX�v��$�;�w��V��Y0�w���T����Oa�k�>��È����$��ҹc������ի/v��vJԟ���t�1el���O�dZ'�n�@����ޭGh4ʦ�p1�����g}vL��7�΄a�u���~$IlQ�X獆C�}le�8�!\�6�p8��x���޿y��&uV�q���_�O��`y�x/�����WXy�k��y���ST589���n~-nC1�:(�HB��6{��j�_57l�{�Z�t�3�`��<�`��:�F�[ɡI~�T��S��H���!�����g�^��{"�"?J��?��B���\Ƃ	�	��Pob��9��`�G�A���p�C�w������d�5�Lf�.�[�pu��~p���zb�T؀Z��կ��Yw����hrj��kf73���ɚã>����֘JqN��n��@Q�H|�V���y �1r����^n
�hĔyӜMӬ�:�KrL����!މ�Q2��_>X,���e�Ёf��+ג�����o��1m2�]��hq�a����+�n���<�p�FdErwf���HA����&`���}@%KN;-������;��x�j����)�D�u�sך��3�sRR�"�Ul�Hv[0��%ֺ�6w�l�؁,'��>o-��#��1^�WH��%�q��sm\rk__Y�X��|�Κ9����Z��2�
6& �L��k�
��K�������C\s.����
{퇄�F�>� �J 2D"�U�'abB!-�A�8h�ТDB�{lN��7���;��L*�I�qRT׫1X�T����#}�j�<�q�6&���ќ��aB� FN�c�A�����#8��PUIɜ�Z �
��,Z�|��o��#�Z�R
hkH�����~FoW�Pe���Qj�������g�����D[�׻���o��b@n&Ц�cX�`�2Ig��\CB����{���p�)�?�Bw�٩��+��rz���n�8�YV7�)�������EC�@0���'}4��͢��TD'Y�f܇?�g.˳_Xr�����l4_�kIoS�|o鍎(�/��	PT-D�:t��x���'^��47��ʅ ����琠�@�ѵEj����89����ŵ���iۉ@��]]u�� �э%M�����J���ݿ��Fq��t%���iY����$��e�1^V����v�U���)"����Y��X8�Lx��/�T�U��@�Ek�nMv�$�-̺��1��=Y���U�FS!����V�*�랽
�h�ËU�Qk��vA"�o�����J��|BXаH��,�,?jU�����m�3~��R����v)M 2�U%'k������&\���$q���ү�Q��נ	ȰJ�遫T:Ea�,OE�"hӿ>'<q����qZ5�0�6f��D��t�|�9X���kU��6�_�`ݶԍ�(�� �N=��ɣ�U�$�)U��G+죮R�3����G�S���f�#B:�=��M�r�����o����h�>�6ocG�jOVo����͹B�/c$���b����8��DH΄E"��}aESf���]JM�E������:�s����S(	"2P�d
r2B/�:+��Q��]O�7��/�#��K��D���hwL�m�j�3
v��b�?x�l��y�J�(�Ψ��w��b�ӊ��/6�����\�ht�� &pJ$fر�����K��㲨�{�W� �?�!���噐$u�i�2���#�ҕ�r|Իh�^�/Ҍ�.U?��fHk�}���Fݩ ��@o�~��N�#���Ts���Gp�jm����Aob�v�B&ϻvQe��+��젤�,&�9���w����	���VE�"�~ӣBȮ9���s'��{p���7��Wي��[a����u��Ӷ4j`̲*����V��N�C�`t½%�%$��!>d`�<
%ц�*k��R��N������%~�>fgч��ב�Z3J���=f�2�/R�y~ai�C�x+)<��D^QT�����v� ����$x�e��g d $[�S�]�H%5�4����Km�8�ÎA<ĵ��ׅ�O�O^̾��Nh;����1�-�V=�H�I�mb�@�e<J�ꉄ�#��w!ca5AC�o��Jٵ\ie����H��UN����|D�
�
}�$�
_��w v/�d�����-D�T�ˡN�IjR&����m�L�H�n9��a�!@�[�bبz�k*.�h�6�ap���h��1���>j�~i��ˬ��%t��Z�IÑ(�[2����;�w#Ue6��sȟז4���I�{6ߴ��7��r��LW`��]Ph�^�bDgf78�n���f��]���:ZH�׆��yVAZ>y�k�oZ�B��\z~�*������Lx�>4�� u^��1�,2Mg�jVH#n"�!RJ�����XA�Ӳ�ߥ*�)��͛�C��"�CD����,՝W���p��ڐdh�&J���&�g&��Ù�ӣT�{PMp�����e��+7�
�edU�V��X������-�Ny��/5����v�>��?~s펺�>C����*^u-{�3g��y��[�
	A�����v�W�J�HI�x ���W�
�5��#f62�J��l%�k�FWB?h��-S�JD����0od+�����0�r�4��\Ht�8��|���:�G̃:A��}�n���[������c>%*o�i�8W���}�ei�%jv5},1,��=#��n�| ��'jx7�-��qJK�k.�r�7�lc�?���ٸO�K� Bj��?�����S�{ͫ���F��[����x��Lgѓ��9�)[3�Ie����,��:����xBS��4¨�p�к�8D�fԛ�r�����Q���5Ǣ5'H�봵+ӗ{�ò��2Q89E�m�������`
p�l�(�M�M��h���(@����;㦰It*�;U�U������j�tb��U����6��.(C��Ui�t��
������۫� 咛�I\s-gΛ�V�w831AhC[�@���&V�?��ڳ�"��nq&�4���4=к;��l�r KJ�dt��zw�<�N��?����R�Fd�5�ە׻e�D���r�"�-�X������+�n���ɧ���RjH|��3���D/�7�Y7��`���g*4+ �5W%^��������>M��Xz�����AQ�.+�|y|���i60�"lK_��y,O�K��u����5�uh����K��9�K�s��r$n���4Ӣ�ѩ��gpOv�%�~{�A���ON9k��F�~��M��m��
�މg��n*�)(��u}b/�u�[--a��w�ӣ���;#4:l�Lj�i��4���t�x�x��17Ux��,��m�A��o�TU*�9JH��9_�� m���B#M������ݫQl��{���?����cB��(E��Kƅ�6�;�;��t. ��zp#?�t�3w@���Z�C�}:�&��˰�D]	z��?3�'v���R�t��8�m�,Q��UI&�j7_���
�,��B�eqr�eo����c�6�v�0���y�J٦)����*���-�۫��v�H�Շ�̮	'��7��>�pk9?�݊b�y&ATO�9.�#(`g��<BS)�y�-}}mwϒa3�)QUyX��A6�F�rD d��{��-��N� �&�S5���JK���Ū������͊u6�G9Nm1��;��v��ؽ";�Ad��/#狄)�f�1£x��Ru����&/g/*|�)����a��5EN��_鍧ø�����_y��q%�ڔlA?�I��L�H|�N�M�ӯ&��~ 76Q���Yj��P��8��#�#�A�#�g_-�������|%�:�q�K�i3`�k�n�~c����X:�4�M%B�����K馞�����	���7�-A�mJ�h�Eٗ����tujϖ��(<^}0z���2ר�&�Т�Pe�|9u�"����n�p��.��q�@���Č��O��a)M+�ieS�3�����! i �>��S�o\��Ѯ����&}#�oݝ���ӪE�L�����]����ItGp�/丸F�����MH�����^BG|ui�b&���bǽo�~g� ���]�����}~kw���v��M�G�ϧ��A��f-����{�������rK�tv�U��,r�ݥ�H�I�������,�\X�$�!
4�A�|6�/4�ysǟ�j}&�w�2�eGj.������2��Y�hvE�T.�3�H���9�1t�t�ٰ��8���ω�>��GvO�2 ���9:A�}џy"%a_P��`�3a���|�2t��!�Hm8ڶ4��C�u��&���t�q�K�ӵ��A��>w`��l}3�����U�k�$7߷K�m���wXQA��:�5�U��Ǥ���gN%�\+7`��@�8Rj(T�<�?�1�����j�L?SOj�X�~�W|	��!Co�|^�K���p�#m�nF�E�s~q�� a���� ��H������䨤� ���L�n��B��,
��!Uh�܃c�M=�1�BHZ��P�M�3nӧ�5PzT
� jx*tW�R����{�g��s��F��k�������ڄ�Ћ��^�U��������!�rE�ra>�U�����l� �U�E�C�S�r;E��:x�j��8A�!��o�3<�9�A�wǷmp�0t������ό�=��X�o�3a��[�E���E�����B��%L��=�R�}�f��D߻�eR�z��ɋ�A�P��ݧ�.�[�cʷ��(hLI��Ȭ�w�=�ii��i��)� 7g8 5����h�v�/��3z�E�e<���L��HO}G �S�hL��X/9�֛�� �&�X���-~vr����ɪ�M��W��A[~�F� �Z Ԯ
������g(���F�Zvk�W��S����m�	�$�C��u��?۸]���
S%�BX��Q��%uR�M2���m����Y��K��_󑼘�B���H������əA��g��E#v���%���.���>�¬�����AlI��B&3D�ۺ�yJc������uX���Em�s�Sx���yY�_�@"ae�]��vY������y�����C{��VQ�d�̚e�m�̪��;����e�����m΁�q0�|2f ��-%�߲��gI�:�pV*�����2r��P��M�xQ�T���B��w�]�en'��֜!t4Ϩ���hW-�G���I�	̻n�K�)�2d�S�H^υ!�c�@�6��)��.�W�V"��c>��>K���+*軙�L �8�:��b\o$����na�
�si������`�9/�c	" k�}J�ڤ D����Z���x����)X�E	�u�[�Yo|>,�)Kښv���%,q.�Fj�W.ȍi��~q��� 
l|�f&�,Q��E{]�&�7���q&^7�X!���
�TF�2��y�v�������W�yD� �,�St�Ho��p~po���",���|⶙���WΕ�x-�����ەq�%�4B��5�D�	�A�w�Qp�uF쨀�$����_?M���<�(&"�s��;3P��C\K�]/)џ��j-q&�{���v_T"%ʃ�CWM� HE��%�
޹_:��H��T��$�& ���e�j=�T��>��Xz�`5�cIy �����1��" ��@DoǨF�$���0�{�<o����uL�Tc��[ub����U64Zg�ys���vxwl�F��0i12EE����a�s`<RR6��/y�7��X�+R�9~�d���v�3�e�X�{� �4L21�ޑ�Aڄk��E�g�Z�c(����h�s�h�X_�,M�?����BP�u�Rz��֜�d�$���C�S�<�k�Y'/��d�o�k�G�%2{�@#aٷ�E��t��ib�#�kR��D��PW_x
Ԟّ��O��B�lа[9��F#��dU6��s���~~�W��-��ߥN9�s4� ��G_�C��'�6����
 G񛺜Ms�9��J8PJ$'%!�oHB�10^�ۙ϶�i�I�\����Gz[�����~m[.BS�BHU#�U`����p�]�S�p=Q��X��L�i��C0o�tv^�9�����Y�Ԙ�kr�5D���{ϛ�v0�:z�e �s���N�k=����s+����+� 7!�!z�c0�<1�=ф�Y���8���p� [�g5%e\2=Ϯ7<�V#�=ճAHP�ld����cp��H��t�'���u�l���n2;1mP��{E�Ҙ�!�:�.P8��@o�7�CIN���J�-��;ϒ찮P�BS��#M5Źs�7����2�FX�#'E�떆!�1���#��i�WY�љ�8\��s�����MAY�ɚ*Z�g�-H�tp��D��e����)X ��]_�&���r�SR��A�����=n�-��]�<PKj$ ���J�j%U���/]\�R!:#U�e͊�!��%�����,�A�o�{0Ic����Ρ�m��
_�#�F8�ݳE�'�sՐU(�J�Dub�^��k��Z:�(�n���I����V����Y+h���s��f97����d��п���pǫ�t�qkm��m�^�d�Ͻ��w-��/w��CR�jkfu)��DΏo�/�x�694Q>�ȼ�����;���C<莜#{è�~$f�蒾������^Ȋ��)8�v���1��b� �RF�!��}�s<�|���]M������5���C���b��ₖx��ko%X ���d�xGG"��	��z�7l�Mb�����Je۫~(�9IM$I^��O��;��ZH��GG��{����o���%�6xp�'��l��n��^F�]���PE���U�c���c��Nk�~`��tD@aS(E�0n;�΄�'��?B	�!�	qB����*�$&NW<	5��]j�
� ��[����ȓ(�(C]���4f>;j��Ke��^�$�87-<�"�oշ"�z]�9���q���7�=���(4߼����3\��X��<�^Z��	��zi@��}�!u�:IZ��>�_;n�sХ��a0']_\4��7�mb�с�a�҉�.x$��d�t(/��h�I��o���Y�{.�Y-��D���O���] Hk�>3��L�܋��Q=*�%t�,��C�"���1L�~�������|�J34��3����J�N�5����ટ�ܷe�u��ߵ��g�,Y��tW��otPu���wu�>���)�T4����xiZ�h�A<u�$�U��e��^9X9ѯg�~*�w;g<�/����R���yW��}��_7�y�ku����-��ef��󒗟}Ԇ�Q�*7����G�����@Q�>ߔ:_�ր>h������K0�s-x�QrkZ�_*�� ?C}�a5 .�3�-eD����8K}>��}ܩ�٣�R�S������R�{ �.`*�z��"r5�g�Ӣ���x�w~G׬�i��ԡ���g�uhM0�"E?i_����r���&���T�F��%�1N=�I� V���!vrO���f�q���Y����L�O��n��QI�,Gh��ŦW�%�HpA2s�?�=����N�OI[��i$W�O������O��j]��< ϊ���r=}[-���X-G;G��;�z����s��|���3yN�K��{�%�H�4������4~,I�2��Jl�A���f��]�&(8pT�x�� ���V����t/<X�o,1� ��XF7��/JZ;����v.�H����F�L+���� A[���(0uo1_���oM������Z�_I�Mh�1%�߲�4m�E��V�P��]��x-���̯���$�8��;E�%#(Z<��uۨ����u�������j,V䛞Q�� �A���޻?8��Q!j9(Q�{^�����"� �з����]7Z�gI��a��P�~?��5��`�k ���q۱�%�������zB�@ܑ�s����ZXw���P��oP���}rp>�
���ͥ#+�D���޽�w��κ�!�8|	��r�l����=���¿U��J��HL
̅�B�oF�=v~���_� ���k���E�0�1o��E�:����5����QWɉ;��)��4 ҆Y��H�$@lpM�j�����IW���-�TMh�/�Q{�Qh���ԵT��_^vϱc�4I�&4�n����d������2�9�+B��i�6���xii�{���Vu���w����ɭPk�� �\O��pv�w�C�r]_�NN��uagTH�.� /��,M(
�U�cCv1IT��-�&�b������$�`�k���ђH��/lb�QK��$������xd�O�������yPYF�7�/��@�����T�ew1�'��$�շ����+T���`#:�}����zu���w'�E�����։ty��|B�$2�JO�w��n\RJ���7���.�4�t��'�	7�$��4��P_���$�m��R$3�itɱ�.�^ow�SkdE+�֭�²�)�ut�x�����@� �m�m��+>X|��P�w��8s���8��tx����?܉vL�t��ʶ������.ڼr�|�
{F�o�����N��@�bÑ��%����8�1Έj��$Q��L�=�s\�&��G(�^f�m��9@���E
�u�>L�=����;ڄ�fJuD��D�r�h���δV7w��3ԎY���$�_�<
hZr�!<w�v����s�ũ�q�b��uT3�hp7�q��Ĵ��������f��m_���:冨w	��}6;�]�
�kۥ0�0k7�˱��Nu����I�� �RQ�� �(0{jWZA~>8�Ws����2�T�XED�S�p
�X�d[r�;�)'ۊ�ǻz,9��at�mKo�@�_M��Q쫥�2��8\��1��)u�yj����R��;�!�j�s�!�y	V���؀�����v�U���tƤm���N��ږ���"���=��}��*�nt�!Ry�~{���i���+8%��������\j���F�����hwWE#4���Qź����'��s�N`���;V�G��2OQ�.p��BwGpK9-��_�r�Kh0�����}c�@=*���$��\\Pe��Ү��3+���A���Ҿs3���h�4R�u���`-��+��|6�g6�c>vJѮ��Z2�z�V�@ř!��b^��2�}萅�"���P9<�2٪բb$P�ֳ�'VVI*JE��D��?�&��������u�,s���lգm�/�&	�ݩnyFi�4}�ZI���e�Q�7����F���kۮ%���}�3�3�M$�tY5nިTF��NS(��[�u]��Y�>0rE�N��-c�3� y���J����1g|�ij��)�C=�Y,j���W�T�S����cb��L�~����+����`�y#cEخ�g���>T8l<A��|���!�v��	Ͻ���Y_�e]�_PI�3hB����t�4��}����O'e��E�|�m~�����9���}��({;��'��Ɩ�D�!̳� �4�j;�O�A����Prڦh���Z�c�t��K@2���l�%<�ڹ)|�'v!�'�E���N\�:R�t %-?���u)�1Y�D�`t~._����q#���7�JHE�
&:�7�>�����fk��cO�Յ<6ydC�����	�us&ʰ�ۃ��a��F�3��vƵ�M(�3�oƭ�|���6.O��҃�d��܆uWf�5�.Tk�^��T�-�c�q�;����4�'��%�v����7z��g����?�q�X�� f7eU��s�LP`���S�@�UY�������g90�|�i�I����qR���g[�\��G�.�,��7��p٘I��?VR��`�6,F���Ԯ�����xK[����n�ff�A�
���3�0؏�ǀݜzڅ��'N(E���ܡ���/`�!�9)uo�t1� �5��.�*i��&n��͋adڹ&iA� X|H�D~����iO]�����̈��p[���b�VIw3��M�מ���˃H�	BcR]1���} �zw�ѕD,�Ia�� q�)_~0"�|�Db�(�(2U!cu���3bՀm2�U2��_���\Æ�?����A;����mD?��a͏��k{e&
.��4u��%�]i��/�5g|�2f�&NC��xcG�F��*���/|x��j�Z�͓2d�
� �}��
:�I�XW��qŹ�xo8=Q�~/˴�G&B��}�w!GV�XHu �O~�6.}��i�m��$�f���]IL��'�΀�6E
ߴ��?6%y��m�e�!�;�/�i�~�� k��AhQ���^*���Z�,���4�Т��5���aG�Q~��w��ڌ��E
iVN@���.�B뙵��e��u%��W/
��716�I�z����S(b���u=U��9�c��C�G�x|(2�6D`m?[�F�H����?���p)�����J��F��7:�O@WY��U��+�N�����}6�kJm�l���+c�uJcux���+5^Θ��}���Ri���v��J��iY�f�6jČ$$���fbv�7}�>�������U�'k �)3��7�]f�{����TN�!�ߗ4|	��������z��f��E5��4T��Yt�Z�V�>"��|̈́�f�'gW���>�B����Z����0��u�U�������zxC_���ygB��.�J���N�꜎5�X�ј�n=b��,h
��Q�*�t��gK$��5�5�	)��K�$ ��<U�-਻I�·X��y\�Hp Yy_�n�tPL����fu-�i�iۯ�TGt-�3�Z�#}WА�K�M��Lzӝ'!����/'['���\�1��F�}�G�{%�ea�zHt����H(la�48-X��zۺ��� #�r��N��2���|M�Z��o�� �,���B�rxd��]�B����1���-X\������>'����i�ý�	��°@5��o�V���2?3�Gk����3���t�/��Vx��1B�W"x����A�Q�1�Tr�ߝ����ݭ�'r�?z%�V=���ꨴ�P5:#mҹ��L!�<�n�&VjI�9���!$�e�"��.p��K��_?_�Ғͼ٩t,�c�v��Ϲ���l��\���,��mEPK.sO�[\�M��=��Gq���_!�B��^������>ֽ}�^e�.�S"@�n��)�c�hu�~�e�)?k�׆���C���t�P�~�n�Į"�~�p��'�LD�Q0e��: P@n'Ƴ*��<�u�΄_��w�{�<�����O�lR��#�U�e�f������{n�fOޑ��F'W,�<��<Z��G���I��������T\ٲ�7`.l�V�+r	��F\��������3D/X�!�-�ߔ<u4��_e��I�u�bZK�J"R^Z��t�I�P�g�?n����ӓ��"�e�����������z��>�H��)��󆒞*��t�rA�J�m�
s��<@��<wTu���c�+��	.\�o����d��(�| ��2 %|��T��x�3��Kgt^���F�石|HmpP\�!\-S5�լ������s�n��~��Z$��9?W\R���0�(�^oL�(�.�,ĝµ��L	1�~�A.���OhK��Q��>nO�d:v��l���;D��9[6^�êH�C��	$����{�tdɿ�G�5諎�q���.^"�jQ]���LFY���YN!�{)�Y��a�`ަc��I[P����ޒN� �����0A�\Y"�վ~��!}C��}�+?��?%���dE�)0<��zЉ�z�/n�����y����YA��o�}��b�"uҖ۷�e�jOM%r�R�W�Ð�\C�o���H罶5���$j;$}����n�(�n�S�jq��:$������s2�m�K;��yZ��َ|D����D�E7�t��^�n�t��r\D���	*L��baBI�}��s�g.���o��q�yBټ� ������,�zF�D����ծLH�Z�֕,"����S^�ù��,w��r��T�*y>��e8�_�
�G�G�<2=
�ћ��o�PUP�c^q�YV"�X��y{�r�\x�l����JdE �yp`+����˻#�u�
'&��Ȱ�c��!���i��tk�&X���� "��J��:v3����0{`]ݳ�IO��ޭ�W_��i��1����Z����k��B�ifį���J��a�t6t����|���&���q�{e͙$j��m��X3Jg�֟s��Q��]bէ�Õ4�Eߖ�)���ݐ��&�w�>�nl����N2Y4^�#����J����Dپi�,8��W��2XT�5F=a-#tsw��[]�.���4��T��*uT��9X�y�H��vL�����1�-:�s��V�N�a��X���\�
9� ��4ޏ�+E�:I����=�Dl14�2<ap�a�O�$?��j��'k�/���l�B�����#.7j���$���%�_N�ӖN�e�����K�uO�Y�J�^�?x�Ɇa�J�w?q�T�n���K�d�jѧ��;MT89�$��6�A���
�O�P��C����'!)�Ciz��e*���J�t��H�.���M��뗏��\=��&���P�͝��&�RM>%J�H�Xe���;������E��22����-T@E��G�ٱ�@��O�T�[~E�1�p�|�H��J��O��7/w�N'���T�1���%|&���0�O�ݒu��g�d
�_�~&��Z��S�V~�
��r�H`����
��˯�F/ٷtN��EH|CS�1���Q��WT�p��};N��MN���R��PXm�=��C~�(�0|W N�(�aIǃk������7D�����킅uc��zu\��������747'��7�ǲ.����ű�5_b�+a�Q.N��tl��@ ���X��<LS��E�����H��>�{�@,���;Q� w���Z�gi�ON�l��SM)����h\�D��BP�q���C��	A�\��X�h����K;����[�#Kب�RJ��~��pH��<�h�#D�aE��e�<d�N�AP����v*Sl�8��z�7*���������u=>s7��5b��N���Bī�1N��d�$�&әa����z%O�ځ��X�G��5�5��b�b��q-�bث�4$��F!8�L��	x?�m5n�bb�O��oCl%�Zx�mD<���I�q{+}�K�U�h��b�s��i���$I՟4|�/�r�u���A��o S�����BqA�p�;��Ky���^}�[�;��qQ���N��(�,�Z��%Pg	x_dX
3�#3^DP/Bf��\��><}�~��&����8T
F2����5t����d1��X�T���l�2��(���3R'ؾ3��M�U�Υ$,�� �;��U�V~1N}��)��L*|&�������	6߿� ���p�=fS��n��tp�=V���~�NK=d�]���E�Z��i�3����)�K�3�[
y�v �o(g���f��a�l�'`���^�|l[<*��=}�B`3�x�G�����{�>Q,K�c�q��:Je��x��L����_q�?�@�����qSQ�O@��f�*��ˤ��2�^{9�v�b=��5�@�l놩3��8��G�4� 9���>3��m���۫n�P�nwW�oQ  ��M�������������],d���z����Q�ᬣx�+'`��w`RI¬�y����,�ω7��q� Q_�H���l������o�^f��"�� �*�J��
�p:�3��%�+�T�ҍ1�9XJ�WX����l��<�dE�j-\]��5�{g	ە�b����� �]�wR��p]�]���*1	
�)���\���Y%�[%#]����Jr�5��߶sm�O����.�'�G�gIͨ�ga�s��?ѭ~Y��*���|�����m��.צ�����(`zmy�J�Է�x��d�2�~��C�"�|�u^��t�Z!�+����Y�%�ђp��L����2X���5�͑��Ҷ@��O��6�8��UΧ��[y
#�1���Z�+܍�?(6�{���4��<G�H�Bl|\?������i!.�Z�&Pl R�@�<0�qK�7��ڽ<�P�2Ӣ1UrF�9N��m9ѕ��}-L��0S9�)��6���v1�f�M��֎�ϙ� �y���r	��l�F5..�ς`�Z8�w7E	 $�
%S�Y(�e	/S�3�=��~�?^�Junk�T�
N��r�3���)�ǭ�N��]Uh��R͸Jo	(+���ȥ�и$�"��ȶ�ps3,�4u����N�d���p�� �k���G�F!�������~����2�5[��3&������1���AL�9�˘ �k��� ����*8V�������;Ouk^�������Y�g^��I�Ƕ�0)�O��Y
*�ڿ&�-hƮ'[�;����u���Q�$ ���F�6�͖v���wIi���Ͱh;+�����r�,|�X1Y&c�^x�&�� �&�	�?�'��g���數â�;�����z��E��g����@F�s�ʔG��}R��9�	خKk����҆5��jؓ��RwͽKg���9���� �?b���m�j��G�� 9�q�h�o�#6��o�)��MF/&�o�%Ia�r���:!F	�44�^vys�^��D$���2��%'�$�O3��!��Cu͓��{!�
Xj������8c�i2�5}�&$��G?���d�*f���o�7�V��k��<�$����z�4����4���������%_ρ%��.kN�sYCpi�T4����k�Mk-�$�C�M�*��#7��?O�q�PV3�~�I�]�n��(f�p����]oa�)��ku�Ԥ�#Ҩ�\$�Z�����9v~�('^2����u,{���я��G�e��D����8x%(X�pt�2`cL�o�dpin��G2�d@�.�b1�3��E6��f�va�vj���J k>c�Y,(gB��/������p6�YZL���k�]tY4�xQa�������>�c�`�C��&m��T�0�0'������3������^X
�8I��2*C�\yy]��Q�v�P����ҭ+���,6c�e{SLl �<���m��]�b&%P��5}��Y��y�s
���Q�~pc��f�n�3�EWz���r:�̆�<��U�L���=:��K�~Ӏ\��M*��ln��yf��$N�3��f��bn��|.�pt�����W�t�·!�B�Z�B���vU���y���Bu��Si5.5>b��+����@�{�w�F��Ee�2��&��\��$�p`�NTp5�?�513fH/�5Kv�8Tt�6$��B�j
���am��H�7w9ȴ/���*�I����Q"���I�E+M�ح��Dw܁�������i��| -f�Gb,:ɕ[�V��d�ˍ��_�ġ�5C���o�a�[�&3����?\��3�V���{+ޥ"��=�&��mM�f*��댖��>�@�U?��Y����v����_w��K���w���2��go٦�S��A�' 0�<�<m�b6�Q��ZJ���R�|n!l�Kw����q�ԟ�k���h��)��ҔIt�݌i�'�>,nª{�2Q.���;�I9��13;W��@Z��|�����!�$�V����'�z-��3���m�3�Fo�^io�-��	_�m@�E*�?dJ���9����d�NY��Zt`fwѻ�y�0(�}R�D5�J��$[�)����E�����Q����P�<>�2�g0�kR��]vOwC(-s��Zǡ}���C� zc,ff�
Daj��5��R^WT��^x*��lc'c�w�[�H��y�,�]'.��;��q�璡3�Ϣ��7^O������� �jՃ4�
N`w{�����p׷�e�;M�����j��Q1��w���}�< ]r��(���e͑
AI{�eSR��Ʀ��0&m\���J���g�v��*�j?��K�-9c�#����q--�Hfkv�����#�NAyp����]�C��#��S����k�,Z��}4��<����l �.!;-�^8,�
�6��Vw��y���u�QYI��J�?3��K����;>�:��Z�H�M��ڠʙ<Ss�����S�"@v��[b�:g~z���d(PB�/��m�����T��r�`O���d����Y>K �l��s�YAϣ�Na�;�#`\��O� o�:��QR�P�$
�u���|���>i_��1�g�hNHT^!9��gF����9n�ޡ�����@�n��%�O/X��}�����İ�ɞ�d�M%֠����ݗ���j�
�jS�VS�.��v�ae��Wz�9�� �oD<��(b{��.Q�~�k'��Zd2�=�!���?����2�_�q�Z4RN�Uȟ��0��l����b���eGrmgE�Qt=�!ꆊF��#��=����R���&�h��͙O�Wm{�,R؄�P�e9��� ���P���R�!���U.G@������[=\i؋'��r�	6S����/�䜨:�ԿgVq/,���yؖ���U�Cֽ>\#I��]��y{���ZQ2ݺH^v��(�> S�}�^=���5A�8�Ȋ�%'e7-�P%%���w�(4zv�n�AI��#աf�&��?�����1�Q�o��ҫ����J����ɧ�|ʛ`�/&'�w�0��B�m`�	q�rm���	� 7�	9�-C��x�S��P���l.�g�b8����ǃLb�Ѫ<����(EO�S�۷�Mdr�[)Ol#�-��c�n�;ェ��n��Oj:��d�J�=�Dc��+�-��"�ft�y���Ls�xJ����눬ŧ�u�{	�����x���_��T(��_N�v�c�,lj�.��{7�a�ͼ�$=���4D3w��W�0@ܠ,��J4�7�8��_9�+C��5�u���)��$� �_A�+Xd%E^�B��k�~�]�Gh�4��bO�|n�z��R�G��"�AuY����y"K�
7�Ǵ��2"U���z���p��$ɒ�܋�/V"�&(���2��D�5��T���:W���Z�����C+�>���r�Ϯ��7{˷��� i��NY/f	H�!\p�VMn�F5��H0J����(�QV�G�LM����90��{W��v墴r�b��\5ˠe{�c���U��Ӱ� �{���7�B��%L%�G�&x[/��uB�<l��T�����}��2p��B9ۖ��P�]�f^a̅���0���_eA	7��eD��{��$e�$��D���+�tg�QƳ�$Jnc��)�n�����+l�3�&\�	$�,i��{�z���Rgac�]#�ZRP7�O�/���0��R���wA/e���o�:<���*�>ʙ+" SyyV��H�%�5;�7�6H��L��H㠳���[�����w���V�^ �#�0-���I�x���� U����vY�[�x�95�J�qGs�N���x_p�cP䤫K�o�,�#�(l=KI��J~q���z�/��p�~�.�`�2ܘҜ7x��׽uM�mֆy<����h��${�,+"�U55a"��͂����㩌�
;o����l�g��B�|�S�Q{�Y6�O�p���32Q��^�2��& 3���X�8���(�e�M�!�~��KF�)�a�K�����ԁ�GwQV�ƾ��b�|6S�!�f�QI�}����/�b����W(`Q�rl�VQXBL]��F�z0���ݚ����[��+(J���+ К����Lph�)�`��������E�T7Ⱦ�B��:��Q��
Ō�{�ST	��f��/�R��a[4}�Xǘ8�-�>��,n�4rU	ʍ�1j�]�Z؆X�L�cЦ�y�c]�//S��qĒ�>24G���ت29�hX�y�x�I��/�2�$ï]�f|�����y�k�g'��Κ��!�����fG��JIh�1 �X��S�~���]G0��a���
hO�U����B|.���Q�������^�Y�8�����o�]
\wXQ��E�&z���;U�C���믋'M՟�#�����c=��[��9�{ ߓ��I�e��dH��o���X�̌0��U��Ca�M-��|QGl�MJ�Ӏ:�x�v$�'�G���^|�8\mE�T�'�w�0e/�<�S�q[ӷ"�S&�OG�p�:���íF�c�qӦ�yL��C��e�O)��c|Kl�Sl'@rFxs�!���[6g��[~���~Y�}Ao<��?�h�Gq}�����}