��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$Rx�y�<��wA�*;�x���@�̦�W�X�fa�M-$u����n~�%���P�$��W��kYَ���P7�?UMfT��q�6�U��k�>����~�\N�(�����X�e���/6U|)�X2pF�]$h���d.���9E��WG��L�X"]�Ad����ľS���8od����e�GT?y	7�������ݵ�^��R�q^]�鍦�����s�ae���h��L��P_���ާ��YЭF���'\��68�b�[����w8�[X��V�F�0͘3����q諵�uW� �h�u\V�?@��_6G�_�*�G���B�絉�f������[�G��U&�����~�F��AׯK1�`c��[<��FY���4I� �#�G��x[X�=�Q1��`��R>(�w����R�O�?����7�,(�H\�#h(W�EH=�������yq��Ѿ��aF����:�U~m<|��.��0=�P/���4ǆ���T(����=��6���t�����n�|lߚ#`�a㝻�h����W���#'�R��2�l-����ìh^_�H��0Ԕ$�;LTaF°릘�+"��Qt���Kٜ4�v������,�=YJ �
�n�gT��^'�B"�����yr�Zo�@8���P�1`	w��m^'��Wp�4W�h�R�'�"�b�SW.�P���jDB�8�� S��ŵ+��=qh7�!,���>_��aj%>���YmK����U�]|�0w��9?6��S!��ל�������U�*��$p2���'���E��%W�_����
ً8�|�Z�~��ۀ��l���"����X�,-�՘��[�#
��r�B�P(f����N�i�������+c�A@�����/y�B�^��
�����"��Q��\�ԑ��ݟ^���(���?��茮h+��sYA�;K �
z9��&��8ϐ�7K���x�����L{ �T�.=�7�-�T��$��C�<��L"��_4�ۇ�:���!��\��%c��+������t�#F1B��v&4�/ X��h����O����<&)���+���9�ޯ��I(
\D���a���q�m��m&x>�2��+��(}��P*6�	O��'���q+)�t�:)��H�.W�ս�i� �V��ۄ@�pl����ݥ��BU����V�C#<Ɇ�����l�1���&�/��'p��e�1f���G��<�Q�k�q��*U��u���������傼���;�Y�I��@w���88I�GG���kV��Z���<�+e��u����oo��~Y�'�UpE�(�=h��"�̼Lt���i.�E./Y|�U�����U|~����o ߤ��6Vy{։>�<���R�����Pݐ��[���ߑ9�@%���rbJ�4���1lQ�����Z��) �YFI1����d��7Q2r���n]k����܉���V�&��&���6^
Ԃl���w�=��Y,ȩi�׊��Z����i.�k�9�OO����$_����rܦZj���<�c^���a�бt�{��K���>�oK��w�&r7�G�-�Q��5^z�K�%0*�c��������CXt��D�|���9:�ћZ�1�`?;��}���1�v�?���ol0��]�zi���0��je T�J��	��U �o�/7E�1� �+w�S��b�X�H�@ƪ߂��ظJ��m\N$�����'�^Y2����2bO 隞��!��mOOӶ#��6!ٖOK	�E���պl��VM�v����/�x����s��eZrxD0i2�s��G�:�[<7�9fE�9>�ڹ�� �Lױ�y�\<��?��I7#���7t�O�-l|��u�0<qBn�X�t*|¶Akg2����`�m�v��+��\��&�^��k|�y�G<X9'���Ct�����6dJ�K"��YZ�@8y�[����g�UJ�hJ�!�~�3�0hS�M`Xp��������u�k`j�+�W��q�O�$R;\�g<�~i�4)1���"H�Mx(�P�xtM����Bmx�钎5��v��f��-�PP/|��pT(	�O
�Kcy�>3f{0��5JC�ʃ��+���0(CY�k����O�>�"��$��Skʚ�I�/�S����&T�c:#ⲗ���jWf��b�Nu�*�����)�2UG��bEq���"���_(�Ύf^y͵�gL�0�7v��
�2٤0��l�#G<��#$F*��-I�H�uW`g�[�Q|��QΑ�q+]����f�?��q�����NI�4Q�{�G�k���u��<�n�z����Ά��D�>���&	��*���c����������>��
�ׂ#Y]f	����rݗI�� bW7�_�-Ζ����LQx�'�J7��)�;�r"2~T|��Q.2T#���e���;�\����5���HW��KBI��V��҈���F��F�*�؋�/�ńK���M駛Z�b{�����"����Z�%�r�u��橇���-��Xv�y`��������`�Tl��X>��.���	e���*���=���+�る2(��6�A�Q��^{�;
M����	��&s���9��r{gȰ���<�b�����!��=��ft�M0���A�E�{ͳ.iV��a���R���Y�nEǠ���'�O0�`����2q�d��hE=s���Տ('�N-2"�A�wc��a��tQ�=��g���yi�e��R4���D;������^�&V?w���I�C�9���
O���O�,j�x�DQ3F���d)f�`���L�����K���m�Q�d��:��	*�g��l�h�=z�R�uhN�p##�����!�FY`��̥�F6 [9�{<\�i.��QբO���
�\�:D]�S2t ����#Y�0K�l>"֧�U,i�$�&bȰZtn�\'�t�k'��F�~��4�@�&��J+Vᥔ%k�s�^��
��A�*���D��(�;��0v`��U��s����)����q�'݆Ȅ"3��J��؎eG'^��eG�7�%��d&��ˁ�`�����c]��i��#��E1���f��n��Lͱ�d�8�2n�-��LO�j2�p7�;By�`�M��C�U��v3��J���٤�;eBc�M|��L��4NP�a�y�� d!�FV؄m���c������$���F5�~��u6l�N��1�.�Ȁc��A���{���q�?��RF۫���5��4��6���0Mg�@0��#��f���g����u�$W��ʢ��~6�;�-	/��S-i��ރ��m�xn�M��X��P0T4��B2��X�C$MO+���Mo�����,�,��xI�ǻ�jW@9�v���ѹ�����𿥏�3FJ�o��Z���̛�ǫo���T
�tX��9�d������`��J*|˽/���he��è��
�ה�_�A�o��;�_�qjFѯڕ�V&�t�)�P�_����)�o!2]0�b����ג�M3}�p*KV�:}K�͜c�Kik��Ga��6N}�;�2�pP#%�-2�g�R�?��-O�<"�1��p֨%�L�����lr�nj.�N�g!���$�}Suw2T�4�"�&�����1��I�m��#���F�O���q��i/5HNj0�����b�v@m��n�J��}�c�aJ	��-9�cw��,�S�$�	u���H����&��V�����d�z�r�cOB�[#��D�=���-���?A���ņ�2,�PFh��n������L^��8�q�φ*R�$����I4^u�����ǸF�z�$S2���g�U�\P7��F�<�;�W[�6w%=3�֬�)<6ԫd��P�����-T���'85k�L�Z�G3]Z��_J�yL���'���)k���2���j�ʑ�K��~��y4H�.�*o{(nV�Da����)�85DB�#�D��I��|s)�·��U�4�:�bax���A�N����h48����!���p1�$����n��)@��Uy���FC򠵫W��梙qDV�PX���r���u6�d�����o�����r8�i���/��y̒�#c䞵p�l�C�kF�����!�b��_t!��Y�)�~�~N���,r}�K���Ҧ;AZ�}:�
9SoR��y���Yŋ��L���qq�Ó1hԞϚ,c:����<� %��_�L1=�� ���&v�u#H;��O��e������ŕ]�E#)�͓g�eK)��Ë+۞!��kI��cX2�?�go�4x�l���ʜ��7�6N>M�̽��^e&.q��FL�����j����OϪJZA.���e�Zө ��J�I�hAQ���]=~j�?̪�c͠��灓[�$?����RqV�}'���7D���&Y��X���O�=�����hI��h�{��z!�ө�$�
v%@vj��4j-[�@�h .�H��o��ԡ�����ZC-�]��aj���d�N�����/;��	����N��	UJ�c85�"��P;�g���ѫS�V]�s��4��f���h�t����\\g5�m��� |�)�dz�uV�1=��K�Q�=~	c�L����-�h��9	X���j����$eoZyVS��,&�u۫������#�IJ��)�����j8LmH�z�Wt��F�	t��ݸ<6ӊ���NR�믛��V�������]���"=Պ�1!~/v��ڲq4���o�?��b�_D��b�����;I4�. 5T�����
�a{
���^�R���Fvg2��OA_qt��,���}kK��u�)J�f;2����&J�見��L��U�R�w���4����=� {P���
�xj|��^��88#��{�mw��m�:j*oƮ[��].DԻ$󀿱���؅8�^;�.oQQ%:J�Y��o��5b��`����	hGIԻ��Z��~<�Y�У���el\3?t�4B����)�f��2F��6�m�#��!"]���(�8�p2+��%�l;�$�Յ�u]��_����3���twW���A��)2��Ш�%���y�R�/$�7�ԏ����r[��'x��v]
���˼��>�C<�^�oEL��n/��>X��J�S���L�b�Xъο~�[]!L���]<ݶ�{�_S���\����C���6��!�B|�c(�J5+�o:���0D#<NP��/x��}^S�թ��P�����(��6=[i,��E�ى���Q٦˻ɏ�A���'�3��8���| I�F����^]�"t��j>��j�u��<H��^ꂙᢠ��&T�ū{x �8��Z���W+�p6p�l}�0��f?�ܺ�h/�km����$��>��ef	 �s[kO�%>��NDT}?T�;A��8���+r͠�Q��$O��iV4D=�C(�}�����3����A��`ю�
��Nx�/^��Ų�p��#�ӄ�~�#��CÎ�©>��I�z]��a�M�'�H���(Q�m�pC��+ܱ��u؃�`��j�n]ҽ�Y[����!d�ۓV䠰�,c=�-����y�Z��)��i)��i<
��ݰ �j_f��xx�I��o1�k1�r��\�hzr.f0��@�m:1���}O�������.����_��عؓX��M�-��f�B)���ut���i�I��"N�i9�-I�j�qB�s/�P=�k���=Ӊ�O�/+���s1O��^�������։{���e�I��:O�K���W�����ʔJ0��i�+�'lb�֕e=&�q�/���d�	���/��Д�[6;䪋:�ｉ�&��M5@v�>E���(�T)�?(,�9�>�O�96�)��JVTpC��e2�%A��Dp���v��T���'�JAЬ�P
���Wv������T��e�w=��+���ǔg�:m�0yW���X|~�O<���.�sd�lțt��3�!v�`��ϫp�?c �d!&J�\pd{�~[JXǀ��^���0��9�'o����ɺ�9��q�^��0��m�J�A����*q�o ��J� ����Ȭ����$�LxJ��X�%�/|_�M��E:o~��XN�������B+�IȘ[�	Z�g��
w��m���g�BA�� ���. 	���"q�7�<�u7'4��\���u�]9�x����^��&m�B��!�.8���Mr��]3�7�$�"�2J**��C,'ڂ���mA�9LJ�?��z _�}`�z�AºnM�F���ܢ}XPi<�B�U1��VNƽ���|k�������K�M�QS}�����GU���MԞC����*�DљR�sOV��7��q�ָn8������7��������xV}��"���������Ds���N���]��Ӟr��g�r���"��wN���{�S���-n�E�����"l�L�s���Բ*��,3ɧ⎱�m�J��޺l������h��Q	�G����"Z�N#Vw̅�p���+0�q6�&����<��+<&�4#��Q�X�����9�1���L7�-j�76�A�	&P�(���Ao��˔l6��R,jejS����/uf}y��0��jj^����Z�N��� R��0,I��d�jd:f܈Q�t0��<�A�l7��*ȊУ+����p
�&.\ע ��U��ɄAٔx�f�2DDOb��RRE���@GB���`�Z>�ɯ�����_
���ah���p�L?fb�(wq�Ӽ�9Da���j�h$�#�#���'�Vm��.�{���!�B���99�	��o۝E,��ꍺƼ�6 �8�c��/�C@7�mR|UK�6�33y���\��a�E4��c�iծN܍ˍ�H��O�s�Y'	iZ�9U�,�k�&$�3�nP(xt=�`HǮ:�W��=g~�B�ڒִ�aᔃ��ȝڀ*���s��=�e�e:3��V����f �ga�[� �q���v�&tϕ�Ub���AQ�p���&�5�O�R�%�YS#�[���s}s0Tg��Z�ٝ�ƪ�S?��~�<���F�f�#;�=�~{�������F���D�-P�"��}�s����F(�J��e���Ϥf2�gף�qs�
��mP��,�Uh��JsD�]�u#W]����ѿÊ@/r�l����^FaY���f��������"����#���)U�4�{s��\ln9��]ӗ��1�B��+�w��,�Q�x�q�`�u������S����Xr�Q[ta��r�Q_/dT�!M� 9��;/�@��M�Z��s��X�j�����7J�Nn�vF��ذhSJdP���t��ᩲ�Ϋ��;�����] \�>��b@z�f�E�P6���54��^��/Rx
<7��lq�[��T�_�IZ������6m8@.߸��)�Wc�T�(1���.�wG��*U��᫣F�`�B5T���nrJd;	��e ��u,M�g˟�B��`��������z�G"!Us��g����!�QU�]0��i(��*� ��*��%s�$��	
�A���E���)�^��D����7�� X����ND���u���O�<E����}A������	�!3�����2��U:�}� ���A;����W�v�Ңh��i�|��ק|L�1�$�Y��S�O�}���3����:��/E�I�1Lޤ�-�^�qNؑ�����~9zG���`1{Ke�f�ݙX$䁆�D�Б��Z:�2J*"�(EI��ʸ�Ui||QE�y��X�T�g%� ZQ�ŋs1;�5�i�G�����J�"]o��K�v�D���qsb�l��FN��3:���f�P�tK���*i�u��[��m���	��|a�d�◗���(b�1���>Ls^�$�8���L�^2���Hs������|Au2H�Յ�MxA��	C�\�aS��rw��f8ڠ �Z�g�o%"�*�7��q�;H��{w�e��u,�C���w�{RG��u��o�(x����R�^|9WO�b�96m�u��jg����'+��w�����=��8��A*���Hx�`��j ol�τ0���>�_kAU�đ�.AY��.x�kla{g�C+�%�