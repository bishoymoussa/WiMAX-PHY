-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
HPKjFOTFexjgm9iB9dIi7x1Ge2qvjQXi9YgE1XdMZvi3RriOUdCsY6zgxDjjevvaK3CUkiFdTf1M
YyVahUuFpR1umxQJ5axU2YNkBoU+AZ1jQnmlqr+zd6ryvY2m2QSHMhl+OH3pga1+9GRu3bG8+whz
TsFmRaj8poOmv6vNPylo/tJU+vnTPP4d1iAbm6Nc/6MU04FrAzR+diAR3J+ho43HJvYDLmyyCMF1
d5GUHfBcS+g+Y37pjafRsulL/hGvhF3fv6mooWfWHJ8H8F7zFMAP+O4mfyfCNqu4rFzS9gsq5uWW
kL73EPnxGRcDsOH0aOFL5JqzO7u+e9h0oLm3nA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4208)
`protect data_block
8DgCEp5Ih5qEtNwPUrdVBX1F0pTB2RSE30Dqv2aMDUXJxxQJmB8lbiv319MofQMbvir99vJXIXmN
bVHPCiHToYRAv7OPbHe1zENunH9Yu4o7Zn6v+lbakWhEMrFsynAYexzIoYLmax2Cns08uGV7lNLw
q/kYNgkArkRmBxVSsxdbc1dyOiQMESX4RknlxZ/YXP454q3++UFF5elGjHx9ztNX14Dzd6wnwwHN
CsesEw86iyeRxcWrdf/IncwTh7xkYViR4h/yb6v8ETYuWBBhrrvNokQSYIjIW1F5H10Y5y7v30/5
xRI5v6NDz2Z/YvEvPgaORizlZ1WLP4sInlWgP3/w6VTt4aIUveGu6pJRMsndpxYn8RPfByqWVEWM
iu6vwQ5Lig6AeuZ4vpg3d+WS7Zr8F20mp1m9jIoL0kgoqYFTImiEvICgayvWsCs3bZhCTGyus39E
SAPYHiU0p3KOQOfNcfM1Wh4f1PHtPUvH0LYf8GHJC3Qo1hsgi5xzKnBD0OYwTDeKQ87+H9A7U1b6
ZvP9X2LH5DJxsTV/BVnoYG3psKEkOpBL1goJ1RR90tGDXaOvkOJOYIiroLWvX6c7ho72fW44ZJ3h
mY5tNgOSIeg1VbhUe5oQSDYqL1vxE+n2M8GvCL3WAxQRBCOOgoeU1c7DPsk0ndLpytDKsRAul9W2
kS8QvptQGDIJ7hleMXEx8a/KKXshEyZSiPXeHay1MFrPvAE7r+D9C+Y7MmacO7V9p2etHTAXD+/d
oXZjVQC9Umm/8BNYixZVxkNU5CrLGAQ7Qp1mw3TZcY1pEhbyK7EoJQj2YtldTcCAe2wOgsLiR6hB
tI5qsB3qZ7gSRAvgNQandjmnbtartzSItmF3w5xZV7/3qz5hAIm52fSfsGPcSpTqLXQq68UaxkN0
SJmoWOtWs1xUXz+KLZq44Dle76WKPZ6CdHubwbiH4fvlbPapWEDtt32vtBnv2yK5afdDeOPZISzm
9DOltDQ46eaHQyYshVmqoIklF2UTpMzdn9q4ztqUsf5kx8PROQsrNbUYJIz4EWY0s8FIHt7F7Sny
Mfo0mXtAdq90o90/aJlD8tlJEFSR+kYBx0hnQp2GGUjt9/IqoPZ80A1pXwKo39EN9ZL+vPqLENEO
Ot5tle+orPDdCTxTmmH1+FdVhUIqkHES2gUNp0xgamoQhSJf+QO9td6QfcuObYGwwmaz/d7bAIaJ
orNaMLv5ScvfxdU2g7737LRMezM/BQT8FXHlxfNn7Gn6DfDSTQhvIWw6Xzek+374Tj8NYCp+fhsl
cOktwr1AEIRVsAxmRfEKtnuztZ0deszU1znRynlJol7idFMRoF1eHDWY7bwJbpQSS2o1QJ/JUI4L
YZ5t275u62N6ZurqW970kIFKfJQPAbJ37ARySlTj9gAn+uI/+QmxO0+URAASAB3VoHuE2UdV8DE2
cOTUqb6NBHy6/DVaJ9c2bGs7jJpGBtp3n+Ayh5BsyAExRLpJYWD4fbi6fAzLkMEVK/En5iffRe+J
ZmaFi6cHAy85mf3Y54WsiHvzW9zcnRixwqcBeqyxARRI0Xe1ONaM+h0bjbJsjRbY1O1Eh3y0U4gm
pgNP5hDL8/L7E4S5VcG2E/e4ggV7oLIb8cw9NEGAgIJhEryyK/Q+01KNAWBn0kOkj+eqg81BNEhl
mRgQrhReTx7t29PE1UoR9VLWUSoxqOzHvyTf7sQG6ta7c0/gIKPhqSsUCX9EKgDz9PfmgcMaqvFm
lUPJfymbL8BIJuxJV9bud7zS52tnnRlxu7zT7T6X5h68kJmp0dEX8CuBBysx2nQ+esn3bOwzOrFA
QrgZoNtz5RSdYGrY5zoowd6Bilc/C6JXLj6+sVfRaH5nzqLn+3ymiFgZPS2qxx7vz1FJY+aftigX
s8jqiIm54KIbozQ+W7/skX0fM/81LqAtBHsnnU7U+ECU2UbbFcG9m5qTddDFF4U9Fo/fK32CBu6g
/J+1oAMdeIN8Vt1JmSs9ia554AYhOgwHy5zx7z2PnaLQeXHkNNV0Dp+20NORSu+bB1gcSK8L811Y
QVvBBJz3tK8+U1FJkY8rbcvThmK5Ue94qe+TETrfJZVXFjzw0KerPZfAfvxi/+n/P+MCPmm/+DS+
ieq1FyenyZhUGmSpZJT0Q9h3zFszy+ruekKekovlLY76REwR0yEM2A5fXSuoxQlE/Aef4xXzonbi
ZWb7SUvluZYSsonO2ion1Mh2o4GOd5RQDznAxeYp1n4kEKTSCves1BumJC6GR95KVRsvyGi5IF/g
bufvywlMr/AZ70guX7RLHfBlZ5CBexPRjJiRtu3d1cvmal7FE8O2SA+X46Zbh2+pdBbefwBPCQU9
TlYN6URmvK24niqJCeurr4TRhH6roM86KlfI01SE/I6QflrNMsAvSwRmFxOUJrvfG7N4+KNa/qJu
SXBl/sNFKooCaPp/df2vP19bvn9V9pYD4rOuJsynxtqYytQw0sjSCpUmrmrqQ4YfBjsUs8cpzdUH
M9h4HjKkpld4FaUzH+9um0yA6BoQXiqCOqwCLRJsVJ5g518conHkmgyNjVC/vTvjnMjjTXUiPjFh
56euUwClJtgF3gn9TDzp3BdADZlfs8PuXJeULg3d4/dLt7QTxVPqa+lIFN2qq0s/IGZUdn70WIk/
DA4Njg4SUI6vAy3whmh0gW223NHEvIVElxJyjLHo5a2qvE76WUhQkEs1Wzua5yoPnnMb39rIlWzh
mGRs459ylCZaXApGsD0uPlPtONDTRGpcT4fuxm6yIgqliPPsLt2a8ETc7SUkstAzbhU5Kp4gpa9J
yHOp51mWKDQxna6LL12x5asnyrcl9PFG7iyfD/vi6ZwdUHcorGqtd8DbjYe24QEXNRtpCxgGGVv0
272q4SXtaCz+BNxjcJiW++xaQL3Pu7c9kUKNOI8ntIBp4tWHXIL94kdLO/Ds1Zi7UCSzpEruxiSb
zTq7ryIk3E7RmQ06N4teUa/GVYGHcSsXW0y7GBokeOmDTQDdl0H0G3KLrLRA60FnPTt6hz9awgAk
+WbptNFZVo2axsEa0mFwSAmFGiQ8oUvufXlV2L2yk+TDy1Nr7V/ySLCHOGYRAry/J6lWQd2tJOCa
9iYWVGN+W1K3uZ2r6AJaOMrr15ZYxfsmoJDHx1AHWjRpNQ5USoA/2kOGkCJmoa1uHYFnmvpd0frg
xdLZ/2WqBO4ktQkoU7p3zUnXYhgVGApCCoo7XQSdfxa1c6fAr64hq7fg9qE2SyMkpeyK8y4/4uw4
8LGJ5r2dHxAsdPA21TSrdxvWdccLl55X8PkRtIfEElgPdUjDjI0qtbLDqvto3ienEbIkZpnvPJHm
Clds1o4QRLCVx1mcuAA2kRL8FfyHDAsqfCo33EEgP4085lf5RCCPDwllbZci2lQaaa2AsDU4U+iy
cFNpfgOsHzMpBsrD0buApFKzrdUb00inHBNcNpuSJcUZj9U0ztBInVx5QGLKkEPiQlbymwP6qXhp
Ze8YemHHtr0kf0UGpn2R8OEzfXylpYQAfwRIC0GTf313h7AiGRiAFN/Hc2gdwzClheieL0ceAS6m
1ru4BJxYubQN61z1orK5oGVr5OdeEhbSkzp8e4EJO4uYF+TaKjYU+Mk4tLKyGVB1aIfXAF7Cpn5k
FKfszWIJnFiwmcMTEWFEipZw5kulQ+2eWHdzetgwH/6eiBZozWW5I11lEnzQ2aXrwxlnuLBm/JQ2
BqQnoOhycbyL2OHYxU0BIBWRuUNrxGmhdpkUxhKnBWTqa3ai5WVhneEFtZfWUFaZ2B+r0SDmjmDg
gms+w4TRrMI+fg67GejALVkBofasUu8bldWetup8HS0owm88qnqwX/g9uhRDPyNsnlwiPdy1+e7s
KPJTNN6gKB+hfo6mqakNmp4SsFO1U1LYjAljy1eXUA3Wth3DCyG2XWD55wPgN2RUUs4ERzPWoFhN
PmM+1ChttCvUFedsejPzEkFWFND5/Peo1JzcNb3R/R4YgJMVtwCABcu7Gy1Rjx+wJvHjCXWiaOhn
49rEVkzfmX2s2nDW1Dy/yhpuLBE68nv0Rf9YozYgb/rK/p24XDq9yIGW0sq63J5SvyDytc5PQH9i
d1Mh2/Qz9qBa0ykMrzykO066Qb9fYv66GzJ0lEpaBmOnOg8vbZrTRWfQ/j+ox0gv8eQtYGvi5hI8
EGcrczsb+ILa3QzuVioRcGtcyroaC5FwEhbiE9KLdCvH0L+lCiXtw0+1tBTPYbliioFwu1KVewYS
YfLP/dL6cIGH8LNi0TJuio8fsOFW32mEhwawrECew468pEWWZodbIL0M3pZYB4LNa9/TRKol1S79
YSUvVMQfPKwblMj7uHO9v8rMcOokq8JeNQSBYtoy8SlLZcrUYOK045qCkNUBElCekCmTl1sbdGsM
M1ZDXsALmJFhDbGV3pEFnQolgSkQAEFqapHogDwzW6uRLBAmq86uVuaUuDwjMGuXyscUK6488+6B
curH+Vy8Y04uOlYBYnI5YpHq5J8V8PELEJRrUdgKZSbn5AJKK/m3NDN/mYclwW6kkh4iy+STvgDi
905ojGC6ae4t+m61S0ytiPHqq6f/w4VvWNQcay3mHyJbLJeLAggDBwCGSAigUsOn390lD8xCYz4p
JIHMDKBMvDm8iombrHJtV1LmF3HmlZKT/o1Abhf77fm6Be8lamN0y3LQhhgeHblNNGY5AF1VhL9S
CrGD4FiJL+17yMVUJVAUTcdaEsPhSv3JXLz4OP4NurJJQV25et/OfKWUQ8Tp0OMU/fdJQY+FE7Up
ZSPDl0/fmaTQ7867uFznsyx1Jz2/HH+WerbD31oJDy5bQFNPBrLydMwPyECLUKhX13FZYPePipne
VtXZHQd3+lx+xv0aea1cnJ/f/QKrdYWHHsFD6JNoD8gkhgYgyomgr8Ctcc3lomR7lPRZmsKCOMDA
ECX7TrNVHAF16eE79dpv/Q49wfv0schzCRlU4NuNjDOcCeN43nm3KnwBi9ex7XhukvHuvbFmWtlT
pboN7jOnyrWlZoEZEZc8dn9me9P8IEs/ki6onwfWKqg/6yrxrW4y/DGU4Y+uDpwCvVOx8ZemZgXN
/3PBoYbtyPWsy9Ga1gZ8FnVGLqkNOOvHgXdh/VJxaR6gj4lQdmC9ca4Q7Kf6YhoWy6OpJDz7YV3M
/spj4Oq2V0I90pgBGITfHtxUGl/BGqWE1VCeW4F5AXWi3Mo9b2bhU9oLs9XhqxzyfpUABP2hxWf+
N7zyWKTKzfu/58Rf1X19jLcrtKiQ0QPMmGVL/Ngdl19dcSfZ0eUdU/3YIiG2bfDAWR4kj3jqVAPy
g7W2eLwpP9/RtQwe0BSYmeCIsbbffyBQ5e1tkTvnvFDlRaRSKxGwfS3u+8F+YVlZHpy2+AAx2eBK
z6oX7L/0Yhac8OROO6O1vSV9k3sTmBFjGKAYGk5yNbUwNqASMH0FMhCi0+7xe5bk82a9N5X4PpMv
Wr5L1jriqZK0+8Wt1YWRRM5srzUj19KNX2ADSuJq7EFjfVjgB4UbwL74XJiZF6CdsxBiCTK/WiY3
ZXZyStW2rdH4+RhoSO4xYRKI6e6vfjZU+8OxCnqVj7Wcd8L5MA0OOS9UyfxqAWo=
`protect end_protected
