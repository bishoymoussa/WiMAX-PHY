-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
uB4jzOjePYzsK4yKv+D0ChXGttonrfA4yv7D431/FdSqnMKrIHXXSSBk78Pq+B3JYi4g5DNoPzJL
ufVJZ7sx72vvkQmX6c9jGUdIyoSX4lfVrvg7+YRuC9MDL2g+Qj8xhYif4xUYCpZ8/X5M63h0lp4L
9Y1xC4lf4rQgxEITFYNzBf4OrymP/s49U/Cn5ZbxKbcGUtXFV1QjoiW6+fS40DkkAUTOghFA+r9e
ZlZtzqKVf1tLhGkwzmK79lVGADUT3Ofuwnhap69gbS5+X3LwX96xJWdqxESuIkYzacIGPQZuJGKi
TGPXrNe2rdoR98FSUEtz/4njIajggwGxGN/zGw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 71328)
`protect data_block
srdBF7gDRJ6B6EI3JbO8hcC15SHJJRcIV6cUGywZlN7yo7TKv0fqm92RbLS+OvEj15qkleWy7gvs
q4B97IGoAx/RF87awYhV6KNoTCiZ510e67GOFw2Ywb8abNe+a7Oo3ERp72BKES69kekiXQdvxSA8
cCAljXwhwqxjXe+N8XrUUHg7bjkjlGwaq2tBWe7bETeXbMcMDDi8ZAvRCQmzJ0lwO7H0tb+sTX8v
TgDzrQ7wLa6GYK3nOHceKgjkizQnG+EyEFvNN2RytueeUIWTs/ayD2Xz/ZLiRvHuu15gkBh21pwK
hITr+cIbtBHZK+V9KVEi7NqWVKFaULjKOOyxNrmzY1v8hJEDmQi22FS7Ir3XEJ0vi0UTbcnliXYK
oArpSSRRY2OcUed2NeoO7FHzp4Em8H22JJOBbIuNQSvhpm3h2vJ8A1KLh2G/JV4qpM3dVz6D8LY/
ovBXkl6s5scPuZBQ2zaQt5uf4UP9e5pR8XhnSr+7820m86UjDI6tY8Rp6PL4+WkZT7ZxK/lrs4mz
XRGAR8KfJDtfdsM2Vq0RSxBFqkU2jRcB12vXBXBxnYysJyxXiiXppTPFVDf2FjI5xqRWfULQ63eY
SjFrc/abAZIVXgznaOX3a06dIm1J9U+yjXZPTrHNsXLKeURNW0+wqU06zgULMyJct6DNhJkH84Ra
UsMeo0zIh86lvFPMj1rn15h5EcdsqnxUYXK4k7i6Lvyvee6FP7w7W7jpdyVgSrC3HqC6mJ8DM6ox
g3d83Tcold1aDoVL7NvQY+q/PXU6Y33ssaqFOaXqQJxXzM8TfmLv4XHFzSUE4WEHuzJzu71SMksL
Ihu0lqoE3aWtJ18pHW09ur2I35NQU79IV/6SDypxOzDN1EBzOReUj061v4gLg8Cy43qUVXm+KnQ+
CDpMHpAUFn+MRaEfLBu36pU4dMiVv9vYF6zhwINT/yLjZe6eUCcnyF62MfiSUeIcytW/3JZH5udV
T0YCiB0zjYX+7/8ZoSn4rdFFUEZtxkZ+AsZpIKKuI9ApSuJSiuFHAwqtSZSRhEcw+yEjVgLhGpLS
xxYFYdWVMsJigEhUHHem6fanNSmuaSIwOPj9Qe2JNUDKAZBUjWVMe3c5Ja9W/vChXhl4doD3SZsp
wtqc+J81V18kO5TU94CNYfeJDpM7FdOCIpy2QHjdM4XBqv4kc9GA/pWD6Lfds4dgr8cv2CBp4nij
P54SHxYNY3UtiKEwlD+hfZzZK5ZX/VzVC0V5La5QJDIWZ0cS+WmYPdU91uvoOMteXRmvOzJ524tX
P0M+NcX88FRm9Ve5Ce84wjfjJh5ZLnlzu1WI2LmFV3J7npTw1mvz+4oGhln4CUjHhcPjAp4IAKvx
PyCb3FtaCdX4RjQNkHQwN1uZDlAp9oEKCtWy1bX7jDywjIYRtlVHwbOQNwI54lTwsG55JLefW6/W
FeyPfXffuUYHr7RazPp9gqx7TZJlnYSTfyjVw4IkSXF9FC3KVBNe56tPQLpazjoWJD8y11je2t2y
joVjZR5w2+6GK1Cgv9fzKaVOH7beejceOJNFkAX3ZCLhtrA9W430O4xyicyK7aMxaktTu7nUnx2H
aCXx+seAAgcD54dT/pkj6E4Ldk1Maqt2tbJr0oGEb6Wsu3ZN+13/DFL0nHEVyiytCytPYN+usL51
FkC/XwUHJtoIL/4uUXU/hFxIRzK0AXOOaHgBUWKxw9l3KzbUW91qdCi5X/FCn/h02G/BKqcpwnwT
gkHR6Vlisw76FK1bAsI2WYPuo8e2P0wtSaIYeV9GHO25iMq+aIJgLfkdZn2kn6/Cmm79xaIgXNKP
Jyi3fJfzJwgRAhKUNQNNFOMT4Op/fHdO+5o9oRI6T5cCPy/1vKW8CXEwRUtO4me70628Pus3dKv6
+bUeY4emSy9HGEpKNZSHGFB73lBFzG/9r0o0bt5hV8wrLR22ojDib7yhziQjjOZRibfGBuojVpaY
oRYltKRAl6tM4Bn8R8fikrGa7f6MUXToFevh5FwD2iDLbLedKonlCjBvCvwB3yZ8jiOlrd4GFiZ9
Eez2ofNGoM+nUUx9TQ2kzyFjLSEDy/CiaG+IgV3tEhOFSiaD2wIYdzY+J9KTjgwxnzD2wzc6Mzht
1lGhtcoVTuCDa+O29vtXPyKe98WTrwclL8v8DuVU9HwpRMvWzQeR6p8zVJoFETdT2SlrRwZgP4Jj
Ops55sTpUYFwyzXC+T/wbqFswa0ozZ1VFZOK58hSkwu5OLRvJLN/zXdAl6RTb3/1Y5NF7/GF2dvK
ehw6xP5ksjA8eWp4DL8KiHkNEFQR/1sLl9WnPV875fcioBqEA4KiY1oSW4SDV63QB0rRqCab47G9
Ii8BpyPscSGoyurXp4z2w3FZdr3pJ6X2wFDpdaS6ujBQvNULq6KVEIuF4MBJ1oGw/j4R7l990Sh4
m4skzqJh8rOrn9rPuc87WBXTevkXfg/Of9Kd0h7tR8cTLmGYjpJ7Ak0fJFV0aZl45zmCM7G/FuW4
/0Aaw2vdjY3L1joaUozl6Z0GJU2tJoawvlJBLsh7S2php0+5mhvk3vE28+GNlqQ4hJkYjC6A6C64
HvbCEW/YIChrhFKfDGbyRYjYONwCO/0j8lVd7ol0sVHScEXUDQmgYLYw6JgJk6sQjl6t90JYj/lk
s9IaJSgYdRI76M0OO5S/RbuM2rQtKLHY0PWJGxi66qzMRsDNE1wT//RgHpOWlVvdgCjizQqex9Zd
80iJYGhxPc0bHQMG6XnhRvGCeXBqILxdr4LBCcuvlNSayX3kPgrtBsKCEJ1mjhY/RMHP8XPdz/i7
athdKz76WGXyzdf1lSIuBVDh+e9AtDLdiKd30Zo8XRlQEaim+RpNKEUs9Zu0N4nm2/pbjyi8sT3D
vrshEuYqfEfZik6+N8OJjJq5VeklvxySXHrZNHSjWGEjZ1TJCHCxFUFW23M2m0Dizwcqoj91xfE6
D27irBe3chT4k831Gn6sgaFdNwYBmsZGkpW8kG7dK7TiQUMjCOGqXkGj7DwCa36QxU/ZtgA5iqfg
iiPiUJSYPE6dEoaO0vHW/Dt+rWa23tpv1thgC8ap+kCaC5U1UmQzPZhIAx8bRJwd7zHPSZnmTpvj
6PcXiF++z96pwcZJvmpC23y+16KYCPpl5uOr/gc/6JbjBIijCJwgPH+YgbDFVju0zEUNuX69IOoi
jRhzNz0iyNUXWtDBqS9e3fFj1t4v+yV7V2uduWzl80NEeLTAJ5z1d5fRCgfnto3QiqEfGwSTBQi8
MZaRcO99WsW2qQbPYf1/0JIBZdoZDNyoEUXseMsbknr/MUUOP2a0r+ei6qB2prBn//PL261yv47A
7yOwyP61JffEfxQKqy9OePnSpIb+Y9Ur76AA7/wIvIiqPkNZDfVN6UEA/xZ4RLs9dxWAzBTDJ9F2
cO4tvvYT3v19689o2TlF+UDDTB3CzjuAHXMEglforD6sPyZiUpmyPS594bV6t2puluoOo3QVZTvl
Y/7vfk9EwZRtSpMeTQaFrKWMxzg6q8sSwp5IvJK6EjF+rwzk8goH+fkgnVwYjMZo2oJnuK5h4tav
3F7m4GZVqy7ONFKsuV+p25zMc3IqUhaWQPl0Eec6a6DThoW1CuNFJ26l3scapUBk+MTLI9SUojby
hxYPyUi0UOqVt9ks5bkFvctASMPCeICWoAz3J8zpejLxcZf+9fvb+GOoZm5jXNB//SvNCCiX31Ra
raFqmx56zzf7rV80Wurz9jCKN37DjglST2eBlSc1OGrba4GHKMgOVaI8bOvi1b07VO9jnaIVdYT5
nmSVyyP9R3pSzqIt/Mj8+PXZmLWHowDiEZFrQpye2t+TkX6TEMGwJVw2jVW3icSdEIqtDiu8R4Ka
YGsGE1ae0DLTSUOfvGD6u9nlV25DTNCyEqMRypeXoaZoO6sUSiG0jUjxVFTsbl6CCGLGeU09Ox1+
9S4fKRzWClrI49TcWwOrY/YLyw9axJeXZZKV67x0RCTht7Bth+/me5GoHAf+3QbXrQzdHiDzr/WL
DM1jqV4aREPEmKHzwMo8C/2hrDABhhOaIxCv6agdp3BHM6pJ/7sZBV4imyb+WVI/J80HPcXQkxCs
L4OLrQqfyFwrftU58S2lTMWIUDHoh+Zx+STYq3U9GBwBWQ7GXykHP5dThvMuniPYH2G2sSkDKTy5
nHpEtWaSmmUzMOmB59PZ6dLYoakSGTrVuTZuSlZkkXMjHwHlSLdGwmcClsEJ2oX+GeyTqhKfBT+T
mhbQQ6Ij25xK+W4TCGLc97UQI3mU+6+hwhF85sklPGs2Lp0Mh6oxC0Bab7hlte+8av3bSdfeQ/J3
88GCCpMY4inILk54Drx6qjY9mDYvAI/nraP9QJLGHThAHzqJ2iMGv7mNmUBEK6SULQWPGTm+c/NA
7/JJV9TM2huDCV/4BKf/XIUeOMnKrk+H1IELzQrjVAQ44EbsqfquSjxrjNnjhR2eMS3w5EN4agnw
Bs94E6W9gCjUEJIApg1A2ogrQJ1uOzwRINKM+xQbfqky1ywGvrphzw3mtePbP4zG894AkYYUISEl
eLV85vXvQ0i3rN1q2I4PFBWOZFpZR0xVlfGIMM/hmVvkm1amN4WTQvr22F55OQbUhAxpGVrFX+7b
crZObiadrC0u7gA5OuD74SwZjNmebMkz5ZJ+aW37rm8bIdz+fhBCIh5Pj2X54dAvCIh8wS73URAL
SHQbcdi73IanE4PkT0/cWLqRPi0Y+ZU2hjBdo2d/kNb+o6IvMofiRZFJ7G3LdpcsaPyg7YGgpYYr
mwEeBAgXS6ee7VS1EkbSuAbkjQw8Q73oHMzjr3y+P697SQ/Vp7HSv720me4ZQ3bn3Py7WeLakdFY
24M1w1gs9pjWxTzmtGUn01swAOFmsWPFkFvqGfRcoAWmK08Z1KLg29iaLsWEyx3l68cmjub7x1ji
QIY5asIyjDnBJ5kiLN/J3Hxn743w3ScyB67pTpHS+I0n1iofB36npjZ73k7eLy7VMOxKPTE7HjEC
gnZ3FLBUe4YHdNmN/svuOQbevFxQxek8Giab7TnPpkXKZe77CJJqNmbT+3zjPs1vjuck+oTbhJIJ
0fTZN/vahpDem9xtNr6LKUxmkEaGA2jGWsMWMBpdCd0M7dFzBnOJGgo772dyJXRlUN5k7kaqJ/8E
kkLI31AXVE1rAxgY+StV34mRO85DPZ5WZZtcYt+0ULBPZgRXP+apjVMw/sZ7ljIIQ4rGhr9ykJr9
sESim2FmQCnU8T/xUIzyASXU8wgQ6uC4xE/OeItJ8T2QQrtrzU8wQDE63V4ymG4TZl+S4bIHimtG
jpl5vkVmC/FQcqvAEFZJgDCS079QT52xjAyg4VuLNIYrBMjC0QrN3j1PtlNSahX5yzJhNB7H9dxR
YOrKWSd3VtHO81YPDwNNUpjZUu0tqWLxldKtgpGCEAR5/GUuFh5pMD52alOfk57Br9senk0D9hcm
/UV8Nob5NoZF4AfGJ2OBw7AqY5WKTu2NL84LjTWmbEsCclVl34U+wJdpHY/BmgvfC92Yg6OqauvD
vLUFNe0KKnu79TCVnhXhIB6GEar0PdZNOVZ0sIZDFqNzU5Tv0zCbpMUAuNpDFKRpbZJVMXHWDt3j
xDCZeUDPMb8F1wRxZDkVeD+aqStCp9hrlUhhvPTd6bdLtoRK25DebcC3NdM1Z1rUfOCTApCodKRv
aYcCUpGTZd/Xuej7SiT0im+/bxlh0bs/WA7GDqd208aaSNgodfFiSmvvwv7eZKUuvGxcwX6pmfot
+fk5DON1IL/agEYAjXlwzRFPVKFjZpLSX1bldGEwWpvyqIiYNoNzq4mzxwfiNCdsVZNp3gRKSyjf
/oigMYYmz+TQeCbJGQqoujiejB1W9JYiK0B/iMNxUJdZVgQT5tok6eVsEYxqZfQ0KIL6YZtBpmcI
1LkJ5ZI7/P34XhKYhVB/VzdWYMcIU6hwQstC3ARLKgu1mfLGalwuaFd5N/K6hdCGH39462zCqNGF
xettgAh4kYw/7Pa2AbZdwRfOOjnxmI1vZ1vnDZ5zb7Kn33Ant5P6Lu2mBoZbjUE8wlTvIaeB6czy
S3OlzyEwL5m3xsrC6y1et8ZBbYjXvoSL1K5XRDgtcYCey/H0iOtnUrptWW7RXsw1OQM8qjj2mDd7
MACFKcOlC4M1E69otDE//yUBPM83zQPh9B2TQaenwE7q0CA85IgQwqARBIcAOccSv67eQto2AwkU
buOOWAgjYTbbxEn4WYj/uiAEqIpmK/gfEEXCK7XFS2ZtU6Lbc1kP1iIgsnj+QvpyZlV+toEzv7/+
jd/wAlTQCcGEBQlyJUfoC7P7ltW+RjLyU6fxpHPv73t/JTaX5h7EycclAza1eDhwJyUsZ2yMn0Hr
2Ya5ImNaEGznOmzSKqFHldVTi/TJmQVaeefU409JB32ChDdUy1xqQHuCX9i3UrzVk3RCxVXD4/ht
Oml4OugNUlqypewJ0E6r/Wsk3EXMKyS73bv5ARK+hUl6yVfXRO1HVWfruSrn9GlHao6HDn4QXD0f
NS3sOrXP5XiGhwRtASdump9t8VPZx4/mc93EiT/mDrwVR7rbIAWtoNXR3raDUjRN96kdF8faMOG/
XGYoqCAm7McoYOtvPaOktV7YuKPSiutbGFWM7yRM8PnbomRLbHcmoOhF48U51zGZ/q1VT20Y6lJH
1xby0uDIL95q4vTnk8CWcPRNXTRDU/yVm03jZ8rrv/iMIlfSrMr7vYrhZTDJNS+RySbYC+3H5quB
VzQ0xrM8jcCpJoEfhC1y9s4/djoYCAHrJXwP6b3mK8axQVNAoswkScwiUJ0yi2fzBA6jKIC2N9dQ
7xzP1VaauMGKZF6sscAJCHoxCGijy9H4y0SCw8HEC02x+gn9/uq2B5IDObYPWkQQ27zE9pDOsA+W
XqAayU1aPvOjvl3nhjmUn1ulSDKTJocXBVJZKMLoMNTjNJvOTxmYqXnxBpsCs/KVi3XpjdOedRwF
WxeLjM4v51v8WsJuwnoWOOpX1fRScvHBkUMs09+5gMy328t59CBt3IOSCk9nG8Gqv/HnV9g+lOKb
Ix/oq6Kx5XkDd9BkZ9bkVppmQSrOr2Ll82pazDM3GZFc61vU5fBUAiUoDrkhz7kBkE57BajCKtAP
6pHuC5SRSJ+765wxT3uGqUnBkunmJXdJQ8B76OC9zc8ietVf/1rA6u19j9vwGd0Y4/0TJi6QfXby
prFasG+CQYEEk6KIUOMEmgRmNeBC2Jco21QMCkIKRgBz/7qmuiSXAmJVpiiP98p6q4OweHhiVZ05
yBOy/oSnvO8Lt8zcd1mDiDHUAJG6hDZh3KN7l/hLYBiNgF5YU2KUZx+s348JMIbyGILwi0mFo/zy
lHUIB5WzZt6w6i/7iwdhkVRJ3PYYrDkmwKvR1D/PU5wuleTHJoYE6uST/bsr9oGkfjeXQUfqWvM7
TCcTCQdsLwtUwit4Rndg1iQhpkEoYvHy+b0KI15JprLYFZcIEWEegJfqvxAUaNY3Tbqev9KiI7Dy
taFzG1CO8GLr4PsPGCFAmiIIebWENOObk3tUIvOpUey6TP1+BSuojcqtnHAlvDlltRM0GfQPdTmo
gOQNZoY0YL7bRRP654GTIqUd//6DEMLg1uRNRtyWUmVjh174KRNfHKLJVo410XqDkclsawbn+3BH
U/HF/t+7jTLsVnqlP/D8Uoz7kNjO0IUSMSAiNbYjX48WLemCsLSKRp4ShqYeevE7zTGWOrgkqBxx
qFnUglJy5Zny3JUTCMRSnEnfsIPRWYC6+8x/VVm8bgmjIBslRZGDvzwlUHdka9Cy7q+0XRmWATaF
WAnoJZrJjSorTT0v4ZxFW+0psp612+Hx8v5+NBaF2HRqOTKaH1dPhFj5/527MEBUbwUWMvWM26GA
yNE/VX6i3uVARVI35fZLj4cym4qy2/eYh+IJwiF4VHykdxm9l6nN1qhaxhOm1IGr5Ta1wL5MAa5E
qwDPTD1TgBE0PyS5W/POIL+kH872XBVt8yzQ1a43fis1w7byDYYITx6smD1yv6VeQcxDTHNrqvLa
pTpuvFT+Fy5IBn43+hFQqoI+UVRQLkfC6cfKFwddOQLpDzbG9Gk9ShQr1ahbQNzOHsEfKIChQoVO
1yccBKfD1QLHdvbfQitwGzgczMCYNKVN+mHPZttu/qdx9BlxBNjWuXtkM3NnNOmtQpgA8BSRL+M5
BR7T0+28DxcIljrCYiEIDcWyz39ZddJu3Sc4YyalABQy7kTp+UVLi3NRWo4v1Ki3L5mJ6As7Bmkz
N2Hqn5wz2tJ2kjzb86KbJtbjSj0zKCI2vBrioEGWa+wp64e07S++xfqi84wCbQ9t0A1UadFOrNK7
cpFhfAwm506WD7oIbOQz1s3U37w0UNmdu4WIY98LqXRhRJrPCHlbRlGpus+/5IkvfxqiFnzGfoF1
lg+3aOF+5xPMe1jei8vcNvOjcIHAfB4uMmzwTwZkBBmO38Io+uJtzquItPgdDSpplrTFT9pBDRnc
tC7kEo952UHNW7FlwXm9Ph8anT+B42boJo2wAjoit3CHR3f9e+IoU7N4vD+c5kNNdorXkQSvRArn
k/hi/zw9Fb200CoDYsrMe72eDXZFM28fS9cLNEartGbTfl3+kC0EX40PsGh0+4C1180ZIdgTR6WQ
LEL0yjb0O0JTuQKegv0dTrEzlmTIN7Mc43xZXHyfuXeWWYSEuftUUylbHUKdSQpKNBcZISChT8o3
btd5krUpguzu2h8Vy4rCoKhoZxHgM2NBZkUkyrCVLLoWA7Eva4F+1Ic7LlX5YIgS3HqzYUJloR8V
saGL7JWprwaqA7Eu0A5iSboqcTkPO4GlkqaPnKSG3vo6g0Eu6urm4cd7bnQ2EjWdYtEWfKBgYzUi
nbTfVL3AsJHqhsE537klmtxVNELVOzcGzpr1pha1rxzKlRx4/hUg/LEG/OONrpjR+uGj9LrpCePG
n6lqOhZed6Sgva3W40OYYmw6T1qsEVjJKtxuCA7Q8VN9HGK3uo8gOTmq6imzMlIQB9ILK4p/Y9Yc
dQh7M2flygB16ZHkLX32o3kJwJlyweox+RAZlWKTajJg+WK43J44WSlUEtWwzAJgmR1BqgYOZyeR
AGDKAY7GUoe+/IatdrqV1DGIjIhqByjytOCOgXIgBDCe9N2laGCv6+iRNLnXhc3jwsQdX+RI/XDp
er9IMid7pg8X9560sHMYmMi5ZZsHaRnnqtoxF+KEv2cB328kIGTuWtJwgOGGbhhVEmJg6kpkefya
vM83iGZ2usGG4ubxlVhWkFudTeg/3rPCM+/ubSTOU0y0UY9vBj+AhqyOSYmFAnaMKAvbUCW/N2hz
LiiFYXmLF/d8n+W4grbkl4bY76WVfeCqEVydvPF5DdcdXf9Wkp8hHpcaGAOxfbQIcBkA7vI45epv
12cxJj08MVoVCEm1m2SEwqaY5d089NRWoBDkXzdEGpCA3WozWYH0uKf55cmju/iBkHqfgcEp+OH/
DdykG+0i7LaiYyi60rOBeluOZ5rbb3LeyozIVGcc/hplBULySlH21whtH5/mTf6qjqzOXhJMwb7m
VBaw0clFoJjM5XGRZGt4nwx/F0rcfsdITP8MU8ILSOYjC3NAn8CgOsUdMKYeZimiaETmkRPdBKk+
ofVCM/H+FXKip5+DSU5UVbEtl8EY85jQQg1dGYpWnu1GsM8UqJURsXguIkZ4HsWkBF4ETs2ZM4BD
ft7cg2pj9PgnVZi6OnsOSWTWTzEaMfiLo0WjMa7bafybHH/zHPj6mKA9d9NWNY0x4GsIiDknpfJn
vFWTyHaJ5ucaX6fNmOZYdoeRMxygjnNOjAtp3LP6VzOqud5OThuVQcVReyJLuV3rnK6zOGhEfflG
92YughpqLEq4nMklH3SozTCdNlx798Q4XJur4uiWho+WOeSL3XSb4bpGevjRgZQ+2cBev+I9loub
iV9CbEo3QQyYtvT37juYxPOvKxLvwRHRHrrpOBqAu24cdkQM2y3SWYxcyyK8n4Ao2+rt7MzS2JIX
oQ3iQw/fCuGVKOpJ8k7hsyNzwIBdEEdNNixfGEq0Z8XvciB+S6X+CWko7n6rKblwjuS9XG1PGitp
OAskOzYCF7iS+hypcQeN2y9c2VyKA4Gg8VSzpUSoniAPM+D2czwzLcXH5k+0eMFgvWlR/ICr4E1E
OEgLA8zoy8knDlCDCfAtDu+aNItOz9nPnjcbI2/9/120/4ClgAa8+fuoRRxhuK//8yFPFD+m+UJe
CtM7icWL+pXMuU5jLugZjXJLhrS3H4JuQ68Ym8YgzThXm9mvdwn7EWR+cHuyXO0PL94CPhhhfXMK
fH7PjRIuEfaDn8sNpY8Jm/rOWpZW3mjGQyx6CRcLOBzREAo+GnRR1oQR9KP12059GmgZLbz0uBSw
yKYBlOmUcKPwppx1/jXqSVmpjD1zQWdcJ1MfGfk68LCYAqZj/0DYF9Y++sspiL2dJYKoPLv8x+mr
CBCTxq22DBUytWm2hWcK3jj6p00g5r1U7FvQLklVMaGmr+MR10dN/LzqhcCvhbw8VWdUN+ZuMGjo
HRtF5TgMjYddKE3FnuuTVMxp0vQg+Vrv88XiinYnVubpsxJXjz4NFOPPOpuYfahdOejRcViK4OkQ
V8LW7pnNhBDvVpfaMRy1OeYzCu6TQYqy3yE0aLj06Iz8s5DM8gy2LMEAoQeO8nKkEE50rSIAgNhl
d5Jt4tp0fugUN2aIJXxGcZR0RghfX3dyItdfEoZeFrfNqyId2HRDw615kbnQ8+8HXPf0iQWqxi0u
BiM9z6V7iX+7ZXOYyVA2zzdY+oNlJWuqvGSA3mwVoQIIeAJ0rejIhsw2cgMwGGErVGv6wrtNp7om
vCXzZu5HURKimxnrYIKLmT3Ms/TG5O8kbujNpterUdBAwD73EB0WNDdA/WL0+wFWeG/otvyr0or0
vFq5awuFHrc+k0PsyqCFUasuJNgdqxkhwEPAWGfVrkP8c9mr+94gg58evrrBUtG5o28ARq2pmGJ9
Nnw0o/fb06U14XNnDnTkiQkGKpiFLDHZ5IC40Ug4BcVIFGgMwtvT/WfAQGcq/DfSzLUgRSZV3h4k
rdawn48Mn+2LlkQTwSFJ83s+DM6jClfsUPUYQ3jno4eEMCM+H30JWVYRy3qn3sOxIAR0D8ExwwmS
9C6m73izKid3Q8PJ+DePaF8VVXo3LXEKU1zcgcIOZsz4bogu9YFsPp+O65PnKwPYqwhhJlMjLF/k
YcT/+6rKdAS/Hjs5obQALOKYCDSlkSK/pK+vMdGNF8Q61AJ+san9c2mkT2irRuZPy06jJBqH3fLM
349/wWyrr3ClLwkLC/AzC413giw1hQN6i0ljfxRQhnHa6CickHFR3pbElxUOllMY800Lce4o7FdT
GQh+/575Cu3TEh8o++o7GnMxKx8hZXS6rYgl9QD1pcsR5xO3Z7D1SK0oWQNSG945z0qkqRdN6k4v
AoZZeFMwtgvCFgi8D11YPMWx/R4uJMQiQF+pL+xZWWNVsqdJ3lUBkLJ/hbcgtPWJsvnpYxjTCo82
Vmo4izmVu8Bq12hsTqdd3OVgM8sKeKGqusGISThVOdIt3cQYsFKoakLuHmgFwcbG+SzEOZ2Gmdg1
0HR2dg8OZ1kv6Te6M3cZeLfiLOciiXeD31YfL4l8zOAtKQVhsiIoBga4gPphjdbu+NPCUyGL1HZJ
YTQ0mvnzhghfaVcW6AkC4RWA8EgXuWyASA/Y2ACGYjdpun9Zc2Rm9UZCxpDph+6P1sxQDZNChqX1
cP/urZbzyYXjLMaeAVhAp8o8mci1gqphV9VLG/5H7qqOVZmEOsY2h/xTva6kluDhJOMW+qvSYYYJ
akt+fQaN6yMcZbwm265kGpKqLxdNhaOUm64GKihOnuSsvSK8+HPOOylEk7nKlrL+UWOs/iZ5Ffue
DNUR1UfCrqpTHt53YX+WqagiMNQ9UFvMy6TDErYFrRZ3U0qeFGMhWYaDlaeW6kyy6pZdnMGWCund
I2Et/uRkL65rSFxgaU8ZvAAxXgqehnPwMshRzbj9VAqChJDEvPTPSD55HF3cFOa5ta98BhEPlahr
v33BnDXSkEZQaDF8Md4q7Ya/RC6NYL1ayXSUUjlvfUCTQQ2RaQJ9nVhCo1smjVt21eKw14jDKNRh
wXoMt5Ki//E+VO4o2U0xL+R+oL4eXPTQp/SGPP7zR0O8vwvVkfB8dUG1382NmxFuNOITePRlCLzV
VinaB6ANfh8ygOCEuK5bdTMXG9G3zRW68IqSR4tQl/8iVjPVo9d8rterFgvrw3oHkQEAjlxSBsTr
ZXC/umQZxYVMsgzuBcss4/MmgoCXAbkkTa6HLuAJVitCeQAK/wvyAf433BWIVpOTzKRh61ehfu2P
tyatIIUuTS/ii5Sier73G+AIhL2vcKonfyiejlsAKLNxkTA4fDds+8vx3V8WoVRVqDVEJfYe1Dbp
ZaUL4kPjy17Cz/LUYmos+lDPpQ0Dx9IjYDbv++5mSbgdnbUP+rymk24CTkL5uTJHe2pZxk4G//77
l7Elos69Vcy1USi289PDqxvhx1RVMpuT5xhTq079mpNbyOd2haBrfBPjtlOTtN4eNaaiOLkVcDcM
NmaSw5a+FHJUd+YXfgKvQofzjZ8CGCdMTiqeajRaLEX+YF37bk2201PE487xAMgT2sckd28tHkVk
UCjVoPWQ5gMw1xENRczFSU5FNE7orf7tvJ2AjlUkIP6bPvYQxMwM3Mv9L/ojPO860ILQ0hRr8D1v
FZi4DivNjuphAG0hoqG4A4Tn1Fgb4NSFej304mZQ11Lkm62ykr45ROi+S4JHuhLgF2qPDFBuUXVX
8Kma/sP6xoQWP3+xi9Q/UWQAEvHy6AW/XG7tFgix8YJaalyvBNb1Htd49+zW+3Z7yNuE0XJy7I66
DcaqMlePt4Zke4rhH5eppheL3xOOg9SkVMmfHvvW8OggTzJSRHYdUnlIUpDChO6vljJSxgK1u43j
V03FMTjeYjRp7OL5+LyP0YVukCjPX1+IVkUh3C+mhlY77OFss7iuwP4WicmSV6ooztOLuIW8YOar
NIvTfCRO86UrjNA/vPlLefOh1zLo2bwR7VkZvAAhsCs5tMJHPmGH0rUaBHTb0DJVJCuIgrz9fEll
DvwJPW23A/ZLTbmlyCf1no2LmsW2YpJhVIlZAYX7N76DAUrOd+BZJRKKETN2WQ5Jh1xYClXcbrg9
UF54VG82/T1YNU1Y6Exq9dC63Khd3mFeSrEa2wrtRX5Ql2zPH7iK3j090IDXHOEBPdyUtNXrLc57
L4o6Ztbkr6RwTjY+QdGOf97mZKjKj7jMSnQmqsDIRC+fWJY+oh2IcCFp065d3oOsNyY7x82hwWye
BVWJqd1iaEDUmu2PBCzEIzxOoOWbhpC70dCOnkU7SxW1rWqf1fPbaArSbmMbxCSppC2NL3drBWDk
vRFPTtdASSREEUnO+gvCgOBz95/j2T3ZY6ms5AoRBytO884FbrcQL5zXsPXaIJIkJbqz+M1iP+3f
RU5X/jIX1+ghUY+bOsxxJMRZxlktoGwlP4e8Symo6Bs24J4NW6COiaKaAL6CAf+wElxDxwswsshC
AqNR/qDV8ZJmyQyiHdEh+v0WXzu1f4xpp0A0vz5as23n68WTxgAVI3ZMnN+fidK9rivL4AkucLQR
ATALlZjOay8d9Pmw8RBhZp1fu1d7+Fq5IO8eDRBPXzo8S1pBsjLQiQhnZxlEVRKjayxLzqVxdCDS
ict5S0PB+8QfLy/VwEN1+GNqMzGb8fZVzccEgrel9Rvb1e32AsCzBggwYp2CVZEvwCMF1i9eLIVc
WO88Izc2fZIgn7k6DqksI+nzee1RGvIKHIQCUtYvFFFP5t/dbjJ3sbCgNOE3WKvBZ1k5z7J1KGmH
8mfx+jgJWvYf0Nq4I7NX6PtV1+RnJ54F15MvveHfj0Jz+JK++eaBp7kJWrrhMy3OPrOGrGo4NTrM
JyVqNyaqsZMYh8Vd07nTeDzld4ktb4lzNXbpOy58jTbA1c08tPu+0iAX1mmWyMwHoqI8H+lioDOA
63JC3tJZ8WcZa5K+lviZI0SX4sAUe8Ev43wkH7oXJzLceMw65NXO7FUTDHSvonHPre3sdd4s0/+Z
304rZe3qLtOZSSpM3WX03csm5tv0fRMkQXUZJCKX7CsbB5eXzrJwwAwq6PGczoJmm09v6ff1C0xR
SJDp6R9wd/97ekMvCdET/6pBPZ2yNd5VJR68NHHcBp0lr0HcvMBR15pt4AtN01hUm28kUmiFOA1w
PxMkGkr0H7IYpjZucjF/hGRSywH4Ko4dtt4BTuURvkjFLR8EGlKezNkd6m/Yu04ciAgLX+wMSNUV
wXaPIlY6if6c7CMAThgR5HMYm9I7jwIE0qqfHu+/PEjt5F55St+mEJRNROhnq2dxxMc+7MXGVVYE
T01Dy9NARGfGJNfyUr/vUhs252t5el6sk8WapurNUM+GeD4FNLA64usBejGoA3W2Hir8vK84jvKH
CzH+CIgqSWD8ivHtcb2Yzu1eB0ueu2VAFELPNlpBaCRNlR6DdETKyoPbq2WSDlJBM757ZgTN1zTG
Pe29jIYkoyX4iXAJqNc1ccDl5nynJ91blZGQgHk5hg0pPSlCXOjX5GyojrGuXoUlXl75bV2KGNYd
H6YSTZbqmTzWbpg7M5GxFkXWFk/zphjNC3DsyD7k50eYspT4Er9tXhe3P9KonNab6XxxaILjDP0G
5Icwk75bb/hVcLJOwNoTTBoNpVShTcUtAbF6nb8NbD5DioyZW5wW9Tv/+zRd4aEbThUp9fJpsQhu
nStQEcHwa4u51n0CPHDU6mGksZv5NpoA88OyYruLPhjNdmuL5GISCydusx0ctiTrk8/WysLMAyLc
cYu7YIHm5pAADr2yUqTVXUsSvX2niLKVwo+ZiyQsip1xHo4D695H9/hRxl3aXHSDFdR20GjrhaN1
RURbsZoTkfq9D8KjvYAkdUMQlO3xsAyZDRMlqcHhtwm5SyvBPNpWNCl4wihmRFAasPv0GFcVjDBq
3vDN/oswT2BngC+RTFpSoLwv88FZPe9g8KthHZ3IEgrTJ/RHVBDMs5aj34ai3/BbPhbUum+hyPnf
tOIJoxBu5SF/Em7YFVzloFCW9He4kdSClSKih4q5P3jaGzecnA9jf1PK75KKJLoWPn7GDxh6wuIW
EljW3KUeI1RA3KfAr58JJxzZvbwpSnRovVRKnB28PwMffWleRv6GIxur+c4IKtJdOPSHk/aW6m98
fUEbUOAzY6bpsq7r2RHC1uTHoF+6QTbDk7o8rGAP2yHZUIbKo3Drae9gmU6RLfYQWFPtFW+Pla3v
5v4vs2jYRjCtDertvFK89tNYh9kkQtzIcWTIDdlCL1xHC/Cs7VLqpwI2FK66H+QKx1d23reD4q5/
yfY+dgLjP/gJGIkIp2XvIhPv5rbcBEZveclZTrSE6Nd3WQpMxYFW00qO6qEI63gl6wCJBdkQesWj
KcSRCwwzLpm0Ey9iNYPZISVSHHnn5OQivXiHaOWB6sMk1qK5pgWNmsEhwKy8UIIv48cXKqoR9VjR
J+wjs+QkIhmZZKuIGq9xI1EZkAC8Zl1SpIPEOpZpzwpl59A3USo5IZi8ctjA4AUELHW8w1luEBXg
QY1CO9zMrcEI5pr+X2qp6HVwYOKU1FuTdkI65lAHTPIBdzYebL3vEHi9BtEqMsRoLp2XWGvVlvnt
hoqEkY5g9ltO0KXJLgN0PJexg9JVhweFJETzsQzZD+nYXNDNojAxmTIDPLkeJg/JiWvgiw7lJnjE
yHxxKbKMqtrLq6afZN9xt5+Iz3n3zxl2u+4e86YdXFPqGSv/g9lxKYD1dEw1nCRTBO89F1wDSjYK
Jx/9/6IGnTdC+43ZmwQHRDkiOqnEjb99Jbsc+i1BuTBOWHnr4y5JBkmjlHGbwTS+6hiVGZrqTxLK
jcet8SeNd9ojUzeXaLKiMAYiHsNFMI1N4Mo2bykyuFby3GxLRH5uoTuAP5DCrPQOHYteJDN4WOKD
0+YBXsADuEXF/AqhWYecWD5l2Mc/LaTbeyubrdaIqG9QD0nniuSG/wXiLHZe5GndkPHB/ko+Bh7Y
MnheX83aKkzirtFxp7Rn2aV/Dgby7XhjIUvDMzCNlXG/Q5XYjFYCtzOBgbtlLNVSBoBn4K5EgvMj
/aQBi8x5Rt75yRgCLMBg9Zx5s6obn9MqipRDN+CJkTKTeQ+6SY+ADMttvr0rLesFEpiZlFG7aVui
EhoK6sA5vcq/dFcbB3hm41usxmQ4/zof4fZ05gIq+rRzAZlaD2tUUlh4SJips7AHrRMHK36b19Rg
SSvKfm/4VjkwgCWFpsT+dB8A452bF5XwfHQzvlaeuUqkIiLvZ9EHX/VzZYG99Rnt07BQBmxH8aPQ
NyFTBdIKWFBcevPKQTRlFWRQF9x797khTgEKHbrfoX2KMSPbE3Ohqq+o9SIa0HnJW2PNprX0LIku
BQvUIjU59rFeBWjPL0Y9JCjpf5blsI7HH81W/h0mhtWC7FTh+t3Rtz6zlAzL5WGAu6K52GFxO+Nn
0g2xoPKApkx4Txm1DkIhchDi1cM8ABeay/B+a8ndE7zo6kr0aeiQ5KqxA2tRw0MZlmbT/JwHS1bs
FB6bBFmVMEyOyjWQA3sKYCNnDAPWXMsX25h1hMr6l+0uRhDi9X5zw/AzI0HZ7mo8hJb2rhY0/6Oq
OhTF1HM+K77qTN8ZusEdaMjl1axcPsUciURlU3CXfUh4Pp8vT+R7b3RT1uvARbf+bLigXCkSb5p/
0gLEclWS2jPhSp+jLKFDohZRjMEl/iF3Zt9LKxwHlfFc6bKrBd/L4TobWuDgXG9dkU4FtpKcUyX7
3kqtVOboolBt3JCHquVZFi7JhBvJvDsUV/7k4scZKVWuDXDx28gXct6lY7c6x3XUXuxH+pbNg4eo
AfTf215X1ljYvuv2IJVDKTwuAmsSIRScH+v30KaX/vELAcLSCRG6/EgAgU2yZb646aiV6osSWkCf
7f/gJrtoqYhWYJETjT3ZCF99IOY32xpN+bMESdZO+EJQxuSU6Mp+WbAJXjVk15mbkTuJVxVZe8E5
OpqSTqOg+/bDJQpn3Tjwkhlqndj7narwZI7FdFuR1WHaHAcXpGZYDtM7YvnwpRU7LvuMhT7SkEW2
Ic4fzUbWuVHaV2Pz0exdr+gnn3ZyvXNO7VCpXKooUEajtVYqXlrFu6BbQo3/y1XXPYfVkjhUh9Nq
TeCT+q26p5kNyBcHfOmR/zMwprZsR4ae4MSShxGEUYI+qvgWdGUHUIsfOPC7tgUC1vAPaQToNamQ
Paxllb8hM34SrT9FdlfxC6C+yCkzctNu7R0xBCupQMOCM+823E6dlSdPdsc4L4gB7MwfTJpRZ4UT
c5zwaD6lCvkcQ6CYE7NpGXgxPzqNnPOa5xNzmF9E59TDkLf3+edkLXWtQvhNKBwN5BJHRyV8c1DN
mnDQD2lZm6kbSQ6zSGG7iOFmaxiY1SZYvHa/M6PcQbTAkSzDDodqY4VX3w7KM2+cpmfN/ZJnJwZH
ZmQpODFp9aAgrO/czGOvcJM9A9FmejknKJI8UmNd6i+g1zaRpZKDpJVlGZoDjXtrdIKV9CdaNU02
I6lRyr/HQERKrmJJ8bi2edzCquStGoaIXKaGcI20EjZfsy7qdC+zMof5y259hFZ3dhk/2UeBvt66
qUqpfT+QWTqgmJ/M0PIvND2Nhe37dYrDVZCuLGZUkjJVlelThrzsw3+Dmj3udAsi3fURm/0vEPjk
JPMN7MybWl1FuYp0lcqAdUsFmnJEGg4NrGdqlHQa0HGZFHlfWu+nToKfpOO6x/1i87zW3tFn1kOb
ulzOGmWQBBmdNNXjY54m/jo4J/VIJr/lvkD5mGj7URZMzPshjDfOX6a7poHXvaPrEKttbsd3QJfD
DE4tAeRk1e2y55zGKo4JNxBBnVBIwMwSH94TSAgf6/zt1p9d7o7Oy+43QdvDnFuqjH5CZRvs4pc2
k6JGeKbqVGlk09kUqPjHz24WCQlGSdZG5IhqJls/fwIBJJSuwUx+2uo6yARHjugigTlRc4O7E6D0
lxM2ZP9lWF8+dsQCvo4Q9Ij+AJp+QJiwPmETfx7Rvpt7zp07a5dUfwzSjyFGQjp2Je7uFPqOVW3w
/09EW7eeX6qjvXnzDPHngrgnx/oyzdBo56AGsRmKdd+K5AOIv/VCvSFLHo24omWri7hfUjTlwDMV
r8ptuw8Wj5OGdEJYDTaInblvFj89zdCU3lwPCMsf5PJEVK9WlocJglegYWwcz8OOcDrtudCWisiB
bgOwh1BdEZV6ln1PC/ZB/3mFGkR1NPgrNDoXu99SSEz1VCu/wJo5OjflDXvKM8C2cVUoisriprno
2DPN1V7RFKwIA8gA1kmCgZCxJEG47PDygqt57ET/IGl5JhCb1wk4G7TKTGaZza16ylF1GbCx1sa7
QXTwTNobYAPjEPX7VEMS9iYD7N+N1Ete6qUlmiixJ0fG2WZ+L5KKgvNaw/s+/vBYArBQgX27KQW6
UhvZpaerFjA+LLRZn/uhR8iHOYLrH1Z5dLpV2ZllLsEw392EYBHRh9yi1VZbmV8p1GDZdWoOFo5t
qkedNYrVd50isbaj/M+GMsy6DbG03HZRVW5O8ZWaFsYR6cr37H5oFrebYp6R1zyCVhpbNJDZ+2FA
p/BitMfGPouQQFjqxTvoN3yne36v2sb4irjFzhS09H+tgh4l/SKRI9LOi5K1JhadST2VCwFb+L5v
y6fgJcAF+Lh87JnGWX2c7p+2+/gjOlzZGG22HwvJkyTwBLmdkTCMBFgyM4lRSupX84wxfyJ74Ahv
OSx1T/kA3VNyJ9jtx9/5JN6I4R/B4xRN/I+3F+Xu+Wc7uAw6O4KuKPq/XvYNwww+Nl7lF06gh35y
N2sTs9T3Rmy2pV2OwtLPxrpGmhKiVFFfOhaWVxC9SMoP3u44lReBLX+CZzS7cD4FF08Uc3KMoV3Z
BJ6xBSw7N/mLhpNNahRnQLO3/OP1oTUNKd0gbaELC0d4LcBaWi+KHfDum1ringUepR44+oRDo5kx
inBHNnbts698BHIwfxnqnQTyNgXS/nn8c93Yr8ZDPuUsKPSABBIhSo2z3dDO5E7whBK1zPQ+2lLu
c8XR3sIIJp8d4CIfCUnmtXjVdPmWxKFgJgKozCyOE13Yl9rdxkGRulJp6996Op/9oRWkBs0bxn0V
7cGgAZEtJlLiBhdqlX+lQEqU4csyS7i2DLoTPWZArYXt1NRHzsJ8JTYFDuMKiIXGfp+7MwtcPztf
7yyjZ8wb9Cx0T2Mzo5lyllkkJWLPHzWKJQ+5K8ixX8SKBsZ99cdHxDPaiFrD78f6v24dsWYa42RQ
7Wu67NjeqEKaNZZ2kQlGQI78TLjUeQ2xT3iPeY3+E0aTXqrBl81aaCIv27Ef/fqUW1b9cXSh/4Co
wckKRiInTANSUn/Db8Z9A43QAg0SxQHSPkJ/d413/gHAbFoc15Tep285zWc3rb736niM4Tqsycdo
6qn+K2ldjRwe4nLdYwoA+GA+J+U9FCcMR9EBbPXL5zKxBxRR8dNWHSOVkiafnXgy3r4+9ZbZt9/L
TSa4nsdKLDBx+Sg/5bK+SYhUb0mhWUlmyyVpTOTLbZZVzH2UqDbR8vlzbNnb2ELQbDT0SRXnWQBH
U1uoySdsCRYRFyHOe9YG5kSV2X5+oQKvvGieHc3Kwd+6nPUIXD5A1WwkChzeHaIiLzwpeCMROdcL
skApLdj0aS8UAsP6GMcMUHCuVSXD+35R4/5uTwOsGmBOaW1ZN05nHWjpVHH4bJeILDgcl3/XJgLu
pt4vTjP+MtohEX6XQAzKHUa7r/7sxWo+lBBoZOU/Je9gGJSJjrtVbtfpPo16klT+qe8JXYBP78+m
r3DLDAprFe5K3g317I3xdgZpiHkAvsEnbl1eto+p1+HYjsZhXDf3Pkb+XgBJHqH2ImYrJL4d3cz3
2YmJYodsY4fW6MfN3oxn5I0Xu6bsKx5kAi205fCusnSKjZE0rMWpqgEf+qSzssSNbIqvSCQ5uZ/T
GB0UwZf7xU+A5fqNAtsIvnJVYcw2JGAvJb0PQ7ouVdOG5S5XjnVYvM7kYLkbk5UhJyLtLPQhR4dQ
cftFnlefHbKH2A0Ec2wD4UiHgq8q0sJBqb4kyI4EJGogx89lKFYhIfnF/Pyx6CAPvwRHYPFAz9dP
3k5A3hKCj1At8sRuRE5KM7Z3PSqG4Lx3Ipxu5zfcIxfj/lfeYmnShOW34Grnt6OW7jQS3qvD9ySj
2cglD+Q2S4ycMD7K8MQu3gaBgyARxYARoz01/UPZ5OqcTBYuczF05NBTTYt5DJOAk/irWWmkiZHq
SCbsa0+qKgr/tKXk2EWRjf15onkzUUZrsTCLBeJCYEnF5b5hcM7KfhTjENCplxfq6jNnJGH7v39r
TlUQBV7YXYpOhgtgaH7fwAPQ9iBBk+afVKM6Y6+mDS+WIexV9VN0kNDBFfdebDCxkNi0atIwqdOM
piB2GvmUv4qQJx1cphkXNmPDDj/+Hec5LcGRvFtVPh7IES03dGVoU23c0Ua24xo2Xs5DS6riMaX7
nqPe1c04kcA0EwEoI2xUadf2UTpeOm3kmkQR6WeXVgSGQlZyro6jAEZL/mfqArv2W19Pxf/z4reB
wOr+2k896ubzbFpuboEhKxf/4/fGmxdov4GaDuEfy0IFPvM+R4NfiNJljiSZ4CFVZNpQcmI47YER
tlnG/+5JOAla3r1uK0FGEVZ+Q9A98KarRgUlLxRvQ+TJjyd1CJdYfJ9WG4fpIiH+p95KOYoXD5Ix
vhJdyItIYrVb8AMrGr2dkic2UeFpYyOq7laZU5nlG37SNbJBAKqckNkOCoSlZXl/mOhd8oBnB2t0
uZxOwGzk35eZXmgOmVpbwJOMsQYN82TNFiVyEQzaGSlD/O8VDjbK7DK8LvLWqVDH8HV1oYo3htDX
DyWXpxTYeNnY314+yZGzaL4QxQ6+eWhrptHZPUNGOQS1v+qFYQwKiNxZYEV8nw4le6uRTAmwJsT4
4Jn219cIiBjXhvguk3HSxZzVofTjZIXG4zY5wScLjz55wPZHrm5Y78pWAVA1hKd4EE4DfMKbqav8
ApvUriPOS3yDIZ9+CXTLHEOR+STZM9wDiLfex+FGCAs7vfqVnQgNhtcChLCqo1uNuV8eWbnfKi2m
7VSQMQiQxk2laqdHZfmNtQnM3KT6/6QvEJoFcV005i7pFnA2CYdkh1Sj3HdURwTb8ICPHiLRahYX
9faTjjbBpI4xa7M0qWwm0W1/fFYQ1TejiQzUqxCOyHPnPOG/yG4iHshRK/Qd0sm0N//c452yv2kc
wGAYPeVYoIJgW+V7oWQK6MzxefppShcWKl/NiBb/eGZBQAQlhYEABlGGu7Kmot1R/+9TLLJ9bfD4
LLp6iKhkb99OAtAuZ5OQdsK/119/njheGXsIfrL1PYTXTZ31dnty6h0yg9HnRXjsj3/DLeXqIB8t
mzg9Sc7EgElR1jpzEqnEsijZWGNmg0FnsMhku6CuM+cN96qfPh2Zw06hvXgULxpQLVEeeAz8uXZY
tZ6Be6OXJsnf5SrjpGoG6eJGDib47AWrecY06/riMEUc5FpjW3LLrJiPIaO8/qN0eySeX4kiLcf4
iIu9F8xqeqSKDUDjilT9EWnK1lGeI23mzSIz1Z4H4UOQmgp0o8CGhqPgng1/HwH/NeL3ZSgma6W+
wal6l/06b8rUJkjGw0IvcObPk2AdEOZaBMcBAnxKHyxx7Kt7BWksCQIxZdUIvEwZWXXc+hXN+Myo
JwMQcEvLk1UmucVhKiRnFU4KNjjygOLumTptVeUUT6LNH4APEMY2Etb3fQvo3rDGIwqr0se7+SED
4kJ5SMvOEiEjo2kywQhpAAfz7Tz/b4CIA7SoLd1UcDufu2x7KFffnoQ2IUBZuFpToYfB1FcSFRgp
58qPypGKzE2QE8xG/DqXphhOQ8Fxm3jeapWXx01D0uvZiIRI7pXnNir1v/g5L5YjK/dbieDAN5b+
u+M0VeupLD+Z1Bu1Q1XhusGBoECL8lcrsxvJbh/Pbz+skxAw26/jKXE8xjfAay0Xv2n9+AxWM7pC
OigURfRtlNUs3lKF4mrMGtHVriLA9iOFK039cvT6N9g1eQ2UYu1yMR6PBGc9lPWJo+X3CJG17Dfd
swHL8GZ5ljTITEAcTWH7W6h78wSM/6OTfI62yBlWAHXwhm/4QMsz0oh2apLYlr1hjWI3+00ydQI1
H/d4swMDdL1DflG23QnDtpj/AKDAtZN5ryCjV/ZWouNiBCvCv5c0ESXfC07aVIMmini2NjFzy7H/
A2E9RAjuJhEt/ungorbNLl2MKUDQtbSzbRNGs826MP7u5Dbz5xe4DGsKs1k1CvukPQSDN/pEWfAr
J+S0Z7BW2/tLCXXYoIneIZ9Svx41PhyICxlzjqUiinHamznbt4UduwB+/T9mEbmSJFyy1dZ2fK2S
hS2FgooZl2eEeNbAba9Kjfk1KfCNt0Djq67jfyNpe8LYoSEpfoLVB/E3s35PqiqlyshlWrHHC9Pm
yQbpW5RS57ZWW/n3Wy7okMTXnguPk1mPTrWtpESGyFHwg2TjYVVno955phrm8XDjB4mzjb998XSE
stxWQNHrwpaAkjaInQQ41+ftDKm8/CWNatmWns4sga6zbnxkT+d7t2+RruMmObXSZ726TyTxn5wB
XlxJFEK+s/sxZMYuhrQCqQeLrG51jp1dTvi9efGH+lN+uwmOHGEcoY5XjiZo2cdT/Cvl6ZzlHvCk
iwGmO0dGX/mBx1Kr3o/W8JktQJlaO+DdaJ16r+hDt1UGpMvVoHUMdwRECNMjsfFq5LwTb3lu8UDi
zO1Dd3Sd4YSfYqRACotjA2hqc04o/PvQ2ttPtyc4N1rp++G0nVrB7ToUpOyn03u5LCyZMKxseVS+
55Ik9tOb0pUfBUMLU/DxEle7ISVhlPrCF2T+bEByvIEUMVxHgc46fBjSYy+csLFD0oY7CAamC10v
BvV3XKn7hmC+L+S3bt7+74B4pBXxxk8cGn51VFAmixQpDhJ5HkX7RspPKm18PRT5Yqs3FgweThLV
Hr37Tr+zTcdxXzr+Nz2saI2NP3nDd1u2rxdUEijhOrD9EXa3/mcYFAlrTpDSuprEm2lrdJOdpBWC
mfUeO5ROXHsjmdV0dV+9ud2QF8JIc71DZiKV5sMMkz9xWSn1ytk9YcXe2wGOgslB0wJ08fQs9cly
1oeuK1Wj0vQXF2IVNMzfhGgTs1IIctX2DxUSorfQVTloKaQimRaO+lEQYIi+xCHXzvrPjigPGbfU
WXyJ5m5TtzGfnZRp5AX5QZOvdUI/k736ArDCPc6kvMvHBiSCGWD9z/6ZE18dt2Tksj/Gahb8Fsmy
v2WDRQ6J3qpjkyKmDkfIqVPPph+1TPcAIKZOLA9QzySIpGV90cwYi8d5lwNof5LG+7bVDfa4+78z
gJ+F5xPyuXh/mZaF7ME5gELuqv8aNf4ImkewgGOHTseihWlouU/XgGJb23UO0oDK2dJhMnTUtgbO
nCDQvJXWIgVumMO9eDHh3j81Cc96BB/i2SmLxUIatRM8K5qvQTIy5wy923If4YQV3rI+3qGOud94
J0dULcj6PvFYgcNoBOR9YekVyh+wiQF/Vz2Tsj/WyXxAR/j+Qj0FuWbL8cYaue6Czpy/LH6+7p9E
qgxqssvX00VlEH0QqXMiAnYct/SwMFZVT0UOYa5XZMdg1nqscyUNvQYCwrVOhPJ1ll1W3d9qCClu
7aDLxZJJqvLbQK+nMr0YXaBZf0OycDzaVwB4E4iezYP7AZ3KBG5gY9D2k4HD8qqhOdUWPAQJjoog
9UpMaUl3gT668Lg7siAZ+a63Ykdk555nXPnrgOU8hH33crhSsJVe+MFNyACOOkhQwYZ5eYDW5rIV
jj5DEihlotKn9UREmcc7c7fjRmVDX0UtmRN+D99trbcc/LPU4D31G7hVqDawsnAVULUn1OFaVUxf
yiCmeM4W2CfU7rozlvPROQXkwVCsRCEYJzgbwWmPdvc+uFmI0w+NKltAy9vGgJlbpkWZVVvHn2PM
Z3zFls/353SAf6cujshjnPP0Z3SIL7tXSE1AaQEMGn14QAcyfC5kmTN+KnN9OeK5SnjrtLrE8/xt
pRLSB1zhPBpT0bAmlDFiJB1J7J8+0QHeuDE3teRWjFIwY3xggDKKy5Wp86GvL5VAW5QSBP/hCKXC
fqZrK47k9vggyRv1zBvRMUp8zYuNYVFJ+/xp0FiERLaebhv/28z6hJ11c9px7GxFQT8NFPAP3X/V
vN79Anf85Lfw1yTS3+fNwxwbGxNFgObMmWRRbWgJxkuTPe0CcI4QVLvujk1kJiHo1jB8oDVNJiP/
9GlkgzfULLl+gFz+6YobAvJRoweX1es5DF1doj5BhAi8K2hNX5zjmS6Ke4v42SKQnbJkCM6Hxz+d
OHy6E3jtR1M742b0AMR9/GyBfUyKKLUpeehVVxE++vkT7yD+M2SzuYzycfVLacKiDyi28xelaQik
1+SMXq1K+b2IFwk8K9XYw5gXa1zgU+18JsWYQ3L5e5cqxKrUw2KSc59aA5SxeUzL6WldU9Bfgx6J
7LJHs49Vk/XQnrF4EcIA8hDcPIHfGEfMC+TiKLeN465uLxVtr1sfZJ76Ykw+FWVypUuOTsk06cI3
lpY9vXxsei16glb7kCXwQi/kY058+z2Wyg5mup2/9R7E0OoK4HewLMiWMOORFbiMWEhBmhwHqy7V
9+GZAEJLgcBxnAgcLmMlUbHzoS8ub09GkACGpRtrLDlFQJNLI6fAb2DzZv5tVK9rTt7k1y52SiqQ
uoVDY/k/JhA0DQsJxMMxmzx1z8s2Mh7tFkNW0jcp17yuvyGBz+T/xZJ5cZ3gQmZc/f9ExkqmVI/T
aoPNyhp24q4/fIYnLpQMY8Y8SBEOnzbqgcq6aJO9jrlYgLQ/TZemdIQeGogmgIgJEfx4F+rOytBe
e2arzQ/Q898jy9QOt2GYXPyrjLDXDx2/Hqc0j6x2diw7yCtGQn9lC8yMlCTkz+evWIjpX4BAaYlR
g7uI7Pb+R6G1iQGIhFuepRqS2MsPzOOq/9NUUeuvlaP5YzeuQ4i5Rk1UnGDyknPvIwyQzNGmMVTy
1QG4sGLdVjCAJAne/bazGuuBMcVsNHfcL7DcyUiVzZg3RwkyiJhGkfHP3LCOICvi06Kxc4RNW67p
AMvC/6v1SA2LZOBLQts+z2fuMPAfTCGyZ02WUitpMMUn6sxi1CMI7li5x2NvGv5liYxACQoIFeMp
YGfCOcBtXREiKbhTYGlOB2CkuaiFY5e+YZfB6/05Otr+VUKeILrPg81pDqN4TWOoO5eVzpn1OizM
dxyaZMtVhTs3gck0/mmAJLj3vbN242kFiKOj34HuiyHmfMDj4apP28ViZDGXL096wbwJ1MNB/lNA
jiqiRWJdBvzbEJ/xhpgZBEIbnhrRByCfF9M3fld7FWv5wrAGlX/ggEiAIkTb2yuY2gz/shDUHYOd
SK7OEfFnIlZ4xp+RhIqSp2fMNHRe6YrVF8JAHcEc3yo3arqC+thYivce9vMf42gnBYpKUwXFBAbO
pvEVqah76pvU3o6Pp/iWp4G9X/21+3H8XjvRUE+hA21hu4stzv0j6gEd95ze2d8T3E3QlsR9XDDa
ysTCo8Sya+1uNyjLvjJYIa8wnHF76Fl43jaadIpjOriBzlcJX0KE+YW+TK3vh4Y3HR1Q3yHg/Gyv
ALDC9oIsAFJrrj+B8UUr2PJqloOGvMbfPcAdaWkT+VdMF9/DUmaa9/bTlX3lQQzAbHvAGj9cMpVH
wNdwW2ctnhmBi8sw2t31PR7hZH9cGPDmktRr78cChX81qqtHeE44vWFXY7dFuvAwLLS/OrRWQ4sU
ivBbAv72PkNhijDqTvoNTW8XnC3ekNb3U6791mTqCLSY0OgBjzgehyR6iZ3NOaHRk4qKYtUPAtr6
KrtyBurh7dwIjcY2Yn2MukYYwR5oq1/u6WppW1huOfO2rzXE/hNhSWHkPmM0deABlGeQFvdh0K6j
sI/G0hHZ5/NY8dLl0M0ORkgatjvPkS8e76FV1Uh/1pgFjHS3pqh2Dywc2wJLnVdgC4rJS80pFyPR
ty9AKKrzbJl7XTpolXX4egrmTMDYpvfbkuCPg4DFGZ0qDE6stVX3x42YgfW5+veBmXoRqEF5ntMU
cIoT96qdbpdxvsoGJGDLxSasnmP8Hn/g6oqXnlZDrN5/ZbY1/E1DS5mcLqryjz3Ka7NGyXbfwZ84
CO5oBxMhx2XRakzyoZ5g8+uRMRORAEm37H/2B+LAg9ogQ95DEV5gkNufvR4yP24PktbnKyp4INif
td9bEGEpsHynThzTJBUcXkiOyQlhmYdf3ndNKu7CwmDcJl0yQoo/+lVFPds3iVD28/yVvM5UaI9q
eqJGN44d59MjonZmbFyID2aSHd6JHuldUN5diTcnMmDzAXKB+PWyh2Wz4VIngf/ZFrAfYzPs3RpM
sYPCiSZaMC12WahWcaNfGpO/ec5JvVp+juoizFx0q5UfBjJID8Rk9qMvjSooV291JIrFYS9DjN/C
oGP6/WDPoEb/ZeiYIAWnDt4cGNoFlKY5UKpnmwZ5lfQxdvOxYl9JkTs6FGbhb8jW/5qOobWXQ6AC
Fwb4Fx4Ny0LBMWBWv01sm30FA/Qbt8QXtFDCUp2liLTErCtqTbtvETocU3rgRVaFUIDLGDzBYvGU
pisPgVnrqDuMIew1Q1P/ENFo6hLqp51QpdHOqaNmNKXQyRJVgwiErskR4ZrrYp+WWU+QP610HhJj
wbQubY2uj8nM4MC8/6RD2bM6xY0lRGiy/w/dUcOuYvvo3ahjACchVyOYDKZAyc/qqijerEpzMdBn
UlL/bpXVgpBtf14So4BRACxN47Qac2ieNbsMl3sVasVzisq7ZrzEgXGXE6WNqAGAdC46/QwU/EF8
hFFSZZpw2ApAzExTWNYe/IG0npXNZncxdGFRsDPpNuDdbIPqeP4CCXU2l3D0TSxwyjN/eT8790JP
jYynZjEB9TJULobCiVI/IQT0+T0/eCBHnWI85LoLnpXPCalfbkyZnjktl0fdyw1qEPpF266SBJQh
xfyUISc17J9IWeFRk+I6UjHhnczwQZJS96jHEYW9lbS5mhl9HiUSCJ4plh9VuqGZUnAHNy4HHqAN
vy8+kaWtfIyYvtksladCY/bSmkByr0dN1GCK/eXP9a2sI5M3mieNTZMoX01+m5/SKvjypiLv8GG1
BZBuUT7+fR2VpuJSNhXbOO8t5R50Jo9FORrZhDz8O8+eKl21jabduMRpn01EUbqEcPPWMy3UtE7c
6I7co4gET0XTMGeKquJPlJxo6L8hMXFDsihoofHLchO3oGcAMy4EGFS2PbCR0tL5ednZJQJwDL9J
yl2lnKLO8r3bPkb/LWxml3xHPtrFUO1xGFdQMsD/wUlu5RjokCBNdOnEWyvQ90TAqvxuw5ju+zdz
lgLRIaENPov855Yqo0DQHm43jcrCh/su2UPTzKMzZG2Hp/JLAfecJKMhQe5chlkzzsmbaNVI7PSE
65jZP8IAC1Hkm4b0GeT7+0MGeJHSuc6KcOWkpwaS7CaIWLvI3xasNAVz+P7OnLd5pFennBH9sdN1
9exEb2ekfp2YrsZgU8HmjQnrl9+XOUk6hB6F7S5EjrULdy6NKErPxo6dRDXg+M9wDA0MBRPLTXbX
dReLDtBMKIHkYYTufLW+h/TVyHGgpEMfRVkMPjuo/L3qrUoD+skFZvixdHpf66+DV2u7kzJv7FAI
YrWHgEH+X8FFL2jdG9v5a6/CNbdKDnBThnbGlAVVtAB8Dc0SwcZco+5AQ6ZDJziy4UlrE0meKrK8
AqaMikCu0Bp8pmleCLp7M27lg7fgVaFtIi5V82u8d5Eu2ZnJycaLjv5T+yRJ0EMBj8WjHCsEU8Nz
+CamUMscG8PjLZHcvPIzJhkfi1cpiWq0lQY+dxx7a8iT9nUrgn336ZSq6rcfvuiZW5bMi8TiaEnj
zvb/zHOR54dBE+blIlx+r1F/zudpDxNnk+e8s0p6RHPIgVjWlbstNWPnd4eUHnxM7sg8zZQwAxcu
Lvqcekz/k4x8iDbUpT6v8xm1PJSvB/Fm5ehpiNwnmEorpWGwG5scD/Stqpdchkt8o0vDWRjC3TmC
cEI8StNA+pW+qzWw6NiuF7owR/VQY7aTfftfiJ0uB4xhX0kqlD6Nem4UjNhimMZ1DktFJqZ8qoim
LdChZrv2kJLl8B9TubgtFmQVtSx15jk/1PLqOVKECiiTzGHKdK2EjEHAs6SnnvFylQVcpclSWT3m
pWrwnpXNNQY3eiFGeOcrK71nz8MC9xAzX/ViGwElraSbuN8BOzchiOOJ3l+BEiBSeB3j68R8oRMS
0Mxyr2FEoxjjxV0od0Cfy602RjT2CNr7TMBQ40YZoNSv2g9IcBWH3EGJx5Z8SxJkPaSFJdTCGXzY
xAXYiNqeq++Ws6Kzc8n3pfUFoauNQEISnbPdRhb/NFAXVgwMPflDaT2NAQFKadGmlwV/55RojKS9
Wgxfotc292M48B7WeoFY+UjHkCwHXW2CB8y1bfmfHwE8pYxEDTSPHhtpup2VkNehVEwmrRAbQhnn
dLt/R8fEdSHIpVUmNOY0WXv15jbL9MpNXVz4WugQhPTM6QxGM4UyUcIzPYV52ZCDwT3NMaN1+oLm
8ky4CX3TXxg4a4KkgicI3Rb8MSVyd2M8L+8a7rKPwVPc/a+GA6LFrAyqxb8jIPU0/eHyYtCyWMDe
j1D2F2h3jujmPbJQLM4xc21ZUddqoi4AxGsYpQ74jRhn2OVmt8VOOy/RJhWzRVRhihwI252oscgW
XTa8HqYWAYWIG+mP9GYXwqnreZMFVNWN1VRn61kQWioadqnGH0Qpnf6jZ5g1aXs26fhA8/xAt6k6
6QdOZ5A0QrMw3rqrBXqRIf1RKRstSBT0523+Ybp+65MslmX+ulEA7GRSDoaqAFbEOmPv6wpkRDId
PafaEbRO9IpXrT5ORPHC0Na26WnKUgA5pJGUbrh7qHuYEh33HhqpBK9eUlftOeF2lxK8Xa45kJad
SNUh2/Opn5eTuntMywrUHoXET3NdAGPJLIm1eoXijaq6UjSSbljF2f1LP7YZnK90DtbMi5wq00UG
vpCw+6sq+kogtBA+P8l3wv3693qFzqJMzcN9G+DWSux16b/dns0zQ3NBAc3ns6L5SD3Vc/G54bi3
HOz0JWxYsyNnQ5sesuXU3A2b6fFf7rtJwysy+vURWnMaFH95SkYurPHeBmEw4XH2jO1r+GJfXbfQ
5sr+wTMXjMsZsh2EVKX5l06tQ2nLqDPhLpl5q2/iA44cEeJSYD+0FnHEMJozOny8HPcyhE/4pgZd
Y/kaYNesykcWeUes5RBGft39VJODacZeEwE2ZyqBSDLnaJH/k7JgTCTaDP9+dazi8pvCqtBloj8j
dn/5lTWeDwsIzhapxA6rjB23u/ZH4o2auRd2V9kZ9al8dxQptvFPr9kuriO443Ol1S4mv+5uD6Gf
RvroodOagJdJslBud6mu4EcmmygNkldaQmUhGOYxu6vszNQnyffLA8eSbLqMCl8GmsYxQEddoeZO
ocjE46CFlj+xXWJfMe5sRKmHJ7UV/Ttj8Y3lPzKVmKiRbVlpD8cgKhUypLhLm24RlA3MKdqZdc+M
Ypcevvl+1nSC8lniqnLKo5HnA4YgNXoMlD2nQacXBHanlf/MpHj538ia/L9YtPmh7HrKYykei9k3
NzxXBumEpqWjN3t7IAmFUfSkNNqVFdvdsFrZPiXEkhv2C2UhDnsG6wHBTMp+jDH+HHSJv8Vs8Ryb
LPTJ+Fas/wz4KWVanjIAQk1pjlBcy6F17rSdaBLjBWBUFMyHU7L4fkHvAdJVjO75kkHTN8BDchx1
qHzKqrhZiKQBG/f9dqzXf767fhMfMJ7VPE6ixN2TzTe9wvI4PnzT8gG6NfW/3HXqSGEIVAqSkxtX
xs6zpvP24LRHJnJ/6+5Fq/I45rdaczwT1ADoHPvrgAggFFU93K8o+undEmSB4sgdyhKFI8w0usAS
0VDGnXZTSioBOYQFG/ib9XHG3VIsH/XgJ7a1RtQNaM/+qCStp1ctjGapB0vpu/A1gwLq6MQ8DXxG
mmNAQQjbCen/PKEXhQgfuY31YLXEXjsjws99dISGjxfBf30bxZKvaumEudgcSeB1TDsLTuc14eN+
7zTzsJpyAXqZq8CXpH2cgJBbBWS8HHbBUgQH95mFHt3RtsNQf7Q5mtGU2sfOtd/Kw+SPS089r/Fx
Rn6HJ/osC5NispUV6fB3oeTEFROLI4LVdOUKoKKMuqjMX4+/qiSdgYiggF3n9o0uFq/gFxBm/eZS
nCAvl3BgBDugy6UdcTOjfOKaouu9aSFFrEVDgY2E7MTICFqgNrC/BJs2+3uxvWffvWCuNwBTyWlE
zM+B5/0YmDj/0iZKl8j1rIvtVHAiMCMKZ/vyfIw7efsdw/yT4daD0HLKEy/MRNHF/xDfls8e+q5d
gvjCAtQIH26wQs6Y2qc6P2tMQi7TZwH9zRO/PBAO8HSbCLATVDjc6KZ1ENGy7V4ppOljdKubW67n
Guu/8T4Zho3t0+i0MUsMadkoYlRFMKoTzqzZKuJvgY0L9YlnVTq8a8Y0krJqiopgnTbE13snLKfD
g9rhvrLaB4KsF30+DEoQVYeLBhvx2rXfaNBgIktvnoFNOKsHNYagxHBkcPSKUHMN/nnsHU/oIwlZ
YIjbDUYzzdSu+gnjqZKwpqQfyq4X+5tEtJwi3BrautOnLe7M9Tad+e3ybNixcKOIxmwxkUOo8rxF
tlfm6q1/LY3vnN7nqTpe8vJXaQUuFKdS73R/mFDdCK3cGDeuUhtT8G1l7NEYMOBMBNEazG/lGY2P
D76lNl9OY9DlbWCqFipCGc9OTqrzbBnInaDKkiWMEUebEI1QmjdCBijhmG9vCXlyzTA8RgsEwFnZ
wvfCyIID8HPbG/zWhQx7OSBOzOO3BM53pX8MkTcYD9hN2PPhT6h8ezMY9DqUMwKVPXwDHxHwTLJJ
14nCIfjuAhEh7bkaaOibNEGQOwtng5YfCWz7W0HAM6FdRdq+eFZVOF5GjnbI0blqPueFxgQsyYoO
+42kQ5ACrF7jdSVjs8qHcbGlnocjAnSIpMzHLJcbY2e72EXlUQYvqhxBTLll+ZpXeZZMYflxPjJl
WmU7OOQMCGffKahqAVsY4PS2dGEdtW+MyLqk+shzBOV2A7SYyFkJO6bpshATJM7M2P02LPJXAzNE
IrMoKiVGtqww2VgSXxBa9FaDKQwQWVIWDzTUALh0OLF+B/JNk+lMj82ed/Eltw76NwdPVE7DKoye
laBHcwwS/QxtOCSgG6EitnqxafdEA9hTKuQXnoiiOpuQamZ3WdoymlCCbnqmXlBxdrd7csKS3X55
x88hUXEj9L7WIpTgj46oLswg+yauEXEJWtRvvtuwel+JLmLRRhV4sMm4o+6f5L2s8gfEiCmLm+he
TTV+ZYIwxmlKBVKJwDo/fSUtiYgZ0NqMiEKKirG1DEHhTfpux0pStzsX/RmtMI/wpz5OHlE3jDUq
C9Omlrgs+2sa5nXAXiYUDe/mwb0jjOZQIXa0L1OQNG1QAVMG5iGEXSaNPuUDkIa4BtJFqgiDbhS5
YrptRb19fBtaTqGsWyWx4pMq7ZIdx1Kev40z8QErPBiomrHC62hEumcBb5qMzmoIsLJ1yYX08t/E
aA2Q9BnGhdM/9UEx1/svueFMoptoyuzCcIMDxhZClIAzIvzeZ44hb0YfmNE9OdU7j/r7qvPAkVkK
x7MRhy+Njw5GC4udGoxJhnEWJLx75VC7BAK6VQjwD23Hl7M48yOb3jUk1C/cAtfQTMdyksrn89AW
KLbHEbwGGxFaNPYXT8z7gGTeVerS0aSoxm/QGu2kf/Av/KBHJFffOEN7M+DioJdZ+7l+whjVSOK8
Qcg5NawNlBLJqtH1rNT5/+LTUH2V9Hvr5dlTJ/sQxvddKymvrf6fbR8HH0H/hfXchWpMaunGuZ//
50YC6yQ/js9XyAPwJR/Br1VJPTWYRbv27K9greWY5KtHpGUlyoQ0Kb/vGW7/vySb4qm56m0K14CQ
mc+WoFnctAGpArYXPky5KO9WKJNdNK4EYcOF2pV55VPkpiJHt/AsybcPVlg/aJfHVSNnGyIwRgeB
koGuK8Rlmd49AY/mbVRM6+vhK1aiaJHh8bYYEh6QaCBoBmiCLDPt61SyLs+lgWOZlBWj4KiuPnVi
aeYie739g/WXpJIoUi9+ZNWZIyw8Io+KWj+a2QT3y8pyRL/RmKRsD206rWowwrlNqPzwLcjpAL5r
uJ4rvYOa+ah/Lz+wpMz4Tpe1/5GvKliYGaVMA59J0dubFKya6jCbfZMLl5PgwhcbcdiH/HzmQyQ3
+Cqr9CCsIV2Rmi7iEaU5tYM5CqT3ZM9iYa0R/J8R71y0MdB+ppKlkJjmyEJDdMiDugg6DTfCxLgV
Y3sorybCdtKkoVvDXFWFu8pxAQjH5klFrsWr4EpudD0wyyi41/Sh8KxuCNhU8OqTHrllIffgYTH4
MiUpT/M/7jGXRoxt/B0VBlehOfILKIx7fJ0Gc6JpLvRubNHSPv4yQ6YR/DrTCRf7Koz0vODksN33
RW0LeesYXJbEZ0WJR4R3HPRHiJT4b3YdMI0Z4N9zfDwpLA592WtyMaLS2k9dTEs80WxC7b8LF7OZ
fsdO/vhAJtqpbYW8nKDBVk/k+el9uEHrKIWI7iGngVlMlTkO+dRj0hGX3eXDqQ0U8KFGdq9N7pK0
2Xqz73BVdwuEjH/MsB3I6HSlxV8t8bAiFdXFu+aCvDwIgGaR0/eI0kX0ZxlNPQyYW6OHd4gIKeMC
2SYP9SUE4Tztl5iOXOqD43ZCgR4Dou87ZpcvAdr36233oLTjIv7fWxCwhlEgRW607oltcgtkdK5k
3ivi9ZXgmsdTtvutnSP/O8Cff/gmCHNzsg4YQWPA2YO1lH/rCVZiMk0jOIN3Vj6UkQTvWN4akrGy
GzSXE/u9OtW+ePNgchJj9EZn1KA4X2vBzVLugeDXyw7AVloIRShkTeEsaie7/9taFhkxgsAcjjwa
G+e/iiBu+gIwQ/6wfSlfjX7vacXvsdiCYTPJA7foxHPEP+PulwWlqga+5796bbry+I/lCemggrd7
pETBHlRux6qIx1Vwrg8zachWpUU9pA3F3S5xAP1x2vBaB1/7reaSMeK+FLMi37iDepxQhvAIKTFs
ozKc8vbpLKJ6WMvDGVaWFM7NSp/LAjFRnCUTPckVImpdPxyW4BW/t1pCirFvDuQ/Kh1kz6paliUQ
+ZNzM2VScJuDgCFS/NaLkstJ5+wxMtsnXwKm3PzM1U9it3UDpsmjZ3w2T+m0bMItTwK7C+eeGdQs
4YKbl9HqMDMUk11XEMl6gFD67TVsUjtDo1o/tA1sCxe6a4V/D2pxZ+ERUl45cnbZYReoWxzid9Ez
uxMAr2edaLg7WvUPFK0/eCVFNEde26OCad3r53SLBSm/2qJSFrKDbYwcjSyia3JI0uZPwl1bfNNh
uJw+mWAEsW/XTe+RwEX4lE01L98XsS9bnjxOOlFQnzsabfb620/uzLmhRK7z90pBzG/kj4h+Dgy7
U4XlNM/AbwkLnC3ygp+4rFlJ48xxvZNSKgdTrXylYuarz0AAWevEy+UIkXd02Wek+67P/y1jB/fh
a8fJCQiU2cY/Pf9MyvfL7PaWIyimjzhQz/HJW1eJumNhJ3VcCrSl7O8DrFbXdsmdzqHKSiub6wXc
r2EDIqlVIT5RMMrVBxwiTKnr92MxNA5IovSajtHUFcfFL0Ehd3/BBS+lHmxfekNK2TXbBTr4onvW
NN8jucDsPPcFQpCnzRdsLPzQSbKbvKBXMdpcIEN0J1nn4FUySuedvMsSsAHyrf4IhIyybf78ynos
y3wervsjXHCKkywLcbwB4bTsWgMjLpdHCeJVxlXWpQwCwdR+sSBsYKtojmIx3iCMsxPINP+BqaTN
l1tOdpDNRn7SAv/HBWXdfrUdWZzGclPb18XJws1HglR6+pvfAbd6VKzxk1rUll6TPoBe2Rpj4uSd
OP369mHnBJBL1bnHYm6fL5vSkrqfCbXE7GKj7AYmEAIjhiVbvRqSJG5sefdrF3fxdLIz/OxN82gf
w20Fbi8i9x2DxPVOL8SA+kNKitFocq7HG0smbr9UO+cx6hZEp7TXBDMjtPPGYL0Zd9a1jty64J4z
jizwTkpyVrMwCjU5xDs+hvSriR1d078aqbwb2DheI5xrMiLoYZC+2Jq0ZcvHARHn+PLZqUyYLNtM
Z6pIvMJahy951nEbh+IsBX01vimi7mkvZkgaz73CUiZxLpnd4UPaRaYgy41bafFfGSVBtNMsh47K
la3kj3HaWPd6fNNzF6OYgU1p/jdKisgl8kQE1G4J2WTRUR1hjH1G1cyIyUhzesGFVqkfbqUQ4aGY
FyrdgFyF58Znhi4gvGCJsdpwhpStc20gw63IItRZKNQ4i8N7Zn8Hle0xHAGHO4JFsrbBMccPHufW
cK87pDHkRooPuk+/lXIea+bF8lYxGxVj7ARXIALTUzqYuTtSC8oDEpnlw6/UDrRpG+Zjj94VMomS
ypg9rgIovg285ri7njhmy5KZ5I0eLP7w/RUuu7KffLHPKhD/jYdGURzroLzHMwckCXyYAjs2fKuF
wYu9RVhZlggidmGuWLKBFeOzOUpnxI7CBqPl26EJoFbJlQgyLWlyLhjt1/IAY8AK591q5304F6Ny
2xebFdsIHjcgy8b+ifVSTTjUb2QINx1BQ4A47cXv9IknAGpptUc9gi9zzN2fvnW+/C1kpGTofU9z
/6CdLgk1SgdcTikIlBWilHJuymwPS7mf4JxxzDzWTDxf0o9d87OOPLn6BXrpBHrKCYhPZOT+q+LP
tDvKf0txUDdeyn3KDGtcIn9xpMJEg1ZsVMx7qYtOlfxss4Nx60nzk+7MC/pArSpDqAlx4xGxYsZY
sILsst3ptZThp3ZuUjaXpD9SppKkjqzdkMaaCi6hFJzOhbpDwhh1vLeM0wB11Cqyk0G16SHVEYSQ
+YWHqNcoh8SNONhqAcl3O3nWSfDTxJDj1PFyUSY3MjXTONRYY6vuNPheQBkw5ti0nYX2nHpI/GIB
FWtiuy+VsH8xkLwDBnYildM1IAxZJzU06S54LX//3tmvRQSD4CttiKFb7F1T97Ju51mdnzCN37kD
ozIOCh/is0voB3BXCxeoZcHDtU36nIoeqKYzt33vyqmemm7Dql2Kc6C3/pxje4Pm+PaJwdjbLgME
eXE8QPv38maHofOzRC7eVCHEs1ND3XHOfsGSomf6opqotErBc/ur4izmT2A4dfnrJcMugm/tjp+r
juzdQj61GQsTNKSkPd1hA/aNgC5e1tL70T+NJbq2GufgG8mDhl377P0pCDXEY0RHvvtSVCJmA17H
/Pzx5Lk3zaDxZz1EYQkAGc1gWCKGv2+Yu8bKHFde6uwUUYKIIqiFNX9GIcZlBIVgDBySsFlOX+MR
D5qw+A8NNXi+4MLBtgnR7PgQEhdNIE4YzqkWW7Zc9Vw+LZ94aQbHFA7F3tTl9JDNbK0nvw3003R1
wVDxE9c7G4px2pWmRPLL6FkoG3z/Z1SIa1iP1W6w1G5+b+X82Rt8k9yWx6CHpmE0hbp/WSfb+ZvQ
cPBqp3b919DL0jU3TlfNq/+70KmtXINj4VFdwbUOseIbtwsA71jMus3LF78vXF2+OZz7puGnp3wF
GjDO49hnxWL7jfdFR2D/GJbX/+zVdTFNGmUSyeOoz2ll8kYj6RZXu1gsSTTJB9WD1iCtpGChP0p/
TOGaK0E9hXE19ySW9fI+kf9LEIDG7YeqxRKNo+uYP3wWNHy+q0qlKh1g7dAiy+DIUUGODYtWTKRN
SPO2fJ99uXXoYhMwxPRymFfPui+oArPonMOIotknwRk0njV9RokXESFelK/ZVrQHvHaLTUUd3L5i
KuQkXKO/+KyxJkuYHUapGzZCqBGLJOj9ksqrOqdduSDowtm/lmUg/68hMnHij9VNyof9CITuzSp4
D703q39MLZV0lU57SSbT/kDOnyxNrJk9NSY17hdOnGIaHsuWfjkaMzcoYIr5OvGSU1cM4QIuR50g
aqjViwiNyJkQyCpD0wukFMB/b2Pt0rRbd7q+wB/RjS8YyMNV3v2HpgxgxyAJUGeZxSR3RpaBzzkC
sagFOwCrQE0zKvniBIcFDC5JhnU/bNSszCm/MzOiYXwh7AM6fVHGB+zxQplKc7iwTazvFyJXAT/W
kZ29RthNs14QeRbgg4oaKLBv6APypQLPGzmZMGClw2MQnrZrs8mgogTvrkso68UUxnohMic1X7up
J/gwrOQPkmd2tGLjVqAea+Hnp0/YybZo/OHqi2/MDCSMC9vVzAK0qwiErXJCm9FuSHcFbhO6c6SW
4yWE6wSlMTenzaVIoJjVJE1ZjKAvylxwtEJ7W9IgkmlgpjYohQNfk0ZEMIaOxBzwzBfkNxT/y7U2
O9kfCwx2sN1sREyV9FqHYfINjECH60lCzjt7qZFPJH/O5Pr4gMk7p57GAFLISKaRPJZ78vUxyC+U
J2Qm1+qE5pm7K8ziCLA6AZU2YOG3aMMW/bOuAZ/LdwcgspkzC6/SIEsOlJavtKMsY+UGRtQPivK6
KSwOzaODIRrTUoC4CqIIgf0CuyobfdafiByBsL2hp8lCxPJe9FdLN/HtDtVtQCr1/p1ReCglVqqL
4E3PzV5s9JMlQjrTMwu3Ks4dHtMF1S+AJcsOam6Qitn27nAA73c7HnA+3pYaVyR1dajOgGgJRW4N
F2dLbRLF7OhYDZSdGrOSnwukXJievZxs00nV5DaVZlfdCwmnMDRESx0R7y6p5q6ozY76HYxlowgH
QZz+tBtMqLK0ZGmGern6qVhAoAbDwHpsB3MQv85VJXdGDq7lQOtBTQpsHlWVJ5zFbn0ScDRGiK+L
f1TeiXJLhcrsurRo4KY1bwJMh0vMjfRGQC/f/gqJHqFArHyg62GsJcnMQDYoW9rtL8RDuyUyaW4t
QAdEuFN5yAorupfsEUweh8gCyIPAJ7F2lisrtI5Ke4kZ0bwItDb/PRbi4pkLgGKly6IDhteXlI/r
TAnkyX4W2D86DgYaEWMUnv9WHAeuuexR0crjiSqhqJqgkwholUKZx4ogG+BrxJ7MMMEGxyjgusHJ
9xfF742+CyDbYPK6f6A/TgCCA4JAGOxLXba6KrebdgDIOEfrDYKCR5JEECEevxMFaS0eCo5WN3o6
XJ5Kr3+6CHhG1C0D4/kTWyhqYWf7Wc8eJ3y+7ot7IoR7R71SuZ8SZwQIQgMRYyhCihLOIC1rTcgJ
+hql4bNk745+XaoV05IMepT+gYvblXje6Slbp9Sh/Xo97XTyp7Al/Zg1tAF42vMcYcuXuEKV9jBh
VsSqfcfsIbp3+VIRI9QThjXF10rdPUcChfyjwDd0yxko4T2OrWf5Ax7Z+qYXN7wjz0OMj4yJss+o
9cxlgMLRilobO1tEztaF7jl1w3n9WvGt0HPjehpuVEtcJ24MYgea6EDbk6GjZQiLRTJgTsr6OIuD
smbKAYM3f135Zua759Gr/ikpJg5T0wbcaz2YTC/QtSB+VlYACKc81wt+B7nYNHiK4+v+6owRXOhv
CAZ+GlNbtwc0fIQpBbbqe8L7jPqcKcZipFqPuOVdchadO+wFnYf8rJg2zIRJUBnago0SEQ+K8IUk
Iel2drxygAS8LCKjX3xSfIcjantjh0ebjVhxJIfsIrmpPZ9aRhmsLlOPY9ZSCtnOmIkfDfZleIFM
QMjRe6h9yNRVErz/w6fOIrQhZxf6nsCQHWq+b7lGv7CiZjkKGsD03WGF3VAhmjfk5VE4Wn6ecgzz
3gcqvtphbYJzV+l/9BiSLYYPS/1fvKvK5txGOvc4ex2ChfPSgeNpzFO64zLCKPdHyv19tMZJYzQD
h3gfXNuHAP9kSu/ZFLWDVaxjnkmNPe3uUfawRpK/6RW1UExQQ+As9qMnwLpTtR3Q0a4JZaH5Qx6B
ZfMuDBrTKbv8bCfFzwNyrW2qUDm18tlUkhgg31IGO7Am7YG68MxR1AvZFSYHzOmWR6HjKbuj+fY5
AapvsVAgVVPVE9p+2n43patJfu93jIsXJtUL7VDteQ9az/fbYXrmX8Gnw+K4LU3YS2zIfpXR+i/O
LRjluLQt2w5wKZ/gubUJek2ug3zVe4N5zOqNWhrsAfrtlzEjBHT3k+xABdjdXYc45PkeUnaRS9sO
3gbNXGaXNyrGuL3Fd+AAsWkI4Vc0x+TK1AsfFcjJmz8ij97mdow1ZaVtPGM9aX4ZVjWPPc+VF7Qo
4smDBA2bXMK3H3iyktTtmX3iteknXbIPhe19QyTNXbiQQ2eZAVrrJCsbZEb6+9kNZy9WKObO1TLZ
KGJaWzAST14VA1GaRpGUQGWWvsxMgZuk1+9aNOQnhusxfQvmaEacGrHQQ78tg7M6yMStkQWnznIO
fXx9yqkgiMgaQ4xNe5CzYVEJ87pTZYn6VlL0xaeHeTht4x6KSIvK7Qt9e5wAOuz4H+Uz+MbzLSRp
no1AA5m7x1R3234wKLGgKCy4lZpN82IBwsPTrhrglVhiFNaYanuBYZIxJxSWcuLgVGkT/UfICDas
uhuu5PvJAuhSWv8dOfSFEavtBQexjCjrb3qETIKd5MvuLoiFAlFt27lUzr/Lqv2sJWrBm+Lo1QzV
XaLs+u951FbbRlw8E2GW/uYLGMPkDapaOzPTiEEYFu10LtbB07GXI8UaQpWmAR3HcpwcLHN/kHnc
Fo2fFvVNiSzL4YR+oLJD5LsfegDYUExL4lKBkWXxE7c9U48aVl9VOWxEnpl7DoX2NqPbf9jT4IXX
gcA8Shc77DhROZQXwd47M+xbDmMnGkrm0/LTkAhnJN/aN9EwXOKYbxKmbAnY7iYZ9GSprhZBxKWW
ZsmYR6k+w61VPmkzQUJmSBFcIv4REno/jx+KkIKq5Une3lNe4kHkoH0XBP5On28WJLPu7BALzIDI
e2/DGHAqVgCzWJvrM3/dd9whuoRn7L/DImFxHQ6Fw/j4qrQPv15FbRBjI4Mi7eO4Dmqz6wBrEQUf
+IPvsM2jFAxQFvpg0QjzGgihtzIK27WoOsyxvUm8qIH/cIVpdJ2ieO/KW4XEasHty3cezGLuJ0Pi
WqtofeqwPSlW7sB4weNLjVbSDsILFsYAdSECZbjLdYupALDQfX3d4VOVeTdTuugAS1sGg+1w9sDg
TmKeCzgtgVPd8DwnY/IoRw61w6PuJJ8aNDL5ZIO9ePlT1Wd0Lwc+Jsxd0n6xcsgfY3J0inIpCb4d
N9Z0KVbwnvnQdF41uDD3SUIJ1o/eww1cLQRe3aNnxvKgi4OkSeImy2bXcwLGX212ahejiHVPqTlt
NUnA58gnDr/fAT18HwFFHPMeVLwy4Nlwkxi90qNsAFgu7B4CN8v8TP40RJDjqeha1nJ0DDAPEdf7
0xuIg+W5N74Ar3LrLM63f2GcwLRlGhH5eaeLEV4mhZ59U9EZ0u4WzFOyrK9co47bFYJNd8jhnb1I
z9a8RywWDFuwemub571l6TinhpDSRK1cQy8Zpik20NwaUkAFUECkSl850WPyi/GHhjEcuVt10Dz1
6XJfl0inyW2/OsZp9jcw5flKW5Nh/61mGO4sVjtax4hEAbtzG2c5a+NrdbhDTGyEKpoYV8bw0UaB
EyJhaX0+Ta6mvb9VJmSO3NpWm/VgM3/fWWHAuZYAuhkE+EGNXhqaInG10s1Wk0PetautNr3flonx
mAwM1smzBzz7Av0eRZbuaVRjuR+dY71q8t52cbR5B9SSeoj7NifQZp5GuqaXTRdJhptkiwS0Tq99
BLrxvwDpBt1l2jLdGbjY0FkWzdSB0aqL+gcHL140l7fa8ytxD+TU+2ZU+yuna3SzivYaEQYI4EU4
VhsTzS5bEy/vCiM4QyazRw88sWEqX0i2gtDql2tEoWd85s0s8ZwLH6R5sKzKKr6zM+MSW4BJ/EKP
tWNEvpPTaGqyO7uBTXq0wY/KrNOr631m/9xpiIn2E9SoS3rLz0nrHgspAaStVL6vjgs4PMWO6WuN
O9VYTzIt0uHVlMmrgv0/Do33xHrk+hPecejtlmUGLqHYxmz4/6szHcOK+Oa7fxZie0HYZOxzrps/
nNikrjKC2IHn7HnhRQlFXfvHuktnA7lQj4j2Z0x8brugSHiuEBsAD19uIL//yuNw2p/4K7B/NhHm
VJygroxUUn0T8kzjnF2wUHvI1bexIVxelT9fe4ePhUSKp63wZusE9iybcgGyGvpyL/0g0GnUeaZI
ITBpB0b+laYZBw1lktevN3M6lyMFpc2Nx3Qics2HfGdIkaUV0Xn6XLlVXCY/blFx5uCGrBleIPnc
KDSXgHrNCpravXKUwwEZMkramTtmvujiZzeE/P+/ZVe5aQc+kuRsbpo9HR6uQisyz/a2XqHpTJ/b
BqJbabyrlaNtmaBdyqgG133LkenGUjLGd/t1QZE1OEiLFvB5lrqxYpyeo+pqeNUqBIZeDdLCfklK
8CECgS3DoyObKmTuhvoC0RMJrW9UklrIeH3uHob6yPAzcmk73xjADI5w7DYQ1xsDMfwkkw4VgQ8Y
MNuUDV6yWkj/J5kkGZJZhsn+OyU3G1l17Q8CNvOaY6uVanlmGAhz8XilYBEQJ7d0SCWt9raVMIS3
jjAuN2hEfc5nKmXFzzNIXvxruoqEPN1DguaP4Dvt+znKz/ufgQQAzOjtTEw0ie0dYaVc1K++5rUB
kdKh67ckq4jtGir0XJf4IzqqSjGPNW9PgiAcBgQQOKatl9O6gV9X2pLjWYB9KL3/dztiaxNDr9C2
UHTaUJ21toXIlNuib0mlTPK3/tja1KfUb0KPK74Nz/zsH2zMxO8G/xJGhWzjePG0syAv87XWirZE
F/Ng5nBZsIXDN8VUGy+8JMUN2x6xLJK8U71HqgmhCnN94N9hxwVkNahBQrn+LLCq/6moMfS+ECYI
pTlE4+45gwqCMKDuoGdop9T4uEyfor5MneB/AvMGDqSHraBOaL9WDQKuZWjc2zjtTRKmJUojG3Qr
bIUkaibqEb3gBOhPaLtuvWuUACZ7d+Foa2/T68lauBQauLByS/BtwBjqNjGfWQfPEXU+wB65EnYX
dAhLv7fF7LqS36+p2CVZM9yE8jtZDhyK0ECaZSIKs+YYYyKWiVC+y2A3hbvzpFRFNI5qy+vUy7uQ
kRNh/VxkifgklroD1xHYb/4I6Tl4Kf48jukIcq3iRqzaG+EIkcUdxlsNcjrG6ijugDJcH0XTEAto
ssz/5nH9js1YkEFVFlbOFf8egeYmOIIpw6brep1+uZ+xUK0E4prBb7uNEw+diR87jY89YoZ6I1fQ
N3eZIlpiNxqzon4Ce2eOfX1tkqpO5AoreA/ixxaklQF5i6YXfc1G7JQff55OATz0MIda4hqv+FKd
SICOBJkqTdbJUEp56/ntffpfw/6RlD5AOdzJqdAG4ci1ny8p/ZGH4gZ2pVsV663uA1jTojcZYexM
5fZHkEtaNOxWXeG4/trDBUh01TJYGjr5BdtY6TYR+QFB59ZoSRBiQB7uBwAhuWjPLjDheMiXCvQx
RvnrKQMf5XXB79pVzL7Lti1KQzvrpYCETRA90oslMGuHOtYQw7fM1bMoDNgBTZKcgg/Tsjdk/dJ8
2g+MiMgKwRUMDg2c3blWPoguqA3Y3CICG2zERF5BAOc1gDvj/v9EfqYh2AliKVJYA03Xs75e9YfZ
B0RImvELvDCG7Rr294+2hWYsGpRho/rqaUdaohnumD/HlVuSIsCBYdf5iSI/Ie8v6BHkPyz3L3hC
SUBoZV+BUAY5ST0/tJmvot+SE4ppppg8K2laikeng5vwv9208PsvZd/qZz4BeVcAGWq5ciTPdqBf
F7W1BBrmVNrrKjtiqjkZmeQd5u+fj4tajFp5O32PLVbEW14DEAUw4sRnn5/nX2CU7YJwW9R1Ce6n
lQfOsowSd9bZuyTKV5N4k9gSZqyyhD/w0kXRZP1/O9VIcZmVtUgQNt7lUTyCjHJv8DQD6LxCB3EY
fEJVc9X/SfDJsQbxo8XfjONg2JxXA66LIfn6oxsHO0qpjv700E76hbLVHVGGMbe+kQupmhwDw/mw
cXCka+YKcxqVjklNVlPtSzk9L3BP99KDCkDprIKjrP1JfikwwLOPr0351/AsE3RjWx8m6YGYKuBO
6D+2tno3gvqgNn4Tlc24HhNRPQzL3ktBoTlC+h30WWjnPifjgqLqEBbNv6EU4nWNX2XCjkGpUi7s
VRG4bVsqeT4GIarKBJKWhwaRKhA40HCZ0BHxIGgk3/1U+JvcqCCr6ahCWu9laXt7YLXuJpHJdGpv
SBomGXDlGky2ytpgkRRaQ96o+nhwAvE1ZzVUq3qwIecpka+H+CKAB1FixjpcBh6c1rMH5aL/6cxh
Nlagp97duYqyToG4HWoTiaDgpbnJWk7lIBZTgN2FQ1pilFyvAz8nnUOJFrHY8+Ym7GtOgYy2fFy0
9ZWQ2/ldRqY1psLWqC/aqv+6Vm48KiveaGN7bzuHDsBxedSVYSW9lSzFLesCynUfmtRGRVlfGaXS
3G3agr7UZsRhnSA/hQKs2jPAyTtpXXz8DE1BS9G5Vv7OOQwv7FfYxlwdOb7GGvqUkLzKkLOdHe7K
bEkxYYrUePQWCO9mFc9T98Z3jn04d2ZHg5UU8paU/kONhnwtYPFQrTvYrud8vmoj2s3oG+c/R/G1
b1k6wuS47Q3njjgXDkbqTYROj7rGY2kIaAFeFD2C3ZF8VMUL4UzqxW9aEVLL3QZxmLIfUxFOolK8
umg9pUsmT+mpnlNYC30kejVL+4skCShr2PEcsppPw1bjD3/u1kIZjVOm1RKfcjZZ5cbizai3Htkt
p7QlZwMHOLzCcdltYiE2xT/zRsltEBfho9W/8BvQtEHiC/zthsR0Z/OnrFFotey3yenRc5n3iWHH
wFCCK5pALeZ7YiW0SO4h08VYu4NPn4FlFmuNiC7FHdq6+PcNPAop/n2PU+ZE3+VYyU4Aj31+WojY
m9MGFylcPGmYcJR7m3Jhh8erxBYHGIq+1PvIp1Yw/rjgtdfSzXq6ii+9nXvtmypNapYPDnD1Njsh
RQLjkhneNHjqVjMHuslrUXccrv3GDTK3bWPZslJ6MKBPa2Io4/WRduojClgqaa9jyp38XHvgQ52Z
p8ohTURx/mHwlzvC0DKxIQnwpTuiYIlU83TTo2ig+KQE0NEGkYBFp5csmpXmfK4ezA1urHDDbkdv
FEDNlFZgdhoCfN/9yMhKBwpqJ7JuhaS22BKPw56jh+Kl4XTPAV1v9aNUAKPE17Qw6iPtBzSPFBKF
QlV94dy2CSqdrTQFYquGMUdAGOAC/BI5Fu5mffPXHdGnz9F1dzbCgWLTRoLoLC+hZS/UfK7el4xH
RKcK3LOhEDybmlZcLdOVgu6/id1+QSmqoykZXK35UaVKkC4zM2j34UhS6kd4jZo/szTRrAqgp29F
pflY0WWyHPA+jeaWgojd6jrR0THktyLWedS+azjAPtsUQMtqEg04dXcGuU+eKMM6MFSOOS5egvs9
5OtK0HHzMlgLfrh2HrhN9sdN2EfpDX6GVDHo27eOjTgZHit2flMrcX3ppZbDj2lU8ZzkzFKS0zUa
4DWYb9n9OV89R0JUPnS8GhQhGo7L8wiUcW0SqjvjUSn26Lifxl3yf29HzDWacLiqudjVNa7kGofk
3sTCyo5anrNZMlPc0KxCBLQFP4HEs7Jzd48IyGlGbA8zUr9ZhVHnTZvPgIfLmU6uPORpsvVuGs0p
OfAn2WctYE5PyZVBr6Fh+1UQhvMQCeNybiNoqZ7BWaSDcK4n1/UuMhSz9ezl1kGSa8aGbhrvsHgY
eg8wmFW9MqWzESPz64FxhSXh4F682CaLCyKL2/jYzmaMc3XKPPF+gaWV14cTYAWPNGeAUqd0lzcw
a6OO1aqJBuo1lmZD25bP6HGXaHh+70iuMJ3PYq731Do4A75IbB4KCi7wMYj5LSMGX7qNvH5jcvZU
uJzG2kro0sFdtqF8us6DLhDw5hXBIHrmpXllEybh4OhKiuN6IPVEnzH2gUR+yIC378CpdN9mVFOk
8IliM21EkLtK/WwJMlbOuXEY8npWwPGRBOymNUkIC3mh7mYYHf1rN5hPC415PrNbKx2QTjbT46U0
ZzGcGEqS9VUX5sB7vk83QPwrrIFTJIgOskEuNbBtfwTnC6aufkUKtj2E4Qz1dqbxxdJuTXjCp7Dp
4JqFhZFnlqfsy+jmO1x1Dh5i3OhZvyqfmPcyp3PEQ7sP35B8Ix30pux7HG3sArbNgJebrzwsbX6Y
0MN0NSj73h0Qq241Rka1pVONwkOF1GMGksHCZiT1dAcM2MJBMo7IYtO0Us73FVqKiuLcZvkt14X4
F3fD1+ltBKLMlHnyMjayjd9I8Fz8djTnoC6YwppFsg8DziyIx04d5ZoDQkRfrjQDBPdo4piXi1yG
vGT6kGi5G3lLfI3c3Ez+B7bvOHvoHIWBUOoz+KNhwPnZRbhfRQyQKL9E6TsQpEmtMVfc+S5GodOl
LUj6OwOytS5AemgxB0TDcSNc8pbnL+K9PLRXD4mOApRgaNZj05Pl7odkSKIa/3te1TGd8xKAm0vU
bwnkmfxw/uH3riW6+GEgtsbgGNhjS5buUi8B3epiXU3BagPJRYQgBxqz4fH+Fe35/86UfFg1EBSO
xkPnTay3f6xDKZGeZSw0fXhPs6ZEZML4BlhzJQSpmzjCmMLX98Nbt1jFpVSJbszBg++x9mvQcEEm
63eU5ykUaJnTZB3vszbSUnnySSU8YwxReOVmdR1vrm+IGuTr0ZJzHNq1LhMIn5KVc6hic7sAIZZj
+Qr/8G8qmpU9uABxhB701Jay9cymBfb8ay1WvHoaaQktBsLY35x4NBpWULP9miAbm+F6XTxUL6Cm
RTvMvNAQIMwl6M+kv4BCjoHSfZMdnBHW9JhBeX3pNRrIJnM91nHYaHcHtvhrXZcgq7GrJsLx4bcX
VWASsD+6LlAiXTlCPlMsFr7ti4Dr7WUWzhI5JaP0AQxElOKIToyosDOH6PB/pDLdLJGxzW8PZcIg
je2C11j0qWsrdmQOBMvy8/P5hy+eXYHzum1CStJzeoqQxZgrzGLxnd+23xueX9adnPMubZATwHEe
eZvz5TLy60DbjEDGsXUS7QrTIKQNH/40xykPuUZnEoyEd7bsru1ZJVs0wSkCEGzLGnsU69ieZiJM
bh5mmDQfGrkEE3ihtIdzYXVIDcq2HHQ6MSsFYFfgQjSRiJ/agdnL8N7KwqZERADLLwwo2C+9SlDg
AzpJ0CLMx1UhPsMH3aC6HT8awWLE8WQOzqoCF1ST4JSCYN+GXAvCy6AbCjfC6y5/xrXICqFwmetD
jbvJ4sp+xuKSTIjKzuyuYt56mXRCmpjF6nMwmsMubF1u4iNo6DYHG+FvL3hDUtBvfJ8c2hAmm8jv
pV9ehHJkX+qQQi8GwxA0iYFHdfWdj9QOn933fH4lZe7DKnZYE6XqmBUhLnn0wypIAuTUXn+LrI1t
F9VBgc0p7oANtK3aTUq9f90QanMrY1VieVCkGtvQn96Cw9UmnPLZavZtAjoJpfkhH5AQiCbbNaQE
RGulwjTr+7P6dfoiWuZg6sfacCY2/GUglQIHaxLLnNeNswVuuzQoL+Mml6U8Z1eF3R4JLS4yNPn3
ybdNCaYLgMXBuXO/eaJQO+TUNBpoLBNRXgnTwfF9rSuB6NdrBmtmF019SwpgBjXGdTSPUVkU6SJX
uc7KmfDd5wY3HpYXtCkhbG1y3RMZh9kloxNuFhqLTKAwlFpCQ5Ow5FK2AxKAIL8zkzDyc4+7L3fH
63ME6WyY6SoebL8SSWElUN7iftQhsyICz9t7T6VtbwkBxz1qaTfLNcLf2GaHBTQdJ+0+J/xki+Xg
0OzHScgkln+BjbOOyB65kOrbg04v/VTAMM7vzQ/201uL0Tc4hG5/t5oNxIlxA2fTyPxJKpQ8NPmO
G4kULFeTiVVojWJJA8/wi68SSF1N6kPQpwISiodBsG7WXCCVHrM7t3RoPa7vznlSJe/+fqaqQXcA
m3caFThrydJHAAflS8bxMNaCwuntEEhjH8OUgLWhHS+EB8bZwjqvrfte5Om5z4T3R5Wu4Vf9XN1h
Ec9wPv9qSHWLNGiRApDvpA+1BSM1GgER1OSxFEOPDG7JOSKmRcOsrZTpHdXGwB3BJofvwU1h9ho0
4/IZxe+zC+uDCuU51DhPur+7vieePWlOvxyXzaZC+zZeCUxDsLfa9IxV8Y+zrcBMprtedJxROUBo
trIHU8EbtFH5onFXCZdMz/JbxYlBemWguMldv8KT6h7yRaGb6f4n8tLW9HzYj8Lz5LeqcFpxFyVi
JFEjOm3rIsFmfJvy7lDqMRmxwcJjuTL4mmwJHXGiKQTyet1oAA59KGG06oPoL/BZ2Y4vonJ2S7cZ
GYdECQCk87vbpOpVinYDoxSLAs5IYncA5YwZrgXP4x5viYv9jaloHEHwR1ardQf6AZUtNKGCx4lI
L1YC8dw9Pa2WWGpiFkpNRjBGnzP4RusxBzx+nmAqljeNZCUnaGx5hRv2eiCb9JjbgEcRdc7RVYSg
2OLfqgkC+fForMmSg8W20yKgGy3FlIYLqQpOZV+EiVIJixI3OJGESiIvIwxCSYVvfyb4ns0VFrSf
cky8O2vRujZuGI+U01FhZtnKdCuHe3QkNrIswO/MwFpQkhAMiHciYzYFHCgHPjSLUxUbBY1ocyJ/
gHSmQ60IctMwiX347iyJ7qvKWFbdvMrfeBwf0/TOu2wH9tRGJ+6ch1JVxAyZ3wKbENxoB1MyJAGw
mk8T3wTYMM+evAdhzaD5SAe3M3oLYBp+/QWnHB8SqYNnnPclAdvmwENXYc4BMXlMeJIBOpAH11nk
uYkI70aDSzyVVe5RESJnX7wTApvzYm+K2SiYIdQWaDuFOPlnVtjwnCTOQmeeVfX5duDTxMnKyIiN
aUsjREPWj6mluyshTXGcY7mA26Z0k3RAi+jv8d6ok2AZDIrJC930couW9cCmDJ1laqIYCQPDlLdQ
Yy1KWJT95AI56deYKu2gAm5lBy7AbQ1Y0U4BoJ2azdHp50vjEOPfOME6ZduSu6IynmYIZPbCj59X
5+vZWoB3R70H+W4UmR+Qkt37PqWqTRnIPc4Os9QJ++3NTf79mMD146iVIc1dWCz7Y7+heT3sJT2W
xjHcqEx51+sSojgLn179jM6nb8wnVMkuFC8cFLo0m4F3hI+cfrReYqPUwnNlIUnIcIveDPprvncw
fro74k8OGQInAzyDOUhhxYqR/eRuiM2r9Z38GSJJbZq2OS4QiQWxSqZ7g5nStrQR/NC5acqor4Yp
P1hSPqZYovHnOeeyWn7ti2IjM8IpB/8BbPKhMhlGYF0i7zLYnVmrhM8lqfMMqRNREVU7U875MXxD
YEqdI69LjojbgLyaNeFNyK3Kr2xjiA5/Axtd/hD4oS/3aBKC3DIVYmPH0ZGPjo1LtIMKGUG0w0pd
dMMAVviab24by5bRhTt5k/nMqS9BFzirFKjsSKr8z/Ib0Yit9vXiWr2gB9X5XvN4EzhMok9LVhN8
ppl3/ydXU7/4lt3rWTJVwgLc8y3v0mY7F8DgoV5O8AZz+DsTKwqnJeOWymXg75A+lrtdvkyYBr0M
pVP/bKdWi8rTPGxNohE+C55Rk8sQhkF7yZa8dSd44ewgnvoARIL+KtzqG1koLOkoZaribSwPS6cC
WTuMijmmWMKzGtbYyownXy8DdrOfMtBMDR3OppkS/l3kb4i6HpbfnfFzQVc4YG7rGOX1OTjeF/Lp
FXYT3JWooObvVYkehSbhJWX0gpL1DV2jIyKYLX6Z01liUje6rMULqBuKkdvPIiMbk74UYtGnAm3I
0tM8zYZ9NkQSBkNxW9B0Xrda0CkO6vzm5HbbiLwEqMZr4gumqbjGC4kRDphFUshHj6OOvSu4fPAM
/Y5E2DdwaODny52ui9qKNs+lJHLVFEVv3eG5ZTlIW+rYu2F46Hy7iKFU8faY/gGpGuzNxoecACLE
TQ1vDCcTw0fqd34Gs4VEBGyAvF4RGFhKZweltHU9iRJQqon6xTZXJfEfLX+ScoUI7bUZbwtqBwzF
nU2CCv8VBkppDQj+FQmuaO6/ncAtY1Vn7i3mY5aA5+2FNyNiJ0mDupTN4KmOQ255aNZnaRYVfevU
gO30sfCZ0ST2m17P39ooI4TXe++NsOUzFKFqA1Z0Rzgj7j4BgzfKqIiMj3V1wxh19JKDRuoHtGlx
11iM/ohQssSj0Ygb62Z3D/rAfZTp5S5zpooYMxzzdoG7LohcZ+337rGrBU06gxWGb3W4/1sBoyWi
aJ5WjsAQ0JqZztnrMDvle3GSOSj8e0obaqX5JrHASeHlfTyV57wc+mXg9f+XnRWDAsOJU5vAlxpB
Mxa0YG9o/zstD9pUxqlu9KukhLlY6QuKSsSNUDCMYFNGUq47sie85VTkxkqOoD9h4FuGe3fDK9AT
l018DQ84eN6/dgUg5BsZmvRhPCTqjdDE/wd5hQepTl+DxlxiD28DdOnZcCrPNjRdCY441//rz45i
ezElHwbOQZIoXzbcIdD3QmhUcSVQD//CSPO3I7Wp2SXcmlQ69L8eQodjm842k/Qbx0XJDTF4XGyr
4dtwlc7oXU4LD9Eli0fI08N2Vr5wVtly2bu+YscowxQDMw5/CuXD0d/vm7rthmgi0wUT5OsWygtY
BvHtqLMY9L9vCQ7u+1gMVS7r3rs+ZaV9d1VH5+LV5L8DzrpHs13EyyqYKzIKb9D2Yi4GS4fcah9z
AiRldyDVIE0cG9paHHcoL8ABdF16G5wacNncPRebpMEwj9TmpQnOgtx+HvPFiGVEWusI1YM/IkQ/
aC6SyQyV6LIcIqiWm0Izx+sCcjPJds9Ev34z3GLguPcd3Dq5xDKJb2HQ2EnDUvu03D6jNWO1lrp7
ERKVYKwh9jUtGyqsiq0vVf62k+bLfUrd3vJ1tR6UBEO4uOkI4mxFPalUUXtFxji/Y0GTBZzsrxtk
zMcjQYcRVXvOCrW6EBUvP31UY3qkjxsn5Kd/Eg78GYSuKQlpJFJjuHIXtW+WvZ7fwwTAmS7qaX7e
btMSNuYARlajq7b5OnkPqJUhrYeehCyj6TN+wSWD9z0sOisbFgTBy34WxKvox0J0a/xpphTFfKBx
yTAjLRGoRkLhL2+2+jvipqY4A9rNEwauVTYLEnUr8amBRaWbSovVXnUAp6uAs8GoQV5Ry8vCevT6
bm51H0j0l+IrqtMHWXqqnQAFoibZwZyH0pzScbiyuCgTFVnXap1Z0nZCgL9sHm5xfnz0AyWFkB1l
z0EDt8f8iN7o0G6IhjYW2Fjz3E5RJJ5rIwDnjm247oV9QO7cvWrXPNozUz9WWeQGwbyf8dZD4s0+
RoT1WkThXgxindjwYzZfEmkwqD0eD+sHHEPXiFn4lkkWFKlFzEYspA6xP6eaoaQeZyq0koY+CACm
1JnLhc8yv1JiDp96Grgc/jcbCI5wObOoRIXAXgJKXXbeeecu/EDc+ew5Ia4dXFASMKAG9mlmCaIu
KiTfOwBNJ+lErrD4GPnlbGBeT3v2E1nHLW1LbI6oe55BYSAxf8BkWLv7mm5gDXT3qXmh68UajM3a
gxh9d9xd/YZTxzGANEVE69c6EfU4LkAZi7fFv5Zb4bNw8CYkwKzcze20BnwkzblWFIuxGkt4L61M
gp97XmZxFZ4Pksx93cMvKiaRA2vO1yq72cLIiyeYK8HS8H8ojLtDis8x3zGQ+lzAvhK2sJJOA/68
fpOYDco3wBLat1Fycru/iKEhbBjbyFNLIE2eWNWof0VYa8kjQETLMLsc6X3TgzFb2qfqSrgBWVy+
ETaxpjQGSoznzaCBEkm12iFVC2tygNmTkfPt03SQUjoj0WALd2mY1yLFX+gC4lqLpOkxAUSAdjMC
7mcKOPTZBV1LnUiB4/BZW5TYF3tGKA2a6/Bgow6Q5cuz6alM8Svg0W5t6gXDA99TFjkiBUzeFjL7
aijFyRBLc0uMJV6dBNOg4B7ZALip46CYghJFgXWuEPZX726UFkgZPwuzsqLn8OFNmU0HY9II7XOa
yJAKJh1rBm0KNdcPXLWfRvL8/0dmvDIc1hbMNVzlhJuRCdUTpjHcZzsHDs9TJMbvnTbZJmGM+nft
Ja4+8wvSlXiEtUVBpfm6IxbYyCLXNW/pEPpca2pjRu2FfXHWDev6q/b71xevB5+S2BvF5D5oEQYd
I8/oeUrcCspSKHOHyMEe47ubKdgEaWuOmG3P7JgoQOzvg0nyv96YhsjIXLMc+U+MW18/5zK/joZq
+zjtAsj+7RFkCtTDux+P47rumGeG5C2i6o2tcqPM0fhX006+yVDKJn5+S7MLhKay6VKmL8Cu/hAw
DaL1nsMXXU97Rs6m6NQ/pz8iNnqrPPtuwO6heatdPrrrVv8c845W0LyDUjo2t0NwjGERHsExqDxG
COpulLr9BUyQlHh48/Lr7+Fx8HIPJLqLuvxOdk6t4bBhZfURRQbX3gT/S/O7AGC7wsQj6bWSCkNn
CRKd7agrWoy31MJOSZn4gzATJMKVZwNgjzJ8vZuragkaD7eNj9aDIGPmXC/ggNro8lF1hlxnAIc/
W6OQUShdmme68W9UdmNrgctFbzeTZ1iuTpcQ7du9f0QzVKNzB7TehZJvnwCWt9Kx8daPDP6Kq+wy
zNTqHu77nKPNfuiyoUuj7Yibqm1579P/gTDRr8G4xX4+aw95Afc1mpFTUoQsUhSjXTVaJ5vTQWRt
OY5BeFUuO/AiT0zuThXFR7ThgwnQEpPfqNkxPFmwWDZ1lgGVAeSMyR/njmYdI3haPW1epU84uGyj
v3cHn1aDfAmtnHxS2h7ImW7wpK2s0a4v583k4uamUYJ5OG4ry0V3AnKoKgZ6SRT2e8dV9ShlltQY
fLDlY0pQR1kWytbwmybjNHcrnjVBMjs1NbeozUf8vhYNjZUQW3+fNQ9izr3kKl45hlw+0Fb6Id3R
4/1jo8GEIJmhPoXX+6/afn/yyK8W41In19yRFethR4Jb+3hc+WA923T/oA4uMMaD971MV9o10+5w
4P52WjrKLVzybaDL7+wYs7w7BQHYxdSU9QHUWeWQAUfrKeH+Ro4M7ZSKx7TW7+YegIyA8XpQDB+h
R3GRvBUXvO7HFzoh1jhD5nWDzaFsHhYdKKVqbk2/fHhzFMeleuWPmiTDpetycg4pf08h1a5Tm8eE
HhMK3iCesf1Pz78+TCcNpipL2Dh7ygHdCOQCiNsAF1RSJ2A6pgX3xNA9+H29SD9ley6psJu47v57
P6Jushe6NLK3DaAJcYvVAl6AyW3grvgPx8AvBIxcOZGAkvrQQ3p6PNsV6zmSCY6I+9TU/lW3Jqhq
EQH4+xQlepxOKmZCh0z/LudSI6nfLUClXW3NmNsTv3WJTNH6cK+eLy5LA2sx3BlVx8tStHVUXzNs
bK2cOuVpFD6ch+v3P8jX/UTkq5O6fThsNC+ogX6DbGdTfO1w96NWgtumFU9GiUQQRX85s0u/imAi
d2dgRTtFoFJmC+bVMwGjLRO7v6f8jdEobPNHXsVUR44sWFxxwjsGcxOzzcrJxQA67k0371jY+5ze
JlvwShKz7osBkInezK0+UUQ7wKlc0ZDO5ompJfFVmTFCdEmwShUpwkOTgo4I4P3jdwS4YCp0mk7w
V7OGjjjvJra7vdChe1i/N6reg7oGGJXwosp1aj8BIYe/bJAEdSMq4mAKWixlGPdnqm8921ZN/xLq
72Sk1nY6qBlbt4UCIts6gheDrBA5hou54zL5w9jn1uzC9q5xO+EV6uncHKygJ9TCY9BF+e3nroCm
KYxSVthrZhg0NwAURUI98TSBagZUtZ/AIMu5Rb2+X2CUlaL+sWM3UXYQxWlJxgYZ6y6CT004W6TT
wXkxYwYYehhuEzzvgeB86vpEcrw06gqcv6rRb1TBU8hgEdf8BeUx/OtfwibymU6ywQFXiKSit1Cl
LK4jfoU27MJldhpBl2PfBeiVKq1FtyPmhpbh1lwgsmAMRADNkEqPwq2D5tZJM2SSULKla+nudNR+
JntQ2k2G9K4UQl5V+f9BiV4i8eQI9sFEy4MPo4Av1rVu0S3OlgrkveEspkyPKI+r509SAXTfp6qY
2Ik0xo/nBX24sPVXRz4fXrihsO+1TYDo0guhGUD7Cyt+yAfpmQdhIrDvLBLCMtLmr78IZMuP4lm7
v7pAK6KO2QGlvG5GRtFVFNk+7nDJynq/E4YB6+F0xR7oElNK2r3XMkMQdXD4b6d0S6jvXbBLQhzP
GqnsKikuSCx6/TLxTxlrGgEh8xGBzGFSKCCG3HCvicaXI57sVSJUhzxMh6FOUx8SLVyENE8L7rCK
r91MlT0lBXW4y//BQrPioi8X9rTWu0OB6yPIzMe3kYAXJNP6BTuP/UpMkpZ9Kf4ba2UjG5VWSYqH
ULRAQbRYZM81zglx9D3GofwKHCp4EGmmM/O2jyfYnluh4MqSKWTfoK4oq3TTD7NfxswZeXEQup/Z
GPicB5NjWG9DhDPQvwehysbCYQA/uAynXYr4TwHgSkRKL+GlNSnqJNThircGMEFFSpsv9iGXYAwM
Ew1XKdTd8PHZ2ibJFJd5UcxBJ8oj2ronW7fMIu8VQmRPWnDq1woClBg/z+BB0S2Hpu5dZvzao7gf
Xhaz3pUkGxZnV3wuIzcmqwsS1MxQH5dQJfLfVtMl1K9AkCMFITjcEaMZMerWS2hFaqDv75Byo3lA
nstmRiAT29iRJs7IGCNxIY8RtCf+bvjAQBUNyY/XkLCNWeIssLh/m+lPmlLvOAfRmjkp+Q1DVGF3
SK6MLBeTuqFeUNFedSIc+/NV3QeZYMn931lBeomA2TS1w7LIp23k58P+UyQzEzmoNLJW9UfrFi9c
UK7gFw8ZRd/p3hhMVspmPho8258o8LpGR65FF81Yaye8xXZKuUtCXujEMpypjn8w6yBlXY53waSY
W9tH9gdBpARfFV/sVPeyFvrGYfnqFNa09jksrnfETX/RQGW48qWDzvtRtU0VcHl7uxXo8OqvGf2+
r7YkKpyyx5f8p5Z8hgVM64jtNu/yDzoxapzG8KJpi7vsY1OHJNrd4SA/MKAdWpMlkdTkXNRRIm4k
e7fgE6FxChQjLMGOwdX4x2F+ZU2SOsOz57jbn9Oa59k+k11YZVnS4ih8Mw9w/bd8a/whiWDJfSRr
rw5v8ZKxMVMHGjlLnPg3/NsOk2v912Lv+maX21Wxi8GnaziKSHTkgVsky7XaKbO6QpByghRWfh99
mY8pRMJl4Ty3iODY35dY4jHnlja5QqXde7g/CzScaQjtPNuawuTvLWr4ftFhKVIrAPmt9lMxtcLh
IgegWYLVBiP9cHwpJXhyXQt5XW9Wauhd8NlW1i0ynW2ve7jR8IEZBH0xzKul9ZyxqsqzhIgJk+jE
TZEGSU/pn6Z/eNlaBM/QJl2Y/0/2fU5a3uoMUgm8SYkntUnRN8A8L4FRvPqLsxX8ciEaM1JIFD4E
GjBqIOo73JlRGts44wCpwdKpyXXDrTvLpvlov0dkKSGh6BKhByytxWjBLzUT+Kac9V5guaB7dYp2
mlFc8eiZR/c1H/Ho4HAhcXQtj+iElr+cDPMJmpKm/Xoe1uygR15G0D+AMBhlXV8/xyHoTX8+r/q0
PdLmBFG8RYP2bLdsh5b3THKMrr3k65x7Dbena5c+UwCpkb2Y7JLhTAJsxQFPZi1e1pR3Sd4hIOvw
4TSZq6aFWYuDvRWvXWzUZ0YXDyYSI8U91H/zZa6haWbrrgXYA9PH4bziGBhqrfZBBv0Akbj2xZRD
rJ0lgpv7j8LscR3JO87/JFTP/eFmUrsU/SW6hhHoo/kwee/sIfmnHmBmN9NZ/vxRGp64kJOa5voj
V7IIwOxlFAF4x8E1HRcYM4WNHmx7UmybsDI3yDmkQ6F6C8uZnNHToapcAaNXuj38syvfj+NHgleh
CSIDrLiKxDnjyiumzqBOLuw9hme8mgHbhLAhwy7WIIet49kZnboC6F7M0aoPZvN4vQ0Zi0HJv2DR
sRyO/tonPCkABEFBk70ocOS/mGoHHOwhuCLpOtjViWyS66gQvzat0ISNbyqtbD+oytRX1n7tRmMT
NCJLkvg8ImRpPavV853Goxg5e10UKpsapuEDYk1E2T4q0I+ouj/PBgjCPRKZU5M8tjHR9DqZD04m
YuXW9C73B2AOAVe9NdF8lPBgmHmYhE7aDdrdLyfiA+i71T9Wd+Ko9TiXxS36TPLDQWxkS16Uex7P
KxrMHC3qGuxhD7T4e3G2DBcHfl56PlEZYN4GgO+RZWgeUD0k+LGa7FuqgRtt+e4olJsP/xuqFXvU
FPJv9O4mc2vKuzjv6fprw4a3ar1YhfPcafovym8jVfj29D3uQ02BY2zNMSkUG2cd9Al/En+oyO2I
HOV2+cdbSvKnrH53hyk2BZ1y+ZTD856WA7GBKJozmm8WdjJ2i5pUOavVZdmJVklGSU/VSf5WkJfM
OpqHTcKECNcAsj6ezdoGXDYA7SSaKa/3FbCVpPZRmiT7QoH+ITmRu/8zBIN0JzB+6iJlgL412cpa
aa8XgG+c/exud83lJTc6IZPbe5GB/0ou1ooMeqCz9/TZU14RQQdiCWbDYRkvmIEtGlosuh5G4QYk
Hfg/FiQeb2QGAR8969lggoVGUQuH6O0Z3ktmMjJQYPtrARlaXqHuXWFBkWe9jotunjIjyt0JxRJo
P+mI/Y9gjWjbutlJm5GG1chn79Ib4NH83W4hlK1vX6xxFNNsgtA0pzxhU56yr6WX2GUSQHvd1qg+
8klBZISPuodOliCVPT/8V/+kx3skKSkZjg47M+5COblWzShrqQQkzKugCrQT/pFVSHqj6h1ekwiZ
sYIzd9fP3zLAl+kbzhdWjNL+c40eAP0oSMYlyvxCbV8o/bu6XbBc0O55hU3O+qeaYI86E5ZJvyy0
3tHW0PYU5Fgry3CyOLWf4nEsO7ocqlJpnCAQZG1N72M/o5p1joSgX0p6tb2ieXiPLDy04+kkQ6+o
NhV6dc2lldVYCp2RRkcdfyYSiwjIiHvt6EJkKIMEpm69cSY0bMVjYdHGReI7yXPxEpjzcjMTbsCV
fKSzP8NwnyRCco23FTKZ0udA9zl0I50YaLW2b0CCZQMXf88wS1A0R1YILoU70ReekvXjZh4G3aKA
LPEJJ9gBqFsKG8BHv1nkVFaDsatRGbPXHeiIhY3WHQls375mHk6CHt44RSu8IIEjUtzAEKmqSYVH
eQ+Eztzft/jXVF4cAh3pElbrFYgDaA9oXxipdIDqWmwzZwcXczxMdVtzKjynXTKJ1G8wH4xfxuTl
1yQV8X+8Kjj7mHQpkVn+cATQaqZBsYlWcAY3QjEgH1pvibwwIiVHI+1yKy2Q+XtVsi+KFTwYYIc+
fDZHzeVLZ2RyqLzeGXHlJ2uCMMoVdk6dxB4exyOT45wdRLdYDgGTlr+VICMW9grZqE3CSz12BiBs
3Cgcq1Xi4jZ3eYz79l62urqhPP/mXnzYRinUNQoBkkTycqxtxKGmW8hEXvWxFWTnaFcaN0lqQNWN
mS63SXxaqUyA4Lp4fl4Bqk/RJA+JD0KLs3OlxT1hX7tmPQnUu1YZ5NcfdyK28aAZbg1K7+zoXYu/
38bTLSYkTYJ9J0AdjGWf+qCYBDxYp0qshH5x5YJRT53X/66r27hA3K6bcwFX4KEVvbyFhowh8lKx
N+A1BbOE9uvdio9HeXW+TPc8Sica1VC5Y58acsfFx2a1q4waes6JNC4t0fhumiqOOILjMLklU53x
wLPAbf05g9jYOGxFkAbHWy2c8mdapToR6aqua5SxlLyGH1dbKGgdD7ULjImApB/unCUxnNMljy3k
cNdJGYpWCfeKD6Gyn3L/ilBpvCMLgngkSDU4PRc8AX0/7kWrvQoNCljqZrhrFQmZ4qONMIXINcMp
jUPFPJwwtBkpyaEgF43fxDyEVuVnX+0AfjalSfbYX7/xooyyqoV2Nikopyqs7TMQKVL+XzlILJNV
oacx3DWJ5iHPcuDtScBKIvC2kG4ou69UecXJQ9Zua1oP0tArO9kBvGaoqQnQQK7TCFPWxIiA2f6q
KCXu3+ZRr2zOzqe82ydROuTD5ShVLLEFnL14K7RrplRqgpVfnthFP69CEkau9Ej564QlfqJoUhn6
neAtNtXP2TrWJ3t6rkA9TszY6T7jQPaOmz0cW3iyP6kZ4mZIynu9VtwA8OMd7j0jf94n31dckWQV
E8IUFsSSh/kpFD8kbJXjlwMUQyFYrPGcvCN7zYq4PNWMWQ+6ESQwwtYGVpD/WKwxw92TCBiBkbSB
rNX025EeJRJ0M6Nm5NZVgdUL3A1NHyM/1zVF07dvrC53/+UbMP2AY5D3TP/gJIQZR1FirwC7ILT2
8b1PH+2x3+1cLrvqJnIpIKz3GRERZs/Ahw4/IPTagioGa89zzf1JJSI5DlerGwzUDP6Wyh3kSrSR
hNqTVBEJNBrml5UGk3sprYVEgvkb2sYBTeR75pJk8PAKXQdLHLbnym271qHjtqcJBITVZw+VokWC
gk6ZsE8xbbvt82oH/4zX7f3Y2E4RuotgwLxoHFdt/r7/c5uDkcHDAbMishFZeJvYTfUPEOmKEbyP
4xjQ4K6MigyIkCmuQMM9yJ6OPD6y84BIF+SeSMLpjLUxCoxx2/y79YQcVjG8BoznWOc2xQ4XxBbP
OhPyd6gkg+QJRaz39Kg3X0cvR3Qj26XDkLUANy5xvqihyKCVUkzjfC52+szFUBovx5Cm2qAGTFqs
qCc9pQfh60wqIkhtbNx0Mo6AYAl+MQMGyaT1ycD3EaSstO4NqJJAS9WVsuvpxJEnq2DuVMOhHiFK
rH/6gT0ZXb7DipChwtjqO+QprNHoPrxLL0tKCpNsG0ZR7jVv6As+4r+NUtrbzG+/uZx+uulCkc38
h75FbvG4KBqMlT3CNlM1auQHIghk9CCMdWW4Xo4yt8DdvTkcYJkJZeQDxq/3T55jTIDNNbMGqPdY
P9BXb99TU9rwoYZb73AJcOieGw0tkbMiFpsICgrmsoKfanBlB1M3Hi6BJbF72zKuelEimAwYaZvf
6ily7NjKNOLN2ey9RCW+ag4eo6FYlJJGfyqtIolEGPkxHYtwUP7kUwnGLzCM6IS0dlAN21oMFqf4
LnN29Uv06LurdahJrIRCQZtn3arbmiiBcrOedAphNZEIuy50MP8yyWZAuwTVOW+IBUbCZfGIQKkh
vE7raVJt7FJdzbuvnLV4HyKcJK5XuaFE30lIaZYLCf9cdWo3nR2y4SubHl/dPuFAgINknMisAnGP
Yy/s0JtFGJvXl6/W9mkI4Ahqe4HUEQIBq8vDS3b2SXCqhFqT3PR+8eEGM1M6o2lcFuxjrHLVlXJe
Bip8wDTSsQyDwjipzXpDoIQAZp/UNvd0xxFVAuw2IqGGl3COGJZu+SrUxzZ2mEnC0MBvEMRk1Zuq
14p3jzeh692lknCuQqccuh2Fs3y7fgy8QmKqJzTg44MwguDf9uBLyzObn04j+H/ZEe9DwpSOSLtR
LtrKUxSEfaUa+YQMZ713qoh77nAJao12Xj1tkZm0LCA1tF9lJjVHnzyqc7hampiRSJILN8+DkrSE
AAulv3qQs/pEMmWahGybQoBfNG/DXpp1FdN6UEQZu1f8UQFUFtt57Nr3c2btEHm0g24DozDf8Xpe
NX/l/MarsgO8up0Fo7XOEd5EmjcXY77AzQFLipX8QTkXmq9zBFtL+/plRInkG8wyGNuErwl80+KY
1meviUp0+8tdoeqejFw2w2CLlIay65R4KU1RdIFNzFmAydqVzAKqgqK03pWZD4cZkGPd6RVDBaKf
PPUe16u+4E69wV6UOfrlfOCV9lalSRVc2QX8Nmr1X6XhoMW9jvfLoWRSce5I/P8R59mNm3wHwG9e
GQ4esV790DWY0xLPs3Jl5bPMLapSh0Ygh50D46zXx00bnvfNxGJa66KvNCfan3RwGCF1a8t64nYo
VepgjxevD9tcmQ/yX6DU/WaDTb/AgkQignwiXudV+r+5X/FW2XLtRRA9Zcfv8kt0seEICd8Np7/E
TqudrlSZr/AqnNaCFsNhgAYZUm7zdLOd2quGrS0eUk0+lfleVi8uutqk1KJrWKindjF1bXfjdKTv
owmpn6jJvJcN2gXy1EP9GyrnGxcTjeXJMl6u7Ic47VKLGAlFC+JMUaagY6YlcWXT1gKbN5yhVQ4c
kGJSO01MQgPWRNCC5fWbeRhzDfyTg7Q461rntW3/3M6kp++HALaPurgMqON/GfQSUoRd8MFGqO8y
4EP5Q8hbJND+tck8s3wrv0SSiDkVGI/i0WsMTzRnjghxyAV/tLxUtmpXoTzOfqeuSGO/4HIWDD4u
lOF6zgCt1S1dotzQt1sD/vTxg01SMi5/0CcGkzYco6JctXFG+Bv3/D2SMSbMNVUHJyd006qZBwBi
M4oj3KYD7C1s4CS5NnJ3i2rg4R+9LGagoLm9zjo/dh5Toq/q8jV+R7OJkZIDVWcUyVElmcmDgzL3
6te87noAjVyZt3cfaNDiQp5k7dDsFpdLD+xd0ijxfB1kPhfMyt89drIJUPCbaPhlLFyL9ZAR0lAP
JgMSRaK92k2Kp7vTTacavWh6QJR+LV5Osoap0DVB9vO27sYj1C3Q3XUZujfrUyQEqPRTCPoq1QxW
Hb8T4aliEt5mStFilF5m2iFXpWaJzhLEQzIfPxNoGaQiGxlsRe7QV27jtYwbWHQRHn1s6ze0iwcC
I+caxpDgPWrjXcggWVi68Jpa4ZDZI0oE5NOsL6ABz2WwDz+GXNPyXoVD+Z8slviTSV93pnCYhnq+
VvfF8oA7Znc+pBySEsns8yRY3oAw16ot6wYAbh7xcD4T5y+Z9M7fiKm3GHKSum68k22FQ5k29d76
dF9gOVN5X8jD1NVQbSZFia9GALV0ARBSWnExlwNcOZ4whHSMv5GnrZ96RuQ1lHJWcExwERzYwcJB
F0Bc31RH1CMFikxoXdagUO+I82eFfAvtHnHi3SG4m5ejSADCZ08VlRm9qUi7hOEJH+JIKK/Vic7o
1HCBhKhiTB5nE/w+aSo3CudH+8KHBg7IiEjqevRvQAKZGcMxTxLTg8xCahzXuJ7fG+OGVkudMBV3
NXXM5UuRaFi/AZZyEJ1eadNYQRMaADtYDpilY9Dxn1Ph4lyRVSoeisVzmwU2S+mrAW/KFjEWsmU+
jDb/m4me4kMzxH8Naf5lgJoQNMpOikZLQFeJFyik4T9byO48bQisFAQwL2O0FpfS3HzIfd1rqomy
fANcMvU8beaScH+VmkelGgY3ktQ2u1HzskSf/g0mQgxVSkCHwV+5TjUaG4GWCJvnOd9OhHQpG9e6
eg7SSqoY3rMKZV7tIGXgzQWSvIiNHulyY+xF/niWT6iPtuYYNVULUM3ZXTdKOKjKp3VftJh1IxeE
TvbgfaglCwWd7Lhp0nF2GHo34cEiC+uW/8jOOP2iznHE/4cj3I0+fY3dr5HWIiOqROimq6yriZ4b
FROjMjP0tbqsnvkYk3/gqU3wrPkwb25CJp9iw5pQMGrjqULSVrvvAK9tArlLfoU+p+qAF3Af9Q1W
6Fngi3N569NKzyvrmT4iXye2j6f/uKHhN1VUP/O5mfbcdFNi0IpwihZ675KZUQKnTN3fP2EBFYab
S6Lfeygg6cUuktvhbkSrsNsIVoWHisR4tyhQoVeMcAhg37WpxwNdGEieNxNG8bz8dqywtvXb8ioG
R1n4gmaUNT+yWhZgWI7BpRD/GYJ+JRJioKrTulTogEM79eMviyO8qOffVqqO0q3AmaC+XfsiKdzi
9w1pTnS7+vypyYMLS9rLZ+51E/9QMu5jbXWH2npweJCNeb+2NmVqGUEJzSU87CD8PnC22CMsWuQL
2Uf9Nq7hTxOUQm/0mdMmlWEjDiKTHuKFToGB7fHfKA3VKC0XazOSsG6APgYbuGXX1WjpdaV8rOG5
9Oy5r1DtwLh7A7cifaP4EaPFeX2kqExbH27pPj7z2HxofxCozVDdFT719yRK2LLHIM2SDO8CHGLn
PmJVWusMvLszPHu2prusIeaucC7nb40QT4rVQ4q1y2SY/4GWca1Ap1i0Yc1wnXjCIoT4hPEaq+MB
zBW8o1aujY3W2XxosxEF7n4xE5YVhS/WnD+p4g3Bb5zhfuk0kVZYpIkgNm5MZ+JFE2JSh11lswGo
+XSG6ft0q/nF7IEaC/G9epFLi6bp5TeOnyL6uOAEnKz5FmZ0WOYuDC5tvcuYHE7vNxzQlXME87ae
wi7TzPx4YMJ5CwPwbEwVxKqzgSTgKyN5Ga2AUNcWDX9PVOK3hjXDwP4nPr4Gjo4fBDkVMibof4S1
Fnz306UjM+Wl8vQILrXUVpXXt16LB+OoBYxBn1SwGASbUGyTwtrXlTq/NK4mDz4JwbW0mdIPhYHQ
S9bdAo2C4X86mFqUG3/ckoef/a7spAXkiAurrvIwbGYXpQM19VfN+AWNq8i3TOxM9wJ+146bZ2eb
Qz6UBFus2vMViS8mRAli1DcX81Q1xvw/eOr+jzlcI6XIF4fWUfSd0F3f2lcNcSxxz6Kah3TJ+fxq
7C72kY/7c8pjgYY3j4se5+Eqw4p9RmcXEW7/Wx6rBN7lDZ/mwRe383GH08x84ySIl5ArjPOvJ0eC
piVDFqRP+giXieTfHg68IMmzwwbXE1WHKrPOUY1JFTKcR6ygVPdMmefK/qeSy3+J1aCN7FpFSGCg
mF8qJrXXQZEE/kDh0QNZBIzZKYvGJI4q67yeGHPa+VskSs3SDoir2H24BoAgiYulVEfszUiqZqVL
Zeb4OeSDwNcUO6NFCmGCV+f3ylmL828p9k8XNs1dh2jWLBoVSx5WBwTY8SWmbFCE1bs+leDowrnh
4/W4TeK/Xka87N2tx0QkC4Tr+8cXkPPHsgHlZUeJn2JWglVPR5m6Oc5bIRf5/53ZXcWZsnKSnp3c
rwqLjvMjvn3Wi3oMaBIdQ9vDd98+9CFUb0QZkPZMRHAHmTw3V6YTbVJAmCe8EGqB1RpJtzBDViBk
HyRQJUsEKJAN13hafFLlmnQ4bxop5XgkSOMq1gDQVMJbKM2OSGinMDp73H9Am9OZ/NSU2Z9n05KV
/9FwQ9pLmXqYDWTLjY1JDoDrEwj3JmUktJBqGaBDt1ktSkq/uvem3+eiJGBQNt+a21/MZpsUZmOi
n5b2ZT4bH2TdcY4/+tORXIFnf1kZLDdy+b+xxxMFavVwhcVYx7nbg9kumTZJU8HoGeV3ZB37m6le
FgomZxhWxMr/eRteM9X8TkoUt09RaQaRkM2SCiYkN7PAGE4WqNCzLZR+/rif6ZqwXQpSnCdI8U4X
7KIidYh3K6HoR3v3qaJ4dCuMxDwxD+CgluFiY74Mmt8Lp/fo3DEYwQhJNxcb66iUez5+X85+Llzw
rZZTUr/xL/Ghe5vqDstc9h7hYSHVTXEtpl8zTl3QjcB6yWrf+kNZbsmGSgkfiqmCuVV+XmzkEL8r
1XkaSaAEoXmw0qB2zAxTxITqmnctS1IiIo5Lj86VQ4rL4pzBaOdxIQ7UBIGUOxAMId8SRVHCcdHd
uUN+ray1q9TY8Ec2KlgH1UZXRIaEX6KPtQ94Kan+cuDHqIXotgsGXK4i9Q6MZ32n9ZjC6PJtxenm
VqX7Jw9dzy7Gv8qVNZVFg57s9dM+FjtqYaynrebcFPvKBzSkEaqVmOpAysOvfDQZHrvu7JEttOve
TJXl/wgnLAjHDRlYR8mlwkHzq87z1OcoPr9IwHt6kElXUY2bNQhhLRWqDJ0WCPnZCVBTwxtn6mLd
CYJA7FgSDRubzbWBZxG2bCCuQU9/m0nu9boc+VkMBV76uHAGONyLjgdqDZ3Kfsj5/yvWF9l4vHel
4fNV+DjktqNVLv2glCthG0vhDpgRlTjncwj0JzamikEG2py6H683JLKlmEs3eH0eBelmWbOIlBWo
T+fGSKNkVQOV2rGoy62Y4SHTsrKa272PEScPc+bsCoikDKwsNEpDXW8mi+diQ7f7DSvOIwWWMD6P
iGCXo7oMFkOPqzp2Cbq/CnXJZPmnIo6i+CZqQ+GSNUkz0+1BHF3Zc/gXCH8ASG0eU7zVkWVXgo+u
Yhzb8VtcHrTZrIBhBOPcnCsHPGUafF6Qlnw5F58obiwebzlZtMxSd4mKyN8J6H2duXXM6lyK73Hu
/mWjnmUIk/lH7gPPn3tEdOSr491A+SmjqY+01OA0KF7teRVyzTlS50Kd+GvaqN0txpVKswiqjg9S
wHLh/z4gAsn2wX+pQfyGrrgtNvV6Pla3QAlgqJONBxSEwykFmjpQiDGJZQz7ChDjxkTDzC1++0jf
ZyZ7pLKQgpZpoDN55y0XWj0IWfoUbHkqLVE+v7p21Z4KcxPsuYGlsfzw5IoHli23WUwJfUwPplec
UtdHHRPJBjQeuXrUq3xPcFzb3m0ElBRTJ6cY1K8gN1ZzQ+mIWMzC46MXMpUB0bM6f9WbHARtjQZj
D5rrHqHtgPhkSV4+lHohvLAeEPeLur4YTChaeWrqUdFKBiJVOKMeSL0r+jrICkB2HWtbme6AY7zj
vId5VkigciN25k29J4DGGSX6HZ4G/H8aOEHzaPCIbcOIJQc1Jxc8c7ksdkX0PtZ4vsJkLN01vFh9
2fD3uaNcxivhbytIhJKgD/c0uRLkbD+2K4wjWL5Zc3b5kaTLT9mI+3ojxpkMUPk+sFzt001c0ekM
ntaaY9+wBykzovkQUwy0yhjKFxvB9sONTTdOuUc2sIqqIB9cUmnAZWV/yQGtE6JXAYjveOr+0ZJF
ISOArRhIuNoXeozfuoj/Am7LGSNgHS7tgixIcHEWgpasEz/slcVZGbQDlBdpa6Adg4R2cuiVi+zC
DFKg11gwOrQKrAqdTqvjfHFe48pRqsBA9VAoXjStGmrMe24tYrHbea8oX5sYcd7CRCQEBD4eT80a
IhMBOpJPLE1T31WHM2sqeEBwtcX17QMU/E5SIgNgzEtrd4Aq4rAJSO/3b85XfDljpXWOOVxiszFr
RpHw5whC5ZSZABT6B7kW/hPpmc8Aq8XVgA79pncKAYEaSVnNqrk+0TdTwyKnEfGfcrmfBHm+Sod8
O1TwJG8eSKLCItQUMHvLdANLLj1Vi1xDsgsVfVXb5Jz4LY46/jBB9foNRCOhgn5/KwuOeBwENyxU
HcZVctRa4tEy900PJgm/cDXBAt9wNusOT1g1BGPgiajBKwsFpUeXcQmyw4cJJ4yeB+WmK1wmtypa
9s7YZkq260/VFxiSn3uPA5uwIIzikqiOD1wMadMwYvkhRe1y4BDtTkr0sSaO++PxaF7Lo+DN4kbF
boLg0F4xKAoze+MhBGdjk9oykZixK6CJ5OgbH3oZJ1ORjxgCCNbW31M6Y9/BcH+u0R7a+yVgi49/
glaTYYEca71Q84nJnoGnENhBUyYPpt4ycly853D9MrURVcqgB+YOPNT0Z2PrrsN2jqefBFEFe+VN
iuF5qtYgtqRVUPxGkMXyyNFKPLgHu52bPUovA44OGz2uYhXfJ/ZJB3kPeMTtsDRknlHcD3EDaW7/
cs9z9wiZa5bRiAZ2JeFK255mCCZNlYR2P8lilMphNj7aT9iEuP+/oB4o3zvAAvhuAyjdDn0SwCLB
+OfYd2FiuSDovHCvsZnBcfkvpBi0SmQKZvO5qXnrh+78TKM2Q/Un0hjmDnI+CFtQ8GulnzMSMjeZ
Zp+idvkjjG2jQmVK9D01KX5pLxEhxJSod3C6Yjqm+sdLqbRN0XdT1pn2O45RCC5Kz+Q/yAaCwaIZ
/0xVrzHkGlRu6T34QzsL5CK1ujxUTycaciNMIF5JORCh5vtM8wVDpFvy6xcDoe+UWkO3i2qiPuCK
5kQ8VEoNx148EFtWoyQiFXm58dbRv/lr/5O4GIZvAWUl6QxzpXWnSo47FcLfpcL6dqdm4hWmiF3k
16Pr1z4LU07iEojgFkBvgqIwIJI81b4YvtSPmTXlNvNbIfpj8r66oBMOQg6pGEDaej4Z820ZrByZ
KpGvPvlfFqKS59xbVywV5vJsBu8RJuz54B01JOxe6tGHRF4KZhACINM282mepjYvIvYmH1gPlKFk
+arQGDE5Q2yqgOwT5QaSte16ti1FmV0bcfhdx/s3ZbUvWYqAUAFy5j4CBFN1YHjqp4+d9Hkk9mDl
Si4THDg7zMROBJ9zGPt+8V7cupSsh4kpAcmJuVaxh9KjxIJmLzELbJueVvkYio5pb1kKRjrnu9kO
nLXyt5BRf48pd2XJ81ky1w64ok/K3oeNoBES7N8+JwSlQ5cbuyIPlLgudjMNiJTt7E0kAMp8F7i6
8QgGfs0ogzZxwsWobI+v2+O8G3nO393HN3Hue+8c2bQwNXuBWFmiUvFudMLtTY+K4/yYrexi1IdK
xyV3n+LmtryipfrCqEYyA4YmDeXu5XBZ7LQWAmkoL9+sQIfthCexWVi9RF2Mo86aSK186+dsVW+C
ey8RWlW6AJArktjka+kx51p+kdgmq43sagl+s6HsKM3qlhwZzaf6+iJ3B8nhmuT8DZYOhChTim2u
khQ5zifeOFb/JGvaX8hmXRhSDPPYrOqoTHeHC56l0ZrFsUY7cC4hnKMxMtYwYGwLHv669lh5a7YW
XOdN2tykCSkMElxvb093kqDOVz7pqY6azRpQWg6UbSctupQHSow3eo1wdpQsTNbOAa4mhG6S3/UH
9TgXp5fVJ5RW1YRqMSPvEqVOM41DnQIhZQiIaPVZDt8rom9MWb/ffAuZh+MSTut76SJkLrX7uVuI
tUtPcu7Ql7qxcwtEvgwoZYLaGJNk8H8OX1UhXr6Qu4wY6SzMGifFpg4E5EL0FzDNtvysjAsvDeMu
4L/KzmByyDkNL9bIVGZKc+Zx4lMxMxrK71vv3/P8+gVWwZxggt4AnQsx4xtUZ5O+wtiUH48l9cwf
z/JpgTttw89Z/bWdkX9EWl9iOgj7SsnH830d6dKhWAazvd1eLCCIwGW4ypp5yfyd+NNpMUnN2caM
fpanY+0s1xrm/mRwW/hNXSWTmUChaUvCpnA9Pk8nTHXN1y7sMBCcF6L25gvueE4grYzShLTRcvIU
j1A/fyTyR1PBEVkh5dTqic/OERh/Oy2EV90huUU66yYqdsw4fVWUlE5KWvy3tm1SoqUZmuNWDtkc
y7HBDRz6+7ZML9oVDpJnOFwHVUsb03hHwOaOHCwJ0FXo4Vam1b+SqKISQH4grKY1hVBh+izZMVfi
fMWW4l/8gzxfDTbKrN/ZcicPbSU7jvOPWaQiOyduKw/j5bNpo2iwDk5cc9Np1727JDTmojBC9rHc
coOcyV3nxKanIBeiNkE/LZjSOCPg47g8bx11ilCaAPz9sd2GCZyuo75siQZO4MhE8fMfdeQ8LSr5
I0jOAOi2/RvBFiwIcwckVFHI4POACmj1a+5AtXk/ChkaxXKNMsREoAe+Liyq1vglWjJtmS3DxzL2
3aB7njFemvKDEGClO7Wkf2hk2js40X/Y1Fj+fUPO6sNd+WRiEj/z5SxRVFq7CkOswRv5khGsSGtc
e95tLl8tmVNjRSWP+1n8b3qUkBnl/ek+aVTBe9M7L5C1kItXneu1x0jCIgMUw0hwBuDmtyNAngTm
3zMWjOCATE1d1tSFwXXYyBrNcbR5qr2bboAFQlh1N4Y7vu7dpUiPdICbLhzaPWmvqtTvcJ1rtngB
KXtaFeLBiAy2Qrt07P5WEgH1MYKTsejCwNDdlagKue2ijI2eMkEQH7HxJsuShs1Vs95kjZ9FoUcA
L1hfkwCDbDgNCT+wURNp3Y+FdnjQwCvIm7o0IwmjIzr+SiuUMqaQpU9JYoQGiWKP8S+iDsb5zIJY
3OfSRaGKfSQVt4ZrqttPVkvkgihZIx6ooNORrTOpJkbcRA6rQbayoGOO63YMpgiypZoT7hB0GaRu
3OYsdDVOmpQTS7VBwj7FQ3ptDWV9uirq03UUYeSc7DHd+zswnJS2KsWY0v/xp/AFOkeGm7TgRBSm
LDqG8HHCLhj9bwH+4CWjlkQPLeD6bXEEmpcCgznPB+A5YJjcEMlB9shekg9KdtLmnkoCVvRzH4F9
OJaPqShr1YP26w9LRg9UDz0YXTm7w4IZPBPyc3ATIz26vKZRmvohdLtq5NDrrLDm90ZUA5xKqkxm
LNcz5HIl3EEMSRyzAH4GenbK9yMen0xlGWCbdcfDCf6kAaot5ZYrS2zAhXx3OROWEQgCtqMLTtIy
gnRcGTfpUM5dDPRZrcqdvlkipk8slYnishwu4YElB9ZCTTQ6NNs+L3PWCJU8js6yPVNxJc+syh0i
pi5Gc2PxBe7maQX4o7V5Mj/0gGbFzz4WRzGAzStpY+7woMy4mVbqlt++YK88m33LhkMtdBbTkDRV
2H3+cK7u1/jrShozpt7iCF7hZReAYF+MfbIyeE+NxzGcsKkiOSOWTYsichK1z2HR6OHsB5si1BS3
NgT1RF/1qP05fP5fVIaULDwKokr2hzRG7GGxSqQCUsZb9VsYoTHGUp9Co8rIDpAm4fwu1iDC5p6H
qEy2k1Vk/GQBS+Cie+V/cE0NHt1c8oh4DoJwSTTWTlY6WEEgi7JKEsddhQdBiyori7KRefinSnVR
T+RvT3Tfa224jFvqdfdTDhnpkWyfu14LQIVT3Ukdy3jrnV5pjmU45Nj21nljX1twm79UXtNwd73P
sQHCMo8t1cXKsMXxmAch3mWEBs4j4omYdXjQvRvA0e/fVK/ffvc9uF4ogYpJh8wpRb9PEMqiYPlS
NluauWR2cyrODCi3ySnHPpPcJGd6o4bA+z77puAK1vObFpqXSC6xXL9kWcpLoKgL71Sk2PaehMwe
nvggo+RViXdCDiqWgA/4L8DRlgyaLGMKPMJR57l/ZCZ1/PjD21tKWsmrJl5OJvVWinDl3N2+cRSk
PFth0jpb/QFBkX6UvSjs80tLBgoS/En3M856VJw5iAk76eYuzyAYFC+JCp7Ny7WqZEbYXCPJELIZ
hrkXww0RGAf02capSq5n3KO7P8zunQbW1Ud7bOBV89/4tPR7yK363N+lYT5cooLbFSCGXZiDYlbP
65SIiUlmSeSGYPd7Qwpi5hMWG+PnSmGsWJy/qWixmgY8nF/ZI/FFMT9Mr5ADZb1D0nVxL2bKXECY
Sg215gaXNqvek+YQGkk3ICL2WvDQsY0htb0vUN02tURHAkLwUcKQjya61ziUpbowdnXVp9Hr4BjQ
ax5MmTyCdV0CjoOPV9/4qkkjuHD3VDg0ZMit11CLeS6cFbXV6AldZlQon2yNKkxKsuxyMNAUF2F9
fG9HT8UgWnjptC82Vb5iMtMMdTZaRa5YLQh61+eP84UEUx1lRApyxB5ucApYehiDBc04GoM1AcC2
3og10DiUQg6PwJsgrHihnKSg4QyJKjEyg386Gxv7myTJN+LRMwnKFR7z2SriPNSTZovEOvXF9zT6
8eT5q4mdEI+P6buNm/YfCMdIjxA7XiV4RvPSgn+dzU1IgzI8bxanISEf988qZeEGfbd2M4sTEGFI
EET6c8W9z4qjQzUh4KRujGgA0vf5fAbC/h5HSDCTHjec/kuIs2TFtqHJr+GgsFT9gpSY2jTzR7DP
hpUId1/pyaSVnr0D7g0iwXZWScnnHuA4mLa9RL2S/r/I4BneL3Oq+IJzMARfT9GMwsSUlcA7XORK
OFqS5tNs35s3tUPMkbDnc2aNVFbmdGQhaHksNZr7xmUCVqLH2MnZ9wZWtGrb00wDPKBXkZ7kVw3u
l6dLHh9lDk3B8KHLyvS5inUHN7v3ZJZeqTQ0vbZV/t/fWr1dJzj6V4p9ok1nY5uu2xAO3ma4KpER
OdkTydX7AWdPdaZrP9ynOnY0PNoIqZzVGd7cFBMHKoKFa0x7/aLmFQdOvjpan2vcYdxIKXu1OS6o
KFRCYMLwac/ZvzxsM8ikDY9TgWiA9KLGsxPOwgz1CJAqDfbULEnudpplh44Fni2VToAUu70Ju0r1
hd88qz60KkK099h9jPFMqytZ1nTdQanNFF4XSXBhlGHKGnygZm1v4dTHU7YcUEsKn1h/JWFKN9uV
Dd4dVFiRUPoJ2K057EcbAF3wnJ9vrtf1r19u2i4cb/yZKIHHSOdngee01jaUorqGcxpWojV4uCuN
NJKhLELqLKODAW0UMPBTWPqU4hB4/n2ngXqwhkUoJPBmktXI9XK3em0UI+aZzTLY744hTjMphang
pvbHwVotGB8hprcECF+WnFD8tzf3zXLsvVddSJSQZBmqzGuIMujtg/BZyFHLpET5lYR250IVXd3l
fHOXICoxjiZ21A9txSJiu9nS9+I807QqvQoUqtdH4wegntL8UVViYM071glelpKT37R7AOm0D7cT
uMUgx2mxjhGNKVADYE9UN55UQjlDkHEVOUs2iqpLbxcQ6j04o+Qe7RvcPnlWWRSGwVbCqVTDMDa2
8cJysKJyaNlw9NobqCI9RMHMhes5ISw/8K5HNTv+hUYF3KTa+jUh5ml8TagLojR52iQNem8vqZrx
vAJBZFaJJWCT4dSPaHOAKAAIOY9IizXdEPp7qPpgJ7OhOFUq2Ldb2xcYf3TlJ6w7Yn4KH6npbx0W
FDq8QOdx2SHZg6lENuu889H9vFag4zVr0zxJSH0d53Rr7VREVlIwqPQ7WjUeyvRDWzlFPl5afzze
dYgl2/iCRV+7BgdoKPhPJeQQRX/Tah6g6ZFlAGttt8L1nVciugPfhYrUGlIS2fxbUa7WPtxqVSx5
gC2xfmToFbNgCTlm9vpe1utLYFbExiMz7qNnsJDlsWLskZSinCVXHXbeRTwny1XBkAMm+KWCICUY
4bjtjfMiqv+xu8vNr6L71kpYO6uQZLW87NiNPJXOOcsZVWniPagt4O1MHYEYLAgXdlR8d118Qj8M
1Gs1yLqMm04vN/meLSHmubnbO8BngYHtdH7bZ1P+rKBdHYyQMbsdtFhjlstY5nfhPaFGoOq4MK7t
kOSnaI2KkYq4FVzHkR33mbYTvtWkKDRY0EJYHmOF6BYjvlgbnkwvd4QYevRQREsdwCKOYEdHsVbj
k+T28ZqrGf0+fapASaiiP2CcX26/igBsYNlVfjJbTQ9gi9+2SsKFmdpYFp9+e0jhI25IDWMT7C4Z
cHnlWJv0zEjdx+SJIbSm9sk9gmAnErlDVJtXx4nPgbPpRaFKQ20vRPBlfT+FtmQOR6Dr+SVjJsGc
qaI2N6Ya6Afir2PREn4LOcxve9wCBaHbkrM41w2q/iBsJp9UIgz5b8C8OgfapnyFoIAxd9Vi+DmA
iggUPZ4jG1XUjE+zhEID7zSVcmzziq/zpsumN69ejAS4+BfgpSCMOsg/8eEgOkn0uTU/DpHOPhw/
zJ0RLSnAqtsAMVJcAKjCm9b/U29vmzZV8BvD9QcbZr79cs6wqRaHyIEvV05MPI4OZCBwubFPR3Xo
Vl0JoyRUPMEVmMwvH2JbVC3Bov5ZGcGIf1+8ZmxeTWIfOIJC4VVoPP1hExyVu6V/jmC5r3n4we9o
ibVGtem+mbMxXwwlKObDUz7CzWCaCEz9bf7azR9NfXUk6X8AUuQ8ts8UlTvOEDtgvNsZ6vCJfohW
i9266unxDznCIbNMfQeIVXFmHmKZOJDnx0VRrYLP/6bzNqokVQom3ppN7/QnyGkjuEqIFDaSi5oB
kAfr4dArzOKdCp957hMeprLuLafolsQ/7Bgk9k0nKsz3FDGe9cCIuJrejOvGFNfVeeBw4hZd/TI6
tD5w4MuVTnTzE5n1akBssjrdlU5qTbavcnmRddj9Z17csR3YgJxbEUJguacFmqyNfLiBtILKRMe3
gGeCDqBP/BvNoIk4ayCuWmIvTtw7/SHDyv/ElUblBM3gTLX96odoYD+xCEaXiUmmtEZKpfFy5KAU
jxRb2574ZLG4P7PawmZGEro2rYRisdm3vgFRFWNXjNyiFsKzeOZ+7+GI4sJh1vJbwi/ql6d+9vP0
/I2Z5DwXy+hr3wG4omqpedqs331e1ELMeB0yBH616ZlX2n8mGFnZw5IQjKASKfzlquQPu0dJ3X/S
DkRDEBghHNreSD+CIWsrQnMnG39sTGQa4aBwQUxiqqFoYWCi566sT/Soyf8pZUVYwj3QAsciswBn
ZF4bshv8czazrwbP/vb2TrSd9mojL+4cB5qI9fQQdp//QVyShjseqW79Yw95St7OAOVfH6xuG0bw
bCEpNiN+QHPrSzCJjhsc7hk+oQ2ocklsGCDhyjeC6bQ/scbyffw71xX378/kFxvfh9D86tB+YTAs
x7GHzt5EJqTWUpV+KZ+O1jNRttkPntV5vk8cl5fUxQ8fLPHJUAVsbSjkghsq8uti8t/GfrHg5p0O
Vik61W6CdUASqShYpUlVwzoajEbP8bwfHrLk1ZSTjDImHAEnJ4g1vPHVcqmVYdjOsLRnu5x4YUNw
JRj32Pu2myRFDS4Vs3A+OO3557jtBOlJN+l85RvkozgcFG3woWZEWTDeYxYX2k940oVxAoo+AMv+
XpZ1OocKDzxjfwvfISpjiCXUYhwFOqqNLP/zmohgW/mnuL/Leedur72boNcEG7eZA/b2YAhsbs1y
TnAoN9zHYTh8o3Ud9M3K1TXoxwLM/iUhjXqMxxathFag0wlTzHqgLlzCOhI5u2mA5y0/uM15kUGD
OgibA0lzdZHG+c4CZp4ZpxKtQjTjZumvBKlw4K31Ml/6viu12S29eakYe6LO3FF47+l3XqBGf1Ah
G907Vo9bM/YzRI8GhiLMqXAPlOwMD/gmJVCrBwkPfHPU3CRNOMZv/4rVWk6IFWx3OSpBnujmWSMC
DnfXC+YxnXiDzjCqp3frZYuvdA6iKfsCLDjaf5oKhTdlyViPMFyzXRGJ72ZNbhwVVxmL6HmCkxvd
KPZY47JzyB6BcCAA7W10IZTDZdvniA/29lcxn3SneWlp9GiGVEnwKvqocE4RUUEIaQCHLgJ3aNdw
We2PVhWPfVvcS8Zeo/m+F6j8RX0PJu1S9cQoEqb0zV8SO+3s7RPjZneVQGlZ8weXrtvlGNxGOTO6
Yuv2PGXqgC0AeroPTh98wQWQCmZEOD3sj8H3wArRolYqbFO9Pi5MDMo4rUedyTLUvwWAMomVKmm4
3tENMqFLsSAG6x0Qt+zCJWXByK26VnN9l+qF60JUCaBBBJR+GVz8MMn7yhQrGhxrpYZZsRnm3oqx
cE1Mgn8N1mxEG8Y4U939eHN40pcLK14rXhJL/pcqiP5unPoQ8EJh6d0dMFqQsTUUcOIVYjCvS12b
Q/CqZxpZctgY1goxDHTxkKuMgGgj7K4uS+YuiO5Fr/ni0GTUzWQS0izzAH7fjznlkeOjTGh0YxhS
vf6lN6sKQFMCbZyNGUJazY1FSjZzSBBJeEaOL/BPivjxBgLyEr72w21JhNOMIR+3BTutfFu9g4W7
WCacMC7T4F1egiicGMJtKTM76HTq1+5SDZr1LVJQCAo5JoDwLIrSd54fIVRyRJ1uAFKqDqn+rS2W
qQuV1+pn/ZeE0e0k4a/Kng5sQIt3wNS3LDwVJYfrD9KitFzn6z1VWKlcNONOV95OkP1C/3fBG9HW
a8ovL9tP3VCzfJJSRvV9ny+c9a9Ul9EokhyriSCWs5kEqfcEiY7acFUHoHODfXW+ZGE/WZnYWE7l
7a/ZRm5aFIOkgDe6Y2PtOuU0+e31/13RjuBxGj2SfqMEB7ArxMvgB9WZb1hZtlYj6QPBU2aLyKV+
n/eSJQ3f15FDDgyQOK94fbkv4GpB1GqR1qqt/Uyfxu9yzb+E1EqF0KS5VoYkAc2O5CTDxJr/twpX
gmArgCG3qtrwJxJO/1LnZcHymIOCoXceNsd6wnRh24i81g4AZjfgADx4sAkKxMdFhTvlBZslpdCj
CzWbi4A835JivLVxeAqbnsWChrnjVEwUOps2jRYARAkW3TuqsYq5QLhcG2N2h/8+JVoJ7sNnIL2Z
yIFAWebS7I5kfzy2JgY46Uv7M9uoovmmUwj6AEMZwppFMfvS3i2L/hQSDUJxb8zOA+iC7XjInx0F
eV+3JipAjLnpjxc+tkDKnJO7UykHYiNHif4jKkxCcGY1aOgeFCFB3Ay/zqjUHLxKX+OlSOL13xh8
A6TcgjJJOzip2GXRSOx84JYpJZVMMVyVqrZXwuU/OM/VOBVxjQy78SYIGb9pvfmDGg1syU7xCi4M
zQUAVs/VawDQOTvzb+3GcA27dXNSuvqpZLMEkRc/ob4xnaxhpznNGJ1XqzuAb32tIlyGu4e5hnKt
Lh/Or0+/jUkth5WCG3o4INmbXreBsYP3mSYgaz+4zS5RGgQh4FgBqFlXSmvG5FyjRlLpwVav6nxX
euWTcWpxi2iFPTkM83qcpotRqHpt3RCCd8bGrKPjNk0xm38GH0a75oPfZjiz0LV+efVQjYtbzPUF
xt70vEZ8k8TMzTtgxxdrwOiqc4sh53kofHbjaK1E/hZ0QmrBTWim56XXq/dOecAFgZKPJr3uHVY3
QzGU/Y1YQzsC7xbfbnDD2OaETL6T50C7gTCeaBbjSf4Q5ATNO9GFX7OnQxYItqdK1rGqVKJYmAYU
a1RV3iCSgvvjkDkZTWfdpQtJ3pKgSzL66Z7bQt05lzgELohWlqmGg0m3w5eyb7YSCSTQqXUVxOOs
BhPMGabAM465j36R7OjaJfltcSrX6c9hYvhOzhkd1XrjhvqOwLu4Oc/B4VOnimv5iggOVnQxuNYh
QFgckVH6GLDbLo9jLAaqnU2ycDuuEv4Bi0FDLf9GFuJ6GJixPfDUvpblswveov39oFgKRmSpLtCM
QVJ1/wFp1Ldgrjrigh1vymt4YA0LfHld4eWDIGRHSZFcSgDCnxW1Y+lOrsb5ZrebqADDM04ZL9VH
pTwVbnYx9d6eECyTPaepJfiu7mkwNcNG8WaV/lL9O1pGPhkYlMW7pHmgspPbMUk5pNwFmXPlgn21
IPjnlOzR2JaTfpeWdD650rXgrkUb56uMjfSe85eJ9xs6wAaGRLo6gPaz8GThRgptltd5ZLa1DN8/
W3uxNWtgk8ywoSLOr+KBwniguzcUnpBRi85od1ijyn9xvf4p6PQp1gHRHO6iwE5TiL579etFsHFv
n/ZBK5PHLWgJUiYuX2H5KHdXEoUg6yT6ei/b3uw4ISF09D4JK0OsAEchRpNh98oY79RulIAm1raO
XxD0maF6BupL4fIq23H7oX/fIbjCEw9GANIV2W6l5WW0DTtybPk2/HlP+Sss2kI+TYBrh0e2Ac2l
AzS3LfAE0Ykd0MOCFdwxp3vYAVG7yuuveQlubvwQUxkSldRTLFX246062+UYhY7J97t3+71t1Leo
8KbxaByZ2LRY2gNqnprusXqw3pN1IvpgHx397n8ssV6lx5KqIAaamkHfSK+dgYr84VYd7+ClPaeg
RdUqOv9cfdZDYjryIgfOjnfsEp9Ek1g7uTDg5jUT4n3Cz7m4qPDeZNsTyFkrm1UEI1T2qylQ4LKk
ptncDcGq7BE1YYEW25OgHkayFzo5TcIFr2dLNtM+NTDWRFbBcusF3SQVi6XBXHOGYZHT6MNCIG8a
FmmmMtESLUKHgGDe4q/0WxSEZaRGbgDCD+RzUGj4H50SlGFps66460ouVJM0O3wfbGbs5iHfvg6i
lzSXR6oMIU9M9HgHK8YYUaROIBN/UCQ3BI59zCWW0Q3a32bwX68T13jk3H2PvtgZJjQJEUj59fMG
BqY8HR0wBvIZj55NR3L7l/09H/OvaU1cwUnjuKtc5yzmmVF2pwby2b9Xo37cZPdgAcaBA0A9axe7
Mx5BHrqR0l70buEA43q3PxqtTH6n8idKRZO4a74ez2dHElCWAAlJzwpDyhf0Zx2IGV7JmXY6e/D7
wPfKgItwvnOrMC7wgrOqIxdSPA/Wa5WN75XNOxlyjPatAh+0drsmT4jQWAPBlJ8+m11+RiTvIqxf
qQlkZ5YP0oxf9R0bGNz+spempeoFQMFEVI/r/BprxxuG56aH+e8KcN3Zx2R218qeXZ7ZyFtw8OIT
BclEOiaAg57jhlCjVjF32BeuS+LYfDivinsyeXhmYLFYVZCVYUcmRQl/Sij3lygsOmx3KK7G8lxo
qK127Hh7aSHgSUO6AMoyrrWs1q4j97TWTwlMq0mw4pWdSlcuX2xCeIyEK24K3MDFirrEczcFx79p
8LR4zuKezBEMFBQFHnJwLzrXiDqoFECZzgJs2Nh0ZaPmsP1VQahGNGHik1XrD76AvCJHgXU8jCPk
0Ic497XLLWEW+ZK65ASoxY5BlIXeRMDeh+6PawCMeZ1DfD9Smt5F4JCR2dGODPe9aBFt0PVzJyYa
UAHkUfbnWdO6JEh2kQWBkQhNeK5hFAqU1udh11R9bU9Fzv5QWUmimEp0PQEOfgB6jLwGm9iprzA8
kUPkcHi3KCMhvkWKGqhaU9tDAkSU9fxlj3H/qnO8nelhuRwXinsdaqex/HRA+1nanj75JICpfgy6
LZStQ1jve/TpHt0el1UMj6c78C5XNYvop8Hfm6bClDi6wCAM71SMBwEcuy1GUqo3ZMcUX+1zlf5h
sc/S+6ZKhcgWh7+GDZs54HwnakMucn99J1EaJyQs+WgsmHT+r7nx4SQDIn8EUC3HE4ff/MZT8P1M
qoA80UrLyIQ/dWuL9Bp7KDWAuERaYs0RhdSVFtI2ZKYdDmaGSGXk642IWHk0P4b6zIxAYmQnsZm5
HpEi7s+Ng2AaOOiICxeDJA+jQ0+UyUYpyfVTIOxVs3AJ5oz5punUeK36bDdsWkAK49VQXg9EA54a
nYrMZivadr2Rtk2qd5/0fLleULT/W66ScH0vIoQVEcX/dSacGx/CiBeDHvRcsPFr4hu+bm1tzf8e
isgx4TelzpUmFUHMitiLD+Wh8GJ52W9CQAddQM679mtJP0bCaXWCdpZxCgfn0KA5r7/TetDNWI0g
ArXx8rbXDDeorGb3Qa8ViobnEwmHEttcNyunW+cXPe/W/czdyG91CPhmMWzr94blWtnvfSlnaGtp
KpZMhicwurgQemDPDZq2ErQKTz7NIP70Ur48enSnNYz4qKOv6m8ctQiAg0qhACoEeKGcy8gnxxCy
eVpBhWKOeCjVxm+K/JSNp6vOW46zzgnFhM8gFcsrbN8sIdFQNUxVS3adbfIljphABOJw/vOLyz9k
vLP6GCYCvgu2jmHv7Q2ZSXwmdbLZL2XjqhN4XLFTEM0fY4yojkGLiDi3TAbqe6WS30w36+kffYw4
ICPM59Fd8g80W2RFNupdNhvIeM3mZK4IQp6sHZN/HQpr/RiOQnABn3iclQ3tNmYMaq3D+MlqCQMK
fSa4SxngOV1R5mWp29yyjFWuf+zad7mtNN97JCFX5a8z0M+xF36z5uOiLbja+rW3beC/e7LwwE+9
3iVfyXS4OE9iKPDCuMlk9jhSKS+JDfJRFGZ+q40ZEfZioxBXOAiH2wSjUR6cZT1tFHV+EZ753FsQ
ewx/aFPa+FeYDIIPpeqJVsoZeh9dp12X4SP/K5z8hqdjJbjigcNEhT6c24yNBxLxSHabBTy9xLAG
gDI+JWrSrMnG1I6xg23bn3SgQ5I6IRREi02kK6lMBk9uHJ4tXTVnHaq/RBgWVoKC78xtqoPSMTeJ
EWIrZkvTfCM1ublB71GDFsZX5jAp7PW6Fd23Bi8wHiNk9ZSPZ6rT42erSGSBXPk+hmHgFro0o4B4
7vjI9E6vF6eDnpahmPuz3Sb0WcTzma2fik8f9fV8L0do9NP1RRfMgnbeQTcRlOmomo1+FF1NQd5h
aZgFtUDCdcbAnhNXcC+IH3+ueobl+fcUV+/hBJCd4+JHoCv1wO41NJXqnF5tqcnwM5HUA4WWVVtc
IkOrd5j0rWSMH/2W+Y+bgGJrGqNzv/7Hns+OF/cpr+Cptrc0XxH94x2Wx8rv+wkWhrpDjBWMS3Ab
2mXcxwxaLNyfRQLDi9FLJamisnd8LvXMGWKoKQGImRpDQHTbp6VkbOKctx5LgjtvD+1cO9X/O5SC
o/4ETZiu0I8Y1U54mLomNn/FOlwN4QdxuplVEwWz+K3zCWweIjYKScr89d4WkeVkQRV7FzRHRMYK
vuwVliP3V0fw8eN4GB9WaBJdZif/4qwGELrDhGLRDhIaMep1FbcCXbJvwAMt+wAWp9btwUMmvyEO
qLahdJjJJv3RsxbMH/lPxKZ/Fc/yCUgubGTzNRFrm74JRW4VbqnjfCZ79Na2GilGF7N5apKlDi3f
zMm5TTWMzSSDiIUV/uS2R6OvzNKCv/gfwcbjZ+B2QEQfUTx4jQw9Xu0Z740h5hVkz7CS9VQbVzit
BySX4SZ2oZn4jGnCYhOWcEtjLpJzPxPp/zDXscGshZCntbK04LoUb1wicE7lCf/6NAHR8J0nMBoC
VXhCzsl8BOORgwSZYerLET/84rod5/bc2oEQLNGBoFNF0CANnwR9IRawL3QCIHQIV8UsRmL+jh4E
1rZGAukaMrqsKvIP+RAr1zswle+aOsde1ntG0sYKCEId6sKnoBFJrWrkjDh7cwEJY2IvaBa4yoEQ
mFek/u5ynCLooyqQLmDowYnthwYzAPYLqYQXvVUxcJnurCzl0MebA0ug0j7n96hrYjTsHppF64+i
8p8ai1y0vMy3ZTruTWQ2RJdG6PywKv0tZP4OMivmU/jrYrUnX41MSMk3y7IQnYroTM8no7hr4UBz
EZhz/jquGgdJoJSWC41U6VrQV7MI0aVeTZ5fMCRBtzjM/Q5ow0OAfh71uOzKRrPJlf3qiOXg8xjA
Z9w2R9qfdrFWvdxh0KUIjrAdxiDheZg6MeeTqi8iPj+6X+s1oGQlgSBhSaobwcTrdCwGZsbpl45W
8Ixb/YlxmaHw3Bjw9VuWW1/KY73FtL+ymV+TvKHQwKvHfiNZq/a5qHMUX+84m9PyKULvuzoMcydS
E905gF75K/psv8N7zsTOJ2o/Wtqn3rim1TkcltXECo3fOMIdvzoZnVuDD6adef7s73SpxQGvNOV7
7oky5+olQH9t66hSoBNXiu92rLQb4pUxmqterwmNqZHBRFS0kXRP+L+rMBCJSiAafu0Hd24/oHlx
WMRkowngvH3fidFTXXM1E6UUZYgTfXX4ee/5lg08GwOsrGKuBL2ANDKQyr+2c4/wYjuIIXLrzHEe
ZC5ryuTxS2KxWaejDskjZKjSl05w+R30nFKGyanpDev9C71a+XcoMUrQQqFuBkOpH6S9W+kjdYdr
LHigKgWp71k5lKTvpQaBIkc9x8RI9dHxwj9DZnT0qbXtb3sulO/EI8IINHi8nBHQOrZSf01kRwFB
nQoWfZis7jkEYJ95dtGU3MBNq43FUAx4fgprI0tFNyAWWcInBukWU0zkahWZOR0JQdoBrYKtN1aK
eS6S8NcqH1rmK3ydlYzpz8fgGsovj1U/C+x91cG+oJ67ZOdnLxveTqkrRc66EcJ44VhC1FptGtJE
17Skx7gCt1DM7Rbg0X8hkbQMfDXd1P7lJ1/DVP+5PFz2I5pgahU6DDlNLJ8dh6XeuEE0J94dDRhZ
s5zU0O9NZSUYv5X3ZfnernmzzUHbuI/dYjFzYVu4D/sSb/+IijoipeJkAQZSEvmPwj9JaO3v/0zE
9XDU538JSFEmue6rgEcAIYtz4yGaesMLrDHQFGYN3dQO8aYlBmG+MbbZPzgkuzpMkRrIRnhlsWD+
IF+r3thFgRoKdLP5fKEZnwR3OcXwO994ziunRaef2ux3BMPdZlONbO1f7Kdy64kME5VmnSyPOehw
ANufN5pH0RX71f27w+I6ITa9n40/4BZLHeKBEyfXwmy5/9ZecCsahKJ/O5+2Em2FGRQjoehHTdd0
qD6M35d2UxhE6B4d2UDBpPVEcE1xmdMo8y5Ch0DiIC748Nr9f+5YHuiQyPT5ByOz5lti0TirAk1+
6bkbENcAb/v7Sc3q1jjhbtVqKxpWDUjIZ0myxHZkdMDFfxcxY41PcXRqk68OT4CAjkVMI6gVLLca
4ve0jg5MzbsbonsHqSxd/XxNhQgoQZa0U7lbmWOaNI26x2Cez9dUitfz7nfL0Y/ET5PxVPd6yp1Z
un3giXKOEJLIp2XVkniiHu2UuaEJqhfnWW1dZifxXT0ZPWYrCwVGxnPWd2nbHbc6Lfx/Rxl+g7FI
tSn/f6w1oSdVGPqNPsNiLye0UYvZ00Oq2wpG9AAXqArfL8wO/4aKTSs6shC/fIHrr5ZdZIdib2eU
uV4CrXvbcVBmKEbLopwSQtcYFOKtMf7lCbOhJWZ4UUk0gvZbpcA01eKjoxCoiO+VwJS1KgvPDbOf
KApWfoZ9Lwvjvt0q0AWeGYaPKxeLFOM8Mavgw+OxHV6tizjVOdzoLOV7jOBxQlftIDNlqQFQdJAM
5zkN+BnHCAn6rd1rKj8ntn+sKcbJy7ZgQi7ukh1/xmBi5STudYgHpLuTh6fB7DGTE8qTgLp95hlm
jJnClLWcq7FR4IiQtcGT8vXF+Gf0y0OWIIBeyJp3Je1vGCcvrCkfhg7bGH+2PWU4YH70pX6kB/Nm
2qfTV/VUC6wabA/IWnaf/FqiWgJnH01lP/s8rELC4Z+focKxkfCJHyB/gm+4wTNbLbZY0/crSgL3
oNQpsx/g29rCgxECFbXKyXFmx0mw0JuUyxn5j3ECR1f48cBFi4MZnUWagtD2mYYdytxTKUwyn4m1
Y9LMvaL0ZbJIh8evIPfX6iKE+mPknpt736OD4hUbXzA7eebThrit+Gl+NyEYORSNgoTjrVCUh2j8
imip6EG/e+VRjQ4/v3tathk3NBWdrWTbNP7Z2aDrQE3c827aJ+7/e6KfWIE5FCa7X7t7JoQypLOe
zHt0Fjn8DEjeR8149oRfZ3n1ow4ySE5Qib5UaKyBIpLkMWbeGISz6WDHYKLq/6bOaA8BtrxJ/rBK
yuXFQQ1lPakhK/4BbkavP8B38e7tkf6Ut0QHiGBzb2m1Z/m+KdonJ8OY3/RKNVIaD2IKcZbYsrqF
Bj9kRzCXjuQ2e6RXY7upKPX0Dxt1VENB+6RvUZM0H1ykBq60dOjV/YjiM2EWH98tVugCkrNEf+7U
MrikwKWRS9WCpFirWRMN/NYb+XhCG4CL9qPhxQLit1QiUeN+Ar9SWuPEm2BOUVKteiQNYUMfzuiG
Z1eNRpKYYfZ0d7+QwvQRLUyU3BSXQd3etF49Mb1QWhmXj/fbypfI97WqaOiEJ9rsL2pZ5t771Fuq
5v3/GdtDWp9gwzQbX1a/Asyvkyb9tbbYl2i6qxY1wMHEVNz17Bc9ncw3ZIwuk9+I4LbJhhR0sx3r
v37O0rP5UQBkzBX3WfnO8qjUJqBuNAvk3jwwIIDp1QS9xqrlhvVez5CEPf9bDKpjw1bE4dJUhEkh
PQKH+CkaXvTw4/QPveyevAh61/z0xIwhQBFiocb55IuPTDlqfkfe6m6sGq4leHrKE4HdOVP1ZsYP
Z4MhUmrGT1GsusN4Z2tJWRyn9TrQrYyYvXMZ1jCm1JpETEMwpeFaLMTYYKeEZGei3lnCm3nEvrWY
OwzzeWK+SiOgKYVoluG5kTphw1MacxmVIuTSqkC54O2xFFd5ho0kdQ9i6j5v2XLuo2Hiy4v3PywM
potO3d2NlW62C5sjN/pfe0lY0rRGlPtKf7avD+kqZXPlR4TDtg5dq90oWITEYFjMGqeF7q0gEQg4
o3zhSulW1Q6lKz+3cCDcS6pL3ZLiB1NhqMz58CbqB2idPh5+oW/s9dZPHR8XEBjsVbIXzU+xDlIN
xKf5PTZoK1AG3bfc2MA8g1C2U3krvhcKnEMZXy3DpPdI6MASFscNuXBCisZDkJ+CmsR73RLXjtYn
sDRP9ugQz2qJ2DREsE//50XlbJIaCpxIz5AGZUEx2L7TLhRX6ONxnv0/CT+PwtSEWJCWBwvZjPwK
jQeTsI7M+2Y74zynsbfV3H2ioZGAwqzNDz8qfWuKOYrYp/+kZxk051QWurugc/O9qGouHlChA/i7
1e4lYkUjf+NUTp/FqGVFaWk64s3s5FxBNbmGStlFdoafURsQlSR+pqMTQTqaiJTckUzhjxcNlTJA
rJumhY/g7eg3ejJnu4y2+yeu7eft1AqUe5g7QQpq0rZi/dw0pCiOMvMUVV+B3FXLOWHxmvLE3Fco
ExkSXe1ndq/BAqKPWHwcQg34yAwLqQCHEx49JBz2ewnhIyFmJFRzTJrCMXq4sIQnuLo5HAXRYvUp
z3oq7PphU85Rgf4LbXCPitt+F0/WVzd0iiNYztzQ97C6TV6UWKsW4IxvxgSNOQy2nHrd4v0Kgwyw
srJTZ1Bfa1yIEktpTpzc/cTlruD/BLQ7mMnLrMbRT+2nd8b3IX+CDVyTVaW8CCcPrUM818Pha5ta
EcC/dWTGc3f3Xe/+fKGK6fO92Jp9STQaMOjUeF873D04/+um/T+U1hkenX6HgiqIMkfTzQHzt06e
7oP+JrRW0Cjnkq/CMHvl5f5uTQaJ4dibnPylN07CJHoNGLsN/tjykbcbcub4r6AsHeAjrhXk527s
vFI/Xn7R3EhlXhjDx91lyddDo4Ygj0tg5S0MiW9OwS8qrmQGP+/fxS79SEIvT2ByjsHZ2/3b7zKb
DRbbIhoiqG+raIiPNJVXZVAgcvZroFsIbKgygfq4sQswjuN9YLLfMTzWD0BwcfReV+wxJslWvAJe
z/zQNE+dAbOi3CwwvrMUSGp5MIe5AECSbE4PlSMp+D2tlJ4g6owyF+nUsHpIOGCPTs6JnxS5plwG
EEeCn4Ved498icuWbx2t4BjUqmXO25G1gVYJktP23FjWiNQVyDGyv8v2O/wefUFw9zD8Z+p01nqd
ElxwpwnnE9TlkPCH4cDslHXoB9zJRMe8vfR2U7jIt7EMe4WLFJRGyQz/tI/I2KXhMd22XmxnXe+u
y92gzl3kf7IezdkNanGOaDoJWQJRBGow6cO40vyQgAeQbKdk8Lc01eTNzKqrjH1rB2xSnl4+nWYm
NRjfPZF3CmHahxameXMR36o3fExpyTBWpTDsGJhgTS6EGzmw24Ph90P1C7IueBxB97Xap+QWWP5n
JD07wJFwGcFmJPUEc06EAoJHb+maOYTDdRm4sCwJbgem9jtG0/G1Sy6cSSiGmywpEo5CFiRQziYf
M0QNVAiVDCqSaEPhRQUdldKiHpo1gS02oyKX86+zWLscNY8BH3RqZoYoJR7pF4LXYmJmWbVyHja7
ej72SpbWwXT/FYUqfQhCkjQkfv9y6kv0fJjn3Dybz1YHFMVfzd4DOhzFXuwjJT7n7mgy25OFTGBh
wHvAvaMiSyNR6omH4juuIkyFktODbZUf8z7UhFs2BfNd1GHwY+pGYcOjaKvrhVNMLL57KERFP5Ja
uejRklYbfeBkWqo3hSa69YNj+zsvG1j6gp6ihVBFNJZvB1szggodP6hhfZc+qq0HwyWifxpy6UN1
Wfo6zdSyDlJ4WhvRqK2wAnJP2TWBbcID9LDjoNokFOGoFv8k5eLUO5SbktUK6X8IuOK7jDxOaADK
eaKzQvapYO5fAhckvM/pvkLVK4Pm5e3yrauPZ/nH+OQRxR10WyUwvqKZwx+2iKzFVIK9c43jy9gM
4XcktgIEsbEKhyqjjxhLJZgkxhzIBkBGC7Y2WZgcHHzMXaJQ9ML/VxCnhOM2ddsrbTwDe3pGCD5D
IQ6hZ+7bNNvHvnx2vVSFb+Z/BPKXZUTqQw5/ix64fLiILkeH19EhsCdDXU+B55oYsngwaHpbpNHh
xExuZvzrD+GSMCI2DIHMM7U3hc52Dlu1C1+pU7n72l4771x48dh3x1TrPiNv1K7VYQP8HtxIlZdn
mVOnw9n+Hg3IZCo+OYO3n90Eqq0EwP9T2nO0iLTOCG3ZuyrkY2/rJoOlZVNK0LgsUbckxc1ncpqa
9IAJRksIuO4b17fB5lQeu94mZYqwazf59bmTmXYbD89UQd+13pc2FzlVukXvW482nY5A/PhwOTh/
hmmzfieXT31KIhPTDDFNUJQZuDOS78aTwJpSviTtEi7m9ggtr2wuT2ttxWKbThi8OfnLz7CcpaCK
8s1utkA8Eis12h2ICcAPM04zmxd3tAUe5Mvp+uQzCUa5PECyap6bTOQbW/JvCfkabbadkjq7rYa5
42kgsnNCkHVUTXbl+dyy4voJu4AFOxGgVbQVkiL9mVawHJMhAD7IrjMIFDS566MBkeOWc73gfOqE
wV8ptGtJlTTB7PCVr0QzGQ9+Dur4bFFuf03baEbWAcpkm77WuawEL5cyVYLpDsgyPqtnQps/5JOX
VpGo4t+QZ8pToOjYzhL5fz+CiUqLotL7Q8VMnqGjEi+j4ihfmfGmFo41BjPt9lMThl7qOSjrC96a
y+IJDP8JOKOavdcQWO8DgrUefZvDZdELzxKemg+AdJnbgX0pGELav1MQTKqPxaDqzgeGoma4WaQG
oVyAYgLg5hAVQ1li8ohH2TtXbUL7CEciqNFFVyz3MFKkS0mJEXqNIcLpI6AX2Dc/XHSKke8u2t8o
DGyEM4KSaMv65pBFyWE4CzZccW43JxuDYHcREfMMdfAQcZrQl/0Q+Q3VdGRjsgxA63woNn4PkTW3
9VE9RPSw2bOFsehXZpl7o7rsRu8MVygUy3jdyb55BCi1UbkK5BqlobftMlAaETp/d4rkRFNsCahQ
SudIzqsCSrb9UeTAqlLiHfdUSgrDaz3CavW4D3F9lqJm5PDljS3COcjRR/jYU+Injhpl2F0TRi9X
R02KyPxSz7BY8NIfzTTUTV13wg0vS8UhAk7M7t3a2NQST754IBQMBQJu/F3L4EKYdLOM01Fq/68D
pI7ql4F4HFQLJE5FUqootZ9KsbOfjp9YGYG2SwPAaz0qT6eVWBXY+cb8bMHHCi0R3UL+I1dIi+Lb
XRtoUVaIDAIC84NVD/1aoD6sJeMqv1aN60ZYzCRPyLeg25FzJN6xO7TfNCMSlNWZ+itEDqdI1qfB
acces4UeQ/o3CogVDn6x7qG8+ESg22XeeQp0mzXh2oqUhm801n46YbfwUmJURVYeao4gq7FyPorb
LFun0IrUGC4fA3Kj4BEVvfGTNFL84Ho4Sowb00Roybl1WnrQhkYdAzdWeRw6pOkAhAaHs7q4peKC
q5htSJfmZBoqMsS7UabuKuEYWWmj3srsXXdPNyqDWdE3ySRczUGtZxUpOb3dh+HIfw7RZdENnPoN
NeS1nYbnBUUGyC3bA5VHLLUI6ZH1BVgZOouud8wH/dCGzFA+KYvDllZ6cXGSGHbg5xJXLcIfg42P
Gg8fySM7ezWs9LnRxTWTvjKPjuWPG1aQX2orvtle14xn2+tFYpRNyJdYdsvsGgAo7O6mQZ9IEN01
0p7kSGyo81KXjABV0k/sJ4eYQGZb4bNobrpiORQuGRD53dreR1BsewV3/KUkpbMWg8z2tmzJYPbc
qnbr/hfs75/fBn9sUPYRFbXAjm22EQyAKv/3CXbDOYo2zfJBibAAvIvP9xSQPqXKuL4/l/lb6734
aNNuuDdUVla92gPHQuMP0zsOzPrbCSLk6J3TSosVaKtuLakO1XTdDx8249JbK72KrPk5pYSxX+g9
IRI+KECwvfWfE81x+V+jWIyhMWDxKhZONhGurlWIfJWrxgVJs9OoGIfLa3EzZNdjNSPf9xeknaA7
cDe8BmWXOgz5Kl8+rlX7I4PFfWB5VHt2p+pa+U1obxTHRoKlfXEyysebBBNdvB0YAJE/arGaaoH9
f8Q61AFfYVNo2K1pbW4Y9E83ZTrCh4TB8VukDUQlf9NP+P4CiL24Ld61/A+ueLJI6OrZop/mWS98
cPm2ibgYVxZFW6ItlcWxzhQieSU9xVyy7LfuVHbi5XUESn2RiZ8Eq5HAIArhW3B9Jkvaqe7o+Kv+
i2NRsNiNO5CpZ2DEePAokhUs/bNB6HO8B/7LajQqK1YAElnvOrZbdAoWvCTqmZ1/itJ4l5qDgyRT
DfIsgx1WgGZFiTgquBWYEWQLu52xkK7wysFsiGZ+EFKagEG1Q++uAlcAhUBtnw/yaUBeEPnz2UvY
OAxKg3yC0qtNKb9ALKAUGbiiDgUnDh1b4dFVHy1dUoLg6Wm96qgiCbR0ovIVdGmK+0Hwo5nFySHa
yTGWo2wq9gf6DYTF+K3FlsM1XuA4R/3NKGTvCa8yhvHVv/sOXYXoklsvho91v4isCjYDuA5TBYz9
kv5trhEUsExqlkz+bbESMo/Rm4HfzcwYZJD8C9xYxsTECP/E+Gxks8c23k7wy0I7lm8mdnoq7vvB
1HqOU9LHGapNN7fGIzXtaVnWZ7AX/+wpqCPo+OX99wGL1rt9NKs3FaQ/jTKVUfo62j/VZ1jBnVhM
RNQrVaWNCjkTT8Sh1DdDkSAdl5rJnBMFYy2lbyJzjKOOmEz/UOQNuse2O8Q9e/cjSdaS+Brxt3bT
2JoSZqwTNiP3d+/WAzDilmHER5oP9zCs3MQzAUI5Tpcg0UgCMINpSMRJ2vOrSh+5ag5mCnB9Ya7u
I7IZx7+VgCtxAYsmeO+Gt4b0sSaDFSGKQGOVwVMdVTkOQ5wCbH6uDP4GRG3T6jduiR4vdbQA6ruz
G7PHAjyyiWS/HfVVOxiRNcNlElEzGeQFL8nCQJzv7/69d/g3O73cJWCLFU8zAEqKFN0oxt5gP8a7
EOzJns4dvXyJfTwVIxD8Y3KSMhs12ZFGmNYNBOnVn1q3smcEgmVD70r/jc9Ge9U2/qi+bN9bc2hF
jpb8tdW50nj37MXj5kzvIPvwwzi3nirTw06ly55iLhwX6nXG8eGWxvTXnfimg6rxWLt0aYNSZqS/
05QtRP9icPFQ0UIE9R8X/hLvKFdqmRV61YGGPNolryF5ON0RhvZuheMWrl3joVx2915/xQ7hrO4D
d7JwbIyVVEq1HvBEwr+xOjrbjYua4+iRtGpkZjGruwRb9xNpVwkPezj7NLklbAwjNYPKBQCsf+HF
dgO9B3xd7kJIz6aNIVnXJnfLKMKHzsYXlJ6qEGj9J9/9wzi5w8f0SaASFCRrN2mX4rp5lu73VF3o
9OQjFM04a9heiYQfvTZIfe383+LENp/ayml7lZAtd4VHqAtns5e5TDv/lDdV5EIDGMzhLysjtQhf
H6pmvzrlt/iBZPcowREp3UgYmGgIYtx/RdkdzAurE3tmcSAMV0/S5CgDz26ZGOWQtipN/frFSxZ9
spOjxaBhrn2gi6lbPDhNlLr/NHlU09yh2uNyxQRAzX9jtjMZHykAeEsWaIJxhtPRvlSp88Y8tyzM
+qGJUtrka7stEEcrUxo/oTis7VKt0O4D0Vw7ge3rBQMOeqDgUFwbdzJZ/EkjirjTpUQ5REdO6wX/
xG7h7yWvRxYPTZtOpaOHdpZB3r4J+Bfhq3tlKS5iLqZCs25zeGYSSXfVVZbK6WdhrlbYrxTLjKlL
NKIsYUxIFCthMNRIveucrH7j5tZkWndNpIeJN4LJTkCQshQzzYPsoVH3Y657H/MEzIAFnhs5R1f0
ceb6uiM1b09bIo2S/Ei9sYab0Fv6SVLRzXnENli6eRapKenyu4IrIYf8LMeI/kTqy9h9WFA3woFt
yPE0Ox7csVeKiTt31Fc1FpQqsVi3lCt6MNCN7XBc/zaJGxqao65nY8PZVuRmQYhD26rVImh7LFgb
mfidSmKxpb5iOG42da7eINKDLgrsJfz5Rh1excoRU8enAgOm1f9J0tcbHMphreufMuB8AyvCPmh4
b4NAnS80gQL3XhDMjdbJYFrPlZdmUADnDeuRHXMdqbUlQ1Q5+Q2jxfSd/AlD0WuthxL/p7iFY650
E9XTvOySfjWK5Hypc0gBtE4VPLwvYiUqdvEu3ZHHptJAkaJ5uu4Ai5BIFRP9dgqxdqt/IY9Z9KV2
j5XBKzyEi/cmAfO7mqZHHHCVAcWFIAC9WX0GjlYv8CTKTJFDBqGjFju5ee63yKavDhDeoSVnjnXC
6VYnc1FCKBBsZo/BVoD8BQPWAHUakAG4h/W6squlupji0nQtNuDHn4rqyR1X4pK1vsDK1nCA2B2W
Ww2flmE3zllb59uXZy6Xw7S30KAjrkv8cw5IbrJL9LhDkDuNB8iV84qhbRrF46GahbrDiN3TsxOZ
UYYMWr2BpSLF35zhNGjw+QBLq5+GnxJ5v3CQ4PHREHrQUa9wCtqtGJp7omd5sfh88nGq4VsGgelV
hbuIH7ypvgBkySp0ooCXk/hTrxCTYtaOlxGP/qFpkH+KhSkWpiI5vUVU1WSFIiBf1Q8Ly64VE+AV
Vs6XJBCteB0dd2kGP/Ds/HfQ/5PdhlyhL2lR2IQjifrGOS8V9bD3sNS1gFFglZXZ2h80I/XoNARn
omRvDszvfx7/Ssis9gTyHFTlcAWXltnlkkIReFLCrUvQ55PPEwnQcZHccCoflcq2zhy0D7yZYgvy
7bngQN+8JywpzORIATmFSHcY1fwymeQut0w2kKV2iLoGwY3CLce7HLlmAZnGdAwDK7ksJvECQIt9
ICtJZb2tYjp2AqFz37HEyfJqhbGZmAbIsJSCrqQf6x81cTIhCvHL8GrHgBKWgDSsZfglzebKTbDb
091FZw+T5Q0NLHPq7L3O2ufk1f8FDTBsM7oma+R+AIJAGg6sGhx1ZvvVyaPFjIMKZnD6cXBSav2e
QwzYtaXS/GEfrjI+iSgufCyts7OEyw/hTg8CiHiSBA8U/fG7tacDtpIoyU7oUAtOb6vAKO+PgRwr
r1xE2ZU33pDoso6qf8Z7k/Jq5qCqQNUs+GV7BjU71i/6Ez7lLkqD+ttu5R7kiIKIgCwuX114cKzs
eUGyXAXxFAk7U56WLmjBx4f4/CvX3GA5CUO2FJ47pJHOp5l0sAIzWk+xT19teyfgWHCbk7VDeVkj
ZQ4qBDZ/Nuhcpye8iytMENJaQVms3aKEEHrw6Q+sIc2XCjnMnovPyA5Gxt9Tk+/iFTSZ1MMe/ll+
w4Ax+As64lsD5U++vAYAhS792TWddC4z7ffdgbxZHbpJeUOVGqExLJlKXOaymr3D8vaJCswFP7RP
UOXwK09AH8vrZm9l9f7xQChtI0ggrDfsWatfmBzNNzAMU7fZsqjrKgPSk/oF/u+aVZNuRg/2fOOS
W90Y6PRXo5ZN6XIrSl/pPeXHIn/s1AvNZ8TVKIgK/uaIq0ZhsdkimDSZ/pVLlrVumnavZA6/OIka
VdsnyDLEodb62s22YjM4GNBjQkkpxsTTvLOnPmLbXaIGxGqHl9+gXXiK1uVAbbUqfIzSsvE2y6vI
j5hBXRrwwd6JLEQYIFP56YdPKu1d+vCghi9I9HAQMv1LZ/45BwXnU6Hwvc6vPty87de3vkOa0vU5
uV11PlLaxuBVPKnW4haD/rJpSEzd9Dmdm+hftoqSeKtVRpMN7RCRtXcFEOP9JqaPN7MOE9BiY8nn
0zmYbpbXpxsPoZ8H24ntguhpTxKifVrPB4wyprdc0a9pHvuSTRu/THvWnYcifv0H94XOnc9Zh6zf
4v5+uWMYj04xMn1seBfUP5WzLW7j6B5U/SRClW2r1jBcu6Xq4qrmNoYQYPeKn2bRLRuI6RW36Pqb
Q46w7jfC5ugOHvERdxWyrNzwck2MhFFfkrqlIvjBMDhTWvzNJM7CZdoJa5fU34YMlY/rYqmoEgzx
rcMtgZNV9AWhRK2hHONFuLAsdLJ23PKAFwaSe/4QrLMrR+u6EtERzZ1aYL3ef7erp6h1VqJ+uaLi
wEgawzW5imx5V1VBattkD2NUTE3v3yGD5fALIuSIbQ7+yz1eNSpZt7Lfw7uVAySTR3Ek0Y2E+irC
/zXObwpeNPqH06YlAeS99TZFZcbAZ8JMtBAUb+Yr9C+6zztIdjDzDt4CsH/JZYr04ZEkSREfYz5E
0h+V9v5kGIZV2+tMwqUXj7+dLPfd5sNRNBf5s4+1nLc65gkO7LjK479CgpYcC1Tz3jeHQl9gxqWw
3dhwEnS8boDlzi3QaUVUsIT3gEPLAepKCa3zROJjOvZbeumgn/0WLro/7ThpcJTJwaw0k6O3Cr2c
j1kqIUC3qmrYjTVD053vf8jNEoxw4bdO9wwbZlCne+bHx5xGui7ruukpmwysupg9qbze4C6il930
Gm6fifceqe4qrI9ssWD7q83oKkyYf2c/pBAqPyV+WLx/6sqR7cgSLvit2VCTwr+n1kjlFqQKHteV
lR4+2aubB/K7IjACrWaW9AbhgEF1Aq5YrFVYgyeIcLFV8gydik2+l8Kt4RKLas7IMeh8I8muBo+D
U401DbPWEay/rm6+u1SLriLS/GcqaBPSVd/3k7p7E3Tx9dqaaDdWAOr/kpLAvE/UIzRnMxjRqwpi
Djwn8u+K5LHwtHqnpfThFHby5QK03hncvEVcjRkpsFc4tKj/SXEwD6CIzl2JmSYmER5UbtG8pPQI
7GnNEsfYCUAz8c06TF+l9ZdKBCTges9Mq2j9MxQqy8ZRw1qAyvSvtl1vw0PButtVjKsx3h5xCvww
R4shBhS0mfTWKjhzlSabqvUPGdcUhtVBA+mCbKaLfV7SbwgwZCDdSgol8jVRt3wDl8GHWYUVjYtz
FTErrKwjAHfUcFhHwfrczbKVYBGLCOJ2AcBOI5AwSUj5/As/gAqAOnPwzHlda9hmKiVByQOjz/F0
233Gp1L0LogQqpPqpVOITGelHjXEaJHXtMaLIjFaEQItUWnz+WbCa0QChYC2VkEU3jlg59l/w5JZ
+VsCLoaG/di7Z+BzWPe4/uk3CelOKqDikQo+6W55ALwcdm4ewvqW59em7LVXdtjRdMHD4BTOoPhV
UefaLb+NHw5Jinyv9AZnWJYMPpwDF9zEY11aQ3sLWGb0z8HxS5wOjalnuzgKx1JD89Va2jo6f3hh
9tPxRJxg9Y1uZtkc5HDTbgTQbGQ9QA1ckYXDaSlXqI2m+OqEY385GFKJXE8L1zbsfi4VJlU21Ks2
nrFjkNdZsGKnWScF8DpLR/Crg371153R9VCTgZ9zawhtFLVa3OixW6DpJKH/pH5CekyWS3jEmb+L
bBUI3bfeapnzjL9Uuq7q72k5osSbIeM2wA2lIVU2P4yHvOfC9ZgdCARySQwPeMPiCSB2ZeDBRlvv
RKsE0ze2+SJwrLiiXQI1yMHw8jCWpAgsK1K75t6s9CNT3drpTPuc9KPkHNRAF6gM05xaWGupGa62
3KzDk/HKJ/AiHl7tkxsXqvFWgYPhunaegqigDtBwV2vG5tJqrV66Q4EupEgZK9WyltCMAuJ1AR8p
3SDb6ShvWDmRUjrfVkIHC/RkmT6i7qQSohBKGDIMBus2DWYPq7dTI9uuP/VujHufFaYBQPlBs1fD
UTvZqONvfPzUVMd7VyM4bNEob4WqH6AKow6k94d4gWXdAJ6tL0L0caAUlTE4VLwLJwFKw7nc5uQy
xUu/CxAflCExmmSMgMBBYclwLAlRCFoihq3S3hbPUGXYxpcro6Kb5hw0aoT2iMMkFCCf14+ECeF2
zeNWNeDjv4vSTd7mgPGTHvWW7Db0YQ2py3vzaPiQR8n0+0K2UqUWGCgFNYruZa6XwBt5Ah/N62kU
/CqnPvuPI//0tU+pa5wE89+xKMYBQdv4zjB5Wnn4dv0rjDOVfFdHEBd5OxUvlCXHSXIemkFwusTh
lcF4MQ3mMYENdW6+mWC7JQ7cpIiFd6qID5EwPCndiizLxqvElm5ahix0iKCJcsQQ/wByDuuTLK6n
m4wZamR4pzjqpVQYgA8wxnQpQkyjG6k4ng5wfWVDya8JvgWf3QxFdyYBdWibnvXQ5rI01mq13pdp
vnubplD6KLbB/x+IM/0boU6kGSVEb05Zpy/waL1B7MvCwWQalHaJWydble/1fKCojKraeWHlWaAY
3Ff2oPwy0oCCAZvQ+uvEgL/wQ23ediyi6DPogb75zOKLHLSq4TJ73YnLA52s1HHGDLmcbwd8J0Xt
PXm/h4KI4xa/Y+JcnGJLnLZBJbqKJ6pbvwBfW+fPGcvDSfbeuC8RYcE+ge/j9xv5NoasQeeRw/Nw
Sgo3/ydAyvwxyJr2xGtjqDrcsUShc7ArmWbfzwXs+ihSMfzi/usQAOPct1kDMjC4ia0umtCEeBWA
QJM2fWNeNgBgqoo8WKs7VQ9wixqsyvQysA2FB75gyDosBgDwKb7bKKLTcUpsSGmAHqAQQVyXscvG
QVQJ+dESvnjMSje+Hll8tsfsPgIEVB/d5i0bWKXIvR6Owaj2p125VJkACG0WL1wvFpU51OKpVeVp
dXMy5Ek45S0pIDz/drXSNK39wJNdwY02Pno7fajPJ9/uRtR3Q1MbieDDVWlkr3/IEc70OOW7UZGT
1CodN0XbqrVFIUrL+94VW11EfE7CLlEmDKFcqeAVDWfvOlK1RoifLxiXj/4vINpnxQjfHZ3urCl3
/VenedNScKcAjjjky8fe/2yZys9B9yXEOTP5C7dJjcWqo6g2FzMGgfn95rGiRRXcRdyBu7+qLHR9
WDmYwmLphnpsHyLv3VLZHRxxbbsdCCBJ5WEwCNNNGXoMgd7fE+l57kzcFHQX5f7QXUd2WBC2lNAp
/8iZUaT2baAAEbMJc69NCRPWJ0sXW9BHznwH33vqBgZbjPZJzATj0XkWD8F9HPPq9ziY1x1uKEwW
0uBngvilcXAxJtmXXPVm7VBaDNLzsK9DB/DUN2CN6M47iOR0ar8DHnnz86j/FsY+ErMbAUed6VW4
8/8R+o1nVUEXtY0q3/DlCuRwd50eiW7mHCxmXoxyf0iDvwFiv3p/32ip4MYllBgLBFWGMTj6jCGv
BtxWWuG8BLn3jY9aoBnT61faoDmMg45tmxhCzefK+fvMH0WR5NwIgYDhOutiD6F48QPB4t/IVbVO
oY9NYZoL9SFhgnanHZoH+DKP17fnD8QFUUwHD1qfzHR2cnZkYFIKDBl12i5wUHjeFK4WVhnFKCMl
cmHg/kJoxX1fiHoT6qh/yv2fjYMJIyPJyxZ6nGJmtefIHwKUzbuAI6b4ddBpPRJTwtorRQB/h/85
d5Yp/c8pMOfEwPVNhhl8J0LUjy3ozuUH2s/2tNTbsj4+8yBACOp33Ilpe40joAzmCo9Q73qIyLix
bmzPoQSwfif7WBWde1pIA7v7uVinp9tAgBhVmdMjrQlMkMyLLY3VwaEVS2ERTBWeNJG7AssqoFbk
AoiuBJpVviXOmo1rEU/N1YCGkJidzK2CrUsvUgr/lJ8YQPiKYNsV3y8+Y/mGtms15fqCtOfwo7u3
AOMQPtIi57mXXMiLGVDWnbU98hztbKcYGwYNprjpaXN094evzUOXhJ4djh/XO9OXIRE7UmdwLeBD
XP3qSgOTNvozy0uAyAza0BBG3a9A7cmHE/Bj36Wm4+T2jQoSdRQrI7JL3Rh3MH3Mmy05EMjlx+34
qdfBTMExR6xfsZ0jC615YF/MH9JTcOxxqYPhPl1Q/r+VEJQDSJHr/lNmcij9kzo1a616OD7kkDUS
eqfot2sZp4bFTdWzwG/4Hg+3cB7rGhW8a5eg7k8r6yb5T8S4MJPpTKu6qTxHPH0FIWEhIID+9vtj
YxxUeYRyLCcqLrZFdNjCDaKgMhb/o/QrpXteFfzCjFbT3yTn/4lZUi0zSGw4OSQ5+1c3hqPvPygd
KvTPyjGaU1SFW1Gntu4C8N9mrBb+tNX6LiMq276aZhC1SPw2J6THv69ySJyr+Ch/fKXWc1cl7jKS
O7snUClge/c1JKFmXunu7bR3GIoO2dLlLPe21qf/b1+Z9haiDjR82BJ+ZAWGZx/adC8QlyAzRlt0
EsMp9a9EWgrUn+3wSoRyAZsIrrIJDO3h1FyL8FN8ozKJBbKDZWRBN4RnqoUXLD3ayNKS+YQBWOLu
2KpllxAEbtHDOvP7pOdUFxHM+X7FibJfFd+4HwMsUBSJSq4MBNJhlKGwgUIM+mO0oqRPF5iI8dh8
3v8Hq2FiWEWTlNizbRei1cKhCWlpCL394CTM0skXmfS4bkh+E7hikpk0TsftoSzkBlhQYHVRbjGp
uG+XEBpyuGwABk7wrwXt2qv1BLqRJG9qwV2XWI9ivWtpyFCU8qjt511K1/TT1u8LAe5w0Nzt4hcB
tu4j/O04DzsppQVHuFJN76d1/0HmZoG80vELUTBszdsLfexWQZM5PlCld49GAZVHzduDRdFx71iM
AdZHFis4DptzHIcCDEHuYDaDP0hvLYlBrkokfQLrv6JxLtOukywb8BBaoKMvWtXMeuRWMFVkGMSX
i5P1Xd4CyDOifSlo/frXl5ViAui7gwUWLvm86FcvrlZC4+0FDRJ5mduZyr5LSb3kKqP2h2Cyai+X
BmWvbxNrpHD7yig5qsFuA0m/6UrNDTWrQ1sneT8OuNfAIJWZIYDSvZb4OLJUS8BJY1xEC7z2XsBY
fqe4bGBGuyynCfBAANwkcd2G+H8xw4AbtcypZMWTlIV39hTJpuaBmlC2tphLhDZjetdYlveb4kl5
nDm4PVuxV74oezuG1BE4ka0QzQfKhOY5VFfhjEunan1qs/sz0UXIxYOzwRZ3riDfwsjMV9BTzhJ9
9BZ8Hlqw9uH6tBsmcldss1eHUhZtPWvlmWMxFxHOR+Pvdj114CBWuz5CLuO8vBwYCrw5a/P/EnVq
2MABIrmjIcrCCY01rXlLJ7eSPkB9ao40pvJSoLvI55hBxs4S8KoLLKQmFGHVp7OPDK1l/qcwI9Jr
7Jh0wtXKPqOOIvUl+Xy+LDz4bkZQP4uErqIse2ZEYd8CUpuql6K909jC9BySdKNuYq92hFpGhjHk
3Judb3qv6VDdbt3asGroeZVTKOtoQAgbzOU5/eDYti3+uO5iD3bVQBZtUJZkUWZq0L0wcRrOMTtZ
zL/gwQ/riwsFB8fAlhZISARx35Th4Okgl97WeLoebaWmxrSYYaPmUVpboyvcuE5ySVvX9opOhDk+
YMD89UuehPACDAQwrkUaeFe6R+xQekq0YV6FzHA6SXRzFoUTbQYEdWd084t8HkH8l/pLqpuIGYpl
NIJ4Rts2u4h7mF6tQhcDXl7MTObzLMLbKZ4eQShO4Nr4I5T66QE1n5QnW5/wz32DzfBeArJfA4fc
tTzAHqPiwyd04m97b+tlaqbNDTz5sLOVo9MrZtPY5EMRDAXCaoXhrVOKhXSxL0HZs1Tp1d/qedGs
sNuS+XNgMtRSQfuFm4xw85sqxs1H9s4STXP3kuq/ZSK9cmad+ypgI18pZsNjH6CG+ZyjphN9z2fs
8jMd9N5ng8TCdGrFq8rRUjjZRjGXEHuOnC8IIgTGmpoPWnhLPAwhVK7/KGpl7M8nP+68DAGFPrzS
hfwqai4mF0q9DNXxNuL5lD/unQdqIvEinCAo1fee8slR8TT7VlCjRgmjhJ7qGcZBukKo9nFymBIp
Q4ivI3e5Cr2p+PdhR7A8tjLu18h4yBjRLyMqyF4oby3nzHReNy+RxXQquYO92VD0U6U/Sk35fTd+
ly07vMxRQp8TP0hXpD7AZfAwiJyDb7IQLVCY2j5mxtIqgBNwBszoNRMxGN9VYRkKkGhhfGCpnJ4V
a6tlQou2T+GUgtYTPShZb7LrROuZt/SV2sMbhdIdroaIK0+to1H3D3YaA9wSVgaxtw07unqgLuVg
zjNKZNbCZmQj+YxA6zhwjLoO0DROVOnKHS2+ychwVisNaIR1xZemmcREGBbM6mUUBhu2KPSI0kRR
fZF5jXpo9AkynzZLP++BDOnwlFU0j/Mvpq64PDcF96AAk6+hgNI++9EXYaAZqojlWDK/w0CnioJO
BevDZI7Lt22yaAoUSy2AOqc1+hUCyeXuYIzUTg3IFQTB6nOeNfNPkpYd1+bbjtJKskctki37Hvmf
IAUoX/LdL4c7iWTPJxxPw1yp5zyPICF/Z42S3I8F5UwcuGAm5lyJTF8DdE+pE78Q1bHUlsk78Quh
hx/mVAIFI+v0Kq6FOXnch/Xh4NASDYuENHWh85QOvhuuANY8L/31HKTniFCBB0cEqB7s5ahCNnSt
CGmrQAkdS+OYDOQLZy0PFBTVlsnmJCdR7pyCdXXpU0MzOGKuzcaFWJQnnx9q0OzyUwubn8WOAT9n
HDoZWuhdbWXQ6dDKn8AWNiN2pXvvj3XuDzRTsgmHlHgp4Daq5MVDoQ/iaFElBfamR+t/300fzsnS
E84L1FJN1XaJKelEod6xyTGAGjTQHeZuheZS2X3BsCkRbNdrjgLI3hcfrPhurjh686Hz4eg8a1Eh
aKsp5CTXfftO3NtA8ytZi1vLDrXiWjFf7xqMIbZwKm1OYc6nDrUmGwemmZWKdoJUVC1qRDprBu93
O6n+fNQXN5O6JcQuta8D4kgIwWFTevE4vDcc2z3HywPCX81kgLHjh/p3anuK26YdDL8b98EFZBql
z6u4zSHSXTpV0AApVmpeYco9C7Jn1Kj1rZf3NJPjSLYqLRq5qmxDAZ0IraN2lVjnNXgKx25zpKPQ
BoJ+PcRmAsWmfXKxWwshvFy0ECHpTWS4aYA7LBu3Xiz/owvGeyHFe4M5Z+6/FPGQiYZ6jZSlu2OI
2g2Zz9W7d9nK8xBomsiTgyM855xjnP9tg+3vjnM1YuuURcO7FSv8bF4Hup9txOi6SEiUhIhI6fBN
0njTOzY3hJeHBrdiHFTC4AIoX0LfBPcygBejHi0B5AKW3KIoFxrfMDdJoZ/PSF970XN0FCqSFieT
8cxt+i50jiYi2xebkSXZBKm+qVyI1ksTLkdkk80eRIPBiLiyUrh5B3haAn2w3OzHQz4q57F2QrVx
3nzWIoGxxTupD9yuGvCsGQNRjgK6iAqaTQ+MU2tOYB1CiRzwWaQmglgAvoqR4XqM+DEkeSX7O7Dj
mS4sLJrOO6BrQMO8bg6vWeMSLeAUU5vLplIFHJqSd8WEs6vWa1+rxcu0WFzaDfIScHDrBcm3ylr6
Ds4q3GV8RRnuvZQ4SWtsb6TXSkPvd1wgQzFjAuDW2jiWo4AHfos8jAQBLaMY723qTgpeg+H5+Cg/
QQBQSVm6ipz9vOA8D9L57RDFaljNZWV1rpUcDo+Cy4g7+fgLYKtGQ53OVNKS9u+53v4G5hVok9L4
onN++ifDsXkii5y/tJphDmQ81uIPaGu4aUYa1RmfTdnHFkGXDfx0ck0qDnJIXsmRBE5sp3JW/6xF
IPaxyt50I6VNxaa0m3QD1zQXwmfp1AvHEY+NqZOvZW/AcucbwZ/GkEf8XxcJkle4ktR1txSeVvwo
L8QkiIUDYOMSw73DLPHwBxKWvmEZ
`protect end_protected
