-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
oKskKVXz7RuqRZVYeUcBUVtO1OJjqpi4Pi1T2sEhWRPGbs8C2kzYFz3s/c1YwtB+deFSfGhyOA7o
S7xwOed1Q5xbxuL7J1AKCwhzH/SM5Qw96BhROqSt/6ONfhtH1O3CmPEqjeADjUOxeoq1t5DhQlOw
xyhA1NWGxOcTSIzJHGM3vYoDfjJ2GTwYQzJ7uDV/wfNNO0rjABlw/81RMR1WpP2Kgk3/k0KALZW6
YpVHY8eaXahhOE/PZcu5psTu3mWJzIWE5Mj6pZ4zckHE/GGAK+8X80fax+dmUiIF8QHq4DuLAk0R
JKBJm6395PkaVPz8uu3HWQUQQDGxU43QANxrFA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 13296)
`protect data_block
qlUdWYrlqOX/h6wL1NQrPq3+c5Svgm0p53dI9G4LABFBIY/HdPylqsmAAzUubAHwX4sV7FCidm9F
tahvVkMgu4/f2GLGL+o8KHER82xEMSWmxq8Yrhagsr1f/u3Fto/RYtug4zP+/5Vi9O61Gou2frp3
y1E8O+Lb0DIv1aFtkh6kZmY9uONe4Uh+K5r8StJaBJmwE6HeKXd4lvICMBxIe4C3Th0ytT4NGBPl
/glHaT79Bj+g6XnGsKdf95tpvVMZjbHdqrwn1FZYfM5WZRuP9zkMx5vUONYgFAVpjDrq5875kZHN
pivIsrGNrmuWGHNImSIyNoKh6BbmhziMYIa8MuZLk9cR9/1ik6YRhWOE0kqZ3qJ4VoDF7x9g2Wym
Z5+3j6HsA4jy5MDDAyqqkXwClcxblhhrb7nJxVR1b79syhvtxpHIo05qpSo9fvLyJeyVWEdJGeOS
k21/H7sA5hu22venMHZ9khB398G76bVEm0N6gteoSSMKWgLr8xxwOQqj6hHQrFITOEH4tCnWDRgk
Zfo+jCIEuDzThszY+m91H8rZiyX1VJyumblF49krYYyo2e/NpIL3o/lLNM+ZE6b9s3Qf2CJq/S3H
pURGe2EOHLiJh6CIO4rTSf3Hr012DO4Dk+0QkmvYRIX9xaONXhGj9z3BoSgjkpBB5hplPy6u6a9g
ZJbMSiUe+tPROsaMyEFgVTVCnh0QPSF0ijqDB5mbZtreH4RjawhrDLOfg7U9xQbXTeHTeCRnLSKf
PsPqaZwU04zhBnIIJl6a9qS2b4z2KaORvbgiwsQu492U18cMdaMnTQVBuZyYmnexC8oR8K7Sdet6
oSfXWhVsEHX48rpj/ip+3gnlT44rNrQA1sC4SZllBNAytkCx8oKlTdZfeHIe6U7gcyyW7k9jbXnu
FHdwcTQDYFU1rWAP7FSZUCC3X8vYlQdvjJUdXrfe6NRzG89qqcvoszSEFX39pfXbyJE3Oe06MfJf
47d35JD0mBBGSNF6JtrCqAGGno1KQ8+p/Pspz+mfQKfsm8FSvPjT0n0KZxJE31bfXi6zmvEhSRWI
JhJKeOqV9Vm9CDlZDNLGpy0CZcMkOar/TL6rMFrSkbV1mhkqabNK31jv11BRTRj2YBofosDy+jhg
jnze0hiA/NxG6IUBRlp+iAXrmIbfQ9RZJLeUX3hAUHKrmgkfrh5zHiJk6nVG0LwvEIrV/10+5NR8
ALqe1/CP8zdXgPyeWNmGDAFxNKVxhujiFG6m4U1UDWcm7yucOgWYGtyrTxLb39EoSgtm5fCKRy01
zj1LAJ97CJpEu/dKcj/3/+EAYyveISaHEQttg4HNrJ6EdYj9ckUGnfbwv/yXQ3p6YCpfXIPLUNn0
u09PWHWOLp56HXZ77R7VTXN8WXcOvhRbPIQuwq5wMocClIta7mBN/Fkcm2VuveArMWvAfM7+67gz
qYdU75kHBJqWbAx7ppDe9VUJWfPHxzkFusbhy4ce8qmJCYqsUlz/QfOzKR2zbNsD+/+Yxzn+friR
HoAOx5UymnUFZKP+Y63sOlmHhdF3A/UbxVQBABS7haxXtMXbMwVudweKh5BB9c3YL81JiSsxvjqD
Xix7Aj94GfC5hCn7DU1yLsFda0qQ72fZA+Sd3GIfr8/zmMMCZtjqaeEQsazj2JhxcvDEj7/k53zQ
qTHXQ3epoPFI8t8nFfldNgvpT5E5oeH+Gt4zjzVwmfifqXeFM/c/0XnzaTvRujroxj/zm1fafVfA
AlKEmg6ROkk0cjSczr6umkjLzgAOJd7AIvApInKn50wa9HE9XsUJIeqmzI1XYDJ7Gs/49x2twQ1t
4w8CltnBL1PvQA/wOR7Pqf2ygU0WuITw3ecLyYsFNPDzhIFQRf9u6aXXWqof5ZcCMir4NIrsNI/O
ShjMiF2dAs0Q/u9/jHmYOw6np+t1RvoD82VOLs6s0Krj/RVogK/F9WeDsJOXiHryWDluG2rwyEB+
0cEr/tzOM5+CvUCUqe2vMl+KaSZwn++BlZAj0LOBDtidak+Mvfi82rcr6fl9ls9uPV5LJKbwrAEb
u4hltOuoXJ3xbu2UQzNfyISK+/Bp/rkf4QZkzi2+yrU7P/mmsyPgQlbaR5oKwykNNOER/Q3Q5U8F
kDAV2D0dmFyiFlhfWthlo/dIUaKVhOl6lHwnIt8UNmajiMLRD4J7zlWaBEhkiE7Voa/lzbbGKKdc
7DQYgnkWAEbgV0ZjpMPdbevQIOPY7JpZAuvunUM/FS0fBSwBa1RmEKaPM/9S86RlNxBlw4dwjlBI
/TaE8QI7fsIkTGd43hM0Nfdfb5ra4xK0ezBQTjPAnJ6VB+tQ1HKp+7j0UIX+XT3TSsLS4Ui7j3DU
FX2og70auqsmhY+CCHNuIIQ9YuwRAGhth8MWARJ3SFU07UYoOx0OkZi4/OtyODzmHQKUaj/mLWox
pYXycntnkPdYPkYoCtde5oD8x0rNpEQTjw5SIN9/UbxvZ6/UjlRbSJta1aIBHhP0i/R9ULLalru5
SL7SBepq9qK6Vl4bH/0XoppACsybSKlBItZS133GWxR8UreKiwh42iWEUkdTKTGBSI5jWveeccUd
xpJAS9U/2u1+ROWKpbxHwsRHk7qL2/A/7BpAA9Nbl1r4VMx4qecemIjR7VbSc4hBzMBqefLF4QsR
DCmFIDLe36v/I2Pf3aa96ugSDBC3m9vDy+zgbOGxl1QHH+e8FfXixjqYlItbDiFYqn3Ey9NKqBbf
5Cz1uu8amV0jUb5ZF3gruXFzINRaya/6gv010ESIq5paXuOMFb9UMX3bFzxJzyhOgcvp4YRrd7M/
3QtDKIyz26t+Pw4Zt7Gw9RNQXN3eY+iR+oG0F5bg3Ku+lFzR0QMpRt4tJt/ToYAV2JvAjgkgB8b+
AkveHjhOpIxjP9PEP39SW296YT3wVkirzUyYB6DfQnK/aSu9SfOVXZPGel3EqMIoBcpayoWZF540
yFducHhvRYuoZUp5OEGi2/FKmUFlcf0LpiSEm4UB1LjPdwzlq+iXEtHlFJBRhWUq2pZN2BrziUdD
cS7quos5QnJRgwhfVXTyi0TY3CFwf0HJYEap+Ey5Px7bgrSfKClCu0tkIjeS7KQNnPcFznwPbl+s
k+Zwo27Z4qn6BiReBvaVMZzQTeKXS+T73kUCGP3qWfEMV56TcBSu4WqCeNSOsBVqsG7Uer4Y8Ky/
IgM1IxnhD6htoKmOmI6Ku9juvjuxhbch3U54Ulf5KxWWWf5wQavZN+kfgbWvZfbQKKiEuhR3JZ8O
fQ1rYkCBWcU2pgFfPG7Hucye81bEm36n+VDIIhjtNLod2l9CmbkFqQCxu6lL+j+KQOT2zKA0sGUP
NziL1SABCKVylQEKWZwJpYbyDXIMyjxrlNPtFx0Nh4r9uYXjgke6yuiNf5HmiuWbCJXpFZGwycIM
5P0S94IQiYXMoBw2jw3sPVpTsxridGHm4FzF8mPsxOAwAx96+ef+bKm+AShM6Tw4K67sT+S0djf/
q1Mr0XYiT3w1pPeVHvOyk13Ivi/ULnJ/wSKZ6rLkMkNBLzQx2sZ6zvQJQEfKPGK66FBLzfVB3YFm
pJaSi+dmetVNyv5z92d8+8pYoY8v7PbEba1Py6BzZT7i4YF0PAi+ns46FIMyOMNIPiUx2VU8aUZl
oqvT6q8cg0zVbCBwZMsaXDQ7unWPg2lXakCBLaOtpGo4j5EjPsWu1tvmTnYxbvUWTDNxmnPYSLH4
A6DS/ezqIK+9DoLshpxHq9m4DuyTHGUp8ozmA3KuRzCmkJnPLzoD/LsfXjA83ULzFM0sYbLK/8U+
ylhUgDvGnT6AvWbpUYtacO0RbCXxCbb/HITZIvUL/adFdJHKV8Y+wygRf7yghe7MG1qGWLrm1CzX
jVldtdjdyF9HnD9qhk2t92ruzXv5D1ow/3QXOkor3y6JEBA1Hd5EHiUh2X9nVMdpUZtbjBFoDV6K
Ju3lFOEKHW4dqwX2tSL1lU+fj4HLFCkvHlXUslaxklsernXq8mXREHfuO29VouDhw534CXAGJf/z
cmohMerbYtIqAgvD4D1oPukOryqBsfR1m5hVjy2DgzM6q+hZe5vY1kDbh/XaOX91JTMoT8BqeMlP
6K6WAmZCfINuFC7x4eLkhJ4Wu15QnZSDjQ7FPt0dnYCLVWPqXA6cd/Tkf+xykj8yNst+N3DyFYz2
f0eSWrmsl7/ZGf2SLYkcF1lBcSVjnIzS1soW3TYFhK8qv1j7Bkdo0NOqaLcWWA7svVXoaM0hMdSC
KzQxRCslzG9UvHlhOFe/59mmzzHQ2IuwC8le+saz0Jx7ooyze4LRuMFOPPd/4E1i+u5kXciwf4G6
dGmI2X/OBMmJ2+KW84tdIoNsTHEpDyIhPp+Kv9+lW+2sMBhgjWqDLBe//JnXLkAYpJInJMRVlmiq
ryS0t7JzTUsV6/pujDCZx0IOg8sCkse31QavHpa0IsOBt1PBTo1Kmkkbs5/H5UdeiOfL/iq8lddt
9CHcyVdY2/tB6L5QdrHlgNR1qqdCak0UARIYnmyezSrDTwEwTPW1gogt55TFWGyI8kw3A8xVo6wV
o7bwAvPAhujpFlmChXfSt2bsbNqXuye4eSnkL4El0YiYGoCwh6aJ1nEfGjR/sux7FD+gD1njUTtB
FoyGPfYiM5MBfA3PlV0dZsRzZjMMzCQ7fzyEqcuxFvkSg48kS+vH6G7AqArqVt0Df5+FIXEc+CkH
2t0maPqutzfutYO2juCJD49/giG2D8/3HYXX5y7IIJrP8VC3yv2W9S+9zUskrdBOE0wwwfHXOtKG
jN842u5g4SHNSbY3BB3PJ6GWWq9657NzRkjZLEUFE6L1/NVbBWRVc0IDnPGAdfYjYDCcMKoHYuHH
RQcW70d0X24xFKh9hGALxiAW0uXWYAejyMhztHCHUsH7EphnJ5dWRX2H9WEfQyXH/GCFRSjkhhIN
k2afCHvjbDhmSe5c1q4P905iSTjLts9V57HmhhBFXXVGlCXGNgPG3gyboFsDn7TONa1x6pPB9i2z
wJ7s7RS7xOlKiJsE3ds3mBCiflrZnm5ZtwmYZ7ON5EdTK+lsvoYRw2yldmidTJrqzcgwGlKF8AZe
IzJ1PhjNaGOjS4KG6WDPofcIIRUyjwMDZ0xEY35QQ05vyNyY5/S4GAaOyruE2fm1MLEoztUDOJX5
QwvgI1ojitdCiGIPBS9sHYPkW+4097xkyqbqF+r4daFPgHWdwwohbuo89fUHQ0h8QJbpeOISoGko
ondRAQSH6RW4mLC+xAXLk3dBSTmHGvtaIM9yar93OAVtSRidCVKMKcduThAAf9nq0yMN5V/2+KBW
jJDDve8A4WAQEeC4KBnpQxQUrEb7q1TAPjkw63OrXM2HJFwwL0QYbVylAy2aWwkVka33zknkWg0P
B4JkgKSunF+6hgOr4MjOcR7Lp/GgIdB2pqGNMwDjdQlND1UZaVttF942yQUb35efLM8f8Lk2o25U
6wMch2+BmANTJcQQslG2qi55W3NS9Sl735huDZh132ZAbtFk1JwjCZZEZTdDcwr9YL5sG3wXvlge
QUiiYr39iiFxg+pazsC1XcBpMwACOvpu9iCfu9H1w0RJ7Wlz8EsWSk1bmDQnG34G8xgYw2HcT4V5
Wk/XPHjYNgnZV9lEdZbwfLdUzNM9q0saO0egfpqmRPt4G/nwdzYSHb3DKQiS9RDuCHbsDWURrvKm
c9FxI4WNA+4gXUNXC/6JJonCGhx1UA/hQ9X2mCJogvr6JxyeDcXrWVAu8EAlUvfpQgSKHCME7SgT
57TrXs7o9Z8UOlTs/BW6idsPvcD9T0wZ78bvNtpYTekY5C0CZk3zHvmoKkwamUHEf7ibNgqU0VuB
K+Aljh8sLyRh/rhHGiOKy0LrW0d5sY5pcnBECo1Tjo0k4S4kSSW9YjfG4QRK98BifOpxLKWlksbV
ONCrSwrhYP8soSl7buWdwMSLR9PFoTM3zEo3WUO9Nbqkoz+k14ZykxUyvvn7LE/QknLOhVcIfFBe
oZZNpG/AzV0OQekesn/A5wkdEtIA1mPOLElsWACSEZZEbOG1zkWAyY5I7+ZuUl8QmWnUOPfJeNqK
uJshFpMdTc+E3/HAFOd7IlsejL2mAL1hZH3sknTfqxa4P4HAsC4pPjeyr/7dndAhHv6pVBLH5usS
iVyHIz12MmkdbdJvACwk0Dklg0Ztv0KiaSYrl34iTz+lGWFLnSTp7f2YO6CNEVEarlCdKVuPk+Rg
BCqAg6e48geDamHU7Wu3c3ZGAtcA0ZWs5e3Zz+VI0dP/g0ujOnDJc+UbeXLZ4468Ce8U9cgJ2xz4
tRr+LPoXzyDM7loJ9LBHw0Zxzhe1PArU+fkL8Ejm1q5HEXopXqcrQ4e0uXuNodqT2WVLXXsvCTO6
U/Bjrk3y7Tpi3lrzCC96n0rfk5yd+7j0D6pjDBPKnzsIUjNiKU1ak9nErbqiP54r34pTI818ZwJV
wktqQrwDw5xc/DRUyY5mlsL5Gh5iF5VuAYDiNpL91WNrmkI0Slvde6fz4/2hLkGAXd6uUULqTfp9
30uVEtNZi8Y5W6g2vUFIxOYv/hqbhWSJgxiIInciDDKowNaffFBQV5hSxEqJF+HATc1h3KAmRHbi
/aw77QwH1yF6lKajjd0QAOjHE217XeSWK3nVZcyV9uJUd1cTiH5hFIgvvhh1eA6shrErbQgwgB4M
lNPEcJOFXNG7zrYQ5z6MeMTkWlI5Jxhp/C8J0wWqypY1IFSuCdEomjH3/Kl9LuGKB+ZIX1RYUxOX
/JARIEv/JlttBxw8NBlqap0YXNN9aHUahVaFaReM3RbIwzX5PRvDgqPO58yFvOHGemQUF3Jc6Dsd
43N2wrIHG5tbxbNW72dt6//GMSCbFQYxueipnq/rdWvOZAfuGVfwH8jFxYtgPi/3HJAruHclCpAs
k9Nb0HWVnfz2uhMXc0PEuMnj7AS0PhabfVYi/IIzmefCa13x6O5iFZQv+q5xizf/xcZ0SE2Al9km
txVKSN80CLIw/B0SGcvqZExA1k6+fiBRJuTeTN5d8fhmNvZXw7plv1+fwx45EcikHdlEljawuqeQ
mfNK2AxHfeXnqhLdc0Yh7j1yN9HFUkDaz+LsXbOjwXeaGhO7Za5NV6IfFBrPzIAtjt/LvyfED/JS
Ddv6KOg8pNHTUIol1Fk6pPskElOTPgvOP6DcUi99RVpugcKtp1gyQnVN2lmLHFvUPQlmZrfrJo0J
VWfrq5Gy46NAE/qk4b3EFUYVNAe8YCSZsyq41h6c4ycSa2z8P7wSedH32wdX8jfuhj1SCKKJ8KBD
cUYusld5evlGE0sfocqEy0+NXpfGPbixNeIlN2k+R9RgpgkE4ASHPZFID/0c125oSXGz3pjIxEee
ZJ9gn1k73SUPJURYvhglJCbEo58fE5QUIMRIWntquycuBLjqWx2oKAVVIquM5gGJWLKHJOv1CmIN
9idU4qbuK/GsFm/+H5zob/SsUrVpgQEqYMOf2DnNsRNj3/jJGEKiF6IN8j6ajz+zbb2E0e/GE6Vf
4ND3qOOS6VqIutF77U9HM/ONVhHx9V6Gpb2DYcmbAqP/kGkdraaiY93r1k6zhwhVu89gXHRTfwi2
RGE1HJfTspJ57uWvfgBAIuWl3m/4Mbpg3T2IMyQTe5uAMgXwDazYhaoTgjViK5b+zKgLASLB9nCU
4ezg8sZfTlGBeEnforK5zwRBVkKtPIqRF03j3z8rgyFNjaCUudjTnng9SAmpBOD4+kh5mpaBRCeL
K92hrAUT+eytBeiJ8Ea0yw7J0jP/Uur9Tu29h5AeVGOdJ2GX2uHiYrHRlkN0ncp8Nd/936n7Rrg+
h9tQINs0hIa05oiY+9GyGWXG2+Ok6TWYtz3l4UNE91sMeWy9fUkCwcSZcFlaBEEolRu/IG9w6pkB
OROOFOIGzCjNLURTyomvB68H/TWTibNuyASUK3kO94eDYtmRhdcs8hqNL7OxacFL1c/xhuuaESa9
JnepJW53EdWTg/+iPzEC7Rb0nfBBfynaHCBchEpMhIGVAQ1b7sk+tB75KaBL0vB2Heo9pSFdG3t0
inulAeUrFLz8xrq8MTUMawZPBjlRpQxPF32szPNBoUHHeqpSI05mdyAzpYWW1R5sVj9HGG5r/p/x
Djg3Okyrq+Lsf0vO8LmVALrq7Ox2akhlt2p4pBTt2J8oR3Y63fgiixu0BlBEpqtnyksSzw6gFnML
1oDRKet2cKyb+StxD9Vs+Ed0yN4lfWn9HZJmq/R0bQuga0weLNvg39i3aO9hg/6I0teI8Blv6iJp
Dnm5fIaeiae21v5Qe6XGApYy6EHGLmvwa5VFLNHyoSJUSXAgZ8Y1gcHAbFd7lAnwO9hWMpkTG4RS
5FurN5At9Zji6gVcYPyf6z0M+Y3uj3yGKP1tIllvkC/vEff8fpJvOmkhP2QZnJhp8DWz4ni141WS
hZotOJ0TGjqwK0w2FyxKSDPaeVtNkyCfZtCrwi6yW2TVuv/mK4YKv15NYk5+O5peavyB6/4mgGwB
XOvunvce7BufnV5J5mkEyZ2IC5BLQrTN8EeRyHxRnGv0YOmv3gsGG87QHDFEj3HYnfL5iqGnVAOU
FIwP2V4uLnpw/LDp2XeC7HH2IlJolOHASailiB0CbbhJwHMB72FgQrGSHKuonbxOobbP9H5eXfbv
BE6Le8vS8SU6IHBV61igYc1zNw3551z8ErBW09H3usni/l95tBCJMf6o4IVmHaOU0s42poPCuHXJ
bKfiGW0qEZPJxJMbtS4IDhEb0gRYNLtGSFoIYqkacjgu+OWBRDtMPryf6rxpRF5SXlJ6zogowotO
8p9qsXBuUbWu4krEs4fx2GCUUFW5WAcHpyvsfdhoBIFG/98eG4r9nVwJR2A2FfLdHzOP+s1dDwTH
No3wL4OikMTkCJsRq5NJRp+5lwEna7CV0VToBWZR/+Q0D2W1OPHaSyn2KpCMGNjd4Ot8y44WQgyg
gMd+kLWatsPW9niF6lxDhC4Z0KaYzL6drHV7ovXVLDdwP13Szstf7bQlXiNBOtUcA0PK15ea/IS5
1jK2SxtDDStEiI4vx1OJgqpacLaExvz4I9ldXXo4ywPxk4djf1kJK+CDveHmgiB5H7rwWPLPl43Y
NlmYJAPcyuWH0piuWIrB34IysENYUSX/FFoh6nLVv3bDe6sKOBtZJASbIjTBlkpXSq4/4aI+egZB
nQKk26NqWr5MZ91oh8AFRHkzSjQe5cBhRxWxbWKHFlOkhzXgsLt887fqIDJm0mDQ8d3CSZ7RnMZA
QLWaqBg9pVShcvJQMgIjkNsdFaxIxAw1eFidAZ2NKk/+xlpdy7aYirMmQMF2woQIoRgqoCCHpogB
JuNVmqpBrwUcC0b/NlygQf5RAWvla+Rky2PGTR3k3xCX7q3fF2QrVAiw4BWu6ib/+/TOQKtvhUb5
EwqHTF4n9pjtdEYxx3CA3+MqJtL94jCer3MupscxsLuXTVRXWuZS09MNdH3wsVcvcetlP+nWNkKL
JMyys0Uu1S0qtr4tEyqD4JpuhmlklSuiGA9s8qkoAORv8psJcHU/+w11f6ePkoExGMGPaNDQ7W3Y
dpY6fNCGKADowauqbpav89sVukerqwqfV9gtpLsI2V/HBiR0SjQ8+N5c/pUy3oPmkt8IZvaw4ILP
hikKzAqwCkHuIwgnn57qtEtxK+BvR+Jk5HVCu/s1sgt9blx4ToP8UWBm+TbgKp7dRXWTO1jilUSs
PinSbHkeh67M+EIuzDyGovv4/j3a9eyiqvLDn6JZ0DaAXiQ+g/Zd+KvR+T3E0rNdtO8UdSGXjhJ6
x+8j62ZWLtP0qMgknxAon9vCqQKqNOEffR1vOuuTICmRaGZ6dPG3Rb8NVWZ+uLgB1oL0ssEOL3Zn
R6HUYLt/AV2z8lK9QtySB0mTc4dfm/bqG/9wwkerRCTW2lG/vnFWwTov+ypZWtWG2hhsE/CHAYZF
5IACRB3Ysi54HgD0Y1cexNqeCg6zCESX9aZBRQAGMjAJeeHuZkZqP02krUx5WUcY+1ZvQhi/FzTH
hvdObYFtC1QVc1XSAICT3z3Oou/d1QK8z7sEu3YYatUlFlqOcaIrMsLqosY1X38fuHqZjQDdKruw
vPLdjfwyFHlziEjts3Nim+RSwjEjVDWFB4Btiea9+2V5tM3dJA3fbvCsZgmAsYpK/KQ+tcpQlTTk
YykaVHrjRHK5UnTbJVx/XPfK5j0g1XC7jPlIqok1V9dfB+0BGXlpTe5XfNfi7tmGWAIn4juedpzB
kh4ZwCmYui3C5wb2slQG0AuAXLpCaCHyx1rC8JCZqfeA/yQZsXKIvvMWpSQQ+pUdDKghbMwIBezN
DDbiM4jVdKF+y6RAUn2D1Ft6bbGEUIGq2MRvDWWX6G0GBD1hXRU11+v2diyeLeDTyxoZTrVLoxR4
unybXp6i0GxGZwzZPbWyOwbyLYUEMR62DxHPpOJVRMdSrajbvGDNBJWuxJrnkni7ydCv0AWSYq8z
TS2YATcrYtfcCYCERqYt1moXk1Kr4KinKVmfXXFooc3TAPCVZU1u3CdA24IKIRUcsAMLH3CBtyrd
fL2E74BI/WtaXJ+orFUn57EtwEDwS1WOhQ1ISwE9tCEe2M+64bAj9EmP8Z3kJ7HHb+LuylQou2Er
pZ4Ul2O7Z+CiYs091o4/xCiVwydqDuEWJG7/ZlU1yR/M8rgKmyqOt0sF15k1CdTDZ7M107eHCPcP
IdNB/pzbhxnlt3wP6NuCnxipnWLxVH4NMwEkDy7+fYYpSaSABWtzvC4GzNSKMM9xbTTaWR0Nunk4
11SRCls7A+jkTFASm30yXZ7Z+2mCMh+p2Jz+T8eG8M7iUln2ei5iEZnuXbL1LYRUGUf2PeF6aoh7
Tl6lbqfOcU5fbdzdJkS/LdJkCE19gTVSGfQS0H9YEWZveIfjKNZgTAGTfwnI13D9pe1CQt8+rvPa
uoTCFWUbupakwZ5WvsqT+KciJ4PI7qqJ2oZ5d6eWNZYRsDCzld9Cqb5eVSgKXBEe+QEVJgCWzkb2
tljj18ZUdlgop7c3As6S8cmI9Apovq7r4z4IVY8EsHB9u6wqIudkeZppy1X/yOyhaSXnwDg3RH6t
t4I5QrfJTRfbEYjcVn9L/FaefHb4MvZ+ujxDKhqxE2m56vgPj8IxXDzGQu5kZrasbopsrBYqomfg
kQtIde/gcTZ6T1pQxEgXn6F4I4MFWRoYkWsb4QS1wNfIhiHstsaeHbeL5NVd5k2VMdX1jzzFGB7e
MRVBzurqCWQJmDnHMmclvM6aaRJ17KKElVOVytx7GnLM8vstr9KUtZBYWhFKpUcs2B0oj6l9dCc3
m3f+LXMdYmvmjcVIoB8RIrM0yOdAnTgntJ7q717rv7dhs3jynP0gy5ZGMampftJxJj08f0tA5h5O
1qq1byYcreTFR9m7c1nc04l1qHQU7xdR/ayf/IkiW8ROlb7+O/nfG9F8MXi5Y+k1uX5z78xrIAlh
0Sj14qS8XK6BT3bL853FjDs3A40tuTTGmBCMr1CKRRsBlhr5SlkC3sD/RL0Xb/dYaBFYygnu+c43
qe8yaNpa7kUxU02z50wnsm4k57UARY+Zzk//COCNBXF8sS03Uu0lVv15XJLvJLuKE1tjrspbwPuk
lTIrMM55qruqPb9V7TctVcKtq5OPBPerxwnDTmxQ+lex+O4jRyQwV90bqObQKtEG0XDIAsd5aCxT
g3L07wEPkZAXW3AvnM99fFcJFawbzvv++8lQB904v8Fbody8SauzZTVaS5yGQxiqk4aZhYj1ieNu
84mysdCz8V1zgq7h77DtFBgD0VYeMWcrAJ2NwQCnBRI81lKel2mVCRVyQQJ6BwTqFYNjboYufhdP
IWVYxXU3/4dxFDIEet3UIBTfMPWLKYoWqLXoYBgtvt9CBYUFqi9+BaaUc16PrxhDKjZKk/RR8hdR
WN08ylgcuB3oZFpq5pCNvNkFPNLFX2kwSRnKzzh0Ip9eqJFgREX/d+i1roiFaXyada7Uz5fyLDf5
odz8kPwNkwgrIag3fyBXD8e6JMrDj5zLWBUXWUqhTV+go/zBAZiBvUooaBm4QhhymTqIFffLTKbA
ignIcnW3ALNNiI90NB+tvc/V5Mli/UhKIUkgnAQT/pdIAIRFvSEulMWv45/rQPg4OleFjNoBZIJp
9b0Vs5/kim0FLqG0KkfyTIAutH2BQTNGLKI9df6OP99K6MvZc7wlu1+SuwQjTqEG7OSnJEStl25K
ALj6vPHBxp4ND31/P84Uv6iSccL2itqsvzsKwF8ybP3nP9oDMTYqusZwjqhJN8olbZYgtnWP7Y/M
2Vz0L7WeS8G+vgEZ5iKc2P+AiZ8B+iZwumyrsC3HheHgpB706QE8sxd18kSfvyjVPXd7LtVdl9/b
ad4RqA29tSUWGYnHdEihO0KrdvnGKEAGNGjfv3QXLGIM0VZJPxN9NrngjY4b1HhgbnsNbp0BiwFP
bM0NXzXIoS4s4sRlJaGOb+VhRlQ4AeJfrbGqR51JBLLSJYbsnOJIR53ppCNqB4+XEyNKmw7WamdZ
L6F/u0e5I7n1FyZzhgjT4T6q1DLJU6ImDye9iZj4GDNblGJ+OtJu7xmViXGV7VCrFj11Zmnh5q1k
qljKv0jlL0qOHd4iJBWY2ojTiSX5Y53ZYgaF4GlN88RMGqj9wS3uWzsU4docAq3GHXHeD0lJ1zdG
Q+w8urIKVguerW1xleuxZrD4bJLLTjLiZwsO3YO4c5OLfiW1SFJCDfVHtpp3cOuZkMamj13+yVqs
B6wQJtcRZWsvsobAbu21UG0dGt12wffKNm4cqImQlidlcpgWIwJFdPKdN87MjQU1/ARzmE1aXoC4
7Lc5CFNKTEZYVh51uG1iHu6gUGSOICgZioxvQkEHud2kXseWMIaNrlFVqGNr++795rN3rXmys3Ut
05p0dxiaMhrN/CPYNbi3QFpY+FqJos1xdH3rWnTogvyO11vRRUfq3JvzOt9YTmxixW8yF4edXfZ3
x3oseM1vGfTBc7cYwGnhzpVc5LfaFHNEKy9JSEui3xuuzVeJZbMJhbgy0Ooc5YlZAbX6HF5WcIyq
XudS0Jzq9bwBCo/g9d2V8EoXOaRztyNYEcdJifJzi1WbeEWVDYmf4/21O7veK35B1Q6d9NJywNWS
97APOMF/i5H89hZ27ZlhEuJnx6EyiGniv9XxWlHd3amm1YO7aLcH6biYIzf7EAc2owJ+DP7o9y3z
QWhgbSwvS7qaT1IUSca6b6yDlVOem4ChF262Xv01+RkuwHEWJUnV3E0SjM+vCFMJY9sfxZ0F0t/P
hcMofN660e6SlFTLm9UngFP9iVEN420EUvaJKS4iAz8CRLHOknDleGnX8V/Ou/jFtaOnmKxZTrng
QoD18hOnPmkQL8icwxUywqeXwZ7CxCmJSBPWLiDp9Z8qGD70bGlWobir0raSgZkbgSU9O3qbeJGQ
mrxA8nm0Salf6thfZwBSJnTJoEWVg9yke2vCFnzb1AHXEPKpVE0m2SGCZj398b/T3htGxWzgm4Qt
PX/PczbiCg66Gk6Zqkm7QsRtLFHdmBBun39KPtOE6vUxUlzSl2lxvEb0zAI+PebtngUZaotxyySs
mL5ZN2pTSYEvjj996ilrqKQjfjSA2AsVWbaDbKvaTlCxQrVpA2hwZQKYbMUfw97PBQcRvVd8jnfS
ywpvcR4XbDg7UDS03QuPTZsT0w5gOKb3DoEENk1VaEE2EqU+NvVMbxlGmgQHXC8GBoD4Lq/xqQpl
S8yyoC9dWXRfi7uLllSi1+YsRmA/UaZ7APiKUoNq++hAVex4bYbnO31oZgp91u+wWp4Q50Wxc9fK
SByYr8/R1caWejcuS7SxZk6v/saf2mNP5jTX14hS6EjpYoK+qWf/3YNS1cIeQC5jwQqWra1OaUEw
8O0LRv49TvdSGbeYt1Nh0jdkV7Ja7NXH8mJYcXfobGqIVQ4zMofGCbzYY56D8fAR/PxhQTdAnQu5
H9xHP0pCRpEFfaDp/BUM7EtsgT9jfqhdDAagdb27Tt7CFuNBIFctM52PbvjqAs5yFP4c9DjzBLAW
vGbyyAfYP2LAOpXYmF91t9MeBV8V10/BtcO2X2Se9KY0ox+UKPifACjUwAfcwOfjW7JccOltdMSM
vxRuEBRpW2+Ns3tbiOwuLo0axTFlt7ehPAMo5WLHBnd/7lEvN0dJAbZd8hDUEQ4ZJcA5aTnm7UUz
8sktKQz2HMlGGvHZihCy9TcrER4vmaEYrsDXvIeY1fFLDZzTtyRXMPLHU8TGQzr5rHWet+npGQ3v
IT0AMjuhOUgMA7iZYDGP1DSCP+aW/tQkonzwtuL0AeyhhEeEDBnMikLoNCt3AmkGajFg4LKtvQ4r
DAOxx8E8tT0keTGzsjjKm0upnEFRfVR/f5xdI5TEyqWMIYbrcUE+e5u7R/A+pWB1WPC/BhIJgd0o
MxlnN/QV0+/MtzALpS58TnxoMKKTgf34LP0gefQQ9CSZAgbAqs6V/bPF4DE4M7QPrZ87/E8ljNXB
mO/8/Lpa4XD3CvIfy3S7MKGKq9IH6B9Itr2AAz991mLdryeghinFqMnN5lyELi+pFEuH1Lw/Y075
vCjfRTjlqIXhxv5b95LjJRSfrgxptp2lvj6VArHAiPe6HihBeKd4uy8pr0uitBcKid0jXHDiSGyQ
mCmeTR7AvoJqvSKqhO59GX7RJJnqGsANThPRcdIn38M1gfsl+dHFEH0ueLC+x7/mR6KSkA0YnXBD
wMHjZqvXsEQvvev27A6g9khtbTFSPBVVR8zlcYzWlZz8vaoZJ2zP5LMh75LHHkA5asIrIGF6AsF2
xZLM0b7KQOks51YP3LmMTipD3CYEU3SwnzXc6MMy53LnEyVcStvVzEOy8XzSOxslXlQEZ9iP9gnM
dJDd9yEolay2CY/gXk9hTvSzK4tFzAptsY373HbgBUISwdWzS20zoNemkcyvCpP7Zh3un5rTX07j
vUj9UFrKAo4uXcyryRkIbnE+rPpXUDTb+/KURY/a0fVyvsAEOx5lR7Sl//Ce3zeNRuvNd1KdJBNI
JJpttnVebn+Ir+OCTSnfiYA3MIjBRc8Ww0YIt7vrHAXewgPrCsH1Yap74UG1SqfGTHe2zaqBp3Uq
5UtYJgOnU4K2wFOpi0VeVPth6gfXKDn5tUCtqWKEStIDBx8Gja4vQipE0noIBAVTzVK+xoMw4fif
5MFr4gmxBjKQZEdFiT7ZdPSX4OH51Ehn7wF5DPIZwXIb/dH8B9P2CnzkiCyotDMvfXyFZylemjIY
QxWfmXJS0QauI8F/bBuiQ5QQhXPJ6P0kPBjk1q8SdnCehdPsqv3iVcZf8nu1KMsBfWKyHYdWcVQB
MwhpVdbRo04PCtaVH5/SDxyCv+Svfg7ylL1GmMQ4iyHONS2C6mQkG2hT9Hr1wj9vIwKo2fAEnhuk
v1ZY58zyd6HVOroXue32/+vCNgw9Bu54vmuCve5psrGRjqtxnG01d1+/liOiH7nJ9FBoJMuJXQ9C
ZnQFm3TdnCViBxf9NLBdgGEDyTE/pHK/6XEgCP1hKfmNyKzo/xnBtlthjkI6Gk85IMCYnarreKer
UfAgIsRwfYMbzlBDD9Z1yPUaIn6Hyb5JJVmopBvjU6rm2EIVKqgbBuzZgLrDXBqdXb54aGbwjT2T
YPTJu1eqGtU2OCztmAFfWlgsHVoEWG1Xo8CbzpBiudSdMPRRX0Lp5OBd9Nauve/A+I82cGpQCRQb
UOM11UsH5EqfGW4//7S+ZjUnyCMY7pGs74YxPJX0MVQ39c9z4i+KGsqj7xlyuGj2QDjtSNJCMQZd
qrho98WbpdxZSnhBDePJeMFs7XlpcQSNLS4Oi3G/+WsH8SE6ro+xYF6a6BUxcl7eFl4p+defgjPN
R3aZdR7HdT8z96LNShpZ9pPgPiMQYpwgw6KhU/zndZfz0hD3AlGbgl+ACQb8xVkIXDAwdETBpDri
lAOc9K02k8xd57zOOq6/plGUspdLvxOhr3+J++dEqMX3yMGs+ZhjwEn/5VhxksPbGY9fh7I43CoA
nn/0N21KGwU2Zyv/nr9SYYnullN9Peb9WcCpaZLGWmcnKBwnCicJuoJQY30NeOKXi/9mRr8Wyo2D
YSLp38qxVmEdqAbvHKE2FnY7CWJMX1X8LjMHT+Z9EFddTBJCOOSvuiD6Jg8SQhqhRYktcnfepxty
4eDUAkNUarmEubVqoee9NJHdcE/1kJILIqeQc4YYohiNNc3SFML50LT6aQ+luAWuS0cQMgD1ng0d
2c/8UqmNsCefb27BbDMNZfxAuhhVSg9u84yIdvmASQd7paHsxItLsgFuSs8aJemBsOOaVHpTxM9b
QbAfuiqUuEF2nRwkiPlIN4f/V3mCq3M3x0GJSOOMGAimB+ErCJgUvIBOc4TJrRL+ipNUM2vEKLwS
3GFH/xKglaIKVQ9ywqHROhAzVEFphk6V8qa/LNnqIkYXBAKm830UMsXaRHNyDPLpKOKbt6Pp5T1W
Phz+fgQgArR0oo/8tbQA0HjzS1rpXXwTIkBqGEhb8Q6B2g4UWXp1HS4+YgtN6S1rDgaYLkO3XlQ6
qN7RxbdpjwzY5HdOZ4V0ylc+oPa74DAGXG8yymlHHo28Q38RwACV4nth8uy9QJl4LyccwT8kOlTo
FlF8GyLZeogGctTA3GjkFirrlUs1q+F4BklTxvQfJ5uc+/3bX2EAiy+GH1nB7B5cdmtaYjc9tMzF
GvKrrOAlt1uvdDhZfHXvGK8QbPp04X9+KF0M19SQg05+nYrDhCVX8KQYs/eDoSvYbGliefHYNxQL
f5siAUPEA3gxQd8SpJ41M4R9l8emGsFPoRTEMOpoRExuVma4V4z4p5HPYcLx1oO22h9S+beha2mW
VnszqpXuid3T0zOFB61YeMpnT0OggjLj6RNh1yizXdMyDpWn5aID7sWLBzo9NjXg4AwmXVLwmHRL
pbnfmXxI5zk3Nptz4CgKZ02VjSdJt/BYAGJtVSz2s0Kg7rf7Klji58E4PNwBaUw943QnJa/YBGr3
ZlOrhLVMFsGRbwzUhhxpFKiMxR/d37Hh7KKLM59DLJtTOK4U0m6K/Cg20G3vuNdyLSDr//NFlAZV
OF4XyCqrcuUF3nlZ98k5r8+rYs0rWy2xtJlr2BlE4UASwMJ/CUKW70suRBVE7oWlPY/Wit/60VPL
ULtytZ5yk5abtmo5v4bma0h1jLtg5GHTD0L3WhZKhiPY9pqNPr9FyoeR5bz4Ojs9yF5SKl7eSwqK
mDGIojECRVwO5pUWLVKxyE33haMytfGyYSZF3S8eVJeVv7J5qCqC++BCQdYdaxfZm28YTKMpsR2g
FDH9gdg69dcEcF+u4P4gDsbzAre++laIaM2s0wlxRcMlJ0j2XWfi5q+KK7T321gNSXB4oIB89pOF
6mLfR0GW4bdt/P8Rg3D6Hs8xTO3QGS8eY8wDSumxn7jg03vcEE9VWdOngF06ne4wLGhIXq7fnEmp
khIcFSkCjCOADQv1lOiQZX1mT4i6Mt8CUlH1Ko13/jZvgzGPENMwMs2sATTULI96rSTbCosoeo/Y
B/K2vYVk5S/tKh/5AmaP0rso6XoYgDHB18QucfSXyQm0sMt1xFHhYPMvc9PslGekeSqs0Q0mEpmB
pHxuqdEpGUtIX+SNBZll32btV3Kvmm30Is37cWdfmEM0q0W5C/klyUY/PQoPBHJTVy7E52EgEFvV
oRSNj4tikTh8ZML+DNBF
`protect end_protected
