��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$Rx�y�<��wA�*;�x���@�̦�W�X�fa�M-$u����n~�%���P�$��W��kYَ���P7�?UMfT��q�6�U��k�>����~�\N�(�����X�e���/6U|)�X2pF�]$h���d.���9E��WG��L�X"]�Ad����ľS���8od����e�GT?y	7�������ݵ�^��R�q^]�鍦�����s�ae���h��L��P_���ާ��YЭF���'\��68�b�[����w8�[X��V�F�0͘3����q諵�uW� �h�u\V�?@��_6G�_�*�G���B�絉�f������[�G��U&�����~�F��AׯK1�`c��[<��FY���4I� �#�G��x[X�=�Q1��`��R>(�w����R�O�?����7�,(�H\�#h(W�EH=�������yq��Ѿ��aF����:�U~m<|��.��0=�P/���4ǆ���T(���C��HL��
}�~�sswMVi� �aȑ��̜C�_yS�9�����w�b����Q����Cܵ�â�8 �h	���4Թ8�^E���(t�������`	��ׇ#jJ���X��TT=��!��cvT-8�B��kx����ni�+�/��.2׻H)Ȕ��};���)9a�ќD�T*/K�G�H�T5�& ��Qn�up%Dw߫�{Ad�&��9"��������d�qd,�
|������`W~=��|;I��~�Uh�#���W�òKr!���-G�� �1ʓƊ�Ԃ���Fb�PlN��y�~!��=/bK��5��
U�^��%�~<?��&��#�\~�ҙ0lQ�r���|3)⸢]��!Tc��H2J���uG�9gC�B�m.����3y�S(�U
�>Z��^����Ѳ����j2p���ou��-�Q��4�ڞ�(edzxr�u�h�ۓBG���?6}���]䊇���{"y8j�ι/���W(]N| ���^^������VaBv;ؾ�<��H
J���l������M�a$�X��>~5�HpIuXZA,��Q��l��]Ta�䓝�4��pFQ0_n�(�g���hs��q.(��E�N� ���ǂ��B�6ݵ,`���!z����=������.We�O�S6߷J��W���e��z�(�7�9mU�<y6���h�l�����&�������;�� �V��=J�����e�u�V�ʏ>�J2��8K5����ַ��{
��˭��fjk�rԟ���j�s�T�#�����FY�8�E7��b!�{�*��A�����aE%9,<mp���%�]�yަ�qТS�q���]TQW1���kht�PV`@�Me��R�/f�M9�>o@|ɑ�M�5��*��R.#�;��9��4MI��~�� j����w���$c�Q�<Q�{1C5^�k�7IΗB5�;�A%�
̝u�����ʺ�F:�]���^��z�X5kȰ��8�}<A�:u����_���+��4�����	=�V��<6�xw�9�t\�N��:��V�$����3��t�G����QPX��솕G�K�#�-�]i���������tr�ߧ� if5T1�k�I#Jds�0s�EbY+U���j���}�6#Ll�!ch�!��X������jբ�/W��K�<0�Y�6t�~H���0��?,BE����I��6��#F]C�t�Yw1�iq�,f�z��m�`�����? T;�5�9�`D��AmMq �6Ј�ok�,�n�޻�I��k,���[�㦢>�v��ӣ���8N��d��{m�w��l��V�G�(�i,*��y�Amх���c�Q�k�'�
�t��	�]A��Q3{Q�+Q����C��6�u���G�T�f�ҹ1�ɂH]@E6֑�Q*(g���kӿ��j���>���K#|�XU���˽:a�