-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
qDkAxLmjjNzIl+AVvI1FgHjU53dx2wBem5tPHop0c4vEjJrkbeSOEsHjflskE5/v5azQ2JeJ0+K8
5AiuKhHfdUk1W+LT54TfL2Uj3RcFJkbnr9HT3azeZFhrw03lNO/RJwTW+1Uk2K5V4jgKf7Q2O2y+
HqmzL7Az06GxdBvlXFwj2ezkFLxwehE/8guztlHlr1DeVuMDZVGGG0Vy9ncXYYz12tVOQwMQztqz
MunErcYGQyR59s4/8ZxXbhN4I8X7Ty2vax2Cz9zmiFfuEqIm3DAqJlLqts9o8DZxGPH4I+7mSJPT
hLowMTp3v4Tvx2/0apDkJnkM+xYPFRwDY001vg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 124960)
`protect data_block
9T9ArzL372LxAjnaaU0PY9QKSxdhxaY09ibEZEdZ3dyVoZIJGmKB4y5PsH6oyL9Srti5RwuZTzxS
ME7qCZqzr1qhB0GewUDwzFFZFCmL9cdZVcvDzYKyyL1KWo+3KwXVFPzwSVFQPQdEDWEU56JFerm9
RG8yajKNn6Pp3QmviatLtzLErNRf+4tnmx9Qcpez+CA156Jw75N3y0t30RKsac/Vt7CCW+Qjghsy
ZUuD3WKx65nOuhPsBs7HwsIUN2ZRR0tvTJQk7ARaVubVWGiO2+NIhTZhY+8bRcF3I/AOYsEhi6WO
f2LEk0TWWw7TIw9C/XV5Tlf1CCFQtXLXgq9PvWXVP32ImJ5PuCTYzVbQ4NqlgVwuouU7Ak4APUGN
0cLmmLOsDMEDWoFk+i71v6hC415Fn5HxdgDv3nkT9cFMYZf+5xvq9Wt3dYOkUfDUnuo9PD/BF8yL
nUBj+KEE1bsuNSdeVBQ0RDyCncXNtWbjpVxAVsVmyK+GUBJ4DCJYzycLd8gEZZnRfyVmy4yuFxJ0
0Igyr2sHuj7zCNseMU4RD9MXTjcUfa+yxkVtp03XCsByAbVi9OSSxYcECCt+rlIlKjxFPhdfv0hz
/0hl6V3OXvVouk52vg4yJhsC8iFSokyfSyF+Wy0nGqyGSezA6FUxulHWAbPYD9dqshOpRDKr2L43
RWYu/ZcsY4aWE/n4mfhQWAQfQo/tT2QfyL5m68iWzIr3zslx+lfaK5GvFZrE8L60iJc91NrifVln
3SW8rnw/iVSpR8I9HqovOOfor3MLXmAUU+1rpA2scYfzgXZ9CDk2p6iQAC1C178EG7T4lAIAFdy9
DK2HWClxVCTxMFvwCFoqmwaJA/Oz/rL31qZa5fiTs+Fc4a8h9siLxlFBXSe4v+W0dRW4YEzNXAYJ
D9T85W3i7U7+LpmaqBp5BbM1J28kA1X6pv2m8udGA0Y4ZFUM1pcDRUR31BeimNk2nkEsUo89Mz/X
feTrgbgax6r7iWUuqXrXmWXazqwGnUTyERqWpbvHnFXHQZ5/xHlVKPmIcwvPJEHNBXnrt6WDQkPo
f5aRsjwdcyGAtD40zCOGBcluJ0p6RuKyuQbGB7InsbHNuRfuwmyIkaMF32zenXI5CbRx5dFFvAVs
bejOtLxxjWuORi21/4wu0oYKz5UkTKYFkOCqClE7HK4N0Pwpi3+vjvlAViVOTFg6FpFtKXPZi8Be
Z2MmfGGmdQy/HCyxPSdmJUnb10trZEdi6PQh8O0SMOSCfrulVMjMe7nE0jJX9XCw7axXB0EOftgf
GFEMVhXKbGniSFQDQqZde2GaxaEdhqm604FPHXLLggDxmmMicPY7KVCgrUn4YbjpmD1GHUeWBzLY
v7aHFYefXFyqFSPka3k7nb1nLqGD786BODtqXwMm/fU9sZ6OAuSvuoGEj9/e5dHcyD94aFCUoFbp
2I1XZ/uLlRm7H6BVscugXhmEfu7SdzmDqeLu5GiOsGc1c3J/AUp6zyfcOcw7inMOP7RBExDQvG/f
RYgil5hapaPf/bm4DvpwU2p1LSaa0TCmR4nBZy2y9fKdI0u9XInYn0TumekeEuhURnUm8cCDaLdG
gbGO2ZS9TcxUSPGGs9GCaDPXWEXxjdt/tbYAlgA+kzPlN64s0CY6X6ayIcZjZgBhWR5rbU+vnZmr
MfsnIlhI7ezJ2d6THL4yAQQrFwRJWWx0r/fBiMIVPlTyQuMWeSBBVNh3uRBikyAAKNP+J0745MQI
UX3kcLB/u1Ycmyd3FiKj6v/gyhQRFt7qoZjHpsbY2LN7OYp+hk8tuP6cOjKdrsr1Ayz2mmd6XaHI
JtoeUeOMWcCZYg4nVB1eG17J1wndvsL6x9NC4QNW7wb7gWcicvJDKPlUbyLp9EXlB/JQuFIdIT8X
S62CZDHBND3Q7h0UTHIQNYc5mqcOCe4+50NH3cxA1n+GL3Qs4+50tivjij/g4A/DdF64n66MAL3i
8Oocie35a2AvZmPKFCrCUUWjYuKKfgy6WKbxVBGrv+98E0dopCFzp9B0Jagf7Mr5V0V+910b5Ou6
lbPxsIF6ewBW5nx9AHQbk/yBrsZC+/F9l4VLk9WCpoTR3yLbFc2Shh59GSLqs8FqDEyU2U4PzMlB
r0gO22DMp5Z9slQqCWqylddbyx2dawrqINrT1rNJOgrhjbMXpSdRJHKgACKt5EVkQIGOnptHukUy
PiUpvikR2PxDZmWdjIyKnZ1wWdXCHPFOO2Linz1nobnMDZ0/gToJg6XnuwWH6V6Y6iLZHEfRB1ST
n0qaLBP0/C42g/Vdq+P2R7c65D72EThdrkAaNHr4VcqZvStiitxGsEFSCH+Mv08qcDSzWwQwcCjA
4I+3TRuzfREYm0Hsw8bIMV6fzpl+Fmmu9mwFo1b0geyBU1Tdnw82alPWqqbCZ0aBe8ycyv2TU+9T
Y87/fzbA3VMg4zdEUr4J2x4F955+HAmfZoHvaHC56mwPc4Ilaga1W2Qe6TldVWOTeJwQ9S9XmCXc
IPnJo4mkzMAONnPfbgbAdnJRElukL1V8tY2ZXJH5qnH8ehReAQvxCvjD85z/yYe4jwShZwmm5HUr
RksMtSc1+P7SVN6ZQWhzdokjJZ0bnX6tWeYgp4KlMBA3Z8mEQOHa1AylpnxZDp/KYODFKX6WRlQ0
mMZhySyHmzLhlNvlCe8wvu87MJpunvM32G9NeXPyDzOnzJk+FW7eT503/yeOoL/AsOUKkK+Rsxhu
wpIkzGWBZkkyh8ouPINqsZCh9YYoDI+FZr8iiY+b1J3FVwAwJSywWe5Blod1yhmsZkIhSA2xonwN
b+RN+dj01HU+Eji7JwRH5kx2BtBTNBs8iYBF9cdMl3n931Jikao0pWFsihA9nTnN5i2W0A2WU35M
A7AY3xdpNJ0/m/FHXZgRAlzVlhZ4Jw5AGN4BSsytBVUl7dZ7Cg+hEW0yXi2S1oclVvAE4sVdc8UR
KYuhISkUN3gBKUvTU9GglAyAuUKzGejj3255VIVHzLknOXjObOrHMx/JIENwro4k5Chdz9zjS1Wr
9RZPa/4DNepMf/phoHBAwJjbm+OjheaOquLz6kQUsy/k1pH2LJ/Ne+bJiAuFLTU5JA4dExIKUWhg
c0jySsdeVT6Pwiv2EMm/sQNMwAiYrR7OPYmURbQTzfHvW4bBYcyZVAwhZCv9P/QYtwcIf1GkJM9r
R9eTf36PCdTE+Xr5kr2vOe8ry91jdfFyQzZoFlvYf+wMDf97aDCEJG01/egE97d878yB0VShcA+6
0+oLnqYrWo9mBoHJWwHkIN8kMFiJwP3BwAb2CcYOPV7T9WnKB1jQ+XUODnJ8Us7Z2ncZwQQkRWhb
euQGHh2zsnOVv/5i/yMw+CX+G2G+kByKgaSrY9PGTvb/H12xEUOBq97x9AoTKivSjXagMAzYFzbs
Xt8/tA9I4T7Dc3FcQXr4CW9+4xtlX/pgV01ap0idMTFJxlsLE9kz6+hJ+ckuPY3jBUJ/ObTfTrol
UieKfuaz5whco0mhMFtUsRKBV5XI99nLooiYBoDbO/ZHJ9vQg82Fx0MuOD/2CcUGBvM9hA8Zsg9d
IX3uHEmku2ocN7jgM3VJYqyRJxb4cCFpVAyDWQ1YNV6A4qUeARiE8bT0RY2EIec+/aK+v/OAEa7a
LnRP6UXV/UrDlxPXk73Rz/JipPgDommNQ7XOKzIUcmSU4gvbFsmMRQ0w7IBjBrQBdnfB+kVRcNrB
GknLi0ouzrXeQK+IIvWKIIAZMkLiaScjQm9ZLXBOiibz7mdslnmI+8WaeCXz0WhVCsqP4PAmkvhN
bCyCvROwbIqSpZbeo1Z2EA6DMXNRmvYFt85b+5Xb+u93dFvPw2zh8NU4XwnDCpCY61woVlW6Z5kv
/0D93rzgXjg6EHo5YPlF5RWCpMpW/K4C7Gems7rvH309G72eknw5e2bxFyPZYqz1/tc2J3KFOelQ
kCNNYs9dOFUuGw6PdXk1KZZHWtUrsHKpeSB44t7a5VBYfRCmNZQcDFwQU3aYaiSzrpkCQI9PQ6Lf
c5zILnWTy1e5J9tBtEjnIJm10VqJWI4lAOIIZtngY7JTBunMdH9fOH07AF9TZheTzhnyA1jQUgRX
TyMNDyzDA15LnVo7utUJ0xJ9IngR5AvY3w76/MjMkOJXY34mE1zAV4o2qBUyHFxNT4EOk56cK7jg
RHbRXwxIn4WEnJRtl+TR0aZgC/O/ICbQ/VpRvSn6qlAFO9y6mfT+QxI7xh9PweEyFAAJdFbClRMc
5zWOeYyOJgCQnNybcodxInTebDlf8u6wu2oyQy7xn6JrSzUJK/Z6+681gIwndXdjXVfhU5lZZg/v
3sUH/pui00lIaP6uSt9Kk9rvebMdtVJ2pNmIl6e9JIHopR83VjlBXeOEu36Yv26uS+gVpB1gbqp6
Mq7ZS11Yxf5Ea2VBgyaIVriWYqdqjjN0Hzr8HpCtTivjb07xHfmG0XxLXuFGWGgT7ZpXi0sf4V4i
BHBkZpvIpkGCnqmOcYnw5/oKFOWQ3/EWw/kCZ+blLzm81IgTROgSIlHA0u+PlBWEVZsBEzAQ01rB
ZO5P7wb+LRIfOxPqNYCLclntnm4Ok6fQ+YOfmY2uLn7GaStyPuIfxlDoS0KTUpr3NLLgOKjWMuAI
7QVtMF9HSv2/F9VIANKL+Dm2ZZTTlT6u9Me6Fcz/tQhtssQpqbUdCmkJdYSo9Fn0CSfOWEh5uEOq
s33xvUFReq2//lUChnY6f8nQyq0bdRxvu7Rjrq77G6QFeFcntkdknxbkTUCq+CyQvc2vNARp1+Jo
cMa1VGas/hJaM7S9OxfMpme7Ft+wKGIiAxffDhlfAltcTngmyx72isw/8xmWEl7GAENrdz6b3kve
xsPoEcXrivhELumAdND5i90Yk00JZmOFmfz2kxJ9JqI7dWiPWACAs6AUXh2hwfA/tUbG8a+7rs13
vnfw2Ra6qB4m0gItpfdiY8oASlv2pzxawFNJiFJbZT1xSRohaiJDakHzXgd32k8DFjg2QuaMcsel
kZ7z1SuVq8K/EMmiAPoIGMEHHyLsFpGh38JArBFec3TteTmFWO0sKvb/s8E0uyM46XQoXsYYAkJV
dYNuQOz4+rM6vDYmQB8+24Irn2qXdhYJY5bfLU9pU745b0/lwScXyXvEuQ025NAch2AK3FD+WfY9
ErbD4F3R/wzGNLfFfeAQ2Mc85eZBwqegYTGnpA/VDjfUmJZeES7u5nRSeafv77w3CUobp59W02pv
O0mg/3L81zwE/evJiRkxuzTEU/JFKY1O4oDhau2InhPBLDm7PuGPW+Z64bUETD8+C65UTGDESKW3
lGNe7YpgWE+Gi6MXP3KLT6yypdFtNnuO55m+fQdWjo8mv81GZQob1KwEEG6eAyR80TNjv3GuhmVp
w74FnEa9Llagi+bGaQRmgfsHoFtSnEVSv4ZwmeEoTgs9d3wbeFvM2/WM2lDpnPHzZ6Qsmc2IwyLC
YqMcXWNdLhvyYSaAEUgfP8bhubnU+Giu98eDqDOakn+Hw/nzcKzVeP9loiVIXWv/DdwdUZoasjTS
IQYa4h8lAFDO8iEDuMvWaqWEEX7ASS1t195ZMt21MrisqM4mJsG7HYCtjao0mMvG+2bF8baWx56E
/oMqRbwf9vXmtuLf55FBaY71TbesB650ynJmLwoS/Ky1+oBftIjKnqnmA+PJBDx8qvlAk3fhq6Rs
vFAdvgKag/+zgVbBUa5UhMhRecWkZyyF5gU2Cg7NRIR5JX4A9X0FvV5iwCa0gs4O4oPKGtIFEGHQ
XC2snU+9kyMcCaxtaOWF5agBWyVmSMWzubc6T2vluh6FwVrPIqdd/huiFeNxxskaQR1r7VZU71XU
bLoW9UbMDx14wxmqmChfghvTaw/vmyy8A3EYKvc4HBWeaYOVsM8WAM1daPyQh9rO3E7EgeYf+i7X
LGj4GHKzAIU351pTPorZhrKBBgifPG47FwjqpvaSp2+w0lWVXHANYXCCZmsaUIECd9b3zfUQlwWZ
ZcmVCvdxbdr+wGJpb0hpsSTtr8VM26YWe7Uw+nETIPiepcuyc8KPo2UdWBKmi3ZT9caqQB2Jl9P4
EOsXFRMv5sQHC7CIfRn3x394pYe7B/9eM/I/CRM8mHiC1quYjbWE7MzTAum9NVgKem3W3cIOD31S
PY3q7HGambouczKG3PJmtOp8UJKRksYh0N8z/PN9WBqtqEBdbwM5HnFKiZKxfQfd+qErH8sa+N70
5Oz+Cg3GUrYRTosyplDk45/4eGre23DF9DsRL8YL5VCe4csDfE3Q9alATx0/a7J2fG1w/5chqXdO
8UjpHP0JlGi3YXqeWLmn7UsrMsPfADgg/9+pDyqcLfWanK72KrVknIiRyFmLbw6og6X96w/JjerT
FqdhC2dWbShwsLuUiG1gOI4DpC1vfxADAj9SLcjs1pU8oKXmdSeRGS/fRaILI5HtCA/aC5/F7f0t
oGOO2Eb+BBxh2e8GDVOPfe3RC1+LRCiv9/n3f5tc86RwoWsVYzzY0jtE2NWBqzi69GvKxV+LpNv/
0xQBmI0ObEZ85yZDRW/k+9vRWqYK76jjRWFHFzZ1X0tXfrcf1oLRdcNokBQJFuZ6SGX0ImkwSPSL
MfbSloeE6Or9BGojJcXJiTh2YYc0wB12Z2PoX4/0ZeSg0DmgRzkvqTJWNTGJXmK0/2xj2prpDn5q
AS969GTbSUZ7+Igtk4JrCu0MnTNEhjN7/UFlSAXQQTAKl8Fp01U8nidqFyBkoORvel8i9CDtZlIj
LEHHXdFRd6QhZg/OMyVPliKu6N/Uc3xns1spezu1ZaNC35btDJbOP7hzgvf8Up5e77d2AUYHftKa
6TxPmX6XcPTAuoyTUTVXTZaADBArUuRzTna+s82ljhe5NnbuVSeH1014D3U/1KDvN67YQFyr1To5
CvN81CJ6gGmtRofDb5Exvide5woW8FVpClA1eQeu6NSZ4bKTlLfUYY2Sxo4twx1VMWUAOr9p9HMw
3ConSTywiuRo0qf1DrA43s9Zst1htby4xoy88mHeMR7bssViwPaA4EO5nFsWKnJFYQAsDYKJAWp/
hiHcK/HYPd+CTTGrSDybavic/+3ysCBgcPjWHEQ3Nx1b5XS2+Uwe50sbmeJg20Z2+TyUYoWufo9D
a4C4VCuPvL9EtgPGdR5mGluFS89gAXaW/VQTzpJdYL0jvZZDeagYbyAgh3IRiYBqxtU2+pZVaQyD
kOO5v9KkigoJzIbJ0aDyu0zq15P0LNO2L4h9UFUXjPyRKL20xbzMaeaey30i3W0yyy0xlQoMOP1y
L9pQxFk+egs5eTf3hYGB9291Ai76DbGLvhfvVyuCjTR3w6ovrbnTBMqhBuY8KThmh5IXIH9ciD8R
9ST/8MhLZwkzxhWo3h3LsAcNVt4LwSy0f55RvELilIdwwhZmX2aBLvhf+9HvlSCO0OhQfd5bbdQ7
AbOUb9CnVzZGTuvHyHNxCYJ2yIaH+Th68Rs1rwlNNaZWTH7cI8gpPFnuzQRinthczbz+mNa07ACj
R82SJYOH0JEBB6B8gSJr99E7ecD4qytIE6+h9aacWqeNmzSJR+wA9rKUtvEdVQaInhN17nIxl0If
aA3jLE6L6kbwf+eq+W8rxTfJI3bN9U2d64Y8Tf8QwfNN1iIrQwWk5pARcfk5VhBUxIgwXXaOFSeA
Q+4BLqYeSaVV78Z2QLQ44FLZHMW6dA4FI+v6t7TfhxaVABxaZKih+j0SUdohT8GeLrh9SQj1ALCx
e0RlcRN862Yq08AMYJH+DyC8B3lkuVtyCS9QSn4BCZkoGPhqcKplh38JYw+PNWr0TwxlSoXhuJLs
69bjxF8D0yWV0zp6GLCBiN1FX762oco+Pj88KDmChVGiOO5mHypP7Gb5UOJGNuAjxcN3/tfGdwMO
y/5BESlWnwmqoKsucsyPyjRmzZD4ECpp4JWWIYt1f4Jh59p153xW0fXfH4rCIemN1OxIS0yPjz3P
cyzVrtXAuntcYjm35U4j2cf7ZjftGIQG4zN3gvwnkginutP8aGyrsJ5rU2z3Xl3XODHA3Bt0bt3e
2avM+zVA4/PqJlXxEjJZxYjBiQb/qfz1P5v4uYAD9e087YUiY601WGEVfIRdWkc5mCwds3r5/eye
/vAeIK8HoOHdMtIDv/roN/X+BsL37zwYmWugUyxhfNsO0JrfUKT0gCPjfHrwJsTrHgbBDwmhv9oJ
GywkcZQnx8VUWFBXC6hGzGNLxjT1wv3ILg0JJ1lXb3W62wLuJ0nBuHz5yy4r87o04qX1RMgBXC2q
YYhDzTxTFl2HZrFs5RQgAn/KkOV6mWi3OmuqdYgBknYalOwQR6eHxslgI/g3hoR7vyYPek2pLWCQ
qdDWri4UKMPSYP+OPyY5FfO6j0sYQa2LRXOEiTFfXHwIHDoEugiuPpEnaIMzov7P2m2RU778uDs2
qzMkGKmelY/KqNk9gF7CNsuy/eWaJzPy3IK39GCJw6vmqdqljJqkeiSFkmJVs6RO6APZblKEWzUc
/IRuoWwDOl7MgV4tvPfij00YJ1UvuyT+DDFY8BKvAmYjhgW9HUiJla6psGEHJ9/qE1ScNiqJ4ZcW
XShocxrOU/dy9bvzXmdrf+TOxZlrAxfkjce6E7yAU9Sp2GALaIHDuP4HG/mHeElaHixnE/eHfwW4
vP5fxDhc8A2er5o7ZUQBtYPpCKry0MQIuphRmwpKi6MJjM6L8Jb/uTfaa95bErZ8EWF49fxdCsWK
0bkRVRA0P252ZIGLBl0QX+F8XM0Pvm0qwmLYKoAn80aq54Nz/iJjzmBao4TDsDrHkKQWtcE5JLuS
K0hUyeVunUo7I1zFT4yXzQwVOFpXe7cC6mb9gsIsQblS+PNShdDSUn7BWnH5ZC8p0cq8J8yK7+Gn
+aVc84AryhaC4b00rdQhsATkDGGuhRTKwGiH0dU+yXF/W6eC8b3VfId3Bv+PlMTHgdrX4fMdjNa3
uuRT21OD3F1wL4eWKY98PNPDl3Auxz74laQgeRfLjlIQa9odLzzLDTCd24lLuE5GM+R4/aPGMtyA
/YZyKJ2bpFte5uA9WdJUmGBw+QDdbc8S7mYcnp/ByO9JSmmAlqZQITP3l+YD9L9RyCS8HXwIM7bj
i9q7OYSqSg2Cs8yUUZMYZcofju/xTHSqtQOLQhdttMc/J3NxqCi7UDCRC0stVZWwnWUhg7fCrwEP
eEoBj6u9Go7h8+hs95AYFEeqdb919V/NaaR3oA2NdbTElkkwYFrBCWfWdEzVDoGPdXLIkGNMoPv2
8lX9N0J1pDwu93NN+mPRxl7BU1m1DP5tdSE7dteSGP1nc97UUSV04KjZwNxSS4JsNVOdTKXhEEPe
LWX/HEnH6YVBc17JJcbznThs1WmPAy8lj0DoRF0pBizutkQcUBpW4E5X5eL/qqlh5a5kUX5pmyYt
PrIMB3MZvozFtYyd22WiPhcfUUZO1xFODuteb5WVMUtBFgEoln/5Kfd3MLLr3af4U8eMNq4fmIWl
gxXgrrMYIhGsqSIzhdgbNEazf8v1gKPox+soVY/gOtjxdiaB7LGX6lajPVlSxmfrei2ts/z33lR6
/mz51KvA/x1YyW1h8wfzx7RRHD2LRnWB/Z+8pVUiEGN27fXezJ2JaO7iCYq2pTOeuKjaHF/EDfAb
/1LHfgX7lMCkJ/cn3b/HDlw/lwtU7Pt5XWhRoWXupFmHoKclkjzCcWPykX1n/6ZBznsT0/Z/fpGX
HCttwwcaWsDdmmCl416puSxIT7WR+YQ43gjZ3Idvm77X0wEsP2Pbb8rAXE/FKOEnXdb1bkXz7eHh
FgqrFJp8mIG31FcBccr2G9kP42D2BAoFVIw6QfIcLFQlgIswd9kJdflzaEIbpe6kl9W4RfIQqd75
1Nn6BZG8kjgJ7GcB6Qh2t6B19XbwbI4l0x63eLNVIx4OiwQ+3jQDfi4MxwGzRbNBdBVP25J7SD/r
5fTmPDm63wi4jWx7IxzMf8T5NuPcTLWhN+xnJTcBsU8sv73ng1yHhYWmQHBJ9NgTWsCET0kgOorN
1uMlcGTfCAU9Ro67J2qgkHnjpmjtQU8g4J9X0RRLTjJTOkBXqDM8WCIPbsmrjb/5mOB717MB3cZw
0L+siqjkpbXcGekmztMQ2xBz/R07/9S9naNAz5tdsh8ySavTe0g5SRaQRm3x6CvDWgJOYptE3+JM
J+W33Flq2NCAd5JNIDSZ6C3pvp/CzVSDU7rOlohGuY7c1LB3MUp52bW87VCf5pZdNl3YIPW1FxKd
XatDG2KPN40nERrCAcBt/QnR7LZyJPq1zTc6VP0VT2nTZ5oT9Or4GMr7dlnTh2Hm0Dua/unFyjY7
O+F9AEpdQztCaPv7XO5vj6j75llp2N0jk/XSs8vPDP3mqbUWLk946DjDzDErcfv+9vnRB3QXji9Q
Z1Kp9ztGmxZcFNXxHK6k0WiixcvoDcsJouqN7Z+NaorLcAkog+Qjl29K0zc5T4ynfkzJ7iNQI/tX
zYhRGQR+c9rOEyGLgN5pjkFUhlvuYPTt0oRH6ZtrRMGDZWzkGIaFBWTv8GXeCY7axwF4/f/icVNM
Ia+GmFMq2YX7EVZIxxISbX91kc/gfRXJFwzSdm45r/n66IHVclanGSv30r510/Hb9O1HePqmXr6F
pfGY/KETwaGgQE4DdR8TCA0KVu5SB0Gat4Bd6OVS9tG8FOo6TBW1Yuozxghrj593txF+U4f6LqjP
muDLmTtxOs0C5n/KzbvTGjyJGTCtsN0OK1zn7qKflqTWkkQgIcn7upRAkwOLMuqbAPsxqXyKy9Cd
sNskAtz8YlR5CQJbB4p2mN2GkU+kZcoB2mxJ5HB2wVybe09vgG4jCOOsFOGHYo0rcKkkJ1R2pZNE
DTQf1GyoW9/UhGvC2yim91BY4wpXokD9yuzjrnkifsmyZWOL23xa14g7X5TINUzMsTY2v/zYr11V
12W2fgr+ouHRpB1dBiyxu0J1zwJ1tZyAW89SuJbhIgXvVdsow5CBqQkUAPmSbuOEvV5Jv10BVZO/
CDBM1vmXSL3q5oN2wPpmJ4o/YkhPpvC1EdtaaUqiW/mVeJBVIzFEVcgydRK2hhR7mHJFXAcWkILR
jRKrGX08iU4nL14YA92ORtZvgOm9URQE4uilFKVNn+0NoI0i4TeLo+t8H0dZ24UjdpL6MfZGiSWZ
dzlPNiQhbS93bFBsS28+IcsgVI9X3TWb1IW56QmBb8OlRo7BrTjOrsH+k4/SWb65POY3wh37fdOb
AHj8LoSCPmmirVlNx5sSGqfUTZLVB+vIisHX2nOaIAf/aNU+aAFRa4RWfBAnG/TOuGxdd+LHWhvw
yUiPt+C9Z/mXI15+vJtowrjj2JakyiLI7unDkkptMEGFm9RXSLutub4I6FDyiyjjjbtsSSaOWNID
N13Dz1A9vnnyMkWxKSUjLb5k9WjPigtlMmlHZcykOhQGxWSF1nBP7cwbiKU8RT0PcJVKni0pbWE4
uHCP62+5VZOCxIJWWe04mfXmqYpZHYyBIS38dDskonSwi5oGlcEZ7MWuXuDKWeiKuinfSq1iTKgp
2hJ65vsFX2cVBeH+/0lJBn7GNo5Bl8OxIYBIg/pUtWs0uZWztE9rr4kaJrIfptK/6SVi4nqf3na9
AFcn5k2QoKgLMOcqgF2pMstGL4WMAZkFry0Vg6H43CXKRArg+U7bxROqVUTLYF6O5yviCqLOj+Z0
BRHvov0roK160TY1AtIfCgrI2uCVknSBduZS0LCKMkvJEteUn/JPbxsUNdO90XzJ1md0Ahqx1wtp
Th84qTCZPtxhyWSrpdt6WOq3hhrmdVjpn1xrMNbfoh7mOkc17LsrUlxITn8D4FZMPAxi/5jpl+ir
d+jGuI87XjwnCbCf14/Q4y50N16l3RjO3BA/qUcmKbnm1H+/LR3a7EdCgH/eEtqe7auPgEH88LJT
Q2/uhOlpettEaJPloxWGryjObx2iYPPebNw9PLIoYOLVe/11oNb2hOaaETtLJHcfb2/lv+YRidRX
/83q91RfMwk+Ucy0BLW1Ck5EJFrGrxMLJc9oUmr2IYID7+21lJn9BNOFmYwyXTy5r8YbEuVQJ6cl
GepKEZtPwzTLYzYgjrwBGOw9u4vmo1POkiCMSskqfasaJY+upgpTY+icQ36peyENUzT12th78EGB
Y0LBpt5kwZxawrYFizWl7C4RA83ydxdiUrJRkOygAm9DJlNpg8dvqm8SK98rRf3KaihwsWpoU1jg
j08TinSIEz1qaATrh0WqNV+454cBsETDnyZ9Lium7cUNy7rIwbOBkTM+LrTae3K2rftgXLx2KWTd
1Wt7h/rdtGDXZ8vEWWa2ZxadYXeNIfUAnL+EMPgkxRqUGttfrrmYX3bWcHUtm3/K7XMr4oQvI+He
UiP3VZecCe8+pOjRhsVJbaBBR58SHN/wG5IOMI50muJSRtVYxMOV7a3HkCHwyAA55mkYEn3SzUih
fd8Ks0teldynyg68K6srNzFml8hTGzNr9Z5Y5QX92DZiKI6836qopV75I0iTIuy92P+TgkGrYXve
WztwZZt4H+YMPTVMssxW6P9PSSyQgGdypGsJQgmZL0Y+QYM/fxvuO5TCEoEqUhMu+e0s6avnAtqR
CDCId6oXX+ZajFYSVzJ9K832fuxk4WrQTEbEgVwL2Swg50Fefs5RllfkQ7IPr+UShBOQNp3dScvx
iQQjRhDeYtmx/6NTNSUW2maqZSMyX3XPH7Os/Rdn7rvloxSuSoKE43zSvFnYXGH3Zc3vdVZyOUI3
RePAseOu3XKJejZWTspZrWSgKTkKasyQyTYKpUUa8a5FfaIeR3AVtPU0xv2jCKLOH9whpUo7ZmVd
i8uWlUPuKOzuifru5FICHOBEHA6SqGsgmCkyMImlZ4FHFVI2RPpOiZaIp6EKjO0FlIAiofkiZmLP
lSjHI27qbAN+E00L4fb00lY7FY5XQ+9srWM2ODxFdq8PW/mlRyZuxCpNurtAC2niMYUrsZiZQKFy
VaMaMsf2KlzxKXM9AeEGX8FTAZsQa+crlO90DLoJWwQ3xljtnx1BetJtmMFUGQ461brJppffhWGF
ERqk3fggHuFJ3po0pEQS77h5qVytTt94D2RQihhrglTWuGCK/zK+EKr+FZF0iTVIS5UdqveBLiXm
tiThyNjDaX0fFkDJFtISOkjsfE50jwq5yAniI7lHixbibay31P3E7rNOJgyqbpYCQQXldfs6MVo+
XN0Yo/9phEO6cDUF2eOu5DxQkPPeGPXHhIRo/C/W8tY9+j28UJpzZ+e7Yk1SjdD2cSbFIhf32JV3
SoDOAxFovfHsbpcqzweBxgC6Kucc4rPZO4nd/plpRUGgWmhRNzGO/x9lx5E7u/7cY2GrRKDRHvGJ
gCJmlxC4U6SED2PDsm598irykMihvp850Cx+lzm47UoZ76cbS/OCIBzgfRhPFZZPEMTdm5VA6x3R
0O9BhzU5YAoRj8t9vbfFd9ISuFFkoapoEB++tQSypaLP2pFTGYDrPQTbppmzjhmA/+XYrd2MIh5e
fR7DR5ECg/KvtB60xIcFNdvVmB0tgov6FtK+2yrWm2PdDISOH1ycnzIqH7EfTX8PrWUJMYiklb5Y
MDdfTAODbpmJlh3r5VtcJQqyoYl7sruxxfniR0hI+L9Zz7THogER6etIqUPHWwNVrBMMYitS9yFx
gBqJhyXnxcjPizSObqF2Q/aDntsH3QytxfJrwOf8ZZd9fby0RUm8+48JZ93/kJ6RFunNSQqM/eKN
uqgpAKkUZEUv6C6j60FzcLlCGPSKVOfQBdZn23/ygX++wVGmeDURJ1/yKTHMhBIR9p2/xMlLgq+q
hp1/7bzQSCcnFHcCThwR6/NOL/nFm3s6RUG/udZa2FFPcLeiyJjRYtuMBCzJpgFza5E2NyT8a8a8
4BzfDSBD32HBjCE+MR4PYpKeQfPIzZHlM2ehWIsGCH8zeNcXe8GUPAyqzhFMCu9xE6uR/mU7oTU8
ywS5PJDFkktduZMYAiNns+i+pGNqw3CpA8Zk598V5eSxQaTs/CSPIm8g194/iWG3s7FtBsQrk+62
Npsr6LacWdUffO1LI4uOD5SWO5goAYQvLpqn313QdB7NEvAp0Pxq7r1xWF/wMUx8yUQRoVztBbnA
pXDwYNW12v2vXbxfm/A4GYgDm8uIiEn3VszDkgqxb171YMlOcodniki/YCM86WxuflsDHD3Yl71v
Hs/DXb1qdpDjjfEMkycqemmbUl6qA1uzZd7AOh+c0+JQlUybg2A7zlxq9nvUCUBMQIITTYAlWWKe
oygIWtPtLbn4pb2kbQ46+7/0pitEcEWOY8ArnMd58LwLZlUPq6SYmJfK1jPUlskUSbLT5jgczedU
o0QSsSRTwlL0ly64dx3keRSSuMUxkoVg/Md+NWedNSTHLDJc0svcfnsUoqnxcEjsyciWyKii8vdP
cBDg3HEGE57jtBqNCMqYhx5WCIGaoeukV8cmXtVyEvmPY+ev1tAeG6JtAJcoYjudbPDVrcETA13+
IbmIlFE+FXXmmi+yjOJuIMQCK+XtwnTqfdQeWSVjsdClj/XvymLYibnssMrkLBM1SSyl/IlYbCLF
Fj8SgcfASlc0mhBDHvZzzJkR9CN1Z8mlhNWgK0Vj8F/4L1PSrFmxUbx4KqTVGODlAa142jK2xl9F
NdN/20m0xkBiiySm0OhCa3w1AvG1KlTD2Ik0vwBnpF7/wTxm82niyDK0fBeQNqcDYtLUzVGZsGGh
kX43VerMmVH7hIoy2yzh2cDEYdG7jsTS4izmxrdxa+kTCraP3UZsnalwfIzEbcmP6ai1bn6GT1H2
P0VrClELxC7muYUlztNqUs9/IiM5hPGb7ZtKBf+HRELphuP9WV+EfPko9ftQ7wM7CA+tMo+JJZbe
0vuSans8YT0PzqpShdxyGhsde7klorTRi94gFp+rJCDOOEQRNh4hMW6faGUb0WDOZ+/K93Qxzx2K
0KsmcFX7ybxXBgxs3ICqJyCyaOmJyWN6jb8C5wsYxxVAa/6bQhxLYGpc3Drd5ChCOeRaRI1tVvlG
wrgapyu3FRImIBwZ4dYDltlyHdS3XZ8dtO0c1Ch8vDJhUgCgPzMu3iMUHsbo46rnZnbsi44wiY2u
yhOD/hfweGvD0P/Kia7utokh9DiHcjcvbmznarzh11WOjQBERm78Hfzhd1u3fuaJ/Mq41vVUjXZC
UCLzAfbd0XIyJqTKKjeDQzeHgntqJ0Xyq27LAXpZfo4yhMrDMPbNbYZUsy+TrvQrLigROLxqgU5x
CGGDEUu0yDE6rM3WBpTmYK6xPUFaLAM4ity7mKcfeX9vikvxf4ocJr8YEzIIzK1Wy5QlpNXOaukG
NpitQ0n5Dh02Ih/krXNS8Q/ljujJM0/Dx9LADBbHZ6Rbk//oWkO/+NS6j6DkB9REvRzGemoV5MvW
T5zdsPBLh5LcBKX40AI1rHXMs9hi6nX0+FlSdiWtgau9iE7RlS9Kq9id90L1npUOLK2a6e76BrFx
FtJpQrNp8BOzJEWXL1xgHJcmDcgfnA/d8YqsHm19AJ5oB/exRlhTATWcRNzMRg+nAvEDvdkO40xv
qsajXfCuYIub+/W40IztuVBte7uE1PfYnbn7gr3/DF+ySTTNQGU7XUpA432NQGK5aUY2qODJ30yK
l0SWHv/2w/nQGYp7LM0PdHMdEqIMypXxpF0QXuQb96UE8mvf5vph3JcyPcniVSL3z82MzYKf4pIl
KMSM5Yyc41Q3ueL3cdrwYTNEBvGCDG+eAqOAsyT5w+hw6+nqa/aek+pJxMJRLRnCmM/YCVicuhxY
jJ0drMfCPisR4vgxzr0IeKLp/AoidBK3c12gK8cM3mBX160/z7RTuN6Qkh56VrD/LPkSmHmyvZem
5RzgC5VvyRCPbdVLdSp9kJQlbm11PGib87S3Mva6Nd/pRU8ajSbx4ENDuZJndYqW2kLC5RqlK1Nd
eM8AoVeh4uhbhfh9SE3Y4pJbGaq17X+qHCCFvUwpQ/iG6AnsQTcwPjNVZKIo2vkc/KBXpX+hjwNm
TuAqBV8blQbeCtAV/l7x9BDQ7ZTWvbyC1Y3KkHTaVh8Jz3S0kY2jI29xeQQfoMtq3rLxwT4+cRbH
oqr0F94yBAxe+ycSPPqMR70PwYVkPDCBZpMdd0clZT2qXxI7OvroZa60yFbwkbpKhnGOSlCW0BD8
/ha1ELgC5UlY88eSSOuaQWIdVaYz4gUC66Qb7Xm0/fgXL0kenEooHOJrdbre8RKS22+A8OBZlfb+
f0C7FIxU3L4HyiQQJQ8EE4lvJiGJngOcrMfR6VUwZZqGIbhX1pcD3kS1PZ/f7MlkKfXOd04qRN5F
bW6rOPtdkYOZrerPrso/aVdlLSW2XuMtwjebEZuOhLsIfKbPsyjQZbFaaZHoH0qoY8r53X4+c7Vr
Y4z5DVBmdco0lYIwpfz5pfGUPQl/UfSWDxLzajMtZ3YaklQpIvEzpZrUBopxyuVOzc6CVqs7FcFn
ih7BjRG3DMPp2d9IMonIR5CYeCbvuhJTxqPMFgQjYWlwe886McXpwI3KSYFLkN3QmHMu9tq9k7Ew
bkB4C5iAmtIeByBK0SVyunHrfYPsDFNtOpqF3YgGhTqUJMqPasd+0F03EMN5gy6swipib8ROlDee
H9I67IwLSpIpSZ2xeAFY3aPhxQy2STUPqLqyxH+dMOB0VUjDlvq1utfV2o2mZEbsS3sKgmgIl4p3
IDT9q49wummp5RsrlZohUJfQQRwGYirSg7xk8hNG1hVr6+WrUgb/qvvUl0jRNrRrbguUuCPyHXKN
7MNzuuHTNerd66t5SOE9zVpkYw3s/D+n2ZXBSKQGGQnMZdBPJz/xPOJez0hZJHcI07mLdSRceYHP
I1U/Z9ZdmwPJHxuMYqpG/D3O6J94OXwf8h+OHUVze3XXDQw/7xpr69QTpl/QS453JksD5AOTvG6H
ibY86pZuZpz2BK0vqBQQWXhc4E1PJye3VKlrjcOC0JqUPK5mHjca+JpQ4YvuXJdELbv61sLoRq4k
V4w6exMiHKlVuVm1N68ilC+khD2Gvp/dq9TVJpEhIF/8vUN1whFlQ3fuzywaCEXJ6zYKwh3PHODA
4WClElgqw3NMXLWu4gqqYJvP6qJ4JSxRhhT9b3aW9U+Mkr90kZIEzlOd22/gQcU17Jowp5LnAmDt
oLlSINONIXCO/Qb5RQQcLAref87rqH9N4faTjnUltEmHx+rGRjq/DhzmBPnoOe+yXhNLmVoHSVRy
nxhVn62Tqryu2B6+CdzjfiJit9f7tuWQaUc2f02qFCoOr/uVlAeQ0bSg6HUQVtGzBdxfmD9hTbmU
b6SKdo4hqNm3x3bTkwS0GB2iWF1sObwyyddh1yO/3HgjDuh5Q+j/m/ZFsMuRoPGBTkAYA5OyQ+fC
TxOSWHeNoUIqqbnK1VPi87/ZZECSDekRUm/MZlk3WEBth1juLtQ3zAAfvXeL6GrBrr66KXw6Hl6G
yWaainSj2FB3bf1ATfwW5eXNu66rp8DB2nazzamh147C+L07PU/iGBBk7WMYyfHKQulE5zN8rGad
ZJgiF/LSFwztfGg/Ke6QGImQMu5QP2XhYV5DWA30Rz2KKQb2ErPknl+YoPUWA8Upq6i3zwlGs4fW
uAjR/I+6cGXvwVix9rb5+UXpU55gBqg49sPcAnFXoWluMNlf/z4FcBWe+3aaT4NW9w+rzIvbh52M
poZeyLGodVlTMGcmif4hrj/lNMNZDNaZc/mGORYey4YtsYUCc7DaPWTuFqgAOZZVY59L2ZPAU3+t
DE9H5Ryi4ooZjkFADIaURXlYNBSuu/spzbqfAWpsbH+TuwUElhJwMAtMvt4Du6Yc8UCI1JXBIXGr
ZuwfoAZVa53oPZqH/lqQxcu8gPoHbu9bGvk7Z+OvuiEcHGjOOBSRG9oVmJCNAOGyi+h5tFZWDyO5
oeIixPLa1KoaGZ2ZyaxgTHIEeM3dZiNoqQNSh7cfD1tK2HmQD32K6v3E3LJjzMD25L5tP4u4uh/v
Z4yEd/KClruGJq9kW5zG3WnVel7evIrn3FGBGEKfqhBU4nIqj/3FFtYKRFtnWeiRKPhPTixksfMM
uI+jhHOcDqMBOJneosa4eYAjUpWM7GXaNXCjy4iTZ9FxhBdTqk8a06p7fveoK5M6e6D9NKkQxyOR
gXBy+Fwq8lIH2M2gxk5BnrOjrDhLEjqVR/rn7faCz0rITJQkl4vnZQofzekD6QvEA/2baeasi8Vq
YeYrxdHUeQr/3/XiRXDqqd4JC3axzB9I/fwy4X8wb8Kl6eNSrCDTH5ozfoDtxtevd1ughE9uz8aa
qJSuDH8LJj181bTAg9Rtpxgs/pilMA+JdOkJne4VRTf3E51jUurSEJPX+ECYJxDY1C6UEJRfbJRp
6SrVEIGhag4d6m5mITO3QcZjri1VbqJo/7PXVKICuOPjEa3D/2a+VLgKSphg8H94cU3RmWvh2INm
C1cRS+1w+AHdzNIIlY9YSh81ZjJy6Jq24G9baKU1QzpU8h1LBI4ZGI+GoCaaOsIzzYS1R/JG8bTq
tjJFFl3Lug9pcuYeiGTaAR78n2VDr8FVxxPZN/4Y8qOc03VxwKy7M2pYEVppsUe0L9rtqslkVrWQ
TblxADhe1xc9lgXgTVP5+33rKG1GGU3b62kcjkFLnBWsc2iv5Q72Y3l8fSGxTOHl0KLHKURnS0az
ULYLbGoLcmJYtJvZHW1nf89mVFbUkFzZgvTNwhB2pJ2He/5cFCQxKcKls+dJklMsabk6jom+/AwL
7bM/NZ4Z6q5By9JbTXdChOtainjC5TjaxfAWyXBZFpU1aX9vtKRW6VEHiK3jvdUuB7FaoLBE4s4s
dnLaVYpZZc3rma8N0mvzpYK6axAaotlSNxtAQYJQt/lBLgWQmFNhVi3qISrx42aq77xS94sF87q0
gT3TNNPmK4S4TK+mWtq5/ekRqklDd+oQx3cxprW3B8A6hKit151QH+OPWbApBKakWRr/X53IsmxN
qgJAjCOTafK8GD7jczC73uSRHsHjtmjSOLYnqmVK+mxU0pNdjG+b/9PnOqf47ba4hF8K85x8ul65
c6UKZwbLjIMEL0M/HBZxEggoT+aaUZIqYl1LedK/h9oi2tkAa8D2dXttOHIR0JR0t6tfWmraG3k2
+vgd7I9Vzhno1VxHNktsJyBuimPH6CGt71bruKYITQeWof9bH0qku8AEo6ymqeTfmWwTDQQ2JGOb
AuM7j5fWZwI8I6aHCyqrmOlceYkOe3+vOpF3Zh+bLd/nTsUfHkNjyGZ1YUxr28yqQmNOoqrBwWf+
lxW/GJtTHbBf3z+dg3zy9TP3QfyxU37bDabw188SU+WE1ymD27Kz7RgdMBrUS41zjJTWcjRQLUZ5
ZdBZ8irH0raxx85w77lEc4vjAwxsq5vp8K6tqOxYd/wMqVSGXppfzPnGHS/ZOHm56H4poM2F9KGC
T94vMpRcltbz9Xe8NqHaKY/DKFhiZRU9YeOn6cpkmXK3AXP6Rovt60LbNCO+SiJ94f5xiwTB1WHo
P4qkIyjKQCmlLN65JLzopQ2l9LlYGR9vCnOHQ0PL5uvmsdP4Rgs8bWttr7EHvEynkqxDnkR418Iy
b/H8AklUO9XmjLD1M0bqW42ZDcTvTP4qmsx8mlNTwaOKZ1p85pSy+bI3PbVKtBG/2n6mkaC6Rxsw
k6cEEVp3zx3w/pASOhpzZq6Wr+6QFZ5rV48YjmdktJBhUe6owyRwSP4ckrcSXpYu69zMI2BLoGVM
3YJouHSuJ+fj4ccIfwHBmZfnoXJLLxi3UEPjqDzkJwcNliCa01qjNm4aCGfBC9L9Ppwf/FErg91p
hAsA4yFPF4gOd41J1zDzLpozfP1X/EkTv0Czyhk3owVgEjpUvC8pzVi4R8Le7Ua2WWMssGpI5jVB
qczjOzzk+Xj7mpsD5HCE0dKe2/lwLQGM5CswFTdZfYIHkQrPXsZ9Zul848McszcaHgF5itKhgfQV
UvgVFVrYKAofuJe44j+/D0QECEyWpM46wSC1oU6PA7cNY8OubeHlGmMa2bo9h/Xxc7IZTfNvp9Y0
4QBOfipyrcQmrmhgYatNNRLEeA8FNYyXdRhRHTKwzBPg+yJWHQ+EqDdP5KVSPwR5aXw6qMtCqeU3
xsjWMKXz2ILAYAc75vxHqWx/vxtIXjm2Oj/g0hdd1EYQuK5/rDVCBZhUFQuvnkQxX7Wyrq32LcP4
HCgROiHuT8pg73gL1jz5lJzYaj/FD/eXWcRAE3RnOQj2EhabIymHyWZkRwAiNBi/z/JSY+hiihJX
zvfVW4RtjO0QUSdJhmnD3Hr+oizV7m76wncscimpDXP5IK1yXD7L8A3K2TxFlWkVzBkfaxKmTt9x
oFO1dnps3EZTNSSTmAkZEieAOmxBNHVaXvTksJpkXWO3OvFCgyjCpPVp2oVm8241QhmyAxeQUtF1
bnCN+d1Jl93a8/3Judsv8ju0h0Dcc+HXrJg9htbbwo3Qhf6ePWFbbrXdLjxGBYdwoQCiN7nQHMrL
1BKIHoCuku6ziWIo5lba2AR0t/sCVavm1l42zKc1iuF9qKOJdFSv6tLXiHaiUghHO6CVDCEzYCAm
LkyBTHKNK44QxR98+uKxkcHZGAifFKNFeMrbS+WeAnHpsYpe66jZu6Eqs/18wHt8oyc3El89OfE4
Lgu9qc2cxghjNUW17maizIugTqtqw1SzgCZl+pUzbq41BU0cb27zeKJumfHUkgagoLry9Z6bVY1/
+k9aTvX4ipNkOpsBQRYcM6+uZcceWfw3XNXgDduLbD16ovAENoMAhteeP7zc2WIH3PgcNVOMKcy9
WE4jAF1ecIlohtu/HtIULRMclNJMEPrxuLMHwYwf9I9yqmtXSxtVy0mXLZWRaq8UJz4cRx7B8giE
pCvyCjXJSKalXkGS4qqLzvkWRbHGXMJWOrrYdVWzC/ePgXs70lHLg2PUd8ADycPDYWHtngWKPK1w
bj/vAW2XVLnai7W1Urw4jTsFwgyOJvraAP/ikHCWlM1tWk7gLo6OMOQc5+4OYhf1qHwzDr++zN1G
uCFfcJElfSYr74+8tL+v4h8eaaNmOnE9rapLCPnpWgRtC29gKtuy6b6AIJq4xrstNZSKFDs84iN8
ZIhF599YWIpP35iIO7PmfBZ2jak3zAIRnpJCc5dATuQ/Jz4B0Za1oOH7w1Zn1VKg5kqym1MyON+n
kP5UPfJwrvDHGDva1lUFtNQjbiotiJvH656xfCRb6YDi0PIDaWSYzbrF8+Rk7m3pnltER/SRM2g9
QHWYwRVDuZXEyzepH8+kiKYRElTNuPXVpU25vab4oyWUZJUN3tHGuOu3a1HlF/eqlN1BbhB78qG9
GJbU9xsqlkiOfIvesQ67ZbzoNPrmrM3gxMtmyd5p6Gt4lrlPg14RqmWUjv6+BSpZ7JyTflGqGN/D
TZc0aqpaLDgtV9wEaH+/j62Vx6oFrQGFYExFgvRrOdgl8wS3izL8/tvcB7/dTq6xloWi5uQWeu1J
zszAWzv2ATmq0uIpjlSYBYimilIKxZ9M6sxl5tYW57QsAzt50OB1jm7WdLuqP6GtzLwWjOJ7U2z2
5WT1W2OMLXfdVTBWWcx6/CvkTsoRcdqDxL7NzINtXs6UO3zm9+0v5q1Vd9JhYidwo/mX3HJ+cWAr
mH8NrUUH58pT1zaLuPqqFH3gUReLoLbV2qFNsrHMLmNYL5Makdi/fCja512ueqy6s0XzBWUl9+Np
nLEwLQMjhBQZ7XukHbDpMyCz5YXLE0xABoKBVh3dhl7jAnVvH21pkb4F674I7yup+GWnWU1i+Grr
7IlFyj2UF7SItg/WThzYN0f3FBO94162soEv3ZEMe7cN0QQOKSVpK7da734R9jEe5mOkSdsAPrJn
uFM6JbWSe1PIlqzz3G6Q4SITFrT2s/pAW0GUfeUcJdcGnNWgKB0dLZJlAnEBMxm/A/CrucH8CV2R
Ypb4XnyilhDniv5wGxWlXubsliaz7s7kWEDZedmnVm/Fx/oRMRQoJHeBcy/108E5kkdibmXNThif
Z5v+V5xya23oBylX5qDkMkfQh1A5HIhIE7xbweZ75fD4GBwbuuN75Sr3AOv952jqwBY2Iqu/bV98
sn/Zq3xOHz0oOV8/aSPATabLX1UAPmhAjvroppc6TzEYKWa6up7Mm2TToI0N0J8txxbvt1QOOFIT
CQAxj3ivalqViUyxSgtP4GV2GI9jwlMEkwascGsq9LcBLN7OmFuX1Qt1TO8SZtJxlkpProkKIrbz
zcDohAOetFq/jgl6yrZaIO+rEFu21MDZt0pfs+ucjnS767HKb1io8SOtsFngtMg2pHAL+P4SzNsn
jhsUrGx560Zbu4Zsv6cQv9Q+BYKo9n6LEeKeIy3zy4t0sTCjXKa02OiQU4zyjhkBe0479NF9WgYL
YriHpsNhr8HiPM05jdbNkdzOBjyuKidX5UO65Ns7jWKmDjN0n+JVgmH7lGx3pDxkcJXOVFSK3uId
Who5BB5JpFBRusA9n1plxDkxjYMe5F3OHWWflGD3YbgHTlmCusqgpQBXNGG10F+7FVPsfo8q04yS
CN0VM70PJm53ntH51q0cKXP1mnhu0fkrAPVaTus7jOvZ7aSq+Xho5dmGJg183DGRCj3fO+fS9A+p
8VaqPSY3xJF8Hj5sMTSS9Sog8Vk4rJg/kMkR1hasRsH278aMZ60zIso1EMoLRUEnxvo7XkfPkhu9
2TC3zpj1c0yFym/sYwaOEpu3v9Ee0TNwy1feINOZDRjSMPvz7qhHhG487eGw04hKb04bcRyJ8y1G
XfmAevUZS8mQE3VE8KQubJ8HL6evrw0xgo22x9UvCWzUVDqANaCjXMk0n/mkO8IBRZKpEK++8eYY
wmP/FzdfEwgxeYr/IBrd4T42KuIkCStHe/2jIP6kQhT94N+RA5czXixMiRs+TJqzVStk9tehLRcq
0J463DY+oIQdFHSf1qJu6awgK+0LadMdlYk7JtCtDTflNz2bqKnqqB4RBmCYHXpgLqq/sKG1BhZm
CdRn7CZ6vZmZBqGXUCOI0nNSBog6k6GSyaTrCYqCcAgBsb1c54k0FxZpnRmzzhZ3uLoLxXsYiUhd
JC4Zy/TyiI+SLgxk3/M7pq/LZxxFiJ7IMpucEBw4CH9AJok0Ns6a2QUH6dafb1yk99RfTJpr2FIb
vZqLWWPlUL3w3QheGspoQDe6XrV9W3UeCUZLTqofNC5gUKmALfOz9QdB5+oUN28ujhiouDC5GBaL
V14yLkaCsCTKqrKJnlOw56p4P64C2IeRVfAITt5NyYHDir8eHOyeeoOCX5N7ogswSOb84nPbKkqY
+ACRvr9wkHTOMEoOjZ1jXsSutMbTCNQqkQBOQqAad4B1/Zu36PLMBVP+xwJK6Qe5A6E8JnNqzdQa
IDNYe/HRdKX7C2SLLJuN6mCkO6HVWOwwU4i8Tk1a3Y44N7us78Eddt80iVGOB3c6mBtkCw5xBHR2
rh8AxOh1kjEfRo4mkffj7y3uyDv52tQW3JSZIb4A1V13CUE1O1JE++aZRHOyjVOsFHkZeDEkKR5Y
7thKS17I9OV3rkIWONoe3tU8HARLqz6mOwlooVtV76nYbXqaHVQXM8UwjPAua96wAwRYGK3vKGjU
IrWBCCjjYhyv0B8SRooAmyh6o5Rg/4KsR7DWngC6RLW5ryYaSyqL/tVlT6/69Igifl5l2N74zlr4
SLT473gViXomN8AT5xGn5VcE/yJWmHdVTltVdtZjDW+zCKwGOzHjjjilhYSWIdsQpTyLG7t+Ciwr
AqkrIq1eJ8AeHlSvMwsVhI4inmXSSUUD9N5I9/GUK8wiMJaZJveUftLgRA7OiO7y3B8V2dwaHVxm
AKUX4zRQeyxPvLFeDX1ZNcktO0tXYO/2euOI4BXQQPBM2ej93h+UMkJ5D0rWug7jZN8LwdEjz8UI
8LHEw/cKvxjAgiFfe5RoN7cI4uKdzAcAjSJJrL5189dq8lpOr+wuln/8pBF03t9rRCmpjbWvbvjF
j/re9cvhcm9NkITT//hIawhhk2n2STEtXsMKknSPl2F82Ig+QnOWQV0TVd9DKirCsySoBUz9FKlP
Da/ChN3rWfUP7hP5b7B/ORL1APFCrXPasYvgnZtPvMGBBHXQdiWCVrAkBAzxAhXC0r68ED5v7X0d
Dg98eTQkp8ohypMAtohWYP/c9vKqnxkdSwsXDUgemfFlfANY22ufiAgt5tu3oa+HBfhDj1SiCQKn
dUbJhpLy3pwTqbcMA8xpY1WukdbrtR5QEg+CdEVH8cMbqVnEHzK0eDBXi/ZVgNloltru/VBVgJ4X
P78+zm5uGKJTuKp46ZJzs8PrI7sVdi2eFoXrDu/gxNg04Gw7GeLm781gZ8G1EWnGBF8yMr6rn/aT
sY8FdGqu6TwHjXAOqv2O2U3yMAOrNdfU0J4MyFUopqHXlM+2YI5L/meoDvf84Mx9Zh5ZRYrto5+Q
vPvBUdMrZD234bvxtCyx60lebRjrxxn2VRlJNHMj/HFKNBDO7XqB4+wMBZz7z63C5zOE7BgkjDCf
mTty9BBKQ7CQmdivYtN17YzL6NpZLWA0mcpLtWu7XJOocTf0okom7m5TnMIPjeyMPaRxP0TDlWIM
1QgKADj9z+LyeiQ578R3kazhBc5BWN6XSd06LxKkpIFCV45RrJQwCAI1BIiNhET5h8I9XHV9rgMf
/HmwqjvkptM4GNGwNDHqdfkMrQX9qO162Fy+UDqx+e7kCanQEDAsk93z+UA6a+R+vOTNwR/YWne2
YEcyEnkrIFw63c/0F/NrhGcGc62NTAKn2snniCwtDTT4ew6DYLEjjq+OT3H1vs1H8janzf4CoZMv
G8v0UQRcGb6iP4oPRKBElrMY2CaFBjclhIzQtYyuBNepwOYEpsiQbN3AWWYBpLtcLlzJOzgCjnS3
AHTLbQXiaKSPG1hCFJx8wqdWKp4ZgjSq0NEIOK7MgJ06X/LzMezIhOyS1vtF2yA3fqFl4EfSLDAb
BoiaNYhIw1c7QOxBG/RFwNBO4D/6336Dl1xNY0xPyRPSAw5qKfOxuhMZjyzKqW67iHEHaMFLAyAb
bjUUGjVHA7ToE350Ju4mOh+5PxVAgdw/pMuG9xPA5DfUXyeNVlowMceObcdzZ/AbWTDRspXt7MM3
/QQa+UaSFhFWHO20wRI9pT3JhxYU3GUXCfP0xTVKkQL2BQFAarXQSIAmNG99wMVpb9GJlnRhogVC
+PFfuwtSycQa66WAmO1GrzocuIA+RykssuFfi6OUI4wJRfPKD/rOKV+ZCiYsWgX5YEf8YF81dzg1
NSiv+bIvPRhMwg8OWT3ipqKp7wrkosiyNOOm4E9zdjpPb8ad0m2n2rpXaHu5HjGWL6SYL0JMQL//
PwHpiO0ErDalsaHqVzt6OThb1YkbRIG8DvKqob2I6wTRmJazC3q3weZf/prjZ1ehnzg7GujVEau9
e3GX82jznlXFLbTUS1wNek3SXMMbkDO7A4B55FuI2yjrjmaIDBJ7F23AOYxdX0mchnlq3kzCZVph
98eAGXwdQ7qQX4NK7+Kk+HvfUEVDJot5dQ4dfzymn+PxD/EY4D++DnvvZpAotEqf/3Zt50PN3Vts
wRO5re4Ck+w0Q/MN5eC3b13tRwc13UOklv2+nKUR1T7L2dBy80WVStmLqN+2g3WBPcaTeqAn0wna
sIG4qhbGqaWFWI5D16tuC7Qk7F5B2rUKq3Qgo+yMQvhAfAs0M4xsEAV96Sa2B6nGWm5/4pOUUMro
LTyqaiFt7Strcdl651gC10kpXwdxS4sr/EyRho6K7AvPeoYGwXoGfAjkx2aoAamcL7gops5ompIT
GwsxbbJbdIXkXF72bLI/SxRw8jSeHx/6tt41VpOcAMHUYfyQBjGjKBA1OGZbIof1gOMbpRngMHBa
cgUdt8J6na5/QQ4EeuwhydY4iXX2/MyMGFXuKfkpX8aYCDvJkGq3btoG1M71ikxIu0CWbOpS/8ER
wRXRg7b5WMYto9ijj/XBWtYypG7mriX0wUBMdx6MfZVuh9BUHxBHcvyhTj1cxYvIX1VspZKT8K+k
gYADKEmqm+/1JAyMa18ZHRaHKCtC1S66zUTdVZhdM8bGoPEgi8aml5DStzVH5hIvapsVehM34N0E
92COXU5Me1EvpgdyP1ZKWNSffm787I8oS/DjdZIrQiVwVxK13xAXWbyKKzjYZvFvhm8/TD1X4BSp
Cx+0ep/uMOQOUwFlS4fzUJqyCPb2ImKW6ZCDhvzmm2gt7AOH7HoB5zlG4dg1gMtsrgt6F1RrO/xT
owjEj3q/EniNAkQqoa4X/5DH3m1MmTwyirGJOhpWPSHd+dWICXLWBt5qW8hICZV0OZ9PN50s2uoJ
XCoce/ta/AamwZfSEgs7auAlcan2Tixs2pCRYx06SnjCC3KcETc2JQUkWVd8s0EF+CcYJb1Xe2KA
G0J9z+u0+OghoXZWsiss1ta33a7NVGlJv76gtz4ZM6TaatBqyjOXQaRxbZcrmDeu9MYhn+Fon7BY
lNSSx0dY4vANUHww9eYtvYB+DdoR98tBb2Eg+BX+xLb3JGa9pBtERHEmpl/KxyIidPZAJ7C1+rcL
iqxIsg1HyC2DbgIdapFcWHaO07Cv2b8PrM+pMeTAj4c+4WrQji3AVjpUwX3IxzvWed9HQNHXEZiV
Icq5otaIS96YCYO2EGd3WrMm7uIBEcXRB2t27NJ2Cy8LUIYF7MGKZIKmKYkPBYTkTMwYHWpjatPZ
+4X7NQ7/8VX9c4WrU7nmaZTFRsZQch4mqbdGrdkNpisX15FzrYSNH/w639hT6YHu4NIOHObdkXLR
heVSgys62Hm1nkXUGf/Qrl4RNVHzv+FGa9JjU+ioj/GoMHsQnXOHk6AKyy/1QGwx7eB3inmVQmC6
h/A/hImPszb+9uhC1KLDExtJNb4g/ClHZhQ0sGk3Yg0VvP1YVRZTSC2pQ+Hfdm1FqV6F0jBXE4Kd
9dWDUCCZaeSjiYuB0rP6RJ3b9axqR+RZG+qCTuNs3yftbRi69TgntF5PrdBQSG9DvwjlY42o944m
XEgl0Xj6TuCOSOMEbXllE2qeM4O6WS/g/NWNKRHTC4jiDB9ZxA1GlVQ4f7pdHbSeK5vftM/Poifo
qe+gOSiXoZRod9eBUZMsJhgqDS8KEgH71auen/rboR/pbfbSamSM10Xb1mt+S50pRWTUTZ/6MFGf
GZPxadJTeuNYJAYe3vwMxK2FXMT2dnzLRpBLaUPP/XENEZIlhip12sPJ2nCsOCjV/6U4eY9VzYKw
mE2ACvX3b8wSmVizuKuM0Ucmxo6j7+ThM2hE9vMuCBvQwrqkk3yYpRJbWi3BcHfm9T2tSy/hgUI/
HLGx1vguOxkycuY5VgGQ39sRc0+6QzNCXWymxKaiI2j+IJy758mWsv8lU6IVvvKaFFRcneEiA7Fn
NMctS93RmrDtye71AeuLmVrfGaTjUdqjwOwaJSC2Ipa7V4MW59c/cuySdd3LFv/mc4jEX7IdhVPr
ijUPuVTecMd70801hvAODxOLCOh0tZX+CjZJXQHbJC3AY6RE1fIi1OYE9zzGI3mo+P7lFiqf2C6l
WwGId9su5ht7cDY6OhJx6Io7GOJoiFBcUp2xB+b4H22MkrCmFGNgBQNf3YFWhmq+4uf107Iz2M1/
0RhvQEQX2Vu1C1mSvBys9BpUcOfld+XsMQOBqFh+jvOvQtIexHY0fb9Ca6XGpLc/io6VRd/kX396
YEglgqy5RGUdmxmjMkUiRLYYswQwdNOhUTxkejJz74bEYzli8rxHbCzYjWIlQCGxjK+7Cr7opbk3
5Z7MYex/ego2dZZKbZeEBpRyWipC4Aftxz3xsu7CyGSvGTECMsSXuzKIIRHJJlNh6vFT6ZIdFMrM
TzquPyXaJKcqMIJdwF4haPSQa8uaqgLW0O9zOCN16CdGg3lsxuHlQTFKlS+Hn0+bI1JPGzfKK1Uj
D+lhisQmonlKDkeStKPqkZw5YJf7PbITd1wxYkHIk4lWIgKOiwVKX5pgXnm+I1xry5EOaqdu67He
8737nNBWW3Ykn9aK5jsTJA0ePqGRY1zyy3fz1rKk9nzB2B5tnmwVUrOK5CHAPN8/3ZESDb6Xfr+J
eEkkpJsZ2wQ5jVpITBtJPUG9Avi8KJyp5E20f+dMo4cYRF6Laheq3EwlHOq65f9m9yAC6dmgs770
htodszzy5sjfAlfX+ulNCi6iIrSu3iIeWdVKeGxtehz+qIaE3liS+D80HlrgQd46BkB7bBT42nQ4
zE73V+WaGmIyVt+WaBxQufYPGlNFE+B1ckeU6PcGfCkLP8FgATDkqZQAmTSKZ19YnayoyCiexskn
u2YQ9gLokzbrJx9pgaV75pABF96DTFU+20xsBg3hBgRpPVFWi67qE81FBSz6/uFifjMGL7aQlcHZ
bMRNewfVg2GYW4j5BZ1/bJtoiYBiBY4HTRG8vp0lvnN2uH23DsYXFNUxn+pL7MF5h4bXDYYPIG+c
HImWB2RN7sNimseEU57YHHZ11nRrcrhmY/rUMXceBQ4iXUU9T1Bn1n0jsy7r4twbZu0HVcw4BLzI
q7UUUrFbw6xOF9Hxppu2hao+a208O8OxGJB62a8s1qK9Dz5EJPrtoyH7axga6f85OXCK+7Ag15CF
UXoacEBzff7EEUD7B4w56A3lhzh+YJ86kCvoFol11+tYNd2+PV2OSiJtJROs26oBs6wEA8Ipj2ni
k5s1BL4968YUDVPIPlbBNRHGMIxNaBH+vkW0qXzYkKOZRDG1p3Guo3vu4ygW/MoOKLCFJIUYThgN
vOl7BaXdTGvefM9aywG4JMeGW1McVi2905LNXJpu6qCkVjzA9lxbluosK78DtHOt5WUOUn8MIpcg
4rniOZF4fdYSDfS5AXEFbnxTFYB4lMa8OxB1/i0Tzdm9s79RG7Z92XCKPVeMwtq6ENSicOGtvRfQ
LIpXo8FpUL3zr9d2Tm28WvZCpSiNeMyDH6SP0TfEGf5j09Se9Wjt8Vi6CmrRUlATVQuIK/7o6W4A
qs1eJi/W/WR2RzD2QRv+pVnuzm0GkUPib4mgoThud/Yjre+uV6J82MvR1+86uJJjdePcvmXwNow5
273WUMBm+MuQvmzuGYqfb2RIjxRTSn+fkBedevgXGHxXYEe8Cv8/0GDVvDH8Uvuj9oMadZOmOuf+
XLCarNztSsca3onBADsK+GJ6eSW7ora+UlfZ+YDjQG/i/4rxuIWVbhotABZyuleZdiIA6Ry+y4Fm
zZVKnSFuD/mZGizFObyaeZzRJp8kNYBweXinpsGRtlIGUhj2PbBjQVXTNnWdbQj7j45eEcktsqkN
yI8dc9DITgBSPAO3FMd294OFn6Bb9xHnYiaWtxv+JPaWyWV90hIlMfPeoMT8ebC+9NLmyAXrJl0z
y3lpxMFZT3TkQO7nG9kqwf90ivSk5FQgfldJk7gobYBJNFhMK9v7OtHZu7HzAVAzpaUF3RAZc/HX
3ujs4NXVAJeXy5bI72HrkIWReSIYKLDER74IIU6kWPa0xmw2c+Tf+rFabZbPKQremTtk318BlSXz
lz1pplwYXkXqPSRSpFd4xYSru6ivs4uFltN+GNc194EfzXvr2jLfyGt0GNaDe+NhRUEwvACbgyvM
uJZNUxigVSk4AXg9XYH3DSXcXnuQ8W1ERk6vLOsRnS0erpaff5HdmzjUZ059JSJl49yvZqjNvALE
A+YBmQvdgZZJu9K7aYOasJVRWuRW0iQ0YprKDP9C6U8tXdYyhM2B/IJ1vpfXhEqC4zx+8421zNPa
DaaV32Ucr2+VdOw9eWqFQZjgyTp3Colz0ZFQe9xZLyq3QVLtftOXaPLziMceR2odwsYpDQX+4xYS
mm70bSi7u6GD3o+B04j6REujYAAhaZVaxJ0TiCl8jzJI7g63ZUEnwYFIoQvf6nlpqSIyAwp/xfW5
7X52mtpTblXPeweJxyiOSqf8oeYi3e5AiscMfaQIpWfhqgzY8i3QlHPzumNl/YIz8n0TesCC7iYW
jA1Ba9w9jHaVt/7XjrHLbqFXiQmS593b52gwt6eZiorlXqVpVfCa4TaSfvFs01zjlA7CgDEVs+Iw
GW/WH6pJNcvZLlROGwi6XvScDhCQcKjz4AjOOUs2Jx5oUmOLVQaLPrGOgSdyWwYJ9I/rSwMT+eGJ
HJN5X9eDFHMv7C9EWzQ+MFJS73dGq5ni1OF/62qoVfl23gYffKETfro4RK3b1Uz/6ZiDkfi1bsY7
aIpdCS+mgqrIxooPQNiq89CwwJODUW9I/p7edeaq+g4aaeCJb6P4i07UpUJEMBwklhEcekaMTJVy
AnKADY6+Ntnd24s4SjCt6KnA7wLTBFOMaH+cnwHwq0gAXfSyTmTYT5XnrTK7+zFDr9xQVoRG+ARz
0HsXQONoyVxPlLmSzZFELToK9GydRlWifENeNBjztKIQOLmT/k6HkeKhurABtX66bj9Ct5WaWC6Y
k4JnOlX6ur9MFaCT3J48sVkRBc3mIuix8n57adEQFWX19M8fVQHpPu1yVeC9iokzbBTWUdvG8/D+
jsKmnTnK4YGTifowqahaxktViRS5bj8zJU5bExbh7p/i/4ioHKzOGsBV36KSDxsDVhfo6qRzmjPT
PS+wIDhWbiNv744Y8uRQ8+LuV/12FHnE4LxoxwXLlW7w+biDck2nd2vEzVEsCepMeDRaC8nuJk6y
lmL8tjtl01nuAiVYZnUEt1ybrNpmYKr5NK572Be4GWI1oCSNA7q0inJmutPAmO/IhXEy0NWWcB/+
HSEbySeTFBekmBUplMaJ8mpVsSi6n+7xYiKhlzptVGhNIaf+MDOjptLNZPPLPABSzFYFNLAMM0SA
xrcGjwDhne4hqtZUYcxZ2k5xTurKamdXzD9wITXi0pPbRNRGKLVrXBgBKrF0t/l6z9BjAFBBYaVL
VBnqcmmCVEfMiygP9BD4+99EEbt8sbe1pKS8aLegdlFTkZ5mBkI7tthnj9DYXXjsdhKCqjLV2htv
mJLCIUALTEudC1cFk8hwrl9G84j30hEMHq047ZBklfL08J5tmOJ+rnRQA05t+dOt2F7jXXREzgep
M8EZhPL8My3RLBMRNEMKxGwXRK/gqN3L/RijfUVNezY8t6Pkh1MKwBC4reDQpeDp8ScBHJX82Jz+
/qC1emBpiYUjt5JaQzq76RuzNfo6edSU9mxzNP/mLXv2rOcBVKok7Hrk4eHDWrBm9LrJlLqPnuIh
vo1D9Jqeqb1JsIzWkcVTjrqKgPBsqbqjCysfHAY+SjsMjTeCb5DjU1KJ5gu58ZLlxnf8dtx0RKrM
s4G9M21ZkcoCb4Phd5idXug41vr4sn4iP4VPOxQhwVhtRCoSCSqJ6WBtA45suAqmsWgzUK2lPP61
rnapuvoTVOg5HC7Aenyesvg2Fk19Q1R9VFtWG+DDDXdtS7Vb585zXJpmOO/6eK1esOxU9nyoISRK
HnQqxxQtYkSHsv8LVhXpR04kMvVXZepCSPWVzg0r4bshhIlxB4cZkfQ+uRSxdM1EogdfqmbznvW4
9esX+SpLRJvJJ8gENvj8Z+6obVWPTYrm6zIyoc8QQGICUYlB1WpLvqOrIJfC6Z35STIUq57Fe0dA
iAc/l7y5wlwuXse+sayX72pOBowt6PMRLaJBnNzVmbqLXHMgsT7mHK1Td9EojQlusZX7xHQmKWgG
+PvuTcGlSpCHRnqguf+HZUwZcQ/G+PACu+op3tYtcX2q33n1+jC/q6nfZKYfYP5is2W4sL3z4Lev
v5DrraVIwmlwr7bTrsVsnf6pPak3WRbXqYM4icAN+XyyO7gvcf/3LE0iBmGeNpsFmM8/zpoVKgeX
Q9yU7ACzlhtP2VPO2ARdInqxZpLSng7F1tnz9FyRlpGXf/ljvREIRJAmnXmWnUhtmFRmaty5+p6J
7olmvR7PRLwPnD91WO1XflW6smPFoLAl7rGkl8D9oaWMzkuqMydW9pjM6XXR/+2W0jKzYHN4QNbl
jAb9VKEIo2yLWPk28eECVxgft2qdqGS0NOR99a0lGzaPXnFkgQ/EZoXtDbDSjRoLnecAdB4Yx/0Z
l5eauwnMZh30pkhea1bEIxXyti0jHUWuHaLtMqqF6Mni6GOhrd9jCPLS8WSkLpOSt/b9KF+duHpb
rl3nD2Kc3gQgfIVJ0/iyrtLNL9QXH8jlDEGWvqbQuEPBYElUKbyUcJE071xo/brIj498rvB06uHs
thitFHB3xziyTvtRqFSls9/TqD1df6XFnhPJRl4JP5PqFku1u++Giej9U+jedmDbOMXxjySqpx0s
92lVKkagEYGl3TXHKhS0Y3/jbnPo3Xub0Vd97lfdDPhRpgP2YiIKzWNsgx4Tr6E5paDUWk9G0JN+
3ixCNtdCaqjcLTlwmbPwe+gS2kW9kwsPxONfXeEcRffYyx3Hhdu5ZuPQCMW+WRrY/qYiXDnT9lIa
JLGypNVlBa9zN4eO5+EskpknF9yzVNXNe3/aiYCvDSUYqNs6+Uj2R9OJWE+WbNaeqOO5nvJdWmJH
FwRHKTVl26+3MtTMvDby2aZXYmTy/zip6RKXgx5jY/SrH3/9VokhnhzOmAlbFQqYcqlJYa/UCWQn
P4kttnJnJE7A1qY+QA92U5yu0zrFc5uwmShd62MDysjv4Idn2uoGglZCYujac/XXSh4i7LDbrxrt
tnFc2Iynbxune65HX0Iahits8WZygJM5rYpze9RXtlkwFtD6K1nN24iv9wjGFw93NXbE022rxIhC
IvpwODsFFEtnrokPiYPWv/SbGFlwGC/7quOc8Ww3CmDGi4RMiWElW8JEeoqRwFpuDch1Bh/zQ/6b
UDYEYTyq56CSY9JgjpWW3eyGLSMG5KWqTeeCcLXgBzHHHs7d1EzhHp2jQ5VsmvIM/0sF4i9hmjlI
nArgu7cwKQ9vgpELTUDUAE8b1mlkWyo4NJbawOy2f7yCcB3lHlc4t6K8zqP9UU3Qzo6HA2wdQ4TM
PzGEyUFEAY2XHz+K/sV9u3dY9g36eTSBAf0dgv04cAnGG2pXG4SDfVNTtKjeYBgKOi4UKLw5sAhN
aOPwCGLzS3p7fVuiw1bYFUvThVk696FNDJKIteL/VAVcJA4H02NeAg6Z3f9xadzu2SLbIT+w1dMm
VFtukRKShV82v6/GWGGkzKNueY4n3lNhuz8z/7t2uG46PSgkeFmEWQK+RKbx9qfofxeTRIhzQEt5
RLtf0RgFCeVyTVZC0K28iHiw5kP9+rXeC2rZOleMPhm/uIHeoE5Qkr7J9BYoi/Z14F4qnqtQQTC8
KqOGUt/keMHeLNmzCbRF0ZlzyQgzEcTF/nTsvMKTDlp+8lUxSZOPBowk1VtyTmrRDEZwHn9ZVZ2K
bfuH7QtEcBUE8yQFhUbQp96fdQqtNAUpQKZZEPKCK3bIjDWbChNljaKAX/L/ushR/WJ5oL2Xqt4q
H0gwJlUgwJ0E4tL477RItbisTqtCz4DLk2AwV/6bk2MAmGxjqfPoNFWPQYcpBee1wIDjiXINXIp3
TPHFTt3l+S2kQK/xCecyI/BkzKddiVxL5B3mBPACi+wHNEtJPzYTiyeHq/8wFMPFodViaLAw2iGD
mMSbf9yto65K2Y6NzdLlArFL0yXU/8wRtZBw7/f7Qtg6gFEk8XDbEAPL/TMxAk61zWGKErwuEwHF
IB8cqp6WTr2RmXXA6ftsoYDU/cad+GEQmVcjt9U+Q2oI5ZtU+FrAdutFM3eq1P/FwdMoG+Yhbawb
OVLGqMcOR10e6tZbYP7TNoGrMAm4vOFQvWiBmhi1KTBtrKkW9FY2kWN6OHOXfN3u5maBOWJUlYOe
33kRPFOj7iVDiYq3+jQEmScICl8L2SVdl6hMCI4Ku+w73BJe7pD7JmsnyUgMLsU7wAqwcfdalotw
9+YVnC4KP38B97vsszLMIUzsCUccLWe/EuOcUydgW2qsP7floH3jIfbR0tJSeu17kJHWQH+SmuRe
0t66moi3i4gUtNwNZr4HfQm/O7tVFqNjgoUl4wwateHQ5Kr1ZVYaUycKk7Zfh7kszES+ACOtCrFl
We85oYx6duWidHV3tuzR4n/08LUKYJeC78RAz8O+U3LciHTTB3EtPewTKLw+6Z7WKftd+FBHS55T
tT+CjE+omMdlWGD778GSVeyz6Ws6ULsHc5Nllhga5/Aros17Ii+Vh8B8Hsd98xx46QbG3sWPxyXr
b9ZjH2QnsgzjF8aawVC1Td4y3uxLEsPL9BLhTSqJxc4adJokMfDr89xguxChywANVGChdcm7Kbsr
t7rbp+xVshFeoyU8qwiW77chw72AeZtu2Aixx+basUdJb+TS4DJgjqO/zIIz8eS1txP105Ol13Ns
w9S0i/bo+yzp2cLyx0NblZL1fsVeROIhLq3HfJLDWiNCSHVWpc/Ar4sE0f10XTQJ4CSNNWy7uOOk
fGV8FeAR2In/aaFVHyafoe32Iv0L/ONxiQe2Zu4El+TDzWFOGvdv5DRODHcUq1QBCvGdJtRxfzv8
KlJxef0gOfN/tA44SMFIYCYFcNNV1OoMwJ08bIsztOCuBX2+B3hYG0lQn1N4juwcc12dSYf+YK0P
pJZmYXAP0uHvYLRkWu2XxPHoaf0RYV6GCSEvaIXusfd/KRX/9gAXqzsc6gl/O4FvJktib+Iloity
EPUVTsrlUM5LxVwkiOY+1mtGGM8B+9Sc29wRSDcuw4pSF8FE/iju/pcC71WSp+359eLxwHBF+1HU
SSJBSgXYaRQFw2lXhXr8pmbVc1K692ZKFed4D+h8n83Ggeh8z2yiPtrEw/oXjZtRI0YnP9zyp3Aj
OI4MQFlKCtLyXgywoRS5PGBHr+EKCN8HgUfjSL6RcKbtNVLPQ728G2DxiRTRZxOz8oSIZ2DR6u5V
Z+fKCqbBywXd740AyHxN5tJdghQtAOdJUXiRhIdZnnchwXQ+RRYKPB3e5mB2kerynsfLK7CeQz5M
zm9s5FhIrLObNlfIFYs8cIdlwmAkXpFkgw9WNTF0+YmgLEW3HDvnFr2gPGQSBTegP8xcl1w6LFm/
uWrf9cTRMzT/VAe6PpIE6JdVzqYGv2QTNqrR5Jn7BF10wOF2xrywHqvgirOa0EdDo7pd5lVfE3jn
m8x7ptGmwsmlfwIbsyT8yf0ibzgNRVRN5CKi2pubvtOaR1SzeGQn66BRL3MF2M/ZgwJl3IuJqfUH
tw0elRTm3cz9rj88gZFBiP9Lh/fwCF1NR4NbtjJK9u8km+GYW/LVMVrjptW3D6ouo5KeJH6j7zsK
eT3JILf624UPWhBEmTT61MIiY7FmVoVrxRMp3KdUOzIDwHwDXc1x1/v/yTW5mp6s1mREVkhsvXmC
8EsKkgJh6lhP1Z1yKNUD9Ug2uiJ1zK4pZ/3OR54sLbiR9qApMUWtrlqtjqVMXXClC4yW0GPjqsze
YO4Fkevd6Iv7XHF88enKbZ7EmR6ZbNyz6dhGj3htueZl3bsjIz8bHA6m448d5mX3c0/OxPy45uvI
WlVziQLu54/yfR/K8Yw54Dr6A2Sc2VNtR0ndObkbQoZnSbb9H9EU8xYn3FIT8rCFjIWBHESk1tDS
R38kXOnPXGC9rGycbZSUJmDYJLIwqWxTe/sxmzIDkRfvZY2DtW4RYzYLoXm1TpXh2sQxUQjwb/eb
iBoTXZuKPdtaRDB7B84VIMe8PPvTr/5kfeFNWvYSytuqwuB1QUJgm2+8XnrjCzwqSCfcv6MAHDX1
sgageceTuRzirxZ5ALcNDB4FW30nzhhmkNVqYnrE/0SP/nKvMTRgAgBi6qVw8VKeYeJlz+SCGpBO
e+yjB26vk5mW6DsSmYa8gGR07xjwPW2MxluLTx1O2J39sAuqiGvsDY6a1PPXL0EobH7mDhbj20ox
S272Iust7H5BvlFuvQSljgQTL+X3bZgqPX/bdtfYDNTEIc5LfPgMzvLAeVbihBq1oNsA1G9CJFty
f3UfsXTmWONC0Uus8FJsEOxJqYi5hu/2xOOUPLkQxgLQEoPnwa4u1f+lSTa34dThCUCmW7NzAyvz
+kCiRnjemnbAOvt5VdLQ2YiVorFQMEncfVEGSRie10zOz2DC9YisPUGDzxEJdWdDyegb70R4O/+P
4jiQ7VyllmxDQ4fxNCthr/GBX9P2vp+IHd6tOM8qTlh6/9IZG9LHF0cdHiyY64sROv8tf/hV+f8n
4yRvCUICwljkE5voOfwyyOA+ki0bCUNms1Vp1BXXeNwFCnE5m08PJjaUF1fM0j/Q0oKueacoi1az
FqmW1DhgssjUaA817v4ffZXT0YopI45SXV18h9vHJjJgvr3B9GpYX3/EVVoEgW953oUtYWFeWG5w
IGpi4pd912A3/+1yoNRmeD59HDN3WFhsmg2nVwzG9P6ZWe0ZNYeFDQOeN1E5aStUSoSPmh8hueic
icmDDP+bTCsSniMxpODPZPbFmuPV/GTgK8uWYWLezvY/RYiqvZiGfiINqt3qVJYTiZzDSVaJr0p/
FsdnnUIB24DrXiSDBLse07P2UzJPj0UkzZgFk/29zB1ZjAVVjWeAlErSBHiAC+JifOXQnT604QwK
z9X/7TfIPslF0bUhyE3Jb8ZFNTWNzHIun0CcMKVB31QOazAFr0wNG77zFs9pNjBucpzV8hYFguR0
UXHyQF9+ukJPoh3rQRHmog8ckfAJ17I894I0TML73tPy0kBtCZ0IL2YYqoUWLLY6iMFIXlUj0uqr
9k5ZRRW77nC3vaog+rpyVcE5VgykudOeaRbSShwrtSu6WfwfE7Ae0ZEK3vN3ggOXyW43Igc8m8mP
E4wNyNeFhEOaojnUQnN+XJYwJ6PcHOpgCi9z4zKcSiceV5rmgnR6nnIYhOlFmcjyfG/3bt0o5jgH
hvfmyvhXoM6GNEfUHr81AiJih6nlAllAsI7Qxv9sCkQnEAhwtQNu1YRiO+vkNtUJQO0TYz8Z94X+
Nn1sybRjPpYhtLi3Zl219YKKD2ddTYveKi7b8wX/tDe/ztwBstaes+232auHouE9vWmpvXzi9/Hx
BhlSf7RA2jA9f4pVd9cMtZWYlaWYbVtINNLujqYbdFSjzo4MQwdREIZj4gjUjIiMUhGqezPsSpkh
mNyqGHuSYRheaYqn0+EwUWlBtIkz1inB8IvXDUHXMhP/UgyEBGjVLUFEyyVWUioDe+NAqfH36Keq
etLNzf7uTwK1ys6HgGpMKxnStS1O6fqVFTH1dil8I1R+93Lb/+H85S/DKl8Js9fkQHK4zo+wq2G6
OpKb5dABt0ZKGW+yYzl9rCmI8pOdmqloemajvyQwKWJngN+tohUelNivwB7NtyH6UUuu/L1Hnn4W
bUW3o+bjiGhBDAa+0ueiom6XgFLkpGAPtfQdxFVHVBuGDioU884kp7k2ivuKbUhSyb1yaJr6DaKX
l8eMmQGC8kIT8aBb+m5AkgFdU4aakGLTMkbrzt7XwtkijzPnZvz+4nfBT9GhuSKyDXz5xWSynlAR
eAumjGlivOwN6i5L8N0GW1zcLtTn1+VSt+qwJNp7yEfgBQxPW1li8i551Cw07SqQVMnm7HUNukUQ
7p0hQi8PJz5hVU+h8u+JgzM9dB8YhLxU9L2RvlBpD58We8qbquZ26ykfTmuMB3vKFeCwty3lzvaE
CxIMt/X5iSx/BP65YxHBTyWM9zJkVgrfoKY6NQhVb0BwTHpxIvUeChRdB+ukupn8cMCQ0PlcoFk0
lQOQxxfoJbcRLiiK1DfS3t1uIou6USzNnwsUNGZCQmr3++23WoMs971KFDlSq7ko2/1Fl7UB6bDH
6jdvElM8djmUEOozj9jlFppyVPMvfJ9RihIT5Ug1UobkCMlrvxWzoi53KH5VHTmOxqSr5gVLLpzQ
eLnBlw0L1s1QVlh5qjmSyhJ+Te5fBprFU7/3OJ9e3oAGp6kAK4oI+KSC6ujP3HYYPl6dOcevDM5z
Nkc82iKcBrK0XfscuPR89x9pkVbKiwn+mIqaAaPPY23DeKHxVs77sBJUndbdJgewN3MBM2yZmo3Q
5eWDrRdD3OxI6wiL0LOsLsQaMbHNEGOJWkQk+Q4yG3nKOSyhZI9sFW4+lBxi5wwDqUGXgYpOpUij
XG3Zjgfk3ol/Bt2e4NRF3e5sQHQ2Ki0q5+xHidfczhee9EUXL5nrxU7uAtp60rDPLfY8ElSHnBEJ
I/4qNTaN7f2H0x3swBM/Dlzhd8iv0ughupdiLzhqpxcFUHFcf47ZHqeni4pbyly+0w53vkjTJ3h8
t2UI8aIQdb0sMLnUrjBAH8QcOzrxGWVodvU8MNYAS4C05qM2leSDy1R0apwTarCvs2+IDdrpyS/9
tEsWsk64MUo4/VhsU8m8cBWS7sKG8TS2amKAxe9EKdrFNkAlhY4H/bmrS53hNbZddcxCi5qBFvGC
udCXTXKg8eL8rHtUXiGDdKG7DlViW4y5c8ymecM6z6X8Y9eY2er512ml/2mrpaNaxhDipgEqowLd
mh7k1gGSWHJd2GeVO9Hi9af1OPE6CLGscqSI6tMxI8XI+02sxuTkMyklRecFoOt7XmVvNuqYnoPI
sRL1cSIln26CAkvlZpdNDEekhptuYWAVtae+GX7KFeYpIjBqUi6QKVNE08qfhVvgTUcEvCg5jI7u
2rko7h0pb9ZwbZgtNC/J0jy1C1QoqPI8tfHySaIk6sqqWaPNjyqnMRNMQ8BkmgrXueQRrwYYPcQP
P+fyDd4wwEKwPw2MBSnj/8/QXk3me3rFn04omEhx8GGPMheaCXLrrH+ZHMWb8ARL4C7oOirraBH1
pjZmbTwd5XyvsD/dpzognezRSx18NTPqMTnvC1xqsS5bs5W0onj4u6VH8u6g/5bAdAtDolYY212w
TTZG9wxJMbvOKQ0n1MYtwlhGdl9x4O2J1bU3R9LIL8i/10ugRBwBIa2DEx8+GBTFY1Y5C5kcw20q
cATYYAY8Lt4vCwYvDnBpjCu5i6eR0euRN8X+plK7Wx9u6Gch/kNmcvSueKtfTynWKPJxixA1VilZ
75uG7w8r2JMsPr0UFEz7V2QS0zCvF0zIK5KH8LCdw/YX2hSkGYZvF3ZSiedQU9lpyMqvPfO0ZJkv
P3Vs7lZjVOe3fqrsEZ+wH9N7o5n49LzYYwr6VWLX9oyjagbxEncPEml43p57SQ7CF18eixq/NmfA
aVAi0U6WKT1W85QrpskPwgDFW8FWtL8x6+rqtXDa+VPCT1ooYkHD6a76E9D3p3P4AeieHHmbHTvX
YwTgn2xQEbp7U0Y/UIKOAUN0Med/UdYySIvIsCQwEOw/aeYU+Q4pJC9QdsVDxcAFwVj7WxeDc8GX
jOc4OFvs0/ehFlLi/WGOtcCUUF23nfi3WRpfLyYrTv9lXb+BZDsMA5Veq+tu9nrHmurcDFZDUWXO
9K6be+kfeAiXxzjNQJr9VQlOiuiDRyifFC6ojEvTSRQgcrshmVg+PhgN0U2jQTYpZmc97TLSA3se
dgcLrpXdoyfgZ4vCOSFSi+stXXWqNVHRoUQDitueqYkrSkAo3LcZHmEfKJ7Vdc7XDpBQLxovz1ml
PewnWHVvHAemxrALnzYOwaEt1gjK4qKmRXEcAliV9XNMi1A+TquMHIfPYfM+iOJBZkz4DYBmq0pn
M8uwK3DN/GUhb3ONRdwCUq6dgt3KCGDlzVbDL73wdpPEoMwcFx9UzGyKIaWvnALT1XDaB7rcgOba
bz+ATwIj6Etu0jxtOBjTNNamGPC4YYRJgh29hNJXM4wPcq2uBscwr16JZ191JHkc+VVYkQcMKAj/
Qh17Z9TiwXicbmHmO435IZjf0THCAHuXmDWQDH3Qwf6tKuOBttfgWCIAS9A988wFFeCwj7ZejedB
YkvBKx/nqKbg/0DOIzDvSAGaX2j1iKk3FYlvTmocCjUBGk6cjhglSnx19lfBLoiXBarg7ZvyDOzF
YIVzo1xNnyqlNPtWi3oai82/v+zuqa0OaZAqgR4KLlpmE5hF3vUjr9SiubQ21oYYi5bohddMfTa5
So8IcfKhBmdiUr1/9miEtV1wRp9N6AOTCzyF3DzdfBqrBifVnQMu7yNsMDQ4w0QZh/nh51VUwbOV
t8FojBy7KhsvnX6ot69o6Mcb9AkXjSzhkFQ4mZvxYdXkyyCmJRVEsCHQE9YO70Ge1WrRF4B3Kruh
zcJIpaNAqbsLgKAz35rLpZv7dIV7tRk6UhsaNKjRKLTmv0QmhrOnwQadOORrvChhxfIMVpXLcW6m
TgqbNNdLOK59+AJC2vf/gzwqPIazBMo325Esesz/PCOH941U1QEDjuCO29TbRWlRVj0x3dxxFke0
pWGRa6ApQdKZ5IySfrHU2qTmnFHGgVF1mmqEbmpgw4OgMtgc2gyAHSGeqrUQqxlQQgExhJ44gZbv
x8L23wLezy6H+MdoR1qXLVIoGa54Y7YrSgrOV8SH1eIcxs+y1mjwBX9jXg95AFK2Yz00IpzT3b4M
vgLSra7P4ZZLCuI5ESwAHCuQ8J+KqokKX62ubdUiTtJf6E/8KUYuRfro43IfkjCKLuIE40brvv5x
EgV8+nGljwDF12IgP14CucnwjoEh9OKWSMRqSsbdWF6ZKf5iMqHcsSj2A1VDcMiT/O1WElHQEpoF
ZHJp6hXZoT1PaSpI2OG6qGdr5iW7WZz8sRf7V7qZw/lXsuWB4eCWH2R5dJYJ3klk/A99qwmCKjwU
Ca8J3eDC99hkln42+FU2LuwqfS/eFKFsZzE8tdh+dNoBEkDAv2TtaniB4yItsm6GOvcp1x/2jXzl
FrKoa14SKdYKXM2QFY6DvMpjnkmKlHmIJgyI/O7GGqi287yU/qDox0RNXAYdrfDX5cPWB/N+ymqH
i3uBVl18kVc394xbcSMQ4tkL1SjlTK9WgdhlzbAilPksH3wsnBuJw+uir+aGRuSliFktzwSx3I7Q
f2EjvS7kTZ+pn2Alu0xWrEwP7spmBZ1UYT0F/IemSKn5v2hFV5W/GXVtdCVZqlHDf4X9tQsCyFMH
zcz9k9NrsjDTtymIVfZ1/w5dhLl190dC1J2633apJUuU0swAwNnqBwOjRz+RTNbLlN8AnfnwNiKg
UDkCKEtIHYF+UREmFtivt0j0q3Ev708Z74UH6mEtZnURMpurX7TL7GqWxeK8PhoKVlyLM/lx6mon
5JXCz8MkrVQB/z6XEQ/ue5kw+SmCCiFjY5td4tUFMB744+jdl8cMSN4N6k3zhB0ll/+otSLc9m1P
/WCvZUQ1Rn/HzHBct0K+Ke9rOF41iq8Hu3JmljooGanVK6NJCCFq9Jjn6ZsANR+x9PpXGZuHVRVM
ojS0HvlURFBUYfQPwcptOGKnmPtjlROzCfpV2vCOK2T+2cLI+TsZT5a0KibcjmUa0DsldrUkjK71
vw28WZWxr8Sq1xgmNdJioyQwUL+XFCKjYkMxR2wZ0A0481QS486Fv7akenU9MCXMDca9jNyCcgKl
yU/mmcf+JDqMJ4wi+X82imlQF5d0got5Cws9bXBJjIMLwLhitFQtwiq7B9ysHzDnFvDsv5IRwper
p9OkZyk4UykfLhyUKaO9dABjP4fKNQ5yV/wJvtGr/rl+XYup5cEFwC3JZ6W17PDhjqHeNU6J0QGU
YBVD3c3Z8VQS+TI0N2lrDvCcU5/ND7C3x+lhyj8SK3m/r8ABDBEKFD9zM/NGJIBsxHFB4m9+USj2
00/VIC5R+UDf4Byb6OYBDHSK5C0rahFs7zIBXdJH/+YXKndd0wa0VdrQOXv+DFnEJli2tzz761hG
pI4VyMIAJlBgDd3wKdp3/tdU3RBNtIXPhZJNQsWkAGFsfWMxDt9UIcGzaQlGOyLQxtEHUciGi93I
mzcOsdAupmZ5H9SiDT99nlNC5jub/+2IR8PUbIPmW1PZtDBfw9CkjjymAYlvWE+Y62J3MwZvYSWc
KzVXcaoz7Y534SD8oMo1O35QQV5dbls9hxa7+WD2wi0EIiB0R4hemA61Ajr/XTwq5BHLk74MXJ+V
PPFi1+BmsokxV1WTwBWsqcErZrc4IIDj3rOeosYWWHEAwqU4TaqTsCifbecFQaeW4cXCpoWElBr2
OVdpGb9Es6U+7y9KbJIkX1elO+muSVQhYRb3J+hfeKm2KchX0+uFByrNp4orfvx6mwCEnKx0qg8n
H8w3jHOHtr4HMVg5xl+LHrkhmpQ+2+ZUxwVoSmT2oZkBoQr/b8eR/RBINF3/jrGtpOaalw37IyMt
/GvujkIFqxmFJl76AxCk0+6KtXwUJDbnEMH6+fv7wFRUupF3c/BGkn0gT7O5tqX7HIcXqi64QMJZ
zsNj1RADXUBFcFnVWhxQ7asMSOmkXn4RthjMrnlIqTPCOB36iIkRhFCf2Nnwn3qglKNe2PVhPnfl
v1zDfa0rtywk9E0+QZr7RuTaqbiHzcKRp7l4+Hj0gyVwq4/3i5bNNOGj6MhXcPZEZVfIr7b/8OJc
EwsQwq+Xv1VxOO5OyS+xF/DB9J7yi/3vM1TeagpjKM20QjwVETRQyn1IZ5rwc8VBlUsaBbarcLFt
LMEVubv5zPE7vANwH1h0RY8HwfTfJdYhP+hxZ12+zC1mbxoRDArSYHPTodf1mAa40GCM9H4KvIx8
BV4XMfDE6s0EAxRVSgD060LUoxwmHdlssWEKVjZxRgpfuZ8r4R3j7cSuiQLlPiQMXIHXyVZ6krQ0
OkxQgW+FGQ1bV8PABU6gGGdW635ZEKmbxFJeX+wOB+w1d4gy0jZb6WBKVoZ6PFseXrlORCXglJAx
w5RfvDxYm/qauh308uJjuFpFXqzyY421f6U3U18zcCgK/OtXIPtj1+Q+F2HW9DPNlY6Eygu4SmD7
hQ4334oao5zr9x8V9O5nCSZ6/BdpGjSkzyQwti+IRoZHuP5LrNebJSpmM1PU9cZVf/E3MDjc4lxa
zO4PtlnK9PnCnafYCirJ1Mn3JwrHHe1Now34h9hqBnMJxSv2kwPHTwcJ5ZWgeBT3AUWl+ayFUfit
FNG2UenzVFotWX2chYYtyNljoUNivti+oySxwynKrQe17cn7+Z9UFRXV/Bn5aWYQnz84LrxdmVhd
EtAcBF9xuoeg1cnBLkBcrJkxFeZx1tXmmaJayb7y6bXdWMQ2ueFJmnIcXHdZGDaV0edwACw6a16t
ZUq1scbdZusuuiuW8VhKJDl5FDuyvi6dyo2ZdF/8NUbCwseUgsQ0+TGUsKRifvCrtHI4Fx3OMdvT
oY0KkW5XTDD/9lg3zzOH7ZcrQAYLCxe37SzocJQfL5x4rZZZh/X0q9+uGNLop+C367LA3cQGEvTH
8TCjGSEu0Ds67SVi4f/9znP/s9hShF9dJDiBFoqbDvWJ8Y785bndYeDRWf2WUopG0shstU71/mfm
jJBvkmyEC1XAux3sYeB3zPB8e6t29/YKW7CYf8jdz7LjCJN9hdT7HGlsuHVGXwRlyGwA578J2df8
gETo+gYvRTD5bZKLCAOP7963L3UFx4UGgWhCJWluSWnl2ugK4sq/uJyIK3VqQbE09YHLJ3+D26Uu
GuC6/+OQStYS0t98RJXwet1fmDX2mEsm6UTqnU6HcyfaWU9cUH4SOsUVT3GN7f1S5gUyv3ruobPm
cEDJ4kxZYOrNWQ3STd8Q3aGGjY2++FGSjSD5jHrAKryJcYG/48rDENP1XPRjX7DBOBa0H2u+b55T
L8FVuTsupUwuzH8phDksKgfUAL4co2U1ziP5sCO1xt8tBuPLx3LqX1w6XXUH4Qnu574I5uK6SJBw
Z9a+udoTMWPhN2upkD/mDXz+wsjGqyvmSmu43MfZvQy7O8q+Pi51w+TpYjzeMkIcgNkq6Yaux9p3
tzQj1eZcVr9TgQBRhSnUGcQbqX5wbLLp36NoVk4/O4W1Wvp92mTFX7PGHY/i6EdFFiXYf4YCI97/
jL/R5MUDs2vZHVlH24SpQhI3upMujzuVuwgyFkfwY46kDYPIItlzsDcHb80O/tUtktmcvvidtxey
HqWOZeeggT/CaTzBrXfBJt5gHEuCELxjthLTbtymPmv0vAXjlYJhCYrcSMpBBx8RlXX4BAMfDpON
MpcUNYG+c1r0Bo7H/iluRoFfAkgFq8G9X0BYhOUL9QP2N6Zqk1dbsO3GbSLQ6PJ2Ij+v7eOTG+4m
83/vMReX5OsbhmPSYwA1f+cnFuyjgVbOyOGFslc5APel82kWuXtOhhW/somBNR0nc2lSjn51DTl2
vqG+86k1qA864dUNzZgTyZUl1qnSwFU6u+eslM+8/9PayxZdTpEMOAul2/fea/i6sk1kg7myWs9Q
wlN6BvAnYe815Igf7WVvXyCc7IWod6N+oH79MFBVZ/QEou/hrbbiTCnolG/V2roV4Es+qOPzD5Ml
aIvABmjBM7GvfM93QErRJyjobNR5xV0V0yw7TK+T4GxZqTiM+VyWOUKDoxg6Dd+secZ9JR0SRMzL
tXDFFmN1OVnTuYYEkkQ5rpUVTnCFXiqaT7c4vHP05AqyA4yQv7kn7GNbR7VjwEfWO5y0f4kPzkvw
CxCmT+YegWRGGOVbd2QI0vW4xMqu1E+iKC184XPN+YvywRkdyWezK/bvfhxYE1AtkyWBlXnHPsS8
ViImxsjELRdzuPmPaxofELrdZABWpL8h294Jd9j71MZyjZJiWjOb1PCzIznS73aAYvwwdea8JYG2
XA/G3gKbCtwgfejVqE0EZDHWToLO56Gj8R9g3OWWzaXla64zQJosRKAa5Disf26LU/uAs1X225In
MHm0pXsgwFXCxmRbpe73gEihPox1xbk0UPVakadBs1yYBrT6F2Ka/dgWTttyEVKojGruJ0uu7S/C
D8HHxSN+m+sJhmi94LtSHawOonNwv7maRNZrvdp4vxr+v295b5RSFIpD+ZfZBPePs4wxqae9p0qr
mN2y2mplXOIF4b99BvZoBu4TK+CJPk4HBj8ATNn34bNOQ8FOfEoxfWpGshJnyN9tuGs/xo1hIks8
ecmB9hQgA+heBUGvRBUpXuKbiHaWV0uLeC445eT7Q1B0WWh2mMkdJJ8Uv0i54Ltrq9NUtF7yehI+
XYm6MupzF9pcMdcepqxjn7bujyIZz9GaMyTEX+uaRediBxq1jwvPDrFNjwpbioqjALKjUU5nA/fU
kfzz189RNH0uhPJFU/RA/JSQaIk79ohvVixa2E8pLaVBg6l9wk0S2lmOFvC7eMiKY9ofDeJ5oQlo
IpBc3p8o1EuH2afdr6LYAKbNMphaGB37qHb/IEeX/+QzkX+dw4vojflV26EsCdSwCb9baYcdTb0e
OX9iZ5P8KMaAwhEbrX29T3KXovixXTtRq++R5wh5vdctXK7mno7FQy1XffcwsqymZk9+pQuWHYzs
kZAhbGZBGvXH+f5OeMCam88mO+04H6qZK5SeO4MJNXVcGSphhQk6PKOz+5k3LPHXkM18EC2gRxGj
rthrCmK08UEHI1zyj7MICvO+jhlgy/oF9vqjWWDXgAfHE7o8PbfHyRvMfwPxVVu1fpD8zo6dZrQv
hfScAn1Ow0io14FP5pUzTh8qEffhF/glUKqo416Ggu6RlkFMYVmIUPzBgH/KT/9ReYwlTnCjL49P
t51kJJQ0xfmleFrU0NmtHbSdRyNzjlr/RjHI86+JzymA1AFOqKlwU3t5xJc1zgj/zjIS48S/Ryr3
23yTq+pRRWByUH6OFXxFlv2w6dCWRurYaiuaODKsXe5Utpz7KLcXUrr4b65Uj03uK/hzDYAIBhtA
qzoXFSp6IXFjbRqYWaXegDZECSgzbaYspzVIBIE8xY5u3Ex1M5Q5jev/5sUjcVSKTuotWmXNPQyP
58LPhI3zcSSVTpYwMG7mNxrQWXc40y/b47y8MCa2Rn3iss6dlSlO/UNljWFQPQq55UuBkUBh5q9e
JgK3HXp+ADcQ0S+0poK7ssMCXcUNt4vQZj72pApEUVQAPMu720QsAJbJqTeBz9hnDP/08cilyMt3
Z/ZG2/lYrQs/DPiUIXXSe7T39cDyHraMH9kW09A6/hJ+wCtN48Op7YggvaEhKHoEeHvLTUg5BfT0
U8c+IQS1qqbc7gGMiDV3K9jVd4utbGYuJGD831ezp1vxByqttxcmKomwy604z47j8zyKk3ojHyOg
IIIiYzMpnHuiAbDombEbi6nzNfJMCKkZCtUTeSvU6Z2+PucR4+fTFyMqeJ7eVBuTS9Gkvjyplpcx
NZRC8TBay6Q7/lY5oTX4Z7CiBLvdZOeiIYlVRJCtDAreIwbVDTUW6gveYdxl7s+creZc3+aYGm4p
tofDVi/377U9FdiG8rxOmlHrhp1gWBJ7gZ/jn8m/OFdT2Ff807aiSQEsAOMxFL1WMG3m65D2lSIR
6OorNwbCmpBMrENar928WoD0bNKKifeOcMMdxnq9Mypdf8Jnu5YN99oprHkYOGcK6Z6e+LyY4owY
wr2bb/ubwrVUPXGUt4cK7rqzsWvVrMUhLR6S0Jj7P0Frg+9jrjcBzkvD1wjEFcmj1D5+kQrYar7G
CgdwVP0UdKgYugIh4kour/sZ+nXUcCuQIonVxV0URYGP570X325pPCinZf0lNesHFwiTUl5PQRFp
xz0Bt7/MoIPklWbaKGmtn2PLnc2XOhlZ3DCK+w6uJrJfTDogc/imKJNcXvq3EgYbo2mdQVal4H34
RRlxfw1jMUGWmWTqy916pfMwH/OaS6ctOjHt1ecorZgyjdHQfnKd8NrxMBB9mY09MWAToj1tnp0/
vNWpZhTnvP21J6nmqA0Ki0t8vxR3EpZBDWETMRe1FiXweYhdpN+TmaSu5Y2AspcxBCXWtbsKfmfB
0aHJySUMQYIDy99mjYWoSrhQMb8ZWjLuLCCrSfUxM6JvYWEeh8Nsa8zu12x4HSaTtUZA1HCmM2iF
5wKYS+W3G+5i1atjdqDHqqdN/2O90AQ1rs7rd1dtPVI2Atc9KhsIpWiS/m59KgdyD/FmDkC601Dy
rr6fhZEwZ/XsFC+o9zv9XiAT2nTfI8fwD2wvQHGV/OklBvXFsacIcftLMAJPIFkntzK8WCpJ/4ia
vdo0pV3VzgAkNKMsnWdhFUimHzap5XngA58BFJgCdv/luNqd7hS/LTG6+1SO45NqO2SCdWIvmD9/
O3yG7Y2lEi5Z+w4JA+gIl3NpbOetoDE4CYFFLk0C/fq7B1waCthvuBuLEkZqWTpM/y3IfyAQrCll
iZDsEoyNJxzm1jJ8g+TQjPZzwKWNAvwAc5lsiXlaMEWqt7J/kORklwU7cO339kuoKCM0Epr0bGA2
YaSaN7Cd6IPEJTHHnLmvpQxuqvs58aJK3c+JvSFihr6y8mB6HV+Y3pwi5LqlGcvQDU9iYkWUr3FH
zk0Uh/BSLnP/4E03AaL2Dy5FPnTM147cI5KWXNPouFy5AQug+0ZgfuubfRDvdHt58GlKcVYvTQR4
eEdvJa2aGOa4udnsy6GM53jDiA0AN5EpE7cQmKe259cg3LtKpgtn9D0kCX/wymX3edjO/Y7Pi58d
Mk99rK+CNejmdBf9vCZRwomV3fVwpWUN/tfjJNnKTq6zRumIqo0nJzhyZ2KPYxoKe1bQg2euE8XE
ilxCDswfkaMn7NMPJ70hp6ASUsXI31WGy2qPtb0HFz3SuLQx2OJvrHMH21/AKMHRCHRb9I6/9nPw
ny3rUBWaJ42SnZgN5huGjwCNMsUqf3+P/jM7iBtnVguxLM+0EgrNOxzlwBUt4mCsxex84TBEw99L
j6w0pV6OPPCnAnJph7MNxcx6YG9NMJMIj31szRS/qCGN/QRDMaZ6gCsH2A0nbibDfTfsXZgBTGxe
QWUfObVCS3QODFFbJKX08CGm2UOAJGxub0OwKeyOytbABofp9YkihPpVhkaZPVc0Cq7un41TB1O6
nMNVdHheEzgq8B5D5kf+cPDmrRTFmG77epWi3af2XTksPd6RZHUobawa63lUDtOWEFG/T7WA7XNf
eN/zw9LPNaqmNZuQ0MbvF7JxADy65LDIYWf1k/noHtlK7rXkya5ClXONLnIp2HPwIkhKLPzsCJDU
4wObouYoIYoFm4f9KCOf/YWsRs2Zowlw2mdFGHYqcMEXAI9aBspKJb/UN3m6GcE5nPU7m4mG17C1
G/rkfC06BxisK3W9sY9JExIrtpGDQ6T2pbJ1ZM8zLBjKzr9Y0yo3JJmuOTWMs0cwKinTIZsbOmq/
KcxCt2pCHQdYnPKhM4Oz/ZuVSbWDYKDeBEoNT2kVAD1ZByHcDC29vEba+P9pu7tI/gMsFwXVBa5K
wuSF7kpP4oN+8fWqfMEwP9ARqC+5/0oW7683hiLHP01yIylBcrFDoRBac7vKS3K9OsJkKuLwwZ+c
Ge1VVF+Cs1D3Ur2VFldJsTS9W00K7vhTcsuYjk5POkfRUJDbJvom1z99EVzQu/EV30lipybR5tz3
dd1YzfdGYHouopTz9d6BSssLXrIuuFpDyeZOT9bSQuSZOZlsN0hYdckOjm5K9eC58+u9N8Zq77vq
CIu5BkH5FBzjoI0vOKggbDcq6OW2ZXUAtsojmt+gSeN8CeiTYBbPHYaTziCmItVOQWt/FhKqPOK3
d3g/1zexTNvHX/rn6ERkiNWUOlpcLjQd1I7WHdwqZ4Sm8TunRAjgyIEow6X54H8LygSJBViGdj5Z
AoRcxr/3KfXdfcqcoJB4hz80+AX7uk24cTDujBgihfk4lxRMCshgzISg5p4APGqix/lADQyHD7tU
1nUYNtf44lc6CVC6/fv7ESYdlNpRKa7x1znJJgeAjfNzT/55drcalPTLR+dN+JholvL9cLJ215/Z
MFx9yoipxa3bfvMCa9oayJa1eYsu8nOjb47nUFzob11RJaH6Ufu1JIPWAEwm86ajtA4yYwW/8Fjk
DDgxJO3L8DQjHmIj4GN6HPXZXMqShLMmMUUk6+l4W7sCGbdYekeqHJ+dDBdwOkT+nqgKTEtR0Y/0
n57eKxpaEV7K3DkbAKiVTNBHe1qb7Mr6E6YS5WcHV8XEa4LaPXjFCzj7R3aLrO8oSSjuQOqdDu6H
GKuKYLChHB2blxvj2Nib+b6FOkEhRyvepvc/EX1vtTXxxIWBBDp+rtPvoBdxGXb8sAUvo7JmvWhV
ojzirye7UihiHpVGEdwejLNsuoNW9IVsfr1y+9CvWBVBgBM2QiF3LjJTXgxfGvDT3CaqT8+9z8+y
VeIO5zLTIdzhyQf/51pReOKQhGAvP2LfFJrauAp0NLLFeYQidd/ihLOens/UTt8LzZJ+o+n157tQ
DtFJHZ97iwv0JhZNVqu6hfIn/dJ8akoSTd8UKGGYlsPCHjQnOBJPOmB87l3g9M+A8TlnQ/Wf7uek
eW25PVgc70O3HhyvrUMwuOFnLAThYoTn1KAVwoUWjcO71nsDHmspFiYrQ/WDxSu0znxRRmjhIpJC
25LjRYhen+fP+IkfQbBhCIEw76vi/Lf4plrQOQWWNeEMkouNTOP183qXABTbyIFozabPmFaoB/fU
x+C+RrPSKASkXg99g86PfIcZAozlaMZ3uUtKgUy6hbWvik6Uk3inemT/k3t/bjex16O5kN+EpyIN
mFnqE4u3f4vR6iSp7yysxQx44UpuggotsWeaGho9bNAF4ncB1j1tIkM5E46A553sBXTQv7c/R/TD
btguYYtQluoGudSzqMkOpw5x6HQOyvKaqJxWwFiDjYuRf4d/cXxlilZUNQnaULqX6dpZnqhk+bhH
JQ30/eg7swEyPZYL5JL6C98qQ8g0571i16EjiEErOMU6HICp1ihiXViRiweZfwZc8ZUW5zBBqfZD
7yf9aGFve7h2GfG62+OpwWP+kn9LCN2DQkrEg8phxhjGMRSyPy3YZO1GUnOk2TaiJtPCywKyI+Xi
17t12fpTVPOZ1KsGKk6H76VLF/XB+cg+aKNrBfFqLlkn4jguslqg/QM4FffGUtR03W0ramC2Bhmv
lejjtUE2a7h5u8XCowKJus+dJLXjWX61mYrbYMVgYqStmulyP9zKXcJmlp1EsLf3K3+xteiprIic
BW87pVWc3rpsK1isqUL7DukRMwGuHoyKyPa0XFyVKuJ9WyMBH0kPVG9RnBR2l4TxEdVr9j9FIkG1
fok4VuKIrYVThGnu55xKUEAhNlOH94BlA/CSUUenpOK6xlnQSgAtYa6BT/SULT4fhVhWUdHRF3kM
mhuCwo3Krbq/6VS7dj3D4ov0/o4F34dIkqty2MbFUxegQ4XoLLGs/aELU99mx/gyC1CG0/GT4AWm
Lj80X981JbTpIKqh3pRgS9jJ6yXzHprpVxyZBjuss2sYObWGeuWClnK4iyqyQ2T9hfpJVOnLGzgT
jsBYnQTJTTWyGqOuBQB3sW3mJIrTutND30RaManwqfFEvvObxsyuEyD0oQgZH7h83UcX+vwatW7d
2oA4e/cMfEWrJLsYFMLXuDrDxVA5vHKd2adGmWy3PEzCiNBi6oo9YIZlYMzob4Aj8wdZz/31Ex4n
mLhyqafQIkAnvaXWC27g9/Xzzt8UmqhUPinm6SDug1MNjlZNiBEqUpeZe9f7mu13odAmdARquQdg
bRLqFo3GX0sfluZ/wAYXOrEpEf/G0jKmlLTwk/pPkfXOhjomXyRyXw6DNVRyxt1mPKKmKdmy0d7B
dYtLTj2z/qVda8J6pHrAGUwhL1LnTKe9gFV214FI4GPC1BecyCne7wK1NSPYSi0h/0JUluo65eNX
02I9tY7u1U5htn0Kj5E7TcUXbFo4eYGwpFSByZCvrT2HSBzHPotjn0lwbWM1rcu2UBqx17Rn78gd
WSeORw3T/7KLqZO9sHH3+pQt6vmI88/KwjSKw8Rd5jRYEKuVpJWnAA6827F3ckfJDeLpGaKipz4U
WPHqu4fvqrJAzq7Xb1gY6tMisqaC2GT4YGYr8qVnj1ls9f4X78+UtzZt3Ax+xB745G3vyehY09vz
tkifAEc/8RJRWbuWPiv0PprPlXaajkpNqwF5gixQqCGb6yxb0bdjLbEy/X8Vr6ZQwrDBmkVTVuKC
5NMV+2Oya8ycAsRYEKrBPgHAcHbvPEf8BOL+9ftkXIcv6vfn1RFLNTWd1O7T+NLyXRuJnOoLxkIM
yqJRUB0VCP4STc2VK/EGtPX3WufsRqvk2ugxRxWxM1Y6o01af1Xy9SWOtASqKVposFgfYAQjZ8RI
uy5TYVsYI9cL74vfAq/bixTdQ+/jvPSV+mgDeJ6VuSyhScPWdbDiUS0SjhGajGrc0PAemHwjH0F7
G+8ckUNfpBtmLCiE8ZdbkyL0s5kqgC7TAeJtJY3aWTWn5ktT3AxxP7j6Zdqdr15pHl+ScN0huLY6
DX+wYcWYoeUFO3v2A1mu4GC6jVzTf6BffEnDskBlZwjPX3nklbpzDQ6On86O4yz/ASuM725OnjeY
jA52MEhwHmyFNYjJ8iyA0kb2J9Tg2RVDFk2c+6o0COimwb0uU5JYO8NTRp76MgFUcHyt6IHY3Qm4
7+11fZm+Jjmiv/lcJ49+60Z4fZAQgVp2qGCZ+vMfZoibZCSWQDUyVb5kWkFbx8W7aiJUrQZMhzF+
rOyKnlleCQs9EDo/AmX/px7Lyfq9YmBpIQvaf4jXDCq36+SylJTZd4Y5dMa2BCJhBilzCLeUXpUR
SWSfzbqnJl7dpnGzndvuXjMr71ZXDu66WMJEQi2/24m5MhKG2wLIGsNgQE5UR//p7G7m0BWq5CCw
/RxU6oqy7a53FPVwHY80TWfPtaa4viQeDGRE46PQVDdmHP+zLhxWiHjeDkAfLhMcAww0husYFiIk
SatonA3RblDotbDUlRtoTtO2knfr1KVvRQR/EuTZpUjC//tBR2QbZso8V1zcZY9+f3auDuS5vsb8
DH2ysdKuZA7/GwNBFnN0VY80Ii2yMR+SFZQlHVl6gRg6d+7F3+USYEuJyNa4IAUvQvvEmtoW5haj
/65l0EVzM9FsFX9V6P7slH32pajSHDmrIbjLlFDwtNu0jwV5vAbCgrHvw65lr3jpvhb3KD/ibR96
jJfl2obq0TNUfODv+yXI5ux61KCY9DNhNyeMxxPaOW0yFSmJymSbldGfB9qckOR6GBaVI/9Slq3w
MGnr7uh1YbvfRQ18yDG9fYZu5Cr/lJp2ECph2LeFHTcOoIggN6gr07ZgP0Yhdf41ru5yr89EP+XM
l1XdCuEE5yyrWwvhKTj8OxgbHTBlulj8z42BT0RST0pos7o4tyNMzJ8mQ4wWD/ALL0IzMjUcrDGX
V+f4/1VyiZcykAUsbCTXKzuUYtNWzt+Xits86kSj/R0nbPqloZSqcQLBt4W15x0LbAv+A8fHpga5
Ym4cmnuMc/J56jXY3b4Pc0D8H3bExQpBsNOUNC9+FshjX7CTI5LADMppS8QEaHqsCGBxHGMz32lR
sWEJrkXyF95vF8Ub1oq2c5Sn2rsgxj7D/vXQsK8qh7FRNbqfYCb1VqxGNnW8BDpDT5tiiu34VkOM
5xGNE+22dOdmm9ymgtXjvsxhRZo5lAkx7yrQ6UzHv+o3D4h9pLB6NZt0LtB4EtOh04xVTxIVecz9
q/5136gHUBwSPngJakmu5KEJLKuE8xDeX1LdVY57AEkdNa2A3jCbmJVdASYqxtY4R6A6hBLkRW1y
kxWAKy3jGZxneXUBWYQUJMNi6pLoxFjEV5jp50MFrhdd8uY4FsfCoWOlj4KIhqUF0oxzEUNLXEf2
BJ+IF8vy8+gMVtvp7Xfb2I8BNCQjRC4NeDHCHIHSIJKLfuoy6Kg4qxvzgUau34UnWlHSGom4oXmA
sWMoHkbyIOcvv2sVvix3rtqtB4sYAGsEhOi3sD2N5jUxtzI03iPU+8YwiUgNCgnc/VKvbeSyTNXP
rdrI1i1W5vClU2U/7bKDxoV1bIJsF1ONe9dBEL8BuRpARqoveQcNr1NIeZ5ycurc1BNjo+djN+pG
MpfLUmK/4oDCWclGOWfJzdXh2M1mhrAZ0kX3x8PTzNOkMd64PBonMUfYkOBrwVq1EZnc5jCQ0Ubf
vGiw1FAB/8IkgaY608ntYQTvDRYiYajFF2ISu7E7qtPh0vEobuBFpzAX3PIme4f6ervu1tWgNeb6
KzmKgtkVbx+Pvb6mNgb68GAP+g1bUzF/IS1T1736R7ybZC8ozlTfJHpQAYX80WxgPhjrk+UrFGpw
rV60yEofkJGyXAHUSQ1GRnO9GTtizAodfKYaaYL2btG6KLv4QU0j9kdQfGQJJttbFmPnnUnEeQhv
Wb12dyoTe8BXXBfSYra9BqvruAWyoRiPOXmbFOFqJZMuFrX12Ad3NgRlqAl7a7D7i3cRGEEREGaU
GmNBv8cOKeHaYY36ynJJoHc6dkM1N/c5fXD3zZmFL5J2MUY/ICvnT+RGtxID/wpeN9nWFYn8QR72
MMPNFhT9/ILjtT86bYgeu9ZkDdStrdVqVW/ElPudl7ToVfLDUYUyKxkOl05IvDGB+GtFXGGr7iTw
mzus7iqBT7L7Bz6oUId/38Gh1ZCn0uYAdBHtNn6Hse9jHX3T25uE3aB3g9AvS+fzW+94GvrVKsBj
hEUZiafXSxBYGrm+p0c+ELG01abG5jwZMvknOqCMkFmZNqSn9zxH+xAjtCsMulY02HZPQHU70ku/
q0rWvvaSdAn1/9O0nEQ+B8O9TbovTvt/0IBI7fTZq5H5fKzpwdDpFtU7a4/X39SC6i0oX0f3U4SY
h5OlaxE6q0R8qvnoj8aDZ2pirV9VehS6wRTzjmQOxpKA3FncSkyyn5hxZAB+RFiONpOl9y7nYm4w
qI7GpZHfWKvz1dtnfWevJPf0ghCCXySQB671IXdjtRZBONHWHgbp/wg4J2jeAjFx1XgEYpFHdSqW
7dD/y69iUjZVRuaQdmuiIDovQAVCVKKPEibCrzDFbcpk0untqN7/N/KUaUXu43ivCC1aRb8fEr1N
kpMwxymAj3QVhO0uYkAco86/ydD/LZGHxyiILHVvfCiSJyAOF/xdN4eZ/58xvOH3uBzxXAIp9k1r
xMF/jUCczuq13sxYHbaVSXdnvbxXNQFsMx0EhZ84dJTk1tzfUZQFGudaOHdChqzddauSD3wrJOE4
3mA6cCarO7YwMAYmuHTsR81ldepFlO+YJu5mKjm4XQOtEteScqRcPMSIhhh7o8kGrJqCzE5oI3vN
eQwGqNzhjkWh2mV2HFghMlRXa89vi5rLKIfqDPPoYL+HwGkXCTD6UJLZGANUgBxwEPX3Ar0e5TaH
2k4MtJcouoWWQ0VAxxHrQ6UxLOZSTag3eRqYTyq9kQHf0zHLStvAmOl1kkBA6I2HPLtuxDs68ZJr
ZsTl/K7BN9lxoJ8lg/ibSWGlXIF1unLlFfsUz9/ya8sFHTlb0syttajTaclSilk6PmYwIxEgFA9B
3hghZNnQDez4DR0iRdmQnNfKF4IK0V8CIhfPQ8meCgXYdk/DXx+DODWdjx0YdzK3fOwjuE9ao0DS
iyrddHdNsxt17itmfQBW7sZxZDI02vy+fF0+3bkN+5bstlbdtwF9QSO8x9zihaU3/+eVIDAZCh1w
OqDaEf7mKCEw1goJ+AkUflFy1utFjoirdzBXSP+k+cCSkQ0028MlysT2VfaZTBcBJGoL/wXE8QeY
I/v9TDScwrWK1P3+4jPT/GmJzuYO5ZpRpyreWRfC8C9IHhqsodKpS5Zvgc/SRaVRd5DNd8o7aolJ
DDUuH3JQHbjKh4wv7ZDlMOK7zP916P0mz12HJtTSOQEOife7sh3deBGUjLAJhIU04vvjtTxq2SgD
veFUmBvvVzh8g7DnTLZfhHWT8GsAzRhQT3Ukn7P6cDwEJr1gVG8471niPIhS+uebs3tqTsL1V60w
yMIBKDhSODMX0jtiAtPb1l3VIiZSBKx08AbBapFcpQ24VYrdl93dRn3v7aBpKKOB2j2AYaZMPfsH
LnqKcQK3hXNgWo6qUukYf+CThbZltYCtetxR0IEwqULkWjkI9MAdc+8e6OSyPlZL+cCJsgmuMx39
q56vwW+96ITE0oaDkQsFcMm9wzT24jso8fBHQarU662rVY9jeIW302lvmBn6xn5+W8h+eJitYy42
sd4AjxaAjz/rNWFo/BEjN/bFzYxusWHNAhHwuVhbFxkKqaJJFDPQGGMEEs+P0k/qPQwM2Ji/S2Yk
f9mD58Kvf53VN5OKtfttDZJJ43uyz3xbLJBsjes5cNm+Jdn/M5Ixj6VFVm1+FS4KtVeSBAmKGhmD
TgjPaCEAKm7eI/ghEP6PHPXhkxdB0zLJEhd5dLQRR+kLA7tt3P4sG0Wf9hSnpSZV0wptdK3AojAi
ye+PawrXwxeJ4oLds5ZQQIJfQl0qRM/TcjhATy1HWVL1wlo/oHE0/glu3BuiZrTFgZIGHsQavtTO
hsc2X7KEgv+lU2T8p/ipZcugxH/UkCx/iAN89I+ZA+ugfEnhI3ibtwN/3UmH2QxXNy2KjXJFrSfV
vNUDVmi+W1gj+kbI8YeKnEckZnX7FMFzG1S5haucqOgVj//OzfURs48Asdyaq3KZSh/R3qW1kyyN
lGr+4FvOwoGI4+68XbSoqaZGvbLtrwr5eavgfJZIQmXIWKHCp9Or1jDcwvfrr562hR80O8QdZt4y
llWyJxUrPY9gFTHrEf2gtIakloaWoI0yNkTjasjSfwqg6D5Hyejsli+6/Xfm8h9OT8XAHMxjGyJb
QmZZMsPnpopi/2rc2fLFBf20P28STg8or1n2MwkjCkyC6ZW8R3kMzGV/Q2zSsCp5+VaaRUwp3xNC
ReiBdATI4eHUgD37MqukfpvYfZza/66tlvxa/bokChtDOeDpqGnQiLe/evjabM0Yv3lSDSttbYhO
1yrphwiYENzT1BogZHxkgSDs55rOO2uPUKzI093H0qk6Zr7lZEH+xOpIyFOUcTKUR6Xt1J/Xvjhb
zK4FXRBc1iWU351RrnSHS9Rsf8u3zPqVA8v+rpLCrW10EAPAjeJvcMx2JnDtqy18a2LI+bQTSNUl
fLqcRcYWce8LEZeg9Bf1Rq6q7pCCXeICR1wwlfue5jCs3xhxxja168Bei/AAp5eqHYRZ3yw/xRiK
9FfKBo5lYYVVpqFCHvWjj930Ct69V4wzc0F6XPGcZgV2rCpNnBwOL9gFAIsVXP+AgQixAYXYABcf
x5EKCR1UXC0zC37JVx+RMMaiWkPgx3tt1VUB5Nb/fc9aCR1FL42kiUugFfvVo0g35sC5YWXjQGqU
hbE1p6cTyWW6JU9kHcKswPJCQ2mijorpXwH2EuWWrYl3HuZXuHWkAQQ+A342HTTqJBXrNubgQrE+
Dnf9fEHU8bn+GB72KbArqPbeLPNKCvDx2ESKDHxeZlH6M7s8ZLfGF9vjyLOTjruhq8Y0/pLju/wg
ZpsJ2jFLE4RoFUvWA3CdDqCM9UB9kYEB2OBnmokEYdXtNpX6iqbOQNGsQ2utXwfwB+MtSjjyGkvQ
5iCmDVsi+kGrAPbxrHeiO0U/gOxFSZeulhASD+rLcb3fnt6MaEoh6Nzh3cBvXxtA1dTCND7yQe19
MTzjz6224dlE7FzpYIFSf0C+WM/LxrFMGAuCUy2ad5K4INZAvjyNFjb1zX5h1us9QTRcM5obFl78
+yNviNIbpPI3H9Tqf9hG2REbQchDMglssWSFXJnyM1ga5XQI6DSNZAJqFC9HK3F1LdLNIXE1rnkn
+byH6gEu0xG5GaWT5e6/H86gUToDtOwdCBNKgoE73wwKdSwvSlw59xMQ2WVBbkI92uGPNUhkVbYe
a4QotSA0FtoQ7xs++KMTwQtaVnEhnnQmE9/LuGxKUhqEjMELHFXSlhX3HlKeP0QoyaMe2ovw1eJl
w/M/QySmYoTQTlB5K+dLB/elsaFrMtAUS7RUCdFBYu/AmmBogpybhNRpOMDpihZ0+GYVwDoYBJAS
lzcdf88USI/KQRkCLP8KBecOzKqnrH/lHDJv8BvYhyAcAO8oqF8K+26xVP6NLJ2BeFtFZF5kMt4X
TkIOiXkwDzeepVrOD5MJLnUixguulevK2i3hc94GnJrIzR5SfKs3YP9cEkq/wwEd9/ApBtdiFBrF
ZtpfXXzUsJtKE6mpGsYuYtPe5NaRpUsZXQBiq/1O266dUWHYNoCYVtH2QS6GyVky6dMxlOD56xnI
uJziWQRMEy/NN/9T8n6HzgIX5PfbgW5usQ2QR7/CERVZZcGyTQG3fD19ORKOC1dxvgdEwrknyZeb
0C/OXEa92mlaMJSlYTSSJJVc87wAXuMAi3g/BPdZCz8JkJN2qK8KuFxHDz0XMieZhh1DPeVgrfH+
1iE3LDp79h5LOKz9SdW0AZ8lIpIYFgUb1R2nopjDIMECq/Wbd83FJBGaNzu3ute8OsB2THHBrpKH
VWDwT2gkDev8l7lZPzwLmxQs+QleRHjKRNF3ifcc2QNFShcYUQFKpdqJLqKGlXjAlwihaa7D1ZB+
ImJUNCzXVVC/2Jg2VNtaVeZoBUYlN0oYHq2wJW8GO7obnTWof+I+maW/2vL17bZkKW34iKQmwKnr
TRg04jL6twBu2NLTkIQM0bCe4uVkZZzwV8OHq+DACEzhkrNxSQRIxkFCuRc8fejEKQ2nisy8XS+W
nj8Ac54b9kmphRWtPgIcntuOFs8EGuc9G2vtJvYnbDJip7kccn1Vyd06O/xTlaaeOjK262USLKYO
K99oM1PWX9g/3rXNP/lUnfEFw8EK8OBeG0kBmJZf82C+1Xh/sJUDt8gtsp/MuJM5C/qhpZF07kg0
FkZDKIGxI7h2kWcJ7Hqa4MmGXBOkt6VvMDRzWjVzbz0OQ4mb5W1CaEYO6jfrp0rgy7hqV6YsNqjO
DIDj/1JLPwrOdluywzOeSIvPvfltl3u7sz8NzTifoPzvPBtJA0LqnEN4c5I1iOzZYbBDnOLGIl2t
ZTUS7YmRZXNN1Kz7+Gb2BqnvDRu/aX6lF8n6PlikYZA9nGSu2e/d+j8yK+xQJ7Z/FWDILyUkYvPL
jyyjWhjXZAxI6ttZqi9ZPnWD5qD+7Ei+fRRVqZVAPoel5SR20T5Y5YvQ1Hdp6jZq7fb90afP/8BE
sFG+WzB9DhDN9VCZULFSYnxx3b2YaD3CyBjZHHnSQAnaJBYHUMKw0TZbczfXo+dl+xFBxw/8TW2s
/hYgvcs/evQOxFHe/yjg7bNpHj1Y/mYK2sMkardQZwf+tNU34I1bI7pz6BGwqnDNgkUmZ+9/ZgkP
AIrohZbHvr567lJvYcJ9C9QXZPw/6R8eCdZPmVEGT4D/BrpvsJvffRnRnQiYakSaqsfjPa/UnQDz
yHhybEaT/sEWCsgRIku5Cj+bS6ylS5WYwBPitzdSsvkzxRWn8lh8LIyJq6DtEgPUrgyhDUkoHpYj
SSKYxPHa+ep//wT+X67IfP1wNuagbodqqKbXXrOKRHrIHsuKeDz0CCP5BIAxNxvbdyxF2cTnud3m
EJ0YJNyKrn/2g1ydfQ2KXTm/Nu+XgGsH797QonvvHNa0k8OD1JkKLjro3MFSQdqUY1s7OEWa1En6
cveVeDHltvNy1kuu9nm6LF3Ih+LoJYwldkuSRwxYAG2eow95r+wYmT5GFEfiSpOwGFrFJOuNWtER
ruh32fFsI9CesopAR9xIqnSpQ0A4mF0ADozYPQsEsQ1NpvPo8wyddvcqHGRpVickmpyJK660XAQD
7YgfezjcFQNRIcggn74F15No5TnE+yYvzgp4QB5adnlMTqeEA5AUzmWEX1srgcue1FUd2mUE4ITd
AJeT6sLzaySBXdrkBSoV7yb77e8gYcPWWtLtK2gY+GT9vRwux0o2W3OACSRZRmOHBagcg2Zind32
Qk+R5LFJ6bOBhur4F01ovLUIf+aYKCZo1UpNWmn/cyzINSt8zRocD7NYGcRQ5GojnnyUdTRYWeP2
VwKoRG3gMxh9nogTO4Sk+fgo0/GWltAKqU+XtTs6q6ilu3Ezo2mZhRxNPtF/E0RbREEusJ+TKjSF
Epo1CyT7MPM8tNfRf6UCDtoh60Nq5S46wbZNMjWUk7isE0/fMfkxqcCJmn/H6XBnwprdauSyv4TS
MmLMxgpi3FAlZTD55Zui2H6Q8wbhTy974CaXltmM9ZXDp/vORp9JlWDzqRaOKE/CENzeqwHYZP93
qZqTlwVf/VDV9dQeaaHs9LTlVDtIQt1mTqx0tVIlsQ8ZjndYDetNJtklCGmmdWWcecRlUwAHyx9l
C6AzBVKHPeKKgWLqdgvgLyeoe/MQfaXWvRa/Oj8voN8WzEqzcr0tz/buSxMQ/1emO1PiJXqRCxlq
OjjQk3ijYLMcnyE2b8Qb+N1crHeeCtYgNLBqAEM9WhHJbNGgDoFIbli1ee9CXCa/4rdNNUK/Yk9T
c+RK2TXC10nQhz124Q+Zu2qQlyZNA32Pwmhc6TTY8HOxzPBWnpwl+VwMoi2VR0fwbUXXpN7VqO6m
SXQBb/yPHN3x2kiVjHaHOJsbjdkeiJoJ8lFJin+mdGKX0mps4eeR8r6XdBQIectoSIsSkr01IlCK
/dEnt5pheFvbLsZf3Cj5CkTk7UJi+YP+wkeCfwLlOYBeWp6QrZy/vH+cjyiyyAm3lk7xl2Qs3qEk
XQvqsivUoNbdQ1Xau7g6JiRykmK+TEVbYiBkUqXfWlOqagwovXhpRCzUcFHyr3BPaXKVUnLCnDMX
4f3qzL/8fkM3yKDw0nKMuuckuVbtP7urQZZPtOK5MDpsf6zLY7aM35zyX24ItmXEUVR9TaK+51cD
fV3RmIHYT8+qSdSYsijsSgnAU6kfnlCUr+vxqqlABbDeShDVRJXP/+Cr7QxcgD13jG0fUUwEv9FG
i11OForNo2YYyy9e+Z1bh8nQmXwiwncxU62g30d/YYlsJMPrGOZMlybYgodYknZwbfq/Qz3zQWjd
RxlIG4idfCH3NRZdAiYgc3BulwESVRncP5CeHZP/GlK8rKgTChrHKTLI6gIotvDxtKjcxrbdB0/d
GVhaD/K43bnVbwqTSOz8fYakxQndW0cH0V52nWttXMAj+y/EcDa5h9Ri+gnSapJnjOmVOUVPv9eq
XTkC6xVO0wZMVY3/cSzM73Niumio4ULTv0RzQ8KRGRiVlRq/6bxNOnwzw+agCi/N6iv0lZg4k3tD
9c4veTmKXPKE5M2b6zJRUS0eL3KMKju7Fk5rocUulFHjM9F5zirbwqZW0R0gZyJwOrFADLlX3J8e
PjKoKQQNSB84cLIzGTvifz7ixxGpOXvjN+coBKBrn2NymlRjJNB7strrjh+E5PpnldwkVfEA+fjz
45F17zwW5DeWGJotORC14PWNdhckG54kRwEPSGet/ppmWeZwPZaLXdJeywUK0a5vQfyT4ZGkKEAu
1TOQnkhXS+ceXvfv1NJC91Ml62wG39XeI42991Iilp6qCfXmVHz48A+c1EAAsPc9JnlSiGLOLwQA
fyvA1ekC6KBAah7/Nr0Hg/GSoBuIha+K07xm2N4RIIczuqjJarXYC6ndvs0ROhcD6vgHn5BtBDvD
Gqg+txvpfTYADhVn7viQjifNWm2IDIsw3xnaXIhwNIaMfb0wrAsbwDzcvhTfKUcoYYbZDIHLBYeQ
2dd2FSsWzTs6Wvm82SnaT5iULfTnPHETE9DvlgbD25e4ftSUAAZeGOKltcdL30vCAUSx/qOBpziV
O+5vy4yYY2OjFE63aiJN6FF791/ZNge84S1XmpQFYyPvcmItj4jGptA3ej0EC5xxwYEcx2nhO00E
WUP3SRr7xq7v3gSpBSqR60lpZHDJjTUC6Q01jM4IfA+CgXdRplxRFsROE1jIX4Hcld3KSO7b/OCn
fEfl+j2AdKSAeJyZIhY9QPSx77/JRx9YvLaQdq6bcproPaE2Sj0hMmCjVYMJcYHL49mK96gR2xiG
hsppA0rfk+IH6TE8XoUBiRvyNVLCh4BCfGZrLPCUKSr3caAWBZFGFQo/CjRo12fM/OaCU3C0KlNC
eUtc/0M/wg1jWU/xeK0ueofGW74ciJlNV2IRKLVEN5LqMf1uEsLRDP2ba5ULfdAtG1HROJ+uCKke
LcjACQnY87odz1A07cY5VvG089l5+9ZBHWkwmKZlEG+WVzW95WlkW4atCfLqgeFDXjXmx0QFqCgZ
bxR3PHSTWdrFQzBwxH4etbjRDjZioA9oXLTxTkfdF2u8s0uZCuxyz04re3QW76XXZsVYwaMOaNSJ
YXcjq4BCvklGeYKGKxzB+cwHND05TpwuoGDtjhoAPSrx0uxqBdw5VhPNnYtkzg3rrsMs5etkHwin
FYGPZcAD51xcza4tZ0HGTVE79uhMoRK4kxLOrmkwq1JmwRGfd6OrHPTopOlzsh1z3CfcmL6Dgy0e
POfgcOKm5xyN5obDBCKMflCUptKU7jzGdcJJtqnp1LK5dgkDYcq0eGWtw+WiFln2deZdOqJHN0+7
3xCmBSuFpmvfNp2YKHWzspE/+9pacjmRcZ2dXNBeKHiF0g2/l6LqkV8kDSVr5GyNaTuswE8oBvS7
7a5c5ifHXMEKWFzXggMJ5xYuBKumkM0HnUx+hQ7DZCA/kECQSi/JP6sAvNENKsnfHIe1VQhl0h3K
Sy3GYc5h+dugmNyBtPPdQyGGryd8qhAg4SnlayRCoQjom4ZE42ZIRTkzeiLSXBbfjRMMtQxv4Bag
FUADqjXJ/tqaPLHYG+/2jBOIvJgiBKp+NDo5aFV6NYC5ibNnvL+F+jcq2JuKB+bIMCPducd/PJpD
XcM1/zo5nI4CUUlUvOTlB8WSvFPRxEAhywgz1d4IkS+6+vQFWixUc7KtbH7JBkIq4pTyr2YFiQ0Y
uNrTpbvpWEiclkaaqbmk6JGaroQQKzWVCWOJhsPD8XrGjOeL/0NGz+01ZmUsRCy1JaS1lequjFU5
UOuxj+z3jKJtT9BBQWgabmDSQJKL8KbkR+MurRwiFsUYJPQ19r4AGIbPNpSkZiGjsg42KO34YE66
iQgew+CvnIq6rc/lyIurajjYYmCSlCHWm/9v/fywlkJeGd51MxfV77+CeWqj5sQ4juYLZsNr4HAb
QDIIWV0/0aXzZ5TkiV15ZQNBE9QCNNiFx+WtfS6TNfrEvPyFj0dsaLnmnX7snw7adapjHCojBqTX
FnNV7zCuXClvLkwPZZr6Ff4xcNz6zo7OrZBTyZhnnAAQMddmlqNj9894ui+h0DOcbnp3n1n36Rup
c2zNjlVmANFv0oDbOKsuaBwJjPNsh/42n+zSJj05w2mUKxDiL235fo47keDzRg+CzWAZ7PPjoBB1
TunaUPyq5YwU9o8GAWRdSjpj9kxg4YyDHKYXwJGBrPIFojz8html3hqQ1OjaZRR3BrTw2a3e8jAV
rxBBMi2GaIlb2mmTUzyzaHXb1/zRQR16ssPJGPTH0T0zmDnwVYSVWc8L54sTvPp6IvKkkX1YNlCN
7d7O8UmNgw4kPlttlZHAt0MNiEy9ecdAo14XShMV6RU7BsiWc4uiVROKuU47Zc8vc1dLvPMXop1e
YB7diV2akXM3hMmtBib5YiVXCdm3TdYP1Dk4dOd02hWrhBbVVGJa+Mwlkb0IaGSIOxHgPrpSVz92
AlMsl8/va1U4ae//uApIHy4j0tfh5YRKAT3z2iFRbjFevCa3qLUjF8muAmp842TAIQMYpJR4N/Lk
7WTXwmPlGotkRXRLEFY6FxAas1JHukK4nxDx9KHWvHRubm9BItz/te+bc6Z7zwvffFvVFxSKgI64
HuzOjMixnKnEUOCHUsnlin93Vi9dEM4/2Up5woxqQ0EE2NbgJSCrUVG2hvam+ELmNXntlOvecNIm
NKJRHCceHUd0Zqgqh4hZxCux6eVmYmBNdvzMmKveTDcWxin2G4k9Vq9frzyfDCyaNVG33ksQ4zrK
FUvdQk9JhKoZkSDeqX5yIDu6cyuVqxLgdG3J8+CteJWoTz7XcmC9WV2qEvKg7m/4m8iimAipljWK
1jumTY1zxHHLNuAWdifsle4pCv/a2aR4zcpu16VOvnVdNsjrqs7dk2ypKQePp/y9Tum/tlsuv/j+
t5q/qSijSW/D123eid/NJe9YaibUvJtpBb2xS+awOhvQ5YOL0sYxPDSb6Avc77quC7lIcJwOu+ci
q5KinpGINbPjns9sNsKd43dKPpgcl7sSizQ870Xg7fFzQZVJX+P6rWNNhiO12GmAwD6XdSEW5C7Y
rXvCzeBytY0S/cqAtbPUiGyFS1hD6wIh+fEw5BCbErf6ZE0r/oIHLtU/b3lX3wD5Y5+Au2h0eRWv
Nl9FJpXZgx0dREvBDos2QyCu2YWPm6uoKSx+giXzPStn9mTa9hYQ+iAtircGKlf3TJ1KbyZlylfY
6bxBrxdFpmZu2dy5aAzOZBGM2Q0dMdHuOWIRPTAzjyFVJh2RfA+e+1dFobb1UgAzDdx3cpNiPCp+
eWJrEiQZb3AxFo0DU58rP7LBjP15ubpmleO4tFHI9tWRjOrrPFDIBfR9NgHd3GzsN/QKaxohyUpk
exP8LVbXzMFmgtPvZU65nL7boA86M3UHKtfi/79qATuh0H1yNT6C6pRRibK7L9Ja9Pc1GWm/+/6+
tHcz15IW4bfp95sFoSt3X6qBa0IlX9ZFYQWzOxYN7t5cn4IVyaCeJ42aJzRY5EU/2VfGTnymWGI3
wdCcFYhcNNvkZS0xDW1Q6OdUHzz700yFTEMOLNHLffvzVdmtKjgkAwzVUCDENU4ekz6msTWSGYOT
3l7pfrnEWDN/n/mOrCWWKC86dp0jGSPPnQHq9ABDMPAjkBpKJhy65Evs7LRgvUJ8LYClhFHgwpBO
DaXHc+uHlr0ymsmLc+3b8ZaHVUjJQ8yDAv4fVCI7QP4+2ojEMKLP/6m6xzdYazVC7xjE/8liqSt7
DRkDCsFU+PJW7uwnf4ZiQnbDVou2d4P6g9jYtOIbrE7WX7ETeILGgVKtn8WAw7vOAXV/zoxChusZ
BR4l05PJSTCfJG4HqzoOwrM8/tMWAUXQAu7f+rWZ4mbeFv1qblCjgKqHHnouv98K8wjXNhbtjqM7
4+vKYPjCkVCT/oVLiu5SDy/s0T8wnRyvr5tQ2MM3wvdsqx0peUGkmoKEyyLbNUUotp4OPnBByYpx
eBSWR1NDzTFgsm9nLmdoa9G+j1jgCxoCf9ae7VVwqHLoGo/27Gt9SVyR7nAPSlUn3yp/DX1P4QZy
0j8GceQfaGUv1WcwoaUgPqLdomwzXnZ6oKISkHLgWLVdJD/xOn9qsnGB82fgBADRfEaGhF8EdKq5
cnPkqYd+672coP0By5y/rnOVQ4ZafK3ELrlWbhWhnusdeUEHwk50Ky2sAQJlug63Mh83X0ftyXp+
oBsKP9DhKwkiTJjonq8Zaa27PxQlpenKD6GBjRjdMVcbFTjoNruVZFMcmtE3qH+w/k+5uyMveVp1
+d4So3nMeeWWldiuog3ltng4hHAoFTARXka384YxqvtoggSfK4D8KB7va3nXbdpmWAaYVG+x7NYo
kwRFj4YqHzvNtbi8UO9qCI0FPqtuSQ/bl9tVc3NgM1m1XnalBAk27Niz+8LtaCZFCKwDabUAJWfL
dS+ybltVIcPPfVuusAZlbrFMG5jo1KLJ6Q4hGT+UkE7hbKZLPzHaREHuBxuoF90hon+9u7XU/l6K
VQdSnM++72kuefF4jc9HEGe26Rnv21He2xA1E46ikazeF92NGYkjp4MKivrlck8b2iJEMoNKzsuP
Uuvsfiw/LilZZrnFM0EOWQGkOsbIbUa262p6eSx3PlN55ylEYqVmAprirEr9Qc6DE8xC1SSAvSbf
bOpNBpIxs9DAn14n3dVABlMAnAnU9IXLTkRnVHn+R0ro6bHaHx1BirtzficMh6vFw+LDaIMTeb/p
OteyXlgHFZ9aCrDuqiY87Xt5Ioc7rq7B6HMNcxpBJmsPLdaDv4PSVGtPLG3bN5PDQQUnNQ5gEfep
WRN5PjqooBh/AA8UQFza3ZaBDlZf3URz6n2jsfQdWJoop2hi99XNPTdkDlRqjHLpWZl3/R5oWtht
TibR636kmpdaO8SmnYJnh2v9V43Ys/J9jaaPI8Hn0P5YxyHvPXGprERJgkDNaHpXXNsw97Fpzof3
32tW+xK1OZvbGb28OhwP6gPifDYBoOLDf5AhXUVnQUG6vT8EL8n8bjT5TR43EDjeKPc+VLPr9WAE
OYD6vvS1+I0OP9D8Vv0mes/rGpRiM5fUMRB2y5T26Dn6Y29fbsConNv77SYuSU3imkWLUstci3cp
Hz2+Bvj5pT59sIQufee0t2nDadRP5abnBlnmRMau1HShZS4SW3gT5L7n2EVaAqGvxeCWyjCX92xI
CI2WmfvtLe24lAJdSW2swVh+xRVaYXZe8uuMQcVcXR6Fj4jrAU8TXhH9JcdbgcSXT214e2mTE7iy
s198JCnId6Dm0m7Rs3Qz71zYVO0fb9wMFEFue7AQG0XjwUqwHjCf85o6Xra2U5mRtExSuwx3nazn
pC/MNN23LpuasHsY0qXUqdhGLYzmofspO7SkNeZWn3maFwXtg6xOIP7P7w7ZUNc4e00P7Fd+SNXs
yFnyvI87IrfYkx+eE6gYN1aakcivOVZ6GkVQ4VXakwloYRDw+JFwIjX1O+rgT6mocEV4XOP0AJGC
oGYHQCwZffOqkYpZ1nNp8TiHG7dtLD2f4ON37Uvj9pMwGM06k/0cQi1NDtNTDsp9Mfz499j5ZPvw
Gvi9DvwJSYR06mICYnNkBfmQm4d1JZsuABEaL2Y9emaa6AW9PW3zQFPIJQcV7mYlfoEDhycoRFKn
yT7mWt5KvKTBD8e+zaFAzBoHm+YzaTwUwGYmKEh2AV1eilmu75zo2mMddRxGVL+AZ23HEH2g6Kr3
7aLuWXTveCGQoVQssdvrQhr9NFLHj/pRpn8rlKRS77l+zA1WDlAtYWMQlILoTvczbvMOYxwcAEM9
H6HFJ4mp3W+OuUgoY6DTQS5BiCfk+llckYay0ViKFgaGgun16wEHpNc5SaxaVWpZc6sdl5KzC9J4
cGknunfVvoTWwPFCe6r9NA9fTPMrAc45SwSMWOyyW7C66Llg8+3/wooRLzx6ZjLOU1evXaxyAtxz
2HubUM4AeBVlLX6K7P4KQKHf5P4Sr1MOPy7YmiVySDSIOjDXR3sMY3jJBFQ0bspzVB02kIvio/Ib
SzCOaTtDNr8krgl0Yt/sP21UpsrNg8TfXdYRxDQGfSD5qmxhgbbyjwqwpvG3Pm0mgfS7cycmlFV4
0D3aazaD1ct9WO5p8dQ/dv6zqn75Gc0BZdk5f+xSHxq4Yekx15IST2ShCjjP6EQw560qp8GA8p43
l2tjU5bCZUDxzaXrYcKHE8pQsah/V6kUbJfFkIor6SBQjEL6c4mGnajSZYimHBJNazynQAMAmDTr
O5apTrzsPEXbq5oy6sVuFnzun/i7JRr5cVh9jWoj7ZkQXVupPVxRxGgxPwEeZ7ocSLjOzAUyk8pN
HiugNL62VwvshnObuOfWCtYljixsfUKV92bUrZbl4pDISSBFm0AoOUwouBnD7TJ0NAxkzmV/+nhp
WMlwOkXwpa4d6MWwh/XuurhxcY20lFsYHtEanMeNmOAI6Gjl7d5gDEjrnEwJLo6ftgwB1SkS5qcD
K6oSdjVJVMQxMi+ALpUxjW2vHDwnrtfamd7J8c1ziHhtEZnDyz7d8PcCBF+76/6Y8b5nEQE0cHbI
nVcmEhFJoSxKjrvhZH8d7eSgaHmjhhkoSwT3SJLvWqUL7v3Kzi7QplSnOtuvccHXtVdGNBMuxTMu
cuz5Fb3ofGXt/uT8b/LD3OCQuSsPnLA/tkbsXSaXTZ8RZW9660hxXuBvj4+DFNd151gyQYsTSWDC
Ozs3TiitZ4vM5ZVfM2GDAWJgOWDkORdnWVEvVPSo9FNvWyz4aLrnRPCFRZAuE4pRzScS+JMa81K1
4RKGtFhn+pCuu6W8bCO3r4f1CLzNgDydVIfXUkuwGImB5x1dJ9QkBkVvKeWOT0nJo3zA6BeO7Qn2
bgceRXfOeXs+muBdmhnuR0fROYxrr4LwOxF3M48qXIPFgB5Z/H7G/ag0qxHFNx9D7MJvA93xJ38e
fiOWcjm0D8kz3r02OwXlbAKEgPcopYNuqTO+34xoBmAxZAbeYnPWB1UsMyTjn9w+E8MXfGvi2fOz
+FwK1aI/ROAg9Ey0R7zQeiRptD75tKjpc6KvxBvTqDkfvh1I2Ccel7hvQCkztJqBosrGu/zLL8zK
dGp1KgDFtCfqToFMxoYyl5mGYlkY3XE8gJI8XV1MLlPq1BJvExy8orAfQ2dZjiqWubkc3Qn8SiNI
PLYiN+S7mCBsozokkmmG7NiFmd+ntM15aMUeOYh3EHPlf7CqPyD6Ma593ig2UvgOY3uj4wapTegq
4FXS7m0oqqiwO5/pDj9tJofG5mwpeA6gkerto9kuVMlYxrSHZx19SbUTaLjAISBKZES8QnE7eT+t
uKqx+Gqr+GaQQbT5pdqcFveyHCaWNqiSLYxOK/qZP087MZr5mPH6xGdTqL7Q2uQ8iEi9OEuFmzKv
6JC1Utn0LSjx0gALreh5vUMyLtfhhCTvtdcEQv02miEQpUDSl+GIMWqqkJsb4oKnf2IvE3+3oZkb
xihnb4TvliMr+o1qCUdYxeqhbJ/tZjpu94SelePOPyOD4BpIW8NuPPOwjnn22w3OP+pwgO9XKQ+f
j00Att7LJvVlx+FQv+tLq3Hr9dOn4V+ClMwq7sf/3eSLJzLWnWAfWfcJuzWvNO4kr3LZOXlCvQoC
+QODk36YrsJFhbnFrHJtTtfGv6nfVY/pjvQcsaF6yv+B2Pu/vqMwlMLPxXvCS96ScQyrXJWLj78a
eI6yIfkzeZz733YRSL+WtvuTBONBVJcRGYcihl2yZ1chTZHEoIdUNlnQH1pC2bM2HYfI81asOeT2
bK+WB10HOZXeV/GvA5u7nJ7TROAqB/clHuHZaBkxZDiYlPXxi2GuQY5SCXF/JMVJ5N+N3XyQ9fIg
BmCcnqaAP6XtBi8H3Wg9wbRwsGyMSQM+HP0mdVAFr+cdrKng9HfyJSZ4BrPRZDqwHDI9/nY4ptmx
83ofimKg/AZexYTH6iPKIP5VLtV8bjJrMuZ9yqLmRRhJyiXLhiEuqrVeruPbJNnM1p3mbBRjeRnk
lkS1+nNx9xUiZMZuyt6L3NYS5Gcufi8R2AEhjM5JCBKTp2v3N5rk8n3Kg8Iv3lDgMeDlvtBaz/I9
5t/LJ5kCGR6bMvztvizlU24QTcDl1h5eOSJG/0AyA5Ql8Z7dw2Tvf7JBQFZmDNkillHEvJYzN52k
7bNQB507MT/kjMKeRe3qVUEGAZaOx8Xsf5oFRlVsNjH5EHhf6SGjPiXh2bAYCFbJhGaV+B3Aw4Cd
0sZW9QqudQTfHo9bSepU3horPQZxGTyQfqolal++NFWBQRwTkGxnpVmDqHPqc2aYYeat4zevdrJR
JIVM/ZY1Nz5xf8j9bsu8ZmhZnjry4O6edZfGLP2XPZJ22VJ5wOY6O7+Gt8DaWYIsXK4gPUM4duH/
6RrkWwq5KW0VrldP+oa5FqLhtb8Pon4WrZu71T8OhPeyNeRQJnEzBw7fRrCWyvpbQpsJch4bK5x9
GsztZuw745lAXGxR9D4Cp0p0VBD5gSSoMDSgN8q56hfSZOHSSB6gnT5VQpH0vJ78jsIIcCHuuS1I
QzuT9sZvNB6JMYbMS5bhZflQoQABe7cRgnG4ZVfyQcq7Rs5h/a5azPDPAHrn4xRJ/nMyZ88qF/6K
/B4BgleyUdOFmmhkbsVudNt/Rzg2Im19FC0QZTea0Tw7zpor2LrWKpbFuhhF5meKHLIgFwDnUEZS
wCVWnzdKrnmpk5CuyCVsq8yZ9PJadrzlg+d+Knc/I7RkDXepJYQCn+qkBDAjM4EnGNYgRGzwFPTa
I1tT8qFIfkILLpnww38IJKmQWu21RMW4YLJgkrFLCQJCdEyLwhuowxT2bQt6iF9NXbX5XlauBKuj
4qCs+eE8O+U6GULPlzirNwh/7B707rDL7iv2Wr7NZVrzZMufLw90SjewJs5/biI7GJrFMzcRrFlh
JdMKDQlB+qNGcrdOoTGW4YiDMc6wuNOh+OYoXKzQ9erDO8uRnQoqTh4jz7LZWjZU+/Pn6NXg6iFF
bZ8Zvij2GdwdLNe+X+oWxAtmFtRHlPW2rm7feG3vT93Zh5bnVPOvICU+L4lJXyctR2P3EuZbvAja
vD9Pr8YJbCCu0aH7FxbdrE55e0XSdqsfwTNGPbVCusQzZMrSc1oMMF5LiKnCJgseAcTO3D3G+25K
VANvOktWy3RckS41W3BBFBYFFqi5qx8AdRrnGxecW+NrAy6VLc2zJxnGW8SlZm/ycrSdKF7YlWDO
CaD92gKffggrHSnOK6zhIt0idveWH5NOqUoTr06BaHZeeIX4lvN87oD/09aQFZBSaDJi+dH5qt+e
7qTdx4o/y6JuojGeeev/aybmph5ZlpvN/GDsosD4jGzYnFiT+vG0SrjktzMWSVWNzJLkFAOMp/E3
14BjEPw1SdGB/qbdcZGFh7aG/O98d5/QlvE8rsFLFhEUfNkSKfpAMhwsOCsUrVu0cxHKE681AwOe
WV/nvEA3YNBHyXWbSyos2D4VTX+UpWyM6PX1ijdMB0hZlgm4hn/Vo0TrnTpFz9tyKDf7pQNvgwcx
lIGU/1hNIVsR1+tSuczOLdY0fmmiD3Sfke6ARgbiAdOPmQ9yDm5NEsFhHBnpmAEQnJLeG+BIxKLr
9+Rpf8Mb0QStGRR35ZxwZyMpOgferZrlbziBPib+rPGBE2EmLsmp5aiDHLpQEsovlziq0EfCMY2n
+fKRvo8dLw3rfCP4wyzYxEQzkzqfBrfZql8vthlnAiZ4Eh3H1FKPolr4GIR5tuSEEbTvxZpBbnbq
A7BBGqfZ8wz5FdnOIy5GK+pTuGY3N7SR7WlmX6+Z4FeIsF8yCCTkS+qKD4mBG4AoJjB75cruNYOz
V8XTDLdHf8jALqjP81DwLjPm8KGhABQtQJqFl5ox/f/70gDTGFw/uTfAviCiYKjBzrgdUQou/jb+
7Do/rteUCQ0YdgGq4FsA5saHMvBRBT1+cXJf/4VLlUlC1a5ZBMRxFl4495WrQeueDcVd+c9rtr+j
1pbr2fPuZhRBov6H0vHy112nZvkSwa781hAuGYZ1F9N35pBtdkQ4PGwUkUdDqVJq4bGT2rD7qB36
icK45jyy8cl101o5fxPBgBXVUNNBDZurb7rGVmWc2DOamk8cC4zYgziwIDoAKaHq811PvX/Jnbyt
dzgqbrPg4jNbD/OK5t8hvY5eoc2b7tJtZ3LriyBdrwKghdzuXmsD9J0vwa4YNZBTo8dVyUfQiCTm
7CkI0F9WmuHg+o0IWWCHSV0EbawSnPTNo1WUd2Ogx4Wj5yYzvuY12v/b7seqTozll5Uc1wMLlD+F
uLvEi9jKBPfFfiMIS+CVJy/OCpTb4LnJC7FR7aOYqAm1tyTZCwA3gBdaajS9BIfqtVb2URKoQgD+
mWqe5NSJh7cofVuUUdkDIp19OS4zKLEB+h+ArGf0IujKUhXIEyZUihGVhNq1RtyQgYiOynvOkZup
PIEP5/ItvsgTz8jwwzwVlVefNPZ95EZ2fOFxbZJe1PnM7aU33ldaSzMjfZpPd07ws54wfIGAoyjg
0YqDPUuEFWYmZmToOsuOK3q9hrPwY0ZR1M8Y5tnt5XP1DeCkzPMSJTYJqMvEgO1q91kUHMyYnjkt
4Xe9uZ69CFEbk566z/X50Dr6mZH9ba3MkNGRsHPjTTLLUyhGsasG0ElAlJts/YWwGLmF6fILrGDf
+2rmfq17yiGHOUW2+y5AIxG+kXDOWmGN+3b/PGOQWY5eu11CY0Ww+FUvY8XJHrv7Sj8yKTP2eO9Y
QA9EMHx8pzmb9Bxm042qUcDnSoRKgQoW5FE3Ru6jNqpZAPwY3YukBMQND7so4hCjtNRStgYcoNFu
NjSTIUDP0SvIkdRmW8SC4diCYCYenP/Q+5tMynI36LcG7LkBfYOkByr/EXn+xillq+mqDus8tmAI
9TeMlxxNOXLwb9Yy2ji4Rrv/u0kI38HxMqiVn9gZkq61M/uIbDBraevI2imeO3EjtiDEapynDeGv
QYilOrURO8ko3Rw6AnC+OL2pebD9yzWJcoy17SkIn4FR4X7AXG6EoEpj4VrWnIJ3jDCoH1SO4S/E
twBXUxxI5jzhK37h90KN1YfSFcF803jKcfGsN4oEfM+fXreC0pT202tfPcJ/2/Pm+MlP5v8mpiNP
EgKs7yVl9UvdF+ucXCbTpmhCkB1lHF9r+L5/r5N05AF9kfQ9qAxvXDVowArmf32ppK96PcxvWIiP
tLU5lirHkio7EjjhWdz09mOmz8CfPfI6voEe843QwQxZ22assxWtRMW8H1n9Ei4HyuhptX6WW71G
EUZLh2DrUInTbHDDT2/k6j/zvLiu+LqzhFsCloHJzhyL2CfKb3SppJG4uuifz1gfWuB6IhhQP1Rc
X0vUY0tHFTtRhMX81dKv+HjagAGtyggnMFuV1/cbJc68FB+zAsoNcZNLkgk5gJDgfpMn+IYPnuXF
mR1Qtsz265vDxHbcr8YIlxPKxCnc0cG+Ui2+5yOjyu4grpSMT7WGzsMmk6QSCWgZCkmncIm3/4H4
u15M0dpcfmoK6w02m3bOGMhqHxD94z/vIQnfZRuRu56ilZCM4iu0eoofWzsXbi735kntB/5L6Hx2
1wOa13dufqJuhryDIZ6nUhf9O2V7JunK3hhwb7Kh8gyioF7IHu6xSK+L7biOqtPVaBhMXkK1JYPN
rwrCl34rYvMkE8HE/y0psOvdvPgNaxVieluYc/gmp89tSNnfcuYApkqoRuiahNe4fENLCRpQ5Pks
jpjk/xpzLQ6jBGltBZEc0iUmQSLTR5YP8OtywSQjtrmdnAgOMQEX0XuDM7jRRdscATm0Lr3YoK60
D2/Jr6nfekiBbylwXon1RxOQitW9UrfOEsvQE0qFo72g3FlrLPv55cllHeWwxG0IskahHIRO7QNu
0NGK+hyNXczY0De/z5cB6hJnnjq6JuZX5B1MSVgoaQeLG/Qc5reRyxFHexY9UDOozVoFeesa7lK7
SonQVeP9kXQI9FzVnrn1WQPP/QzNiF6ANR335M4xM/tq4LiiNPfiOT056t8sHb9YFzKxKUxNNWVl
dEHwF9hZcL9IFG4JQC+rB+44z504ap0tdAhOXmTeA1gAuUcgMtlAzDy/v2C9p3Doz7Hit0ogj06h
KSUZgGosHGz0J6qp6E7BWWIdQ9vt4TQPpRAfuZekfO8x1ouz4miEKhMxi+JohbooyftbZ+MsX5gY
Gg7pMzdbSXeGAWhoOsCcE8tuHoR5WEXHL1KpcCi2FeLXC5NbAkLcTg3q1bABpQn8tXdtjEOQep8S
+FG23fCdVycAmO6NjZpGSp5Vn3G8KcI8um3laPyR99CecfM0bLMseD25wGVtGfd9NJiFSwFBAeII
zA+pqiGA0/+YYsUb7ztrOPlyTbLcqnhrvrgFqfrQdmvuSE8lKwh/cikfkLJ8w9EoZkmZsGNyHgwT
a7g7S11G4SrqZQMd4ZWyrinvz+KsYW9v5WjyWd/e/Q+LnqwBZFZNrMbZdje2Gphnkl/1aCe441uG
z5+WWWuNBTUVKOZGQYAb+xBLvARqHSYL8wChI9sb6UrnYlXkHULgFgpgIAaz8kexzlvXUXSk0nb1
m+M2nSYQ9YZY3KbNSnSYYEFCqits/U0ovEW5Uqt4xgGvzNlP6vaZc2Xo9a+ysJAcxgSapkLo1lob
6TgTvdA8Nn8T+kZwxwsQbW7c93+YG5B77ki1znO52X1YzkGbiSQpg3h53BwKFD7BVItBAHqNxsU8
FqxslxPsgKy3I2XqPraFFauPbN4kIsrTLX/mwgxemufA2DhUj7iANqade89CA/OOamhW8LarLK2F
JRig+cwgFqP3ALiWhDYdKyigJY9tXioSnjvo17ysg0VRPRekoev0WrsTEaWon1djjoyZk1QsdzgX
5MZKbgPIoMf0ZsGZrR/fVEIN6UQaqh2LHd8Jr40sYsU4ywDWgND6ZXdt7iAbd6jTXgi1SptJN46A
2tYQ9msxj89m6A6a1o+nEfBgBfYlxOTrTKaXZ+avaoLRfMSzHX8AHNgUd2sy4zRdvWZjddiZ/8un
Ndf/WYqhdYu/FXNLRy9u36BovgMauJX2QkjRq/Kp8NGdqUOyxPyLxhc6RkIOFK7aEKDAyjGiepGt
ugqblr0s+OETi82Kgs9xYqaPBTief5CVvsyRukc7O3BdKR8AhklqB0jvkNX0CwzqMDrUUTIH2w27
UfLl6gt1Y171KFQ4kx5xMrTwszhfsl+KL65wzoQgA3ZP0grUWNpNIAK4k5DKUH67Qaj667UNEMZN
Dlv2U5mSrxDY2/dvCHe8DGAiLdFF/BV/DkEvoMpLX0TlHA8QEnwwOfeCcksJtFqC7yXrsPnZgipo
zBOqi4vLCoKjj8Uxc7i+dQeoe6bIsyXEKBtNFlVS1vhijUsPIu9w7ZQYJYgTb1Qnn3Ca6J3rZvKU
Uj4HAGmw1GskJVAy8l9r/fyRwAweLrINQtbTUIT526gjhGAEdL7roDQIAFmKYNSjFpTy/EtSiCe5
DsyQDSHaS4DJVprfObAuNIRUcrVU1Ou73/76OUl3EbMEQViebs5P8T8wb2F7WTj8GIZryRimZiji
Av4HvkexPfXoJBEl0PE7wsT+NFndYKQZOF7krKwcNdJEWZ/6z3f8RHlsj6iHpc6jmbu3d2m1nxRZ
ZQl93CCGhZRBm5eEdzm/AvMkarCVTigU3GrV31UqTGKgGQGyEeuPjJtdJShiXNA8JomtGK7Cqxb9
P24nLoFHjmETBZy6jEXjkrBd+oNKy5+dgxRsiYYa5ycctUSuFr93E02OlBYGaf/QWH7+zhwDTg8Z
NSNd1Fc7+loTNZR88wnGauCBdkb8fBcfSxhinkbKRK4agxBLRBIfCTsP1IfRekcOUqiEi6T/EGHK
2f8oftJuD5QzMiB+8k/mPbvWM9J4jxYJKc/hq5gCnzgxJbtHb8q711ndME8DpPriSzf81KmLm0SR
cv3NAiC5pMbN7k8MhNqmkMU3++d2hEBW9cqEwvfef8Ozc3RuSf1ahwLZ5wgRFgbmvtfbbbJ/MGpm
WN3Bj3d3lrKX4pV36qYpS6/32ORFxp2T6i1CDo9gW7WULc0jdzX9rmnCkirhvfJpBu+JT9hr21Fr
tGnmIu/wO1ihVCBava/rh4xHnZSGQc08ypqQ3CbBz0pcV2NzC2AJSndU7gE6qSvdUi+gkBkUrulv
l5c+WePNtGZt8kVmZtlq8GDYq8h0YciJmTwKIjO9DmYyxLQisabJIBjiIAHU4wisaQAdJX1E8jOg
9qF5hBSRj2JFmDheG5duzqkvQHALgd219slLP+a2HaA3jV4flFErw30Y9sP15gwWSsjyYVo3+D9e
X8wPNoO95mVyVVhhNIbMMeOo+x0Ym/i+fU0QhVEZVk3VBF0CTZq/vb+P8+I2E0yRdipMpQdpPUnZ
8DK9I18ue0Iwn1JVj+EsUA7JUa+T5cFRNeHuY7kYcca4xCiTsXtTsMYIJNIC8DmIZ4E3+kHSjhgm
7l6BG0XU5XaRN67I4zNj7vLrlJIJCT4TBK+9+NSy6FDxnzo0RIVuEXN/LcKSGlqZ9baf5Ex73Khw
+0xKNv+ZyoR8a+q7+plnhiUT3eBHUawh2ZHa2NT8MeHlnDyMHalYP16wln8YcIKaEcf0MT+gVY6K
52B+vqmZ5N7xxVqbZJREB1dSGjWiOFBo5cFbOpQKtg6bz3YmsWKpclTshOH1iT/W0fJ8ynh3BKFR
qB7dkKd3lluxdc8FiC3v546bmWJ5WCIhCBuqx3Gunjk8TuMQPd/zNAnRFmhimFe+uhZgEfVzSaH+
nisQjHVuH5xHCGfZp+JFW86OyWBwmHWXww8ZwCjAIhQh70k23WYxZHRfNjw/e1wzADphyiAxxo4C
kyMNGS7+Ssv2tXMED/Zz0RVsbrVqV9h7OIXQKVSbVEspkwu0O0DgAzZmma4RZ+W4mVXeVCWw8Kfq
pacrC/Zaz9Z0QHIA2CpmgyXDDAuIYHQgfQsY8inYrS6jt/q/OoQUNtJESVRMXzB9reTsfTtWDpPa
Vm0Kcg1wrDMD+yo28OOBQSmMRT6FVsaY6mYwhaG6D2SQlVZlS1xGjc5iZ5PXjR8ykscDOdrNGFjd
YRE7gO8BxN4Z7+1nawGe6+bFtfjwJh45kTDe94qLXwKTYlemKq7EXpSpOOT9MVEYamODv/RzZYA3
xnEfZ/d6VVJn6L/yiZHRhBvrK2SBSOyjuMvIQGzy6nLWAxh/q46Zhy9FV/jh7K5NZrNrQyZndYCW
yzOOtrTg6sc5tZph98NgBe6WomH0TratlZD1Ex2f/GICMGZin9esmqMo+Y2kntQLW+WRBU+/ehML
BrO86TdfbUk0LbrnsBzQ04F74vBzlSKbESslbzZqzz8aOodtM2Ob+Tow5v9xNr3+frOQ53fH/uRR
QmdujxltPNWar65lGmk13bRSzFG8gUZkwPbH3tF6RrnAP3K78ausdjpkPByNeIUxJ82B/I3vd6cm
WTn/0Y68SD3dGajbvll+oarcLF7ewBhWvjvqG2D4pnxbn1391/b8DvuhvS3ARz8YqQ5vCY75ExRl
HEBKuS/wW4AuI4YnroIPcSNXXr9esxmw0sBYYMYrUrCuIieAzFEo1IYci1HUqnpUZMw1KrxofeCA
z7Qrgw/hAK3fMjKsv4XLq7tKo8/82hgz9kDlbhQDiTkapA7tv7xJ8USMI//CvdkkC9ELxP7FXTe2
0y5FT0+G8NO0jE52jEAdwnZwvdkHQXKIRytAiuTBcIuJk63GiumptZ3MfMcnoEY8WFPGd0dg/q+9
Xx41yvjzCU1AnLss1rHQ0TsMSXxPROui5Scescdo2VLgd+wVl9XVJx6dnxmdtBFIMavIxIU5zr6a
T5IYfVllrwnkmWfFLQsuGKW6lk/1w7EdqmeXz6d+hoYPzL3xocbDdKVw6lgSc3DGZOhl9pRY22zk
H//R+Ah9CT7MEXI4Qzp81tPVwHWHiDLpbRR/9m20TcYFc5esU5bQHE7zqSfU6QzMjtb8RGPGHuSw
RgjbsX/fG6k5dzNZip+phywP9bpsy9nAPXXpA8Qnvj58RH1Avf0q4iMJUtg+/gPB3AsE1mlRcZk/
JuEBq+FuLkyFJGHyXJnu0oZxh+6czv0VX5vvn+EPyEviAwLAtCrLS+emosTl1e4d71PfsOCxHOZt
6gL+jI9Lqx6QN6fNy9EIipVUp+Lzt6IeN13ty7z3vBgFsmfXc58imZ8jbtGBy6Kd2xeri4O941UA
QWieQ+lUYQQALiTvqjXRsgz5qitU7uqdQkPaxFHBlUCLJXP/FY4FQ1nD9lYVJcxwLC75AGNPF1iq
ompxxuYhTxUHiR4SQCjriqZfxWHCxENeR27QYDfQpAb6w/SW7GT+lIWwlKx3vjXjHiOIJXX4uk4r
ZBTgsHQCpO3lf8gg2YVGnlsNG5e0DoR5WtiiEiVQMwUCaZgh1GasWz5bkvGTBgRPT+HG5ZoINY2F
gY+mNeZqJW+LpaQoRie+VRYSYA/ezuDYRRZ7JDWQXltgLQ6sFLsQy+tGNV1JQ1OY/qi+o8nHkTSx
N2NjObMb5o7YnP5M+CB8QXmUOKwsFehctFUyMryWs3XQEPExwTUEs3BYqiiVTvY2hzO2wLscjyj/
3VefUN1057KwIyqNtKLNF+8Lvh8+GRLC8revmPpZt0WzjRiw1bhXVhjlikQpVXgU+Y8nFMbW56aY
UqkzDRU27k7lGoqpLdb7slEo1oiDHRIuzf1qgjipiNiw1uMiqsSoZgkMEa4hWTKrrtPOjePJjDki
bLa8YmU1xMtvbmFLE0rFVuvJbHqEWTlYV4kY4fLnq8yJGsHMmL3ddw5Li69sOP4FsZTOM11Fgy1X
1B8vHqN6pKeUcrYTirmTfM0G0Z/clWJBIBvguI8fROK3Cj4okWx+mctHay7mwtNunzTUmUFFOBGm
EeVaF4jEkGf3Fnj13laQ30jTbz9J0bOrjMvmrOGuZ9anjMety9zZbpdL1x22kMShr4+hZ8G0NrgI
/ChJtxr2e7/DMeyzgqt+rPo7MEIIa3bu60Dp+oauSNzN5qyFJuQJdROL+mYuCjbvUWjD0q3BE8BN
LOw7A0BJp9LIOC4sB1jRxHrXdgCK1JwAEC1eXYHo43ovYIcMms4n34gCe0EGu69lxEWvcj9jGd07
M2zCN26X96w6rkpog3MQujkKBvaB1SWvDV1PzXKTUXzt5s6D+fdTyVUfIYbPqF0pPP96LyR96aHG
GmI/TZA5AIqSA/b1clrrZEA9rVAUf4wNxHbUUZDz4FuFkX6ogGXJOrUGWI0bvPc08woRQMDDdTnI
JNkFxIiZJuwsvolCzZPHxlA0lnV/F//fbaQJ/onFEbDKah/rRVBl/u5YHV0aOcjd8w96S3uQjFHb
e8HEONPXQYAcVw6pVqlMaobuDu/5j5iGNy1T0DVJWjHO+QZWcwyECRHdTnZkCJH4ZehOJlNh9wRR
7hXZX7ub12mnytQuuXjBwks3ONu+5Nt8luPDNbf+EKGdbOflT8Fgx+YsX9p2zcAtqrDZSZydEb+U
1oOOWzSRW/ev0KODOEN/wboLeQnz4WaISZIEL3ksKFKjoFAKEhNGEN1MwHQAOhfjXSv4QN1LrceX
CTu125cQA0qk2fkwWScgQXwOIf8VGq35t0NJMoZs+CjbgIwN0NrzZY58QBDeLoL63UGBTnHmletP
vgxqsl3PsIvz09D93k9jvEVsW32aDyG7hhsnoT/c26v7A1A7iPMct7FIwaPSU1y9aKOrLaQQeKyx
50+MZpuyK29LWFOZDAiYhb+SltJMspa4RlZaTEgiZkkK3LtMUWeYgZOGHe+WF8RWluqLtlzFcj9h
1ywkwEd5pJJKamzB5nmb/2FrNIPj9TnE+SgjL4f+BUOuWYIbsuJqch2XMDwmP38tg6wulj2iCiVy
P8mqd1Fxo3GyIaHwxMMcDDWgoJyfQMdWT7cjIndaqqxPJi4h/sDM9BIH40THAPBVM6A6dDAztRYA
SSt1u9F3MutcuwC4qqothPiqSz0w/tfOOcydjCSy3ZQN/iHarhxkDLpLfbnTF4xwI2yD0t7rNF7D
dl6mo0z/JqyYAnDiz3pU6LEsOZIyVsdWbue7pyLMWmjhnRPumFSU8ui3LgI2RJ+fhaaz/Px18yWL
Eo5pc3EJD7rgrAzw7YLUu4ZXQgqBYV+/fHguEKzwZW+U0e6Gf+fd0a/FcPpBb2dE5WRMqQ/0hjqG
rZJaBeyj46gYZkK8K9/9vT6hKxldmSq/oCynrgalbTUy09wI6Rrlfql3ZPSleKr9ZCaaZHJhzkJy
8BMWQiwCu+CcQS/iyXSeEY3DibkPoI5EgTvZMiJya/dnZzw/APBiAqwEoGsDET1i86alc7bd528O
aNNDHt1ADbjihv4LYrDyxsVg146xTadmKIrEq1P28DdlCMLPMQMSlWWRQdLQjokl011ggtGK7utl
HGPpyFJHCHIHKyc1j8Zr1KJuLLhNgdSIyW1+xCJiFY5aSvfIkvEyppeT/cpd0sN+MxvjatAqH6He
w938HN95aHmsqgymkIceECpJe/j9FuRPBZGtFGnBLhzl4yWAY2b8jS1XGhYpK/fsKiB6uydrSoCr
FFwh7M3Ab8R7mjEmSxJ/vofS6yf/qn4Og6ZiymdJNBtTVRGyYGzertXG70EHqQc5f8dOL9Sjwtdy
fi4OgqNOPpFWP5Ei6TAhZLmqdWQYHq00SI9K3dt5ofSeDYWaRNLkpnAfXdGQw+2QtnFAX/Qf3Ejb
onmDNWhRB95FuYumjXOm6uICs0TizELc/9gWhiziZCGuUaZ0G12WDfEy5aPmYp1aJ3OlmaQHMwBv
93JO63+mXaVvxfTk7PhnExiuDUKYMms5LpnwNNWDiYsgcIyjrwo5ShrIGU2sqKLnbMJxsSAkHKEW
CD2Yb8ha3dGQ+u4CFdpXOtYKs3hgoVzbPV8yUq44OlNx4bzmpQlfS4m3tqABWnq3LsBS0QzdOA+U
zkvDzx4xJTRpQ60LfBq89QR1wTz1tcaLgNv70+s5E4u0fyjx3RTcmyw6PhZ5AtevYDK1HLlMNbAW
6OVY2Uc6h804PgSjM7q6V8euPYv9/4CcUuatCWEGLcQNMR1yUolXxZQxzMw5fWoDHp9/ZsmDxng5
zgE4YCeC5ggiPSvWMhM6LmdW0pqRrZWQ+kddsty1aukZbcoJYKGE6WQlhRDKVOMMxntwZzD0uMzU
tipR9IN3zqCdf/gUIdYZ6kU3liEadZ3gja/3FBX8Jx0RprUoJ3OYhnLPOivv8Tkuq+51/Zczdwas
Umhw4Mak2ImiZocwNTiaNguBKgAEA7tAyXOs2mCrgQjO3jQIzIi+mN9B+h/5tQ+kGT0gtSxFEioe
GT4CtYdU4lD3dF6sROOLR1anNYztBt2ywpEDuOOiIMTGrT3ry6iMzp4GuUVRmTUeO/TucvydS0fW
vWCD2cLPpS6wjie9kns8kNu6qv4Zv2c8w2KZEx8r25CswTznc8PQAxmR/mDNih+rRZoIkcyW3CFL
SqRc4c5vJASe9vSzoB7fc1MDUKLphOyLKjOcahP6cnx83dhpdToALl8ejkzwiInrBLM/G7vzV1Ng
2bsGb/2eytIB1535w4N89eKc5VwpIzo0e5th9h+F+Ua58B5jd9j38s/EBvZPx5sceWy5uqonBFYy
4MTSNnByPBklU2vvFVfma2AUxjqCodn0vixmuhvN3uHXCVYHXYl/0Lef/Ufu5SZNLFUdoO2BYYyf
RIilBYU14P01+yVuIB0fINCGfL3+4wTCjgkOIL4dspR6c9Kh5AoSiUXIT95murMixtTgpxFWf56v
UzHLLpktUEuefypvQAJWM05JImHGCVbRwqSOpCm1O1hsmplrRcnXWhGCzw6vgpbbdgVC2V4a0NDr
ClCOvbg1R7nggdlp2mGHUxAEVsNyYUpYMmxMzf2nkTtAG5yHJOhWtfb7bs3ZMBtaLSa8+qD+MRmN
Iz1u9JQcsxvbZRNpP2qmfUxlHsjkW0lTLlGm7eCwx3zbX9Yv/j1IfXVJErA2JJ5TWhVCRu+kjCAL
XuAluEcmXmqar593J3/UcQYTGhgfwnrirjDzpKchC0GTdh4oAdQV7dbFhHeiE3YVKqNtSftzMeWd
IZpg1YkiB/f6pzFwgFlsMKHikMm2jz/QV95tgVtAnjExJU4gyhkHLNGDLHNugXc4KSIZ+3gtjXNO
NFeCoYYXaOUqT/6ZKgWHfllyGmYenBMCOcXN+rI03jy1cEte2XgnwFc2um9p5+Q2LCRxHudQ0gHx
lfXRWMBFgay+q3OMafmsNoFx0OhgPzakfhkXc28S9n8+kg/BPFPeQVuVkQjolvkZIa7+SpgNmZdq
dNC0ILh9b4b0sQr9Wcs5wyqvDGd4Pm2n0Z4fbFX5GI0OLVAaigYFyRDE1nElaYai5iIEWml+OT8k
eNVXj8d0i2uBKzrppgoSchAUZJOHxjqxiRDBZw9lGaDml8VGF2MSvt+6T8HqVIDF6+Eg9c6GU3nG
y0ASsfa4J6AQpYtnJpEaF2VA3gY/ZZ0YPAfQ8Wdrr1X2GnR66yTEY3RUDHbSYbI5/RoYD1xjuHQT
t8pW9LEx+zsVqpsrR/r2RBEh5RxVojaSyi3YqRc2Wt6Aw3lbAo5NfTS/rTeOwttMQJiQ1fXRRrA7
vJ4f+DqGuH6bJEsmwbIscHpga8Xobt5l7UMMIz2px+DpKamQzK0edQcWRFFE5oun3wpilnNTMXoV
KM87liHNHmHZyx5icNV0F7vv7gyyz6MZIs8C+srOtJj5E/U7uje7FS0L5Pr5D0gg/JlkPNUruBDg
4Ld8CieFoW349DMJOUev9hoMlr8TrUc+ZcVIZKwI2hr6oSEDrzwYSlcxQMU5qFQ5oNY8mztIT1ko
cyHRcJboZGm+UyDCWuguMEpjfxXLdgwAsyCOlNjsnPNABmpWUdm02XHgWK70PrjMf7ulEqIDvuT9
5JHSLRYxdejpN1ccnxTpnt2NsLxZkYORoPt5Lv2DxpzaIOp9XLsxVEw9cyx2EwMB+KenJwK1w9m6
ZT06ZtLh1R3FAo9T1znJhkMmVKNbEgNwr65uiYvDILZn1Q9m8CtscaOAkbeuOgJbHM+lxBeQKQ3w
PlAeb66p6jX2cQb88Ct47dQaLu65wZkSqntRkSm4Irwp8x3Kzch9eCfhKa3HyMvdaVtzpqDM2pJE
HJQktlv8Jl3xSr8ahRecByo6Bm2vLuZL1CR21PMa7dDNOKHEgwL/fm3v7aRZwrMWWQkwMTeJwyIJ
PByD93AXiRymTkC/vz4Rkc2zK0IV6CnVwib+3zbEqtjG3gsnVWXTAUVdq3+sHFjaqBiOk3Bk9ZoZ
Co+YTmgYoPSMpXkENARXzrsYFyX5k7ZPy00DeU9vGSU6Ac4l3IO3Q9ZNuAD0ZusLoDwVgHZacqNP
H7wTRiuFtobp79JCepb1tL+wgb3Arj0MCuZamzY5/24vABbS0Fy9kTOhHnbpRjtk3nrvX8PyHZG1
ShXlBNO+ubuFOr2m4ZXAyQIfsk2TF7F9N87VR1F+MNgL4hlcyFYTPWr85dhFMt0zNtzmqFXxJZuJ
+BUihS6c1Bs0ZoxKWbWu8mD+ayYNG7N7bgIOB7Akr+ekXEkRauIZ0KgfZ29YcGd6JxiCoJaRvka0
F7zUz23E/Og66Z/fuZw/5Bm4ZYnoaLK+NrdH0TqPx8uq3g3FccCpdOrb/zFHWiRZ0m4mAgVANwxs
SEPQ+rIzvGlLqGk859Anv6K4N+WNyuDHqpq5CqpTUFQdNCAAPbKQkGdW0L4k1T6IKsNq/IO4JUYv
Qt2znBuVB7Sa23aMcBq65TAx6q8KhBoh/A8iRewnoi7ICx1j8wykBLlSRt/3tTSaOWATD9N+HGpM
71yqMNtJEoTCYAkC/q+0ruRTVBPN3jHVFOnm8btzdv98VPK9Eo1ZMvGqhdL96RrxWXhTQScGw6Gn
Q3l5cHIwz3qGKwpL+3ZDsTPN1yyscD+K61fu85c14F8nbYbgeiShoZFE1c9kL9FxvV8MbxENiTNx
nZT9JcuDj3AAjGagbWJyYH9jO0YWIUwJUoxXrTH3w7RIXJt8WXf07lDof2c0UsJC3VoxAOS7XbAq
DL23TOOUPzVtfzxomIxm+37CvLb1km9+rShOhFJAU3r64hEdrdLCMj/OFnLrTUHTqMVpVTCg1Agg
d5rpUuUQRfh8eOuHpOiGWAKE5vHkrQqGRND7Qbbq7LqlgKlMI3sB9/+jPyMrS/mO4BfiLn992Tvy
WL3yrE8UxbyXuYevWioCXZTFPfxlhfIaoIZeQSXdAU6JJ0tXcpKtXYo+V3YqhPEgjLXysCrQHuLl
2tmIggNjLUMU8tFCA4jaWlMhV7QMjLDakaafF+G4QEVRysGdBIzZhlxagSEo8deX9QsQ854g7Z2P
op5wN1LbE/M0irfI24FbUKVtFXHC+tGv9ZZHmfKVjx3VMMEOSUHr041EK9SHnudb35kw8Cn59c03
aSTVN3I84FUikJBfdKgk6rL2/x1d82AatoUaZ9vy29b2WFbWMQELuZldL2BetcN4a+Pcvrm/638l
cSbzfAIE14q9w7cdag9pZm5awgu+l5VOm7N/wuLWFbGFrYR+vJ2DjCyj5vs5vxhiLuDFaIArFSkU
33n4W4cX31mbSg0BYR18US5SamUpOwUZ90WpKR+Ivj3kdjAMtGOd7NUwtWcJ5h9a8yZfcdUlV1Q3
4QS1cDx6WmL6qyDXYdTUMXIY/wAQlCh2LABg457GWTk16f6kzxDWxSIaBL6jPo4TrATzXKEp8oeY
Ke/m2aRPSJCzPZ/1zTHYiiQRjpSkhfmlv3Uq33ilGRFo0ptOy3bdIKyXZlRnTGaXZfUzDQMLXlAX
erhlph/bsgB92XIzQ12jd/IQq+cA54IpbmQBcUm9OugAnkHEqp4pZLhjgHBbZgvn32O1vOJjJB5k
SU5ab51xdqKVYUMd/OKU5N9NGsWA8hC/7UL1QUEIeL2sjJq8cXNfSGMN47TbZr3EJSu1Y4FBuX7w
UVSHnrPpxWe5p/JbN7Y1lJXtoeL0dofYkfEHKxQ48nAy3paOJp2gsF0mz/wmu8F+POxK5bVo6k5l
pR6pwflOuK0wWe680/2v1VunprTZEuPyULNoQq6q77dRVJ9io7B/tJBvb8S9BCpMBW6TcgnH6nUO
LCGTW4jXsTGusIxabYBPv6SNRjdzMXJ0VQACG6A7JObKLBLoG5Sz62REHwGrv/xCeUEb2kYDLvXh
sE1ouWP0BRE3XI6Cfg0tzXoW1+8WZGykJ/O3ZOD3gQq6VpIa3CV0oUyhjyLzeFz99BR6TvgY3BuN
CKd6m3+P9+4CgAakPvXcm542Z7RdOWbqLkvslUa782Fa8j5TRhIWYOx0IpZiops1pBCB2ggWrfEz
Kujjc2YCWYbqY5P3lIqU0M7egsuXOPX7SKcWKXoUPHjh4xp8IdwbXtUl37nf5I0j6jhC4gDIygEx
1Yzl5wMINcEZrJe1A9+nH+NofGmZ16PwxdwZZLh2DzNfea3V8Lg0ydJCu96JXau8AKPx6pV3kq7B
idswvRIztyCxlkOHjS5C5jQDG9s6rcCkF5i+Ws8CwCNihlswpLSZkcLJZ5GyBig/mSwoREK6ZNGO
PMMDEnu0ZrJXPstHmHxpl5asGBiaLurrewubyTdbFueVcDv1pTlT9BHf+YC+r+f8bOM6PcwVzlf2
D5oqiLUocfmvWuiAg/PWdqZaAVxhHm3QTQ6XEuLSk6Ixk5J/aWjRVCSGT+4q5eZPZGr0VhwFyR27
zbiS9VYxJXwBV8LSSpgTvPiBC/Imm3sLMDGWtob3M4GI/2L/opdIjr5IwmoXxhCizDyehgJj9QIS
Pvu51BMhh3zt+Y542AHLI1zR+/TBVKMN8DOii0aIh6oaiH02cmnqPgBfjz0z8JhTCifabyixyFx7
CQPJF29Qri5m4856l8X8iOZkwXBynrnboqrZJJtJmfpBl14FY9JNbsLmsS65BR9goCz24PQ47Imt
1yykreULMqSr+llmzfGvRW6SRfg035JKii8+1Q0U03URTylapB1JgXIl0C2mqCGXj8uH3hjScZXf
A/asXE0DJEzh4NFJom0hpzzmbm+EinwQJ8VwBWQq/53Ln0tmIDX/YFdHn4IlVG183NpX5xuIdTIg
k9qSzeWxOWyrk329lzGw9kmICpEq54Z0+6G0E10ABUXycOLddrosuEwVXHztc6NTqMeruK0bZW1e
lUu/7OxTlo5pSC58cd36PWgk1MId3W6e9W4wD9hQD4YPolTVdbbe+sIe0IqsUKvTZAnHog6rCZby
/EvXy9zwDdI0fK3rwKef4j0Fvb0fBLk8ZnC4ehVQgrMKredBPR2JCf23yT9A6TZF7LXlBFXIK/y5
uHZB6CLOcOuYVfHR2vX+2gMB+UtzMaxELrltaLt/+df1j+eEF2xInbkmZEPv1/LSDAFNru/AvLbv
W0FbJSz30fYkp9htogBAARqkt19kCBv+WqANpVf5Q/ryXNyLjB6uaYdAhn1jF/K1RufrHd2TVO32
H/m0aJaJE/qOPI8xiLE6apeJeyhHw5FXOBGT6R9JtZeXhu/ebt3B5wCbnkyK6QpKC4jmkxv+mXff
lTJTsGHALkXxCGm7TiPg5sgivp+q7L+u0Rp33CDJDDoiI9HJNfjJchq5gBEKHqqajsIN44DFgwKf
JnedRLCdK9QghD6Naz4JEv/N8YPzTWaVALaTaGaV9p9hXhaHrxrkgHkkaUjPZfH1sCjUijUq1KLR
bKSeul2MvBidd6SCs2vE/wV7Qc810bTTx2a32CAOO/y9NuLaNxVkAyvWcWCWtZxoOexExA8Zdnun
k7qOihNau/e3K/MNlm1Xa8itOT+9yV/nV1v/rkine2KHy+e+b18UIYx9ZOa5lWaT/aZaUkM7SF9L
z2xQdubQTT32GqxK6EkliWOd1upGT09YdKcKHtEfRd0sGuOnHyYERJSJ3dDkvXS1fTrX2hEtK1GS
c+VfqLxDp9mg5X5ZXm3GV4BWLWZyJOIB4U5qhpmKsNHpWsHPAygC7J7DsAiXaM2UMSEIjTmuT1n/
kYVvFEzMA4x+SONUb0dvT8DeFctqpT+Yp7S7LxTVtvL05CFqtBDs6qJ7N6cVy5ONDKT/PsFRotPK
a/EZDFsZnnM5g3aWEyYb8l1eEB1tN2hNDZFuEHZ+60rxkasFfGO6q10aq5csviqMICK1PelCF/sX
DBWzvJ/EbkA1+R2KmPu3NdDhvnC75v3TJk9iU9cGW/sMtVwPuWcGEY4X0KD21TW6mwkKWoAeZUEq
T9qcKfEArWA4hUm9ZfRxL9GKxGVodSfcALdtEyIZOootzqO93fKyEAMRERA3Aw7C7FR7OwcsLDC6
Z2so7C5zU18qDKXowqnYMSv5/QgpIkEX+BwsyQe3N7MVSBh9SPRnkWGvsopKuWZboc95vJY7JOga
6a+ZowXzTeNhxrRsxHx63J1ydZyrhPpH2uQUL8Bhl5ayXuNoJsBk5fhAKZqc+sS1+1bkOlyKIgWe
wOtYVXPz9+Gt66gBTMLvBhNKtXC7mzAnSH1/ZkGQm1Rxpwxp9JS32iWN/2/+RvtEaWf1aeA6TGY9
LVAE8+8+aJBHzh3fIakpNDLW2Ep6jKSTc7CzJsPUXgNcrQ8HxHe8/Ehk3ma1ToKClpzyTV8fhk4c
VDZCiGa2z1M2Dsn2maqCBmbgo2Fl+9YbuFOFCut0lWObM5gPRw3Er1bE9e5lrujXBmxvJkWfoEwm
xindRFPHG0npHhVbkAw/EpHdQhUcLyAVDmrzgK4WoDRsOgkDMs5H9LkZHjT3Mq5gkTlaK3OrraxD
K/aySiVHJ4b1NP/nApv71MiF9cKcxiXUrV3J+K01LM+GuoU43/oNkmH44+BLbbTZNhrbJUJgGmWU
CuvlwxtMrLVsdxXQ4hWGH0ohRJzAEEsecKdccgfmbfg0g8PRO6fVMqK6+FyhLSJ7vf34keKoF6qh
L6XZAahw8DZ8CZgaF1o6oRktbcZtZEZw+ULhwC7Y9dK5J+dCpBaVlB2GViyPjBCkJgTmQftU2PkR
f6rDuTDXx0GRfr10EecNfe3B8p67ZA2UfG61zalEPoZbxjf6sebBPFu/tZKFElq8c/T8m91WCxJH
vN/+8tbIx2X7AByvKuMeaSuW2xI5Lt63IIgcVFHT1cjL/Ay5/CK4KrK/XFn26gOKDAzUukF7oTVc
YC5Kk+Ju2QrkyjevNAcIirhtQcB5+R9XuQXiu1NgJZ53nMatb77FRN+e3ep42eYcbZnBU6pfxQrc
rZd2jaBO0ej8/7kGj1qS+3HwrEniuob9rAapvJm1GaWRBaILf0ZwWQLgpLqxn9dR+lLSQy7XALM7
9qSAV/OU3cAdZzRqtHfrPMQ93ZsIpuIBvHWeY1SKj+DbyRdSdq4RCeYrId87VfnvEPICqhH0Bf12
LJqFytU2NA93a55PvIzVo6LsiQvq2DlGWWbNgxW/BOfKWs8Sgb9ow9XACgiPIpQYITrn724TvHMy
9e1oIOJEJHS6PPXqAPp9yYY6US0R2xNGYj+/TQoqA5GMWIR6TRyzWOXGfhRjsJp7F6ltw4xC55pC
NkSuyL+7nLVTaRl6gM+9nLlLA6jFxWR9hlpAjDm3K+dF7+Tb86GbPv0Zv/+eTp4HY/e6mEgghh7J
PfuCABNNNuiRV5k4rQg+pOb8QMTagR49Wvn4Y0+NF7vdc392YI6tv+9LC7IcMD4K1IdOFZ3EcFH7
Lg+E2J94mAk4c7SU3SMeNAI03Nt5O2WJKPpG6UlmN9Rqks8KhuvO6vJCdl1u9+lPX/x41hoxJKPd
34AlKGpMOYyBQWaRRfAvLPvez4GxH78S1n1qJATO4Uu2EoX0E0fv/rz73KLv6EPnRinQYO0jqCHj
wbCjDqreOY3odcDnOcN34cP7dQjjZSqM4fYYHTuGAhS209j9BS9+ox4gGsfUMW7/BF6DjH8mmk2s
eW5gpJl9pq+p8Zs9N+TynChmCFRn0y9HCzqFCB384o1QsvWI1u0CsB8B4lSs/XVeh2pIzrDk12Wq
acPSDSpvYBdDCQm7xbOUo1IUvA3rWN1XBl5Ka67Y5f5LIFYLqP0azWpS7E2o///Bt7DqkjSRk09K
+3mm2xhui4lIvJ5tBwvPQAW0SJFVRm39+lLtZ0Z9wG8UNhcotoHDxaTmx4ynZgohKmg2dx/h7bt1
WO7xObC3lW2Rkzuyl8YAcWHOLaDJE5jK5O9SYqD0h0eeqWGGEJp4z8baJTBuTT2kjLhMCrxfBTrT
Z6SJVkV1rQ3PZZSVL6YKgvKeUH27sKQMP/DolvIbGbJ/vFnKC/t+XZlTQFGAhMyFamOi/7IVoL7H
aY9TLTuK6BGf4UEAP+aLKTaYSeBiZ6kUSkRRugEBO1JmPSAYcBwSJtwIcgBTAeSpi01zvFUyrcnE
HxFQYSAFrVsIJ8/cB27UV7x0TSf1fKffIw2yCeIdYVzqZKk3SSC26Dh9ZQm9OS/21e+P9bw1ffWe
dn5VQG2uYnNv66RC5qM63sjHb0RU+7cCxAxo+DbJ9Pvp4RmBXA1D4ylq2YGQGGVV3dWbuH2R0Emx
Abjk98W739nYITgXkSQAnv3sR3nHHxXVXcLBsRidd7XkSwGyWBQFMqIriMa8v3Vty8v480CTXKn8
2eEoUAw1JmW7d1jIQfqb9jIa749STXxgnKPeBQOe3jY5b/fkAieWpdL4INDItFXX0On/1tf2pV0T
dO7pM4GMogIoDIt0qZr3UDoSITcDlBoKhlMHpr9g1d11pEtFbKWFg5hjg6oKFYDhJfeBz5gErr+i
HAQDhAkKZDXsCn76lAe+nQr+CGGB6Xg0lds/BhemQ+yof4oC6xk1zQSXcsrdyL5WvSn3OOvlgZYL
w3mYrlvMgIYQ0bxI07A8yGtRM857kvAS4bBFd4Mb6gHX2IdipILWiWLwdEaT/J0Sd/19BFskf1bO
rg4IiXpu7AlG5EWnVGMPk9csO5TASI3xAenDTqhmhGnJ1crnkoI/ijghzzb2wo23e/h1oM8asgFF
p5zp44J77z+CJvO9RrU6MZC+5uwbsuh0fDK0s0Z4shbTH5Aim2KZXfzJGuwpqKoyoaNS7JfabhMI
yto1GkasmZaFj53aGoyl/W7Gf9PA71NEPK2W6NSTxxok9RrcCSDhuV8fM84OOWRJpa9E2K1SaiSC
Jk+/D7nqCZUKfxtQ+esOpeALluoYlAx/HmtWu71tlcBNKdfsYI0JH+26Gu980r1lAPY8/TcllgK1
PHAwv6eKNUo1HOVJWXIWtHv7eqo4ucJ6RZVWD8FwuYGQfMq47rL0tNrkv7IlQgLIuKPuCbPumeRh
cIotN75QEN+eFdEbaKAwlnmKM4I/7yhA3KJ/XkbglCT3A5XdUUhtTTujKSjjEEvnYc4ck309XeLH
yIeaOToOU/OOi1COfQR34qE752NVx+fjtWUB/rpatgqDZ21o5ZY3NqGoHzvfotmYNSlB6+ZRhiiq
dTLRVWgaxfdc/n8QhfQ2Cy8p2dOIMBTOEWv5fiOMsyIKZrDa2ksDT8XcSuJwe479jCB7ghVRaDVB
TZz45osfQ3GxJOp4cBdt1lIcJlPqY/cPSBtRMCxv9LGtgCDH84Be949WKW1In/CBpin/xxsjeskm
hhygYPuSu8rJRtlHYh6G9Cf2vrorVs2GZ0MSKxX/NcqQ2sdGsRLMR8ruoe8Xmu+9mIynxqNSN6eP
PWJhiojFAYOm4bx2uKrVYyfw0Dy5VO/OA6McrUSTMj2id2bidgcphFqxxWrjGyFT5MhNpucrbD3w
RIbrOC02uYggvHtg+wJOyN6K9ndTW7iwT1+6/+HRJGrj10qAEqu4eS3Xnq+teMmeIAZch5mEfFTw
3J1osOHLhqYzBp+iyNjRNX90UxO7CMvDGuN5JfpoMpxYnQuX2fVlpXjTx+s1cxy0GiOn7NdutAZy
ghvOKDWOIbaw6t4HsdD2pbpz22rg2nQxdIaeJo7d9hTeHsqdm7hBvj1XmwqS9+nMdYTNyI2HRFK3
5LoTymLe8KvS8roOkoAdusz1tzqN/8cvYCFlRTeOSLk/sMekVmMrS9frUZbeHYDAFIfQxYTKB6WM
FGFBdoFvwip9QZIxn/dcNSHvJDruXSiI2p9rsVp36jl4IqfCe5LkT6c0h2naFITEHD6ATwJEr/58
lMVIRLsybhjTjBr06b38l+cJl8EA/lgFguSw1rkf1/+571s5dm4Q7dh3fQdTOtqKqj9Mphsx3mSE
UHWU3alwGk7S6Z+pdv7FxF85klgxAga+W3/oOv3R8Q6XiNByMxOM2cTGHq0KcE2Q9rVXXIhliS4W
7q5ru25PZWqXChuSholViKT7AJxyNPDKQG8RVWNqY6SGxY5o3MATylxtGLI3wWUizKwd81G7bKRc
3q1h0id7VrqwczyiHfYdfbxj8lf1gO3WJiD2yJOa8LRwYdGFf+8ZxOf6H86szPVNGb+JZsY4KldR
l2RKk5jQsZy7JpO38IyRnL3Z4DYcLeNxzwF5r2m2U1Sxg8L8iFTDn49CU/woe1xYTopAC3ISmfIm
2BZDl065iuZHLqc+Ab017z+NjMvkP7qHhCEDJV/UCbSjDSY+H0Xivl++l+/nD/XzX76nSqeNkHuI
o9Y6irWSkA25qZSNXrQWlP8gixDHykgngdS7hs9DCj/JEpJIQ1AGp25E9nfZLTlXvXqVT2/mg6rU
pNwFwqCIYOtXvTvEoBNFT9bSz31OeFXBl+DFa/E2bmaWFOTflpjpLIybU/nc6rQ5ogvvR8hlHzFf
F8MvhbMXf4HU3KOERZIGYtoyFjP+xPEX3OcM8NYLUXBZU4ABFxxXJEWrHi/vPdOvvmo7W47dzKgl
uhTjKs4gHYdcKw0svbORwOLZHTnh2HFyqxByfQqtv/pVNUiyi0hvUkcwHDFqB+xDkWx3ikYdvpE0
8mfSemBy3GvqTpD+gLQxFfVexC/oB2SpSNSW/JCfY1B1H2/HJZyeYb/qdAleTSnrA23u7QJg8dcl
b5hvsz2QncMP2rvZ0p15xWfqXplrTIg3biss73T5EwjYaT9ZFhf/35eunvU+7if8raAiM087Nacc
gl4XCqN2XeqlNEHnI9TMubVM82Nzk1NDzx31IHG9su4gK880w37n0dMN9o2AZHtYw1gboTmWqTQn
nzbn4r+r7zVawXULe7BFCrn30OkT15ZUVKIfNsuDYTrn1O8rTsv5agJlD1dtvnOu96GmqoZMGL8P
P25Tz6ODlJ9NAlCtm0SJhc9c2FKUQ3FwwAd+ngToxSzf7MDu2Y1gNxeZJwOAUQA9ISlH5l8Ix/U8
tJlq790RcTSdYzjMG0z7PsXfMG3Sv9NbhXZ1fmt+tXAIsUgaaDtPhM1xzRSRgLbZbvEc+iu4bIXg
kdwDfvNL7La0VC46mNANN6oBD/Xhn5GoBzEuZyy3X+eNPIR0X6pDq3B9L//Tu0sR+Xy22sYdeF7k
V2GKnunwsNEfih7EfLgQug0pgcWUg1LhWcadxItrbc9CH4fXP7oDgb8jPkyOKYiyJl52RLzuYKaz
ewdKsV/ZymEwee7zz6NtNgxHIaPyC0AJUhmSlHRuID2uHPDAfQ3aibVredapbtTZvB76SRIp9Yxr
HhreZJQMILfuWJ2zVaAaeAovynNQI26JYLxVbAICbtmMQSQ3zxXe0YdjwqpITLC4xCWa6lelXC5c
fhMTIiWwvbSNxM2Ndl0XpAdF7ZP/42pJ6jXMNzb2BMfinuJuOGWJ7TiD/5PPRfFLYfPLEH3oQCIY
yu+Bp/Yf/2eHmGIJ7xF7DVdxrubU6Rbo/i/SQaG4gbx47hW4FibMbo08Lsui9E3VZrMHthpPq9pB
Yc04twvrAf9r1Ih7dn4+o5u3sMN8RM3xemOIoXIhOg4O4/Jdi3JiRFcEEq1KffQHXdCXmfzqVT/m
tOIi8oyDl14LIa1qkpnbUrQx6pqfHFVsfcH/9q36NgSl0ujKgJEU/yPU93XOV/J3nStrgaelOKbX
idTIMhrdeIGgzy6KunERAEOXQ3/yjUZGTcC+Q3768hTStPPuujwBy26iIeZ2JK8XWK1/rfvfSGw9
MiIk2wxpTfIHMPUuB57MXtuAI4o/gZKQEJU6DqalOJ7kxenvBWz0qC7cksD49Kc33PFkby+xXaGS
n6BRucElFKPPKxGFQ/mvzDSnD+JZ5EGK0QXo4GkrzjmKiVeDdWtJcCQiWeOPC58cW7pfyTMa6IgK
Nm+6o1o7NxqqqiD4PNGfj2Y1EsW1TLJN7LmfiBBUpz3K9VChxv3nugZNICt+aT+5jX851YXDMg7I
RTfJXlgna00rHTOxgXF8Plob/mJ74sohv7i9B8xcwAuIBGEoIAJIAk2/4tRT1Cp2NJsS/ltEf9zI
hZRHdVtXvUpdNZfhel3gO3pDJVWc9Ia2XYkCGtwnVto3Kv1Ot96wRYUVP1GYZSNO1BIu4ohN+D0E
+PVT8mXVflkqmxDYRg4hTc+Tpenrl/8CxzDRO5HR/8xCDYN+Q27EFdlvzSj1PozdZWRUwVVcekCD
4nDL+nn4MZydU1RQRd6r1VCXm3CdO5C3MOAjLKdJclhQI84azRzNJFqZuZzTm0cxBw5uBvpns5dQ
GrcrSN5ebMogpcjXzysIOkmfqEHv8EGRKfTFygYLHJRFM5kaHaA+QYYFAKbRytNZJqYg+0skbaLx
Oc4aCsmP+elf4FKb5nDMw5uqFjuPIcIlTjCx3+Xf0BRMAAYNlPGg1hDnazLSLZfSjq80o+vjX0du
PwD5YWxvI8368Tz7E8QKOFBzb2yy5vmeks/0tvKks+Sqs2BBCf4AW4YM3wHilhpVTtWPbJdefKni
Hq4KdSnhlldOAKJJkSHQgj6ndPU2xn2FZoBNeTHXfl8HmkEpCes9041EcbSPHOPdUnxpisJZkJhg
klvtxz/Ujw45NgqoUhlNzapCrOZi2OTpw6e6GcCsQT5lpksjFUEHyd2cD9OabbJA1Q5wKqx/XZKa
U5rttF9n/HiYuzOUXTKB4zQCUa1Kv0skYhgHjgiu50cWwrsmTTPPlLPGLdm7vWjgIkjkIjQhTPyf
dr4sR/9U4rmlgvY4zjnEkw33GYeqrocK9xTUIHVmcIU3W9B49QtY6tSaFedVAmlcyKlK19ReJ24H
4wPVgtqfjwYs2J1UHNdshS5FXj0cMlQ/Moh1UnP9BmrFwv2A3z4ZJVjVjEvv/YfZFh42vr73ias4
25YAX1QMOBYFKtuQffTPMYUO38VGoMwUwxByV68Sj8+Ni7V4TUJgAQZVUrhyJD9UnmITQ3MVHdR+
mqdxWnppc78W4vp9crCYrH6XdEd/JB25MZWQEJBo2qJ69kiBWL/zBnx6xZC3WQg6zOWYRJhHxr7n
nI3JaGqQOpBYCyaau1z6ddzHHaKhspbZE5UNsOUgawGf5bWXQsLY7aDuHvAcABY94Bt0Kecd6jBg
CPu4GQeSNzmne2X1Zjs/Vx2Y1izEiXliPi6T1mA9ymzKt3xIw3A9fgLaWSYu6LWn0HMRou1FzmQN
m1JtOWNAqSP5MBMTMoZzb1gGzlvr7FgSi0GK43VfK34CmwV8N5G/THzmU1frliXtWlkLsh74l/ni
Sx5zPFFsFwBSdm8VUd0J/KDMRjO1amzxrKjmBN32gMOwpqDssV0bQhe1Ffq4tnYidgREvdB1UbSy
q4R3UfXxy6KTJm5yqSlEOiQY8sQGqFBFI+yfa9x+9Z4mGby+L18hMPZ7/n1uDfBPH67TBtWcVWr4
3vFgsp9WzcoaQ5IWfBvW1X0qPMzt8KPGo+Ss6niiXZ3wjfhjeV43hTGO5wHXtJQgZnR2EiToYtXj
k5pCGk7AGB+YdH6ed+loIstOLt29u37lX/AuLF4/kE8x2RETOOFt//NX0E5CnOZvdqrhc13jOSt6
KFZTfQ1BmoT8yCguXXdsscydLg/FchcdIAUFyXMiIzqQBxoYChuxnkndddj5GcN+9IGqq31yXXcb
A7QYM/FvIIGA1vwhOPOWai4jnOdZxB/ipAdxaMLU1Bq5pZWSn/E5epH65y+TpdaWaVuBBFF3T+ph
t4eCwXKZcqWbPqYbNhFPqyUjJ03eX2OyBnu1Mt/YURnQLavLWRZDhHf0iXCOAbkBPJxgNUK2+L6V
u/a6LS8ytdZ1O0yfjJ54YvH0W158UAzm+j91z+un65ZB61oJYIwb74ufAqvVVnqw+UtJoQh0sM6K
gnxTuxy2yLgET8FBIc+ViVapotSfFtM9MO99jQ5GUVXF6nLkJXXsJhqnjcktS619SLEDNwX/kikU
RaG22ymo2zJuonR1cADCGISXczsjqG9dg+keNFwvRP/0+s2v5j+ux9a28iybDpTBxthiu+yYEOP9
kajA7ECCmuslAOqx3F6Xbs+U/x2ONGrNx+HZtOW93Pe4BMWElHEJZ6gGLIvtUjSabotLEGK5DZTq
t+QBGpgeDlI66tmpJiCir9uLPIxNuS7l+4nEIGH/UR7YooDMJuR8IdYucqsS+tMDFWo252yuFwcm
xuOf6vnGuTwCBY2g0CJfHzzxu5le4RADT8PhrtnqAGoK5W6s0eSs1ocYHnBZRolgqni5zKw+I7Zz
1eb815QEfMi0S1IbcnjTxyplYZMmmcS5qHwCWtrRq68OO6GWXvP5MqfVFUY5ZIVyXFX+IdfjkUDa
ulHP1bzT2t15MynwYIW5zudqtEx5SYK6rrtTd4HBr5D/vV4+x0SXGTy98vQocx5fpNYOtsmX0gmT
fhoa0tsO7NwsMeues72tSNY+jRhxOJtMrkUwtF3H1OAxwOntcuAInPg3j0QRi4mq8XA5xk1+AT49
NMU83LYNrxzB1qt5uhta5k6Wg/lYotN+eokEY3G6bbf0gbjxsTgywpaVQpeKehRL9bKM9SS7nP/g
0YDlCogaPS7U/zoPcQF5JzjW70AYefaf9C4ND2NQmPgjzOhzTKCjWNPFRTonNmsQIfeSiNurTwqs
qQja0mLdIP8+xB59htXhrQNqsCgmIfucBA7DSLXyls7MGj+wDWk/MJ34oBI6d7BvFshpekh3yIjZ
nXmVyoxP48AFFxfv8iRTmW9vv7779zOr4JG1GsiiTmhiODFgZjfPQqz0ti0uSPczY0K0Miij0OhY
ThdBh9daXAR+mlDou4I+UKvr3Ic68hy8nAZk5czxPJyyw+V8/y8ikHOYB8rtzjeQd4m8Z6uUQYnj
2QGOGTmQmqLMMKQ1oMsV4yBxIGEsDsw0jt6IVrPDLdvJbaHKwhGzO1quaSXc0PKiZnY5E4vSzrdY
3OsTkxO47tmsXLgzoxDjPfZKs/2iHmHed/H1ait19QCWJYYWgH1Efw7rONzMJjusfJYJdTnqwy1A
hflENYOxoCNmi06jCxQnBElcyVAl0fuZcz3h0IajhrZf4WpMnCXICF+d1gZ+cYuaZIhaXaG1ZvTY
a/hZpb9yUgfxJmmE5oWGYQeRv/1EcgKEqqgTOrYaZYRNNpmoWIFpFz8UHevKClrPwRu/nH37xJgU
u2pPxRo9aK0kG3nCDMw8A1ClDNdDWxEB5HTmeCnCNticgx31tA3oLPPLHG/oAt0w0r7/kV6qx8Bz
7ZsbG1WzhA/MpFL8TWiB1PherM72n9HOjUN1oZW3bXY5Pz7CvNMEs+kfGXaOynqmnABBKXuW+i0m
hRyr3nTgwXmULjAovP0myiHkMmVC/D50NE0WNrGYz3d+VVOkKsZIleQisvnJZpnxPV+mamoiKo24
wnWst7fEnPm2etp1E1m7tzGAcRN6+7M8G9ENJS4JEVFsV4Q0GS+P6UojxUNely0txwpKmaJqVKKB
Z1RxZgwzI6og5x9VJMReJolfb+mJh3OO0+/wjzyenG9XZ4DW5TpBC1vDsj/mWy+IgKerwUWaO/xt
Mt36unlA2tT4LBCKdiRVe4OL2Vd5o8+ECPvcVkGK2iTIWZAzTsFZqYzTRpEXCV5rmztQt/lkwVis
Usv+7NM2W0HweOBoKPy1BOo92GP2wieCzkAbckRlMidsBdVHle+i/1tBetKm693UwNrBS4RWsn5K
gn+mbhd3m7bLYUiedzDr/tnlc4JXZnjsBqtoTAfIzN0O+5cgdTtLCFcGzNs/aAhyKA9uuZwUPNZG
2Yit60LnpAdamPJvn3iaEjXw/tgH27/lLQ9bRQy/p2FDg3x/o/UunKrbwRXTr/k2057LqHlnxODS
+9pVExDbcWFU8jkN4Lvu9uIY7JvIzyhVskak+iZB0jJdyGSNiLFHC6kSBRtiAmZNPjbFrOLnAuw+
Hy3lQZCraCt7rCq/dYR706sIksIhwJS8YeKDz2EKvjBl7oAGDAXeMnHw0d8WmNyOwmq72bBJMsbB
329HF18OL4sDiyz2Cj9drteC+Aj/DJF2MNTRc6nxQGF7xLNv5wuUiv64LbERdcll7094HqGYVxZo
b5nCvJ4Bre0A0C8IXTDvmb15YZaMz/ny5CTytAj5vVg3c6hO+nMh5dR9Mtyxz3aeSUevmNCjHfZL
cFAcDTdbl/7p3aMUYAesF6gWACuWtx2Xbs0M7StW+jyKBCLzuXqtfqVjxslwpaaMz0un1Cw+BWTH
/8yBl8q3ybm6gqJsXR81aZVdfE5UmGljuTDVnuZnePTVLL1aNNojS5fbbDWY2AbO/4wuCsSoKm0n
sk0+fk/QuTwzsKoaO9qcbpn5y9riYpWL6GFFESxD5pNsNSnX0O4RTDZYZZO1cBMWXdCutl+iwuPA
Zmfntx+wE22SORB0rMBJ2tqspouMD+sabveC/sbV1lrfSNjg4JyPGuMJtWAQ8GjzpMrr83m1ITHR
glzeskh8FbYcLUWkGpxc4r3MmKvxojoF9mwFrYEZIV2y8wxgY7ae4CtYkoT72c7LGls5Y3vKBRtF
PX5KgvBfqXSoF+Ym1KHuOYp5uFjzNDE2ZnUdRRUzLQg8rIrStAUei8B2FM1nYVIP5HjEPt0/h4fG
IbIRU/Xpf70ZirCLvQrV59LzRZbvBjZl2JXZwS+4e7TO6Wu47mDUi7/g1H3m50tiNatYS36VpJTP
G3c7eu3wlyZ66moBCzIsQz9WA+DaDd6TiJV06sQHYQ0LlpON7haoSbsPi9mtqjFlhoEV0MX9rXPr
Ady3hKgSnu+ZOvy67RIvhWJthdwC47g/6lwj9dfOOni/m9ITuzM3+YNh3PMy3Vs71Dl2BsZwAws7
sObDGxacQQQaKDjs+RJnzhe31Oih8mGvIBHwAyc2IbtFNFiSr38KRNK6ffkjbvsZdlC92+Rt2Fe6
hLljKXJ16vMOw2RSSQF1KQ4IT8gYaJ0daD/2AiOCayCcqT7x1AbiOwbJT7Qy2V+L9/KBKLfqMu68
S6ww7kasuqKl0ea67lcAFJI49WQlX7auhkAm8b2iHeOrYXkCljA/MoXpolyu63lVRUFhOIBQxInT
b9bSHh7agmQwan7YTViykFs2CMUgEnIdQfIVAFGtidfLm5Ve4hm0zPs2BJtN2ZrOP86lYA4xGsN2
yRkMTNQndf6V8+0bXLXuRX/Vx77ijoL4s2gH6tcf3Y+DFai5l9Owu+tPjc9phfk4AMom2laMTpHs
Qr9PupEJJPU3a0NtqTkegPPVZBpo+MqUkg6A6Bz19O/pkkhJ+LMaE46d9UBWqyKeWkrymd8+0j2o
QrUG/GAlZU1VXUe3QU5JzZw/OnrJqbgcPNl+NeEHUi4zURwSlfbO49j6wSyGgVjlBQx38fco3REK
CQ1ehf2rKBDDNP5GjQIos9K/Rd5CX4e7nTy/ocN1a8Nln0ZOtyddWbywX3Xs6O49Q5+qXXdA2Imu
Bg7jtuVlgajW+h0/na4LorWwVb6t7pV6k8W0lK5qSchmaehrmohI+Ng5/6V/NgWmSyqi3Y7T4pLX
oiiY2K2oWpOcqeCmVd/fMzdrH/5WOctX4y//XlGqFWyfbaXu5W37+n0KAZhL0zTsYOw9AE8H2yWB
/8q4DvYUTp8PciQUMV2McxnM6Wb4LUxyCeGLaVCTVpbrdVJGfQl6LCvejh5GOIcU8fq51erypfzQ
A++2+fDK9A5JOA7iTBWg8AoMLUVKiFFb/+QcGqP46V4tsHWrq41hRJ4fj/7BpJoe/BqMxa7+IQK6
rHf/XtdKpN24QAfHBUwmc0l5SFpPXtcL8vZjk/5wj+ropdMMwVqCt4pz6GbSZ5sapBI7fkEbljTP
rndUZor6GldaA8Z60Me5oNMtlqM/JlFBvDu9dTUNFZ3wTL6oBBMkpGazAHlNAQJCz/CkDSiqdCTs
sqDluRtgdonxeL8v37KVwAmKGeGa1onsYsYtRA7bsw4IMorVZF6fEI9KcNr/suZ3adhqHe8YPlmH
tGEQT99Kq+pqWP5B/lBLZvzzAe3Mt1CXHn3YxirDnx0W8gUtMvYy2sjHqpIBaNEvPbTJRO/OxXDg
s3KgCGwkjoj1Ay1BzAEdccMR8pfiFcs9ssZvD3I9RDy/DcTI8QVBg+xgXJj8TfC0n7iDzMS8g2tJ
A9IECT60RjiyiojKvbPbsAfIYbi+ZIxnHyA6Pj7yiXShNabSp0LR0s+jm0TzMnktBwSs8/MzkmzR
evbDZ4c4ZSoZpCsvlNfdMel/mx+bmtXm0r/PQrZgnlpF192IQWNddM6NoGKQzKEVmvOZ8Mi59Eg0
17PIwFGoWqrPGuOyGd+1ceoqoTNRuiReAlMw/R5ludtUE/XFMCy+9xDT7cJHLIlrSw4PZ8S1jDR0
VsDAC4CgRkg2uJqyqsdIXXZgMxHqlMwuM6WCCFOuMrzM6RaoOOYScRm7bs+Rs/PcOMWQhw+82E98
gmUQU8YZWTjE3+tCFWZZSX2F8RAD9gazI49TO7yarOqrUpv72DjxlTSPIWQEzrOLrd0qHJ0q/zHy
uH9kvx13xmSqj68MeIq2Q4RXlVDaYCFMyol6BEtPQRv8cQTQVvO7uDdM/Kmopj8YhBor9srwP8f7
dF/8y2Yhz03z6IS/W3N/EHx+upTFEJDlSAPkpHJVzuzFo+8YELyNOUfak04kIuocsOrVL5GwqjR9
0+PGHL3S5G2yVLZhWZCGXWoZq43caPMDc9c0+2QiBCDX1Fa7vSHv4zDzDv8PVodiBsIX4wxRnU8r
1CQHMqr9/pC1g6ER5YdUVzQ8EnDrEHexuQo+sxgI6RdtXLv25/eAk0ihIDg8423vzRdnQIHhthw+
K9+WqZUJtfRFqfPWz+IB5zgw6zk4T+M6YVwmIGvDNX3VN27PSHILs3rYKjUE7lbb3CiZOLrrI3hJ
bJ4rgnDsdt48imB5NCTwv/3PMMypDhyYomUgfwddJdrRPCOKViCWDZxYTPlkXecOHRXb05Rz95xb
MXqqClnkhAVDN2p1n9XHllKTSPWqUiYuTKCVD1ox9QswDAKl9ia6nCdpaUqY3JfzqYyPRt2jvKSx
vPtijwvV7zGbo+lMaZc/26k+DA/BSVb508tJqY+e+Bd84nruwqnDq39b/3qNG5z0mzs3wthE4G4g
jmUAdXnBc4JsJWx7M9F3IC3UVGko6LmM7N3XiM8MXyqOz5s4NxU97zcU/QUbXIux8oD4RATFDlJk
5N7UOLkD7SEY3mcso/8frRGfRN8k5/Gbm1Dk79feDNzIUNbkWrtp7uIn5JfJtP2puJKYkuEZgJ1g
idS1qskP04cxX0m2cFxYy9hx5kmIIcq7ynnxMqDX+PUMF5zWtEFgJI+LUtTSBuid2zXhQlk+0jTI
4KTzP0bu88l5KpBYZQIm5GtPt2iKl4DXL7t0+v8oSIJnOkN6sAeicXUk/f8ZILUTpaIh2nP0cDTh
fobxE4uW+RYSesAOTLIdupe92mCxE8Y6Apvy5Vw4hrMcWyLdcfSKNmx17BOKnvnHllcpkr7r0Ucw
1yVgNhbecdqv1+zTjMOiVKOJKc8c1v9RIsyO5fj59zUnv3Qn0MuOLy9fAjupLSCXASOL1/b+OLTI
+EE8pGl+UhIBUvqP5Hq6i/ey7fKrl8oNXDdIT1M7XZHNlX6l4q+osW4LbyY3FlfG0eEVegCTwGMt
rpDCGpqdZc44s/kYUezIujfdq56+4OkT8s25aBC0P2+ELlfwr6FZ1CdiikrFHETrlfa38/aUwqPh
YKx/B9OUY5JxAdMBbdH/edGakyOS+XWYLhvHSdQq0AQz5oWQYAJj33YInkjuOyL1j3S8rkAAbc+j
vxnwNFt5CFr3MHoxCfw1art3KPwp/T5cX4WjWBfc80K9nFSE/DAaPNYAINCWPytpqOCTZKaoysTs
OiFuK3UQNc8ayEk0+tmezBTGOSF5UvALltggRPRWuC5QKLjcWr+qIUIVVMrqQuA2Pb5ThPBbb44i
0wfUqymG2sZXVKsr4A+exG9SfHcNUpKXCxlLNPXrwb7va0L13BFq5C+UKWF6xrFqgNeUkFbhjGhN
WHlk+8b2sqd9rsoeP0IBz0bWnAKTW0Fn4AJiStoruorlR0E7HOxT3QssxTV/NVBGMTHl6mDAneTg
XEO8mEHQYZIg+miGM4fYPPnA3lnNIuZndI4wjlE0bvvagCxzWbmjYkeJwtgnRT8SdmlnOaD96kJG
ekfRtosYAK8uZlOlUfJkqz5eohGVH25XGreCPzqME3SZnHneUzyDjJjvMQ/iaD9DZeguJ5UWzUrj
Y7FB0b1jkA0+2fORj6KI3BQPjCRUhQtA5Vpekn8X7vvh0gsSmNjnYyINGhBhYmzWVx5GXfhXKMeC
ZnRsUj9xWF4JgMkQ+NvA9X9kQZ4CzFPw3NUiti4Y+mQq1duQJxcBxvteaYaNShe2u6EeR2XF60TV
/nu/VsCUrsWR2Hum/aEtjKiuJS1fOfGzUbsMF8tLbRrom3quhUf5shBd1oGme91qy9PjdEIT8WGh
D3YTmW7sDlISNz4weEVAFBN2rqJhtwYdAdwX60Xh/kO2CA4VDevmRFy+564XeD2PpGlKEAWnDzy4
/mjI+Xs1wY3/OzyW45YilRuXaeEsHMTXmJ9MY8sTejvua3Vqj/GB4Ujlj+xdeFHWNqWOSPF5vou7
VhcJra9mmaorw8pkh/LEQXxpRhyPJgJFEZOWv1EMKcRiD1wyoiQk+kgCmFzaiFPFOmQ2/U9y6A88
Oz+wQWygt4eDm/wt7uDMo4UnSqVYYC5v1HjgIS5Npo8A7kJHpPJkpMbARKY6TEZYzAPgfj+iJ4c7
8+l9SIKTLkXgs+Syo9TKyVqrmkxFdQ3qrldK7siX0DNwHmRlmLi7NtQAbV/9lnzQImz8Q2Zg9prA
J/gDqApS37iyg6Zy3Vx/RKUxjXsiJkKf091DNoJCtFEdlUSGAEIY98hxrXtuGdw6sCzMkK7HKPQF
WOrHGW9BOmqnE8oPvd2G97JkkiMEulSm04BNYlCYuB1C3CkTdnOYEO5iVr7Ug+8iiXfFT1uxFsrz
vD1YFD+8+4m2JaUjrgVb1gB78alm4i+vagRdOMlrWNQVcuw4oJvcLA7WP5pqobe1Kva+rRVGqmas
slKfbnoRNayhITzbzy8iSlPR6dSTXuD5Z+OX7rHlNx/G0E6xOxqjcDBgg3jqnoT5vMsslDljFodI
xUClqq1eC1BpUkDvkkq75SwiiBi/SivNsrFcj6DBxgU3enGICZtK2zi2ye1XHmRUMOC66cr5RdKA
nAURInqZK1UEe9QWYh0UdpdfxRBawkbLYYaCbRq0dHkefw/sUMCr2iqGNunQ8CgrMTXKu1IIwOw7
vqWoGPXUSarTGoinOQYx1QcXOSYiMSkhGUMxWqjs/qWnjAemSeqaF5a9JcDsSzdwOETFA9wZnE3f
M+c3LQPKrSllknIaEyzYUkifTGz0NxpzAGJccdq5Zf4SzSTrYZEZ0H4xhVnyiH9NlluuC5S5tk8d
5d0SMfWirCPuDy2/kKzcUL4myc5sQZQ+sa/O0/5vLVc7wGCip23GZNCzBtiUdapphNkCk6skwjv6
bautGSEEXxDJ4TZ7vq7VyH2j8kiJ30pplvNpVjuoSoM+1Rgt/NVhtkbxpPyIQE1GzqAPOCjREd7v
yyZizVc4arnwsDfUYwLbjvG4tPuW5lAUsSwfYC+lLz2UDC6nlWHgwhpaQtI8lNoA/TWhUpPmLtax
fNcEH0AnSH2K5STCON2yPA6EMgwbDDag3fd10Uj9wtcx10TR/sr92+Kbp+z6newv/mF7oxKwN9By
uE91T/gbGExCV1STjSLfedez/oWs5aAA03mhNxq1p0rkAGSbewHd4psmdMmuU3mS9inaun+HUNZ6
IAzjyc2+RS13eIRRoQQ3tmkjtS09Oz4O52iQSDO0vZh5wGCRuFoJyuTiUgeXnRg4jGlAS33rm5ac
zuZGyeypvqEhCsLBjI63dFJiJKnbT8S3RSuIe9+Uk0v390EPmeAb4+QvWnk1VEULTSd4/A4wbDsf
xxkIO3RtPvEK43R6JeXVfCq2/MZMnHH/OE8ji6LO54CPuQlIdNtHfRbzzI6W4J5IayA9Xj3PYIiR
eSqLAZDSz7sjcrOFM7Rlte5fWBMKSqfDP8gQZJVfwrh/qLY1l8ZulWR+yxibBGdRBOZO164Zoy0t
seqadaVLt0soJw0GEoDGnT+ik3bYb4nbLGCnBv0Dm1FvfzOw2CJbj5GNOvnpOp1Rjn9p+pfoHz60
wXSeuN1WF7fLFxhTaWSSPuZ4uoZlWVlu0ytnr6vlYUa+MF6V966OkelGHe2J6V+AgVXXMEIKPRqF
l0vyFesjlMWG952/Shxags6VtleUeLBzncFbXzmRWDzrOy1Nj+Q7TNHqPMQHM4MWxEQxLVew6wQs
MGEh4/bUy5P4XZB8YywIN/1bYAkWB+5WQgqYc7aOUH1bcDXC1XwYv6L6zh5OM8ZHVen+zO65RNVG
l81f4NreJIcwULLDxukB6gGpq8Q+/fjFQhzW5V55V4jnhnU/66rhYpNZB0T7YFXiCFj5EeY2y1o0
39WeSBQqtjuoKXRtRs9jpLybA1gZRb9kXCLmxPizbG/GBS0D7DaxQU/DGaW4ykfAKhORLU/rYz7A
GoRGmxa8sd4xobyNHY1rgLAh8eTGBfxKTIlujAEz61ze0tV7hBrCwozC5tytFP0C17MAeb/9STzy
/CqJIykW9+8Lf3UsZ2NW6JIBkE9DOcaKHSHnsa4jdJqK/8HT3rnEADinJ7vdSzV4QjV1eHtQt3q2
dyotKiRwZz9xgl7te3478uCgzFXtb/EBJKq/pDJFWylvZNHFLuAaKf8lzqmk9dWlfO9dbR4qHW6C
MmJF3EiPXZ+Dk0ESoY0NV80DLrYFuxfvrBEdJlq4FOtybQGSrs1hfoe6RYgk/jBtFdqxMp73RHx3
fNcIWu5UpehajBdRNtIpASonnlF57rCq8sL7MBTuYg6PAZYR3IG2gA4qXQ0LiNIkDO61jZz2Dpw2
rDVUjfoRuPk2Qz0GEL1IPfrogKJp7me1IUauQkCMbKSThTgNvG/xOuXXIOtVE6BhYjG5DKOi1WPs
72BYTaucRThQzg5qU1nvJ3CaWC5mXINn7yzLiZv/JJS2xl7TYLZpATn0o1Wr/+Jqrdbgv7LVj0tx
H40pRG8COtfpjiewEj7V5VoZO3nDr1/ojSCiDzgmm7N1y2Y+NZ7umHcLc+l6mztVMPvHH/o3t9RR
1gr2UszljgN3zbFBSgc/1LEkXXo0GSHRUnBM3SRLukKLmdxBu6DRFcs11jq1LxJAT/Jjv/JkITjx
vGTKjvfP4B2/KsJvqjVdNJyOtM96S6YndOUdgB2CT2uE+42/n+2csWvil3AbHXMPGRtbSuJztL5N
m1qnx4u+f8U8gMWxSgMm9Y8zOPY+jHcCVPja4Y0ZURJhLJF+D5E7nFIeZikNr9fZT63ixWogJ/+v
ixwyjYLO83OZMwpUecRitc/lh62hC6MFH1x92VltiA1A2lhR9THfL00XWT/TVIfAqPNJoyfI98iC
3bN6OYcpIc+K6Zf59y6AxoqRsAhIesJ7MEu9KOm6WRHsINztkOQ7UIkhv5c7u00dLhCc2PhmIMrG
zpymDtSEsC/AIgNcEeQMT5f/v/kvvfC5WXiJVW3IQuaoYSRfK+QyVdyF39LciC9/X6ouMJajBFH6
JekzVZN1SbCd522652v2xZJ0r6+HFGhoN8RNFueVNsvPk3+vB2WA872jzGf55ZvZU3cROTKkWJ5V
B2Tw9E+WY/JslvQVxMiYvYNDKKLPcOwWjWnddw5WtR0yxpgSDLa5nkPuQix0PpwWyEiArLlr+tHQ
+P2uN+/RUFvG/yiTwavzkpZZ4rl2aoTI6qSOaIh53GdDyzpj/VXhv1WQwgfdLDy2vPGc30KFf8p5
jm2X23nbmcrP9IjksGH7W/4aT19j5ymsVDsPoo/snklWdwH0HUsej02I69+OBVAn/Yvbu1680wo9
EGB6q6enSfdb41TqIhzgCfA8TukKJZWM77GGzVVf5kzaxCzSSdsMrda9wNZ8OttnnreMr7b5/dg+
pX8Vui39lyVu5uW86XBTmmhkyR33RbzVEu1t7qBLxplDQJFpWEQVxk7uJMtTHIi5Z28b2YRVAJFg
R5NjRHkdXyxDzTy5VRR5nHSttL9nye6j2BQ7vUX3GCTQyZDGwPFSDrlAXGqLfpEFwCA3k25BNilE
pfplwYU6Y7Nyp7sGE+3zxv+nqyEhk86Bk8NsRAgknYQlG3TG+XE0+AP4ZSzAxK4M46mTvuAOshBP
UrejYallCQcpNJnqMgz5oOas8UdM/Rvtq/VRiayJ+mei15xTGet6ggGuGZtpAVVEGZtxYPPVJRWx
QHhNnt6E8b8PXCIkbA1uZadyeBnGJD984YtgkkF5x2QjRzsNfDjF+7fQ6AbfgmgAI8Yw8AMhuTr3
QTmTc+KO3Qi5lMxH3PRaqQwvaHWYMQytxfl4UP+8xgV1VxiOv6umB1O1sDHPafXWZngaz3M9EG5Y
l5m9bQq/b1PUnzDNVeiNZLPAMvhtsckJzUCnEshJn/7D1N+2UyjAWIZt/ithepD06SbHdWmPf9bD
8zTp1RS4Z8hzmL3ZRU9WOuuzqXn/yVeGXn7KPTdqSVV5uoKsxAQzNbvujiIftFQO91PCQYygtHW6
17Qrwpxs8DsApXHYpSvKdy/bA1v7JQSNnQmGjzNrG6WWLXxOKe++dMv1qa+UPwz8HbN82AwzOph9
JejCbISwT1MMC4ncfo916nSL6+ZwQrAY0rOC4rwL5sXHZAE+tj7Jy4jje9yjN2U8iTlaS56UhGsB
Cy3a/ACkf1c6wO0SDIVbCAlS7M6uyku1yPCKKQfRPwifr3TGTK4N2SNrUTfCLDrjMW9reZMPbOx+
J1GWUVlIXd0ucZMd7BHKA5fEQbivVxJmB4J9F5ZJ8CYqeJcDluyRMTZ8ZaTFR/Y3L/sinsMwWag7
CIqg84J2D4FR0LY3sxe0W40ia6//Bq9KwL7pFjqaL/tnYFFXKm0l2y1oEhcILpwHId3F1NmMecYA
fEfxQko5gm/0aOBSDyPxatp/TUkUoZRHoFV/lvD7qK/Vojalbf7AXwVu1VZ3emq9DjqH4gJcIOUx
MZjzoHS7Fi7fxAN7GF3m1pJX0vieMuK8svCHD6T44q/VpnpigwXJdAVYiuBtwosRz23KStGqR/Oe
eZTC+6GuiYrI/wQQh+jwASNgZJj7O4qH8ufXnAp2n00Zn9/sJhD9B7YM55OoXvmQhzA/FOUbqrvy
oTyCFBbqmyh5rU8ebJtykutjoVhRysPKSvNydoK0IxYeHvLQeoap1bP6zS24kUyPKnN92VC6apJc
rZXzjTu7E3INELvSvMXTr00P7DkNsXhMqlZlQ6S7KLKD/NdQ3m/KKuR1JV3LH1w+cMg7uKrxBpCw
FHVB5F8Jxf7/6YoPvbupXeEzdmLiq9haiHkBWKdD/q+TS7bB6xYGBii3gDrg3U8gjAX583l3BI9P
zs1DKVRyft5bOPYuQZE8D6Sl0wQQc86O58wn41mOG5uf696v/LScF2NoaA5ZutGpnFPpCu4fWpDv
LDiEn3K0gCEUueKHTIj2nqaXTWUFhymPKPAnop/cGLnm2KD9vGZQz7gIJpStXPiWEoCDBrgooWk2
/V2hsZ1anOowNq/1LlOafqvw6g0QbAo0nao9Ig2zYMUSW4kcuyp5TsX+YVdZ2YUDI/x9ygjlzz6P
KjIi2fUKstJmJsdMNFk6r0SOqyLujc3h76MFvoDo8cllyCUQyHdrUfeK9+gD3lhZ4lqKFdqb3mbC
yalOtNLRPggi6HLtSRRTBg8AHUlcmImCbkU5l9iMBAKg4Pe7KfEtbQXmpV7T7w7b+3KRw5a13V1x
G7YTL0amdeohTS+WY5KnuI4RWPdp6QwWVusr2W14CYbA/nMMLmc53e79uEOLn4RUf26hzxN558wO
zcpi++IN3WASAnM+GSKaVJQTD2Z/i8wLWx4pUjAyeZbpTKQ3m9TLLXXN10S12Kx+FGXk2293Tlqq
ko9eP5BvtBn8eCjFy1sPoeyW7SxSmXfvyyfnL/DkBQYQjPKK4jC9yF8I3GuNTusO716YYN1CR56u
5fLxQdgolLdK+JaTPUM8AHdnsUdum0/iZ4sZLSRboj5rycdug0gV7CDjc2MLB8zLkhGwpdfQ5icW
4C/adZw4rIO5BnomOCJGgPKaM8qpi/bwYqeHD/4UxDL5f1RpM/TrdXQhBodr+dDBweYhxFADXJr4
XJVBeuKF0zJGMVLCZUgomhWD8nKshNSThbDr19UA5fXYUdHJa8AlxQYoQH976XRx1Yrm2GYb/+J6
infzwR0zBhQY6JIHKp5sP0LLip9rwoEof/zGZMwafilr/1LWZgq2rRv5EnVXJk+7T2U3XMgJ+cf/
HUFuTwgk5wnqiPGac1NpT9rwS6zQeerjoCBfmbT3YLmdGxURjGD+LqCo1yPkk6ZUc4OZjf2+l9am
VHVWvq9YWy3o3rMNzlRaJBOCyOF1o9Kijiz/SEtO16kNAoVDC1SbG5/781xbt4kmLf2HM4aR+G3N
z8lwjSGDfPgidYAd0HJI1pTgN0OrluLmlO9b4+07gR0uN45dhwckE6McJDNwDNQB1eANVUXn/e0P
JeNoSl7ilHe/ko8mDtmFbzk3DXt8MLAg21Yr0Xz6OVg+gNHsIilxsPTZf4K/SyIyXfzAfl6R43XL
aJPyW4eZNd3lpH1Sjot6qW1/ftYF7S5v8BLZTfLnaciqTnRniKHJtZSzwOn90+f8+mdY2FdOzzmx
rfPRq1Re0Qj98YhHnwC0FKa7qmOwM5AKnm3vW2sMoL6Ar3Q8V0MsyUvakqfqB4pcxcffnXl9k244
f1nLfQX1rdZWIaVpvK0nfdWEPRL6vDzbMXaVxaJCzbmm8q+zi0eizYcFAerR7/TAAH6Y8EYc1uxN
xI7IXe4+eEOlb6+6Lf7GRgSqm6pvad5smvXILsb+c205jWPAFSRb6O2afpTAS67wjb3tg+GF/z+o
I2rMobmA7cjuvdgWAJ6g2YRIMikGzUqVI4PZQ5wVvLEk3gL0aFFRj+/grzBK6TihSkK5byVRHWo3
3tBvHzTcL8jYOFZWI8F63Dd3pwkT2W6pzRh8MlmAlvXdZp9pT9DoYoIAiCslGpDccxByNkfMegn1
Hz87vfDOoevmwIHrh2/svyUmm/U8bXtuhxxUoTf0KMvw+3m07ETs0a5wa3iEGh/bnaa9p15rbcKO
8Ivzal/amudo7kupEOQjUyxg26MSnlQcHm1I80LR1ncZ0wTAvLLmRJ3XvkUYGjoUeCKlHO6S/72f
6YJZa+HM+fg0cF1b3WqesS9D6XpMEeICQHV+nx6zSSQUrp/r7JyTFsgTVCWeoluU3frYn9s3Un7S
pQ/u8Cd2uFi5pK27BaBTaQL2mEB+bV5DjhDRuAb4hxn4bRio7B5df46v/Dkyay3kFJe2FP5Ev5kU
MedrJmB41eHClqluAskt0OnAXDqWTpqNivh9dzTplSS7LDPeLxaMMgPdKS9vbsgL3COwN9zTupsD
/JdG8ku7FHMtIn9O3YtH/HmUHQU01zcgnhWf4CmyDt1AvbHpKIyv8CbmBWEkOVxTr7kULyjFDoez
HVEvdTB8wHLaX4oPS0Sn7TN9bwcuyvLhZ9PxdrTO8zyWL917uM8syjH6Q97fGrDRYq0qhma9E4mZ
Lclq9era0Yw1RnlqQW+5TGtS40PUwGSY78+57AhJCG58Lzglq7csNkpSsn/UdL3pUcZy/sHFg5nm
xfds2A7Y7UNQzdvzPDz3qHOdu4ayl1W8wnDc9fR0ggmh2fFRmB1wBySxOwED6bnO1Xi1lu/ZpNTj
1KWmLxlRATH9p2X8tXlrFX9LaGqleJx2qXGQxvmy242U+gsFITbSEBVaMOg/56QLIv1dlvlYkOP5
G+PhCUaXnY0HDtXD4kOKSetIDu2s5U0Wp3R7iv3zwVCcWtcpXC/9Eg2IR0N8ND97ZdGRf26i67F1
+3lx1GD2giEqrYi1r8KoQkNYOtMQJ4Cqi6SlFbScsyFOey/0ZqrMiH9J2J1UfWv6LwpWJQ3Yqzvl
d1R1CDE4z3Ci1LH5KLSiDARI33KRpS51FsnQk+HyDspJNajKmRZAGsYlQM2EIQ+PzSDPQlcGbo/p
1kWbThDi2v7VdI+Zguf/dcOJkOAAbkF9EFIIkfKmKXUY6VZQVgBHYmCKt1esN2DMiqYhN+ltw4tZ
XSBUzvB+960I7FSaTo8gKTu1OQt/kQiddUNw54ztrHyN4/eYvNzSyxWlA615XSNqyGeK9AIlCVEj
vP1c1fBvV+/iQENY90qkI4wCfLtaNYJB06iqs8pMZDFI8XcHbKJWUkQVY23/kFYJEclcAeSH4ai4
V4TvgDhqOhj8dHmNUfXYZ6PWHhKaW6F06m/3mTKRDlKO8uaZXXXqIkVJ8NpO6dQS1sHRvvSOum0Q
Gw9h3z3TePB0oNcmHAkns1gZBzSZojsq3Xp7MdCkescou7yvCcz7oJBPYFgzV//1AGcr5sOEMqmE
IgEbvXMJ4t7mobzY4KEH4Im78oDiOKKC9BFC9vxZ+PS4LXwkezvw4smrIFv6oLXJDb9SMiac5R0x
ShT1ZPXvsSfxCHp0CK+sfhe7DzYHPKLJSea9iIDVYT39WreVi4b98Q1OPYAnGGtLqMRnvTa4VWB3
PS2+7BZ6scsDprWmJgsxycjdDnoHuITN7LMCZMrcij6MHX1lDcPdmOfIjhi1c/UTfysPPdf2GVAv
dUOwLZOMl+rEu3L/lrvQPPBEiHf8thjiKqN5df+JUKF9f9grpMqPNfD94H7/EO9+9rGO/X4KNKu/
0kqJXCdR/raj8xdgybJurb+FI6lt3UOOgwC6RwhxfH83X4TDP5T8EkIuabhvA1J4YblZmBcPz83P
DtHgFm72u1e8/0HWxMmbiABTISRzFCftNM89TKA2GJxyKSCPyQdogWx38Wns9kcPont5V600ooDn
bsrjOfFQdwGQmpK9LmjJ6ikiHov3yFHscDsfdWKUfImCCLdsvtHyIWSVOIXNGyEDHst6zTomkEaq
z4P9uKpVbstht9CUkOmB0d5rplOS1E09hDkS0OPjU8THT/8DR62drZEcGpsnx9DXtgMnIl2dmJp1
dynvBDbjmGVPUaBFGaOmYHfewgdFLR1tuuToZBJGPOE5Hbem0ar4FO2wMGgR1YdLBMTdFPuXWEVs
AA9PMR8pHxGsJDPmYLDjER7dN5MZeTgNWoBq2Q1Ynzzqj7HaheAZZoA1FBC/wU5cq2gB+adfh+8x
apcl5LO4CRGLcP4ZbrFRGGW4waMQzwmDUS2JyA4HfFxrmZ3tCoJKoB4GanVAHbjH0NV9SMozkzxc
XWd4vSqUFEon4iR3KathM9aDEPTS9Vx5Qj6apH4wtfCO0+/E7DZXkwgC01SuGUFWnFOoS1ls+yLD
z1EGc0jAqYLsgSdwwGZcFjTUE0oH1rOEwoN0NLl8Aga3A645292JhFj/Eez6WWpO8FJzmup+k4Z8
PZkcrIywl501hQwam+G1D0zz3lv653ykRgJL6BrU3xUmVDoEZzU/+wqEGnhpj7C5T6V4K3vwjsky
SzFxKzd9vS3mu23e7kVwYQGS2xSkIPv0L8XLVYQ6461IqLs7lxTU/yNDq/o3AhFc7mcJzglgr25I
cw66ospFIdJYv8F5XCdUziKjLK2NGb8rKBV/C0tOETn4GC1xIL+VqyhqhZJ14lV4JiLzzxm79yZE
izepTOqo0FFI3lnyi6N/HuUr4X36lSWy1VbnFJ2UWiLVBRb2mbLkjOoV5qJNseHKU87XT8Dhjm2c
0xiNN2u3LnFPXAcMxVPCZxOfyORGSC3MxwIY+hy+I3RpuacBf76OeoZbTOodUzpkB9vYpfuCUiw5
mu0bIWi8B9JEJyuMPqWMNVZ00o9+Pz9V6kPxj6+gVJ9FzRQ3nUECvXVFxaUPqUIs5m2yD7BeBQu2
nOVS9EkkLx18OrOZzrCW5aMRDkVy/QCbwFYjM9OtIQIZsNFjsQhjBpbflRvuirH1df87+jmRxLYr
1xgDPir9olF0ouB1OrA/viRWjpmPA0wdhEQISgnOEj938gWmEUQXP9AiJO2CMZteOaEb19Ghd8Nv
zAkCPQdhDnW0PtMxv14Ln2MzA/hcsoXWeA4+48kNeR8zLAXs6+bc5e5cIX0mXISVqkCbwyjIdsY0
TjodBehcZM/hD/te4UUVVomoQcWJn/ikDoQVi0j1xXmgEVLPI3G9i/ATBObE8Y0xn9jadlO0Lo3g
tY9Epzd38apB7AiBrrdxavDoM/gzMnY9STVGcacOoDYSmI6XIGToHTbOUPK/5gcfxnOoP6OgSRsf
FtNXlF9XliDLmU/ANg+Z0NzypXzFE4tLC9vFlk7vox4TxDgADNi2S2MFOhTJAbEr7/ZTwwx3N0pk
jhezTrFaXARwcrMYBdXpOtD7LozFK7BrE/phACZXcP7yv0NiCCiwl9QMIwVKFE1aAGcydLhjRU5w
ii/nWgIqba5Xnei+P0WGNxQf0VjPuiM6XZ4oT0CXe2tKeDHNnnsYVhhwIuixexMvyrm00GwaNmio
7BwPT7WZeN/smWC8qygeppRdHQkx95AGnRLKIUfzinmRkarmpHvICXSFIWb3Khp0mEjHTm3Whk2U
imfqzmyAzBDqyAuimI9J7Mxn94PTWDgzTGkW+enslTEynMSzj83c0++FkpDV1RIogSBkVSdcSaIC
26K5c/2nGMPRQyLd0Bfax4bjrexQUlGfldOaVwgzUo9+0XBT8cEykjlnEXYMWJmoin6WumTxJDf0
o8fmZQpjLcXxo/RSFZMLdr7RvI4zeffMP11Ymhw50aGDY5aieacl9r47mZeYnr/gvowRrFDIzmBd
K7XAi0uVb6lCQMy7TCqDAZ9mw130Fk4dTN/DHI8IbiqCi9ozgvFXcPgS4MM6ICWQ2x29A6sU64iE
837SzDZiXVE+rDqwC3PXlaUzTrLyGP9AcWbd4woRFr2ggVILbtDGIJiNHOLfIHQCyQGx1pL7r4v6
grAkx2akC6XHAAGhCBMONPtp0+lwNmwmIbwSwbVQWZ3tKVQodGqDUNuofejsT/Eqbsn/GdjaV18b
gJeImmm/6qxGcw7KBvTderU0vb819DWSnuAD9aalfWIOIfBAyIG3i/WdsVwuOnG9wicN3/uw36wC
lNtkwbawrtj3IajBtijYfZ3Zqlx47/37vogV7P39KigL5UKJFm63lYQIFDDM3LCTTCq/W2zRGdq0
xfLu7IoSPXSxyVlEkdfxAc75X180xKVBGb5706FZ3bp5dPQ6NMOANrEp1KvX6HMh/PVjtNUMxLiM
tS7ZwxCft3mxFDB0ETXEJNVpN4oY47OK5dm/ReYVcCSY1pR966ZpI2JuGyUfhCqPp1YuHsuodJ2R
OWt7GzGTx0X0X7fO/3yiErqiNdLRWdkol59xY+bf7UZzz6/jljKGxRkk/8fdVV0jiDTFNFMkfcqt
m20GNxkf6w+JBEyhf7fzjWKgnmM96Tzl3IepmFZFkRInbWBUJSs7iGHbc3+eBZjcnSqqyY5YgXnN
X4Bve1Q4nipQXFbrgQi+4Ko4QR997MjMIxQbOxTX0wX5uYKodwkxdD457Hpwn80pznc8QvBJnFH7
wWcKjIR9C/UPBlIML0NkKtVYLfEsD0o7isRnDu5GUKKgc/azCPH5iEKl0fu8JsemJxkFaxxCYD/z
H/OWltPJe3HdRtyqq+ZPb3fCGOs9QlW3A7hteQXjmf+WTNZxug71awpDfyotiYnApajUFQaFIUjX
IUk37Hg9gGOwvTER6dfmKlE8MNekMPsXBILe48gX76imBIiNFhpX3hWbmHpVYJZLqXawrPNDAjXa
Dr5qft00hzA+pChc3HYgK3tElTCPg8APiOV13dRih6gsDDH8UnYPuskvxhvabZhplbtUtjPF817Q
brHkRJtNKX3swDb2ZXz4RLRchhuXO7PwcEvgtx5ZLCBWttuCOlmkoN6/L4JEitFfu5mLlbUm4bDx
BbecHr88vKEPdrgnSsqyNg21zL2zF4pNRkEiaVre+YH3DaIPb0goxTI1oNPEAUJ0uzaciFOaDf3u
ae1YbOM37D/4A/Gb5lJqQUoQ1TIBlxagrPV58jZuxeIrX+gTsdGfYcG/YAp2zDNbD0Hi0wzdEr25
WfqW3EDO1Y+THMX5+TvX8uHZz7Lt/SlKIYzTnRA9zaf4jyzBGWSdvu6Kddvxsvf6XSEq27ylzedb
rb1ZuT/xnUwV21lE6DauJlvJwKQhcWXM2DJdsZPFwm2ZhbHLgibg18wj9s9ToVTdBsLzTsTZb4Iv
dkqqyR7MLtNDBhwVzBezC2U2pDBYTCcZeecrENKPbKv3tBw/piSlJCTR+9QpJIOCH8dj4Vx1KXLe
LyliXaemxjy3T1eCdrj3JQ6ED3ub1F2StMqcrEV9XGzt3i8G1o5fd1dbM8nuNqMdXoyY+dlDU+TA
WcwTypwroMi59PepeSTUvh1CmdJpe4R6ud4XjeFX+cgjS6WWA7pmRz6H2JwzxpGknnHBCNp/YlAs
eRGMCA+q0s3G03uxYkk/MRdvBUa4qQLX53r2RUN5Sd5y/DtObkb5YIP56LhYgT6eQUUg4v+Zyvnm
q3m6ZAFIgxNPn0s+uCCeHQ4uPI92f1bctsqmICgtBxC2DZN5hsFXHpYCvPL8vmZq5ATHc1BKDYp7
j/V8IEaA6sBRUveASEMHh0QcVA2+gklfU2E1DcEm/XbHr7nvyS4aushH5pUrpwrEpC1/qS3QKFlx
C7RUzNRpfw8Piq1yLxNTWLiCSGjYRSGGcsUk/iwRgmwv92zbdbPQtSOpNMGLaiGG/ecLYngBptdx
ZTsBUpGpPNYQ9I39OSriABrbFYbExSF30oIVpOkUrKs3xCu1I7aIW/53zyd53qKM9TWJfRuaeCr9
9/B/3jZj8pCxLkA7nJLsq7dYaCS5uHn6/vPYyqvXQRQOVzEsOAIeokr+DdvJIYpYkShgA8f0qvZr
zcX7QcylEFc2vHxJdO4IdHY5X2qiJbpBshZMRe142O29UH84yebowRjVc5is+DpKV4IZydeIxkCS
9Sy+vLp7YH7IFAPDw9A0+YafToTibEDpJRlWFWCHc0YZHnIIV//HYKgowVuRHFMaVuLRTLLoTVsT
t05AgOQ3+LH8SWiGDE1garYYzmfpGtkS3xHz2/nhE1vRUsuAApr4/Au4eRKX4IeVbDIbdP3pwv+V
yQteCSWSJhvWrtFdLhkiutsYDQY8+15/F3swpX6dX3glkyKWoOAL1BH1zS+idhUttbJf1/77BmpO
DI8KITJ7VQpI7HlvCBDswg5XM1cEPb68vX2t0Z7w12ORCudxwjKhuYDAmpKM+jDx5hLVl3r1F2DQ
PMc73so8Ma+RbC9GVXW+SkEbV5Hq8BRuotSEkcz1Nxfc//DFuKfJ4Kbb8YUQahT+17Mmm3/EFjgz
LFikDOn0nko+a0Eklm+NA/DNaNjYI/TOad1nuMOJqvU1mysH5sStIxqAQhsVLJPKn92PpzV5i2yc
uvb4/F4QxgL+hS9VoxDT0J1it8e9g8xXtZ3I8LoxULjMvEkprLi++waHqSpwZrB+3mrzgHV1/sAJ
pphS5uyE85taOy1fFEFwB28VRwn1HKr39hWPMRmO9fPwsDh2QIMTP8o7cCF7mQeGzT/blrubHubS
0dCAdW9WSENvWz3rr8ivcHGaMnOhMx1rgy6Z3baZe7iTvx/qXKmLJM3pJmj82w+lx9n3WxevjxX0
CjUIa3Wtfh0dktCazKH9OlNrtKhE2fNYf5f4NcHkf2McWzz7FMpWOx2CdzPc98rmiKDgNMyQeGDd
jhqPEEigFRLC1Hymj7rtbGabIO49bS95/eOcxaHiFnTlAPdvS/xIRDcOZGgheHKAOLeGiIZxNn2K
1RCiZ5JnIo2r9mNDB7qn932c3/5lWMifDz1rm+TbtjVZj+uLQc3+sdref1/Vy/8vFP/Lr8c9MdtD
qjeY5MW340VRfUGu7vsopXNIus2cXqTC6SDVNqmFqr0s3JFa587JG7aTb8v1kVsR/cbfju8OqjJ3
qQ6N8w8OchuokNlV+vyCJ1qpgXq5tSCqhrAU0Wd1akMIm0l///uyKeWYzKDcNPceaVnMQ91UFgio
dfsLoV1PWDYPiiyZq8dqKMpi+SaTbt9Lu6Q5b04yzO6Hc6bKgYyzJgQQAb+WzqEswtOgcQbIRP7S
CdJo18X/wRZICVxj5zfo+/V+bhsOuqduPO41rRLTseX1gZmluwTi6MaDsiviwO7jGa5/lYNYHkPx
PhnZBIXsTv0UgbU4+Wl6JYUDccj8f3l9iOyM3I+ui4pZSzOhpq/Ln9E3XGJAXdPmcDqBzQgPs0kg
4ssxbZi9Md7JNUC/joTCbdBS/2ikg3EnMNAJ1mg94IGUnwyW9Ve/Bqvm/88luYi8x5uZC3Qqln/I
iQIOKbMpUyYMp0vWulT3A2wVCjGduxroMp1yIB5lj2wnG8MmNVSeRsI8f+xvW4RlQocAC58XxGra
cJYULe30emS4THLNvhG9EVaVF6Cs6mtSm8RoyPBMMiTxnM7N4cxdwj0SVipC4x/GZ70oIdjDStf/
2VH4LoQBVNhIJm8uZ9eILjc3TEZ3hxOn2j5E/xkTWy1epk7yLlMh9PdGpoVxYRPNEZjKRtw2Mvw3
H/cwZC+w49fGn9m8soGSNBL3ULnTAGxKw467oe2PhaGC3fol15CQEwg22SaULBI2DB2MuyocPix0
A2A1lcmW1vq55Lc4s7mtm4omx5zi4UGLeoHmuDyNQp6OAW1IflotOf46oYnLA/pxgCeOZVwdYMjI
gAhCJy6untPMJP6WvmuBKpYe+91kTwFi6vws9Xa6WrOgiYaKmDrBEX3zKjF/IitNQVX1dL2v5VqY
QOb4jBbGHTbHp/qvRLP4U0M9b+SIHR1LDL7PZDM0L6THfHEwrKJNN2vJj+Ths5NSP/S3/aUKR5Lg
sIyoBVnXtfr5Hy0ESfIb2nokVyVB8zU1m8EonTIx3RdSYAFnhua4YTHSLSyppp4G7urfUbwg7/ic
DzwhlYeRWHGXqv34S24nFBLgOrg1iEC5Ex9/OjHPF68Lgx8EJLnKZ84lz69NSooQee2NTTOLZFLI
cLjVBbP8/3ohKQNfSO+R1TM8mUN8tVAIPSLjIZaJ+UCO9fx0RToRzsZXSyf5dmFrqTmg0sKqUUWp
yAwgqDoz1M5fb3GbX4D/VhfI3ypMHOotzLo/hpjHpI15MD6LUjNRQXzZUOrlWw38WPuJCkxPoQyv
VoRebB5R4YAIOcr7PMvDA+EnXRueWDuQFiH5z4nZBbNqk5zPC8/ccuuBnCk+kRzRYgv0H7R9HEPz
D4A8HjnGp+zS2v2Py1ifj41++DxAPBibrHtYVbOdaLB7Wd+w6MemDDVYSCiS27HH94prfvBzuv79
kysaOxx2TTy5BGVtZF5gLdU95bdpBg29KpD9hyLKkXmRrojb959IoC7HlUXKPSzZgTYCkHQGcLR2
9roJzHOnUd37mGLhM4MQkihlRsySpqPJxLOph+2bB29lo76cbLXT/m513pc61/viPUuOMu2T1NDp
gBvCwnRT0tJ0Dqt8tq63NGw8dw+7IHmNIZE+IbrJNst1mCqZdCMlLl/R9Z/LhOAZGnkqn+RK3Qvf
GgyXbTfRLZVHpLgOpOx32n7k5hYznsgI5ZmfA1akIzYogER3Csl2wC2wFhGq2vf6ICN1VzMwPZZN
I0lwKKg/YH0HMARpHEU1uBbd9R2e1QcNuqGDQdahdrgD4t3foPNVvbbmhhOEps+Zy9G8d4Zs045z
IzrYfjc+rCHimEysg8A8h0GwXk2MMkphBmSKaBNpg8TStp0yKcnFvzDxLdwYDDR7Q2+W76Pcn0eB
91E2u9aG3XuvW1Qy0y0U36MvEIknO+6kVjb2BXqeQT1+kxPajsDPRHQw1lp6Z5+9GRYmEK1fO3WK
pCM601uQXfjUlEEnKuwALWLys0f2i4ODsGssOAAF6N2rRgCKMCOt3tCZDevyMGyOFoA0w5LFuQez
pisuQOweEV8lbVLF26y/1INktxQ5vPOFbGGFbvIKR2dJ1J0ZIFguzvi8ghws2zYBg6Ldy1so4+st
FZOM1fwwg4gLcHzY1IWvVa9G5+tf5F6grcZdL9LnqfpR4bo3/hXDbvaz2n30MnVS3OmugEpG+JTW
BvIppeVHLA/gP+CMgxaeZZ4TeHn4KNak/0Wmt1lSf4Mm07VOl+jlliIUnsIlszxLUw+wq55GEPEd
lOK6Xv2MBkV3lhS+BtBQ2UATmeF68wLzvBIONYppLNLZw0iu0yM3bPzxlINUX59HsDFThnKRMY4y
ditNxSQrt3OOhPrU4m6hB8Kx2xkDOgPdB8dyZVo/v0Lwt/wGMS3mp+6ksSujzL1k/7q8PqsWHFCD
pue/KOcpTMHuE4I34CTSuVrkg/Kf0xyqKN+lNDpwmIlOuQCzFyT3iAbgl5OxMAg+gR2oLOwRK54C
DKdZfo12+rizjO8OKCShkd0dBHAfL8Y2R+JGGB2AhnGc1fyWwEjU3Vbs1A+1sa0jcMNII8JEJcgc
GpKYnn3cUbVRy7HHyN332O8kTsNEstwAN87Lg5Hc02u6J4KK8z6Q/S00plmGAZKKMcpYjUBlBQA/
uiAg+u1bVtvDuXWgm+coVZE8/KwSpLd/xB1pmTrSLpL4ROACJCcOdZ4XLnj8Ble7dNcq8ib2o11z
/LqpgHm7y8i8fgA5vo9qh6XmIMV7qobX4MlwRb77Z+ErZ/TBVK/2ey8LvHC0KN8VypH229H9KAjg
wf8oqHnQJXREyiKAhTiu77eXZ6GUeienP+2hC7HkNb8hvgk69wG+XKox/WqZbWyD9xrlc9HhVxO6
5DzCxY1sJBH4fztEhiCRGjtZBv7ZUIf+yumAvi7MyhCosu+9Dk/2Fc3xVCM7F6Jef1Et4z//vj91
jltsL7gTDdvNrLonx0ncQMJjQhtJxYuvGEjFjBueFJVeEvpFfkT1H1rA+rd1GKB/XGuUNuUxmD28
RITVolmNfHTses5ZNzpeKsaeZk4IethOLGEo272FvwFkOFbeXPquCjw/p/vvrvvjqOPY3GXlx4so
7gHS/rtcQEMNI+qwQRI3RBUheJTc00vgt2SSoTLF91LuOZvj5PdKebMPYBi1NWs11Abv9ufRaNMq
KkIDAimb2VbvRxHsyTjl1SgxvK/6UA5z4ZiM9tpDfL/5TFsAUFLpzLEGdwOsvY45KxD4dPM3Eh60
/zJaHkhf3UfpnXRIooWOSlgPFChg1jIyz6OypiPOj6/+nJ2lVxVZKzDeLRuIznoiZsljb6ulTPj2
kdECs8U4It1gNDueZgr1VbqWxv9vNHwHpQs50pZNodNyZt70PimZ/R0UeVBAWjzoFjRgyYugwmrk
Svz4WL0tE8WcmS/JhuJQXmjh5cG8wq+wKjVPLsHH8QhilAm2oNhezQthEMExit28Lz9ib95cIs5o
AvvSQPMXv9FvyzLvS9crh9jF5pzzd1/NcGacwQiMUmL3KMoF1qlD+8iHWhGfVDbgrK2c36q6K9eh
Vn+H5EvSxSZOQNt4SRbdK9EAJs/CWLYcnUG7WfPv+dlpJvzmhs60j8wM4Daabk5g4CK5UEApa35T
V/rKTgaAE69ObO6C+JcRdwVma9Shb9a26RVOI4sI+noQ0BnskMDN5dwxj4Psj2y+OA288YMLiW1v
RIgjqemC1GBHqbvoPc0dOaVsRviSNOMfiIXsfvzo/Kqnm7rkLZeEYW6XAtfIBGTnmcqkshoretAY
yqkszmbamFzMYOSZ9qsTBOUK2OqgCKwZmxtnvVJxBsxSXRnXRWI7t0qTqVMNirhVUyPAJf2Pbf/Z
oSciTMV1kYz4jlvsT4bf4RXy9oXFMWNyPDbGQzkTunnyip94d5+b82AgqBYmFDsHBjqtQrwHa/AY
7cV9aQo2sqdC9jiqwLqY6K09logMCmyXU4pw2zTqxLnIlcpI3p575YYrPszBntTbCHS3GRr62zgj
ii7guCrlPEwdN0WgRgfL//7VrA+3hFVIQB5cSds81Xwzco13RmjjNdcvBjdeH8SnztPtdnV9lt1I
d537Lol1/YS25wAk2iBfy63Utf2h8er8NOyRh8ccgxp1M2VBlOlWNMRNux5EmIkZuBJhcwDL0vzO
IR6t1FFSFsw2dOBKI0HDLphcXIRHtatkhFowkYiRw1ZfO23euJDwE1E6/Qh4792Q/49UwNE6TBcA
1Ze99Disoc5o37xMaSxJhC7Gx/DO2qTd2IaeKIjq6L0Gyhd9HjZutYKyIpHRWEX4uCbxyX4YJ6mC
Ime05FsG+rTJkX94lJb2ETty4X8YG4Xpjb/8fPioZ6FL94a1S3+ALonmTwqNG78K4iJRnR2R7YDW
dEvgdSiirGPLncFVHlNhWI7MARfTIaF/xU872fCED7bnz0/3K8BvhX84G+aTYTz2OYyW/cudoV/Z
ECYdWNOzWpmgO1HmkiEZBbJ2yA01Ivbf2IU2thVM4KvsAIN19izH0IgdoDZTLQdbENhHAKSGaoOM
YLcrJekMNHcQ+eYbdsaQ+uVlbPl/EBEQdT7Nd5BG2poDxP3R8MwAgDaMdqIJxOabK+aqIRoa4H0W
9cjDWHXAi8796wiZ5A3cYtfr2aePhvy2CKgH1s1a1MWTycpFnwOyDzLKVK20XP2qmlbev9il6lhq
1JeNkS9rUU+nIta7pQdQz6Ri2RsKaSiLeU4UPZgMIrql47lnso89HgigxRIywHbOad4b0zdkiUhL
+Qe2urf7DTY75AFFcWyUdpNFU9p0cKHUlDqwQLkQdqWTkWSNvtljPhgoqRgSYCWaOT+Q4jXTnMZK
eIE5nDYpHTs/MVJhAC9JuvoCOehpemcEz5zxdol89fszXacsTDjcrXjlBhsX0KCk111bueZQEPrf
TeJp32sB3ZTM4o9cHY7q7HRqjIow0xpKZ8jCZkTvPfA0NmIb5FzC5YYwbSdI+8GxBv+3JklmAzri
JApHdp12aH7A9DlsiU2gYRKsihhME5DeLeGAqW0qH9lXXixmE6N5OvMRu3f/S+myWo2QJDI/Dbc4
3KI8K0uGVW4DuL7BJpZLkxffduHpWAZKL+T3FkielMFmg+LWA82AdtQcNLcx8bS3btg1up8DlAbQ
RlAt0dZVIVh/VWk6BXc3qbTu8quFRBbbjbKGgtsqUvcXWEYzCZU6Khh+zQ0GdxtZ9Z3cxNXEnMDB
LGFVCNULsFSfGjRVgRT8t5BWhwID+gAl039BHvrhioCtNY6Ons5fzBOfv5bN/41jgtghJ4pq5ki9
5EjBgUkv30OHL6vDZfwH47ydanNEUW8G2+JLpJJQW19TGxsc4KCkR4OW2RA9rJoBuCmvlnA3CEnV
+IYrDNK/bXnaop3adhu3EayLyw7lgtKHr0DrR+hTdM4AAlk3YjiLQs3ZUSjaxCr97ETkCpWZO3MI
i66iyj7DqSCpKA0Y05wGbrh+OqiontqJoZGVoZxjEu01bUi3sJ44ag4kebtUhihdqDX237BmSaw+
D3Z7zf2ZfVg2TEUifBrCxsrvyz1MVOy7m/A1brYUOKNjcI4zjzQQr0fSxCVTyG3VV0XEbDQda9Qa
ZMP3kKflIaYJhkO6JWUDhtDNEv2d3+RzWZiH72VhB208fVbjgEhJDHNgWPF8fAOqH4NZRsg7eqbb
UfwV6W/tBAfhVeyxF28KzJDTty3pPUAqLtfOEg4/6E0JMD1tdh0EpqH95rXpTJqYH745JcIf8AaT
kScv42kZM6mA6TP8BmiWl/rHbHSMo2je3rDkC83LcTaQB6rEoZiTmJWfG4MtgPvuKCDJb8+wOdh7
9x7QF2keyLLm2Q1spgVILS1BxqwgFYVxWIL+nyJiOPFLBZUiYHftvv0XZLq1vJR+yh1QSN3H4jA6
N10Vvbgr0iXiGCu4czD85gjlzIcmy0a3vNrSBsBhENmOeat/os2bDu8YROVmtxQMJXKkGGAg6OZT
5o8rEKG54Mcto9b63mnvgbvxTKrFLh9X75d5fA7UALHsCq9Aw5WZRPtm0ANj2gALldLfvwabgVNv
ASZheY4sE0hnLfyAd7o7gTl0s1geY8Ko+WwAZ/DuthUnI3sxlesxfmog33RJ3MBFrhn+DizTQGOZ
H5TdQV8RYFUTIUN1hfhJSsQqnRmuamgyNdo2v88m11jDTd3e04SKU/RD0CtEFNKJkiluNhys15/N
kH/Cu0GS9j8VVFMyhk8R4DhScjN7kUBfiC8UjWseWBQFymv65epZ0/E37I5xTj8oWaIo0MTproLH
YfDNpe6/lRK1dBJGieemcYR35Yo05frR/Sin67MMYR59g0s3LNbwS5P+vwzikd9wSREUfNhzudaH
VQlcR4Lu2fE55fdbLWllctuTosB8PB126Q6sA9JDgdAPq+3mIJ0OH6tlKNxkg2G77ppmyDBYCzZU
ygJ17i5w1gUnpzChvsUQKuSLBCdXf2MRG//5UKmwNjVdgv3ZAxbVoR4dN9IHdblDvnePB4izQgId
vBnGAmyqGVhLAXbBXMHEyXDNMuvPZpiUwSMBUGJr0m5e3U4nKLdeMo8LUSATCNvp7v8/9QCersUv
tU0fatl9qopsP3asscirfCthy9L0A8hMC52jc7oWe9zGkRSIrJu7h3yJ3hV/SZw36BHpolYUACqk
oyx47sn1AgSAx1YAP0rhKViwH/uX5z9xfDYwLLwW/tKMDRsLah34VqarCjjLPwhvbcGz9kEaoSXw
nC0OkzJAXAhbCPa64OqUrxH4DyB0wxo4OIWm1LTFIKpCdWewBLaButiUfCdExQwEKsrv8BSXkO8v
l1txpUViQLANI/nrtJ78g0OuD9QusqUSHR+iiKeZpwg7QJaPomIVfarnf3usZulzY6HV+SU5YB8i
8miUFLoK9Yp1HgoR7hFYV8zJKvf3yNUc7QpBk21zmojaJ083wCiXJuiUqEwu0BRB+cx4JAFfBs8U
fyXdbGezmRxdVqFjNDqpiKIMc5caW0T/e5LhyfbTbzzBgaX1mhaeGzFDPAWcnCGZUEUXHQ5glEF4
tFUOsN2wNeEZUQbE1p7NPrl/ab6a/U+DNoZvz4ZV7Xhq9I3qQesxenZmkDzIvYlBa1xWJEPQTQfO
aW1yhvLYZyYPlXFXEI/pEAXx7RhWEMidqP2Pmu1SIypna3yQnoYOFz3PI/juJ6bUGrvNlRxtnWah
4yft1lN3HTOLNmlrqLex4SPyomuw4K1tqZyVS65BlbePfPttKk+O5Kk1DhPEcIx3d2/daXUsu+ml
C0CRBLVpXHMqEUSwBWF940F5lnioxU4HghCo/4BPiE3cTjoV1z0qI+vZPtI3djqh7R0JsB1s4Ll7
U5cyfj1/1qtagwbnsSsyjPjhI3YWTAOQ1bKrPU8fVQZejBwH4Kh3yebKHvzXz7ZMWfnu0EdlFcCA
cknwrE62aRrYYhiX0TWpXWdNBfCZFVYnxhsVC8SWi313zvmgiIFyXPznO6zwHQeC5NcQ5dzNTvWL
t0RbKdxBSL0XeB80wWKp0qS+huBzXUGtJquOij6tpMrO0jZpItbcYr3iFNrn0H+IGh2V3DhMaJVV
z4Gf5EPccTrdXDlr8DjfXZ6vPCpsypLLKp/Ez/6/4u1T6BJnRqTdAzdy49XxwLTmqjRRDGsnst9g
+XbJZpwqv4v1wpiAKFjoURu/sxVyURNQCSKDFlyRpzdw3Jh0iGtnYTixbFRrTOzQEwohphg5i5KI
buu0liTC12+uzzKejc4O5ZgyAcAfW0LmW3hQR04LWJJZ7RoeyYpvd4e5qxghl3TWrCNXWcFtaRwT
exUfr4Mz4Ob6/O5ZB16Hf0BSJbjBAVg0V7AZlexBTJaWMMR/hgX5LRhYJBjzJGMGGAaM1rniyaZN
NgzU9z1UzuSPcoVtDhCOfovj2lo26UrqhLq7lgiR3R8OltDdgNYpKYktempquCDwjz2Jq4fYrEF5
MUJ/7zb1lbYpyTv+RP7BqdCOqSGQl60lcjehMaFJaD12iqe2ZRJ8qiEa9/HO6H3e6DOhzbRWKmjQ
Vod3KPf3kjwgEiRacxNvRSXdGqPPvOXdxVkvw2/1fopCEKTv6D5OAIFBT9vyO9oEQNFJtU521wO9
SkIicL+B4dkjIsCHLLSKx5dKjtuoMlPyVG7g4QZ5Xufof6ciZMsmHLEIF12iGesyWyKhGda3d7/t
Hlpc+0CjpuOQE5YGzb94ZkjcTVznWFRczc2Avo0YvwtoaxGRAzr7nCP2OyHC7gTQQ/rhtY6aPXN3
a0e9IF8mS2KHp1VFbjWWPP5+Vjc790eL2VvHbKfm9lGsYJ95cAQk5kDDsSXQjwB8lV8goCQIcmQ3
xjYsK3VlJmOEiLg512dY19cdiirnZ3DQPKImMorbGZciuQa1aTzR91D8YgTwSnqFZr2dM4ajjubj
qBJZdtlzOuXCt9UZQk1017kx6drnXt8IxnEATFnEYFZzSwT4xMRmql0uDXNEIw3QOdx6rRx6+Rxc
6nRRZVMlv/EhnKktsZ2DXDgBu7I3XYx56R4YWCmpLNl2P5C5dTe8XGc2NPAocm57ZzVLD0jg0A2G
+6WL/ka75zVwkyr2T9kMd1U0sujQHzLthxx20y/ra1gjujaSTGVDKYmQmJmxdmhiBT+lJYH9rHHc
Z8ilZXkZKosHqnV+XF3Rq9J4GD0JnWXC8F590ykJK7UVMPZ/8n+PDCx1nw5x5mCfCm+Yyot6BB/t
4BpZrqp/3bgvpEu9/aV8Sq6vf4pX79+xmKBh9nFjdckyzjVBqZlqcG8Di7DBkCdbjkA+GvZFpqoJ
snap2VptnXozlWMfK8InaVQWaGfGquTMfaynmCaEbbP/8qU+k17SMCC8j1bF/qfeZQsjJ6zfRi6s
FDO0kNjjtOV4bgaJCwLJbPfVYd0+nhB10hskFVqKAHz5rhNR5A+OCE7z/XbdBAs8BJeequnfwoBb
2MUNTLrXHiDnvtwOZMu3PHVkSN5gDNC1qwoNjQ0cUZL2F0OgqIwEKQ23q1/3dm2X1i97gngoCc5J
jh7knnBS5sml71oa3xmLVJOqa/u3ygX2mIZyORMajX0WP7AgSIIoC0ylWVdnfam4n/n9gxgPWhQ8
A3h1rjugcYKoXdcFFmm85LJUfgULTTckdSk9QjfupdK+7uDSGMKp4lxUlLFap5ODH8Hg3BBNvGED
DiIfvAYdgYO5iE7ZJ2y2YZoeyxVPRVk5aY9VyXkqqMog9aeyHf6HmJaLAnIYzY4Nboe6ivrrn3ES
aECG7iqOF8U59RMIdwD/9Pub773NCSAkCs3aKg/fCogUXQtVloUgc8ZTKA9l4Wo9NSoDu9ukfTKr
KyEbwIL2b1xVCxlVtWiV1BULHn+V0V8BDQMi952ThCfi7zmKcGTrZXPVao/Dy5pCbsPjUwP22igG
ymBPkip1682NDhhOpFnQiczVwLYzcIwZzFPTmqFh/3H2GBd9qUqxkmOtuJO1EXikSOMA1uErRsmU
YPzZpEowsUtlAw58mz7k8v4FIIpQsdmqG0D3zhq9uT48j4ZOZh9foz4V6842RElnT3ZO39eQhZi1
jnI3sXJq4sCy78j7huxuvQg/0fC9ixI7cNNlfH4w33wn8zVKyVzoHmA4xe15YTrzZp0Qnlj+fbe7
bzUq0STPTicrc/mfrXgVbXcR8vHt3dSX0k9+zeikuFjQsWYFqEBfrjOSqgRMNmCHEmwv6/2LALYt
m7cwqyFEAdcPOUbXmFf3cWweZSoSak6Hr/I5K0VpApGe4hyWlGSstroz3Qof/k9fECkMXnIo9d9T
59oUCy+fjSOoRIpRd9iltl4Rn7+z18JN7ZWxWNiha5hbP8sriLtIeuKIMH2Obr8FuE0p0754S1jO
M/4aX8Gi1FRnsF6RHcv2eV3mM5L4/WP9M9OEglht7UwKEYdAHGIkI9yGDAyt6tyXk34kCQ4VYKsO
5IEW1RkaFqucDjPXkWqEkH82xzh4lQyy3sr9cQPJlyvXPEtNgVZe3Xrt7mAfvgPPG5AM4hXGaeLY
bek/pOekqzLWbMsCoc6p7Dw5BJ2PXRyze45tjWE+GDBZDu0NX+i8+HOS7P6GmI90S8svmaDCnNqW
2m3GYKDo+r9XUW3ZB/QRBUX5w+tkCMHb9Amv2+2rkQBJGlBh6S5S13MOz/MSQ9+8IO7SNkvZQLNd
euGO75dAOVadpwkSDSt4oAHxzy2jM3Dr+W6LLTKb+6dQxklh802SRuWM7ds6VjGlJf7l9yGMlPGo
ICy/4th+QizUDcrhXdSLFlAThN73jATzU2VTU4TBswpT5UdUfSAXqTuEoXdZuBSy47e4QqOj3+g3
wZOcP1duSBUDsylHSIlJXuv5LF/ugpeBPVEC48RBALevOpno07wNK5g0zEp1eKtMh2YKlWvAXVD8
DQu65CjkBLm/fKleOvmNMhlyfkgL166oMseLvlxDVbPTRDdPquxSjZvSRRn/xhzyhJK08O86orEH
WtIexUhKnHYrKjEupVanP1lnq3JRbKLEPJU7KBPWOwRzNBpU9MvGxgG/cHlCY8AZTzyP/rhWj0lL
fBrOzW+rbVXUDC/hiHAB0TqgqDXC7YtfvUeOzLz9jaKnUZTDpRvQqBnrwfMzNRrw1BSLHbWPAC0r
/zvhhJj2evTX28ikXUBzP845xb8+FMgSEWFw413HIPvLB0pB+0x5uJlp5MEuoviGXAXlkW6n2j6A
JSlxxeA6rzcOFQCGgHpUA/kqNc6Ca+8QwyufkweW55jnum3gT/2g3f/XXMUzm9PohYG1rjTUOPfl
IK6Qa4SKXS2QRTGNMVip2xe17d3zuJ0lGZSxjHcTTX1sZQGIE6mBYrOxjq0KdvTlvIbKF0Qrsu2K
gjb2UeXsLFqiz6wWkoUktOh7CewofcqhVYKXg3EazYmximETNMkD5B7cuF6Ed7jb+23V6vw1h5bO
KADcRhW3u1AHwWfBcLkTs22Hjq0nS0AhWRWLc6GZ+VwItkTvDX8cl7Djt3A6qzzrVvE7JGvqkG6H
u/5at9GMl7NR+y84j3aq1KEqXfiKuLNFKtIUHWyKPjAvO2e+MewiRp/AnpxjWABsrxs8GkVrZRK/
SG2vzSipGb9gyTvVH2m6PoGhTaUrATUxV+FnhDwrycvk/CYfB7dTeQ/uJI6VEvix5+f3K/HFeDUn
jAK6VfpaR+h8ePsixogiZnP8wAay2kNgCatlhPDH0RSzncermGVPxBgieF+huCBi5EfE+yrCmp8z
IKzXmQRvKYJMbFzLsaJ3rn3jgyPEAFhKu1noAdBJ39l2z2b5gkicUwTJizFTl/dKwStrhN+WTbDP
zjkW2pT5LU4udSfRXV29wdRzv4NZDcaxPg7YBRK9h4/ggoKHfDrkTbO0y8GMoUYBa7Q1Amu6PZzP
8XqtTgKbQBRdg1eTa3CAU8lvbPpDEP0T97Kydn9bEPm4Hjz+BmwxyNtC3p39y22bk7pIGrDnc9uA
Ggxgotw8AuQNlzVCr1PYWnGFnZBLxaXdKqrPBb7EBwH7s9XhoaCPcOfmp+jhimhdEXS/tkv3AZLI
Ne3PXNTxy2BVoYdAbGOTGh4gPVUFgTlGg7l8Z5i626X4dGUb5c+cinNn3+2wezCkhkvWvkRmHint
6hxPCm/QHNuLxuy/SwuNepXa4KPcSDREC8LnD2Q+AoPm90DY/aRRp4arnrq6gelmP1oaY+JsqA4B
9Xpd5qLWSZzcu/iQNrXJzR35ItxKyIhhjl0DkMCfTXL4Ng4q0PBQ5roOEsN0E/RMaMc2prAILWo/
pWEKqiZPvZQ3GGObMxB3Cx2d+eWNs+tTrdpsizTcbr7LBwqdLhgk2TsiUJyhSzvQ7mJe7KZ31+TD
JorSHmdpzdeEGenRWPMELlEJ+bB81AIDVlUxI1hMOS7chOz9VvOcfSlrqb++r6JxrMa/koB2cF9m
sfIkiKwwRHcOqs2t2DPblu1w6CJgmMAB88z/5ZeAHvhN7zI6s6ULeuWYoD/B2ovZOBu5MxmSWDkF
umdY1MHO+uG+PMSZKEDCIkc2OWEPdYHFLBwodctETBe/bQZZ8LRjprPf1q/Y8WEyUIySrFxlgsiO
4o1OkXLM+oaDw83ayBcG0TNlDWARJ2tfvqF+jE+AGteVamvIrBuQ/qEFIexx0+CZnedCYA5GAaa2
LdceKiVoFmPjm1wbofJ/dDCBKay9TudZ2+abOqqsEOHmDv8BgEGwf+wKx+rVxfaQ65fATokvJ4Kf
I8r/6XEUb/8/aa/VyEmXHH99JDwCM8F98pjO3BaJojK4fxrl0t8NLjmbc+SZR5QaFRmV0yLDMLD+
cqCb0BvyAOFuatSK5OsqtYvIeyo1LmsXzk/lkRqcK41zEEVjzC9RwMVAzNpV4GDCcTqjD84p+l0D
zWlgqxxBizQoXE41ycgle7qfF+s40nv/coDzP/otB10Z9vHhzCfVacBrJ3ritaWcMbasaMlM5fXw
fJkkBV+KFXIlRzLlOSP7LtLp/OaWRxfeAn+6U+LQPBpTU3R5ZvFLFFMZ9MkvniWLNi9bk7fzF9bq
rEvDlNboRy8Lqc6WpVXDfGu0XF956PgIZ1Uin9+66xq7i+GgSK5sBuNY/pfT/PdcYfGyw2KO3XpL
BnFJeIyBY0D02rlBNRSP5OCwAXd9k2EF+djstpyZVMJOCR2MKV+d37++/lcfD5bdc4iw915DXiWm
o7UoVE3Jy3h/fACSuC4zy77XN+iRDwbTgWkGp9K3PsburVdejWp1wekuwL+EMc11A5lPGcKyxL9p
YnKEifV11gJ7dGxmSXHaaqyfp3YF1LHEXS1BFF5tMFUlmK8991QQApAZvvL3AgLFZV9uXqTWwMYW
232K/X3iHQQKemwmhS1WqewmniR94KKwYgKfq9wx+nA6D0Rjlzawf/B78UYmom1kij4svz6p/+Ny
My1equ7mtzxSbcCfF1fNZyyTHBcKSxwNUc3tPy5LsRyG91sFqG32ab+AVL4UrR2Y00Y8i6Aj0GpO
E38/VBYEdO3TIbolIEN702cZ4/s3nkMxjuOX6Si1X19HfUWOK2CHwJbH8xEWn7NAf11eCWfBPw+w
mipRu29VVmsTqTzJtQrV1kJ00+HxNcqJAx8KTgVHB7SAmwQq9LDWQXVujiAttP4AC8ns7Vvav/nu
XDQSH8Gd+Bs0sclusK76ta8uCyw+OTz1H0URXZ+pgZNlPvbscA9MioxyIaVp0N0tBVdJ1gaJ144v
dR4EvVY/ouIrLmSzSqQgF/8qz3YFn9NSveKHjAzGPjy8KJZZww78HgE/H02XJW4/CbQel2RaWfAA
d+LlUat2vDL+bacFRhURaKz2P+EgVvfkLXj5U7aUpQMGdAEvb0aXq26NziKxdR2amj3r/odtI4yE
zsHLXJJFUixYqOkwq8LESjDLKo8jNen+pi9gaDxMXdZNxj+BdYV3BIRht2j8NZZbVKHahpgtyDKu
l7tEG5sixwgrLEQkbzG99ctr38e19QEyFHTa7HuOQPr3w9aiZFKtmLrXPQwZlDBwHTQZ2kJEiC8G
AqhsWK+G2za7uXBDc4AzPuJ/KAkWLrXyxuXctS4hajKIk/+KsZZz15QMichzO+Mi6ypugexJ4fT1
TKWa3f2Jm4/VfrasFfCX+DeHo2Y1GtikoF2wUDRcShZJTGGtBlnzaIm9Zc1+Jd5ltezOwZcegTZD
P7mf9MFbhT7jb+zp3/zXCHODkpOODtTahR9akAFwJeVeEtg3oojRObViHaCn3udc+V5sSEa+oIAj
7NEGS+Lvbxl4It86dvq7+4cfheDg7aoRrlvF9nxvilwxSrY23IJu2Xzw8gR4xWjDHvtZF8TRTTiZ
FuaHrQqnAhuX36npxsNjzSaHuaEJBB5m2SdURcDW0HkqlQwmwvDpXN1JMy3FJuTBZKhqWp5dm/vl
eYEJb6rl51GpFLYuk6Y53QCDRf4vhz6xfV7WHa88QCujO3Ud3Ijw1M25e2VO327M7xlqJkHNjDoq
HeEub8Q6plQqSC+mn1SIbhfftAgOiNG/euHC3LTjyDGPE5culGNcZHAqpnlLbXHtC+R9L0SvHbjt
cErr21IeT8naOl06tK4v9z0wH54a2qErHEVNeOaCM+CkhVQk5q3E4A02iwrASuJm2hIxV43nK1jc
ianZ+mRrTo8d842bGcvDDitqc1sGe+pET8nmke/cJs2cM6R2b8iAuNBPeEWXKzFslfXJbXuBp313
XUQhAOEitAXAEe/HhxgnFQbO2QfKKzXj3XIUV34328hNri8aqfkIIi1yfV5mUxEVFcnjo2+mPmCh
jW+0RNEZnBXySx7ywsO2+CLuqOh1Gsz7xySf3Exgs5gC658uCWInEZ4MrB/varwyUfXXs0GOSE5T
LD6vmyKeQIj3B9skcQhq96WsIHnJmeXXmYKv8rKZc/CNBN3cYoW/+J+Pea5gF59kT9emvCUKSDGb
jVRLGWUvgn+pAAXzjay2Lvu2eg+Uk7P5cOroXUvH7z6UJUvJft8BJW8W4k5o40sI716DPYJGeJFW
2hEXZkxVkmfXUz7x0STUFxpYtZDjtYuY4ZhVCNZnXxjfHjnv9bqByx0YZwXetSQFDraYkD0Nl+ea
JTtxyyROeqTfPXvMnW0IeIM9DbGUvHv8odMLNb6cGtkKsRkRcEmCrgjf2o5B+9H4JedqnWDVlvHt
7gISlIsPtTrqgwOe1wE6NTOcoxmt9fOzVn6hJa0/P+jZCqHuk+a79r0FRgqEtN1zodRF++wZ7gMz
kLYx5T2VJm36wCI4U34gx2j+02+wVONiO3sXZJlo36raKJwB13mlk6cZq+hJ1IeTTtbhH/9Nepqk
ck+J/m0Q3v8EVghczUDY0I/CHwhjw/nv3bK9GxYAPjm0gCu/WZBixFILuagH4enOcKKkzjrNB0vG
ptWeRfqHsemacks6gn16J/Qihm84pR3WkXot6FQ2JHLmv9ttt7z9DxH/gkZdyk3xVmvzK7e4eZS7
mlhlUVQPbP8LRHSbWFQzSldX8YeDjzpIFxUSob+1qoRsmOKbiDX3Q6ZLUWW+IQA2rosa4tv/SQms
nHTbLvk+Yinj47MasdD2EvYpd2TwvEMBtU3sNKex/6nG/8lhuQoiOHJ2clOi4Ia/7aDuy3U6NS8X
FUhykdjG1PFNY/8KV0hRk5iEyDG20boBWxTx+lPLOSBLLDF/Q6PVJSzK1V3KAaiX2IKMYaVaa7Jx
vaTx5n0DfpCp3Ih2iYDYcHKA913TUsdEPFhc7kUprxpdRW8R93/iTKMVskhOypJJqYH2QHByEHZa
gfOeStEdD3qtFi1tdHOEkuXXbeD67pO9wyw7Fq+mIKzeeEqGNrjdqcdWj86roEHxRp4w33YKBXNU
4REtwG3seWcaj7CO5ZaHtBnUXOt38GEhoT9aeS/Cs+FiZBLHTpdNYTN7/r8rMcsY7HTLhlkQQNVQ
s76iINVvOXH9nY5mZHHhP9k6t1jGjgSz5Tv6KvCEZwfNjOjdyVwErS/N0CvLAwugNQLDAuudxQi8
vJNNkaLzXF7nJ7TaKnFiEWIdjikIOLZqycBWVxC8W6/hMGzbHIi/wP6FkgNrs2mgGMab5WsiAuI1
JYfH9CatXYBLVBfQN03lxRPFt/VhNOh8XIxifVmW8EMr5qO0fIhLQigqwXYJOZWL1h8bgH0DQH6x
a87GBsbCCneHB0Dl7w41766BAOw77zxNsN+3qHnqmQ/3P6F48rUbu9Hi9BnYVW6H8kWKSlZRrAE1
jShr0pTYRboSZFaHIv6XgSLGCEH2tWoh2s24tMttWCI7TZ/KP+UiOdkUszTnSJ93JZ0uu6bmKGfy
g5bsY6VrO8wWwIOc20o4vnOCFjMacZUp3HFRA3nvlsW0ytHX5wTc+qHaih18v2PG7jsl96M9HDZz
ziTHq5pRi6aVto8CsAxKBGCI1/JnUmoJgcin4Mys4QoksDzNDZ2j8Jt9zIpWdXZGOw10L5OjBBJt
tTLe5Klshse6e/z18qX1aicLWPR46oM/UOxZfWKCyXDgC1vcybXjl4yTwIk9CsoHv3cSoesyVlTl
39iFfvwK/ynG6T0zwbp/Yo7ji4swBGrhfYcUHmeNwROWDKfwlhqrVW90dT1HbDbKWZPZNMzP3gx+
tsWdybp0DUXNqpK+knSjqikWdRm/dMSpZyPGzfPqIZ8mHGglvnGqv9//DQ9q23TZVjRKlfpJ7X2y
0MqVZz/zWu124O1mIaWJjV9+ykBIpLw+n/hArvbF9wk0ApAoFjyUet+Gon+g2s/O92Vsbkke611u
JMcpMyQZ04GXGWBHLFoWSQzcL7AUTR/QhYOU5optXGYcx3yUecQE4S92tDzfoXk6i1SZjQsFa4s2
yVM7HJu8zaoPZSTsuU6ZROZW3FuMkdkGqhKZ6mfXtYLzZobIfu1caxZdLH9JM/SW9itYxxR49voL
MFHHmacASLhMtS6vXm2MP6MTGbs7R+bG+yKE0RklF7piSJ8LODZ2g/tcI4o3qOqcDyf6lHro+J51
UYT8odgTecVGCBB83Psm9u1QgZwKyc5JoyQAnUcEx3hs0iULnyVHjLrE/HozUEQRJcYCkmQfcxOQ
FiioXAdU6ezT9z6CKq4OTV+7ua0SPnECF4Q7OVedfRkaZ1SuCMVJMR6nM46jJOxU9l0jRqlj9C9j
1m65qv9zr5sqbrNgOFQ72+fQVVBlQofU5Bkauwj1qE3YEsB8TFk5b97/bd4Rop1ol0eDObFTRKTr
L2WeLgQFy069PAcjSy2hUPHiW+D5L/mB5FW3cB+QraRuEfy8LcvycbG1qZWQ84cBBW+8ZFzfylNt
crAIvpl1Qo6pMudxPCUhFUdYn2vvY70jtju52VC47PQzWboJ9TI7RaTeCYS/vCaMpEMzOB0YOKOb
U6yA6ssZpssuM3tSUNQkx5Aj23lnFW1kjNLlaJNtxUmD8jyw43B5awby+93kf1hTgLX3g5Q+a/Qg
CdBYuDL4sT6/HQZ+UjE7AJ5lNMQswl2WLcPilJAL8gXNKGd+yEyC44F6Z9Ft9XaGx8G9EqQUmKdA
kb7wEijbx1b55CEe0QDOCYGXF4fNVoZlw3Pl1oZkD561NefQD397HZKDfGhOpK+FGjcTVCOSGi8S
hav8448lalO5zrTatyD0UiOSvae6CFHyj/EW8FZwMtEafwz1zcNwPT/Q0+1PQGR2kzHchqkcgu0x
KbeAq3khzxfsPklm0L7DiHifhswTpQluWj9cZXW8tmZYrep5UIwtcbMgrYzSjXnQ0uT4Py2DkpO0
SK/nbr8h+lweoQjlP03sHzeYzI3GA8fIaRrbZGfts4WPL//2iRgBPsq70EdF8TmoGTodr0fKR2Ss
WtrwMZRVzpz7jkVZZC6saCA9+F5HxzFO7h7h08GF50bVdOus7Gu0VKfdOGyZELQrTlevTI44Cbt3
PN/JWUJn+x278vhRpyTJUsY2DdqBGvYnq6Smwf2F9JAho1WUgjd/hKbF3rUnl1gzBgfr01szjj+s
Ua8ADTqSsr/XXGHeVEIhupnCoco6msr5Q1dOHnkRv8gVDOfnbJ0ZX2gKLIGcqukei1JyQZN1oTU2
+RLI7DMum7YD6sSukxbkKYGUJICx7I/yd/LcC3aGqtX7SiMCcAW2omB8YCAMONf3+91MTd9eQXBf
PzdahFjce+MGVsNIB6+CAJazoDg6clIJe39zn52iiwm/hOlW9LO0SNILu6W1Na91zfI85lqpaPdJ
yvg4xbo+0oNqVSAk7BwlxdiC94sSKttPuN6tAlB9ZYtXkjf6D2PkYHa8XjsgxY1tLUy5EBJnG11i
MgEhebAZ3+dADumLn3jT7LsVYQ5+aZy7b158XVV30q/OuG3ZgbBnKoTJaW5FEuNKBPb6RbkqUOT5
dZ3Rkw9SQUI3jJ6a7FKZniEnhMeKBSuXNReCjcCifec6hppJ+X4D6lxpng+bZzhuZqn4RgUzLlnM
qd1BUcJE0WqocJtlIgkckcENzwCfNB2Ir059Hblylr+2CpwBcPUkZuh+ge1hU5YVSrAtCPMIQh6N
t50DEry8AnexRIPCmBsWIgeRGEBn1npCwOxWUm/cDv3dLdIzqaKYJ/M7dZc0hJMHMLLV7mjbgosR
lAQw8Wb+B+Zp4lN9Q0hZ68dborHH0T/SatSEJd8gkxXHRD6bWjmRxexm6tA5nHgrlw/1Pz63ZoAM
X4y7VXJrzs8BuObKAvEKeQS6E3UJTEdS5CCCvAd5HoygGu5Nk6bcXxQKv0TlMHtNc62NFNK/X8U4
Wskel5i2ibanWycrNAc6gdFBrIdY1R/9mMaJ3mWjgkn2PoLj5FqaxeWKyMUvf7pHShnGFsTHw0Ac
AvuiidB3Q7mbs+qWm7ibgtzRl4bzOn9K22NyGT2DXxRNhM5fHo+R7m0IsWgWyU6ihuqWEMF+4MON
z0TyIx1tO8ez6AAJtavLqwlEFSQWr6mr4C7xrPkaDs4iKyOSMrrCdhmclQYPHzjnaTKE1IJesWRL
LaQk+SOfQVP3tParXXEYvqsG7d5+Mt5W2cS4bBLcTV832tc7j5+PKSEtdXT4lPLA49R+ELt+9tUi
64QFflNjC1VkSLzZ+UEhilXZTLnxJi9nUVnwVMFDZ4Cgqd8mkvAiLWD2Z0xhIc+tIoIwKG/aGMOB
flAlh2SZ6FIkLlhAV8SaW0GbSGGAgnD+zd/wfeBHpYR4fNQqq/13jxtwPlVick9e8pKLOwKqiAHT
G1F4Be/DL/ElX4BOF3uZrbzmlkMuzkZ52DRUG9jV6f8FiQOjGx9nnLscxk/xUbGmiT6MAGWOvSCY
rczQv1UhDDz3m0NuJ6S8yMYm48tVbkzogg+bfZkm/1YIL3bfCR2IyRccgwQyI9MmoaMOyyudHNfw
e+LwLExi5CiCcd5TdwcJEv8Y5qjr/eVoEbi3nnWDrTQBPDduzHIooD5BEBs55xnz1k/edD0t9F/t
NwHYuys0C0dYau/SHYa8NjBibr02qy3qOOXkqsrUa12enOANOeXtTe6W5sb5EjjmzrpMcMJWPuIi
9sjhk6WrzYzyFEpjNfB/EDUvqPhlAAvkigeKtnIbRXIR2yBztnoQe3lsINKn6o6/tGOTcn+/WHB1
6P/07+GdS4KsbiwPUDRAveWmolBcdhLsJp4wDWlu0foVoqdzClZebSgFhbbnCz1oIl4cKgFvj+X3
smAoOP5T3e9sfwRc4qcUM4SllBRvyeSbCQU8XHxgzNtWUAiN0Xj/6GTF2xrzyBPbsbqw4Dg+PI7z
3fsBJABilK+o6Pqj51DBUDLh53U6rWbsvjj6i7bJiWDR+04fZT/S5m9LCkgMXFjtDfHBy4jcLSem
9Knd9MIZsXCRfXLXFxvITcE/EOSR7TsT6LyKvv0laNFNzKoU8+bZSFGan9FqGptfpEl4gZEvVKsO
ACKf7r5MuqzXCnT91WrXII7FWWbVFQAiKneSP4TcZT+UQh/A88BGWZVmPK0ETBT0fho6JTdiQl8p
pNIFMWCot6zoKRDd7XFRzegSbylPbfepdpzAK5Ca60uv1bcWAgWoAUezhBQKwSKeLxA/poPNKcfG
Mj9uYtmtQOE5Z4YqyDoWtjSxrUAWKpWWDOWX4Xiw/ZPtjrGejVKRAYuPDhhrTBLq1OXksYCF9F2I
1GTmAA5FmsU1D39xTNAjmX1oFFwx+uQLZI8LcMj4QgfHzxlL0duWMel3vIoNT5mq1XZt1R5x/SJ3
mOyvhqIDyN9BpqrdDgOSPNouoAIb4wKOGaHflSTXCCyyHAwjEDvUqm/W7d2U7GgX0g+S+QZk9Tz3
qRhUAESsdKlPPLlNC3ngJJeYYZvFMZdqbtnIDNQkUYHn7//gLNew7S63p9yXZmoobXd22Ul0UEqx
vo84ter+E9UnIYmdwWyIqphD6vi5Wnp8+CbHHZeqy+u0SX/T/3ZBnxrwTykYy2c98hnEZ5cmLseD
/M9zEg55+1CL5168MBfYh7lB8EfNvED2N+gm+lgr3hzHqBmNe7sUD8Rtug+tH7V/xAeHvRfurgaZ
ysP4IW39Ceq/XV6PTyNouBfl1D1P2SlKX2hRVcBXMQeQxzgKvv6vkyqAiHlzAepm6GjdSvfrQ2IV
FltSO4LwjpeaOgd3jKQhJ09fQLxZRGn30efrB7pdR4+YsZExkmzXI4ektvCw8Y+AqJ/5D8J/eeT0
+CCbZfbJXk0p3/y/h595ZS7oSk41JhtKfU05RBaClKHEUEoMJKS1pTISPkzgzC6LCqGu51c56WUZ
Vgp+PKHWYwCTWRH6RAmsotRfT8WFJLNhcz5zzJ2YrGG1AI9i3/fMohIHFc9DCN1G0H/OKy1oV6ez
2fAr+FgwFPAaJK+NRfv9PPKzLeqosj4PtRK7fAGZOaF4dwIfokAAg6aCtWcg2xIVmrCGjbEeQ1AH
gSd5ppnAtZTnVpLGKgSRiC077WpoX1bZnorsKpwu3NRVy1H1I9b695OGuybDfoxoXv8I8QZtfK74
ERxZiY2cACoyZg0ZLEIVEY8JaOmRxWIJmAQqWpOBJCimR7bpSDcXWl7HANY+nY8vlXadAYm0zDs/
IZHqelQjobAaeYXRPEZGUgGrPY3gzjLyIAuFF0ncIn59pPAt9uMu3qGQ2GOkARWawe32/vFuYVkI
DFD7glOS+oo9W8tJNybSvOU+R+0wTp8QFvvOvD4XsrJ4ZZh/0pbBiN0WtGxcZzLXjFS120+BcCnX
/AG8u1KZkRNpAmgnNkFSmOfwcZkWplRoUYkp1DxQ4nVOiDLb435b1hmlUDQv1XPHcFxWckA1xbx1
d0CBjugh7tQ5dd6B0P1Q8n6iqa+qKRLJlphzSXnnlIXMZ30zDxBJC9Tq1PSKo9PCiHECw6ZfHHLU
TeGYtDd/caVi06dpNEhDCwGPww42/OQL3C+1UPO2q+4RhufTPOegL5S4T/hIKiAf2cLq/Ll9PGcV
oJHE84YOTDUL6mfKuHNcCyVTX+fcNw0Cim8oJfAHOPxwuiEOPQQjhZecRQRvy3EV1fcWnmYmGpWr
gJ63yjZFyI4CFePoSmki2tT/t7pUcg7wi3IFBB+kfhBVBgp1oWeKJ4XtBfa3Ex35bS4tyLxQSsq2
YSRXD4isjnIe+sLgmoD8bYakrk+bHIzT9UKvn6Paa4bskDkymN5SlBPw+5a7tZ0TbhNitb0UukX2
nhYmxNVIiT7Z5AjTAH6cwG1+1WfrlbTu/fd3z+hhDMnnaycWSVAbOpjRZimZhg7+FhmfrXD9/1zE
sUmB0NSslPfd1bY5uBcbTy5EHpJQaVfVyJjZWiR34K5/mNwM1uLVX/FV/oKPooYykmr4veC1ztlb
cVJOEG4d0n81Cg/eoMHuOPKvl1JWDGJIETSG9YKJz+tKKNRlJgdfJi7WpL4lYog3t+3q9vQRhKLH
ZJ6pY1mgVnQpb5oeEMNf51NMQoHnKvFJu0T19tJb8wuv5ZXOJ/yC8aa5iUlZE0qD8CdKR/9OnKZu
+KcLv779WVxSQzlZ5+oeyEGmTAlzh6tzInYL65XWEu4JwSfMAFSaf4Vd6653o5uPNR/jEIalX4+4
rnAN+GA7F2YfQUqW2NVj5N+Lz/XKA4/UhrCIuRzg7QK/OztZhieYEWkQrstimS5/OX1lgRv1nwiU
5ePJ/w8y9XwkUu88SBNKNq6WEy4mCXaXg5FreZtsITJPuWK2X05FK1D6+CLo8BiXOkOWKEEy4xV2
3wDJ4AM295ACKSNzBA7wwa5UvQJi+WSWVbNGqcBQvA6Qw0B8Z2iKGw3K8TGeSjFGon8O9NHQ3xtQ
JMU6ENwu6/PSpzdzggjTu8xrafO1isddeAqy4hm7wf5b+uGqclWany3HjDrM7CjUmQXjsDvnDrN9
JKvdpVb9wwrjCzbFB/4oTfEpXeDUz0zmVfjjJ7jsyAwFH7Omfm60oG0IMB0zOAAs3OIj7zKOlr1s
Rp0WUyciUUdXOrjHuqhz0UOJAU0jrWIt40gHno3DGFYTQ4UFA06HL7TqE/xhxmJmlYU/Ra3oyhnd
i8YTGB6h21QXf6HgBFVh5fb1N5Kzub13mKwEXrFRQls5olucjl77i2BjK9GuRvTTbIJCCVdCN+de
2FcAgm1VJZaa+ZkqCpezkqiDpCu6oZxrrcK572a5R1+cNeAOSGIOcsgCcRXkH77p1OlEq7zAwhsP
kO73JjVCSLEKxqK2b6Nz85m2W5fuOXEWql85kdaz6ikUEpKeXSMyCS47Pf3q7B7Ld2z5bmr0h4cP
PQ8z/bvb/H1Tz7J3PbzH3RL1Ybja8t0LweCpH9/Mn0i1JPhFsto05fKga6Ak8BIE8gikj842dAsB
wPgK7r+i6ZwZJq62Ns8CDQNudzE/+5Eph+XmFWe+76TXwsMOl/YNg8s02U/PiihXdeTg9IpEfO3q
qa3OJ352B26o4rK9eL5GCUspLJ1sO/wOvwtsOzzNmEw+iw1KqE9NxcsLW6Mys80jumwHOcjfDLn/
982Orm3/jmDSbFoaWU2poIo7BYWk5/c+BHp1blXRicSWEgbKaK/xRtkbSBybTD7j8UC1vz1Ruhf9
3tCnhABKOyuDkWURlmHJI7hgS9eigFrN/h8KUGmWfVZhEAv7K1Cv7VK0uGDfT5+xAvHP3mIBoxQR
BejNs4qGlj5l5sWwlXxLZ2q22ac5BpvZXN1OXVVuaQ5xNQVkgHb75XU2LAiVKbrYW4qJdh03aKXJ
cAZWBEguP7AWAs2YD5ejxkD2HP9z1TlY/4/eYOovxn9DQN52x0JODOv34kaibm4Y6dcSHhYHA1GI
vqmY65i5a+yEjNCXontzdmgIf5MuqQxkrE7U+noA71ijAB1nw+tzsT+A1XKRCiInaqUZCqfqphhl
H9A6aFXqMafGr026IVxVD179SR/9/ZNIPTGVVsg+n1zPrjyrSimNNW8xP3EopQ0LDEjrcYSAb2mc
oFvj1RvvXg/BnREVgcv8LwBcRSt9plkqU0HVTk3OYm/LXKwu4rH8gLQIHrJIuj2EtyYznW5wNyyD
If4tcSq+ydHSsGgQG46ZXdwt5ykZOzmZ5OWBJKImAOTAzJ3/f0at9uwMZjUOCSNdj8gL7/oBU8DE
4iT+tzogBsGcTLH3aYWiO1Nn447VdInSjrYhyremvsXH4aKfnMwDiRXxa29EYApaTnAtLv7MQvtS
IcF3fY1aABa0Yob1T8AHVfRSN7eOZiDTilbiOiPa67j/QMW7vcugW64YCMSOQvZM/RL4ZkqN3IoH
Ozv/jIouGFH3TM7iMQWcqGCJdSKwdVBJO07zd7/aFv/lza0NyAXMMnAPnW7xyT0MpW2juIW4FcL4
SaDh/fgoPJiNdK+XxC/88q5NGcl/6irxTg8S3mP7SWzo/a7GC7rvgCKIJAIo3Ywne40EEPXGOvk6
PMQPrGncKN00QmIIulJI7wzjDmi7H4JI5fMKQzwUojmMWwy42AP8fSIUaLim3BP5oCAHYcsraYBB
jbcq3ozrZnU68y3ZeeWWATgRMooQw/Cr8lj9IdTxK1EPeR+Bq2TOVetd0dbivTGW1GqpZxiA6WMW
zMhiLOg4T7+EpWKkOSgQsODhteB4sRnD4coNhd8qyl991va0Jo20FxfUTkDBa8QAHlKWy/APbzet
6i05Ko1yg8Gwe99s8oShs2XXtOem6XRLWpB4k6KC7H4I3wZTDeyNZsM6RjKqC7H9h515CHQDgn5J
/Fq2rNa7ft0xafwNh6FQWh9Zj/nduZJEp7wxLXnATiNuxV+6zWiXAQc8S20agfgdZQl48JHOhV3Y
0+oziNTucBAQx72uEOy9SzuuT1BWH46SsSU2I68bhMvizqGt7YkiPe7FxeGPWQ7I7tUeAMsYP/TF
zNr9ZWv47mjjpHShPG+1h3dOy3bfmhl2zBIcfXjS2IQGtw7ULKscYCbY1rRxb3mmaZe3V33fDhyr
48haa8PVJuSnc2eTs3R7ZdxQycYzuwnGux9v22CSutDkYixQItLPw2ucNBj9k3LLpTtF6dTph8dE
dSBuN38+e71VnDrQmeUAs6tO+oK1h26k3KqdCsGBHHD+1yqgtMs6cWCVLPtODSj0zkpXx9UARrbq
Bad7Mx3pXW88B2/13zk3KGvSFQn3h7k/Z3wnpDSwUAjDsAa/wnnctbp4GRSOsOQdtT8WeaQ87aLf
mvezZEYsDAgseOUwAfj/GfdnThEh4cVdUCs4YeymEGI91nk8IA3zGMscQlEctfQmOLIxLOQ+5DPb
u9FgWMqyrbIuZ1mBGWHSzNEAcEKW3tAJS01bPaSOoFae+9AH0MMPGv4jq6DRcUOh4Kkoekaat7es
TYhPjkSBwtep+1rN9P9bjuj8mp4EXVfGZJeYanVapU8KDqS4LImB1rAiGB7qVKm1ZeXhA0rJ2T9u
5KSDH038O3lOQtU5htP96d4/t186iayopgr5tw2srrnsZ05trHbUUHmf3I5yEOIxf9G24obGQxWH
I2toi0WoGEmhdwbP1jcRHw4S2fkgPGuSW3cNXaBKgyEcAVSml8Qp5Wb4VotNU/HuKVL91uREU0hD
rBIngOj7svuTbYrbdLZU2uAKVOyjtK0XdUm5Sh88tKv63ZoHbBaZMWt/+KsOwkZJ8Wm8r1F5FcfS
9aWWYd3NZtVAp4sbyf1x9cUODFOHCkDNLdciY0fpfUZE0RWt23CI6xAZHhT0EAj98VDX8p6sr+7q
5Wks5+jy96rIIRG5NpsLwY22kY94aODNebzRy5/gnQt8qr9f96b2ao6SptretMMYrGSX2NvHh7l3
uDG1o/zoUvviQRPZU5YDIfxaw+GPfGsntTvK+6DdpSWCSIl6Q0+9qpzHJMpKoFWSs3iJZFLKK59A
rf4re0FfKuo6kZBFD9MskftqpkfFuwweSCHW+Q53EuLUfYSrqbnmYWAbBhRkJiKcEidwhpDu8IJt
dzX/9XwbeHUFnqDf1GNgHnNezr++i10CTX99W8JLBAiuGD55u1fjRoqBteO77+imGjX1umsLkgwM
M0djGFLeHOvJhUFZclDCirYArV2gfb9vMxXZdB0ssbbUUrtd0HCNvtGVDDEKhLRCUs702x5YwvSO
2H8WC9dL1Tl5pwVPU1yAh+83UL9YEKZ8oWJRSGp9uc2aS5WGbvm8NzBnxwi1jVmqIbG2eYE1lANZ
cHmcOwcbCsKEsaf2+XLMJE8GF6/BiHLzEl84RvYnOaeG7OFtDz5RVWmq9UN+r7QMhD8YJMD1tNC7
YrbXpt+9LAPj/fKryoJiv2NfVXDenemQcJPzA1PcfCQajq2yjbEc696XcQBimgSPWAwajcwPuJul
w/2F4ZLpQKKua0DxpembzuDkzd6gctxW90akqtl6DP5c54HHc2wosF6Zlh8u1h165Ioya2BUJxb1
i7RQvdnGqD3BuplzSieZP6F+DvwLn/wlf4s+O/SinsrbDM5ikET/lka6MamPUnK1KPcOXNBOS+7L
AunBu4GKeJhvqGK4KDEfnfLH5+a+qVzTs3sGB1uy0IiOGx8Gwkja0n2pi4jefF8PI6yp7Ohp2E0H
8ks+iYfQdB2KKIqPUZGlI9JfJW2GtEs4nodxVx6XoH9hQ+1EsoHP0H1G+Rva9HQVE/xKBZajE7l8
B8mSnvyQY0POdNH95L4Nor7qFfP3ODrgNoRbe/R8Xek1sDDq6YNSqopnXKQI6twwt+wr0xmmplBB
PkK7HpWDCwAPnu6vkMcgkRAHTH4CIcKmrMVnplPp/h52uheaPmeWxr0Azsx8pMFKkfedoVyZTa1T
bXb/8iLL8v8HoU14PiQSlLeqCpbsmeIplNTwaw0oYIz6D6vc6f/53MhBSkEeooyT7xs5ay65EKB4
iA53hKqB0rr33qOVI0sSDO/BkIFrLvQixeaFr4kGva4u2TExSmG/sWuK7eUtdFJpvLd09vTBELNV
0vw5NXiyuOmulIhLNUQRYFACkhOyxsOy4g5nba7vRbYE6wNvS+KlzuqKZBGpWcCiCXUK6xIP8GMF
ulUa34Qo7pNnhqx7zqcgGZQQzkoF3uGVuCK5SzNk7lR7JE1zWINPkrJoxO4OZ1EmZkg1CHf1CV5T
Uy1rV+Q7FOlZydyGnwEBo1IJECkqpw/uk0vnKblVblbWiEi4sO+KUMXHGSLULQfOfaQOrExD1HuJ
ROngzd26+REIGuP4zjDr9FhJcTrGhYZgrHf/VQiG1gVxZ8iYhhz5zrM+EC4cKzJh3IPZKl6qmKgK
tsJd1z6bS2LKDMkJkd1UKyZLEOhCvJF1t2Rn4GdOtTh2dSaS1T9gQT9UvJntibMPeuSyx0Uvl/Lk
bEbLVaeV0D2VJ2yHgFPn5M8Y195NQU1RTWWXSb8cL+OGU603v8Bv4WvVkpNNpheuomGqLCO+bYps
O+TpjsUVphHgw2nJ6DKpEY1lF6arIR+FJs3QHoMsjaLM64QqpANilqZXUtUglUqcz3L7ii/W8ZKc
Y1btZJWAmKwmEU9qnaQpUwFRGXGBznsoUkw0K8lpMvb3rn9vdW8LQxo3GB0vXZQenPgMp7NhRSBu
sqFkCwhXFgBPbKU5h7Ja8IcjLEflcFUB6dcJnsNjbkKboN/0KG5YWsICZGZpxFfWv+qiDpAAri3q
Gd6XsESfDAdV85Y4ehmqBlOqqbNjXpMI+9M2RN7YkUuZaouNnnthR1udGOFK3livp4/AqKIobV1y
UahCumcQhpyctYyTXZFhg7GJ/EAykopaOZForEd2vGGJXx9uScrr4HeG7OvdCZ1bOoM3mc//qhwq
2ReSHkGiUAcJ998QRaXEdO+LjJKVods8K7eT5Z0kCmqojlWfHxn/SHaHgX/3w4kYz0yN/exzMr0m
4m/AlaQF0OQV+5uiC/j7Fvk5PmxAriVQj8zeCVSgIx4U04VaRu9EvVbDMeimMeXBuJtyLcbsVh/Z
G9R5joDZrucPIwN1F67SUcDo2DDH8cnltC9Y4trSJXw5eX7NdPo4sMZVPJnGFNgvfAcEZiUoGaAZ
PCD/1fQnKXINVrhRmAPh9rKIMbA+ws03J0upfUtRgj1VjnvFGATuwPvz0mD8JT4p4KZ3G01TFj/y
h7FI+avtJbvHpS5h0ljU7JlJN8wIW3Zl1DLefws8BAGN8OzdrZCQxFdnjGZ6kIpNCsX94xvmXCqM
g6KPYz6kLoRHx6uROI0COnQacock7nVPIB317gRszkwfNHfRmpSfUkI0o0bjZ2yY5QymmI1chbk6
eB3/w2SK4IXVrUTN2WYWOW2DAi5Y5osJeB0bU9gCklPibkSyNR7DwTcrkyY5dTK978MfqUBSqejw
SE/sM6G0ZqgmE+0ZIowLdcIDWvRU/1nE4FOMyAYsEyEWJk9bQHUWo0ihz5s4m7ZUtg9Bjf8bVYJK
CT2xY0Q//e72qU0zCiztVoP6gDTaQKB96naUBBHoz9Unu/TJmIzomFEUAgkrZZlz/7hM/3beS8Ng
1VHQ+Wif62lZv5R5VftNpCZPzLHqI/BP2PJ14Eh6S9nwlE8nDdh+F0fUevZD8AK8oaJ4LcGK+F6Q
wljk3wM85+dvV/v4CvlduFF4o2Vr7WaUwXnv0OkSICxn1kxWoDbpWU+u7tHwQjmjPfxf/Pw9qVLj
7twn5o/djHm5EMiNEh+KdCCifWsGuCCUt0X35A1fOoRkzD8aQhgTxK+tml39omqz/YXglAVGaAO+
PWiWOPHTPjKkqUDbB4IbhdLICbqoHPKHn2GfHwsoRAfQ6HvWkoqbPhUeDh3VkiQJuq7x387jOM2s
3fXKpcJb4xetX567dm3DieXxSurKJ/g7S1kOnl0Yl+EKnViPdSmUdKQ8IwOvHiwKEYxn7GLLZNU9
cbyFrkWwipwh0LTDUVb8Znv8VDpAPpFMXWeb6eqq8Y+7WapiQAT1IM6tjZp9wMRDAElCBzalTniF
4DbYIJSjYdFVIG+PESzD92apQQUHfuKbDsyi1t5JkFLj2eskzu2fXvoz4TdB4XgTOt22AZqHohhI
gID4uI8Yw4ncmZmPKKTLdIB3sDgnRkB0sLJ7cO3P5fZWMvSW/EaBAAsuTcajQzFLCyRZwlEY2P0X
GfeTD6Iklfc7K+pwp614PHetePYGs1S1+2OdZ2b7KPNgHUgGvaxgtwGR+lsXGFM/3mXpemRp/qLX
2IgWPY7wsEoaFG6U/VzBYeCb140fDkdc0+A4wudqn6ShSx/aLM5rqf36bv66VQdsYiZP4NBRTfZI
fO4RHZF9OfXW9J+NmvJQrpAlY8F+mDpr2x+JGrO9ZigrmzCGOpPcUFFc/Ni/kcyb1XYEEToJgeP0
1767/V00RaGwRWgTD9f2qLjE8V7dVbQvjc2gqRU73dS9MThvuAkshY8GiqVfTKWztlofxF6ntLHL
Aqz2ILMfbZisd58wHABc59AIA8GNTt9mFzR1xIvksgm9PvmcVeCJlQPSd0tMCh2lQc5Qkb1QzVdV
CMI3ErnzultYaJdA+OB6R5nEqZa3Uw03nAyKWTjjpufGWy71AIrjqIMchrjVtVYrr29uZJk7hMlT
FWnUGXDUYqGO/8yLSeAyLex0TFmLwv+PutxalsWtzfenFwFKR0j+X+6QYh+CXdvgWP3RsGK9zC/5
fUgBkV0gKA0a38mOFGPa0UH3DNCFWmJHmjUbsjB/rHmKwPYZDKWCv4s5eQZ1kqcwvT2SShJHtoyJ
6GMTTmirBNV49bdvEPBfm8RN9MfSQgViw45y7eV2VW1oJbHqe9wfLPC6wfIeztcsMvljUTJLlETk
53UCVpxEc97pp87hl90tp6+0rcrV+0gaHbpencwDVxWjrdgJLG6T+LR7DQp7ce3Fhe0UgLFM+efl
ljwITn+sXCkfBnLYuz9ZPrBANNRNMqOPK+dj6puyB6EtayytESNiCT0ys9shnhbaJy6p/0+wB0RJ
lQe6NY1cBK6wlbRrwVNr8cXV12EPjDJyQ9kYu5KQEUs36DAAMtSyAlKhW6HjMHNe7Y3U2IqE37Ab
g0zMwdKfePF/u0wvqR6BYyzQ2dYCNDKPOHAu8ugwD0IGaMZd/q3Y2bWMj4SBd1lZfcrW2LKf+2V7
oAivWlB15aTpIM6B8G1aMqQKYHcDjxH8rzy043z4/As5xZcQRTCGQq+NNsneHuFLg9NPiOIkgnbz
sWfvEnSbSeUzowyFFfFcy8qPA7j1JrQvxbOWtAyesZytRWTuSshkorI0DtNXqofQenQgrnvgtNMZ
jTPlwgNMDUWqbrdc2su4D85Ad5SuIrkLC9O7gtBHFN0qsn7stk8wdlwI/nJV4xharrz2IkRnqlc+
gc3yWyJBbKq8AhoMkJsNqJrikIRhKbkze2oJmxzMF469J0YhmHK4cqlPSDOxm5YfhsKzAdAHw9IY
OSySZU1cgfd+Kv7hHfWgUckPLRJ4387kYn6IQVaKgSfy36nn6crNeafsKDpNY4go/JXDuzvGSxMe
Td6UsrXsDg6WcQDyYlUXf1DoLu/ALQ3nGi2V54Jl8WeVIepxndV79w8fAg2bYTVvbAOqO5fPvOEO
BvvuggZ7I4HppvyzqMAt0ET4UMI6sm3m8vTUWGgEuHaOrHoRGch8TV+SFIMa4NPyX1dJuRwifr11
LUVA4NwZ18278C9VYkar719VLQqXeL13LRK+Ye6XJhbbrkUF33D2Zwg/fMfFjsbvOuZSRlFuVxF2
4vc8YkJ5QLajaeI/9Vg0Mzb/ttFX7VSgUkiRc4YKiiCk2BOCRuk6ryEyxUn3Mu8iXO1kPpFiwk4L
DFySXNzB77h/eZChfvz7nJSeXx2262xYzMC+w/TewwJUYrB3k9gzydfTtpvNqSuWxLHOwSn0dmbV
RxFJp7gqwDc30epBFTycQ6vSnHRynPSlixD25sfKKFmJMdte4+czCV2dE9fDe6YzGlO7S+0Um/+3
RUXGsTAsBH+KW4OIZU01sh4oto2zR7n23b4lWj5Yb8pd9XyjvUZkQ+/EpTRE8xuPlcIBQdPcGXNu
7u9ac/ATZTVZ6RThuFbjtHceXWf3u4k69Ja62BBxOeEUOKg/ADJvDpVUaZVaPop51MXbjtCBU+y+
xjyX2myXLK98M+yy9oe9q8+ZpCRpU1UK/aNvgFyN7CZqjbP3ZSKY+vUr/rE5/wzMpJ+3/gY2PJHh
NI6jIYGXfsZ6zGyCk4Lx55qCf7rchPseNUYpYC9fdCuUlZQqmJ55OHPJkmfPCCU4G3eZO75dxKAs
twDQV2o72Fi+7E3of0iWELmmgB3FhCtRkxMH4P3cw0UMJc+T445MD1acrQQFpjwGkcvWJM/Oi+cT
aMyImEuU4aKStwtm2NvTqM51EASgnzD+s4LR24BaVYIYVVEpR9/DMJ8fbgMUhivkuf7tzjB/f8o8
i/iLg7sATXn4FopqGBpL4/33lc7K8CID4Mw/LLJf0VsYPp11nvcHPnIH3vlav2w4daP919B5S6Kv
asj8cuocaP0a6uR1JtL2syqk5om8sw0wuasuJVh70USE5nduxAnvgM8tr1CXxL/lyi2KqC2NLNVc
dxkpcw50DcryL0pABbqJw5gMROxEBTPVhgcocUHW279LCDPHq7B0WGd6G06pzbBib4CxhE4TMspD
RvmLzB1LlxFz9LdkL9w0Jgj4SU7w+D74TTdcXLuldJ0kp+M+NpQD8v84T3uZ159lzdoqETq1e7ln
9loCFg0LLKv44C+34hlUFScZCBB8cyEcoTCYd9uqTkolUA6ioKiXQG0pRgeiG6cm6wwftzXy/5ae
UJdGbml4vU9ZLzVfvt5mA9asrzLu6XrTirjcGjgMRj8N9Wv6rIyEq6ODurBPwZHrf0U2Iv46MnCK
b3oUsXo8suBG4/0Y0VxcCplF+e2OeucTCZ5QyKGtOvzxie0WSGBh/HsYYizVoXk958k95b3sbpCS
Qc7RugEHx739DgPz68Us8+tooYsu9/6n7eAPB1X1m3nSOAGgZIv7hae6ZRSgYeUu/WIXOt0AKUG6
72u4d6g3GzHL8GL9bZbF2u2s/cYflDCBqnkHW5xiWDiBza1Eakz28gHJlkJfwLfSmj39UUKOoI/6
ralBY1n+3w+9h1I4wXr58wWDPnsw9QkQgUHrLcv4CjMcnN0PIh3HS3kVagiY7mvMgFYXEOKXn5bK
S1fNJfr12vpMSikt3DwKLvr2R/oURXj5LlA0U5JxUxqf0wEVOocz+S2u51kY2PDhkW0aZ23JWcQ8
22Fs+OtH6zXmcOADtbbsgm0i7oMJUBL0dAeuP+SF7TPlP6FJnAWXnCwUH47P5Y5sPr+ToyW/LqTe
V9gGFn08EQ61msX5iCs8BNPFZCDniUX+gdjMvxn7fBYRN9F+Pu/Kc4hYUF5jrauuUfCAA7iGx0UW
atiwYt24B3y6VX6+kfgzJlGgiWMigqghYZv2Sccfp0i5nG8Q+EXtJw6c/g4GEGvjX3v/kYoRPQof
WdvvN+NCOUH7/g8bHzpxs3bDIfqQmquKAqTgnj8xNE4lrszfXAIMamgRUIWDm5Fp9p/RN9YvPgqx
R/7D8m2s6iJnya5s59iIN5OSxj9zvG77xEZL9F7bVwH8Bd5gHogUKfrpBUGH3WsDWv6tgPlIaCi6
U/ZOyet5AtPOGWzfKnxIlqOCTIn9ZzLB7Cz2MtF204I1huQkmy3z5iOCYjuCu9prGo+AAYzEqweH
c1h/1KseXZAyCW/n8n3wUAeuHRJr3sosoDGeiMjE3xS4iym4XmROXsLA74xtZI2gTXPFZVuJ/CG/
pT0ifaJKCB0JZ92kNtIxm/MuPI125U9BVAERPCA5oPEJ13ODIdVW8K3jNLo7vShbct6rCX0Psp9r
XiH7X3iBQ73cp5BZTWVEuC2Lb6bFcmRBC9NtjlZPemKZteKw6Kt8JQA92wNckV/FyUtGuYA1XAbf
woj0Hkp9AqXNFcDwlVlqGhXFVs1IaDOQqKWeeEJr4cbx/oXw16Tp1uINa3b5TLxNU5B+tiRwLaMK
C+5sBqi5VDgwLrXkORZU6vcLIrSUhDEkkSeCQpYqhv9BFACUyJDWnw3TwhPsTmLDujAXORMUQpwy
zhxLWUaVK2bI3h5+sGv6rsPCzzsIMk7n4bmmpF2hKc++sz3e8yj4K6X8UapwLkmuz3yv17/EfyAe
AXZdj7LU1UyY5Z1qNPqofVL8uW9eYOEEeUJOWTRpcUGQ2iQk+k1U38y/ZAlVF3DhXQkb4wLzQP86
loWkYrElZNgTgLn6cZ3SJh/8BTSUW0pywsi+UExPdz7JwOu0b0gLCHy+RdYmC9a3Tp446spidOk8
hWXJxY+jaOEUmLW99YoCw1GGug/LIQxRr/Bml5Ir/sB8e+B7ATmZ4jjrkj6N8DaEmv6OZprx1aZY
VZOoYy4y2ixJmlPAyvu7pTM9CuBeyl0fdazBzg4t9jxjYudohGw4FK76mCgt69bg9Y1ZCEtgYHkZ
WljouBSlbVZTr1T/8mItxdzBB+R8PI7/eHfAmmysXvOIeyXlvCDZM4f1p6eUF7hK1tRvJ0m2qrlL
01hpsJuE9F85IKe82zkIx6vSNOKKjgxHP45OmkyqbstvU3pLnnpmurHm/rpjqkNrjwWnBZXW0zLq
0zPNhFDJZ/fIwvdeumEysERcEA0X350VWLEDgHAUDRzM9M9M48MByLpaaRyQuCPazjQT4TgMt+Zs
d4ulfSTdyKTf5AYmHueBWxEB5h7S1uDO6oa7os6WjeqDR951AgcKivKx5uj5M6YqwaYkwBMxRUO9
ZVoq/z5A6+zXIfv3bwS0wHo8iOSEIArEVVeYPvCx3aAej2sF9LPEjAwkWRS9peKf0UvEZW3+U8Xx
WRIq6r/p8hwbieNLE/oMkyTIy30ssDcIT5D+feqng/mR9T14lgdTkqP2WHfXQK3GhkCNJHPPyKdQ
FIaCl4+hHhEafrKihiGk7b2t8xIkOg4JZjb0asSa+QlD8XF9TAWmpkXO8OzwPw5FKPOFo6+Cn5oX
AI7YF08C+CUokuxPjwbSyqsJ4mnL5TkQ1kavbldwHP8HqQeV+CJuQpHrLK5XOboAuNbkRYwQJ6vZ
tFVa9NLXPhnyQwrqGnH+s5B6G5HiBlBeZfX+vByVtbRezYX+3NGmhWQIvpF6lUOMBiRJLzjGmAIm
COV+4MEDeZJipB2VjdRJhkjh/QRFucn2mCHAdDwxQvcYdohF1ueOCWFLAdPjHrDZWX11nmOjrRO/
MTmIx5uboo7XZSzV1tFRSNjt9dy9ZPePea/3KDNlpA4FVwJrRWtaWq2uFZJOEQkordswouXGA/X+
ZbcRcbtX2Jx7tOdZGiTVvQswmNN6PQk3tTMPdTfPh+2v6c6K9UQuom07DdylJEip0mIo0pYrADN1
3H4aYryOm7A8sgKnNfLeIR7KxtAJEbIkkzCqGRkTs4AC4BFzmp3uY5SeLwZXwqmQtlTX83nJdqiF
q//0OlNzWqB6+OWd+i6C6BdrvtxtpQvEG78fKM46qA0zMUfSKDBqEeiTQEgNKJO40v3FavOTRrsV
Aigglf2wdeZ4iMqsfbeUBd4echyu7GE5DR5b+a4lEo/S/UIr+CL+4cOn/AlRixICMfnGd7+6qxOJ
DA2Lh6PrWg2k1m4Cyk8FTfxSondDiyr0ltz6q2uw4HmiEE6GW4uvo1rx8gw4O4FAwHCd4SDSxFUg
q0m55xN3U8R/OvmHtffwjpJfbMUEi9SrM39qvkURIBMI4FMCcvkrXf+Vpt+eUsC/mTUQs/R21FEx
+PLyolPrAWx9Ek/PlfSGLQ6WHzQ8NUHO+CMuxhIf4NGKhTyaRRmWGjx/oeHWfv8FeR8TA9OvuRQZ
3KcaybME4OrIsVFFCLaphYj6CL4tVeYQud5bwW2b6G8ssGHzIsVAZP4GA5EJATSyBdMrY+NSp/LL
AzRnkJfbgZmK3AYnhqftMOTlV/s15kSW6UX5AqLgnBxiCaH3+13b6/8h7N6OfYu2/UlZ9rjhqsiT
mrJqXKrYoweIqlC2d9SohEiWm1s0pYYhu8QyJ9EM6mk4nxqJoxW/Enxlu0TA3QnarWzufZ6udWC+
ZAVl0vS+pWw8XvUaJbOBXqwaho8wn/r3HEIPxR5Y8MqlD0LbkrDwkeJpvZ+NhJ2iRVgFO7jFm3pv
H2e1eu0cGl+OYUJfC2qsQewUGDyEamWoms0wJB9DyjYzdyicGmpx549hoHczA0MiGZ6WGSUH5KHt
ibfTJaREcTpORYhvZhDjlQHA9+cIKnwjLbCW1DtW6b5yTZkI3PFfp3sNqLmxgZQfQ0jdJOxBgsTQ
tuaCWF3Cb8EXEGeP/wvK2/SSMKu3cgwjQfkHUviaPpx8id4UOzUopjNxmHK+ZeqqxYIxoNMfJKsL
qA9E+Bj8XMsbBRA+XS8BsPQUgMn91pQaUG9Mhv6oSByzhN1foijym7Sg89AU0J0ITU7dnRBjCDK4
sVAhqgABmb2MwZkNvwY+m3UwHS/DH6dWlmODDufVlrpOFhC62m6FGLddOnf8uISwXp5XHy7bXGNb
Is3xBfzfWUza/XbM9lJYVWJj/FL4ngDuhwol8Y7zI2fvQbPD6l0XS6pptbtP0aSils38q8tqWJT3
erncOEovvhTaMGBmKcX8IlpyseS1IMCUI7b/sUc4Tc4BFeOTWSPsVLNQ9h/NAkSY+gDBngD+ajYH
jcBEvRVC8VloMBmX4KRFFryh1r23GYE+5bCRw/NpSiDmSeZxEPywzcz+0HZzT/3wFt2/PlWNsPJo
veMLKanH/vx7wop0JuDcTXbiRc+MonvsujI9EUgO9x+HM8lWrt3bY26gYgeUahmaSBasy+z85Dcg
Pd1YBxhNPzdu5hqP96hknVK1tLaU3cjMQjfik/Xlwgu4RF3w7K9wtKCMREV1lsAKea5/VpWsTAKz
Fmk+ucHXvcxtWWwjJaE7PKckeVyB2uFi1QW3WfGgW5DuRW/N1zY4hBFKqz1uvCVFQxXa2eW8vxLQ
8sqarKLYQF9zNTl6JmhWruCaRqJpgcYNWgw8fjc5eprzRiNVsP8WXV/e8MFGJXjEsUiu9iPeRCK5
uxyeUYuWFLiIR6f2WD8H9n7NAsy4g6C0EU0rSVIEaWvuEwu7RrhVEY/qXk3GeNbRYiXR0nQLMvUC
YlCLMNCMrQHUCzZexSvaXnjwGG/21OfcABwolP4fGmcldYyR6BMY1FSrHw/YRkxSBs79RHojYOVu
fwf9bsfOn0s7mnRFO+62vf4vRlCx+i1JpHYp9+Cjdqq5ogu0KJE6ZgAkyn4p/VNdJl41LWK25Y1I
HX7rVjP2kki41/atXzJ2lMVyZ01HwJGas0aNFvnhNw3EWt6YOzm38qchDrGVqgGwUgW12p5AMx6g
WPuuJfSsRGZ+F3fyJgFgTJuwo5LMdFNThN/QOT42qRWeWGP28sdTd8RLwOqG/I7oFCMJsrZ8vnoP
r7nav8sobM+eKgAnZcWv1ZKgCcCCOB/pSLeEfDM62A/APoxUomoDAovIEA36kj2H/PlXIlu+jxhm
dr2Dh3ETLVCh60vV1BrmegE+Y3E11+YAUDl9i+tYr3qhPl+izlYWYJvf1yj71zNFB2TaMsGWbim8
vu8IEXdsia0orjUS73N6f8UgfIsYirI2YVUK43039JWnMyZ0BfLZyw4mmqNJK9ZprCeVin/qMjMN
BcwU4N7JPclpp6URK22ok/owozaEb4drcz7Zy0cTqLjOmA8I0b0yyrCgqRXMx9qR2oFgiw1IzC9C
cs+kGJQfZdTDxFewVkGzD6lc6aFgPIjisfR2IrKGhPiC7Gat5BF5GIlxfHyj/R2ZtUwk244PrgiY
XkQpBkdFhfZiBLRfR1AOD/t7Ylg9wErL5Rwy30RY0N1BX+5ExbOLQL4e2/fTKeXAcpkjvewEbXo4
rOXQA2DqaO9Ga7pkjb6YaT1sVSuMizzW8Cccusab/6hoYO4z+fmBDFX0Xw2hAOlo/L3cmc880t4N
sENOCKz8ZwDO6I2RhBUq9FPoNFvnpfUPGi7sRlAgMyBCfx5hDjbLh5ksn0msw31ZpAy8SBgj55+4
Y8onZgtC8yEyn7pTxtCPpm0DUiDtQ57ZROoXdN4p7WEyMJv9tm5y7bjvo3o0AcLj26KzvsNBcqCG
Qdtd6P+dWTyHxzELM4+XcG/fab+0F6ozQ9h2RreG+/b+F7Ed/VwScegaVS4LPRzoj15ScEOfZ1MV
eBh0d4Q86bWhKb+nb+y52QkLUxu1LSI00EivfjKe+tdlsz2jCvKLIGy9E/TPQ5KVCkfM0BtzdHQo
CZJqoFnbJGal169pSIdlqUDlKLVjJh2alowc3dUIqotkxQK6UYjCbuktxJ9xfaN5xQMDzzcl6YLl
GzvbT4LiN9P/fIwzASh3xXfZcabknen9upNUqCU1r2yHwn8ZCROBTlrZvfpiLQXZNgLr8zaRmENX
tOJs2GZ1DDaFslYMpjb18L4G5KQK3adWFm6L/GbNGyFUxviHJTNFcfsC2/MIFwirMH0utO61bweb
UJ+bwomNvcYjuJn93EkhZGJ2QGjKX6aRaYm1Q0VGhzjsfq8QpliA73IeewkEz0ajyHQc//9AZuud
Y6ypbCtSiI0c7vvn/QYCQJr/iI9Sul2R7iVL8Cmb9fIdBLzdj+JE7g9cyQELz0sDH1Y+Sw2Bd+yb
FR3RsRxEfu3YzI/I8xAbvMmHlCYQAbP7Vkhp8RongaI1ZryVyitY6mxnyr6lUpJTPVuHtNpYwhWH
HZ5A4Szd30uBiaDHIqiaqr7/Mp1y27RrFi3hrJgY/EPWFzY+n0jFqJtUU2Vt3p0ZExMoRGPaysaz
+yDfuQpWg6OIXVJnvrHLTOm0tD1+28DRBxl2Jwz7WZObQck7ASDCriR4OnJqbqGBN1+yci5xjBTl
54xe/Y/NDFlwLeyIwHr4d3sX4RermDE3qjAvB4UavaGzUT1HfEqVH1nZastmME0DQ7u3fBf7Uc9D
Qkgx4Rj8ko5gaVF/pzyW9ej8x3PEicCthyEiwwbzorI70Rw8Iv1gTNh8lX3Tur8Ej91NgIdtaVtv
vNqxVDwa7zXA63KL/F4wqW013M3ICeNbwUmxnxDOnHwZWds9da7SELv89n34F3FGyQiQtLWxAYd3
jeLS+DMjLATlD1ApS1G5WgNxCkMPKh7uz8XaNQyeewm4Lgk6uBycMVkf5MNng7e22HmiXRzvuKHV
lg9FzAxkdajCtZnAY++xXK2aTn6SW9OWxWQU1TKdQGHvmnh4EZI1J1aymErKTX16DBEMSFXTLRKa
w9/xfj3BGCc+yDqavG4YtlYscOs4L1jFylwzkPLId+Xzs2/HCQfvS1tkW9Ruv4HYZxOotTHkb6s+
TaMiEUg8D60gNpnCdmlAOKdHVNxc0iGh2dso/xRj/ncp4iDDGP9qFmDTIuojOIlBVuDNLpn1mgc8
pCZiEDO2h54UgoYeNRAe+OA7hZeg0JNoM6xaKMmSnS4Tp34CusmHGAHILTifImdk+Xs84SBS5bhf
8BR6WtTEjAiHzbzJUod4Yxknp9Q8vgERQXCYPuAU2OCxOnitkLRRZ41yALuR6m3IIXmGYmE8Dq+h
KUKVl3e9P1Q3p10Vb8jGqZfOZ+8sywOR4NXx+LtuJ7mfC67vcE/Y7NjG2ZhMY9BdsJCsJj4y0Czg
Z9/9hhFvtxNLDjFGdbpq3lZixOPYGue0J2uB/YEVq+cE8ckGpUs0TpmW+j4xUcF76hTcyVrAemkk
eAFq6sDBGQjEy0N0e9VFocyC6JIrKiXDGdLWXiZxh07sIiUGEjP2oNurmsZXXLGeiI7pxuzMDiEB
mYctH9hFr3jHMFxKGuoLYUYgRFfU5gc28iNsapxiiTEwYRYcBrcp5hQHXDF/uwC6wERNNrrAIWg3
nL3LMAjLMsJSelRuAXq83h3kXV0uzcXaZl31r8T5wpTtSMwvNhPWa8mVJibGx0gDpnWZYYQm4ih6
31B5p0qnPq9KZJ9nSf/9pkxcykndqLhiEwAJdDT0DCk8Nbu8xebI30Wd95hoTlKrp2Al0u9I6Xx/
8Kw5XFM2CMN5814mwPLxbYr1ufcQC1dqSvQ7G+ocremC7fj/ejdSuZ+jtpLtsMq5An9ujTSbgTb4
GRPz4pQTOUr4nh3lxXyBPRD9wO7/yBjgSV9HelM5YpN6v3X/E6Qjy694Qh1L9vZegySnMP9kzEs0
g4ZBD33sGD+/U1tsS03ZFAllTIB/tmHEhCNBKYlTwRxL+sL5nv2ALvMJ9Y9D6cPCgcqyTllTAWwO
AnPGx1qbpoC5u8E+3MkfXJzIjXKe1akd2MndAHYiwMe5QKqjP+OugFyUorTZMc+NrgjW1QE6nQIM
6Rd1XAeno7d+TH29nNrvyS5sCnOSZkShR4cCqis+hbX/qXu79mitOFzxLLApZkGZI+uDDprm9qcF
dog7Z/pyTwVSwIdnOSlkLOGgKqf/9tvVvI6eqa00U6DWvx7JVNI4pP4OSL9XEMwbPynWsBNlFeIa
IoGFLiDYaIdwrAFICRbsQHcJsAFczZHHVDuhAzeWNTKgZZeinOhMN1dFnzhRDfM6Ago800j9Hnex
3XYHM8ZcvUZycxBD+q3dmGU03Xw6BDrIWOxnT0WqHzWBJDube3jLoUyGUpC20tnyM+tV1sx54iV8
nuLvSmJEQwdtzuiAV0+ORQ5TXDv6uJbAa+JEP7sA90dI6G3eRM4l1HQvtqsvkjW673XNEbQvD1YE
VE01OGpdk4N/5TmllNOUOFdCwh0tbptqzJnuS49bXMFLbpMtdFXCosUoWXFCS3cggnuuiCS64I3/
+5pq5nXMRbH0DGa4RzK9JWfVy6kdo4AUCE10QkE28TJ29FanzU90kGkiO2s9JGylTYYP1EJ7UdKe
Rbs98BJ3a89fyAGqq1UeS41PT0X0cMJsopIrv9Vkt1RP1TlB4B9B6DUqTQnNDTEgvD+PGOXRHGOA
l1XCVzYBI36aeNxxblg2A2IsW1iHZjCkFAf+N6cotDUqz93MAO8L4F2RvscveZjThjdM4TlsycEx
DCrqEUSDc23dxXCh1bQb6R3J1tVTXFT4dRkURcjqH9EG1mfZ+TqG+/nGab311rDaT0gnc4t7NFpm
x5MxHBClJFHZtMmawpobDIYgFRPT8uDsxXB8EymoeOaYdiDR6KKk8rC2Liys08RWlj7M9H2hViSP
HFUXr5dvhFxLV1bESBz0BvoUAl17nP1cL42WNmqj/g0OFjq80qtCaSwZqaZWmAOuYImpKcrVgoeh
hbebWgBvbmiY4tLTdrjckkA6oEJdhIp3ll+iyW+rOmdmpyc09Ip/Pvsnt6wrY14z0xiLJCsMTDei
iT15k+ZQeyfSdOYK+Lphigbq62fTRJWhKPQaPnROPEpLCZ/UXjdtTEDHMbiW1GdcjQeim6SinPJn
VPsePUpXNUPysQLuC4u8Wv7C9GSpSg47Hp+Anq5CGDpjkWQ4Gn0FwDOcgpf6RmY66Y5j3QtKtr60
Q3eOic8HDxHEFivE3hDqNwqFgghatQihwuCEYBuHGBnRzsJ6Ua0MOfpb2xAV16x4ged1CrjuzuT5
pjgJVY0LEbtfvYnEzWE2oe81b1obY5szBGvCQSfbmz398p9vihUOzSM2xiImkNglalA2Jlrz9tzb
FesCOBoK7xl1OHSHW7ddF92A+ef7Gi8hw17jvMqca2wGp9vII7+Dg7tZCfWxUvIXqd7l0AKLZ6p2
YFdtFVpvCr6hMyOXcmbGTWhpUfMwgm8XmDteJW4y5dbvESwXaMI6O4k4iAq1wZa9BCeXNHemTWug
qlFtaNzpHXCxyINrH/0YcnhecR37iT6KW/3Iah3bYk3WSkpw8Elj2PnuRVFq6Px/Fj2KHbu5Zksg
peRzw+mS3pURq3rlgyiKZ9uE41JxQ9iA5u7XtcWTb94Nv5+j92VZobc+CK8aWV5s7tGusy6VSyIf
gzUT5BIdpcvLYwsief74VbiRLmn9j4qx8OM2AgYlI+ZXx8vlQVFclxurzRG3myECzhAhItXlEEzc
PhnSU0VIRECvi1gaN5dKQb3fOdfGyFjyk2qrtOo0+0hKHXfN+J+v7mLfeUGnUGhbaqzbFo4LkKnV
6ZoTNlhD9wES3I6KXgts9Yym7xtiQRFl8PjEq6gTxgC7bbER4nzYBpCmxB2RWMCjGZikhc2qBuHw
F8zc7LE1IwvPeZocxnzOE+7lwZt5beBRWlYl6txbyk9V6CIt+s6iZUQigz6brzjwGj+7ERBKBDPY
geLSmPbkAjx+plZ9TaJfay5Dbylx+XvWmMIBZGIAeSk21AT4TZdLrej8Coc2xn4zZjWD5UBkelXZ
y4J40L99hGbnf4vXYbNQxJACvx/rfOjWxo32V/P6eZ2ravdPFDNO0RgP1fL8PV/mZ/2gB779uHMR
lmdpR3Mm6JfHIC7Cvvk7h2g219QxbBbu4ddbnoD2Lcd5CVWuIuLir+a90Dl+APtt7GxVm9LC2K0f
7uK2z0OQ6BtxlDmgrtAaEgpx7mDJhezPw+NCccHgjyZqS+G5utMGOVX+cCBeiuGgJKaENQTrqy11
pEzVNP9YEtH8CjJwUnKIIMOw7pj3k/ptK7WLglUTcUiaBV6BAAB90+PMeKCX8GC7K4q35ANswPJy
BqtRZq68Dzd4T6I1xlSxCTgI036pq2ikxHP9sqmW5BbX3wQbNPJZYM2xbYSdDXum785zrWJS51oI
RfgqIOsssyA1GCQne5qY4Lv7mm1Ka5P+MjlLgPYrtRh+JG7r+sWoNffOKN2i5VV3kTLXkKjc2iUD
H8MyxIHRaACOYKo9HbN8XrnwX7r8WjoJEKUxu9e7GlXLGuKuD2I5HJBN46T0/ACWVgIvDcxmvBq8
B6bnq3tlj4x185x8iZC7ezyir2n8FJNgzxxsJqfeC2rDprugdYT226aQM5G5Npop952DgVML9p4B
jq6/+EShmjxZfKt4/CNF7xNcIqSRSy3LWI2JPc9GydTBZJChgPUCIO8qZCiwtgFopW0u9esK+8I+
yfvWLN9FCtG5GsksDdDgvgpWFmZC+QfoN1JajeGhiV5sDgD81o/R1kbqVvSuhxBVZIddgnpp/KYz
AA7j1zxa5msCZ8VzsclddKDi+mHT7UpTYvcgSzc+uc9KCf8/M3EUW6hTbhnJoWeW5/KvMFhKluOV
c3zpnBUxeHi8yXW83YQjcxXMqT9ApStUNot90urdOyrVB6ugM05Wk5FCHMAFGQaA2daWAi8azjJ7
A7V2xokjngesqW//t9b+mAWC3Y11kddXMOxKfBHdFPRDq/xmllM3AAfXNdAjMPsPBuUX1txhB4F5
jzC2yvPHXmna6hu213Cs0Jlf7blVWG6USa9RgMmHtDvEf0eGTtfbN+mnSAwdfzYJVvnLvznZTNQk
AqNdP91G7uuMKQBLhZH66RsvWVyWvPk8fP/EVlR2IRxZ6D3SNmw1sICYvgcz2TZgs4iaCwJW+gE9
1oNOa04ubtsOGn3j4ozSK8nzNr5JjhsZvChQJ5zXN3zR00ppQmpv7C606CPxjE2UOJaLT5oljBbn
0nqmb/P817MI6mU798LWXfOCMX+KCREGekm1lpGqlmplK2LentDZyS4RdPsfLMLGFomU6eqRm3Es
v5RdcTlDYncKpLeUdZNSbsypGHgNpOBiXHAs2PQfJCGJDLYXfNQoI+cQNNgJm5GGmr/qpzJWtrzT
zjuodmH5nExK7G3oTVOADCf5jkYVGbUkm2s3p1femB4x2TabJkpZJNMJSBXPUy8vAeL1L2lYQTFL
wiY9e8OQIqHjePLAJbgHcla5uKb1oMvfkLqtJpH4wtLvAFv3ts8DpYYlCow94SB9czCYrGbo1WSZ
+6hqOv3GIAE48o9xmdbJJ8tYwMr1WKjrfC3m9BW8G3VNoSlM3FDHqbyGy6Kd5Vsrc6DPPa3n19mQ
BY+Cs+LgR+J4IN6nOvZBkwGrT9YfAfaeyOtVq4FG2xbQVojQGHg02kSXcMKBBMrhLBy52gOp+i8D
ixThaSudvgCXJS6IXNi6WUYp8Rgvh0pcqVRMVfeZRHBb9Pki58IDE0UNabkfc9gZB5ebcFS0bc7x
G30E4d1c65zo9j/bPiJZkebPQhSaJpKZJKKcBUOzhPoJgj4tXxmJ2jsO4ZwPDD+pw4a3fw91lZLC
zQl4v7RnTi4a452glbbT7A++x9BSWsRwx35EFf7lsPd/1kHvhxGOGDuy15cT4ZJo3mYPtwzrFvRg
xCCVgm9xaC01LcWx5O4orw5hqZcFYTjPF6hiRPdCI5dkdQ1UfrsPeDD9FtbGAlDejSmzL/0P6Qu5
YVjRc9nkq1sk+pFEFk6SgTh9QPu9aJFB44TyX3gvOS+GQrYmbDWwPbOsDyuOH5/7MFq4f2d2lxko
U3y1EvRo+0EX5Gvut1WNRxX+lnX7vaFc4wIXmA0P06dV+UO+hk0xkCOqp8Wm6lHNzMNJN1wtEQKm
7ZxZn5lnPHCqpZdvle1pa4Yb+gMherb+lvEjtc42ZQp/XgPrWhtKLtDaTe6hbBam9kliVJjujN0A
J4QNqGLdFF2LHmK/K6URQ1pxzlRnBzkUaUselFUqlBCkAV9i0VVcyA324xYKpugdtMpyYepDzowR
S1iaIFVbr+dtaPsDfKrg4sDIfZdHBNYJ83j+YQGDHOSEvfTWAbe8JIP5bfwXleRasG6vgFSExkZG
tgjdntM35lyj8sf+1XKD+tuMEymEZFja8PAhWXK5BnvZnODQ+HiIwKuR3Mpz5WXYCpn3nMensDEq
KDrO3sENxpI3ZeELRdKGCQnKReDZW1AAxsVx0Os93TCie3Z2BS2GM+X9YxLIJmp+CL0vSsqcbr9P
POsyYoOQLC74xXncgmNauxHoodUKVG7AETlEdzIUqxupJe/qsezreiKZuFgj1Q9tDE1Y6ec+T8bh
aIQ4B7ZpU5Q5BBDtg9eyq4MfDem3A5WPEN1/mCDgKwsZFwWCr+YmzrCGYmkqJXynWgCUFRrvJ11k
m6DYPr5ZXzblk+EywLUFQV1VsAJNgXleC5cT4M4DPlqp2n0zGkrjSCrZUXTCaieTnO7S2AkCZGme
S6DAWj7sAu28iDNQOQ9Dhbipj9hTm7s4BpkctI05X8bpo+69XIWI1lhr/jtCr8yNDCMky2ktkcH4
XuKUdiwP/IONTO99jPgXsHXCxXZiez2vgdg/DLULBqKhN9swDYzpGS2iVvDmb5G7w//5J9r6BIu4
tBOaycN75CXJLGlDliCmPJfDYSwbSMn6sO+5BJYoKMnDczrwWcEdnS/M3kHbD+U7iZBdz6HaMmrD
ugFGDPUZqNL8g9HvDPJrbRQ5Ztb5sWM/dvmcLMtf6XrKbhfJM4WSGXxZo94dmSjIq5yBt9g4iCaM
YFV1G3CZQ//IlLnIjKIdhSw2GD64AeEhEfLbDFZFgv7obKSUgGA3g6dPydtTPN1O/jZ4tvnQRl3X
kba5SFm6MGL1vkk4hK10wwuk+IhHVcoaoINl/C4wCaqR1XpVDLMpqVyuEJCe1WJazhIiHyjLlyOe
yiWJ9d4/uVHjpwWBL0f+PvJvhRNr4jqWhc8bkMdfuQ5dSRZg0lL7WBVgx+aHilXcHHEk/Z2/QkJI
OG3oVcJ0uPnM25impccbrtSWvLWErZunTYGavsL3rJtRxDcf7xMY/gufbWhSjx+JUFnUI4ZH3lwd
c70Bp8EWI/Bq6ZGkCV1bUe4d275bAnY9qyVEJ6z5opNmXtaXfzZ6rhMcqqdzJ4fz8LjaE/L0zS/e
wZ+ivRxWtXOWAmqSjmUmD2Fa3W1mAZgJtbAKoUkBR6rpdtYWd9Utcl6ET+Gu8iyM1YYDoKkavnIV
ogvPP2curXrko2SSLgv+KuPvDH498/v2cP8K2F0CalL8M5JswHsNFukpsuPmWRyKjSLQEDgN39Fb
MM8nIu97b41a2qqtDjBtoaEemx51WCXD667va/vXedySieP5WBYNl3Z6jsP5Oaaa8T3dv31O9O0A
QXtsT7Ka63itOMuDOGwNnOnFlKBRMkEm2ommGmpH/1TsqeAs/7MlaXSIs5uK9YQFOA4h00PXdiGh
cp7cvB5jRoDM8Wr/fRnHhQOVhvLSI64yAWrfTuE9gM/zup2BBIc3/5psnxLNVDCmHqGBi4aVty5w
LkN9nAc6g3uBy/jUm2w9v5bnMq1ePPlPi45gjd4v6Wownu4bJLJv4U6g2GKpFEzT/jUfle5DelWo
TFptPmR1XUmdbZUh4Q4kOj4/7e5+VeiBSyBjBU4+D4va3PukOwFHUHAsgsI4/BJwKYt0FYIZxqIT
jHaEZbsMyD7nFh16w2blpWMkIou9YXM6orQLsSIo+FwwVR0YbOtJ5NSGep+wDxUKvPOZg00HtCgZ
wm0Jo9WVJETtwBY+k1g0fkVPT7RdcGh7PGAnklKlR26tAoa68/iItNjSYgF0obLhitf5bk02SQ0s
WKQdvHgdzynFJ7Guq2slIC861ifnumUOHjvRKXVcnoaENnkeW67xmdNCZny+YI5Vw2KOn63XRjpm
3kbGQsmTuCGU7L+m5vKCzKTnTi7XHy/ouZ6m8eDs1hkiW+E4UFtGWqh0Q+Mz/tZgwUX4K7F8DdOV
Z/sQy44qtSkqQ4CLuknGuRQ28JtGjRYXHreGqgoIpjkuoMO62ID+hnm8LZ+VJToT0jk8PaV1OhbQ
a8FH8rx1Mx3xueu36EfUdUQEpxL+tL6yXZFRK3XuQwO7jypJL/Uu30zLrKIM9Ty2vfDN5wUkxElX
DvJvl6gVPq/GK0sQlPeQ8WQE2++sfRztftie3K+6bvz+b0EHXgQs0jV6zSWdXF9JdXEJ3zxYLuyd
rrPp6oisHLiTp2T4Hd2jaVAg4p9I/lZzW0NJa2OlzldYawoajcXZwEDOAswmGrhg/+Guihey1Rrc
usRBjuaqUnhleh6WIY6DpevZI5VjU5YISS02asBtHa3Huhtc+lqpHjykKcNFYwQUolgvmt6/H2f8
w0/Uk6XJEPwsIl15CE2ULvV7iKTya6Kg0RlH6KRbjfAXkMc2jbiG+/w37r6hhUlv/rBUCLtrsxpP
Fbxq6c0LH0FntcPAjXYKsTQR7kAw+l5oOFgAwO9M2HMHXve/8bW2/q3SQRjW3uSt0Wvg/2gGraJI
5WlsdcakhgX1Wpq/yTPJYBsiKCp8AWT+0k1pfITGqkfoXgxoLZoavwzTCbKbN3eteWzdOunbQ6j4
xosuOshjco2qvxmLmoN9MwUCmwNYONoN7iOVoMTLPgSSq+K3fLz9sM+Mz8MoG3/kx1YR6d3JciGP
rvBZ5/QCXbi+Yl1JPAHqrU1uaXsD99p6bLITpUMa+3xX5TuYwkH0mCxa6ueCjgoOHomUX3IlDmmt
BSX4LP3XAZmFFccBmTBppLf84jvm+riE3nbMgiEZGfWz2PjRtZTSvb9pdRWRh92EjYTDoC9t31+Q
vtNEvB9qQNBL9/RjdaYnZ+XWHo2F3XmXYe3hI+DGQe5IUim5g7XNGa8LhIkWbH56d0S7F4/9kBEd
H5JHRgIvZn39trJAJzG3BhFPyqZbrRGHCkBbfxxMinScjzDB6VHBdAaO55wlu3Dmtq+NV5pgbLrk
vp0qptiA43HSbuCSRBeNDkDYRuxUDQJ2DnrEDVFWgAn1AfxZ7uMhx9d/v3do1RbCa2P+OmmpUq6u
sIomXbeWBLrqwtCeWB52GU/YxVFXTqfoF0NLLXcSVm5AwKcrpjHpbsP/7RDvTWRDwmU37p8VCiTs
1+g4yeoeI0Jk4SypEzKnsCylU/VlfmgVzexcj05j0IQNLDrKGyfzOZ/VwLYJpJjBeJTC7xH638by
Vwquiaf6UgRBnLO//6D64uvEXOj43YMicOZRuTTK7CmmQ8JgDE4DKYfTX4F0ZsO3VlHvwd04yIwC
/7duNDKi5T+LQZektkGP6i95UlVPP8eGEty/+ciygs1HuPj8OtCZLxbMQmrcCXHY+mso9n43NAHr
ecqLkK54Na679OTALxjM8XeuXWu+dQcFJCb7/qIWwgmqIB7SPYtAhuDYKYyEgpXnoLS8EfPSDIPM
xDPvvCEafut//5M5cyKGN9NHi4aaxq7+eAEEeEU+261jX6Tj8EAB2/dXbhjkWIsXzbULMCmlmYlK
mNpU1GICw0lmAzULzSJaCFxP2Z4StYiuUEZeK8vooqeslv8n9uJlNiYMzo0GATpEB9SOsnnM5HMu
qWDuaT6hDV9ywUMVuv5kwdWGkeUTdeGEYyOfaORGMW1C684f/7NgQWFkML0JJdbAgNw5By81mBeQ
mskKYYoBYZ+bSbTpMWikFOFVoD2J1gbLTQ1pDyLE15Q+e+KTrgmqvmTu7uoD4EDcfIJGmd3ZyRip
vTXZhu3G/259lwE5WLFC17c4SElLQGaHnne53QdX0Ln6bSWtJckynNOXErZlSuiKgleo7j0Mkhku
ylaYYFxUoD4fKAibY8jUrsmtqLOu4vYKRayEUXWM15onmJQxSEUfjSK1UGDp2IMpSMU0e/W5eFPT
aCTIVpPXgHCLLs2dfrFrgS1FigFEzppsrtLz0cYdhVmnmbCkYgFAyr48x3TQGNu17V/PbZ0KR4D7
vzP0pz1Z/6WlQgSvrSTc8Bpc4Av9Z0kgzGcbAuiAkZJTIfgQQ8tebkgiQPE0T0kt6NOuCWWpUS5t
awQVk8sfgIUDcistjUrJF52PlAh4KLSG1aEZcf2cbyDK7wnWmynWKcNsNvffM37iLjAiDeBTX+VF
Jp4nLwEys7bQVDsieHyq0E9yQ8mQUXWiSe5U2ty+tUu/JwvEtXMWni9qkIi/NEZXG3/8GMZOvMJM
Dp1q7FebapzUUOq/BTSVywG80AQX6+uh1jX4LSBlUD4Q5Hk+bCL+LTQtbXUKTpuP4X4GGRktYJiF
DpCj1bk9Ub3u6bfh1U+4ypz1bUWGYS9delfq87o5VzsiZUcog9LBawUuVKC8uyFebwI/MMVe0hW3
V5Ycyc5R817FWGS7J6ICrLIDh3dw6fP0/aOGFEkvVHVDMO2zoXmmTPu4caYIPzn8gyXnoH8Cpy61
jDyJAfwU9EkhDJkQ612c1Tng/qSNl6qGP9Z2Hat8y0rDYgxayK+M8cZaPfLQTNhIEonacfuBR6nq
rCFxaIF4FlKhOZKDyuqVs9IHnXxQzCciTM6pGOjBBlmLJiJQDFXMnlbTXQwvRPxWwAM8NoSuQ8xz
ig3luR9753TwfAIl+uPnCFqpPWBopZA0rgRqI30DyjNQAgZB+fZjmYccirAbfBENRWz/eBgFRr3C
N++neKViheC4mbnguuuMY4DmHXU8h3TkST5jyA5Ar8zOTCZSjY7kcfgcqk6LhjwdpQ9hAOYRHkls
1G19Rkx+wsObfjEeSrYb9obNp5qjiGKlCqKRp/Id9gug0haIKY89rFS1nqVyhorrOcR9JYDNQddd
3ebIwVDSkI13CjUof/3m8AWFNefWaWWfaB7YpEdGONiY/OY+IfKsE3Rxe94MmFbU8HEF3N7XK0al
i45hM9cPLQckNbYXpE5kRMt7deWIFSpWoJKfQ/WcQakHk9HYSDDi8mR8de9d+oqf17uNfFEYuJX8
a0Hc6eDgW+89wnoyrplPFYmT9nkH03QxqfbuoZQwnUG8MTiAeaZWfj+ZrycwAAffL9pMM1KheS+o
vXit9UZ7tOdtboVKidKq/pvwjq+vFok8gN2jdB/3I1HSn41l028zMW3BH2dOzf3LlJVtN2qu9aaA
rxPi6rhaVa7dN+YzZ7PfzhYCq/qcB2t3LkgPb1p/wIPI3fg7w34rFzUVqo8cI5rMQmE8dxHtJQtt
OosnkRCTGM2eVfuVMXMJBLQSbEQubXnHuo9uVqbKocsp2MZGA8OpOEfNlUXzEePGiL+LLhctassz
zqcGho61W/klbplZiqg2SBiyZEr+j67xYHTYKc+VrXE1Z0ep8IxYeBMK3HBgWr2w2ZmXGtRsc8Ic
D80jzsRIOv4DCL5ciY5sQunwUun1Ayf51r1EwKR7ID09K+NoB+TdpaLMJRA5o0YNTAxFBmzbp9XM
TSWOrPx7oAnZGgQgH5UQZXaB51iM6KFyOvtXY79SLZyekQzIaKQi9+WEnkMEEnI5dBmg4JwQa6yR
uB/S2iMFsxkzzT5QOfNgkuqEAtzahK0SDd61fwqQhgQ79/rRGd2ud1DZ78h1jpLsnkfc3UFCP5Lb
F47IgVonB5RRKqyFV4IBi82ZbeqFkRtKyDvyjhYvCcp38QtFRnoNV18zCKLD+KsnQTnAlHU9nMAm
ReZcFYkiyLLa0nPBMCIMi6DHX3QeQmlw7pUX+7Y72opbnsm6othc6PbdPaNnlFfhkmdd+E3yO4BP
r8mVKx8z+qTAGfF8HpNyHbTZicXQPlk3gk1g9GBeOOy2mQHeCPX/sOtCjTXguZwmPOXBlLqpclZW
apQRWc6aw9PUbPL89Jzp4+4ObSAP3P3xIaSIXnHvwMBf1Enn0muvYn1b6M9c+jTW0pbV6OfOzG0g
wATHOhmeh8Qdg0D6gK80HaPS6t5lHoF2zK78DLsRUP0jmU1QKYldZgRWb8DzQ/Ga622qk9L4xzxE
OkYKTLf2r1cKGYoUq+tJ74p50pNK1nhMjdouRNNS0Ca2DSWlX7rhoGP4p8pzYYH4eGSIvhvHF0vx
b9lgxNqdUgctT8ExRJ/ENhA/V/CxTv59PN89byTV67OvEggHpO/LrfBboeQtsrKpuj6iAx2xOxyD
8UnxsAvyN/sEtHeQujkPDZYB99F14DDKv9UlHB1FxgFLwRhLWtKathpY6kp5GI0m63v9qLrxSLS3
UuIV11fcLL+I7BAv+x5v3KTg73vsxFIS7zgJoLbssgvd1exnbDGA5R/I4RQrVcg1Ch3RLfRmqqea
/DCG/7qdv2WHmp9wV+SelaeMiG2HmQtORGLaNxMhrWh+5rk3X8fxanVnDLNWC0VZnYPXm3SXl+FV
RPSNs367u2K//bbL523rhtqDH4tiMIPXScnWf1jf7AZSUyvmZczlf4XXUCthaEhibqLWPQ7f7fKD
vVEjuWtC8981GyLZyQBFSLkh82UT6AaqGiS8/EeIhy7reEryDU/Jd+OCKV1d3MavOWCEbNPDvq21
agoAAO6Srqp/QcgKyGz/jqRxovin8vpL43YMdV/VPRYp4tZmMBzamTLGgsdd+5vvR5ymkbuJD1Q5
8UwygBqv/3kAdERCS2CUe7jtFZKKbfs65jHhZBMxjPAz/kBkj2Liyvg9+RWT7xmOfQXod5qa+E5c
eDuzJCS8WgVe77KdctB3jfetI8NoMBLuVzpKqwCRrLvMgsf2WrprC93oSoNMAKn/s8vEDPsDTkCA
OwRmFHqjgoIjekSwTxZ8ixxAwNVPhzgysNK44+VQWRr5sQf4aJZOenmDsuRRv8/+6D5MJLzA1N05
5wG5K7eCW137NPXsNs2uH5U9lkgLQe83AnYPmirlzwPeIIl9SUvDUEdQA/k0tUIGICPN0851tWx3
pbI1SjxNMhn4Ng/NuEWfehYYvEFOG1+JApTmGaJPYYzW2QA+Oxez4hzo5bkorfCHjqgtbrfNpBtT
0tEDKfof++BjTfPsGIalv9J7W1Gf/Dq+ocTMG1CH+6dQE5OSNfPZybztkbyN/LK7sOeFoZC1pX6S
ZjjjSCcT4M0I+ZoJFO+xJAS89Bp+D964wy7g0bm39kBWRKgUyMPerEZEMXyhi2RFLlKKvC3NU/k2
OEkft55r077OOFZk48EC/vEZlYjoYzu2vr7twEgM62UXwC/aXWOE3HgYWBD+BpOeTOrurnt6xHJz
Vps4pzI0h+15IoS9wVzyNMjJK78hg03dBxdXaXVU6VGWI4p7gk9BwDwTz5he0ybYVqUOnKPOXdor
jO9hAAmUcCmAuoX5rMAxwZgyiUVa4Un2JGefE5+zjfjyNIJu4HY3jo32ligbJ1LWAnIYCFJItYjP
K3MCz8JfgDAhliR/ejTZq+xJWgtSjep34FXC7r9L3rgV5NsPMML5pmj6n0KrnX0gWdV3NtULsSKb
vELE18QnppkEJS5s6fpozh9CCzoJis9iI9MM/ueXlVhcZkvpMohoXlPiZhq/RCqMUKYJ+rgjLKFJ
b6MCrLSqakU4nc0uQcwtwGn0r37vLNRR0uVA0UwVtTL3vJy+XrRo0PYcBExvVeRaekq1nuH10/I8
ArsEKexx+sT3Pq3m5iFP0fHTHK2sQMgr9u2qiKTz29bs51v8z9VuQSEu5U4NjNOrE45+C6GJIUvF
f3/YlwNoDYGClxlbMEKBHEafy8Nz/3zgNNG/auMwP1q0JBrvo94cn89ykk6w6U4QL3aJB+CSMIk/
W+zz8T+o9abO+XTsWHx92L1DBh5jW0vegmGQBya93CaxAYnOUGU4kqNs59gDD3FJYa88qoiB4WS3
/UT+8ExYU64+9vgBGnbq7e4qz0oUo654hWM8+xRmpH+6DwrEqq9tZpJ9Bin8XPNkwIQuHq69JfRR
moijenSR7zy1C5cP6+c1BDqKe0hF6xP4PI6bkyq8ZEU/YhvonmgWTnsys8rZZE4jNxsaQOHmm87H
dauyJHuk1wbx4tcIzGgl8Ov6511RHIjF6zUOX5CDhiib6Q/czM/Bbjtymi9wYsRKu+8wNkXSjtqD
bmfBmWD7J3Xa+HX3gFWcwCCuK/ewpZTI7u8/48IEBXoDSKZh/ZMvf9EGfwwTtUUIKVeRYU6M4wkP
o/C9Onwl/mMdqp9IZ0KefzK5ekO9RRRVKV3Fad7MbHB8SLA64eg4H6YKeV9Sc1uS+ZajKHHGyp9Q
fGeM3rWQYySWSHf7RRC2A45ghcPwX/GT2ID4dnnmW/TpT0LHxWWzzmOhQJhR2AdjyJDVKMxk5+8C
A5aWTfX7/sykiDDT5mhcK4kTqoBPB2qqUcvCmo64Vsutcfpn489Wm5lK8G/6L+VU68tqs4Jv3CnF
X+3w9sia7p9KKauRfgdC1nEewN4Qydw6g9vIwUR9yx8d3uns4NTF2qL7YQTFOrazbxMEm6C19/Qv
AfmuqTzYQ2rfiqgAYszjSHMD4ABSnWIXWhx2m5rg8ZdlJCcFLBEksp+fcSJgbPHEwjdbJI8ZwN/f
NSoraS8m+Cp4vQan5xaipZ3hbMpV7ehTiCqy4Ehd0aKIex5wF3dBeJroMA+8e14RI07h0bx0scPp
9yhU5m1cHiN+b1V62nLfCLkFHoU/C0AHZkvoHLFead33Lcl11m7LUSTqHWgnXtgtf6Z/TLvqN88s
KVS65bLbVFxIiH/BnHPesB7IO+4CCjkobEhoPjogZXg2jmTggNv2yhjyFA3bZqT1HZJBno4/GgdL
AIPpwKnrzS/8F15qzNny++MWh/WD7A+FLAx8PVEX4AYVsYaziTbW6BgZvTbXJOGeT4mSmeBx9lRQ
w78aJBRQo7ouU0EA/6B6gcfvm8sJgjy8OxAHGsH8BsGeAcpZO5M16AkAEHZ2grczsOecm6jRO/kd
rwAVmJDN5MLfQvu8Vt20nKOof9x5CTEiXFdoPdW62gUNvNL+B0zYDdaKTV92XwmlfRC4elGI6vgM
s7UJCHF0j52KHnbjxlpExL9bmvAEirREzq8JD3UKfd8WBgOR35pN/z4vFr45anzdLVDlop0Bj8/D
98TnNdlRJJh5DmACBmahNjta6BxymX0aeXAvvxqrLATAGHYvlCQiwufgbshNjDXUX2lMz2nV+Wy/
ZNBEn1Euwc3Lh73J9Z9AvU+DSHCdkabQD6Dp8xdQDhh3JbBC7ahc+I0vp09uuspC6Q+I3MT2PlDG
tBDaRBQj/tvyP6aqFqrbj3Pv/dc1aCwZKMD6IrMlRnyzDwb6gFhw7pG8rskJ/oypys7qr5JLttCG
gtZ/SfU8IHbtt3NdRHPGaY607hGv5KdkD57LMR7+Vo68RA2ycNaSjwwwqmyWBunVyT4n8KSIMfmd
UrcknWwNzQdoFRnEs03jSwXE+IFRe5QwLBNk7biLEmNJnz2jn3La/rAQa14PpgGs2VB5XKxf3thZ
xMR1ZeKGevONKaAU+RFB2rD2cwxXNZfFP6oQ0sC4MxV4nSA7iO4Mc5qXvphML5qd+5rQOMoupp3C
nl5OoGS8PHGuf374O51ykPQQuAzcemcybTggtKJbHmzmvmV6slgl0pGTto3RR2mm/x3gl8QJ6VZq
hcNcqlMAUnMiov3QQYeFrHyWiKIujReqN76VR36TocB0UIPtPieroGyfMS+PAVNLlOuzMN1IEW+f
Pi/QA79Km32UCDDHLihlqgz6EHZohblXUtnw6MgzfJG3VgH7yt4nwZXcoQgv+NbThpC7XU5vlwe6
MplaxE+OyskzLh4oi+XA/IffNoDIrtemTElId9bXt/qJOzetGWE6840OhqDEK3TP4HB/Y38bpdCO
4icAgyoRxLunIom8Fd+B8hIwZhdJoozcVubdHkH7O4JHpzDzq73kLqg7UE7ettGBm52f+9mUmiml
VQCHGDIkbcyF407lqduyq05sPh9GMYDTzIAhqomBqM7oHdlQ3NzwKhLgJKflBPX8L0LIFbjFZYp2
o1cXwMVGEAQX9H6LGcjHOuLDB/CmInG4jZ5Oe9tEQ7yThtoW2tY5yiwlCgK3tj8bT5+M/NMBs9KM
Wt8LU7tKYVH9dxsNTR7QAFUpsZaFJiU7B0igZzsST0NCKFoNNM4SZEXeFPpeMW46KgeOy65PolZy
Vg1CUc4gyOpQNaFs5NmR9JukgRnR37syG93M4QOyAbIIQthw6YjVWHcuPzPWy9ruU7MPKnp8p/i3
0E5Ukl2H+xpEnj6Z9aJIhMK/888vsw67nT5iYTIX7ta1EwanjNJ0CT+ThFVCqE5n9YMVBezEI9CO
BsHA8AIk9SoRSKUJXJEu5VL00eLaETUJYlbCx2TSAIHvKxZ/pyTkvTFUCw2chtk2CMIZaPLm0t3B
yf+D4dTBbbwuCNp87W65NdoNrJoEDAv0bGxq8qa/XbteNyZ64cpiiWGuFOGeMDaCe3GebmyPOTc/
SvRdGPnmT6b4y9NCzHJbTFWtbC5lceu4RqSHqPx1D0Gp6NTrE7GYSxKeeP06K6gE/47kL7lA42Ud
d8D0xSTQYzkS13spveQ7xuJC9wtj7dvarwQ70PBZfuj+1gx6KJ0iCGJLp4Jwz9xVnTU5c2s8w9hu
xYpwcmVLMmpPYW5Kb1gn4IyWd276n1G6/DKqXDuvRO1Z7SHnb/UbJ38UwMjz7nUxIGI3yxLHjceg
TRz56/hczCfz7xl3FmOeRFUwSVM2bKbQWHiK6NRR+Srxmv0IdNutHO0GuFh6puyDq8qATcOY6uFc
RzdmVC6JCIVrL7ZXBIPi1R/mAN1PFT+E8W7kIgYF2Xugzjqv1IeTv46L/bOZ9IXy846YwEpB9Ejw
zz0DqUfTJZaHLWA6rJQoEudJlPG77KDstCMYojyMTx7hFZQcs93DXYvLTz/xhbjlp/HQwQ1XBFyz
/SrfeSuQmm5qGLvVHhVbeyzygTx8+pEcWvyIHE3bLLDBXUEijJ/RDuN1yYbdMI4VJjExPZ8Odb+/
GzEPGa4y++5JCpcntoRkcIT90GRLNYDUGa39FoeHSFGEjDrjDOOLROTV5pnc5gGLmYrrsqUmtRxx
b63fU6vsghY88goxxKC7UQ==
`protect end_protected
