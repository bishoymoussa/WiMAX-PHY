-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
AtbsopqLne7/cZXKYxn8CJajVOG4uDJIuy7DmOIn0xBY+4zbBqiiyEzvki2T6q92nOe/vv9sIdoB
v7ZF0VjOfAg7Xs4AJ8LsxnsBLubXGDfpWL5EXBkgy4SMmPz/gM+UctovjQ5XG4GDarEUOQsqKicH
k4dRRknHi4lU7BUDFI66kQaPx5Ed6XqA6EHUbUFBCFaSzs5BQZS/hlwCtWHK/poC9bIX5H/8sDSB
bVwI//Ajkp5aS6uwVuYj/32JmLkCbIprc/x2PKnTq4Eg9hFIkjKozHs0ua5lOg9p5FqPiNFNx8jp
W1Clp2vgsY1A5a+u2/Snb6XiTkIxfyvlWMIVlg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 91552)
`protect data_block
9gFSMOL4tpFA/3EXGuFsoCKumK2vftclYa8xeHFiFbaaQfM3OIPScOaprGJN2dYCS+RJQ1kc6mVl
9FBJKeXBrlkGbI2n9LAtFasLL/8v+76Ba8VU7bmJHgoPcCT0xkY8HUbGJ0GrG+igQtWcGB6Y+PEq
aNUO5OHjGB0/1550o06LibOeOHcog7m/xJ7TUDIDh7XpvSAgwx1jWtWs2E+336M3hsDunkVub52j
OnCsQnpjcE0Kz5RUE+HoIvyL4Jwx+imT4T8FU4nqDpM3ruCo6ZxDEs9eFC3iL/ehlNZ3/2URp3JV
oDhNoAcQgewFfFlYzqYdvapp6oPaIQMRuXCOke+WqN/WZZHu1G588Ew6+AR+hBw1vwPI3j4NtTOw
gM3vPnVOLXAO4aNkdqbuXrfT0LPFyvpD7nsz8X8VEUa3/q6s28JGOfFvj7yRcYgDla4ptbW7XBAi
/BXhcS2JVC1njxzG951WbtuYM+1QAvIycB2wqoPcGM7qTPWNR+Ce3oGxV3XIRrxqEgJ5TNYQCxzE
q956Wp/kgVRjaKdUBZhN5nTC88NsRGXwv6K8GtSSPJnW9/CGhCMfFwcL9Zl4tYM4demtknats+Ly
NG+YqyR+YuQUIq3n40/EFOX6aY+wbnBj8M9Bcb2PFRz62uI1Qb/Y4hCQfQTv7BuUkt+7Ct0ZGP1l
0+W4Uy0NktWyl9OK7j+9JgJDbcVGhZxpFJdnBSFmxV5+7mdMQJGG+VAbmxpaBqfB1ifjbUEhRSEt
4uySaNob0AKI2V42e+9a0TANum9m8YvI+ZdyI4uxhP8S5fa10cdqLNQ64xUTmpCaeipiEvxgiKdM
NP8xHKeUZ1RlR9Oj55EOnUVwGBVRb7PPzrh5lvEpEne4cBYy8eMRHcbeJ3RkP9Al7ar6ErQG/05B
9SjhiOZYZFmmb1LflkkxMMsMgv0rNZ6CJonzTPBu1FZ3zO57Pk6ugDrOlLFAL0h1GNq2hdlbpaxs
MLvsWOwWh9jUot2O9K1nEt29PINyJGqw/qDOoOAB6khCHs4IJyKjtq8Yc+pcv66xwFdUZfuJWxo0
bjjhsUTKB5aKbOZkGrVKVbV35fjtzlzsfLDpLBzqQ75Jc1jPdtD9vwvT/6xhigb6FNS2a5bD7iEb
Fbu8qgs1VD+tGMNPYUl4MAzl9aWeGE4fQUHHW79gPLYqBipVZgnZQMs8L1721JnkcsgikEzRJbJE
82TF3KY60jbKnscQEL7qQrv9dcpSP2hpKBX4Zq0F1b5mo88zPUPNmdyVpAALkMbfCnLkc7MOkes5
w1Jn1Wiy00L6dFgLPDBQjCBQc9idt7WPst/Hd+sQrijceAKrtyjFMleHKd/ltKmLkJ13Cwt26xw0
u4+sl/SI4J1+g1+OZDws1kKLD3YwCuCqBKiGBgGIVY6vQVTQWl0O9vhwOmiSdKlZAR+kkAS3IDbH
1zEd4/+x/XwY3+1qr8WswiOjoCZT3E6wJiX+XxsQEpql7200b37wH+yZF0ccHgKEn0obc0SYGH2s
npjk9NXuZSDrXg66xvOtSBSOqbcAPD3GUDxIN+fSKwlqf0w1R29BhIoqfzGkt7SYvglM+GqQcX3p
Q2fC6y0duH+bI+jx1XPkOS0VHk2AH3EiqPv9WlAdAqMqF+25QPQMRENa4l0HIuWFoye0dXlGDB+d
XTiKfve5Dp/6BNGrq/Eifi6lQM+fJWBDJKmY7gslngd37t0P+FY87znMXCUp+0acLs64ly1SQLJK
py3QKx51wOhQDcRZccKA50Vzkdhj8yyFmMFiWEKsBlMhlLkcK6KHfe+jgxxIszrtTiwK4aB4l1Ma
iGTPpMRPZKBcLAQNm5Tbk33GRvVHx+vMnOSU17A4MSMb/ImdDIWPvPzJwf1/GYyEjrPd3wvzCMVd
r1dh/H6dRVQXd69MpTKjNZewDpsnTrlS/+gQmdxuwuSFWZEzcoftzG3S4H+9vIbeEFA26fqpke4z
t/zbXzU4IO9qHm33CF086pMkqkaYSOX/3DtR6EAgVt+g0P2hGl/YXtaCIrqo/B7SjA3nvrNXn84R
NFARRzhrcJa/TKoLdZ0q7B2icBuf5e5n16v8hxnfxxJXMQC2pJBgtEYszdR03y9dfPTUhfYl4Gxp
ZuNRWEH3/2iXgakrVSFlsoWLlJoC/AljN1BMEJDMgYhvclye8jzYtQsnjXL1hEOJoOX/jfFjPdIX
L3o5LTTS4TN0wMLxnhrFaG+uoNgqBFT4ajBbKf9+NARllcoQqJ3N2e3QOxvPQHX3UorpZwPp1Ejc
uf3ll/ix2XMV4KE2St00cHAQ0OoOMQaCMdqhCLuSptItMnIVkmZzdTZSAwpFb1m2tU8Y6k5pz1YU
lmLmpg+djNdZ8GOsUd8BDXUT1+yE39ZbIJEYEHhwRIgK6sQun8yKBWNsvMA5mXbexCz0n2gp6GOW
KxY5GT2Y+2lrN1mLAyFjpcOtC8AF/pVw4IWdiv2pkFFG8skEog0W70eqlTmR0ewCxTNDtC2Z3JhE
NGf/rVxBNmOp4Vi/melY/KKzXruJoGtpdBi9PamM1gUS7Qx+ZZJWduIOEB57vQmi2WT+OCcb6AyN
d/zvbWXZrmK3YyHcYI9beF8AhgxMfiiMJZywJWz47OQlxX4vNYNYrxMx2fLUGnB2n7H2ZyjgNRTc
ruotRQtyfNm22j1iBJef+zVTRAZi0rXAbjN0R7x0NRQqTJDVXbnu/bGSSnS+pRp6Z6JJABiloOGh
KvCyAu520/SPMkSwIPRRhMAiO6c5bXKsW3FpGHc7hwKUw/TC1yONq72M71Pjdn62CY4d/HdJpe+6
EsXr7CwFubQgrRwCPRthDmS5TvNS43Iu+KsZ0kAexgzy46MKkyDnFKaQEASOqpPqtK2xXck29GFM
b4xJINV16rWpdno4UdL6/WUlHeam84wA/xjVBiZ+uIJ0MTmIshUXNZoENtcv7zC0w/o0ocxyiCnr
QHwVkGwrcTTARKIsx3Z/OOAluU2ZXNB2ayIRkM58eEdw7TEz+hRn8T3T3bzOSGyI/iyG7Wfo0ej6
YB6YuoOtYBPtlPmH+KfGx32Ry8v7uBzmVrPuRTwLQYJ7J389N3wm+lCGFlfSA+W0XGjCWkzx5g1a
lUAz49x9YzLeU7sFs5QM6sCTn/c2rBA3DNaQQD8ml9jrCcqP4LM/00CUTQld7cTIovlnOo4MsoxS
noXRSJoXusNMzvdmLWex8kYdAEtOZY1QZLvtIcm/WvW58HV54zX8/8TF6BIEvjBkOTTI5qSt6Rrf
sXzqOeu0309vkC6C4aGfKuukSlJKPI5BpkuFcZaFN2pEgpTA8qSuN5Aw7+vxKuqLlLWopm66Hluv
/O5vNyyZFrLOKCsR9II2JMBAFVygboWyRiOgxslwNIc99I9yUnU9Qxt0NUD3g+A3zFJQZ3dRJW2M
C9yahtFlt+CSN5w01lkAWGEhbGZfAfI6oIkr7CslQC/FraZ/YwxuwUqtlriPc9gDwTg2xiJlqldA
/9A4RdZJ5o0Vz1Yiv2YWMhG3AhEo9Y60PTl3TI/3qpxMl3uVVDk3jACilWOrJTo5M+bXU2lbiZ/X
zFuPNa8st2Nt9fsyM4saNbwJPphh1gWRYVhqNmEWeqZsBfbXXuIiklefKzu7FXRQ7Pqb0TFRO98m
HFmL3I1eBHzzUgS5i/YeZ060T0AjjFEh4pBbSj9g5CC0uZ1EpEswrUONmquaquifCEP5/KYFOiza
sLhA/FInFzUieocfpQRqMla/wCvUdotylfk9eBtBBc0jo6ehvIXurVVU8MEA4lYoC9uIgS0uPpiX
bQ5OgJmJeA6+r0LgSnOeq2EscYQjrwzJtLJ5GQVAEStuS6Ds1xZ9UrDmDXSzqHHpVzGUcsU6vkms
p8shZ9pfJ46I488ysltBEu2lKB/CdBpUErfIhOQ+OnWn2zur6YnQJO+XGZ5M35EAYFMRTQsPTQOn
Zf0FUPci654cAuEyb09DiPAkVPl8GSB4kueqjI37LG5NBrvi1SPx9ODJh5DauRvSlNDxEgoc0/lc
w7rpJQtPWokIv+gQhFcndv2KiV2MATwlOZo6hocGtqUk2U66+7ran5D4dEFSusk8R8273/uBvPds
Eq7eLr2Lf57b7Ma6SS/sS8TtejOvZkKpUuuheljjtmOZ2sum0GXjFFSe78HUnmQ0IDmHX+WJZPW8
8jYD9wMu+hALy4CC+62EYNeRn5EPfS2/W9S2RfglsE66ZtUXHxFQKHgdIsO9snquc5fOG24oMXBs
eKGpkK/+enqLt2D5aqiey/nyC4IbBL/nWlvR2AR3HSW3j01bYuPT+ZnvxlwLxYzUEcCMnTsEeHm2
760qqhyHWfsP1kqPKjZYPkMa9BQdpZIYdJl2afKLK+hDBSPFvsVNl44qvRWK0w4rujpMWFwWAA9g
Q1fvvvrjUeFLFN/AbpixA94dj3x/gWJf324/1mM7PnWSTEDqQBnDRxA4ZGO1evSkqa8y2qbdDnIu
HlqAR10e5GHkjXh5dAGUALs+hqAsnrv5c7jAn3Ria+FGWOevhqZENI6lp0laNYaDHSiO2viZQuYM
fFR0Oqz1gX/IZRXgrTcFa5POKr+cANYRxAB5X15FJxbb1PgZV0+KuPBzKKD5+ib2ec9s+BzkExZR
SVCVtXPDFnCXzTP8hFbXPFH+EYKUEH6BG6rwS6fUr3vBXzTSORr+nSN2GTJHFMi7F3E2oMJJzMru
ATtjMmNIvhE0wbCObrydGtaJXpSQJGAA7b4rYAjXF/nnpCSbwGQ4Ko5u0MlddmigERIupBh4e0rS
WBFSfZLll++eBRt2pbglS3yFZDQCLRNyNnCqreuWZuK1ACCghkxYqs3zNLIJQ4l7RbJ9cJ5A5ie3
67bD4rWhtdO9q8ogkHqX5vgEC5w8CDiafiAStR2kVsimkUp+q9kpUPmGl6s5QXAk76HJhlIWzT9P
7eq/AFs7ibnNFmzvVOPHwZY6UopxemklQ3GoDgAxu5ZdbIihKNjVr8OlKV63DNlNQc1Em8hdHCe9
ulq8Tvmduxq8iCc+FSF0i33HlhRkAn7U4OkKBqTBqM+8c96YeOioi/fPs17mOH4vIs6mTqyNCJ/V
UlBf/wAPF4Z8N6TOSOVlBiT3S0Bxf/cWKz+7OatU56GcUJLqTt7iesNhxnghleD4e1mgmp6lV1r7
wSWemezIwj83qfGPwTLTff3S+uO/Tq5ngYx0ys6+3VBdI1yN2TYD12gDYCPDkiKSA2jWYP1mhzmY
D7qM78L+Fo1iH+UxqWdc/6e7y8fB9Ubzai/lW1vLZLBLx8dpsR54FXTe/OSfDWaz9U1+XYRiF+zn
ynzmMkSl2SUV3LfPzQzwLcYDfviHnXAtNAJ3atf/jTgbz6vBXwBywHwoBm7be6pZhImqcwbI6+kr
nnOOsahbLS3i2QfJXkXsf5Zf5Eceu1upI0BKyUS6Ki4QGx71pEy+RwPcQDVG1iad23GnUSKBV20j
53FTe5angkImN5nBCuNyjXZezOWNKPOIG7IPEXxff/kitPn094ruJayJtLaxSVsRTkCp/5roy2z5
jPwSKSJURJ6E/BHqiKYdSkhJ+93+1PsgKLRDM/GxulGt+wsjDmrPVwiDZ60AsK08agnmo61/iys6
AkW1AY3qjC+EECh3l/pBD5olEcsL2gFFwOVpfubDAKKDovyj8yKYnd/l0XH+ZCBWWfDRlwaGL/Rw
j/sE1RCwpkvCTZ7Y1BJSYewR9986BQp4Als6ZT/VftYpldSZNG69zFUEhrBFWGPO0mWWinjha41w
G02+SUvqaqcyID5FLsstKEKHb50YTYlBOlsk7gya3TAhxzCdM90W6o8J8l5ro173xhmlWgoqXiIP
OzkWKoK8o5huef92+riXmUJXE+eF6vhPZQKy05hdP/sWLfCdbpC9p52s7xHStuIanUrBdl6CyP6Y
fH446N9fvzBwCLWeitF2oyy76D5qWMZRTkSiOWQtXL15D5OJ4tabxkgnYKmlHIv0F+LJ3lA0+3dU
A0FGRYYgaCX/UOagumVCZroZi+S759tSEJK4Yl9t3VyVeZk9nc2Zw3Bk+o2Tj0abXDQ3MS1EWbrz
ZOFTjBnRDCaOKN6D7uGUqgluON2hhJ+dF47eRYv/9v8LuEGJzgM0RtDQWxXgV1OoiwXpa+OKekeG
Jwyan2CAAhd7OUt+HKdOPsQXCUa/miVsJ2Tms6VwesTJIx9Qd+dWfb5TkQTzcGu2aUOTwrHFTCFy
DtG8eXyJQc5GwltHKYFGzPQmgwIrZu1v+sb3kz2zX0W+jiu1+hADuoecm8SmtYAGE9uqmrTXyXNC
GO9yaxSEUQud4PS110aMcNbVJl/jiACH2RO3trDRg9fQBkpTzrkxJnckDveDq8qfrRzmyLvE6Ed6
3KtnKR4XJiaSomoHr7lOxWe1YN4NdTeOswsDP0RQ3Jne/g4GnB1aF55V3Y3KV3l7oHil+qRQq8v5
kpVpjpFiIeiFxaRwMa13jFuqb7zICM3mm//eOHTgvOOVrCr0PKU0pgGXTYjMv/t6Z2wuDhdsdiEl
cr5b66HYfD1HrCmo1kRPhM4x+ytdlfeQy4V8iy1JkBeR4wG/FO3uDMw59vKsxHFN/QEoaP5sDjZG
EKXGS1WIpZwi2iKfBYZOZ9ukhByXNA0FjwNv2p4DfrCzUHx8YyUx0cr4+yQu4KuPcY3jMPMiTgAm
dXKy+lPPm5eeQEwdDKxfchjRhN8Y+BKrFhtnKQkO/1OzfBOwsl/AquBPvWOy19Kb6RH/g68YNk8K
UREJpuKGhXp3JXQU0rZ+efVaQOK0DRWTqEGLO/DO3l33a+ELdhnbVCDZbYVP3Uxmg+7oHGqrUc8i
/tOCj8zPj8H8EF/JKYPGFke5510+FZcr/YW8fZ+F1u3Dmjjbp3E802Vu2shiKOplLe/KCalGmoqM
f3XFS+AGdBuqo33v0TsGK0WKFZMvBKiBNgtl1bPlA+Zw4XG6jq5ddLfGhBbr+OiOMn0TeSN/e/cz
3mN++d/H3m3pzD5WCsGwmsgYCJ9TRg4gpqPKaJBScjEWgFX+S7BEytQU3oW0lpYKaXjvq4sGnxPM
pgJtcdyX/lKbiM63eMao6bsGH2yXcaVcgBHEjd0Mizomp5dNeBIMqkW+F8KrRqDr33i3ZA+lqdzI
idHNaevKeQ9noBPuO+l9hxEjxbJtWnAr0vy2O0quIlXwm5Qys4p2aPk867pyhiXo8mGT7y7Q+oQd
gv//mryVt+bNnPHm5rEnlnbCKAxxvoCtuWkAsqNFrzSoX8rUTBVX9Nmf2fjzFkwdw9tr3gXCRQpc
oMdrk5sH+l6O7M0KtuqYI7w5xHdIQdcjv7fYH5svJTlr5DyRtgUUTgETMnOWpfoSnRcyOmOe1b4b
e4cQkUEfaryoOllLdLAkAoj1uuKRvUAyeWnJMGggcwoNekUj93D/PsDAAThG2Wh9C7GHLELBKIii
GmSu5k96DRiTaT+mdyICzuW/zk/poICZ36rCB9tGrX3X3cPXUqOWP8XSmR3BSRViqCR05JsqL3u4
hkxAgGoV100LiADr8w9EWtZlLjNhbIDEljvEFp4O9qGo+T5wKgz9kc43ThCjxr8dOQYdjOg+/bJx
0RLzJYmjC79lb3XYuK3vjc8SMxzGzQwZ1MOIPRmS/8xHQj+m6npTq4QY/XiKFpOQm/Oxs8LlYg/h
vHLrwpdf7jKTh6kw2av7r8wAZFPCMVlAYyEXs8rZAfow//+rNjdbNXYF/zEqVI3n/klEEIIfnslQ
C/abcGGJnkJ5a1RiXL9CELV7ZxX/QK+v2PvytlQxYKXLC7GOqAwpyE04gDJ6qTQozJuDJ2C6/3fh
XpErC83QBI8/0lulHFrmB3prrq7rGSJQVVhA0G2BKYZiwHTWb+RsRWGayLCpC5GSfoA+05NN49Mo
8961ywaAHw1CMWKi84nfxIGWUVV8QrCVeEjl+TxgIPOEUdoFJ7G7Y3D4TXq7FJcT49Tn/+JYTP6U
XnIWbmcZH52zsqpazBdrTPjeFsKUu8WxuFr74MWCg+IatVLyNYdvj2XpebE5ayB7esYpMQP6SSq0
qXTlOE6wira3ektIJ3PHOKPktwsGKcBL1U5qcyY8djlD4Uvx5oLNAq81XiwuAUTQOXMZ+unH13nC
psloWVtmomUBItBtvhQ6PFRKZ5ZV+vvpI0PUCdrz7ueYGNV9aeo8WyIjC03/swBEi1T+KJIHd4CY
55JVQw1K1STPyoMnIZNGFOzzVrBJJHcC4A1H/gF2msiFGRe2+ZMLY9HORyvB4D0WxMTlwZaTkn2z
J9W9KzIGMWRurKtMXVlq5DRkJFmOfyt9NNi4+I9a+pVL6pE4gP2ezn4wag5PohZKNMlIoKF09f+a
JmPLkAb+bG8eyp6AZ/2UZYcewA4UoEO4uGJlHNoIy/N+0abUd3dh7nZ8O6Lu7Unc0XeKZbCvipGB
lR79W0EBE3uj3FOtoJO1kzWugcAD9TtrGMW25Sa6xMyQRd/HhSWbi5mE3G3GKpgrw3zZy9Vyg7bq
gYObXRRFE27i3JUqC70jZ94Ko+S7CEbmfYj3sIRxm1LZ69HtahgNxzd4rRK/VjufRN5evqQj88us
hrUCjYvg6y6PW/7dtmt5V011WG/nLYUnHRZOu9cYiNaq4JRAKPuJ5Uuf8TH5ciQ1eVfb8VqpXalr
Fg9CDkQhEihyORwIvAkYfutrh03rJ53B03kQtIkbhMRBFJJ6jHjyKK5DSRh5qVJ/gYYMkqzv/BCM
3ULwQALD/s5ofi1aQE+epGHTp5lkrw0otFUkxCk3U/SZKxOsU99LuhZ+PTzCyOJoomHgAmxxSnIW
txy4UsbcqFfeG+XivYhVMV98Gd+Lye0VblErw4x31tUzU8ga0WzRQLUAVji6TjepSq3eMOVcKMeC
Zuz8vUbunpVc16hSgee5IIEMjKWoorRU9L3UIBZ49xHZuTkcQQ/LvxvfoXElxonQQdiL47CiHaCl
Al7HRDcK60C58IrkIewJcPxVDc9eZI31TBxh9EKfoHKgicochjhoyX0y/rYArtt5E8XJU74Gintb
NlXl3jzTayBc9DKTvtjsUPOu0423p+abZoqpUaPgKAV3LQBuGzF0rlg1YZo9OSrqNpwJHI+qxCNR
rn7C1Y2ZieMg6RRET9z9MpnDGyH0T1IiHVCvMG5FSOHRxHHmfjgRfPV1ycGVEHa5vVWW4FBMLqsj
gMC98H/g3HXD1jTRNkJJH1qA83IRGjwPC3rXzRlxAwXxlmitegv3oWi2gZkFTHUZnRLvZ0YYU6Ay
L35BQaprrgBmNG+lwDhpg+E4P/q1J01boRC3qL4oBt8W23/iw20A5kSne7xqz9MaRZsVgU2sa8GK
iPrYfzmHLfuCS/0rxx/eIXWFBcMIvRkLC7CdD6Hzy073U1CMJc+y8xZG8g9Offw3LtV6XYBY6ASs
isdI/dun8CSwTyvIenN/0WHqriStPLKqq6HP940oVSlUfSbVtk7tyLEu3TEyO+kMGrw6FeJ+jhNz
YGyUm+xqz6fzco0OyqPxEOYiJYJmNXA9cpqHcqyWJe9Ca5JORXeHPF6O5RpFxYyI6H9JM9lqne3b
Et6tcTlf9aPCHtQ8wXG9ABK+/Q4TDzmltkc4x+aYeVoJMU+FtwvYdP2K2BWs5IPY0gmNgIX6dkna
Z4nGr7i3O5OzKNWAufxMvX/dA7JCpXNgrvaA0egzGCKE7it9MpoDZ7Un6JVW/K2HYBF9KQzwQwjr
4VEDz+sCGi9nN60vYVT8mi2Dg0PGUSmw7g8zbqHjmRZvJOnFwy36GJrWDlw/SxT55mbAE6KJv3OO
zz5w4aqK73Veiik320nJzQGi1nhgSVFBSOYhr+6nAZaB8n73uavWjgLsdAZ8ezZmCD8XIK/UiYxx
rTmnz9s0WYj0bWmxN3DYQWOp3ebcMMIIvBWWfJoahgY1yPixgT3jKF2X/5xAf6CognrDLLmKf9IH
1OWAGvOqT+2Yxxat7KoabAIvh4co79Pj528oCahysN1Ldh9vTImr7dnsWfiPxFpN8kv9HTqEKS/m
2N1fFaeppGQt5eHbkiGPSARdFLeKOm601c10i4JRc4j2y/stTApHpQSnCJLb0UgAfnHdEaKk8Uhv
T8HpDX5fllJSMUfxQsfMPomWnfhTrw7jlzpbMz682CkXbVoAuY27r0IoDXPh4U8js8JHsU6YkUql
PPHYhxECwce0RRO3fEzuj/k7Wj+aYCbzq+nXlQhTp6heTjsOLRyPARIKQis+uUQYzAqmyDi+ElSd
IkkuzR6QjQjnKvplYyxTnpQFhpE2EFrZsmcy/aZa9BQuEfHXwv9lYX//KXOiNl7WGJBp8gUh5rtu
vzCMBRIa4+mdHIHEHoukaUBaMRkeGV22xBflpY8xgI3lD9JUEhTglRDAoCeUFnKx/pskiK19M+XH
0CVkI9TDBN3/N37AjGgOuatVcICMvvzwAYyn8odTVw4yfUHSkpSrEmUtSQ/EfKE3lX+0piMF1tg4
Z7JzSUZuby9o4yRcH13ydUYWNlzxIcU7Jgs/Xc69ZoHPn2J6BvWhyX6l8m8jwi/Y4Xp9gzX5eWIa
DJRpyN7HMGtQtA4mG1v+8A062SEVp5Wl8PVAc4WPqahwmvVhxm5UqVpIrN3guF+ZRpu/KTHRiovg
05lkUHtz2/LBU4JZdqzySM7h5C5Z9S2JM4VMXdQ1zvrySi6bGuN82XylZaX6gDOuoNuMjOo5qIkp
fMUACS0VNzITneSmr1kitUjyra0rG7PldUZs3i8XzFF+qUmHV0exShTXAk/DcdeN+Y/EGWluie7z
CQnvrKIo40/3fWdVUv+qyvDpqfHR9tw1nACWPAL2GDrgtABFZLGBgqO2ESsZKtRnDGokvRmWF5by
yS2wUxFqN370YnB27mp8pPC1AjsQvpkg51lUadAcPm/O68ZRQRk5SpsJiCsWnyWABIOm84UjWcop
+UjyWjvKRN85J91AquYkiwtG6G1MIqq6EJlk8VEK9LoKyD53boLHh1ySQYDgqFBtVnE8LRPQtbr9
6dK78VtPuUiU+0RJqOT+ugOMIJnHRIaewYSB7vqTMcl6SG7lqcpz9cVi8ved5Zz7SW2t/lS2Pom3
X/ao4f/uz0JYpIdcpcgaFEzTMlV13+QWyyPh4HYyC5btU9I/RQy8YRGjB2P4Q6ULeUkknIQuRNq0
3ij7YG9TcdKzYDQ3IgozwGRgTRpHQMem2jcF1fmuibL6CjycWGeZ0WKbc5zvMB9/O8vPBYDAIkE6
M1Gs0SUS6mfwmx/ZJHs8ga/XOIWRCGDvZbLhba9x2gulaG2KxQ3NSkqG4vdTRuk+kKHgEWc08p/X
9113KTuPU1eFSNuFGeWyIln//Wf1XI69Q0t5Fjj8gKwyR/gu6k+CLvCC13HkSkLV7dR42YBrQJv3
bfdLL8h1e2nSfG2k9GtJql/Yc2Py3LpkRWdq8/OdwMKUviThPh9ca2PM6pUkSiOblv4QY0h0tfwD
YgJ3lZKmp57+qMrMF6G6hRpohxWogtpNohwcnaFri7bmxDiMUZ1kdBdPnDzrMJhjBBgoOv2ASUnb
HoYIGN7nurPLiqn9BvCTnxHlyoTZ+swFIdHeAS8NOp/+YJJl9+7KX+KRMNipegire+Z31qh7/3Mr
F1e7aDb3bHWkWSpvv60UZxriLNaM/gm9o//mTKGVheAs9Y2PQHUhMUGnzT/uUiBt9UIRu+cGq6h2
iCAv+z8gzKFFGRoqlMJnVNrVxJ3wTkAfLsZA7R+0XnRkulgFAUHHN1jLBMBOhYfbOYF+rhAE2ktG
uhIl5wO6mieYt33jzpnuN+9HDAkRSmRXdOBwcnziYlybMSZcS/V5RwYDDzuTygSNWHQ5t6X3iYE0
7IDMwvNgrfwv+oCVp/TXC0wbod6tO0CP+gRR1iguvo6GzuEwXFzYuRIn19J4wl2Jn9BFGPHGqiNb
oB60pe/F16kBSEvGgbJk83NLmGZV8l+Xwwhr2xo+FZfV0Suz3dkohCvzA1CFZxtNSgp1h9qoCPWN
swARArY1LygVSfmWFhUEu4yNXlTOjJKOXoIrF2qaiq+6Y1uhV94+yLA4L3+FpQZCRsPj/t1BUgvm
iu46O0FZVxZdt+uqJzZd3zi3rO8wVIFOMwD78ND3uWaKvvtdNIY5lz8JdJmj4Cb8qZEpDc4CXTWx
c81MN/om871hNtc40oLNF1g9kCkCMeL86b9aOOVzWYhKrGf2jU+g0bzdnttkDPoJhABGScom+LYh
7g+/aWgfWlUTUEWg8NZajq7wGWkxjh5LPOQCngjf81ZZnXAPJu24y86oGdVxen8/WTr7Ke0jh4ek
FdH+LeMW79V9UHLHnMf3w8Zn5zbE5zCKUO73+eORgi6LtpcMa8WWxHFNmSFLrVMv3y52vvkum+TP
u5Mf2/bbFPT+0giluXJLp/tBhezKYbH/Z3/6MfJ9yYQ4bJAJqwucsrINyWlB2r21iXNhZyvI6Zjd
j25tsa9ngDtwMoO3aq89BrkboTKSrGEwaH3zNAMih/ScWr5rxmv9jOYe3FS7m+5uKKuWb7Oy1jU5
IhUv0Go0WhLtpPpIcOF0B53maUScqSv0seFJrKi7vU1hcDtXPMBUObiRDFCfPQY9kT1getCbZiNR
84NsS/eFqgxaOrCeyeOVAjeSiRZ/ioVOCv5prXminAHY6ZTWqmvi+7if0HfjvX3Speq5bAtCFub4
3IgXnPkSw2mAyxOfvOJzwIEajc5udYhJXBC10v1509Tpfx4IkW4BHtxrAvaKCy/KTN9O+r2HFjy8
zK8wm9CODRfC1qBz4WYHDlYuVRsVnzM5pHe3yDbbfV59uAm+So+xamP4GKlBS5DIYsL1uzVXQtMY
qtjMk2bg1UKWkNBpebsX8SDzv6/5s9CPK+ELmmf+PhfKorqvYdugsnQUbLlLK2Lae67cHGrTV/op
Wm3V3otMzU8pkxFc0L6cecaEJuhssOL/6I3+jtIWzTj70PNlSukQgQwuAuxqLh9Q7VXW4K8ZYk5Z
po72vIe1mr7BeHhy+7HrKtx7cjSJPvjC1YwMk+9tnZYnK1pZJ9zVpvcBCLPlG/1+aWp/xtm2IR/i
v3YavIC2n5nWonCqzLqDM5XOMlf9dldGq0Mq27odwIqG+9o2c56k6d1FuHgFdWv1tfKbbUewsugZ
tU1j8q/uCAOyq475wTTNnb5YydOVdi1/OKAUwxoaESx4Iv4BOoqFNa4HMrbxiRG/7APNYG80aDLe
pzcGGGOyqS0ASrX+MDGG0Xk4grQ9OJoWer2edTNtxsj7jAZhKhAhyFjrP8jo77nW1cVuvjNEMTuj
qUkx+Yq6PU59Dw51flhUOyvWkVHZumfcozQ1WYA4364IkO42w+De0n1PAbYGbQNFkcGD3P5gkczr
IEM4Yj9hZmXvN0LZlnwlWrpA8O9k0Zhvc3bxu7b6F57m5g9c2HR+aRXztfAP4jmH03rY7MrEpyIE
xArpe6QjMNnhvR30qMiEWg1WDxTl92uzvqlNkC350949t9uwxsNYiiOQzCcPAriqRV330pYqWbJh
6EbCIuTEhGyxDx4wnsPHroDN/fizllTAuNY/UQkNWvPqFPNm1XzrbglvafKa9Z8yuvyR/3qi8U3v
xK91Z8xpWmXJ9IPRGY5fVmcYGV7GW34b6Y34AF9toJNzILWQIbEE7fMTSN3yLn3RctzeV7CKGs1V
uuEmRFTyikEar3R38/eO/NBu72s2qmoAPomifFk10U+DNrNHBDf21TUbN3PslWiV56wcf4LUVmTO
aDTDJOnaCX1DDBhI6URS6Om9P6rozixCw+kD84mvD4/ta4/AMxHJVV6n7+U+J0NzWKHx24Ewncm4
FqsJeoSFYi/I/MDwEQ+jGpAYezNG53dWDIw4ZHgrAndUH7mqxID8yzDftQo9pTOmsjguutxrb3b8
ZO1u1gQ6I3z5wqZqhreS3bQnniti6B7eAtCQhiv/aWCbUIQwBEDZTEdVIaDMwOveb1a6PfWVXceg
DCb7iNr78nYTWH4Dl7AcZj1K/JzmZuoQE/lDWfo7EXaVJxtzJJiDSClXjoScxJInDHRlDNMY/crn
FJ7YvXxwDe40le84dr0RFGaIHkxxD5hS/3d8++Y/1vWmduo3bpNHH34xQF56Nya+YDKkSz6qqD0c
dBj1NkvRwqHMCKfJvX8EUOjuZGQxRZQFjMgpaRdPCcYbCz3YqnKE/xASfKSRECUTMgfNRZ6/Qfzq
abPP/7lfiKACdzlvukDVf5vr0eO8Bf3oKfvbN0hw9lLsPyztiIZ780VH2OsKfSBJadS+W7fstNfc
0MlWY4EV6IV8lNvpbnEnbtJxx7B8t5Vz6UEmTOIXitYcdGixjjzaGFqXFR7aMg6QlziOqRWTnnj+
L15dn1mE3UGNaXqvjHUIiHx1DC901UVZghTyTtmcWH+6GfUyY5+/SncIGPZ2h40Y16wYHKPLpkiI
d7XU5MRLfoJARWpS4Ap0YKYLtzGC3xcwyGeNxtb09xC7whDqJ+uIGSGJytvBrCeVopZOe9Wj3Wic
YZeqrILKmA77BMkAZPHcXv1BreTJ1sA7nWFkxt8u1U0oMWxLqdRoVHl5gkFxFisTx7JOqnrLrTwS
44htKGBDF4lyQoxzenPU6caVOJ2jHHyd+IwdpD+z5jIh3iy9XeI9KCJHue8Yzu7Eux5fzlgewPl5
wVQEDYHVyKAMmX5WbDKSwOkzxo7qC1lWYKgKLYM41bLcZlvqNES9rMShrm+bzRUQhdTCAavEFF0L
6i917XI1EIVxA+LQVkq3D4CuXdr20UfPM9DDW6dm+LZwN0ZoSR7U6vSDOBYCw1Y+gteDV/BOkDaN
nDdQOgoUXCQy6kVgPMfoT0hdnTG/I/dcfmO1ESp85UddwulOZ7yJqERnryM1FmRq4hwtdw76GVY0
ciWQSxbtUREPs88JoRYCU+Q3lmKOwX3WKx2HagyZPIR6vphOOFcXjzNGKFB/cwyzc1gnXXO1VJWY
jY4q1hkKtvKhRj4TDaG6mab8b3tiY9wdnyMqm015iYkcLn+ojJzN1q92IxDDrix3HptA+bowVEj0
ron1Gq4kZ42S5ixyAU0U7LVID0rJFOj1/9kk+QBxcgNKg8P0nt6jd6OecxjSFyUF3Lc6QJP5c1Jl
KhsBN3Sdwfk6AAr6S/YWJPFqbTJiw45vTKJgOwfztLTRWjTNFLWqF0jMFgMKZJknpwrvLaB0b2zo
ouCDmDCI6Dy4df46r9Ym8RQPdSTIZ+/ax3bFZJ5eHuYkWVp8/wiQwanWtPQt+56bfckiuB3ygVxO
dk+jUC+s8LHnSGSewEzYomn283Si9Gm7SxQ9pqpwbTfvdBB7LF4LTeS8YZ3gsz6Nbdqi596PUrrr
N+xdJhlmZyeAJ7r5AUqDxShUOMTR15hRuekgpkjhjz0ayNz0Mzm0lAjqLvenSHGPxz/xobZvfsiX
0hLWD0YlMVRgokgM2zShYaAvBw2CKw+K6ziFjj/EbfTh8wVcJBCOixQJKbtk3dPoP8YGTlRW6mu+
Krgo2yyP0YnpE35DgenljGp+kLt8M34F29EwJV5/aCGrXVqoQ21mb/g0kw5+FvivCd8xtJBMjwjr
eay1slAV5kav//BpFmES5PBPXJfk9f2jEowJSAkGifyC+iV3hf1Q7mH/zNbLEPqzgYYrJwmoa8Lw
oVp9aBuJfg9+NSXZeL5zAMUfcMJl3lQGuSzz5DKIxkXjYwzy+e4nF9dvycvTWVHp2kWumqqfMVFR
MMbFJ8mAHhMg0ELsEmcSq0mDKx2sMsBXqYWbOiUdgffFYzB3JRAvWxxerQtr3x7G/2e3yTXwPoIY
K8Wu6hEPj3ePVRUq1P90O/4YNAPw8MioK5EWYBpuzau8ECrzV6taio6D75Q5JvldiSo6oPPXdFb4
eeWMoDgoyuiTyUgsYjbWCg3oFyV+5oxC2znISPReC/EzmtQknvXn/stsj2xEegbgfYPqIon7Et+o
fWdRtJ8gCjw988iXX7DKyGgbwT/rtTZOGcU/nKvN+bknMoICnEzsPKezMjHBTKNA+yY1mR44Lywj
tw8KjpIXiefE+tfU82Sq8iluuELxnwT541Lv1EkeCRz5sx1+VB7ZRikLMiy+eiBasQNxckThRYiE
icJKjD+63NjXYj+jvs+KSfzKoQAZiqM8+APIAubdAeG+Ux1ErMmV/xiGBM8Rf9Yg4q6rdSVV7UIu
Gz3s6evYfjHuIQ8Y2Rsr2UzGv3qyfKdsEF6OkjGMX11bcthKQO0knNMzJjRzijJNejFbqJBXdDny
x5D8kJk7LorSKNv2V0mnTx1wKKsL/ZfEyBMJfOY1/rbY85hZ8ZcCjsQ0J7nFjXHieTza+Xuq5+iU
dDj/2Z7wePyXg0iCxn34LSM/XzsNuTavvUlt9a339Olo21Z5QVBbxpjDaYPJqKAyFooIbW+vVRWw
IsP2lqvAc8pyFDBhUTs3NxWy7mGZDWamn/hErIYRfhaL3ldLkNdnHLK3ZbqrBpe59PW7Jg2BGXVy
mJJMjmM2Mv70w3ZxEqTtpTTfQrYWij6oU5bJsnig7x3rlZHMjY6nk7YL+bAv8nhsFbwUA8WLxXAB
ozIq3i+auCYQYsVg7oSK1le/MLHtAhsxeiDOK3BZ4e4MePGk6Z5C1usLhXCLf14z9tpK6ahalpaX
5+IqHX6WLoVI576eVSsAai15bTHtMiAtwrqnqqiapWqTmZ+L4Hi1AtVSCKBXpKyakGgjS0WweZ0z
3IQEhJEYLODWEcJ5rGVzPQbLBB8VMfRoUWS17v8yjjs8e/Ozhp7dOkLX8ulygcaBaB8oHFxUD6xi
nLJamsrqtYCOp9GFK4VFD+HFzOq6FI0WLfQ0pjX8lxRYzqBVqIpgIwTlaeZmDi1RWRZANayWY1Uw
4RTNaVmU1se9EJxbomVO9A9XinvCNt2OlS+lRoJOL5ZsQpG/4iAeEbcS8wCeic1AzRRIBHE95XhS
jLekHfAT4qxP9ulIU3SxRF4X/DGx5oxb0JrnHBkiulp0vVyBxF/9u5AUVD2nXtTrSv2kTCgw2iHR
0b8PG1pVaedpjwRIRrNYRd5uUMxkwJawQL92wJEA6FhYZqaOu4a9MsJLWHm6DMWBW9arTlzCejWQ
54EmCQWgtA0lcNGWYnSXxcPwmSy1/+P2s+KjxeCBAM2m4cuNnWIal/WA7YxKHVLrERw/ssP16Jow
+tqFPbw0G3kWvHXqfujM819nIBYq4nUP5xK8akf5X0YgTmUxN70HhdU6dbBauDXfkwPRwcrWvqcy
f7FPtz0cm87iqk93rum5hTWqyCnJzc/OzYEjkh4cjolIeZl8QCjJmf5fr/RsH/rAgB74pnt0DnGR
UKtaJ7mPPg+gXFRGxyfwhJUp45lKEX56Gw5ZW54FXBI19mnvnOzUCtjQQYZDr/vv/xf3QOwJfq2k
MzaLMn9fD+jrPE3w76tj6vgZWVcrNFBvo2m8PxPT6yh8j83C+DGxzQfgJd/EB2LdqwZr+JbENiIM
cwVNbG/G1WoIcXGiFMKwEtKFR72kQMO32SCpSPI2zujH9i/uyQb5hBEUJN2EhnBSQC/fIs9XIocX
DojL1yiIn6wkIA4UvHFSoeJ+RDWGvgYryLDf65yPhs1Y53KxknrsEiNg8K/xi+V3twVJzVn059wm
VTIhJUzh0DOIlTV8bahJ25XY87UNzRk55dkngafkG+cBrhVzUAh5uXFWxWae3xKQ0akLyLF+WidT
SXuwTrlk01yoKr2LTG5BpCQTbbOen7JKJFFiH7P8GBNOd20ERfrBtXLxse2DdSbU7p+vBqJEEHIl
eEoNONhhzO2AIGzOR0znMxeB3SpUWrNf2nNWbUKf/T14sYLUy9Hr75S5q1uHzc1jknZtK8h/AdU/
ymFYG2+5EEA0WUs+HKKtj/sNX8LLDy1Qy1k4mRF9OtiU0/ePu8XGTEnqU4nM3SCruD73sN9mDVvu
PHRzM2BS3AaoNf1ouYqEKCARMiFVSx/Im8dvD+729BO7UTtDfxn09G5HOcKEJdIE6UlU1EV5y/K0
+qroskDdMyg2uZfxG5cDAOIeNtoHl+4vSuKh8K2zF+uixJBlmPrITZXl/6By4eS5I45q92/KBWmn
Tq1ela16T6w5PGrbNM8erx/83u4WK4/Ee+mMoNlV4MbWfYDGCaKLG4tUIqv7bSPt9kMWoR/V8KyK
kQLmG63rBUt7kG4NdNC5WC6VNkSvazl8dhySrAByWImbXrqWElSsweWma2GV2w893LSxWrLMWmqX
GVRSRg9TZJmudTsQaBTkq9ERrZlG4Y8R3zLnt3TGRVO4Ph+HG4SP+c8f7cy+fxIAXQ3O9NvXe0wx
uhjU2vHP0NWd2ZTmnDKN5SWddNRhV3CzRxrXHNFE8dLVJQuaKqq+8iz6/TKtLv1hxieay6n4L0YF
UJH3nsF69qtEWEk8h7lU66ltzrPInU+RhX7CrSxyBtwU85s73z6vYD687ergACKvBTJLDLXl9JVd
S7KLxPB2efsPo+pCno4JTg/kDFaoE8Ld8z0STE8IeQQMH+rk0Ogyp7eiaCJfMUPsATYV51NMU+w7
lKEwE7B7lxTORm+XGivMpmhMq4jPjkr1gzUPO0xrVRuQtcbVwK+sAMyT+G7IFFW1kOqbitC/nbVX
v7tUvWUTnnDujQngIl5ViwJmbOq41L0w2TU4vSvTj+B8KE6+7plSs8s3+RJhid9J/nj3zz3VD5Vs
vI1XL8322JHcirqGc4z0lfHu0Uks97fP90cNyQM+8GqPIsos0R95+JzBP/qUaPe1UgGFSvWJzwma
vmXYg6IsobAZk892EvNASNzdDGy2Aob5ps1hl0Jy7rY3ERWKACMGRoiDMcU5w7BgICh4HxYvX+SF
LO5xKgrsfH4WpszWOAmFSu/8TWGLzRFcEagX0ImE5SQd9+lkUQ7O7+2AXCJbfaE3S9YP+6uJ9tFs
HBs37gVsZi1sjy6irSd89boa4by5KGXNHQMlCVjir5VmK7IEH1FE8blcFPFwog7gpG7jHFqx+oMO
IBewk9JvNJx+pCdSCiNeS4wW/UXJAcwv3a4Rpzt1cfw55LiG45723oCvETY7RDswTUD7iKMCl5k3
4xXwN4BS1n+HQdynfwOEOEKHDPxXQd7LkOtchbAJxEU1dGHV/+SPg5+YHWYA6AZGpbCgyCGlxihj
GdmHQMeQRclA4SCQVoQ9uldZkSdnTqdajd8x5eG3dt8+jdr4TqsD1R/wdOKfpg5tysRNgLm7lksY
JHO1kisA0Z8GakR7VKNRuELwO+WS0KwiHsRgptNMI5wbWDkQ6qlcKZstw+wKUX7ojlS7neOPIguW
DbQkh3geTTJXWe+bJjOqsiTO7ziezeZxOOjCVNYuJRsfBj/brKSBmfPboMSWW0zgjH4J4+lzHaOJ
gGw63cIClwRkcnI8uLkagVJOulKOWZZyy/gRZFVJRI7qChxqtU+aBYhsDnkeExkysZrjhIGt4yss
MTBj/bo+4gm0+1T6ucaVQDEP1WdwGFEd6/69RPdSKLdu8Jm1dBKHU23bRSMLhcaRaWDTDJDVGWPI
3/028ipXMReeZigiXSzOLvN8jCmS7BNLJwE0s+oqtxMZAY7KKuxk9usQho+Y3FRmXAGTAbfUPSyP
LP/8lg2oxgEHR8yVgENuG3iH7XUUDcpwE0kYCuSGauCnPNQiS68WIdYNZuXZzsAkWHKFx72SFrfj
8QBOJy6TqgeImDZN+B6ls8UapwYfeujEiR1Qz1zeX1yVmGOsi23rsWUEf14aLDQ+lkEbmdey/tPG
oKADc691gtXeBuDEro38kqUeHlme9ndvLzEbE51drVpZZFs/gXodMUsgl/PkT/cjL73WsHVWEuFi
rBR/xEUR7pF0PiZrpXoankNzrGnKYouLIocx88ITqdR3eLFZV5AlRw/NapY7Mm31vCDQq9X/y234
hBWZMDmzb3PvWGqyyta3bKWIpO1rkb0c2SROqBifuCKTLN0ckzeKw+fY9SOLcYk45btfDpbcD2ci
UWX6ZFaFbAPAa8qYySHFDaniDnZqNTSmdFTEEs1+U+vBw28YrIQknzWcd4F4R6+0/bHRVFcNc7yQ
W1OAs1O4mE5iv0Fa6XjKuoD9g8KkcifJ/noW1NB9jJJh394iqjffCUIOiwPv7krAS9pNdUL/ZZKP
5Yk6Pkv8o7AJIbmV2Tm8Y9U69sIWBH56hkbKm/PCPB2N5kXPNEy7ylqvYEXou20qN5/uhO+nZ9+j
JguGmRnW+dYL+pPaFid2jDZRQw5bNmMobV4jkEGwLWRDuwRQuU1GP0P2Kky/KdQBmAMXO0ZVfTUW
Hdf31wmi2fz26OOxp3QGvY6eLMiZjCkFhNT9hEdYcdMDE78lzlqpV+W3Tet+gNCFrVSCiYPhW9XP
fOThn+cFaaO9jeOzP2te69XOjYuw1Wz1vM0TWTvs5Vds4Fc/y3weDs4tMp1l3Ww0JG50sZSlaqZe
JPMfv3TyrEM+pUklZLkMWFu214C3aCDjDB5+2N1unrLXO+kXobnWcQ5VmRGLutiP0Z3dC5UlKMxd
HvkKUzK2JhKjaVSogCJUfG6BiJOCE6M5pxSy2ZrClSsjpBNJtct2UkCYt0DriROUgbpYm14J3xJW
64r8HqGoPxgDKrgGCL/0FgDB47ih1X1Vkve+0bAPCgVFldKAWdnp8Edc3WqLcdHMdOblPuAvttSy
U/B10XQo54KXEAw/R7PDgUAFLBWBGUCpQOJV3ACT3ZbwUK/rhbLXNZTkz47Dpm8Lw7gm3mA6m+QM
ouxMqoSh0sKgPDGWHTTc3peGQupazX/5LUZajJzdoPAfTII+C1kuTIqBlZtQzZDW1ThSuGOLSGrs
RpnRx2Iq/39yXtveyRjDEroERpDatxCxwntDogRLTp2T+ffwP9gyUeO/8JwG/wqi2QKSe6OBdcwO
ehiGVRZKK9D6HS2C22g5WzTDrjQeFsVHqGk+VkjwbZ4r0/BLa8q5wYDlg8i0E7k0y3RyIvk2Cl9k
B436KsoJNvGew2ZIk2p/Aa5wCvjRI9+qeL41Fumkw+0A0FQFQasGtwOhaqg0h3MwvX3YMnPueXGm
zUjpg8OzYftnQEpNRVjW559oFM/oHfzj2/Cj2ulBBGJaViIkPbIusFwksWy2jrb6xrO6RlqtgWt2
nozDZHGq85tjMevkHbS+/NlfuwP68iwPVylHCgSeWPz6kSlA27b5dlJQ0jirrrOH+lcfud7C+dgo
a+OBXPAp+001esZVC32lPIxnYJhAJjEnL56vr41T2q3ltMovUig03HMcddV87KerkzJyKG8PnBal
dsH32Y8iRh6CbwtnnHJUM1Pge5JFQNYG/mLEbZ/2fGvaEJDatHw6oPnqhsh7VK6VjTCKLkOgwVv4
7nxBGpGkaXoHIaxkUOgWk+LJWU7yLXxEn1cQmGNPP5CJuC7OdFecDOp22Ua+7pXP1J5Joy6/4dGC
U4do6LqlfZ5z1YBFTlhaGsuFJQVtLtVLTNUSLeZEBKQHuOMWDSuOntQxgCsG46Pvi/gvZCt6Eg1e
OGTzJXHbNmAZ+Hb0gpuswYDRyT7DY7V0KKcw7JXFA1dvQfLzRVNIS0hFZ4ldXHhnZvfhtH5+o4lE
geCTXcMflYL9YZsnOXf+GVoHL5+9XJrhq4TX1lTJq0mPdby+GyTd8sgjPrUJnJnm4Dxq2g9SaWbV
irNQiCV0zWjT0s8oNS8qXtsqOTNiFmRbiaJeg45SqGcQvQI59Yc4wX4x3o7XeqFubDk0saKpAC01
w254xJPdjz16HVviIhu3u5onKSH1wliwb+a1BEhWR8RKULIRqNzQKGK0SGpQt8CzGdpWOZyg+fut
2asxH9Z438pvdkPbJmWCSp+cVtcexCqL8+cYsgAoSxTQ55PvsfyIpglnmztS4LsKJ/NLV+SRr8vw
xliOcuQSVDeTCZqXCyCyN7qlU+TOnI0tuBmmey7N2dFVFxsW9y9rcp8Ao41th0jzGCx4+uDAgMME
t1gY4RUbBxZQJlnIbR1ih1Qswz7LIJq/vVfAZ1/On4wB3RcD0dFd0VS1uIltmuKw8yVRHlXNYAho
NS19sEuZMtgkxjmRdVe+yBuF/Sk1Zc44B5PPLE03DLjgRU6RjvCZ1B0vdpVgSFEH9EBETBeEvtFO
F8IZsPdzmyXZ4m6CHedO0nG7/k3z/6nAfveCw1Oa5QUmjraDi5dLVaowRYieYqWkPb8fxzPaeTi+
+Rlg/OvbRUrnllnq1MN1JkmmTwWJlDGKdsGTBYQQCQX6x7/SMNqIqIGfCblYcCF7sziB35MtCGV6
bT7R4Y+2wsHjigc/e4UjFkF/Pg2nNJ1874EuSn2AO39iavNVFXteBgU2Jc4k2S8nvFfXxUrFM6bY
eOGs9wQwZm2Ghkszir/LvXtK5wCBePmbqxvuav0ZBJ39N6zm5fCN7nDj5mQFLgkKbytgOCzuZ9av
rfbo+QTfxGyolvTXRkIs7rZOdBlDAViLBgFZwLN91dzNqwlH7VtYTp6h/28IP+qNZ+lJ8aMwwQLo
8U/mKqcHJIvmLU0VSrb23wgIim/BBw8HGAThM4shKwylXPxh4PDofY00GZkDQ06eNSttDXGBYynA
dISzOnKmneFNeHoax7t7qdB0LV2oj57/mUAw+6U6+EiaAm7unTG+K1GvB5S+OhsnL/2Y/qqTYGMY
mP6+8CnvKIlBtvCbKuFu7v4lTavrJdz199/ECmTIo1X+g1zRcHZ1AYzLjXS0peKDdxWJLF9vixHg
KgHYHyOww+ngKv5pRIu2C2+ZyGJvKiLGcPwVb+e8i4cBv4TTGgY227pT34BGOiEPTbtY9lvbR9/1
TepcuckBkUc0cQLXRPb/rnjOuKOgfMwhxoy3DC9p+/b2kDN32FCK7sOAV547lXRW6ukgn4oY26Sd
+BjUn9DCIP+IAoz4ViDffNNLDjrmN/yuV3EVGGdMVvvjkGGGNJfPyd5ycCfANXDzkcjMAmX7y77J
QYCXEsZF0rK49fbelmNsd05waL3e1R6nlxz+uJEwt0Hbweu5wHt0oeWbBaFv9sLqNritnPkDQi2Z
S0q0niLAZVsNx/RkGqToLG6JZxPoliBLMeAKqWouDu5c9UmviLMxXhbXXvGCW0QV7w29x3sTwgsd
ptxJp0Nn88AVrVC3Ap/Z9M/rySdRbj9A/wVo3yKCYBTWmb+rMm2JxWJZLaKvi7mzA847D2fN7h/m
PqasVaPwvy4byuLJkHb+0nojRMJX2irxVr7Cj6prdeI9j8F0CJULVtPIYDIxB6Ap2UXv/2oF0nKu
CQeZTrS5iUAZ/rzUS0m0SjvBlrtgZEeBMFc+1tXAkf+7tR36diPcsowFEUp5mL5ZRGPkq7z8xZeS
rCZc1JuQ6z/OFD1jKAmrGYhoxnMLEhqN2vc2zbq+8uZMRfNzMz+fEbpA/SAQPl1hYZMpDVFhFGFu
1mXu5Y2EIrb6NBMVyHwGSL2iNT9kL8fyuXCsY90agJ/Dh6Rlx7LYX/TW1EJVZu/UXYtx8P4+HCJP
fVDwaYZo6Q1jQeNOphbDwud57/QX2TDzon/6H4Y9sEI3pPGtQIRWr/ZJrCbQwJoYxe3koSP6TC9b
byhZVyS4+HvrKrh3V2Q62VA1j9IsfSwHsJhSDJweqEtBVGLq0l7ln7wzqegxiAdxtw+AKIct5/xX
LtNz99w2teR38ePj7J2jEaBStIxfjYxwI1eWDAuc10waDF2kxvhXZb+BrAfIVqrY/6jak+Qn9yIu
FMTTtnkBPdUbQqZvnfBNIUMIXOUjaq4y3W+jO+eLtyLy//H0ST0NGY1rH3tl1kvpLGDcoW7frz3i
aQdy0QJe39DD4u5OeX4jzpgBFGsJ5KOmya9QDu1hoc4pr9SiromNhjiQb7JQYjTpZqFM4XbC7eO/
armHIlyWGaIszFGqqc4eygmwXyZ1qVkBS7InAXKAMeRIUpgqzuVVKtEOzinecVJaF04D0Ey4LSlz
/oYMu/+rXBz34pRJdj4ibjdKrSqafA4a0jrMkuf1EZ+5VC7u+FokGNvZw64McuPzw8R4Z1k9bHz8
pWkOThZ3ufJwWgqFJu8P0ixQeD3+Mwx9HrgalRPA3EdGKjlPgsV32ffm2bZqhsExh3IQbc/mPV9a
hKT40oQ4fxq8pLwIEkeWh4hp33DbW4STE2XYxXEHEslu9IGUuA4sYjXPyLpFDBdX65xLGU59p6kg
I/lFm2XpziuxubQcqokcVfsNndk50zhcvY156BjMh0Fm1Y4H0h3IJ3f29WUNEr0RE749RFOH2ca3
cnRCWGzZp2VmLvq3+S2QaeRaA8ebGXvjWzA7KQTPGLDQWua74ltSbs3p9rmPCNwCjxmL5GvkVMNh
7w6ufKLlhmT4NlN/a4xXK88CQO37tPh9nVZtDhDKjhYsEu/QTTxKsnSjPLaaS2pbSpb6vevyIosA
nod1ynt1BpcDQvUhrE0G5hBYN6/UlPRTIO+n+z5VTTy7F5WNfXCsbIi3+sOCZmpBW+DjNzeMvT5m
wz/UtofcRTd2hsW19ttf0mWXDgJLRETHF5GjjNuo99D3RQbUdzYuKm1Oaefqr8zx26/3vckyoiZQ
f5tynPqAX3BGHhR1oS5f4S+R2njAm9mBHgYCuP0uTuntn/RIYEHDFRvN1PTXJzAu+nil089v1iuu
1HGIaNxSYr/7nIsuq5tDltolPfsn4c5p6TyN+kTi4kzb3WAahdGlJwlw8IC0FKwBk8jg/4yH2iPC
0xt8HtPhpSNhiniqy1h69utGEQmB0XVbMw4RFrPXU7vInNS7gpykgKV5Ea4bxUaQXr+uYxaHJ76i
vcAbAKt6FJnBO+iCjeirXO+T07P/OyBWE+EFQuzWWQCqhRX9vls/wfY4EvpxAJzuUQVD+VBU/vyt
ZdtlUBPugHAjkzFnt7LaJoOnBt9Q2EvlWbCleXlWLf9qGHGp31X7AQO/gwQFD00MniMwVUcIlhfb
1b5etDCvdqICvBStGPWQ6xfcpYRy2jDnFj/9B/T1VCfFqtIVLDttCxh5T9e96rj7+OhvwJlN1zJG
4POu+Ccdax3tAbiIbyZ56/NykFoEo6VCCdeNup2+i/n3r37OxK716EWQIZZKj/gN+fuLn/Bp/LTn
i1SBt32a6hVY7AiWMHGm3vDzIKAN5ekFVmvmD9M1khkBaGtDIE9DWcqi45GVQKe/BNtuvYsDmWAN
GK0gHqX74qPLSKSs28wNcjgHsO0682lU4tigqCRP1yzFZ29qJn9CWjiOlgFvZN58ug6T9SIxq5GE
GojVnWRKY36CnB2J4N9NxIo7te2/x6hOIPK/nficfSUWRIhx7neNtGydmhj/6OXXbSSnuj8UpE/N
//qXfT+e7FTiPH76A4Dt4W15gduiuk5oY1/yDTSuUjdavu9Z9QolxBPGD3TQiqiSDBP5K5IJEpfT
9Sfv9GdMtL/gtuAX4AGOIu8yYepALHb62oQNWAsw9DfaPu8OI7n6dCiVCySTeFd1ZNkhVvZfMa/r
Uwt4UmPlfSfNdIQ5h0jlIu3gBf+V+Gc8Dwr8W5Go0xy5jPE2J1PAGJ83+Gsv8exBTQZGpwNRa8wY
Tr2o9x6Shl7XCm9HlZAciKdSMgkEylx+44tm7NnHe2fS0yhBpeFc1jFcdCG452dL1pUayKfGocj7
7QdfDb/lVy/YWUphd6MB6lYLbsfBfdTi48Q9aMg9neMP1R3wMk/WfD3teO6XOtVETGpU5YaARg8J
pbJxrLW5hue51PMOXBDH7T/ayaJJHn8fBeAGDyUGRxSH6/7yf0gx/zifznWe4bB3VAcX2LRgH3BW
ZIt4O6wvoI/1ITFE5gSUCMiO/JXgUucU+hwL693xv5lcO8MP/+uJV4wK9Wfze5WonfKq07couiGY
pFf8fuEy3bgG/dBvCCdBBF29G65NSlJMOYbWqOLFrrwNN2922sHZtFBxPtJUlrPRd97Qvb57gMaR
SsvEvw2a3FJQeLCVsfcs56U4itwuooLuoyA1Qc4Uzsg7JOe7F2yJDxGO6dkg12ichL/n9EHN0nHz
bVrN8RSytsj9tvy7/Ch7c3JNOmTl8IY0tUMHXoKFrfZUw+qvZZiKyO5g0X0jvPdXpu4inuY0lXYZ
aefPVb6RAtcyEgpwagKnJ6Uuf8WALyI0yl16Pa+TuPXu0p97Lb/zXCPsOyz6jrhrjSYUVRUh9WcN
e7t8EexmvKqenEH4OeDVKv5q2EWCw9mF58jeDKluro2BINpL+BFRmoAtNhj7e1JrizbNPf1X16EU
53lkxADJhWrJeffj9NWZXTxgjQLCCqsNtZmxj3jtw6Cg+jokCSa8+t62ObtVLTRLc1L98Shctwrx
/oz5AHxT5FKOb9FqeMPDat/9WYkDzM0a4eB0NaqxnNs30uN8Pba04Z+Uafuj6C21p+4g/zY+JUBV
9XL6EhhM1wC7DlwzBCjA7MW5pcXycAUCxQYM6qiG1HI+1UsD4oIJ6aaH00cn5vilt6SKoF/UPMOO
dIEuVSsRV+GlvqxLtRhUYiz8p05RnP/VNcEqisYtidyhujfSZ/R7pIC40TlAGsswGpRb8qitBPWf
GRRRHK+hjIhGA6ElnWoHLYRXnd1hZzSr2MXViXHK526u+vcvHbKo2g9G9qqQQUGl3gylMs28riDG
WsYlYKB5xC2YaQ61L6udvMJWdYwkbZ4TWK93Cr2MJx/KBMxbTwrJczl9huREQaaygWy6MGTlFWqZ
Cx7cHKj34bafn8LELPqUQakj3AWQmBiBhMejq9a9rriuzOv24Hxfvps+xqJDZhhC/rK5AuMQXh3s
Hn7Xxt2o9d2cri9k84/yCz+dj9t8uog+h7W74WFQZEB0OjRtsQLdiSchxoAW9cAPb2QaiT7iG3T/
yIX3OG/so+qAUCqcsi+JfPydnmWAaqS5S2PNDVjiYwM/1pNnq/NMQnr2VWGYj19XI8ruSPZgnqqY
UUKvVYUw4wHyXHnaAjTIm45HdoxbSDk+xsKIMCIq676It5M8Kf0BXVjXRrvRjy7ya4aqmno/DRu+
LAixyyunY+RGMpQIatI/gWc2WEMmFx7zBUVogpZikP1LHsUUQ1mZcT74cfZow6I6bOaezuNIMq3G
R7ZmJ51K/1p136u1GHj3qpRTYfaYPyUfyo9+vL2auDlZIpCyheVthJPje7mA4smjFm/1eDZk+oWs
gniFS0EL9syd4xvWlphmnj21pRPpmLmOZnyyiAKLQGB0tb25eEwEC9V+i6TUtyZc6aQ1O8yWpLhu
ji/QaDnuDGzmj/4Eo56zXJ5CxMplVgmWNabXCoSrlqW/CuDBPt0lnejt7sUTocFfexgSjeup2B2c
QUjN0zsaJbPOon9XZ0okhYnehTbcM1OViOPkvNxDOq4M4Afejpvz6E0UQa8/8gSN3P4je6DJMRCV
gG1CxXEYs7E0JefOfiqtzH90j9lqEVnjDh258HIgzhwRQTTJQdbtTvMpy1b+iSMB2QdvSI1rstkV
bVtAMmE+hSMlPYPIJwhNLQ1+UBgNBdKkyoctCfvQBCAO6U4zKz+UcNNRK3gJRznl9kVCaezyBSz0
QfjfiHx0ZzW5xUqcJgolz6vcBRySU3DXxtzeK2b4hxjNQg9vfHU53Ly8wvNpIP0IucWlvQMpaJZc
d/7OX6vMlobEs+EckU+Df/PQBhS2/32MxO4Am0xI6XInYh1ZYg8eWvtsY2LP43qvQD2oMe/al9i+
n7sfnZZD4+xWtTdhyHv/gZpGydHiMekazEPfHb3OiP+qL6XPt0noameVLupLIEyaXa1mnimnBkDO
/vJyHq10szPt1sMJboERfN52hbGm6mjn4cCouHoOWSqCTsR87o+FMJctcxQk8RmzT3sq6fh1+eHn
h5hiNkMqq/O6dUbZVYrH44eBuy5bvCk8mCvIoPfedhdHhuVRmWigszzTKyc90E6ej7UfhKD7V7S7
oLwbvBEOmZQqItH5xH/chMsV5fEqY1P+2dY6z49kUIgkmN6gvB+GehcYrGdEPAoE6xgyNxX6QGyb
fKCCuNVxdjoMdsdF0k7NfY556erhybHgy830CEY4EZstVRkkskSfJXk6PQPLdrRRhQTnUmK/YV+k
aF4I7sj2gduzbbGAFADrs7tQ9xQhpQc1jeoffUdsG5UcQqB6ls2ItrRORxWileHshAWBgiYvGrAh
2q+o7xsWx8fviS8OkZ5yHPPs4/dy9f7sk/nJ3yl/cHghp3qjNY0mmPUg+4A9R9jNbF4dtoENDsCV
QJICz4RFEb/1QKAa6rR6FmdOo6XcXH/g4vvTjDKH0tTeOQo9/AGZqrgUl2LC0Totp3vn7rMYC1Z3
dBeAHmLihjISjJfE14knK1ITY5GT95PZFtDVb+BeYS193tBaatbd+Urr6zhTZq2ffZ4mg2lbwJyg
Wn1qXuTm0rrbesqdXBzXqBxqmIRo1Beo/x9m/qt6w6Q0nBSJmeNvUpv+QlQGWhF1RxePk+mDQAv2
yQvS6j7x9y9GizMX3BLA4CNGLbluQamY9ZHkMTOjNOXXf+1Gyi9Vy5s89kiW9zK0QaUadZvhNSHt
/grUDmFltNxAAApsLMMDJ4EkpwJ/Jogdhi2ZDD2mglc0f4brbbqIi1JDsw8ISUrA75IddLs7Q/AY
3UASJVEKM8XN9azrhe8bScr9WkThsjGCX14b2Eh4145OLx/RSqpnpoOqi9LYDj+1DbkFlGn9reuj
O1My14IoM1l0PKrjF0dzm8LGfu3/ft+pSYQwQ/1jsDllXstTjm4nzRWYym7bi8cjmGDQ39GjRdwf
7iCwDSYsHQ/ScExHu2iEzcdjoMaBtK7rh0CU/cGG9Xv/a4nN07W9pv8K9rbJwLzV3yVy7DHnOQvG
LYcNQsriP0Ppnytz6Ykz5MF55u9W/D6bdXOGgESgJyH/s8YCsoXpJEWqZOlMlr6VB1D2nszbP9KR
MZS74kmUgbMgk5X1Q7c12wUFMqRPpiLU1ZEJKpcX1NV45FV/8qz/oRnwtkz/tqSD6O3CgDQPWiYn
cwpJc/801nnuO9HBi0RXiHYak11LHcrDZUcjDZZM3D7FlTJfpgy0+qvCtDUEWr4CMK+IsV6/Cjh3
sSMTJTdmjEC2LRFDik+2P36NBj35xfCJiu5Mq/sij3mASgn8DiA42M2qMgpFTX60G1J8WXCIchpq
7tHKx0aUejb2j0xer1vaY6GbRvLafzivNC6l4FyY2hRff0FJrYPS6t+wizZzvgCVup3I0oI/3ZuC
skbjaFEk0g4VIRDbGafHz6P1HLbV4HCuNtLfcaB95PDxNhSgs2OWeScKqful8hHQkWWokagxU1O0
T37ntzNxFI+F0x0dpGaBDA3vt5LAFPu1JqheTINuyhTzz10zcoWz32yJBgIN6QegYwa5PU6e+Q1c
qaFl0xhwFY/Mnt8jy1J2rPAd3qtUFLp62g4yd3OPldW+r0/t9s6xv2AdgxByn2vOhx4PUpVE3+sy
YhxhBcjtolEOs5uOjZ6OQ7A+kCyDhy4/fAx165Ln4O1qM5tpafOUyVMNVWwuXdaUgVMMGqIc+Ywd
c4GYxr1gCJ+BT1tob8htw4HByIVvlbpD+511bX97GqVPpjRCOwJNwn082606CvNJMQt3TU60KAuv
IhKPCvTMLE8OmgKiH1Zli405EOIw3IyVG0I3IuNKDKIdgzMqHPBfE2bkz2scMB0GWUXk73ZAQW8o
sqMZk6M116ZS2woneQb5gorbgVum8+07+ciDPTPG8VUg3jrIWzT56K/5m8NZdNeUbWAad4MkVW0x
JjdL4x+5LeADmIjWjDOU+lCThpj3thcU7ZZexxuRkmtOULnzcF+fr6rydMYk2OyxgYgG2NYos+qH
bJgjErAuh9BjRoxSvEx+XdrKl+8RRRl3JIBe4r1kkukMQ+u94AbEBBVjo6TB0gnmMzlmeS0rPsmP
znuwHFI02VIS6qi12s1O0few2CINdfYf4Ost6C4x++UBkt1d4S/tMfdFaNjEix3lGaCahcBBaWpv
Bn6LLk45fPNo87Gpx4swabxrZgJ/RbN8YyDo/PWZcyLFGS8RSDcEKWXwHcyzrNJhfvYKXL0kBF7w
b3S7Kuy6LSE+mVgS+oSZRHo0lgrHsDCD8m+yDbifDzPZAJCweighbHzNcyY7bq/8TG7p13sIdcup
/OpabBvHbw8QkVC+szTk1+sp6lKN7TfuX7ktE+7wuvxhzrLGQoMR9npsRvKpBy2wrBMYnDLIhy+F
iB/r3dw8MPw1wuSFMNIDzyfMwrsas+oUoEbqTCaYcwWNIrCDfKMov1YYEI3GIkX9Wrzd6SlLPFzZ
cHbzcSbcntC6aBBYeNOZCBFy4j+YcB04vg0dm+qOrU4kKnVwt4jFbl/Emp+hke+Pp8m7I/JbE2/L
iU+LXBRMp/GizeIFgi7Icv70mswjhrESHNsRk1xlgPFgs6nKNWzceyMylW8sEvAbRyDMFMcOgMTs
PxzvBwLHg8iBHF04TKV1y0YWgxVp2FKFk75Q+df/cTjzBboYO4eJtgnI1sqpjg6f5tdAc4gggY6y
Zkn1/U1w9Xkhd0+RZ4Gw2kH7O6DpoUHP2ANk/xk4HQ3B/TpMbkDLUddD2dSRnV2GnEirhdC40czh
sL9bHLYocmvjaui8sfQ4LJdRR/tlSWfzNI8+wE+tJX3cNhpanmV0q5LAbgedVH3NXuHvpU/YgcUr
cARctcC3KPYVbI/pLKiM3uInwiOXjnJTCQWOSn91jolYqzx1/mFC+KmOof+hyTIluJwlzuDqUcGA
hkuYMQGA4ZfgyFoILxz1MTH8Ob9L+j7K4THdUyezvIK1ZKXK54els7QwRI/MFIylsZ0Ba3IFsSYN
rDPxobSvpvYop2nICp1qeNDJDCOmX0KTaoqTNZ0JuahJLecIWv27rCvRK3O/QTZ69nBL1Q0F9KlR
XbsiE3GXSummOpxL7OST+2lNjp6GwwMx/zOb9dNIJvOKHxt1fX3j9Icme8qIXUntGhS3LOHejMaX
wqaMX1pK6WrJ1ND0VoP7yM7Ta1jwwhBQ2S6ScH2zbFWGs86vlUlTllx5iIMC3E0MfWFknr48FNC5
PtJK8VJxlRpniH61yR4Iu7oP6F9kM7dDpFJeFysP/fnssLvmRHFHD7W5oXUbBZrJoXibHCC87ll+
7zhnUCBXXauLZtsLZ2blHjLxUIbzhB8WvyhysCngCTYR1j4XV1jw8Ebmckiq0/C5wBvgSVl6plLi
QjX7yWqAVJxa3A0/KVwJ6gWY4fVVf974Riv5ncWwBnmI4PPWMEqJ/pWP8a2vK4r0kOfp7EGOL16u
X38+mjtMHvtGc83HRRST9f/iZkPYyry87Q3Cm7BHrg47oSQ2WZbwRZVdP2vU+TSrCvGtARyFTMLd
0xC9UqkO10d/LUv6qf91ZKuft4dqSdULC9AJ3CERJpBR1FvdcjoKvYJx+I9NnF6kZYVgsWlS3Fvj
0YiJwdWBrB/l777GKd5DnCUt7R61yNO9wXTotlFkwawjz82Q8+TwyuNQwZPYYJPuUQvKpVhAtMqz
TATtc7TMRecm8czKRXERn4e0Ddg2Y7uNTvJQiNse4MnM4ZWC4Ol0ISpXU9ib0gam3G8bbPbXYrRx
4jBUjsFKdkRIAa7dM3BIFDeigBnVqavLFaTuOUC4bMPR8P8u1VGL9okfHUiii60mUVyQsN8ava3v
nNXCOYnFY3ZdzrZGBypMF2SyqusMdZQbSHseFTy5EVgWgSnjGimIIaP0HlrjDTB+eUWAyqYaiTnx
QTFrDC1rLxE4l7nHHl/zts9IxlfonJhZJx/HgSHR5+68WIJonW2Rjn6ppP0yfKiWwhb5wp0bW3hT
qn3Emspp0MPo2iigA2P9s6KADk1Jjw3GZd1EqMjXO58rha5mGtwFtZ/zuKDCaT64itzjX+Bm575/
QfuIGFkomM7GuhZF1W8GYPvuAMKVdTMnSXwI4sgbx+AF5kAJeg/x+qKWnLXD2nBmACKr6wOSj7Dx
x6xGfXwnJusWbnJEvpRFNvyDsh8IUL8+EIy4EdbL+eizmAZRMb0IcUivisORT9gvMBtKyWQypulI
j1uDEIbrpd0srKrZNOztfV63wmr3SMSSLR1UWopf6dia4UjELaxYW2b9pE0fTZBr4m3RE5qmk6Ab
8W9Urql5x24J3zaGqo5lqK1Us/mZg1UUieyyjTmjQJo4eLZWDZ70YaUCfq6j8LfU50ifqXwO/Hhb
z/TKEtXBsEcyWtNSCCY1SNSNGg/uXdXh8ZBvGZSurJ/5KYdfcanQnC6DVfM1RoNi7caCOcDZqtlL
xvWotiKm8x2Z3ltZ+gnoyrW3SAssFEhfyghnoK7behQjDhA9C1eKXDfF83suny8zPOUtJvwWOj8t
H5S+YZUuHXBx5caCE4m3HWQRhxPCKS6F3imDrVZchhtQariCoyP8DAVBeXxk9V0j7YudzY9G6YZi
cG4HoPvZIqZIvli5DFNrCept9i/C0ZH0LCH3KOk0QDg/rJy+maMdVhumd5K26weJgimz+obzTE9z
Fn9EnaP3sauRbnIZjlnqXWNSGz72Yhf09Hnffth4luyR0vc9MP9RwXmYCxJoiX6/3v2e1UF076Of
ybuzag4WSfbS7aZE4ZwIbaL2g7Te4fOFnFqTjR7jmVOPDkqAgKxrhEkh3GBYYOTHeulPO07VJCmX
pQjMr+lZ04XnQNTs+vJNV2wYHStKtp5zKpV1zPMa7VDYXzoDktaSBOlZmb6rkRHGDXY4Tf1Swls0
5nM9r06wl+GBvlc30sMpIDNb8TYUTL1m2REMiAk/To9QN6T+DIWzYxFuzXI1lA/R5lSTy/PFtqLa
NH0X59n7zx2JhQ4NFNsV8KT4eIiyWnW4v77ridyNhvV+9L8xv7DLOaSANwK+XqK57KJxphK4PGlV
tXuzEm66xZXwelJLEdPeMVoaCt6Vf2WjSaEkTZtXAfyQ+S8flmAG++ClopJbpcREzVcsbIU0cUjp
/YlxHa4A0VARIhJYE13vVwilyDGWpNa4XNNS9HHmyKY/TSGJdee/PVrHE6Q/0GQskVGXL1klKVPF
RgCXe5JGzadC7muZTqaBLQZXgAnVHh4FZwbejpp9ZY81xr/DFMsBZBcrY26kmuG57ZmFNgA487vi
9N8+uFCGq71dwIunqK7BLjlYcQAxjFL4hk0jzsBb8dhbxscUIstQ/mr1MgrOEBEUy24vDds4ibaq
4t8EM0iVmKRL3s4KJnkbT88e43aBBIN5oY0FTmovvE1C3OX66f8ly3W9ULV7h+eGv2ZfpBCsEQXY
qYXIexym38rgqEJttQ+NTbVp9F9TNqlVbiXjlhrPSVM2Pt4dnaJba1QD+tXH5kdzwZ5v8iu3a38H
BLp3CjoNkTJFM7K6Ze1gcGhcTkkcc9mJYhGK4SFXCIYY8PRO5Vni5QN0Xrz/0JOzDsYeCmNux4qW
Cg+svxEePCRkX/QVtmjdfcr5afYuH2m0QG3X58/FvPswrEyOo8mbmElpYMjVQjace9foNZJBqE4n
Qt5AeY6ydPuYYvW857uMSvFIyTAOSNIwgy9+CTiHxqLv+16zJq4yjmtLgGQMnbLD2a81QZjytdIC
eRBAvNGi/22PzZBDSnHJWQPd9kuH1dloKQEiLcBOlKvxFSOKzrqJUOnsTvgkcscYXepQu//B/nix
bOTAwPmwSQeYY4K9MrBHj870ayrB8RpRGN0R2ioc9J64NQ3TDxCxzCx+a4kVqF77WJfD9y26/ad+
tjMEHIW9rRru2w37CY8G3cRToyph/9Wb9l8G/qx9097egdgtxaCIjHL/FPamK3T1UPpgf9P4ktrn
UffCH4T3PrlqIYQiOfoH0m3xmkHMKQ539pudECeOQ03aI4jY73yzNpMUW8xZWAEOQ0yhUUvyHbe/
ESzVdPNQKfqwJbG5zSEcq7eAUjxHcSYRo4FAR0IlIW5XZGgb5FJHCvtXgTHMC361gny8yCHEpLBF
CE/+Gs5nmR/HFtaHXJQi26sA1qvLWgit4WBnw6OOBmAaSBTTvGr4VD6KSLxxNvqnDoO7o4cGMS6d
tyFFkNwnWlMvmeb0qbMvG5g5mqL6L0DzeIb16lz/+KiiSOU4IAVcEIC0F0GmvoF8LrlckD3SWAwS
6fyE62jBKoA/Y270mBNeIyGbirL0q2x/18H0xIkZxKpFigHu+yQizk4ywxKmnD/4ZCF4ahf6VXvQ
2Exzj1t7AHWRXY6NG+dTfTCLCkmeYE6G63JticLBSx/sqjARlivH2eHvjqu4Seu+zxen2dezXZUj
5nfzkSbm4tSOXbWyLd8PGaQAhWpm4xHtVXrNr35UeoXEtUbRkwsM+JtY3jIssPtHxWD2i3CEAgyr
+rSybCw6YLfUfJhFRRdwyedKlAQcJxnj0ox0NO7rDatKWW4DAiVpeDZ/K7Q5XpB0k990bcBTNVNs
2n4FFM98VE8nMiplCPX5uspI/QS9gNvqoA4lTH/SdMwT11HUv1U1z4x+qHb7oNwekQpula9ZsCJN
U8rfduI9FFv06R7lIY26KuGcgZivMPGNfhHDVa4HwSDYDoEO8VHhWKYp+p7xW2C51DZbmeH2Kefz
z3lomzXYZ4HP+SWcv5hY10DyIHnfY78X696tOkC5jVZtj0hECBm84Jqibw+2PhoDPmvvaPl+yYNC
fXSosC2ujfSjGm8LpM/bSTSS8mZRx1KL9vjtSHl7kmVj5T8qw9amdlQCvWT9X2q/gOybsoQsByGi
GkuUkBUJVx/pkAT/lraqvEoFXObxwyqE1GUZe5sRhuRL0m5ek2rXZduECbCQnOesQ8QE3lHuGbey
z7xDwnfWSjLXZenl8t+FRfrunx1nFAqbKD8iVhDctCbczig5ts7eOjgGQMndE8svrG9Ln+enqleM
7JDA4p9ekaOFj7C5XHNBg25egsRKMYpJVi7CdesZBE+P2ZIqHJ+q1GLmhS9GRFPwTT8zUAbn3j5a
KDYZHMqjNihhFgcXY2mp1H8VTk8yNJeB5Fm8CDWe4cgwvtvSHnQ9vnWBgLkORK9TEcgPp06sMdVW
Wy1UkAuUwm+2ymQ2FNm0EH8HqsQ/KMWXAnRGjGj0/bOd2CnqM6wuVVRqN+8dHqoW3657+UvlJInP
ySU82phzFnPsWWEG5iBwdeuGSM0iJB/7/eP3tpLy/IGfGEtdJWoPQZ5leiRSqRTFINdsPgudP7ck
M4+d91ykOFBUTQ0qqRtwzz0XDa2+283oT9rySKQLCZdev773zcRoll9cCo7Nb6KnDL1EsoezhcTV
vrgPw+72mMNuisJY5kkXoEls0iKSqNxE4ypDYbgxyc841zfmQ+csGoRfqcN0Hg1O01XUXSbGxVH8
sTluzNMpxmywyieFO3PYKQvvjSEuNK24sVSXW0vpM5vKU4BYFdnbM4FnFclj1a/Oi7WZNMYvKQCo
QUbpJemnw1iXZ7A/hXUoGJF3VFY9WqgyZ4OIssplrPc2wa35fkzeaABEOhoiBQjvMe5vFcp+/Po0
4ax6DkKtxgLRpW3RSr/vgXKVeqKD7p8/qPDCebiooObqsc5lxIIBrfU5S1iYpgaZXWYmka+C9qUV
dQduwngDpR55MHfk9sj6VR7TPSZbAm+Fj0QUO6one0VeehqUHF/ZhfZQdfl7TS8MPTv/wC6UP+2j
zAa6IDwfjV9busQwBPXkWtIN1cZd9ODzSZtBvZdevdFJf+epJkM1yb2Vp57ucn6x3vm3vwChr2WK
McLYny6RlawN06cfvcyp8vYuKAQ4EtJ22gaReyBoSoTEnRyiozuGbKAI/0Uf+UFdHDSgtCTVdCMs
RKzN38sKMcw9jKjCa2mDu/rvONVMGIydq/SNgiRAbZb7aRfWTStPRh1b3rtQPkAPlFr+m3jrXJPZ
8CNRVr8RuA+2DcLn6V0/UED6rlK024CqroQJQlAteTUXgyBQRXKLDSoqwvSChAE1A4FC7EnE8iqL
5pTDop6CN8cTFV0gK3YpIbFVhZj8AJytzxnYNoRQZaZq13B6IX2Us2CPh6SM3KdMVj39cWbiCw+2
2g4VwZWBDyvRkYPEC2Qg1HTf0Q08vqKlCRSYqV5bm+owXtq/KeaOs9w4pEmNlKt1JUG7ukfpOvfX
mxBxM119qdGlJD30W08ZTk90l0NcASKJgXfTdg0+YUCKOcXHPfxDLc0V5cwazpg24/YHaOkPtdI8
QODTeBV1wM/stjp6/KxmlM8NxAJQ3ZnPPRN7nWtY/LhwV8V5twjfRIBtpGzQagU5ZmkHHxALQytQ
QqVd5pyeY0ZOZnGQjoOAuzHzPQw8PKXW2B+ITey+q84+M6vtSG7WejiZ3UoQXBnzhAk9z75hXKHJ
/+VWLcULAsDlxpHBs5sMRPW0T3H8U/3TrrDvQcFVJ8cioQ3gtG5THXV4sKU6+CxjkRHwamVYzXdq
O1AV2AxrDuhSFfihI5f6ZTQxxqzBa1Ime1HdBKlEMwQ8W4CQa1r6T4NxnBCyKZbU85fHcumDPKzj
zmaT6RxtBIJhlsJ5HMfFDfx+eslWOnwN7t7X2nKHjz7XayU1UvPbGThzUYF4Ncj/gO8Ci5u883fK
5ikFjiG60E0MvZY2I99flkN7vd4EnX9PRGLPMdmk5NPePLUnyBLYOr/GiwhvsnWqisaYdtoHeEWn
S0vLrUZ5tcaZy2r3PFsdp9hVrsX/AK2B98XeeUrh/4uP2c3rA1veUGHl92WW0c2yOkSqLqlCfZ3+
kQADO0Hx+Zsfn6NS/2A2Bf32iVzrbBIWsS4T51J/lEeSKsbA6PEvWlVhvtsfXrj/1BrtvB3L/IhT
h3FB+ak4qxkQf3Zqp01fqFodmVt2y+BbzGQT0H8ZFb68dg36+J4ETHgXLlshtoqv+Av3CgaOGGB7
8PIvA1PzxWrFeu0O6rC1Q+yEpot0WCqMI+ktBhdVvygTQBLbCwCpWtBjekmNFurEAwXsLzlnDqRZ
f0De6aRY5waHcwS84GP/niX4zdPuXAfrQsyzuZqerZKr+tKwmdAzESL6OYazs5DXKcyFdrhpQzzF
lOM8GiAXEc/Ii7J+RcOciwLR4f/DbbOgEJ2KtlYKVjPOr9DPFTO+RqMQhXTEl7zDeViebWpgj7i7
D4Y84Aju8UQe805tHcIs4RS/w6NrGPxL8P2b461neXHXJRPaijBxfABZZZmheaGBQh+uFr6pKL2W
r42HOgZRJMzOOyA61ix5Nowx0YbeK8EIVD+JvRxTGlTA5iRUXaMO4dBbPVcyg/XgIJkGBxr1Eu/E
WkHFjRkvmAespCL5xg0/v63BGKh4p89Ngb3ERpQBJi0QW56NntJd5QlKSf+frMVBAMxAIMS5KShV
JyJ5fntBU0Q2ttvxgN32wWsKk2ObagWHTkL6zkteCz4gBjF75A/xr2PUsAAhv6YCv/agOmBuKX/+
VwU2dkC1mbXjOlX+Pvf1mjRrsR2NZpOWcLbX0bu/X8K+zR3PjdKMjLiVKVTLi2VP7nEeEW8IGQXd
PMHY/l/9l1ChavCDhNoHk4j5KmONY0S+PhbasI3cP8qh9oWZGwe8wNHr89weqfkXbYybZ0Y5JIaZ
qBflpgVEP8QYIJ3lQ6NKD6F0Z9KaJ9wQqHqSYaUCgtEcCwzbFkt6LoSkVa/G6rS7NmIAOsOQXcHp
62/T8PeuL1AV3kkpjWvl7ZkAlurVsiSV6+yVV/RycO/QEDIS1BVydnFBmegpJcT1sHqJZunWqM+c
oiAb9LycKSbJt7vddeyiwDaaJNtBL6XppmgmQ8O7r2T+S5rMMTj3NmY+XFSJPctPVGTcULtRvh5b
8n7to4A1bna3Mm3OsaK8gZfvoC3dBugHxPiuFFGVZrdCo8LyCRZlPEzpQlFLJCSVp/egxYsoKK7r
+FweTmTaYLEEtb66BPyx9ddkTDDJRqqVZzihh2HkEdkyqCV0a0Tp4fDYbROyk4d/Pnh8fVESWtvh
4Us9lku4eDPRvmlgiFUnU6mmbvkSKcjAspz7A2qqc4GvBCij2yC/xK0ybAvwQOiUHcxgc+wEVtyR
qFfl2SNsmxUJi2y893shhpjCN1ZzAmikG2JBIq0tMtX5b3gv30rgnA1uyo7WYIi58z8GK4RTtxvG
3OxztJb1K5FAGNNSj8X5XAfkC0UdICs6Sv+kIl1K1BXkw3KweMJ+SSjUjVaUnLHGZyuwSKGfKJ5+
gJgPB1ayYKk2sXj35RR9DYcyaUfoBmH+NtItF6tWuRIfKyDrgpFsDAnnjJj4ZSicURzIZdakiWf0
h0yas5uQb/rV/ac2c/g3MDZv8Qe4eC9+Ex/btLFuKQT6XSlnQtwCBQgvg+Kw5YICvO0FnRUePVjS
mzMUGC1lYVH2AWjVTCpFUzo05HvB9fmLU7Fby4S+Aj3m5NihNEViJRQkXtZKv76agpXDuzdozyIW
IhGXa4Kw2T05Q51dPyG4xddVQonLL3wlQRxAI9Z5NHJ/tP6GFHwVP5ZKkueGFlnDO0usq44cSmj7
fbF3xUIMekJlEDLlCUDmtcjZ9G8nezBfgeWvSi4UQafhLqisHbudNzFwLXiH/Btf2wbgoCDLf2Lk
PATnFKlSgAh09wfuVmp+z1OBTjHXC8dABY9FXW+ogrJAob0uWBNKZdh385vLG/PvECLIEJtJ0Gtw
Pi9ur8Ox24I/dZUTWI6+G7w0SD/XvsZ8QqmPIHNe+OgBfnRbk0VBSZHUcpdCBGsIvzmz24t4of8q
Eh5Q2XYTRo7pUu6fiJnLkw6WWjPbxoKJ/ZgjyqvjDYGGdFFyGh7VOMVTdujkMgoSEIhTj/Glz4+F
TXzjgPkKY+STVUSTunXYC8uQ2OsMA9oZf8XuWqWwPoTOA3feoBe1TliuC/txjjXhiPrmTYg+MCv+
SWlpQ1AmkkBwOnaHZSHJOfCXEJ/8rQZPU+o8koZRveuAVWBjLg+REwZL3gbGYJ1xWFxJmsLV157m
ls86dCuzn3sKgdpYSgJ5nyqvHq/iyTCRj75Djoh9rsCt/bXfarKvTYUDKUgJqOmGTaGZ8BVCVFEQ
HUt61M5SLz7ZRx7upG1pOotyoKb68x7p6iw3oHOLVJpZPaAstAUl8BZrKAPqCSDFNBChGj8NBb3L
xfur3lagrZszN7g4u+0B3ES2FO06q6MlMnqnGQ4Ji3NxF7vcX4Uf6/wt+R9YS3u+FrCelBiIhg9g
YTH7HKuQC19JUcy2LJdB9WKaiq8/Akz1Dxzbi6JWb2XVldRwGtFX0lEaFH1rLetpxZnHW1iTXR27
dhy1RPYVuV8/9tlYQZTAAJAUivVsaWxLfhEfUdebGQilDVwgEAJnFUTuvwYRORa6FpOZPTzNZbO7
VIZbPfg2/zCLkgqxnVhVzIfNAAwX8Jcwt2lXOT2GFOUmziTVNis+D5Kvg0F7rFNQ1oiNObCVpDYn
HtbvqsK4U8AbagWM4MioOeFJ3vSsRvo8IiaOdFsh46QqrWxmmAb5rX54QYatAIuImurj39ExtZxJ
5kjeBrbJn57dONUgfkacNTjm1hudoVyfB/0JWNa6NLnYvQlQd61mrSYDOVJX3Dl/AdAKFXhbA40/
ebbH540pctiCkQ3TY7ckSIUhD/RHFH/j+y8eztkjkq4/ddxGvXB1ASUMC+e50sqjlgHOQnIRV8W1
Xw/gzWT6S5KW2M8FB3w1k/3B9LpaN7V2ZSDlxnNvbQ5CapLZW+qQIuN9LGYHXLViDXBRNZNgWrAz
HrISZs+bI9XcqYe+7KzK18UhKV4qC9RhB3QRwyNRKvEeVUjB3LJnZa4+jGQ7Sl0/z+fXjvzml5r9
gmGRs/8pTwGdwKa/u+d2dfCQG2Z4YTLUJKzeKJmAy24e/kxDS1TI4FHqOJZudYG1U16PSuxvJ7TG
3Lb2+LHej+1JN8CR7/kcghR+y1JqtXEke6YLNlpsPaCDWbOrcacHcHUHZ6CXOk5LAd/cP4cC9GXG
zO/d8HQyJlZRQstWHS9zz9bh67iNn3T9wmwk/VYxBybx35lFf29x3P228dM8YHbAGnwQ2/B5zzRf
y/RMiykgaPZbbdX9Bzrrq/XHoyw7DFRj7ilFAfh8knOmSFvWfttNxb8j2aERVOa2Selr/s5mOmCA
IIyhAsFmpyD8psTs1LV8HaSF7sblnlLyzaogLiC579ey0buACCXvJQNGQpBY4vMQ8PaUZP1HnS9N
Xo/x8mTrCV2gWEz/uRPpsqx1+s/U/b+6OwTUqbYxbcxwaOwlx2bRgmdGG/9xHyx5U/f3TfRLaNZa
hbbisFLRRX1Wmn/Mchqoxcu/96jRQquweVHiE2PKsYnOjQZs1Fze+/kE7OpwljAuZn9ed6qO8Jye
9vOYqOxz+KISNfTOjfH6a7BIW28MsVJU2qFZIlCayEaGcJLzFT8OIqcUeJRMb+t8Bk6VKWO8W4Ox
JsHZz4rL7QMq+ArrVCdaYdNIhdkYUxg9iEVIDtu2PsV5GqHkRtE5mFT+Ef/2SSBpPEmCOxEWY7WE
WpU6l5XyFXRz4HTq4EShaQEYAjucSBinEBAJ7wD+fl3qKO0xtmZZ19dP6HAUqUhl31hfxsvB8Mz9
8TbkVA71m9hHSVvNkjtmzrgwQR9wqKatW8f8fvBO50JGFWKaMdgfzaU8xelWjkAjLp6OEE+n+3en
JwvwCChoAHDQzKxC3qUnNCz70dghYq2dA2CVzcwAX9xmXJmULg2UiAGOaPhyXd7nJJTmYqXuhToD
ZBzf4AOVX7EiQR3FUoQKuctvQHLvS2rW9/sI5dv2Pt6ggP//f4j+7oDIQ2p/Z/JcTANkcsgHZkaY
v02kQkMk6tv3OTbFFThwnyzOhep+QMUf4udU3DLpqRVGqShKWCmzdzedj3+gt/nG6CSruDb7xWpp
MtsmFt5cEjUPHMhKFyP8CXw0G1tS4Y7Lps+sTgGtbPRqVItB44QfeA5OPBbZ2SkdWSqAQfptp9i0
Ro3bUHHBL88cujaIlNmvhJmAzfRODcDOIhwVqDwM+yj2ddCO3UlevHJcif32SVDw97S1RoDqESoo
bAavFfiWOfn5diiAdnHjlbTsXJAO+kZQ+OcJ2PM9CIpbBsIZF7cmCRufCJj+FU10KqdYzVd0UaGC
6ro1R4kMOJznBW7KFNfSopAuD6FyHBUpSGVrYvXmqiFkrxmmxF5Rf0xPt0T5vdDcLvQX56MI7p38
0J6PXJrArW3R36vnI4x4WSz2AJeh0X2M5UAkkcYnOob/u/FDKo3fBolMk+jb0pjTP/0Y+hNHXp7B
Y40Lm39Z3glbv3YslLn1rR35sX4JnaCqLYOp/bufUpuDiUQgAd2+T0ekBup9qeFxL4Y1Dt0yzX9p
VCZiMhMPgejZtDjM0V1vMIby9riXSKeFq2hlK3YHPqoAiJcpjHSX1BRWckLyYJflqKhSyzicJESZ
8yoMpjNi+FJoLtQoYyT0IUPG299Lf5zBxEt8bE3P0qBLIgDzw5kAuRceYr0m6UjH02x+g9SV5JJz
bSIzhHjmjosN7Le6RWic0HS5mBAd+GTaqN+7j6dU00aBaE5qPUvTVPy0MvltnDgBRQlzmEYE2jSj
G4uCmYQgzs3I0wBOyNR88K1uNie5dXxN5zuPxPXZFuQToK/mMknN1jgXR4PIEcnD/WbUI44eCD6n
tZPaGM7YyuLuQ4tM87lQz9zwuU/DkvPh2Mrrozj7Zp0V/pRlhMsIygABCnkZawWkwA9ef6p7Z2en
53Q8adVi2vLnjdcg+9p6+ry9Ag/pKf052kXQ2g6oO9kxW9LSb3yfIvytHzQ9uNJZ5Ix5+bAaWg8R
rWsgJCRjZ81oljpYeD/ixVX+FnV1ebU66UtnSUO8jbq0UZKJcuhORS707RAanYRqu9n51Jspajia
2ZaRZOXRV0IJNfrR9gR3hTc5HrHjCnVWO/0EmozdjTvhjwAzA0K0hWKLu5MtLhq+1IGUBPKJ35XW
+m21oycnraFIOzkpMHmm0QnS+NEheM43OSoI9bG09++Tu+k6P7745XEoOyMHtsGPWxJlE8FSmv1W
EvgginXAI7gfKaBNuZ/iOLkrqW6n8XnaHT/PIRDF2LFhlwjwfT6yiZXugHE9U5s2gM2Cvc3xsKr+
/DD74G8B+Knt7FDC1fKbBNb6jgrnAOr7lBEJnwiTShhdA0NJY2Pw5AJU+PNNHDJkKqhRElsj8t5S
+70uETjLVCXflwN8nx52jHhKCyqb2H8Si1oCKdT8lCnLaS8AO8eCh40Tv4QnWO9ZyuxoK/qPpp/r
B5bivFuDjj2comkF+9ySjqn7QvxIBz9ChwqzSCPEIE8CL6OP9QhtY545PacbE58iMrBG3WdiMnRZ
LqX7Kn1+PauFK9h0lN7aHBIFM/dwBuArKy0q8kgrAfiuvhwhQGvmLpsXWaS9iF2NUv1X9QR9h4VD
neN3i2H6IEdXjS+Ob8F9cOpwXUS1/z5eOyNWbCg2uoUylhPI6i6EvcUL0ly5xtwjvltVXDtpgzaK
0I8mRUOkfyDkInmSOMTLktw4Pa6VLNJgJtvAsr3VSWmE0Ab+V+RX1KIHaG6sZayDA594dkn+4dYw
1gl7VwAyYp51qGRB68NmsURTYJhc9+IP8uc/o/32If3sAvC/ZtaVvsJP/+wzIK7tn4pECLPIwmZ3
978xcCG1TB8cIz9s/ypbt7s90RLn6DpOEVEMBUrlquZQLOF5E4D+vyPcRUgo/dwka4qcWBlC81F4
ex5OyuledCWciy0jSwzZe2viwgRX4+RPdYrYzxOJUFe/OxWNCdFBDDye3/7Ii7bG8ciyWXVeFJEx
0ZK2EAD2ztwXoWKKZdJLh6Gv3JRKQUpVt7Bqj8X3fQMh18fOvUsZ9B4kkc1z1WSOYmxkMONaNt2V
8e2zn8nhv1DBaQrjAuqCaMjG+5oQmC2VheBNz/dYdx5AzO6N2z6ivYvRgt/G/gc7zE1TyqLPnky0
rafb9iFAP/49r4Bm/7jIuUOeVRJtVi9N2tAJSgkdQP0LV7z5YBQItbdFeIuDlurb9jdnunCxJf3f
wQIxsyuP/rYv0A7J2Qv1Q8T3W/JgHZFNIemPiJy7hcYfU+AuMPw0q2rvZhlUXmFtFkdfalOO7OcJ
chX5r/wwPkg2eGU1i+mIUC5GKotEsFS8iD37sCnPYtp/wBKpj80339XtMzMS0ai98KKgri9iMoaE
fvFnT1KFQoO1r9t2loLsT3vAKJVMI6JVjRuMHCfoy2qt9nE06X7l+/9Gh70Kqq3X0LPYMxjaH7wl
sgpGshoLE523RK6kSeEyyw6gXXVXZhVLtz82oQvohw4AKuR+KqUAmxz7fFO5d8p08KO2XXpKnFQU
UofZY4f3o50NBEcZBXA96ep6E299rY3PnmWJObNsOqkp3YeYOH4Q03UbVHKUood9378aDPx7PmHK
SsO3JK4nGEF0r2Sl3cnRjr2+utf8K0fvfIw8zZ9sgXZkSsiqltVkG0skjIuODLhFZeiz098i2Zau
1SPhxmAry6Kql3KQbSIxVLdOWoWHptPxm4W7jTgRB9goib9Ab/NzYHsVQHI1rrF6h7sLRKYIqu5S
Rgw5uFEBa6/QC6UVaAvev7MZhW+/b6WY7JDYkWsHPMQesXFy3ZE4e5qq/zbRxEzH13lvX/xW10TS
dvP4WwpXmU9LFb9hQYcHq6o1nqQxf0FMk7FZcdJ0MIk6TEKoNOmButoay1IjVmOxXLVt3k+PkboW
6EofaBX7vEP2yuVZ44OmHd1egUWO6SLjG1JbgrqdIyxXUm9PfCQuI4T2x0eP4b6pIKmWmwFd7SBf
7+iG9aZfxByUjmhV7KM9joSe2dyq8dPjsEwX/Nm5fv+4VEE+WQ4kheHnPYDicCUraEaeSbwcS2LF
bcGwSO+e2lTHkzmJ40JfWrErUHYkm9DKV3eM09TCbDhfg/Xzp+FPu4TUjL3Q6+pxtkHFcftH1Mvn
PG75p9sPpSV6yI0CKBV2SyW/RlgNRjH1XZVS3C42+U0JAdVIKETcI2Q6mRbUPv57CsuQujlwkch/
Gzcclmn7Ln1FLghLYY/+S9ctVUPAkZR/aJRJqXCdH8wSDiboxBrGhlLLsTcqO54C+2+5BL3QeLI2
9nmdB9A38XnYNgj674/C8uTdSv9DhL7VG54oflxkS8knm2lKqISxBwv6wrlfYzXNG+/q3/3OZV3M
nbA4G5c+mkZg74RaEAUB93Z4zmIGre4R7i9WAca44X3H5OYeQlvomvOiEwYxRisTK93JCtxfalfM
lugXy4HEdoZoEe3vzl/dRcBei118qxGaAjgV8RDyQw2BwHlVujwXaOC4UfxViQzQ/bpZrXPYCw22
3rkEQSIs1IHSJTZZSbepO9PHLpUECu8sMprbO28heE+FpAtSBdWuPLbt+CWmUZnzjbGVv57VJfaa
teDx5kEYwrYkIPXHcKyYAS9vouImQVNAPuL9S/zfhe1/KxS+sG1KBsS6Mlnvxv7+FzxYt4pL3rD2
k6GjIRqg/cHEYNlLCpwz52bdRVbaRp73/YYC84Xm7O1L6cBFmJRxybgQnSPhPl8XeCfphyjR1kbi
e9ck+FFEaXrmvxU18EiD5Kmufj5GIe8kJI1uy3VlIcWUtOBu7xzOwbd0mwbXNsTKQ6RaxE3ISG1J
+mFU8jUmHgUBIuTexHcFyE/2PACqIUTa6UdZ0Nd78d0gv4HH8sHV1+b+kaktdzuCvUjCpiTQgjA7
ovmGZokAg+A2bgmdsUUoVjAzGlLcPQ1oSbahRCVU7jODjNFAxMf+d4q46T3osLjUOBGVYbSAPAWc
RQ0C/J3zQ92KSTH14BsRecjkgl7sQmNy87KuOzRSE744B/HvtRVGm2AaQQfvIH5aXA1g3bVoTkyI
pTXayqdFEphEwDlQ4J6/clC6t+W/wfrkRuHqzSytETlkvJ6PpWRAnF71dNaxMiwr9R5uWYMh+Yi+
2DD23NgLxa1Bysxa1a9DF8yQOAMVbNNKb6ho3y2e0y8t+qf4qHlS1pJ/A0kaOSpiruwLOtfrotlD
1CHirpbHYYW3cxNG8K01ZwU4XxpAN+zJVFpNYdX4ygIseKBQ1cvnPkqmnPfwnZ9wjSKynqN56+Ml
V84l5PsRM5MkWOFJpyOfOZphso8A60nCHqQl4R6jbOujraFT/gwFBxkhNnRFKUASrsM1Zlas5WNC
rnCQ/sMvfEs32VOzhFh+077Sz2GeWHWy+UA90NdNzo6vdO85GrFrrAzSqtf42LB9p0aDNFSz6gbM
sVC6n8bVpJCZ03mdww9nuMnUeevGepvrjsaRLrDdbnernPW8O4ZbA/YA8EUOBfTfOGVNDxQROgee
hQjL5CYj4hI7bia2seqnShA3zyUxi0ZCgy7zTkw5tATUMlTwmdTszXLsiaN2J/5/OK+PcPSOIdyn
pDwogdff4QGj2SHItglfQvWa+5JiEAP78CQfOg6Z91OlDHoRHz4Y/QPgT+gYnedgCt0QzmJu3u82
mkw2RZnTkbv8FgjyE6i35+TtHJYzHoa7g9new9GxWIVAqoHhqHhxfXAjDh7cqS8VyLU2Sj3FkfSx
QQunI7pWIus+osLv1ykGix8p/VtpIfTRZG53UBXYOhBchTDGMMaiWobk1xsGKwL3XhYs/0I+Rizp
rA+spfVFl1dS2IgC5i0PqxdKkO3bv0xZFKDYsUUQAPVKLde0Hs5zyLqcDC+rmHE1aayd1uFILJWI
/MOqdIfd6wW1L++UTSr5seTSeeTvG4PpEQWOjepk1nLosQPmv9uFjt7pFBCXQTbOiRH1HNI01+I/
WtMm5ZgT8AHQHoHPo+8agmNEnXHj6kh91y1gk1LFR4x4Vo+znLgxsID8TsKHlDayGg27KCkYAd1h
BhucBIVLTufkknkVsJTq2vzZlwCPHtazp365/pZIX0tuoX3CtjKBLdyn72F0YRBkN79/i2oeebSw
JRHwpwaQK4Pc5oDIV6ktiksVb+AyGautJuPt4sE+mrX2efSy4x9zxOF7TDGzE/shYnCCLTUq4mBH
ezCmtyNklRrM42ZqQ+PHiTzNRO+i2XSbPU9qc/k7X2+tQshsF9Shu1VJU4yd5E90rjy9DYfxz4yx
huDske6SJWNhKPScVodwtjFjqKND2nRMWP2v0I9/OSQgTKtG8QrHpbhKhgRy+qkaHn7bCjT2W0pp
4FiOESMwxW30khtthCTusw7+BxAMjCQpCK/9gDUR8FWGbwjvOp1T3W6V01cebUwL+yMUJu+NMIjU
9aqZy4I6aQlViiFKBTIK/BTqnHNdZyx25+ZDFHkqV7fNHR7nGjAj9mohIfzczqGUJ3PWItQAyYgF
/Wuu8Gb1flIEwjsN9DVU21uKpzY3hzzFqFsODZMQcQuSywh3Oq5d3Jxy/yruINVNVWPZ6OhK5RtO
zA5jRDlazPT44wj2D89OXZWupM3nN7/o3OkLmgXPU/qwDz72pHSQVHv2edrOSz0Wg5qrpDwgg/7f
YAYSyl9Am3tE7HnVAz7VYxfcpLQInnpQwXvWnTAMKsC+l1+ewXREvhfbF3CV3C2r8ldWJRMmlMby
fKIQHrqkwQa6oFyPyKqTV3RM65uUzFdNdJOGgWawHj+8Zfec8DxgFwB0z8WKVau1ujeqfCF18Sw7
/JA80Lnb4hQj2F1Evg8/+YZ5n5PKqu4a0P5106k2p1A7WNtJJ9Kwa8mkByWydBUL4ZL4uv+n7DqN
ISx2B1QzmuBpvE1tRwLs4qi1Zv/PIdEv/3zrJ6W46AEn3SFMsQf/rM1ImZeKwqhiYnmBCPnUjgNt
v5EeleP+Hs7NC9pi8XyLCblegt/K6wwGP7weN5t86gR3nAP4c5BGlXLilquv0JxDCuUUVMuddMJ3
0LeYAQv+IsaFvGx6PRUKnoSQJLbzr2tZ4URmhhWeZS9eISBsHfCEPQzJPdjg4hrFMZO7W6B8MmxK
hS0iQ9K60Yo+rxr2REv248OPrjb5qikeqnrU2MLXN/jI/XEMlfXO664xtvVMV+UHrZzYzh3Tcpie
jleL8BLeCgs2IrEduzhFzicLhbrEysCuO1UIOgnUE0rYAFWFpDEuGrxOmmFQGiHZYkh/9f+939mU
MItwiGDfzILj72l1eIirnS/9Xaa2IQDpm5MlFvWKf7mNjqrTJLUHhSQL4o1t/tedn77SEqsW+I05
ujS9cThiuiULwRLUyy+kbe0ljxxIYNOagH/cd8L47XmfNS+dmUe4L9A1CMLC61D63A5VIDsc1aW7
55t3n1oW/RuijKOfQeuwv8AaiqTAh11XS/S2PGIdaM0YZ/rdWqFmke2k7OetiVadmi2dtMNdatwP
D9BWHcxIQx8+wWviqFAXc00dHIMdSSTdwY8XF/Gyk8pjRY0i4W0UfTbAb/pBhgslTpfeKwVqvvbb
nmm/5VEbQyYi8Q3cDIuwgY1zsvDAVxLYJjI3oQl0bW9EE2l5zouohpeyuRT4s7vgtwLNeUfbehzN
NYJwTvSp52SdrgpzbNCr0M/SSjVl0TxwqN5+98B5kXp1e+ibsMVZ1rb+EP3XT2zwTC5kIC8DesFq
izzhdz8Vkn5cMLS9I7VcLugJd6cGW9yQETtIH/GE4dgFz7u6U7aYaS5JFGFKvDc9pxGSfzMGozhi
VBbDpwly4s6x8u3DbkJ3MwT+xD7/ilUicgG8wTvXizHPFKdzOlw+GdepvvY3SlnljReofA8Uk/6L
np8bvbfi8tVtVMlitzbcIsXbj+YYjSi1D/O8XCBEuIX8fXvpUEb7Hn0gW741KX9c/3VLuF47/NfI
x9GeiX2H3IXaoqVLHj7QasOxjifNRCRTMOUkhsDZbKFOzbazQlvgLB1HcN8N+kf9RzxvdjDdt8mJ
DcAz7Nnkt8QMd18hg7CbufEGaR1ABP0xz3cbNT7mMkVdnvGvwtGCwOfRGUpdVxmjNRrb7DDkY2/5
J/rX33wafz8d6mkb9KusWTpX0TJaD11g0ts2eX8iWSIBi4JC0mAce0R/6a6EkommZ6Ta90Rop4Wu
9xOmINR3jpoci97i6n9ZakyKa6AK4utHUbWTjjwFXvqT09nl4MKq5JYOH9iVJNurEqh9XcRymw6/
08/aALI8CJRRnmuWxpwxHfJgnab9MpN9X4HWXyCWzHCZKwWBWUzHgmkKh6gCTg4HtuRkg5bju0TY
G6AqWni+brpzvMLJARSYuM/6aHgvYJ/u9IeZCid2wv3gUUbNB0KXShbSyazYVddCyytozdfrQtrr
7W8gQzC7E/Vzgxab4miNjvCNiADzJ4Nk+5SrbaWI8VMS/pYflHo/01dJ9peSsvCA40svrADEPHkV
p8u5GyVNTMCSQ1KzdluBVDJafaVpNrCqK83Tx6rAl1ckzDDIqGOGALwlKTl8yEU8+8JFbuKTsS4S
HbWTHuYk6YGr1Xx+LljLe+ysTxK0uaOjEm8nBXnoyWs1PNjpydVrV+vTnlbrOAxEj1InDJv9dX7U
6QvbrBip4QM4yLxtGLI5hEzkM/cEi+5xWJnuLmdxwaxtQAOqE/xhfBEVMr1BsDSA2ugVi4DX/JkR
/HPfhys0Te1slk75ktdIMZLZmp7LKk3ZAiPJoQRJMfZxKbyTpm06hlPGJqlHxAUu8EOJ4MW6Z+12
nyJjnZJoAMwlitlx+0cjTZjvx4IQhb6jjQdAkq7C0zfoxb1vBlD0qa9AlJejwUwbP4koLaBJ0gVq
8jasfbHko8B54oaRspjPS8r0C1gr6HOSQ3M1oY80CelgPdOfefidMZ+ffWornCZmjIWVDZ55aHbV
M8ZVjd4btrwE8KzvLiy7BYTyRqrXFnnxT58xBPP+toxZLKbu5CC5fi0crQuLjgPtoTAXKn7Q+6A/
UwYcp4yoK9xWSmLijoUtFvW9cWMHYN4SDgy8cVNlw/e+FdIN8Hra0OLwOe74kqYGYqyRwTN6reoi
SiFoOIKtkaC9vz2KWUxQFMhuvil84e8yolk0hYhR9L3cgSIdO/P61jHsLpPSpyYyzfjrwg+5ue0V
bcUs/e2RM2i0MHqB0WqLgREjxRVMI20LCZ/5mYO6BXc3rSgGBbrMZxyvFXvPDU5S8WeoT+TIk9cH
JSIusFOlDtgVNA1l8ldYcouZgIM+Q2TFExawuBfVMF9dYBUAV76Vg14S8WB8wEachK4b0TIANLO9
/37Alfs8U9luK6eJORkhVeiR8UDQjKE7x32lwYs4XuKPCojT3Gsrvbv1km4TeHwv/r7W02bBNUQg
vFsy5UgyaWoIILAOzwKnk/PPnRCDLqVLj91tmV6AzkpBwvRQlfZYWq/tfXgOF7w6StYlE4PI5U5z
7YvQ4ksGrUD+JJrQkDC9/vbERZDL3ea2QRqZk9acvLfE0F5br53f0dKLNNvXKFdEc58uig5uo2h1
CX+j0BCXfm8/MtX7HEChmNdqb+/hQOIF5b6P0AmCTLlW+0TVMkEk9akDe30f6/EpkJOdtR8O4C7W
eHe8vMxOcpAyWm2QnUNAEiuRr8JlLSPCb1pFsjGojqXSj/D9tZwasWMa/5FiUMW+IjJMenub6vbt
BDjSdVpd5RBObq0Qm36zsOEg7Z1if3Nt9E02vGvHtSfD9CEqG0Zqdj5gWa3DPUgkkrptVEpKzjKC
+RwYwIovBOgl0sW5RjS6RSeron9BcsppeeXCTpSXKH0weDkEPlFmZ23M0iJvzBPk57BbfdbE7Lt3
S860/9g0hjdcFwELCeY4tL2VjjngSo8H++2VBCkWNRc5SYQbTwLfOy6duf7AXZx+UrIWk3lqChOy
nt7pVxPfsOIuYlzpzPrH1aJTJ1rDbGagjq5ltrTSG1S8CVEnyGycRh1rEm1JLmKTvGi7RG/FMcPS
ynn1Ol5/bR5SEy0594OVuIZWvt6aMsEo8UqRBiF9OzPrmHeY5RDdeyjs4vETn7Zd62pFTqbkRl06
mUyp35QcQPfjtInWnKJ78td4mtuhWBbUgSISb6EDY3kmhCbP6jPpUGZGonjdK+Vd7hFDSsq0V65Y
PjjIW8ec3fNyQO3Sklun3LEjUXNZPYguLPZC6Go2gYj3DqfqJx0ToIXgeZhrtLT4XY8xZZdIQPxG
browJnZumMQaXhW1Ba0FlRRUW/7zg+hXW3OXVtLAfs78guE0oY/PGZukRRGodQObcmGkm0BC65oq
ZDgCHdgOfjd86QOtfYhoM1//KjVAlcYUBSilECQ37ierZBoZYNvuYyf7T7jgtkM9alDP9FPphv5k
t9e3JA+FUcnw3rVf5ipB1fEcHTVCTUkI061ddWf14Kc0Qzn7tMPTsYCusDq8LzQdE9Q2lKa99MY3
MOOwdiLaK4dP+mx3uWk1BPgvjLpkC6aJOj/sfV10MY4cQc7uM1YqP+AWPeJZv/aznFmVLrqTEXpl
nXj5F/bxeRI0tTs5fdPs3/qzdbfxkJyjTjqm3x8AxOCdS2TI6oB5VpHnRXa1W7cWck3Oy/JazOLQ
AyjMl7Octd7Bgr5D7he+VgAyJYBDHnQNPv0NsT4qlayfWDHH+TeQMP1KbcutySiufyJ1CYxUIRE0
waeXJbbzVyndguv6L7ZljYQwUfV0p35eL2DSbHlewRhd4xIaRNpsrG3rV1kt+hiPv6Ajzw2yEkoK
xWxC0aCIL538OPbUFuatU7OuHJ6kmeyyF8a/OiCXSm53v8qtJ8lLuqhPEO5e1zwc+441uIh4kdI4
jPbB/tGrFSTttAlNFfSRvJso0FN3xFDgkOxQi7n6jStYBxKYQTApqV2aZQx9un4Pj7YCcUp3eaii
ijceeF6jlOBxgwBfxaZpqHy5cgIAGHGLKHwUWnpbR2ziHEDsww/g2iTVMx6FvdiKo9DM5z0CZ3yY
ktONBLVCVv3oE+4K37HP+N9zx2YicraOPqGK2DWJ1UPTr/A6lFWxBJdat1OJDmWFz1Ek8tDM5j3O
vFWniRtM66VArP/ijJEYkqSdCh6PERkeGRxn9lakWtmlb2PWvMh1LwhDqRFBize6QNCrpZRAyqbJ
ncy4zSDpZnXS+8wW/XdzUtPXZ/yO+yRVWEFmMox3c28TUtFo8WuBfKIWT63ynXZi7MuvY6V9Sowl
rmGB9zai/I6JbtFalN7DGSroHGwFqt+6frXkKcjqbwNiaaHykArCyLHKzGV0qhht7AFQA/aDhqiC
JismrPvHpma96rAvWb5q2j2givAt98R2/a9Pt66XQNrdq/+wvIFr9VgLD826gqhNJf33/HDmvovh
AyDtMdo9R+pQpGZDJihNw/k7AMG5TpnO07+JvmSShhKRPqp24iuuV7DgUQ3dioEaCOhDLQobBY3p
jGVNcyTllM9pP8CY/j19A4Vmep6QKMm8ALy6P8Z5DvX1g8MqlvadzhwIGu4Ss9QY5ey5ldBC6F9h
mQZ51CtP6+dIxhH7Kxb6hRE3NedCk+s0yLwQBefxumnh7AXvnJqcUfcpM0rwKeFyi7A5fAcyksvU
D8JSuY8huH70SukUQ4i/2NlfjSlWlqiTfXyoB8zYOsD9G0daV9Gv4ElnQeuAtdpy4nT5IZVpECiV
69xHOGasoFm5vF/AJ4Ob4Nu8YXA2GFHgfbT8CQHXCuu8TyLL8+xr352ta2HAIK0TR+C1YGGyujfU
d0acbquZG5ZI6hBhOsOMNnsnt1zGRD5T5UzxPfKRDSDYkqJpvSkv6k0HP6vCyZw8BwpkwZSDKFjr
ZBVeKr09WWKuo53yvGhILPUBg9DE+CFVqQak/AjPHsD6f8xAQOw1y6LgcUbxsorZ3uEx47GEpfHa
XAJW94OyPkJPlXV2H7qj+kR0kyPhsxcCOiy2OOpmcEAmNgAY+tggwBRYyUtvbw4cpZsEF+cugeJr
WGptmyiWNGsFCiDAYLK5dak51610iVTnXiC6TsOizGAVaWHzpWYg5jCQxD9JVmE/o9Smhfq9BuVB
Pkcr2x6W/ToGM9vhro1u3LsmA1DXzLFrbI+nPjuLS9ZSVE+B9C0v2zgocNjCzbYXnoD7/67pLhdp
xQgQj+y5kTPQ3eYfIN7jyPmoyAoaMnk5ojT0l1LtpUK/MwNoDK4aBL3cktHe0VHH5Vg6FqOGvLT2
JX8L1HVL0JaNXzvweMcNCmoLUSyDkA9pVpI4QGUGzU37VjD1TVAF3HItqIsnYHoojaVerXOaJ4aM
J3g16/kA6Q/BWbhOuu0dM3o9najHqO/8iUVPVHEvZTcIhz49EEfs2ibY0m3RVpQCXhwVJRkzMg4s
hLn70Nf0vPjmyIzMMrgXJQ0lqjPsjgcGg2xsS9IKjHeQx1ycbJPEcuPwBPeGvBH+QATotL17C0E5
Nu4OHJ+zEv5ayaV+GKdSU9xDWjT1FDNu6iUZs1wPF4k/NempC5ZKg+I+NKQgVrpym1FXCTSDQ5WD
j7HDGWqNvomRI9c7e3h2M7bk+E8eIdcvGg6Ve3YxyYfA1Ui3pdT+sx4/LfqB2UFkoFTUBtVsqfoA
0dIayXmCbTHnQ9+5uQsJtfKLdFbMY4XJs2pxfcOOJM5ixUMYHMxJLE6FrpVAFrx8vTYZANCQN2/I
Mg/GNiatboW7CdwOcUdHidp2NHHb0sfvzWiajSyKiCnjXqT7zM/cBGAuEcxAFZdNTjbRKgK7SpX0
nWAsvCT59ySMzH0oHkPHA+/P8HipJ84DJDLynb0LjMBLj0whvXeugkUOUhjCSZSCUCCpSc1BycSB
4RBvH3dvq+gAK9H4KFYUZbTK5b1yyQ/+WGos1SOw3pFk/nK3EWgAx4rXbkTi+adMCcgM4+Hl6Gul
N+YpggBfH7Wblrg7NZ3xfT158GK8Entob8pdCsUFsp0t5Uzgv/np1QO+R/sFqdUyDZJKogJSSAu5
RjFaA7Tg4MMPeK1VebZgjV4PfWslFwfwVA/rdYbuKmtqJ67ZFUa0HIOQpo5QJvYeSZ3dt5yV0ehQ
Q+3t56niYCSzYscL3ZXKxfkncVBgQWmhbD02WWCQw3Vi+QN6xMGOzyk05dD6NzwGISIk/og6Sl42
dCr23YA2VD9rOQcF8pSxCoiqTGT0eEGbIMjleenDZ6TWyBBpeYd99NqzWIfsJ3R5LuH1EYPKNDa0
uOwrCe8NXauUk0dlZSan4yf/brp6zMGTlo5rEr2tE606ntTxXbnonL5Qsmn1kM1uDKNHjRwZD/kj
3zFEZ29NmJZ/9meOdb3ZHPHEOpM3RbHSfYg+NQFYA9uSTlVA4v7pe/PzgbFfhewhejaK7KQbjWk9
TvdHR0JZNaRe6D+QKU0Igrr4gP+NZfkvBzBNJlysbkH128ooh0aKe6bbq48zrBkCNZbUiWt8xmrE
RxEwiT0N+CF0kR4KSfODi4cmL6Vf5jGq2YtvJ/0BdhhycppgmII43k/eq8fusxNraz8L0Gf0z+Nw
EoZ9ls145o54ff2npTLWwBDHUBdtyvkqfcSFa8j++do4smw8R8Q98m/PW83BFgww/PYKvjvS2CjS
F9X//0rWOqQXpnLSJ85ABN0mMf/0kCnXKBAZrePzAMXBBHL6Wenf6g8Ipz2B4C/K1BIX3js+Uucx
wVK5a+BlT2vhsq0kjasQzoSaV1ycKpnAVg3YFnr/9ru2+4vP3OIJLluhurCD7jWe7yiLa6zA3PRG
AhQaEwsRwtMK6rz8mUH47iBR7pvT0GRMk00RaWP5034oySTazl5mfJK9pCCpw1i560VBFw/vT8IN
4h6Ii9KJqf9v+XdBlYxPonkFA8PVGvU7VLXC4UkM3A57+AgdBIDgW9SlM24XnO2X9y93wSCgw5qn
gWg/4UjGJapxTmdle/AgqYF8YLy+34ok5p7iLQIC/3S2ABb0Uy6W12qwsaCJDQbQedwgl6Ohihux
T3pntB8UFaU5sygyn5Mo1QFWA1cdAV9u2K0JfgOcQOSETgwP5KhUx48eS4ZxUF5ungtMBLjHJtOP
9uj0r3/aaT7YCyQuOCOnqLHHQbfFhT9772Zq8rIYRfCM33rnOTVWG/qK71sJEX1F58kIPFHqU69Y
qN3wm0n+uexMU/6pDs1XjBl/zXUXj3D3w0RwA98EVE/kfWXr5sFUmnWYgHfT1+L6h7sKhMiptN0N
otiesM0Qaue8VY2UzFsrGJ6lc85+0dkY6AhRTw87LhWsrBKRkE5IJPbJxpg97th9HNRnoPufBZQQ
Qbe71bkiRIaF/Msgbpo37gFDD0j706y9ilK9KuWNsygW1iIMtrUMqv7125Aw0qW3m5nly7/TN/Rd
jmh6AO7J4GoGnoDHVhaKeWJOgMz5kueuCnAkKNsfw533gvZbJVhaMrhnuXeRfOGh2PNXoSweNbiH
Nck0xWheTemBbcsw8Z9eBxiAbU7g5HQqlW3JSHgz/8HY7ldzyHGNwMMidlltgoquRmcjlbNlH9XO
R9mSifAfF2leFqEWBrkPr9yEpqxwpgRG3N5l9BUSEJ1sr79zzHqbFquyF7ngy9S7x994VCs2Gqsp
Li4g6XQAagMvaeospKFNBBNl9CAfaL0EsaQFD+7dt9t55/rtXQvmtwvazqvtwRR+wdK9pp20y2Re
EXbfOEVhPXCOgvyS+b5m3AePqdu26uuHGuktC5tD4e5RmKMJ+g1pkW5tGzj7auhDA5FJlRtu10/P
G9IPnpPgldqCw0NLppolDm48MjCaZJi4UXiqaHADJz7Iur4oCgqyDNC2U7Tedf+TOlegwpDW2rlL
1kK7WNyEAR7hsblHCyU/imd4W7BVL0dATqMKplBn1YF79V2St0O6Cg5rrJxDiX3gNdkZqYIh/Jip
dIvoGCC96h1QqE7dyMEW6cURG0U7cm8FLNbBuD4idZlL7lw4JU6XVQBaTfs9WG5icaKHAgTOR9ab
ZXaZrZ+LY6t63dm6zsS2QgkMFkWRg9hCIzIe4l/w9elPQ2fk1FYZQ0myQm6Px8dfZnMasSVa4oML
1EfJCqax2b0QwaebkXdaM3j8AxOE0Poom3d41JsZlbmYPcqUO1arKt1StR0Hz4R+68eEHbmnB3YC
6js3+SfOdI5Al3uIEQezXoxIZd9A/giWO5Wh2BsUvArCJr8GCfqVTckBWCKn1LWrXro3vQfTQD26
pMR1p1hbgc/gPujIEBUh95VPztMSgtJCazREX4wjCRlMTR5KsNJYmp4mmn+AAC4XEzYdGq7XJIkE
LxeGI+J1+U0q+2VlqetyNl4XjtoqML7VyJBKCV+MaRnU7EsAObi4D3vbbtHUS0OYCPjONiogflim
YKJC18bwru4Dj8wW8qZgguTzG4n5ChhraK9d0k8RIN8g3IYPTfcf7muhGKuJgFpo9w0oPI5vuYW8
d6q9HaHX7Wthq66rZV6dkdo5MbL0wKJkjlGazZ/VHUCuQ1rCXS7vrtx1nFkASKSNeptvCGwSbVqY
kxkHwlMcM1otYQSQ4wdaphX7eA2qj42ta6VgFirHo17YncaKn8fd87FPQo6RaADKLrU7zRW5EaGK
Pyfkr4/AG6PK6PeW02VDNlmJA4rCE2MiQ/Z5sbRm8RL63+8U2GCsOdk3l7koisx1k8vqJPqGtbdl
Thu4Mb4nuUZEkpCz4tM6rqGEv1c7aSjT1G3jbUWR79JcQuM7482uXRKInN9HMKgKpfbbiHV58Oio
rHr6k1Z2rTXZE10QRN7umycbwEUAsHfpJfU42xY651tXu5TFvi4RqMVkkEqYYSs2Tq7h9QELFnFP
56bheaiLwj05VLrX8QXviMYxIN8wuyaZps0dnBDTkcGaMFbE0ulA/cd0DR//0gNEDY9LBYkp+DeW
ZuleHGOhsZoeHh+fL3AbS/Nif3Sghgrb7Ds3EpC/bLQuKglC5Cz6aJy9p/RCZCPiRKyos15LEOiI
XPGLsEFqXvau6KGT/9H933SXycS0RW5bsOvmikUXBRoOjuGLjGnxKhtXIKT/CdNZMjSSG3HPqzrv
EraMPb17w7A/tlED6DwlhIIsqQTx9miHjrXcrbgGYdKKPWm4mN9DyP7Tw2imR+VI41vzFF6lwXPm
PlI4/jdWgjhqAmk1K0IgKWvqMmmxioHnTLrFWljUh1CMNZsrcH94XEkLMqS8ioHEYgxTnnGZI43L
Re0QSB2uhyS4cuvGoOYohFt2sRKyhy7wBeMlf6fwVN6WwG42dsSx6G53ooxUZS7jlbbz1x8IXGkn
7km6tFNP3yZcuG6+G7+IGTol7ZrWKmfM58s6jgVv5JNTa5K44/HklDK0nLvmk2cJ6Xj91RKAFs6M
Hk4wip+TrgDNGwefueOV5TfdbAdExxCkCamyOdGDk7BRSEUYO95xnkbSy7Akwv8ukgdZgY7wgRxc
9IvEWu9Tz9tDHgY8qMZUu7wGJc6Ps7svtn3WNkYRcYlbHLsi4iJ0XxZpDcYnwqoApvEE1QdWc5KG
nqWRiALCf1RCaI+OMdaXnXefn/ScEhFIHHv53cIofRx1hlhwG0PbnxjArEsDjbxl7iTlFilwLPdC
vYQ2yVEW2GkyX5dR+7x0qodfoQV11/VXDqbzl3NcA3cpwKr0QwfHUtX6B8bmunlE2vNbzNNPeicN
4QRfFfNS9XG6MahKHdtN2w7CbB4aw7aFiDO/nd/rNmL62BhBAqtdXeZ9nEH1Ojtq6Qf3NxDshjzI
7mU5VXt/jTHzPv5JKdsX0QkHxOPVawB6tJmXMqsb+DNqEF8TF8JNz/H5D/uq70boaJRI6Llw76tS
Nz88wer/3D+kJ466IHKBnQR/Thl0f+DS0XgMDjC1ArNY68TzcELk84Oc2WjEZVdboqSQmCZyKzJ7
OtCFCezOki1cMOHUeE2WQVOAFU0xG/HCkWH83jI3dkKjCD6RgjhFsAu0mQnYxu4a5DU8SoWHFfyk
mz3+cOPQ+COraZz9AFkn8J6+urUHbSNTMvHvj8/UHaS1w+gsU4l8dfAUoCGiAXQhQ9nH/GyuXJq+
lvJTWikDN2CwXVpIy41QZNI0kQBRU54WDoHZH0STl6syVK9SJ2ijMspm4MEpkY+xIl6EQoNi8yQS
emGZqKDp1zc/azmXA+iqFziCp7yeI5/4H9dPVRjnXLNWlaZgbymfSQstJOzcjxNl+aCa7ZPfuJqj
5/7FtPz5FkzZNBSxoyQSBXF8J6YPm5zqg7StHLmJxFtu3o7zdtQgxnxXczV4qZawGzdfvdCIDhwJ
/eXO1CMB5MmwlXHkwJ+9GLg+9vBWbyr/+SXnnTu+Q0nTkGyM+8RyYuMXM4K1Jik0ul+eB7W6hClR
3tqNfJ4XxnCUpsTA6hkwUqOCKoArfm1g5qT/VnQ9IYCB/nXsD7aLQk4D3N4HMHAORzAhWW/fa8xo
HZw8ne1BToURSU29+EnIzPR4n14IopvcIKrbfWjqRnNgNpD/Hs9DlLLtRwfw0+DpKcFBWOjgn/aH
tC9zoQ4RYQ0Rj55+Zy1Em6qmojcRrBwrhdMHwP5+TQ72gXGLdD/bCmeOwSU3gwl7q57YnkV9rsBB
sa4Cvan3t1ysrwOJC8l+onm1ZVdCa6B3cGMWbqNwDd63ndVPEFNUbJPld++Qev59uA/YR8O9o+0o
SMqj+XJXlt19vdnGDhU0lnbw9svkRLiaku/RtTe2u2Df90n2HKEOW/+Bx53bTSSX317n+WjziDwE
ybSuql0hPBLwtI2WHfXDBs/K9FvYeOmTXGS6bSLHhyDlevFabej8yNw/v0jYWPDEXd4ofXl81N/F
swIjRSc4UKWrjmh1dIAziu/LKjHESjvdpYJo0saoi+LGcrcUk3grk1PDdBuWaJ51YJPBKphUVKNx
oMDphxAFsFrwYeKn47IbQhmg2lC2Uum6iz3dQon3Nobbfd3jZPFFgV2FN/dKky3O7vnjFXrtzSVp
VCPLNzmZ0hXwI9zmASlUiJ2CO8QU+xmssUMi+Yai4IYu3qPwuZgrprpDG80DNb0MJcTy1pSZM6ds
m16hjThVMkp9yfN/0HH8xmTtvJzrGC71JVtuj1ULCwHKSi+9Ng7f16QPyIYiND5Qu+NXzvpJlYBJ
inPOaJ2Wfpfuco1AoFgfbt4ItdO/zu7Dnl4FNV/ygHFgZ/6P25geXMqprg0H526oF4leUki+W2rv
kBDB6DbmuZ/Y66nw0GQR0VMTpyCT8tT7mjqGNKI0EuhtX2nxdZnkRMVKKkjo5rAqPosqq1VNWaNw
wrKSVjxnJEaGa8C90Hikq2u4ZGdS6EuAff/at1kntPibDFkzNiyH5FXaY2cjdsYOSVmFljHiixwu
TH+BIPM6n4LyeYtzAO72XRBcugeYJkMFlmFXOu41S6rsTFVXOWN8HqZNOjS4e9zgE8MrIF7vqCkf
rOLoJwlM2sCrJv/E9h6oGG2ir2P9ZeWrp2rG8YC8qZpbNPzwMvNaVyq16GW5eQEFZ/jKFNGMjS70
iH3V6ih5CLAjhoSW3vLCt9R8XMCUFfOFlKRpF3sP7EgWP1KvoH21P4SpK3f69Giv3rlaQr44qMxa
kARdbmQPzdmJczHNFQX2rycjeB007CA5VafcHxoSxrrZAu4vN+ai26IAzlcdmJjFQRhOxeCk1sx6
QaVaoqglRzPKjC09gm4dE+9Fu64KQN31TzYsY3GrwNeVfSIEgr39/oULmdxed2aRaHlfM/XhC6Zi
K6BdQT21XlfL7POVCzixEEBP+BNTbuGp69geWgFNsRjh6PXuf4QMkgn8PJfoXKOme9C5lu72D/wt
Uga/PZc7cNYyZYM4PhLBUDup+aDvuGuakbdWBFg/VNJ60uuCHzah5t4xeYzN1QjD6CLFlLM6/Acb
oeZnCXlZKcs9zqJXa+jU/sZ1O+c/h4hUuh2XfLOemdxHuw9U/nwkoXihSn9vx18h9WHkGuTdrVfB
gPpBEPcfX0SzhOVkDPE2IuIawkk34onlzcmDCvckPLCNY5j5tYgYTtvwucVCDphJ0c3q8IOwdiVS
vuNIohKWTtcmzWji9jWOYkhxtgCSw4ebrn+X+80cdUevlduc9hH6tVG6VlgsYobWR5EIazjJkKCO
mAdF9MyGxNrg4cAe5Ij0xH8Yz/m4Q5WX2dC8xj8TaTD2YlTBVbvE3f1u7vfLyszLWlM7Eng7FJ6J
4blAjueolz3u0gVmCfSvKA0QCViIQKNnTT1c6HO+L/8dsn9t58pA2kM9zKtpO30hdnkf25WLWOxr
chNxBUvhTcy8uKJqPx0beAvotnj8cVCyqKSQXtKquobYuWtoqJQ6KeYoq8P4DQNexCPkSkPm9BG5
f6p0gV2i0sGbuo//N/M5Ib4giO2/AnAV7UNoB5hf7Gif68zIcn189dEg7mkTtOPOgpjHVsbPxCEf
F6IuHe/5H3fDJrLxyVwfMFoiaIGiJJldxtmSAP6TBEauXWhX2oQUhAWcA3uW3WmJ7G16aNcT8yHV
8HLnh3DhFYN2tqILPyrWGk7U+eUT/lP71Li9HQ9c08pe03gzPgrdutjKjGLC5ZwgC0xbesl9GxRk
PT8RZZDFWCmUYeKmZVm4hF3FBHnVefiZWNzSfVywrhJBl6L3e0rHDj/GOQAZOQWhXRxuvEoJFnSA
git8dICe+PtpR/W7A72AOACzZ8u/A9NpNEVbgMrVauXu1lvrXhWsLrVILKSKZr6fgpOkOiVD/tAm
/+hKhlz+Z1jON4mRhy8tjn6mxH1JKXcOVnuGMVZhLAJNRV+B4k+11BO0ZIsXtAd5kN7WL5QdlFVW
S5jP71LVj9Td5RUEsPUdbj4QHB9Rt0RAMnZJ9FgLPDqHQHJ5grEM4VXeaNWZ23hvQ2gU5iqLmVEm
P2RNmEfSNwnblwbjuhfJxyTFL0FhKLZfLijrviX7UErNcVwkBuYq5EUCB6Y0QtRsdjq7w4euDibB
Nc05hkfObAohxrlrlmpp0Ewu+P0OzrhSD9nKJuG5K0D/jYKci31ylrje+oIUQSHZuHwrVI0Lxujh
RmLYW3OoGXX7bW+/3PFZESwM8bQW2uFYKNufeuNw9X3DPXrtnQa8cxmdq4N4q1NL/jB81eGPOk3d
6FGI8I5Pw8ipeOa4ei4F7xTdgPuH/b7hrJliSnjh3SMh3TrM0iWfCMcn2Y0pwXFCJf08d+WEdCyD
pWhR0NI8+MHmFHMIqv3GjkBS0ZHj0Z/zYiHWiyNPZz5rArlMMmUh0MZs8hT7hlk3jptTEs5YxyOq
rUZCnMSOJbOFIZhUA8lp2yioITKEhdiTXne69YIXrPArzADRli94qkcsqFM8bQeNziXEFfbh1AUr
4gv9KjFJxGoiOs+AAMJ12SC9vmAhzp8I4EI8U/HwQAQB5U2RgN8arv2GdJBmv3hSzlit+FVrBzdR
kL7bV90XfbmjsWdFRQ5YBHiTiA758650x2tB+wZ2f+Ofgk5LTlq/b6IJMVgY4GB7X2UpPGgg628S
D7SWwOxFHEG4T111YEuuQJ0LIdXtj7kgRdZAd+xExsy7pQ0GfhjycbeHUGmGbbC0siGFoza1wnS1
LH/ClbatMetl9O55QGJOp6PrkXAC6IUbZDRufpaq3y5hsLWzfhtQ7uPZjZgj4FGBx28qK+U3VfOR
bdU7Xa2IVdYGyFTpvswCEr5genXJu2BtydZmmG+e/Po5iTsSJyl74i1HkuosJK5/mAyjXGGRBukG
tZv4961f7qF4w2b8hEUDdjM2NUuuW+aJl8dgJubD3ypsGIpihoROHcuYGwRt17Iuu6dZq/for7RS
VFaaEhe0TpSpk1irHNWlHhwXLiZ86NtbvxyVcEOFhdr91Og154IGBjkEHtKmN6DZ3dB6Hf7VXaRU
Ft2M3TNHvfwAELh0vaASgFvLXF48erjrC+lSF120wOyUxulT85Wiq2F6dMI9cjn1Zmxcr3L94JJB
OiPKtwLEMru59Xsp6wAXs/bI2nW7KrfZCPmg2uhvmyhIf3Ay4IO26R1X18QnA8N9/T1pvgOrkuna
1tuB1Tf0jyPjPMO5t9mOD8zb7H4zcRlUAPinExpiR9i8Iwuij1ESnOkS15Cun4fW7CPFj9OMYdWi
SmM/7qXsbJEit2kdAMcbrSm7gGa11Jz2yQU4fiEEdvHzCbiWNdnl9RakrgIQPGaxbVFYY1WxoK22
kdXMs9vki3fBt20GdZBaWD31JnFH40dbNRBtLTVuMkhrHanjLugrc8Pl7G5JcqcT6pBtah9Dnx/L
93NGIhNn2UukAEOU56+U2A1fL/qqsY57YmnmhnRY803JfATOoL7T64y2RTyZ306mPO4l3fH85f3w
rOAwLVumGyRYUIyUWCLdH45al/1R8fDLE9lmVPInrCQ+oOwb1i2vr4haTn2lBkQffHcoyAC9uAkG
YHGj512kI3zQgVO3LqUNWuZ0qW5HOjB7jbFZdoK9EEnkS7Kzb6IM2/ggyI88ROsrZtkQ1RMDqsLO
W+MDTfcq39z2ESFuQLwCt2CH4s9eM4ltrDOtWj5d7DrPrNrKzjlVQ4OCIpGcawinNsg53P88gDjL
IzDCfcDcl6Q0SVu5mlgoNwJmlmzwn4F2KiuVGe4xNmoJuRcUw0mSFF1XL4wt0yWlZIKX6hKAMgLn
z9WdMwcnbByVztQVe/3k/9+zKibkr8Vqb7eLHMz9pSkD4OagR1EHE61QpQUU7b6OFaOv5bjZddev
XS1Xw2QG+pL5G5BcPlgbRJylLmGJVxhepvNl+xYkK+Izv6htEEvm7grsgU6GVWSd4ltz8hfFbjRp
3h25XcboYv3sGIobysN5sOb6XRMDqo8Np8bvXzevjYIPTxpI75yvTUOY9DOnf4b4qGMpfHnsYBER
yc8Dz4dtTmZpnnioVJlZ+kkcxtMKhFOFbow/RIwx5EgoXjDC9sVyHH+HRsqvHJJrybxjG4viMwx4
ZN+BvpDJ9VcY1OzJjoHVIFiew4clKpVJi925oZ45ZvGrHNFO+Y/rG53n4kDTzjIMdgeYdP1y/LbX
Ngnt9PeKYKP6YHBB30FxUiLENj6Es2cp6t109VYnScnSmks0t7RcYoyboC7f3EGjub0UjjsgAU3N
C0PTUEvDUeZ/fnI1YwpaemCd8bmsHvxao7S1PHjC9TELDqihon674FoLXgyfZ2oEdE1/9On6TBjT
Cln1UBf/QoaqwMts8rZDLGnGZ0xcfIR8//bdBJQ8lvGSTAo0udDKBgtS4LXu1KvQfdidWW/D1EWt
pDUYTX5nhpnTZ7oFffrV7IattNqz+bG7fMai4V50Ibh7tF7zlUArKZ+QfMd6Po8osBV74CTY1Rvf
t2b6oeAGDjpuLj1gDHOsU4lt4H1C3Ea9OL+JSv4xdyZyVz/OFvpuRcyNj2fHEpng/UcNmIyVqccj
duexHDMXeK91Y2GdQ7UNt8ec8ADlcyLTL0L4bbEGETDv+EBE9zqiPvPuAfX9gnSJCq51CpQiwgfR
Hqbbv0RH0HApX2w8hO5fhyZ9Nj/2x2pqpUZKN7CRpulrkuFNUB0wRrhmvf8pgxIrh1OT5IGG8ERR
LOutueZrH3lRCfWdFnsey9vG0yMT1kfRqMFJzHmC8EUof6atKUWuLDBeJQoqah8S9xMSGNezCSP9
LJkm2UG4+mzzdXnOr14bepkjz7MF3iHIuyFrnObW1yGjpxEjolztfHfwdsPCxOGALcx63N2qVDor
2QLTjQLEdmKJ8mrgoKE+YooqN+paojicOZ2CWX/nZUj/SoH0GSe+SbCgHzQ1joZ6wcUbONoHnJj0
a5VwMU9kespX57zKyY7grgBZsut9W039SpZCrs+80o813tPWhlG0uULoH5Gs+nrBgsDsFf5hqoEQ
QHC84iIc8IGI5GSbdK0FMNjuA0r903gHB1pnMpIqgKp2OgnVexV+cswLgNXXi51IcSBea6pNxkTb
Dj+nH1J+bdnHBAcOyULCj8uk/sG8FZ4kzMR6x10gWtU5elSWGCQ3ik31HFt7AYYkULhuMsGXG0nZ
TYSFGZkg1H04EINUPdEBggygvtmUe3mUoGajXayWrPh+QKNTTuw1oUx+daXKEx3HCpQq1lNk7iHl
9EDltP2MJKSnpzvdMtyW2V9WX2heXIrm5isBSG9SP3oa1k0oNzP850LlLI1ROYHO2qnLN9og8lrL
8nXWWf//jPLuELmfJD8ZQqScpAOGypQbiOGXyupfqCcGdbExTNh8w8EaVDfsfyTdadOIhJXJDi4J
LnfHCh02FzFiA9hRhhruGUimS/Sr7+jP5nStsGtTtdcooegQiv9QXEcs62ARuHeRhq40bbLG0LmY
1IcwQ1PxkaDmu1B7exG/yjpxpOkV+BWaSFlXf2+vbz4HlRNqngqoKw1Fs1ivclaYx9I/NIlV+hNo
FnTZwSPO0lS/QddKRX9eGCG/N9q0gIYkJ+ymvsHS5+Sy5LjL+xZl3IoiKYH5HniU8CR4Nq4Hyxp6
fKprkmy9q78cEdZsa/5JbxPfy+AvCzr45k+jXAHZAr56qJEU62cJSlxtiitOo0Ralsc6XWIL16sT
pNEPJqOs+rrD+B12NSbAAO8KornqOmHsJYGoGrKr28rcHzp7vGm+d7IwwJqK/WNN6/kt+J37TU+p
UQJjGYbYmJZBSZ8nbEd7ixPCsfqUYy8+HP/ehGRi/y8Gepj/o/U6a6Ys+ScRYpf6gnePQ2r1i/Lz
c0HtWkSq0gB044HIpbnPqy/sztQ300ttIlr8fe8i6vU9VJAoeBq+vdMaFwnP31ityfioIkFB8xxy
AGQmFrc4HhSEF8CcxIZ2bDufpt74QzDhqLgUgHJLcPPxjgqNOTh3JrBO5gbfzo2DYiyIq8OAskyP
vImWoLHMw+7gLhWuboiQGDYea0MJM0ZksXXAvUmEUAp6cUNOeMBhqq5d5I7CO9Xd+4x5pfyt/owQ
Uz554WUSFDjVk/at/dcPN6pPv4txJj+Qre71LHAJkIZJIIZyu8VuRF1f5bfQn2NOm0Bnk1WJ4BJ8
KJMUtt0n1RcLtworAIf0LiXKxOowatBcjI225kxHOeAtoDeuR6ARYNvlhtsZoYpG0qDyTCIkM0Dd
uXH5wVvShRjMySOFxWRMmv1lnxC6fbacxw3F/Ns6ckslNnThjQTYle7rKGAu3es7/OFjXBe0HGd9
r8sKsa+pWttnayAO+1aEf79f7Eb4bm6UlYvtmRNQsTHfAyM77FJ8Hs8RKl6eyUZ7+KBeNeX6ec7s
cd0ocvZ9lCrCUgnf/jXLjbtDFhx3Dm6kMLnVDgqPpV2QDsHQmo7sTS2qI6WQKP3Oa4YMudgYA32Z
zn0kl9N78O7hrH7S6FarDVKUkcwMeX+fueXF0H8slN51EjLKBoKz04oUzGmKiixfDYx9nnSq7U25
bUB8Yw5yWnBkTzRTv/4HvgJtV91WC5hnkxr9R0gGnc6c0/5bZSobR39ROLjhl96KNEnHlymsCmWZ
dS/tuh1a40fJs6hRZjUBerbMzjiNP4K5ux05PFG3YQ6O5+VRuIGe/FjLS+fTBLMCP43RWqL8Nyyn
aJS/tDKtj4qrp7vovO/AHZFhHD8/zYly5OcQnb/gRPTKcsKRR9HUGkTKWlY3ikGMSuS8kaNw8iTD
IxfreQi/zDCzDlfpF/vzMcs4URpjnOSq0A56zjJDGuWc+HE7x+qLpn6mQvcnclu6vh/Xcke5OL21
3i6aA8MV8vhAf6+6d6F8F6bTVaIOz11mGKw3HJg3jhER3E2NpWA//yt9t7TVty7L6WJmAEmHZvrC
IMRkh3exjXMczCezcNa2BxmDByt7BKphSRYH/gldMyLNHMUocdwZdwf5v9MI+JM1Bm5fU1ASexrD
xTErYzU0ZJg2fGgp4KME0cpME163GGlxO9kzN1U0TjWyZs4AxE1p85nAmJ9zHJHkFqC/E1sfmF/R
t1Ic/UwoqdIcXmbCgg7ZOVjqjAovJuVszKBL/wVz0tVBTeG/pP2GPHucrB1dtj8JBsyMU4tQDLVk
tvbTZ0pNzhmiQvCO3Ize2LU+yxEQ+twqIadJW7sOTgAnqTuMG8jcH3ow2K8T+Mgh5PQ1R8wcuCqN
Ro+2QSgR4Dy5Cz4wZDfFOmzLdvFHHiQRsRpd2Tq4pTrNRxADAN8teyr/+gP+aNgXd4muu5tzouAx
Gtbj7w+N+WUu4wJHWXn5mu/GvONG2uf0TvXc+5BQBxTAJLUgDGpPzWI6RJR11hkYPrOWrA19DcUp
azf5klhY3wN5EO7jGKJC3IrsyGE8Bm2XWy3NsYmY3QfdW8FwvWeVila00TYBUy22svE22XfVm89p
YyDYYCH5VhtjaT5JVUkvRZjmcwmy3w51jug8w1PmlV6UIMepicQb+JLNIBqLUscQcloryMOm/Uj+
vgQTMzNlHN76AzFdbx4dr+KPZ5xQL2RQc4QxxiuMz2BondEa1Xtmmz0fpz23qYRdl/oX1IIzVEGE
tS2/ywtl6zqvhZe0UyOejmsLURBUA0JSKOeTuXHCMb6DovjONrD0gAvnH6Yt8u3TrR6rVjH1DIFc
COBnLVTvaLVJGZbUPUVgqxB/YqGUNgG5zLHqwji1mAln1WcHip+keqodRBNmeTgPIcwThf6DIbEg
cjrcxUiYjZ873zgA1pxzSBXRwPGJdliy97ZJjxpSTWJf9CGBW4RPxTluD0d/kFsxU0aLe2fAL8h0
K3NGYw/s52Ug8AYgRB9rxOuWQJEo+gq7UDEk1VTpe0ZgOV/XjNrvlaMfVr04evZIcvW1QwYbnwKk
VrK9sheEjyhfBSmV9bEMnHvgxqkjnt3Xj75xuJCl+DIaQ2V/d7nAWDP4XfrVqSqWjJBm/ZpJrVJ9
4OKgKrutfEPNHFTdFmY3bMP5pYyajxqOtqR6o+KhD+jV1trdyz3TmN6WqXNYIgRrX698jDw4Vsw3
PTugotZxGCL3hvbs4GaQWut4l0XobL2yEStyRRSnkrSvZOgt1X95eWTP2ySVwpjyJmFYg93a+4ZI
1oafInLeKVX+1s5TnGw6T161tXzFJ3Qdp8+mlRPXtygskFisDrRkyc/sC15jcynj9rzarBWsFQxy
k9WXJgZZ4pvN6QRuq/un7UmRRN08OpQi0nmZf78sGmd+vjowwVjU1j80YXbIIz5FtConaMspqFF+
igZeZwWg9x8l2I3eoPab5gpt/53O54gpfyv9ibdlz+gsKT0+GI3RDeF1xjpKzYlqVD+KeNFSrtq9
6SLOtgN3pu6g02KmG8tag63t/ypUg0xfcAgoWJIuJpD9DqwW+KwZRTnv+YVvM48gfqriUupbT4jq
sxWSxIKWQWOLON5/KL81vvkr+j97hDI+QX62mQ1afyLNImqnGY/cqPSoReHz8GTa1ia9u5MLoSRT
t8Ui+wlr8OV4c6ouovCX29JXFK3aBTzxjhug59MLytkTWGJ09fX/dyrxeaFCfJPkC3woLOwjs7UT
ATE8kJu8Enx8b9AktaY9pSLjFcK3eK3Htbz8GLampcB28vs7+hc06Bw2ZpxCrtns/UlByLdRjiwu
mCCYmTpWXPz+gzu+4XQk+fmv6DVveoCcK8JVY3qP76upQGghSJTqGYcKVof7hUmDB1DQ/Q03dCpp
whME4wjJ+meInA4/qiQus3UfTeBdzFdqXdVYlC7xhIVx7pWVD62QUObFrVQflFZKVhcREQkdPeLh
Ar/P9Jy1WF9DVkM97kxubrvukF86qUQOzO/I/LiiDRZcQJzysDnIy9tPrA3E5v7dSinQ16mlzCHI
3FQoRfRN9ecbKNcJ04MJ3U27hsuYEE4BHvroJksIg5QBlw/orWTwzGGDbQQL+fxzPiv5hgp9S+LJ
RBWQ8SrErD8wyyE1idwBFLWiLvvmJfhynC9ZZmOIDb1IftSxKQEflNxRMlX5A6+nuh0FAN6A/vKn
femHi1daL8iludioHFtyxQUUrBJDawXuAuxqvZnlj6AfEKW0jrAnDO9VcDRP7uVqADDAkrTZZ6EN
rUITqd3ryBu0qT/0CUolSFEEqpiKFoieHp2R2xV4kA8LruFjSLsFcTGsQLQwLcrmAJHPRaCZl5z1
jlilMqXGjj6UT6ecWH8/v5Mi2y8NTxZPm2LXWZonoCfReILNgxV+rYQ455fIQZGg7W79OzxtqUUA
Kgt5CXjaZUe5RdbYLxJ3F5FSbhwQZ6gfKcNaOlsd85V/q+G2FvbIt6Rq+B4kG5pW5f4B8De7Zsoj
OcU3QxKAibdediRF95l6zV+KEyQ/PSoSZVMNzZP64zH4IDdhWzrY7reapvjTAEyl1ZDn5w8cl9Kx
0Xcy19h07C4ZNiSSqkj0TezTJUNY9IcF5BrbJo8z5/5I6GWoO/Fq9HJOV5bXgNRfMw/z6ZS0+Rfj
CvF0dSrSuTAKD4OWUAjR8gy4qKNOrV5DtmxW8yu2VhM+paWv0NSZ7Mcybq0LPt4Lhy2Q1VS49V5f
Ge8oqIP7iUKxbQBVOyIs2B1n9QQJG+H//Scahn2J8rZAWf+EstRiprCM6qhI5bBfEtmKm8GkGoIC
MnZJYLIkoWE4fbaGqqe+zUXxiqDdL4LNGz4/kbzlwMeVHOC4AhOV8fxZxCp97DSB0O5GHLq4BsQY
W3PHyb2RR2Aarg5oaMrY8zPIgyDRI5oT/2OxUq9zIXCRwPNsd3N4X0IbFKb+ikLmGzwrrp3WGc5G
wSshhZVZYh2enHyCGEqbT1DeRKkIYy9ZkDBpgbs54YerGMcl5c31e2ei0Gzz3hK95EY5tQ9GDqlE
xKpRlSSilwJ7ZfplIHOPMVrtJ/NxJil5x8NCyjyRS/FScIdElBIbLiFtQVsHmWhZ+G6dlBpRRwtV
oubGMMqkdnJCBl//70ncqsHCQVurM4dXpMd2K1ix1KdKUwHqSy2zqJTwqnGOEhOHe8qwL2V29qsG
WbmCbx2vxKlfCLYiAQXP9KCNA6glRXMaaesS7WcekfYa5cBZENSOtbn0WqQGlST+3wX4W5NcmMT0
Cd2aVxc+5MoOseccV7pr3iguXXyuWsR+gycxgr45ctmiufHC6fIu8vuWxl4zmXXjXJcJDF+/KKwo
FdVscD8DCtS0DPYjp+44/qDWmGgWbCBP+kcmSxaTQp2DbvD9OnQTDTSOeiXrf/4sBIPynAXkwTBO
vXjsjauZoA9nh/Cs327xHlSwaCd6CZGWSw5AMv+x8hKc237hnQgj5GewPxLV6Kqru32ZU0Lbu/eU
oG+lTWb7F4r1qJhIwjI2JcIFYO5683ghrytoRXJntLIqvSsfCvKoybQ3aWiAYPsQyYLRZle60uBP
YmhxDHNNpAnth1rrGrot/yp7e48+fwgcgqlHjprOXs0a/cDXApqRD7dDq5rUlPN5Y9284cqFqnUH
A8/zqa4emqTqctPkGN0On4G8Qqm17DyXIb6BRSqERd1idKLnivLWpgG2qb5GEpVnWikFCReudYxC
aNLmb6uF1VDVe5rXJyvmToZs73zMoTEUx9Prt1QMLECRKxjhNQlLAjtcmTToUh5a8Z6Uv7kSvOQW
fK4RiSTz7EHydb5F81WrRNRMZE1KRDQSczAzpIysUejWXwTA/xMQQaqBPWeYJzleNtVIaCspooAG
fmY7wGOugtbtOolSU4T7qTVuII7tdKu4aMSj8MUW0A8Ll8E9jR3ZulgZ9eQFg9r8OiRBpZOZ9dxR
aUFGJG2q6uetIUqTB2RgGOQ0+sij8KTlzRYbnoViEEmOvL1VOKtBB8fe6OiwjDq4KZ9Nk5gBVbxJ
JCrYStfjn58+6OggWSPiOczS+PxOFMvLlhULn/fdQXsS2xTUGnjdGFGzETxQqSma+vIRhVnAgb6m
nX2ljbvPuxIbs1aA5bEMGaXhDQ7/JjJpe0dFdTxpUKvfYjvVf2dg3CYjcjTBygm2HIAOJI5K9+GY
JRKnZFtCQYFfO3j5Aelpqq7laCT6j3/c28yksMKimdgxBZ6h9LnsjCXCL3NVJWhvZotbjiJIMxVC
DLB/nVar4WmNxbVZpjhWwDHZDMGoN47sSEKE9nuyFFLam4Q++sWhe+yfjyBTjfaioPNnaVJqj7pd
nKmj5ZLAvoSChxuuozOXKqAIpkOaiUFL+iInWgK2iCmRc5HWas1q5Cy1JKaTpd6iLsgkO/oCgNep
PIHsz5Fat+CaGcKcCZfCDtjlM2/HwBOMGnn0AnvzJEFAJpbLG9ec9MGmYohTPLx5VFQrexCibzq/
3IPPYcTNywDcI5jKtkfKW7/qo9XHGNaPuKHGvotS7cnOF/jjhlFygIBbjrUxNFqTKQelgJeNF7zW
wLyZZiFemNPusaHkFaWflT4QMBjeJl3MRPuHea2fLEMvA92fF7tud4QA3IrObDjvFDaFyH8KzjwI
o/iR7uXWpQGoiAhOQhuVRuZDBPIDxGZ9f4Viy7AuBv/m14FER65fOBtdSfhFFuvSHrf5ciC4F1Jd
gHSp09hdMIFovhtsKu4+95zR0SLJfb9Gww2qhfzYU81CUlYT1kNsXisUEnWy2JVOyUe911HuB9YH
mcE/hbbecKXyLiOHAXpS9c4UTqX2dyTQQakUEwP9oZTJCrdpshfjyZNDp108t9bp4vqF4STDznuK
0eykR83ezHdsnMpdEDUc8vI8li2h73MwKwo3Z5UnoWVNep7wSed49tIdmbOVBFhejp0hElqsop9g
r/sDhS8r2P62gVKh9ma1yzz7gXIX8HOvLH+Wpf7+8VH15FtEjZxq8aJMkWlp/dIKcXWyYXqzRtOT
MgXqBAa4s6VMpF7I3KgGOaZiCAKZX8hVpTJ3D3JbG8BBRcv3Aqwo21npvrNxfdXaNoYNTcZt8Xbt
txargAtQvS/zfROUQ5WZOLOh76gk0AinkINSXxHWY5XiyW7diS83oSLQCYlb96KYKpnZ3Ls1Evfx
E/2pN8KCbtG13xUbHcw6DNf7uGAtgiIZpggDaQY/5ri9MH9dmS1OVTnBFflac2AZRGsBKioVYzs6
ZEEm9jW3Bfox7lhKKMh6jU9O+ORIGgn+g826YXLHYN1ErcUdasldDQ69JB6KQVkNi+oxHe0wYpd4
fustdVpzKhwsvGCHcrz8Vr3kIMJ5Uh3hIGtCISCsnG7iK+wdPhNmHeAeMkMTcmbyaB+TZr13DJwL
6O0HI6xhh6FiG+WxHfr8vODPdmzBX2s9b9eR2KjLsHqb9G0XgBRF0pPkKdDCskr3W0HAK59L1YJp
n99uFEbXKM4XiODPljhp8t88ubNA9GBifcmvDn9OZcoi5SLJOVHcSD1hAbjfAzMChtVXJ0CSfVwr
JjCC+7bE4l4IUEY/DDjp5/WgBPhwL+liSQUBLl8janSaVKMn+DWPfabVGP5fXSKC88bGAhjvwRuH
vDd7VbaO7BT3mgBqT8+Cq/6c+0yVP0i7fYl8csaxzN5EqDAEWnJYp107+8EJsk3yuWPFpT0LfFWD
u4Mx7ng99w0+O39a6gJW+jGaykPXFz7HdI+ezc4je/SnM5Sf2u78OheQOzDPERKeVkXTAQpPvBhv
I6AbVD7rxEdEoXMZwsNYWGBnTO5BQquBlkTO5eJzwKjY4u9hJR4VzVQHqe7YsTT12C9BpO3RBfDL
c6gzhOUDimQKklnkdzU1uUZZnVcC8CNUVfUvnSa/7efMuMCh8xRbDJjremJn8GQXh/yadmoX6CJs
jiD0+dGNUAt7Hv/5yVasf4ZUysCxRQvB2NxzbG6oqKhxM7QgnGxY1D8oQYtQ9WeR2S8VYxO9PBjz
BYh4XYJUsEHVwnJLWYMoncRSkOzP2F5pIOYCsk6vDIjQmywQRcDJYxo+q4wn7N9J6Om2WQD84GKz
qHHNYdtZcVvgsTglKnidmPqzvrJSG610Ayh552Hk66W2KEidEOIgUOPy9weJFaVWxy52Vjr0aTQo
nOZtzNaBl2i9nKgKZYuMy8Rcii+ZCSlAQozMX8HRzJjxCTyK53S0aor5Yg2v+Vaoms9IfWdmUXnC
350oJJ0HYqaZtF5r0sNNBNKTQC9giKQ4YByFncgp20KQ0drOd7apfLlAYRSzNYQaxEehXpuMhJ3K
amgjIpvZQggPrP+odNTl06vnuw72aK0vd1JYBFNRGdCR40ChPp7EBtjso/3hHhvMpFENOMfmqQG7
62ZAGbVIP2QXaAw2Y3O4pvcKBL6wWI0s3DBtYZ1Ah5OziY+9Ap3VIpWOk7sYCqzQfMzZZFYz0fcl
JbRq0P7TmPm8fcIka6gdG4E+D6S5xQEF66l2mdcktr+nKNtuZfKSOs7wiM7xY7cJAHvEo+7wQqRw
ZgBQ4KRLYBUkFzHc5Ref031sKS/BAuVgfVaZS2VpX+OWiqk1DSGafbVj65P4+8dvvTfxrR3nIL/o
u0NI0V68+urEYgb4kvcqBXUMFJYhwHo3VFK9dXr5PgaWirdofSjxNi+Vf7dPfb92jvHR4Gl0XQSB
3EoTWCrY26aM6nmrnMGswKOkdWqny73NEEfxE3LCoLNPTd+m0fnUYOVSKyBMwvWCJvbBwFEUS2V8
5IT9xW3QYe95nqLkqmYNL6SjTBlvRPp5S5045eX1nCR+pxTHHJK7kwzo5uT77nY8/5YwIyfVnlAy
Ahx20IxBph7Eb2D0StY2v5PhfDZwiSVzQhnwkjB5H4jSCjf5JfYQcZzYwanPk6tIR+v6Xw4BthNI
yLf18nk08SM11Qfs2AUivIBkS1yBz4gddeik4mGTl0Vt6MWLYVVQuqWTQquRlL78YuVsThIKfc88
sDDlBgje376GGUcY+t3rcgS5T5nNe1QViXQzNLL9+1H9ZMzdtyKpKwxfacVpnOlfauRubiHSTbXy
SUbl40OXOlrIBw+iwhqq/AGCXAR2ZxNug19V03SQhKik1d7dvsO/cviNYT0w88jmKrL4KdeKJzZg
rmdcpJRoxgMPhCuRFbSXPTHi0FCuv7PD7tpqGHxSyhXiU0RwJVH0CmzIHEO23HAriL7AOKEMCQ+j
FXmBEjlw6Y6/BKtkjLXUYYFGd2EyYgIRffq3MwzXMZ+Yvvt3j4xpK1axM+qEYwWTTxp7TKGDZ7k0
+JHyT3k4Wz5NSRe1tNUkM8Cz2a/iu6dm8QzhbGe4Oo4pZNUJdIxC0pLvOfe65GvEhmrbJ7JMtTxN
W421mGjqLfdbJCVfcufKD2WVSL4JG4vNmgZadgl39TLT4Aoz0P+K40iUmFbSoIHLaKXPjTI2AwKq
R3G60yvPmb4dYHLouOz8qCKHPfbZd3oDE/ttTbuoYfSVml4UbkE5vddKHqWr0p6e97/wp2+CZFuw
vjK1UOzO5XPb1ydmv8YnySbdSBbmTxe8U/K86QnCRmXDqvnearLDHAE3vzGEqYNhXvQKe01LyYCC
g9PIZ1bK2yTpwBMAK/eYgc3c/HyNXJRyaxfj/vvqiOElxJYa3cublJAURbLd1U9MJx42zLNNAo0o
8Yjl9QPkRBaEk0rqksVtt9pMcMasKv8/z3kveSFSzi0NY7f/TB1ax6hB6Cfw70vzhmk2rAiQVUq+
P3MQypBW2YwOYeDZwnsksKHH6O4HitKMZ76VRvjizTlQKBA5JmwNrS1bVA2Z0fRzByVVfG6FIzRA
XB7oRVJH9YwBM37NXHnrUfb5ESFuBSQYUeD7dUH8WnM175s7aje+va1LQ1cVZaVEieabKeBkZE/T
Ije3hgxcfYuf4j6zoe0UQ8tafoN+YIr2sXEaJXaUKvmqViy0f+9vI3K6hGk6eSeTbXTMy3AEQstP
qZmDHOGZRSMcVgDdwAxDPh9bAB/O4Nc3DV6RYHYw6/pE49Oczced9g0SHYSJ+MBiFMMuXNwafaGY
wBcV87YeqO0ZtXn2Sl/59+jaC7faECShtg0xGqDzxMuUmj+HM7L0vr1I4x8tIzLJ1g6IahhPNqzJ
HppROsf9U0RaB0w/Gh1avJJyc8rr5qdf+wW6adVRoyW0oqxEsBdJS218rmmYEtr2XxkZUaD9RIZA
Uf4UlC5ndX0t4bni5vXfW2n4VJSeCtKLjPcrKcMjJVT19BPHvIlrJsLFXJBZiWL/6UEnSq5ftBbR
rbcD5FFu1GbteYdZbZKmWJlFUE13wZ1yfqoWYxalHuUYX6xgL1sYzCUP1sN1p/rlWW0cONrGjcyG
uUgmdF3mFD/tZCwRbyj84Hc3AhSvIkjBhTM4RXBJsdY8rW+gLR2hNvN0WchA3aA9bmePcEgIlejY
kTj3RUSAjUKs2BGAT+gwnD3TBcHgtJjhkVbNfFj49LXjuWuT2uqHoO2/5HNiSumxdUEgdLnUhRk6
cgOHGPyxduhTZC/pv8WdF+bqlvfkrUUbYAKPGnWb64VDdUXwXeE5kZ+y3cuVRgPq6ZVgAOZUYhRa
e941sJFmXx9fFZLPtHH4mhvux3ZrgcrtdnAwpPSmlWvZTtsN0z/37AHnAwNPEmQV69J3mmvExYBZ
7xvyoO3UejNgSoVhNm7gkWLxqqWZZvNBxefUDlWlmjGme8bsZBjryGaA7w44AL72EFYjXJrWPWcq
af5qdtIahaQBd17S0CBWOmkYzb3sfvKCAJitA455QDy4ocGYSDE9gLAyGok+yJhChZ/nKeAxPrBT
vAKtZjN8zgSOscLMKaLpDkbX+IE7thS3KAIWLdXLnPiLFK5JAkIchsl9hwNKex2Y4orviwdqOXf7
q1gtIOS2reAAtSH/ZSdYOKAcN9soPm/SNYGN1Pv4A+esnQ0NVxWCiwPdqJEuSBIc7K7LyZZrS5om
x18wjYWuvms67ErXeeXQLD9xBzn42/Rw7iUVBwanIsdfaiHvp9APA8jxaqgwuGNMmyFx6vS9oVUd
OYRyHCKGqhkc+iXe2CYQPqZ5Elb466tNTU7RMVPjlEL//nQo4VvJEsD1QlQaCyvsYURzfwYYVy6U
fMPSuiQ3DxF10FEg7pZeYqwZ6QQaU1tTkW/kETuSg0LnWNsIc/uxfRWXxaC//Ip7cpLkPP2snzks
WoJ1z8d1vJJpJtgNmVCYoWPPOSS7BTmPGOcrfm+aYOtQ3M9hzZmnZWyxmrHA31OpHXk6S5qSlaGN
Gc3/pJjKXzISPdLqIHMua1jz8w0lRLvOwkNS3EdVYkTv0sM6kN/C3hOkjuGK5F/6C0TKhag2wO6k
jNqCcVIS28fatoGTzvpsC9+tzfwWVr8j3WvR75Lxc4wHAzsSgmgB6uepU+n0hCdWwryDep7RylT3
c4mFBGri1bMYBe44f9hDhNwJEOzogcZrBB8fHVElhNsTIgzZndjvFEbRC4c18uXExe1gPQZ2AU9X
jDHBgbC6vYmV6CSSZu4nBCe6tgctWA4KdCeqD2YCQ1ilwnym8bXTToWLPjGV7wySoKnDOzF4Uf68
Rl1uCi6Qy61b+NlJnkk0zJdkQ/MuV9rdjj0Wvmm06okTwGBGnGAaW+Dg6ajIWvIGljTC6i0LFRDS
IE0HXzoDyHiH4LRBeH2wvYVXzhcuC1TqCRpFmE83O8eqGt3i+CzhqO2HBclGmIGJbKTZOEjqPdHf
u5UjS9KRtiPm315ySUc9iU7yOIZ7S6ali6x/z7Ea2BHT5XMq3O8vAKiyysLFOXXkIRbUNjIX5yyk
p8Qb7oHYwHzAK2fn8rC/p0L2whnvukRryUIaHgqNai2mrkbyxBO2BDXJy/3NTikX1WXDJJcMsiix
F33xTHgYHwdgmc4k91CqtJokGvAOJQ4qjdmBexlMDYToWDi9kf81cRoraXKolCNaveGMKHQYa019
n/qWm5neP1Bt3g/a3iL8Qk4zrgfHW++9+MDH0krAL9olO7mTN63hi40OYdJ2Peo/DCISXVE97DuQ
XRGIf+cMPFCYIA44UoqfMThRpxyjaYbiltk7IyqUTWssnfz+oxKw8t298BwvoyhxCe+iWR2iHrw7
n6NIrRaAxje50etlC784G6pLrDjGygg8pBs15M7yRgGYPv3Ue8KX9EzCTCIarin5gl6fIKMQeTiU
nA9nPZMz0dySZa5qrLTnz2wNae2r59oXDgYL0cscAKTAvXdV14PvbdV34ERsoxTB0UR2ygB18c4k
RDDr0C+kQ4iOQCRQc7H60EDZ3ZqjeYx1YSadQKZqD4fcsJ+72SrFs4Fad0i/j/JurC6Q9Gx0sLzR
N1/usuljtKLX8Ssm2EPPPTNuffkUARgz2mLiblIcrwI6anvRHS5xKEtS4DSXoADV6odZ6DlfP9QK
jnu+55LDsL1WS10nW+o240Ytx1cqVAphfGJb3sVWig/yToLJBto6UPkAR6TDHNupdsQytJ4etTfX
gR2R35SwbAnkmnwnCY/ShPqpDZoA5A13AHBESVUSm5AdC0SdchVfcmUk0QmMArnRaQgL7HaV8IPN
oDJzBKkQohJsNJ2qgYI81fbYas2RFXK4BcQXsVuCf5GTz9XilVEacCUI9lIPK31p4vCGplEFf6og
Jna4jKIWm1EgaKbDaJkc+kqKf7WOvP3DfXOHW9F6O1pp8Uy58ptESSLn361sbptuqDFDwjr4M9ol
QwOjU7s1ncuz2u7bIojS1KQRfgVIHmFpWdwGcCImEF6zi74D6D9mHdb6awYCqY6+D8qsBmTSq1ZZ
XDwBY8O4LXQOrF6gndd32mh6Kpfpjds6NyBx9sjA7FXOu7brnfqJOR/o8zmoLvjqp22hJTGrNZOS
4t5PtQm4UD//L0ariVKHroBh5bdkq9Fqd7dIwaTl7QMjsd8YI5373A1n17I0l/dbfVvlgkZxS9+K
KhlRLByDUI2nwAHPVZGJjp9IITz5COMFqP9VhDFRYc9gW4XEdfbWaLL1UfMKl/VuuQGtiio+j2I7
Jvm/Nkx/KF97nkex/0MNiQAQfcEq51oPYYJTxOW9ddLNODtH+1zc2WC6zsJ9W2O2A2Vrv4w065U7
gfib17bIDg8kPtj9eeQnNcbFBnhjqihB7l78E9KL3Plc/Gyj9IrFOF8mDUx/gEHqjL31Ydwxbxnp
u9MoxmCG0FFQmPkyqBouyvmcGYtDcEpZa6BVLYsNU264BZ2B+z4hztctQQQwyyUZWZ6d2u7PUMTj
H/lpOT2S0fBWSBKLsTgpEU+U6FO4o1wJKXNKzmFaDZKbRaQn651oja7kWHSsQmHP+mNnv48bSLCH
ZaED7BF/vS41btuMNH1pyX0JnUtJkun2QYogmfEfUR0a+BFhWoOYU9o0w+zw+xfVQ8RCt7EeC16w
McLFCPt0TYCyc6FuCLhmDLy4ogh70LKl8rWwQpe/yv//PGVYSCY52/ooyltW/2J96r4nJJ4BQHYz
HaH0hYHX2/KPqm8ypxmq14lqL9SWW0j3ndsciyM+jHBr4OZjVVL8fodgck47ZcJTxDpKo+KHlcnv
K395Yk+LmEY05Cfw51Bn7nZoZevrlUDA1MCZvlRJTywUur1N2EBboPr5waYx7j5hVt2cPyOcaJ21
AWzwMYvyXxMefKs3X2SGLQuN79G/M2vQUJuoNZRLg0HU2pEsSJA+2yLFjf3NysRl8zwmcc3tsPfH
uJm8lc6/o8At3in0v3YlCoJFV3XGD/tM5QGPSixbwG1nyBtFDYAALmPoyfoOtgrv92IUncCJ0ktc
1h3F1xo+6MFcTRs6L7UzuEnwumziO2Xdym9K0ZnN9oh1wDUxUtMI6DU5JXNTFkkiCQ4rCdyTgnUX
Dp6qXGbWzqRR/4H3rNA7fpn/LUi1a12svC2ZmAxKzax5wvEoOhctWQ9/y4r13ICpDk7NzikrvEb2
XlUwdACLc/eWqH7KDqugZHWoRQ3Ye89sfAgSYfFAxxT8I3BAcDhCQVNdUfd5aMxDVNWm164HpdLd
Z3YuvYJyBR+kynf/7DD0t/WzXlEbqGB4I2XWMrlSwx7NCpPigiuwm6Bjq3zfcOVCUNAU0RpHN5+b
K7cjdchXgwGPAXfLrGy/pV41X607vpz4zpTLBneze774oXjPP4qtykiNRXWUVeOTDNMe//qUb7oJ
S/s7bXmBUsv8rqSNL8CQV4ovBvGsL+/57BuGXeOWBa3PrRsh08EEpX/4MWieIcm7dTwcFLI1aTW6
TSHBfxzVKEBJRiYPGkI+WMCGo3dfk1AcV+HejNfKeSoRO4hmCf7vtoUn+jXFflBo80QKpHVZwN07
jyQIhLp3NdaWN4R/3O7MT/ZoZ44fU5Qg4hqjQhGtJ2AhPjmVGtKNtBJVoDhygRuzpDiy+lGG5Jfy
0N0bsBfqFAOMz5jP9S0zkiL3NfEtbrV96E+fJfvP11MWBDyTo3Dy1/jzlnuWD1xR/+Zqr9m0nC7K
qGketWvoqfRItTTLkuAb83irgZu9zxi6rXnSUs5xEzE9up5uLc353LGjuIYdKdsrZddCfAKBaqMF
EXGIu6R4Qwv5XjR7Al4hmXd35hpwP6x8lJE81S/DV1IxWFTOzvMaagSUPBWZcmu+hpSdoqWAINTQ
qCERKgiIKqN03cRsrP4d+toHaq5ek0PKJpExLZpKXNbw9k956kJRN2VFI2jppq/kmpvuWekVZNEd
WkC4/mYT9G2r3yfzbUv2x9U4Wd0ch3wxtmHBWjxt7bJb0hN4xh/XeJPUl3xQBv9aA3hKYYNEl/bj
p9HHX8FZ7hC+VD0VjqdPOODzPJ5AEH3sRQf2E4W/lzS4CR7u86vnCFBQ0sxhhu9GfI1NsbcF0w2v
msH0rftlO2Lypd/vHtV321rwwa5hakKW1G/hnYT8Mhk/fzFBODBk9Pu3pHiElzr8UeibdAnIzZFO
gjiC3vdHlgl9on2jfvOb/LwmSN4dCe35khy7gHWE3oBFcKRVbAZUgNIeubESAMJXZUcmxLl+n1F0
v8sIOSDMiwepU66k6OfPvsGuaRmMZRrb1ey1mRx9yGdL7iN79cel4TBmmZcFOKNq+Zxb2YsylI65
h0M7m2U6wZuNfd0kjghLO06TgQiJvMTG1NtVVHKS6+Tnq3Ud/tYkKNKatlQ0HN0zbpPbGQTgqNgm
6/wawJx6HEBCdoRYwrTxPLfdwUq4RLJ4GO1VN1BnW6HOe+/JEFlBukQ9jFOw4/d/yla7XmSrxGfx
sjBY0UDVSaPZ/e+tWn7jK2BU77jX3EsSEOJDfU+6CbzihrpMLFjQAZuDHbamIeDy6X8O4P3e++yq
+mfI9L0Eu5soaF9zLKfXcnC7NxDg3vFxvTo/AFuLUKS9+oUEvkPQ35osyzHwFeSLR3hl98J5z7lu
dDCy9IqIDvUxudf2kvgPrDJkyxyZgpue11bJk6aDz9GBUgKidsrf3q/FQlpqULhb4xzs9atTSMra
8mZ70JZDOran/5RfM3OyuvkHUlx21ssP+rYWsIHtaeCRs35HHmZwhStPZDMken7TTtI4rkji7gVY
zhAksu1QpaFrKimE9HCBwos/c1a19iQhYxZhREeEUdMy0uCAhjWSGbUewJ6TVX5eRaAoGWMsya86
9vInQeXo6XsQTNgc0verWBGMN2ASpZuM4rb88eRkw8tCg+J2Lxy6cbK8RYs5ZxuU/WVi7J7hTJVi
lKpgDDCTJRhvUKV49YPLUj6c30l7mPzZomqsuQufoeLFtL35EixXjZ/EHdSCddr54ndm6MYi8LXs
W4OnQLK4jE3F8cyLVmj+h1lVOQvLesKFfXebBH1RDLKb0ovvGzfNv+9EvpL2Fd/qzsx0k0I76WiI
9iOG7+zEzX7rACbo5YiZrhuq9fKat4WLBc8st2CkCtYl86UhuMfXATRY0f1GS2hpaJ9sNu1P9XYZ
421InFTM+w+8+TUaZ/PBwa4/Yi/BnYWXvOSndj4rBQz5C4vgtWWULrVN8pVWLL0t7aULuTePfRfJ
x/rVIixSx0pktiV4zVayfbDflUaMBBmax3joWvuE00JFXs6yZLnM5VBXhXe5ZCCo7cvo7OJse1I4
1uC1vXmsK5Tc5m8lkteZNpxsz/crVM/KqIsbm+SPWl+QmiomXt4gDrIzKjtxzMXMzkOYAhYYnxfa
/bxWEBMKJSTwuWmbFDl+YoMQS3hWjjBczAtk2qOxIUfB/6jXr3JNqaxhIDYo4AX4v1rob0SjtbCQ
rUPsNC7khscF/dzcWB7QRprOUaOroPd6aTeNrt+MnW/QqEkYBNqTgkWLU+jqvySSyIWoEh0mlp8m
03y83oUDZMRZxDRTADH0LA+3r7SE0Q1LkO4zTWbeT3d4gULd76prDpTXPur54yQTalu2xNr1hzUB
8TQUyQPOYEAyRa7A0fwMILclFYHytN2SR/2rnNW1AS/Cp08h8pDuHR8ivp4oVbFBKYR6v4dX4u6P
UPrbDcJ5oPePCfaL0sl2PF6l1tgC2qPuIPZvaoF09KXMq/gBVXlTilSOOtsrNrCk0RVqEG6nyO1u
ddViPiaPEdoo/pzsJvxTwT3zI6clG2BlS6BGBzChtpN12Jr5UPrXDhr7Y3ZWoXVnPqh2xhvN7T1v
Q+XsugGXPIlH2wzhrS3K/oRaSppfSDXUFW7/oBZAMHtPZI+VZCzx9Z5Mn0Gi03d61d7Q8hjiEuxS
hat3lLR0lzCUsUoO5hBqj2Awq/qPkiTfSq0WkAWjUJVUT5Ido4mlUJSChmCX/kAYkz9VwXzwDi9S
QDzQkK+mKRg3TpGWOu1ZvsGYjBRuA2OdhJilkb/sEh+Q8K39VpkRDJAplsqFIxc+VNrkcctSfZGn
n6tFQIX1SfUXJbPuBpzlKR4gqhu9IbW6ThTPW0RS2izFuiAFZyFPrhAjvjLNzLzn41wONWs2H6BE
4MkMhR+7MZl6hEycoNx9cXtj41ZZPB/hMTc11nFryvQMIobZZ2icNES+BBY2ZnC+KP2IdLjIRAfn
q4Q4BreMryq7n4eU5orj+icoetdaQNgxV4scjSczAzJKJMBSGziXrJO1XbeOjsi7nH3Tao+fuNl7
b84ZCUsvoxQyIXyHBOAVYUWRSEQ7SzqPjxyUhpTWi0lOCU/4c83rtgK6M/UYtlCe1cNEKAsQTY68
MlDpHtppaKLDV2KuvCqq3JqCfgyIfo1B4iVyxJQXEDSKqBzYFGJU+TkuHFhieNb9c6XUJaRoklC2
k+33L4P81KrM29gqOevxI4+sHCu1OlRtcBnXQLUpEgCfVzJ1w5njwEFXBm93oQuvrqseLeOwnuw0
kJxziCwhl2G5cnx9zad2KPFcy9rxwKLik8/b7TiFQhIVCYw7wgK4aR9HYCBcIvOftipr/oBfp7pr
BMealuDtV1AebWZKAZ1JzTSsjU3/QcwezhZwekpaL+03G+eDfaaEYBOxYJE94ZEIErFb07eP8bkC
cCM1ozNZaeyiEqt2wv0KC5sLKWEgLRHWaSYIPh73yVVQLVYrD1Rgi3lJR9Au2QSyFeiWE9x6pSRj
nARW+TlJVTBARKvx5jBQ6KOIpAZ1xeht3qQOWUxT2TmEKHRQ6yxb27bfbHxXzpNLfk3eBIyJ8JUY
dsfcqAWVW9wFkwVP3P9AdufoMiWnEzmvZdh2Fulla0a/F2guzyWCpMSvjEEZdGaJwVLQk6epVJHn
dzNqkalB/098RL6LpDSztQUCPCuCcCTOyRCSMj4u+fCZ+Y0WtproglWb6nEMjhtQzmCt3bloHjB1
xwJHhVk5gyCn79+Iwrx05g6GoqmaPH7ll0lUQkEsPyEyRIXrLt32NSfO3JYBjABIleiXKBDi8a/f
dp+urPSJKSpnxvQF8S/GihI6Ygf5MIGt/MSo3n8G6jSp9bzio+8Glftt80UNgjBeanlBfRKPwRyw
lV4WIJVHRGjafIYEjI+rv58OsTAeRvYUJax4DIGfaKtRTuQEGffBr60xn6iyyz3mhyuPhE2Xs4Sr
xTCXl8N7Qq9TLIyFjXBt4CBLbz3vV+DZjfQQ0QiBiRucR19fvPiBd6d4ak+z4jzaL76VBoNfdC9o
W1S2Lzy3CIr62+ZksS/g0lDmmCM4rqvhp1pMbvMWY63Gim/SuvTQlKl33s2YNLZGT4rPrVWgQmSh
LCFKP7QmAxNrofYsql3ibTVBTMTGRfpoHwZvJhGHzDTU41XloideX8/jY3fh3hPbctGZJTgGbhze
kj5OAk3wbkd9lgyIKJrMOc0C2ncJyfPCp+LuMAx30PYAYYlNqvMS9eCIjcMJCsBVUFA3YABaRrQ+
CWvz5o0YSg2blRTAvPiGFeHJqgfmOHkEfZkEY7nv2TN1oir6yIIzXMIjK4ft3q16MEytlJ61qLUC
JnxFR5UQ6iP/co7SV0XjDbV0WpRkgjAsmL3ChXjbxMwbNpJOLSa0wKw6ce/BsWqUyEH4Au22Kp4T
/jK+8ILFT49p83e5cq/EcZoOovq00CgifNPZsH2EGsmu53Nfo/VK4D08+blU2idNknaEwRxN/CW4
OdEZlTsBq2pCHkbf2GPG2wTxCTvDAujCpaxveDQtv/CW6miPsO+IKifnN1o/oEuXi4lKspy90YXS
SREUm9GjL5o64ieeKQI9rJ9+DPr3DZf73rSWUdEgxqh/gogtZVzb0kPZ9tjsMPrSRXzePp9wCr2h
mCJBVsMsqedXiS035CZs7DX/0fivg1RZzjRGwdyLdMQA6vifupUVuJJa+siagd3guhorobX+wj8Y
237ondH1HjH61AmTPksA6R9QiX5/DM0ZZemdxgFD8//kiAoRoiydVFmC9LYaQebNYOtw7uqihxqS
9j0E2QVRNXREf/JCav/3aCpxEfUWScbinJbz+Vnn2Yu0xrAp+eNBBTV5Zm5iGqvhGx15+JVPoV0M
W/GXHVxkWm/Kj1sBuUjG5M7TVab5mLeuQ39vciUJ+cX3YLy/9IuZ8wx5SRxrJnXCych1piQJqLA1
dzDiHZeGfQgqOZcAkqPQFKSStdgD0wRhQKNT0m5UrcC3DkoU6bVf7awHQnLTK791+pGJWmttrIdq
wOV8wLfAkxcspPlrUQEdY98vmPxxr8uW0NfIufKdkHLaH8LerM9/2yNT8Vj9BXHpKwZJnsZIIMjo
LlLfc6Fmq9F6xKPV3Sv0ZFaIoHA67K5Cq7qvXCnxeoZtV8lcfxd7rIYQIM751ZIGa86X3VjvIHfh
Gq0Drvf4qnxtShw9yrge3lMZVgueWJKcN4Rl8/5g8MhaYwW6YzELwE/5SfUaundbJwoNWw0NUHM4
uJW7NmLAiwT1mVz/G3K3mk+5czIKfDe+2H/W6tuVK3SBDbNYzCa3mq3UnpVczfiTpIGkJwhoxjWv
9g9lE3ZFplmzCoY6FLHYXqM5pSHAebdfLzUBBFEmlyx0MgotHR0V1lbc3NnkAr6Ny4uNyiWSDVh4
xWw0nNeunK3lFfVJOXK4Vo9zIzhMPmZkd/dL3bDgTrmdGeaYqsbG6mQqYd4Dn73sfMTrbV9AMDzY
QYCEj0/MBiH4jOafZ02NOuzM9u5uzg93MUr5xPGDflbNyNPIfrRBrNmvornlJsx5urCF8Uq9mO8b
kgCiLpwpYro7COwk8MkONiBMDjlawUug7XxXMoss0JyhBKxK/7K/xHANtW/xOmwRLnYnvOZww3r0
JO6jTHMENmM+WP54F5GxXcC/0nUmXNjA4TFXt0Dt4nAHn5EV+iX/tUkPc5INAZ9PltSesftTyfa7
dINM6IP1VhzQhksTl56tJrZnhHs8+eIIZOpiPprh6q5hW8DxMz0JOkvaUzpDcQ9lg6/0/F98SmsR
8RX6S/D0RB1uJvbuQeEeMsmRuEhDFKDfmOdpR31W2VE2BNiQWAWPqNOsOFs1KxO4qalHeJR0RnzJ
x+L1HT9n7pcmiD/G1K52LG8e3oSaeo4aZjVo8TLZGv20jrhJiF0lfxVb5twhRuGdmfnVw7EG1GtD
c3Kbt4TrBFR2R83EvYrMUrYR7kS8RqH11XV3CBZWJZc/OOMpl5VOT6LX2OUoQkVA1pk6w5AkNW4k
UMNYcvTUnygk2oNcI1mb1/Tc6/M+WWAw43khilgKsCg6MpTg+I70wl8aWRE+FVx0LK5CZ9nM1npP
zPsm6AP9Qo28mIMGyfl3k4KxMnFC9R8Ps+HrtEajRwavqXloYETmYb2KTfGDLRSli+UiqHv/neXX
uZWnG4HG78Rw918H7s/rH7/KL4rgskBTVWFI0l3nMK7iGKK7PR2sLkloRFlMBmvye65eLfuxrjiX
BZ3KS2Dtib6zzeBioqjsLjSXLJHSMLCqBfHiWqjODOZPNqWTtuTtrxWDRQv8E3bC0XcW6JIgPlot
6bMi2euHXrQ9HW/GelKwUNGJQGiGEvT+RLPu9BKQvd/P8lo+5S14IDvXzD5QDhWCYLm24h6+Y0+Z
mwdHd0L4c+JSW1Hef5MbNQ+m/lQqvlipyYeOT7zHODD9HFhTzU59j2lCwlPTB6sUOqNAMdf+OtKb
M2ub0GqZxGcrTOCs4nBjFL+SKMiWw4wxr34Lr9J7gluvczqSSJfeUbZul/s6KXYAdo1EHhJyzFsC
79WFpZjcoW2M/O3JhSCweUvL1KeQIquhpAgUifH37lWXAWyJSR4LtjrusHztsDffZXujV60NerQA
MSG7vD44Jh442Qe0OzeuTwP/wh2CYM4B8UJQhEeV05+ZBxMymuTr88WejVdZPmVB4O9emZd1FWTW
gQFRJbTY/JH0YyVrVOOs7iADyJWASMgdOBjWYKuQloj6d9GxnZ6rRlH2tVDFeM0bRMxKxOaer/rm
yhMVjjvj69XrEJaqk7qgUorGURopFcJ6CNE6pg5OjkOLECocDNYOU1X8Zq0EcF9yl31vY3d/OpOI
NfnXwINloHRKm/ov4OUfm9O8U23GxqVPXaHE5Cl5+69Po9cVPguyX82vEJ+FWm6WtUjgpX27H2Qp
dqC0I77kLjDD3Cn7SjfPJfAtc0GDFMovibLirW2yWQScWbAirFA7lmMmcxsItT/gVuXC8o0Cg4Md
9DS2U6268v2rgNavLFBLbX4NCU/eeIv/ItbxaXyYtxVIUonTTfXYP3ioZq7AK9WaZhFtUoJ+YCi8
8bdbt4N43AHvOEbuU17+zwL+msBlNUiUJVeA30MdNmkifJ9PVuCHsvN8rKlxgCerreerEfAKyftZ
Oq7LvK4TTbFGbvY1r4lwqWGm+3FPwwZhkGTF9UVFeG55yUDjvAXczFCoqWj2GZpxQvxhcIk5SLk3
RU+dlflzecAf5PWqwD+jPaepp9Lz6KxmR8z46QYRihFbT2Au2bfqgVAqwwSIbbF7Kn7FbV3+9E7M
AsnqZPiVPxGCK0FvaVKt+6byc20yAQeXd7ns3h69eR0VmPZ+1OxJpNsO05X5ajg4C1BNNfH+pJIy
IaULyhN1lQg0tUBgGYPuE0hkepQKHoJ/t3H8fzgHxbYO/YHngoyeDiVwIXxnbo87lQMj+nSIutGY
u0NQGh747ujjNQfPlQ1LSbwgO+Nu9PZ84/YJuQ7wWgCtTqM4gE+35DobaCCkXKjWzPU2/E2j3fsa
+IBvhBRS5Be25wMeXL/gx8sHl/kBfO379fV8lmUu/VXBwGxcWPWdru9zHGjDHubfjqBpE264SOA5
wizAB+BwF3YQZBGPUfwlJXnRNIu++ai1K8TJiqe0/Hhc0UY5datsjhZjMBhHOdzBTkjmR/Pt7iiv
LII2OvY0l4S5MEu3TMllU/fVPowg9S627vL8KWICPufWBACisnHrHFNc1hX6YG8w9FfW0C8paMC/
S5Gt1U1yivmfRe3fMrXjAkxBhqS5B2gvjlR8SYrXiG2E8UqpvBjQmeqw5K27S2xFptCF82AoNJIt
cdkVDCd49lVrwN3LyAQlwhEe/PB7S3g3eZsSGY50BumoX7MA/tgfPwPX2UOlKMtQoqlCjrPcZFDt
o5TwWh/ffACM+mdIhNXY1ldESczXvh3tOW2fv2mpKQR4Vj1WJJ7w9peAH9Nr1aXq+3bXlGPeD4fs
mkZMO6ZvZcPl56pcIOy+4s/vF4mOOSg+rFXYz/+OSB6SYkKbESrztch05g534GLvDZbyxaJV0e7A
0AZn6C082V+CelvLymIjth9cMPLTRTOPLa+fxmEzN2XjQxJ4HpLed7q0yQl3LByU/j/RQWVwTCkg
Cymv/nbcTwR0e8vpOTaEEMzFCfLIGT2lvEJgOw6l16ve3inO74W6l37ByyHIS+RoxfO4h97xCIp5
4yPp19/CXmiHA0gHPyU32b4sG7HmSrqEI6sApYgC+j6NxMHx6Qdfk4Z7Bka+5uLnlJWGWxpjB5nb
F7TZn72gwbuR+sKrzP+VaEa1Iyl+C/Y1wi22S8OJ8eapoDVGKgb7oMucO20GbJ+2kkBhYL9LpN4f
qOS0Ta7gn3F9wJBBho/o/SDt9mN85oC7bFfljWiNbIETgS7UxML0DXOIncJWSWGE9b7IQLbQa/o6
ABMfOmLkefl7spX3VQKy6Q0iViFzeJ4RnSm+szdWe5RNjwFa1eVX41N8eJo2X+082f9KRjZuD2K0
NK59ChQ8A3Ww6Cpy4j+6ezHOi8Pk33VKJMHIb7/KPG3Qfgzp2Hpsuhvp9eAEOmgZfluO7XKdSiAl
vWZCSBqkLq+Hp5Qqv/D8BPog0bsHzbI1Xgm6SEWmoNdAZWIuRy4k6AWWtKRmkmrcBuLzZ35YFGeK
2CURjUt1vGn4GN9hC3AMhVI3Yq229MkgaEWwSfjGjykRm8jg/G+fOBiUJpgAxge4BovHRHInzJA+
UXyBMpsbjy80+ucGUGF0SpydGJjSijpTbhgusLJDrDj3JsCQBHgztL5r1ZGYfAg/wUUXVN7NFYJm
A99beK05W7bTfNHPq0DUR6T36eEqPfUfZFXEVmJF8uXk7YTtNOHrblXGhxOsLbpljtkSfSIgBtvv
r4KWfSeVVKLlrEiy45pmpAkcPze/PZ6q4BYMWDM+zmLH1YfRKHKc/R+kPnZA2JMEv14QNhVC2HVe
VeB7fNbQWOCrEKhHfYsHI3AZLn2DelmQfyXBAKAee8jD9OsYU0onDze8Nq0OO69xZKA4mYmj03fD
xzW4SrppK+AaeQPhI9zWn/Cblif54HjPpxqXA0f40WQeNYZ+8fYy5PCFXan+q1Ov39+KkyJv/avy
IOnpc0NKILW7IW1apRqr7A6G5xmWZk5HOXsbpcea4D3MhXOcBOvnkWESJtf0b7sl6Th6x+41i9XK
/znnYIy6y5RJrGpnSvp1D3wAzFKJP9cRj9/+XIAWi2rp6ZCp+pqrMmpoCe9FyxR2IBaQ7w3tOsaY
+/ES7m/oaIyxyPhvo7XSH/1oxK+OQi18JN8DIP3ph8gcFvfwJC+RP2eRraEz08xiPN/3MOHjqsQi
4/Rya/d4+YJIfBsV6zM3RJvpLJOveyXyNb3yCdFRyOcv05FXtX5K3NVsMl6cNF0DWP94GIsAapNq
dVZbvJiNLTiamdmoomEL2yF8lvoGQKiDcNKvN7w6S15tZ7Yk18yLReww3HNoulNz9eY4qQuXmKOn
zTteIHwnaJyJHOKCj21dfrZGBZc6UQIdvAPo1lgdiMCsgtmLCxJUN1goq6jo6FFbKkyupz6w51co
p8+JBQcy/NDT9BbVbGBGtK1kwc6OSqt56tPYwDI5DBNiXeUgY1eRXv6ZpLfFrzMna/2CBiUzuNzv
E33Wp9WVYzJ5rJgJWf9W0pb2QtxcW/ughEYNVX+gklB+rCPll+reSesY/VhyTlsgGfFfgVDPBF1H
zGejstC0Ik5VGi6NT7g4pvAO95XIg1eZDbwygtb2W+WIXOZwrIl3oqgVdkrhVlGyaj0atdWmITlS
MlZlK4zJ9ShFU5Job7WYaq7EDVwIpGD+rOL2qYCAQt1eqqSrQJgBlcwbyFcTKep46UMfXeGJrxCD
EZE4u4OHj6ZWW0dNUCigSEZCuqo0H+UIArm/Bx683+RimLVpEaWwCDyu3nnDN7ZelEnxwODpiPdN
wxuqjFz7f1C/adwWHSBuJe29QIm7udrdODgaykgEbjKID3WOOn8ws+IT9Wg2RAxApNBnzcoJlc9l
gLM32nTRSvIG6H3juLtKMzlqbqVtUJU1jKv3dPoww+hsT7F9rI22XbcxH7eUoRkkUBboA6rnbBEG
L1elcmLw44KaKaKHLwJ9SBqp9WvP89fI0Bk2esRIor1k594spwTF0QFHNbwfwvMTEHcjWxoAqbi7
XrFFyGGGeVmIC3Y3zTwjXhlRiMbq3K15BzlqgdqdExhfE8ZAPaeI83s1oVDZbbI3Tfmhtyl/t6Yr
Lb0AU99k1oaB6du/nlTYPGCyPdAeKuF+x1DrLQNmPMfu3XMr+bkIeEun+CV2LsUtzHEa3wRK1JB+
7SXinQBmgZluM17NwmigVBrV0dtnPSOZ5PIALgKMQE3G1lKAc2EdFlSeLLC8Oc/d7UZPJPUbOzBo
LLD1uWSRAmHOvS6BBWHYaMw3ON2UvQZVukEFnXOLQnK9WfdIgFDCMKTuYz41365OUbW4VLtVkPzv
7h+dJoM7eW7jiPcW7/LzUwGYpA+2+Y+AX+igvDqJ3UNRV+IYWFbizNMcIZ9TbXPwPo8hyHzEH2QW
I6TPWtVZRNoBfQwBFjU6Qp6dgMzUuBNlMNiFXd7GtYM3mY5AcZ0DjoUmIR0fmtO+8oVPmL569Xfc
Df0aNXk1+2ZB1bRM5xBWMNIysHiQy+0LVNhBKltSEIXkfTfladdVHLkt/AlM6ppExWETVhEs0gB3
iNhwt+Tng59cJ/b4NCQZdqA5gTWIfxdug9W/vOFIVQOLK50M9QWUsSMu1XSB6d2/FgygsJGY2pAv
p/BL+SPL4nOSrOmlmCGBx+Aex6PqTtjItX99ByKuf5tjLu98eVaVTRL2iWxLk2M3P7NxaMtyUp/D
x8G8NW7EQC1S8CANKAebDv33d8Dw970BEQnAIE+68CR7fs9k2XQywK/IZS/7956kAakORslBl0Zm
7FhhYBJGgzE4u5HiHTl95fXlrtKFfOIOr1j/y5XFUUwOoxJdHMp5LSXwq9kCIsYwLDskmD6g3hEk
NpPZn9WTpsv1j/KJn+RmTY7EaPolUkQ0bjMI4F9vVtdn52hQP1a0lICUO3oBd4Rast2RwmtiSKyJ
jC5Gdc8+h1mIXTf7ExqnJu7QaDmdXd4zyhP94J9fxxK8YkKfpCtkeGqwebUEl2trLLv19FAehR8t
ci44+ritDi6KTh3sAvfbmJH8Dhkqd+GXIuOSpraT0RSzOIVcVAW5qLFgqDotVYeHYGYWTn3pEaUN
pPz5UU152UjclPSWP+LJzjamVh7UOkARq2ln9h/whDz1rnWK5hCSxo2dcze26URGstjdIB42tmDJ
PfeNaZ4SVQL1F7vRK/PjQHQi9vYSaRRnCBWH//MuuPurUkdxyGxY/FY4M70E3bi9Qp/PWDmVKRvF
wWxCG2lexpv9smQhXwTGtQmZMXuU65oP/h3i2biQHHwJxCh8/kwOxMkuOQKuKYje4EuMc3w8e5fi
WzZFOChrfNQ1qkDTA1yPtRf3lWT+xJ5bTxXcjC4uAP3H1hO/Or4AIBvlu+YHzlRhdlnahf5m4yXu
vMIbTm6yIuqZNE+c8d2okikB0qkfN2PjHWWLEC03UR/LxgNLrCaltm86GNq6DH+8JROZeNjijkCB
WAFX9h0rxH9dZFuPOgWi8ogkCnEBFZrxK8eq8NuCLFJK2kkTy3Pzv7L6+l5qO9N1EEudcvl92rXg
7hfEz1RfFniyTaBnS0pu9LFKF2m/7yZnzpXrX7gnNi9pqa9KyqWA7y0WGhlnGxK79vd4MN2bPozI
HAQBZW8yb98boDMPiH+eaTZ7XwF/jLFxttspOFCz09zs8Sbj8f8aoFOO5+MJtlrASKiEbIagJDUM
yU1Q3D6HpcQAqb8aTIDIsa7PSX4/2HG/tOnX76b8bcIhM0sbwNLgadtnQH5vrPfX6n2aRp5rbBju
ZRFhn1KrBOCchnX4qEHK9xzhOHLxadbHbA0xPyZLA4Q7nNKmM01FykawbGzkDbtjw1ci/PJd/1hC
eJn+8YtvInizrOqkovjaohoc69s5TwiQfj3vWyYxQB0L7VHFPrtn0EbSfBBzroPDwFuBiJ6j/SLM
tSkFdg6QSpzi66hHwHAMEjVNEp6ftUcFJ/cHLquOMY8fNtfQ/cOdCe7jAi2HmK9C++XAs5L7qDmO
I0xmuahC6dF1reUntf1yCOxH1ZNWSdi1VYb878XbFnp5OXDGwRbbGVjsm3FjLuPUjDWqUa9a11yt
n/T+Qwmy6KrRx/tUiapNWLIpIcoY9F5yCuCfv2ZEi3GduIglvV8XagMV1d3TgqG1AGchUhull5DX
lSzzLHv17T8lsehTDHvZnVkFv6tOoE1yOJPin2cNNp7yBceynl/4X8gVrn0vWUoZwJKoY9l4Jw9q
ErLo/n7DIckqdDtMZxL6U1EQdc51+xmGpAEV0yl7eAHoW+EJBmzTge5tJDgD1cUVztyhcvMwRK/3
BSYE0pf5+P494YG00BkYWO8eA/uqS23zHIlGkVxlO8bLaAA1YQml4IEYUEJeMmEIhTWhuCQeMwM9
QJUmYQBmiWZMB/eG3MlhgOKBSYJ/BALfQJBbXOqlJ0rPRDORppVRmamQD1UbacEJRTDwwt90JGi9
DSXTfZ18MZq1mS6Q8GRelT9rYh1WWWSipefIyiVm5qlslPYkAmzx0v5IpzhxjgjZBTrKGPo7pDKY
fMQxRK0MsSagMA6O7VqMOH1HbGM6pANPXbW1IWrytBIVGI5bxampt2+0RW8Vly/w+xGHTCPNAMuV
RRaqgmJFAUGgoNi670QFLbylV2zlgHs9YdgbnssjL0B9ji5Jscc3VWQKYXa2O52z9xLiccARkByu
GeYrbHeqegbMzOdKaR/F5alESMfazgtyTK3sRKb5q5AX8N/PM7LQ6tsM6ruXTn62FASrrXeeDO2/
9StnSfzapZ1/INBMbiEv21/92RDrXMAsqyj1Q5fgiHDkUXVwdAvv90EYoCfXW2LwuPjmi7jr4BS1
pesC/XaJAg1GbTOUKJje1VmiM2Tux2a/lyeEiYKLt3qt0LH1e19lweSkUc+rAcOfW6RJtyTNzhjR
+DXCh2qJIWwJ9HWS1120DFrImYTN2+Ml3KqvorBCPJrBlEdf9kqplf6sQPrTtOTcvtJCDOIVaOYx
EILPJynx+WgCNGnIUynQMidioqDNeDSn+mNxVwQ7sAaWUEznPAPprRnxaYDVdHqm2b+m3OY9xVji
d4EydcM04N9hrh2H1Ycq02vaLC2VuiNrs/bmh8YVtIBpwd0jwQtIGCtbptSer7Y9/iy9E1OnMcsB
/qsXdcBAIFro5I9hxdH4veThhiQGYTpP2rj824NQ2H5SxGm+hvYeKdcUwhuDsXMAoRYPo0RdVXqQ
20FIewWdNjbGwOhIzS8YYvWqfjdKVB4CtLq71IBn15PEcTw6w2WUU5W8xSuDN4nkI/7Nsy0cVnTD
H8CwJ8kUR9IvNGNEliJ3UGJAfriNKWZwlHSHJuaCczr7HAgcpmO8oaz1AjgPNZGteLqeqU+CUMrk
yQJV2q8DUJBKNzORSeNDuZsU9ibPQiR55Sj0H9dYwbGuT28zI9J9aowSCEGViEzk5iNHiv0Hf+YQ
ynBcIUnmuC/lMfHsdONcEVPvRDMR29q4QjBP0Wbl7oX4QAqKFEupk+7quJcD6TpmBmDNmvvYYZtt
XstBt08be0Uv3W5Lx0TflfqvhFPXVQxcNlJ8gYtdEVNRp8gJFnPqJ/NL/VtjUp/SMpxjlSPtgjDV
XMreQoicGdDpJqeqT1oIoYe8G2sc3C2qectGUvCZ/KHAps7VdLyUn8rCKBy1QbWeALvQ02mm2Vyc
LshKPhwg8kH/+TuHC6FYpqsSj2iLgFV/iRdQ7ksgVbwqFDY74NOnx6bduqU5FLQrEL7tWvK+Zcdw
1PjrZSigyQ/KPDggetFM1tpVDDi4opcNWtzg8ssQ93J592Ju+WeI7PQlStWPnIT5ux4lbz1nSS7g
p1s1V/cnudeaX2izjXXNPP8JnyOLJsZjQ3HCbNvnAGf16kSj5SbSEKySCc1GgYu+nBOZnEKhl0Bh
0s7AmBv7OrpL0u8swPeJjuUibTcAXoedoNb9BmTgemGrluDOzcV081issu8/IUyZOWm9O4KfCAxE
t9mUw1AL0cZeGNeBgvOu3VyxQgIfU8bEeVyaM0d60usSPh18MIzE9mwx0ehFbcUPiH/sz3szltOs
TgEbB83q0a0IXx49ZYq8W+NoOqlXVcbHuN38V4aPWBkG8yMGfBcD7pZRgKs8ca3ZuvJSWQ7p3+zM
tuDVFsNM/5DB4jtTEoGRcK0B9BbQl55BHOMKsH1QEVh68xZTrX33PqGca8TB47VYsdpnYOu2YcIZ
L7rf5jo3+OiYf60u3eWRdLd4txZSgDs0+8D3+dhR74Wv6M30U7UYEX8nXJ92a4sSrBHdvCkULGRf
OfBo/wpe585854PW0un9g3L2JPnw0pR/m/1qHVkqgkha+vjTp8JalFT2JOPbMVeGp3jgXPsRaCY7
YEas3I1KfRBybqFF7vkUMTs/FC3i9hHxWtBG+2yHb+llitt1QenfTDal6RIJ8yeZIMeM8JjwYiKt
yGtyHn180M77XtCZXzOP9S/DCisHJX03B9Rmh4z1JyrW74A6JMOpD50HYweDZBOYl+w8GKU+OFRr
JcB3zsQHwBbygxvSYTXth1bUFYWpBoz/AFbjlPJOYrsRIFYK05H8MFU7iUWXfv32PK39ynndf7p+
cNOIvqRioDuUGytBJF4ALyM5JXDANb3EJEIBBKlVD1tjqQfu88F71Y5uC69SqcbfAtbSWePvl2xa
0qJ5KeqsKkgBF2JlKcO2pLAJB5n1nK3qmfQS/dDj7LHBZ4y1umK2amCUoaN4wLy3yy93aB9cDyLY
SDalgJqyYZEe1A6YcGm0XcGIs7Q/6xPBD7E62RfOgoJoOcnF6vvrSyb4Rh1cqjRGDEtbFBlH/p9M
J1/eecGzFdCZiTuFBvVob2EZTodMEWpvg6eDWL3sj1jpnjquWj0KwDLTCqYY5g7fWML/g4kQ+PwX
LxCHOvCRvbuym8dE6vqoFpWeEOVwKutEZRhvx3PM4ENbz01io8XIEK6Uo6uklVzHxXgzboRYdWLY
qJexfFIAlBJ/+yE7GZlHpvQVFZvIE6HCoo/3wEkvgG8FeBFpqjebE3U2a6at8xUzUFm0qoBYenlQ
RT9wvJWIyjtAIwTmw2O7S3C4CHPq6P+AthPy7k7PxmlTHxHNb+jvMDGePBqkYwVcoEwPCJCnL+fv
3lt67Igt2GmM9ZiyKQadgh2zJ0lNyKhiHael3O6jEZTIVCfaKUwj61cYLI1me/TSxfh2y+yzPkDT
eiUnKlkg1ZWhsXWwZwhNT/RgZpFDHGN3qjEf8PNZUHCe+GpSdgNmsoRndbDzX7udTzSMb37faFaf
D/6WYzrOqdXEUIV4R5WgcC4qh3Asxv5/1UsmyNpaGKk+IVeOXwgTOhCnNfz/QP+mzvHqhUJyLLNI
1+6ONzNUIlPf47EwtDJw0Gr+bm4pT3ZekZMmnNpJFje796Z6h9lqKQv7Oh1zt61KG8EJS/AC3Rzi
MjOG7+WcfG7/1Nvn81NmWtom4hlNGJpZO9lHTQbYaQeRuPNZcZIFY9j7Hv1KL8Vg3+0DMw/h8F88
nMMTHE4Z/o+yPJE6Dexk1g0OZ3Fy8X1LO2wwCqzWyb2/Ur2AsQ6HYote/JUUQtN9peXFtCRw9Imn
1vTMFPbIiHZlbR6e14/mGQMlAbsjukm9HOJ76fP6S6/lwu4eq29cXOqcOQD1FL8JsWxeX0V2WGCa
B/lq2yf2YFu0Wo2PW8R8xq7TCIkexF6wybd911KL/iT0U+ziYRFBPSt0SYyRoHNoKxwrgsAPk0+1
+ZhqTrTeIWRAGmU/CM+Eay6G3VFoMWmWORJU475lqIhZc5EsnAi8i4GOsBFeQZzanpgyx/1Spt7Q
jkQ0+LwUqYTWqjBV9vPnQfIudqJXdh05+CO6P2FtuVmkvD482qv4MZasgsmCy1m9GOyP+Qzy7oXj
nSZgNJDfsg9vbIkhxTkw9Iyx3Yrmndzv/8LO/CcLhHrpjFwTIsuUL0oiPwHdyWsO7togFDcTVaXy
JLn0mVWsqJjyJOhKK6OEoBOopIHJwPxHLlyU0/RmAVYF4Awq6FKLUKq8QlIVBdEu4EdfHAuxasYt
WheVdgWA2n9bzIGrBbOT40W64wcljBSHzSMPVz3dqdEKlkdWNhz3RP7f8XT/Ll63iMJb7w6Yt0ei
UPJ5cS15LZJGx8WcO0QDirlv8z1lHcjDM/qfPEiqfsCUWatPggCiS79hYf8TmPuqOCT8j/TXgDde
xP7x3tG01oormwDVFKwXuRurcn+BxgjhYNxN/PQzHrnxz6Gj0XcI4Sg+bJ2+A1ZNfFDOmt+3vHL7
iQjBUIIHUOqWOAk1vv6Dp+tXkD32DVRLzbGDUN5uvk93PAP5zqwVDhQT287ngDIYPYEYzkdxcf7O
VsXUPYyeVQSYwwvIy+EC/n3Q29wQmeHJJaj9FGyyYDhn5Y+skdIOy0N2YX/QrJ6g6pGK8Sh/RLq1
u0z1qvUzwqq+ECceiovYKePRkwl9kDU4iMjH90IWggF5bFvaOhQrmQKC2Z3xu2O6Ubg8XsSUaXC7
NmKErk2xqw6S3jpIzFa6BvgBQOoDUpyj5I1s1nObKf5VpB0Ga+KrGYtY2S2Y5gGWxov2gwsmOU4z
JRwhpYAARfd64v/VfA1mOWMn2U4/y6Khslc/583QlHXFBnT6FpLQJXTIjKlC/If4JFQiORMQpGWW
EL+4nodAS0tZSmrM8vKrDM0spv5wtnjjopL/arnQb6l6PKjUtDop6AetOeX555Z6mAWG3BgHlVxb
7aHv6lm/ZT9z0PXQNr/RXV1AKeMSZLmqfYB1FFPGetc4TlfajYR4TscsdUgji+8Me+gyrV0pjb5t
Eylbtu7IxlyoN3T+cYWfYWm5FBx7ssuH7zo7f/n+bku7sGBJhVyg8SSLKUIkBAkc/8vc5+g4h0cz
2Bzhg/iCdH2x9SK8V9gzIXDOytGZpUbOJoiTECiJWvEn2VsZOlXMuUE1JIbVIv83XQiJIdURSsSf
5FQVMJKuwDim5I0rayToZZn6KKyoX4zGqnZt4f4Wsl7+wJsDNC1danyiwRvnmTAD9GeTWf5DvHwf
fcoKSqPkKMzRSGOERGAPsfAPWThgUxJ8kwah37Hq9sXANCZBb3H+Yp2mOM4x8xRknwFdV6uJYsSM
8xxiUtNUXFa8BtodZu9J2g5cvGr8qv6vwEImXlJ0VHnWJWHEjNqI2qgCIXt+aAr9vIaMOB/sXvt7
ewbsoSZJkBC6Sj7AynuqwkuR9KHFmMyW/PyQ5/3/GXUxiSLb8kViYryCp8ILGY6bYf0v8dlvew/l
TX6AtARH9JjIbOaH38t9Jy+t4cWGMOrb9e9cMLZblg2obEvgLpdu3cLzrLZAFEkmJxnTmKJ5P+24
LNwfntmR63E6FgUT98MKr5dU6jRMLOnyMw9286Q4S44N515VXLATn6cGhb6ZoIN4Ddy+IedREkOa
hncy5bM5JYoth+gYuVy7SaffwsTeseATW7BsEsMstIHfyY2FPSKICOEOvNoQTzbEu9gWmYSSnYku
7Q3hsL5RzrpBoz4e8PqWQDFiK8kox75hyt4qrrN7HmR6eGJhTbFdGLQX51V9PaaDJj1Qg1l2l/BT
zb+cqHdZfUK2iXtgpOo1QBugl6V7bbXgEhLm9rFpzl87Oy0ju9AOGQurKXPm3RVpz1w1CedaffJm
ly259q1ut6rJLQii49Kw8rsaYwJ5odCGoyOHtwz69upClnkiArrJFEhw0GJeURlmBqtObkE4gR9y
y6e5DqDFtqUeh01WgBYFq56oLi9oV40rQcPjvduwNSHX98PY3getuATKldQDPfT5vKFA/lfP/9XR
WjkHm+3lEujOQOAhGkZTKzjji+F97elnLF0THcfpvsXhHXK49oDTwIgHEXmEPnxFgxVcLv1HYmAe
FuqCM73ex8o2NtoAcoiEvxgA1iGOPurXfAy1VCKYifwMOlypy8mQoMuGspvwVM6C5OO6/6IuM11z
XbEvAQsqbkfQVLmprxH9C0B3jx2O24kPnbmcyiQ6G+G1qZuXkyHr3NBcLDLotZQ/vt/uH8SPiydr
dFOccmtC53sI9vdvmR8Hf3WIGb6qw8a8xL1uze3n151K7Kh/ArvkYzTh6HORLWncyh9BTaz7Efi4
jdLHVdJ1VUiBI7pLsQHo6Nq+SzrrKibatvozdU7CMhqN8hxgatXJmvACxaS4tiJUFNY23DysHHT0
On1VzZbTrIYmAmLRlV0w2OexqyJ1oIoe8v7ehtVvDUVD7CeSTLL248mdJs0GyukwG3HCs4TcIhrr
gKAc0Y6VoI6oKd7vKh/rCgZqhV7FfnJvpjiJPXbNjQC14MVXb0mMr6FQ72C3BBwH/NC9Z0PqvNfO
IsYiQTufwheXGEdxz65Le2vixxAX/TRu0w1NKBROwbk/qFmcWiOvS0yWonylsob46/4NhybWnD9Z
guGQnLT+3KKTtmmDsYoac09LKpVLWbrtKZKe3kBsnYs5UXEXXgDIZ/I6tlT1qIBUjyAyG29sIiKC
Qp/s4v8iM3tqR4vPBJqz2+EM4Cd1Te9fu7McnKn0fzlpraHgTmcFeSZ8bkJPqJv6e22pOFMIGBin
Iw+IwUFoS4Qat85XR1S0+CuqWqeXtLFG11FDLn6NiHg01/qnrnV/xSgfdBhedRikuQJ7iwwxiHRS
Z3mL9uvPGfudocgPhW+rp4Og0OImMUnn/PRzArk+2jHCmbimv8B6a3qV590sCRmx6jwsuVFVxvuF
a/4pOSbVZjebjt9NQ4t5FNFYFO7xt2iUbav1PvhEan9WSnSew132uXBu1EFCzKFKYfuGi/QDUBqZ
iASy4BM1f4EkIadvErS+95Clt7s6dlq/We+LDo5BhNFM0GcBVAqY6bErUQMltZmD9CZcZUkUn/5e
vKWY8IwC86e9AsxOAAb/wFUbBS+2ZlAcfNcWR2tYQpbCbYHMRdZ1gKZ3g+kq6kKReeo9d2sZJWny
2UIkz3CxCbnRnTY+fkqHlD1STnpNapWHi10Z3hepYH2Y9xhik32FhsHb+VgnDyZbPM/NG8a6uaux
m9HLmw5YHDcaHisDJYkg7eMtlMrS3Hi66CTZsozP/0prpy5iBEJ4nk3KNSe6zz5mbsmohl9GIc9f
3FHhMd4bDhO0Ljfh4jhEps5eDNJCCHMXIbCGXpElskCE77qFlRrJSBO7b0nIwUjtpWR1i5Pi1zv2
jkEG2W6J9aVUMfz7gsIGt/49TKVdnk4sYLAIO5XVoVJ6/+W/D25rsL+d/AwCyd4bIXJOSq7nAaYe
yMJkSZ8+6g/fXrPtKvOjuxuFZvy+LvzaT9tXTHuZmH+74QvV889tW9OmyILCb4wPeEM4xqWB9K+Q
WyVRb31PD/YGtH30aNSYsyq8mYrT58kXV+hYIU5DrJW3bNq1D91qfsgTIWbrKl8pMFiYvUWqIZ/k
N5NoMcfw/pqNwC/Nq5MbGz7w0Y6oIQdJ8Xswc0qoqnrQwb10IXaLYIE/A7VbViNZnoM1iS7dsaHs
rDqQ21ueQ5rtCNYlMvNSRk2C51hjNpgcKHnNK9dYc/pb3xEyO0NKBfvCi4pF9cKGsFiJLhbZ/Jum
xbMytOYAJx/rZHGqF1Bz0aP8wI1X6vAQGpyfwaQ1yVlzQKAoWtYSYZnVYdldCWXpCzGEVrhBINpM
MRXEGa3ssF/J5PE2L2iXu3m+SfqLdeC0f04VzEGuZ7YCpWnFhL++eHNhhwzmZ01OhkF08MHbwph8
V8Nr46Jg/s+gBNJNY5WwBIKWj4klj2ixzWD10l+9wlxbdjn30okzLcBBt7AatYFXpROCpChUzXT8
s43qFIDQnmjBPrrfhi2L8pE2IjJuVWGAkC6CP+OJEePeWJWGnk60qXMGHxdPFF6R13c9z7WhdeRh
Y/0XObd8OTv9RMIHBf+/6wC6SzQAzeU2U55JaPUC4HLMBsSFmK6+xxJPszeoYVB6NXh0uFOAgIjk
c7bM6R/17AoDjx+Isb82YNmmVUZMW+Jsg3K8HWvhgCRaxt1rptCTYTeGjiqm8GJkz0GO1+cdFJYa
NkCLA06EW+q/bzzEoJw8xTyH47jB/LNa6I9dXwlO+tUnCu5WMVcPI2bxfoTmv64YoARS/0r75QZZ
16yv20TtORahHhwQX71DpT4eOLKC07NE8P34GEScvgNaZrr6ViWR9VOH6kvX5tJnG5vam89H1jNf
jMb61N2PajMh+CVsKHkcrPjr2mwFtuD2PUKkRKtxVsBPziUQhGz+NSv0F4KeGibfBVx/5aYVby0Y
g+z+bL4ydwYBNbCOfeN4ODDIY0QhVbW/oVu531gc4S7tYMpkFD+A+9QA8gTqqNyzoHGxyjSl/eOi
fZ5RXE6h9+P22bJlWisH12Yj9k6eHejY+9pD5JpUat1+wa0T69Z4jkJJugB0gP5dvgo9RJ4hnRdU
pYeSlP/3BUql0yfj7KOSfK2pUrRH+4X4AGjn/d/iX/Qh4gqbrfHNIX1ysEB1PicGPTx8NPXNlbri
/DkfUx6Z2qfkjvp7wCV0r8VSkb1T5+6NswujHy7EsRZ2mbTwGoY5MrHq6RULR78+TzVSKVjMCnlB
qgoAIrVZwLOkBS7I1291A8KfSI3+HsFb/Ws7dLlEzjtXGdC42bUePqKxtFVdt8lElEldV0bNTmal
0UNxypRMsIIzJqM71hMk8WQq8nQaiw0zhHnxwKEN56lhqx9Md4IZxuNvjIGOcjw20Uh3C9QkK07b
z4CEjvERFM6u7bTHdyg6TI2mxl9VivRzQaX/vDogbMFLmOhYXXgLhzXFbERbNzfA2FjqQxMIuSVo
+kYTKq9djW2+rDAXhZEC07UXQdzmfwofUGOwWCtNAAJZosLI1j4pioQjUwPPB39HC99UO0/J1iN8
wyDIc1LgTmnehAv2FPu9mNs2YgQgHa3CwcRC+bgFxAg979VrmVCe5S5LlWhNYCyl6c+p0fj5r0jA
FDDXp9hhPFkyczZCY6jJLCWYljGfjiCulfBfapj+kSAouNxqwK4dgiQeNUbXmvHzya/9TWIa8L4G
m1wAskV04GFgNxhBbtAaYn6IXXVBXj1y3RlLTgiXZmA3gZYvDm2peS7fh7UPsHIH0EV4wG9iP+DA
TV0jechqfi+b3oRO5RiAlSReu8tJuKaUHdnAIuY4LyaTNyZPhiGHYvZ6jVceMA6ghYhtBIsanMln
IYnUugZLyDA+SuJVqFtes0h1QA3MK+V8HV37OCtu5uGC1wjUvVSNIH9sRfDRIosyGi3EEnClS4nR
ExFCT0gKeAcBp8uBinbvGmjrj73RD5bqvgi+19jKMzwDuMwdAgkYoa3/E6YsObjX8ToJvdiYNS7G
vbR+At7lt6ADd8+Aa/6tDKspmtP0KBF8P/4ruVdbeoG8Ss8eYJkH+1aA6VDuARZ0BQJHJF98pQGq
PjsjQiwnDabsmE1cOSS2HiG1ZwxOQAX+XyUwAahncec9i0xmyetO2T6oY3VUJxMHMz5MUZuilE43
jujKi8/XwH8eSs0EwO8Amrp+JB1VG97+WGhYD+fqB+rER+I3yugK7ghehybXuNRSO0DGxzSFlWlx
kCheOGuQPx+lOrZMeOJ/kWWlxLpc8vgoHsroSeqDp+3Vj+w9l5FiEa9RI9AbB56N1CQhICnR5VOE
c+IAdbjh8hA6TZwdeiYP8yVuCiTMkzyhkz16Vs9sIJLWuToG5Y9e9kaQOQ25UZYCg3faCgrPRq5p
i05Ms5VowxAl7dSb38R3Wpoh3tkEHTEhpRJpWmz9mqOmh4SMWVsdT4zePtyWeD0eB1sCNX4Q89JD
22lehJfAT7X6mCPqdzbbe+AJHcRwG7/ftofkHt9ZVJHkcTMotSI68XlgdNXbaNcankMh3Lvmq6JE
1ASq7mn/Sik5kL/sKk+RVN0waD5JbRk41UtMJVIMkUosjZT8Y6V+hsuX/0nRMHFXRerPRgqWvZ4v
dkEqhElPXUzRWHhNYmkBkKd/sEQQfzCwUC2YpNJhOClX58L2IrG6dNpuIP5lcDhFxxI8pgmtxmrF
YT9d6aUIXc5fD+wqiJ9qPNfvBSTRr7x3OyOc6ll0U18nYKtU+/vUSMZwlcl17rUqYbHokp+TIOzI
YS5fYufegZssmcE6U3pLsISIWAkTdRwUqIllV0EKUHNrkaxeo7wP4f7c12susiOyLaHZxOt2XRMN
RWU9BnE/izoaj+aBSiiS42n6rYp78cDtFYCMxS4TQiEHvJBhPyUZTIZaVac4pxtI73cdT3VQTBbz
vV9Qk59a2XMMuqnEvojAthggheF+UfN6tWI7imDq1qYNhFo9v3EmTEdQzKiQm1QKay/toKxtMVSo
hnR/E2osLUMtaQVkaL+0DJQC6evC8OqVSplh2CA2xihJ82uaOAWyHTlP3a8d3tnzRs1ZJF5uqY2j
DXcvUXYHPjTksUSekCVuGFzLr4jjKBEw4ScR9CNFMCoIPpjxkoUdiKMh9YYZ2n9V+HLmELRmSGKJ
9dWs280JQw+REZAVVGwoV+xLotzMVxBKkQ/CBzb2Hgs3D8Z30qq19rRs41UXeVl4gkPD4FejIZRr
Sh2UdWndvAT8fNeZEGwp95O0YRp8fS9QiLN7wl16/92PxXvhve/ZZgQN4HYXvpRVr70DJWHTg/Ea
35JBrHqJ0MzL8m4dxw4JVfC+tkMVzQAq3DEZgUzc5/lCM/B5OORS2TlJrWP7+aMICYpS11EMN29y
gWzgQIb3uBNPwY3J+xJT/jAjeJ1sVl69UTUZaWcf/cwbvrz55AabRDLPjk3/qBa+BjpJaFlbltGp
YClyRiK3sW/CfVxq4pRsiQS8h4sMTQByREKMXjlZJm4gYO4rMfKQuIqR6GcEZ9/K9+wbAuavMvXj
oHEX4IjyeqOkldhuYr1wp9Oo8wDqLhnayo7Z10xi6+QXEnWRUvvjVaGyg4BsaKMi6h84E/d7VEDq
1te7PY+NHedSGuF5Zs/wJEA5Ut1rvRIqqgTwtDX0zj2PW8sTklE9oQ7PHqdkDOuy23LsA+Slx7YQ
DJ2TcYreRCNH1kiu4Y01nbax4sgp2Qd8MwMotMn6Dq6MtOVeO0Mtu9aLJKpSZkkK9lxgK3hN4aSI
4ubZju55tFdQ4HIDhiDncRtkuBl+GqDVvyFuvpHEKJiIiGfM2j4c/a434PiUipChah60nb0AjT+g
ZjySsppMUGIXYAr1Z9ZoSg1WaCW7pqPfqQQUZgL/wdwCEAuG1XciS2/0hijj9BkAzK5/QJT+4hQH
cVCR/zznvK1keEmNNoyGB1pcPww2nVDERFbT0qVzWufPjQYhPnozI+czDSmC/AOm6ea2ziUh//ym
5t2B08Lbg+l+1XYDr+Q4/e8kV2qrR8snovA1f5Wc+/jZRdyZCIqdSx6ZThTrJT4GLgNInc1WEA9H
qUGrwmZZ97Hsb3PFw6UlN53/iqCmxc5J3w7nqK0HnKkDPzZfEFmAMdiYTgbWHoM3a8zuQne4IA3R
ze3CbgO2ivF+iyRnZ1HL+8KobGfB5UGMizKjADmkjPndVtzIxADp3SfL45lG1m3mlFHSiLoCeccc
Qdak073FX5E47EEi4naRsuRCBA4gUOYwKBJ4RTwxJB9N10G5SzdezAmbugBaD/wKzFOci+O8oBM0
MCro+25gV95d5zu12G1457QMmJ0uberEiRgD7nbBPrz93BO5u0Tqemoa0wqjneIaRxPACZC50x7P
Lsx0qsPSS0o1iVmwDoJe+RB8Z/9BDkVjF0wuTsJPUqMWCVrfRD4LpY+Qb6RKxu78IE4JFWZMhQvg
ly9zcTel5p02GOm8FCYhyYOy+0A2DJJcbugvVUJcsdSvhaEYPI6mVKntGBzHYT8RCh+ece1eXDfu
L56FlFEuzo9UfmYlDwoUqx+fIV64EM+FN+TEZXmNPK9W5uZAb0mIcCCGXZ2UiR62tyRYu/IziQuq
kHeTbwm0SHZmboIvIgnZKC8BNCK5CYNSSxzeiaYj1JR9n2QJFdl/RomQ3vKHOHNbbrv1247ck1dL
eswEzyG7axrUh+2mQMwXCqsxcP1/TA8DjPXXp4Nj/2oREryaafzVPgvSf8YHVStDKTXrvfkXLYN8
yFvApQLuDQzmIcjv3PdLX1VPN4HV41qNikKJEHYfRhVmz6LJ6FHtul4lMg+qcrXlbK0+Aq6ww6YR
LDN5waythgSol7LfUrxNuzklnH2pUjiF2tdgRFbTJPiEje8rpwhHSdzFlWiyjEkFPE6rPXHWY/Ca
fR2lvyEMzv+KuqQQtGHGg+4Ujywbb0dq4NUX7rj72+AB80xq9fDVbYBn9zzeM06/4qtH+tMUMgf9
OW3eC1FdyohI/QRv3K5w1MZ2GfikaHSE28r5abytzACWpK7Or66o8E9du/o3NlzWC9IMqkC/OorT
1gChDS0gYgy65N/ZxSF3FYT+ek2uBio1J36LuSl/FBY6HB58pJkCL1e2G5vxTy9WSGcD9bo5orKe
GiXZUAt0VWoyOQZVzvSlkMRTWkpwMZtSBLUHRGS3eg2TWC6b7F1qzE8xr6B730VoYNKBxiOB0I/E
Bl1y6PlZdTWft2GNLg882UEfpDgxZER1+zd4pTudkyNrfuERokswOj6FtbHmi+1GDzamHc18SylJ
U3I6NDkw+ckFfpFXjajnCPL6R8Te9v/p/LAoIzgPj+zCd/TrxIZaM8t2THEiI4DQldkUbqwj9pbs
RzBvImCcptG0BERQOpjKMdCzykJjpYxgIOC9/6Rk7tiS3RqKl/yw4OiLa/evacDbrc40uzk6nCfh
wFx0yWeNpL5i65sY++Bi9CkInAIjEGP+Jj8O32XF5xbBE26EGGPAmbzux3gzJD/mipwOxu9Byu4P
+x3NPTc20IMaXZulBgUps3Nw34DcElJoBNbrtvse0GO7r6Cwb/GrvT3Fj7Xij+feDS4BxL9bjEZg
JoaUNgT9chEmFCwQGFvFfoOFK9X6sY5f7ROyzmWjOUaRPCTdQCPTQjqxqlkg5UvsKubDfBIDCgG2
8aQGGQMtHflE0h91IqfXjibsbcEUJ9BPTAnbHFPQtH2Am57qxJFFZ224VEb/4DCfj4C+H5p8cktD
t+ZvCvd78R/qirmwx+tdiF4Hrg6SKGZBstrVgd1Uw2DHXM1hG+bbo/uolzINEXKEqb2QVwMdTMav
Gevyo5/UYd6Yox9GR/IejfeqIJ4rPTkPSjGlWRzRB7hjpi46qgZKouNK4O1JgshTry7dIzbri1sB
ZdJC3s3gRYl99LnIlhI9xw31GgeDqgeWPljxWj46ARWu8PJv1EZc9aUh9onDsEMIFoIM0PsJIEpT
KAkLepvd03sVhkz396Cq2ARR7fSCS8r3/GBbGQwng/6PBKo/5N9xHS/mBLCbVnDhIso4eGO6d8gg
7g5mYYnGljJ6LkfuR7n6XaGp82dpy6LSLeUAYuLK11p3QgPuF7s/PBTZWYvsh8D5FKYr4gms0Ms5
w7X3vDtwWM/lHkK1XnQD9jknjUCTX1qZ3xGuVw9jiH/aTwGbPLol5v+06eBYRZLFvAV894b+tBQd
PT9iTLHCBeTihelzupv4L5QkshswTGvLzQngFmlYiOeko4hOPuOhTKyLaBXIikmC3u5Bd+ct1CzW
YGofuMfBbeIVIr2+FGjmJB6IuWSVHa0ScjwSwGj2xDkId//USi470hMfszWjgZRP+Ryh8rESyx7Q
yBpH7dpxHUg4K1AI+CJRUb/YdN5Nm6ruf+AgYujhmv6eN2j3LECuwDf/moo6V21oZATP9FLYOrZK
pgoyGTN5rFQrSmvpy8lnCkaCDnlWfrCk7r1OsljvDnRM77shoxReIJIFG8ZOmeoX4txkfhZUqiaK
7Fub0UGAckM15Us8LWX16eli8iKFVGaFKxDE5tD1Y9vcc8bMLjqZxoyW7NJdfP/Zb5VZBdRWRT6F
6mUgLIW2HPpY7JElMNHQR4GCov+ZDiH2PZVqSwMwbSshL8cjmC5Y0qoEJIYX/xnato7yA5gc3zGx
X2wmRm8ubP1z67gXmDq9f1CZ9NuDpFHgSaSFEvU8z65u2i70qkjQN7CbTQeYfV6r4FUDhp/ByvtM
wFFkqVPBFo1s8JJykBrzsDPBy4T1nilfDE8Zyk9N0O6seFSVARn+pe72i97BUAdxVuwqUevUnx86
T7GQnC51sZZGB34IJVf2vbGGiJcdlMj95KDb0hBLI2oS6Hwm3aU4DE258+ApHaogGCYoXrUmqK6P
S6XTqgsIwkOpzgz507Vw5Y8BzEiFZzqVVntTHGUuF2bFrsNJCsm2E1Qx8gfA6UiTBBlRFoAxMjug
UN820hyJ0govDfz1tzuir1J2opPXid6A1oMWm4vRXnbLIVS5V9UF0eT8+mcq0TromMbpM5ORXJ7p
lZ8YhzinwthwDe+eoKBv2OXPaHB1tvdm+ow6SBSN+kdC6GARUsrUdIeFANK27cXiiRNWjTSPOY6e
rvr6db7uUhcvXx8HwM1nQkvEJooGEISsLv+O0k6oycqpRH1UEgQpQ5MWzIRtKXai+cYyx+BhnWdf
TjVvYFRLDvJiCMvZW3HEMWZf5T3g7ezyQ1Kv4Z9uh5bDuo9SUSoe3iD6LBVws6C7zPXye+l081j2
zbBZQnaWfL0jHdTwcW2UNoiGVzJjN7+2aluixD+SP2mDyu2MOA1w1dYfUgfp9R7YjAC25g5ypXYj
LLytKXdWkFXv0AJF9Exv8KLRP2A66QFVmnyjeRB3kkzg3YYrqoDcOTz3/3ZaSo/wPh8Qq4djxljA
FjZFPGvHViAscFof8UchfYZjQkeQy9myX4xgkJMKZwlsMv+9rpew68dh0K0hjdhnFxKMMqGnO1Op
8740R39UCIu4wwTGMSt+ut08MqTMZOTD8QQ999PtqyHLHWAUt6zcDT6vBAbzdKHxw1hR2i30zZCQ
c4I4r3SWc9ESuPdBktI2l8GHuFooJKKGd32VNU4lkZR76VOyywvw0yvhPYtGl7M+R/9Sgo4bWZsw
URgkN5kqfrbC96BaHMGRkmVdBZYprOD5dNbQUF6Qq7i8pOvMPGNw2XBrL3/ytlq4z+2aQc1PBCbE
kf88eFf1+lTBx1Zkc+9XIk7ciHusTfMcYhdYxQ6P23iOj2GMLo4OlYmjs8ZlEW0dJQFL/aZ0O72q
IeMdI/stDnr2aYr6thZKg4KqRSfEEXurfbDN14rVohIEByth+AJOQis2cHjjCE9AzopjrsKKAmZR
EyIprzUmuGE3JqmEEY4S7zHaIahAuUYcO0x4GM7TNFl3KouUgAPyZntW6F+Pxebu0KZxRKaHvt2s
ackQ9jOjvIEe3il8DFkHpmH9XJEXG6w7sXaliF4lEYnr+pvHC4neN1C4PXOYWIunr2UtT+9nvSxk
6tAG7MerA98kUuJQZROHJzJgIjkvnzuGzLSaSylLumJirZ5gPGDUtsIS9NAw/uS1139DS+UPYzYG
w8x8cnOkgLibLgu1OAqotkj2hAsWDv40scEKwkn5qdie5cpLWZpX4pIT2EvaK2r+eBEsNeWfD3Dl
m83zlw7KnRGw2/F59rPENnxqHJ93RzNhvyQRyvm2NYi0Bi1HpVvlktiA+E2HyVeEKOUXInsLFRyJ
MAJRo8GrD31Po8PRozFP8r1Rk131MlETqiq3zHUGnTt+1yGEHKCrYCfR7vPAI9j4sd/rq4j85M60
Xn9HfL8UqSGsyfr1aGR+0D4CCGFHFu6nWT/GdAHD/HCs7CDVuUBZeFEYiaN/SLdbhoDauwmNshXC
vCNMVTfhYJ92BZPJMF8piQ174RMHQt/B7Gr10gkHiwVsTPDbo9RHx4ISdhOfY7DoJ4K7zLWpdHHF
4THETyRmSOCl2e59jsVKsoSsC9eC0e4ygLYpbEICrG3gK+mwNdbLvqZzhLKl0M6LFPzT4Pppcohv
LddXZ+QVTzUsT0N3KjztJCmGJrLU2rtsc+K7y6HC4/lvefCHwKqHiY4z2lVsW0V0fTFi5ckwKUFk
GzFHqJzjHYASz/hT/6izMdA4DW5+klUycFYgh1sdoiP54+AodSaz371Sruuf1k38WDMbgCXMzqht
cMX+M7Vl1QvLZcwMZN2/RQOwmslRfA33R3MAikLg8VgzjlLCqIK/1YZOz3QRM2MVK1MKyuf+NvK1
k49YfalsWZnmIvmCGebfUqm8zkR1Hq9slnRMRerQGtJgfRcPgB5OgrJAdJiXZnNmRwnGn4hvOxGI
X/hYymJ/HnNBby91ZyX1VIqHDWkUAA1h1iqYem4+0L4sVy6VyVFidJENPbStZCLmnU51kv4M7HBP
SVMXkvNbh+3EyeQ5OJM/pfAgDh9XPjYVBhAjMVCNknJEZgMwgw32MoO7Qh/BlaLXKJ+ownWMGv0U
E5DH2U5zdfqlwHbD3zVCUMTK+Gsdif9Gf8wMIOwy0hYS+ewSNukZ8oi+zLLd/SBjsB2PvosmyVbe
cVPTnRfQyQaCMqfa+e4CsqnxYF33FgL8gj+vkQ4hwPuIP/tAgWefNUt8II1jMMp9o7CKCsByCLmm
9FCpdAM2PEzSB+uRs8w5JwILGIX5HI7xFO0Gl/FtbIJp0gBkYMJfGiNDxxLUuwovgUyAwgHmjGrP
HEr7jwmCnDZg+R5ox2uGz9i/NVD4DD7Lr8YsH5rR2aWf13jfMFprslj+1/vCCrJ/jxT9Gwb6KfNu
dpgave4S+4hzAnEnaCkAh3+7nWfqJqb9be0cdyuNyDetzOz7gCluSb2Wt6FyVkh2LV65P69l73Xv
K1X95xSEDcYfjY5gNfjID+hh4X6u2ZhQDTkC8j3O3+zFDMrULMe5LZIm/8ZZ3rtpRQsQIU9sATeL
UXahm+uDgN+Rfae0KVzIuo3JAjK8dmeqn9XJmUb7+WbiRKQeQA5rKhhIgGlDlJT2bYcyg9QbngEo
oplToNBg2M/tFmhEEAYxFdUu8PYj6c3KlYaZNGM9KgkdmYqWbzj1zE26enx5ijcSdSt35FbiJrPQ
6yL5tHWQFPtVUVzWr9JO90wZCbRylolOQGPS2m2HS3OVduVS7XhibV7QnSycnehZNemrCp1ySnJN
a85yjV9lTWAGtKy+wYb3AFNTnuryrO1O6rDw0IxUI2GIG86+W9YTpODk24htm5ABaZLowqPlNx2S
UeVLDRRyuy368NE6VO+6/MThHcnBw7yh4dSJorDwqiqavNX3FnWTqVHkoiQxgEY3H1L+LmL7kVVf
2ksO1pquVCfQBcyOCQhZvhVvj47EhRoy+IT+n/G52+xPBzcx9+OISJpbR1lNhcbMz5NfEjLr8QCI
BWQOdiXRVvrRuaWIjZQsuq4dvEhHYQjGbqSrWrl205rMA4SVAYMRDgm2XdKCzGznHL++26osfCAS
wiiWwemc41207GsGimVMZxpcfvrTDneBumMBY5MlYYdiKNe5B/HLk73hlFFH+y14KsqUDe5l52VM
6jvg1EKY+r9iZU92+OOAlvRh8h9MWNHBi2RePt/iDkmZfCEaoHMLmBYEffk5iXyWVRwjqRyQ4Yqo
ZNikJ+tztWlTeuFPPtEaCOM3EWekT/swsZTOVfpJLBWGmCs12u/LweAwl0u/5hYISyfP5ugXbtoo
0X34UxQme52pJi9cMpyYjmfuOQ80CqLi5Ld8hwVi+B2rpxYoNqRjVexuR0bvm1Ecl73zyCPnQp0r
vCpCONwQ5oBScwl4RzVI+ZL52BodPTDHqWS0W81Kg1ivYlmK1Ctk3qpdYamGapnleDiA9k6Z+LtM
V5cEY/vWOvWFQnrdKKuN7NBA+Bgo6xVRsYi+jLxd82D+aAkb4Wz0XuUvZLTCBc4d2PEof52O7tTo
xmKZjehKqO205FEG7ZPBa/aWmP/SU1rvvt5Y83PtYbIbfq748XiGg9kCQTbyLSWG2nC2SLR9H+VG
NOr9dmeC93wnhO8uGDFEaOSwKspNx3jcWOw/urSyYoN6T6L/WiTw8Lz1vku5J9OUILaiF8WIXMks
wG1pWZVKPp/669K1xmrPFZULdBqoTLML+xpKJjZURnACLsPiDi62u6Ouc9cT6kCMX6D7sfCkrB3h
nfr5FH9Czjfqjuct/OPqsbweIuv7rINTb9NY8hXmys+h0YD8/U6TyJLMOmLcmOdgx/CdqrvUK8NF
oYBJqAmVVWkr6JQHGTgr68YCinlvuvy1XGb4q8/MEPW1WfwQHDAdIDnY2Fxo+wt/gMETHoQQHAlN
sE3BAFIphReAhMKMoy/iOPwwHf6w68iX7ci3Kt59Y7sV1T3vGj17yf4a57KRSYrHDALnLoCk/g90
k+IfrI6jQOkAel4vMgSm7vM+HdQvbtHVzAMurPTg8eTR3bEqxv6UooC8h5/hmKn7YzZdMQnyseXH
xFulBIzFNnqhoDiURMNUc9RQIGq2jp4UzGR1uy/JLLXxXSqIs52YBBEsKbb09a8jsxSrmbROK9zR
stSa0BT6TePvECa0sXkK1ceiUwGDhooRXm5dLrKR+P5ROZEIWXC9OHbZJX6H30K5X0832MrNPh2q
DOEpi3IK2gyIHpdf4rnmmdDioQJL+UqaUfSkH8Bc+UVhRKcKEIbZTPpEh/OOG1L+nuNBu+G/hVbm
bC5E1hqQp6k5KEtklaaMFlhXlohg8l2YJn+yJfo5hJG1Ak2veUdZdYmbGsZ9qVlG/jazEHG28sGA
JNIYZdI3Z0JpImSVP4T+3eLE615unoBdigjy68+ZZfPTEyEcvxKE8lGgJeyxwlDfwcSe9OZ/YNv9
nAmotgfJ/wvMvQy8DY005nxa1d4R9pGe4TY/C53aOmGwAeMdEFdcGeI7OMVSJ5SQgZXGZ5i/YP2p
u0E0YiF4rv2HPZcVHeDR3C7Fcc3kW7wXOgwS9FbNsDKJ78XZOigQCAmh5cZfUtSNtnQU1ceB3CRO
4t4qUBvInKiN6QG0oyjykR8cnt4f5mT0M/sQLPojf57nzuHOIq49wTFNiP4o+1Q4RJd6NbWv45ub
IKgB76ydnZI8e/ejJ1gvOawLgihhB57aSdz3RV/JD2RUzhar5wsVXxpv97SjRCJX5G5qDYUyUCgu
okZdpaD9y1VudX+g6jmbNPOdphEVlSXeENsKMu8ToF2wqS31G1YqWzwo8Q4y1XyO6x34Qetww3uQ
WpIXa1Q4pvIcDM1es9g6/AbzATDp1rU2ZBKQIT7jNJfSq8F6hyfKKf59v/UOozAmM9n+LMEzdYOA
H36wD7L+DcDctN44+s+pTP+LKNpkDCKODt3uG+gIygBgCzu9q9tI945RXV773s0wTnXgd/0khert
pepi013M8oGAYZ8O1UfeYRudnUpA0+cLsZNbYGAAMg1lIVFwzlbXE0EKKQZe1bMTmMXRe8/owwc0
gpHso2Sae+AgOQArDmnB8Bub4KTezE2fnJqotvzx0xhsmrCY/voA0+hSeNTxuOBb6XecF5GG8P1i
dBWEFge40Eft7QjZQDHEKfMfHnrtJTnv1pDUrkZc7nU+2joiagmsCy+5x1dsm5mSVeCkwtFOrqH5
Sa5xjLenLPoq7aIuO3QAPD/EkXh82oYGDOLNff04UpNpgdYuwqP1FYb3dtadt3aXYHQnn7SKYKmp
bPOZu/yohrL9Ui7gVn/IPWlwVDfYWFVZbkQp5SowB4udELgseVmbsmElqWjY1WeIOqqF7hYap0FN
vFflIyGHqbLkVC7eqggVWax/0OOShWUOQnWqCjm9UKA5ZIjgopeQ1fCkOQbSeiUGRAZTG/qktxud
PcrFv+emnibrJbknyKc7NHBmS6BsP7m+CPLEJNoeGnHq+gZtTQ3jRlggF5jXFucf0rsL9jreDPtA
Fk35ojtRnznOAI6Q7GpizYZozMykPi8cYf9/l5lv1UzBH9w2dmfG0y31KcpFAPi38Cb9ZRrHXke0
fncEWgPJ7l7OrztAj9pcil85HFj6lXyxHn9d+TSoYgV6NH4zMQMuX/h+ixPXXPsco1VC3otfYKYO
sKrvQfWQjGcG3c+34FzUBgPk7IgWvA417WqcidwIICOmfQDUxvKvq7H5A15QrbEg+patI2BfVKvA
ESFyzTkYEAa8xG1VR9dkzAqGx2n+NKUG+W8G3iK1Z1j3sPi7j9MtSc1WrwguIK33VrH3ndy7HOmZ
bXbYyjM6LTQjyorgOHXVrWa+50QjO/S2/sI9dq9PdpkkCwPlZV6xBEInq86YWTdZP32811EM4sF4
PC1PxD+sSKZ/fYZUEEBmT64a1BegnzhesFpvzMRDKeHChXsVOqEvsyrZ/dldRcEBurTE4z3T9awL
cRGWNRQ16TUXOrl9gt96TWx04/kXyhwNr/r2i/O7ZZWpCJQeB8oMZMa3vpcVq8SZ1VVmZNOZkNkx
VhMHTU8ge/LglVl4bRkMUHOECITwMWpUYFi/mDxWWFCtt8CQwpVIAJjddcK1ibOqKbftSYwHkS4h
YW6HAu67+TAmptcFatYeAO+Iy7CG8yfc3y/QUEOFlrpyvEGpDhvXMxmckkAaKTBfHeM8NW/MIs7A
GmdiOOg1xmwcHCy+ft40YVSU0Nwurf4NBqfVEdrSIPxGYHJELNW47ROz9uoxZm5dGF58m+glLoWl
3wxRbLVbZ8eX5M0y9RZ4mjutHEqmvGO34BI+xJuUjYlUWKTN3wKY+eHDISNKkVGFArNrpRRymYfm
7HWmhX0Ox8rCXdvn1h9dreR1RL05DK6u4Dc0opc6aYGgOda/WkaGTnIv/2CXtkktKYsYEZgzkApL
0DSI9kn1wuVyjeyUmV5EUcmeRMlWJd6vjroUa3qoz9pDNcE4s0UzVXc0VAkndktmwAs9ghMd3gVH
b8IqfCybBgbp9Kh3gzc0P3UoOn9Dy5QI7pcIdSPKNqAGFnKn5yC8usSZGmaPRw+I0EM8jr+kLcg5
F2w0XshC4cHdSwHLWxljQmys23WuZE0WlTnxQc3b3TdWyroqhrLXVtwN9vPAulK0H295huI8j9bo
cf0hhu8NgiTYfP2AK0OLDdgATAyjJKqyaLh+w3Snr+vCSeKhz556j77ZZaLg7WU6ehcYLb1SsOvr
0GT4CfAzHDGeTN2UXMZqJ3UQRKjYSewkmjsaXGzXUPUjOAASMAb39n1DX9sATBy0eDgD2iDEFAqk
T3Ow+U99/RaJmOj/EPgMNxP3Q/blvjrpIhO3FagE9chjF6n7yHWXFr0FBsJgZ5l2LEDMMLj5VBSc
xQk1rmxomKTRLbiDo7hOQ1gb7+Me4aVj6d4t+IYIX+jpNCyGdXIm7WphZp5h4gh23+Ql9WTvpUTB
QTaZINEThcLvYwSoJN1LlUU8ZttzEAqcLcUAc1xbRFf/o/pBzjGNMIyb1LE1XetaM9THQJl9Ba4n
ZMmNxh71FLok886HVP3mBqixSRMAVNApP5yFoMqw/9RROWKRFv+3hnooOIdHAApf+hGuuKZ8gY4z
NbqPnF/hffljzuA3/bSqfkG3rBZ6aLJU25LIWRF4QSHjsz7Mhh9xJ0u7vfy3ncdXRnQaGVwX8tn8
70qBhIRipOIBAUv7gbQ+3mkzQ9wuSstVqSXUYjbegaJYmIkZYFzjeENrZ60TCwR4K13Db/nKzWwU
8BjBP1dkUIXgc4DpSJFUQPmudOlJv5Xu35kTjVBO/j+at4zpfKk5Oe6mNUxCz/2qrkWdaQzn2QhW
JIVp8ADU6/Xt0reTwSCBrMRX1+XNK+orXqOfagiT7s2T/BVB6GjXNED3vP1y/9EVT1R6OopFBLco
wwNHiBwY5ScwROZFzYjZa69PnqBjwRoU43fsmn4ymRd+cLuapZln9tO9aCd1Ck53dObj23uFBAx9
ubzsr7QSiEJrDXvfTBOS1wTXatc5TEV6SCoMbCmULusKyJ6pW0+QbkppvVyxsm86TfdhkZodMAyx
knAvRqoHJV5BtjY/QF0+L7PEFlpGjvTpk/B5DqCG61AJRJKFFNNn08LIcwcinF8ODAmBNfugZj5z
bFLGIMtj2bRnrJ5TfgWyGaz6VXNwmOqGq8U45uZP+gpiVX94gzi7uzDmqzYtOu1Q8o0E2eO9Ma/V
V7ld5C2p3N3kNRXdMdusaoFJh17A00jijGLpO50Ky3fSKclaNPcwSKRv6OSao/EVQz6wFAMrNnN6
vJUhSOtK9AJKcyLufS71G12IeTWy3POg+T0IXk9pn19y3YVQX0MU+976qu/NN1NTrZD8s6B9/Cj9
PA2gqV6A8ZFIZRlusiYnV1jLbZltswjO5r+8iSh2bKE4NC8MlLWg85oHbe/yNH8Dmv1Cd8KQ7uGf
Qin/A5ODfMa7QdaTihQ9SMx49qqDdJxJDjzPNWV50OOTHaKhFvQceNuyNG5V0aA7469VKVeQzX2x
RGCYe2fX4xi2FmhwnDwd6RUtcLCxGOUERM/8NI4fRror8Ok0ZAbhPZ3X4XTiiSI3kojgBZd1SAtV
w64Uc4MSripMUdHquzMpAaakT9iHnY7Xt6MeIGAWoctwEVaFURfIojF0UIBpgHfVRmPhHArgmAbf
uojxQ+o5zkb+odBomRIUJ3Zw7SCpXS+8GUf4S6SVlBlKL1ZfJqaraoPWTVDNN7uceue95XsHDKBT
0kI0bUjKofOcdw4X9VirRmsUwSWB2Vc6Stjl+NeafiMs6kmrWM3IyBv6R2v1sogi8jrtEcVMBCvG
jDjui8nCAFOw/VFubFczWH8Ou8ioA3KrVR8CPlmB3W06v6AR2Q4kd2c+L60R4mZHKS6YDOJ3qmDe
TvFDJ0A6szxi6DlT6qnxWKPbibwVas4CM9TKGwskznAPYIsD6rrrszrP1KEiszw7TxyN8ZPpQFJw
H5ovABzsWWyFrnjohLsh/T6et871DSQnM+Gn82mR7FHErfPtjeRp2UWrCefSnd2UrghDV0tTpbX1
WxGWLDluQbcpMwHsLPID74oEstH6KjN23svKkGEqHI/ILfPcGmw6LdsQvHFHIp9RKEB6d2E3DkEm
Vk0TuWxgYgbAT6eOtp09CTiEdTLr5KH+f8DJXNIgDrjqpWM0zAfmxEWlCzORs+4BXZRK2GLf+b58
e/22FE9Djtkl2FmowMNfYzjcS166ZCScl/ACIBaGnyGpXyyjF/LC8sNF7cvmj0TseBL2YjGUlbm6
NNswhv6mlMbtnJDpi3XI6xDmUb/wtZSajttpWZydoIj+aWFWW9DlCHv5TXZXt893m1Gh/6qQu0gg
DeL0t7XZ+6HbIM02Fs/7I1n/Jd1+jQbYKp66HmbdOdYacSUZMUfGXSx1/tz52EabcN5Nn5bDIzAM
pKy9ncLfpOrHydHZdLiA2elnDSPUUUi7OoEGWnI4YdQMtw5YaLJEAAqv3iqdE3qA0Yf2JowcTwcP
pbOwGWQaGBxLnQy0oYC8T/zy6y9LBvJiTyTGwt1qyJLF807yompPAUJvZtVgDs5FDGAdmfhTfZXu
rGd72QZEANFL+nbMDK8HbsLfiat/6gsQdkcJUE/Gf9Io3n9S9hd86Aq55EXtmobkurW79mBgRAk2
xm697+4T3XA6VAoSrMI3m3EUUzPH5qEnK1+xC8xRG0trESAs7/HmUZ5rm56jJcQlgD6asL51ehFU
ykhRN4nTYGKUIlsNWScqThZrbI5xhJvGw9dz6cojRHiA/x4n6pgNBGSFumbV5OMMCu7VOqB+WMlM
mkML5wsZYNMgUocQqrdax4XXu93lStfeQ3THOJAFigHl+B4Ct9abk8mPxFWP7h6dyYrqlEraEKIZ
YIhTevnU4pBV+tGTnjFQjUschBLUOgseGHKhjBAUjx2aWlsu0y9krIWg6QWiOzFN5vGdo0nxdAX3
ym34fi5WM0dehUf0x2p8xUpC7uWYVIKVU2FAxrK2V6p2jnOeVDpZ6d39TV9F9h585R+16e2GaxME
RdTVZSlZJ3uuH8b1QSxcqqW0tozQkHef114K0cQ/by6vQH5s/1ldk9WTj/isP/ep6QEsnwuwVUhn
YKjg/SS7J0Hzd13ncVdxRf/e52DJmjzal8zpdB0cI/HeVIULV1IZXqKi6zIDUbivCka7AshXPVE7
wpsLL2aDhiJ4pVI904kZrzFjyZ9oUgEyta23JBc/w1fKz/0Nuor5LbOOD9eNqUvToiAQXT1gHVNb
6NuYHoifmNAxIzlZ87OXtllhc28g8HXJj5tVmGkly8yhBtr5TdZzBaFlSTh08bT7o/y8fFUbWgjs
cSLFaLbftCas3OhpQseEPgUbfPi+sJn/vIjPoo1/03vTSTpSCJIkSXrV+Q7oRgxOU79dzVwGyP1X
/3s+Z48YHffxIRHlVKWIpLDjUYfpXY7E6p818EC0TCoy4W+Z+RPViIYf5Df8owEaYFRS1GokuJAL
k86atI9HlMLEZ2gviI50cjDbDEDLJpwHpVsnc81+/wV5KHQlj1jAHeNisnHKSsuIL3sw5KkQCoYG
RWRb6wgR5ECRvSPsa5NBcy1YDTKYs0ZbQCeE+Zm3fkC9cPcUaZjvF3goum3pUUK9dGr0alXY1/I9
1gsj4y+qe8lyU89ulP5ihyDxJWxF4hp0SDjueGXITwv9GyFdqWO1jX+EMMZu669ldHCBG/kPHTzH
FsE6ATAyC5uavQKN+Ew2ZidD1oYPjjDxFYPX0s70PMfAek7BsXe0Yp6LrgFR/2XDKUD3GHsPS0nc
sxmGf0srLqJ+f7D4YFQmIJ5P4U488BidYo3WwakNrV+cpPbWsN/RtxSTtVphnyU8ZAvVGMiJQsLL
FeKb9kgoHFjr37fTyaabDjZW+yWNFKKe+phIF7nlL0D9EenfDiPlqlvRjiQeKxBz99PVaF1rjXCW
nf4uoZsGZuf0gX1Cgf3acy6/b0u/6izeFnYrx0fKSZc4Y9VILIMJpg5IAvPvA6xLb7oht/xM3owE
wKiHELKOV43hOnw81tSSsqxvQOagQ83esX9/y4bjx5YNEtckM0XjeUJdnKpkZ39T9q6BSoy2wCsu
W8La0PFM5DhiwqCE9qsfrFhsa/fpryMSikzQ3RGe9vznig/2pZNE8gYj8CD7Tx/oDNvZ/9yeMwFn
NphHexPaUejGfwFU226nFTYYkqMjAqpcMTeVWNW23q+WfbvYVYxGRGqAy0psOhAJMIg+v4tTAJnp
9HI7i+raMH36EgxcNB4KAt6gOOcY9mFTtsYQODHG5X65Ekkc9ypuFvGTavCtLOi3lVWYAxzJPa7p
3edZ+FF+6cX/+j407b74XCRTr29o55U9xKT8hh3FwwiWZNtr/HBUdwDr/EKvXFpMX8Ec/jBQ8GRX
VeEblFJBnsh+PVsB//2aQUS4A6ZXpV6ARg9pNQgLbZxCaMVXbbvwoNGW5myrrm0IZn/qmyPVpeXb
6LvBj+DVJol7XWCZrZ9Dm5JZSZ0dy18Pu6Aj1HCx6VqoWAHcoIGB5iV1f6vY3jiQlvzml30hTHak
3uBvFAjf9GcrRGJdtoBcWTZyrWrLTk/F5Yhp6EuQluasCwj0eRntdGqtLuT4m9c276hmTFwFCKlg
iu+cphp56L4TW+2D3qRITSRQA7pDL2m3Tc4raNIDSQtUPAUzbgsZaeiVTPa3IhMqkE17J8uzyKNK
DjHg/p5xUDHbRHRwG8RpZgUH0+rM6zuRukWKI7rFoY+04VHamhIJI9DKDRqvvEjD1wJcNb/958Cy
8+zw1OAFw9CUfk1axvdt9oGfcapto6RTcJfhJh8Zr8pDEu16R8o2NlfjVKBsXwEcyDbRzdabbRsN
w8eNJgqS1XS2oIExrAR620tksvqcCWssralAQg4lhOBKtkJtkItMJJbsNvKY1Psot0GrvOHfDfMb
9LC2rFIAqLq8cmMwYT/hG+ns5Mkhcm5jpr5bs5Jp9CM+VoNQfrSLl1AeqeAKKDnTPSHhVj3rBoMO
4rDwwr9G/1+kRieGlnipbwCJyTOFZWxqqqriioz2hqdg33xVcvyYxn3d6bGEB87lv6Popkns8Zdw
B8PA7hvpiGzwdy85278JTWzqet0aw93Ab4XEynAcuM+EDy4JLwv/quRDaJZYYN6J6R9PdILVHPUH
P1r8fCrieeyvPksuFIAy0z2o4twyoRKemaOraSODdTnPjtwBh7xrtfIw9/jsOl14r1CbxRqedv7o
/3bPFIGEjTTFeq7lW5xdbLAaOfjCdcjpf9BUnnZv4qF83bLGR16ZAFVvDEFQtohWvGkC64fgrnw1
PpvtR4jm9sUBO0/vHkP8HgKax9hWawqXmGpNtEjxmhYOUiV4xGPwz2YKMbuUuok2iwWC0QzErwcJ
3Ev+1k4LJBndVOtxBrNOjjEefdfqT5lpHfzmDlk2sqdADZdCZx2658JwY6DCNBjGD8bX6/Wk5+UE
LSQW7DJoB04s15qx3fXXon5qRhiusTM/XDqqlC79b/xsIMTjB3XW5ezpGl7p0JI7p5kPatWDldUI
LPguuxP8h3Q5eGU19lYgyosIAaLD20t2UtBgs2N0zyS1doWU7LVLPucwYxSSr7fTTeKVZ9WK45ah
vgnIG1Gk1KT3SwawdMPH2XIYSI8JXfFlA5dLOt1dJMFy0sNPnfNzgDXDTAdW2oRCXKaI0bhEj4CW
WItUi/wgNLm4FZlHqYY+yHlem3sCzqa/qPvyc5CW7nbQbq0FBiOZRNKP0OkmBF5iJxkCnWItakKP
yjXEzQeefH9ps69FaHLM1jVqKbioLuLMg/8X94PXW16KnUe6D1mAGPKROqZ0/T8YrmOeBGqll7Zx
dsbux5E1Mwh8iltxIl/B416vqCRH+127FAJRMEMyRm46QyIy+SxvwV5yx9mGVsgrpFgf1RHEQ/4B
ktlZAI1dU1ZEAr74VIwuiI/BFnnHrc9bqPNytLpkdkkrz+8D1b9BfQLEBpvAmyvsV5L+S+gZ5yje
uHWkJDji30jLX3za5l8eGp6tYra6c6x7MEqS/mp2/A2xGIJ1pJY4kBmv0bvBcMObGBaBJdKjjwhc
t1iVuQxxr6Z0RVh2lm+p9OR4Zxvx1/MxzwUBfxEkAxDsXwCLehBlK6RtcJz33Tk81cp1by8T8zz/
k5Fv7ThYjAjS1srZHiRTjk15gXMJ7oGQCYEfNtnkusNejM7PCTdJiAKvR+fco0VH4TM0rR3Y9Bz1
PdMXxyKgvnY2735TZwRmk6hFQBsrhaMFoTi2EkwXKiqeo641QhcVXsSpWhOzCdVKbmYgx9C+I3Jw
r2BMP6uqXZcg5Fts3ck+vswU7UloittoSlOafGIDG3AZ5y9YcUUO1r2y+vuKu6jMFn+8NmVG+HGm
at+aJtYzBUSE9IlJ8Kaq0uA5RmH7PHP+CV6Em4vRmKIGKq6ljCDabfFgOl4ss+UDy+gBGop1vf7V
QdJIbKi6Sk7KqBJK4pna266lTc0o6EUBF4BTMbc/IlRF+47qgDnDmwBkS5MKNk286Cww7X1q6tw9
Zkgo57mJO0IxDX4ha5rXe2TdEbFcR9irAyVj/cGiDNG70u9rHNxrAkRQJmNvIgKXEx8GXFpDUnpq
bdmndHFOJYgSvCSDbKRWmxX4iJl6XNQxzNpajPYOu0mEJZSfCdM4YiVz4NtrEFeGTjggRG2s3Umb
LcAWh70ZF5tniRroERXov4R0w7pk9uQ0KHor0rVlmyp+Ck4WA5KjcPp3zAl42Xa/dWYBSY/fSe5N
LFY8te0tfnpJuHhcGusKHgNHjOsb30XAjzVLdJDrkaeYeCiE7mbftDph+jgtTesh5s2oFBuonUYr
ynhkj9HZ5cVZ2dF7CiMoY25UbNV2qFDWXWdKkUvqChpj2A+y4RITPIkILXxDyGa9l7bwPAJ1avuS
C9GldgCUTxyVN337Z107XI6IMFXDjwpiltcAtITMrfgQCmEwpzkkLvFUCXgmdASqILwPjAQ34GMW
ATiMxyGdM0/PD6gBXHqNukdg2QcHLIdUMfsJOAsV7JwcT2VV1abTJLYWXAEjwtu6N5CzsogbWjd9
tDODHpV6wmDy5vymRFmMVJYppVCYP8nF0zbpEgk0CMnmmMUSUjNwpEIfvyBZOb6MWDPrxDatcPR2
VsG+DjSr4KUdxHeaYMzECb0YAi2Tz1kM8ea+wxFDwlimF2aikmEb8Tg82HPjXKMfDfrNlHwnhJ1s
9QUwHiO/mEvaF6F1c1AYnVHRpUR4k2j42JGNQr1XyNEkRWaAEJQrh5gFI7Rq7RKQLzlTwZjqFU4o
Eti4dvYxtKTMGz6xVJ+Fc8j/MxuufN/DfEH9SxcLecn1PYLTCti/uYTOCsjpGqeZQnVbkPyjOtsm
VlLI2U472CtWv8KTppH68y8dmFTVlwavOWclBvpX29v9wuR/8X7t0Yxtcti8WmhubmAgJpyj8nTM
0HateDwD8AFnZBnuZ0y1O/c1ALGyY6O8AtieIEjxzzWwg6uguaTwUSlE/j8MVWV2Cj+oV0yk+6lQ
y7qkJsrzXHENhXSxZNkH7a1rVBMc9QRbwr8P7/xGiVPKctnTObbiRTPxwP94MdwJrN+yLdy8fGDI
SXWwYdPzLGOMDZoDaQgQAu9EBlGNCYQlUwwF17kGJCwqcifu6im0R6Ko0K5mQtTMScfCNFBCKWeJ
4uS4qmtzQURSo8o3pTBUinnQmJ5cwwOzjGT5Ks12twRLjeQXXIEKxOoBD7SQZ1TGj5rYQzRhlNzR
uzgrjcR/bQmpXGZZmK0FYYXhyG0oO5IUfzhvNeUAAfGAzyjSj65oluXrw+uHIE6b8T+9c36Jj0kT
8v6LGxNiNkxJ+t8eQs1HLq5mxW5dHc+GDZeA5HtYRmIu16u9uIz4CE/gWohlHIwW+8khkOjBpPH2
DEZVmRvacAwJDPTeC0OPRJ1hLTxpBI2kNyQm4N5rzG2v3rNPJZOVFBbQRwh9hdwDTPEAQRHidH+w
AiZI0FPec2MoflrU4OtlGUJ4Uss+QGeHfB9hVO0qyyEDWvseawVuqXMMXpj8Famox8s3wchfFvEU
T8NvCAGFi6XGCLIndFYaDOOcjrGT1T391opActI9CcfjCB77wAf/zWPX+FyFn1pXmQZWgGu6DLFO
rEHvx2jHurZrDO71YJVoo28g9VGaE9PHmJvZKxk5SLOXxXsXXkNkgnksq+rv8igMownhMd8MMufV
L1D390lleIrHYe3p1R8nr1QpsyXaYrx3vuXMfxnqmGuWRzbhiU7NeOsu2T3q6JJNQcySaG2POnDZ
8je3EXBE84upBoOHT3rUFRc+b0WGIKvOv5QMtLolfB4e2JWLlmVJprfBym8eIe5A83BVjMxjlUB8
aGSmzlkmp6OcLChWUsrEb5imdJcVK9ho9grsLLZ2wO8QQejmaD97ech1PZ8/f0INTwIkBwqnTxZX
KCtU8hzIPRKsK1nm4fUjHlCIA1KPC3A7d+F0BgzaE5tRJ2pdsD6LoaYtxm4zFOIFkM7yBALnpsVw
2c2SwOLzbRHztjciB65+yU1pjxgOaULIq+aOLmQTAeAiIv6vP/q1EvnWS5ZvcxeAWksDiIKTPX5B
3Vk09JLrzr0b0wJVdG3OtReColOTsLOIq6cIGObDwCGyUdy5l+x/GIRvwSkRL25MiaeWIGw1d8lk
F8yYd3Pkcdqq6qpP5PHfwwhNwiy7699XTl/6rT7jMIShVavC75TP+v9XrCCisduiNe4lF5GPK+wo
0AYhzil+Af2e8ScKOF3oeAXJBMonff4RvzxVV96EsTRra3hbcdtw3yiH+gm3q+pBxIn35Xy8dKMy
JoKTSS3drxPT0zQ1yt6RbMc44IQw3QrTqqxuNERPKG9omN+rM4f56LwrGBnrNzZZOWJ2MuUqXsXT
JT59/mjw0AadKTZel/6cT8iVALYW85Qk3SSOJ9D/tD146f8EfCcZT3Nvb0kevBTWip7F6bEYBhNU
9TudiwblF14JFLb9Fi0ntMCuF/YgIp8kZzZn7i6w90W8o2BjDV63+qVzz/gKzevMJmPGSdiugLiO
BEkOnvZxhrvBXWEoHpRuvFtVLJy4beDTkPJ7W48W+IpSzdYxrBVzhOf8VIzBg+mfziIbthfTT/bY
93fz88QRlUR1Qn3Xv6OxQRg/aYPiSJYeYDsKdy1qZhYaOvoN4rBlfp9bcCZa9N/ohEPX9yAriuwB
RrTpkwO0v1bGyMUuk7TprY5dKGjDBuAwFEDMgRuCCsYdqKlZinY1Ay7c7eL3Q+MsLrRQpB8wAIzm
5E0EREW4jyxdYsHF7XhlEbUo0PS8wGFkTvC4erQIuDw6Hq2Pyxr5bGb199Gnr6JdC3ztFVL+8XQr
9O9PHFZpfxzVTqUTBPPWSd6TE2G1UEI7DkQLSZQWvbT9FuwGyryf8ptE90ilvOpKD6hAfvIT7oAc
tAP23GOoCCyzwI70VIuySmq6xBWieBPQU09FTR1hLnSQs8aZY/D5C7yujR1bJWN/c/L2tvuc2zOY
ZBgTb1e9JIxZXIDQAX/8KJ7Kf29X7etFkXZ3/oRLjX3BDTUEbniDzWmuKMpItlNenTxAsg8RvqYq
7/fW0OR++8fjxXQojpqrhi0Ce9IVlotPQdPTapuff/PO+xamdfGlDqpXaI6M5cp+zDZl3ZSTffMx
QBCgqyGLmQ8YJixR5O1PbKuWUiq1d+l3Y4BgkV9UkeMaS2S78aLSBrfrfLtRyM8bAxTRWxaYO5iY
1MjJ4tA3S65Hs4LUK7jkpjlaTqISZRA+qpk1ucXyVHmRM8PjfWSqcXn9gD9Gk3H6uoXQWCEjUw5i
XBT6WWv31sKH/YmdrEqV8wF0b7RkHTAjJPh3VWHMt8Cry9A2vYYkEsV6C0830xsCesAbQkvI94MC
a7XgMV7/K8Hab/TRrcQhsDOzOoMnFyRPugn6Ngn3wP9LHLjqnK0/Ujs7jZedgvc0GIs6rfQyDG1+
cUYNidgEq3SBQeVL11XiD53utB0B+JFwrcZx61jBDcEngTj1q70yQ/dPsvs6rijhfHOnZK98W4eH
nYlLOck0Tuk4umShRjwR0YoqMzryQh1DqNNaoDGKeOVPMGUJjcs4Y7DfRqW1jlXugwAZqL6wKOyh
noM7V9AI4sAQl0DktpCi9H+R25FdNaMp1JuDVngTjDIuTBn9hoxmo3VuwgM9AzgGiD2T9MRqeD01
/XGm8PXgbOy1pLTv2VS6D8OksuscfZaICUxTaINyD41AvGOMxyPaJNTQFEZQEfv6ttUTPKEFBe63
Lnv2oBbAlpx3IHAdmQ5sZytdp2z73pup44HtGcDly1FcFvkKi3HMomo7XwJVgYTzTNutoUQjaIbj
kbIzDeEOQ/WX0m6dcgqQLs1kmHApNTwQKJrzlsnPD2NEHBtUvg0jjBTQNWJ8KqA9APUZ7Gd+UbHr
8I2HO0Fn7/w0ohPaCfIUar/tMa9w09AR6BoXtAFv2tr7Ij6IShgZYJ79pMgsuIiD/W66B4wFBvJf
7eukj8ZJp5DwqRceudgeS1jDX7fETppv7E3aSENFaBv/dZBaNErlBi/yFdwzIHKrcS1ScU27iVz+
WcbtJry+QJTz5vQZkis7d6FatMoh4OhkXwct0nlq3MVV1nv970crLcFku1tgpHMZwCbsoLUNnzob
Rt72FC11urwtgFdxH4sF7LJHqpBZ1g/+Zgf8aRTmuAms0FHlzj2je4KZ/alLKBJDH56vd4IWwXli
GKm8LFCORQ99kewqS8IvHc/34ADaOnvlj1bQy52qv1q1TXK8/KaRIyKnGWXGlwfykAXXo5E3PAgV
kGrU+p6CEUdhVVMyedTRRr8A/pk5SIfY4Iie5gzdUjT5QlEnE8IoVdFOIB0fkeC3VLf5xXf2lEqb
wn0fE/PmmaxExUkd4B+dce1XXwCmbFTzZhC7xP56TfxQ7ztIp605DV8mcTk5ak15D+H4JZwGbi2Z
pdEFYKZrqCjTAh+7R/YlYssSmRQiqoYYtBaLNNcn5oTnVO9HWP4olRcqlL9qmYhMW8g9xz6LotMw
h0c9h3SauaC88AvY77At1xQVqm/c1HN0znRuqDKtMNyLE5zz7dD+F6KAryo64WXv7nFmZ5UJl9Pg
VcB4rWsXy2DZTIdjrQWKfFsAlexAHqcI812QIamg49815Qjc9tFIPzoSC51ATVHCcR73bEYeDShV
0SHPpErAb1BDgvyYO/gZUCxAjlU5Xw7Q8/yxPUx+oteYp72biPHoRR7URDfvKH5GRKQnUb4i9Vrg
jyjet7Zy/ggfPkSRgXY04zck0SCEElD3XSJRH/Ktb+vJtQt8gtNd5R4QXYkWCh06jvGaBv6Ha1Cb
f1YcWdPKvHZitwELP4fpSQ7Jm1ILEyTRLaZXrtZ3wqr4hfG5PaHBfuXwFJuRPmdgk17xOlGw7ut3
LjN+1+IcI5OV0G+tinvO4NYem3MTqVAB5ba8pLJqKrmUcVQctnrS0COmlFx1joU8+PFZLELdzakP
SE4p9Pe9lkkidbSixPtGenp61do6Kh38h5Q2+G/+pjrNYlMLJ6+dps8oIuUm3Xqyq2BPoVGWoRx7
gwB8zW4C4q2Fl/DbVHnd2HY15IQvB0Uw1MBuxFy8Nj7pxVn1pG8X+juEPLplouL8VK/hni394ggz
72DUc6/eDmBksWiCRwQEtzJh8xVsJLJWDVuDjRPigs9TBghlCTu7+yxTSmh2OsMuOALY93Xvi0zG
iPWlfHHBjwb3Z8BBjRYiOWIZtRhTcXhhq1NuKcvQ0SK4uNdcXv0BH/SqKZG4voMdl04t9TiS8uzq
l9so1xkMZqXokecvL5JE2h7JmlLVyA9pFy3GrfnFm9plIznh6sLThVdb9YY0pw4zQN6BylbPZLZ0
PPsM3M96Y7e9XnYNj2Ujq1sr/mi1aOCV1F4ZiXnsyghvIGdOd28XiUlVEJawCVSdbJcqYUSOz8XZ
Edui0Z/Q0EEYWqlqDO0pk4jQdUI7CeWneA6ppRaD+A7CpsGWEyuPV++p4asz1oRaWe+JDtY5FIRG
QTeLsm5uDRYafcNRfiqiju9q5ncSAk0n14p7KMTpaazJLTSa4Zot0efanKUGrKhggphR6W/yKALT
Wl40c+fnMBe7lednFCntFAlAlg9BSQ08rcKFLdwGnEfStvpnFpdDPiZmkRVMcUC9WUdvc6C2wam5
/YE1ReBUJTCrsT+sq+sZGj4QOyPcncJMQmgvra/fSnL4mcx0qsofCfNmczhKy5oDfHEQP0BAv3lh
0tpHbsaqfBwvg/soZOzvDcWSUqGfJ/dPyN0gm8kaMZzETmAVrHZwzIyWXRz1sOWN4ULs9Hw1FqFv
scmgnyCu3eu3Nh4RYr8cPEnf3nJtONv1TsffFFiewyZL3yw0M2HOiQcQnF2X3FoqKP0oqrmjg6Ai
+HFmkvpfafEqwqSC/4HYrLbvvORYro0arcrYy5oC6cZfSdhPoWumIQJcASZzdlw7gLCuD37GDAU9
HsKqCoGFX5qUQq5T7zSaAEadzUHbeH+u/ItnDx85AvfWHjvvA+MDnDuh4T7vXMNtcPcR7QqLjYbb
9v5bQBucTq3UYavPAocfT55NLwItrrbhyAsO+SsgO3yYmjIOSXmThj2NA8JnOUsGfTbst9RD09HH
NYlIYgBsjoWE7YuRc/v/hG/UBiRo+sDdq/WkCHOmJ8aR0uGy6JuhURAiNXGdWu+wxtokquT9ufLf
ymRFYBNG3Ua2H6X71rJFxk5t0AzIuZ448R5b5nDIngAOf+VfRxvnmY9wE+z0ezvmEeMKVjwDWCQO
cIybjbRD3Uf55o4UaAaB2pFIil493Ds+mmKp9g832IT9SdVf6WNj36oxrsj6wBWLE6ZKXAJwSn9v
c1AaoaDFPcqfvU0b5bW3XBNss2kXxlynHvL80sq7lqVyRvzmn1KG8cE/JcTRv1bUntueLcqF92gD
NWAjQpXhkO/UH2SuzohTmri01EaLnjir6tSr6lDynzQP4umlJMcC0Ev+Dp7k+QCo38MFj1VbUKbx
1SinxGLTNwaImQ==
`protect end_protected
