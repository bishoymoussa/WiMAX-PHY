��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$Rx�y�<��wA�*;�x���@�̦�W�X�fa�M-$u����n~�%���P�$��W��kYَ���P7�?UMfT��q�6�U��k�>����~�\N�(�����X�e���/6U|)�X2pF�]$h���d.���9E��WG��L�X"]�Ad����ľS���8od����e�GT?y	7�������ݵ�^��R�q^]�鍦�����s�ae���h��L��P_���ާ��YЭF���'\��68�b�[����w8�[X��V�F�0͘3����q諵�uW� �h�u\V�?@��_6G�_�*�G���B�絉�f������[�G��U&�����~�F��AׯK1�`c��[<��FY���4I� �#�G��x[X�=�Q1��`��R>(�w����R�O�?����7�,(�H\�#h(W�EH=�������yq��Ѿ��aF����:�U~m<|��.��0=�P/���4ǆ���T(����q�v���I�ɿ����Q�,q�&t�Xy�/t<R������^�� ni�ś�;H��*R$��Sp.��54m�끸<����6�� /lb�:een�,��Y����������S<W������E�L�K
�^GS����>�u�!}?�m���ﶛ��.�+r���q�gf=h�ٕ���w���r���H���u���~��!p�΁���`�K�,�>���\�A6�B7�0�1[�?N�V���Ń"�Z<^��({%��?�Xg<�-�CqL�[�!�ҌX��
�77!=-�B�jL��f�w��o�Q䊡"�����7Z=+� �&',v�恿,��+�
e(�n���	>�smnHCm��(3���wԷP�[���'�~+td�����wԡF����Y�dw�ܗWZ���L����"jӄ��_2�������ɣ��F6�8�V��s�,H�]�pK+b�g��DR��2���jNG����,i���m���d��r�"0�;Z.���cx7����y������K��Z�/~ޱ��1��p+H}���vY��^��9l����t"�%�|����$ɱ�i��m���x*�?�I޳�\d��Ϙ���I(��˟X����0�����8%�����oa�ϴ 1w�H ?wΉ
���������JA/�������v`V����J�s<N瑺�n�����-�3�Z�wgp���n(����N{�Het%�]�,����[�a�����xoQ��}�� S�%3�}\�����x�-JA$�{f��/����F�jf��v��ƶ����S]Q���{>�ǟ�3��%T�6��BxKK���p��Ϫ�b��>0�0A=W����;x����R_�n�_/�$y�kwÞ��3���P.}��&@��:P���:�;܈��������9|:��v�\Q
(��t��g�Q*��h�n��G�MvZ������&)<#�p+���^X��'��dp��<��0?�,K�c�E~�?��!��\LWå_]�8a%-)�~Us��a��������@Wp��Վ�L��Twrо_����SK��)�Fh����"@�-�uW�D�d�J1�{��	��9r�%�lo� WK�R��o��y�!���sQ��1r�����],�N�l��2.@�N�N!�}E������k��N�UL�n~ө$#d�����|��d��!*�[�e�������
|���ؤ��5�Ȥ�h�^���T�(Q�(��U=e y	N�ֱ�Q7}��\c�� ϭ}s܊����W��[.:���&,�;��cil��WO7�J�?���+����?��x�q���_����`����;�7�8+9�>�v-����[���I�>�Gd|�>{�T	=ib> ����>3d�Ij[���R<���]��3�0�n�ݚ\s�Q6H��oۻ���TÃ����)4��dlch�o��4j������U�%�4L�������;z&�Q:�7�Ms����;<%Zwf[�1H��'���9�6�m�h�З�gO5�"s��N�y�'�N~������O΁���^�?	|O+��<NoY�a��o�<C������5w/EL�м�{#-g 5�B�y�S�a��o��)m��$"���f�/*^�(�/2Rь��KA�Y|�:<9�	��j9jC��,�M���^��q����>���v�K�wtZҰ|]v��V�æe�R'�:��^�C�*�k���K[h�����[�H��$
��j�l�ԕ���;6Ϥ�
]�7|��#�:h�_'�v�V,��&[MC f�jD<�������I��,N2�S<�'�9K�譗����V�|R�;�;b`�WJ���%7�Z��8�ʍw?�m�?o1Y�VPA����%�]����n��2����,�U#n�;�Etsd��X���ᵗ��c_����#
Fs�{�X�bֵ'��-��*�E�kz ��|fR
�X8�ʗ�C�T@�������ɤF�nl�) ^�g���x�K�I���	�0��,���T�Naѻ�n�KpM1hp@���(C�����w��W�x����UP+)����j��0�i��AL>���*�)0!1
F�<_tO`��҄k�	���;�������H	�QڪN���0讒#Gp��ń=j��,_Ȝ4
�9����h'Wr/O�Z$���޵�g�5��AkM|����Jaw�:Vi 2YȆ�O�� \ύ��lo!|-8.L��^�C��\��"xyAT��
>�}�,M�����Vr�S6�㽪�ׂ�C��:��w�QQFВ��>�{WmO��.ϙ��n�d��Fͧ%�NZ��'A���C=�
R[�Yط~�F�� ���# �N�%��!n���u�Z� �!i�&3�&#i6f���#^����o3Ml�T��{=��lk���6�D�������T�&�d\�T(Ƒ<�u�(ݍ�����6E��g��)����e����3V���Q�4�>�xb3+T	�'�p��nH�}���e�Y����7:۹v'�]�P�{%���h�;���0�i:�:�����b-5���9���P�R^TҲR�a_gN� G���:Xާ����ݺ��1�/w,x�qT>  V���B|&{C1c y��<�cA����6�=,jm�<�33mB�м$�d������p��hZ#BMQ�垨�霊��g@b�_��j�e��A�d�C���*�u),K�:p��@70�A=��@Tn���*6�t��ƚ�cz$囱#� 90��Vh�3�8�
{?��"�R�
�j~��!��]@VyF��y`����{.���(�>�����e5x���h�X\<��R0�Y3��@�,���B%-���>������ Z��D�)�lDe��ێ�Y�A�6p�)�̊���#Vo!�pD���v_�a�x��� �c���]��^�m.p�q8c%�����w���_���ǖùa�97tk3���G����,���M_]�	S�#��E����z�P4ӓrH#Z=������N�yh�.�̍��68)��rKJ���優L��N�`�^]�G��	�ϊ�m�V��C��l�1j����df�X���[����-��h�z'f�R�̸�(mSym���b9�Ђ+(�\��J����:K�	����?&\}:ñ7�8�qy韖��!c������-~q����ȯe���E?���J=wr_�
�I1gE�u��aC�Ϸ�9�	��1��+ҥ#V�@�2-T���"�Տ�Ӊ�"K��f��F6ֲ��	�d�fk��*��(�<S(X觻���-��D���r6�x�8{~~q��B:�_������9ҠmZ��6peh���]V�D=�!IUOY����M�IQ��k�E�z�O�Po��9�b�	���(9o���P㘐�K�<���J_��X[���&Cы�Z��2�AҲx3�~ 4KD�#v�&\�	��UP��2��6��C��ߎ��a��F��VY�\;��ߨq�h�'��cKT����N2\�3���z�S���B�嫲�-1� �����M��9G�봴vzw��Ճ=Cg�	�&$��o����L#�P�����̟�o]��W�Ps����w���ǲ(jG%uj��h����8�]~�� �gbK�E�g2ܘ�,��!�#tEtq����9x4�UA4��"J?�9WX�s&�[hω��"����F���� ���;���ꗨ�>fޓ+ǖ����H	~4�U]Qz�ُ%�8KoiM�����$vI�^�K���q<����Q�y�9��*n��n�SQvQ��G��̃e�m�k%�M���B�Bn�o�Ǿ�B�5	^W�����Z�͜jK{rjۣ��M��=M{�ۙ�_�,�Jy��7%H����Lz�!�#Kp�X����m+��j�D���2�/%3�~ ���g�h?O�߀���`)Aw/4-�
�tSV��@��Ǧ��Jz֘nF��FH �5 ��-�nQ8*-�ҡ�3!�S�����J̠R�
�>�|�i�frA5��ְ�����)1MШqC��t_���&���|� u�#�Bu���,�B�\���<T��@������,U�� Ql��2I.�uh�.yAr��O�#�t��^���h:<qdhо�]�v���=�?��Ĉk��Ҕ暻{څ��9�����@�����M����P�"-�a�i����1Tr����3V��H���9!��w��pD+��H��l�i�����'�<S�`_�+�*y�s�!Imˈ�KU�A�
 \�jQ��9�����%��n�U�:C��Na[P}-���.���PN~n��Fw����V��� �-ocK�x�0u���[&��r���1L�k���2���̼�g\\�w����j"�����1xEH�9�z&�M��b<?<�27���FHT�j��	�^�R�ߠ��;n/S�j��1d�Ds�m��l ��c˹X.�"���/���ň�s���՜�0%5g*�+�*�KX2
�2J�\,��%�і&���#�$��^�4�4��GW|�1��Uku�3�B�붕� �?�?�*�5;�T�D�c>fz[�������G�r8��������;���`v�,+�h��Q`��݌��������A��	-��M�%v3
.�����"%�ߛ�K%�c���DU�\h��S��ammgG��`L��rziL@�AxQ�:҆ʩ�ܴ *h��=�3�+��K��C�yUkPB���*O4��89X`��[�B���®#@��O ;*�D������.�VӔ΅@B�Q{��pj��y��4xB_)A���Rp ��P��eH�+�`�6��� �̠"��Fg'�܇ʹ����Y�`Q+�\��@�'M
yg�޴�����S0�W�O�#n{���e�5�%+�g���I��f"ws��v������I�T�Wl���{��������~�����ɒP�RUzh}�[GܐW�nf�����@���F�w��Oȉ�����h��N��2����������L��ja�,)/ =�}���g6�uե��7�tl���!�;g�����n�!=�R�T��E���K�A�-�	�Tf�����n�