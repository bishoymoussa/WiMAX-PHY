��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$Rx�y�<��wA�*;�x���@�̦�W�X�fa�M-$u����n~�%���P�$��W��kYَ���P7�?UMfT��q�6�U��k�>����~�\N�(�����X�e���/6U|)�X2pF�]$h���d.���9E��WG��L�X"]�Ad����ľS���8od����e�GT?y	7�������ݵ�^��R�q^]�鍦�����s�ae���h��L��P_���ާ��YЭF���'\��68�b�[����w8�[X��V�F�0͘3����q諵�uW� �h�u\V�?@��_6G�_�*�G���B�絉�f������[�G��U&�����~�F��AׯK1�`c��[<��FY���4I� �#�G��x[X�=�Q1��`��R>(�w����R�O�?����7�,(�H\�#h(W�EH=�������yq��Ѿ��aF����:�U~m<|��.��0=�P/���4ǆ���T(����!Z?^M,!��F&ea�[@lb�BY�H}X%�/��7���Z�B�y6��z�O����A�W�U��C�ݨ�<����s-ur_������u��E����ߕ�ͺ¸�K����lq}���?-��K���h5eP}���~���d�۷J�o�-��#�p��NH��0��9M�]�F|&��R��˹(���Ud��%jj���v��I�{��n�J@Zi��&S�!��2z]�G_����y����*�v���
hI`2z����В ���T8\��4��(�����Em�JM��I��.�D9m^��V�2�W[h}1���LJh�jޤ�<�w(2��a��/ �nG"��	]:^�%*��ʲ��V�}���Q����A.H#�����L�|�Ƴ�V��[׊/cS��f�?>N�S�{��h�剹
�UY �^&���asR�;�l��'�V��x�f��4���f��!#|N��N�sGtB��V��lJʠ�kWI��*}�:��|�Wrl?�RZ#unReO"`�-b��t�D$S��و_K%�M�u,�w00�#�+bfg�xL��c�n,=��_Xq��dE1���N*�mn^`ᑞ���m�y����ј�ChD���[��M���%�IX�]p�CC�X:����a�y�6쫇,������������H{���JA�"�x)����o��� c�.+Bѩ!�n}��ػNã�9! Ϛ�el��-����&�7�C��vVZ��bfc!��DӃ�m_:-ʡɊ�kV��Wq`b��Ar�@����ަ� ��݆rF��m�d�L��� N܇�JL�!�9�����1�`�o�\+յ��D־��|�DI�W�*~�0.��<ƠFB�c�s�f���ܩ��?��>a�-4SU:�{k�7�ğӯ�qQz�ԛF�������5��1J��@�G3P�&0��f� _���L�h�9h0
y�����H_����\1�@�Q���p]����?Z�Hlu�dy��zl�#0��p��3;M�vhkP�IR�L���{t��J"Ov6��@��M�!�.E%��;���Ed8۪��C�Z�	h٭��oz��=�9?�m�*�?�����z-�l"�{u��4^ɬ8_q�o9�W���-�M6�Ƿ�P:��-�T٥�a��b�q�>�;�rn/��s���J�0�m����!�R�>�F������i�D���$6e=j��(�Y�sgYҾn\S�"c{'O�����P������w���:�Q3o�Y�AL��ꪒ0�U�	3h����NH���E ux2}���'������w����;�4])�8_�o���PY��[hK�f?�.�x7�@�Q��m(Z��tyߢ5�ܨ����-h~S��ѢY�Tl;ظg����/Եe
�KA�5O���~7��u���2M>#�J�N�4���8�<��N>A��gzg�"�e\��e�~\U	b> �pi�H�Ho"�},g�]:�*�=
i5�f�B�׻�8�)n��)�oV$�ovibN})2SI��'����;ȷ7��fF��h\��N
����V%$"Q$��nɟ���
p]QuVb+C���gi��$&���.9wr�{��<i�y?`k���3��c���d	%\��TS���&!��S�B����N�fi|��ȏ@�U&��2(բ�Ʊ$ ]�x���U�.C���y������U�D�����N$��Ma���%h{�^knv������$[z���8I���x�DMaQ�L����4���ڬ���?�T�O���ڐE�4�.])�;(��5�y'��:��W�@+m������uf�|y�( L��qX1[�I��e�;����e�.T~�^ھ�@�f����9;j S�g�)�r�w�33�:��@�7��]����@a˷(2Xy�W�z���x�ǵ�k6�g�o*�&I5�(�XFX7">�৅�.��������S_Y�ௌ%7��A[���rOj�o�'��߹�C��PH�5��I�[������v��hK��ϫo ���7��b�m�/ZF�wR�kZ�izRG���j4�i_��r��*�+� �c1.����H:\��[�,Gp�t�Te�w��VzG.�?�ib�
I��g���hq	���q��LZL��m�1�|�nݸK�H=��]�H'����I@/��~AXԵ�W��('�x�V,��ȳ�gP��=�sU��{�5���}�%��Oٞ����#'Ĵ��'M��1XQ׊4M%^w�"W�۠�1XO)-�v`,|�o���?A?�t���@�y��!�ѐ�=
).�F�z:�L�$����H2�ŨD��H�Ĉ���j��u��4���%0���8a�Ś0z�i�J�Fa�}�]��H>�Aen)�.�>��v�a�s�!zF��z4�P�"�^��(���etx_.��V3��R�Ac�D���Z�e�)5jEi띮�m��c�m����z�$=�q�w̓����g7���)KD�ʯV�$	�rX��2�l�l�Y�>@iЧ$t�%���XLдVt��>��suc5�ʼ��#c��"�}'1�����}Ox�z�Ӫ��
�p,��[�
E-�h�+���Q���f���q�B����f�%О��w�� �l9�9$������4Ê2:G���IMb�L��T��� �����x�f1^�e���r��-�.,N����B���Ӓ��?�`���V��݋[MXѵ�q`���~`��w�Ⴡ��P�0�S��l7J�(F�E�u��#��v���V
:I�EA}�����:���u���FtQ��D~�����vOC4Z����E"�l!I�H��R�^ٿ��"NA����;}F�W��-Zj�4�f��T
���r��(����/��ߓP����a;_��@���v^�i�-��������t���(:̜ _�:2���/��"̵����W���R��W;8��,�3�+��ş��,SK~d�x��0�j��5�')I����� �mYݘ]���Ez���́��A���2Z~�>C���K�d�I��l�'DZ)+�D�eݣ��ёlB�I=�U�/Ly���֌�Ϋ�2�I^3vP���u����>�w0��)�ǽf�C��#�Į�[&1���\|����E��F@NK⊴C}~`���%�n�/Y~��G*t�}{��r�jϏ��&���`@��<�p[�;/F��k+���e�W�{U��
��,GF8��d�>�6����~��J�aq؈2��צ��z0[��Q�/�_��ұ���k'?�P�+��i���*�b�۞+���zݷ�F�b���̲M(U��\���E1dG*[@̾�E�L��_{��t]][�^�t,(兺�4#B�J�� /�(&q,Q�~��DB=[�~I2�>�+�Z���
Ŗ����
`k���5k�R��0��G� 9+-}τ�W-�U1�a�y��,W(��'��'�^8Z���{"z����D�']Mn-
����lp
��Y��[`z��u�,��ʩӃ4+���o�ȉ�8R1�IB��&����>��߽z����k��{��A:�<���66X��"��7�E�]���3���K���HAY�Mt�F��n�¡A�5�y�c�}n����oO!�Z�V�7�9�,��� l��3���F(gu�a�X)����zY���h`�w.�aF{�t���k������M���rJ]Dz���-�a�h*c��V�c��Rde/#%�Bx�0���:
&��[}�o�u�4������׈M�aӅL�o�v1@��oު��Y�X����54��2j3��D\���Ep��ɑ�|��I�jt���ǁȇڪ���IR��������c�}���0R;ӷjnŹ+�Mvu���"��"� �9�j����)�ƿ�X�}>۫6�$�+�����f��~b�R�l+г��˶"�Z�|Ǽt[�b|ʬd�Qq��e?}�V��_-���W���p�D�y���
�O�.�ƨ�V�+��?����vl�LB���@k�~��H�t_�R�=����/�gSi�:ְ�L�J �#���r�}����D��L�Q7/w�Y�]�1ν���i�Ӂ��v��ȶ��Q��&���Ä%]���}�r;˷
�)�)~�d���(�.l�fG�O� d���+�[I��O���98l���9�xp{� 7N�����>�̔S¼�~�S`�N\^E���l6�8�씈�'���i^=][)���h��c������o'�=Z��4׎c�~O.����y6��b�Z��Rs^??��jP�-~���� ��rB2�L�"	.�h��}�!.�z~*�^s�m͠���P���c �1��q�|N��eT�g�������	���,��H|�.ȸ��'����m>��b���z�W�>�볤��w�S.2ɔ��&��@ΨM�v�#2��4�5�
���V�s�ţ]�<�a�= ��C��.��}�Ҵ���T_�t]YY����b�M	�Ӊ�@>��	�ы&��2)-G0 �w��gk����y���~Nb6�ݘ� 	!v��G�Ë�k"|Ѧ���8*f��Y���U=���O���h~N������y��J��0���h����V�͇���t�0�~5G�n��ŏ-�M������@sܒUP�zkmꑻ��'j �(�������9�@q	
�锘���c��Q�K η��>��{���i�'X*�4ޜ$CG�O�+)���[Im����������6g� ����O_����%�r/X�h4v�:�̵	$�(���V��M ���u���3}8��}�2�B�bM�YW�j��8,�U�"�<��a���Ü�w�l$'�0-�PF�S��3���l�<�qj7ԼI>� �?������I��?��J*�ƒxr�<g�<v����RS��A���6�	����)J��/��!��i� /���ld�jg�>豈�V��5�B ߫ ��ڿ3
��ҕ/�+�iu �ξ?z���ȶr�t�����>!�W��={��LPy� ���n�40���$-zޏX����>�"Qr5���Jj;ȳ�~�Ɓ�s���(uc�l�YЮ(�5�{�H�Hz�L4��#'mL��� M�
~���Dgx�@d��!��蝮�F+}�h�����?���j#��(&����w����_w���X����&?�Y�0x̎�߫�ょPD�1��m�[[ �Z�|����0�~]W%��+na�K�Lc�e�ьX�Xe�0-r�'�W�-\ �Wy��X;����x��q��;��s��e�1���#Z�f)�C�3���&`�MI��Z�&������!�Ϗ"{ժզ�D�CXJ7@�lMr�m~�[Y��A��_�>�a �>6�=A�5b�I4]vnh�$��r�oh@�1*��m�v��C��)�CCUJU��MRP�\o�����Y�����5����f��5m�����π­��L��x�h�綑aM���G-n�t��6��~�+�&ZG�"�,�f����K+��7�	O!��UxwK^U�
�!	�l�|�s�K��}��,��Bėp���M4.��A���P�X���C�?�u�@�u��%oA�ٮy�������l"d�W���6d��`4)��6CЉ�f���B����u?��&�4���C�a\Q̾p�m����zQ��5e1Z�B�26ٽy'~�٣��G��.���"���5����,����t	��4ԻȰ�����mxz���-ID>���E���?�k`��'~�fȘ�u+)[`D#��^���9��)���h���3��I%���F��)r!
�ykQ�;Dm('��ݯ-sQ_�t��ޕ��Yb�����r<���PVJ�A��[��5�]^�~O/����)��=G?���F��GS<.��\$}tS��Z���.y|�q����P�69�9&6r�H]�̤u��0dm��-wm��i�=!��s*��<k;�_n8`���Ho��eè�����zҟ���B"�f�.�\��(T<��z���ç��'��2{,�2SV��~�[�\��5�a�̝�5do[���j"x���H1�h�+�61�/�F�.�x�q��#�l�,�!�Y`N�9������ �4vޓ7��:�ڮA�^��R~V�U��w��Y�L� D�Q�G�$�6��s�+�$T�� 3�ʫ@3T��e���m�x����Z9�����s�;і{G��Ô�u���׿�mn�{����>n�"Qsk0������ng�tT�4gA�fr�%�'"b1&����1�K�켫$��%�{nฒ�&K������G�����4&^-A�+�l�Z/\�q�pW��!fbO|�6-}r�GG��Bч�*`E�CN�nU�:��A��t2�i�π��楮�ev���ݪ9����X��n����/P$�\S�;�\��!�I mٹ{�o��kS!�s�3b6��Ǒ:bώ)�>�����	�C���?��?>$>I9��"
���Z�y�y�����_NU&�9��b�O��r�Ѥw[������Sr�~�Zaú�fLsl������,��#!�b@ٜ`�I	]bS��J\O�ɜ+�ɱ�Q�JѶ��hR�-�?�9�ۭ|Y���CU�9x �b*��(YS���V���u��t"Z���^�ß2��@D��dH|]���:��|�W�(��d�͒�c���&Zĝ1�)��h:1}�iPR#��f����� �i�G�r��.9rJ����=!抃&i��م+�0o��FE1�$� ¿es��3	�EYy�㼹���=���u�m~Db])�ԻfD�[�rش�.��	�z��wH`��u̗�0_�k�;{d�4� 0"���BBK~�=��bR��;�R���X�M��\��7�(*��~�*�b��o�l��(�2�̗�(��Ш#E�����Ou'�FK):��Ss��K��o���@���8���z��V�&'R��^�2��dS�ɎQ�u�SÁ2���2q�W�7�qHJ:�b���Зݧ�~�H+tn/y�fz፪��3�F�mR=W��]�<wu���Y�N�3�>��f���D���Y/�ǚ�m�o>=$ٗ
�L��5Tk����uxɭo��˦5@�"�p&JM�����W�͋������ܜ�ʹI��6�
��ߝ�qďb���L&���v�{���N��FȦ��\Sw����i�NXkK�����fz��%����#��,���?�<~t�zvu&u�]����[���}�-�؄�٘rU]�K�c�\�%��8�c�	�����E{��Y'޹�j����b]Lʶ����� ��0�4�v]2A�E��"�xk��"9;ó݄R�6�#�:�b�X��I�.��>��?��e�9V|M��97��I��t9/�6/ܢ8,���k�Z����
;���Duk���@Ֆ���W��Njm���P��e��P?��\��)U⫿��FD"�:B�5���#�½�ı %��=(�0���Z�79�Q�au���q>�Ü:[�o���]��h4���ҺeR0�g�?L�2M��L�^�v;ɲ�Y��4�F������6��<h7Q��.Z�
:�*
��N�0�:�)�`r�l��p܋%��:y��}��������*#>c�����L����B"��Q0��&j���e�H�NYF5�2ggq�*Z�8Y��)/��{���r- �_���/+e^����Y���X���p���s����e�*���������!�Uyh���x�[��$ȓ�O�FhF̀V�"p�O����9�o,H*H�v&�Y��,߶�k�Vٳg7äҪ�9�=� 5����SE�����!x�d�s����y@h��k~հ�<
�+���c�S�8Y?����Z��@���K���LLi&�9�E�\X�P�e���uC0�ܤa�Z��FqO�+Q�}h���?�ZT.JC�Y�g������k:)s�F���h��Nu�6{o�+�@��FO;e�Z�S�x-� ��U�H!�D;�أ,&�z�����+�R��'&-CR3���](.�}��r\�I!� 7dn=���X.()��$�Ov��˶��@� ����z`�;�x��g:��(��#"���~��]���Q��p��ՃO�۰ :��e3�*�`ȼ�2�Ԏ�H^AL2��A�%S�U��G�!$Ø���F���+Gܬ⩹=v:� �_�ξ9%�,3��Ĥ���\��C�
��& X������ۥ}�7HF�vb！�����?Y��d�fN����r�[G7��\�r��N�����]�a����) ���f_8���յ���pԻ�Y=�R�-���b��/�oxg|����y��q;�1q�����X��((�\��O�	��	�L�����<ɣ&;ϼ�e�s�<�	İ|�Q&�ZM68e]�����f�#S�5���(��T.nj�p'E�8�K� �3�^w���bj��ּGg��GE�1�%�VŚ�������6���1���ؒ��g(	�:��C��Ӟ��6�U(�)�=�х�V�h~����u�F}�m��X��3*c��j9��v�ݚi�>�2�����ڜ$MX�V�<$BIs%�ď�������s_�b>�0/�5��:f����������
j4�����T�e�N�T��2�DϺ�Tc�� �yf��A�Xѫa�e�[x� ,�g^S`2&��