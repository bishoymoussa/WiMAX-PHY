-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
brQ5frQquvlXEkCiRXYEmvm3/hJfbZYrqg0zN179v/RSM6enVcr8qmNhYi5Bu5rUuwbIlxbUlOnD
q/CM9IwlOXHWmtT6S5Yig0x+BrdkOTjONBa/0Yo6dImlnETumzvaeOukW0WvwfwHsQHEGO4gIurk
6QcJOyeF0vOWN7Hc0hdSn4ByCzOQj3w8IN3CRkpCavnkC/llsb3dfPif8xIW/7KuOKC26g+9Vhjc
tAQocyWTVcktba+Mwf19ygSdNobLdx5yyO+ne8qqpkw1d+4YYkIXGxk3d45BXf84xA8aIvIKpN69
pvLcya0p3TQ+QwSCcrcqScMJfieYGCNEvGVutA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 47136)
`protect data_block
k99qODGOnQHMRQUFK1Dm3WGESH/hxIoFqgW4uCpQk4ASghpJGfMXq1Bz8WzgzRXLqkGoFbifHO0U
cHPQFdEsmVL6RuY5eaxYgOp/OVv0oMnvUNFwC2W/mFD/d44f1epZPE7eiigAltsQukDTkdi01axj
EtnifB7qg6ay7gnLxlw63MBmuo0TH5HmefvGFUH2//vClpRLTyhpNNyq6s0sMpLgPv8gtdSrBIol
INbV9UbUXbtU0Ij/HkFxCuoBNc/eeot3NM2CIs0mspVXYAWApISm5GDC/lpiTrtyvVe4pzTyvscW
jvimz6AFMAiiMAKomMy/W3ygjW8G20sBtanbf6eXPYibDp9VOY8ZILh6qVFgW1/OKghZLjOw1u9N
Fl5z6NIwqIiFkCuzjHfAW4M8m3QXmfLnjax1sjzRpc6nLyfUDY4h+tzZrDc7UnqVhGbhZLnbcdPM
MZaLCJHHjPsw5Ijm+iHTQ0EIxj9KTVvw2ISslRW9Ta9UCXLMGMUz+oLBEwd2Yknrj9GrdipvtM5Z
DHmIa9c+iC3KW2AsLsCXDbjFtZlzejgb3J7pwY/PAlgj2p19yHiREJEh0by369N5gIs/6h3R4zuR
B1Lz/MEfynkN7YQ6h2D93yfKisUhHDacQapo7PsSVPO5nQYRihuAHj9MNIMmzgORrNJVKAGCCHVN
0H+7C7L19mMNYNgC4iAO0ukzEdSuHFULHl78UR2GUv1jNV0/XR9EXYd7anxOWHMhVsB8LaYASxHm
X7tI+S2kEhp/VZ14dyxSK+777WDaLxsLkLvWToW8k9xRCAuQTF4H43yD8bNnBY6UEDEwsGUCj4oC
+8Yu73FuHCFNvOJUCex5svEsDIn1ZIJ06wxtTOA7KnDu8ueVtQdEnA42NNdK0JhzLJBXi6jOPBNe
LhU42mUsSQnl4B0g4ee0DVjSQQKjRDU288hu/qIca8DllL7+KqG+LvetCWptYDX9j+aZsfA5pK+X
szEAmonLWnbrFYjEXORjrnMAKKPniTCHoiDVytkg+dtcBVDG1PLqGZJO6xpoPg5BM+KuuuyblUxZ
AfpoOlqHF4gABt5prf2VY9HyhGGR6/pAVYrUiN1JgR5j6yfHTtuXI9GiwLNEbh5U13bgAOOL/Mhf
0R14v/zS8oQ5Yl+auGEpQc9Y6/U+5+8fmPNtN9u4kolneph1tE3gXuvx0UzdVrHfLKeq9Qw1iUFS
MCeHLOjhCIfxfdNBmIX0KzNLNU42qqPlzp3VSHBbBhR349mY7ytlZJSUUxdvuvXTa+P+jgoJUXDw
AYVwl2oFtLSWaujoc8ROYNDaVsFQDZ6pPNr6LS4ejMeVlKMJYm/6mPRVtd2IENaKMuDwbpu8bscc
k2RCwlu4piHnyhAixBQtLTQYB8GWrA66O+dzEjvE3nPOH4EUxGQzN1cEDTXp5T1dlb2H4LKrXMYa
lJEhWs/Mip4xC4upn7OTcTu4ynBjek42wuhHbK/i+vOWX0Ptkst+8HVQ0LmQCASrLgef76cVLEg7
aoJEST9gZKVBOKUBKHi6pLTgtLBOoRuilm91VKOvhoWSaMgzrRsLJlsuZ+G0jQh2IMxyN0baNPEx
tYd5CxIWbdncJ8Kj4xFHfGJrx6kwnGxtU9Lg0zKABOrIDq3p2O68j5309MyYbsud6kInhU/7pJnv
z3R0/LtZaPP4kTbTMqsCh5epg7jpiicXp7ylop7RIh7Gb1mjG9OcylSzUE1XVgM2sb9wOU4OgVl7
2MjokTecDzKCG6pH3pSkfggVJqFbDMPLI1j6Exrg1KPEVebRVIK90I+/9EL/34SVI7h0AqKP9dlN
ndWyrQFV6lVfUYS+Cshm2KoUzTKPITGvRHKssz5ZTil8GSsMcUudjbwe83l63+r7AKN6dKofHuDU
naDb7fsjTTjfgl9yi8cw3Bd6sOPJmOWTqo5Rj5OGjlU6H73/e/8rUz+OeL7lNteo0RiDy6HeEBCq
tbIW2V3sHjdSCUnrnlRNlqZgaJR74OcvDLhXz9yfYN+7Q0PosYCTpLe5tXLyj01YJ0gQ4tn4AuNG
OELqedm7ku7F3Sy5oh34v5TBMfIOQmG/quwdifA/yc0eCcfUHss14XX0SiWuOsOF9mEGTBhRHtCy
GKWe9Egwdtz4J2PZduWm714ghvJuQb3dfXj7fOSx5qlLImNgAiqZLrsYHm10XeYQ6Ra0Nn/0ztAT
gQ2+25pNL8VFBd510KnpvKEjU3nyHNvOqrQjx16U+SNcfFx8Qfz7h5DG8HGnQqRdOj5dVHRWz/TM
xABAZDNrsxt5XPF2nWhYzrnpLa4B9aP6F0BoNzrUJxzAe/cbBs65aEid00oYHXVcFM1Zs0kP5/AM
0o1GmAJ3IrConJFLoSVea51PXza76JVmOOQzv0X7uN7aivXhLu4U3Mkf8OeGwz6pvhmbHOi45IA4
nO9NsMXIqL2kR2rZpFXM3eOLjbTgAp8DO5nZPUbDmI8vJ6CAqK1UvqA9aDbYMyr/FhOuP5uV+pGa
XudbPtP+1AmdZoytJ/9qgBwfjmWdnu/dbLFq6N1A2z6szEXDd0T6MvD5td1Iy7yHtw3m9hyLwijb
vQa0vfIrn62nT2lVNwKKB++aUw5gmZopCJe7a/GNw43C360ZpW8i0lvS9SsWQRTlLsKKFd31XBwb
jQVq+FFKshf7QBFQUGZW5Q8A5B3cjX+Md4jlSYIcbu6oXYI1gMHn5SoPSx0tOMKXM7l3TRACsjQg
wkEgh77nCwvwonCN5R6hM3T2BkImkF5icSDZfEro4agpf+jujR4n6ReCP9Ou0TUT79cX4b2r2y8n
t9jdiEKZ82xqQyi3MSgcNgOHsAEiTMyHh6Y34vZTrM5sNU/ELT4eT5DnShT0t/c7lahcGj8ndTlP
KNu4kLMOrzUxZH8l/DjkowiboVjOIsMjfb/lEkcqwcIYqQXY4mK7AvMnzKcldt9/X0uvWVvzI+GU
9T6ZaOlBa4jdG94UweLC3egyZbIgWx9Gth/25SZDPuQbUzdxujoaV9k7VNPdNgIUGHG3h7i2EKpn
EnwYxAFXBTt1SRznPcKJcCaej1ushfYvYk8V+1yrKVIrXV02TQuRagRDRNlfj2EsgyP3012poyy9
uo1x21U7XlP4M3EpaVtXefDo9DzSy0nBv5FVu9cXufWm64hItsX/4QrjLOrFmp98xd50CKtvEqPQ
Mhrc7w6O9g3SwGeB+16zrglw6Siv0d4BEnpL6Gtp7RS8fi2HQDwZ6yBmEPAHExM38Zdrw0T0R0QA
Jm/51Eq44BfBZFbCzDsiN0FDItlgN9n3awBy6yFemyw7hwHh97400Vc6m0NgefnmiEOjJbzgs5Nr
aQQLlOkO0TYKOdiZ5uctMvQwkowSTWPKeEmSt27rKuZxOVxPZz1tGxNhGJ3X7NcZn00M/tspXfRg
YTs+EDdDfk6RGA1bpk1Sct4L4vqksZgtHU0sIbJ0kAef6bJFo+kyRjdcn592lM6IBhQRQvbrwzpl
RoAUogUrIHXhMIDMpo+g10ACNl8yko6n3EAUqkm2ANz5WaXAStdGB8s+4lA7N8ZZ7HHaD6oNWSSs
U+ttNYK2ASU47/2L5ROppTi+2xVReJqfN63z4vvwmi/Zvlwdxx2+KmepwXr73xp4SjbJ+4i4H8T0
qwjNkJHC66VUxSwMc9YUwWmyzDk0NJiVywEwksW+v6qZWsbtCkh5YTimzegTidF0YcXGnAR/93CX
/CdrHh+DhOoWaf0HLWrIV6D5E5aEDy0DAeEXonluEix6lWPLasFTwvZ4J2iCQ0rLYXUW+6aUBekL
d9ReMovUdAh8/HLRbc70rOWM7EuAD+WQhvJbZPxr87t3DYs/Vy/OqFqMq4MQSzKWDhK8oJF2YCkA
DTR0CfNSUDFzYYBrwwxbODfmRFpYBEIQ/Qp+hl4pLJ9eqgbu1WsDTrn5eNF2281QCqpNMVOd2v0I
KvFvIr+DQ/H9qPuwz0omCeWQPIFHVOx5GW3A/eSWplUkxwd4P88VbspQoUpw2xId0Td4qYWxbZgI
vFWoyDLNbvBBrdgb/WxfNXW2wkF8oSXP+rAfK4qAQjlJ7JVGlWBZ+AjZmmddiBpydsOu/s9rgjwc
ec8NSIEZg1CABv9IuvzGhLmrLJgUp26RxUuvePv9B5y0tZSKeZolyDkpp8PzsCOIedcxMaebU2FF
d9olc/n7dD2ix2W7P2+chzCw+Os55Snc6lIt5xVNVewUZy0LkwhkiJv566P/lhy7wDevDPsGjPBF
akQxX3aXUvhRmtsyk/AbGVdzj5NRiJtHMDl/TxkNEtWxRIyrqI0pl0CY8I8Xktl/WgLgsW9u3TiQ
GccxudbwHQEVpgeFV3k4Sq/Sb1wmWgoNYd8i98tNcliQpXOH0P7tNvx2IrAqFAZCedV1kLprA+rT
hv51rNmZAjsIh0BcFwtwnd63EJRTr0gT+DnMWojGNpyAHwK0W70/fVYesefPQ1eYi2yub10+5aAh
wa3drKjHlzqCRqvkgHBB3CqA8YSg0GDqcXB4uptHpnyME5QEQqvTFez60ay2jUh3y+e9UFKj3Yhg
dbnJYeCouciD3Iz/P/MsG2KOQ3noFUVYDxChXmCThbdzOPipzGqPTTpYA9uZE4VF5d7Fxq98zqrF
5J0Lyle8MeTiotnW9PIzaQsiOx6Sw346AiUTkqqIrYH0IJV1IuET7sxXj7kFCiVP7MzhrHdn7mJJ
HidwMnjZaXoS+r5oK+XgVTVPINeDyLQ/wlPxJ+zZphQkveMeMa4QBnn5Z7S8ADK+drvy61jrKnbQ
thIjiJcjzSPdSRqbg5J2iWnh6wNDgMIG0XjSmvJn4k5b/WeougT8RBhpxafE5mQP9rOyC2hXhEop
/qi4nRZm3XiUhZpZFHcJmLyJmRN7ej/34NCPGPiKCq+3q1tTsvh+pD15UJ+pHOVft76s/VdOdKSp
PdpnfeGAKoejwySXFco9aoM/L6o6PJT6LYgIgEauvzd8TZYTCirXwfXFg8Cjt1IVyR/OICPL1Yom
DStGs9cYHafi58bUbllhl0TD83fklA6BqWjoUvUSW8pLrp/eJCWXkqWcByxOSr7k3DD0OxmjhRFc
y5a1faTvbLFDvx68fOJRJomtOMcuZg8/izS6kj4fRXB8jE1wyMWr1DUPuAFkirpzqM1ABHX6OAOL
H9VZ+4PSMxjDq7ftkyj0IzEJ5UX3uwdVJz94WymXJaCJF3Ve7XPfGGuVe1c8isQ7h7LkdvSl4XdB
GeH5B+wf3poVN5tZoPUEAS9qvrvGZkvWjCxpF+vvllEyiv+Na6XRkOafxGOkAVn8sBUkNjngCzUl
vrs1WPLhF9hyn0fG9QPenbWAJsMsL2S3UVh58055ZSIlVxHFfQL/N4diJYwlNYjlEQJVFT4y9UVt
EgDqF5TFVSQl4p0jU/JTTN7nRTw8tGs6NIwGUdhahuwdIQCGdDXbWeakyZIU8xqZs8QjMZ1Zj6Ns
6gjJV44iDYStWWbaVGVIn2eZDczyUlHEXSZhAaA7w+3jomPcGp3Jm6A3rOKZVNmzlSsro9B6lnuf
MdZvNv5JKR03it6OsqGyWP6p3OQc2hXzpOjIaQewMg5KmZh8Ew6KoS410GE96cGK8wDTh/mNwdWo
RAtVEZTbYV/5FE6gWXgXLtacODym9cv1htKAScERrhRwDHuRhR33vpHzhGFlxgN1gR6F+nsEVPXY
OMozEwgy8FCN0aiczdaKhcEq8xw0A+C080SOnFR1H1BcyDtXP1yV52vzkUdt1H05+t7WHuK1V49B
wnziqewW0CZX/M7fZ2fWD95h7EDh+17BUO/lU5pgFbWeXmT2UN0SkCD6UhBjel+cXaZqk8BakG/w
foIXrtfcJvwpxU4C/F46iryWrHND9kWgAzWeBKwl/1Mv/6ib4xwb0toe5REg7qhhEW0OguucZXld
aZOq2Lqf3Gmu4QII5NIVmIlic7BD9Lp9TTmJ1t7CL3Ra3LsTFnXd6SQjzl3343bH9BKqwBqmx4if
SeeNtP3CQXFt6jULgYxEGnXh0pFAjym8rRNRwyhEQxSlrdhKxoHIZjdJ0DQK0RPp1AdWazbszpol
ggdlNG9cMU9uBXO+o/Sq/Dkmadj7muLlsEfJKcfOKVcjKZFRlQM0U2ev6jSHvYbLF9QzVDTj/857
vGSyfthKlIjWnENL0HNvNXvz5cL9rEbiw1Mpv6NHXHzumz1vUd/3wtkmzvWEEDTlTQG6TMRe/Cyz
KUmfrTMpoCd1JYWh2WbjKGM6DdLJ+Twn3ve+w5GedGpUoghtBI/g2lrMQzVNLXW/QR1vUnFqHAzs
kSVAd9Edl7eAcAIHwFiwXWgbMkaFo1YDWnXx8mLrMDl2TW093m17wE/cbD/i9iVOHGNk2LU41XwZ
sHT8ba9d0lRC0pmGtuhYQnidH/UjfqCbr8CDDk6Aoe5705RxmoYifNpJCijAI2X4mSSgJ7EPeKHI
N3gGx4VIcg6FVGDTj+Xw5jb5hXSs0/nNZgVpAXjnkoeQN09uVAfFLzUySWIoQLe0rh+PoL4btjJ/
r5LgIKmv9U5i5eVXgpnEQahbrlnFY5KrtR4YccbfDzR2DEpgC3fkcfc/9gfMOAQqpIk0dZhbnzGp
CbEKFCxajO1bukq+HJegQ6VdvhLP51tUzNgVI62mYgsfoAfXC+X2WsTn981UJdKT053rqHPSiQ6j
NhtnOKPWLcjBXQ9nFCRKfxj+DP+UdVeERkvVwF3nWAKwCZSW/lJlLwN1VXYe01JpGR0zSkL90IFj
p7PjTRmWM2+qkIs9n4qLGEBojI0nuyZMBUhJKazrzJILW6s+GHWAk38mxHoHk9kcJLbQrA4m+omG
KsbuP63gPbnBug8mBfDbERrxLm/7iYqY0E1QF51ICqCO6yp6pspYrl7Snymg0TfTNfNw/rLgeiVC
dBkG4d1HAfng5LfSBxbxjNgVcbEPeSi87nKwgMF+ltet4ZpQGcL/grOCrYPOft9PRrfN8MrGDH2D
T+4snlOPSzWSusZtzU/AWBU99CGklRn165z+Kr3ThncrYAq+nkpDEAH3/AWb2oUZcEhfDN+A+BiK
F7EABSU0I1K0YBWKbfnBz9SzjafhbVlAqWqht3l15QTaXl2WW5RJHLNfJiuF/31pEIF/YwHCWeoj
11X4S8IYfvk7C4YLEGWtfqmzHQeDBXE1VpUAI/wm7f008qmDqKSkN8ZRZ73sAMgqSyhWldbqpAb9
j3EAprl3s6JiWJ7644bjqUyTwzQWXsvo86CedZQHgKZX2jMhnG6oTLSwlDDZq8bDc4C4kyIoKhfS
C3ZMpptH79Jt/Y+jg54rPy8GMmfQeg1G+MbS8gVIP0nxB5mmHvrgs3BZiIzY2XMkbv9+wS0YiE5S
6sCw/q7mcAZ5hwbYXQksXqf3Io2uLPnpt2IHNekn1MphB+FYIUA0Rabs0Gaoq/dZCSbGlc8UYO+j
QJV0i0DvIaIFNeUhZL3GV7XmnqzyMvQq6V6my984tZqK5Tp8ATIr50yE1J3ibTBapYmr0K95Vdt+
IKISRdRpT3VQXo2AVJZYT8LLlBvJmoi9kQRYzlEivw/6ag7WWgct5aHsqeOvvhgdAIFuHDPoOHmo
dOPEra/NE91v90QmL16j6VnAiHyiTL/dTqCSw4Kc787RNqSoM0tTv5LgfxaJTywIxkA2yvwXPE4V
vCz83PEZtKFSFY7UUm7Rx7gPB9AwhtGqTeYgPxT7qNKOkV1b7oEFUrfaPI842nuOtUfMx+31XsB+
mpbwAzgS8uFInO7uGdoJdbmGYw1uzZsxWW4rhE4x9+OhH8bcbZjy9j4B2vClbwqW1IgcmCm+cF3k
C1O6iv1nDfaFmK98xNILbhkDRCA0A2ah+K5mcjwvIKkR/QeUuE0aS2fJiz4BANadul2N6LeRZuC2
gL4M1oNFXT8EQ1joN9/qcF9h1yGLkujimOuLUGz+gFEjn2CasQZY70FG/mOeQw7vq/G31Kr4HIdz
WtT/IZpkcnuxgYmAFJr7ZmLvU7L/1W4fC7tgLIIUtDXtEpIwJQgn52zyG9tLIm12pZpCaEUSnHqA
OOKJ/MgT0fkVttkqoiuFw4Y2apSsh+5nfeA143bsixp0GoGDSvyKcgpSLy9kh8p6BE//C0OwYu6W
NxnVM620SWjk95orqSDeFr8EdkVw6Pi2N3GoVnLNDP81WQ7BWO6SngQEkEHlKz8k1p+Nyl2yVfRC
HrE0n2xtTf2GUgE5erZNC3BmQTDsIcUkYbh8rwpuc9O6FnFB1hY8vuovdd9pqYtb82R13OVdXcfq
cGww+e5huTR2MKsLJSUirRpy0/hSdcFRSTQRm+jvY095qCUaX5ljVxIfhgR338vIP8pDPjC+scog
CJfoVMW0jz7qrXNFR4cj2rs+0IA3YTZQ52wJBhYHl3lrgUBfLsEpJBbqO/NEek5udD73Rie/PS4T
WRMEgsQGa3MBB0qpqstu8aAWpkKfEGJJMp86JueV1jvJlBP3Hy7ZI3qxcTE0vrGalSYwiImw0vb9
Xy7tRqGk7j8GDNk5+ER4JtbNHZkaZ3mJLltobzOIu5pLV3WbZsOL148TJ1nb5Ib2gv3TOyWn/Fcj
h5WFEToGb8WFxyZiDeJTOjOLhS8p1kdW9miXknlw8SLq1PTm45ask6Y1pJxfaZ8nlcA3zVEzNf/k
zO4wIMjtl8IqfBX4oo2Um4EbLNxR31zC2xnorFwUB0Pig0meYfuu8KvCppja1L65D246FBkv82Xi
rCewz1D+tH84d2IZv/nyatMKCoiuuYkgqSsQtQ3z28umfmeTgpEViwkeukQcEcWCsgf24QqUnm4P
cUfrxX8mfrufgRQphpmCv/PT+TRaHgFXttiBziJjIFIwDVa5danNjPxo/g9nu5s1Qo8xynPs17xy
cFfapyhKw0e3MxLdR8WGNOKF1xWAkyEJMJkTx2m5avwPNFZ2g6/9yN6OwehgHRCVKdFxTyX4XM6z
v3RidmkQY+582dt70gQMYcxfc+X+KYNuStVacimRTsaoh/eLbWqsaN3Rtxxe/qFeh5ew/+0fAjq1
PvU9S7abWfZmIlshJkj7+bMK29NwBvoTkUVSMK0rfZx30OKYDR2zXBWv4BkE2bVb38isvZKRNx3l
ZYFIJZOtNF8m5SrpFmFcuE1C79XLIHYju1Ov4F1iXqWJPM2WNsy1i3KkvUCPPtW3H+d6DCRG+xx+
weMUuK9PhrYBaj2IkCmMK2McMUNLN9jEXdvG11MbQg9xf9ZqrE0n35siCwukmHUyqZCm7/nYDyXf
1BiYP/v4UKW6OE7bfjPBq07Y2baMoeOykjGn6Gal2MmeFdI3wDAzfj4vI/P2SVkvqt5kIhssmL63
kt+PCzp32l1Nr05eErfL819oqwE7aHZjXCxlSHYnVbfQsMuWnbJJFDmR6vk78bKb0AsJxvWoDEYz
E33aufA6MweYwttTSb+y+aK0w0IG68lS4fJNLXlcHDX5rsJHZW0ukKSq5CHQH+jo2MfzVDPNik1z
Mcu8zLqEzxIwH9pYiAnjVlOSaYS54eI8SzPwJA4sdBn8Fx6M6NGaahBrk3mzDWtzUdgyJ451ViHt
ctU2q/jgBGeAlIG3JtioAxM8pGEomx29MIRy5x9SS5X3fO9rDJneZeFN/N5s4YqloEwFiY47YRCl
bUnmNGkepLi6avcTPgHgd1DN/IwUNRlWD81vFgsLoOAKtCR57oE9k0A5TLWU5ulT0nwYpG81F4Yo
YUdE+/6YYtyP/IEJmgqSTM1pUxamgN0MJdlJwZNM0HY+nFWAZ3dKCDhPOI1KjL3G7v9LJJ0XYwWV
NpZ0ZsG0+4atDeJW7i2zUpeLh5QCRXQFTs5+RtXcknnJTrM3x+a5aiDdA+mW7ONT3NV36VEE/de3
AiEQxdsrhmx4QyXZBBpAJy3eQp5CUv4yvzQUfDDbmGSwu7xB7MM/yCcC8sgx7H8jOpIRGdZUu3YG
d/5a/0ZeVRHePKQhRfcbdoVuwMh4ECs+ekmjk3E4+LnoX5ee82efX2SzDPmnh6+k/KBZyd3khY/F
ayz8JeHXiyQoE108Xj4wk3LsdS/rtm3VlxvHZhL/ymtH/l+Oees8w8hRuVvsEBzCkGLGVEUKfA6e
8NFGWP5RsRAYYgSVI9lfqG0p7qdEUNfUj61XdpU7B67VV+LiHAX3hLI2doPIltk8qzT+8zOUR4vQ
q+uPVn9qNrLaFBkItkVO9iS9cbWCYNjisubMO43phZVpGgRcaZchVIWUHm4TgVdAJMVMrBnI90gc
n9TIlmGLCRqGRwxpsikQeQHQDIljouABQvDPcUxx5g96da0Sx59QqKKW8HhYiWJO+9XmKQ/jWhph
ayFgWjpbgWvt4VXiMCeTxL/oHjtxI7eNKN7Fn0NndkMK8Is/bdG5VN2p0bwyztuDsPROp/z/bYjs
7DVdVw0eP5VVTBnheQKxOOU5B3DK9V3/+pXeuSYExVpq8A4xJf8ujVaPB4yslNwmdhcLUeHn8iBK
zr11OMIXsz+1KZHJc5Wc71IWUYkCQSZxO8Cu4xOzw/M1obGb0HyuLHFRkV8RGnrOujQ5pzZIYboJ
lVYbOKXufOffRLX4E3OPyhRoQyl2h1GbMFmLjRdoOW7xmZBW+0qmoKRp53E0q9A3VaC39LJ1NTUV
Yb4H9bjAGtJxedjszlztRfgt2G1H/vPJ2W3Wwmn1AU1Lk0X09++cuUU5/DMsUciSL0r+sRZUdJq6
EJJ2G7EafEEXA4XpSxdDuP4YWsM/Ied/INUn8rCMEkt/Dj/38R0gUSUSfg4jED4YFHB50ZjRhAug
zlroxKPV0dHYu4MVgRpwkokQLux27R1s1Jg02TWq3pgT/0v+dtXF0wLXxW4y2PvrK7NgGpF1vwqC
kxAHHG7tMjg0NTJbtn2PWzaiMXp5iSd/qAT1QqKqLqJ5vq473p0SZK4AoDoIGxQqkPm46MPFUhoM
5phqsLH7MCKtaU0+vrd0vdRCAgfymkdWY979TdkIULj3BrZa5Iy4YClny9JA4p6Icma779FshA0J
rR01n8m4x3s+sbV5E9gukN5wa6CiragVidBp8+TBuHYz+oA471Tr/Ht9C/LqWJVjJsPT9H6JSxZt
jXzLopYhrjFIFbKZqxf4HgTTTTaa51O/A8JoZjzH5pbB8SvwsOQsOSrB6nJQAPCRRRgbO6bhHn0O
EWF2phikvQtE5iAERINVgQrCT2vb917WdTWHC4Hvl0FJwxHqDQDZqcS235VxXxyASJ9yoi2qJwip
LVJTau944g0Rzjz2L7FgQQ7sLp1MfgTytYnhCyOc05V5wLrBaiMdIoYkZz2UmvwGdyecH7MhtLxi
MU7TbSbPh0a1vdctku3xXSf3jJ5S0WtAg8YHvqq5brGMXfsmt1zFGOMbM8pM0808xFfzqtOY2vzc
HNowv/aR2w5/ym4aEUyAKCEbgUiRsGfnJYH/TEk1XwqO9/J3oRHDY/pP89mZpYAaWeYyV/UQ08p5
ilMmEeg2FfytzVe4ClNBcJPd/iiOdkdp/6kkyoDO8LulxwLVMJhuOU3BcrEwu7rRzUnM3PIKbQbx
AoiCKGZRodoo1Qz7669a8oF59UJ17BrCEpzqpHP5TgBOQCEqEJgN2AmnjwuUYfHMeQTwaZOWBNp/
2NT8UVzyrOQdSL9L1lW8ff7Ru6q0AgcLpq/MwuALIs2o54Z7lxNYCxkF9kmLYcICXRO4qL17XOfD
vcSL3VY9FgppsfvRh4+F2lBCKy61yGpErli+q9olLHhrCOwC58N9k5RXCTYincm9Ph6eiaaUCL5u
jEyw9NiAAkXbuITiiuU0ov2O5oDvCrZobgVS/+TjQFySNlzdgds8efu0qAgHW2OSflXCsOqMhcGs
uBLAjkwTspyr52OfAz2/CV0p5nJW0R1WczqeCwGM79v8Kabx3V1de1BUkx0zk3iZliKbUjLM5U+Z
RyUTwiC7Zk1UB1BRrn98BaCoE/0glu9ZcGCEvNeyeic7SURfG8PBKKlrXZAKW5ME2rhsTLtEv9ab
AuA9g/iAtctQY74JT4UaVkOxSa1ofGBJnJgSkZlglf9RcmE6UwQLlZMB08Y3MdlU3B6rst0Sz0oY
rh6bQNbhW2LmClubMInL/nw/39WyK/IvzrZQWHRBjXat6k1Y97mjRDKr/OdgIyNISES8ujkbYbco
bhD/PhdBI/oep+/o/3cJ4VOSB67xIQMW8YqYhmZ6rB1VWjBJjTWgfTnONtgKLI1PUMfzvuCJROhq
AaxkeC+fmFGBNI7lRocKg8/lJfqRK4s9zGGvFawhGkY95r8MHQNinhVEVqLEAQyXJdJoyPg8NRRu
qEmNyo7/m6a2pS921WevBtIwslpGWZUUPMTHVSB91tHZOzWxo7+F+jQYy/c8DoLpZK2NAOAqvWWZ
Xju2asTIC+drzMg8OINPx50+7MlSQR4nrGEVbtkv1DWI7jZWw0w7Q7zS8T9DgS3c3zIQqUB3C2TU
2bLZN5lsLGbFhaT03cpxADaghSZIxZ4uFuLDBRNl3rv+rlInnCPMj6adokTxuHKIvKirbLaXLlbH
9TmPX8bbsngVmM/MAUv9z18EiOXTfoGdi00C0UkTlOMgMpTRQu6ww4LKm9B3+zDGLy0O+14Sp/jt
ZEr5DQKsY96O4GsUkuf3QC9cHQt9EZDxrB3OxJmpK/7N01SsnXNb/sW9rMQagqZH03hSxSkwIChE
BaRis686kjDWpICjlrq29rnbwbRlFExAmOVks+sdnlwwBez7b+9ikAvY0tjuIRcnRI2HNnW8abq0
V9Tzj+p80hJKaCK1i0qMUS7mDGjZ9dH/k/KPjPOej/hdgLcwNdh2ycZQTMeLI729VB8r+LTr4qFF
WIoo8NDqMmCyjSVKsKfEXOwdYt3SQeq5lmHUMkNLHbPVLf9u3YoV60/taInheAttd3fvjPMSLNkM
T46ui5vi+hVLATru3iu4Aaot8dw0n8DM7LTsQnM7ziie/i+ZjVErpSqX7kYioX1ECJXmZRIXuduA
HrAYB9D1wbqJzrhaMlALR+UriESzZSjQMB3ZZYCzqqdjiDK6esC2V3SMUF1B3FK2kSKapzF4F0oN
RlEtau3D3X4XF4/41vp976e8JfloFT11PIV3IFKoxvateV+5XuOEFW6yniW1+JKWJFMdFzks+ZNh
THqJfBmExdlSF+c27IqtZSZbCQNz7w4kfR5I/3tomNVrVlnszVEJ4hgbO9TDOHUAw99c0usSP6Lq
D+xM/JFiTQrtjFTeyfXDZvBOwe61fD3LXLJCumpIo9/ctO0HORLupOxJ1GLNQYKR8wpM/pRPt5XS
bLy+oHzX2nZTF1nk574+/lcX8kURJMHFImrRRa/2xdi4rIcOVHCsMEeIHHnJ8ZNY08i57LGu6szT
G+VTQFbGM4pW02jdPxtMTl3iKC5tNYPk7KtoN1p7haShTQAweqpX2yLI5o3JXDfqMAcEVMqf2AfW
ZTdPn14l8k3jE2CyrdZCaIfRC8km6+RAmoUT6PQvNJYHj/otyVyC3++E7qqpxanQQa0dm1S/xQ87
n87C/g15FrxKfmzCcag+08e32twwFoSiJtLziL+EMXdaf132Fy/Qjt8f3PK7wwB1IN0tdCuPOCM8
I5d0DcqHBwd+zooTlHBP55Jkv92E3LKQ8LJXeRFlvG7qVdUUkvoR8MPrkyo6OP+bu6wPtT+HKkYF
i0T5Rkf0L68UPsURNMXlPyZdFSJX2sTAk7fSYtwI93Xx/ngB9++tR/RjD3ByeulQVKpAjG8a83WD
7HAUV5PukppBn2KXmIqR+XlXs4hwgk3gkJcjtp/P/iqSadqg06fx729fNzaXnaHgIaP//IBE+6gG
GyNovwlfSaoXO/vdFllj61JDSXybKpQ/7MI2vYjMRYD68L1IVF33azyu0ByrCgvklc270YENK3r6
waBf/+y2qLKpOIeHqlweu+IjiAzOaDTmzeCe1095xx0rvGh7RHNSFdRmNFN41t5R1JZsEU7N+GMT
jfOJV4Zl6IX2ZXMh1eqXCrJD+SrzqBPGWNStZC6n79btCGKaUEMuukMSy4faYfeRmeaV6HVaXNUh
ElhmdzGfiU2wS4M7NDAZWWMlw6pc7Hk+aEgXh+ywTL2xAGPTVUCPYC8eQEz0xn3c/TveOcrQdEim
HywM0mjbNNdmjhgCjIkX4Hr2U/dr7jwWHf2BPdtcynxXntNFo1kqkQU4EMXHUi6q0GrReMdzyxLe
ERy889yQSOY6KUCrslOZsKAIeQCkrvs2SW20zcWQeOQPjYfZ/sb/++8o0S/iJUAKyzetMtkvYswW
twzzXO1SnJveB97tJrtfLutQCcOpmCTH8lXnhpiRychL66RhLyn5F1YArr77Ny9U1ny6Q+BAp8S4
PwOsMjzFyZIXaBXqms/Vjj7iHY32R1uUZ1i4zxtwaOMMvld3nwSYDRQSi9US5d0PXyMqJsqcD9yv
+Efap3x/11pSMoEZRUkzNBJJFmlUld2/LBYciK0Fp+YCRzhdAiUrsXttDVGKEmyynKuv4POrIugx
UWjFaqfskElvfOrSm5cbWgA4Il2oUlgrjWzCzfQCMwMXbMILD/cZgn+1b8pXR2SjmpdADSA4dHKa
D3kJheC+WZulFpVb0H6PUW6bq/p31yrn6IMqIlWvz5I9euDxMCZO1y/xclMnLOvBukoVBabzu1an
yIPxhAw7FSndezFkYQkcYlrrL2xdMwN9Qpk/WfguoofIx2HzZ54ZM7W/srowOLWyGZB0Qoki1JwP
SHTCGj3opDFGbzF+J+RFsx6A8wGXH2Z8dUmIRf6XfdvgEkIgQqhYKCh0GQXF6MTCuCf35DaBWJtk
Q/2M/CeKLTUfcMe3QFyI/HoNhbyV3uAxq8X7ZV9WOdoIFpSFcie2S6+FiTgPdt2FeMlSgLEGi80s
GVVgiUebvDBcf15OqNBsdwuO3RtyKB47nCxLc8MbzdVQfA7rH7RKH23bw8oiRbuQV4C4i09TLheo
dkDhNU3QpBxoYlCo7UKA+PwNZs1fHRWMmpTsrFq1TtzzWVMZFHFh7qLDzoLGCzvc7Qfgm3TPQzvc
SY4EWuv7xPrajKMjDcLK4RhjIvgDoeiVBfPJo0G7mMuwxYeB+hHEQiWFhtItdA8O6Z+sLa4cXwjV
I8UIzN56ra1RS8UZpmilaVN01hc2mE8MLJY69TBn9sxQJT7PlVgtawb8WrQSp54hy6f1WUZMf4zE
ty6demF8HZufLMtSg0Xlh7G5NguEOVUYgiHZaeLF2nmMS2BscYpoPImEW9pnqnkB0oNsdFWuiR23
MLsO9cStWBKEpI64OYCYy8n209a9n5uGyDy4H41rCf0vmEMaMUE019HCCd1vL6n15y901PXXX1LR
tYEiNHDM8aJcL379aKKNLubWbL4vWPZe23HJfzAK54hplWHKKmml46L1LDjkdhFEilwmr/BpRVQQ
XOLoTSCwYWaRi8958yDSNzpsGoJTNuVOUD2cXrUgfCnouyWZG834BZ+yHKAJmBuTDFhTh2psoIbl
rfHNSXWoEcZGihhNXWxd+taXGuHt//nqTjfuWT2pFwvcsfZJvB5xx079JMqH+jSvpTTg4eP7Dfsh
xn+Hda+FFQghNdLmS6ZBXqNUmC/2WgqBL4VkQTwOdbXvXITjPT3MN5bDJLK40yPmmgtsebat8koZ
MF3IGomAAeR8pNfcTgjeNH84jfq5erW7NliyzBSBQ4OQ6GQuYUQKsa+u4ZDTehzb3dd9WLBgNbB9
BODi4Lw1J09kpCUXCUNURjWF8vrbv268zYGzsvKzxS/x35IXzLGM7kPEhQL/c08+eDpv11rT/OoF
lZtemmbxLAeQGkAmgAhkx06zGuHpA3E2SWcfINfB02fqLZefOh9JDOc1TX31s706nUYW2wN1Q059
fFjDYUZqrFwMeczMfTEpg/gwVYSO+HLWjyVOCbEKsAEsZyoC8KRnxHvqQzyAZZUo0Om+qgZlOgrQ
E29PJeCXg5ePKd79j3yFSGpHd9+7Pmf0k3ps2XNCgGTqfnkrXWUzaS65+I0Ywr1Aj9XC6wURScKH
aGe/XbyKNrBGKBeEO2Q/JxJfnDDATHIilJP7g+Eff8OwgofvQppoOBnOpcWJNhDoL1xRjAUP6TaJ
70+w/f3YIW3XC77Ja5z9F+wc3ktdAQ3Jc3zap9IrTCO1q4uTdyUsyrWUonhhFAl0KGBExmBeP84H
sRNY4k+Z571Jw4DwUtYXRV0DDe6vfYDiudN7dNL8pghf9vEL+JvMyw11q2j4h75UbF3hEljzpImG
maCV3qOXsA3Rl6SZxNDkopUtucs+isDf4VD1Q4vqzcFy7UKWl2SxdHqgI/XvCOtwMKCnh2dbu360
m0ZLCVtudtDWaa1QKoqQC5SKzQzTrO8knRmIUDoZt8lGsFZHkvy2YW8GlxDJFN0Gcy3gcgF1OInr
Q/1viP32QnzsfYkTdvJMRh12BmzLQjYOeCVNNo6mpnd8O5Fxdqz23OXqeTfr8Y94il3w9jZbs6bj
u8CF1KbBAw3f4obYhgKZV/yNsoASRsuV1fa7wrBhlxeQmbG88IWq9pN2kJWK23h2ZH6AfQzA6nQJ
06Bi789pRygqI7cKz3Drs/0RQQVbkIuVvpejx0yHjYH2tVQrZqSkb9aFeUX69xbYQUuheRLbsjg+
oHa8v+knGtmPwEf398AZUFlIL3i8kcV2xwuZJhnonENTlBT0Q/wq0FLIJcqCpNLVnu8aGLV/+QZL
EMdoZSlCOl7sh1/aD40rPuL400YkSwf2IUqOudk7BNAWuNdksbK9vCMZmEoaU2WUwzdHL4t89kTA
jOPArxs7261LkTd9aOPOFmXcwpQAKJ/e0+bZrA15AhMlnTZsBdOAicbjXLCAQWdodY925P6qwWxh
4uRrfW3UhIAqTgWFs2tdFxCPBnZsNvV1TLjVSH0VGSD/DYAV95ULLjcyIMuR8rDzTwYdY5tb3VTC
xU8M3C33AlbMLRaLcNBnh15eL8t+d8TKN3Xm/rrpMYR2WlfU5MJk+qxNVU8wQY5D3MQmr1RlyUQf
UNfq+Gdced++rn7xsO/4zyFfBWfALLm//qbvAB5AgCFMpRp92gik/0A59eHSylj+gjBPjgR+mxIK
NGNI8sydn3n7EkXnf0USv04LSpJL/JlWRbIvvGmX73zgf5ZJV4epfWw1D71BN1RGoR37WQVdYAui
seha05fSisRJY5aaC+HKtq6L+Fth8C6pWi0GCbSWlITRpqrbZyltKkSFqeCFdL/v+Dmb/DuhTCuv
3FzWKV0A6EpVlaxhMcVLf5jSNwO9XwyruiotxQXwm2mJFMHm0MEqRFj67QWG3BQz4Shwo80mRSVw
PFlLkjcPvUZo2Z60cftavq1DSPUQLBzkGtknEhO4b7h8G0Hu+nOSclrdQi0O0E5nHv7gaGGCtnW7
EXoQNmXi5fM2NtoZ0XPbMWF77jS40XLCIQkZ9flavxhnAf3wyZf141pWLio7bLYGXysRk1ngXRDt
j2Gn7UNCksStWXDJPl5PQ3VGN87VpJpdsyh33T7c75VltNcYJXH/NsC5bh7CXxGnZ2kW5ZdCABmS
2SymleevdHlDh5XmFUPvIBl+c6cZdkfoxGniBZPtDE1+BzzMgm7L+TNaKnjmoAubZ62pOjfEA42L
ErNUHpg5AEy2Gq8oTTaYX3AKS70D5grT7YXbiDSPe2Y49gptXeUhySkyiLrdH6GWETFq8I+Hrvcf
RUz3aWxYk6gA37H6ztbmDZNV39NCSLoqHNZZVNJLY40hsuHXoJhx6PsS31f1sXDygvm0oSEZkDWG
ZNx+pokMzpAZPVThZgFvKDpiX+9n4SYZ9KwV5pGUo+4Wjigc3M2Pq+uQmqLU3qGOFBSkI7h1AcK3
1pczWrluLHY7MrLUFG4ipLCyzpEMMs294HDEsS46JmYZ5GKq2ufcgtNHh6ms5MVHXapHgKAFqYKw
B3fjEYI/7/gLQ9cEsXnijLle7RifRXY/09WYvchMpNJwT3ZPwePUlU91gsVjX23enrRt1GDIuKmQ
ibICW6iN49g5xT4tUUG8Q/P5aMZnR0plowerz5o7JK0rmzsz0PmmzCFGCsMwiZtofyBNTw46pmkW
PnB76sbzaFmvsNIC464cqYLIOak/Bs17+eGsvWIfFgZ/aPmoNwUs6LgMOlg0KgBumYEC/au0w8Fk
sWue+RlqQUB2FYBeYlL7fp+64c6nnTN6b+qrWKk7zk7zY8dBsqZuj56cwYWdCh2i+TmWdzCrY1eu
gZdKXi8BbhJTjgXDObY6/37ifypRtGJg7CFCtxFyu9birC+MBW+NxGgwo2JfRUuUtqClKDR3dhoD
rSUWoI0HG03CPn0RwYAyq4H+zVnvTsRD3OJuc7O0NcIbbkh0EbNZGYr65OEV/tT5q9YaUdqKdBsX
QzFM293oQfmzdYe89yoxRjwseZSO/PX38Ezx2YJbm+S2b2XCTOO0IziM2N43sZVhfwxtxBeTb/97
vl3nCJbUjR8t5Az167BmEgyMbS9xZPJPm1bvaigtDUlZQImBcg7CtMa8Q9DjZh+2fjk6q0YZhw1K
UE1VgMoUXQr3UXktFPVWH4kiJawsFS5Q5+l6ZUkqyBVEpXwawarxGpF3zabk+6m1In6eqGsVHoJB
2F8WHWvNfnmoyceh+v/DKkK/FfoAV8o7GJUs0EuaLEYt5Qe2Gnue88m3epu0hkTawnMogJsriFN9
zbDvCgGMdjZfiSp0p7dmxujD83LQ5FOE99I+5lDsgy9qNYJiiXDa4dlvhZUE7BJSooQaTldg5bRD
XQQA6t5vXu8LEog5BENLghZ6D+Gvm2knFHdV7LC5pgSrAWWSqf8GQNebBoUfdasL03bRUukUCTQI
sttYRvDJinL3bM2bT5AopWOIvxszalYGQrGlY2KcFPPis3uMiBx1TnQb2sBLg6dv6eH3gqnRD+iI
lDxezL1I/AhqHUo3dT2mkfyhRcWvAX+QoZv63od5DnYcDM5v0M2ESTyQGE5S5U0Css/PPshVBvgW
qmifnvViI+ZfyiNr2Dmste2xL2goYOUXyncJnafMOXUXE8oGBEumxHNuDheEkvnwqjSL0MvSw1rQ
uvNKYhTqUFiM5dZbOREfB1ffOrb7zdWKeFWxu8FePsV0GbX+F5mXEj5UvkXvfmXd+8tCGomG/Nb/
vLwAl8nUZ8k8GoLSYoFw3BPwSe3DEMUc+yldgc7SGEqAfNLzsOBSxdjny+SUF+DGHP3ce2Pw9tNv
jU0SrmtiDwY0yY8X7sxQbWZU7w++xwIsiOVi3U3Y9gkXtcYDYEnPnJGdNTG9nbUgecSSRp6KC0+w
Z+PluNbVJ4JChWJrpb+3P2tTS1ujthKf6p9ANKscYyGlbPulNlgAjqfe/mtGYOHLcq5jImLXhZKd
kDuhQJMYndikLzh+AbDkvDI+RNdm+ildBMW5/Hu7GTT577tySPgsmICWHeiuaZ1S7QB7jRrA9zwF
1PzX92Nkjhx3luGYo+lV7DZGOoxqEQvdxTEyIxdzzbWQeJJ3lgeaJb/xly7SMnYbOY323l5m0jQO
n4mjFZn8T35gvbz7l0lLbPooQ2KJyimnUo1a4UbkJtMyekPWxImQ95KbwqAW4m/h2tG3xfCF/Jpq
45BExS5EpGqPVsEp6AMy3WZCCqzjJ0Qcl17bOPxmSTzQWfv31MWarI1VSm6gweozpRViKRQ9zZxW
qSTNatmMqRmFbvpcSVA51KodmtnpWi142ZYJCbkDeSeuUJ+SEvenk3Ck3kW94N7T/hmclGmPukd6
CQ+RBplEQFgwGQBt0REIk8p2XDICpl4CAWvYCjVHZGDm6YnZ5teLrQuSbz0J7vs/QTd8+XC/VHZD
A5RM1X05SDY7BGqk2PSMB9H/makf1qXeLR735K5BSuqBwJWTZmtj5w6GniqdePAw62LKpVREqWyv
QSOfuSldeo6/0jy9hUqV/AGOz6bVERqQPAsQ/RKpCoEbEAg73zvi47hdblA/TBVBuCZoo8kwTEZX
ZutKFLAdcuXwo+FTFyCduTBc2AiwVyDMwzThdg5eqv4QgsulVqnQ1PYwP7YeoubhviqXZnwNA2BB
JSj7a/SIRTfIA1KMo41dUQbb7a9zHJDbXVWsJhJrGAYfOU1X5mdXosBqF/nBG8g0WNn/Kx26sqvC
CQdsMyOLjmRwE8a1P2a1oUeIy8fdn4qA+rcI8UjvWSY9HfQkC/4pUF9hhO4L7hOF2uQQVdsysnEq
q9nG0g54JP7tPYBW0GKVL6dRCwi7dV9wjJ9hgNd8oHw0ORAizrH37N+LF1GpeGwgn7wzxUTwKH7Y
oeDe4+EEo8e+YIL50cIMup/UC7gqIQd6X1KVdJSmHIF0bMHUV3d7r6baQf7wcgjjZ+rzzadPc8IN
ilu627ExOmuGB1JgSYQP/HSgwz4oYVPy8z87lWg+s1bOrZ42gp/a06NC7iQ0OnF2RxMirFS0PMmA
jaldvpymBj/EondRb1eR+pKjzEEvhhHwZJK9vqw8CFKofCCVozINs9xWLcEi3/j+Aos/dPhVXZ7F
PRC5Ieuz9MhVpFL6dIdPJ3O7DnsUxgh7I2SQfkYU23VWSqGXSH/a/fnFsx9JtsNEcel71HY7XyBu
wGr9ClKkdbfSnU09Ox0YBsPXRReGKFg1NtPXrwq/LjCwgQMHzm9p338mUhhLcW+NSVXEUhY9o1O5
QHqJb+m65QT/TltmlPouE3CP/HQ1jWKTPbaXETGylz2bfIZOuBpxbNUn3BZFsFvWV1pAjnIOxm5H
Bcz+WnLfxu0ZpO14KpljEdgn8WCrwcB/S+caQRlqQQ9VUBJF5uq/5VU3w+C8+jRHxGI1oIyvmizO
vLrT84HoFYBiEED3W6l7oYbBWQla1xeyWyfRYK3AuLPB/ZSI6EdPUFSf5WnOwu/t4ImOgE7tiBqR
RXNjjJZ8r9XTMUw+/sQkcN8aXKDsyOE8xk8TnRuRTwFYH/YusCs+4kiYMriuAr1BfBI0aJBQZQM9
NIViMwLmMYs09Du+eKH0lqNUySnZBdO5XVIGHzrI2iJJ418oqnF9Mc7+VxntK/cHfOUYdZXo1GGf
hC1DDUUWzQPL2+xEXWdYLcbKK20oodFlgWJ14s7a/ml3vyOj09cmjlV/wwx3nrpQGN8hOUolDyi+
tFWRqUHsZTTxkDVRRfi4ICn+GHBkFyqiGsX/iRdMm5VVjZZcRKkkTsgqsgxe3xlQMfFqHoLt2U6p
N9k7bM/V5KjoKvKfS7ls6NNH/sITAZiVROrQmv11hhwu7PdgPQXg9dp33Z2GFbUK6XWx1QdJh4Iw
uDNuOggvf41P+rHq+iW3ItFosJNJesB6Nozza8HgWDM4qgr+Oi5x89Xu/19n+wcr5onQfwn50twU
QIKIPeNjXtdvGpcahQHDPcSXYpL4sMCdPP3RHJunAwqRQnfiFEbtHpaUpx6TlW6j2MM+oIXWQJxl
grBmzw5JZlh9WcGpYMcl64b6OX5BptShIgjR9PiDxGwaoS6ehrl1LflWwdZXy2fN0v8jIfljddHy
1rnrMiNcVwx0eYaVj5AqzqVqq8q8daaay+uajxfLdwIaOw035C7YtkA1naAj+4XQm+G9s48XSzo5
e2IpqCmOMDL6sQxCyp9Ei3PYI07mka67ICigZzoIL/ZdHvzEUmdfAimV6+3WkNumb7ycE42izQSu
ItPc+qMrviqs4gvfZqyyrXYGjUJreWKQIR554hap4wZdezB6RDnezyuAr7pfYei50b+qD4+ViPfi
dFKLyBdnFdfsWmFAclJE7sFlSxln7dTkUogER7F4OGAa8qVO2WR4eLIcwNBOn+Najm9WIjsI7wBd
V05xob2Bzlse6ecllR0EmlCDne+Hcvk3dSKtwtm2t5sWR4gKmtsL+OVigYESWzIKuDki+IBXckJF
EtSb1GRxmUDek2CAT3ol2njLGwleJ1Q5SILhCUHCuC4UetZd9g+3srNnJXABVNYG1brd51/TXgUx
FGSYmbe3YzlL7LVkFtx7+NN0uKvjC+aA8LXdr+Bm1kC6Vh0UwSjn/8TcCULLnZL2s0ZgMwSac4yf
9jsMhimQVfXopIqvKjQRacvogiBpMCGV0IOo/nWzmoCm5AKkYpTgUo3alyml4zVrBfDSYgYNwP6b
BjD0pnbwsFE+bXwVrBxQDEoaSQwQ3zYxa3nM2Tq/aY6zTovAhoCmN2b6XBBd+9vCRJaqplJlyU86
equV1HeJ3C2NBVuqVZAONnXKcriokHXs4qZP6SxYK6pqUkW9ZQxahiDb9co7j8Bdc5UYvurE9xLb
H8HNcYsAK4LpN+wDZOMd7bo0ua2ainUaLGQ/JwuQhMefK2hxtxpwhJz7oMCVZmHPY483F/mrVBxN
aLxM9AQBm7yd/lwlTT5vGk9gAQ1ylTjPC8YhHlA7DidDVhtbSjJQCZMY5siPxJeEVnLeIsMlR16l
My1mLGUbKLnWxWzb7OQLlT0P3d1BxPQvNN1v2VcMAMn6FXS8X5Lb81ymVc///vpZLf3wWWkQAba2
jDbrkkD8XHMN7Q+mYb96kNBlP+bsdIOE1gZop4ozfvlYgd8ZcayQTA8OHUkI5P/Y3zep7qsS/Gn+
VmabPiHtWW0GPelyK1wXNCjkripre3Bnq57mYhXIqnXYSbv2WmlViQPfTgSUbGE6ZbeLyXBxi4Bq
p3RhZ+Z0CWOVvaXRWKu+N0sTZS31RBbbGhZMCunNrUL00nI2/pu3qV0S6eIKcvN5KN+7C8+GEk25
7wBWqRdPVtNCjFgNCNcYa+gLE9y23TqydFRHX0v+Z+GKTR2Ji9YhPHuj/n4FCgr0UIanh2LD21U2
f9bESAyZ9BF3j5ZDYIsb4OePW2zdm9HUgMphkVJ+hzAESWRxRR2t7MZ3Y5is5pzGLtOULAAoY+F6
n8eET9bqMLsuGT8XmyZ1J+J/yLKfFMs2UsXpNBTEwbmVOpQzzwalnRpOYDjFIFHRttDGrTnUmKPW
AdDUzey8fk4oK2wGCzl1o4mNp5nKx5k9SgZMu5Kwl+hcKyVVa9V1dAvUjG2G9zZQEjc9uwhYtRDW
YVIM7F2g8A88+kFkDMqHH8jHcOzYq0BokR78jB5vA3Tam+n91PvciinKC6tBy7QVjlSB3IcYuvXi
0zTKEAPDib1Se6kthxBJ9Aaku0SCmZe2FLfJdLeQYc6TqWMIJEoRcSOoxtvS+GIPXjgB/GIbiUA9
DmAke5KXdNgqEY7NcJdPRi45X8vr8/zF67DWfpdcGOqk1rsTYA+NlyOKdLMDxoU3yzznEIas3+NX
ZH+Ze1Hi/jrmKHf58CD+b10LnYDr6/VRs8cP5Y5TnRkrPtJi/RjifUiVfB3sPHl272FEli86A7iF
dUWm+RVpbrNZ/GL0UWJdjINXH0WGQzYdvk2G/vi7XMDq0e3enkfer882ykAe+yCxMmk4xM7LuT0v
IfqAXxGP6kIABEkDTUce561nohosfoAJNOmEnAO1A3+r0iVq7tu5Obk7Q3PElC3/6yJ9bVotEvm5
v7Ct5KWsSGVtOdFEGVyVdKVrRY2MDc6GJEMPNEIBowZeiwZCY1J1lRm8kebBPJ2dsDePcfJlySxh
/1ZY+eUZbuWKcj85XsmKXtDHahgemXS30aFiNzxWAo+6R10J+Jc0AtDSNg5meFnJ1xS4bsuOVkzd
A+vcxm0/y4S7G0JMaAihJ0F+fO2wMvN9PcSYov5HaNjqiHz95p4k53lFdWsmAbs/1uITsbZj6hlT
h8gW+L0HiiHlIDwa/2Yo87Xe14QlAJUjyF4vRkXaIp2vyz1DMOaiEy7OMRwKxN2pqtxR3qLjNfEo
nJtAPLeah5PkFP7tAjKjzBKFH6gLylxu8fHgEl2h1Uk2HeqKPO+CHwEI8Um6zbgRDp4Q7duZB+0y
/rz/4arIdXR2WwJyrPACvzDRkpwinviORMY/Plyx3rXXy+4uCLhAqGDiX2jnDXwCz1hZQx3R4oad
wZ2H+Rb8pLlk23UwybYFipk9xipf0HhIQG5sA0i81rSFQh219X2PnhDkSDoJbAnmkxVXuyd3f8QB
jm46bDNEqsm13cvn3CgSzwu+2f4eM722AJXinf9J7FWgTRVAcBVja1/oYeR1g1TeLrhFoAC9gzW/
z5I+0Ue2PNAEU9aI22GzHqq3cGtmENYenWihIz+HI2ff1HYWoJ0OmFyl9yuiRKVH/puotS4DIHLN
vSIRrxXgmm5ULVBxWKGtDSGfApVaxZoW00nyJL0RHqE4cNe/Ii46K+94r90qCftdWIzz2mrfpgJm
FAYuQzyRX6BeDQizrZGemx6pjutbxfihgXm7v9LSK7PjfzvPDdgWTlCVglD99fHRHbqeX86V/3zB
q4iAUu0FGAyA07G/4ZMFUJbSX6Mq4v5L+h3icty6yfbqPpFaWwAVj9/6sTgbHliSYJDLHyVWrcFF
Vg8MVAv0ujaUlLGtWhCCO20HNfUNOXdKRl2AVzyAUNggaoEAiKbJWNkXhYPy2o4Fu2KhK2Crl+zF
qlOQegunai3b4u7pRqX8X/M0p2a6h83LV1w64hgoSUFSTLixOW3W6jVSRWTo+t8PCqLnBwYlhNls
YXZTHgfJbCVRX1myCS8X6inUs0NZXYiBu82CmHwq4jvwSQ2atZqGvIbSJKL7WsRzTUMHUStEA5Mk
wf0g8zUs83xNRSplevzUe+OGiku3f0k0Dcl06vDJP7KBO20GCmxA6qr81XCAlIK2K2TKxY8r6gkQ
XMDE5KUYZdlGwuLi8z9J8gPRCU62apqEyoaPS8Oyr3tgjYJBJLfl7FtfvKthOW/uqcFV6y7qdP8L
71Lle8qW4BcBOPHxKKazxc87EL8kIVSR01Taq5Zzu8PY8LWbPii6oxCvBYBjiKH8FiYAA2GCpwuX
ycqecNVmEszndmDgldZ1/b1kFi4UhW7bO27KMzqdmlbUWrqSDpTVjLP2Ow6OVzGi1BQiY+MTcOT+
hP85EtYfpSaERqc0KSKg/VNplYxY9ldjN2kUpSenqK7EHrPJNe/MS/+5E8A5vErwtejKhXob0UIY
kf4/mmdTcQYLotxW5NCJbc4qGgv8/btbFO3NZ5x8XbBeLkKVUhODdSas32kZmUEWLxr18hr0GFAM
ESpCzEnOZ2L7zoqalrr6YOXXk9VXyOWo10lb8En6KB8ukeq8r69N/+fG1fRAVbzIyRdnnssgjiWR
wNA/0S50Lh4TE0ee3TU5JVlUHrhBgo5oKnIOtdTJc8vRDdAQlIgBjNhq1qmUPpGwz3vqWHJA/G3a
Lv99MjizEE0hVbt0JmOb5Av/JdOO86FeDBb9ABfRvqGVodQSKhv4F59WBfxWfMEKLUjOBcvx9tbs
jFs9R8tGvwD5DVI4lWPqSBw900g5as6ssmjDr+ETrk+/mpyYOfM980iGkdw2jvkBe5mLQAZaoqfJ
cEFm7cmBDymFDkMq6oD2C4WvGv4+GdAYdQVW7BOKc5SwyhenYNgRSwJg8SR5y0s3S0/prmfCNbuf
CrpvAOPSDt7KCdUnaYSbNN+JgD24to3jnwE/NLYRSLUEwXi3HKxuzijNpkhkJN4OT8v+v/B++UHQ
VfUORjQ5bi5x13E73ytdP3MW/f8txuQqOeBpbMNDVHeOjNkwUFVDzCPE2g+ywpuUpLO6H8WgvXfC
8gOmyJctvzYWWUIQuMv5JzlYeW3HCnmaXk/Onl6GSbq1+eOA/7lDn1FWGHriin/L8NbdP4UEvwBS
cgwP3jqaR/MAnc35qp6IIPACEJIEF5+IM+auYNrl/OJw1aiTIgtgpevIjLKixkPFJmuNV1MXr5uk
9tXiRiIM67Djr9e8zT5sW4qbjUm2LphE+Rp9OT4NnDVcMU7rzRDYAdpldy492c0Zkri4r8gTeWbp
CDaoLWDcArenSoF0OPccPeQWHVJoJAafe8cX2lp7sLjYsmD42Khb52LsmdQK/Qi+utFCHR4CJ2uj
sIs8GZN1qcbYIFpr6NNnzrMnyhlZfl999uViueUlD/wMzruSZCsa80TcQRcGQtxFOjI9baL5XmOZ
PCL2WDft9A0veZnKdEVwU7J+R1ZafbX5+0HUC7zh49f4AT4UNb3kNJQI3tqzZDST4DicxmaXXvzt
KPhEGN94qbDZb8uM03MgfrIuJj7vCwX6RR7F0XPxFB/IatFoLQrRiV3eTmiQkXP9vBc36qPO3TDQ
4vfjJ3zdtD3m36eZeQMCM8Y9bMZLF1TyLdc04qoiaLPW1mPQT3a3QmQX3QfO+brlf9EC5X35xmzm
wF4OGxkM7hT2+B6tofOyh7GLLAMQbzaromXmXgELIDHzJYtOKokxUOX+ed74cj91eoW2J8/7SJEK
z0qsmx5tUH6qNWooqMTDq004NLiDoonKO/OsJTN0o0i7xeDw2wTYI171J50TvsXWGnAq5IafO9N7
sHOi3/6ysAZCFFG2xA7miDOXUdfXSPhsiPi2S5Z/vFnwG6YvDy1U/+Gal4qcNfsZaglviwIpvz61
k57j2NzcjlXnskssBkGiRzCvpWyfhN5Oybe5hxniUTIVlTqwjoes2okzUxZNPn4bLgzTceR+YzmK
eokTqTaJgqLQYqMAihb4hC/Y6+KTXZI6ORXx5pqQyf7eQ2vDCrAuKLN0LSUGRFgytufD4+4jDpMa
NOIzKQ8tChtRul2gK0OYqIIcvZHfaUIe2ZxcB7uVH2aZj6NkXp5Ho3Sqf7rdH0F4UmHSMCTgpoZt
D0nFiHxoO+m8egFHUq7HEU09NdyN70ZMiIvoaDe7gPgV98dvXw7gP7hn0Ak6htP3eJYuGbTkk/hw
VmPB4lpt8K64HnJP6APxPhsyvDRFdR6/Mtdr7OWYB3XpWrDAjc1gFWxF8gOwJJcpoNkG4xkMGLQC
aTOTrE/WywdwgnUM/Yz8V3BVQ2N0IyXvTFcccifDmfZ2/50guQASWc0NYNMfMk+8QiMi6Vyeev9S
i5ltOxtY/aDQP70Ue4TujtaOnZUVwgh2sBRCEx3lPSLuxfQ7mrP4NJRIJPV8krmIL4oORfmcH964
5Z33jcArdJCsfq172HVmQYaJvGAmjsYH0mNFPb18u3OvMrNsHOW0vT8z9f+OikonG36VeJBkFaDK
tFoE8DR9uwjqZL8mL+V/jZYN2+CmPCB70LpTCoTZp+13GL2E2plu8Bt0p6cEiAqM1IVRNkZzYNV6
IFRot7M5sjBCslU4ahop04MtQX9gOgX2zLZmfG8DAhE8D2R6EDXbUM4Z6g7okCTxV35chPSXI8yh
0zhGnkNfH4FDRTUcqz6VjOQMZcH0s+rpEUBhiAu34NjpHMSChrHGeGgwEcr5nw2JTxGS/46Cpuas
U5a+hvwmtMWeIByFZeujWWxANdqUhieXdk2PiDl5Lj2oHiBrnqKYXc/K3iqB9FGLQT9DP0Eg8pgf
jqmqveQKRvno5KmGuP4jXewbkrtv4f9tdHrpEBIevaq86GsBLwcdxo7SQ5YO8Kb3XSeH7TOa5hhQ
SVgDeVTcei+j9UCEMxyb1lDlUyDgBJ/2nWV6DdqO9TzJid6/X96rj0iGu4FBes1TNOeh5chezgJo
NSx6pYZjzVGe+fQj8FKQLBPpI+fTWPlKsPbliSIW6o+uz0ElwmqVxsYrpp5+9dOEosuLvdOlEqAo
VVqtFM7x6JvxPrR+TIOT6nQ2nxuN7IHzsHoiUc3XSxiLze+m8CVvG/YfjNQ6IZy0tkzdW4gARnbz
lOg1wrTk2ZR30+PBRtkJgACvmXdmmv55oDfR4sz5YzNs+kMSxVunZ8chV19v135eAGwyaQY4ldm7
uBvQUAihcM+qyDiDvbzt/gQ52EP9k2vMJd1+LiAfASTSKUTmwKw8F8Fo9AkBN1oG8XEr2oTOAXdw
PFv0sE46nzaDOLCoAC/XO9V2Vj6sV/p9L8mWQ0bYD/hEKd9OkA+Lnd4vOWRiBRtqoG1ipD8pSRns
ceaBzW+CqmXpx6vZZHEYsm+bPj7Ipl0njZu4wNuvKiNRtbmyqcJVXsue95Aibv0ieURDr40TjfmN
r8yDpVjGxDqdR8ZHVq/hRZoUVxJlk+BQi+fskCqPL5nJRdoFgBnYX/RaSmMqG1SIhqViLE/FJB2t
/+JV1wymm1BG3CfUiTgQvBaBnJdwmVBR9mpfAv46rB6liDNlqwf2GnyauEMxZMR3i/b3nRKEhd1B
RRccdn4EjA3IQdl1VClOdFb+Ygz3zOxiRI3wJ4DnnLtg116Pz957frQbu7/iaxFMGQiQPy/CeZRI
13LX/3xh54J93oSdCqb4+wyJmZBEeQjEB/twsXPQIPzvNwGgQSPYvxZhefqabtkoeNYxHmR9lHUm
jWL0/KQayfFBOrTW/b7uQ3wsUOyEghlszAZDS/Ya1QuC+8K4OvslmNmiBTUG+AlHbyvSGTEWyXP+
3cSfOy/aaTcToW2FXYUtZt2rD7OZkBQ4/UylirYWRkAkj4E1s3AlSZSvMypFD3EKESrLL/b+3v4K
4o8akXZdTwmgDPGiqTwDbWbUhsm5SJVtOJsy7+piWX3lJqwP7ilK/H3leGwNVPr1jefxzTYNT8Mn
hGk0pAUMbF29gUI7jBeSFA4dwRTKr6ipjAeHpGP5Y3B7v7iYOBjykL/xaXGluAYhbTLZSWXicBLy
JjjTh8ofVCRsxIg2U2B4T63JOUmMvK0WTWdvNCiRL+HhNtqtzNekekPzXL3QqR8fjimxyBsgZg+G
amu/lhLcLbQ5K8VU21rtpumaCMaQAHVQEF7JcOgaVYAS4e5KjiMEffLznr4/sRhqyKRNp2oi9FGI
m1elu/cPqAKVbXKOeWmuuXBz8wp6VRl3w1frEe7EVajBc8KYGO5r6S4s9ny1TOjg2TQzpyAfCJky
C7ZaPsR3et4XHh/7nh1wpZLgFXnMiqEVwJIdfrApkTZdmRl9Ple8NoPeJtZcafxs/sMDBTpjGu5o
HssMGZJZ61UVtGBRMd8KE+WXW8Qoqblu9T/PCJfrD9CJpqAaPoh7iMI/zB7Ofwhp14GnzCqcDqJo
F/y7v0Gig4hYKDjVL4mgpKvSpVt+nnvi7VMZIewB7wzcPx/+VaXuFdQleMi7YWVPbyMVQnXrJHpW
oZlzeg5YDh/3cvs52XyY0qIyfQKpoSfIrWCNxU7Am2oGRbc56ZQc1++6Dt1LjTZJxW30MJrJlOwe
fL9s5WHJ/8B1ey9CfNnqEMIkEc5mkX1Y/ckwLraVjA8XmU4qTJtm2/OIK6WN1MIfmPT5WS2Vxe9f
iJaP4KxCTLLcWaARa8OefUmKtmfoaGRxhyHoUJsITt6IkJWJ+EAGyuYF3ELCDhYO6/SvUK8TBCYK
sokX6kNrwDzWEYOawQY9gDzOixD5HBIvID6YiwdlxoyXh+ZOdthOXzC4d4eMdvyNSpJpIE0OSiRi
dkO3GGena5+l4dnVrNWf4i4jqSje9zjUe3cOELezS3u9/Nn2LPhATFU+dsc4IYo3SSjxWWZlZXN1
LEdQl2VC9dkkBz7XVW/eMH8782uewR5hX69Yazo88Bw377QvxfynEtH+571EY4T+Ni0sEf9Q/xTm
qNni1EPrmnG3kXYuTxNHnLFudvH0tM/PR7KLjeapvhg7Vm2ociEkDYr5jLTC3v9MbvSzmRsN8WSV
eOuIKHyTGHWLoJHV1iPEG7ZSqSfyeUmZjm4ZMfQXsVFzpcqg8zgHf3c7al9i/nsHc7Y4VB82yXME
s4Wvw1swyIDD2GJCLODmNDPSs22rZy6U7pODpy8gCZMCazeXEKnm1VIdV4Fz9LbASiWjskR985BJ
Bwqq8RRzozzjJ1DwWGN/H5q7cK3rA2QQVpk+POvxYGkhtiiawwAmKrcHnxzMyUWbQjPLBM/Og50B
3XTXW+q6nFOh865gRIfpTEGb4he8kmqwanZDURChCRAp2xU2ALriXPoTYP+aIT2HbAkdtwOOVe7+
576oDJIi+xautpLQDJjuD8Jy5msnGmnUdcFwIG2z90fyDCwK++PLc9tEZTE582UmmZ2aljjgYGTY
qBfGAPMrgfaY/3LRiET1fZ/zo4u7Zs12/ThNSOoYRoLA/exRm4KJyUbNQCoL0m4m4Mpsn2wDIjfE
ugYeZ/SjovIX0mpDR4D8jIPu8+X7oDQr6K0caFhdjAC1KtNDY4DQbJIJXSIfsFMN+yi+g/ZrSP55
ND7RhRbXxz26mjIGg/W2asKX0mtlamQRftksdEPkDF5OpMA/SYmMU3kxOmIPNzr/a5rb02qG56ru
heNoJDzUTIGQtBdsTs1WH9Mv6SDayjaPI/i3nRm9PK7BDxhPokp54NvEGHgY8plsLuOsG2aBfpBO
frhcNlDepXbeS4ls5TZlBhkBvU89/LsGSKNGKg3svGVDHMHH/movGwBcCSr1lQnlYgsopcKRV1LS
YKZ4PoywaXy41m2konq0bAf/Kq1jlTA+4Wg4vD19wcoMrVimSrfiyZBlQj0pW/JwMqsBu8oTNFq+
vgW1htFRvzfx/U0KfxMUuGbC15mC3WaBPLnwn8Mnr5VlRGRbcWRnzzv0pURlGroQzZPm5qq/07qJ
7Nh8IS+KUZmJ91/usk0c7+2bahIAj1ccD8XhAYZXmORhNdEH1PFqhA9memeAWjSxq9YswaIecax+
Ukf2FlO8WagjcTCFtvCBJHo9okJy14NX6enorXpBocZrgW1to3a6FMFSQxusSC2YZWqWZkJ8O+bW
JOc5Q6PJZSoCC4w5/oxDZIgs+ZNBnKFcVpmUxHDO3ouMYnaKCjGQkLXI4b6ws9yKNIDCoHiuTMan
LfGeLLK70h5OVwZI/VhVWzWFJPYahvE9noF4fDvDGhhrmVYB6diHyrRExkSvU7adVfpJOWPtlxm2
dr0G4MyJQQEwdN5c8lJzqwInmYOK7s2T62U12buPxkY8xEiEOOYtDSlNJ6AaScgHKod/fl2zdLeH
WLRD5lPPC+hCqN7m+BOSwO0ITrmcXg2rtqslq4CC7xvG251uXxc9kDM+Py2q6WyC+HOpgS19N0XT
IueXD/RBjOeR21pQw15gKaXD/SDKKAFgXVVdbOPaa71UNN1T+yMk6+mzGi+1EHVYIxj9va41H8Ad
VR5zxRIWcSAkugtsxIn51R8ZDC/MqlYF0UlqqkLSmjQgKl5JOc4QcmcNkUgC4+T6YTBPAQeC1Une
j4vP979RVmzjo8oUlINEkhbBbpRtl2xLKNL1ZsRoN+lFZdevEWcLyYElDGkfSQYloRFWiCUuXgFS
AWHd1zcuEr6brb+jvDZquX1c5lTeVsewyXtHJG4KyFAXPUVJbSZBQ4Z9KOjV6oUCxySlCE/7EPCf
5i/ZmB/rNL2dgvi3lqHAPaCBZKP4l14h5Q7xWy/rueU4l7bXh0Ix2vb+AtBk08lqR1UVvcS+cd0G
R6Iz2sY2CGRFt9lV1OzLTH4m4Ua3Ub2HsPhV6Qr5ma/oKyMuVlC3oFjzhOefN9HXfNN/zt+2da4A
twPDDLk5p2aV+AuCLgRqz4UdYSc93f/YwcTNqLxTb+pWzaVQ+FeZHdwh0vPa+gbv5uHIBtE/MMOR
BuB/spQ1UaWUkTU5+/iXQz9PfE52cziUFgeeqz98+C1VsJ2c9Wukz204fNmrVypuDdn3Z9DAw/D+
67tXvlFFZXBt/JMNggqT582r28V9N91GbIiX1eTObaN7iDPd0/8zVJPfXh1fPF/XkBC8qHcWglh0
zqVI90efdohgJ18MY0sHJB8ZOIawwNkxM4quOc9hQFlVUg8qfSWrcw7QFu4ugfrJF/fMMICeWIFN
KlKNHeLV7VqjMD4kizQ+dz/AvMBlcHGuJ1vZHzn/pLfxkVrTO4Arz6qTySAMbTC6BBsAO31HdFBu
gxQsZMvAMDhhjYFhtPTB0jOIpj+ZF0jxFaPiHA+7WdzIMd9dTbK80WQPVUaW5ZUFcSOefpsBWZKg
O3uPN1aWBXrme810mHdgWKoor0ZwYILr7QOIDrcfHnhLizlQJv4h8/y0WyN8OaDZ3vsNopc8kEvT
UOLV3C2B8RVY4UF4fMFmWohuOcfXmP74A2WI+XMic5vO7+9cWdBzyfQagcRV+fgfRLqRCFVWAu+A
EHVkjRgI7StFL76GRVuJglp9LCpxjJYdkBKGYmywDTWqez2Wj1KeC+xHAUuqX1pdB8FqhyDY8qJQ
wbCz0fRwxmYUVUz40iWwMhPMF9nzJM3gZff+u488AHWO8fC6kDQYkh/zyKQ06+TZ2EKIsTpTmuAq
8naje3W/VT3DhPqtEfXBL078mcvE8xMK1zg55+yT8nJDvIAeupofW4IcUVw4OcduNJQIvXa4ctb4
0Ed8yYpHyrPznTWHdK+Kuuu6QYXntFY+qNK97g7OECn9zYYIRoymN3Bhc/FycvIDT8xo37vC5E0A
xa+b/uaeWyn0h05i9zz1qkh9Qa5OkFvcUCHzMNepQAPBlbI+U2Nx3N2nmNaT708jspqFjbHKP2O/
+tEXaxSemxKQv2OUwiheEGfOiRDXexQLaadf2Rbnm9u3u3Tst6xxfMqGKJKvAj/PhmMDv6tEcEl1
fWpG5P/HEruYHoPSZOf+bFvLiANEZCOpQ9TfyzpiKMJdHUBjoFhd2xQwOVudohsmDyAYWsb440rz
sezJ6qPY0AKpv5Fzs8AW5LOt3eb/vLwNQXLZOAMbxNNY5BrCFODdDO+z2gPZiXVKccHDISrODW9D
cQJb2LIG0jLGCQZOkub5ZAhgz9i7JFT8InGELyKggBsuk7TCvMUzaqcDBWw9YF5vYnaTVJ4yT2bb
M9ep8ZVbq6tBca/30hGGz3iMV4HLOzpCVnzIk3veBvIFM18psbEPZG4VO3Ie7nnYCkmnaGiKMeNb
Fvh3ZG5zCeEpl0qD89i6T2qBqqmnN1yApP4n9xu/7iZN7PqurgcTmG99keqjzdLXN24ck5J0ZOuK
VDsj6ceQvqPvlZBFk8bmidL4zh4S/3zK2GxMmMOTkUEL1NTtFHBLBYu4v/9Le+N4fPbtm/XPU0GJ
RcVW0/lQhU9MrbraJsux8wAGRKAT4m+iOxGM/AzDKklcyy19nSmxed0HAjs/IoraVsbfx8GYdrTu
1tRb7p7YNkCPrDjTAM2fgD+awJRP2T/Xdauqr6S3sJZvui2adZslPJnWQAGiZrclpCJJByo61gCE
2QZddH/9Rx/KhgrU6tLAvp1GImt/rH2T7xENf5rK+KfbIizE88baeSuZxZm0qAcVokRqMdlGbSaG
abD0bizD8vfaq9W/Ic1YzSVp06g+cLCg0b3m5Pi0c6x+xFAnZZ7lZJ8/gO+KMt3AB5fsew2wRvYN
qvhSZ7MzBssWuNO9rm+fbFA2eH2DQI75Le2YHTKQLufGBGbd9AUUvHdVhFIdqPg7FzMSrg9AdvXg
ZQhNxrgjTQmvLcfZke87UjrOV2aylYxcZWmO2HKDBK13ki/iPVtHaIYSugCnt8ibq8qODJ1ojmDx
hU29RJoQuKNZTRJqS/+p8lf8LBpNbe9yESYPG0QU7CNBZOdqJkAJ3//dJNpL/SaEj31n4zt5vW9a
/NLTfIONrOzzqIv1Qe4s/dPPO5YcqTF83YAVcBejwteYXsdbCNEIvLP9R1g7sNKQE2Sm9OEDYtaJ
aeeMjVl1FqHe/IL+BVLQmJrQT78at7DSWtVglF9ko11Dpp9PKbgMUEWd1Yv/vP0MjdmusiWDiFo1
4S7mLof2D8K67LzYMtfcG//sgTg+/yWJdq+cxvg1jA53bNfnlVqI9wqY+Y4FDpUYszAy0zTrFAYs
f5r8ZdAB+ryaxgXEZNwsRl6MeQIke/wSmM3pJeheS3AbXDGXEbhsOCtvUZbgM9nNXEPw9+p1eO7/
wcTOMK1syzQeTA9YNboctRTcooi1NvBDf0gY3XXlnzXWTMoEm5uAuG1x6nv5jOBMe9YORI/QkmoX
FvJTbNVT93i1tmdNZ1qNDqC2F23CLJ4S9pW93NxCk5FSefnpyGT+gbQ6F0t5vZLWyNndzZT1lCCq
OdLp+i2ibvTAi6wckdWTymZW4vkVfBw4895YfnEAAnPXLpwek/YuV1v35mcph6N1zt1zfwZoaufT
OZrXqwENAnYqxDbp9P1cF0qPH6v3oRNIGv7DdPZmhKK9fR+P+7pHgIRkeMcCrJroPqEYW49SdEfS
C3o0OoTGk79enGDCuzwwIuuWXhJRyBZ0Nb0Q/tNh574DGb+OKMXYa2hWhUS0mO/j6Opo8gfKF0QY
DUjc4ooobo7g/20cCLGNBtWdS8wH/bmi0/sVSRe4+TpZJol56yATI3f09OfwfNcWqVihRMeJV4XC
050UU3zUIwdNyQg7G0up1H15sPv33w2FrG8Mg/faH/X9snOJ83N/L0OorkCMyEsuX5nfnlxmAcMR
2ZxhVs9ZPxOmrEvBaJ0CZiJBzAy1keYq1p4hn+M2dmtF9LGdiAfu9isjjdi8kxOIFytOa7hcS2+M
WEssmbi71wDU5UHG5grv7FczUTr5NR0TCBmudLsN7QWtPsVsVl1gnfbSs9I8BrBbcjcdeH02Hy4P
JoO4rKsLZ1UZVK3ouHV9m1ws5wPR/b1bmREzaOE05xIMaBAyMQkYTFCaUTFUVeK6fNceToO6l8ou
woqc/o7KJWiitmmV9u2PC1QsqvtegZFyuqOT+kQWegDEbzstZeuIrm0HF9APDusl7czBCoACriq0
UEL/Xu4UcafQtfeKttEC4rbYhHop9d104SsgAw7KPJbKNgmd3Tns29LE5PffQHivuhLvHRgVibJy
ZyScU3WUu+l273uPnJK0thjy0bG/2iCVNwqNRxmx1KvnqWTDwtL4fK7T7qmnur9ULDvrulg8LE/t
1CNlIIZ/3NpJ0qcVXccvFeU0TmPs7mtyvpflyV5oCheL7Rw50xzZqFDcJ4oGmm/19verrQJKz38u
oC6TN10a7d6zaMZTKbFdjhCp2vcUUowJ9W3jcwr5TIzy02u50YnIVdP7Z8nP8oOFWu7R/HKLbmLX
mZGkoidVyc2LmfBmkCTrFtyBfSguDnazYET63ElTsLFioOGgFMv32Zuzx0kt0R34qBiJ1EzQoQc4
Mp9sKwtOn9yBvPZcXs7DdlPwLJvHi7JrCoahOf+uc1q9wXQhUYMY9ZRGw3VIBnX1l5/rcxIB3UwU
b044z5PqKoejC/9tts9tR7g7jo0EIEVYGWMXqHk4GvwdEFwleXGVkhqRzjfAkdA4+nipCtYxvHsc
vP0pO5mll34uAA7jbx9ruzTQ+McwLRFEdr81Xi2xtlbGL10GzasecVz863F3B182q3WbvysjV7lr
R3mblhgTupNPgBz8NM6sloipgS7UhOmONVAoEIXJDb1Lz7H2x29mAFnyXCYcDpET9G6licJ3+MdJ
iagdFvTcgf2OREGFAoC3+WnLAiapPULiUJXLJPZ4zZh+3n20yujzJ2zjmokKkrzC8tiro8nQWE7v
F+aAq7dG4XvUgvRWIpjaoTOYkjKTjzOsAXMylQGHSbJ5jIyyNxn3Airwn5WxWDihtQn3kaVq80Kz
ikx+xw9pjw1NTFo40H25zAJ8IYU0szgAz5CT7u8p12Q+rnz3n7/mxVM27M+Hml1cZmSbWrLjePuH
EGSHqV7REIUCwRpGT4hzsKwXy2Noe115k3uNh0cJyu5Q+ZpA7pdqPhVApdOkUoMx21DqiQjNtLwX
co5g7Hfjwsh5ct0f8JvNM9F0e4/D6UxB2gInU/fovTaQiq/P/dgRn0di9NXa57HBxhLpI18bwoBE
K0OW8hoP/ANYeiQk7wQ+9QzwMQXSROI/0aQLXzIb+2OCi62sY/iNHryWvD4BDqFrixrwbRNT5Ujm
PIZL8wpbv0FTFtqIIvJNPHfPo8OO7s1Sirik8kSaPvoDNGPyXtXW+FTtDtPEmbWhH0eznY6lEz3P
kHsk2fV7tZQQFks7neCa4cC0lQ0kladzSd5r+wxZGVXIGZ4RjsoI7A5+cNzc1T/OLs2pgpLAfg5w
emRpJesds7G2spiJTagOt5sWvPTwQ7HyL2IquNJFEjv9v+Xyayzd3QI9lXUoh4Mv2NFOEh6hU22a
XF9gNtZsTAt3hctMkksTP7hxpweoFYcMIy8JwNBjHvBIFFx5OpLiKmDP6EcupjaQe73B9/1/iY0E
o/Vwg3ZYLHG00OXDc85xTNVaD3BIzPtEJ9794NapLyFeyAosDS1gJOZWt/xvoIc87awRlkLKeMSS
kM84o/Uj5Tio0Zvsc9vwMvnEl+0ATnVLRw5FzSyB/OXaK9ecn5g7JUsslzTKuCMuFNPnCegZ1JmX
EWy2/v20RL8HTCrYd/n78jjGZxCUX5uvKQYORQ8D+2edNQlKr5TFjHqXJB06l48loAjOQOOyq06H
jrjKIsU5FXOAeFRW3s71Kbo5AOithiarcmoy6Ir4mEkdSYkLfgNs8u5k4jlUcQ+SvhkuPHFVbAaF
nFPxQ7O0IhCc9sTnQoekHbhYdcMl2OZxUoNLttTvrI/rSpS6FjnMMBeiuFCCU1FEOHQJYhYFrrm+
5N6NeOMpGp+hLEuTJHJ1lDpgJZkQbtOiw0AQbfQdVik7EGdzbT9MooEFez+4vrjqaMM2LTRWEA1D
qZ18nEU821Ar/nUGlWczFIEqJpB3AeqiFafA19uqDNIiYQGo+fiLv9OnIk5X+t+eJE/KBGd4mG17
QMkySCE/D/aW9FJTvlG4TzP2LFi5B94jKWrrl5xz2XZAl6+ltIf/ACat6bvVYGInDTo2auPZK4dw
PTLwb/j4+VxUL8UA9FvdrqG4zO3SBR39Gw+bER7zoJD+/2U9W/YKII8F2YXlBRFuWljRJ+ypvExM
M81yyH7s7XFILp3JBMGIKxr/jqocWGtVGJnWo/y1M8UphVKrlKThSbHZVU+HyilYnTookUZgaFr1
dmhSnixJww/qLfiTQqfxkNBVmzIwJQcF7M+/Vjjaob3DLmfnZqQ3YWUIT7yIoHQFNlOcchlRHMmm
pZG9WBsdWgQ6voq0nPOnCBPXb4nu3xHGVhG+ZL3GmDnd7ondauXtMMxuSCfjtiNeF80iTaZtzNa/
cf2ulz7gWnR7q8F+h4buGQ636xhuqeWQSiWENCvUHPwH0ZMT20cvuX91UJW0n7g5vX3RM8ceUcR9
9tMcT5jBX3uqlKIpc47idAuQKKy/RSmZqQWm6Z1Wq6e/f7qvqLwx4PjjsDRcHGjPIn9Mml2AQXAM
AzaSlfy30ojlwSTIm0OR6eyrrEMS4vmLVbXfUZHgrKbSUB546h73sxMwEoTTczaMs918Ufgor4F4
NM8TzYdQXzjf2RYGGHHen+eg+UpciurOSYPduJTxGAmnzCDNM2pxiRGZltLMIWEowXFqgNQ6OgeD
o0UlHrRuYhDL7uGt6yWKFlcAGigasSrJBLltQ2K2hWQj3hJL94ZyCF5HxG7iHLDQL6Xi9ywcoFTo
NV0/rcMYyIMTbUQ5EOzMthf08E75+Ywkkdx4/6rNmxgf93KP3qio7A4iFDNacDUyb72UFXzevKR1
LxD5YlBPd/OO6kOQgpzdpb696h/e4l4Ec9+4Hi7YrFrbghsdNXHVgdo+l/IiZsjl2lc6tnn3TtcE
MIaCwHzDR+uKo7ZOumUh82wOEnvM4Z5ooRO58wVgpU6K3MveqkWZWSh/2WaiklIHIfw2SUiP/b3T
4saRQMvtcoCMZFCtZiMIgCGdRzfcF7MalXBULkFmg+DZpunkLrOG9QbsroQdIgQXvcQAREN4Pl9k
BI1CsPJKWtLcd+pU3h9ev/v2rGiAeCPomQlxW4jEWhW2UIEjoolNqf1k/vF9OD/x49FhAo9N942u
YLgVRshwIvON0FdxsJzWL1POWzH5qDK8f6rrJQy32PiReA8VaQycDCXYDfz8l5fXirwRzIo94E9i
eFls9dMWBPIFWqRKIR+AFvv1BLroXFlbOEbZxfKgT8lzhVZW7tK6sCvzoVZFCJnkos28eIOor1Mo
jEyOg90Ctz++4qCWlqm51Bwg5jvEVVgABDn6g/xgFl30VF/vhhgJ9rwKb65gP+UPQUgixaTbWSIH
5SPRLood9R7TiObE01SY47wb7pDIyvZgz0KQK0breVwJlUcV+GiK7Apt8FNo2pSNXl07WukCodIG
RmjJw386Auh3oh53fuFBi1HL4M1PpZgIkZ3uT3kEFbFr4o/IfjytblqQU8Vm06HYaWf5P14vFjfP
NdAZ4vyBa72lm027fKFiVwZyi/99MSZ49exWsQa5IVuTdVikxDeiDfl6LfTbJXARy2A2AxwsC0v4
LNIuheNWD3dtNi1vOxZ5CHFb9iYj0aP4nl1yWwP/lpYVJxar87B9zHZ4fD0ccWgO8IisU3Q3Xwbi
bsjppQtXnwCd45lrF1+8a0ETjjs71twf8iu+abUxaojAF6686DnNwcyopRcs5pkCndUT1tV8K9it
7Oulq+9y7hvQ2zbpcrxQhFFkgY8nb/XJGlZqZSvKYMO7g4YCHohdl+SvVjDUlGdJjjks6g/JRYEz
7JuVzTkoa0RLVAegt+WnRA2CFIGEsgeHAdaOuouGMuPmOZpXrAvePSMwWiRgaXt1fmLSUb+9QiBt
5I38YvA3Fr4WDHzxjulIEAIc2pZiIIv0dPczNrNkmFQv9eyyoP+LI8JPjyAgskSsIwqMljcXQk/d
gbli+EhFexCE0KcBsLWhldKrQEuBW5QBOSamcJC7XrHMgpfFU+ATGbRQ5OWC2H+QGYWlc3u3LRz3
XPxypcq5HWMfvxyxpkd6n/84sTwpfTm/ftm5GZDhOnSQ+pR/cAg70I5dctC38JI/9b5GGFjcmi2/
7wkNPxc6Thra8/AvvQ3TsDmtwfEqt5yyKLYL6N3dMf7J/XFHRl2YvOo5lT0RA3xDhsTeEEYvHQC6
8KrNPp3niDwSbMYejMyX7THH6Idz2S8Drs+BvmWRnMJMF6rsrfoPktoklmH0w7ZLAMz6Ia3qUDkW
qwkPr81QnZplMC9xIzdm67FltPFWYV2VBIysxVQ4nePCMPhd/YoiUhD1i96cX02jXEpBAfHTZgJh
HOROW1qTfu/mb32OBlrsyD9fFVTmqNyzQolts2SClSEAVj23D5+Q6Qebiz/WVzyZFn1O2GsaCUvX
4y5FYKcdQQfk8JbFcWYI+vvjw/n7PZYszuDgzjZVzzMwnRlNWHyVARePfbrj0dEiHoDXBVEyHisM
FWtUKIn4H5mGjo7IKjR3qoJ1P/LmxK3ZQuCc0sNETCqVBYV4qo5gfjlsEq8ZlPjKKvvstnMGE6e8
y2FUWiUSFTzbL6m5KxaLM4OrY3s5FStujhmsyeGThYUvlbNogXoMdIPAa8kaeV6RmnCAdo137aS3
LGPxJ/zNky6O1CrrCmDiRKDpPYKJifjuPYSFhOci2w+UVXD739oWwfd6ZwwvxVDigKmkxncLiJ8Y
cT/lFFIJGkJwMDna5THoM+C14qBKpxkpFza2sXj9NgZZCneXfGSXbLZs6Qi2rclHgtaR87EE7SGD
VkOK8jpo+WsIrLkHJwGdl8a2hPovQE9ccOFig+dGCFydTPjXvYaR6z7l3syNxCMR/f7S4WC3n0HG
IBeH3v3HBHSETd0uUUovP6+MMzxWg4lIIcrx+cvXWZE6vslDbUOLUCQOB4PljyuccVb6iRht2OEe
t2C7CY8wWw9sz9ClYC9zyBxnH3HTyCt4ufw26qNyR7VAmCw/o28Fwf41zDTW/TYvBoI23w9BfY90
ESiyeVGX9ip2dwDA0rw3SD/c+8vrgcU3AQr+nIFRL++forPMbS6sEqKZmscZ2qtpVv1I5AJmba1Y
WwgRENRvnIWEkdFrj2XXeK3AbsU+VLTZqrQ7mPpEfnmkFEwTHC5X3dxPSqRFXxEhPIYzPy0hADXm
XoJKxcs9ElmI7G8UTxivxPO7UVpEoZMEd4JF+eMLPOf/YFZC7a2EqS+RWlgLHQdyU2evWTDPzeA7
2K/Mi1FO3Sl+edLsIflv3uYa3xmp9pVe8DWYID2+R6KvMuBDjptS0aYbSGFkfNxB8f5uaScHerxl
m/jejpKWca/6s1t8BpqL0YLq2iGNa0qa8A3XrNKn7u41n+BU5mUazqzM69H89u19G5zg4chpCQdC
Mq/lpww4da8dPxrvkuMKaxoCdlqwDXPWqYQzd29sAOdo75COzH9RrLyaRfa/lXKUHfsE72f/ja78
LbWFIGjSpl4ciwJ1jRpncZDRWB8/q44p/pd4XV0Y5PApuRyPG9taICg4A/z/2P0XTT5CYrjCSt2y
b+dQti3KmRs+Th43AVMdE0dpghbpV0pMDIXw7wZ7YdO84f7jxds3XAYAr1/y/bvefZNjXhx2rgMC
pqqQO1mH65ko/RMGzts2bVs7kfL+2NrhG8mv0Lx+fKZovz+AV/1BPGdFv5MDosrk0xysZ2SkpQKW
FGcd3CGxT+rmIMyYpEBkr2D31MQDM8yH5phorkRQm6Dma4mCtqagJLQOaTlnTviUrKCM16LaJ5DD
bh9IUlLRtewjcSIeGwppn+6QduRjtZRp0+QTqAqW2NP6F1SVptd/VLQ0ktZYxp3HdmDVE/Tlnrc4
PKb/Tla9TM/pLwiy+taXI2syMInRcJ7Qvr0IyhO9hqh9C3LQq8L2QIgwn9FOX24rFHuyzpeh42jF
+37YIlY26A5ctfWbg6i1YXPwdE+tJnAOtOWovaA2ev903pR3rq+DzqdSd34FZmO6yvFzKLjKFhZF
D0TgID7tO5agbI/M3JyBmEMVACJs8mULnQUSWSbiYADKs6PZH+zgalObcZMayiq9RtrfvIbSRh8N
ZnMeqLzbWappMVrDP9OvKMciwPGwJCBWqbPdqYn+0BNRG4rF+p91//+sMyuTj9cz70nTQ6eQ5X9y
MYnHJNxsuH6WU4MTfH/PTBSf5dhMjB+tD4pesRtm5F9nMZcZWycV62/jvAKA6Xwy7AdXxKOTURi7
95qDt8Z2NpeSHRlFNpRV6bvPIJM3aTq1YWa6GqOBlzBxnBUPq7DpFXawyAh0/5v8OGB9LSXwWiCl
NP9qQ0CxtWw3HdHU7uVRquEelh807PvwhbYarUI+uAvhZ0TKm671Qd3jMmKWXn2zAwqUmT7fjIOt
YSyvqYaVSRp3SLneRdATjMBOTnjKjdbkFm56Pibuq18Y/jWYgJcI6EJUL3EcNq6srLSFZAZf4610
QTzDLPzwqyZdCi52wT88JFjYf8kVzxS5VELTIjz3HE4ZM+xCT3GHhFLDmAtpkzop8/9HrBFQWXBw
/F0I7REY6rG8cvv9xvG8YIAG2ub2uHDgQaOktj2k3Qan+fbNs/748ilUrHd1+DAfkBwbIU9BaM4K
rlgju38OGyC4X9CFWjLET0RUDLD/pPBFURBRYqePd1KlRZm5WsVStJAs8x/rM8IM32OOzmk2uzNo
xVESCm3wL5a8W1IlZ4mvZ3e/mV+oni+l8jgpgwYr4zhQ9NuTwip5AJ3LywUXfZsT0fZ8TEkK+RzT
p9qZw+nQRChQy6ujx6ivxHdURjZHWgmx3MBIynYgONzBqLYo5Vfl/uPwX88XjmJXu9gKfya6oIL3
xws6N9wjRG5gCg051kBLRaYZPq03+BuC7eF09ISYfoenDko//9R73jDviKhpmLmzPxxPk5PJyUGA
B+6gQ5ZFEkj+TGUuIvcW0UILSHUYjY/mpbzpwrJ5BQWB8LoTAXrZFKpY1lpUfZZRgAyuKGiiAeYB
bnHxbHxDSF/8F4+ab4WG3UljqR9mwhcsQnfw7TeprOhmXgVH1X7BulQiDcrsvachvXi9Wzfm2ajG
ylyTd6sroEdxfZu8kunLcyXtziDLIQ5F3TPDNUpe43JfTrTWwNa5mHPY1+Mrzs4F8HUFfpT3vH3f
LIiU/mZSxILCjZ98iYSyEEsthsVyN3xXMczfqejBS4LrxqS3iYZSPkYoXCF2VqN2lWWFBUd50ZIC
2bJlSpOqOYtHkaqms6IyG8qcn67fyK/4gZbpQtRVoJV5Ebl9t4m7kQZQ8WadJQsUjsi4wrkhEL9V
PIseFb665Licba/AxcYlC2qjqoTB6RBpJTO1AWpTHuEkqEnE/FUkN9h5X23OeVvvjCx51WU2Lwqe
Sc3nxdn+ebx4iKtu9Bvk4r+PF7Aw1n86EYDFCx0dAhBxfG1xIYketWMScVfoW/swSsxm+VD9moib
BlsWmSVHFzWB71l1ouZR1Ltrua3ct6uoSOcMn7kp84ctzrkSwqrDpQJxk0kDrscEbYb5NR5ZB58g
lwFMOg+CdiclKFBg016YYdMuHCvOhvHdnNR+OWrPW12w09bw9gdMZpap616U+94Zm2LKcxqE8I0i
uyD7WWsEL9RxXVtebVIjEzv+bVm8Svf5doCO5cUSF0DjwvwmJTrbLmmRwGP14Hn1IMAmP+iVAvPU
fWPQWr+aZeYgoyfD4DIClYGJl26UVptd5TYEusjILf88VFhLvWkBiXt7sCIpU6hA6HEWFqhzzmYP
UaY/zRzhRU3E6Owqm8GyAmVkTTKk5JlRvSjD75lM5/Gfo5HJlK/2wdp/j+PWehsC/2abJFf8cRqX
eQ4vNLMpIz7bO4Z7cf+Mx60wc+Tb4fxz23oHrk6ud9laErPWlS7y+RsayZemiSeVMTd+//TZhRod
YEZoKP5fTu2bfIICjedWYsqzG0j4IauxKyIkgTTuR+G1V+D8I4VffIG9LLweXKM+WPwljv0tItqH
ghTNyr42ixdbyJ2ImoNuJgc32VwgACl6YFAQ1JRtR/Qx7wIZPS2w7XPW9dOKRwva8yBrEbdf9VId
yueigDLxJZCv6+OZc7KdTI0anl4YeHYa9+pOIg38ibYOE8u2DTXjyZ5FccvzGhgTlx3WOtbd0MiI
PYXT37ToHjBpjUdSfKoTK40t/OwMlbosNK9g9WnVPwBkgGoUlZvlm5sBp1UZVEIfgF+NAvyXJ8h+
sA5aWGiztj9SlM/Fol2KYAc/JLHSxTPjbDVKT4+mJNoYtUnkNIf2RGnp1WNuugnRLgf3hoE+HCJS
eLh5pmZR407Qb8HRJnfsanwP2PvkHsURdI/mis4iCHab09rh505VyIheM0gIK+v+LXANSp66pfgU
8FZ4pAt9U+zegK1TASNCpJ/7uURLKvgQ7/mcFH1kVJcQi5Cl369yDEbIIWqkAtMISVAI5p7ADeJ6
JxPf//vPCLDnWFmmzZPPnIh1dy+MrRq/VvBSjubDZ6n6tLqEMtdh7JxuTeuzF7aGOfJMovamMaoQ
LyMkh7FhAdD+3UMIE3WPmIFhbZBxsF9mnAbyI/rlgSu2iMfpQMC6VNs1TOXL4FvAv4nRPZoIpXGW
IYY+G00Cho7d+3bsHWeI2L9WJnEbsCrcwlCtWwJbTuPI7dcwg79AHF72yrz9yCVjKI83QrEOJ8ZI
DlPtwFNUeNTmnEZXI+9xBBYVAYlJ0nq8eC9itcxJKcydoD83MJTOMEAaxGA3NKNlt7Qqyxv5jmIl
kI/Qzj+Etq/mm/q3GB54+uITEgDtQuqfbJ5b+201dvEMzVTx+e4rrbai+aQ9FOWIg0ZjQ7wbhGIV
bPkDZb7yNTKf7GegIjtgfag3NgOhmfl5c422VnVAhxxgAgOFP+v7xeaAvP6gAYQsF+G+t0dF9D4Q
dyif1uHS+9iC/iFSjBhaImEC2pKficnlMpZ+1CpqwZVw26r24vMYVptZ9bIsDl/47cy2M9UtXcNf
oPk0VbEjndfMm9az21ZdZRy/eoe3uB32UgEBRXf98PKFUHtPKeXgXp10h2bBTeBtkuILvgQKsjQ7
IQBUAB3QHkvNF4cYZCluezNBJANnFekZYkxYC1tkCSylBDoq0En2AOUUCnm3MydU5qx79I2t/gNE
a1QYWD12QnX6nQ8MDFzHy8vkJXfNoI83YN7hXNRY9LYSbbSiIVKDKJjR+wq4OJVCgcEapA8f1KJo
l08nZwOhTmkr9NcOi2xJZqIUx+vSuPoRj7BhsY+qqcOi0P2RSd0mEQNybWSdpulMBdKra5aMPShR
vTM/JcT6NK1Kd+IFa5fW7TktPwOzN89QN0RdnlOhESabM5urxyTui/LXTo7x7+aXmsSJzRfF3pAJ
2s6KhQpjLmXIl7RjxE6PG/yvaj3V8KnuDX7USBlH2X3dtJHpXHiIb7hL+g97SXQo+Gtok29hnEKj
dfX2lyfaiLS3+53C7lU/OZNcMEmokjfKcyS/0sQyaPHvctGGirFYMPWi8MUF1uziZxvB7ybReR9d
r1Bl1OUJuy3xqN7nfwnLMXMKvGgAXO8dtIbb3kBWlV845QKf5XHc6f99tre93zKSFa9lKRMidemM
LglG7it8WXK855F458BZIofJ01V/Y7oZ9Hxlh6cmwoyReD86VJX4gg8h3WQboe0Kh8YW+UAZ6TX2
fIK++BCUQ9n5acmeMFQJ6VJS5/PKhSkvMQtVou7iX/L9qJv2d/cHGIMy87LvFYwW9CURg6Qloyz8
GV71b6G/1cKXcvTVFYrlEtjN7jmTMFnlUYQpdM36uLUW+YbUT4LaOcIKlqGkPRmYr+ChI8wuuLaA
DseYsdPzPg9oAg0p4ELPeqIpTSCzx8flJl1k9UyvvKApgu0sjrdEx6oTiv1/BIn2Lgnc+cy6XKzu
r8CtVrWj+TslwIwjjBF2Hzuv3OXc4hG5wgthYYNkxCV3NkPdYlc+NwmWe/K6er0j+0Grazs8L5KY
hWjKP28VNmiFEkC6mZRqQQPbCykluJyBZYynmpFFajOUTRcRtsYqeAMniHwUerbCqMK6n1DcE5MT
WHBAnYI4NNKkhcunt+eXjNQFgJjEVTb0njZa3K/T7RiFArZffqB3sAeJW4OLOOoBYeK0c+gKaQka
brxVJAyqv2OWWTAtypSe5HmA4qk80ybrpgtBkcrCbssrtGQySYt8nVOtSpkAzM7j6UH24Jat/CvJ
ned6+iH+4HjjWPmnDh67AzqzsPbu4mJRLptUVqQEK1hNmDiLz9lodw4A3Gio0oEMikWnDZyeDndx
QIgHGsPQzU+uR/xWwmFe1oWt4kES62je6jFSC1k13y5v7+pJH/GGqO1XJ/SAAhUj6rtJD6WTmzk8
04zHHq618+xa19JT5L/ukg4GsPY2UqWgbbT1N/FRxMUSAzCeTDgqek3o8YiEKWHNhfG9oWfxkyTs
4xKHZ8lJ8+7g5fLuCFdlfy8arUmgFDr1GBD7+YQeglFd3GRKA7tw9E5lkkk36DnSBSyQFYQ7GMos
BdnP1rU+WYVsaPS1ctWCGLQNsc7WbMTwje6Td9h7wXBXZQQFXsvQFg+TgWXaye/PIriTF97HMt2B
M4k2DbqpBsUyorp90pHGtXNV3I5ea2fmnWzCcg05OxnAeURKA/87hL05RPfkN3Av4uci+8Kz4pYc
VkkmtenpMW3bfnylXeUmNeU2+5GAZt+c1TcpWT1v13FPuYoNOe2KAfA1dkA9WOTB7hEdhnvqA+xM
WCOBVeCalNQ8IKb6dk384HCcoknSvODhy204CpwYbxAEEm4J4RUBZ8f5g/RNAgeP6UFJnhmFc/9F
L5ggwCfV99gHBSD/JQNrzgi/PAcYVRQ1HU+GAhwG9AgpZjN7iyCXmdHBvdcnYgRU0HejliAueu7z
u9Fib0JuQG5YAtoTGUJq2UT89x9uvFb3y5kw9c4DWl+TgQKatFWAziVbqm/+cE+lJ1pdo7cp+9fj
gjpiGQOJ4qFTNaDVQZrAZd2GgAfwnTyJdA7dunIfqwkZw7vmS7C1cXlH/LSjCbyiqrnqwgrSUy+a
f49q8w72rAmLZ3kXBLlBAiX7pv7orVFMhYNNzNJiiuUa7oR/8MaHwh5nL2QBOhKtSTD+lAMvKyYk
r6gpW78VWo5xgLifvIPRZ+//eNvbIZT+FpvJD9/85JWv2vVe1lL+RL4mXlL0pPtXbUqNH46LSu9c
Cs8lWvIJrZERGPqX6YLYpXcPLoBXBGhOfJgrt/gt7L4UhpdEKMXXSfTcDllSwasC4hqm6cqK+oKe
ueJqbaDkUp2utJB5U0Oa0AXaeZwhkreW8+9yPN65pb0xb5oCiaqwKvb5KwCvqO8fY0T2YXxQYBmb
pIkSGFbiz/1WMheGsyuGap/xJPG+QCRJJG1RPtxTewAdoNQEGEnSAaiQNZXqoXAS7Fp/cFbacqwX
JkBIZC7DyixQ8qu79RNI49M5sNec5XIf8SLRDAf+JfzQSyJxq4IbVX+R4C/TDODD8IGfD+yUltbI
m07GY6ULPa2T890tHA0S3HJ9Sr0jt1I4c23oZF2lntfRVlHppyNYvLt2iQd5b6uvwMKUB/BegVNx
cpckZP7vicxo3CNXP2CJ1G3o+dpzSq9qv2lkDn8Sxl5XlufHcIjBChbyo+fmQkSXgS/YqMUaOL0z
vXOto/yXWh6Ayjp+4C+NnZiTQBKisAsdhlgtE5ehwkUuKJs48lUGMXZnN1Unvoe6CoR0D7mfnhvb
W86GFrHfp/DUgoSQZwdj/iVRQ3NAheulM7BbI4IqzZM2VBA5eorsCzBOVrBjyiRIdQV//SGGgOUa
i8bswYz9CgzvSs4YmyRvrBFtzClvVT4KJybdeXApNp8P9C7qHcOM+d3vlhmjEX+E861mGh71RdKi
BdXQvIhL3FkCX+3BrxvlqebFsUN9z5+fMSfdfwK1pCK5LWw83OqO7OHvDZB45qRiwbg4yPf4xsgJ
gpZ++wcZWiKSIDXh/QPD4t3c1PmHqqQg4Qpuk3RixU4BMxY193lwmCGa36OIC8BWYfYz6vysf1Mk
4cDrARFzshhiSRZZbR8zcHA71fIAkcbsJvkSzvHF6Fdof2+6JmaCF2H4QQl83x5o0OuhskKgi8X5
AJrJpIhXz4r9zEfw3FHm2732dRSLwMXEHCxu1HOegNs/o5itSulqIiVqih5c2tkRmzD8zSsE/A1s
7XI5c0DYhN2XZbI4HZH2iBKIfqJLJDz/YnjtqxOYGFORf792LZO9fx7sdBZqpT1bZbE0TyMSbXC8
LpWGlLk53M1BTdDqfd7Ziz6rmPQ/Obzg1j6iMjwGaz06cXBatdUW8nuJg7+CGUFNof7GqxPlPhFS
XrUNShWAIqNpS9lIWl6GdLvDUPx3halWV2RJUK5QYZE1s63M/DNtsatjXkwCD/telcDVrzbYFZV7
oz9zm4lMlsZfjQ11IoKOrrKUKMOijFlg/h0ZzDVBPCuSaLWZ/QaHSrQ2sDZV8cFDwnZqPhxLw1xu
h7ei5DCoLFRCproKoqRPqhGvRErHVEJbjNBBaReYmyh2AG1LuPFaO8qgWVrAm1WFuQfxomh07yLx
1VdgzL0BkFFCfbXo9bBWBfdtNZO6KGm9cWDp7XRSW3UWgieYof+LlY1Xuwg8+hymf5/9q1pHGRv0
I9+xi6+yxlNQSBC2UTvfm0olNEjHt/LuUjt7eYcTBfVtx+4u3fs0NEJ+FE8S2lNLXiiG0GSHGgHh
5bt8j+QJssviO6/UWLhP+fwWkZFBvtNSGv77RC8FMHyUXvrisy5K/kaefccy+hzM+rnsqa6jGd4e
qZaTTR6dd/gwG16RKdLbNxXIkgsyJYh3FL3QRRThv695Sr8y4kguTBw70RfHylAwrChp1oIhC3ts
vXwJtX3qv3zE9pRXrsgSMh5HCM2zD/ojFYqkiF57Bh/Kpt2JUthj7emKA28UWb5uX/PcS/XlRdhH
SwiInE01JDOemZCIgITbLu7Ksj/91yyUkBUjUXxOYrMCfcPpSiz8uh8t44M+jz21DlTEYJd1cyM5
cg2LIOs2yXDFGSTGyQHb5XPtzX+l5gWnKj1S5mSdGJqSW5kg9o95KPoqSx17RgMwingRBrs0Gkss
bpSifPgtvz6H/6dz+zQmONVNQE3gY28q81lp1AdHburVFq4GIGqjLnjJltW6BXJI78weOAHBZxDL
+GAwyPJRV7SicTJxHPZDauUjPVOkKnQuZai5hlUuigq3qZEp66EkAs6Wmcy3nXBA7LnGvuhEPFH1
fZLfJPg5HPnkb5AQaeeJtiwyWcKk0ziQs0moq/E2aKKDS7gHIHjpVQDdSUjoJeg8Y6c5QF5/KJz6
aMm4iwiwT2fhkf44E5kq69nx4skpYijLxZKkegZphj/G1FDhUCSlO/R+GRBvKRwfFwsC8iVdV8zR
XlwLBc9x1uGvFDMsM7Y0yCSHb6KcoH7dUaG0P8H7N6Y4ayokO0uGrR894CUCTSsPR9rb55vyVHjs
6BPzuMT/RjQRChDBNVjx9wnAkHYp2+bOeIIevGsc/yRMFkh4KzPB1QIB2au+amau0tscfQxGnLBS
Iezm6bIZeACVnym1dv1uSZMMEr+jgYZswRBZxIVFzfMK6pySRInCCGBl9b1SxSzvrjxYYwMuFnu4
OvVYGodCqiZTjI++DLNXj+EpI+VreaRrRY8IWglxGuw5ezon8AiPVKISNpPRRp/B/7YU/dVXYdAD
bSSIwkcpMddyv3ygGv54phnbRpRvVi9OKXAMgnnW4VfRzJNagLJZ7+nyF1Cz84fFqWXZU+m7aUhK
g+ayKZocG5VukbdJ7SF7qHDqAup+aV9j2cZYp0vBvU20YXwFDuv46AdQPd0dihkrK4+hbSBnS+ox
r6gmdI9XZ6LlUVIUjD4IGWERhli5GRu2GgjRNGOhIt3TvrvxfQTJyQoEeScN4rIqC+N2wGBwhV2k
GY+pu9BjHQ3Jq0PWD2vUxdYdBaIMPG40a4xF5ryCntK4asHjuPnXuDuXOLLLgPVxF9cmwqaWflza
482mUbqxtII3Cu1mLJv4Ne3c8mysGEomixh/mDdpT/RDYFf53irSsVah4WRdO9UA3ykBNAJ78FAT
LvsgbvSWjC/zyxcbz/ygS/Pko1i/9Rnj58O50hkzqzDndMPWnDbxILs07f1SrSqO6Jqjpx0KxNaI
BjxjXfvTWDQea+UQtiiTeFCNhPCH6nv+WZII6zAD/S/cnLJu/T+sCl/fAKZN4qAnt6oXBBhjKNvm
FPQz24qikhOEFz/NDdO57Q/wkLKkK3kAvj/tW9Q+F0dVlzHojN57gZCedCyh7YfSGDLq//a1MbA3
70SMIp27MCC1xGsOBuCGGWWqz5m2QS0FhcWC/A1BqUeJt2v6gibM3UHX4XkAJX/BqIAx3V9I1a31
+HGssp0E3F8/dUOwXBRQl4VzRkOfF7CuYiKehKOknW89McWbdpVCg4GrZLOzf0lwpicr4R+kSIq/
7Y4X8U8eHwQI91OvwLpqGi+xvcEv+cLipo0xnZMkj6KWTWhdPQlY0tjAEssnPjpb2VctrL2jaRJI
Kl1Hl9MTTxaQbtBG+Xe3qBfKEuznCFw5aPVTNowfs8dgXcZlJJAv9loijGW6vqo4hwd/LjLG4qB3
SswZve3u8mUI4wMKF0dIbAZ95q2NEsGfFE9RpeBi8Do30LtyQm7DFritXGrNaR49FSiJmtOhJKtY
A1Lb1sd48xv6GCwUeEF2/7IdHwJNjbQ93SSW6fBkFfCO8MZciqrK5wYuF06cF3ahX/qeFUdlIws3
UoduHJrrI11DtOmMRaNQTC9tE4l6Tzr51Y0uM6a5FY+o+nFRA5rdaIwD9h2KhicJ/Hbqz3Cr4VZh
3kjJgMcaFSRLbpf8h+n4Pu8TjFk7O3Icv0qVgItraWQ1ofwuVnzRblQnZb9Mk9MiV6dKX3S8e8y7
o+0IYVDt5Bdtfkcs1D+Jh0VkxRbVepSryl6nj9V/JbsmbzZrccdCbPyXXTWSq8Bbw7zmdxRJVgfK
VJEdVcW776YPq+pmyH+5sKDM25tfAJTpiOEbGisf0CIyZPhhOFvP8r+Zw8a5qpsyftR5m1g4dzX8
HJuAAINCxfe0PHAkC6QurCThr1KRBnVyh3bpIirgqWmsNeLghGvA3wu85TTn9qTim82cgV9gjVXm
byCFy0CqR6sUiSrquas8XoNTYptznCqIWARiuMKg8Yjz/mTQriwGMZ0CpoVNdR2laX0Bl4Czy8gb
Q2cRy95zz00i3WrC5RmUq5jG8pvIzNDHSvdwXJRUUrC9GENSvzk3rIdTA9EET+qvDJW3MrHyZDVD
84ldetz5H1NEXLwPUcOyn0k/79/8xEqemxw047wmUrcRSB2R0PNbGF5jI5dYwnrCKGg33b1NNh2Y
9bvhqMh0BWR6nFI8LI9IyW3vMFRh4ansFBFDASteKVkgBPiTs5fCjnMN0IHtKTtIkmPsDttPzMyT
8Jm277FrZwdWbQsoqMUsARDakMzQhpwr9m5oTL9j2aLFuwdAggUigZqIG9CBnptSKuaeZIMFdP7L
PIgXOKL2YdyoUBL5dxhSehoeOXSmpVTgxEallrnYGhKljecHnQ7Yr+MIsUxpTvgSptb3pzZ0yfv8
XC/jL/MavC8jRSbr9uNJgotMJYKtp4Mcc99C8a9WmVAjNO1XdXUjmT0ACQvCAPjNwXMBr5UYUFuz
mxswVELtHbZVoawAJqXlgsTMFdfIpM16jjjqp9eJjsJLBwz6SQwvgtMM8dJs3jM5lO+P6K8o9g02
IVE2OBmnBf15JAYLsEHalyOiTvr8aj45NW4AlMwxoCTqxrm0Ffdw1YB/3cASRVIqvUhNiXOEkufg
/zdrL+qTbr/E7mwZLlF17SU8q9jtDKUYCDdipK+Qa9YDh7FL3XK5iuTmY8+Ps97sEjgHHuudZGpe
4GHMz2MJsVMArr9tAstN0zoidgJOTniOXwfllRLBqYoH0SJnxHtuMuPYywgtSE2wCAAoYjyZRTSd
iikCBQWBfyvDR41T55goQTy5WLWt9YxMoi/lQCKtIiDdS1lv3Opf3ESGPMDKNGRBgVuqgOw3Q37+
w0//VCYpOGd8SNT0gyYA+dFbJNUak5V0zJm9ZNd1cih6lTrAb9bC84Hyi+67QVI9D58oaHaxrL8z
lHHuyMMwRb+W1Govx0WDvDPUx7YFopB6R1RHGvechFmv0vZeKbpAQ6gJbxUT14VNVuOV+8HPMYg6
C+iTOr3rvwKxmo2xTgblcINDGfypxTdMhStEcJkJ/d0NQjYR1r8U8Q/bjZC7UfOwz7BjoIDiDh2A
IjljPHH+Fmsi+L9xsjZr8EFDtc0sO346B+ERJMhd2x8jcCmuhIary2clmd2W5o12QNqz9A657Wq+
Psrxefu+GkzAdYyFz7M4zl+QE9QIQwmJB8oftDvCbEUtIQcxL1cjWIHnZ6yLUMsVOUZnRiranqhD
5reddRxhcn42WCH2VGaEH0FPM153u2lDXFE+nFrDU6CY1xFQI8mIbYSnq2JhmdIMuQ5wuMV0QRWn
2FYDj0jW93GY/CQYVPFgT6/UAGYOFefqu5BoRXVeyyMIJ7SWx+juS++8Z27br1AX57nqskHbf6BY
/7WWEGtJHYtdvJCLtWOGt9PF8Rj/rwoYlpXeihUPLXioas1Zm1EgUUzx5hrn5PimENMdRoGIPuZC
XoLFJXUCBoIl3b3MYS7hUsogS2pKFrFhrvhMLuAHO43ogWFoDwOE3krApHj5GEsvSmIJEU8NnZ0K
oMUl29oZpG/nSB20Pujhr6JbEoCpu4vTUGG1rnK2EaZfkRyHxo7MTwWxQPuott5ciDIMkYkAy1bo
KHdvr/Cr0ernRhRfkrWPATW9u3sbs/4sNNTz0QWojLVCc+DBJOCSBhbeb7XzHKWC9i1h5sGkzqiT
mzii9H+qb0MycMgIksuSdMK0em8YJQuqDar1K7N+RT4W6O/LkTChGxN1vJ8dVYKaRAMXNbD07r4d
ESia7zlg4txjiFr+HEEHm2BxNS7j/2Q/HXXbVMPTK1+1LRpGqUjIVgtEPCH+wzM4DFSEIRvVF4Pd
GPYRMnrFfRc5qH5VCaKcvFqJIQ605/TwEBtEJP9u/06WCoUCWccfFE/oOFs2q61qViMO2vJeLsOA
yVq2KWschbuxR14zwBoFL4JitlZgK+LsCWS4Ehfy54gCLfjxcyKmsoy6P4X7ftNg86tSShtwh3F1
ky4s4HAUKO3pn49YyL+A8kPQf63dD8/dfxT2CFS4sPT4H3//ivtFiBu/zi+EUcyZQMZbQpzYDp/8
2O/9rRlreP/NF4rxCs9kNeU32iMGwdP7zu7n91JdiXnfNN7ayRdVG4ZI5Zoo+ylIkF8JdtAypmUs
0FehjaAk1eVDsyeHUSvub3bM1kZX11hEwVhAsQ1hQxUdCzAGt+mFH3U0G3zNB5BdsTaeDcv0mGEv
rpM9yrGxPOteyhGLlNBGfqxiyUyxXeJtUbGiyq3W7t2gxq4Kr+PBQf3MUQq42+mtDRchf9ymtcvQ
OzNrocn7f7ZhFwP2twOf6ROxeb6GfAbFFupXIGf6LtW02UHHDzBwtujFmTnHOPcVVEfkyExu6B0Y
3bxl7IYq87R/ufLYIdcXEVxwEkXCOsbNAK8RfJgpaEwzIN/Db58VmjhYLo8/K3rb7DXY5kRYf380
IIVmBAW2WVTzHlmYR49lDbjl48QYf5XtR5Fl489HZlMivPurtAhsRLBYVEB/2gKYHyP7dqc1iFHF
rHsg2eQ0NEuKhQyZf48oV0FosEBiaUORxHMz2Qb+xRN4CxLOsTpf+VNcmzpZMTDw8HnMAHnBhpuk
RoR52ppGobX+FZTmZ1c6zsn+S/93pxGu4zXVeFeQbCqfJXChy7PNAzV2InzN3zf5HnXEvM58E1MR
Bpg2T7Pu8ZJLlwxU1+34SArgPVuFGkdGYWMRqfwfHVbdx1UZRsVz8qurGob/SecM+zPDOR5pB70E
zLISR33bfb2SP0DYSp90Lz4VNNVJBDFWqxa1y9ww/BqGG8juNWxXRKV9Y9KFS2fcDfjvSoFAnqET
f5vJn2QOIyvnmRFMvp0dmQy/RGf5PCrPPwm8dc0fAOhaXimahoPDRegQkhzeYMRw7n25BGwskExl
dxxkV9I6jnh1xaauodpT5ZrJ5qv0yvSOvV7gqqOCu2gWtBBiGmzsqBNW6NWWsI3jdvQKR8jPvOQi
qTf0o0OAuU3fTchbFn44vMOBYrQJoR724uOki3fJiBuUvDmovD1WN3ZEXCo3AHLpZ7tYhDGbTqHj
H08BpbTXBl1NiiRg6EYw2WyaCZ6lwuvFY6jrGa/jMMQLoKQH3kZS0pwsjBdChPiMxilhsd97a2JT
OGaXVRUocbOQhBJMqM9/Hr1jjBnqxsPxRT1zldYBHYNbSaDpLlq1LMS+cTp92OJorglaaLIXzXoW
m6uCmrSJgiWXKWQslAmuGtEx04T26jIlCvAsYnE80BczcAJN24J7Je3fnWob+bVlZtpOeQQRMD7x
w+0b+jDnhnD9NZQjDvNM+Fj2YCIzB0sYNu46noZTpZVeigEdw3TVkEIwmOu7SDUFqn1uRmM51HCW
YTULotd7aYrBmKnQTVQgwb31aQCAaYdBRg1dOXIoAJXH6RScsgSIkf7n5NKHtRaBShGJvre5VmUh
zC5wY89lJU+uM8r5kLjtIsuuZDjk5tR/PZK198eSc4ipNKWrLT9mRTNzVyq81QUJt6TC3gxxg2iE
pJZ77bb1DVpjeiUlIG9mXJxqGeOdTQqL5630mVhw+u4CSHyxWjFXo38s3a+M0Mircc2EjMOhvUEj
h6K2+U0dsSguMV1cgt4e9g1RlJwcH9t+rWeY1Jrt0Ig2dVHFHBP1nNYNaPIHCQrXAUoNDq6+ZBQz
OAnTO7yzjDUHM1jBmFaioDuhCM8SNB4sNxUhu+1sVTT+OK3Brd+Y9FFRezPRcmeazKFhuocFIvhT
WwSOUPzToS76m+vKfn0Ez6Qlp8mk+qRH96g3eDjtkrIrOK6yFDZj39kWq7EpOQe+EBNPVEs0/uyr
EIS1+fhnNIZ//YiJA2AM8/kXJCf5DsSxO1b1NXqot4Hr7ufM9IfoQVDY1w6vV3BjRr0k+EU2gvFO
lRC7znsGqCr32iwbscVwe9uAbIX1FFeOiM4aEZ+ZF4ZUlGQbEMInYVVOoH2YnEf9I3Tkgld3yRy7
LuQDDsKaMyDmza/Pgjod0mV8QNqHykDNHIpccFJFi+TwcRtBBBtQWNQjdGxluWueQaKwxCKSoTmP
CQt3P1lel7N2xgBPJt8gIZuhPEH7MXPgasb5XFN6qpXs5K2H3UP4ScHIrbIrFJguG7HDLzKxm/Yl
rpr9qyTQiZnwDYPzSS3hm9sNGgiqPo+keTsAUKwYIVwvYIcACig+78BR0mhGPmCClr6fjrzadWO7
XIpPT1pULmTS9PG2IJPuX46fVtMBQn2Gu9xd3b9vQHMWT/a29xnPJHAKDoWR80giJGNyY/MRxEyP
TAyMhwm3iOu+TGH2wvVVHddkE3kCJ/px4b4HKKdZ+ph5BytmvSnkxpuqAL5clzmEF2ORNubAMUdz
yoaVIUZLCh+zxdtVKfFyz2EukfjJNGbelaiUdI3emGJR9UTh2Wl771oVciii+ED8tg2yYI0rQNbl
gNGdWzIAieHMFxWa3DdKBoqXzkvTXf94FWENAvQwQldnofSsulVljYVov5mk5hsr2LUSvlu0Z+gX
D8kjxNoIwU9X72Xw74MQWxqCd29zQdSmf6HBEhc4a2OG7pDDWETpXrV49wEfjMe97MIJA4nHF4PB
Q6X32lNkEa2F6zyRhVU6aEPXqBVYlCiaWcjw1cD8QythsgxDBOKnyiCU9cBOSQxP66XlEcpvkHYF
+KlC8cr4O7kheuIhng4o/cfzvpxsW3bP+oTLrIyT8lP+9fAo0kxLmFBDQe12/jx9a42HvgPja+54
wwSUpPWgrukmgeedJNJYmfDpcSXyqKrLpJo9lPfka/79dXYNv/rMWEBw3eiLASzs+rnDf668ZFki
a6PUcD9EAff100abUD6xE6LHqY2dN3F7mIp0YMccIRG0+rhqJrIHnYRb8D4up8DpV/6kS3LiIsvn
cxTP4nMYYoKzougVSxsfrQP98zHGi+c3+oOVKctV7c1huyGpIfshqKNZk5IakftZlK2LEFykW2hY
ZsHMPaSy21k/8D+B3VnIDTlvjvBGwbXCr01kZqaIpEiUXPl5t5x7rW1Ybaz2vhABNv9+E/9DmKz9
i90Fql3w352CGJ5D6TNq8i9/do5041wPpSbzY0EGZi6auiVAAyr/opzlpOmXKEmoMV/7gymhv79X
g6zC69sevKNJVW710L7VrIbIacVT1aB0KpfQlHKHgCV+WC4TY6BWN9pei/xNaKUE+paG4aZhsshs
Oc57nhmAIJBAnBtreb+L0XOFau/tw5YyRoHY73H0r/BThNrx3xuWrWxPFMNqlHCt8PThalXG5QoZ
UGsAUtQK6naorpp/BRnbZNyDeaSs7Z0kK56RE3lmZYlbHBBX85SJLya3S5rOdH90A21RFN3EX7Sd
OA/NWQl1BML8HIKGSuhPZrZbMRF2T9ZvjfOiSx7BR27ExninRkZPVHRtQt5A+2u8FrZvhAVaDCJv
t3BrY+IpXoXBVXFB80MD3f4bjmEiKgRU0sFmAYgi2ovOaGgI+AHjRtxR2+tukfKJPGAyxH/DIyjB
eI6IWfLcGu2e8XqDJTbb1ZhukjY+uOeJ4qr7Vb/APj9mdIBeSDOB1kyY6Wlq0+I+AhiMIHhhgvl2
KxKnMz8xLOaJcpnn1sopy0K9jhL84BgTYv0XkHjt48XWR9S5QGmn+KLS4gpRdZdl8zxY1tbj4/26
1OqCyDAd747G/ovtv5OH6bV0PG1TAjlbre0ZTGu0OfXvI4mM+ZH7OMsuLFB/LOECiXxGGC/IjN3o
KbZ+m4WVgfVfvuENzOZ2D4ru02WXVCkltWgBN8cakDQLyvuOzvEYnwZULn47tMTuywsfZUpiLT4x
Uo/Eh3qqd0e0owsPt0KniVarmFs1pj/jkIXWYw81y6Yl0avcWgjxuiUMz5PB/BGhI594xFR/Gy7v
9Cz974jEsN+feHvl93F58DhkMkYduIoV+RO8V46IjQdEsZGWSR/ITZwjXR9wzDFkbXo1/WSHdEo2
U/bdYdClml0ngpSEsT5KPA/QD0zVNli7+YlJfHMdC0BG2eGJ5xrmR+lV9vHDUA5anHX+Gw2cb+uZ
fIMQfoZMkYTdjKCKCqzpsloN+L27vZJq8gFUJ/iaNd5Y3mF06DEwXAQ/PNjKhOsoAJVXE3rAgwhs
XszGsX+rux+sIRGtZHli8bH2GEJJZOamQ/NiXUXIAUZCoA62yTjmxawXEDuGU2pd2+gzlQOPyM69
8Wop0UVnJIrqckuSxEWj8rpRTHwxtuMwv7laVYgPCfnl3VTz0fF+CHJlxyeblTfoZ3NSVcsHdXnN
VMLWYABHzAppRwugs0zVTnxnrezydmjquMjKPXKtVUU9x4iUCseOY6s8cnh4ntFqnHT2mLQCxJXt
MjYA8ThGw5cOmCgOpcvWFAYzoV0PWtKk73gned87A0qoxrdrOfmfoQjjvuEKoHBBAXZW1UHjn8Jx
OLjA2Xi6cV9R6dtmkMsKyzBCTWy3Tyl8IfSRinOl+ma4VhWGg1lD5OqFojzSx95RIoTjnGZqNB9p
MUi1unWCCu0k9UW1qdA4V3vIht/1k+2y4vtcrhQwC2bvvtqNboSny3bk8O9y+OaFJbUoHYodtvQ8
1vRcFGX/4s8QCVc841+H9hhGXFDde9yEShQf0kDToVDuhrzdjz0Mx1YjQ4JdZLNQRUR33tLhEcTt
GZWJCWg3fxkiQbv7/TsecmyAxKqdZ7QC5EFfyXAfgTKghEHHtByQCRrfIy9d9vgwXsTgS+5kRx4T
NxnG9PWE6oJMexhE+pGjm1kHyHr67zpeviIxbUWzMhPFlckHivwFPW2/Pb3775e3+taqxYJ635zj
+PoPW7VY+UQ+w5JRgmxs8tVWJXIt3T/gDpjLgnJmzq9rbFRROzu/m+OfbHE+c6FsYb8A5evh6fkm
u50aPY6yz2924dsRLSAmyeQCzsbQeoCjzu+X4Z16Xw2bSS+Dy6Adzp7HWX+87em4bZ1BiBJrc4MW
z9lUwBJi00RDuCdmJ4GqqyhttvC9/aKA039V1DOIkrE80E/BNH+LjT5Vp1stHoOHd1tcrj4hqLBq
awtmqygMhtuqdqpnK3QiJkfUvex0gv5D6sfBT63/UmBfByRVDSWilH+QW4a0iAPGcDh00csnpoe2
7qsNMdiWmD6jNW/jHSisd/1HIwIhoY6Ia6Ncz460XJQMaqvQ5tqPIoU2L16isOiNaRKlCbJ3GuU8
jvqN55naF3eoSy4PFEtPeAxB0Ca3n8FMm5EO3svNvy4hRNNEX0Lk3MIJCP1zavhYkWwtLb1WQjiQ
KsutPXo1GS0aCGksTAoH1gvHjCBMgGTlmfYaWmcVqrl0V1N8wmLa0ZboXQ9xIkqEk5AM3KsW4YcF
rXS0I7J40fu3SagqqfJLdg51POSEjWHaZhYpHj0OtnMTsym9kiQChTzqaDq5tIOa0Cn0Of1sjUNj
yWbrbRT9rpPiEjFHjOapLfo6xgNqoJwxK5xmTd733rm8l2br9oD1FoP+y4qm6wZhSHHBcWdYKp/5
SenbkcEfF1lcdLTN9N/tj42y/gwVu9YNoOnWCrOWthJNUdH3+7+HvcnGkKegB1wKcQ3v4Ce3xvJH
bxa8izmRwWtNofxTFLMExkPcsTs1BbFpN4xtbUvClInWgxPdueoXDEGCHO4iqRmzD/kA/jLNRtCi
rny1B4D/8BIW5jaHG15rWhao6eFjk7fZVB7LJTLQn/bLvTp8x7my+ONiQ8Q6X+8ktLZWYyZK8AaD
2x/U0wD5hQpLmHYfn1IOPsBcxX2BNIkb+yYwUXTJzI/Qu4dZnbmIHVKjmuhsthl79grFyTJ1aJPy
Ltga022mXLC9bc79lDzDlvOpsEh5BXmelq8SiubrZsSEK91IMPvSJbvyCXtYCxFe9QCVt3FcH4bs
EUrhSLgOV67pQ9giXrKscyYjKP5YSzmZXFiX2lSuRuO0AD8/Fr6vQ1cy4Kk/MnjgPg//ZVmKamVv
sHBahkCesPfUuZqF9/0IuKrbd2I0reKou4asx8fvRA39mPg23XiwpBll+mJl+KZyfOBp57nO9JnY
UHqoNq3FCI4Pd8uhWl5/Wq1G7S/1E+pxZ0uWOi/bjXRf5KLBdwDIzLDL4/qL2jb+C8+uXmwGB41o
eBReUU+8nKxmzaHzTaM1xgxUbqBRtCa/3Fs9P1Ii91rmUPTHjWISaeY6GKBjh+ag28RnIRVeVpZp
+itWApR7nO9q1q48jFfcRT78dmNv+ML+uauq7I933uiOdBQBrL7NVo7wmXMR/oyVdAQpoqcpBYdZ
djdpGjzX6V83cS+FZawfsxa0LdNZyDasCMXHdewhPhlImXVVkYvAFlNDDIlt0CAfaGSnDWcME/hZ
W4a27j9kvOaU34ESFRaUo9xvVbI5DIyBtQ7Y+ECevN/tyTiyLXhg9mgz7GeCBexjZrSf8+23FPal
fmY4JVZTnpZHn6of8bnjJSNvnIg07pcl20V+OCdOZ1zqxDzBHnJC9jO3ln3V2seILiqzWkvflcZV
HoaTi5Sgdl/LgCF1Xc4Ce3Bql4et7DKnqqr0AxPE7CmmA9PwgUOcwtXVploJGL8q2L/012LWs+SL
p6MuyaT8IqPLFK9iWF7JpOMQy/m5LE9lvdFIhEt91ryCfIK2+civudNW2ozc9k+Al8N8YGQKjeu4
TOmn9FWXNyD30B44CYpa4Av+4/26o2FvRQDmG0RkdHCw4g39BQr5dFIoGKnwcoh6MMuxeu2pBY5Y
70MSLV7LNZebuG0ady1xS/irC9RL8wOJdF/ivhvCAgPQVlvHbWNigBHckx6bg+9rj2bh5wcZFAdd
nSCqwW3vkYVHQ7rKoZ8E5prJ+M6NKx8YXhe8Ac8fLEJKY9CsRebG17cCrk8oqe+rejwe/x5RoByb
S27eo4LhAgtPWYiWgAp1W+cr+k4z3qI/V7CTfg7PgNUVznSGuNDCZI56xtpXzAt452vam4/39NYO
nykP/OTDfo4+Tn6kabCQ2XzqzTWAAmW8X2+jOPcnSCfO98YuqFt+m5gjiUqSDKHJR1pG/fPxOtnR
ObczOpNl90bYnSVzVODgJeCJqNUu1Ge4ydOO1a9+kaN22ahB2pl6hDRbGDpLLdmdDqOZka7wemTa
jlqvjh9PluqrWYWP0BkhzlYh9ix6C8XCwyzSSs0bl6kxHSHmqdfq2qY2GibPq652Fgk4FmocI8+T
Eq+/A5lCWxnRx/zu0qFZVWgsHq3moZkBVggqzz1eXvRyu+dXtftzrmO81C+1f504l3ULDHG+XVr/
UdSxTFCLP4n/nVYmGkPMuH0iC8RdpIT899ps0JYELafizAgt24G0nFHSrE1BppLyAkBjieTUkWEm
hilFwJO5kuWlaNI/AuFvNqT8vwpRhoQ4ng/LuAecs5yZlBVr6a8b0sp3BSFh3HOfd3ib5/UBbrgu
shqX0hobfHLQ2BpDZFTMH1GwaX9j5WmyXhekg1Who7r5lQXDf5PcDWobi2hP3Ru/NoUFPRJ+SKHw
jdY/khiOBNV/irLr28PFyGjFn1x1XT0p/N/rWkfhaE632tGfidcHxVB7RVYEmQahZSNAw+I4rPJu
YE0uosWNu4scEzM2HTyiPBHyK6uOj/J6VkqTc+kLW9aBpUlEKaQRt3+ojDcaXvf6xkAfVVCVbAyO
nNUl3YdLiUlHE+ofzBUOTGBnFEVJeOtGLNkHsH1Ggn/VkStoqYqxFHbAr59y8nLQKgxLN/ncWwuL
57YZU3n3VlUq1zfDSnulo098k5c71xksz3xTS9ikPbHOIhEU3tyfA//hSoZxKckB6o0B6owFQ3gk
zhDmmPyVkWFwgZCj0WoJAIxvh1JKLaKWJSDBpDYsP0EEooAegG3b2y11Uarajs0iaFNKG1nzlT5G
K2K3AzWSpfFkiiJ/gHisLWRbd2FTa2dWe5uvPt1CXzc+TGIuXI6RBYKxXTWd9pj9wbk6zyhsJ13Q
qWn1Yds+3Oo/trm9NC+rdIPQYYI/9iZGfyW3u09H2x7Wf83nGmillNTd0gafLJkJel+qaBRsi78L
clMKmj5DwmkS/mT1MN2DOvmi2VmJVuAQ8TqboDGonZQeb8uWioudwit50Ts3em0h5GXb8Y8KLrz0
0TY0WginXi6gte5XoPIqalgDYsAQN37aQBxdDRUIUbh0jVO9gsvpfElmqEP/R9AhCq7N9ar9AVKT
fM12oTQJDmGlrXb0H+WK0lG+RjAyorIhV2uiyY3FG/09vwNnyMTSis1bLtkiZvUPpjF/xvb6FrLY
vXoG3tKuBfIUrhWIKsafuWKWtbQwt4xsz+Vp5xZ+MNBfiNpky3+DX7Y/NXMjEmtDTJBRajbBj+jP
4tm0k0wuqaO6/B21tUxz9fxtn80JQRCxYPlSkUELdxZ5fcag5PjaYDo9f/LfIhmwrcVZHmeHUs48
irSG5h9ziuv8sa+DXJppBnAp5I+TlEAu/gWy3n0HGEiDpUqWr9mRtCl7AOa5ILceTYbh+V7wJVJK
KafKdTDDxdqai68hiDYZ1k4MkyjDvMhoLisclSrK6hCnPz6t00MZeRPj9SDMrdUw9l2/Miec8wPI
PC2mAoxT2ivSDkgKS0R0QVaUWkh8LGjZNHsMcEIijChpOSdMTHAfNvdO231eGFYH9kq1N8+DzA8r
yPY24oxLJgjw6o9pqfc45VWqtt8FkKEronMniDW/BeV9mjH+9L8pQbij8tAV/ImgkMcNADe2jDK6
9SD1Ptl1YobG7IeyLLEVu25v37LOMHBTWR18MH2C7EpzZzw3a3o/zOAvJ28WUzNfEMbUIza9EZT/
72jeuhzZ/HGe4TmKTTXXKJO6VTXTZWyBKzZdYlpKEttUtUVfPQLPI4YYfQSxzQ+aQb7LPPY9XpUj
PpOjuJEaFKE62PyZhmlQYuOYPlEEWdYNPdX6UUEQJRAQ8bs+r2XzyQj6HtfUSbRwukjeGBx6NsQk
1389/PixKOUwiuo57Z7TUHY1ZGfEIwZtN4x2z22gQzoJsT2I/6dUg2mgdh7Pr991MpLKkqiDmAgS
tWG/ViuJE5CHBZPLUG0S6gmwZJlyYF/644CRo+H6wAxn6UHgOe/Z7cgQeziIV0tb4dkwHjuB4KuL
bJq+Zp246JM8YjFEJcdIG6IcyudcPE2GliINTpsnNQDcgYF9vnAJRlFHRt+Mmw7O+bkB5fUVXbfq
sG1E09lUoZa2J0DkIrAeSuv79B4Scs7jc9uZiIoxgtS+QA9Z2oeecFG8f1P09kbzeYNk7vRMl6/P
8K3QKYGnw7M4JP9OX6WeoPWu06pSIoERzG29UuKmcemPSlHl8gN/3de8ylPiwuANyJAGIWkSUZrL
s8F13nEk83SKUXXlqzqMMkHoCf/VNiFM2I/zyy0tRBOVoi4ZWHA2DMmiel4IMiltIUssuDCa0uim
phWKNKUWAXzGf+CDmdvqdTUMKXBrYI1qB36lq75F9D7lEcpPOBBd23QtMLtCBpDlQuWmFd7V2nBi
zU883Z2P9zinNf/vY4UkNey7NwPDiVD+WBNnOc2xJJ43nYjkvsMVDAFjZSfunt/7vKtqbgWC85y6
QfwWayFAwfp0/qoyC23majot9DtLjbDruXIBWR725atwKLPYy0Zlb8rqV/2Tbc1nh2njvtOTqC0B
/3e/lHRRU9CTDN93Ji6btVx4x7UWteqzywPoJDqHJybXBqZtcz9cYZiR/vg5j1fSv35CnPWSVnrw
qgb7PeAkyhFWCCZPdjU4BVx5OlDI7q3nJEyVy7Kwg3wMwc8Yd3UA91JzB+Bz2bFmWqJpxWwE4yEn
VmgPvnqu9EB7ANwj+9v6MvuTRve6kwqaVi4Up3OLvgHiRpBBVrYBtKM/HiOmi2brqqEEYUM+1iU9
rod/xoqXBewOK97C9fovA3E14eYgN6c76P2bUbOY5PeiFlwdSKrwX95ZpaRDCBMH8oYaOFwcUtN8
YE41w94Gps1jMwRk3RRSrB8DcDamva5vuc+bBLUou6IvUmMxQLBJo6g/TbHIomoxoWkd8WS9XcVN
ynjGwfEaZMG3OcTzDZavlBXGb/DC0pzDUSD4QFSpUuXRCVY/fQY2ye6DAI6lsNkBaMuhp9/ygdif
UXfuEWrazfkIItbmMGOjapSMfQiG86fDvGUy3FeVajyJ140Kw01eudu56WP2lpH/ELXoDy7l2QZV
MovuwYrGgrb5dFeLRLh4zYw6b35W70z6ndRc6r7+Nek1IWp/gUYdn7ylqoabnCa5ALshbT+maMHu
AtAjQ4Pa9e5lM5pyRFjgAJzQHX7E5xM8QFE8+vkWUuiMKSYukny9SK2erEfayX9C7l68PW1C3ojw
aM26j+dpCRN0vDGvWgx4FPMXvMUOujY1+c+ya79PX7xE810l379f86em4fhuEHAy7fGtHqPLXBvx
XReH4ANcO1V+Cdzr9zb5YGk1F6JiBKISisJ++72ABUmNO24tFq0jHLLIJiDZlT2GflfC7XiFhfst
X6YpQVYjMugxp4LGle1DTICJZ2t7Xd98AePCtsVHMxjE7TSkoi76n4qFXjTZJVGUcBedC+vPYASJ
zcXrNppLlXftCjQyXkS/3hvcPXPuhpJNRm1p6mE+tHn//TUpGgF1TZbb5BGHpASxrDRbRXuVuto0
3Iprq5W1hdBEKky3s1Pn4xmXsHwsHF3kLO2vBTbMYklRsNktM2Sk89EQCn37LlsbbkIUWiMdT6GI
4ZOO5ugphA9cYXLR+0348K3tdi4tZo+j++gFxCiIe76dWcOwSGjqgsM6msc8IDoqYo1KRrLFVUTg
ZzFTYED7wjb3OrXg8EY/OiyCN+OWXSwzcaDeJTK+7XdhwK/1Zx32Kki8eMbyT7hTII8vemuKF5eO
yiqqrKCHLSQTpl40Rn2bk+AjjAveZwwBPZOFK4rpkrtQ5XbH+HkbItTNu8qNlMMdhRY8/W4vlXci
P7MRl51a3+rAN6XWxgyhQ0ARugNAoQ87+IKARj2I46hshhs+moyoCzyvloQZ5wUXhK1GJSY6LVFr
9s7B4x+m7/JDUNIfZCVoVbddp0xnrvZd1y1s5dvscH03XqRxyDZZ0fRKDpCCB7AxPFpjt0tODI6V
WXnON93W5SPxREG+UjpS3smEvI/kCMcYFz2XF5d8qiHE6LxFt2Kb633txO5rDq+Vw6Fhc7PD
`protect end_protected
