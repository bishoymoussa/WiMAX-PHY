-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
piIYy/6XPGSV0xgE00l3jm+WnsieQWxzpQlrW2Z376mt16W12n/yyy2lWguF865DL9N3P29mqL1G
YzdNpGR5rwd71Y6KjhDLpDryZrmetvwHosN0MHSsQ7GXUJmgKz24eeiH9hWlb9usQ6qT0PbxKKKJ
E3Ip6f3NFii5pWmWcyg3cFjDGA+syy+FvTLJbrgY6Sxn5Ad2cirEk7qn0gPX1fFf2sLrlgJiUOMb
Eu1Uy2kp1wxGb50Io+Ipz2S7Xaambj5N6UIAX+3jv4ZXP1JmYaJNT7Qif/ZXnMlhaGIBth6oixBH
FZGNN/1Y2LuctQlP3lVylPX8jnpZom/bIjdDJg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6208)
`protect data_block
qw0f0wbOQsKAD8S+vHpY2ZSpr8QtWHqL1EQJ6pGrrlw0kgEuUcbNfoBnbOkwDYiFpiW3CoLd0d9Q
fn06GtkdreogTAJHxqJOkl6JCpRgpWqlAx1WpPanzQt/ZZEgqHl/5c0llnMy5qi4MDrSpotOijPd
AMKohY+ls8LVrcPRT59fXfe5gsKQVXTxOoY0WQId2jazU8QOKLk/vnb5Bt+32/PTAhrWkeN2WXzs
AirWiztpgItnBNJYGGv93DoFJCDALEY6uIy8RRjzszYupZWWnaIjGswtESe7c8CX8rpCJZVtyJCW
6SHrMTU4RVza8mHoiGEDt53hizC6RDQzh4Dne7xfu191lK4USOsddVJ9Wp+u746IsNprmiXS/e8s
D4Lv/DmQWuUy/q5fRE/gZ3OHobur09fWXwaOcJ2tqaLl7URto3BamIXmLtlabdGqQaRrf7sgkSd+
qUjLRvf8RyNoPr896pDQdqVblcS4UL3kPAVgQP1XbR214tVMNel6jLueI1bdqFLwZ/+DI7v8vTYE
c70tXNu1uOo5Yh9/pPVXU3yDu7l8PNTTTs0cJKYtW5fBIeG914FI7bq9hTV69up+R1JYmNt5f8SY
sUeiK7ZZ1DziS1i1tUtJTAZhsM6SeJqqVDVLC78ow/AARl3SrQvxBEkFNW2I7p/9flLtCPz8NEc3
OEMkguSmdilqjA4d48JmXul6f1jHV8+Zp3c6cwjKiCeWhp3ISoiqxegrdQlZqCTIic00d6sEdu3M
pR3toNTq3xfS0IJq5Qv79AvVSdltuEuqtGglpjsQii1tfxut+TEKZlxeoqS6oJeE+XKp263foUJ2
MTjFqwJ47tqUkoaw2n6faOmF4KymX4bBqQuOTV9galdpUHzlZpxK4lPUTCy8SU+g7bfS3vaOuYQ9
gA3z+hVrvWy82PndcTWG1ffCwDBqxqlr8gnUOxdlsBg8bnud6qbM1znIZvtfc4jxLfyixM/CD3H/
yt4bAkFL/t51YV+L6QG5U4WoW+SObwvhxPyk8WFnrlqrccULSfeMMGYbJMEO+jFhJM0ZIoFJrB8q
Wca+HoAszm0ha7zoT8RyNYZq3MFeaxWgmSa6WJ1yM5wT4HmFg4eWy9nfrCoArNPVG5liWEWoz+cv
G+QJTtabb/HDzo6If4csd41aYHk4uhmsoVdbNzCnl/XmuAFLuS7ogx5RhckvmHXNVyVyzi954qfA
wN0deFonSR+wOZRo8ju9ilQ3F8H90AzW5d1pB9zZ1KkfX8SGn9H2ZIWDGuQbrvpKHjAOd971ePTb
quJdDZ0+bTtBlDMAZ9P7sgfy03bOlQB1Z5595bujy9DLAuITgEJu7ec0eQqhbgrzISJFq0mmjLqp
5n+QgHN60tzpl5OvhtD6y/B7g6efVjExiDdFrWkfbrgfUPLPXuZW9fkb3kL8AFbSS8iMWPw0N7DK
hjVSAPfzcTmB09xFLW4lgJCqiO+fCVzySg6JDIM5mvgiA9zo3S9gg/s8GIy01zXMJRLSUq1dtykG
KEtxeEg68hrPEFxDwuRn6P8qTYD+gtR0k13B7jqfEKnNKDiv5IVMGw54t8WRNWUBjIw2AEnFGlU6
EgYoH3dR2o4X8FERjESsOufydjElPxr86/n2NXMKEQy8XIOypgRs7GdA7OEH2nz5yDyVYGlAKlul
O+WhDxEIc8hI+D82dZFGsTST/v6u1p+WwV8uPq2Mu6rQpK1iz8Jj0kix3Z2TrREXEADRnHo0FM0s
sQqU9jjhok31yfsC3OfGdwUaP3w4sSlKKgM4OHRiUbQBmSI6L8QrXggrjCQCcX3NIiv6MDV3OwdX
gM4i7M5Q+S/N6BlbqfetG1JBmztUsRWTPpzkf0yELpBZ1DqvPdEZTgz7AfW49JTmg2kSL+AV/X72
tSpSwEgJvLisXD7HzwH9NQRpM1KwZY6fcrtF5dveZF059U3DrY42l5lYoEgGFJBqH6U/SIK1P5wA
x2ZCN83jCOBZzVXZlGJ/OFGjAwEIiafeLEmggin+1M9ABG58nGF2iab3XHxbvTA+En+E3fYZXatN
dvRaple3irNt9L6E6/bQPDtrL5n5oWRV9DzW0kZsZ6VqoPpzqvidiGTSAgllwhaU44F1/4YhBBkr
b3lz6E5KLZTwO0Jki0gPz7SGmgtQycZVsLkfCww81Z2zW3OjOjo6/WXUeY4lc6JeTUG0aWXay2Ne
r7ZiFSZ+BZd7CdcRk4gsSvI8jHNphrESbSnx7B+XH5zWTIaC+j/mHOwXmsA/5KmXzUvZkJSDQq5J
KW50m6QSNSjsMfz3+DRiZ1OOKI+2OHK0Urpbg2Bpsy0u1InluMFkax+2qm8L0tmfL7lJEzc21JSu
ABSHy0kv1MeFTlSzgfNqC6nTRdaTO+TE/apweSv8lhCUpH8yNkfCm3+EhAD9Lm+HSE158eUtaJtI
Bg+WXpvfBQ8gnAHOB1h5/TbOL1Rq1v11vHRlCh4wA254sUWk1wfd3SRleYq+0gyZKo5BqJcWt1+z
86QRwQo7dqSZCKtiijt+oQEnccCIAjPR2p4QESQCVc4CK1SiW4F6eZ8xBWddZd2TYLs0e1YFo1WA
O4X/pnO4Ofc4jNPQKFagKjAHVPggDR3TV/iQEDpfgtqJy92FIDmUSnHMved8Xt9wkJC43yJ+9qk7
xnaRbahW2mvfc5SYdBDS/STupRwh1d1xvrn7WR5ZXFK69YkZEtX+UZuSFBKUg3Bz1R4Dfq1Y9ghr
gmW3Z+GZqtSYbMc2jIWUd6eDu3Lff0uWe1GIot1H8h519qkM4dW/kxfOJM6qF1BLIPoNEQgHVapC
RxTMzDqSoLgzWzwfCRnIov0nWtJ6rYWGV//xBG7yboJxVVXEE8Z8uvb84TH7nfAwrLoIl6gafwtp
t6/SBleCBsgCinwis4+sWcFLli3gzi/NFh2BIBNqyVZhyIEhuR1fevJ1ndGxgVvV7fOrZkykMXK2
oY4DVDBT1hKlPDLrvjEe/mo531xWFge0O+lmkWcY5SWQy7mnZ+rKpXRjROo7JKxpjw1t9lp9hx3c
1bt9Qj96bNgknsWcjlL7vdkRLVRNqwmnGCII/uJt/2EGHwQYcnKSycz7JKEX6FBNjtj7Q8Ce3lxD
cJmsEunCTHQJvG2DGLAtzVBziE/kilYaBvq3gry3VFVfBJFgCHRX1P4NapzqAA9nEW3WJd+OKxwQ
fm1Y7MDAuPcN30sI/SCosdYCDHqvjMtevrsghA/W25zr58R6on4eyUv3CoPcPoYgFe1yaM8jgz9O
RmIH9e1N638ZxXav9sIdRwGTKzccvnJK74Z4+HTym8lfx/CJDYhqSVQ29KUSKw9ncpEg01WCCtZ4
Pi/eiBJGWph8u+BA5sef7R8veYxq9+6YG/q59ogFqpuJC6XmL1JRGBX6v2zLfp50/2ASCdnugQfG
QGZ9/lTBtl5Wix0BEPtEXpcJOhB0VWe+dZ8iizNq8yKsNenrC+7mhsqQvN94j/GtAYif/AMa1nxU
a4+Pb+MZVrlCk5SNXXrRBWEx8/RelpGDcTEAtkfmNWyboos7SQt6M0fG2IGid7VwTIwME0qr7M9/
QQVrizqisvIpUoMahtUQAlGUIUhVJbV4wIEuWgGIlZ+wfatb0rZX5Whh9e3C0MCUigwmnybrnnd7
+rlHUiSBrTtG3UJ3ZTP1Cs+puLsmpuw6aQRGfdsr1KY62KtJzFXp0dFRBRH+Fqk9NJKd2xxWR5a8
6mZzA/HtIKIDy4+v2y4wP5VJAbn9Wt9OufmF55jjmhMskDcV2ML5rAby/nNXTwP5OV7DkUkGSsu7
qMOp6/Il/tJZLoJcc91lqHjv1dE8WbLU236bG52Ve8jyEu4g9aEgy9fe3qQ9SgfjrFl3gC1XU5yA
Eri/QCc36jSRLej3U9+H9aGQieAJ7a7zNI8TUA9+SD1C+ERiqVxkD4mMovb+XT7SP7QJ7HCH0SYZ
wMUqXZOKUlQNdKgP/NYnUOb1ZcM5Nh+T/K/AVT1WstArqA0bbmwFPqlDtuuYZw7tG7VmwGSLbHUg
yifTFb2EHgBV94hn/kyAAQbjR4xChRFmu5Z8rZbwW8RgbeLsS2t39zgtAUNqX+eVSW3VFJ1iUZzH
M/NkkDH5f+QOC3wSIhBD3/lVpN7CuzO+bxMFiOSw76d2qW0EN9ruB/DQwceGrcpaIicXZ6xRUr5Z
9ASJOO84HgCHdz9cfrrw9udvrUKJsq4/KIgKqyOdBN1eSy+39ZVtsG18sf+r4uJXiwmasY0Eks52
551ODXJ0YzRGhEnaXnHJmtK8uOYR+BlvwQ3rh13+ahcZ+Zu1xCCojpxWVIEo3dKjMHfaMkXnM29C
DKJd4FAWSF/vHpUrLi5RX0kZynrO/eoOJPfcaHaTvOko4AMAJ64xAlbTr3gb3dgP4e8XEQNrv3zn
zhroN+/8Ow6kg3EIRnKsbpgmDR8yXjCatH2n/QtdSNOtWOimnokXP5Xc7CbIiv/nl0X8t6kFGeO1
yxOTQnyQ6CqqrUiAtCI8gKrzPYguBV6moNWmYvnjl5qcEV6InQwpSkoCZ8Tc9sgJXfGNgy4HEHL5
m60KJXmFfQnBGlO9z0WbGvO1IxMZ0hTx08ApYddviLJLoxzTx/WsPAEmYeL8hvagJfoU42/S/6/k
ImyINDjfYEP8LnJq6TnJDrfcw14hfdDvTGGqKDR0Fxbey/xfIbdY98/GWx9QVfalaumsHpjWhroV
NxdCRWyj9mR7KLhxr/dSgySdClqExdWaf7HnRXGgJWUhBMrlzM4ZqIixeryw9UUAnlEmQx+PUMU/
PHoqT78ClQqOkx/NsofnyXmfjGMBQI7F7JbHwMGdYBUkX1IRkjO7wBruTewlzclEyhH+/ltE4GlW
KVT1wUbKspHCSvMRB8BqjpHrcGRBKj4hLxhGqF8f80uwX3Y5fNXz5raX9ybUPMO2icsnOlYxVmRD
U1G6B8RsZCBmu9URKuda77KU7DvmUncrbG373mqIskSUFGiIjWeNbkH4hEPqoOcMc6t/1mTFf8/9
CAkpkHA93CahE9cq83UNAjn49kE2QrQG03u+xvKpyzd/00EXe5XY+ApYviOnc7A+d3xCU07f3q2d
KROGJ5QxA0/MOjEsTCdAry7yHpbFd2JalM7FtWXR0r0DoxtNb007thNJB62ILwOF99wQOFp7Pqje
VwZqJEcHbjNnJmTR0utjjnG/sNksWyr4tParQG03O+FMLC3ArwJXASGgdNOJb9o9T/ae95T8rkx0
7kvnqedofg3opwDNCpIRzPKhzhwwNZiwdeQnhXDqy70OTIMxmetp97oFZ/LYkwkgik85eq1MJUot
Bpr1/jGguPqWs4OeqBITWvsFworiD8U2enQzh552fiGkmczoGSObQXTbNSF9+kZBBVIQjwk+eS29
vEy7xB54gqAz5VlbJ/O66XYX760sgOdY8Xbweavp6w3sTSFjffkB5Y2DjpzoVLqU0JufzG9k+cxU
WnBO8Fc+R+hqa2CWWiww/lF93hNbvn+cASDeJHKMifikyU02C9iEkN8K0T7gkQc8+FSjLOEDbCrD
OUEr8L3x+jMioBewW2DbmgHA5xMtAOUoL/Cho98djTyycXATvk2dbfouAKrPFnPX01jLPyXBYrqf
nClm0q2u0dvuv/CnJXqVpyxUwNEy/zU84MVciQZMAuaJ6g3abkZnYRcv6zkjGEQiZjdsbE8204is
XNMLobyW7dTQMLrMBg08xQiQ6WufEuuAC9J2cFwMDLqma6HdqAwy2jjSBzCGiNDBVXQQ4/wrcIgs
vyAQJSmr5on6DU/L3eDJKnJPFHMBIkuEYV8rKDfOM1r5uIwW0P2BukK26w+QBVYvRXLCNqJEGtCI
OAYJZR7CYIkGsz2sbT0NIzoxIyJ5D4sUWMc8MfyJwRs8U3p73kMd6GgOxnbHMx25maOi1ZIAmuWW
MPVHbuDt44dvEgta0g3Gncfi5hqXlY5Bx8oWpiLwawQjCZGQKFUDaMRgs8UxAgjSZcwWAPC1PblW
/A9JCEbCwD1SHY0ZsDdED1D/e4mlwWdNmKe0BBPla/vrrW0vQGD+4OzLrmmcTn/vd+koSm5VsOiy
1maAls9AZFy5XDef5HREXP3v+6wft9PwfpkzxavsIrZd1xG0IftGi/CS8DgmEw9sNjAO9CZURdxS
C8xVhymiQ3mQIHxWU9DHJEx1lFhUQslojcPi3pJjqXxPo7OAV4fwaSrMCIWa1J88hL3d3lgofYrp
NbZTpSIYQBtshspaiKyl2bxGpp30VRbU4vGubQO+T9cSAs3xTjR7qe4j7FcDPgq3NPb5D3ERIRqA
SBWGv93YN7cHd+daf/nIxPNk93HSdPhBgLFTPULyy4YERy7L0NLYqRayFroclXMFBbwTdMhjMmIy
PM1lGhI33YJWD/xapMu1hsZfXT2qLacX8blUwMF3URa0oq+NjdFfx3Zdnh/lZlJaXV86pM5bHe8W
jQsgReeRMHcohiDUBrB44oCJBMlbxKprFgdj/K1KSqWj08dGBZGD7DZ5d9h3MU+YBBz4pAMEI1x6
vjHB4PX859tgMA5xNR+aGNRzJiVqQs9sVb6eZCxwJVY/EiM4w8K7Sw/YoDM+CE/tnoZWu/0V3Mdx
KN4xv4qDKY58RWLncDmbG/OMReHLsGYIT4fyFV9fAFh3TbHpnzDGvAbk7Ma1FBsIFa3DNZbulHOD
hmkTMSnYtMwHorBhFXeGB9SFYMmGy+uMal+K7vL355tZDWoJxNACjzE0EaGlwOwobKLiRw4DjyDo
ML5fwSwvZ+LIB/mNocazyjBJwTjnCG8YaA4Gc1Y9xtaKunuoTgMJjJR+xQS+ZfwNHGW9s/P0GyaK
FtF0/ZMT3mfqaBnfaY13M217QLcNQBxXKUbxo1NQu0hbIxQHRBOogJ58Nn/dNgQOu1St57Pb5xTm
0jcmLij4VvUP5PYjYL/aUgDiPdQVmedpBNfwEOM9of1gzyO7leglsFojtAXHqn6t/okw8TBECnBn
yVS4qCiuz6WSIbwnuyUlqOHXPb3rB7XKMVqP9iLqrpSQFW74P3cu9lJinmAVyvPO07rxU/b1eMxl
R5eBhzPff3XqaqsjGP4G+MqYxl2diXVGGyMjPKlvCYkaK57l89gaA7r+lU2Ll6U1GfVq0srReK3m
JKjYECpnZH4sQU9rraOUG4OOXF+A98TZQUetxXm4hM+bfUA09bLesSgSUfe3SqeyXsnF6/e3e+UC
PIMUcy5vvIXlq3nYtLRA6mUJ7VkW5HocUremXHnhths3TrH0G7WCRLa2PYOfnSj+KsELMlkM04Ws
DANPxXx8sIAijCHchlXTkZ4vvdUTTU7tlGHEqHYvHFRxjHHafkhUk4M0vemrOJmmwrE2N5sWlg0D
nOyoZsLpLA+0PG3m5/mYjzKRr6pxZLV1Z+Jid0qNNfEA50gzbyPlUWnHkXotz+ghR5lw2jhrd5it
vcRELVMOgJ3D1+ucEDkUF99DgaNwVUFNjhpY3oldsi40JbZ+9Qds6UCDBBmn0vnRGmsZoenCAIg+
cxQjJ0ZcS0q+v27g0onuqHVFzfxsqVrRz6wUWzRQTQczbmOBD3aCDAkUp9IK20/bqWHBqWjuVI7L
7k37mmdbJg8FBlP8mVAtVxQg/2RUIwjG0qUOhbUYli5vHkgtX1t1Qmz1ul7elgrK0n3alQp/zHTc
mTAalktNix4A9/cC+sx6s647rxVCB6k7Zx2MvR+olNSD+UINsmrq3kw0FrAJQdsihQLEHq3cJwry
rBE6+Ir94F440O0zqko5TBj6tiK6FqqB2++EHGUpnPG8EtQkHmLBrMa9tZVWVP8cZdJrev4Jecyc
OsweOYpIIvyWGNrFU6gKxrwrhRWfJpkM6JZcMgg2EqfnZMvZ93nc2/0zn9jYms+7ja5sPhEqkksS
jpycHI1fvXoVu+RdEjZSk0U8v2h7xGIF3JzR6ZQkCKRrrSOCcA/7jcYsv6kslb1WmslMjZz3HjZf
slaLjoPXcImWo0vm/BZdhvnSkWSE9CWFkERrDQ1idz1DwbY7DNPftfg3a9DMeO/ofWt4iWhsYsVD
Z1FzfE/m0+vLp983e21Wh3F18CVSFbPMEKnhtcyHgqyVDljDVMEQhoGTCHxkWsMuelvwY7xA2dKP
xtJNS/aKByqxP/Y4n2hCELsJbj5Nkkx+YjzUMkpjkYA+St493vNxbViCru3r0SpbugaxE7YY7K5t
QL0C10HFm7UAbnYuhZ4UrMe1vDbSU9rS9GPd6sGSBS3actX//s+YdVUl1o855oOGB99tOg==
`protect end_protected
