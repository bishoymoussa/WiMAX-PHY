-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
rnxl9FtH5pLbbhnDtCQYTXNTcqDnw41Lfy7MI2Wyj6O878WwvOTKWH8Pa8v06gJZvHx/BXptgUyX
U2nARCKVR9utGhSvDcgHEsAntUkVficYK2MlGonrcd/790WILD+Qk86P1GzsJJMYwUKm/MA+HXM8
C43zjd5MPEM8/RsqVtEIA+rehhvVdmU+FT4l2tSZF1wEls/SDV51DzlZyNWqVT9b8OU7HWzRlwc6
vmTR5I0ISZOJn5Z7Vm7+F3H8Afm/cLbY88gj3xlC5KhR8XyM4LFs4mHgfgqYhoZZovsjhJX9UppI
i0PIjPNYXT3OovXMOk2o1AwQYviu09M90m79Rg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 71328)
`protect data_block
cCtK5K3BNboVaTx6lQ+l0ouAFmI8eHSLGAsnhk2Nve9hiATjx5meX/KMhwZWfzplFfsdpKMmShlf
UN1bbKP28ME7kC+QzHBpJtdNCCsj/x2dG9kBN+dBGjndQgtcVYmZkMsIQNkup40tCqfTngweuKJ3
Lu2XX7Qk1Hyyfldap73naKZyTCN38RMz1K+sb3sKphNuOLm9ps2XUf1PJ48h/7QqJnS5I04dRS++
JjlNZn2yFKeUdOyRb46ed+KxtbvcVF589Lgv9v4BqsDiyYNjkCyWRa8KHABnxY6GZzkJwiFThkCD
HVWPdvCmsnA7ZJa3dJRdjugvmY5OVJB9m/F26Hwhp0qZx6vrtpyKd5fB+JOm73QhM3EjZHd7TyZK
o+YgaQAjOot2aXKJ2qem3IDBx3pzcZjHQbYsqSeeX93iAUjt2hOYgx+ykh6LEaSyis8TTTkPOmOj
Xp3rhWhM7fq+QVpdfojhfmCf/ObbHEf0J1uYCWb6pJsMwsSOYp5zOxF45ZsXysQMmTugG31iR0zn
5g4nHIEWLdbfemy5JJeYUwAX9B+dQDSlR0YgdF9XstPZa2ifnQQ+i9NpMXUTZba6WVRyX6Y2lZ10
VJ4h/gpMFuQpwDJcXXLjSenNjz5rdmbFO4gTNQDIL6EeczL0nOGhDICL35wBCuR6n9HAbPxA9oge
+hCsrXLfdEcNkaHdIKfVI3ePThleiRtvtCy1GKnVsmKG0XXREt9mnR4vQNiKaJFGpESG/lgfDnlK
qYEdMg1VntSVbF0gUseMbDFHqxrYqEg85G0p9bQZtAPXW8ixtoJXuGe18869Fa4Ni3T4+pPC0x4/
RDjBPX18jXabtjCir83wfFQS74+SPt/afpZZYzae14uBIFOjh5Dkwc6TAWmN96oVwR0WSn9vM7CY
hWwiD26N+9+JC9GdtuUaDGO4hOqmhQUcnBR9UXaECnbMNLetY6+HY9Id0giPpIXi8VWJ1PEanA7h
xl9BMFH0u5r9l1FfitASNkQNyN9E7CQ/OelcKNOm98glnZjByjc/xjFa04/LXxXVdsCyrhReWUw0
sbm7WX/aMae3Y/QSSOfTGk/XDNEOOlt6OxvKae3tJLudrDBn6WiwiuseOHynA+fTEM8Tbmv8kYE9
IKZnCizfz2NnS2F+xZEQlfWk7UkrU2pr2x97AUCdsRWsRSdscKaMXofuCOkR14MmZ8q2fibs8iBW
vQEfshHahyQ/IriJ2+rYL48AGoTZGGMyCg2EqbaiSFhZfCy6uAyTrLBjcT8vx3EFZuwXG4bYAILV
D862lke+fzjrWnc3yzTb6S8IdI9Ig8nmcqJJ5bCf+D0WoIqCw2maWSpyFo8TfDDGLOV7JMFGGCLf
OS3yw04PfrP730tN1RVGIt2TQmzzfPpwVWSr/ND2hxUctOqoWStdFSyfb49HcLo2iSAvRWk7qW8J
WnbtVnOG41eXadXiUIK+xsjkXn5s5fF347YRF9Jw2pbx0ndloHeAKk+S+9uRBq9tLzqaAJbq7H3a
xz+pm5dGjqrEq1iaibOkV7jPLlg+jb2o1mBUUPpyEnu9nTgMYSN7WRMnhy5msqRj75zzc3znUxOE
4gKxsMPUyzA2KaaWsmtYWdcDt2V4eMig/KaQm45P4vNNI1DbIfVbTnX9ZBYr3No45+AhWxUlOtnU
PKYWkpluGAkrEoa5CU88BvXeC8n8vdmOAdRRNx30oz6n5c98CLpem0g6x7MFkuL25/yw8SaDVH0c
JW4gnw+7N7mpZYFznnTnIdLmwoUhQHhXGvHCCMfPRwQ0sjerVprjzpMAWOKb6r+zKGlE5snCquTu
ft8/HF6P1AnpfI8lE/3GOMMr6srbk2+NOK8IYetRIWQQD5boWPffWqKbNT/SE/rslpjU+uXyyA/I
XpF2/1QTOw1JcmOUINcAzaEG20aYG/MiofVSCYja5NDi2elWh2coXFfegTEiRsxLBJSHyoH3/1YO
a8KCOqFZ44pTGo7JjKO9xRvhl+cp26mKT+VS9xMB5+r0jTyTMyTa3cvA8DA3lwHhde8EVz/hrYe/
5/bKWSjPv6QHscQBuJZdF9hhpaesPMwZPvb3ZwoVHNS16DVe4+mHF2zraedDLLhvZMyFYIRb4Gpw
V5JGnsi0NNaKYxlumQwqbR3VpANfUpQaNx3PsYO2Txqc8VJcoTSvRVuPWfYJFQKXlQc7ksyJ0qCV
UJhVu391QuQiugRvV5p9K4FUTTAVTf4dYdwlrBYlqsDJIIF3InyVU84Hsoz4UjE/iFx8l1/wNh/y
rmY9UIAghqcwlBOX40tj/KVwkYlEPMqwJk48uNm7pL+IASUWumy/jXKrfoUpmGz/TsV3YNr59/AO
b4RRqQRWLgD+P9qCliVH/3ZaU7gF9cVtNqFr13W70DQw3ubb/QxDRgU7bn2AufYirKiRmy5jsL8V
nFuy+3jMNssEPlwsQQ/dZAfHuujObOA4lXznnws/63r5xSVFHDcp9SeLrzXdLh6bArj418qnWPSi
+DQaf6TCL+42TZOMTL97K2mSWHqy2458dnMNiocG8iTeokRqPr3gwG5NCDoO8j06bfXZw69hds+g
ExWwYLxBTuYwSAKGd6sIva3wtPVc3/ykNBOGxSKnWJFFRtHz6bsitePRmaYxn6hjFOSc71iKEeMo
wppwJICkzTqSEhEI3Okk0nH7EYXlYTcnchpchGz8/3t80/XHJ3iJr/XICbU+o9ntnQRbBw5zWy0x
MpLLtjdC/Hy42Po0zvxUo2Yx/QDxMXtNg0h6pRLLMXb6KN20mrPgD7JibO8VVUKTWPgy68/Gl0b+
zvdpNhWucBs/VYuV9kozyPh0WCROQMIMaZ2KFtMLzrfdnn2f3lIDFP6SVw8QjRG9dJmm55N4Zt6d
zmRGb34Jrudd6Oxhwaqq1KLAK99/ibf3ME/oCcVTHt21by1xdMYP31CUGG+gRVr8JTyFJ8ev3S+Q
wxt9d697aFcM/LRo05uO3zMsUxtRm92HSOzxlg9mLWB+VielDQSpLXO2p3oSb3x9pboSI/ned2Jn
kQ6aGNJbz+AIfDsOf6/Cp15RhK9CrSoj/2Hcj2l0Fw8jVuTIyu9nE4B7rbYutzzTnIxxHHCUv0bK
vk92fU4np7j9Ky1jCvDP3kTgfj+lEt7h/y6n4yjL7RvBWn+9KKKp6NAvyVOHwUOxKsrvnRCbDX0j
vX5VRrfZBVX2YAtmegDuhM4NFcaR9VTOUfq2kqulahdpPaHtdheEcz/ZSFkbmv82cLeeKkdZgA8r
rF3x6Qd15BEV0U1Y3JHatHqvTgqw4wDGii/7n6sZKiZ07REqhgCMYuGrl4U84s3SrCpZxt3wzSbk
SqB0r1KZ5zehzzkkyGeuLdiBJSrgNEeX4LOoZNzn0KF18Y0P5n6aH00FGos7LiJlc/8Van2hde0p
Y31eQm2Zmd1Y/aIFVxQeLzNE4DnjG8VvWiyYpzMICjyIP4h34b/pwpL6d8bt2SoAQ3UGtl9R99C2
66zzhnk6tyjePTKvn3GhbbtDAuHZC+Mwkt3yVSUYNtOx/Hazdz1fPzrO9KQ3BVfkJhKthuSgDN8N
ckmybo6jsiSH6lOQGdsGhCrBwDvNc0ud40TyhEI6Eg7E9jcWL4iRPFRwXit5Xby9wWNbcUjHPgDn
EWRO7Z8U2vXNz9CG7snwvVIIoYq6Wp3BzNg2qtz+IuyhZUDdu6/WK1YZWgu422yyQjcMa0N9fKJG
6YtNW521OaByi8und1K7CT52QxP2Yq8IYcBmAiyB3NJy0Nk6JuOL9puhtupc/Qe4Ir37zqAmLNgB
PyIjn1vXTEjZnArHcPzGR20tn0YJIQ+R5eG4uJ4S7/nCiwfmlY/wUXFHI9X5o33IEWUb1eWedg9/
KwVgmuDMenSeikQs0IfoMomuQioPhFvj/pQduDJ1VitgowBu3pbrTbYV6AxydHCeTqNu6WvusIQT
T0VbOTQR9EeT+RJ7hEVv4AaDOb/FeSm6QJkcUvyAhsX9/dHxX2Fq6cZ999psK3Sl5X2TvPTL0xls
LVtpVLpNENno37KAXATPZXWCnicN07fy445x+Zt6ipWdKFGDKPPOtX+uwuZHccMTv5j9mdRwcIwP
mF0o4z76UHpLg1Cr2M+B2hra13xt+HZEx07eWA06Zs1ULMFkxSSYCTG5tjLhFFtNCbhSvL290mZt
245bnB1hQ215igkOdPgQjgJX6wsPOgLMPpZKD5CXXlYbGeJYuFbECZZMs3qHHdJo1LCu3wPGkvr3
873OCs2fKm321ovJdissqDnopkCvPCukuyektNU4zWqhC576nuYTvuxTctI2jWU5Auniz4HJJtBY
1fFPYFj1BrbO0UHwpsobHr+kknQbMaqoHKTuL3LpXUe+tW7SaFOFbZtin0dg3Q2QJ2Q5BLBbeAA8
VoEnXOoQ/C0la2rV2uWsdW39lCMSCDVpuVGMdApgctjqSCnhXLddyt+Wr9xhfMXm3Z5I+7lHNTxz
IHku9bC4mzRzNKdrQQg7qMmKfqfQVfaW0knpbWYz05mRPSOTrnBnJGYZYWQdFt1XOJts0yXDd7Ou
wFjICILYNqCHu8nJxKB2TOmtRbpXa6t4qCKCcZtwevUeSVtvAwNSRhjH61+gHK0F9Uxng11Vt8Kj
UR2zWD5b7dsWoafG7s0t1UIVB0FKkFWmLCO/lzSD87WLDbpEujerrCj2s8fbMYACVgVShMF7nvnv
KVWXVhSehsYcNKspYrP34dpdVX7ck0eD2VqDzvkor+gHWQ/oO6J9CqjQbyVcVloB+HJvbwWu+UoA
GH+zjG+Miw8PAYVLZZ7e9GaIdpEM/ErUUNv/qB0PUoN1rzkr2hm5QvwoH/XC2K8iltKtGBW3GHY+
cbGoSQov5K4IfVrDLjSxWkP0WrtgiFO2Rhluv+cTMYprgI8th4iLC+fq1q1JbnXzUgEuE++8+sT+
bg5IA4b8mo69caqb2IevyHRxNAoKNmJnMBMuEdOd+bVWFXXfLqjxymNWJ3iV80Z1HVxMQ2g6SMEK
ClZ/+dmVaZyKbVdRYwwuJbqCZoneSc6clDdz3Mjr+xVuU7eFpM8WarYJPq3WCXiOMCnxYVfbQZJF
8fyTMRpJPgehm6Eo2VfoBO0nFgdHU7f5o8dLrfX3eHZH4dVxRghbPHk/uqQ73fdpC9oetAODV1gN
g4uDD1MfmNXS1yzQUu+4sc+4MJb+7LyjwSGV2lZfgP6FSrhG+PlX1Flv6fixCiQERVEIECgQ94WU
NmAHGv4It4ravxUJR1swePVdwpiHZElXPhR4hH9E5ylEJiIAZGFItIuy5Q/0/w72kBx8E2IKKHO+
wUytSMfSI9mST2r48cRgJZE5NkZQWQXod/oMXafiBpybswG/aSe6UMcHB2a24eSjtz2OM++7xUDX
Vt618vmP+ulLY4Q67l9bzYMRTW9p/XuI1J0GFFLv/CIFkcGGebMHam+XFbWcfpk9r2gfeSsLEht6
AD6wzcZemrP0eWPaSnwlMZedYz/fTlexy2+l8pLyR5jlt1hjwFN2NrHiuVW/KbR/N/SooK0vfKnZ
I86Ij/vrmQJiwW4PKHVyyHhGij9ZDkC/4TXxAU0PSGbGZpyJA8fqFZJJTMkCkdiWgVzvRv1W9n/v
G8pUkEJXQ3pwN2pmVM66oxzZ0b/WdT0xSqvMkTgvn41wP0uP2SjBgqqmVQFr3p2dYI678dDrM8cy
lvL8WsaiLgJLSMKJjN57OHr1fV/ZNdN9HzovVOHi1SVAtE2mG6Q7RRtJztElAq9R5RKv9yUqJeX4
wK5EAVB3sSVWbzsKhIRzYtGkaEdFkvY6U93ilCjfVgKjA6c1+m8qKtH/xHLGsm3gfUR1+Ldj1KD+
MNJbMyqSaSu24px1QBO37fmTQShPoUCmJdf/njsHOK4bzM+51ARnwtOC4UodDSu8PMmahGnZ+UVr
MTvk6RQbQhyecllEfGRl1gHrVuplmG7dJ9SXaAtRc6pfh8kYD82Oyz7zJRTpsMSTnpT/AIJ7fEKF
UKDFKkA8IuPI44l0i428sUIA+S1xWAiy6+3C3+g6GnqJNMzkxdYKyT0qJV+aNN1dfLYP4X7iH5eI
7ussovqHoct/xuA28HOyjnC/TVFG87Rkfx76Cw+iRjeLh8aPM2EvhJbvV57KBS0Ve+jRZdUKkBgw
v3MISjs5sT6e0HLJWRTHJltO+xcpl9K4Ltd46LzJ9cblGPof/BQNCKO8i58RLJrpWqYsvrNDZY7e
pxJtsyry4iosy2Bd+S87h/ly9OPyxU0/aYEoSIsVJM1fFk4vLOshxpClbpgGB7Yqn3lLfdmrZZrn
FmR/ovgQzcunO0WW5ZPB/NbEr0oWcfiYNyhCmN5mkF7LvWa75fe36ojCVBrrjvgFrToq9sLa3shb
iVE/5kWIYE9jQ58doFSp4me+KMf+hd2NF2IMVnMn6690E6dumocq7g1H/i/zEpKra/ZmL5bEWO3E
nNxUaP4/D+dHuXAmhWu5HnvVfe0bbja59K7xjG6SxdnfgTyMs8Iyal4SXOva4vQSfeKRC5eGizne
a13NBdjl06QzfjTTV1sXYuPaLofd6bcgok9hOke63TJd/V/5Al0ZYA+lEO8hpKCNarZGvr1S1JXT
KeJx7SN0TktK+cUAY+d410j2TOSg9PQORkXBg8V6F+NYVKV4jMtg8JVMM0hiZemE6QHr4dMqd+e2
ooLnIBwbQzEYOG6RrcpzSWWr7o8hd5HwWPGoAOnwmZf7Z+uvzUYDDsM8jC/IzsjjWybdPziQH19r
LewEAKIvEPvWBGjyt49LN7g/+TdFi2qy6sT8kBuf9HPNDGUHcQWDZZLouLQzt4a6VKVnIhfAwtiG
vT4WChL9/gkyfq5btjF0YDDNx6K6NynHzKlmSj6npKkXLueYBUOPgVRxsY8LHQIPY0zKn13Iidik
XlnrwVbeT5jMhxdv1pS4wyQO2Z2eyvMND0NBkWP9nRb1C/ya4qPkZntSkqk7PjyaFu2Kgxknr8L6
RppU5wbgDpZjGfxBjq8z3sTW5jofXVp/4QxVOKzBt4i0rP8w1tKTtyRmzpMpQRLIknwru8LB5xON
Ia5wS6xVpqo1Ll8YwcaTg4EmJeNyzQyYB4k9nIN/A1u1kbZ5D8GWw0NQAg8/e3TR00JcYTpXd2YW
Z4QcCoFND6QOziMjTcX32WEa/R3KlM4nQJsTpUZdR/pktU6xbwWogThazxpT3r7WZQHfZ0obwDy0
wVbL5RI1iLW232Q7v5dV0/W45WUFmt99xEpiKp3XtDirNZeVr5GQU7r2yK2EUoZX7h9fYFeGN72G
zaN37yWX1re/Lma3MA5qAX8b14CjbaLIGg1jHOF6hpb7YLytM9F/PYmO4AueBxoYqo/H1uyrJD/o
nN7HBMWflrnBXdS/urg9chtuEXC97rD7UefhL9thj0iZBGhERSqihw2SNvoMEewy2uJEzl4s177E
wqaBO51EREfrcZs9wwqjQFudtuUcPTO0jUzq37dZ9aBZ2XeReEzLORwv24ti2HiOm84h2Y+YLw80
HRAKgmu1mxLyeu7oAI6ZlI4wqEm2i1ofQod2lFnr3SodJMC0Oxv6/kLTkFQv269F+XL9cZygv1as
cxOcOtgWeUwrOAzvdq2Uf6sokkEwbSfEaq89IVYgnkj/MmKk262q7/DF6jarpt9gq4bAehTt4Lob
F9GSdq6HuDUF8AndvG7YrTqmQwfpH+aMXAtFYF6Z+BCt+Z8cFcKTi6GvRQV2nzsNnZgihQod4EKA
aYIwhb6qw4t7c0Rnu4eB+uLQzEffSiGUm70i1JZkKaYMP13D83FhtVaXkL42MgppDwp884oc2CwD
nIFCZfW/hT6cQfcFNo0vd0TQM73o7hKEsvvFB/IHz50nNJn0ogWlyJNzYAlA4PcgrgyuGivehwpo
Lg33egPz6BF8DQNmQG8KcGJNZbDW/OFxoWw144QbH9qDcgwbxNOfE94ltVtOuhLKHo4NzC89OByG
ayX/fWbOKt2Q36X7+ZplUuN63yD3L0DUK2GSKUIaYxQPNwdjWqvc+arL6OpBhDrsTzA5vrAZu4f3
4wkyzGldVbYFHDO/0ccBxb1AetrScsGk4FfBmYnpKP/Giu2H3Ee7XymAsI6q/RAUJ6CxWGo+lwTs
5l2v+njm274OTahYawzAXflDeM0RBGdsdYRiLxHW/65K6Gb5+tVhj7I4Njvk3ddWeCJatJIYJ47z
slJ8tjwLnsqiaMDhiHqVJ14hKXIZYsY3NBVyqLvHHG2bv6VJ12NnmtIn22tznNp4dn4OXf+LFRCz
isfC6AwyWR4jGhpTCoaC5OC3ORAo77AE5uEcizXUx7d/HITOZ3ITCwGCXQoM/kntz25zvtL9kiC0
PTIT6GkbRUplYJGaqbqD2n7tItLYwi19D0cLQD+r0r9eeZuv0T2LW5tuJrPZyJIHBo494r59U5MU
stb5ECPQvJP8fk9wt1QFel5gX68k7TzWlPqUiJ0wzLbbY+kVB8svHZ1HZEtbrE0XUJHruMWHIIjS
w7O2aYd+vHehk2txp9Ug6WY7MdiInViv2V/SwwcfNRd66dofB4YmIUt/0F4ewE2NKtOHPVN4kRa/
r1ke0ErmK4I7mp9XJBcHAtRuOnzUmQ/4zLrwD/2+/mpVLDRefulMfeZe0THNDkdUk3PG0Vz6X/sV
23/EOWxNgWjNp8TAQWxIx2ifxXARcWshsfmApkVyNFvip8TqDro9TlXP0zxw2MqZKPtuEYm7Pr0B
LyMgsnTG23Xlonk5VvThd4sEooKfq4hoGyMMNWTInhpmh01EkVutpBiOnmetghD49a4oar3MdP80
JT+NQ8t328YBIwSnZ3X9v1Xe0tahvopKx9W2COWKh4FfRVFOF5mbllf76+WewYH43xkTvqd4rtp8
6nUkpXAmcCLJWEVEPd/4DiQVoj9fi44LtTLa1Wpn7TsFdbekz1VYgyr2HF/PFzYRpiEimZGoe8kb
oBmQOH2Q4BDt03xL/xBiuxBVg90rZ9fhwKv2HIcBGF1rI2S6+XCOYXlEhF5PS3pi6FfTpsuP1Un9
WpK1s4f7jwhKIqXETwq6VzcxnA1YRyVZ8zX+BfUQxxJM2D9BSOCmCzgd1WtpLVZfMyAfERVh/Rmj
LVhuTF2AMfK/81BHG3o1bl0qxqFQ5eIQM0Ns8XKnXlJy5siwuu5jOZqffz3hEpmZjKr7noUEXmUC
0PtOzUAxL8ZQyg2rz2R75lOk+FjSNeUX+7EkPb8whuO3DdNTFkNWbb4v90S+0l9KQlYTwklnTir5
8SRiple8i3AeGKJcJI9F6cQrEmRgf3QQI9l5qlducLe7MisfBZk8kxxW3clxCFgO/3qZZA/9nEgv
uakbbCWX2WqkYUYhfgiRA7W9Y2t4egoGVfOiQTUNR7M0MUiwrTPwhfa7Kx//dsSRgsAPYtX7f6iB
hKVfUwgalmG6QD1H3IRWSv7ny8qDvqPO1QW+wWIGbghnlwjS1WVB1WnuPro0SqoV0hFZTmfZQW6R
YMKF4xLB2qm22w8dfMqpbu4GlqDsKgB9RtNl5OMuTMhEub6/DXbUTZXL5+XD9iQc0EmO/Fmxzhk1
nTSZ3FlYwvI1tHm6pTFirEsVm4KqiryS4keq+pXqz6DkLWiE3MQY70KP4wWIlnZYg2xHY7qfk10P
FysI8aT6/BB7GLhZI9EE2Sy5OJYv5j4okRt/j8XcdxXW4c7IFGBG2D1yUyYMPD/U2oEns2xI9vGG
TrVFgv0GzfM/F/sQQodJaFS1L0r6SLAMqK3Aao85vW6tJkacMH6gZUpxoZIqxV5Ss4hieNjMDm4x
8llGv3MqKAGhVIfx+GFiJH9XjV8rKXY9/VFYpRlatbzVzGXxLbpuNn8m6jc9RPwxEZ5kzRoo2pZc
sv+Ty2pD9k8nTqE+iGfKmRCweVOmYS2vU3Rru2x+ukRul4ajzoAbUKi8zClSk3K+fARFB/Ns7Szg
EIoymiCSNrv4pl4V703wNbiWkrrBBNEXWNdTypawi+1kk2jPsSKVMEVmnRjR3w2InPuCUho3Ldc9
AvZ/JOAKGGUebOR/xM2UDVyt1ZwJ4qEpO3kpowLgL7PiCL7HrXJdti/XY3c0TqP5Jc25RKOuv+1t
L8LbmbYgfWIrx9747Vt5cQX4hyZf1iqbiezMYX4gpxeLWDqwT/0wlRk/+vYCMAIj1Xq2NxtUf+GF
P4NnFT2fFvMZpR1iJ35kJwrHc5IlMvUKNjQVNcCLjMg8hY7+AP+AhqfLDAqqVt0wTUsDRSM+UsFf
wFZ4EVLe3IA4ukBLbVK42+5Eg23ETbLulrspZNcnIAI3eS/UihDFacagBomPpW8bnv7LCw7hefox
vHrC9T96x36vFBoctsFN4jWLMaszyF352a70VNnxIjo2SBmMO699dhWSBJrXkUk+n+fg4JqanwNI
FbAUY/G8oAg0gHN3Jwt1BpeX2nc79BB7sL8sKynVyyx+WAzN4KkGuOPpy5ZqIoM/ihosc3om6pBr
tP2/HRMGFmQlHibTjbJykvN+V5LD1H/NjnoFuZJuIgSZziXUS3EoanreeQm500E+ukVKyqtPmmag
Wl6bMdBTqoIU1ZgKO//bDPqF+i0ax7/lGZnknQ5Jp4QAuepd+RIRtmqK9KZXIvudfXGnE+l7Sv60
qQ466x9fFEm4RrGh+yRQ3i2otOOmGkavq1FqkKba01m3RkiKEJIGK84J0py0Q/q7NFIlG5W9nk/B
DcRDTRC72OuiN5z5t9Y5Z2vyZBkwyohtZ26FsnXRlWtvD4d4muErUAsaI1AIff7yBD3c8GjZKf84
EzAZkWA0COmFJQQQHL0T6QbeAWIDdO1sdWwCVCmOxDQsKoQ8E1hGBrKduyEQAGgsTrbAgeOQiCRZ
49uTxGMRDrNVXqHLvlaqZCkNLXGqaqfvtmObWV7tiIIaEyRbIZSuCYD3VYWzs2DJoOtF+Xq7y40c
uI4l811h52yPg3GPruwU+/tPvpkoqkYW22ah3YlJ6vAeLpXgygRmY/URgk4MFfPdJkWksbxQUIL9
GGzd+/uH+9K3nChFP/MR5Pk40cx7vJQNmjkHDE0rNW8canAKsLWsLcrb9yNoLJ10yC4kwi0Lj6Ix
TUWi+2GX3J8G1n0k6l+52ir1N6ppSs5QEioQ/09+/xWgSSWWTHNF1ZAwRRWDEvWyBfTArJ5NvL7E
BLO2mEqFQYM7+/7geFyRl6Zo+wHVTEUYoCaslxzJ3ZfBGsRhBNbnIa5vcO1Qyv0Vl13Fb7r6zbNy
TY+qBkWCex+q/40FoKcBOBfEepaSzomlig5ub8+BNPoX/bFd2cOvGVBG2Ht5+X8CEoSIGGC0jTT9
Z8VUnev94kuy+3cQf3KVhcjQpZSoa10J3Mh8y+rSDyUDGmi3Qdgu3yWPZtJEIhfXp+7xTue4zqXG
Svsy6rpvcImzSse/aedFshnIaqoWiXCaZe8Upnm1k58mhIM3hPWLwE+AFv4O7xJhVly56mTsGab/
/lAPRDUH6vpycVpY+j1W5XDyqsL411H7jH5q5ppd6rz9KtGpz55rsqXneKktH39VLXpvIPVZYUqa
oeqqApe9dh2wRTKK+Le60K2n+NaRkOujdaPVkopcIKRvI6H7KeJ80Tc1s9qf+OkHxQBYEf/+G4Gs
GRUwGwDyf7gggao07Q8Uf5TAOK4MAXIZrg8DuYMbzlJoizUN5DkHepu1NyqlRvAlK/5zEWSIqqpT
X1CBl9T7bXW35R4HTkEzosQrIiJ+wpK/abeYq6pHbBHObmmFToPyX523Fw31aTp6Ttfq3S6VhsWW
Tt+nfSE8PG++Uu7hejKtbS2IA1cyXEPVPE4z8onD5KnDkALhBF4ATGn4IZ6HJihpWVAxwRbiAvr9
uOildw/TzhS1ZxuXHrgQI0ahHQ9ik2y6fB5yo8HZUuoq0VK5zTR2R63F/lWOa4+aYZFR0ujgwDli
T9FoY/npPhPXGLiEyKgAwxZ96TerkTKLWES368jMbLap7voeSCXlMtYwgQjpmvy7l/lf5aIT8pWh
gi94KS2EG1GYjCkEHlkToBpUW5hoFVTXBMRty4r+8jqxeKrZuOrDxS5NWB+0Gy8guLO01L3kp+1/
TFb0Qj3y/BujqfA2OucRhoCVS4UFZQ3O8UK6CTi/P+zdUufr7LsyA6mdDAgedGOy4rdtSbPR7uga
r2KA2ma2v+iKtTUEIpPrfJBhojgojaJzyvQyNQpP6wZiQxwzx/CHitsrRxrgbpwVSQ9nQvfID4mh
x4pseXMfhugDRNVmAd6AbTcvUhl6rmNnLQuY6SsBZr+vGxViyZWa6ENL9tQemKmqQWDT1XFzBD0y
yS3H4WtW/+Csvqwt7uIFd5gHMSxMMm6K7FHFufObZTbtWFVcHhdjmCLLjJzKIXw7YcQnyVuQVdVv
HyWkv3oabbAuxRJ8RamK7qWs5vYashaLTuY4PjPwhL2fQHvLhmB7lySTK8f+51Cnone6iBqSoyVD
VhNpCArg2SRXErcvc7jkx6lM0AS2F8qCvwEM+2wA+G57SaNAsaLHc/xgI0uIooOP6fgxwTG2kNsK
yIUgu8a9asZ74QAOyXIXmz9gQuU8z87yUBI6sYwqsylW2z5QacPPAt15s6q3McyVbsMGwMp9vuW+
cS1xRjpgo4TdUG4B4DcC4y0CPm6QhkC+IOQD0Lq8rHe7jJgR3s08B4VOzMY5yBTCmVzA+0bu1thN
PDw94HgXFR6AZqAUxGESUmkSrmPvYi6eB7bOzWLEENyjUiHix3e1423qX4/I7ZY1cR62L76KQM2z
RaaWPx9jQoCd5qDZiMXF8z8SV2xLViIiJn79Z8b/xMOEPK/V4VFQ20KHJBu+9/LNuIh10VkTTcIt
QMd4ZG7Dk117J602EYik0UBfjNpiL9hPSbwf5mG9tYYYuiKzrU5DNGDJDL9YYuFSpQNB5UQmT13/
W+DNSqP1FKdmy6Lep+6HrhSfSoSxjtZKEAozymp2oVJuFUdLdAWnuNciXGsM5gURBbRjXBLbtdKr
e903e+8ZOwQqIii5PqoW20dtvgFC0oB7jizHYXGIf0s+v++x90MOV4CK3dz7GFOoXZJAZD6GL3dt
Uxc2HCJVXLh5Zwsdwm9M/NXgLZoym81N2yj4452Df6CgB+iuxUsMeV3Ui+mMAssjBRDJJI0OQMjl
N5VcAxIxQCQep6KNOYPk+jSLwO2WQBahuSh5B1NRk8pZOsCbTfOEWMLeIHEK4lejKdVHN/Grj2da
55wnmLaUrOGX5Ez/WIzvXQr5ytuEPyXOqnE70cQdXuTnJL/kjHm+hOyLBf/45gwKaiIsC+xXSZr+
mGecXZ8+VKRoahEDlzr4k1HkBvXe27Z5XfSN1OfNcSaNMc5xOqsbTjNHJgYwUJbD2oU3tzYBv0UL
eLvn89X8au6NRdLQEvm6W5q9GQIoNOK3ID5ebYJ6dhINCj3gl9QWu2snNXgWlpTEYy8kZW0lbece
/QWQYKHwsVAIAk7Kq8/V8QOlj0iQiQZCwICafOBn6IovOFcSdMSOqv0DojOhXC82q9NEKcnSxqvn
0SVeQMRlbTZSW4G7f4fCnVDEMRnN9GJbaqT8ciM0lVrNgqscPDoxkWgsk5SDdzrvMDYoJRx/328Q
p0tuCUMsRJmcbpz3QqboINK+vzE7zfA+DfptDrGeAJ4O4nFA+3JvanZn8yqWVHS2ImJkBNK8MR/1
QC9MBBhmYUVyxQ5ANbNBu2A77kd4m7rhj4kXb/ZyOwaOW/+DvX3fjHmLD9jQxFUrJdKe12KIWi+d
aCSnQ1xTee+LBQ4xu4ADPPzTz8UUatpSIVba7OcQww52VRxyqBJaXYQrCXF4gmETQgTzBYXf4LlS
1N3xQyZe7pBHsgJfBFaTg9NeTY2VSeovlkYsQylT1lx5PxMyvaldovAhSTMKH6L2l+En9WAn7CxM
fgJTMFTYlc9lpHlcOZEUR+kRf/f5OrTTyaG+WUyNrJxltPJrh0VcSfWxShMqeRVyPM9ar6eT54BG
7L5xadm3xQaAgUDBDZGouffEKEy+KbohkgIQ2R5mj8iA5e1N22pepGxgSH3CoqYKxKMd55Nshnee
DgcjlyNkxJXlthXQ3pfREQafm/ocscaOVPN7032/x8GoJbRq8pVQmfxcaPTr354HxKbvXt1yZT13
VztYOxIaRfKbapBXt4sTtodekba+ElFr8UgX6D8zlW55nv8lqNEaBenLrMbSVWMPHr3uY59orBR6
l6qbFCDYgXxu++hvECA6LGcxFtOSOX16FUIsw54PVK1oO+hKv2q8tzqNYFjyFz4tRVkih5xSmjYI
9ali12NLmRT+IxGD6QSecQAfquvj5OCDJj+96bLsP4xs0hw5g8yZa2VK0v/vHoIjQAs+rEa76vNo
l+pujnJCYmWbJN5xfrynqFCxdiFY7qs0dJ5iKEaVqj8yfk9ImHCBOnc2IxiIxIu1eNRXBDe9vJ0x
22F8pKy9V9fosYENtInNJNanGoJNWTy/0NGJ9iWuin9rdQ9wY2BAQXTonCMhNPLgfUic/MaUfY2q
dSnrlgJz4n5RvVc74V9RfRJVNeBL3QKZ5zmfVq5BR7X0+Rcj4CvIH4PnOfapewVRV/8nYACmyAon
3UsiPpwAMsKtUh3d30D9sZPYR4Ll2DM0pb3wmTJrxlraQprQ2CTat21ztlug5/H9F98+xt2gbAST
j0XhfRkEYNkPIykcqPvkjq3Lq6LmzHijiWsxRWbxL7k21UIV2v++f4kIjBD1pJY7BoiJ55cQ5iz7
VWhwj3NRID+jKiPfRulESZyqLNf7qYhfkyegIlwBFWXtrwQHggr3bcfhLAHxKUJilFJRPKdOlhK4
/YZPh+SuVfkUbmk/JQAgjZGD6g3xscnaHVXnrJFPblQBs6UKm5BDFa2fIvt+Z2pKtmsdjobBMPP9
SQvvCm/4cwat3gLV54so+VYRFO2Mlp6FysCMe1fj+TllklZM0pw5itMS27Vp84rCc4dN3w7ysYrL
3IQ7RX75RGvdz+ublnpPOp0Mrky2DoU63BfoXWhBmGuPPKdJ+K2qgHdKhhyXqoGd4KoRqBar7nW0
8MsI5+VDNNDa/HniQG1Ogh7dVTFqCw0veohJUQmOYSxuwrl4jrQcQaNqrQFo0V24Ft9N9ry5jiaY
fc0uP+kF8fdHynu29tfjhu7bYwU50UenlJ7E9Y8TKhJpt4+T9EwnOaTEq3j92M4eaem17D3gkmSy
t7qnyKjw4xJz7vMx595fFaU5Bse/rfMdzj7lLuALPYy/i+EJ7xA8O43q047H5AZHnY9u3R1PWsAk
wphiEAxZ8rBYapgB7JuK6468qZ4OpA5K+WChS02XMkD8xPYNq2ur/hDj5Xtg4Mu0jjPb6ijo6zyY
CloAw5Ze8y+gG/BAXYyMm6jcde7rMhkNjhbQBUiNiZNrQa1d9wE2klgU4wRNN+YLS/h6KHts5Eob
4DvNcs9qW0uhsjLTllAircvthu5uq2YsB7bCiiYqBpSEjoP5wjc2WQxOj97ftziAbcNt7aV9mQ5+
gqvOn95aAlcPVp03BiEkKGQ5etCskE135rnRtnXQfiKvgvveLYprJl8pPd7yL8kNVn+OWhXtIIH7
WvQ2lg6dwUT/uW5yyCejwJiIo7ytRIfEAHCQMOzBl+I9yfatQyRu2laxcx3vlVZpkXmzJhnIN6Ng
ivfl5HEd6FIXX/NTbXxtJ7NbdPJHjKnaTvWhoAmETpvV/ShGMY5t7u+OayRwhrv4VP7cDZBxxIZ5
tX4bukX548XklDrkNEwlSnrnqHJ6wkm4bthgmUUITEwXA6mt+4dzMVnvjYr3ve2/uO3IqD7u66xl
b1Gz8ffl4zuFbPpnlwZzrF92Vb0VkfQUzB4Lq+htQh4N/MskZFmk4DUxSR3i420pvkz335W1TN6Y
aVtQ00TUSkr16GdC8XGynFNPzVYUEvoCb5cd4GO+BjcQXfbefbyGVWrxGbuT3alU+9Wky/+LjcVK
gJRXjR3uPWjYoDjQiMsqf+eCNIyuGmoSuvv5jl0kkoQiahjDecLitwNJ4iFn7qD3+k9vH0T9aXpy
kGywZAUHQ277lMGzJNplTiytFwz79VvPWEZFHN0+HjRfogrd2xnz7hW48GcGnWF6Q4s0tGPYs5Fv
qH8+F3zMl1sYFRxtBe3YnveM5is/jg2AZDCG0qaQ4ZEqGRq585qZspFvcFSqTdHeJshAoqGLSwvv
v6RXqlepjXBIrIMOyg43Yj8xgn5tYyz8jxMkYqXdlAdbHkopIOr7xK9oF+oYVMeaaSXazCaI9VXH
9To/D3JgDwtDuvQRMRzRUWgHyVFvd2nnfpqVB362wV0R8j/klL2YxjPovuPuVOeHX+1aPkdwJnM+
A6hpFNabnJTI8dOjInxXzH0izoXRZO49BzPW0n0VYQxfBGIlGRa8YhiyBc7mSMCLDWSLmISbtKqi
UkdHD8J8xpPV1D8apxKRkcNNPvCZgqpXSdJtfm3QaHcwpRzJKvyqH7ooXPG3+Ux0B0V58YC1FnYv
VYz1dybtBJ5KqTj6M9t6HIt78G/b109aswP281GRfeJ1SKyv+6aMa4JrLgKZXU4IHPCCwnhzQ3Xx
zVPxRiR62sDCEcfsnkRooMy5afAFmuYb9oJ+tKApMSP6DytVO2h5kjazVyE0og8qyWEvbHM/JrpA
zXLnYf5ERXW5Mfx5eDH9q+NsbytIi34T+88/E6xIoUg5+6tHPqc2n8hubzG6FNBQozF5WCs7ZtWm
KyINLT6Vl0qKU6+gI/ZHz93tTAqqRRKo08d7Sl0BRFGRwpnDP6U1HKCJkhkdxYXtyd0JKjIRS6vY
qP4PSdqpXOgXEnHQAt4TDtkDtv2Q+PD5Z6fauaLhDx2c87lfISnF5bwMrNt4YBm+g4N8L6r/XDwG
GmClZmwOincHvPeGq7l5gNJglYuwYQ+hNjXqDkowPAwDNjXLbbinYDdzI9cPjhkV4JWE+MeVFdPn
s1i37mFOROMPPZ6k1gQfpjjf6KvxFkAxsZdiUNcaLVHaQba4SSoz5PPwYw78Q2m1/9zVsT0+sjfe
aU0Dh3NxfcnbcAkI5UfAvPrN0wchOlr4OlIgWGdZJThSFwrdCobZR9WYL+ARviTGKgSnChYXAOE8
aljqCKr448YHngSHlpe8g/iOQCbHCeVMOsfCRbm0N10yyeHQlGDyE4LrX5Fgc3el+CXpe3fzRNQH
kmIY1OJaJeMO5fBLrgaXi0SLykdB91r4twpsGgG7zXwJ1elbq9qCIJzqZnDy7QmaDE4qB1+XQfs/
kepukHEII5mPAHH0orjK96qjIL0w8aWQVpdVHY8nGeZ0kG+BG73zU+ZP/6zWvaMlrerSTMWXw28d
1y/DqfQL+eEfddDnEa4UxS0TnmOgbpDIfSsREGqrH0G41YpDVupEyjBZG8SrNquhKlWHmXLTHDhV
RISLD0XZw4Zc5XLc382DxpMzF83a2s9uIjQlklT3hYgVBlUFT0Z2EdzpM6k0mXrzrxbBURhyi7Bw
D8TjCLEFBt5ICeFWYJKeH7lyMx3qRvbdBdnf2nzAhXV6tS+SYd4LPW1y/dTLK6NnfAaF4lqtTSL3
W6sZlEqC74FdHtb0xbgYvokjRwmzOVg/XVUgDmFaWmRERmv/B6/JMaSY4x5e7LlrR5m5ncCv+p7P
ZF4xVnRVAH63E9JoqxJcJMKfRh35XaGXyy6CYY1aPMDD4rwJD9TVt0m91lVPIxtwwaRYbJEdXfYj
J4l2phhWgovn0s0Yvidr7gsvKCMV9s6OUysYVebdgfNkZiJ3MMhEv+HkTyNjWQXqjYP52j5fFOQY
r5b1gqQq0pNvDBYsknXbFs5QkYYRvQugLd9b0s/9fznVwON1IMbTJOur+Eal1rftuLJgMmMygTQ8
CLO+pvPPTB9iW4m0m9f9aa9zwZR7n/tso7LcRsyU7lKammTVs84fMVmbwYiDC3pjv/WBm3PIuham
vf1IapgK1p9yToiqOcTQXcjNRwXwERkZt/bwCSBVigy8vcx4h6g7uDCtFcI/3pxqECEoqhztJH97
Epzk3NxnA3SzMIjgix194P2bw9vAwJGvoiSNCcGqU2FtOssWqbMVYMpnC38zPZS+8EHdTgbvHfEz
PnWaG7SGIrShzaw5oLWFwnpvYowoI+JO9JEP9QzxAgPoEooZpwi7y1G6Gfp2tbZu2fo1kaRfuvUz
6esqGP2u/lpgZFECbjcsHQmKvgqNePt/TOGHev8FCotqwM+sfni4lnr+r5bRYBPmKeb7XUQ/7Iu9
9crHYMfoXpfZetwlKu11ngaT/TYV98PEg49OtDi3RA27285oBwI6exqF26kbRr0s2wYtAVOVMAJl
1U1+ScR+8BwKsAXYq5X9jk5X5aKlMgS3D02DSpixn7fAk+iOFKyeG9N1zjBGsM5IMS+FzCwlx8l+
HoXjpHmFjWPsdH/o3L2c7HCVMovbLIzkrbvlRkZI3CNWl/wmKOU1MeMiWqY9/W71UhH/za4UVY9h
sWKKX7J/Quej1+1rXZBKtQWUkQcSXRrUafE3IMIdUbcDeVOtHI+9uNzJaRpIj2iGgJVhWGeTT25f
O66eUEn+5OBogYAT0L26kTsffagHeFBDBE0hDjO1/PKCjRtq/8nHxjljRD9VaUKXSk33j1gGukyw
gmYEKfd6ZZAFI09X5yezGEibM2/lrZlhYNUYJ/gQWiSKnM2j0hxqe2vZrZ8W7yd6zsQkjHJeVXeW
Daidp7ATdvT7zrTDkoJeSBhJ8sz9j2iIlftn4rj6ibiTxhTLRNhKMTn95iqkAZOLZWyWPQ6nsc3A
XCfiaRBWjHURHFEO3JqmiaR69ejdf7N8V3HOKDLTZuw3U7NgEWq9Ps9Oo+vEMnOAScibmvQnM1NB
yq8my7FUlE7ZqmIdl5Ylagpf0uOMX5ZhNkXLG0G4O0tG/qgBQ5zoO/A1fv5pRXNyVTaTHsT9GXAX
bxiFqTbJhBfKep6/y+0S2V5t1ERUSc5jjdCEXTAd2pJydzmjCCBL35GjVuXSRHJwWc8meWJ113tu
52eb+qNg0crvfraqqXLR0iZgm8DKPNtiL4WAQqeLKyh/ikQY7DXWhJvxyOigUTtfc6Zf5P3+cPX8
BjEwmQlaA0vfUfo2VltAXi/K14ZL43nEG2MVCjhRNhRmGjcUr6e6NGEs8GCMKoQ1QCK6Ytw9xT+c
ZD/qZJxbDaXIT7Yy7f7wf7uqFb8gWZN9c3qBlFVR+JKPCh5Y2kv9MCCAovpNLB6U2IMgVu5KpQId
KIodQz1vrjYPK2hhfcO+O/CDZPctlrwm4ZIFg/o8bcVrOQCloyTuYNUzFi98Y+MvNEzaOaItA4r1
+/Cga/ibXuOnLPfnzHHk3pSl0oXBdD1ah4AClnY4Il6Gg7Uwpe811ksmWCXKp0zyuufOppuGDNv9
8uLa5Z8J+9DBEdJzEh95aZzzTJ+fg2CjPaHjCX80WjEN4rSNclIOiFFbYQFRMI7O+XPXE318Nq0z
hlsB01FgyaCeJAA++DqxABZ7XlsxzCuyxam/vNQK1y8HIqAqlPgZrk56v5Tu4Jaeg3tP9PbDMi/U
6AJzZoJBsxWE5q//4ArhChwjixfu3Ywhcm+1yQ4ubW6ZTgkkiV6UjA/ma/skD5DZYKSDFlPknnQQ
jKUIBm6f4CO+5gpYTqPuECWaIkdkZjhuF62U28lfymcPaQikBYphSz8/10NOw4p3ZI/ZvwUNhXQV
hB426sgCer4QLkOEMHj8PS+g/pBUSdqCXnSZ4xm/sHrbaDEJlp6aCMey/FebTHfJlqgdrhU5x5tQ
V+2dyJAp7W90gwtAdpYsEJ4S0DMO1kFgjXoGvK8StHwEYgWCIcPdRn40x717q3G5ZlN6GuksZP1o
xdigDkTwiJNm9Wap9uT6/mkTQ4DeUSNHsJb6OUbIIZAaFSiWgAZsqq+GdN+qT1NrM7S7fGi7gPjW
apCiEv7EkDzfy8luzDmct37T3LXmnARywlGVEhlw598aLq3Jf0Id4cMFS9r9YKXco6+uLODjntus
ibOhX9RaU/id/LKMLFx9DKPDhASQM7LVDDVCOAbXe4saCnw1kalMedO+KmoXVhP3jV4t5tqw3AXk
s1IWXXWtH2jUECg2PNhAZoLIcm7LR74WEblkHm+T9tSk4xwdJ0SseYuj2f//+1/6IrtfmjT0Gqj+
3EpL5i2sqEPfcPC4CcdFbM8jCiDptaFa5r2/gBXI+f8vSktDHe8isSZpV3hW1F/bxU4zPccswt0/
koUwPzARVwPAXlVA9qG8x8IFmJcEgjKYBlhFXPMB7f07QFqkh6LyYAuYSnEGl//Hr6uLETDSWmCA
nq2xAukGR+iab7bImccgRUIv786zBfzTCqDQXzOv4k4FCa72CdLul5o1WS8LEcGlT4msevmq9UGL
cNqjF9blv1pMspc2i731aIrzQUUYg+u2/MD9RC+6ruKhbXkV1d3OjXijsfQx/Y/0kJCkVf5Ql70W
DRMtTumNW35ADBtr2tERKDjVK8N819ogc1xRAD73VPbxtgUM0W3bzpslA68J+c3JUCkulQIpohVC
itIez2YkKXBBNAT4PWGs1yZANNFyIkmn/G40Xxxluom7Lmnt7Ixpz+PMNiF12is9L46DFMXTe3jC
FkHrCKL4TNwDHqY0XyI9carN27NMMFyjPdqwWVTSUB/qqysVsrv5LWqEKuky0UobKlVzyBSvv1Wy
zV4PgL71gb0RfzscpYSt4/lvJR//wRYOqNfipEcYVhCbyvdF9rIpv0SQSJtdauTZRazUJXCMgIcP
royxzPaLUi7/hnxD3HmkLytjH2u3dF1LeVZdLB18enl9pOQ5YSNI3yuxhCnnQG1hck3HfGuTr6a6
wSvWzz97DTDuGXmomKgSjgeHqHdi4lHhuY00ErUL81ZSPsS1Oidf27FKxY48lJk1BlEzzqBnoxno
6TrjMaBUvLfT9RAfzJTD/cUcuphv+DKmfEac09il60HYC+fUQfrOGZYXkwtVZ+81bWFEdVYTdH4k
rOiMqY+K63aohHZxG1rplYDoDVDeIFwjbxj7BJRQS7xyb08U36nE//LmPle9A5nXve8UftoBeGvH
vAZ5npa2yE9PV6xdUOhLHiJuq6cATfCc0WfD94dQX0qu6C96cXjSN7Vx1xKkFgJo12G/2e/WkOgb
zDQESDuUJgGlxY1xlUAUCJNjlI5jRG6BKqnVpe8CixsIU3rYG/AFQoQ9FTxjLlqYUEzadDNIffxI
VqsN8P3SQiW67arddUUahpN9KgtPQPQiUVY3iCGMtGhrxe5GgG3Gz0oTTHKrGZy1I5vnT7bkUAHw
GATX9CXZD9zaVyGz9FwdRZYmQv3uOAD4E71VFgRj5B2j1nF1DQeo5uFI5JEkz2r3THezVFlpmZxH
/7jq4WYO9DPWwl66mYBiNalGJZFGOeiCoLhGknkRYWoInArD0HYvgpzkd+B4kTJZwjqVUXaL4oC1
agiWodF36xOnDY6RmUAlPE2Lh3awP+Z6gLT7guBXSF47A8A3r5yfKZ1D0YwtszgEvslNmoVosvZe
xhJsgu+cZO5ecCul6UBjLa8ZEYkowEPrHmYh+I0Ta18eLfWWg02/eNJVEBwVrHYcSI+8vAOViwYf
WlzJmV0yKONr0Xt/7EhAR+Ae+NTRxqTD7wmneeNPBnqgbjMldUsHd8f9X87y9sqMvDYs0TBvBmQE
AZ1EiSymlA+BOuVmRBD5GS/NJoIBRKhFZ1hrwMMgVHiw6FtBmCoWB6JKN25bKQpkgx2ZR+bfDiot
Sur+HgzptxbJ+dqnLi5S3lY7kReX57AuKJjGmcYggdasmtEN3+uoQqnz0OTddXVT40nfofsCmWxi
Y7c4f8HuaAXMiECVZsXCepRBtMmDOw2iCn6Yy4ynncqZp+PVOazfzx47UgeElD3nlIfwHDMyL6M7
zeCyxhnj16nFeiYF9Q5859GX7u2HeWqvppox3VqMA/nYnzV7w0xzNyjnfVLr2VFk8wZPkbnYwFSV
hwwtEO4jbbHiMpT/oLnrmPPABXf9YWSCL9IpQHKedgzeLPD0hLLp52a8yumi4YgpjQhyenuttxrK
T6Semf0dyqCJ0Z4AYRuXls1n/X5sMP+m5B+Vs3DONH5fBCS5vMefGaoydUU0ogeHycEyrHMciE4b
fGhJ2HgmmTO6OAUuyxveDoim51MVr9akDbgKJyxQcVZH0YHty538Vk36JCU93KR6CXUguIy/YefQ
qepmjvaDkjOt0GXHGd4280ezlh1+hB+f/a4JDQmGaa7gJPIFrzEnBNFCYSy9jacpCloX0h1nH/i6
G+qND9yu1xF0kRm6AthRpi9qGbotfdId8X5JTJSZYrMVguAdvWXVZYsCbbCCntP2Drm33wkq2hms
4UugdPPaoLLy91lt6USjYeI43deLrNk/Wd8RhcCGgEfVQe6Pz09HiYCOD7cMg+I/nBO30aT6kr0M
AmsCPW6x+GD57RpT0GsoAKC04+zHcbdBitAuqLvXxeCAe/KV5rv+P00GcKrhMR4srDrnggtksI7w
CM1W94gDXO0OP665HUAayhtYDsnQj+Qv0bj/4uHO44blVFzKTmrqspNTmIug8omEr7RpKFRD9DsW
d8ybyApXBipeKnB8iZav1s3TlzyHim1k8+sjoUfgMdnk/JBoH+33KB1Guzgk+7Tu333EB4K+UPwl
MSXeQfSNn4JO2lJl0/m09HfpbMtVE2d1Qp1fPQjYIdXIAez1s9Zq5+Rx2Z295YbUfjZFouEgkdis
N3U/dTK1i87SVZ3CedVyoiH2tll8NNcw5DNCgC8A+efchycD9q0snWEjXKL6Kcgg+u0o/KBBlqXD
wMKrnX1zPfwcR3S95QjEU6ecV3102bL51VaZJUILAWrYhGc8DX5be5PsJsbW3moI+XDUOpJBQjQU
G4JEM2Y7MX9S9ioUL0WyUdngWJxCOaOZeCOxmK5OVXYf+dFzaC/abKndk3vY1ZPQT2YlMRilt571
zszShz5PsKG++g5OqLtcgrPAjGQ4SJ+/G7lAmuqCxqHGNQl1QndJrvMtW/noxelmD4hAnmySkRK/
F8X8HcB8H+JcDyNTVaPIHF4kALXrltVbk/6NAIlkhzGVfjKklA+Zj9Aies98ZVeRWaycvYa6hE86
uGhWkmr/ZtkFjXq2yc25mLytjStNwkHvRMAuYwHpYQZ7KiW/HW/2fpBvCo6sKa+Fk0B6srvoSpCY
nyF55S3UwgPkzRt+GSM9BXSMJ8eW0FM1TQ/N7jgK6cCyBm1Bp/AvDGzSU6rv5orSsC8uNwe8lYzY
3VkT/WiKGaO6QdC0q8BEoU6omhP7Xaakts85qDJLLevZZApRJJmsgjdcj2mBrnkJhfsVxJY0HWFp
lUJKnOAaHGeuz02gz45Mm+CcMj+aFowGXkbFveNbejaRFDi6z4Jhr6ITfS7czzcNP6z3KA/Hpf3t
6nPzsAqFYdiPGDp+Vc/b8l4B0qV4/XdUP0ig8lhBQEPZ6TYF+zE0cNIOKJZih5R0eAsI80w2PaaM
LvCklriOqSxdZ/r/zXzKGEnpwWFlH6iDkCdLWubsZ6ikmymmyOnz5dvlOBZLm7tIwfA6nPk/ZH+P
CsRqbebDti0oiBqPuaJhXuqZaK5JB4Lh5MGzSVc/jNTxpnXzy2MyKp7ZlLWgjIDDich/bQgkYdmy
5r3UHkZQLA4lrzsKqANVNfY83hgZZl7Qq+BH8dZIWKTDEAG4Td3sUqueCcp/4z2jUMp4jw6e0Nyi
YdZEvZDXq1ymChHrVrhXHWCXmE3x+5Gr71iohiA2uQpPjDTZbabnf4nv8p1QprGR94KQhauRstRH
ZLNOmJLNBH7i+SSN4X+KYjk6mS+G9eCRVtiDxFlRUKJmghcII8RVcKM/zpjpUu+rfhKWiLTMQIe2
tE7OEsYBD4KIkfBWB+C4XrEHYY3A5zR0cw497nG2bXr163C5gTK1xeON2uSd227amolQ1bRVGOvB
jOrqQLJUoeBzHJ9RqoNXWZzqxM/19H4Ldm+XT/9eHavsKM+5uOm+AnI4LpACj9l4BygynZYz8Fl7
KtjRuxd5kJgKCHYc87rRsXag/zjcYLBAgbVZko1H7nv8u/w0NFThOTA3mgfhbCTBrgoaAl2GiVH8
sWcQfkRJH0Y27juqkOn5v+ejtcmKPILdCdH8LC1aUAKSgvNFVXBr/gtH4aMu/a/B13CLQLOgRlwP
Z89cBhBILZqCsTiKMqaiOafpJKheq1aIgw9TcB3nqMYJ+qki0KMZxjcD/9aSRyZLF+1A1rey1Bdn
tE5hKvG9N0q5YtV8CM9Lo4xVoIAbvra751jBWS0O3sDcL4D8ZhuDUa/8BPNsnxH23MLcxKlRh42S
0b/jykcfiRf3GvzN+N0nuhS3aVi4i3aWNbBQJCjhXXq4bLLI837fAzXRcE9xhifZNyxzeRCp4hj4
oCy3XFXNqLawV6F4GzRS0Z5pNtEc0rNZdhhA/iEwMmmGQbOVJaIRTMxZxB9zoIg5cHUzp5pPReHP
V3FxZjXiM7/nyFzpKqYmvrUdq3znEMuN2lRjkeQluSOvRPPL8um20/pF+dUy4acBVNX8XtWXfAbX
XsRbDkxj8or39k8b2rJPcKN9ZjRVC11Dm+h/2Ns8+WMVZWas0lre0JNkoJiaUfYVLkDXVyJktbs1
Hz7cOM72y4z1Zz9wq1XdzyN2OXJFNvyD9ylv8fslI8h+i/Oblys4oa8/yEOmqqYuWrGsA+/hCd1f
GwRi9QE/wohERFIaBzkmllkJIFE1LBDzhLuBsUVZhjZX1vubXsqxjJLHDIzMvDQSGBX8ODRXYMD8
ktvdJweTt7zWSLEiVyW2wyw5MjxJYdg2d0hBE/QiWL7sWlE6+Pm8G3qtzIAeu3saXiY2T/MVkIOU
gKUt/aJylo01mfHxH5842SUB30R1hzYjkeBWi6ASzUCBUVW10SH/fce7YH9hl6d8bsKM7TjDa12i
8ovC7U5P2I28JM5bA39tWJzK4Etj+Y7WyOoECrMvtQYpn8iXgKBtf3hx5t47MuAaz5kletfZknmG
scc9uLvWmdc/cJGpZSb96ajxeGfF2qJUjewFpUnD4/8acdqxCz15ZNCpoUsGUTXG9zlfg94qx9uq
e/oEvdh6TMcC09PzRdNS2NXtd/Wn9CxmHwu7Ki06mE7TP2gFybEgA2cWMKTOtBHOy0DbSULV2vXq
2YGO+4+IcbTP0Pvl4mkTg9woDtj3Gy25dda1HEeG7w2OmkmKAwht5m34hXAsiWzw0YdRMbfwYdz1
TVAWawH7v6jFuy5y/FSUykSR1+SHwL6BuJOqY5aNbhSqusijqUjR4zo7a5NLcTu5CgudIS2gLgom
7A3CqIT79OSFQg63gbTaA9cpurT+rlE4uTgsHNqmJmhyS8BdtcPHIdCLDxGL0E/ijdP1jxYnPWWA
WSOW7+Fzk0phGUEAC/F14xg8GHUDzoQZlJ3FIMGpe7OynFkp+Ezgmu6kXqv89ipGqjDfHel76oP7
O0W7/kGN1yfghc6IgsSFNy/w7cbSnw5O2jS4j1Xrf9f0jmuJJGx4KLIKnl3uNOi15pi6E7ACjtcn
w0fQTLQB8DLV38c/1XaUtHyXDTW6sWaVHoOoFunIaxhq4EpAUHxXyQQ88q0gmyDVDItq+jlAHs0u
5EGM2vnkSknl44WVcQ/8j+QzA1+JUN6iyevKvQa+f2VgNYcORwYCHk4LbunMHvh2aIJ7TxkFCXoR
VDgb1L+d8mYKMgTSsCwmN7gc2ZMmog2zbWkze38/o2yOAljj4Z4fKWLf/qdGR7TwhKbpI4XCTSzO
oK2RApIFcdRpVoTehtOWY8iMWva7UPuxZ7PZKMJRHdi1rHq+68wt+LObqvvPokHWmouM7xdni1bU
6Egp5Bj1DcwpUGfa977KDwrIRDUwIIhjod7qecjDBRcls/M/uvI3xw5SUWsAWvBkDZqooKd6PpEO
zbUk82bJqVXqr5alzUHPdzYN0FnK4Z1NYXKD5kav5FWUgikGSEcjbBxYLKq2KtcGQAcOGMvS6kvZ
IZNkQGCPV7zfqbGFdwifL2CzFysLoCjRzZvEPUj4WMY8uumlSj2+SHz1H0r2BfEm75ERjTqpJexm
AKLeijeuLXD0hoRp9/ELUsnQW5Qtf5upeoQ1jrzeB5UUY82v+GoWStyoi0JBe7VfbDuSWDG5ehDY
elAfPRERBZvtBf8OiqXrUZpsSWryiu5x9+/0sy5lT6Eck2R87i+jfaPa8DCmZpiGIMvgQBMSqy8H
MBN0wUX2DtYSr5ZgsAPo7M5RDVUu0V90cr6eySY8GxMNd/go1rcGFHXhFZACUY+Q8Sfqch080VPG
CIQK+lrD9Z6EaxX2a9Kq/vH2FwkYP24hfygsWqlmbsIp+Wvq2D/u2U/EZuJyf2T0m4uVZzzEJKLG
4PZ7CPh/NFLtVUgkZYsbDJTuKrKpOvhBO8FkhCDqY9/eNlQyTsl3unPgctsp+lRmAR8tqa6XggfQ
JaIrhpoMM+aLItYE2GTBLbd7nqBIjGeZYv5nzJ+GG53BEyQIysz5NSGzDBK4XuHA6aZJ8ZxP7pzN
KyxynbpesazQoF9rNu1rdKgEHZDGSO7SLLYe85TO9UIwNVr4WO+lE+1JmoIiYj/Skaik7BSgkfgm
I9L46zu7RuVdCoY/Ruu+8SfrPpPBijJFNvh6Osxuw/Tpm8COqIGVzofXflD/3NFw7mTjeOHelM1i
bQGYyMx+MR2yML6TUZJeY4mP+QANXRcWqlJc25HeZDaBPtEB4pi+SYcRA79zYSURkZPBu+Q9Zbry
5AAUJBsfbHPsigCu08wtYlfF0ED5MFBBpMRI8rtzdDW6MJOY+pU11N4W6LffOcA2YmbN0E9H5FH0
VqFKNzx4gTyTvo3M4/PHVZ1+qZSiedv0eGS8P7fJ5ZikfSX/f83f/kG94DiZN+Lxo8VvORpNluF4
U2ZS1q+0tV1mKSRVylJiiqSnzpEM/nK6CDbx0jYcAQEoU2Wi7NwBEy3XSTT9hDE7iVwt3MGQ9Y88
Lt3iGZSXLHZFMRG1ipluOOcxdOaQU4o4TyxCUGjBYKe6+T8H/zkUlYpl+hdlhQNjzfE58PKIZAkL
TGdsDyv1SP0iUTUi6xCN91ar2N+HxCg1qBGaGQxyBCCXeF426RyYF0QvcSkxJSNXWGOyA6kASQ6W
AQGWsUFWGAdJYPy1THBerXpJF2Byl5VwQGRTiOCiYCFKSr7CdrIgf4V/M6GeYkeLXIyvbz3x7LE2
VTYMF4Ow/JHqqzs7LPrT+2RbzGQF/oPELT6Grn9w3TuQLasoFwmtD8rnLxmwj+PT6dfkRqnpegAm
8pufd7ZDzqPAWoKSv6Yot5/5ecNQn2nHmRxiQaMOGxKKL0f/B3KV+aeySMC20ldPPDmlXblFzPhk
E/g2UhcHw8lngwXHfngES01zIGXwpi87fiRC17IzdDKwqo62fUWlG+Yzs6AvOuyJSRoo0h1vrUQT
t1tXBpOCNnnKT2KB2VwPOsNWKcnoJXihvRcSUMrSvVtFJtH9h8rGucNnqMmBQ0Z21877wJBg3x/g
KIyakt5inXOKWP5AlXoBgk948FzxqeIP1W7B0ny2+ANgm+/W4Jsz9qevbC1s/iWXCe8EX1X8ycYU
vFdAk0fyeM6OKdB8ApI3TPnXlX4jd9EC9byEaBNIi7axTrou3zMIyOJgeXlUPdPrugORf9CTVapu
P8+IFWiAGry+7MJoMG9F1h8LUr+AlFo5g69U4Odd3bp/qX29ICyT4uRLdRShg+wCp44UTay0FAaH
ZHZphnRkQ/nZW+eMkl2cOXj9iszdNGw2HzzhzTIIHEKfAyUJ9dNH6tCnmDyC+H05dJW1SUv7FTnt
L4wWoN8I9yOkSXSYw6dS9/44YOVa+sTWdKXjWh4J2YDph0F/norMKEhO7qLZP3hSA6XhOiw8FQI2
v+fOkf1NGJDbQaL2b4rs2m/h4Wn1iyIiDf4oxvGD20xUdTnqaSuv1TDmjpwMjXK1wj//uXHqTQA8
IxUeZbdssV1rYq3xnS/LmK+J3QroRo+fLzUp/GArMawY7ImSS89gY+cpVvGcmKCMnyuUQlHc4MGG
TyvPoGNpJc04RXOD4bbzrhkC+G0F3vBy4fXo8Gom7wUEP1MUTbcS/YdjPqINmLWV3ecXT1i3G7aJ
xvRQOQwua/o/rXem0BYhEbFfth9KuLYMruyO5iwAoCC6QH3K7d/c5OR0wCUbAyevBn+BVyb3pMTX
r47ZrKajO/aZCA/LgmyePDP/JhYD/h1l3zxg/9LpY4DX6cqQTLTZ4AsFR0EE/HvvdKwDMWBHW9hg
KQMbDJb9K2UllA+rSD6VAUJhohcvmQA8k73WCB2GDUsaL/LJb24UQjUVboUP+tuplSMJ8SBmPnMK
Li539Y89wuxAJq1JVZpvZAD14R/Pnz4LCSl/8uXmkZwUAfxay/+I0x9I/YjN1srSslM32ichztGh
1i2LLZ8gGpgWZw4YeM1qlL/wwmDbekYhP7msfwdLUe9n9KGrh0sWpvhCtJlBLMv2sMbGp4W0OVRq
EHRr0iyOeMBqzbtHZkBY4zS2TZY+UatXF3JqbKMmpQp63U46nmAi+HOh5/p+9MvugIV8kJLvoj6G
X5GjVLDM5YTLsJGnk1t7FHa0b4rkPd4Q+rcs1ncz6edLzumUrkNkTCeci1DdFHrd/zi6zM+UvqX6
LwH5rM0MSoIkBmBh+j/zJ9oUHO6mGZXjzTD0/UL0Ah669hvv0Nivy/1sJL/1BwCpieopx+aIJjPi
Xy0TG8rHnE+udpKZHwFdTVdbOZRubNlMsbAL5OyNlgKjAuyXgY+ijIlaVsFZAt6lhKyl0cEfW4V8
ibPg0MY+VlN6pDecfuYRoPl5iB13HBPVjHJPtP4EIpBIURIh4zQ7DjQTgTlV56C4lzf2YcxTkKJ+
H0hEGX6e87ilZhen2LxyXmm8PMW5DrrC+FjPtzyY/F1MAp6c+MbXpKcXkfEUn4YXQ/6ppMyODhU6
31xYGC+YRlL9ftjEfjT9G/ami4AKfoBoR/79Xl+nhzxq9o5N47V8xlbRPEmbCqF3NCE6PRTPcRb9
fq42VbDCmT03d3Sazc7xei3wfLgtS+v5idOkjWFS9COssVHLfrH3+TTIP9SN2Bw9YyrbOD43wX/B
dz55sC+uL4ftIiHAs/28+pmu8CdOZxqVf4dGSmRVCePFrbDSAOpHi2qdCMCj1KkH5KulSBXI3qI5
WyNOkURamjr7foT1K/rANMEHx3ZCfVXGhMLrNGrOlioW6SUKg2vnkrs31j6VQWM1IQGng40223F3
fNVsv1te9Os1Dpma8d1/OSjaMUcLr2l34LFpNjTEhiKoFJuewJNWTMFITKlUotqKZY/BPNv3saVW
ygjxwQ6ENO4AheX3MVx7VhNU0CnWeLU4jiHFd6PzffsxcQM652ZTf8gLMARcy8V8DWedJkVud8b/
tVqa5YeAQFb2xdZgWG4ytI5IYAikR4docQak9kHMvXhDv79X/zFevodhi75QGz7iNkXalpS4aPEu
LSWoqMPzVnAoTzbN3sWHVD4m01SUH8b/L23i+OXHPLjSBfEgbZzazPU+aUO1PyG3WFrASewPT5uK
5sDMli0JfdleUkStdt5vz4JByu3XN6uk4IOybnkoW2e+smFdstIeRJwXOpbgcEFKm3Qt6410PsWo
YTSyUTFf1Yeyor6zGmGgXffavT00hDqLi4huGclR9D1QRAVUh6KjwFWcG8xHdQRpnI9fZacf2ZXW
H9UAYEFKETwKN10zJgQ7m51Nfyq5mt5ISQ8O43Kr9W2OWWztqv+cbdSIsktbwYp4mfsbOty0xV/r
qnMLsqwK35G4FWKPAa3wFEx6i0UxCCwAZQMgLn/JriYgeC/fICQ17GwQrA/Gyf1hRsNLhLBdHWiR
Deca5O2a/p8Hu6iV+9cYdVZTeasawwqNH97JLBhXdNuLaksPr1NkvDX4dDp5qmnEKVg99gXwLKxe
rQi2oGRhQgqHLL3mPnHnJ+okyhiz6E3vhTHUqzaU+YL019JtTOqGuPpJ+Sv8KwWoybtkmf8Jxpg8
45SHCGKpc8LEK73cHAM4pMwbGvbmf7sM/RBX9hzngfeP8JfPk1C4/KAKJCOXvqwR5JYJgQlQ3hHn
UBUP7nw0JxC2amN95hBFCVUiXsOr5Td1mG2kEozAnXWeihwYOUTj3OFmm4WUEEW1Vv6zRkfvW6dT
1a1dJedS9xxETvUpIscb/JjTpYxickOJ79p9Jg4/OcXDkctq9qZhnmriBO3tK66tmMWcQ4QEC63j
Kw19+8lcf21BXkh3rlzpEtKz2bVjYj6nZNkYi5/jGYhqEYWIHZyWxctpyxFfIbGl63AtsizES9xY
OwqWoXkeDaazzZpqRD9J7W9rcQJV7aXCAfibMXFydvvxxYQf6VSqzNz7s5hQRLhWbJp6396zT/9p
O3H/JPB2D06JMf1JAShK0QIm2zZ4n7kyCFKoyVo8/LXLzcPfWfzeGt1aGoToXlwmX5mvesiyhiBo
KW4DGR+yUcTU+ubGEYHR7e7PcAU+eBvzWppKZMYbVfeaxmQP2hdF0eFZxQanVij9rg8Hnj6fO/oj
cOTT3wXCDoJ3ROVsIMwNOKsJLLcFJmNgyOhlMsj8k9nr+Jowzkez7JT9lMxkroqbywll+DrbW8Hu
HEwho8JM5lnB9Mkt96Q97pBIiRLuuXFoc3hU0WYDI/hE7SDqkkvG7qg1R5eD9PUBjAzHphM5hhKI
kFY+352jTofKhEpD9HURQTYJMNwHMJUgveONem2OEaZpkM08cG2oKddSJTQ6uRkhEaPfYymWIkzk
JD4vvX+VYiOq6BroKP9NMHtpsGRu6ATyn51aHoOoSgF8zjuBtJ9WIdXUqE1wgFoFmx6Q6GFVdlto
sgH/n07/7cGoL4iMLRKY8DOdeAMgb5PzxG8HgIDFbNadz2G6ZcqCk1wNUJUTs5YA6EZJd1mM0aSL
MMeX+OVCjh6g4gH4gm9Pf+VuW3NHTHOq1k4NoOnQ9xhhpevzCsfshostlP2ix+Ka5VWSITfQOK8K
upskKkG2I5/D7SJxRnowcZlAU60wsQPDbqcnRm1qio8ax3ifPm6Ds3wuaojPgRkqfd2UEjQapQB9
pX6BpLnNiKCYMGEhSERdBWLJK+I3Ysf8BR4jAabaOAFY/lyyIxgorJGXWcIb9AERhTvZCfoNPNPQ
wurHFWR3YC+4UBn3kBivYbpMXVSZuD/39Hagm/AjF7NZZ4xVlNf7Qi6Iwhg84A/kOfBm3cpLVXQe
WZtcG5o+u5CcEhPTYswwn2aM/PU2qsKHcE9a8JiMeY/M5V5KVU3tRlfqj3VPNF1AlxZZIKjE1cBc
i4jO02b7vmAYARwPGS4sEz840CvEyqAZrtnqPaHaLNPVLeLCNDID1cBsA7M4SYUh43yUrElYHBTa
6DFYqRA6ObB1cN/tSaI7EjcrT31RN5zALbpSK/akG3TatU0IB6ET3pLmpnKTUPOtkjfB3IgXOuc2
hKLVH2vA2ZXhrOdZK9eVo4AKdJZkdZ50+wv3YEDUQuWujQ+jTaXfOntbG0pAS9rFBy3DXnpaexTa
pZT1aSGWKY0oYhgFXwQ8d/2+qo9hiuGFtlIF1MICA3QarsyT3fnzY9K4mI9Mf4sBmly5/RFGEVMX
+jaSGRoUEwpjscuoC87npuh6m7st079npzYbRYZ1Zhhx6TMrpquRT6FE2fV740efT623RZXEg/JD
K+54SRsSQ5DjfamrA5nM31v+hb6ynDuA4iIt5tKu1yqyAV+WweRM/ynBFJ7AciamzEiTs30wlqNF
LlY8K3CREboHvkZ3QA+yX2gDdpNbFz5aYe3y3F/krkXwSm/Xl1aqc5o551invDy2Vh37HmQzCd4e
UtgALFtuPj/gSTcT7+kF/iG98ZWWbr3g3BiR6w949iZrr1lGInjf2tCVWJ35+QTrx4KhDQklGBfC
wSNtGELpf/WB41ZOTnQ3EhWzk/dSCXpEjRzhZbmlZC+mEDYhJNGxOefwRcaThePLUBAf9xn80sfH
A6m9euFb1g5wbK7dyW2bLaDYG5wLvV0zrhNGciM/F+l7gYCAgC/pgxdOQKB0G7WLdIpLlYFNfJg9
NkYBg5zZ/IEE4JvuOKVLjItW1hgoK63K9oUrJ1L0/tdhywwkSvyI4VTmVSw5gwUgfjRkgvpDTY0U
afSUKs/72cqwLj/EexF6WY7zAQUJfxMWnNxe4IpVYXqeHbQ9lzdmhfBZpAWRdlHZqlgtJIZX5dSu
vDWpO2gZUGISyTVFKdF8/9fOBKIr/MSoHOsPA4c3Syi0A0iyD+MoJltVKMiO/2B5pruDvZ8j0uTt
tfmf9Vc9PMQRXl6xn+Kl+E8zJhdKsj6Yg1s8QkjIwO0xid6P5VPqf0cHKjR4vu08m41UShggtQ5h
WEWWl2Gz8PaVa3kHStZ45nZM2cGUocyiu4+KK+NokuKWpwkeQ3ihqUBRt/n+mBcd5juFar5ONFzy
CWV85KVPInu3VyIx2q+DUdgmVh4YUpsFZ6HVGAQfa6DBqJ5ejksUFXU6dBN3BdZKIeEFM4wbfxyG
bm4VXa+IRzus9nI2tx4+k8TbJtyMT4Fon31+c44doibAjCcnfRcqD0RgluaRbQYg/9BR0/FIXY/x
esUQfeE0zPfQmtCa4GYiqckWzcxTCv7RFwkIVaQq4dzKOqxQk9sodxRC0w2QRKvvRONumwb4JDEq
vw/27NXvFbkMJq7RwmsQHs1EJYnpr67lOCf0K+JQaJCkGN8X8huAuKFAkthowtevHdpY515z3+q/
xyYeR42zEqGHwC/gw8XgPNVceVemkwqciQFKs323CQ5OdNCwJeRJns2QK05vN7ih3RmnAU3K7AbX
ZGzt4ht/pD3L1bGsIEc0J1QEHU4btv4p9TNgqBsl5dtVOU+c1TR0WDgtrpMh9iJC/qzCwrMNmF6d
L6j8utaeD2slWQat6nR5Sc5BoNKpR1m9RKlr7sd8Lg8alVEDSnIPajheaPXxILTdOe0bJe3LcDqx
fJyRBhP9IjbIZULrXnL0odRDRDSyv4dRgecnGZK3MjUg6kW16FeUUbnEzUmlnaAxfnCtNNOgO7UW
V/WwKWZPLrL6KzomUOn1n62BGkiWzHNvzkok0p2OB2ZCj5I2QEfSt7Rob8REHYcKbAKqgin2ur8L
dwzHXy0XFwZvYSiLHkLPXGUcoM9RZ1iDe0PIJsrBOsigE1l4qB91YVNH8nnDw/3ZOLwymWq6AhiC
EyfeN5IWuuDCBR2bXpEVVmx6G1Ftr7XJzS3ENlqKtNQPPv9dKFaY3eNdjXnYVPgbhWi7TM9zCvmC
YI3UQzGHhqx9K6ZEOlZ5EptMWvYiPQdm9Rc8obaN691WcroDlgZp967ECDYqEuY7NZzMUDKuPx8L
/jCROUBP/EB20BkkLu4nKKMD74dAu82pZiZL5A+Z+YxQZHSEPUpZUqMfKCohFhctyPBbgS5+LryJ
YV8EKzPkySf3nlFcnQkQ/g4+1sm4vCXu5juYkzPNWgnPlZFLX+9y8BiGkyQ+IwRglFIYtoGMzYg5
eTVIUPoSIgkSSBmLDeYGuOXiQN0f42XTjXyo+UmVW7ymwvOBp9ypYEn1yD5IG/geldSdLWVqteHg
8q0+ZjGcE9V1ai407W4EAjhEZ2o7jHhmC6EkunUhws4jtr6NDEweT5U5R+GFhaDUIqK0HnWVhCaX
jVx6WotpsqwzQAc5ZPUGnb6SsalyYluMJFrNIPcNU3VocQ9lUmBLgzZmWWAEBn2vF/ZW/J/Cs16z
U4tUWoLqQw5NQEzlMp0xURZGmpU3pwMjjcCoRQV2+gujQymSFP7pRgOd6pI9J5RUBlcNJgPFIovd
ZTPxhVqt6XJfK7jClwuUuPbP5IffZb9ZkS5n7glguWTk5GZP4YJQ76GlqJQ/ePMDU9bsoGpzCkDq
h4BInRc0RHECPYez5qOcJrcP5Qop61e7tSPPi4L1eGbHXcw1PXvDFNZ1X3+cLHb8nWN1xpFEazOI
bMlE2bvit9/QheYpLzvV7HfJXPHWsLYGS93/TgFKlqOA8n3n8SszTXVIxsWtAiO0oQulalTKt4BO
qFAPpn///0Nh38bUwdrSBNJkkfCYd122ttWUiw+QzuFvLWxCdANuA2ck/o5Oi8dZMcunKdB2tVSI
mRDn48fBprxR69HYFXNaVmfvI9dPFWo0HXAAivsAelNqOrlgeIHcJuonYpuxPP0EZLyftKN8Nxwr
uro/yf4+R2gV/q1tVqYe1iVf4559LDYMCLzPrC9UBNSOLAxSJGJjGUaZm9aqtaEHzb7T935g3v38
9GAR3zGQiKKjtXAVQBsN/P58U7oCX7WOmAxn7SQ/dXeFHC/RCuvAt5Ge6xF1LFJ5LomhWnx76JhO
5CX82eqF9fNFI63jCv/7h4WCzLfB5ZVLNhL9bVlMj6UoGy+a8S7aXo7AoJyRGLC5BBOb5jUL3IOj
ciJG/AdZpOSFdAxV48XJmSz7TY424zH02cb9W58jEImPgovpahrzCXPgw+fFRWGI9wDKZ+kUy50N
zEvZ6eO+Hb82pcDqyxfIxq/11bsI+Lg8h/1OG3Kbs9bTiCfN4s/J5DDk0++9BvEUmsdJ/haM+ip7
PCXBq7S3Vxrl8QIE0PyapcZeucqhFXf2vQaYX3sFJ+QqFOeyB+5XJXWwzrT57aIs/SkVBSN2t7nD
af1MZZ048rVVPmLH564etC/r5xK4jVXYCeHYU8HR9UOIt0cMmF7//dJjkqcTNdiCInX7y80W9XGf
FU9vYr22Jy+Q0OmFIO3qDerWyfW9iZLWoXMh90ct4eLDdDlDGT9xipQ0k0iEOkJktHLxCrrpAtwf
oCw1uw5mwORxa19EwLgvv5kdLrcvpIVlHwbjvFoS2vyqpcvkjI6WxBqpZeDKM3cZ5A3HLxJ5Il5l
nPtN2Pos5iDXAHHRBeEPdxBQfl0q1Nz2g1KweKUrLSsPDiVzMfsPwTF6La0xFfvA5X2f1+sAjfyP
LQPE1gTF/kP6wik5xemvUOnJWaZpFLLwJobD2rRuSBte1RF6KQjXAiAPdXTbjutF+nXFMg3EUjFD
JwGyK2ECV7Mf6ctNVeIWnbAiksffX41ARK89dNUNfdzcLmoqgf//Sl0E5O1pIR+6c6yfSATfBuvJ
d+H3LD5F5WGy+L6/LROWsKbixgpfApHKFtYlvcnyGcnDDF5N62X6Vzsfav2DATvyd7wwYoSak2oS
R7Lz9tYronYrLTF+eQy1T20nE/kNiRPyFhiCHu0fUMl9jVj9QPAn93KzrGI5//SHF4Jp9+erPuCb
IPSsU8qmBx90+BFWHehMw0Rk9CniFLCKSn+EFZ3q7y0dozW7gGHouiCCD7xsXwpXopvc8FkKiTpN
Q9Y77myINGypulx9qGdGQR4cSAOIUsODNohbsO9Oq5amt2KzE3qX/85DcfXeQkiVSNvVf4DrFS6M
GRTBAkjYUCC9dD3+ll7/n8NTLUF1hkgPLyqI6zxBc63x1FAaijtBp0fD8h+5NMCTHrh/lU5ZxhdI
GcqTZflo/QaRkjvEEDfdO0AyVOdcN20PVRvcmDTVUa5bkZTpb1Vm94y7eWT1J1Petk1lVF7b3wrF
96OXbjy8GWQ9oxZjHEjSipGX1xZZuOZGMg2/Qva4EjiPknJX/rMX6hfC4AemZqOwXHJDU404DLrx
FadCwib6zOHU7eEwNrkgWSQYdDkIZY8cgEz6bGFMpirCcbYcN3VpmCMru8zP814hZb3CQH+0OV7I
UgkweMx8u9ThDhtCtEqH21R2UNMJfNsluGVNmCNsxOkz96t0KaKJB8C/sZov/ttpwS45ssDhhdlR
VVb090Lb6+aSiZO0KuGP7jXmZdZTP+w0ZPtaKnxl0StYfB6kNJnbiXn19P+Ltpww+y2YwiRzAgQm
QyDqAvT77nIzDjXiC+49TMc/l3nan16vfYsDylV/AV6OyA5w+sCVEduI9s5yWEWlKFym82O2yHiE
7Dbpqu6oVX5abNTmDT5ar/ycXeEclFHkRNYSCC9o7OtfExWZxD0kZLL2VaiNFjdtsKreetXv+Grf
GgzmdstaaMR4VCdV2QlM8zAzeoqAj1kH17oP79a77TdDTc3GogWKoKJZ8kX1OJMtzvmlY257Pclc
ht9tTWvKT2Vdz3u++v1kxnu072c9AaMyCHYvs/srrS4ejxVApgwitTP4Rqb/wx5f6VxMKpGLO896
0URqJjDPtgVwFyDAsbBce1lFXzoniOVhGffEmK/cQe0KilfLCAKHXkU0gACLILSfCuXkRnlHg/8g
/PnLJLEAVK366JWlDW/E9BgC3DEL5cy+TL3/Q4f/HNpZ3HVpTC/DGmfeEhZtGwoxmy3kowtnoDPU
LtS3yBDbj4KRY6AeGQ8FTY2el/GX9ErHJPCE+jUwPtbC+BvqQQZcGJ/O0PcwExAemnuA+MXIxVAp
NM9Mdy0q0vBCu2vU5NyiCQ+/3F+wkFvVN1khIuKhvYClZg320/Ob5LfE4nRcGEqgVDCZoCA8//qS
aA2rpj+Lo49zn5gtS5L9uEXGEqJVz9H7eyhSde0DX5/aCXc5OQQAsjxkJsG0zqpV2FAC2nWNXaqF
gzn+OBwqztrd4+CszXwCm7bsV5bEO0aMAVOhbsL3VTMi5XEjfr9/18rZlJ6j/XH1DRnwRX1cFq0k
YCvOLIZvXEW41qXIbiJU3ptDwipDwjjgn1yx9nL1Iu0cy/mUsT5+oFnFEJelEo0FjIwiKyIa9AaX
o88ZhcyWCVtXYpCup9/rD3Zh51ffBqKASDMHV6+g67Ze3puM+hVHUNcuYyWx3iYFw5ZdfD475QSe
aqaNLHSo6nRXKkosJ6+cFi8YxEKX/gV61xkv8fT38E2pshguFyypawnVzJ57HKo1gKJF5bazFbXj
5XEMRCtmGqtZ5iS8EsIqHTOk2J8f7FSkSsjSoEPTmK5wccmWB9krqAKghvhRT9IH2sQyNkahZf2V
SfrQyTkmNw++aTYbwxWTnsyOP+MNznEOT5ULNbdF0NkOFjq6NraXl7gU4YIJyaLZ2ffctxAAuKQ8
HIAZ6R9sfZ3PeBqhkeje3DoC3L+CgI0MmKymovr991J7uIzh5aYGKoO6uTTmvK6a62/XhiATcOTR
hJnGfqSL9q7Nhwva/FsCMb/d/XYX6zYcAovGxK3Y1Jbgu+z4tuB5WgsEZ9akEARAB2VsbXqEtwwM
HrMpKg2Hv8Kt3+kFahowFxlpMHVcYjTa62ZOY/FDPew1PLmUE09oAmNR6nX9Im2oNgxvLT2rHp9j
ox4h7R0AToIHut5O+gjl/XsK//Jz114ODagkSKunoNAjTuXD/TUW9TQZ4Ier9rHNuPI8VLkBW+0p
a+h4pxXMzCEmG5s7GQ/IORc7lkMIpwG6TBAP7rdSEeFjNMTghyxaSH6NM1+omEBic38APmnTLlFO
UxgNylg+tt6r0aJQqBXUz8ZJfSncaKTEcxOgI11VeulrzG6TUDtFPi8HBQ3JQ9xkuEjWvmryxCQj
XqGiZMKQ7eI6Qsazfr3MZZExi643bHR9Vw2nh8Yw1I0dhAsqZ3PvXMyJF0x80Rv3PbMVIphhN/Uc
OIWgkfvkXWkVQVKxRWVA/vNsA65tlra5xR0zdhnB5fYjLcSFvy5nsd68xwg6yQo/3B7cXyUftV3B
rnYeW1dAkrf2mEW2cERGkUQmbjgyzD4ZNq9b2mlgnIxgTTcNWWTTrDGdX3QHKdLOIOwp7jXvL2yd
1zT2ab4PYUjQY5OUWoR+uvOuG3lfGWBoVOj8dN8xmUOrCO8irAOwPHyfVsevbGspzrg4KegzLBhL
Py8xqZmcgk1pikk/vt5IpGyxI0VeZQu1i376LvT+mjFTolQzLsT9Paf16Bnr6/whU7Z3v/eeK4em
P2ojRtBuGLImcCZ8xMpafCMSEioJXRrvV0DG/8w48TbzK3YBwDVJMLOpXCk+n4Z+bvi8wg9HdlvY
2s+ynquTCJ/VAD80UOR6dF9TtWQf+pQr7zqDLg5QQ0Ii3N6xoqALwIbXB/kOXupaCpUgJDgFEs2p
/3QL92FzzVhDA47iHX0BAn2YCWvt2Lpmirh5Nmc1tV8qY3te/hA2F/1KgFDkwAJMwz0z7bVD2TN3
fznxE3iUFOMbVXBTMSgKXw7kAG0BbjsJnEYRdzNbp2f4q/fR4PCF4BtPrmoi9cDKvH81s5mzlkhj
uDUDnjR7LBSVZZd3h48v3Qm6g9HHpcdqKghOWbq5rZpRVKKi8COXPto9//rzXDjK80d+s1Pv/B9u
9KVruby2ER0xZdSc4e25jM8R+NWdJRxGZN3SnW7AKeHtx8MhdQ4RMCTjnQchmGRamD+WaM4nRJna
qDRKZoI0uIN/uNleEFUPivyrbfkLhIG1WbZltqcOAJfcw52Yy5y8f9wpLf6L3e2/XVpwxldYqhKL
0UbFaDT51nB1hjbvI9M+5acITuvVqGM1e+K5WsCiUzaieS2kblUWfMjlQKAdAA0SXDGjEhsGMFyB
vWXlZiTWeBx6eksIp/RjBfmn/ZhfGFpuVEjT24e+gX87cxFB06vw7d5ovGYxmfjZjwy1s0WOCCNK
kIOC1YNcdoBqo1+Wg726DqickixVrj4rSPqVfPex4Xj3TgyISnPhsB8aooBbSFK7C/Ub7NLs1Tks
rza+6AlpPATQpgO0gophACeycxgIOWgF3valG+h9j5m1vNtY7tNr2t1Rxgf4ac6BwbdIMooOizjU
c+nM9N4Irz0X9tWar9mUgakyyyVEoTCmXvxTS+KTQ0292ZQ+Vu0QYaiXG14ASgevCroPuQhGY6Zc
EF4N3IrY797xoxkpOPdsE4fzKIdqAdsBP/NEDebwUfZV3205qNIIMDDyn5WpmFLpaxb58PoOqvjk
BmtGuknc1T9yR09HHk3BIPkob9lz8arzMztjVp0aSjZBrtsBp0V+NEO0JnfGmSkgPjIYSmxykmdX
09ZLQyWLK+KNZnJC0bGcfwddLESEsZR4LS4QXeVjMCjMF09iG6eNu6DBGMMi9Rid/uUbCvnV9Oi+
EfYO4EPkdJieCGTLGviQPAb6RCKVUQjJK9tc/DqsWLsnX3VZca9zkdzcE4KjE1JjD8FEcllvWzfg
5iaFJ7RCf8/fO3fa1qyAJkaKhuu5rX3a92r1nxerokrOhuNabzVywwOng6xHUzzZ7KsaYPFeYGxX
GrbA4sSV/JGTZpjyaN1xm4HCvKfqjuf1XPlN+FZWmmuiisAWKQE9spDIiNUP3EwCwrCDO+1yWCUH
J5kfPkWe/RMwMEAlgYYTqgK/I+oYVocbgYLVJhs2+IkSbIvUIVipujiVrSQChb08jJpj2PM563AL
6uNDrcsSEo+N07LEyHBLqH+JyDzIvL9Fpd29T/0f84GKXB4A46jsKX/J/UoG7iPy59rphll4rcym
lgOagjwcTAgjBGhV3FxMIt59UEjN88tZQ83eH3RREWEMr6Wa23QVjQngjz3V/CXryVWqhVZ21a5A
pN4OudJUaMlxT8P/16JNDsEU+Qmlnl9UZULmavojvt7Xd0LMTGWyFj8GKZBuSplVS+9yaKXsVQZn
JdcbTBol1/TedK3bPP1+EgbNuMU/YTpKL7N5IWnbmcUQY5I2qrVPZuU0lJO4wPEu9Opb8rcs6yS5
Pm3LZ1DYQlhyrP2yEuBRXnT4ThioRwCnfcA1yfipA4gw9zHpLDfTuJIweueAO6EGTq0Pf3iOl2km
NaINQanzby7UB6N2QIKvWk1T/0ubVrlYfU+lLR/3mXCOGLJXhI7JGXSVHuYtTxWMmK5K3ypckDAr
BhKrBs2wzB/4hiXQD9eW6iffpSl7yQLAHGjq7bkKE+DS4foYIZkpPWIj4co85pim74PqOhN0WmMf
vCWEDsqs+w74Qox44A0UZ6AEfk+zX1t+2quRhLBktZ7wUQSJgskx55MNEymQIynJv9JkBoPs2Wv+
Yq4HjXEcOXaIACoI0PMtm4xtgPNHnwdzg44qleYSUAGQpBD+PxrZ9RJCMgg/ipeufWXiVDuIS8Tk
rfLk7x4gAP3Hu0lOcXSmjDrW1QZrqDbrMqkMoWgDmSNeFtkGCDiwkPkAaFT1Fjh8e6+2ZOJD8KGy
40RDjGSxbl1sJaF2H2JD2XLzLhFb4/jZfKz1d6PHR5Dgyq//gaHb7ccnP/z+pGiZ3MF1RK4UzNs9
P5eRM8OBQj1CVyouN6U/bXCbo/4sg/G1eXWlqwzmC6zO/vVdAmnRBtcjOhv6j233cQRFBEW3PPVS
vraqvUpfqdzwNjoT1KDxGNRchuE4dgH24vw/3AbLaul5Ncay96LTu2bHZJI9pxjXIbNcqIgM6Ycs
DWan3cGZm9HKCB1vR8/Tb31GGX9voB16c+H/WnrcryyVr2Z0ZgSLUl2nsuewKZoYa5Hh22I0ZmeB
B0zji1pN77fpczuOTNnzxGUu2joNJBbLIpse7AQ/f534EYFtQ33+uqZ4Mi+xX3evpqB4ac2oVDnz
ItJ91awma6KF6qRrxlFXvey0Vb0RHJwhyU4wvnYNUebVtRDZAfAz4ATdeGdsPCG7caz/tGfEIF+e
obLSShRMJwYoOX+f+X3ITexNu0NzrPQI9cXeTqRKm0i1YHdOKgkGvgxWZ3nFBP+LqTdWmcMF6MUU
HpbXJqWKoNY4UwJBTzVOizeM0P//XnjH/KYgqDye8DdEFN2mgd2rmw0PyDN2mwzZrhrpT5s4lqUs
d6d8f/ZY4XK9svJ8RWxGA0UzHbxTV1BI3dPyFYf7fwzbbICXqOL13s52llVYZX+a2RZdicVCIC6c
8SEzAjFEUYLxoCybY6UIWOvaXEvO6Gb/OGPpqZeixQedqAp/xkCqOyT5IqugGc9LiNscGArjRmFf
lZEVFC/WMp80hx3JTQxR4AQWjxfHRkMLrwZMk3zVIS5uoF2S3pmTZyXVFhhR4gZWXySnJRAGlNWh
Q9naWqqvkq7TFg8IxqEVyyUiRA2itJx1KJKZXLte61HLgQ6seNjw9RO2SsW+BM4MeJLCOi5zNon6
qjnrHaGrpVKTgC+l/W6XYZ7+s0mZXoAtq3Mlvcl/VwKNYeko+T0CrIfF+6TCWWm4nygNaPqjU+ev
3DQnfpLgp0I+Z4t9N35C0z2GzRrtxx8+7P+RWFzmO6I7FYKSBlQrdUKmeH6Pt9EXVtCkLqQaHs3s
0vvIT5ah4WU0dP402xhNOyGkxFutnHnH/jPbT+purEHeT1TLV/K5tS+DqH8SFnlaZbv7XAtEoF9p
nVOWKPi9oGNZQECtZyQHk6c0XV7uzx57osuVMZHjVqqwh8S0e0LX6GjOEn7ToiK0fCjTHD4/Fu3K
1NwP9zB6MbXecWvo7yeoiBBVCtZ3EB0ogl+X9dKoJpt2JfshPnpfQ+pcYME3zOtcCljKGrvmgEt+
4cRzgXkjZF7TDQONjma58vJRNfzw8NDpe9xUzIqEZQr99QsMOm9AlaZoSbcBAvbChyFJfly0FWSz
cJtMk748uKe4T6IN/8TdhfJB/vXswu53Z7Pzpk+wpxx0+2p0SB8BgF+eWQw3fpCo37TmpocoJuUw
rtTse9RQbeHnLAEztcF0yLs4wbh0B+pUjUNNFXO04TbJZOSxr8ioMeLNft+eVrn3nPEPdaYCoX95
XFF4q9RvSjYwdGfc2Jct6D6Z54WYGEs3/uA9f5rBRnHeMRUjm9C8ioBNVk0Uz2Kib6c533hBnp5B
hs5jUtGcUs+7KcqFG6gRSapaVUfX28C7wtanP4l+1czdHqw7fPnFmW25uKuU06OaJDXu7tH/6yII
IG6f3zys5muVUnDhtJ3qhv8E881MzLIMUy0KwfY6jgyBxi3nD/LsSQDUGmlJPfPvYdd4DhxbFw9A
ya54BLgrZcdarsQ4jRCARjmocEE48X2gqTo/WwXRj876/mmatlDv1wlJuNe2DUlxtFKVtZ2whVsV
RIs9CF7NpiTSg0AxMRRn0q25hYYPKRx/98i7ZmZdjEmqedCBYOKkrDxBi4mp2bbLTfeh4exLJBwt
wqpsli8yHomeXsm5sCTuZXrRfXu7i/7Borgaa5hkr/P/XaqSOkMkykS/pO2siJ3X0QPyRWp+DzhP
S6/gKpzyLgmMW4M8Ck0GYt4bhfzTaH4VVWoUEvaTF09X//dFaORu0q6Lt3LAaHvuGbVg1ARAbJiR
9I2hJNuwVwYvmqJrs/XMZKGS2faVlzIYL8xxUZqNHqdHs22tFfHGGyyzjnmq5MB23CPnsjsJyyNC
jeIC9uhduN57GDWiLPzFTs/9vj8Q8Ese58Htrz/Jl6P53no5l0gmbVl50OoUdrJ/i61prBcZWNLQ
WNdqzIs76tw2yXNh+tzoIXdqDJ2yBgczewYRghEaSD1NGGA3fUU0eFOvyfZuS9qNoQAvam1ZLdhm
VcwzKbdUguJH4c5SwNPyxMryg51CRO4SyHkJlFK1spNmtTp7LouzplkEt6gxdKVDrtiRj9/UF9Ya
GwLDVY6s0U+sjqAigF4S0OVAm+k9oIl87MmpogY38U7vcoe9AGlDegKrkSrBzKAcUacpIpI5QzSS
YpnbMx7o2912FR+aNq8DR4YMbjxTmmJe8Fdv0aZZXxhOjn3NMi7tlWQIw0Y4rSSIhmFJj4h9FMf7
FFMIL25Se/iauQRVoLyIJXVzodRUxmNULEJGiWbzzmXwjO/XwNFBLMNORNpns35b3ar6JVcC1GvN
bIrOUNTUK88rWx88oNkorF+rU59Sb9Ypkv81Ek31BGkS+dCkQJR+oEiflY4lQSZS5B/rh0x/8O3+
BIp2L3AgxCgrzZPhDvO1yy01aFhn6d+lzrx3xsqO65Q9VRuwe+Xf/SGTl1tN9bjsRWi35340yMOQ
cJO+41dxUcbCD2P3QzvyyB9ns6qKAi3jaYx7xwYukjpfrdRKZ/5XQlrE2YChU2u8Ta+uuRJMHm6l
ehsVWrVT9gjRsIg2efQrCUu1LqPAXdv86GyzBz8cKa+k2XJn1oLuQ6CKbObhRIQU0lojcyqF47h8
dQ5tEMu4vtk45i6XpalZzvNwSmeAKAnyQVxZGfHwbOw4jZWnhZyFkjHCuD/MrtNrCyLAriT4Xb/w
2qzF4VIArXbjGUZd07VgUxjZcNqx+82vDuEm5dClPYAQ9Y73wyfSzWZ7OwfV6gNzLpOtYU1H5qBv
MrO6yDSY60ezn6TLQPSz5TPSJmtp3UwkdHYNjr2IT3aGnlfopZtyl4oGsOrAHK2VHHv/S+BiOP8/
q+gyIyAQybi+fcquiObxYG2DtUM50Dp9y+1wldjfhTYN9P0EaUl0lcWwSg6/5ptiO4g2yfyQpKjy
W5FnIJeko59j2UklJqGGaLjVl+X0ANTthTOFvR2p8FgVryPHNZI/yKP2EKGqZ0KeR3Z0ffDsKjhv
GpGwdpjNndT/dPWuDDutffjs/0mH5b2YL+fl7OyKlM+byIqAaRwY5B15o3IjfMqMOtD2PHPzq7yp
ChsBlL9J1feaDCSqDDP2w1FWxGLH6m5zQ0TCHOaSJbtLQqgMc+Re1IdHA3ye7ZXpcBxafDAq/kU4
I/fSjnuTm4FBrcazeU8zhZymV/9apvykFVZar8Yke0zjH0d3+q/NLe2jc/Y/zoemMlf5oMovUcev
U+l1nOUOx+Bqpice5RyR2UiUO31u/cU2ZsPnZNcm8f3yywgJgL9JDvXJMrSkDYVbYq9fUblbaJqo
X5HctM2xbY31u6VW79KkD1jlfq9O+A4tdZ8OQ+B/WVsna7iN5xpK6QFD0u9kaZ8/OWpRLu1SwzlW
JjHJ7yb8dVIiagUl2Nhezej/QyALC414X0UTt22lpgJCewBKs9eSPJwx99lN+3d4FUFHG11U+Ek1
itio8WCnvQ0Wr1/dKfMax0lbaU0GF1OEET/HD0JHoeAsdLDXQiHJUJ00MINoCOkRR7R8gAek5JwO
f/ElKYHA5wPmD84Do4+zAVqhr7xSbc+XqmxZ/nnacK5XdAanJSU+Nd6kZbvkTS8j2bn/el+4tsGa
XdtuvrCKzN6w6ivOkK0uCSuPvKI86/Sj1tUtZJM8iGqP3xXDB1RDXXy6++/ASWrSzCHdXBOd9Ofb
hdaeQauIPTYRVqDgB3Siu8mXBrwWN8GIJ8SmzT6UgXt/ZHgy4vZPxtaIgjELkyBQlD3IAYSd2MHD
457hQ0HJ+0OvalW1Ev3C9QmIFaoMubR+/GVpMDxA5WpQtA0dR3TGIY+fliJKuCA3bTmIr+11817N
h4wfHLMG8qYD6HDvtvSMmsb8cBARxipqVA4g+yMCYNPMJd2NvoVdvqbZ+/yKXaIdftIYsN7/Qgam
78wt7b/vogpA4nkRIhdb1eESbJKl/ghUHN3LT09LshvQNipQNrfquUIP3pLCckT35xDbIiEVybd8
fGJlgNy7x0HgdwlZmEnw7/o4GpjlexXILal4AoF7wPOw8EtJqhOr547McJ5/l3sDHSvR7fjdRwKz
M83SItmBCETdxL/Omha8cpciTXuEmzRT60xfSY+t7JzTF5cdVQwWY7s43D051VAM3PnYyvyYwGgv
FDvld13mMaJdz8lbHCLOElyxDdHEWHcZFDk3/sAS/lEbSu1Ce19HrhZOmKLYLq1qbR/Mtuy0aFiR
2OYSELHB4G2FT/Tzj+9Dp/P5YrRTN9euoxVf0M+aly3MjhyLrF1PpA3elFGIT4jhSPMxpMTzjYSQ
Gq+LTNUbHi7Cj5pNuwgKd0H6anAR+ID0e9anZk8o85ZtY28gDkPjF72s99MGBj9dBBuH5l8WoVVr
wAubfnMWQPEvonTMPiKsfFGEQg5+D9MMUx3ianjkJTJszSyPxBBRAJ2pHjQOSW4fSfmA1Uy1vsbd
sLH+dV050skBJ/yzT838kUHBlaQHjNeVgVYTpc5ugskO9p1VfAXjKFwdRGw8xPFmPQL9AQFFJLOa
Mmv8ZBzl5PldwKh5URGmcntzdQn97JBZuCcsBjJtPFjGVTJLQsh9cWdXBRoNnyYNyrEZ25v9PwFy
VmDw+l1ND24iysg7LkvMx1mpQUxXBHIQe1XsvNMLDNkU/FtK6MwlHcN5z9BMi5HmqyPURPmZNITB
wGQp5gQ+pOoFeb2nVVqyUXMa6UYsyM0gbAf9uCngMlv2VExcD6ObfvZ21FSvBL5gZVpfXo7DDHx2
0BR08J9KZmi+5CRRs0QuvPU76AUijSxEI1yZIpVwKpGtPnDusJkoEYrvObgZK+csKbrh3pHM+vBl
Yfy1TOyZ8qR1Vv9gwhhiRwKvxosnr7UD6DIytaTy7PEnNop4ia8qZFtwlBcWFk0g8MSLNve23Omo
Y+sh0an+A8rUFybVJtqH9tY9ejkG1DI3E6FuSgixW2NwFWXmuR7KxVbfaSVqFFKDwxIWIelPyPiD
e2cUYLUhJoBxSzR7XTZGPGX9LQhioOMnNpJ41aSt9dWlWScQlWZzg4zpXTm1zBH8harChaBuoXTt
CJCxLKmQiRdYgpKO+GkjXpT6OaJODc5YWbbOrdTdEloULzdjsjQbMG4l3EZP0b8EFIZpRT90sk5A
azhLoWjGwGQem2YVzBK8o7ZYIpgPWXUSkkbsrKqJ9MBPZQ5yv/qOsSBzfZIabfwxiRL3rhDeaEoT
H8UyZBGJtwVrDJTZfvGG5qDGPLbXKW+BZi7vO/Kwua2iehRxybJargVJNOQFh78PvuSP9zhSukK7
xkTfGn32jdrd85snHjstn34ntei7DQrH4TISglLTtOwvBp+Okks8K4HdIdERfVczFjmjnlalSTcL
5i+tcST7FrmsMbA0NblYcN6jb3jbLwkW9Xo8+tqlWaQPv5VBFO1Q72KB0bLCVpbo69MKZRs0OuuC
ciahyuvU/riXBIoqH7zXvgprZc34NkcVz+LjEE8uUqHm4jeQbAqM5/aJH5FTiAyjqjsKMmf+OpBg
H2pUGR8y1w3cMkXpdHYm7HDHjvoXAR0GhAAVWUkmG99XKFwPwIJ8mQas/EVcKtz0hOxOIU37IOYn
K70JrYRlDh4lqEhnxFCX/Yk5k582uD/phR3+6Ah2ql7WxOCRzubdY88BRV1sfbjecWvwAZ43esJj
PdBJyAYmx1ykjw4AZMWyz1jNW58hzUDQLDyRLSSD1w+ZCVEstoDSsih5cT3+EURLMHSeFrB32N2k
LqRFlf7Oe7l+9eNPdbrHnyufec0pjRsj8J68Ix4/EE8hk/ZsuvZ4OFt/wojP7JFjlJ6IncvWP9+e
7CcY4bNmeK+6BKZ8YDZtXgnY36+LClZgbXH4ONgz9smcswG9Ow52aWX0CZaGAojmUixLa/slskjB
5Z3Y/p8ARarP3sicj43yEUNIOb7FX9+VAR+zd7XUyhVC2C7qQavk5/gfHZPMRkCC7wch4xDrJ1vz
SsQ0TD8I1zRpim+oXFGAi8/we6/WvSXD4WM1qn4Y+HMC3absVa9G6zONzaCAyyRNWAvPfzlEyF3P
dKpseGNPM19DXjDGJJZKtHHO3iCDICWuNqJQx5SCvh2j8tTw/fKNki5DPSHWx/RSYDOQriF2qrzu
4HWfrmpyDB7WYY8ugklksGnw4mN1ItjiZmyZSimGmWS2NZ7ZaZ5brfNJ3h/QJf02SM9zx6nANGrX
/U/KXcS0MySkfKpbC7NTqV6kLQkM20TEHod1BFGg/HaJ9hyEGZ9PTPYwew1x9GuVvrNECyUW76H8
jDXhxH1l7xTEjfp7b+jyy3/wkfl1FrmfGO3659RdlTiM7t2xCYLN7X/3lOghzxaf7622pR9ZOheI
KJ7Dy4Pg6GBlzCrd2zNaCU9lgpnw6uXW4izDMvUL7vB7qgxfGi0GKQN4x7Th9CYo9jvrFhMHypD6
d2w7q9Jf3rQ+XfvTyGdhhRNjES4gd1Bk+rTqPddCY9Bpb6Y0/G9tL0Gbhj7eRvd8jV5pPdBjlW9D
d3mxZVrYBfbQa4glNywjF1YLV+YfmvCHhECeUtcDOKxL32ppj8PlbivyyfIiJy6Uo/Dm1XBfFVpj
YFiELn127lsW3Xy4bZF+aU1qci78eM+UN0rSuz+xmq4iefL5SO4f4miFDOAGGFArygSM+Beheo81
SmwAZFniqE6lhF22y6RHfC+7/5H26l9tNB7EI3pfIDKCuBDGs9Z6qjx6bGS9nYEyOYj2ql6lEMA8
dSbGQphofnzlecDwqIY1JJvPeNtHJqA3z67ucSSBBSnOQuiZx45QXs3D2l2YnsXSm41pR4BBVJtj
47HVMhYOA+01uEeA8XDo7LAiRdAWLLpQU55IZrUSKQURKjNJzwhRL3+k/54TFUe69fd92+6fMiJQ
6vxyepBXtRYidWqG6edY8V4NcQhNFNIgEN27B6WImQivN8DfIsOnO1GPjFifg5R74tAvsmzQd1tP
0aYjrr/gITE4C0i5dqB69PStfulfPAt/zhRa0KD2IORX4BXLzjBofmquutJrem+p6JLyn3KREy1L
61TaIGaohcO4ZkP5NrlLocsJplH9ba+njQmW0LmNRT+JaGhIikoO766ZGjC8VwOs/1WAdwknTtZJ
PQvnsblt/WkWVoRcv2tfoJXFuEHTc6Y4cP5i7iKKzympEtc4lKEXqRz9gwsHpZ9eJjC5gXUazSYO
8qopkYV2E5sYgoYpXQPg9bxuLC97l/s8sWJU438B4AmxlDqej9Mbw2uTXWS5Ax1Knfr94PEMz+Qu
XtrTJIvx1wMwvNJI7HPT7r3RD11d90Fx8LwvejxEF2vIwC/Qd0lvd2Ft2TqQbwRwIDik7BN64qB2
Wu/VllvlHGdspZ98kdc+va6RHqhnoprlzWJ63DnZg3uC+nwqDlEYDqLUaTFRQV4eagQ/ySFQ35zS
F+fj92Fslb7UHVOHgs3DOuPhZOvngqEo2xDPj1iZHX/c2smhCSyRoO6Id2xr7e2dRP1a+R/KP2mX
zqGpn+ViRbr0ardxoO1ILaXneUee1uEvXijzDV7MEtsxp9Q9vD97F5HItteVoDlFWuRy1A/Gxkw1
PFgW+ZL124bx16K7T6HJvP4VzWJE6RcyOkVlNuS9lQ8lsdf7oSxQLwjcyW6xQNSopMc6Ts1aVb+J
ile+xhb3hrU4gs/4+/dAC5uPSL8tUtZAN3Naf+Z1HllK3aBnZyfVzrf3C9tTV/MPrT4EYr36wsYQ
zV+x7HKbcmnHN7NhFk0fjERGOEnITNXqpO1qXtsf1K4G85iDrm14LSNMoXb8MmtEml7moM8UjilW
7sDZq5K96VbzmFfvXm1E8dPgUMcCyZcYEARBV5hj6N04PMfGMGPzm8ORzqCTIc1B4T79nRsrC71A
VY0vcUIAUMkBGzC02vHccusl/uM3ANVbWKiBSIUWXkyR3zMMCS4od5D1GJmq3Aq28XtigJpw/G8I
xdnGt659Agdh/uZv+N1brObXGrcVDz6Ti0ehyYNVNdP4h+pf9Fy9dACPUM5tYn5WIdN5knXFKH5r
Z5X7JCoL0jKp+2H2QK+/GW2Uvsr6InnM7QphJmzshYo/ZpsLBLkUGr45bdSp9QKrflbqpCRSfJbg
I0ez5tkjb6doYzzuwh9JRdRD+SrECIx8P0+WetqgldnhsKZ0l10G7yBYGQYYB1Gy0IwRI3QpaKLp
meibER7nU/1MHYRMoYq4IBmbUe1D1pRcj6V5ebDsa0lJMlx5Qi4/10vdxx9BnHeHwdZGVNKbiOpO
dR97pls1YcqtkkzK84TUTg75hj7OwVxp0Vw2dQqj0iLChCE5woNmTflEzTmha79jhdxrnl0RGmKI
z37Kb714bEd4A3o9EoVQef32G84/GDbshF8NGdGtFHSE9d2umdrrJAan7YerEvN/+J3SgKLqXyyz
tKA0B2dq2fjUyztnf57noNHG0+Lc5gcylWaLMnx4Ni7Hiy/bKa4tgMQfQH0XZuBuBJbUaGkfkvLz
RhVgaNCidf74RwhNiJKLNwxKZf13faQEBBy2MTAJs/XswgeKuRszKbG9dOqrJn13obn2TVRvS1LF
BvU50Ta4DUDdsUD4BHyQXwrI+0bJ9vrb3DqfU4ByzNpfqJRYWmsrNabtfpPVfMv7TMYXuJ9Ye1z7
zK+eENNhHUmgZ6fkWUROyH0swiTkD+4UfX2EOeb8O4TVtiRdaKE9nwPax7SG7Hwx9DnAVoJ/OIML
nm0ecH8iq39+p39brRXvRnR0wK/rj36SOvZEG5gKuvoZTYA1xPmUv5aBxxWZcZW3hjqBboPbxX30
JOwpoB1EewoeFJOtsHHg6ZQOdd1p9PnsiNE+0bDw9Sze+kYAOpXLNMBlKWs3cq2pF9grhSkjWIac
6yLGsmhbUQmbKvXK6eZ4qwr71eVny4AOJzi1l6G6dYkpbwxa5P26E97x38pM417GBTSvex3MCjs3
xi1DmzpH3PK3tYqd96Duvo+Wrg0nEh5BsuyLA3ATOeRxkZtPlwVxaCjXUswSvu7SBycjLv+TJYP+
jU9JI3C4EieatagNsUQQ1+4GJb9Vj1lwOMTs+v+EWolrJ7BXMpplbhIWAu5na3yPagmX6Xn9Fp/b
mi5d70cO6GX1yd5fhOAegdCem0uW5gLd6pxr1js059OiZPsBOoIv+xbZCISbyNx0gsnzdT2wIF/z
2r9KKeoPWK14bF5pF0HXdYrKHZ4wwxpZUcIYPf+Td5LQKbnBgDnZvsbi6YJyrS0KaVJEyqkPW3wO
tS7E2O+5afi/xuQJDprCRe7grRc4QmRiJmFKsn9sWz7wj2eAWwt8CXk98GTSIWaloQ4OMmZosZaP
2tKkgalaXfbcbhiZ01GGjWGWAiWmjkKbf8a9IaMUBV6spTBy1Nr9qa7XU/N71DbcBCYZe9LzKIrJ
ALYRn+2OrchqS3uLticIQDjlW8NwSSzZ97YFOI+hZkMJcgRB0dFtwxw7i+tAZ3kmp1EMDDlE9x2Q
FtHWlKkcqglW+pJOb/CTGdJQ97LXqfWyW0Kjyah9Z+Hv2M0GwNkHr0Jj+Bk3X64POd5ksNSSXd4n
mMofkPP3oxLC+d8HX4bFPktsPYjp8zs7a7VWnX1KWKtmJMdOnzEG3GY3raACf4JYZhrLDEXJcfgM
rErUawWY0m7B+QVlSJTclEYzZU0BZoGpdiSKStzX89aS0rVaQKSmJtQWphUt3rEtv87WxxrHvfgB
iZuIY8VLuHzI6yLJlUZ2cHLqU8Q5TYyTpqwE+MxSWYMP8Sq8W/lChuXFC+OsxmTc7zBcc24cFkSD
zP+43gWFQGkkvP+ybpOwXxujExCg7HfXes31LL7AabP11cJcwrOmS65dto5Ix5m4sDYBQXZOySXD
HcmkmoikqB1Q0NDZB0Xql/hfXqZkUmKRbblLjSpNJPgBy5O920R0fkSQzzhF7X/tFTmsMQtIA6I2
2lpbEKjlX4QHh7A6Wq0YxvihUD6FW2amnxmua5WjtCAnrLwQM4vKB/SkFDAhPqD2HEAuTOc+6mIN
a5cE5PdLCWYg1G1IyTo1VdfxSNIjD40GbzTjFrKheewNqNJywahEXaVmi32CQrxc0eum7MP3kEmA
FuUfv5HpAz++q1t5M5ydnRGfr0mB/iJ1FHm2yVij3TVegYf+5KQbYejIxdDiRvpD2tz0KPMzQANS
LO4uq2cFDbyv9JtOqiROejxQwyHlsyiAtVdth5+d/gEe6QqeDuoLinJlY6bnKepHmzh9Zir128vD
4baizmyI8UMSrkhC9zjrFujh6GvGmOwf9de3vA2Dvf84q6RpsK+hPx5JuYVT2tzmqAxyYhVuo2Cz
RiDJCjF0GnZxY0DGoyspFe46LgJE2u+Bz0gD8Jax5Bk3wp346lFjsQelY/spbdY9siNLuAov3Zxz
xOpIP1vwUiyYTFbXv68TwFEspVweBJ1vGwrK3sTmniGHb1RC37rlqtK10OjFUJCNo+pIBI2i+Vmb
nDOnhCXAp+Z+ba4mQmgo+WX1xmzam7RgT7FJRn6nmmoJd287UhYKyEQIMpqdqMxaeHQEAPL5VP4z
P9qp5TZ+1h62IuTbk2OjDKyBnruk4WJeSERo8XAgIGpO5kVyXlA1lETH8hnuicQx8GM+rVxNdlHB
96l9zYNuoDbS7Q5RAf9xJjt437XwzSjOubBhF9wSMPlTxlB7SqQ0a7hRtIxHwZ7dsK2ccwY6YN8I
AIoQp5tKZTMbFljFZXo1lI5dq/mu/pzwCHcRRR9kPyBiOh3laYCWJ6TCntpnqvijUU/nmER4exAk
ZGRe1gHCQAKBKTh5mV/K7o/Hlw3MOb+0wTnV1+UI95Bd+xcrYmSY+ixps7D2Utzldqmq5uM/ZYyX
YsUaio+qxWu0V9rE9h77+TozxtzHk5NSgkv+kNQopY9u/OvvK0K4iZz14xoaPfvXr1mInUZcUgF9
wYFzcRGYnXYkS0KUXemGHwWJ14a94hvEccZWCSmXACMBvrmCGI9XTOT3aSXciDuUCGiNJ1xnHx55
tpBcHpJgXc7W2ULZaV1ve2YYZv0xlY+5MxLJK/wv3tpMx+4o6+dn++cojDPtc9FoEDgrYd87IZE1
ZoxVwRnPmZz48xE8qvT1pFBvoXnuNyR+fGeoUT/zmL7FDujn+KcgDcbzYO0wVD5qAYal/1AUMTRD
ROiHvN6Y9xNiiHjTUgTA5mvrGIKR2nt5RdI26MEu0waAoMbpj9TQ8GVMpWnV14T2G0ID0SWgLm+A
bGJfXDtU+pyc4ju9bQ4/Iahd7NjkM44CM2svRJ7QnSFF5m6clNXEz7YRIDmDdaiwNQ6ns24v49Jz
8rDwficGI6WMWA1XUnCzCBjdKhMQB5/FndF9mtz/DK8Izv32aVG5G0vfiakR6YJnGnEpmyqPvwFd
O6WNFFKeeM2ZUsjtf4rpT//smN2gh6jJAU22Tng/N6yLx2GNIHWZtyVSqOx6wxHw2QrQX0SeEi5j
V8lmNQ2znQzp3S/gTn2MGpVNnud+qO4VVk+YrhfQsnUtYtiNMKfa5v+bz6YZwWaLc1flX3x7ksMm
HUkpzvxzxVBmag8PGy7tLz16YqsafQjSjB+hSHiqLPnmtbn5X9VU3YmcdtVN9ipo1nyUDE17V/6K
gJZ0fSW12ezyT+oEI7JglIwO/ODryXU51i8EhWlbM3BDtUFHwTzpvDtN5O38lDZvY27mujn5zhry
B0dZGPpLXHuFGjpwSwCU/Rv5Jv2Cf/QwTbiazxBwoJtGCGX9+warFg1LNiWi7huL2xuy0EzYVhxd
LBFj6ggy+0K0HCXHKwDbhXSZm4YaBlPvPX66rXsaOhFhhce6uzb6/vNX5A8Ubok6HkTkW2uvx486
dUaeWnexSWJ8TdW4oqCgM/a4tAVtzzB/bokxey/NMa14HmuUxwUnNcOxhrAXnnvClCslWqsYh7zN
youYxiCDkAQz+z/BpYOf/WXS46o057PGUozwuLWFc9k9+QHMNQHqzm5MLZAx+HFllemeoCqQP+XZ
jEYcAZ+8ADTTnBnOftoJTpbGWvUBW/0JgCDClS49Vjlk3yn3juQeIhpMyacT2SL/p5SVbl0k8/kc
vgKRBX1H+N83MD/NzWPgJo8nNQVS2cz00CEC50DjsG+UPk3HWJUpIHEKFwaM+iR0UU8GIVFnLkx4
XhHf3Wntiv5PPre060yVBIlND9CexL59jlaH0plBOpdFYT7BsKEvPc+mMNogi3onYLFDu0qUdHEx
9zUVeXKKG/dYQNg22QnKBhc+tPLvM0Ljz+Z4YldXETf/QkjNygxeinTy5KmA1KqcdGRGPXuk1YIx
MgFE0nWQdRTRQpkaOXiAMcATMGouYW+0jtYc+clyg6GPGwkuNgB3TrBFkGTrNmBAXxRIRcfksm/U
vD1RZAodvTg9dRpTMXHJs0YIiscbd6YBmY33ffwSYcmaUu23t17ip8PcOJwydjyS9sqPJMgTz1p+
7ohYjdoUCJjCZy5hJ9WXTeLwqczTUB20sbK/aQL2KAPgi6CZIttgLR8vuQ4DNnEy6JYmGtRcAV/q
cMLUdjEaFL1yifs5pQe+WKd3qUR7A3UgX8HMpk5p/HIn0Rc+gUTfXm+2BBAJp/vUeKCfJmBppkO7
ObGH3MnntxmRQ61GE9JidhZv53nR8b3XzvLtoY0AmlLI0a6s2tCAuqW3eOG7CJYo04dd2YQ8z8tR
ft0tJDc+1gYsbrB2ujLmlE6pdVP7DLXSWPkIjMacVlWntEDNv4A2d1ZHWvQG+CKoh/GhbAhFGFa7
vzj6j3xgdaKbfEG9qH1kbl+4SoBqaiGEXjkfR6XIU6SByHcQ08JeIP1gLnIVXKO+4Ldi32Ai5qiA
+SNJlxfDB8vNM+DB5t/2kyInFMn8GJgUshNcfKoc4/8OQrR+LmJOr1ya46LPnF17wTHHb2qISGyC
v5iaUYgDqUaAo13Hx5wozMEcYDVl1BuJTYiRLtT5uV5h+AAM5far7DfLDxhCKvczfs1sTjH1wXy7
WPf0IvYPr8Fi+1zfWMw6dRTlFOmvjhtMnd9FhdWECKGTcgFCWBgWZQCHzpmLtfL2lNPhHKQRu+ii
RhkyHdwQ2ONucWOV3h4QxmhbI3QCie6L06x5Zlf485QhlRzqTNuBfExjdXLyWqVtX3FJIvju+Sq7
tG/9W1yjmQmBKYdfbnkX3cZB8Vd38FEKvNGvSWvHz4IpavVp9usSeS/UxEttTTavfdf0YYGHVNAA
zSQK6RK2+ZZQRkJqunLuh9oFZV8bNY7tvXWnF4AMO4Ximn7kFQk9XbCKxp0zyJ4h4yMnRw29Pyka
mJ4YvPpkwnTJYFxvlHBCIzVnD7dUq6nTVEwodSkMXhJIs2XqFJQ/wItiBe7TCQDT3hWNmkn7IsKV
+rxM2FZZbMc/zrVKI18xBnguhtVl8YYs9PvNy21SF2vE59yzBWg8nRM96F/0XcJVen7btWTVcrYq
lXFtaj5nsuZcpWPBEgrXdAZPG2syb1HcS/s8PvS2ChDpaoDwOs94LfGjO5PBwomlCDW9ttHen2fB
McoXJQ+RyvaTmvLA5rm3rVYJK27AahQq7NxDUDe33Z5A/EQDKPf6HtfZgk2viMJdJSOw9gWTMKW1
jM6zUycqvt0EzpzbT6czYwQ9EcUj4rzroy+zCGuO3SJLXcL51QvDLAzR+XfW1g4GAHd5d71GQo+o
/g8ljaxtVe1PnuPAkBKp9pKfdbf2BUUuK8Gih/N6x25rQXBxYGIp8L1aeREZ1mNga+4StPBRilbL
U8EwYK2TXogzzrnPs0VCC/Efm75sSQ6N7OiYMz1UB+WvjI+wsWvzNjfkYre0JcAnok+/b7HL/a28
DPBHhSxJC7TH/gYSEItbf1RxXUlLGQnoFsLzPsDFIm6sxn7TDOm4wop5ZcC1S0vlXU09V8cH084H
Z31AZ5qZkwhleMSWdTqFDPQbBSc/2xg2IOx+OVtF/TkaZvUdIpdhz0+kSpB9SHeRttnLKYN0it1y
79Td02QIlqjw2jIPKDsFiwnCcH+U5PlOJBxh0t/CQBQWQ/b6OaXVJOcI2etafjZG65baq/5kv44P
s4wUHtimO/++Mb7tQvWTGKmObY+Ja1MnbES9Vax3o4bvEtanM8oeVdx8sT6Opmm0qFtys5phA9+H
IEppJOdp62D9vW4I1EyjKMjlscKbONVSOZxcGLOtM/7Hb9gW8flKFp7911ghq3Jf5nTx8VrBp+28
2XmuLdBX0QzMmxSl4pjLxVxNtbZgAw6tSqzoNExdqtPXDAlKElM/WkVy2DdQHGyh4//+wSYNXr47
eP5LGDFL2AePcvrbqpjJuBzNZU7wPrGP0Se/fpYCs9OVdj6cQZBfLOODZg0kDh0hoteYG25XDtgV
Kb/+Kb567L3fE/0VJHmCMnuQMeDHJVDxjJ33XuZBbsL/eRGFhoxueEtYqTKNU9go41pIOwbi+YOw
It8VA3ks8m18YCHb1zXeUq6cStnnBOY8KVh1moORQSAQeS8PnvcW56Y2h4YzSBQM1XW3V0mPYsAZ
3br/jNtsvZ8fxBr3lrvADbCNm+tuZ67oZWA5DKrixY4/yj2XklO0tKGn3SEapItyeeKoSYD6Tv1Z
UfUEtHJbVDBiWo2loe5Y4iTPZ1+FOGxhRd40lfBjwRMhHiKpB8776BcOXxLSUCjfHN7jSeFRoScb
wP7QIYyRc2NsMd0EBZN10YCu0sphgFfNjZNN4KFSxEUnTpbSTVye8dchpyc1ulLdDIZ2ySG0EYk9
xwf7UHyQl0XZEp+af6lfWK5qdeJxWMJt0hPb8dzvOunuePoACaZKcTne7k5GyNeJUueY2uC+dhaC
DV+4bsRiY7LmnnmhWfem+pZfAOEc0JNabK/f5WXDBpB/0VbS2JtCYVfCrLPPwfPN6MPMtBVzYgRG
+Yl9FCrqDeGODoE2y2pFcjobuAubEQlrnLVbsh+6Z6ehmPXmfvcxGpCiCLBOpzIouRVjxh1pJVU9
0fNLy0KLuy2M9GI4cYAXg6AWixjx99+UbDBYKPY+tiJgDHb8s0wKle0AIzgL8IU9iOONBpp3nYst
ITy/zugldf76tUcH/MYhjhZ2+DG+gaSzEVG7iCzAKdf2NQDM9fBJ8KfmEKG/Iih88FweOXdCgbR5
erybvU0I/vJWaG7fZ9ZO4zB5wxoL22CaFSELpTs6PKHckXLheGq08X81b1YL6IIyP4FpCE3XyAg8
GniiA8taeZNEFoxrebd8cS6d3+v5g55vTX0ljYwKFqe0SGFFipfTrwfQYnL5WKb4Ker128ss62Xg
HQIPbPGVJr8XAzn3oupMLmG7L65WYLmhdAulq6McupghW2r0OBuD2wxFIsDNBvwSw6IEEOSZBCaB
98cVmIJmlCxR9GSMQ9mwT7+Xiwzf8JQzNFlBhAp/WyvtevOOLfJbvxcow3UXJsMriTdyLIXiEWBK
rN8PAiBY+QLv9Yln0J6CYAINYARMijL9EBrzVqFULv09JuDbSAoNFwPGclIong1kN+Sx4rEedMKe
7ZP+zgnxGOL6VQU04NAB/WxMYLYPzs9LCmJjm2ksyjnAch2tRtE31b0iUILv5Nv8dKL+EidIYPRc
qIPI88ARWUPo1K9YYlt8f7CdLJYVNQNH+v+lX2rhf3n+I8oppnxWw7FyQYEAW0QtdidcsYjwX9Iz
ESGTBSOnlpRhKaZGIKGp+M3V/XDq+/Qps7qbULJDYHhr7mwXHT8kS11JoCHuMU3zIpbPokdV5GTA
Q3wAkkVbZcCs3n5gf/G9iBlRlZwP2EJrgGNEzghlE+92hHdCvZvVmZzZyAaYVfj2roFqrhoJSIhZ
hFfG9ifquf/PQ4v4yirD0W7AWz74EAPLw6odMMYNk3+9h5ElX6+77BOWBgpb8Z+0VWLUob9NCnAF
ZTv+sA6XPzw6y6e+d3pns3SmrMG6KDAKu3JDAiBoM00KE/KBWqTQQFIEIOxzR9LV/cHpihc3/dtz
Fl/du1aDp6SkNthFXyr6p4JHdeoRqWGsVK0bzV+IhAFKxkCxdn2lP4gRaqV0JEXL5Y7A2jq+UP3c
c/ywEGIQyYJGslyWY4kygb64KbBRSDo8A62dC0BS9Fi3OJHmN8q6M5tK8SBtMHMZn2ZFq/VsdFVs
tRbni4sOPRJA/rR0JacbCegFm/fLoB6taKmcklXTSdc1NfCwjg8DnbYe58zTMa3Mqpx0s2WgSaAr
+fdj6r/9b4VJbZItGuNU6dCi7vXeKwuPJ8vYhVyY+c9sA3+oyGyc1paM8WlFrDyHYsjA0ek8vsS8
lAW6iz3Qj+3ULWd393JVka98DHZGrB6+2kJUnZz6ULKzCUgqyXWm5jU0emnao68FVvfoP9UbV20b
Z2R0EIN77NiVg6Ij30go23s061iA/QaJm/UYctE6+uRi7y6m9PqQJp57aGDyrk0AP1fls8JxgnNm
OMw96DLX3jsYJnAQiXahCKx2RVdlU65NCCn+HKi5e/YjhB5ec2OUoPg+0sC596ra/tVL4xGgu1dY
DYkFzo7rudyRMg0d6St3HjxtVpAj+7pCyRvSqHOygaTpD8QFY8y5xEO2AwJ21EPtNPxRcAMGoIk8
EWdBraQX4xEPsA4i8WFxtCC5Q3zFewN4pMobg/dyiupmwlYNjLKjdANz19zeZnLezuhddrzg/Xo8
gKoNgci/EBnbGR207pUk/vBJMUIHYeHszFnBMxJ9Pdp1e9yFibTCdXhl3GKOelKRb2xVgB3WLfBI
ixjeAEVWO9aHb6w/lk2mpwtiVh3GY/Eqg4lDECpNJCGqWRDSD956avqcHaM7sPDZsvCX7WukNZuZ
k/ubOYHJq0JuCq+6bE1pphKNwQ76xJ+OJbNcYmw1vwVhZqQmY9WXm8/cFqqv+2OKo6SuGdMXlEGB
Bxwq6hAzytq7xZ1B6nigWc2/CXLdAw6ebTJizYfbfZj2aOkhblbXKlCYk3DCegqh80SJE9eZ+9vR
Ea8f+hgY2n1x6JdU16HS119ebJnTnvBIZl3QhMg27qkKbAXSZiYk6CYHaRW13siLz85sAzK5J0V5
eJikMzdmSIM2E/G9i9h3Qqeno4Y3aVAcpVT8cRHiY4XQ9cLa7+8l+wHIzAROBkgv9oRa8MdpFLIA
xkkAmVf4sExVb0cPkwuWTa+FQdyL9M2fOiAZ2XJYZ80/81ULc00/iHAeGojgWoLUrA7wYx3ktMjn
/AcwZXlQe4Eu1rDzO0Mb/Ntd0exLedhhNHt2PGChxQeQibfT+Ywr424yhCqDHAdqwomIy7umSpFU
/XTxEdvI8bww8AdSiO56ia2dWcZ4H8FAn6fT/F6rcWvybjs9gOyegSKDJUhutv5uGNGqrIUd4RFd
GZXmS/qh8HevSVHLV0HkRcH+QMXTc1xyotJ7CoecIeMVDkVHOEVTUV0SmxrlkeztgfiLxMiyfgqS
WBJnQM/kEuh7X7Cw9IDmEeWm/G+QNvVwy6aacMQAhSI76AZdp3SwS5JMEAejVmPQpFMUOZkfpkTx
kiFVnjfeRaNbxtIYpICbkwrfEZ+F6eIfy+YH4+hlCM3oatGOrHUnKxw2DRbLgQB5VepCLTxhW7Qs
7qj4AzLKGO8JMsLL3v/pZyEuMEHhSKBl3EZFe8pw/Bbv74nakJPgANjKHxAvRB53xDY7+gnZYEXl
jDKxJbAq1qbp4R71PJuRiG0nWAk2oQQIdRzRJTLoEQzz+9VCX71n7eKU30dCY5bK56gfBOV8QSz5
S16iMxddSTu83t9zwqUGOD9fGnSQSBDAOOMCuSvxB+p2zaEhauQnvju+TNJvh3VqRtyMzlZpmEaM
4YMkbeHi09j+jZg8UZUS9MaaQqokq7hqJXv/EuBla5F94VOWPmxrHuaEmvyUi5+I53J/hEbSGiIs
Qp2iLVHwf3OLzSQ/L5uJ9wPLHvTN/xRVFNaSdPUogDNeYVMkG34o5/eKfLG4mggXQphZJBio3ADC
ps8rK4O5LPHnC/QXe2TmKgKOXBnYncI94oSgRabpFIgZow248croa8RzlaaqOnaADDlz19Izl3lS
ZM6xtus7SFCkZ2mlQieFsi7UeLuxKX73PvTzbAG3Qv1DJgAVSNsN1y21aPGXfy6DZwn8xsqAc0AC
mryRCql8Wqe3n7PGjDpU5RB3NKbN+CzV735LmmYL3Ft0nd6p9MFEUXOgdAK1hL5SXclemD5Usa7C
36ms/NR1zjk8+Q3puq77k5Bso8C4toJHxBUvKowdtkX1YCEt0Uc3vlHm2iSaQE3ebrCX/RhIB9A5
0+V034YFFGJkd7guLsEaOXbPjPxThJIl3p5SYun4h29h9ZZjC65fgdaa7zrNk126UifldaxUIpTy
eA2ClphhVjz+kb6mHW05pDMEU8U7khkuB+jp/bhx57XVo46WMMC6TiPWclHjcXDvMFsGkgwpP/4a
NoIomzAYRM6sUT6ewb8Zc8GZXoYkFcVgKEh54ZPiXkLxQ3v8X9ZV7JIiaw2jGWSbhuAfb7qlxRAT
BnNmW4DfNaNKhu69lIrTTgoSwIu1QWQEfcjz+rLbqr6JN3Bat+BVctoxeP8KcZPNiHEkoa6i4gyy
oS+HOIHI+DItqii2dhlzv6UmsrIJO1VL5YAqvgvCNieVk20s9MGl8ZJeHXdomkgmv3+UQcUhL+PP
BXLmpVxwe+BKW4Y+5IKyXwAxPW9pxxNUtcliasi+Jgh9ae5ya4FTJMIqiAG6Azo3VCpsvHyLkzdC
WjYEY8ZK/YxaGqnZG4zmh+fF1jlmk3uEJStuj7j2Wa91BMxODrUkwRsj89q3FDn/wdgdPFSTmiUf
gCjAKlAG6RYOyKPSDXWkmYIOuISZVlTjrM7EV/DQMnfY4JyPbAc1dn41fUXTct8bOzj8PdFwfIb/
MyjDS/uNFw+yLqt7HG60cOvT8InIgRuF+Vh48pE5FrKHSY+boR9p5VnV+9qsib/Uasuj39DW9ghg
Z96QEQaKG1MdmrlXQpYY1Qqmjl7dcEYngyBoa7VPxLDVKXICvh1RevWjC3gqfKwQuv8Q9suNftNu
5WEKb4PMUmoSdvTLYdG/8ZfDV9f6NrXR5kUA/fHAhsWvuT4X/8ERVOze7DQw8/nKtHDfr2RYhILB
oOF2kCYVWmjmP8HeVjRZs+WGbMNejITCMt0CzRhCLsONUot+blpl8WnhHgV+9cunCww6Bn+mvysS
o5Y6ndcCpTm264aen4Dz0GCMiDGI0dI75z+syrOTdZ3d1SLPfKO8opRDALH3qy3wIzAUgnsyq5pi
qO4PAP/u5DDwXWmB+ZbuaE1YAD1lPl3XF8RMviLnADYRcAMenACgMz09WJrEOmVyul6PYZdrx4lq
oJh5ohqNAda8UUOwen/IxW6TcYvS7tOTVrRMRsaW/dkE/QaIAEUlpJYCE+KV9m/JE3HSwr83tYOI
5uLFwMTAgr/2IEJ/zPupM6gnkCctdVD7w6FhiPIEu0suIWhTQPo3ZkI8p0A0PpQQ8kqwOsvVLKTh
xhoanm6TJx78zWV0b56WPLJWfKSP98SLlxFvYENwVuhWaP6tLg4i3lEHX/hfk4Wnj4f5KQ4PJsYF
kMxINpepoFgwF2LQiuKfR5P+uI3KaOrTGRfwkDjpumxt91Vu6YZOt3TchQBl/pIHnye8HluvEE4M
kEpaQ5TEbu+gr9YDagA/XeVJn1PJCOoT5CeAHIPCMZCcT4uieA/gX/ARuvcLECI22V6pj3J5STHT
EFamTQ0NdH2CKJh6CAEJ3vRsHMVWJuKKGiTp0rKn/Eaf3qFCSkj6wl8sqKUAg0DclraDPWiMpTRK
sx1QcIO6tFaq51gTDhN4hAMJC/FdXGpom44HY1hCEqsW6/I1rWSiN+lxQg9vGlzlhjk8MzQvjk4z
UtKHYhDQPNRMmKqwk3/Bfncktnudg9pMEamIDwOXNKK8VAUaeGlk6gUDiF3k80WuKsaYmmZ8ozXR
gHwM2bKh89OCGHcvC28QZX8J7TmPtirKCr/VuSd420ry/uzUDEnZRUc3nmZmI/nteZF0c8Enys6a
v36lLChJjnofBz/EHC//gYy4IpjwXTdI3qD/tisSm6jYpa91F8W1xfXaN0yannkXmlWOzqZQKJD0
+TYrAsnB4sfGTDRPdV8HjqBPPFzwpDifUNb1ruRh//l2VsV5Xo0zTX8IGgHByDZ/MVwO082+LRRc
TgOa4Dj3+lNo6b4KKteYb6MUhovtF6sCx1MFoRIgRtRaFPabTQ6+6pDVa4fn3jLKTCsOnaziRBP7
/Vh2UZdwnHMwMy2jsjvPcdpf1FKCDBcw8dh3mJkXN/OAR3Qr2+pZfOINH09m8kuYlPKS1oCudGD1
41qwIf5TPdE4ylD9JSOqzk0Yan0Dx4JsXRe/Z4JddxptkZQg2Rfab6FJ1bS5wjf7gb61wcnUKDfj
4p7U/yAjFHq+UJsWn4KwSMqrC3RYJm4EGax4YOHd4SiLgRJqN0rEwpbJ1RCvjE3vNB/oTOnJpVyh
u8c0BcUshgD7u/zd556U33TVGHxoK/LcgXsBPY138lns1pbKkVvKzNbznQicgR1Wf7sGFxG5M4mS
V6fp+6g9VCNH4hKXoUSz+80q6r4pVrw+A0NyqCPk6TtoSjmSppPX9Ct7K/vvudMgQQ9KDq1HQkwk
P4/fbR3VQDOAedDi3sxsjIn6d00Y8ZXH9cU1eLxfQ47wLd+4FSG41rY3ojNb5uerHGcaQ8QnKSEa
5Eb3NRVEf5b7kKKL1F837oTNsFCSLlEhCDsrERTQBi+HAoaPbDW5ELHIQESRB9prZx3jDM7fsbd+
eXz/PDl9E6v5CKOd7ErYLvYgi3yxap1jKDARJJl73bfAuLcH2s4j2SyR0nnncGSGGcNiEhbwpPn+
Jx5hEAqWMMw3TRUTM+L2fmX90ujHJUdQFIkKntrlxeTWKCgAVnG1/G4qKQM0JZ9I5RsR0+GL/Pmi
Sa4xK0J7rJ9CuGE1ymgfIUtz7cwvxIKK541pApnLvwR3sNGBcOjPS0txBAK16twfdg62TBXfQ95D
LeeauFJkGa8R06GoM6xCjstYEWbjOhAi8CO5bdEzq0PCjPElCM+uhsk6RiKy5QZTGSrbmdm60YpW
D4D54A8wHOAr7LJ1clfUqd5kPH3BXJv85/3XzjZRQr3nOcctSMMeE+seVDGjvdOdkLJFpbJeow6v
lq2v+RbMDAyqBn5wH1koAcAuIqyt39jscViNUvRbPfOKNzyEwxkn+FsGwqIsYXLL3nMdPmp6ET59
SybOmx3506MPWOAR1Vkicr9g+AQ+odanaMfvOd1sNUjIiU8ToteqeeI0MS5QT5VHRSXpHC5UZszz
XLvkTkMM3rYrohigkqkyrIiFJdR9/1M9kJP2RaE1NAqDkJ5Jy8pRkhv1XyAfiVBQPOMSmutxwpmo
sk+SI+dsHrobtzfp/d6sf05zJyhKPUqervppt3Kmey3zLCny0c7hF3KsRO0oAUGR8DGy2KvdGWN7
jgJDuds5aakkyVlodaFrw/DfMoPEez1NuhRwOv4XFEBqIoP1P1y8JLd7T5ve4RMfNRSdYtORv3KY
gLBuYVMXcwNp5SYqaM6CO2C5SE5y7kSatnhRHq2BD2XZ0oaYEJXXyjGnkJPg5xMEJ20tq/ESS/KO
EiI5WkOVhTUpGgim3UakohcYj8iy4xdr3YjbJ8341oCrjQZS7PMlNg0n+fXZWr9qEYl/ZoLq4tij
IM4EkBUYQ64xFzxE+7X5Fr/pUuIRqpdANU7X6rpSHYEMLjm2HmH0qoJt0cCO/TgN/pMY0/mwCgyK
k+DHjtQrPH7e+17uQA4mzo2HsmVCqYM6+XF30RrG6Zmcm9l6PKRl5sogjB/oE5gLOTynsvbWsh8k
kH4a6kA+lEx0k6DJlsnT9fMO0V9MonIywMEq46YhqoIFn7LJ2G4TPvF5v7ry9aEyQ+pAuQTpsw97
T2mDCm9iFacmBiaXHQarssLJhZwLt0aSEId8u9qZtEU1oKDtss/7f7G2hL+zZ0i8i6Lq/fhYqANp
a+IdkmZQss6Ab3WMFzkYXeEgYhZkuc2865DMhMmKHSzjnMayS4ABugOPRivGKfNeRkNQhvk8pW+Z
b63QJ1ASioEK2bxQ1YbQey4N31Ul5OgMFHjWccj+qSLCTq5pzHYZJhvjf9ScITnQ3NdAA0WuKLi9
tbD0kYqyvNgtCqJzvt8J+pJn6egfy6U7qVPbYKUxLU66rbT/4+Di74l4UViEw6lXAiG8i9Sf9cWI
/fl3Hn1OPvsxG2YPnSJmVByKEt5N2bxH72gdF/05oH/Wemss/x0HxyKhtvxNhygXsE16FZcng6lC
QMdSXBy23IDlBhyOzSrL53OBMQLrPpIyXH0C6q2L2EQny5bZVjGaMD1a/83bXc6XKNQAoL0nf9UI
zLY/8Dj0PfH+JIPFJpyg/lKouWk+8l9ekUJ5gGzm7lfErGEA7RAx5vPhZEzoFteYcQls/WpMi18V
isTK9PEVebsiXwZphk/f4zuVuDHi2ivdmDzIjOtFom+xo92ZV16tqdTSsQcCrsbMzfYA5Nb+sek9
/rKTJkONu+GDI94GKsHsF3cqhCJAdHtWybxQ2hbMou4itPn767n/NxS7u/xrQE4HMAuRlX82FXUK
Czdd9XtphbSMCV8QiNA8ZYPvnced/kANPWpVbEVFB3JoKSsDMDySBscpPtIFvDuhKemtieKFCD6s
SFlT4kT6LksxuCmauidAzK2kggZ262Stj1wWW2ALJo/lmHFSzZs7chXrOEMP4Z1C3Qb8kS4Yazvk
KiVdiicQWRXZ6mU2u3sCKi+7zroVS/gK0jLy4Euncsj8q2OFbHnn56KZ0eM21o8EXOK/7M+COZ2n
oNIE2eFqru2ks5OaO2xPxm2Ipv2RuzJHyka4TZHcXq/Jxsi+sMgEeQQ4QFsX3iRlHrE8S2jw/LBw
nu2r1F4MBBMoljy6wUCuEbZZ2xxP/cgFO3Om5R+TQzUsPWowyPJzmK4Qcp3xalJfIqZKTa4iL2OA
Gby3+Zv8yA/6raKnqRgGdfvbHbShLz0fuLzDVIfJZwTcJzjD7eiTgHx9Jdwwxuj+Hpwy2qypg7lB
g+JYxB7d6NZlu2Av9ur0twXlNFsoKmnukLYytDPJh5lHNexyqEBKrhRluu6JSN0A7GCJ6MKytCz6
T8nhzL2ODKqklJTjAbiVdPOwTmi5dryyLHdvCumAR3zXmarytH7IcPlHjc79UBnTuDouAhnVr9i1
H0wzCYWHNZMRl6JEeALAtoMUn1J3F+9ciTr98EMVYOZMz0Z9ro4xYsZrstbnUZx9FuaPoHcTYLpX
kbBsiDjrtSuOP+ohekehLXzzxLQNJ2UD81UOf0QjUxOC8bxQAMfOwnqc3A/4zu12FGtGSs2PXRd0
/F2EbbMs8cqYPHP8PW0MYBqPW7jkWPK5wTjuOnSXDbcIHUxTzyZ4l/0yHDga1SUeW6b714FGHOQ7
0zQ8w0ZlwiD7ZVo457ABI/6dOFuZe+JJIfxTQvgVlOkJFmbZ5cVzNeBczIJ+r+0MBiNVVzjpdcPD
/hJY29MZECM5hP8f07YHUYnatE33508HhbNEGtJ1nIGYdEzVks8EwbsuH+zcg86bIobNvsI2KRp6
TuhRpcE6yUU1QV++TDUxSO5xusT0U0mYDxCYdz9YhivssQEXX5a7ymwG0v07hNJAUEnZIWqJccBe
ft4WxD34ngqoQrcoojolxXB5Je+G01QP7kCvYDr7aHTrMdJWzkYA1ywlWBW0u1RpVL/AowZ2ubdR
kbRXHbpjB4Z7LZk9EamT5HOGDWtXRorFzFgRA+X76PRK2N1ectAgFxC1FOzC1zZntw0n7vEv6lZI
+lDxcQVU08B90iRE3qT9pvBHWcu+k+7Gpn+AKAo8L51Q523K/JHyz0N2cFyZPO98ZkHKA5iAHRbR
6yaVkCC5Q6drfrkssSDGvxQT0Z3qzrhgbZ1x49aTIS5uO5ppmxcWlTxIaUhXksLncrbiy5MQsft5
Xembv2CIZY8Qgz15w9fduS+qo2FZFU9a8zVOpRcdSM8Quzr3l+WD4xoaoyjEe3cGkbtDxp+8Iwik
6VWQuy56KLEjepk/Vu62fYOFzuriSOc4GhCENt2S9Ut7qwTmhiKf15G2MxLUwlixsHFJ7ig4hmzh
LioF3P7cpD3Xo4Xa4N17I0hWI2A9/8CFYAxy2j7odLUsn+lodfYtr8p8qDue6TKMjMxqi2xQ8F3Q
q4DfVVG2oYOvwHO9isCZ4V5JVdhVJwkxtAlprgpjsDLVUC+a+IXHfvtfjjgkXjnZf/x3BZNrHkWn
9WxaJ1GneBvVoKQXvv3Gc8goysKGLs7m1mqdw0U7rQqgIVnQimPpsYM+n1Fmat33rSU36RoAUTjV
4mp08V0GWCz33CqGeF2WskKG0/DSsuRhZ0LIGXmasWVRpMwwe6zCSp1JHgydGSQfts85Ypau3Znu
9T4TD9Nsz3+WCRnxiUmr6Avf5uUBp+43uNjcN2z4uehzr0wACEVqnDRGQxJLj6xnH5yKnoCoGULx
qeRtpE3a7gi8RGtPEPdQ+dMCYlduo4T1F+DX2haeXOGTNn2n3h+F96r7B7cOFU07Dj3jGqNamtJY
Cek+qcyFzMFj93qBcRl6KetIOT0/BIwOy+9VhZMzaiT7tWGuYi74c7TYKF19MEScT+D9qSQnXzID
6TU4sLCOiaURZUhptB1/49WPF1ZVlYjzkuaidZ7WNMIkMUCXBDES5PK35KUJ5/ylkSZGynvaDuro
TvJmpF5uN7Y1veld6gMADw/v3i0ael0emniNTGwjPKvWi5VX4KWCDc5zCH2E2uNTwod2r4V3I0lE
qwxjqpr4VEVREgPJax/g0dJwA3VdFOwwAVxNN6KebW8iT3Qs0O8sOPKVtGKdhL+doOViYeV0CXOz
fPAuEUGbQeI/Oh6EhkhyvSTagZrAeRVAotU7tX5aV93SsNj5BbRGjg9yHW3noS8VX0NDMbA9XiH+
AbbHKDSMlXAQWmWV23EJDfKB85C6hp0Y2Kr03gpoHVSkopHp+qb8FY975iclAQKNEZW/P1rybZNP
Mp1KRmrkS8C0EsUrQqAlAiCAZMp2thDsnv4/Ec3QHoYTB6zxaNQ/mAgtGEXQ/MerdsFRzRHootmB
3vBDjMgl+uyWapAXLgIX/5VHHmRJYmKzrc30iFXJRegn/bEub2MXsrzwmTrO/hwFAdH1Kzo5iYyE
iP/l3girVv8bwlPpdVuu6woi7CPd3C1ovzoC6I5uNA4nL1aGBilnyB5m4eLA2AmIeznsWxomEbeJ
Ot/DiIBOhQ7WUdVqdPbTElJHn5heZLp9C+XFaIPCWcwWDCAX99alIINsPKCgFZDADm0NItc/cYXJ
YBWKi4IYMy6W4gt8+iKrV3pyntjyfCJfVAKYAvc+UJKeeLMPpQwCVyKmhNDPnhEUpDPMqwYLBmN6
Y853Jvrd9QmRC7ja+DRQ/PWGMHzRRbdfnVvbluZDpdcpma2175qOhqVzMAPwZWuBne+PU5iDIcHB
RUQEu+s2AvjbsEZibok7L2Fq91Ir10hQJt27ValO3Wrfyw6Iz52Wd5a57D29ZQaAXwdWn2Y+iz2L
a/fIybpBgqSHBWF4oGgOSQeZqYUq2YsoOdhVTpmKcB4O9l7IwYHWkfHfo9DlBiwbR0aL2W1viHRy
ADsIwOkOpukjaNS/NwXrWghiZydUhTYeDcdEeiBAGA+6q6jkI0trfcM3xAP1cHV1o0uxV/x+ermC
vdqEl8MI0iBPumc8Q8Y3Z2+MlR7D6GSI15mWWt0fk1+WycfRePHNPdPHuPn1m9k+xmgO64IgllzB
26qHqr1gQEOpSfswMwBX5nW/ANP5WRk5iR5VksE0k80aCrZwSsf7kQC9ubAeiZBwhSEtr4e+h8vg
9fMw2jXFNgRzb4ACGyBgI9yCXtcnCihw/cI0mmub9x121WzWO8t+ntclG9oKEW4IYvimAVbJJS0A
veJRyGVbixDOXOH3ARCBkb053x8orry+wScT4M8QmmKW9Dl9orfLWXGeh6Cy2446LoryhbpgaADk
QRO46ISkXdlup9Dqa/41wsO6bl8KKfldfnxFe++sv4IJScvj7cceR1mJIqY0riJSnrKBDBdooUAh
W/+bwmSD664WiLX07H+jyhHloR3kR/4qk+mGU0pNFCQkeBe2x1s/Dj83aSxyAwa1hdvnfdy8pTlK
oMEHH+GorWXZtgvusO6FmBgj9R1ciJ4+fv6jYF64iwLA0ELzMohY5B+iw/6fo3hTdJdN29UFP7qN
SxKmA1wD5vSWWq8V5KVXUy6OgTyxbXtNIuggFH5PbO5N5mvQC/BjPvjmD2I0c3amWXwJn0bPLmiF
cAareBDYWkdpTS+aqjWMzeQEcicZikTB5eZ/EKdwJYc92gb1GOv7c36RO82GubBPj9jo21KgbbGU
xqZiLnegxW4LXqA5lnU6DZvyTulWAFo8yuAKedrRcpFcHMijXDNuxe0/WX6yg734KRkgPy3pwz2y
irVZDjOQiN/URZzjEyJBa0Fq4hnIVLy2jrGhDxgeCwhFsudoIpYQ8gsTzN81MM/1Scfb3OIAlTJx
XctnRuHd006n/1Yf50hc8br4wwc//um00lWFR7HJXcgGjnbserspb/DGS1deKJ4ZMb9axCpi3CzL
+IKOSw2Hq8Hnf4RL687bMqu3pe5LqDM2qPTBK7mhKTQAmvlPg49zdMBWZO6EtWK6nMQWxvAslNjy
u167oWBbkLPfldwBxzBnf53SIXQC663ul4QfyFuIxYbrFGzbh+upcXD/0srOzKXFEy6VXwyaA/7e
znmOh4AKqIp54C6QvDSTihrYNic7PQbPIRCkVeUHqux1B1jZExqPI4DmVsTgeP/MYcro6YuMrj2f
DQX1b6sbbvKqo6yWIr1IJ20WSDh697UmKnF3oA3mCU7C/D3L0D1WNlqXwS9sPYim2rGY4WCPTQL8
GV99nEbLGnNC2aU+tNSBA73FE5pwkijxqHtsk3MCIMaiRSGE727AN5tAwrwif7B6JVDLA8hPKdv7
kbvuwcGnfnvSGX5a198RwfATifnUpu4pCz/hgh0C5+IHFm2hj1mxdcz02H2jdCznEDqJ75m5g0b6
stylEJEUn6IeWl640bpN7PcHx7TE7j+9MnLJV8VmqgwiliJGuu4byzVGcJP4YVqJuMLJy5t4YqOY
mADNt3dIe52nYEyFKWTBFjb6iCgkxOidEgY45f1CngFGsYuc45naNrJjSUrFsbs4lsWOnjAbsk0N
I/SEysC/P/TXvDIfHnixheVHisij6uaYa7AOE0MAhc7f8qxP037UUAQF7ztqYfabkBoRluYnpk/1
4TxxI6CpnNgDC5Y8a3FhSq1f1A2uOBb0EQf+ekWfzjwdM2JVf+o2sQUA5BAeyHNTBiJvrI6w2hTb
ja9dOJm5dP3kGgckP/GYb73SUVNHn56AiwYLH6Y9hl8ns66AjppbfrdtJYuNRSxRuGNajwGMpOGx
PIxykT5X4DWQ+rDJQVh/5HqhhJTg32Lox7b2DB7F1V/I+jJxDcRxtENaHRAziz2SfJtWt75xU8vx
pgSQycatw2fF/gf/QXGeb7bQcSlyBpZdXQldaxJRIXzRszBSfvrXRfTfjMDhofEPKbn8AWDuCdH0
N3/KAcZPsiA9O3ibykUrEvyd4X+Z4vuNkQtafEAO0v216ugbVEm2elj0TqeoWUZ2SRP/ZdnhnMdJ
XmJgTskXJ6LIlWtu6vG2mtH99q9ywuGmEa8cntLZchXDBGLK+RdHPExf7W+LxeFJeNgHMzxc5k7P
CtKUeeUpop754pV9W4/pAwYAFPk2Ps6J+8EIm0sskw4ieLa6vfeB1AVGGMRe0AiJ4aw1pyNq+U0P
rqtfdxNFSE3MQGz23gtJ3TgO4HVcpKscT7k8VddTZflYuHM4dirHfuhIoaimW/N3tAgsazULTKqQ
5VCYaOAY2YvpmVz9hvM7rOEy+KVFKdnum0gtoECQzMuVxBNGLnLiVJ3fhmqWOqxK5aaf0Qtt4AQ/
aP1qoNhREKyo0RjMUeR4ADTymLDv8MJVWHxdsQuA8h3M3syB8Qs1lg0Uqdd1NEVPI67MOS0lqudr
ImatAYlbDM910nWEBDhYeh+H2SCy+tG3UISiiqWNPQ63rRb5MKMnzGhOUcog0fTdPJhUVxOGfGy3
P5mqOONfRxu2T5iivaWnyjDAqVh6tySY4xe4nU1yk6bpzytO1XeS76155IrJFwFM+NnxosLSMnVW
bmuT/uZUKuVsJ7LY3VdUAaoyAILiTA2OgbE5khYkz/vCtxL32EbbjFu3ltpbpLTxC2Mo2lGNKgDg
aiiF61urz3RcgRhhCKTvPqcrvPnN2xdc/d3tANd0FW2Aw2L09rrXvbSuGLOiKe41X0Inp/+18oJB
Yp8YKTjBF+2c0ZTzU6qZnJYF0pwGxdq/cAv1KyBUTXv1U/EsqFhLWCpyyIXM3n0jiWDfA09xeiVP
WJbTfef8tcfOtt77KRYdhO1SllKm1QHWM5a9tCXGBDFF+B1+ubA14TU4Sw3/uB9vjVrf3djLlXdN
mePDN1KWv/B5Yp0v4PqQy/omTmB6Imu3TrTdcLGpU6S112Rb7OevmreobrDIzSPvPXMfiZ6o78ft
KzZxniQyiCBmOWXC+OwNQJSokm3ODbFmW8nsne1u0eZXRKm5IkwYqndFD+/soEk+QRAyuWNxaAbo
bX7tRZJVZ52Rz1VR+wu7+/bGEwoK58AfkegzdV/ozzxB8pGaBZRd7dnlv3sw6EzkmteLYUpFQLwm
sSYEtI+BXDEsRGIJEE1cTa7rSSlFJrnexf7pfFEEa0B8zf7PXkdziNkToDmnnC5NVvyawSr9mg70
cm6ucjgu+DCN0izPNMyR/xV72vYaHTKOhAmK1LqAtOOLjZ1Jg28yUOjdIhcKYPKxKt5DpP9p3mi6
NDEgiKYh600M8smj08N/688jhFqsRfzqactNIuTFtUBXXpuYkmO3+xuauFPEoPB9fpp1z7ImunA/
DpWECGDJ8EW0mu9kfmXbWt/ZSYjhmFRIlum1Zxp3Y7EcxSw2sctApoTMJh4EN2X2+IvLJqoxkgiq
E8Wi4kC+eEJ2dfY1wuQKRvVvAWAMzmFjaw5HZrDzag9jxfN1XCPmHreiSPweTNOhohVzYwc6Jt62
vKW9D75ljBMMFpZL70Zz4SDZUdO/h372Hn7HY2GHoG5t88ZeY4Au1yLEzf31g3SIPjNaztc/FrFY
cftakBpUgz13qpVvtk/NM4iCksnqODEMgT5UY/G4vNAMPB0IClxJ+fScAtCiysz7IUhu09zoLV3n
LTOnbyWRql7fRsihAABFfbbVZBlKfbr8rKhGoSMIjzfodbOUkK/xtrikWnmAqimMMjxgjR4cN8xt
pBh+koLQaQuKDMHj+LkpcCeF+oaz3I/yNnnUq40FPnzxJB9p7yoAT42Gnnk8a2v6yy+dGz79ELXv
+gM2cxLgjlxDkohsnSAY7RMQeCjePQ1chyxmfKEzuOnEr9O5qwgw4+jxzBrkjWJmoW1LEOeRrfMU
ZDTuzgT9YslW9I9T/qvDlMmypG3o1pN5EuAge8/fJGLbEhRTWo5Sb8EkU2wThBWt4ojjA42qCDIp
8kDBArZdbeYOpXxaphwKl0vC0idE6qDDAcp7cGExgzvOsXifPrWu3Juhr/Zg459UEHh8EDorSjd+
PSY7MVUrE6CD5brORbwJGMH0hfPEyni1IkUeKxxgDUnR8IGJhvlVwymQrRmDq42gs01xA1TX4TzU
t3tDJi3Zfis6Osu9a7qkbhJA72Oc52FZQoen2zOtfdwHgr60pDapRmp3eZ/NWbV5dABDh7HgZhyH
Jn0CPCQnzhfDwFBeiMzmB26WUfWD4ygj6j72PHZMKVCBTrHpQnCwDdNsYB60MhzaHlCqwhyzsNvL
tb/BmmeDElez59LmTJ4vetljDOM3/VNYHVHgfGahILqhIDE1F+APNB21OB5L/R0xkZHh4SLzymLt
z9K3ZIRClij8VTXPH+//y4O3CeOKpx29xYVjl6WIDG5aGPxBY4jYAypCwXYT10Pih0W3YpW5EGel
4uhxZQSs63vFsqu90MZNHxfQ5z/IeGwGX0IDQgh7QPUbwXv50MIvcUkniuLRRw8T/rsatqoGROdx
b0+tRAKHj6tNBjCik1PipxTA0xp7r+D5Iuu0Wuf22qjODJNZiily6/I5SlEzM1AnY8M2Mqy5lAhw
BuhhOSnyUntW5owo41/rKthWoDLQvd84bV9XRdP0p4nE3r32nS2HSZjpi46NQDmjHtBWNAFcTaz8
uD9LQGC7R/EpX+aNqA2xsy/i2RU9HEK8VnBill8hDdTVbUytH/iyD8ofHmTVUdl1c7JakGgXL4dk
HZz+uk/A2PXStoo0COfprGSkBhQc3Hn3Qd9KZXlMUp/XnBZTSudZ1QPSq8jlK4N73j+hB7lc57g1
pnaVetVZ/3HHQ6KqD6f68Jt6K2ptmvuN4QEd9nRMhXErHL9RyMEX+XihgzmeSABNu/G4uTs35zoo
y5iDOTp+Wdt/YFNA5F490QYdM8njbkS+EyFbC/rshK+tKUQ0tY7G54hEAFebpRWvKx1XRyGOrq+K
GL6Xb+Bti9BhlL7zCXYNE/sW7pgLrk+M7Z94p+TYSc5tE/ARHov09g9v+XFOyNO4C/HdBsTJjNVo
nnoGOwVa+DBv0a8Z+Q6VoPshmrq1MXujAIIvY/JqoWzC47OVBNHYQhFldCLII5yO6JiXca3CzEyx
I7jYfZPQ7G9mKyv4sfolNXC4S6lpUux1vkMy3bupBfD8HEICvqfD78wFSol0uDnyfeFDkRN2xfJb
hfF0Jr0mC0GsyUppTO5FkMcosPnx3zkNFRhts6gkuJDSSGCKtM5PV9Z3Z9GFCgHqzQDt5Ldtgce0
DgJnTz1nwlLx1GGSgOES9rDRO55tVDVGd4hpLaLVM0vc7e5EgtGkKP1A8Wf598vsrKkyktrDrr81
OWhhXSNirCbZ57eHPttlRTf/QUTv9l8Pm2IbenbWmKJbtv5NkJNouCuyZZvqdoJWiUFv2fjIeHG5
Gsei1TDpFHvUrKXla2Dr/gc/59GLLWs7RrTCN+dEefgOgub+c6D2fYLXpEKM0v7fu5WgLdGM4m1c
6ejjIsk30saan6sDto2GH25x8S5+3uhjC7AQPnFzUFEgV9R7jYnueP6xTkkscx64gv0DTv3aodne
93hmSfVYR1w9Xvtw7xSN6QNxYrn2Il8Rp4Yx4/00gRhjkMmHdZ+YkSyPQUlztfpflOIz98K9G7hW
JTYqSADcNd1FVgU2QuWGkU/Q1ehn2TCKyT3xw23Pvp73pUGz0hinPZ5ICKe7C1t15PaHbyUPK0rz
kaNLskkel+tGSj7VbAukqAYgYzCcXILpY4yPl3HB7PIsMkvypjB3HYkJ+1QsTgHPhdaQfLDBaR6W
qLtEC5re+/Uu5PhaVBt/JlSGz8g1fVaS81XFm3Q5kvLjGiwJVH8NBbZTtjADO8HidGaNyhx5u3JL
k8ePsR7ICuxVPqp9Ogp0Uhu6807FLxTauS3jkaPoIOhgrVBSMGIQ7rbmqYDlZTVj9rhEwIdVG5hE
NFH+J+VY176mC3mtD1NwJW8oHDf6qvKUAUwnNlb8xkVkS6M2GcJ5sHTCY41JsgFI87HJK2CZzaDo
xxBGNB8kZ16S1cHqveDdrOgX4jjfrP9TDn+czZOLv0+G6JkbKfudeCGgZTkeHvrVaS93WVjr4Ae5
NapOr06xUcbAKMPWyQEMGpZJSXGLb946ezxU6YJK+17Fn1QSFtXR9PZSE1jOOAVFerQ57FkgCcQc
cI0o1+pfUT0FmpcxXWJv+n4eu3Xvd9s3IF/96IjpnqkhqhsK4XbseJ+bsyMClEbsIYoF2qjvxAC7
JqlWVnTFK8SERducoFyXOk2EueO1tmB9L/L4bHYBU7vkpwSkwQxRLAVgbNY7+nhnTd2DablesC83
Kjx8Dw8XB+Z4R75LR5R8TNxoPya/qMHTI285R+2ljASZFY2N/bOiY2+ZO7FsJp4nhcot+cHicoTX
aBxuTEyV1ZlW3XEIiGGD2qG4xwJ77CytF474e2brBhg+PBDpJyOSU9Td7ibAljI2o11lJfUx5zlH
QfpPzbbR+jC9LlF0ihkTz37+O/KtPQnFGpOUwjdPA3/yC/z+NYtSyY5YP8d+1J3Ss8nrJfT9vOKi
PfxZ5bRlu/ulojG1qyAAuOvlleNyiHsG6EeuxGZpc5/XMawW5EyjeUTw32OssYunaTEUm9HFWpvS
ah/u8nERQN2tScpHxioDB6MuULZF8+n0XafxL1o9LEi142xNWdsZmbmE5JRu0PTi8noy5w5sA7T/
KYa8Rj3yXzP9v9qKihbxBXgdH5gQMvJnBD2UL/9gD5ziRhi8bgA8NurqXDydmF5LaF8QR+uDmhXg
6QvULL1qSsPOJ6VwmkvKJhryyB/IAw1ZXuf/wFtquLM9DHhTER9wOe6JSlx3Bq6D0qoG2m7i9jJ2
f0LRK6IYU9fccLbgQZV0NxvIc+7GMdZKa+3IGOO1wcotepAT8QilJtEeBLPmFIJcE/9wd6U1nidS
ZNceHaI/gntw+tuORVvMhUdwEKY8SgWVo1bf6aYJUfxgg0cxIREcw7jiHawvaO/3/GXaWzyPMfco
vonM8spRtWD2HiUaUPbp71qSAFrzoijPUZGFkx5/OHxW5q2Svt7ACaIDUhc/hqJE/w1UbH1MX+kM
FeTiirIPlnEULOOlUV5nKl9ykFArX6zaM9YQYO/ZIgUwNhteeTJjEhYeP9dCF3WDPtntLknmHYEW
XqUct53wRwJMOZdiUanEyHkwu8YOART1K8cCuvDL+lOCMZ6XRwIKmQ85zSiTGW9hGUMlET6+7Mc1
d9yZO5/ZSp6qDQemrccP2GHXHpTtEpLBe8VcUk3wuzntO75JOiuuwfA+gZLiLLIJY/eJX1VoMV3i
EoVUwMIjk2hOFKLWcYVpJa5lOgRowHHWIHVPAUSOMrI0jfotOHU+g72tkNP4oyml470zgQRGzhwE
vos7nsDtFkwdwapehi+QJ1xxFU38gvjq9wHxhgBDsk3n1PF1NW5Emwo6ZhKiECEwD7XRiPb9CIi7
O6eJqhvfg7pd7MlIBb6PHadYeubZN5/MzxSWqBlXR16cB1+1as4q0DRBTcu48yok4/j/B+yL2yBP
1FFdpbhnsHucHLJMxmXqVQQ1ARWgtw27bAnO3Iad49IyKE1NCu0vP0aRdfuubIjVLJN2Il9HnP94
ipTVs3Mv4jT/5Au8jP5YvXpDuoNg9HxZI1dOIYyZM6supjLAIeliBG1xv3YXOya0bwyMCB6xlDwl
fI4TOGConGBMiEW1dOZhwJA8zxEeUx4e1WkpU1h68eql9/aVxsLpVohEqZYGu/0VwFo9+UcC8fN6
BXw/uIWQRCX4GBgqvQ/zPMf7Otv0WYcNNFuso72+8oP+QcHaja0yBWkZX5a8mhvcae1YRxUN0183
jjBma+cqmXTHW4wKwPVEvICr6Y4mpYkP7KRgOeVKU9PiJ4hQbY1JVZn2fSppk2qTOajC6kDPm3xf
QzUwDpjHnUVnQIafbje2TckpOq/jUaVN+vcSMJlgOCGGp69S5h4fF1+vy+npv4Nw+f273C+bSMyU
BGg7EkPQem3s8lQx/CvwAx6GM+T1ozhsP7KUZi1H0/eTfrIS8Uia5SytNIyATNKxKFzw51TC3XDc
fBrRL9Cj3ja4BoPpEXMGl3JmXYUbo/nHIIy+R2ne6SQQr84W2Dz0Z2w9pNQdhMhR/yOwgzPthbvk
OgOeBxezf8CVJq1A9mjynWDr2hLm+sCZvBuQKpIKeQYLtI2fHHs6F4cLyBTdrdI9kom1ihwiAE5H
wzKDZNEMjQ6UWHAhSwUEwcCFfXEAtmIGwnzfwwlSV9w5qVnITR2tpNNA+oeMao1ItLqa0sgpa2RI
fFnxvPr5pv2Vro24QOKIZBWOvFBkjVTx2PJKNK7N39pEDUhnKfTdYDcGkJ0rPS1vxcHgnIPC/VeX
3O2nN5Z15wyy+usWVb75syKQ31M3O1BMLNsRFoWs34Y3XqDbMaBd7SRd5rZBwy4YI3G9Ab+CUJIk
XJD21atmpJw1F32XuCf1iLvaAekfAecJc0n1gUdqVIeqojNJEhmc1GA9t17y/wPpeZdOSg037rQw
CvkCGicP0jCyroYmLoD9CNMpfJxE+vL4mGzmDjUfkSgxwL6jljGMyUSboSEtMaY7ZsQ+JSBYgDST
0jdc1hTZT0QxvcMwc8AVFORowIdFXA99E58Bw80l0m7F1Nd1zbW6DdHxNuRM2mQDM7VM4DmVvalg
bvWEKiQMBKEmzZKb7/knH2xY1cZZxH7kLHj0qL4SlPigRwdXg11eDb3wPiYPudVFG89PW4QSAx0x
UCmXimkk2PuUw0mWkd3elCcNgG9opffZLRtXiYPZTS/4+7VOelwcTSyNPGfF777+6TZ5niAjc+MJ
eQSlM/wF9/3OGdssa1Tk9RRb1rrrsQl+zvY66L0mDGZubOoy4wHi0N/V2d4iiGHtIa9b/6CleBRR
Q9GEw+OLOrUeHABYY/e8q2m1cwFJxamS2GijyQz1c1qLsrwI5lSCKu3JvpZLk5lzNFcRLw2Yt21J
HE1fw3PkZP09n2dkxArJf/WB72BQRxEhoiTrMB2PkijGbyYmOrSrkofmBCHXBaYjEHniMFReiCHL
e3vT8OBeKzwtyZeTJksScXcCnAkYl7vcGGJ0n1L4ha/phlDH3RpiUmhtEh0o4RwnXYJVkf+VlzlQ
lG3SG9tm98CiLBt2C9Qwjje/xOzpa6OlqsQxiPU6EPTwFJ1DQZS/YyVqpDRLBuiEQ0RRqBIvqujb
WUWHHlbCsgegUks+aNeqZupKm5VO/PrpWPFIdaMOW58YZUYHVBr8pmvuSAOYjRWpZjLBo/4w05KW
OALOcTTtfzMD5yJRbPOsNR1xhJZAxUAvKBeu/PVoRK1X0WNWSJk/AaUZkZPQxBVEy96Mvr/UaBEk
SJn7SGtS9TXTKTwAtvy9ba1rFe7iqYOWkCbAlZUJsqeBBYR1s3IJxVNGMaJ2DAahpc1zYXgb/hOh
EDzmaoIozeerVsPx1XT4P11bcc8ECKxoV1V4TvSO2Lzes5Xz7MxUNm6qlSve0sjDZ79LH48CMx2n
IJ4IePmFfd5iQBbZ992nDIMneMDs6kLa7EgCEU0RrUuTmDmGb8a1xUYSQQbg0ipx+vP05SqzvAH2
/09QcT38WJVwfsNYSCUZqybld/cXpLq4jt2KFALpK74gANSFGdRRKojDYRZED5p8Pga6AgBKTRkw
1X7o12QwfbP24w69FOF0DyV+vEOKgPjaeU+AVEoPaWMZNPtougkyIgyuFBaIgWPIpAoqk8xjKzJ+
1GS+ygzKrxeDVcTtbbXSA6HGFtFl2jptc13uvhInpmx4CaCXFOkUtUd2QmEZuOaRzOtZLNK1RWzE
X1dySAdDWEmOk03MupE9wQ4LASdGn8p6eMBPGZC/JP3KtkLIpLr92FKBkvJ1F9wGyHYbaD4vim7b
tK4FbLivZecWkZZpdWkYj44qJDYns+wSInoIjJ8bOmsRvP+yFD8ZNXd6wEsYoOetnbK/8e4mXGN7
W6TgtnebZ5KNcbQklmMeZcWZfXF1iMIUaKbW59mNbCuQ1QFAwfyfS8is83G62QLtQ90JvtY6xnVR
zHoNHV0G44dDlPYu2XiiS9h1ZAVhibDZ1pEfk+l+ZRm9d68F2DPnksQX0ZVM8qrcjpK2zHhM5x7b
7DtWtFeRTpiM8QvOaDUV+qgsa5Ba007LMnWW3IoVoh6yGQ2DDjf6/aFNXdHtbf7oB4w8r4Ac8iYM
mDOLqPrAIB5fjJsrE/ZRH9ZQ5pYVmR92ApPW5IYcFDq8EEZ23TWvVGdTXLHl947d49iEK4r5IWv0
WrDJzKNH7I2NLqG/uF1CJJz/eN/m5j41NQIQjopBQXeRgmHigaV7r86o3ibSrIHgy6iQ00lQOUcw
JhsqhrrZsxhqDSQdTgP6nzfyWC/U1MFsnPzIC1s6q4InxBS/ppQWBJfkMSTerdr/DGLzc22O71QN
/FH/SeX9dI4Q0mLdxQzemQU6A78OvU2AQFafiTQ3YHGetCdj1z0qfkwS48/dipD/81r+mjYAKPVO
g+WfLy8vzNiiEdos/B1raYVhZ4r/zMco7f39eEkptiZQqRFVRQqr708qCZXdUXDix5TygVVl/drM
SDHWLrMz19qQU4+PmzGYp6rQNSbi20bIzlfvsNBa93L/o09HCN3jzaFM1c/+2eS96z37hV07pEHZ
AVSnID5lGlONCbW336mMVnuIQdcApqhsv50CUBabZ5vWP00FEGwX2iwE9j/HHuGNIgia7xj6r5Ap
+aOG4lh3mu4HFVb8RGaivtMfQVEabTgIuPCgvP5P0g7rC0LT1SXWwScLaZwsKJO8Y0jizAKmn382
HeZzSWSUx29U3U1ASrYPJvCVElAgM4XeT0UDUZUT4uT7Jgu/Bu+aLZwvNJF9hS+Wz9MyFDasFY4Y
lU81tR/Puz0NeG3ECFClFplI+U6Q2YEM1snPyrZSgSO/xQvtgtCW0niXsgSeSrHRBbhzXo/dm36b
Dbwu71C6gcUPkoJRiAKXT6Ks2jvjs0BHCR9o2wEhLvmEvgpNMx8tp3/51WXznST5Fkzt+gM2cKzu
GD57gexbkacLDerjCuR4VHxP4qoz6sUfviau3HlqjUo6ql0oqZb6c1sxDAu+QBjDy38EK0FibzrO
r2cNGyCVX4nWawsxKR8OGED1mh9EQ8XZhdY006xA+S49VJNxqA9vN/Nh3fxck4UvJEqVpyj0iXy0
2zTtzZXr9TQGBVnDmdKjNfaRnyYzQMdSvAWH3Tnouk65izVW93GetygcEN3MY6ERkycBVlrplwdo
P5LKPzPQjzKB6C50DTN+PLz38bZ2+lg0aFG56WFNRUv4k6IS/uEfITeAEoiJAUf7bEzo96Onl42J
z2YNj3q3kemg4mAZc4teZrWxtbfpD1j2Z47GWAvUGAodIovEjS6kqyzpcNrrINWCLYTPKcLhPe94
QxZ5tSGQXknsK4Q2IAoozYzm5eMxpGORJ2wg0+EKeomR/23rZTl1iesK5BgM627SASc8k26ePbSY
cHsR3YEpPUTY7L7yPxGTB1IvDM89dJJ/dH2swU/yxBBqvL1+tR6tgJSXw0IdtXR3UnT3uAD5NY/j
msZbeCbjjR6YdOqUHThKO7s2/lBRPqqqz/hhRswfQAIU2m3Ke8CuuQn+abVqSx5bMl4Vo99II94m
vc1a832LvQ4Caloj2o0jy8g8XdSjl0FOhlnKJ8DWd0e6Di4/ayVg+17SDNyRtgSPJzYhhanA1qBK
5I1m8DosJR9E6Ma2eBEI7MoA0sGbNjkgwmq1eAzILH9dH3/AcbclagoLEeuiwviuUIGRAaEttzs7
suzlXUkHh5EpSG6F12kL+6EVgSJPulgQDFhYFIBgN3E3w13XvCYXQxZkCiGguTecwytnDLDe3bdo
FJRNH3WhWUpo2mEyqa6o1TW2yREEYhz2a6tXrU8WW7cR7HJu6jxe2gqcibTopBlDEZdH3bExkCin
miDGsB9hP+JoPzqONxLjHI9zMOkzb+XTYU1quGHOR2UYTWJJmoDWVK2swxU/1ZXI0GaKOIQNLXt8
wfEVUYEFszMq4PdKva+VFT5jSsaSKZX8zfjFf9/9/Kz3dvF8yaZ4q4xK2EKpq8K2dy+zIxXXDJcu
+xPYxBKR/SxhMTHgTPFzeKklGdVTMCrRaWHJFQ5pqw6IMOzSVDHFBkYucL5ZkbAT/fccE9ZWxCu/
5J6yWj6nxm30kCluo7kSX7cdIFvY012rc0vOLyrWd0DHE7Rwc5y1Uhgj0ymnGVTmMhfKa2Zu7J54
cz9iIWtvW4iWPgWYTtQCPLzLmq2fxAWBjkUNhYJ9H+r+FTK90qp0qa68Lo85MYo8Sbw73Ol+xSFH
FdHJUhf2Gdego9dvRwWyTQpY22hnC5y7IlLRwrrGEoWazlXNZiFHJUpprESH1Uxhgcl4Q8uJVztr
rkB93SlzqodWQfi0wcBknB3rIlNGNEV6fGWykxqDSEQhwCj2aDLACrH/OXGOUmMkw1LGH/s0yjbo
jQfjSmcSwhtpUTAxzZSJXruQQB3PLCViPWoJwsk9XgVBOH+LuRymot6Wqq4GLJ5paKCqSTZfVZuY
ROzf0WkmhSxUpYbHxCi7iRcc7HBC0mBYd9bAfmt5YLpmB3nRCXphNGARH7LppXIUiiaslJodiiuR
GroBDgXP6C7jdSdEvSv3dA5PMoMc+uwacFP9XguJZAsGTuf5ZBT5tRCRRj3l++wawMZ06wS/npLw
3fyduP/zvMdv7XPb6T0wd2/02BgXqEeCCZcw5kGNKT/M+Bn18g2Q8A0jwXiBgOQn6dPk2huBXDso
4S69D6O50ukonNFxXnsMA/PuAsbSodvFMqAwhp0DC12o5nrg79QlnVs+Zjj2AQgZVnYQSfcNXb43
ZMONh71zHjggNlqbTc8J8vEvb8s+CTCwi3XtuKrqSIK1Pm8iSvWcRJl67BdCepXPYtPP33QT8IO/
yadNArQHS4vz0xWzPpr+ASQ8wuekXi/A1RFNxHl7hJ4y1KS0i1An6QOotbdMZecq/R8XX+uaqtmE
lf/BAi1h+CAtFaFxfsRL7S01JC7AIKkTWcAF3vw9obVFscr7hRmCIQ/Ve8N9EXW1flFBqNionBcJ
Ytkm535xzM1MHPwAwiOsRVkOn1Xw4a6mk15YHUZ6fnyrxinhzApEYlnWS3gjAr3Xb7AYDa1aL+jQ
JlL0ERj541JXctrdgF8JN/fpdd5HFVzfQ85eeRqXCulsy/ZuHZ/DflOLkt37Kd/DxR0vvkJtH167
UkKsGTVShNlx97jP3J3tlEVUUhPIoDUlS8s30VUW+JcaeAxT7GglAByf3a+rtzM0RtqzUKoAzwto
RH+h6zRNv1EqKoyDfpF9OdpqDrJHffa/0ttdfXNIrtbgIGxGVnyXiqNrFnK2+OXwm3kFnYn5eadg
fulGtvUSNDGUK7gT76EPsCWJXV37JcL0QTeL4zZ885/CypJLl83hxjnHQj5HJpbaMiW9eMJWHCKR
EkS5WywnmZtKrHrIGy/zEyGYVHnBQrI07JlA9Bu9qJrSbDlg/68NWjpMhgA2T4qEqzWQNWH4+tMe
DPavcfGEcy5r62aCzPBWSAUGBPDpwk+bOyrXaemAMMXEWpoJVxbiP9U8kDfo56NlMc9BRZxvrv1e
N+fDVuznAldOyOmWcZv8qZvE2Di+TQpNge6r7pZvBC0PN/IQ47MKkd6T7lnxqlCnkLIZ4a0J8vrk
sNpgWNGEzpbHizaMRJzerzCQViE3ZMJ469Mji4+kNUjXDaUsDo5T8vteUm+cfb9IHDatDo7brl6O
Uq5xS/ZTHR1+nMtI1uX1f/dZ3onMqceJubxV5z4DrkEWxr9cukCgo9gJHqctgMI8HOvCEpfxTw1+
e9dEwti21Uanth1tISWrkzc0V35vK3ILd+zMGkWjn14ATghFkLPsNtN1Frwhh2UlwDut0ogg1biu
6KYr70+SqeMtpcV4sZC6X2jkGOuZwghj/Yq3RDxjlE601SRaeor95iaAxG65zlPiEAytJLEDhs5T
X5SKdUR75iTu8r9FocI7tr7ZhgTbK9cI75/Ki1Q+1WGsGB2bestdqhz5uSYDwzq0DE4aCc99me9W
3cpisZo1eS3npSyqkCuiB86EnQ5SnksirSkfY8va4ps2wo/tDaVgh/2Rd6qtYSTv8plCE2jiftXz
6Op/3LzCgLwc1UVK6LjhG9gEET2t74nLEXbjHqeiTlaJGKQqqqpUSdUxzgPnHYvoSs3UwLzUFkdL
dWz8tVV5h9+cU4+3bo7zXgFZETeQAA7O1FGbohZepbi0Ez9YSzaVE0GWbgcXIF+TLcGxBWuNjnYG
htUMt8BfmY+yGa6gQM28j36wy1oWafpPxt1zTJk2coAKFKfOdwgNildYZM2winuIkW6MbVLJnmdY
RSAKqcDm59Bf0OJT6vRVjRdO+zZyjOhUg1WOg3W//zu1Y1WsehAXMehctN+kAiW3WbDyjpdrvXZl
w7PWLi3Zv6NZ7BB+a6c5gtcxApvoeq8Kn+PliVVw+n7LuzEsyvYeg9yAjeU8AHdVAX0cFyWoc0d7
OywNDyMF9JS7vkH8AOisnCqq84MxbIzBQDyLvI7scLTw8E0u5ov/TlP07y4QxX5ChGVPtjO8TGty
0khpT6JdD4lPVaq9l6Omw1/8Y/TXwBq4355HY1yCxDPxvJLGnVoeXO89UM7mUhO/fnYvRqA5Oly4
77ISHjkQfbaeRN5fMdekw3IRVe/wq42c82Zi4zfusHexQoNIps9/4/L81KNkT3eYuivLzxfkMpHZ
/9oSVl0fc9ZQcEO35EvTuuhFiJy+/2WoUWum/CHxak1n54y63t8H5HRlztPiFP+8xObIRe6oMOKX
HWPsf96ZVFmI2tJKj/+T7cCX4DRvQUItplkaMdFlOCuivNSi7pyCzqFEKu1JT5p4hPt32lG3dLm9
YQGaSFU7iYz6OBFG0cF6Of2bFpU+h3MjGddagLY4jq7HT5HBRCx0JwSOX+cp7jcm1MirCahMuUTv
GIoifemFk+jgJah9sSS7Hb/JDcNL2nvY9VsWV5IFX0UMLLVeDpkTHgqE6m6yENns4BGZOSJQDMZb
duOmZI+oB3QZSfIv8bbYvP931Zu4x9Xwo7xgvAqKImFhIP8O1PmfSYP9xDuJpsH6GVHb0ONPVhp4
o2TwyBXAX6Dr6s/vfoGWloZ4x9DLfegr9n53obfjr2f/36udvpYd2dfe5xLDXbD9QNBZwINcguAc
BcuAJ9EbQYKMa8fq6z/ThpfyDaIZcYMu2nDTsYdgghZK8kmELtnUvzF60YkLdUDpB8XjfPtESrv5
UJq3ANDCuYLDkEE81pe7rf7jp1tUkdCSC2yzoFgi9JKKV4E9A2Y6/Sl4tt+JICD692RaAsRhoRx4
EJUSQldmmm5/6GWwyfE4S1P6jLyK4hcAsYSHdOBD6dALVi47QX2H4i0dXvUB3CN9ksLdiXa0KjmJ
ueXHFU6Q5fi0163VKfwT7bmT246H6iYm/W98tbGk9vQpRATDEC5uLXq4yDrZUKeiGYGbRrKqZ/H9
rB/ZVVIeTzThaC82sxWoyEvLZc4o3Rs9BC6mN5TOyA27V7q2jy78VRV9nRdWO1b2N9EAuf19BxCt
cAk5Piv48ogmxOsLXT4Z1KH9Kapx2USkpNfsKBnqB3GviEElyJLz3D0No4MgY4sE1yrM4VZY2Hm4
5LSBqYUDag+EOo9vnsGNEmxXZ3EN42Rgm5WuUZIasqKwhf31R9BL4kvYinfMz5yvH3/+zMUlz1Cg
A1nOS0gcYgX7qmdzwXJ/OYo/tWiSAw/D1ymuiLuzCwbRESO0+5KxrhirVObB361DzkLJL8J9mtiN
gnTxp5OV5JTv0aE7FqiM+SizHrytVvcgxlKg/LIwqMuB+bEUYjliPEf6cD1L4WAQwr7nlz6zgAei
pN2aJ6+6r5AC2KZTzXjrV1/c23Q+6OUnnU2Uhtg5lwGLo6df15tjX0dfOOKyJ5ncfG4bE3+C9jv0
83+PFOGpCtt3dKWMrTYpmdEFJR8AevXkMFCk2YaikcyDyBjKCtfkkPLhU3LHvktCdW/79ve1VNob
lvdugRpEZGAQkheUr1KM0HVIl+Z0dljRIf/r/6l8b2B4OhhQCQfTRF1zmeNye5vQU/SUs3zmKwBi
cNmSdaPnBepdFoQWb1HkE20PDAPDwy1NZVnNIztiPwvenDEPAYcJNzbqxhtjmXaT30jqqBNGdrvm
mZwWbo1xICRqAtPt65NpqCJEUUoQxEaIXo6tdpd/Kqllj43JSqTPQ0EQBfXJMimOC2Vmk6Q1JAw5
ZcMUtu5FYDKIVUQ0b46PNIyS5p+Anc5xMxK2+lRNPLAq41h9ekl63tr2ksSN+O2+Ac8ULN9oKvhz
yfnb9mclX+zj6vk7du736/QZ37qmkVtCF/aYMnfDnohlsDk6uNJQG7BugSgqrHM/2h6uyTleqNeX
8RIU0FZGAbxRkULKaEKhHXubNBUcArxfHzkTX4eMy+Gv8qMXDeu+9CNdtmr4XVslHUZVMaBFdEFR
rRGUJUvaxO6/EwUJRTERn0OjkbkwDHuiWQvjmi8JhssbbunFoxT/e62uOuYd9hepxq4RjGbTHKdA
6EeHglxxMtTmJBa4sPwxg1YHTAHg8KRu1KqSRfIqxkUUk3uOwAi77ueMhnsp+vv98hDt6clIlEVd
wKfXpOCeJ05yXtq2FslrDk++5WIIYIOh2YyoBD96rPfbG9IJDyumrgmAzMrDRGiyMnaTxczzZY7Z
uUtoogX1hqQnLAvYsZL6zVpRTwIHIE1BBe7znSD9Jw3vLtMqv0ry7tKTXxxyXocIyNEooth2qNmE
cWP2KBAsT3+bBtK2H/ha+AVXi14c0voGAzN/i5pSWZS1R6sW5xZ/kCsDhB/yqm/aAV/YEwJLoLtY
SWhAJEt7BecYLR/zp62kkRtxbwjvvLcN8yX6kN4GDzugqVCsZMDx/q6C6BLYFjrJNqHe2+bEs+bx
5f1U6GYSiJdvJJLh4GVt3dkzCPW1mVdxeeo+9TgMYzewuj4xRNvwl78O81WcrJuHHg2dUlzhB8Nj
/2Fo3CJNem/iSDWYuWbZuPjrqensbIfhGuEbcfVxMPvXaan7qWvR3hpasn4ERXL7fKPOJom4C65g
+DAo+mzQnXU+2ux503zlE7MgXz96yY2wzjwQb7ar3Nb4GVRGI3Ntids8rkg6ruPoa5CVKUk6jpuW
tjqjF88emI20FKbi3JRYCS7S6sQnQNgDV5BKrV0WeBQlJgALy9h5W9xEEkydwOvCyfgqJY5PJKEn
h2NR0mzMa5CLoCJKcqMR7lkK1oPjpk8DMbPGGdg98XK0VbLwseb8qUzHpTmhx4JAKlLwGxMadkfa
bdZT/n68oEGv1BXDFGoeji3UQsZs+yuUnvdrhbXFp4GtYbvlTgMjQtNV2FyHPmaejWcDy2Mp64Ha
T3iq8Nu94HoFerPMiM+3B5ssS+OI97QcxzdMzOEtTum1guDYTxeUqDBz/fmM0FdgLAdWatHeJ5PW
mgCjw4gOZ/RBVdQt3tMDb6iVEz73UOHJPByBgsRhlj+T2z0ENYtKK68x1kIFLajeMz50KJSxbYp7
ngOjUO49Hiv9mS22TrhyXhtrH8VOOPpLvuhoYqkfqPi1fo2Mp+NUXpGBvjm26o3rOXtj1qesicOH
E4y5h0HUd9TEZZSj1FO02QNwdHKKWYN+PEpkkaybQkI7o8N6hO5DEWh+TIn4FAhudyW/JvkNBlaL
nEh/2nK97B3keNDr4XvKc92uKCjXv3IraLpOyTUMz8NdGbKnvMa2G8ITm8mXLfyet3ppCxy1Qz2r
hk0durh5/OTpl4xQnFVl0BTPq/hfhCy6skeJD4AQGEQK/IT9plBdzzaZ6q8s4t5mm66Xsi8q0Bcz
SyBKOIgvZN6hPpCnuNHuNzNIL6oH93q8plBqbsepDpMMxbyYPUJNf7PipuaTZrCk+nWGtaKfNnnL
y50/x2ecRfOVs9HHpJrG7QxIsXKUKOUJAokWppTqWqwlpRkyZm0aol+p0jFK6xGH8P22yk/g0Zpm
XeDWv4mBUNE0LCmogcLcSciT+b786/LB9YyliU6M+56EdYimozxI9hnVWTlsMPgX8a+1XYljMuth
GgI3NukqnJ4qa0PcaakEmEHLrEnD6F2fxsjhb5rO6L3QIK3RxUHFrcTUANr2G6Xa0IE+AxSftHGV
j36efGbItGklmClgp1fRSe63N2zhP/BuUM4jsSNzWklkZ5ByBMnfPviIpnwZd0SIis2APzXqmbtJ
NflL2qY7DS7rzzHhind0skbDAYod5GN6/rLwZ3UlLrSU0/rGTmmfD9eyNcjiP5ZibNCERDIgNVTR
d6e8R7ctfWNRHtcXcdoTatj3UgR9/7gxsxwgQ7jqBZ/n+I74bSXAWHs9rey1v3XhIcti4yXB3IIr
+xi2lbtIHUHkHL409cQywWge+cLNJichlJ+QA+2sS6DWAP+TeOl0fWOe7aQZ09q8AlzQDcgO5kVO
ESJ5bazV1VOkG646KKgxr4zCX3wMWUKVi9NR2pR5FQanPOEspe99GGqmPKj2L7IiuUopAPI/FvyV
fEhWJe0ywpI0ibodtB0nfEJq7ULzk5C3kwz2XPGIYZH1RRilMLu/PVhWiSv2a1qPtUO/D54cLs5H
IOsFA3iPHSrFTMqwK4XtIUvv93HR0C4wmnJGPUK6K0+hN8I9CIcytHPIZYjKsqFuumIOcBO8kIYU
DIxmIlg0vLtrFu+FCJNZzMXWVQDJxnFUlvxE7HVhmL4G+OfKLcT7eGI1XGP8SmLoGeWepJvQ6PXW
5J9r0Hr3JgXKyCXPjjOq1xDhmivUZc9SDjBBk63ofy/gkeH7cv91mML24fouFUyvzm4luwmwsel/
IeWAqjLVKXjwVm7nyy1m1bMmyH6x2WBHBPN55bLPhdT0nUMP1Ktm3F5rd60fwgkPtPgeopzrBwUF
mSWqk/RohIScG6NpswQSSoTezrCg4CWiXQYaq3CE7WirPoYGH8BHXhSyWT+ZtZNT0e4WtJOwjA/P
hUy538YHYK0Y4233l4EijrskPdM+MHULLlq0OSjY7QRwKa6B9WEXzNXwZeaZ5BSqZFk0to8XQor3
O218euMWqbrg8x3/QshFk+TbLl51HXgX0Kw6BLWMGF11v7/5WGZzgdhh3C7aROG/C9JPNP5Yayf2
rABqBdqaUJmPZ+5Eqq/f9krJ9HBKKFKre9mzNyAfmzJlzHm6vWNhrToYDEVaN4NEMQpb/DyCIvZH
xvlJ35caGtAYt8m7t9zbEWRO2zf3g+nvnd0wcmcJpNESw176aqKNCAarVIjpg/oszJCar1TqCVU5
9/D2VM70EGBdw5TtSPwgPa4wZYyn5U0mLHem5q0y366/kzBnnaMXCPaKmcrjg4vPvOWUZ8aJPy6N
a7jeLmyF7ubnToFfyUmd6uLNH/xJNzm+cGTxIROF4OxTTRBP0W4FTjNHKmxa+R/dIidMw/K8q3Wj
fkgIK8z4ruLivr0px26UpElkJJIzdb0YOY7/+DRQYamc4XcJLM1tU8Vqme52iodyvbnSBv56mqXY
THzTN4w7ARqSxtdkiQ49jNVNfDGYOZeCwZqjB2C20/fR5fX8oPNDKCpNQjngaKzgh6RzMK6mudKt
6VglT7bR7WBI84XI7Jv9EzqPIQxU2S9u8/EXJ+RMRraeLHmesgMGlpWKN9fJ/uMTpvzV1CRxDbDE
WLgRDG7itbqck700guALtDwCGsW8ihdQzwjpQpsOOTkKAUNXZy7jnjkME6iFfWllg2G5guZVrglz
86ryZQo6g36BC3l088sI/dXtn9pgD0BGslHhSj7CQbEl7V9DLMTD8lFrDPVJVMk+pPkvqR0Y9F9L
QJrxUJtIgdEm0+RCGfo24Kk8tRz75NBHwZLUo3iIDmGfXxXEWoFnR2Jg8MpOg+BWoGave3tobwnO
IYBxn9xyO2EF4vS9oocdOpmGSCvKY5VYysgXwSiD+FT6Y43Mg48QcX/z7mo3C+P3JyhAWsgLmUxo
ynUPgzNSFA1QPgFvnYkSUTRLjMuLHrdbrGLwkoZymtCTcvuUh89HM7tPuTJg9Ielnpc74825GxP6
VdBng0ubpd1yVJ20Dy0BC8Q/u9xCL21MW8VGOot+g21zO39uVDim3x15AlDUsOUTx98LpGN415yY
9mHDOJnnIIGGGUALFPqPtA+pg2UIHTkcpz9pMt4JZajJFClwTy9KcBWmDYm3bDemvDt1blyaWBpb
2P4VAami/fKrd82p3T43UK4BK65UcIepCwiHDJDsp3TCTODSQvXONJpp3WPnaEiYNj3nVS4WuBpa
hKmDr4a36Ucwwb6NUeBrXBSSFQ6RZvMUJKnkXlCKqJAji6R1kAG8da9j5yE+KBX+mHEJLrzWGpCG
NYZ48i67I/KNzM2ByOuarVWRQ2n5g57ejHAtzD7LrEocyT5EvWc5pg1nUUwVLjyEk5fFCTQS/SPy
gwzSul8e+QtnqOgCZApFgdDflFSIwhu9BXtr7/NlIYtfNw92o0qO55sql/UF5r0ZHOJ2kllUKjZP
i92HeJ/kbbpwMYnOQVSwvyzmRA/bpd1BKyD0dDY/weyE6Hw1kLhzvjobAJ9XaA4tx8ar1j6S4Wu3
O6ZZRc1vo72NfGsCvDtsiz9OzaVQKoSnxIUJnnxAh1Ub2gBhEvv72UkAqiNpuiQZG1cZ97+VrxNN
LDt8+RxqgbnTfh9W19NnE22tuA9+v7eIUHkJLQe/dYT8F/gJTy+yKn6kzFtt6B4cz59tVlcctxK6
+oOSn/AhFNPv0TsGd3AUV3N2xOkzAjQx7xl8M3gaFukU8JU+TFrmYXDMe1D/5+CLKPmd3o2gCsf+
QvAIB61TjfPQXnGZJyG3z6s6dmSpz3JNpGuYJJgLhCOSv49NVBLMQzy3Cx3PYHxWSXAYL3gZZmXO
Gebgxi8GvTQ9xu10WM6D/c057F4OzFUivzMLMauFcuRBoh0ARgmet9nfc1JtUAxyWoBSf7rg3Kmo
kg8Ly4eRjxAIpah3x62iOjWa9FxN6u7EOQ0R4o1tnxECsx1o3tmCz0/PMqQv5bdE65dXJLxG+hMS
1klDwVfnlHHpV76OsoovplmFRDYxeVQ94wkdBJ/2p+VeT0++JTO2t2s6K5sTfrm4lDV+oTl3gnbi
lZRYBDTWZ/rFzNrorsR2n9xZ094LuPxXHHdDSJTBMiqirjSjiufGooLZxL/7IGPPJHfqSO+j/b5R
W1Zohdlcm/yswuHGV07rRtpQgu5Od4sZ1/eZDFEdbKqyBJDrjZSjJrxR/n7vZ2tphcz2mE7pP/sZ
SpMpdk3EWh7z4154JXl8+86UaoC5NmZlD3sdJc3Vxw4NK2ogZcBjfZE0z+Dgbl937v9jVkzeFSVZ
UQwT7eNZUdIP4DBYpPsLWO9JATsrMUbb2rS5N227lNB2feb9Jq6v7YY4JkepphxzzQZV50a1k8K+
Daqk+S9v1HHKoPSupSkxPI+DpzDZfHWImnU+fFrCKQuWTk/M0A93iufwItNpjTx63LHAIsih6U0v
FJ2+7StHwZPtqQ6RXu+KfOcwO+K1AUvSGFW/h3IWXramifUNOdx/B2EGZtFC0962f5AAvZobaTe1
l/Na3/kQU5DmRj7uAKkHh2t9Wd5tQDW2IQXBJIqzUr7xXl01WnBQ9fdFT8PwcV8wyCQIFWCNG6ww
bcZEbYLwAOQ56ITVfl2v166QY1MMAgRX43LrsUhjKd6gxcThjMhU0AmuSmIm78ywTMkqKFzFy25l
vPeq/vHoQonMq5fof06XSOnwApcqQWwvhplqepfH+DNszeK1Nb9Dg6E3Q3G0p0kMQb2CuDqMxA2o
vFSAwahextjDPG4utpWG+EF2A/t2e7MYlP+3MK75qpI5YlM9bV85HGpCnE7RmwtGLbf6Dgk7eJjX
xY3EyTIOmTw6Iu+vocYJg09q+4+DrB76i8NVlOjWekz3TufjJ6mDK3ekQ0fsx9r9SLobIbftWdft
eDWDEh8lyq7b5UxXgKlMumxivcWN73FTDzzihURcSb9ZJcb82Xx+qiWqp1VRJUXg2Se8zWB/jEl/
Ll+7ur1fE0LCmeOx44DaUIhYdmRSjvuPzqcfgjQZy7EQNxYo/OkZ5lxStPsqeNTIiQ6YbWGzjkKG
se6toOsorq5lUBsrzrUsQLEgSOHswl43fy4FuQ0tmuzaLi4CVTgCvDWmiGRlbVSNEcv47+Wqb7s6
DPoX86Ht5vcPxlI/mNuZXWjE06uQw7nY2GTXvzRmlfn0zGVCBGFMjHC8ThU3VfYH6kt47tbiTEST
MsvRDD8vKbtREgiJuYmlz/30NTJVPFh3LWYD55Nst7UqujLlqVTqKu76ZD7srXK2MVoxRhu0IIa5
FFeoMy9ZUUGB+iwaYDIOahc5Qv4UnTsiiLAu6RVnOeIXz//CIhOq7GkaaN1aDIRQHJexBUKbOfCS
Z7Kr+RFN9R6hLFzurjovXvWfIFSv9z6PkEFhFkBkqQyXTez2Koydp1W5cwNxAV0HSSpGuAWqM1L+
poXwvUZ8dHFNeyZ7D6Ojw64C22mrJTYbbsh7g+pJ0MHZfLFyOvt3Penv3k4ff7visBUhfgr+Ky8b
+uk/KT5ERqPzysbTJ+WiLDj4EsNB3dJi7gbOlJeiWIGXK4k0JBrUdgKNWa3qZ3qkYgS0KCTqj2qF
ZJ2+/CHR2FzcdjeRt3HbzdsoI6GqDs9y2oow4SC5g16qpxEBT8EbVPi+PGDQ+bOvzjT0HabfsdwH
GiXxc8EriYHsnW2dBxCITC4x+h/qqSDFdOgrLeezj/y8aHVwWV3Wq+m8rERKgOavV5PGIm91uZAZ
65/NYcgqlQNzlk0VYL/iainmMu5h76GdH+YS5rIODyhjUeQkNdS+GwJMdHfdL79ge7I0W6SPUiuA
UwuyJ8f6PhmBZdnq5eDJxNhr5cZ/mMsUbDfNnrwVeUPQ413H5JAke1K7LZ6N6X3Z5FpXnOigUeyS
NAf7xdpAbM74t/tqcTxiq3C9ielOqlv3a+3K4O/HX098qzdgKqBuL34oJSrR2NjyP29KHI2ZKBrI
6ZSkwaCY4Fww88zvseOEyBI13162pcVNRUtY30XNUH6vIFwzmuLDML0o2A5FlTpbXq2z2yugdUtY
p4x2K55JuyRCsrkO76nbyA2MrLA3j/1bbxPq/iCskVWx0FWJO0Wv/U59HRq2PoCtmyZ34IuctLoN
AN9lHSLtueIwgKf7CtXVa4yNXnPs/CNiRLm5lrIvfK8vCZ67N9s+jSvSU+bR/YJluvhAv944Es52
Xrwh7RZ48Htnao32RtRDie71hK1RpipfdRGEflGCfLuIaDhxOm6Y+6612u6bCFr5YHLrh+1FDi0x
MYHYBc5z6gPgmN5O2T2Y8qL58fzFGaW3QINs/dNWWOr2US3cFRnZm1vhomVNuCJY4m2FjSPziHAk
5L0VEvs5M8sZVV/gtedYaVCFxzrXqx8tFjLWSvNavKlCrcmbjSI0b/OPqWS++A+2d9rUdvauSSAR
slY/6MOCVFvmSwj1W6RqeD1Hd9PanTmitr+9tymC1/a0rN0W+TrVbF1dqH6Ud9P9jcVEVURFzUOk
qWDzB88DgutJvqPFBpXHh9eUyvWFS9ZDBchDUYc6FUul4uUAGqywZ6LO3xHhsNSt2FIdNXZwlxC+
cKPWlF85FneM9f8xnLgoboe1rfd3CwJy2AjI8KXIwU8cSiyueG/kNu3hrjDnfbXsShRAuy8t11vL
ueuFWbQGA7OFwLbXXDJkYl9jgVOx5bYQ97+YzukATckPH26e5pnRcJTXav/W6O+HleF9Xux8ugGL
r3JyMBXiWCKl79fspnagLPqgljUKoZ6uiAzmOtZJCbtdsltKEnlpO68kc1T5ApnColcnI+/dDV1Z
6DAF/cAh8vGNckRdm0Ui0jUkHPSutYCLmuTFhX+RejrHI5u7elm8b/BBZ99Fo/HK5sukYaxMz7Ng
j44px+uMBy3DEOdOeu+LM/Uk4qEEuXliK0PQDqs+w0JKUN6+5eEnOBYCuo+jx2+dHoqMiYKaXoja
DE6nNLUVCmF9SDUabW/AkCPBkI5Llk5I+cLPzt74LcZSjdGXeFWhK+fkPl9YkVaFwZLNqAd5VzWX
P0nNkqPqfB5KzqxfKrTGKvVFZUGuCp1Gui9HJJPuKeIdVjbL2tlG7YdJbpmsoP3lGCSh00KiOfkL
KiyEZUPzaJqjvsc/nk27g/eX+i8m0h4YHcuKd2CBHfSh9l0Z9WmX4QKYX2jYwL4KG/3Pl4A69Me2
lkCXjXRrTqDFMXGJftk330kWgen8IakXkDP2AF3JBAMIUFkzkFtE7RDLVgJJQhfv7KlB0SbZqTKT
rX5xEvs7OGX5KgJN86yBjRXN7PrADqi/RhbXSFx8qveXf0tfzMju7DTq7ML7dUjdhUIy6xMRfx81
ewIEKIx2XJBbLj1UuOmkg9W0Onxp+kCiWiQ+nehKNStgBYlhp5SCHExLLpV511Vomp2zfBBgUL5z
UjKQF22ohkksEJuYYCs0t+A1AHIJwl+3ahDmqRq998gbo6VgKvGHAFcTP/rxj2eYrSbNTkAbhzgP
eTDxw/L4EmGJyyKqfOThMwiyUKKGfxDK7/27HTknR+nYq9b3ZuDjT7RTKkZ2cmcCzy1108KuXHVh
lAuCVpSs+CX/pEt6oOqSTvLLh93WJAqutC/J03ihetKvOPmuMP7yHl1F16HaNv5WP4b5yuKi95T7
pKVMhhFV0kDIAnYfkmkL96GcaRAztDlGG9bggf6rkxcJrAn+xPjP3IcpRx7c/bwZEsgsO8p7eFn5
uGHcWx1OYdLSJBBL4E1wYp5OF5YHJYVGugRRQ6q1/v0LXnBaBchTFE7FMkqebnLLfxTq8Lu0EaiS
RR3/K0MawEh4TCr5L/ZM7e+FupG0fFZEBnVPeEaw4cw6gXmStlwOAI+JnER00mV1GID6fB9AJ7c0
mgb1qWBWeHeMX9apljDcyNF6aYLYuHP924wSQjH8wtyp3JPeoDNEAPi8Oxsvc0sa7k1gDPvxohlL
fDLLncCtCUg1fmZQXIzCLla4cj2ssC+q8xHfEiqBva/YAfrC6AErMmlj7KYaZyGzeoUTRzuCtDEE
56TTrNo/QgMW/DXwqGZfXeXgpmHOgmRjDcrBW0YVjSBruZYQtdc7zqpnS8GQJrM/T4P759sWDfMt
VsAPjkJJgF+Rd1SVLVD9lOkCjnngrSn1Gc38tRtqkhIOmNQtj4lCTXuFc83emT5fk7j7TomA/NMy
77XlOYewr5CSVL9hribLUumzIunAiUh18R8vpdkqsMgjzt9IsksTojeDQwuOYWxsAq7cYXy2bSzx
zl9KAc9sXo/TcMqubykDc+MfLZfhsReKYGIAWOqp/ZznwnutO2qp+I519kFZiDar6Cw2aaEXlgHH
v4SvRsbntvtCacmM/0Vn1ZhEZ24b6bMbI2hG5BK+w+zsNyf7ME7lbd3pW2xVgZAniDDKBFG38fcx
z75+/BVnwJpGQ/7Cd1FG7JsPKyruGBqLNLVj1pBvlb3SbFC0Dom42uDJT279oGwlXC56915YrZX4
BB8d8DE4OQ+SwSI73fi6YyPkQm7STyXe3K61I/F91a5kn+nijiZxKs8rfeo5+QSkIJbImbI1c4rn
whfCtCSyps756g1KZjGrKrzswMOoBDfa+5aA2BaB2QCE3su6vgZo+xwZw+eN//spGoJ4CYTMsqQq
rkPwv0vZnEndbnlOMqVJWm1ZOW2XS/eTD/eVqrM/lNtyr239e+pP/DptQ9/VP+RDAMU/eEe1ehM4
langS2uik5nIIUGA4H6z4xA5Gauju3Vi52EnNX6wvE8X5eg9iFFzlOXcTq9dX9yeqXAL0VdE3SMX
hdNi8cBWBBjCMV1k895ku26Pa03rZ8I92K+jdrhikROjIWuDircDjbzp/S3bUsyYmpNgmOBrK74H
9t5dIftnBX+p2Sqd+8G3HCDYzjgm9JIqM6XmPU0HYkqNDMQ/rJQjcgwI2st9uHcM3Gcv8eX9C9Ab
tZZvSZuALL2tHWN4Ev8oeZjK16d4VDw1HEnEoz0U3MxTN0N+lbbsS6R0rKdN71tu1rlt/TToeJ60
v1i6WsT/rYLwY+2605IPx/hWqVBGQfLD2ww2tKYw3c+M1ujF0kE3pYSrpN44RWbbH+ia5ItWVAts
oI5cyvug4J7b3alJSzhDfdc2rapUWPMZDYRu77jCEl6mDn7kdIy9UBAEP9HbgmvcY3J3izeb23mG
DeGLv2NDWD1pgQpuIM7NGn3nid9aeYnUTZ2FJyIgTy0Rf/Ts7z6s6SXn9qE6CZP1Ehcv3Do9P2Cr
BDD+DO6MuZZqhenZX4mW69+GcAUvazZjmaTC/LjO+9e3qM0flmA2RJiIkZIu/dWIo22C6xsa9Jgv
/fQjB9/PS7ad4s9XooUYJJNxIN0gp66G6tx/8z5AXjbU1dEdB/TveoJ0uJsrEzzPUOyR+vw+c6PB
FzUHrpuwn4EHQui6+Mlpt0rvMnSsZ2OmtoMvdX8gl5e67USrAH1CI56sQs3DBs0r7hxVrUF1Oov8
RYUZnFccz6LOQ/oLY3KwlEwnwR3JmuB1kEvbMRUglmVqA8ZcZ+Vxc6dvyJIS1I9jH21VO0Z57lhX
SZBxA48XwEvaYppNi/cru/OWPArnkj6tri7ME0Rua1bl8jn8bcclE579+MgrwITOt5JtLR1XR3Xx
umh/5mxk3E0wtTRrIvvkypaQr2iEezAUAWPN1ToZM1HMEfl83p2xp54IfVprZPv3uC24DEEFPSTZ
KxUeZUyex975B9+Naate0qEVaonFvLDBfUjntYNhxfK/ajLtTJ06opmqNPrc4235klJ66fM/OaUt
VTCIvsgcUxa3/0K897uu5nnrcTMsb2qT+jv3Rfy38qSvwZmdBqUxs+gmPYnMLBIpwvXq7GLkwefV
zfMRag1y6tUtbxHv7ZvRZOXrd/aCMA3n92S7PT5FWlyj9YWhOLn+ghqHyGvF9s1f8VmZeq57VamG
tT/faO9cz+U/YDrUridENdMgMjzASVV8AHODjV/g6g5qy6fR4pyBq8j662I7i6iay+WeZaqjV6Na
tex6Px9wH45SP2m2XG5vbuulUK8TCGcxkmtn4kYcBcr3aen25/FKaJau4+WMi/iyc8rsvCzFTfZH
YAbhVLOVB4/DO9kBqIfHZUruZgfXBLQ5rovnUxcAx8MBuUMcYZO1QmbCuaisUOFGMAUkpcZ+9hEF
YLR9n0xdI2PgSQw3wMN3E/V7PT8icI+CB/ECWq4/KeBRy5Rn4mw+kEDQJOVAIA5cp9N1NIb/Pa8M
nldFUDu+SK/0r5SYLDwEyhsbaCN94YUkq+H+kU7gqKnxK9wnhzY77uKCtFQwNT3Hz0XQ0K4HuNe/
+hX1AjtjwcXf7iorX4en3vkHFrdgX/itmGLzGqEMyh+0+DXHkL4WA+NF5UqDztH0tnTvlwSf/YHw
yDPzQ1VfETmd7gFiJdirJ0up10YA2qJfn+9BRh/os3M7x9aEEaE4C7r4M/xIeI7wNPmUxJhrxLwc
E1k3vjPAgzH+myCnk7uwUpxpi4gOER68deEoO3jwWxvagr8w0Rvk6l9+aasefdmRwPofH/zwPJMp
FCrjAf6VrHZs/hwyxI7Dx/9/Ek1/wq6HVk1m2em46tc46E9+bjA6MxPMWrmvWFxYTQCZC/yoyUJm
4hJrE8LSrQDf89Tec83/LmMPC6YvHOYLR3CmqVJni1p1E84yLAa+s+5TV5YBHJCg0wtRDlLvZC6E
GF287MB0nmHVwneBOZIib42w/Le1tcxxY0YHBxtV6CQzQttLEGojSh6lp/LweCQw/MeCABmBHbEj
D3pVCx1KxWjEDXuE/28F6+8CDm0TegeThyc/gQ+pbzRzh9VywTD73wz3J02Hq/KjtmuKH66XBIe5
ZZb2ant1S5iIwOlVAHGqSUEaOTymYPj4nOeplCDH3YlRbVegu59XnK8tB42HRCpbbjOD7+wFqVUb
XX147qeQ/Kgfw8DHFBxCcNL/Fj03OZwYziyUHGSaJppxP5o6yfh4A79t7cvULQ3F7dWhQpy2sSXS
r4MmZ27FIZWHIczn/XEUeSAwZNGaMZIf/g7cNLnyAtMThX3EAR0+sgo9BHVhAWmd7wwbeGEWaVgL
7l/4M5Sn+7oUbaC8Gum297PddO8r/iqfrtaRhYih+OEu3QWGu27Hd37kz+8YQ6JeBVqCEWynW/1Z
xifohzHQM8tg0hj/61ebFRseXsxKsU7o3rTMHk7TJXSHf51f98yD8F8IcvD0gEEZ7UpqSR8rCUYG
dAlS1vcSrv3ON/nnWUe10ZxV/+M/ZWohQTB0/9X2sTKwRDAib9MPWa44bdmfh3PC8di0K8t38Ct/
cyyywmBVBGE7pSjx70JaNk8WTj6J/EWpZadkdTNCnFJxKiJ5h7CivdBU5y1Tq987jRN/IoOX0ILC
U8SQ5wKLCYNPaNOFthYejuaHi08aTz9ufkbeyLulquwHsh2XsKCjlWTLUzOl2U4qqfCQja3pfo2X
n6y3ffw56bHpQ7jbxICGlaxM2oaVjH5QCLIHhkJ7fxBSU6xrEyG/tDcUuCCyZut4JovTpSiv9PKZ
uHYy5KsHoNaP6BpvjgnNhSNt6YUOxVTW5AoZDQv4wd99dwcXZcVQWMygCdh1Ez33yU4fDAruP5M8
Vr6zsx8quXFkDcWwQEsn04K4vIWknCaTeXWHF7hNgiBNGJhlTBZ4NTMRpGhjFxWKjcRkUT59RdQn
lcNrcVFLLUVoJ2+TC6oOABgSisCFDeOEEWwOOnJaSYMOHOcvYYPpzBBSgc6Wm7zwJRSNifZjE7Ay
3ytx/6x9jiH3Dph1vLbU1N9ZC3vkWDEvdV2Dxeh9E14a3TgSG6cNsgJdZOB5PgOMCJjoZzhQHQxp
c+MpZpbSPMG90WIPwsU9B9XsNR5dIG2hfWIf+pB7NjdleNVLJkHe6oydAdo/zPPvXiM88OF8Sdv9
t4p77QrfPR/7FbLaKU9iHNUeoejVXM1CQtzgxW4lqKFtdSMZkO7HOzsC7d78ECPXoOMMxpL9f33r
jZkS78iFeJd0X7nsjIFoXEUBUd9C2TTljwgDzO4HHaHlN81MttcfCLUvAkgiUr2476iLT+MXnK2+
d/qoM19LqPzKoFhpoSfMnBT/DyMzr/ptOlTWjW7fngio7hoQirNFH6tF+cZIuMkp3qwIheT6Wqlb
LMPbAsnPVPg6U/bjj3njAUD6cVya
`protect end_protected
