-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
k99Yh8yTDGTh+04VBQ/2RF8ukV5rc5bgsjnVKHfhWkOqgr1/Z8PlH0/4f3ooy4laP6MuZxVIEj3R
yjyLFtLx1LqpojcP4XJHBWnjtlxIPf0LPOb7la8DpCjtO4PmOrczqymWHLr6bfkbBH5rrbNvA3XT
GHuVKCpKTOcJ/0H9i1hAs2Q1iTnLvH5ye8T6QXwDgUzc8ScPa5whhUhCapNR7ClXQtL00y0YJUid
KBeVMJJAOlFKg5A6jKpqgs27tqyOVANmP9sK/GYnqMjE+jY+pJblgHVUAgWclsEao5GI3LcStjo+
Dt6ZRVba6Cmc2MJAlSzf68edbSCC0xpXKDqyyg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6656)
`protect data_block
rgN6CWbKp2WiDftPrPNiF/Py0AwdMqI0goA7HAhdqgZt8z0ujF8b4wJC8gb6CTIhn83KU/WseNa4
P3NW1B5mIMp5GexpyUht146AlnCzBeWG8q00AxvEgonQhnN9dkD9v+zDrF4qhgEz9/p18XOsuGbh
Y91jXNZgMydk4+dfqe1iJnpsIQAxKDfMRy0SaUI879cNkNvp3tw9ZoFNH64XVnlVGFqvu6tQn5ud
ZhXXOuvytxkH11maEf9JdM33PIzxJK8xzMEnr+gjswumbczoM46BoalcIlHXMesBCBunbeLQG7bE
8bgpsv0kGd4+wuvGJ2zLqTf1LpaLlcNjL4KBXBKrexkS6dyG/cN7LbeKIJJliTHuyLwIZZ8oB+5a
rYVsi02Iu+MWzxo6JaYSls5rxwhgi35lzFums5kJXPWrvZRvJoTjhPQefZVb/wg4dzZuBg7C1K7t
4PEceLm9L7GtDpRgqLhmKAk5/341fl1mcZ/9PPONu+RTr58n6Bw16aUaBIFOT+CN8uLAovaFwOMk
GQBIYIgP7vzNd20iNRcOrmHylDMPsv5js6uA6c+kEDrmchlFAZ698Ay3AVRsktFj703guco6YT8F
4CdXgta1pEjAr3/bq5piHUkTo6DXFIjUZrmVIYfp+dHOhwlAyLYL/TrW06byigtvllTN0uQSWuVA
WdI8U24oI+b7CGIBm7HoFoLBjTD7Lq2lExSak4R+i8IX3oWlYeX76fDi+qrpHEDHm1myHviKTY1y
YJMvbCO7UTVumVvaXlv1119Fo2BJLIYwAyhzLKDvNvMpLfqdWw9xImHYxYDrhS420ofCyZ1e/M4s
Dl8a4x0BOQRH0uAs4FMGIp7vXBgZxGHC+cLHHiR1aUqe+dxvHnJL5E/NB4Xyx1wbu9QrcbQhMFFH
Voe6vMfrqyvOoI07OqQ/Yo2eKDvwZYWJQ3VLQwMejaJECDSBnhUARHMBpjA6NShJZ1evqc+M0rVN
E2KDYajCrdU7HIGAU9Hc9JWbhii+KRW06VDlIoxlqg/BFr3jJ/QJNHIRnh+MZOXWDwEf1BYaVywk
YhohNoXwO3SVcm2J74G/6xy627Ly1eXMqsvI7ToQKnGX3bOQxuay7QVSMyLZNxum5uWsWD/ij66y
gbyNJUgshnVkX5d7A8KuDsXAPe6qOWlM/ZyjjAxhCR1UXIvCVV+0wLk3uBumIBfSXnbTfkNzQtwq
ZnwHvs5qobt50DrYVYPRj7Ey6crPxQzEMYhUA/8U64fvjqj7w3TyKgmVVAM+f/UCmZdrEacEfQcl
SHRUwV5AGs4XL5kMEcJjBg4Oab5PabOudbELDDahEcK8iDhWTBS9JeRAO4ZAvccqSjeqyKuFyvDU
63ewyXWvTftt9a9OuvHwADerdqRwGqBDwEscskMBg9ecsyIj+BKYpswGPz05Mr0KzYq+Olcu+e/u
oTE+hwoYPNojd3ZrZnUDalV9PRWnOR+UlFfmmAuYTfAH0GlLqFdnf7GVoLAiav5j5bHj/DLpjWJI
232mHEGAFOxWkEf6BYhWAfw3BzwCotyczNyA9dE76stPsxKuF7fMjO8a8TDTw2NdqTKdmOadrkfh
3n9nIiwL7onYsdPus7C2Are/y0Vv9di+LgxwSpBjGX+wFyhI2bUYW/3q5WU8xOXKFlLlL/xa8yIH
ZRStRXlBJuJPp+mZodxpB3iE24nbWkQhYN/6VenRuj+gd/oybsov0p+1pVYj3leQnfZZpf4FAuM8
ifrYxrnttquvj2qZlQZuV/WzBtAJ443FSJu9mohWouWoSZ2KogURBkMkFfFmDvJzXv3ZkItvpaOH
ZbhsQblU94w8h5UujzksBc1msAmv2Gd+ipWMbfozoOarpCQRpFwKCZq6wiqUQmBYjhdIQmzfCnd0
ba7zPiGkzOVts8LAvv2kjsOGttt7N7yQxkAlms/EQp65IDU2GWAxzHBlWZFEX3m8HA7O073jeMv4
X3fEkoNrfvTP6MbWYvlfu6EjBJCesGfyvf/0E93hN9DTLRC4r/zCaa0wXeVO+BnbNFYZo1HwhrVy
zdAaehuCq/ITx1qwGwaEcfhmTMOKBdbBb4fuRE3Me2Nc24DD63agsIT6hrC14ZdFMMhr9PK25jcT
spA+aEmLfCB3WVeQNP456DAotCliyTwBDQX4ymRKObRp545xkZZk3ZTFjUVziv6tVNhWQIUnH2fc
1xKXPXXjRJjxuO9rI6THJWXaYmLzG2vPXUemLT7TnJKzAWmxSuu7SEB9QMcSmguGTDVT4RLuA29N
uA1EqoWTTTSVBYF+Nc2YRWXfwBphP5L8tNsxYU2/5FTHg7PZsiUSe5QyVbRnGx0O3AqPBZFlqFfW
knWnrea00HQJmC3BQtCyeHrHKzYGJgsytW/vXjhfVEd9Pd3obqkZKrVRzHolBOQUsuHy3Jvmokfp
echG7ydnG3R1P/DTPsCJa+OB6kYSrArq1y1bYWMdM5G2Gtb8I/ELDrpXBP3CLV+c7COYUPSEFTYh
ruxulbQpskn8NtpPtsuOy1NwcLgI5YHR5ZLp7wzOkt6MvlFIYySeQbqdgGi7ylCBoogotCGl2y1J
Og7GRUjxmRea/kQjoGsioDiOo40FqDTncGgHr53uFBraVK2E/4gIaDQFYa4GrQpDTdVBvL/1omfy
kjrB/Fav9dmiYGXSu5KA1qTrhuVEbfFUbXlSXwz2yOHZGvpyzmds5W+6ZiOdG0bOCkdNodEQgZyX
noxKgfMKfJrV40s08FRRGesEpG2/yMA7IuuXewQ9J1sQ93A4MkyWW/vE1wG48fBEFWqY2kxoz8sc
aA4IDjRIG8G30fkepUdlQ6oaSbwnY20RBphAH1civBpVGPAWz6PzC2wdAT1ngOW/5kIhu6ZRyjLk
cif4Qw6U0euPIhhCwBkOpWzxOZg2j1b+Jyeo0XrjyLx7f96bggobpOl+usgtU07KwjtGXSYy92kr
5BZSHxcXWkwTHC4wgfAnzzLa42zxjB0A+wck5wgjh2jKTX07I3nwBl7Tx0181LjHwSVNZztQRMbi
T9tgeInNH8YIkw7TAdZ1sbjYFy6Cseo0AshLEv/HdrAwyCSQ8lv7aXEVEBMoXyVOFj7MDFGTmATU
fU44vKnfFXPID4afoHdDIk1wKjyqZsDID3YIxiI4IIghAluqZr3jigLjuuU7CO1qIu0CkCMgfJsr
KAYMQ4DYncOTNHoF8TL9YGGKN/ZtYvP+TzftBHHG6Rh1cNJGrD1yCOdyyxY5J2EN7/XON4qCB65W
wVXXiz2zaJuLOnCmG95Sfx2FFXEQvQ+7xrS088STxljil1olp5nQNC5IcPXXPE5XfN7A1TOf+Cdd
z29CZ0kP00eyg7lUtmnCPW8T0iOJXN/zxlrfYP+yzDNvXmWZ5/5kOFxUjiWtQRzbpn8ih8XgriP2
ohHGk8VPcaWKsokFD6sjY8gCKLDofJpKag283IvSAEkTvYdgub90VOjahqkz4CSPdGDJufAEVVLZ
Tk/LWMf4kfZG3rshQ3CIBsXQyqIkE+p2vkA4Yv0ZZyiPPbK+/HlgUxcjDy2f2vTIcliOeaihiyZn
Ur1vRAr8kvgz4kGaCXI6j3oDj4Guq2286/gDKbP7FbNbGvZLoB/aHwSBSUAwEWSwOyntqtgAyGnT
CpA8OIo/2DNg6EPdIfXH9Gehaz4AJ9QfECANlAWTcIChWXyVOlyzyQZjaze0APCAZ7cqBs1hMb3J
uqXxWeeNnv2lzW1Jsjvzd1NcWZv3sEvnsY0j6JpHBo3/I9+xwR1ahEsrXcjJhN6VugZGO7A01VWP
kMqr12Ut5+pcMl5Bh2wS+A78KGPjQKgvyySRJz4MzoL1rXYf3iALxpGDhJ03ATZ9GO/vroWY/z1f
YtP0g/f4Q03szLtoveH+r6IKVfcMWQfUv59WxUckpReXoMhFiaspHSUXH85KcV1BxhZ6KGM/W+xm
kO8uCgWUCiPVCzlgTKRW6EO+UAsS8OKzxxOHU6ARptx+vAd2Y/UVUiHQ+yZroCvVvUXDl48BDIsv
I7/hvKP+al6+ksUxHZ47Aq6NT8Z4lWWE3O7qdanQ0NHoNlZCTUgNrCHLpAxAmILPWkppIWx2CCib
YT/1sUR7Q7oP/h3drbSJwkjNmr5htpMAo7CXECzFyqvL8t57eND895Urk7CxMeiAkbqOxOGzegZj
SsiAiNl4sfga8+V13jCfhHshr1iNA80aVaoE6RCMF9Ba3oQJZf38bx0PoGqd4TPR1pF0a5VYY2xf
arIVvK4liuzjvx4K7AHJM8k41zm1w3no96yg/XoBbllSmt1I/VIwHvXmGh3lW+Ms5w90CEMavGyn
WqUy88FSilE5+Eya5J3rbVNooEuSvc6ZCkZjlUGg/OLSmP2baimNlpuVM45q4XLnGGhKEJFAQ8BI
pHOMtZVQn8KYU+tnAVpLcKvylG0Vl/BeCwaXnBLWYr8qBrP+Wi/GwyvdcWiuhWv5czBw/1AMiRLo
rp9pdTuxzIOtkJfzoi0TUwCL1efNc5JKtPhhqhkuwa1jflIrYkn8moTPQzmtsrDeML5M1sxQb8mc
NbOk1z1rw/1yFWF7XayZ6gcXouADKqOjPy2jf6WIi8lxmWFzVzTdDnj5/H59LDSBx6zgLparIgyD
Z54WD6PYZSUb6+hDn6gXs8GjTWfsf4i4Vh47f2Qn9Ebhj0DFLxipvip/mJ3dUZhD6OG06yGph50S
MZLFJZuHvbl0MGFqrWYEGg1prgIoa6KXq4G2LWTn+9AmpmYOygipWRNwEp/QOwDlPvULO6s/a+R2
8DQFbxJ4eqsYGh0qOExi0gjHHGoCOQyVjDZJQj81UbGWHyond/b/lbt/hmO+BP8SrRej0TGxXuDC
eKNz5P8Gw+aIdT9jrj/f2Dx+hAe7CbSpJmU/gXAKbmjyu3Kn7nkB1E32nzmeZtArPPEaqwSpsAHX
ke5tJacT1VqojelaS99NbAlp+Fu2EMPfxIjD6mq0VzAQDeNX+c7ihW0AYa34np4OLZwgMGn0amSs
XydhkaKYpzxvi7niK+JhcaMTpQzuVyeePh2rlj59bK9vbYwMxaV059lImXFljG9A878DGsVW10Ut
BwZpUb5kNkCGN5ktFHhA9AtXcyMlV8jzK1dB8eNPmUAESL3kVue2qP8SheRZ8msjqDTFEbGXXmpd
yvrj1cMKg0ONb1GH8juDcweS3X7RnzuJbVKqPnLMR9ZRZIwVZWhiPM4GT9WDFxxeY6fsUaHHtF52
71AMECTKB3EwyQF6zz22/Mj0nyBLKEhgyeGei3JVvL1AYixQawBfbtkRin01sdhhcgJZfZZA9Tcj
GZFPRDqzoDFa2CHQvp5H16AMU7PkduWmG/3K8QCug5Mp1/pFpsjhyfKl6JLbPPQB3g+GVZLgM62N
+J0i+bG5vIyqlDBL0VykiQZtYNme9FAge1UUskZ2jzHhZkb7n6lPeLEmH8i+3zrkpXrt+q+33Npu
UlO1SLnkMcZkl5mdsUXAtxehQx9t7RbhenZHgcodV0CFzH0aMA6fjnvhXchwyX0/zxa2O7tgwLI2
+1bSfL4rMTnLi6IYqLeNu8pHtRGPtZSBVLU+z+c1/8gtK+yNm3nq0VimXFWFjLAoAi2hAZYNEAGc
RhUQMeyolAeXEgAjqfJiZOJjstFNyv/bF6sMsbcX2AaZ412O2pCOOnmULA+JuGicCSOM4vD3CQBs
8s+4XuCBQzHWInr0oszRCoUL9df1MFpA+CGCRBBWgVBTqLfFSUWQW7ke8QnIxnfdROlyzLN62iUC
x0khGlvXcx7LI3JvzoiA6OqgcRX8m3V0rDk9CaDJpmiaIrR+PPLKxYZv70yBS1isxOFkSnvkZumI
tj6QcfwtRnc0xqyyISOlInxxVaBKqz8HczAZozry4PXgInR9nwsMCy0UBxB7PTgr5mqJpx48GbDg
ME/qaA/vVDUQrul1Agw0TNCpdlWLN2mT7ngVceblUcF67RS1KWAUF1ga2Q540Wv+XQgkEavyJobo
72C/6y8saEe4zh0/z+yhGpk61m+xmMbCJhsPW83D1QcjnzoUW2m9P9VP8Rr18ErWoUMAS8ElXkxq
/Ea32ASg/DA6Dhhm4MBqZy3DekP/QqmieudUyfGH+DfA7JkptgCUiknrzzeDLGdXcYwysqWKUpEX
FYPtm5jqFNhNIOhfJ4UcaL6SRhlltt4yr6lP0EbMSFP0nw53btZEbEaiQ8YNZTlZVpiz8ba1xA/+
If/WaA0LpBb8NdNL8BaCMqY81/81BjiDB4eBdLZS1wvHPV0fBsvpG/Lw2HCxMyjUKlpd79ONXxcC
T4qHUn6a4JhtKfVKkp17PYPAy7+cKdQfeHu+43Zz+lgizcepWffO+4zHKcWC6rjM00RrMIzYoXxT
6AetUu0mK2D36iMiro70nsekaUtJzhAsae9dd0DZMJwr3v9shHaD8vCwItKyL9fE188qxKcEEoGF
jkpvtn08TxaETunsHQ5yMn8nB9bng+i0LVnaWhGJ+fc5gBKpln82qdQW1CiD3+yDGZFg8wrDbD9w
t9BzVG/zg3pIr+a++nkBrvl+zoikiRza1j8L2yT6HziEidyQxXaIEo8xlyQwZ+fKtuDKPD0uOjbB
Pt08z2tj2J0Ym3PoovnN6SPCmCifrYjFX58R34vpdaZMVNy/r2fgpr6uG0vi/9XJq4nd7GJTvQws
Fd1A7J3r1Q1bJtUDR04RmV8nDiPBJ3YtXWLVsPaURa7jTQ97UxVlq5omHL32Z8Cb7LnaVvpNA+Fl
OVB9GPKBAvpAJgofmFIlJMCXXf0ywJux6BVJGFMnx7RE9SwLMb2FEYiM3CR3LjRZkWrJ5i4axOSP
GYaxUtBNBD7FJN7ZqVq5UDE6gcooOVvARBj1E9ORRstR+Ust54ZP5xBW3cX4Im6vOxGDL7DfL0hF
u4zg5WTuzv1sP+QP4pbDwviENMjdHLRQq79ztXWG9/fflYjOjO3lVIigQlKRyUUuYhDQ0n8a0tmb
qAVgwFOEKHjYyWfi/j+uJUfmudL98dZeVXWDpf8drvYSDLw22KhRh9ZVT2TR1m6eGhCQOVb8i8wK
/BCQPfkqDaXJsip/0WWbgv04DahiHCPML1jccauF8i9j3eZGBJv9ydhxRTPi+yLeMy5uJi/iM56A
GyBl3jUqPhwH1FZiEkZnWQb1KKr4PWBrN3FVm9anwJPfoA+Mxkm8lZdG7HdHj+xLvRX8qMpQLpeH
INTYAZI3gud8XUumGehzxAGEzQnoExNRXIFt8JQbAlrzNUVRp6fjzZn67KYHvozB5Wfxj+uyQa6/
jPHTnAHQ/q4B6+2tyyN/2+tRTAzrVr0IRvYpwir/AY10wWSU6snUbBNPfM3LLJJ6NbPFjgog1k2Q
luSAEtnPSq3Vk0GKT8lQWZT9hNn5Pau59YyGqjuJM0WW+umYhL0hG5XMTnLlMcmEplvFUNf3ADPA
3PGdJAEEKBKD/kGjJfprAMzMTyDqNWlqRpJEfjgihB8LD6Socabg76DKLkzK+hlZC8Ej+fisNwGx
MNZxfQLRUfbW7BmW6AOxRHmY39EG6XWJMIsqTIEH5TJKuqRwYYlUcHD25Isda3wgnEiY0NGFClUi
MhoUQ4TbGgmRd3kZjQrN7qgE3m5GqIjAaGs9YS3uF5M6v0WF5LcCSoaZasCIBnaEB2WRxvUylPJW
B8nvEjdiAv6K7I8S4R+a4xLU6OVpmoP5BOsyhnAl/kAGYEcOQCk9h/PHZyH+OiutrowgHshjcuwd
Lh94VsJu1nNtjSGwPt1GXhRpWgnjLz7k4Wm8qwkfkRuz9Ev+omRjbFNyxTtKxtmbLxTW7FodlTT1
uCEuO5Lyr0Nw3vlwOXfIgJHzLy/lC31tjXn8wTLPd/2xhEd0Ech3iGjm0Qn1P1NnATNTdl4zgiDr
aMqmSXJ0MexHMJ0LIyXDWL2my9Z+rDkok63kkrztR9WQuDk6yFwQjRryXVm8gi2NX3mdUO5yooQa
2c9dx5d0rXVAz0SivWD4YvPu4orYHTwtSYSbD7z2NiVq9QhtjIbLXG756Cv3Ie2S8DWhr2bR8ont
5BGrnHgSO32kA5VzhsbF5wHA87sTiaAyVE8cy1lR0us8AXY4fe7mGUaY771XEeGXlWCcepf6dTKa
U7Cbp2G3G4qzCWFUU65XQIyDq7ct4pERrMpmbnnnrTdgu4SL1AkCPFBFXKe29IwwuplYMyonI3Jq
lKjKBZMSA/51scVvyvD0UYsIf4Okc1/oPQIswSiAa3NCwRw++kfe6otqF9OjcvYWmAbb06wUEp5X
eon23S1ez/FMcSvzAGqZDEJ/HKbnvJJn5Q1D4lJRmNYrTL4sLK119Doh6CWzJmrhbzqCWm8Q/ZL8
d/L1FdXNeCRpy988BV5atzw4oId74sClSjA932Ko/dHxRVpun+6WOnQO85j+uqfGgJyuyBMd0Pxf
BuNbH1WwrVNqnn+ppW7y9xHfh5pfJ3KO1bQDEyIwb0koTOwhi+SVRsi/lKgrjT7EYoxuQrnjdZtr
IycHhV3lkFDht47B0415/CStLaH0mP/vS+z86bBPsEPL3FN5JlSYC3YcznuwpbkweDwaUWbwEmw/
ebACxCqqNv0QbcrzePGhnbwOknXpdvaQxOQeDfAXE0styoTXBt0P1Q0oG02RcSBd5SxBjq631RbH
nEsyzY6gHMzWPDdyqH93j6ux4w4VYHkXnvcD9XsN8VP5Q+3PrYBRsCmJOuE/BURgK1virNyXH1d+
cCOr7ELXrlSeirwE+VerhMVX1w21afgaAF3Poda0Ct2su4UhdBLRq1vDr+5ZJOiTZAfl85sS+roa
DFx4XXuPb2RAnM+DpyWYlRD0sOJe/OPTfBUM6wG9jzuYwuoF6HFuDrJqhts=
`protect end_protected
