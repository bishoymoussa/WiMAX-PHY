��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$Rx�y�<��wA�*;�x���@�̦�W�X�fa�M-$u����n~�%���P�$��W��kYَ���P7�?UMfT��q�6�U��k�>����~�\N�(�����X�e���/6U|)�X2pF�]$h���d.���9E��WG��L�X"]�Ad����ľS���8od����e�GT?y	7�������ݵ�^��R�q^]�鍦�����s�ae���h��L��P_���ާ��YЭF���'\��68�b�[����w8�[X��V�F�0͘3����q諵�uW� �h�u\V�?@��_6G�_�*�G���B�絉�f������[�G��U&�����~�F��AׯK1�`c��[<��FY���4I� �#�G��x[X�=�Q1��`��R>(�w����R�O�?����7�,(�H\�#h(W�EH=�������yq��Ѿ��aF����:�U~m<|��.��0=�P/���4ǆ���T(���q|�Y�|���/��S���>�*��#�@\ڑa2}�E�e��'/�v�ֆr���pz�ᮆ��HQ����:\�4�7� �P�t+>�	i�"�w:Q�o�Zb�4��n�ЄP�	�0����s��	S]�.��� ���0+��b��$�-�Q��P�8^���1&�`��kBO����6]���fg�u���L���b�FQ~�������L�8���f>W�R�m�f6/[
Z%���k�3���ф��Hg�ll�CWu���b�0���K�$��J����)�V Eci�Z2�G`?��4�G�A[�@<;���ڶ�'��u�'����o�)������n�u��WLc7
��B�����`�e�DV���~��� �����߸�F3��i�s$_{q5�{F�	U�̘��;��y�t;�я�z@�tL����/g���u�wj����#O%֖2��ht��X��L	W�_2`��|��6���m����!�kF�Ld�<�b �y��v��	y�������?��H'[/��3����|�~�a[�J_Oѷ��욿"i~��Lf�nLg��k�E���K$���gm�y��^�7��X���!8�C`��+� W�B��z���*��|<��WE��q�Pa@�ʹ����j+��$d��e�r�_Z�CAf���ӻy�\�XSkG����Hm[̌үd���wZ�l'��E��U�ɰ����vI�p'E�1?6�,{t����><{cx��-H^k?̉��W� M<��ʜU�Z`�^�<X� ���f�5��7��7�Г��6ۓ⍳��0���Lp`]l��m�3�����U82�l��b�^.�zL���5�~� ��
�i�#�%M���k��o�պ��HY�d������fq��O��X/%�F+��dk\2Yz9�'r��Z��U�jjؚ��p����$�4)茨�%�\�Y�p������r�_>��P�.:jڃ�K��4���xw�;�ɬ}䲻���	iX����l`v=�d�]�D��_<
�~��|�"ҽ�����ik?ރ@�3ذ�<�M��%�O!��ȴ�<t��8���P��U�*�oiZ�#˖c�M�F��z���tއ�S8�&��xCd�N6A��}?�P�����[���b�� ��+�����_s�c���͂��k������8��m���V���H �r*]Qc�8��tf+p�I# -��w8A��2z������T���̼cՓv��B�k��ÈX�۰�܇cQ�t��ą�|+�FL$l�J ts�j�h���a"M��򐧠���AgKd�B*U��r���?�F��Ta�Žಬ�ႌ�r��L0d��U�{"bs�E�UF�I��v\��n0�C*��jZ��	�ɷ�Q}�u$t�RaJNr���q&긆��K�Sp���?@>,&^<�fl�Fs��N�PYrcԿ�Bۖ�_��G�ܞ�����n�63��c�7�Gb��R