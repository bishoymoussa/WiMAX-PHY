��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$Rx�y�<��wA�*;�x���@�̦�W�X�fa�M-$u����n~�%���P�$��W��kYَ���P7�?UMfT��q�6�U��k�>����~�\N�(�����X�e���/6U|)�X2pF�]$h���d.���9E��WG��L�X"]�Ad����ľS���8od����e�GT?y	7�������ݵ�^��R�q^]�鍦�����s�ae���h��L��P_���ާ��YЭF���'\��68�b�[����w8�[X��V�F�0͘3����q諵�uW� �h�u\V�?@��_6G�_�*�G���B�絉�f������[�G��U&�����~�F��AׯK1�`c��[<��FY���4I� �#�G��x[X�=�Q1��`��R>(�w����R�O�?����7�,(�H\�#h(W�EH=�������yq��Ѿ��aF����:�U~m<|��.��0=�P/���4ǆ���T(����!Z?^M,!8�B7��m�E��8LJP����<�7l��?Vl����V�-��x{�T�Tx� &�~]_���H��-0���� #J�IO��n;�z�}�jЄ�f����!�E�T�y/��~�T��M�m~֫�4��s��ASCA�1�`�iC��jt��6����?"&|�U�]�ko��#U-f>�2�DagL����Hfuʛα9��u�h��v�k�-u�z���v,��V�\���eܔIM*�C������W:]]c�����Z��Z���^����CΗ$(�}aLg�%�t�X�[�]�fՀl��y�C�2pvuC�Ԙ�0���Pخx���ݶ�'-'��=��P5i�����`Ru�9�(e����O�Z��e���~�./�.�8_��(�*��1,�=yt���^����R/_d���hƱ��� ���b�Z��$e�*W��Y��Ai�>�ؓ¾�VH�kh�ƅk�X~�'�`d� �o�3g�7Q"쾧���`0-��@<E���|��U?�O��oc�Ϩ�od{��/�\�1�2
� ��3(��Ə*V�f~&ǠP��l;����3w�x�{�J�+���],�3���<Ե�8�w;~�ƓD@C^�p^��.��Н�Fte�����7OsD��÷�%�~$�7ҷ��L�@yKS��9(�*�,ݝ�G �ʪ.��{;��O��;q�i`vK��7O1'xS��yP����P��Z�g���A��<�5��m��׳�Ȩ�jv�oaj��|2�d�t OAz	t���L���f#P$�v��V*7}i����T½�ϵDY��V��2΀(��y����|��Z#Ԫ�4�Wd
�(P����o:(->?`?*�n��At	M}�=��$/>�6�{��y��l�:;<~���O�?���~�Z�d�>���"���¥�4�K��.�펞�^���@*1���nv�5h��E�/X^����u�P�Ӕh�v&}m2ځ��6�	�vu����}i�}셶�%~����@���h�4xVH�#W�K|͇��cwf��Ꮒ�Z�دܢ���B���,�.���^4�bG\�V)��`��$E�g7W����(e9G�3s62�����wD�v�V%�i��;�\"c�Nɫ0���,�~<oW��թ����A�n0���G���#��lk�~,!��>pͼx�d����DqSX-�F���q�Q/�X�I�'�O �)�x41ڊ*[D��#����0��:=_
h3������/��$�GȄX����E�:��z��_��0/EkD��+8����3ǎ�<�P�+zA�5 <)gŗ8	G6{�^��\�S`��߄���!Hfi���M���D%b���q}����k{�f�'�O�҇���`�r�=���>�����.�o+����Etq�{m~��t�Wgn��g;D~*�Ҏ+�r�D��.�r�������`2M��4��,$��˹#" ��`%ӯ��bGA�nai˕E������P�>��|��g�e���k�{��K9��Q 4��#G��U�#��0q�2���("�BvL�����T2�Y��;�H�f�Y�	 #�=�5:ɵ�o֊iڅ?bH��{�܇5�C�v{N��6�9�Z�-���#��.s�-!�'��Q��)%��`Vh���D��\����&Qz�M{����:
2Ĥ�ڝlԧ��<E�눶;���H݌+��ʠ����з��p�K��	��KM
��Wa��?�6�o@a���3����'c�����ǵ���T{{�����u=��0��a�ݟJg���ޥ��d���5T�AfI�lj�-M�΄[�lOD����V{�}�i��HP!��b*����L����Y����9{Kxv4�}���_����F��c7�߁4I��HM#���Z��p���-��;��]AuA��zu@��6 d�/@��e��L��ŋ㬐J��8ɏ����'��t;��hu-���R4�w�~f�6���>V2:@�cP"���,6��ĹI���LlI�ƹ<���!In-�[��啝�]�c*D=2�����+����h�p���]j�Ŵ6��э�����Ϟ`�u�2������ʂU�`��ͤ�Y�g(�ӃW��+���:���쯒��$L0a����>�,�����5���DwW;�3T��?��g���7�.�z�+B�{%P��
y��Վv�"������P����w0H$?'��g���i ����(~M%��}cB����T��>��s��aC�B��lt�C��c������5�gB�h�Z	(�ü�f�m4�����s[�����4�,�D&�҆���J,�n���\�� ��q}��6M��)L�%�h���nÒ7(�eQk�0���4�Z9jެYY�W��y�ti[G��T���D��A��Y��@��V�C�1<k2d��7��:��v�q���؟h��(�l�/���y5�ȇ6L��YS�S'�(����o�uLg��JHbj�C��=�y��釗l'W�e���Zh㹩�c�A.�QWC����(�^Z�7uޞ�-�$��a3�ވ��Mu(��p�����<n���+﴾��w�V���Z�4z�]8��7
�e,~�������P�<o���n��-�ԅp
F
1���5PWFB<��c/�����T�^c�;�C�meMaV�O�+��Z�7G�jx���n��}ASTՖ00g�?�NK�r���H
B.a�"�P``�1F�w$M11`��0u-���z���cj�ϖ���qG�Wq���k�}\��r��;�{���ԅ�Rg�0���h~eM���~/aȣ!�`��6�`�^\Ք�^��m̄z���T�A���Q��~��dZ;�+X�(�8��Cy~�4� {R!-� ��Ifb|^60��T.���MiVHZq��z���M��3�i[��k#�l���Z���|�����#> cu����t|]�K<�ge��S��H���-�F�����D��,g��Yz�h�k閴���kykUx��L])��U�����/-t��Ք�:��wX]�m�U�<���g�b�+��#L`A.���.s��%i��APl�_x�L��&7�ñ4��%�3ZdׁA��*M)h�1��Fg�X9���B����@l=K�7��Ņ.�q`>��_�w�~��!���&I-65e�u�[��Fw FH|��Sd���т�#�
�yD֚�%҅��Ig��h�����y\=w����n�3��*���|�3�����)�S�T1�{guW�����Qy0A�ugj�a��8���<C
����	��ٙR0���Vqr�%�Iޖ��ju����7e��� �_���R~8�)��m�i8��&�H	�Fn�@}�n�t���Nڂ)Q��Ɛ�.��Y��'��-�px��!���u�P�L3	6�=�Hr9}�A��_���� �)>���gst�����|G�1�;��� �I6!̆�ܐ����?���L�����<>�����[�݁�"`�� ��`4#�)�拮�P	Ҋ>�Z���T�S�h���[u��b����
�h��ȌGQ�/`�mb�ҋϺ�pM@��F����EH�[�R����y�|@Ē����	�(&�VԺ1ůxey�*i^����u���P�8X��+�vӺ�/��J��2�1���v�X��Xa(J�L�
<��EJ7d'Ʌkf�!ػ�y����}�M�f��Қ��g�9���Y���W�	
9m�J@�AS,�AA�8Ao�`�޺l=�o��:	�X"80C��)N8EP�?��>�c��A��\�?>�d�!���6棨ݺ2��:��2��X�5��fA�iI�e5[���d5������R���6�P��=/5şpBh=13x��k��`�c��Ɛ�T���o�cdU�����>�s�������n`a�kU���5����	�����W���d��AKf셺��$5�rKR�Y�d�w-ji�E�\Dx�gXm��$^w=���nD%�� ��}J�ɏ��rIL�w-�+d���l<8������ b��Uf_��mH������m���i���ǐ���y�;Bxƅ���wj��$��N@�r§�3�8+�^����f�RJI=�6�㑴Q��r����F$�K�X\�0p���*�`�.��&y�e�:���F-_�v�9R��]�[ 	�&��6)dP��#��������dU2��x@�����KB[�p��$A�֒���	w��|�G@�$i$�k@0�s��{�خ��T;��|5"~��=D�V�>��B�-�`��_�b�qM�`���]B7�f>����O��C' ̄<�erK�S�n�}������ޜV^�����^>Vu��U��-M��@�>�<�9n֔�#8ysr�O���y��dhm9e{]��:\wN��ӁJ����e슾N���w,ܝ瑟��QL���*�,���eR�BoĞa�
I��š�K�O�o��-���;�b�����6@�,�SbZ|�t�����9iАEQe�4`i����-�K[���p� J��]��	#{+B+��#�e���[=��F=�� =k�O�R��Z����Tn�x�^���f�䷪�6>C׈�U�`�;���҆�D�zB0��k�vp�wwJ�\ߞ^���}��5ݘ�N}X�v��d��s<�/@gs��4��Q�PF�Ps_A���!�����<�yc�_5u��=6�P�C@C5�-�TT�~�k�����B�*7��E�G�U(TR>�8�.S6�h}6�lé��iY�2�8HDb|�I��!��m���$`�C��J��Z����&��O��)�ٴ��V��=6@�^��WX��/ng1�D���mг�HAfB�e�@��ܡ�@'�v�fw��ͥ��V9��~|��{µ�Տ���Oa������Ա��	���n��ĺO��'�G�K��,�D^�:��ءs#�3�!#���7�} �6��C��;l������آ��S�C}��{	p�.\ 7ŚP�r�(���hصg��br�V�/��
��7 )@C�$�&�)|I|�y)l��L^�l7Ʀ�CُK�*�:۶�D��=OB(p��5��@�KV�ˉAK�]"v@ �
���r�C���_�$$�\���0���Y�z)��X���T4�"!B�.�Ut��&�'���Ln����t;f�.��s`+;�K�ɓ!�c�t�l2�"yD�M��?�	�2O�#�k�b�<+�bѪ�ݢ��W6�����`�Q�0��6���S����a���������Qlyn9���{գ/(�5.�n}����]TH5P"�ӿfK06z�h����A�n��U�:7�N��1��9����憐/��O"4n~Z���ΐ��Mʍ�������`��p]v�N#�<�t�l�9�`4@�����ef�xp�����VbcN|����G�O�[b���5o����ң�{e0�#?kH���W�
/=��q�;v��2��\�_{<�2�u�8m-��8��IdI��G\�b��#ךYrvA�zi���i�����<Ц�#7��oz�]⺃�]�2V����ԁ`�S=횡�����O�@I��7��w���0���}!y��.^W��$2'���i �#O�$�3�� �˰�n��.���g<c�������.�,�Z   D�K�,7�x���`Aq�M�&�D'A�W����m~����^e�-^7"\\�\��#�I69�����U
�y��o�F.�3-��cac���'V@dlƲ��%���[\�;��Q0��̨��&�M�p<bvz�_��U����m����t��=�����n����Np
��).k4Γ�� ���2���15s���
F��-Z�-#,�����k�qd�l$�l�d����N*��|�C����/"�B"�������L��̩���M�:,��-�q�$'��+C�����m�l�Xf�ӓ���G�@0�q1qЃ��;�-�QT�
�^:]X��@jw ��O`�Շ����v�Y�,��mL(� 0a^!Y�|���Q��j�����i`9������X� ��|��yq�c��$�ə�'�~|��1��� ' ?�UI9�K�_�M��`I֫�~�I}��<�gYV�z�O�] �4��M�Y�-��<��|��y8�ނ\z�\�������-��y�Ʈ%DrSa����=,�x1�:g>����SV�ָ߳��(sݍ(�~�\ �4X+�}�ٳ��3�ό})�e):ߑ{�['Qi�`�߯~ى1/�̲q<�#�۬��<��ʀ�jq���H�o2�r=���ш%�e섆�B�Nivh�`G�wS�nH��������RA�T��h�!��^��M�6���<d6k.�x7)j�u���1����%\�穽3���_��`RsaB��J���9��xX+��@�q�������62U�R��:;1�C��K��fPv� 4T�t��O�|������˞�q�5�+�R����3����^7S,A2��
��pQ,��/���/��*��nW�����9Ad���]��$*,���Yb=��t�
�����[�N��U)��z'�Q�;Ӆ)�@�O�!DHh�OEX�W9&oE�f)�]�34�O�zzK�Vݖs����^�U�-���zѠ�WC;t��['��h���E�Mfͭ��f㓫��-����kl�r��,#H��@(C2�(ǞT\Isa '�8ty��L�������x�DR��� ��ߵM9�����6�ʔ۹��3��TE�q)�������h��PVl�������P�vJ���7>g���HU�2s���`��y�<�2�b6�j>�:d�г�����-݆��O�(�5��Y��G�b�q������v>�I��_,�*vuF�>��
)�/�_��
G�w�g ;&�%!���=���l 4Ѱp3�}Cې3��3&ߜ�z
��?&�!A9��E0� ��g�C~}aac�y��ř��0�ò�n��v_����[�p�#j�'Y��g������rl.N��҂*O�Y�ȏ��XaMr������5�~�KW��{˭0Z�Ar�o��,h�k�1E�Tr�C杈~"�����BKrn�����^m��[��{2j}XgB��7��r2j
66ڄy�j�XbkH����ưR;:�W{�bw��ن6���Ht�����7�y�3�?ͮ�P�`�k0� ����n�BgH��-"�����_2�����ǖ�H�%���e%���VY��#E����V�YKN<x��Q��=�2�cS�tP`��!P��\(��JUSJ�2�^=��)��C����x�:^{��޳��9�m�2DlJ��Ł;����O?��\dn�-��"�����ྼw�2'~ZQ�����Za�<c�_���>̴��'�h4��e갛�{9�M5+>W:�7�T�g����f����x�����y�V� �-��f��N�E���E��+ҭ}��Fsg��$�y߬q��q��2j��*H�(z�A<��h+G�Ï)MUh�A�k���Y�l��Zt��\���; N�X��p�_D�
�sN��E��)�6���sf.٧�Y��}�����O�87�P��db*�%:��ܘz��~hP�����j�i�m�(���|�orb�ᏻچ=� {�n��=~��@��&n��Y�/7U����t���I�7�
\.	�w��B�H�