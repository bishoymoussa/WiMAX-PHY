��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$Rx�y�<��wA�*;�x���@�̦�W�X�fa�M-$u����n~�%���P�$��W��kYَ���P7�?UMfT��q�6�U��k�>����~�\N�(�����X�e���/6U|)�X2pF�]$h���d.���9E�	�IN�f"�\��e�z�y�b�����Oo2�?�qˁ'�͜k-�K�P|����y:����3�l�d���bl��ˢ_�d���kx�rq�mh�MذM�`aS�.�DW�mS�9���Y��+�>��!��!�T�uOB���,��\L�7m�O��W���6����'���j)n_�I����2:��$�K�2�Sʫ��l ��!���{�l����.�j4�	��很�̢=�����N��s���s5���_�R�>����ТP .W;������	�"�מԫ�����]�#7@O+?�⡾�Ԫ���e�O�\A�	�ͼ���ƹ�d�	@�nQ˰��E؁Bf���|D_�%au�-�'���w�*%��"AM$w�*���S����EV���+S��'���93��ح�;` �a��Y�����_���f+��AJ2�sz�}mJ����
H��� UYVy*�V��d=�[���� f�B����_���a��6��#����%VwW3�t��:�o�\$(^�E"�~�b$F��N�@,I:M����e=� G��X?/0:6F �b�nm�-\z�13�cx+X	;�?�LJ��n��iWk�:���r���~+�v�,\�
v��߁D�!�^��
9�8�V�G�.,Nu�.j���wپ������vy��}'qhU�l�h3i4� ���xmf�UԂ���ӳI��������G �A�/j�����q�p�����]HJ8�/�e��ǧ���L��bE��9'7�+sz����E�8)�2o_-���S��{Wq���g����U6���c�<�{�����%�0��5i1D^ř�5��;�����+�M�7�`Kq�׻��U�M���* �R���0��i*��/�k�2A���,J��-�X���1�<S7��?3��X���pT4˶���0�^ޞ�/2`|�\W��uD��3li���6S��i�����g�{�qvE*}�51��F�va��O�ײ��Y�	���XC�(�/�t�	*EUz&�����7�,Q攀+��WD]q��>���uC-ŉv��-�����3|T�$�.�>�" 	A�� �J�9Ï�<2дh�[�J:f^�Ÿl��L��y]k��Z_eʹd�P��}{��$ӹ���L?L!�|A�Ӊ��Y}ZQ25�����h���o�)�|N�y�%+?lb5��wP�x�P�V �"�S0���4ù��6����n.)u}�)�R��v���~�7��je��@2�\���V(je@�Gê�	[��q����n*�������<[GZpk9D��-Tݎ�>r�X� DX � �m�H�� ��L(F�BT�KHr�si/cb�3�1�_)�zAY�o`��?�!X���7OJz��Σ\J��$$��Ṟ��>ث��JW��b��(<j	��|��
�u���/��4ʛՈ�6�vd�!3.�6%ˏ`qU$���w���|B�t��Uj�8%��GK�߳2B�9GE��Nݨ������&�B��]c�:�˷��O��Ř'����]� 8v)�?e4G���ԋ�	.��gRqOɛ_l^��4(�.�x/�P�2���"C�]b�_LO����!�p�'�W���֤�R���M؏?񎙮˹	(���,^�O-Vh��1���Lf��ф���3GΘ���� ӯ'�P0�lD��8�@'ɀ�e�+&�A@��o��le�SB�נ3O��$�qh�#��x���K�WO�����sm4�N�����i�&��������G�a'4J���C~�Fw��x"p@:��%b-_A�Y�ա����24ȧ+�(/��
,���U�O��r:9�C�6���aLG�\u��6��f�j��Y�/�FP��RzC��I����dQO��?�2y�Y��/U �xF���t#�D3,ˑ��[�%6 ���yKg�h�x���y|F-���3�U�H��ٙ��j��x?��p�$��,Ŀc8UT����L�b��­�$	���)���<z٤{d l߽`�	�{���?#�5���֛��Ǘ�q�p0S��Վ�\w38���[7S��o���g�#�R��(V����ڱ��rM�I�\�TΑ�0$��-�##�w�A-���KY�I�;-�Cf�������߀�	RFiw�|-�]B���d���L�������E4�V[*Mv֤QK�xW�Tn�c��.$�L⩾�=���yq�3���=:��v
9Z�(X���
�laY-ۊ6۽���jx�QgӠ���������kY������Xh��4Wbi�1m����dA��}��|,�t��FM�a+V�(�P�(�(����ݏ�UuV���� �vMF<������L�C�,!単��J�$Q�s��\W �;)C[=n�t���zz����isp�Y�S�ۚ.W���C�p�\���%�n;4���eu̰���Z�^�}K������M$W#��L�j�Mr ��
����e�ev�� '�O�i�C6A�v��1ou��|<M�'�`׷�I����Y�r�ݲ�'����|G�@�EM^O��fǊ5 ����g�\����X] ���\I$�H �M��͡�CJ{1�	�	%'"��#�f�d�}2y��`��UvA1�iɕ�p�� >�4�XKCl
�4�P'�J~���J�hy?�TiTTPe�(>��?�n�[O�s��Hʲ�3���C
Y���5/׵[�e8��P�� %�Z���a���,�qc]�S�}�Z(������ds�|��8x�Ո)8���5�2�SX"��|?��	`!�:�ẙnlꁬ[�K����'������il��LO��4��u@ ���#�D����K�ʌ"����as�u����י�L����35=Q�ܒ~�Z�
� ?�q��t����9��,���aߧ �of��}�٬4�ܴ˨�	7���9��Y�ut:h��%�:qò�r�*��z�Jʔۗ�;2vؑ��x�����=:|�V[���vQ�:�%h�4�Z���R�/ۤaf��W$n�����+㏯dQ��!#),�Y���F���*K���`q�&S�����U6��g�NY�lr��%��\h��$�bY2\�dnk�Z^���F[��?�w�)	h�B qb�wV�o�K�,)�6&�6�Տ��}E15� &bř�&�%\V Zl�0İ�fI�ͳ�K~JBt<�[s^�ߓFc��#`ЬN�f�B��,,�]�5��(��\l���C1�vH8P$M�e��������Ǒ����.�b�#&bc>S>��W�Ih�?�Z+eJ��P1��ūR��4avg�oڪ��=F���½ЧI�(����H� ��Y�S4o�l�#�o��9�0y[�H�J(6��,B�y�ƼB%f:d��8bF��
��Δ��0|�HG곪X= 3���O���"��eV��K�Q8�����sL1�I�]Ղ��N�addcZ�qp$)	'�V�Dhˁ��z��N�0���`�y㐉w10<����aI��i�N��A��zN�:�Y�����r��G2qE���d�8F�	sl�*"��X����1����v�Q/xmY��a�M�G��;x�Jp8IJu��l�Qg�$_c�x挀��֚�P!�W��'��:Go����ҹ�f�U����vP2A�ݹ��e�k�ԝx4xƥ(�J ��Z2̐��*L���׃��<4N`�\E&�[�fC�}�ډ;��g���I
�wK@�W��u��/�2^�A�	��trd��,` C<O���w��D��d��g���u��kB��'���	Cl��O�U�ۭ��7�p� <�W��ǚ��c����&� r�_5��c�����D{�ɮ4�b�U�o~3��&b�p�6���e��Un΋$�ؼ�/��)�aasI�m�+{�y,C�?�)5X�e�2�:Y�Pa�-�.@P�Uy�}�� �$�jC��<Gc�?X�}�/�ΝDݭh����G�#�o#j�����dy�VL�
\��pAQ*����r��`��1����4�3u����ڤ�=���^�
RD�6�)���l���&ˮە.Z)�H?P��q�U���3�c5��4�����D��/Х�*dtP_��__�#��N�v��z�wk�:�
&�$ ��s²��]Ҷr�B��o|�e+%�}�$�Z�=ܐ�Y��
|�C���8:$�;��3�]�~ �����֫�LJբ<���O|��ms���aE7g�|i�-׋��r�m$@�At���63�����g�P��X��P��0}з�S��̂(�^�-�+��>������J�{�_����t/{���L��Oʡ���u�"��d��6�w&x<_�X"+
-��s��BfJ���v5�����K
�z��VY���mp��1� ��K�y�b!L]�VQ�3h�!e�D�L��:�Qv2�����:�1�?�Ũ�43Yj�Z/i��Y=Z�F$� �oсZ8J&_�9Nx������lG$an�_X��/�2N���GŸ�'"7r�-7��`=,�+1ّ�Bq�UPRw�7���]s9�U�̀2�&��*
�E'��y�����Sb7��l7�FP��*`:6~��Z�?��˒�	J<�r)����4r�{,��c�2:[���_�Xϯ�?�A�8����SOK��J�>��.cԲԤ���\���ܕ�."Ȳ��:��%
����E��{�"%��S�E��B�9;��ǽ�]���f��8vd����~M��<�\'m�Dy�	7AB��Q���9�NQ�}u)8:��|K������h.\�5o�^�X����75��F}+޵:�=�.�CT�p8���箺�i5ybBI��U�)+!3���\�ib�K*�b�~�􏁷L#�+�k�-�1G��M2����Ư,p�0�9�5��PeJ����j�J�J��U�%�ZV9��D[��Fx,׬�����;�J��}�?M�[z�~����2h��x��<N�I��D��mp��"��Hv���Ǳ�BEjS�*
`�_�6Av�S�(���d�	o�%����C�{���C�5��m�Z����t���|֝G�Y��(vN
��j�:��G��1����\��L�����Z��z��:����Dࡴ�hJ��]T�&��������AL�����'Z�l�O%�����D�[��%2���N���S1pc�]�&��6S4�%'��.�ld����P�t�y��X�eI��.��A	.9{*p�N�r ������f��>ğ�<���9��{��������ԴB77�Ƞo��; ��5иp�Nv�meo9Z�+y��? �]�DLG����+
��f9/�� �S�ʽ�22�lO�����=�0Zݤj��]��h��Y�l��rTٛ���x{p��{Ϧ�KH����������	}��v��n	
x��Z��wE���~J�cd�b�]m����	Pe�[�+�o��õ	�RrSU:�ti['�Il��L�'
���=cs"���e��Ҽ�RS�|��Y��k%"��:�O�fl��2y���G�1L`{�ez4�NM��Ni��%�3��S�9�R�a�2���cRo4��Z߽�ˍ�U ��~�gMsw}w�o��^G)J��W�d��\�'X��|s��ƽm�^"S�r�ϤN�%��kL����[�UQ����p��[x8�:ֺ�l?`x�J5M����9ȑ�RKn�&�}pu`�e�>��i��B����#2έ
]���e��0F]Y�fi�,�	�U�1u���>=��G U6�*'l#�N�.�8h����U�٘Q��X�:���{���χX]����1�Y�H��Ǳ�ڍ �W�OSW��UPW$=ۺ�+�kD:���20Od|O�	n��dL���?Ab�i�(R� ?�^z���"��$��"�A�`+���P��jX�SR�>&�O�%�q�����C��-2�g<�Y ��r��r�Jʴ��:��2~�@R�����U�~���'0��Z��h474�e3�O'��W�$�v�y�zY~���E��~�~�㾼�Ç��lS��DN~���4�D����Ϳ�1���|P��� P$��&�=���B�Dȅ"[��ƈN�T�r�mƗ7�ξ���A�;���`B\ft��"J<Ŧ���g�`�W0N�	a�h'B	��Bi��W�%v��RV�;������7��'����{x��"���y��Ŷh ���� ��)S��'��H����^�%Oi��B����J�$�avMt8X�<�{��YL���Afm�CuG�D��U>(��Kf�H�������'_�����b���o���W�89�̸�����~�p�#�I얻��l�M����8���D�S�j���1�:6�Zpk��yG�
�o�,g�7��o���7�q�}+́�fb��bߘ�=>0Y�k?����dd�_�� �lS|��	5��0�IY�����3�iU���:(�A	 �����	e����~@�]�Z�����Yl%N�	�����o��_"��U߄�b��_�J.���#�xlo��w��N��%(�>v�z�b-T_���_.P�AA�f��^� 0�%���2��2�����8ݴ<�*E@30��[:������]u�ĸc�w�'xU;��_'�q���5+���gm���Z�G<����a��V��S����0N�M$>=��k������$���3r��I�ǭ��� ॣ�l���[����0��;?����R�u�#��	=O�;�!��iP��%
��:>q�r(o}|�P�]QM�c�G}�)C��8ż��J4���v��B��g�I3G�����џ������$l��`G4�@�����Q�:�'��$[���o��R�m�]ӿ�4H��Y���A�����q�"4�Cq��"��C5[��؃R&���Q��m���r�aO�:;����N�9e�?p!m��fv�tҔ�kx���7�n��Mi���u��K�3"*��/�f�:=���sY��K��r���a;��7�F���J��cS�hFғg	�r����ұWg�CP!Nz?���P��c�#<��*�o�d���T=©=t�Y����t-����H�{�ȥ�����.~�kXY	-��)B@��'�#~�C)t���&q �����uF��D�!^�IC�u��Ԭ��FĈ/T|ߧL	l�|Ռ. -l��h1^p6��5Ӓ�V�������K�c�!�&$������L����l�x2���O�ڕq�2�.#˿��{�QZK�NȆ�s�,����KV���� [�~]RZ,��Q�9�ѷq�� kh��a�A�% ��[�3d���$ؠ�N�w�|}��S� �U4��n!Y%��ၫu��	#K{+�A����y=�V^)�ڔ���F���x.�V��kΖ<�Ǿ�q�G�tk%v��S�g�݇9M�<�g~��<{�^�6`	
��GF|��c���1jr2 %�ҕ�M$�ͳ��P����"1S���Sw��j�#����s�H�Ӂ�tD.�=Ͻ*��iǔ=V��q ��/��r�a�a�^��cO-����c��HD��녣vV�O�e�q�!MM��}l����%��W'��EPσ�w�ۅ���H�[�m��T�a���0M ��Nv�i�D�ɍ�1�K���|K=�6�锇�	ۅpغ-"p�ׅ�]$1����:^^�B;n*2�P˖EoW��XZJ����n2��i�Ö�����@�� Be<���Ch_������G�!x�I��G�U��o��?|�?�u��ͱ��T*0�BH4ON3'�|�?�_Fd��+pA�����e2�����r�j$�U!� �����"fhb�
�f*���lW���fg�q̠5�_&�>M�]X:�s�1E�����}�Ѓ�E��T9�!\��rg��;�h?j!U��*�u:�DMy���봜7�;�L�P>��d�G��H������F	߷ٙF`	"H%�z��`\�@[��SlI����A�^4܋��Z�Ȏ�oO�J+�q+mټJ��^nի��B���`�{�P��CX:�/��l�ԱMʛof�ԋO?!������u?��N&5�W֪�-[S�<�u�)e���9+�Eb&,+�b���(�0x6D������Y���mJ���Kʿe���H�Wc�����!�e�vx�fۋ��37�[g?y�k�/63��% *&]Ŋ'�=�{�CUsi'Ϛ	-d$Il
 ���I�<cr�^=pt<��D6�6�ݠ��v��p�p�����\� �27��$tI��Xl�!
�*�\r��
�J�Ҵ�x�h��[F^�$j�j�u�z��z�[wJrkp�!i�;-|�0��$��'8�O Jm��*����<��sq3�LiΊ���ѰDͿ��y5�Ѩt]MSյc�Uࣻ�����iE��:�Ŵj��e<��EK���o�cF��i0{�徏�:�w0y�+�Z�8E��޷!)�L�[���V@fF^G�WK���]i*�Kvt`7h�BA3R��f��Zhs`���G/��D嵙�.�S������f��I;�w)Z��xM��?����^$N	 ����!��
�L���R�깵������-Ё6���<�W������,W�^VQv�#�ө�G�ڗ=��/ٮ��g}�l��4V�V&�ɩfM3�]Ri��c5����Z�����v�[�w��a�k.�7�H
̈��g��]d�y�O�H�6����{���[&�@J"��4[2�_�}c�`��Sn�W��W���T����xu����o���@���=����
�Q�������!����kfQ����@�^_���wͨrxa�	
�7�9Ig@�ԉT$��Ǘ�͘��RM�F��(���v��np�;��Q�Y�����D'��n2��nP��pƦ��_�7cv��W!��A
���ͳ�	V��(v���*K��+R�C�!��JM�}�0�J�R �8������D�\b�r�tʥ�<BiـLI�FZ�_���v�o�X�4��C�rѬ+��0�*������~�Z��x�[�H�E(��I�D���T�;�����[��'����(����\�Zz�^�}�p׆S�Oڿ��T˦���޿%���tNj3B���q��Gڤ�UE�|5wHl���Ȗ�`�T�C�_g���[��Tr�C����~�6o���-�a՞X�#�uzf
6���C�+"�E��NO�p7gCH��� 
���Ş"�sN�|y��P����,�<�\g��.�q7)�O���$�R�N�9� ֻ5Qu�����\}e�pV�^�Y�	|J3hB�!���3�t=���js�	��J��HK�9�L�-�3_8���p�õ�$N����ߙ�xѤ���b5,�"Bz�B��	�,BU-�W-�m~�"d�:�$+j# S w�W}U��--YҜb���إ���<?��j?ȥa��Ab��L����G�o����'D_��eͻv6����`�Oj*�0�|��0��8��2��%��΢p��DԴ�{:w	 ����`y�A�
���q+�;80�7�`o�������'
I2Q��?	�"��䒠����9O����¨����$t����9f����Z<�B����cK.pbk������_~�d����"�_Q�q]~K���G��o��sI�@�V�"��K�;?z��`S�W�L��{��++*Ќ,r�	���Kn�t��Q6�E� �� (��i��{Z��+��&�����=�"{L��R
��N/��S�< ���f�"؇�2y̲_���|�x*��� ��&'Aø6�o���%dg0�����ZM�A<lF� �]������\.A���ŧi���9/x�i�M�h�h"o��'�#~{��-�R�v��@Q�-�Ew;�b(l��O�b
�����u����tkEFu !d����w8_ �'�@ ���]6�O��=���0[�![ ����;��J�=���ѧ�룑�}��ޔp|x�n.���eD�O.8i�C;A)�gB��[��X$ ����}��Tq�p�WqZ�)nG��A����ԁ���O�.炜��wh���m\Tn�W����9Lo�R:�����y�'��S1m�׸�!9�b<��_$wb�WMY[�&�6���&M_�r� ��w"�4o�j�2ڕ���s5U�&-�!�;�����U~u���+�QSۯ��@bt�k��n�-��نԗz�_o�^h��A ~x�d�7��Y��)O9"!�͐&���������L�ߝI/��l���H��-3��ױ�^�eХTZ�St׶����m��1��A��6����a9{�d��^I=�8�?��p��l��ڵ����t�R2Lm���m�A��� �F����o�9�%1�.�ԯ2���g����6�
H�=�`�S�?9�}�^�,���ƃ��u��s���6Q5u�f	�
u�N�Z]�ӫx��;OuۉmF�e��F�oh���/`�N,���q���~�[��Q��F0\:�F���!��Lb��M<���iGZxE�����p�B��e�rX3�|ĉ����G�p>�+:��&��4����ː��zs�6!ߟ�K_���.�Hf=��`4��\-`�yL�E�I�謐�B��������I�22�6P�6az����B����R��6����Z2g�k�D/��E&����M��Xn�\���?��&|z��ظ�l1Dh�9�N)��eew����2�,��1y�d���2.[�QP�Q�����1CT��N�y��NLW{�W�h1�-]�lUh��VA̳��Mpz���'��r�4��Z`��]����,�,'�q�a�:G^��8~�2�{ *�ݻ����ӵ5��a��ېn	�Y�ídqne�"���/b���F���R�[��,|y���0����M���%�~��� ÷��x��i�N�?Л�����4��*�J����x����<�P	�/?����p�J����� �!��r�9�R^΄2U�������]��U���yX�)B�Z/�����Y����Gl>d^,{>�v�s6��%��,$UK����s!鵼S�nH͆3Ne�.;cU	{��{�x<m�>`,��*ԉ��uݨ�x�^fn�G$^����d�ُ͚V�_��!��,	1�城v�ǋIQ���ː��fS�30�r�iQG�?�t�5O���e&;6_�[P��1g��������,������g��:׳apR�eުr���_y���'	Q�i	<���e�q^��0�u��خ8�+��a���� =���ϑ� �N����aQ���?e���H#��6F�LT�938��y��8����><�P�\�Jo��X3Kp@RQ�,q�젴�����НL��R���Ŝ�-�+�n2& ����P���ܹ���)ֽ3[�/�H�닲���V�d,�myh�D3C�\`��j�kÇ���c����`K�s���^1*¾s�S��UQ&�����o�����A��*lRD_�0p�I"�vRO��#�o���]k��O`1s�4���l���͖Va�Uh�L~�0(r��J�#{�b����}$�W�Y^`�)'F]<#�	��.\�5	�TqPt:|Z$6?Ռ����(��ܥq@l�B�_�yB2{���=�I?����u�.��*<��g	l+U|m�f�Z@�������n�^a�i��֗�t�ƥ`���/�+�T�?kvJ��%�8�,*;[�#��J�YL@ꄷ�Q.����T���i�+a�Ʀ�Qԫ�f6��h\a{�rWcI�yQ�Iʥ�d5�a�(	k�M�p#U��Ų���TC:_1��g;��C��"F)k[��A ]�ĩ%����6�+_��.���7ƔofD y_�~�k7"�s ��>�s9�4� �I�E�Ń�I6$��`٠l�/��?߿�5�R�Sc�C:�1
�q��Y������~���}���P[���h2�Sڻ[�Q���Q�=��ɍc�J���wS9�$�����iz&��H��f�X�qD��ү��A!��#A�=���E��T;1��#���7��(���s�	I ��p����YMؕ��pJ��i���g�k��������N]ƪ��'/)�'ǻG��ZL�.ٹ�U�����v�..�:��Ջ$\]:�CZ/S�oGo�[��~�ċ8�T+Y�P�����a�{B ��ק �^�@,hOa�� �gћ��c�3B��v��l@��;SS?k7��#��(|F��W �7��]NXP�It�S�d�R�1.n}	�0�$R<=�-�g��&&
�Wc036�xC�����t�(�/��x>�K��A��R��yhzx�7`�X����j1���ا�ao���+s�܄���\e��]S��� ��M����HX�@c�������PSti����}.M:�͞��W���ۜ9���Z�{?��U��NU*sUp�8�%���Tk��k����Ŕ�����B���ͅ�Li��-��rzK=�iLJe�y�@�o����<�F�XJ������V:�l<12O�|?����;X��;^F5[ ��l�Nl�i��W�~�����o��4z[V:w���^Z����)Yj�Q%���%��|	��D�V�h���2�U��Ƕ�������lҐ�*��u��N��O�#�4�lG�<P$�*��Ԫ��{���P��h��"!0�ϧ�@��nS!��V&�<��wO���c��Ћ��k^�A��}_n�_G��aW��&W�Wp�x����D?���q��)0�EZ���R�f�T�E��РƆ�q�����Z�/�L��c]C������'�-�S���B��U/,9%�)��Uj-E�H7�nF:[�<�y�[��P0�+����3o��K� ���ƥ��uV;C��nQ���?�������̵0kH���ע/Q�b����І�[Փ�rE�\�d���Y��e'�Af��#�#�"�i]�9~��ڋR�M�)˥�Q�[x�$�@@��x
�y�h��]C^��$���<���:枤��	:�1�
+j+ �ê��I%�Ul�t����Q�Ď���y�D�z����%�&��J��-.�O��<~�x4�
�$X'E[�)�� f���������v�a���;E$S�a���K�	��Oa�0����pj��Ob�9. h��n�f�>��+�@�U��1�������v��~I���e�4?�����o��Ǉj�%��Dm)��"k����m��L$��̥��E��kk?�)�7��H�M�af�,�0W
`������p��<�FMhG��T�-q�Z��-ބ�i��z�����0I�5�$���#��4��7��',��`b�B/d����ο��{�^3н�(� Yܮ  ���p�weZ��NV�N.�fdt�t�����q�-~�kd�][�
@[��^��j��T��U�2q��Q��zv$oӷ�N'nFI ��
��0\4�b۱.��Q���1k�d��b�Ӌ�:*��^ZN.m�=:ɒL��v�����V������
���N����,-�Y���!��c��y���ζݷ#�b!�"x�~��yd)�� �sQ���7�3P��<�DoE�(�ʋ�̌��Ky��0�:bZ�G�%Qϔ���9o(�4'��Cd�+%I`��o��Z9�Θ��Y�fL^=O���sw�3�;P� �~�k���u��>%�K�
�AX�ͺ�X�_K�}����&9aW�%4K�n�yWD+f�ӷ��Uܧ �,��2%�S�f���6��&�B�Djމ�Ã�O�Mh�6�	fĜ*��<���,��W�������� E�Y���;���h҄>1��x�.L)&�����k6
��Sӓ�7(�S@���	��\�\��/��f���:!Y#�P�K�g�H I�9l�t����kE;G�9:Ǡzr���4�ײ���Y��^a��x����.�E�DB���n�`C*��SL�q�0X����+!���C-�L׃f�S6?|�P�u\%f(U�ُ�/U�B���#lq���d4շ�p�����msHR��"��C��u��!"^Yj��.w)8�[B└R~�l�(]z��ӑ��+zݚ�(&���5�}�����c�9�*���������j�׀)B8W��f����( a7ȫr����j��As���K�;��B3;�M�{�*f�R��z�3s����n�Wr
ҙ���N��7�R����E����1?�aYF�'c���0��lUj)��݊?=�.�� ���-�"^ZÈ��6P�5�\/��A�\��g�ޔ'SMG�,����Z`H�QPM�Sh܌� B��N�r��D��]{�G�^�ך�ŝ�I��o7A�I����gFpM6V�a�oPzh����M�ؾ_N�R˯8�q��Mr#
|fq8�N�Ɨ�v:t��TQ}��~J�Sc�V�w�z�2���p�pS�0�ߣ[h��{fA\��'l��
��d�]�:�{M���	���$�V1=��g��Z�T�7:	m�h<(7�rp�"?�M]�����a���]��� H���4���gn�x���컶J�#ûܣj�4�n4_��x���]/��9�<��j|=���Ƥ��K/�=G��׃�Ϻ��$>��V�p��gV��eڀ�-��h��'�uU����G�*24�糟6������_�0�S�4�h�N�k.��k�sv���&�TZ")0ꕠ��О��g�g�ڵϬ>T�JRm�GƁF�X��D�����V�3�ķ��E0��'A�����o��h0���ݙ���/�T���%���x�VI��@��5;�����]>Ŝa�k�
��D����;�v�R�h� ��d@d�\�����!��^���
����2��h��Ę�l�}U��?g��8?��=��X���@+r7�1��!ث�	N�? k�Kgu�����Ó����R����ǣ����'6�O�/C�E�򘣧OQ	�1����X^+S%� �u7��jL� jw��g^&�y�@�:�� 8K�\�Q��z�,��i!�xF>����ɾ۞����"ûQ��vG��\�V�`���G��O��>�uؒ�������t?�Ts~�Nz�-�ӽ���,����5��K玜�[ϕw�"�@�wU��{	se�ET�@]ocQj�W�EV�9����L��V�����z��>�f�?TN�l��;���v+π��]�z`Q��9���9]GG�dӪBS�+ﺵu`�N8cֱ��q�� W���]o��T��~&pY\��3PH�A`SkR��q.]�f�{�۔0�_�Y��N���5�+/&re	Z�+J�z�.�?�t�ߝ.�f1*׻�T7�c���������[2ƞ��0*9�B�/W��v��|�X��W�zݦ�Y�VZx�0�_�!�,��wZ������wU������E�@�rDZ��7����c%�ı�����͑��&���:��.�v���=
[Z�L�EǴ�[�uHQ�L��H� AE|��Ax\�6��	P�S�be��̯}�OK�Gqs�9�ȞZ���u�����l��Dq��)俎ݠ���E4�+��p[:0O�Q��#��ڝP�6����~�����C�a�2Q�����Uͧ���t4�	�E
�i��3۝�l���͔�g���>��
$�룤�aO8VVrC푳(������������c�"F>�+�nC�%�.ϛV2�D�mp8�o�d�ĝzDq�&&��>���0�\���0���=�{�~Sd��G���}��F�<[�JY����N�D<�����&VtX�Hđt:|���tODO�Jh�h�b&�raxS�����I�k� �Wh?�z������_v+F$c� A��zo(���Y#r����xȞH��LsM�4X��W�o�N����O��POB`�W�z�.x����|���dzC��4�}�bۼ|AnS_Uky8�*�N�y	W��hC�JO�y�@E�E�SX/ⅿ��䲔/DL���0��LE*�CP�'eKf9�=�F(4��J�� _��J-���ssġ���ڿe�+����/_\���`�j�^�.w��'m��T9�.
*� �0��z�������u�����<����^������{X��G����<�fm �3D�#���X�k*E�s��~޻QP��{�P��(P�(!��>�)����-\��Z��27�ƨ,SJ� *3Q�K�8�j4�w��� ���ڝۧmޱ�O v�@�)51�N���\K��yj��s�%����3�WlN�/����f�M��Q�5�~���$����0��M�	�6�:%T�f�JSɪ�w�EJS資��M�+ ���2��E-q*,�܉i%-�>���A���Y�؂�u�߭��Q��i&��������\Oq�s�����N�U;��kp�������,T�㺃N~]��'L�`�l1��I։$��W�Ĭϸzrm�k������wp.����(g|�R�/dH%R��
T$����0�����"����*���,���� OS�GE��� sYm+9��c�r�� ؟RG���U�!�����}S]�+�P�Oq�����F�;ԗ��sK�M�6#����8w�F k���y.�<�V������T|v)g����[d6�7�^Yax��W��?bz%E,���R#+*b6�4�`e�Y�Y�Wр!�z�����u7^�F�c��>X?G:<�O�!������:&����V���:*y�>�h^��ɣ PO�.�3����yqh����0Q�%��M��C>�r�ARܪ	��z�Kg�^�u ��)�'��"��HA*~�t�ظ|��j�"��y)6A�_�����nL����Q�G�<�;VY�|��XCRn�ՙg��+����Lu��?��+Y��_�� �?�ʼ�L=�T�J�ϯڅ�w���(��OMe��k�p"�w{ S��)��
�P��O	�����"z}3T|@��Uґ�ㄋc_�~@�n���e7�m�.N��^��^V�P�]��6׎m�;� 9�p0a���R����*J%��۳��>ƨ�|�8�d�R���c��Fp����;����P1�"��]���'���_�����x��)����R([�'s6��z��D9�`�?o-�On'���P�%�t f0	҆�O\ˣ��)����;β�Em�u7��ϵ�c.��<"�^79IꔸU�JA��G���F������n�����ƛ�{I[{8FTm�&_�{[�bT�d߇W�-�����S;V���w�V]K+�r�g� 4�!������$z����	�v�]��D��wX)���Gk{Q�݈݃��^��7�6st�� &� W�E1�B�G��dc���)�#@�뛍,5��	��!��"�Cg���SE�Ū�q�*,AgZ�d�v�Q�r�>4�����W,w�a/�R<�9�;��Զ�gl�V��m�}��	�4~#d;$Q(d����U�~Z��
����/������WEZ5?�����
p��=��#ƣ2�ڛ�t�2������ңу����4�A5���~V�ª�u�G�tcf����Jkj-��E
ͱۨk�������+�j�� Z9_���������sR?����u�#�ɜ7�g~lDt)���Y��|^��j���V����H��b�SS@� =��Zb~�_�W+ �G,f=H壁z_�by�fd��H�?Y�7�P��ck]��z�b�08^/�'�3�Y����;.ԏ�[��Y�T��}�L�6��:�Q1�FE�����+ކi�n	���T����Xr?;�~7�T�4��v�"�XEF.�2,&9�CC��dgkf'"X.�
FC��=M�����������.���!�\�<\�& �X5QO�������L"��C("�l*l�4#����?�`����@R�\��q�NKec��)�DZ:-Ŧ���y��B�S�p��HMq:��"�֊71���\U��8HJ����3����xWcJg���%�˕��_- D�q��{��-�-��`�7>Kz3�=ϙ+T\�����a���:�"^��
-X�2�4[!,�!+�bOɆ�s���L�|�L��8ĒvU?`;�w�L���&��A�b�$4�axN�<��-��)�d�ń�+:@���I���QҚp�iA�d�5� ���92�4����Cŷ�J�Ok������+@G��kY�BkW�N0����K�98���v�dl��A>��t�m����	���<K�Y>́%��?.+O���Y����E%6@WҪ1��5������H����z�Ø��ܵ}�i�ː���=��f)����t&�>�i�0!l^Y�,�XAܙ���#4P�i1��;�q�g�A�z��E��K�o?�{=5[d�~�Џ���T�� ���8(�~˴F&e?2��" `7��T�K)�
c/?�#=��/oTt�ǖIҵ��_��f2��¤"7��XÆ�̌WQb�C��ۣ��(�2x�`�o�M�q�(GL�����M>�&�Mo�cz�9�<2ٯ�H�A�� ��}~��g�U�K�uo�=J��������C���^�V�YZХT*�<��Թf�e9X^L=B6��W0�F�yaJRFA��B��v�Ög}W}aW�nZ�WS����	9ɋv&�c/�P�6���e�F���n��s�kݔj]��="n�	:m��2Uqm�缀�2t��P-����y0׭���e��[6*��7�{��8�:L�n��aFn��K
���Pe�k�:���?boef��q礻���9U���@}:$��E������������V���%�t���	Px
R$�n�~$j	'���px�Y��FV�k���2�վ��Ƅ�FH�1Ԇ��^��Llz��[���[���5fzS�)�O#�w&�δ�6�M5�C�>W�d�x6]��������Ozn�f
Z��{�5���!�=��@jgw�r��<�tgV����H����x�ӻ3֚���Z��3�(����,�dϵTB@p�Ԯt���
�����}�����h�b��"�:ףC�b���簅q���d�����6��r����e�g�M±+k�ͧ��$¯�Z/��`���\J��K�����Y��]kc`(�.4���1}A���LJӄ�E�dI��>�G[E,���GI*���qد�� l78c	ߠQ��Hr �X`��.],)Cő���&� �29�����Z�c&콣 ��1�����;�)��_������Yd��txI�����g�:n�~2�0:<�l-E�u]�#^����./����VE]��t��v��\>��5)��pZ�괺j14�j*�:�c�:����3y������\���q���2q��	5/dC,���<�}��,-�g�:�a�ȯQ��9��\�}eK/~$�H�7ł�/(И
Kn�d���ſ��/Q��5�xf�,���|a�C��v�͗>��JA���mR��Mn�ׄ�#D�y��
�x�k�l��v�3��WĦ��w�č���CB�84 ;�,#�������\�oGx#鄴��S�`�G	�hP��`t�k4!}8�9����ȉ߳��?F�4��XF�s����=���L��0���A{.��r���y�➝G�n�'}�}�S������r"~�x�l�m\�x�)r�#7�'�\�����>\�՘�(S3K��IY��n��UcJ�,"�[�V[�if�`��y�*�b[��
qp^����a�Cz��}wxćm�L�F�^	u�����g�`�������d!�f>�כ�"#�D���#�S�#]I���ߞΏW'WF��C�w��R�Y����K�����A�2�@#��#j�T�xn�hQ%�ƕ2�x�*����f�������G����=�Mປ�q[�v����r��ZS��[ �h�Z��1L����]�J5��)�ƴ��g����PJ�O�UnJ��)<�Ȕ�/Ͷ"KО�m6��Z�L}<�@m�K�ugA�p��:P���Go��<?5
�ɂʼN`��  :k�Ţ�LŻ
���S1���V-��	���T��DN� >`��_�P�)�S�/}�����?����6tRL�UK�SaWG��-6��h��i�64�����r�3�^�PMx��[4�H{|��Ɏ)s���W�ᕛ�߯�r�Df���X��[%;I�d\���m3�1=(x�q���="�|�E�N�=�:Q$C\�E�9���#=5Y�� 9�l�Jb�g����D��=*Տ� ��JMCY������kno�I�7�Rk}A��E�*y�Ϩ]����L�
&�W���-bL��p���ʽ�w 6�z�����
�GY�!�ně����G���(dE�W��}�@�R��aQ���4���oW��� 8�rpc�\����+�=���NY`��|n���o!U>.nH.b���t��3���&PV�ȭ�!#Qn�_Z�;R���	��Ŵ�uTpMk�!��/�I �$�thDB?���p�9Ж��S�)�d�gZ�q��Au�x{�����
@�Ko~������������܂�%Ƌ�|܏�Qы1;j<VCwL�%����_��p	�c٬/����H0F����l*h��;�XP-�0^��*�N��Sqy���0��x0��zz��ϴ���a��ktŞ|?|���hf��L�������ȵ'V����c��-ǚ��1�Y�ŏSV�]/������Z����)uu(Hh?a:�ٿ��Y�8��ܑ�4�2�pT�������\�L}{ҿ�?X���Kp�l��}����Kq�<��G�`#%�X'bEox��;�ױ���V�O�_�Df�W���3��C�m�!E��UO/��@}W7ϭFPaOF��3�2�0/C�
%�OӉn���1D0����Q$��W��S�4�Nݯj�>�"aU�K��Cp����,�cW�Z���l�0�\%����tS`��U)��4�D���l����%�n����W<.��K�_�è��(��+\�Z�΋�3b)�o�)~�%�a�c�@N;�\����z����-?{��o�/,07�̺o<!��@J�Zr��G)�Ud�D0>�Y�ҕ��G�}IV��~�E����x���.W�A�l��OѨν�cژ�x���S5���[^x�^>��$z� U���!}m��ϜB��i��>4Mr�|�^��D`ͣzݲ+�kE(��`C�rIT���=d`��cXx���A�K��K� <�㎤f�ޕ.j�^���Bȩ줺_�l�;�b���IRِ�n�.�y͡��n�2�����3XT>��q�.&��< J�FDP��~�H�r
��x2��s��s����ŉu�m[�e`�Ť44zX�4��c�3�}�إd���F� =�?�:G]I�k\Mx���K�=Ο?oz�ewq��g�9����]Cû�}̻g�x�����>��h8�/+��|Z\wvdS&���Su�J��8�tla=����V�O�%��ּ��=�j��4��xȊ�A��f*��g��,�X�qU�
U�dΓ�����L���c�̡8f_~�?{�7��j ���Q�F 5��<���rn�`8lG�N8�h~� v��L�������9��ZWYo�B�%��㈂��>YH�����X��%�:����P�Q���f�%��� �+N-�g��$�p�Y:�T�b���U����Q���hZP�X�z!w	%�dc��R�7=`̛-?�x��1S���aS2:�Z�{)�"a���[et�xdXiF�����n�y�&&B������D�m���#�dcx�ެ��[�-J,G%$s%��6y7�DY�fb|oUm���K.ld]T�n�Y^=W)/��`k��=��@�'��#���J�⮲(���j�xCc"�]M�?G�:{�P�N��[�7z������;X�߁ӥ(i���&j"��=��K���]L�(�Y��_��66L���(H�I�	G_54�P�4���:=v��	59��xe	�� �,���L�Ë��-�01��?WA�I��D
�}T�s+/�cPl��i[D�oR�Jf���6��(�H�g��q9.�Z����:aԁ��4 ��bM��s	����	ev�l�t<��e�L(	v��f'!"��,�}W�e�k�q��V5���vQ/�ux`�+Ox�gs�g����H��9��޹$t|A�O�x��F
�uR-��bI��7t�Y���u�ьuhP�U
���rL^�3�w�5!�׼~,���6�"�n?���P� Ocx��p��<wB3��,9aΆd�����҈/��|�$9R݆{�D��4
�������\�@8U��\r�}�`���0�j���G���;��4�>��$�ܓ���M+�L��U���g�o���3����մ����$8P�nD�;�Y��Lm��%9�6gX��Ʊ^�@<Z�W"$��Դ4�0�o9E�h���� &�ı�
��:;"h�G�C�G��!�ġG�1�j&a	���r���T~�7���@�P���hӥ8f���QR�o��2[Χ\V�*�*D2�(�����57oו[�b� �ҸQ�K0�R
)+5`.�8H��c�}�R6�QS�R�ō!�m�g���������2� �w���(�O*YX��<} ������Y"-uN�;)k%͖�i5~�2�!v�1����;y�.�o��ý� aFH��?�	����hL5l��E�E��e	�͉�ŷ���|G2yN���$Z��=�R*�/���}t�E��,( /�uxϧ���?x�D�'C�[>�8J�[�Ǻ�*�X����U��G�cGMl���l����]Уt��l,������1��,�l4(\g�ƾn���.�z2;���_"O�c?iסi�����-�8��hf�>�[���O/�D	���)J��+F�(|�uGZ�W�t��5����o��Ҕ��/�Jq+�H��{�����E��):���z���*��V4�=��LTPb��-�D%Ly���(?��ڧϭ�;����R�Ӿ���ߍJ���1Q_!vX����u�g	��铲~���gKǉ�i��N�N�z+�ys|F��K#j�y�$g)$��a�ؐ� ���V2�o@ۚIH[�g�Qx��Sζ�Ճ��T*	�o�a��W$�i1�����gv�Z���X����
j��q��k�*�w�\A�	�T���*����6K�"t�q�TgkFO��/ꥄ5���\���L�	6J.�}}�2L(Q[��`�'8G�����Z�SQ����'��㬐] �N~Q/f]�h�E�FW@��]I�fx�����g
�qXq��Ò���tg=�[����I׵>�AI��
f�	��碦L}"|n�t�Lk��5_Q"��	@o�9ڼ���cϔ!��(����B��o���{
:S��ɶi� ��g���'�ޗ� s�c'�C�"E��l���Y�``�
<�������]�d�+v��ͷf�=�qq�G�_'�U�5��zQD6��	�?���d��b��-aV
�̸�������Wzg��K84�뾝�#�=�t�i�'B+ގFM����s7@M�N%��z�E�w�>=� �k`�1���?��N��dhܪ��#dʖ��˺:\�X'o�,�91
���pz�tU������<P.��Iv)����5�����3nz�j|�(�A�h{�"�N�mؾЛm�8V�X�!6N	R������VWt���z�X�k��{hڽT�x\�}\�`A�Ӵ�)��[�*"�H�A4x��*�"��{8Y��q��������� ���͸�U��dr ��M�I8?�oVUp��V,���/�m⬥�־f�B�M�OP�G�x��\�]=��[z����k�c_;�@��V�,!���gJ�hQu���T���K6@)p)�8��Guߢ����~xc�F���F�?�iWC�cT@�����t��5Ǒܥ��$3�$[�2��L�X�_&а.��k|V�:�L��|��D�*�X���q����/(H�����,xAq���ʳ�G�VQ�K w�Q+���!B�}Бv�^��mWGkV�*?��JY�Kb��X�_ĵx��$�Ρa1E)W�9rf�j�jB��*����P��:�F�	z�,u�El[�'"�ĲU�h[wu���i<�8jA�DB��cO�>�Q?�'�������(�N�Ϝ��������j��o[�?�����BPA����J���^g�h}��k�	hʆ��Tbs/��v�|�g�<Ö��`v��!�K�'��V���{��^ٯogd�"�e&���P�x��oo@��m��C^��b���)�D���V<�d?�@[ԢAg�,�e�nUdfgW�A]ϒ��Bs��{Y�Բ��vu�S��qj���_�>�E��J*W xDjU,A���Y�HlU	��Īoh�f=F�8R���d�#$��eQ�GӺ���@���Kri?M��d��\^"v��H���n��Ӻ�B��KZÔ�JOj���Eʆ횶�z鵧�����Ж��]����.��y����M��ż�Z �L���e�:�>B��P��5\Bp?a�py�m�vcݘ5V���J�u�����j�%���Ж��_*�5$�w	�e߀ ��$eQa����:�\�w��A�\�����3C
a�2��Xs����%��F�1���h�3�_����gMOJ�������,ڣ �'U����
9my!��I\��5�"��P� ������q�"mהUbd�Qf|�e���˶��y��������)���C._�I+��ĄsE� 1��."�Te�Ɇz`�<�1b��^�@�Zu� ���C�?㓖�dn>�<`�+[/�Ap1)�^n����O4��l
��d8��&��;��ߖR��l�����9z���������T+섖��y>��8tKZ���u���}z����3-�+��.C<ꃊ!��g��LQ9��,�P}?T�a'l	��#��]�ͶTu��4p?7� 5����q�&���x�`�|G�M��aRH	���]/��W4��eS�D���_T����;
)J~�M |�N;И�S����-R TA�7�g]@��W�F ��]�'A�D�l<�t�hJ��qMԦ�$2��lDl�zG���,�6I8Heo�Nt3���w�-� 8w�5��#Eݒ���"��1�X�����W?���c�x$)>����n>H�i_�X�P@@���!�)��-.�q�8W>鋃l��9.L��%p�������LXm�(=�$��;�R+�iJ�����'N���#~x�W�|���6)X���e�Uf�Cx;��K�C�u�R8�WF�/��1P�V{z]��{I�vh!_�o���enB<p��!oҪ��}6Sγ8�|S7Uv����Y�,�r�u�����z���E'�3|C����ޏ���;N��;�G������3廥Ұ
�LǍ�������r@aXǣ��\ۃ<��Zc���#�h������C�
��F��Ӗ'V)���"����t���y�����J���<�#Y��C��/a��ԣp,�E�ܼ��P�ź�5\��X�J��q7�Lz��,�]rvV3�̛��e�L���]4�!�����9�R�/���^���و57�*�������7��֚%x��eqJ*u���kŘ��8�������t�\�*+�;����|�1d������:H�a>5f&a�FdJ���l�d�j*{!��X�WB��3N<V\<��_W*{-)��ͥ׬�i�%�m�8��6<I�-|Gmw��n�jX69 [�����a��N�=��fv޳�T�
ьw9�@���g�h���)vtd8� ԯ���ث��$|�E
�_;�]��9�y!�âN��X���	�o�eY�
�ӃI��~��@�������� �.���Ef;=Bu;zWf����OŵZV)���bb�'�)�	�Y3��`�G�I�Ev�w�)�{��O�2��랃���u�&����Ts0��#�*r��Dr	���?}k&|�$.�ew��*e�u��q�z���l��j?��kȕ.>0��1 [t��C�nAS�pY�f)yA1�I&+������Vf�X��0ݚ$�Ŕ����n�}I�L��Owd�E�y���ҏ���
���e�?K�Rg�Ҁ�� C��2�"�t�y�+���K�:������Ѣ����eJ�j��y�U.�J�1\����৫�1[=A�:_�(Q�cW�Ze<Jib�tLC��0�����?�"�.��r
�a�#�r1B}�w����/�i4���L/^n�&|񓰌P�c_!!}���8C8��h�,YF�av��j�ͼx�:/;�{ ���%K�!
�MC����f^��(���avk0�}�k��u/��z�9��ύo��&��͎ʣ�9���d9.���0�\PQBͶ�i�R��j���{"D��/��m@��`�;wm
� �y��!^�������^���{(p�e�8�(����F�U�}�(w$9]�h��$��2���\m��Hd�R�k���NnM~�R�|���Ƃ��etV@�~fyڂ�(���.0W���P�S�*�B{Y��ޏ�K
腁橛�K�d�<wrl.k*����)Ƙ'SBzL�K��!�>���xy�/M�ӥĐ��G�+J�/S݃���l�s�1�(~����o��7,$�-����W$4R�	p�ʘ�l�b��a�Q!�w=�'Z&u��LGP���!ݗ�#A���a�T��Cܷ㥵Ҏ>sd�����ҙ导[ �b� �b��� �H�͒/\V�(�·��}��>�*��>��M�;�f	����7����EڋB��ph;�/� 5�97O��c�ɼoED��X��T�QQw��cq��X�ef��5��"�0�7��X�q'h��_�wqo�_��k4�!�y�(������l�J�}��51.�24"���*�hS,��!g�:����X��{�=��\J����+ꇶ�����@Gͪo�ҬU"�L��i�f�F�Iڔ����Y���HeQ�*Ax���3&���x���|��[�VY�P��Ț�x��9EU	�J����L�՗3�"H�͸�/?���g��N�#z�q��d9� �b��1���
�`m��7��m�U��q�ݬ�A�^�ET 3J�;�/?�=��s���a���i(�zW�bFe��1�,�����_?Y���D�P4�0~2�&b�j�$�䏲A���:��!�+� ��i�R�&�4�mp���sH��1�Q2k��cNk����.Yq��IA��<��K��3�����}�C�04D����Җ�ާ\VDS��3�cg=�=\K3�����R ��yA/ȭ��'|C��{Y����\ G���ps	��?����"���|��`�=���KNǰ�$����N|��-E��.��s9�U1���&>ȸ�[�{d '�o��g��p�'˪�
��o���t�g[�J��������_ISft��;H,gdy�g�5�Y�҂���f�����%���')FƠ\F������(�MF��^$Z�9J��<{�g���#��������Ps^����g'��G��rı�0/7��_�FRD����:4����i@7nk!,e.�}��U��`��b|�A�ѠW?#	^1J6��D\�geq]��x���q�:֦���tHN��aDA�=��\��#�驆=pԶ��~�%s�&�6R��2���Lr xc؆a.�S>��q���.3h>�2�O5�5,�w�l�=�\7�� �3J1[�7۰��K���UC?-��k��r���6�ݢ��,�Δ��Π� �� ��M>q�m�E�X�%	q�T��K���������I��.���9�-��T{���>x�7=V�!#��!L�ji�e������fL�n�HBZ�w{�;]Q�#����˳nN�M2�@��AF�]5w���º^���y�q
�2�a�h @]��Bc��r��J��e�<� �ks��4f�{��2�;����f_Ix��|xҠ�I���X�T�2$8��,����Z����:I���`݂�V>_ȱpK�^e�����y9�(�H��%�By�0p�=���PP��M"A_1"�5f�8��vhx<�؏+p��E�e�A�y�����7��<�gs:�Ys�Y^�'A��o4=�=$g�fvD'ըV������n
(����g �BQ�Q��<�SE����9�c!m:eצ�V�ZA��'�� ��*�P��N�������<OG�R8mY:��k>�*�m5���(��n��k���h�;��`�gj8T��D0��!�����mF��Ah�/���"jI|����ݲ�@�$	m�[C(�꫅8ԝ"F�����W�ѽ[��;�D�q�F��r�?>���g����g*�i�>��w턼df"<:4H��:[{��0ߚ��8�E%�I�b��{p+h�G4�,���/�Ƈ��nx!R��n���[�d>�,���R$XTc��xӒ����5`�������Щ.ҳ�����,�p������9�<ܡ5��K._��q�s?Q����\�	ڶKM+D��(��#��4*�q�I�Io��M���{�@�]Qcrp n����܊�\?&����χ��x��zL��ipA�S�� ��1�LN6n��)]_$�4���v}v|7jHZ@��9����x �R��I�FCC�'��L/l���?���WE�Es����h�e�ȾU/��C�f���i3X6�ġ][�=�-�/����V{�e6�cw�1醃�d�:�������ݟZ�]w���5�X�1(�g<�'��w�ݨ�sD@e�шf�4�@�kH�[����I�U+������9�{��^�5�׻4d�����]��1K��Ωd�W��b��f�MܺR^���X7l�,�k�V����|����*=�8LX����ǯ�0~��]uQR�ز�4��#Lh
"+cI�,�H�'�GvO=�{�&.�p�ǜۉ'J��� �X���v_f] �@��w?�[�/�pM��4\Ob/��3�b����n��P�wS�-�lG��Z��G� ���8�z�}˸�Bg�_��w�*������Α�'e�N��\r|3/~[�B�~{RFu��mDY�@̻��N���3΃�'٤�?��@����䬲\D,E�/�8��.o��H��KQ�t8%�� �ڙ\�Qt�{D�mY�c����Q7ŕ#;�c�c�Q���I�2�2�k�
�b�����������΄��K�&l� �P<���ry�P�xF\!k	��ا�[�&.��}fM�x��:iG���W&mKyCĺ�uܞ�;�:���F$����F�HK��U=7r ���<��u���� ��r�P�c-��R�x8@�T�FܶKI0��]��b@k�J�k�	]���ԗ-��X��0^��}�;@wu5TddEr��D6��'h>�eA��d]��X�ą�������X�*��w��ţx�_�W�v��Efc2��c���?���]j�9�����ߪ��͠'���E�{�W�.����p�a���I��ܛ�Ih:����z�1����"�i/�� .��;׼�y��)!��Y��A}���pL�V*�{�,ʬ���_��+���o;v����߁H��{v��_dM�#�>)���0�?��Rb�O�0�Ǽ�߮�� G�60�g�mE�я���s��*���g��A��1�0Kq�r0�&�f��M�;�	��0{� }��ϛ�F7u�>ʶoW��#�'[LtB��:bU�&�����"'2<�� x���E��@#��[��)�c�@���k2�x�q�0+m�[��Ϭ���ħ�nlsV8����/o�a<r������������lg氥�#M-l[͊�j9�N�![�S���0e�o$���vq�y|���fU�z�g>Z���U�${�	��m��4BN˰���1F�c���E.F�"��~��#Ca� �9��G^�ᰛ�h�2C+���42B��0���3Y�G=�@�����e#hH�4����eju���Y06j��O�S)���^\F��?��s��hy���'H�Pl�~��H�
�/��Q��u��xil��`�F�:5�t�Ȧ���~�s0#�XLS47�����ٳM4�����o�&w��ph�yT%����^�R��3H^`׽G�_2%l�fW�qfj�=c	��=�l&	`�4�K����0!����\9,���|,���=5�}������"��؞U2��B��Z���P��+�w'E��0����o'�1&4C�Z
���l婯H�1�<=,�Uۋdx<�i�IbT��|�A��p��,�'��bS뀦n^"�;�����=�%����S��4*>����?�ؔ�*���2�F]7� �KU�k7)Wi��-��o~\T�L�ֈ�{+�9�m�N�<Q���P#��xx��n��kZR�v��ڂ�_�Iۮ�.~����hݼxWL��)Ve�4���5S�����d��E&�7���P,��"y ��.���9VA�o>�L��[L�U�í*2g���+C:b��<����$��c=�r��/0#�l�9b�+$'���D�N��4�O�X3��>& \�d�*�v�Ȼ���ٻ�Da橄��%��S��q�~4^Ŋ�U�K��A�&����j�ubU#�������Vb�z@NGJ��
�VHO0�^c{$����H�(W]	��O$�(�g�w^%h
�Fe\hK1�� ���q"&��/��*�\���PK�d9%C&��%���J̃m��|&%U�g�Iu`�FM��SϏ�Ba�ә`ዅ�%��޻A��h'.����XH����m����"v�YE�T�@���|�$��4�QQ�ҏ:߈
�c���x���aZH�8J�g��Q8����&�z�l��[����� ����e�h��F�l���ȄW�|�v6�ޭ��X�
��S'���[�ƭ��8R�!W����&��9�ۻ@�N̼�Ӧ3�T��WI��=�s7���J۞�V|�:m�ԟ�MB�{3�x���x$�Z��7�I(я6����W����
:�s��%��̖�94���3J�衭�zx:�Mc>��XQ6l�0��*��1�?�;+��p@�R��E���`�v�������F�r��L��"͔�}��3�B!D��<�s@ݥj�OZȾn��ʐ��+��6�K�N�Mh`�1v�R���ǶB��1M��@n�V����27_Y�����T!W𨣀2u(�����.�
���l*L���N@o��V���v���60���i�Y|�\ó��߅��t�U�� K���f��s�nf�=�6�lQeپz��?cg�I&�v?����@�Bl�}1>KO���+�dw.&�c��^�1$v�m�-����Y+)X@��ŕ� (�� j/H�[~:��$p�D�7^�GE�|�*�]Z��� �/�����1�"r/���ƻY5�j��y�9�¨B�|a�9�2%U@�7)X�͆�`2������u9�DP���Pe�����q���[b�ԇ��xL�k�k�]R�m�*E��Cpt!�q�ȑ��}��xFr1��F6����8�C��:2�%�n"Wh�����B����f��X;ǅ��]����H90��Ա" O���� ksO���T�s�$3?�?���V���!�����8ڻ�7+p�s�Ǧ��n���&��Yej�k鯫�9�������)�k�ICМso,㶃ǆ�6:C�*��PV�.I�7&�Q����Fq��BvE��@H,����K�����ԡg�9F;X
�O�1��Q*žFp\F������w��T�ql����>zn���6r�xSc�ҵ����k���yk���QdM��W$�c��X_�IYD&"�39�Z����4?�����\�7��S˪�&�*���b1�4�����.�h�Lh���"�/s��,�n���=�\ ��CfTW}�z!Sp�Up!$�)S���C�+��:,�o���X;n��p����آpU-�_׳�PP�v1|[���0d�ׄ�ku�2d��c.�kt.����[��y�Mr^C�ǰ�,/BqG��zy��0ː)E����iD�pu~舜72z9MC��H�z�
�c��G,��K��,=��π��ա��S��cǯ��2	���7��LI/P�����/�vHhV
�@xT���0ܣ\xS��P�r����(��V�=7df��� (��'s����=Y�֩W�&�N>�N(�}5�[�
T�qU��cP;8Y��CFmf���a��dlGL�]�[��ը�F��QT�k�.��d��"��4��#14f/��ö��v|����!V<,�~��|��S��he-]65Yk�g�V��Uqˀ��wm���"�ew��A�}_ڨ�	��p��7��:�g	G=aG$��d�S3�	�A~PV	� �z�@������h"fq�M�4J����~�I��;~�k��C���>��~�����LT�k܂���;�MF����ެ������/�^��"6��	��2g�'��o�^4���}������PZ�ݱ��(u(�q�� LD%'8/	�i�������7|e,>�P��2������D=C����<�G>]_��=���X|��z)�ya���4 E����_����>��Z,��Rw�X�zN?�m��Ҧ @�6^!�P|O�k2I	���S��ՆV<�ty�{SOV�z��~n�9<�<?)����,]�1n���H�k�5 I� ��W�s�t�N4��ωqR�^�0M�M>�tk_��ݔ�W�,XRDȱ������}�kA�.U|�3 �QV]�w`����d�-^�&س�G��1�M^3:lE���A�ݏ7ǀg����>�!��¬�4E���F���cOg@��Ԉ=v�t���	[H�j�yȈ�52C���N���hC=�8����������
�WS3iܑ,5M�c�o���*=���w�e����wѬºh'\�y��l�o���mDM�o������/T�!�.I�H�_҂�(5~�VJ㻳���e����-.��!�� �����{���X���8JgHDS���A7:4����������&���Ӥ�CO��N�yZ=$�~\%�L��H��/O�e��#N�o^��]��]J��wl^�e�+�S����U��y��}��v�������"�s�\X��=M&��/�TP�C	P�o,�!��5���AwL���Zf�Xl>���i��ʃ��?������}��.]\�����2��?�?Ac*-��o�N�@겉�]ΣN�o~�´S z�������	Yd^g6b����+C��	�l��6��2-��.�lGtl0;M��@�F�8fb��C�-4��B�X���ے0�,t	�w{SD6-l�����x1����w4��z��2Ġ9��®��%����6ҳ��M���C�o�<ݽ��+U߻�k�w���X������y*�AI�_��)�|+���z��H��8]N�.���3#��J�B\5�6���h{�Q����{^�p<AD��]���y}�+���O�e��h�[����$(�I^��( * 06G)�MWj����y��(j�8�)���a��=�cM�K�;��+����T��.��0�h��1'����[�3ˮ�*<n��Ǡ1"TAHU�r?6��-���}��{JH�A8}��3T,�&����.N% ]��)2x�8rJ�zM���Au�ޔ����'n����\��s�R�j9���phv�x?����!BΓr��i�;&�=�*��ƑI~Iɻ�!E��nn&'!AJI���.w�/�|�I�NNd�j�l�k��ϰG�f���� ���)�pMB�1�YoJ�q�Qqg~����
�s��._E1r,W_V����z��/%��1<�F,�^)�M�?�� ɳ�z�&�Kd{��<2l��ŕ���;6~D����}����}n*��A8I�V����o&���C��QLܳC>�Ud���/�}Vk3��y`Ȧ�����T-�M]ױ1��VOk%�M\+�}W��Ψq���5�ٽ�ŵ�~ڗ0����ǉ��CW���'�e��)Bܚ\Ȯ:�&�l�h-�V)�"=e2���r���I�MYL�lJ��)�x�*A��Q�-�Y7�"��3F�~��·�q�d�w��qB'�]z�g���WD菀v��� �D��N���2&���Q_�y�'��,a�wa�z����20L �a�о��yτ�0L��-4�jR |c4��1�1��'�/�qKۀj��+D��K�ͼ/g楷VCy�۠��%�D�?f�g���58��V��/v��t���wO�{���5�8{��~{%��r����&�3���.�0%�d@��%�a�|�D�^�9L� �y���vm~Y؝�+�G��<h,%�����Z���iI�7��}v��rҖP���h������(�Q���� �T=�l��]���H���-�95!�����ЋG-Ñ��i��d��%��p����`���n)^t����F����>.S���qC;���,2���Q���'7Ê���\�(av<�#� G;:��WK��ʦ7`���..!�ɽ���+ꡩ��B�z�t�Z�k�>o7ä!�6=�������kY��#4����:+q�,2�LZ��txh����f.��w��]"H`Q�ep%	6�W.\9lm�8w�o@�35sf�^�^!V3w���R5�B�]z���zyܥg'�2nZm�ױG��״�|�
N��ob!P�G'����v��2��-ý���cd���q?�PZ�r���OcTh4Y�����ϣ��4�nRA^�z@ �T�?L����4��w;�?�����p�����"����P��_Q��MӡH�Cv9n l�c*p��K!~���xR ��\�����M��j�y� M��O��l�GN��|��?hk�6����|��"?Y�t3p�i_�g�ɠE�(�$㻣j%r�XE'$7B��xA�����{8 ��t�$��UBVL�z�u���W�tz��M��:F}�����9��O��G_��P�e����N����L���U����P&W���f�A �"h�B�B�U���t`�z�{��@�n��I3'���bY�M��t0�"b���]lk���&eY�3�]\.���H����p��;ˉDy^�d��:jKO��!��,n|�ΰʖ��1kx�q"˘�P^��(b�Oa��4]T�@�D��/��&��j���"l�x��D�V��3�BDYw>0�����.3��W�k��@*�P8��7A�Xlp���Y[ չ�FԜ���|Z ��@����Ђ�C�Dhc��h���2��.������G�����A~�Z���Gq73�y�ƍ�tl��-����YȪ��&0��	fB����\��*���1F"�
c�>`�¯#KI\���q+����J��م�*�F/n&)�0�s�F�U2� �|��p�쥏 3�,�"�Rmx+�
��#f�̱�w;d"N\�+TY������u%�)�1���JU�2���"�����n�T�'�^����q�ͨ6#˲@�h� pf��Ao<'û���
HL���m*5�j�@��d�i72r�=}��3'`>#��]�52Y����f�ߣ�vXE��OD�+T�"ш��.�/~r{S�7_;���R�ΰg�a�b����q�-�(,���0�g�p��z�%��ѐ�m�[@��	��Ӣ��(V~ϷpE���1o�����y8Et����i�Ů�t+����3Q���n��1�}��)�Cv,�����m��]Vx�t������؂�a��(������W�A�*h�g.�CXd���4�%&Z��&5�!�D�mO��n�6��,�*#�3>�8$��Ӱ[*cr*����O'�
��n��5M�Z}�x���~���[��nH�����DL�
���(���Pu��a��<��7�q1ނ�0����8*�[��DV5s��^1n��L�d�	����z����@��$R�G��`�ڰx�L[�v�HOM�)3?�UZ���/E�%z�c<��T�X���t��$��������U�N�1�� m9��:���Ij� �L��ֹ�r���k����b����kkT;T�ê5$
~���d*x�!�R�����5�!�"��1A�]�ԯ.���[W`A�d��(4)M8g|��`ܥh��q��d�XD.�J��!
�l=���X�,@ Bm�K�?JD��2�~`�ɶ��\/�Y�;�D�ˋ��׾�l�����?~�O���.:~�A���^�3�]s �8�=Q</����,��,'~i��x�����bHb�%���.@���r�����4������	��(e1���k�m�;ʈ_?��Jy�4��c9�+���߱o2���sR��2�NwG8�'M���O���e[)PA�a�S����)o����#l�-/Tj��95�>'e+*X��rv�Gn���g��W�;�7�4l4b�Ye��T����ܭ�-�E�ɼp�8��r| �.A��%����W��{r�!�.6ܞ���s-s.y�#�隌q{�r���~Ug_�Ǧ{�ŠX�](S�=D{;쯴����n�iZ��A�����
��9#��®D�ܙ�h��N��t���0��u�Ps��]����+����eұ}���Nkc���*�rQ /�������(�8}c����Fy��1�cB�+�oA=�������RS3@��C��\�a9 Մ�(ן�Ny��;��X�_��RGiOqO%��2��Q�;E�g�)1cXwM|sQ�Hʡ�?��g��;GC�p`�CZ�Hb:LLsgh��YZ�+	�wf3�����MȨ �k����j�:kBF�'dX��0`������eB��tG�N4���zw�1�w�<�*�s��U�£~IJ�Rf���-o�Aܠ#*�iK�¤J�0��KN���N�
�H/z	k�Oi���,�Y�^�K��ݐ����%.�?���#�'�Я*��x^6d���a{C=
M��]7G ���\Ϣ U$�U��˕���CM!e	��ƀY�]�$���.�~�D]]�a�����ܠ��v�W!��˸ki{^��.(������7r�k7�E�e2~[�A��U#Hx K��wx������Q���������Z�6}~�Y �/�C�a�%���A
�%x���ulB���¬��
Nb.����*J>�Y�S���ON�% v_�ҿ�~U�J^�Cg�:��$g۲�-y���/-ꂛ��]��F�j�V��5�)J��[Ke��D�k�� �{<�#�������0��¢�^� �JP_m`��.tW8�q��mS6� ���ޜS����!����)!��:�?�X�Oc�Xjzhh�Sw�Y��v$:�.6z�o�ؽ�Q��	M��b�ˊ�g>XZH��?�B�6��i�a�Y����C^��] �s��9�2rR�\��<�J,j/:U̫:!�m}�|PBF"n��3)��NZ7� ]���c߬���_ ���9"(��(bZ_P 0t�\M*e�&vn���'���媪~�\��5����_~��ӈ_��Yy��2��&�*�^Ʃr{ժ�خ�+����$Q+����~���0F�AV=��5��$�P2����Ͻ�m ��Uk0�I�K ���F�����ߛ�,�1Hs�O�`�k<=�f�q ��D�}��qr&�u����<�w"��dW��m���Mb-�;�L�u�=�_��TY�0��Z�-2���ؿ��'
"�"���d���@V��'ΩQ-�kGa��&���3Z��#�<Ù���V�2C��pu�{���&�8�H8Nu�g���Sț6(yWÕ`���@ �9���(@_�B� |R
�Đ�$�Z�":�T��s���UZ���N�_�&²%�,$�kͳ�����ܱc�Y�K�q�t^��D�Ը�+*��1}�|���.�g�N
~��w��ݧ�r�����L�qo���#����P��[��}C*���vLѐ$����D �k�`h G�^�ɤI�̜4��W�w�^�����t�c�I��K��ǯz^^���.���2E\�LҚ��^���JBI����,+��"H��5TQ_63�#��
V��hv�����O�L�P�<\Py�.�|��L�2ЛY�Z>�&�w �iF�-�r��@1��&��?��9E������\HC�I��U��,+a�`g|��������Ћ-S/�Oi��h@8VCT���/�]��&�q������T��_�Fs�11��w��K/b�n���/&2�(�V��tZ�	n�LU`�DH��S�=��mK�_(�Ө��A���T*o���<����O�<�MGU^?R�5��u���Jk{*|n��k���4NL��!QbY��4��K(�����X�/6G�d��i鐃�mZm��@�w���r?آ��^�t�L'�5d�E@��5m1I���������W�g`O:A��nm��#H��s؊����[���6o�z�Aԯ��I;Zrݢ"�d����A�6	{3�K���z�5���[\m�z��1�:y�h��clZM���;���~B��A���r0+'�]�����΀���N�Q��2^�ܚ�-�枘�w���?I�,ds�W�k'M�����}�
���{��)@��r��!����-�St�{�	<�^em���'��-���*�Ғ��ښ���ƞ,�7g-Qvђ��r?��9��쩄x��4���L�A����
t֐�T�oӜO[���&Uh%���ѾO�F�c���0�P!u���:�4�w�-� }D�F����w��.�y��_}��{�3��'FT=:y�7�+�Vw.@l��jfVR��->��%@�q�i��}M���jl��|���ߦT�S��1�Ҏl�~�����*�e�^7v+�y�\�Q�
�|V�|�ϙv�N�֘n��b�h�
yήztga���@���	�uW�c�4`�}�a6�tvN�5Z�����>v:bp[�-�V���\ja�O$jsD�`ѹC���w�7��X4�QȢ��_�u*A�Z��@!����Z�8z)�{~���f���)�aM�C�.��/ᳲ�кa��1z�Jf��-�l�	a�~|���襽/��W�`ED�h���n�`�k��\�z�j��Z�n.��v����s���#V��I=�j�(E��vzR��[6p�[0;����D[��_�� v{C�e6�\�(�K&�"�.e�oɩ�CwN�?l��gn��a1�}u���;z�����u���L��&�����p���D���d��c@��������ӫ*�
��ea=ĳz������=<���r���F�O.��O�J����t�2l?wܛ(��T&�R%0( �VJ�k�3�R6,�j��LS���Zm|����70(+	 �G6��j���ɖqى���������mg7�/ei��;���	���W���E��(k���HmԁJ��Ǡ0䈭I ��^�=���4�&��_�%��wg��݌�[�3j�X������У�A��_������1s�&�ҽ��:^l�A�|�qJ0;�����n�MU���.:�����0m�&�)��^��z1#�����M`�L�,��u�	���'B?�Ӻ��o}=չ�W�v)~���OP]�����Y��Z �w���mK�R�덦A��'�F��,�י(J5�`%����˙�8����$YJ�ɝ�<�J�g����[�Q�5c��l{�=|���.���x�.������K-!j[
� �ںd��i�)}%�_����H��M�WVߴtއ�C�{Ieuh�E�^qu�O�l�Bf��� ����9M-1����'���؆i�j�o�h@�p#؅�D?R��*��2[.��:�>|�8���#7&U����Z�]!kn63��T�X>w��PG��w>��mx���T��8l�i�	�G�Z��f�����d�:�f�
�"�ۍ�P�J�ѽ�jy`g���e����n��4^~�@��5��Rv��y��K���3ˡI	x4��ͪ�ab�FA��Q3�"~�V�~��1����P��Z�J�8�R[)��E\�*gQ�F���2"0}�G�AĻ��#�������:m�% ڦf|I����Ϟ��/y0��I�/4���Y��}|Sx���ֈ*� ��h�}p'lW�����	�87��ϕ�1�K)h�N	�,Q��c�\yͥP�M���<�_X�K���J7�����F,���/�L��X�<kD����M�k��v�k�r���2�%<q�un��Ť{�W��[#_��YV��-D��%�.������~��f��C����$"�afXS\D�H�C�RL��T�:��ӻ^D��A�ABʲ���K�¯��߽�^���MpD��X�#4�}H�{@�YQ{>8�E��K�:�.��!�ajO�Ќ��AA}�B������
vB[{V&�n���oF����ǘQA{��b�Eu5:���˞��k!`N��)vʀd�+_���GmU���@��Q��+4�ZC�}�|�,Uә�{�Rm�eW�PD�3ң���D�1>�M/Ш��A9����w6�ZBp/4F�WO�?�|��z)40
h�%���e����uU���3��g�i��<0�ꌊ/pci�fI ��B��Vߥ���Uq�p�.���v����$�Z�CW��h_J�9�xZ.'�_��^��y�qԉQ`�!��P':�H�ަ�uL�[=��T�˽Q���#}��މ�
bL7���'O���d���B�{�er]�h���z�������`�g2����o�86h���j~E�W�c|�Q`%�g��z�Ş0_s�t1��sA�]��$���鰫.6I.�vj��B��O��>*��$��S>�pݿ�a|(
1�����m�|7��Pǋ�B7����`��]����^j#�td��Q.G95>VX ���ƉQ��,��Vt݌��\�9��1�V�������K���V�;�h"v��@�܄[��zwߒU(�6�-�Zi-ɨK��}5bV �Q��R�^wߢys��XR
�D��q]&C��w"�Ͷ�eS'�{� sc�~w�觺�n�Ⱥ�# @o���ޫu��Oyl��]k<$�F���5x'e�=�L����>f�ttxh��m{���C���H}������������m'�nl�|;>�a�������P+�}h,�[��p</;Vg(��#�XI�������Z`��nC�:�wd�rî�R��.��@�\t��]5t��~a�I$Fp�駘��i�)s��Z�7���ܭ�sF���C�'.���wm�I�Fɢ8�vB�n�f�m\iŃ�q�rN[�B�ۡ��0�й�	-��Zx}P�U0+d;݇_��Q�f���G&B���)�~85zv=K�hd�6�0J2`��g���_�9��7(Ql�	���77��;z���S��V:�)���/�����<]�ٞ
��5�3�v��p°1�r�9��E%k�c��?fJ%_X��,����fA��8V�5*���_��cK?Q�Z6�{�������[�^290-z�n8�A��u H.�詪��T`L�A�Qg��[6c+��}"M��O�0��ZCd��h��}*񩭉�4��I&�L�4�⩻�>:��R�����d$�
�����+��3�6�1м�k�S>&�����0��l3���ރ��R8ޡ���rȒt��=�쑂g7��%���A&"��bqC��颍^y��W9d�qZ�X�K��s8Q�����Uɔ�z'#��nh�@f��Gf�P��a��
�5H�e��yjW�ܶ2���D��Y	�|kZ��؉��l72bK����d�ȵ"�7;�M�R�
O
��[��Ϫ%α��kXkWf�YH��+�E����/D҈]팿_=�k�a�	s�\aJ�ί�ԟI�e���������O38%^���;ƹQ[�ǃyl8��س�K/�Y��E�	�����ȉ�)	���o�TE�qNG۱O�E���.ol�A��x���"`Z׈��^rY(��h�"L�ʽ��L,M{K�ޭEu�����Km�
�w�q߬!���a�H8����ͺ�_���K������w�[*�+s��T�+��(���q;$)�;@ue^GZ�~�W?����{e�O�J�����g����=��|:Q���]4�-M�.E9y�����/dV�1��'^Z�K(���KF�y���c�����~W�U˺���TƤ���*��yT�`5�, �HG4�F���`���nbߧ��k���
�<�]s6|g�Vj+f�8urޯN�M��>����em>�����w���d�w,)K�C��<�
 ׺��&��h�5��;2~��g����q�ˏdw|`Y��#����' �G��y�_LI��G=�f�uy�������<�Q�'ЭN�I���~���e����F΅v���ǫ��UH�h}�7D�TU�	�:4gHC_�88���?����h4���)Q��j<�ͲysC��u�5�ݪ�7�YD���UR�rfU����3=�V�Hm(�?��_['���!��Vލʅ+/_P��x)l!/ߜ-7�)\s��\������NE"زU�����WR�h9+$r��!�h�_����[�FR��8�&��=�� m�~�9�R9�C�X��9(��\<�9��� /�R�����:z�1 c�@�_�/�Mĝ{��	�(��&���_�p�̘��������e��S��Uނ��07Z�� �r�a���6�/iƦv��eIE��r�AUC�������wp���΢��G[�!�(�F��^���W������!�r�/ pt1`��w�����(Y�5s���ZfF|�Qpoж`v6;-G'x�33��qd�ؒ��'��sr��=��q���k+�G�S)��u�ݙ�V�h��������o�~o$#��0AI)��^�/6q���ګt��q�i�y��]��H��W4����#�]���lBn�\����R2��F��i?S��Ch&���-�.����A�z�J�j�S��4�};(QU�T�SБ��s�+N;��X�_)�ܒP�Z�������hBLBTf��t��D"��-�6tE�7��Q��ٽ׾�N��eBI�i��j�yn���Qp.O�[��< c�ʥ"������E
�����1���6!����,�Cs���^0�׈䟒����G'!q�Nu��)XoF�xy9�?���p��/�_�meq�����W��MY��T�DLj���䬝�*�P	�Ө4bb�d3�Oe���M���< ����!��0�s]����;�f�eriς���1u�C��uH�[��L��,�c)���p���H�9Kn�I8 k�O%�r�v&�:�`��B,F��?j���a�rYZ"��a���	�,��DWd���e�i�B��B켁1�u��^��.	7p_�@��R}
���U%�>������%�}�j���Q3aJ�kq�lЖ4��TgLrEN���-6���y��4�l��h�$C�>颇�w:�=�O�����o�'ZR�ԇXwZ�JA�4F0��%��]�	?Ȥ��O�$a�]�=�@���ǽ��si��/e�~���Ir�B����wS���Nf�P�=(���/F�p�H����3�j��/�'XN�i�8��C��F) �U��8Y��r�Ua
Y�F�� g�IE3��-uÛj����O��.�h���ܥ�f�%C�n�C�${�f�Z׺�}��:�����o������xI�MU2!�\
������4�	�d��ƹ��ε��KP��	���~�ֽ�g�{��x0UJ�ˤI�de)�Uׅ��˷���	��·5%��P��=�Q��X��y�*�L0�fݹl�P����@f�2��k�lN��SM���M��o!� �>�ڸ�?ZD)�
�N!�;���d���?H9�B�V�Ć�́&�7�_<����{_�W�ؔ4^�pֽo�0Y���s䁧�����F2�ο��E�z��p��Y,땛6�<7\�4x��)��*˹8r�L���Ht�B}R��B�I�$fO*ڎ��c&�d�	�4V�;&��(�wR4O��5��LL�}�D6�A��}�ʽ4<�< 8�/�.ސ�K� PF��c;��l7�\x�6�xl���i*�W��C�M�"b����7����A�xo�tNiy���M�_�'���w���!��&�F�AN;�~FK��>#a\��`��H(3!��X�6��d���$n� �q�Vd���`U5�F�9�*%&����n �6���t��]��CU�0�;��<�u�Y��Us����d�#济�#����aeF����A�8VFԭwU���`���ܺ�X�3� �B>�5�;Ѹ���:��
u���ws�.'������L��r��o&3?E&z�<�
A�iG��.�w�����oCR��-�S��d1x�<��j�|Ę��U�}��u^h�_�}������Zf9�T*;Blf���9
��lu�_�r\yX��j���zax���`�27?֫���뽹.		A6��m��Q���_9�C5�(�wy�j��~@�MxD��˔�b�,>�n��DJ�LX䀸�9��1�AT~K�Nc��Nӕ^0���킡�[\0Ux�)/�7Z�oJ�]�D( ��+��fh`��
�o\��Spc[��V�,s9�����:��d4,��F�FT���Ir	j�%t ��i
K2�sa8���ة��S�ZsH۬O�)O4���D� g�Q
��!��.�r���b��M~�d-��f��`{ъ87�-���#����9�&�/�y6�r=�tt֤�=��i�E���"`��;QJ��mKd=Y��4 ϒFQl;f��N�O+>Y����U�":������$�����ޜH U�>����L,m���(躄׳����Wv�K�ƣ�6IK����%v��+�Q�/���'e�[	��d��((0���ھ�z'�t9�ǡNEĜ]�-SkO����
�x���`tR�͆�s��m��X�,��Y.`�%=`f�W�gӳ|���P��[�˥��ji�Dl<�S�������ܓ|�MW"I� ڸ�0�ʈ����NZlb�s�S��\:��R��8�� R9����k!�Q�)xȞ����n���adT�������'�C1q&��&��@���@��^��o��[6��h�K�&ʒ1��j"E��H}�;���S���P)�[w~�a� h+��<��ɜ�u����
b��2X�'M�]V�<w��;��k�)^�.;N�H�*�V�n�cơP_�mRa����8F�A߹�T�&�V�8��+=�&/��ӝ���n/�7�@@oQ�+�(�{�4��G�h"�n�^k���ʸ��"pN.��i{����W�@�΅~(��v+[��h�n�yS8��\�$O�N�h�JK	Nt58q��Dq���A���B#{����6����J�[^4xxWA��\�?����^!T�`G��*�]�|����c��I�G�99�z;�pcr�SZ���Fh�o�j�I�ǃ�2�,�	�6~O��2�L���������ݢT��^����P��B�l�I<x����3Vhy�T�Ț�n,	vr���>EJ8���{J�l�͇B���EJd�h˭�dO��J�K���o�	k��+=�q �ڨ�M:��7�Ͻ]�@e�k���m��s �<1������������WE����m_�9Aü��p]�юD�|8�������UH�6�BTztXc���R��-��'�OuJ�P�M:�~j��K;���sϨ� ��;�$����4��b"|��N�m"���dO�cfxfV����,�����SX���W�X(�,�ѵ ��5�q���p^�+�i����+Գ�g�&����W���¹�d���g��̊�Y-����Fů�"�Ѩ�Y���Ss��Ra[�㱑$�"u�*W�;Η�?s����X�a��q�1���a�5��˴��P�چ���3M���A.k��vo^����o���<:�q�������^��1�v��"��c\Cҹ�|��Sg'���5U�}c��w��!oAn�j�n�*�7Z�l�[U�Z�S�M��ݛ*�'=۪�g�7M�`�]��2`�е^/���~�^���m�����j�{�h�����j(=��������٩5R ����`Bi��/�!�.��SE��;���&���]w[ �������C�@�����u\U<~s���>�qz����i2# �`z`;�� 2�|��45hf�ب�n�b8aIr��	0�ӆcF�Sp�x��q��.���jE<j��{
���*��	�60��d\S�J�ǵ�V�a.<u�i��_X��[����O��ֶT�{�[��}�0�ԔX���(#t��e*���`���K{�q`%�lr���d�z���2:#J��8s�/>��e�x��1j�}���ƌF-_hN�r�B�C�����Q@�e �L�2f�>�O�	���]Н�l�u)+63�Y�2�~W�H�9���6�=�� r[�� #�x���� �E�kV��֟���y���wo�C�/g���I3r�C��X��nViS�p�Գ�r�	�z�������в	��#�Z� x^��v[�	�K�0p Tv� �G׾c�%y8O�(�C:/t��3ty���MH̒�	p�����r�	���U�;e���5^��:]��s�FTt�\�eb�x��2X.I1�'��p4{���g��`�گ�Ψ��l�A�nĈA|� ����a	���H�-�B��A�~�
d��J����t,�)	�I��;9w�?T�G��$�9\. �=m��P8����=f�9��Y{w���n�>��`�p�BG�g���p��]�-�HĈ�Y�g#����gش��%k��`�D!��]��%)�X����Ћ3��C�H侵��[�#ɏ��c�67�t�C��ȿ������_B�K�i���F��mwQ�!�|���1�M��=&�Rې������%r][M��k�bX1���B���a���t�	�@dM︜����b;~���sz�'~��~2s!6_�ۮ?H��#��=^�8~��w��d��z��I��Ku]����Z���v鿁�H4�=g�Q#TMdL�0�IFmw|HgJ:P�k)x�� ��p�S
�.w��.�?�C?���U2��o!�7"+�ވ	�Bnb���Bc'k�� �Iͭ��<L\F�<v#��g�q|x���riO]�����&�*�Ѡ�Vܣ�N2��7�"�+Z�=y9��]�`�iCD�����%D���P/��_�feM_,_���:v��4��7�Y�H�p�=ǗLe��B���hI�l_ ��^?��D�G���+P�D�Î�.�t�
~oC����uK��4J�������z�,!5�!K�/J�VG_a��a�i��w1�j��k_�-��37;����o�����nN6� �\���s1�plWbPq a��c\���!Q�(�^�임��W<�9��_��`48��zY2�Q P�����2�;U2��Mb4�o���hr�p2nB���%�[ʜ�<S�G;]�ꖼ@���/1y��kg?���yV��E�}榬(��g���/O�����R�;�@�@}��������^��