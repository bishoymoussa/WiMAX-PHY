-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
fZ9G2G7XNlHJHNOpusriaApj2X42mP8GQe5FyIVjhfsuGv9fgVrZMFsgWFPjyYwNaYzM7y8JKm/a
Vxpsh3qVAxBvla/C1hO+YfoSXD5IDEHZwzmxfJMQNYlqLMMQfDdgiXQFViafoJdasINFqRiIMEia
XsnGIiHPYVkDd1Jq4qFwjcM0M4hKisu9aIyhIRWCjyCs6SE4ox3z9znbPSChqsrb3j62Mf3MIX/m
24ydiJasS+/srvK8m7UofjC31AlDW1VWeWhgcWwJEdaGXxbGD56vTpFcP1aNJFgSsxu5Nf4z1IAe
xDFqOV0nDH1BuNTsP+oJvXUP9qhPePBHzg5Tbg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 26880)
`protect data_block
cZxXxCa2NxRWewMO0AuAgA1N6MsxAx+mCjgFuZfb3ADMom3BwzDv/5VhiAWr/jGaD2tuzWfdSt1a
hMSfi84C4i1B1cypRmpDmCLi13GOyx7GQARLaf5y1zP7CmMNK0x8/A0H2FZZMfHSggPB50Ykq/D4
Vx8yao4yGrAdwwgMOtVBltXJPFLzqZkysjntZ5ZcdtOW5GgCXSmiQWWbpzDH44Abn0T2dwFNZeN+
/NmHmLfDeM+rvVefpFR2zKYB5ehqtSS71E1EvSlCXQlY78mWhl+URS0Ilk92MwHrxLxqVGTYtcat
jbka7fD3EWrWr1L08kUebIUQp1ma5W006TuFq2vNVvYH6Sylt349ZXKnK2adUjxNPyLoQ55g0eP2
S+fu19XH0iuvzgmhVPVFF1zS9E/eaKKZ/y6SNr4nupuUoF2r4rokA98ubLsbIfklBDQjU7MDdXqU
j1oQHnFldCCn4PfLDtfnjikQzVXFZnDWJ9RTkR7NCSm/IPRT6PgIA8un7nKkCoAwwsPQ/opv0byg
UCKDWZTbqRV8VuBoknmcj8xcwFsOr+NfOK5bGUyPuoSrXj+L3vZrkljh55cD5iJPvmbOfwUSDaSw
CzQ2jl/i6EpOFtc+czSDVXFdFjmpkridn93VxmB9TUMLeoKO8TxRjGlGX0Z/88gmbybV0PGFPEMH
gJwIa1bRC16LX+ADsvLBCa3HF5bhLwIkCk3q4XqH24+AvnmLX1/QuCafwZW5O5VMLIZ+lTpttmf2
Y2qYOVoalks6TR1W434TTuKwlQ7QGfevkeu8rdJj0jffr0WLY7iWg+QV/5r6o+s4aPhSx85lMyD2
8xptQYeRbejfqQ0ZzeFyO7D8R9ZwKv3alfR0lP0C/gK3MPUvcefYD0FiA5AtOhvkTnHHl2ZpAqZf
yRWp3J7fr70OBwxiw8BzYKFXav+8TvMejPc8Om67tcRpDzeptJadrzwTH2NphKV4T2Ml/3eRT/O5
f46dQBVy7BEFtQlk0a7y2OotGE2pmC5FVcPlRD+E0EWCQomSD2G8z+lr1QNlk6ZlnH/MnQWWzr5B
B1pIkkrpF9WOnq+Y1oFW64U9j3sDZ7OdJ1k2dO+LQtJvie07fEShsOOGCigUK6th4bD2yHCCOdu7
YqSiLf8DRaa5LNJjACTl1z+UXgQBsy1PyE5tfZDb68b01+5levB8ZIGdgKdX7mSjlBarOKDzld5g
5HbEVaAAX/++em+jS1nK2e999hUZsL2j+1DRiGAM7cT9p5GOXg5ZRQMKgMr7uFDjvcNi/VTQWh17
lCYqwX7aXJY4knHywbghTwNflA7x5w7KYQFX/M5dNMzTVJhSZFqhKFRt4M5qctNig3UtQzyRRY0Y
lGpmngKKANFIkIY+y/y5wAawxryBXzm7GAZjtv5M9S1gtlkH1kS/Qso1ZCKjPiQ++3sUjTRwE/VA
rwBO763JVKsHANv178A5wHiTF6BiyjTW+qIJmDFArSvjDayiXTINLMeMZMd+dXpwI2yupsl1Z7IF
x7lwgAtY6JAg5sDAzLNSSPSyHtu9Q2nA8yr7c0eHQcawac3hqVhj+OTSUaXMbw1bvDFElRuzrkgZ
Fxt5LGwSSOBaUmHn5tw9UErJqe3hvYZfHT2zwudGH95kv7Aj+PxyIaPhbrUGS9SBUHV6mK3A4LJG
H25wbyub/Zswe9L0ST7mbvhXcO9lNgdJmHYVhlnSDecMw2ehdsGQCpxbOiUYjzQcKxe8TYe8S6gp
gA0U9F5EoEVnz26RXc9GuMw45ZmGRM65hgeKR/rRakaDuXygj3lQDMW9s3QhiFgKPsvcwyVsj66Y
uH+QGN0Uz0y6qfn4Aq0Onz3MrFVFyD5clnDscwZDe96EDHc9W9jlwpyDyOh/haS+j+cRi8+vgonn
kf+vHPWI1bySv/mN+QtIgOx/oV2sKuejxixxfMowGkuron6Qw/QRJdiY8H6N5t7mr11PBK9ZtFvJ
1yRAfjOpjB+BF6Yelj0ha0K2L6X5ypfprQqAAybFNAiSO3hecm4d2AHVmQPY7q8N+B+Hk4y8zzo2
5DUoJoUUEVCfDbrmF8cs6E065zSWtjNLPZ71O8cuwovcmDP84cl1ibEHCav5oCVuTjKjIX/o//zR
M7HodOlEEHPjcauDREURSa9c1vl2EURH1HtLq2r92/cjzMjH+EHwBy8EJqj+oaLxfjG1zwd/0zK4
bGDM6cAVbBgbx5hGKuzTiQMmphBfO1PGp3cqogFnoBJicdYSyhRUyph9Kholy6q0FALyL33S0Ypq
k9I/M4YVb+NUsIgOuyBxMUybNznahteq7qjMMjJnNnFIwmRhE4heLVBvLcyARbrKbC88Tq6Qj6pQ
g6XGvwfLYzb8ssf+JBmw9KLnwFzCKpzFX/u2+X0N/bhV/9YUhtu35R5WajDVXRI9BKQA2nheQ1fx
OlWQR8/gaxfv1C0S7sS/prHhCqxvtBGBeTVFrVNCMz/T4SOqKNhFIZGVGtImIAD50SuZ00XQN4Rk
MbxSTDa+hTSdwYmtl+ona8lIIqsH6vE8vGnn8TndIvG+R34AjrfNPqK4AmgSW7lS7AxCDcK02tZc
0p/drjNJbkgCKS097ixcebcx+J68TM8oy8m3uJMIZG3qTsnCszl0/9eHIPxqZ4fzE3AFpDZRICKR
CM2T1Skl28Y91fEKZGsLi/hHEjqdgsZbAh/YfoX37lFoNLUiQF3/NZzEU3UT6bEePvA5Gtr1K16I
EUidvQ4wIHK7IMM7HIEY5g2RfVN352I0YEBdySaexqW7aPyJyZKS974WATyUB6M6SCYAjDxrs7TO
AS+Jbn9TLB9DKZC73/w4vip/7JO0TVBcToNA+I8duubXrxllwF+Cur2jvbTW6VaS2pKqHcein2wF
/QCy3OYXtic4mDAjkz/xJY/Nc309X9XBNBwgL1EN6B3FuZn1nRl3xed9IgKAedH/4ktNkoYH8tIl
YWGsiMiC4/aI4xmOh5qAQBzSiwW1W7CcKMIyahjJotJQd0bYSH6sQip2luLFpXcMbAPwxAESMJ0x
G8SMypretGGidG/WbGWKuArTB6GI0qV/xZ/ahQe5t7Rc3R7qMuh4W0cHn2h8Bi13e8TnIf8Cu9mf
tTLn6cmimKiA0CX4e/j42Ev3b1IAhu7zRaM5ZMJHy9A117af3DV35DVbf14VCSLVqndK48FI9iRU
CDAQIQC2WL81bnW/jPKK4MGA76rJkK5Yk7IZ933oOoGf40OPDfpvBkhOiJkrOdPqtm2QTI2HcwGE
BRDnHt1mjVpIyYZ+nuLkXeWwftXWbcsCWtQ5vjxWh9nmuVZLHt0w1twA1HsQNzg0hmnZ4dZxMulZ
CFKhoS+ddQjHh08IvosTiGwgaeLEmbL5rZ1qbwWE3Mf8gfVXzfCeLbpFh3FcBdJANgACz8Qu6SPT
a/ygl56xQWxjFoc3UjYKzMsqoiyS5qq1L7tK4xkipqd1SmBAfgc3+9EGmZnPl/NC9d/Usu+2ZJeO
T9Kg/AcL+5y9HNoTRqR5G/XDVJhgOqCURYmT3jO9WlKyc45xf4Qic9op2lhBN/sCrTUhFbpL1amT
/yRtxZ3Mp/FooSrDjvdZZDOXQw1MZP3NJ6FfW90tLW1fBuuSR2pfslXeG4pVCVov/RG/ERGhcPKf
UnyleLa4Yv1u85hK3ZGyJSPTouTgGzdSlJ0wNeeGzwPwN3jHPnheNKV/nlZcuNp8+VjydYiCbesV
9TkhK9G7RWNUwx+ZQq+O4DPYX9J9HeotWKYo0LshxbHvAiktpZYdJGyPHhaXDb9FMZM3m1X2huNe
WDScFNF+4fFgY7ttIr0H501bTbEakk/2zV999tFgVsPj3NBH5VqmKgtgjbm8asPxhkhd8nR+iw3Z
BQOyeY7BMBYpKo/oDy+8hjZbouEWdCsM6V9gF1I9BRujFv8I1JsvhT7RPkLcMNNOP0KGZLgZmqGv
aCjSGOw6eh1qc/FiGNhXIZzXXhEqxvEZniMuxJ3VBOSuWKIEJAhSDXmBdyTkZPZchK6lz2E+HBDp
DEP2J1XRGjVWuH2fSk4LSxV1geiF/20Pb6ampVaod0qmZQHJxH90tgnCnWO9sqFKfMgxwnD0LEA9
wS7MT5sVKE1+yVN8WEV4CV4WhveDFzNNMsOFCcNAiIAtd4iW1iErjDTW0unQ7MKwsx8Od425qn3q
IvZ8+JK0zwrVJMum+xwp/Dz3RBfVuT/KINwViui4OlE/UWsvUmAZIh6U2tueuyNqpKff9ebaG1u7
YwSlW1ZkUMBiGVFfalDxCMJ5kyXg/4AxGhTDtKcjEJ/MDO4iXkuz1W51WEnnf9thpfNHBmWs5C7D
/Jx8QW0SwHQdnBZ+y9layqV36xJ05o0izffZtU3nbQNMO2S+k0JetK1Od68kZbbhWxQah1qQtCyF
q5+nzMzG6cumT2I87JmPu89z82/jRUh8zmf6Bbviv9EPnE5jMPqjfK5dCX7Z0IdHmvGQD4fUtt9O
so2/lQs9d5xsh+YjeDA1AAqj+EbKQfYI86Jve/PXuGUMgtBOXxBVZvkd75LAGiGg0LtRQcf4R56T
9ZgXlgyshz3p32YI+gdewBUw8td/nQ8OP9eB8WSbrg2qybfiVlzstEmOrvCzZGf+hbcDCEn72XgD
7fjmwExeNYqGz5zkeiI8dZMZrSTVoMNevxOnpVniaoWs5ES9D3NlTSQK3mKPEAy9E8UlblA8/CJj
KIjpcNJmeM9W4GyWdXhV+w+FvXUBvK34WW7HsaXDQUQo6oaFyn8apS7p5CqkmsH+YDEjQkzdhEJY
0otTF5VONd6D/yi+XvbMUDP8rRmTSviGRyLw3YF5EVqNl2hsMUhAIxc+c5yeK3XLqbFQ73rgaj0n
E57bsovY3AbLH2dzt2TYn/3dptch5hRmeBmY1OLXh+cL73zhWhxUgo91XfFzvNRVplVaxn8pgUi0
jMgpr2LqoCmHYLxMmUv/dzw172MJ9LCIf0jvwv35Oxk7N/6ZeMaZEzpbaUXx9CqWgD6LNHb4cSxO
Q0IGGWIMf3uOqngp885J4wYqvANtgqzoQ8X83V8bTB0utPWPmpMcgSlznOQlft7HeAVNhG7yAwYD
h+l2DGP+xoHyQ+qF9DfCN6kBWdCyQN9rAJDio9KJhGXemQO+BPiNwNNdyZK9hdNhz3iuIwc0TKCv
rodmMHSz2vzmCIfzgWkxOw/MtdaV79yYb93CUG0fZ3pZDYi3HR9ZzD+Ub7F+Vj/9o5YfnY+MzFrT
6AF0PEWse9mD0+anM+bImuoZQqnZp9t95kU4J2G+A+DhIXNRGOP8cO2o1YEOe7pFzHL4d7cUpKBm
Bl5mmIW1+A62Sw54zWLV9NEL6s/hrkq9NV8wfsi5ibF6gpzIqk271yk35mA+304yp+oLgQMdePax
8H0VhCd/OuCplDh65hhvKYnprdcl30U56wCc73NdUL/AGNJuhhynzcwqsgA8HBenJB0X3NhWEjKG
0D9PTD6SnqXByq+G2h/A0Q7vzL5tVEIuMCOI0HckXKgR8A/+sm6nVIIRK0Ttd0LApOjkUCo/sd2R
4ZDBk3KEqeNSbU34gFS9lVoM/XohP2ghTRA733qCLyuTt5DSTKKaiWj4oa2Cyzn1sMKxQrEdysdr
Y7qQPcOskm9hPh/0SbfiLRxfM/CRYceCIUxdoqxzHSNgdzjtHblF2txLYM/wEGRUpkiiZzOdfsEK
DMJhQ50J5lmfvqVjW6gFCXy7b38z9meKJVRbBb6yfaZcKAiXFrIlJHhrSkquF0bmGq3uGHsX1FCR
P141r0l6pt5rGFsu9lcvmej/TlNdtDl85KAY+VCmBhiLSl4ak2bBjSLigUp/+MVQCe/zIPvhYnNZ
/iR6SmSNV6gAaNjmyjwHmtSXKMKi7nAIqwa2vw92lzGuZsoaAOoTNNVmSLYgn4MVLfmgUzjRtbjx
cJgDAcfNTb+0bUZBiexqDtD9d/MhOvbBrUC6i2a1OsYvrpaRry0/f6vcXOse3Z9Zs0WvpdYumBYY
xsZBupSsiPCrQMJ6uhPt8y50mEXm7ZVNGmsXpR8FT1LAJclbgZ9tiKwCIYlb1AhP30mTghrMjWCv
6CjoEAsOcGEEIm23VkpSBeqKcPXi7uAKAIO2dLjo1tGfZsD0fHeus+R1eegNZxzAuzCBaZXebiT4
L096JxpUPBNyxHwHi1jmMhK51cX89j+mFQh31zLrP658QaKHr+FmuIuNkmUOlYlGLUf6OG0O4IZc
rtTANg8KnQphgu8IazzzsX2wKy9HBWbYE/isWLMFXxLbxFvtCitCyb+QTyEG0DQ9JDzvuYZ0Cbzx
/KG4lu00xtG70gSmFxS2gTD00uM+XtT9So3a3winiKdJfQjcw/U/LZ6oAWmPjE1/57Eh0MDq7JKq
XCwwWM5RaMr+99tbJ0QyizrWaQiUjXw7pyXa0IdLMTAxGVOc8potJc/Qsk5ZY+qydUH1948X5HXy
oTxXDyf/6yePuPutNRLbZhGJiNQtngMoWYGHjOw93ExE2c8ux706/2zjm46CayipZQ3ucvZWx7u5
Zyp3mXsTLQCdbR9bPOPGnE5SQSojgDJwYQjNu5DeWz93Qnx3QTnOwptZcy0jnJZjV3mCN8HEcqrF
Nl/u+JccxLixTfDr0oYgNAwRG8J+5siTNdD4EUQ4eaCXS2oWfMoWHwGROsZz1aL68WtHWg2VK5nO
X62Gt6n7/o14WLp+tEPOmC8ygz92K4QpXLqfjevbA25mTJKSq+wSwUlJHv++LGnwen5r7odsMktW
EohohNe9kp0IBN6xyKxfYm7DHh4rjsfPXG8sjnpm3SYmVnvhuSdb1XRfK85tVixLvAvRFVyv9utu
E3nsmfhm6Ikbsav9w/NxHpQ2lZnOtmOPH9l5TzacXbeOfmd6GlENjV9hBGs9SB58+o52+KPjNHoM
MjYjhV+mVf5mqFGTlp/oaE8/60wGGucrb7ka0M7sIOBLabar8HndOFyvQQr7kfocqciD3uD7R0NJ
dpFS88u9dID8lxEGyPUq2gGwRWX6DoNr1OYf2cwLT6WBtdVFoWKIUTbNXbkxTnsq+qqD+9b4H/zL
jfnZ2PviB4CAy/YDM0rEXrlrYegDPEiqQBRba8ZqW/nwRwWnP41+6FiZUBHcZMyz0mhB0j4F1EHp
2HHwFnDuETwQ4mpOuTgBZz/uDE3pYUOXY31TBFlLJNZltf3n3BWIlRhsGe6OBXdy8fEHJ8VHfqqo
3CKSnBhpwLjr5mnHjGD3+/GCliLRZWxH0usBiq5LsMiI8cebxquLIyCkkBt++OQyg44Soh6m3bPN
2F8PRUfB3iwkJIZI2Wwrz7JhaXUjApGRMexGb/mzIkH9mfzk9oG4hEhWjLuUinH52cw7YncIOOPf
C/9XbyXVCFZLzC0EnGJ93MZxTYeRGGcSjy6EP/3xdFzPmKvSvA9M91BVLOE4xgZLbPPdhWkx0Sv7
euyx4dGErndJLGJTjdVfooiD0PEtiHiau2VDKoj1y656TQ+7TEkg5ftVILCKWMnehXICUHNzczCj
eyIWUnpHBrpHWjQqNgSHofEDYnTEpRjdBOfMhzB2Wbb5twSD95Dqu1DyiEHxwi41yFtES90jeCNm
GEq/2VhO605VgNUBGpFXTj0Qjeo4UJKZ2J8NUtRXk8K6rHPqmEM/yfaYOU6UZ2w6vDeMcoS0WhU7
Mnwk6GErCy+OajaCUH6jvapHNkHZb5WKU2BUgpKdvl1ylSFgSnwRFOZELmPH9/Uz+SUffIUDlnRv
lBlMx16t4i2jhUI7dfyr9ZITPJF9TAAhtrBX/F5+DmvQmCIgVWDu4OSkYjCez88ibwy6KTTG0Gfo
8UVj+O15UNJk4kiTybRU65Wo4qEVsAjsazzhaYLAY5hvwwi34mmcrOdis7vD0On9dvA2dcqht752
av+ifpEyy5/WFeVsrGgToVtq1fVNGvGvLdMcBNXGUZxsDEqPmsAsJDi4601cbVZIWoPpmazLMmXj
01O3M1fxI9a58PQi7/lMKzV+UeY0luFOFBud/t9jKDpkGZx9Fwl1H4Keh4BZgoCbq4CJ/Xqk4L/w
8GNmbV7qwyJKeTZ2i0+0+y2mkIIDvk8wEhMYW7gj4lyTjihsVUeDPzxWZyjFXTxVtVDoJpUAtLHe
y2Or0UGC+UGFA3Tnvtlu5uii7vQTrW6h/4gLAHCp8fdlrKRmLAdyH6HnZz/VgIOQB8tQAfZJPnjc
qt8y3m0gFlwces0nD53JYiasa8VMH66QXTr2YGjbNfrvk0vqbmG+ko1zrRtbrCSkxgxwR85oBzZw
kRMgURIE4pnXNmv9sXUMmmWIm0h/Y1/iX1c43X4PlpJawZH3jaH8liK0qWYUW73Z09o+taemJFSw
Wn0l0k/ZD6PF/06Y7G6DiS9Qv/Qe49zrcelv1TMLs5sS2VlrnVUFK+2QfE64gL3JJBhwbDNdFLf6
xGV+SYFuTKGXl0H5eVvzTup1Kg9lO6HfDtoFLcESrtwK4BzYEJvk2gKmhxGprH9k0kaJcWr//myg
0CeRL3EziPqruPykOMhkyurtwMCp2gxCi2rePmlOpsia8YP2I7yl+kC3j6y8Y1q/cR7+kIZO+2YL
4Hka/IrCJKrhN2R1SZ19t1Cm+vtQAbzJb8hq2Fjl4IGCbsksMmvd+wW4NSBvUndWV0vYdt4TaGXN
+GN7NMosPkUi4p/dGoFREYNGG5wE+8m0lCj7EuaY4oHbZ7DjaDw6xan6o/+VLww2xZuTQarVejT0
2OCUGs7AI6sDGEMVvGkBnhG/rSz9etvtoAFny7XLSKjy0H2MAixAjRwRKWVG+SqnME1DeE9j4blP
XQzgr4ghBZegK8/G6o6eL+JwqK1ctuiGvhvcoEQwJJwfbcgfk3DAqd/IlPIFQF9fk78uWKDwNI3r
LAj8VHXuepCq/RPqyEMhB1SNu9eCh/ZQmzdnT7HhsqbJdcb4MkfDjP8gIBNyaM8r8HzJ3gdsrwuW
G+eEZW3FfXNJMJs4y03JS2dSgiqub4j4inkmbskJXBA4nldghzhworwE/TiFIpMSpper3K9ezKhc
Ds1tSKlx8jUqFkK89X49ZsK/NrNL5KBy9w4fNiZarhVOYJHKtied6wuHJm5lVGI5uXBQMM0KudTi
B5y9ykzmeM7kR0NhPaA+4EjtzsbAGKBOqMwF3HZkQV+MfuKCoBFSGJXSGJI7/Kw+nkNESMMcLiWk
bD/oJ2zj/YCMLb+B/5DG8asITD6ZSUl1eCVEN4kvlwNorcFfgxw5rrL5LWZDCZGP6yf37B6kMJU/
oJgV9TidLTriSOYetDRO7PsEy1AzOv7TWA7NRf9UNe3LI6S1k81dhz7yk5o4uPKWzoqqKyaqjeEZ
mup0y347Y7LdTHDRrBcPou+cG6UAuzErAN0z27C4jK+RcTt3UTUIEE04GrIPEdJy9PVNADKPhLnu
v/V5V2MDT9S7OtbcZuulD4lUEZlxtQtlNjKPfVJW3r5/5QNA2fbXx8U7v/5WgewJdA6wI1+iR/RH
eWHX6c1JiVnBEfz/d1q8d25nxWkY4W/jGsBsBYQRtkjYkxSrbO1Hhz1Ms+Mk9Pt2vLanROhV/fXU
b2Y8uXaVr9UCe3O0eddGNuY/T2SU82mYd4wEWXDRosZ+n73zMIanHSmru/IkSsLzuMEqAdzuZPoB
oSmZ3WgvTj1imBw8lJy/WD/Guc2OmJB6kI+XzTbtDIYYyhinqGoaw7q509oxfzf1CAKqv0e/QEFI
6kE52q9YLnPiMBWumMipWGC9WNQGTL37jBFuXRLJX9ZqwZa587sAitNB9JWc0LyxGZYMdkYzF1jW
2bd6V6vB9yNKCp5ziRbJfDmEnIPJ/WHaTragO7z8e1Vc0hdbPopalA8EsJ1KHVf03YrZ6cSlpyky
72tHEPHUuAR+tuNk2ZPOg8SE/Kz22IqdZ6KIXabtJpYCNISR9drEnB1cwFXlZpnv93OpCHJz/R0i
9MGFkW+cTJocRcNPigtbYPAZ/oiDplcDbAR2lmWA30zOv46PaXfjYTwmg2bi7bax3TeIISTIW304
3xLnu7Eeg1GYkGRmn2w3K3HCsElGs1Srl+q5ezd2m90lhEF9bDPTfW1Sz6m2hHpKjqVYzHdVqudr
U2H8MieWmD9fL4bGlA4+DcwIpAhYmOlbENf5h871eAv7brLqhoqfj8xurT9FmsU/MYtSu/YLyWmk
7LiaOPbN8yeB1j7QEeNBkY1IYXq4wM9G4MiYP1gxbWzupmqEp5B3AsNWTioImlu0HzWcnOOTk9qf
5Fd0nhW8IW0E/JGwB268N263n+Gv32P1TW5KuAJi3OtOO+q0XgPe0nFyuaeGizqg0O4nteVszslG
+tiu8U96fFWDhwWclj6q9EVJYiaZPXQQdwYb+o3cbLO/zI8HjqevuEvUrlaIIzkb1592qsAVngaY
STcLOZCSVTJtt/mo7tjq0LfvykmOcVl6O+JBWyyoxiT7W5IN9ky3cqLEMqLGClbxV5gAfV+nXInN
Vdog4VYRnfoWEKfL9rr09/Uqy9P1f2FUR5yWYw2500Rh6O4Qbe8Gf1U+/zJmjbSYr54Ydhw3nuKu
Wp2Jn/qrDxBu8QRGqJ7kte+h7MSdOeKZEMy/o4HgpQkPGJU6HMfhptY4i5PpSXGr0lL578BzsN/A
uLzqS4sXxvlIUPkmuZekK4hsT/cStf30U5tn4iluFh/SkPaJqqWfMLi0nYGV8JvLvYeu6YQi8fcs
PL2PW3q+TuwOLV61ASyfXZzok/LQZMda0kA6zudnbnh7Bq7/IiWwXxLy5B9ebujPW71qMCYzQBtZ
PWGcJCGzJbX40voaCBmJxdPfJkqJZSzb8vbht+O6tX+hoHXpZKhWiyOBIZXngGoTtxhwBI0M/jCG
W3N7UkMno1Py/+jbsM2MRpq2R6j9UbATcok9A2uhPAVL3KEi1D+bw2lEphr4vCR++usjzrYNFNRl
/wiakH5btop33Gf2aRLaCaHE2a1lgiP+SC5SdaKX3wuw3EMRTbCPYRrsMoa8MHBpjHBAWGfCYeTm
IZkqdUo8uOZToO4rkg8eeNG2AMOEc8OpbRGm+Vc5/J/LnH+VDnwmp0LOh7aCZhQu4w4lDO/bUnrO
CFOmYBl90n/BX1wNoSAmM47xCOqTyUeiLpKCsshB1E1LxGGzY5rLvmsk0nkD49QclJyefn7j9QsC
zlBHlivDMLs4eepH01Rhe0tv00X/Clgw34oKRjfGissp6l75LK4/XSf654DFB26gwf2KjCMcSFR+
nslZSOhbbLlJmRdu5QZi6Pa+WyOjgD6lW3dfuQs/5clt4epgNAZ+vt8nItQoCn2Q7FJkbvGKb2jU
Nzp1iY7bUVMIjmWBJk/cg+lgGtRKyNgVtXW9HeVnKeUjWeoetRiGwDJyo8xq0OhCENUyCp0p2pSr
2fch7RmeMr5+rLGQdFAbte7fvpEqljn5+YZQuEESzvFR2naSVNPxfrIbP9tsc816yjASOnrlLccE
y8AtjFKkE+OmsnWRGNju35bZD6c2Z8XSmnepa90SM3s4ArzcuSBLWt8fvTpEtUlsaa9zSWb4qJ4E
PR0nQ/EgB7QGjHLqph5RGQEcSeoxOX44d0BWeWdobf3IJMxerJvp9ZsHH+pEQqaCchBzpF/0/0Si
xwAPFWJK4+1yfg1Sqcos6/cZnBj7EjNVHNLkUv6mIHzLfKm91vPch5WaY7ulWQsmqs8UmHaMyRHU
U4NZAXaIaAQTP6POC/urDrawUtGWiLLnF5OCUvia3YHDMMumZ2ULDQPUeJwyx3qxv2SRr87N1CCQ
1r/QPKErAKB3H85Ct+O9Jx2R6nJQnLxlCv1n2hGgXExdNyldPT6GsTjZS24bDAjdMAjtrJDzbZzY
afDggmcuLshfKT6cyzz1o9YY+6seqfh4ygLDHWfzHm7HSklgdgxCNWZzlni+mPsxTkB48i1lok+V
XEGao1Mdc39S3QZwRPrkCFo+v5TA7c6I8gnpiyvNM3lsQxaDYRUEtRKWszrJNLOwVOc2sdQK7YI5
JWa7O7xzgd4xB88XyNkb+/pIrjZCjaV4ru/LJvS4GfaPewR7emgmIllfg79EbH+pCR7kLX/vPSN5
eK+2D92RweLJUb2OxXMeDNEKVHNVM9cNWqCCFcJCI9MidPcCoQc45xiG0bIF+0TMUB/kftM+Eile
I4dG8YFPIfXtaUw5c87hH1sFCCU0H/mPy4v+0cwbYAz8vuecWRCNFfTtMmdqK6y/JpEn2zzJ4H/v
Oph2YqmNi9d6IBlZd8XkBzNszV2tiNpU66s0a4p7Ka/u/pRECjd1fuNG5OdUXPcj9lJkDs0Uqwci
cyiNyC+I4HvppBIu7LqXDN8C2kxhobjwYXgij69J4ybcb97p5QjRNi1SXjYM/dLG1GaH5rHZiN8M
JGWBC2YvYzqvUvbLVZtliBEUh8UW/fhNeX7r2V4sTLdUlY7dIs09e0c/9ZRVA6hHQF6Ecwu7wn5U
f6cl3Ezkoyr+AjA48BaV0ictzdbLpn5iuV46JGvBL980ZUpIbwezC8AkEm24PHpC2YfmEGdpWqYN
QO3rFxNcP2SrUj2mqezEQSzg+cOsqBJlU5d48WmFVP+xw9jC9d7nWjC06+eppgrjUMoRKgH2WK/l
ySeUNCtfyLobHfA2epNCXzSnuo/8gMpXSDndm1Rm9PBehg2ZQnPhSm8R5V9KndhnLVtTvdabxUJf
Z0M+osCpZN32AaNBEoNi5H27qWukEOU1eL1qg3NjoJXXLsoLWOJjXJ4tQXXilRzKZzV+iWBy8ros
eVnfPiRqIgjtwM0j6J1CbdeJj7gozxwt37WDq8HD4oFadKxGoPhlqKZP/Ze2Jdw81V8QCpBIQwLx
fn+8cq4ZHssJA+HKq8X4E0r25xbZDNgfQoHjovRRyWSiyTjTVkKYtqLyQZw8XDK2BA7okgofuf0F
xzWtNddKOuH4TeB7f5cQev+d1kh3pLxvO+xGx8Sv22zlS30guuDgztwsR7izYCYAg84YIpjfFFG4
z+5OujqHb+ocDR0OIplCVMUfS84QEI96wsAiOamcYLFGiMvWiEJePm3av549WSUJO3YkOAObNEcr
VhOkcm4h5pbTN1wTMNafPa4uDKyIb8MxQVlcVxwPjga6jeNz+vBPFPmA7roo80y+BLZrCq99h5KS
Xu5B52bEXjTgjr2cvPxASBplow6YtQpN/yQDhxYS69D6wn5jVoXcHpPfIjfV3bPj+tID5xPKUl1M
/89OKeeS8zG0LDcZdaExCl63J/0I3Qt667jE1ZiNN1nIP6x/ei6+GxGVHjMlRNGJOHtAXdPsJ5Oz
1UsphJJbo1cCTUzBS4j2z9EbuVnrOI1kop48HMfDLF+td9/L5fV56wiqsWHtzBhHnh16QyEPN6wC
Q2BO96iuhIINQV431aIYZVqW+yJlJCLPgRUrsliQVFJAqnp+V0G7DZQDcHloeDcfE1wva33+ex2W
vcqsC5UxI3g02ietteaR8z4beUnAtjpBX2vBDAjOh206m6Xt768aWedhTzyJXfT/5GzOzE4yd6Zm
AVIMrKEErkM9WA/J4u0iHasRweSIj1a+niBn/7/Z9fQlYwW+v7zlNyHlqYj9PNB91Lw2hN+Brfkc
+ZbgZ1kVJAgpbXi/S4V8MxVyE5jvZmhHe2NZIDUHcKkCRKVIfMlEIxoYD2hEQUggptru3FwHNOkb
TziKqViKAlJmkhDUL2A4+YTsP4J8yjcqPGYuvcu6lsdNbcQc67F75dQyPon/kiOMPzR81bYHwkUy
WD78Eit4xDpSzDMNao4i7kkxnHAjWY2ASZl9dLNCPCtFK09Amx+Rdyq/2aSjg9rbkdQMOexNUnyJ
4Jn+ROiUCFWHVELCKKBsOuc9USsjTSc/JQcYBPxcxZs2HgqHmkMs3ryBO99z0BpQrDu7YK9hlWoi
dyp+yMOigq+6IhPOXwKjEqrQM+StKLVcIMkVq45TO0hj2kYQaZ6PM4Mt8ZPDnPqET009B/HJPG/L
ObIMB9ss3Q8l4dcXpeMWL8QHk3uZZ5UXVM1W/XvGzTv7pj8eB0dYX8ng+iX6vPRirgdT/6p5Nyto
umJXznGMK2BrzMSG7py5DVScBi9UNCKTrUjGOYTBRzj9Olar1kNj/hEWC6Tx9Ln6Lu54Ka4zP65N
JSZMbOa5g+OvFJimZFUdPfHqe7XLDr9kgJPEqoxYBJtXT/ch8mHyg+uZUV959U0ItAdqeYf+G16T
Rggn6lB7udYRgmlZssRhuPa89tT4eQ3hbw3IPgpT1BowKzNoj8Nd8dm5/r2lwp+3HlXWrKmjzK0g
ip/HULLQ+MrLr/4lFkHz4FCWJQgHtVgvWALEqcPIARxBMF1fjLw1bwVf8jmTpjOroYjzkWcb3Wgg
Ie4Q796VWnS5TdJ3gufiOdR+BR3IXlLpbg8IYTWWgvBEuVdj9L5imY6V39Y1WD/SLmrscGexxWvn
uCH5F9ILVIVAZF9JokDPI9lIrbxJkfilXqmdKNmRwY361mzwALt6C9f6TYchtTF3OHX896LFCwHu
PHc6/os5xbbHS6J8k2xv5gjJniZvopLDcxweD0v3pFv6hydhKwLuLILXtjjkncgwKFnzMvI+hoNc
xfNVSlIyFy46TdD1cXzjed8pwqmEnL/6wJuYrSihfVtRZkn09dgHOAqjILh3V8QxjtXIx4gDhm2B
YUEd7X3ChA6+B/2gFCHTBDrJQab/nH84xcls90/PhSVysLBxggiwCcX8ANRN5rUn7QceYUw69WHq
xNT3zDgQCSQ6Rtp7GUsV9bxOiLfxJMJYxuSgAIBy018qk9xIKcFMhK3uz5utEHvzdvhPcF/V69WY
Ho1afS7sHjyiITyBK55D91/DBQ5m5nWDvi63AVRvaM0hS4gmY/UqoI674TpHKpiRYMuJ8+6PfkwQ
Tg3pzSQEhJMwGtfJ01vzwIo1F9fupdhc5JtUg8Qyr/VYyt57SsDjLYVs1D10yMZ9qcygoYs4la5f
nXB4tTcv6XjMGgVdgx8AU2wzUpah6QFgqHx9pRrc7XFD9j3UgU3FW/6SXZ/RxSRlNHYckUY1NOYp
doSQRZLq3Ll4Qva/jc/jBoO8MKLLCB5f2fUs69IKPKpBcEdSDNMPfXxaneoP4UNCAsB8xZakBF4i
o0DA/keLTd43p9YHQwXX1RdbeJ0RbVkUBQHbf/F8BDG3PWexrCiQHS9o8Edlamgm7LajOMjPQyFR
RPfDHLQjRN/B7gQKKMwaOdy5XZp4eAgisbRkzdzjsDSWYAxK5nZ16g/B2fq0EFqKYE8/cy85RNIR
Ue2N73Ki1B0IbEB6G6ckr93R3uD1Lq7Y+GuMrRPcfk8/m0jQ5PVFYpwq/gfBBvTKofh9dnSWjtUL
rtDC+xMO71b0JV8YWf6DVP0AdFZcrtherZ51wd6HG0f1OlMTezGDClKYQLDyKYcZDY1NUXnofxxY
THiPVqfb1FoG/J/ineuM5pGK9ccLzAzDvdMVytqVZV45H1dS5PKCZGxWXnOc+VPDtpC5tzLVahex
CpaSi+xfPh7pxC+0HFinJVe5nIfi/jxaBgmo/JVOkvCZRDs1b0SocqdEYgSuMQpuxV1CyN1Og7fH
RlI6s86pXQZ0hhfnY1lmZ3Jt2vNU31vSqlY7sdNbdqLDv3LGNGBj2tzQHuCah8ra44sqyUcuPWvx
zElgGBJRIC6vCJHngSyyk6Zfw4440+UTynhccwZhBIrCE1CYxyVhdc/y/+af0ufaSiT/a6++AKst
05YZ/25tfZdoZHcA/bQMViU3fml5J10XyeSQbcmd9xs5kzuf88GeQ11eiFKZstOjpEEAgK/RCsq0
E2zZf4VXU5XINa/iIpbkzCd5lkvcz4efmJnJJCbllDUlNpx0HpthywtXmFeYyzSYE9v9ILEYak2R
5BKYr/afw4WAPIuGNQ8VjlHR9OBkPbEAG+d1AT+ZA4yhBWKZ4fnlj0Xs18bpuay/2v7vuPxOUvr8
ajY7MWuMIstGm0MP87WhTqjK8SLfbShF+BDRDrAy7wja8i+i89RI1lUJHoYvcf1yWD5K3ZVI2wru
XxSIWj2Mg2hTLbwUFeMhi5UFyxEY4yZ4zMncxE4TyQloGyFD6myMtvNrwE51PuDcH0ry55TQdTlO
F1FLDMOEWpw+2D3kwOKctM/fdAzrzmU5Rkc/ga73T/vT3QhkgrLduuGKxNgGbbpfTywgJPogMgsE
vUmuRiU0ayvWFkbNBMDofuTUqxpuv1xB2GW3CLtT3TshNyZgFKrwlVn0V+YtSlHy2wB7tMJiXrcB
dR2skk9EkX0Y16x/UNzvGpbfcVgbwGEyTua22hzUT6h59Zb7sE0L9D7t9Amh56PyKyb7XljVop7H
OM8s81ox/jR/vQrvEVazrplRzD3xxarCbcVkmPLdTPsp1Yt2CaCCKjXrv7W0CZ9YDeYEnNt2gw1D
v+BTxLs7QutFmUrJRy95GnK32kZEcvyegMV/KJSdlM7SHiVWIdKd5REf3oIzSiCWflvPYWVASpPH
92YoXm6xBdX9pxY9vwF8qON6erCcgy66sO5ii12pZ/ygOHip13+VchwZKSxwp+ZtT9/2oGLO003U
Og4yBsoOROcwYTTCNUZnxitGZRafusogall6A2sGNQAKGmDc2gFKkeBMh253JB9lCKKIk0f+Lcfk
Rob9EjN0VbjqbABKIpguytkU6GIZZPjLfKvJJ2J+ZnTUX2bDykobW9bGR0QVWPqE8NGwWk0Wm5y6
fW3oM81bTZpeSoVQPgUx6I9eS8ESGpCX7NgZdTOvXLjXmpYgbrbV527/1x+XXBZLwZFbn11ZAaQ4
iGRaMlGzYDhfHhXh8y8ln2XQ9BqDqBGYDChnc/axjejyput00DDUhB8/Qd/ZHcyjPtS6BU+EPZ3w
ZFKqujI24AbLPVjhvvUO7XHgnkPW3WgDJqrGSGGnCKiHSFbmDxISDJ7v19MfqNeNAwxLm8CEb1Hx
JlPt2vWsr3ypTQdSvcSINqUvg8wioQ9aKSlnUWC8Lb+N7Wql4RXkReY5UtlsFGVjdPistECxLBsU
hr0EY8jo6MFsYBDcTAE2rGg+zqVMt78v6AhPJeVopKWVzD0Dgju5Q78fyH91ahIH29boCJIo90yc
jHW23IB6m3Ucem504OMdAnefwJqidXtR3rk8AjenvNfh/X0LURRemtD6XaDimlJjvUFC9bzdE4Fl
TL+3EwiVQL7dAZIi8FibAR/4QwPTHqCdgRodn6HN5KzPRJVFcZ7ZDU64/a5QxIfAxLUp5RGAOSmb
kxtDb/6XTbqjgoLx1Q8h+MU8OGCEk6IBsEcDxOMldwux+1/x3G7KDItMAQOwoQb0pGyjqDU0ysA9
c6/gpAyCe4/PS/w6nZcneo8F4+ytpu/u/AwRiJKeLW/anFUxzG9vP+8kr0INYlOpMZmuQd9nUIWe
40Xbm5XJbG7cl6LchrbWwBzP/2KaSuhbAqT2Bjp98iu16gZ2WKwL7l5kxUooDvYGu4fXJWa5rBoL
PxIdNVJ0rokhaS2a5GiTXV4imsmF/0NxOqTllbxjGtPHd7FTLLuc9hDKn4jZjFp+YXUWBwnTXhfF
RgH7hB9ds90yCWMIAjFbSI0/2lDzVzeDCYNdOZgKvG2rzZzdUX3sBnWEa3/joK0mgS3undIBczz9
oCpO5tpYBxaWWaMJqKYsxpvCYVHuzkRUX/tIJy1eyr+M6sgt/zNieHS/sU8zVHQ1jZVxyF2/MhfM
GODogwhYiH6okJ3VHASA1oRXP3Lt3XdY653Jb+lA/sP0domNeoL4IHsOUr7b0Fee2QGHKU/ef+D0
1j9d/SDam1Gf+KNlECtppR8qfmad35kbAYXXdmJ1j3l4AlCe00riEo20TXYnbrirAhSddwKAB4fW
xpKScwAerLFDH2tfu0zvQ/4WyScgVg4z07LCXU3tb6Vk4msxXF7AlRR0Xda9G3ZcF/Ucor7SaXhL
geBG/sLmdMK+AofjXRWZV7ew/6cWVUX/+Os4be14RoJk6R0FyIltZtT/hd61ij5Pt7U1nqEvAmjP
6tZhJRCrenBjnacI7C+v165Hk7toJQEp00ct6veA1HFT0BEbVHXB65woGWAP8r9n3noisgpLAbiC
cqacJbmW5XGL+w85/uwBX4S8hM9k/OdAfxTWOere1HdDAfjPK4oQjgcp0NdXUIIwdvK1ly5gvrnC
lCs70rHGZ5XwyALytzmbpGl36Dwo4zOreUPlTMobPssXCD9Kstury2UP9Tx2SktQiEs1BiCQ7f+j
i+jFi9jNr2/1gRMDKpo/PTfywCXYq7fhEZVevJGKjnskb847EmDi0G2ldzCyhivcHVncbngmvYlG
/+2/PusneFSfUoXEGf+BDDMDYVvkCz6bq4efGA9tL4yOJjhOgPRDe5Uy9J1Y9JyboYXWPR9isash
WKumX/IcE+2D0luveLbH2O+yG6FCtBPDeBvVFx6BhPJ3czqc/M6hW0raGJSzbNQh0X7rV7kaZ5vZ
2dpoYeexvfwZ4lkyS8ngMugxeQif2agIdkV1U/ib/OhvUOFFRXxVJD6+rqm4fsz+s+E9llP8BIc0
V49vY+19mgWc7ZIhpG1Icn6R5kDTvKrPqtzgjb63bxLUKlPXmbh7L4LkiHzEtv5pKboFUNACT9o8
6Mgjh1vX6Tn+E/LneJwzENRHfVTy5+gsvO4sYAdSAMKysKRc9WWVPYctaMx5CUSybAP6NLKxTufa
bqtdjwKoFDgnowfKOE7iMYVfXuwXNqiFxvbML08pytRfzI/gz6P45EjQx2wsp2v3OPTySBUwlyvi
AMTSQpr1zC4ix9IfOkBUgn8kWqEODUKoBvA37ohgbFefo6k7Y1oQLWYOHucQYfX6seR8vzWooz/K
vzqYh2/Y3u9EPMz9ezdvIqFMUwJFLR9ELImjOrTi9N0lOjGzIlQqDt5jwmojUbjbg2LJEsc9q78m
3zCEt7KIByLTJNAnB3qztsNACV7lwV2dF77TvEnrbN1SvwJSed8NHi899CrrFe+oOPGLarMfa9xY
LUFVJ/xbYnNnITxAllqqX1eEsPCMTxL/jhe63TI2re5mvqTfRuqTiiA07kGIpoiIBKe2xttFPxH4
p+kAnjUVWQWhkfGWgsWGW6DQJuiGHNhFskb9Z02oke58DuEd5DvQt0+WiEs5w5brHdwikvQOCKrW
f2aIg9wGZchdSH3RKZj0UNXBiMfYij5k0zOlOxrg/UGnESxJzI4NV3sPe9jmgCV3HkQWvwp+/AZx
i4e9ToDhR+T+EZ4qWPdjDHzf9EnQtTOzbsZq9Hai/ZoHTjyrazh0BVJay8cUb+WjSXGK+RNo1Ed6
qx6rw0ah+RRy59IAmOETQRlHFQlpJAKU3PxuUwmLqR+btUy4dAqkBRaDjnY88sFv12oMbZyaZt9f
leedZ/+DFU0EocLcQg2s/2Br+j3nG3PklCUeV7pzDwJ4JPYWYGYuYxMOjIsUmv8Y5DieJtB9/Szq
jP9XVNNUOWhLMVdbyrxjv0stXmCsoOJHw5mF8bqyVEc0w+wzX6j4z73vO+SLwpwGcgcDNoOPesNa
EkyDRxjum1C8kHbW7l0Oyc9ZwAXBl252YNclW33dAnKPOLvng95qXhDcWCSJMULHWtJh8rt53mDn
Yrw3yogLuuBlgWWhkLHNiEIxQDFhk3+ZLQMXDAVmxRDnHCKLjqWOl6z9KPO4CK9I9ZPQfwGkAWSP
bH6ub3C1xfFIxV3qylVd45aXgGhiLm69rt6UEt08VYDkcWDw6ysT8TGBl3Z9claZQEagydaE55yO
E+vpe1dlEdA+zYI0sdy9kv0ArnPXdKW/q9BsA1icuw5G1nSNq8VOrRMEEM9x0hxtinK+u9PNvFIu
yI0sd3B+Sl2o2mzeKd26aCS2w0jzaR3nZdl/wNzZ7UsunWDl+DkiPGYsU4lXoNjKfXFKn448SgnY
SHiJ/beFsy58nMDZbl+c7r3BveDYW493J02xiLY0l4oT7CY00+aJnTXj0s3CexJChZLcDmtle/pW
WmCvzbWgsBWhbDd1dHA+K5lrSInUE2WCAW4ClaMKTXkDUNZZjj6JikuHTH9JgmxZvRKUbbJruQsd
aOaTAb8SdAIYrMkASubhpzwjGlJC5NR8dxfeZmTaoh356762POihTOfUI+jEgLocYaPTyGE9QsTK
DEsumcESnrlkieQ3fN1jtYdrvGMiktJdk0K+c2kqj+xvczFqlgrR+PzYO33aavnPEDpkena13Squ
xoWjJndDvEtJ0SequbLPDMgeit94PwIAjleEfz5zAyReh0S1EjUCBzbE4Xoh3lcaJPCazVgBXDZ4
g/jEXuss5BkPCfpvIWu6TjdRQX9lue9+mWG4Q2cyTlezF0epuveexxntCvQ57cjYUa258BHB1Gty
bGw9gRXUNc9KiKuqiWzN1PgG54jr8RCNIKmRSBNbXc3Wv3MNhtcQHkhZhN0EqwzfWRpW0JRLAgp0
jhrCfqG8T9Kz8TIcPQRO9DwVUt1Si84o1bS+8aNlQNcwPW1GZNLVh8KjqrTYXN7EAZZQA8rJBKGI
VosWK87jA3hRrlgQcbAzZsHKP7J1w8gC7qeaNrB1eXiOskVzqyGsAeGHxmXVTY9UFKsJPwo7GtL1
hidBLE/8GDgSnEsYQtl7o5qGQpY/A8zLUVjQCXMKJLGyAlVEsn0H3eKC8JiMXdMIqLG2QYIPdEIp
p7olh+dSaOFiWhOMjVyn82h8u2Fv/lZLJTNrxGlnB7JihPmtiDBplTgiiZGE4+GIuh65mBula6wC
ZTcw2uFUxUtQwVARltieakBNPDuAgNuxQbSjT4bwp3QjmZxYn/WJHFmPvK0bSfkci79W9cleK13c
76K1KocnUnuJjQaG9OKJ4p8XAXLAUsfJdc9OXqcutoQggkE9MuNvIABLJmc0uvVtE3nh/XYKYmLQ
RREWVCsNYp4iOJW8nEXU0hshHsecVAp6rh4USr5y7WYvyLsRrSQ57AwbCIixR5v9lICRRUVOrgdk
8Kp+GSJxJIVkS1My4gukdq6WQkA1djNV1QjC2iF3CUvUUtydk7AcuPj8JeDeB+tAxGKPI1IEK85l
+DWfQDb/pv54MYKZzZ0BhvzpB48cb4uWPFS4sOks3OmmWO45zOyLJehg6cpIzdIPrCte+OUsWtv6
bkJ/CmfWtPlRdwj63U29oj/jtacMSkG1IkC/4ye06lxhLz+38nrhh4l6MUowgB25RVByk5MtuIMT
rdEYUOVzeJiIUef6U8TTZU5nzchOsHZZRzrXj1qsu7AKAWpz21mLVzOo1HjDUbCJmFkZOhUe50de
loliRGK6rWY1CollS/gn3ia3IN1/t9n+9+XNX4hsXiRBQT6us2xWEIP/1xBhEyG3yV4SyJaPPXDj
JGdyHvScI1FxShKHdmE7ThtV9mBOf7WRPDZcNe3iKQV9ZkH7HNIeRyXXzu8dXa+iBNMEMSbn5cun
9z7IGyNDXCOgVVDMXPwVjr/P9llueB3N+ITffeJsDCuaXDCkWY6lVyGwuifIBObCMQ0hAdTgk6vF
9fwgLkdCdI6Qm+D3dNTXePpBmc8QAubjzZLbybC7SWIszHQHRGtJTdKW9ea3HqBfRXe6nRhTAOXo
XaMhwPZqvPbju/0Yl6BfpGbkGwffuxZLdzOP1ZnfKaxXZ+quvvxSApRWmlzYiDjftk03iX/qYTis
4D38VgZZudxqqGEmvjdxD9q9V4TBkkjBgL6Lf8L4310i9jC7lS9KSNPK41lmIQ4Ngdx7tHX3XFu0
68WIEkFZmYLqSuDT68oF+uk3ZVlIANmwzB9h0ID+iCgvVjWgeKm/TI7fJQviEX1DTltPULuJYo3r
6Bj55VsKbvvNl8uRZHK/hNtjFjXn3BpMDjLshUuQ+1jcFdQoIAdZz0jrTLGk6JbHdSKtyR8nh9/U
exdnQj9Czx3n2LXDzcKalEKz6ZynWCv7GNJetXCFEot7cqM4NJi6wgG9OVEoi9Be1VZvyrgMnQJX
V9kHMceNyfrkEeDRfsi4x8XwlQpoHhXxefwdMemkzfiOb2kWszZT0oErmiV8TP+ivTaIcAP7yhC3
us7H92j85D0bTj1V6GX6FZiBa3AgSMotoE9T8CGWRsaKU1KDh6Caddpn2l7PFDoJid+Twz/d09WC
gBvLJBXyJxscY4kutrlr/uHMbGd83rNxtczodMD9jzSlwYxLZkF7qdHt9HV6KT5Jk8YFPdmzl+8s
AhZY8De4c6TR9xx3nHxqQLk15Han8v6/JMFD3ACvRFGoay4u0mmykaz/6jcOKVbshXDF9fQk0nv5
0Rm5yzuLvj87W/9c1Je2iEIyxDnd0UpeCWcTtD1PbsjXs5/nz49PcM6hD08GMyLBdRmq0qxvG+Y8
o3fLzX+DALQ0kGMGpwik59RN/6wuIKhSzC8B3px5t0MwflkRMPg/Z/H/aCLbae9HEV8bAezCvCL8
K++3F5Ru+SHHVGOP6Ia9U8u+tPXcs4QBMJ/E8ddp6/z+sWN1K8iwCXUqAeMJPXx/9fIKtMswXRgM
4ViKWab13j+Mejdnyz+S/2qQ8SFI3P1Km+xzdmnMbDz3uZ2p4W2mXRp/Rios6S9/3uh7fJGbvbjq
XmwKJCmhByqXwRGAARvC7HXM7GHEITr4K2293Pwa/lTplp5kZKESP4hRwsZpxdD48Pb4mkROd6jk
qDVRoLMDGb259zXgvn9WvCj4WscLgdo6+VxJHJ7BnW8DvMzT6yBfHBBL8eA6qzIeegaR+8ppsQ6b
sNdNNRwZYULEbRkK18V059zmkVnMtu+ixwodj+YwwV++9BYeG7rhf/FeHV4zJwYX8+9Z7l38fQcO
jU6nGGwAVcQ8Zajbm42l3avdFUleVkUDsSm3A9z02GTCoUkgfPM2Lavd8ErCRA8SnII0z/KSIpdO
2hTB1L99qI+SntxmS4c7Ml6JUf+930hgKn8NPs+1PYSM15AuwZmeWbibQB6rYTJc9oDgcwyTYfJV
FEU8b5HHp4B4ljKaCK3wxFkqc6kHIPyGGt3y5pouQ3OfbaZADF2GwZhi9yRU+XQOP54dnvsReKwV
fXUnqJZg/g/DZsRLEhaqXZNbsiOlX3BnJJSscCqAnpkkJc0fY6HO9NyL/J0tV7Pq6nu1JCP75FkW
VAnTSqCkuANPdllUC9aCHRckl7NAv+P57psjKHUugL98yPr5etPADMdWIEb6+BUo6UEnXVrpLP3O
ApgC0reqQxHSG5j4vOtyrM2kM6m520lmUtzZiv0C85YceCJOXQsxOBTmo6Ti242DIiNLd3bq8yXI
5VlhEYYL8rWq+RW8zSA85O2L/dU/TJZ0fPH2r1rA1D3TkzXQmL5EYymjTHRsnE1cJorVCYRiWmQD
ySGO/5ukTnO3sWOT3qor7GVXA1jyfJxXcxIrg1eW62L6lt9ii1YN6R7LayXSY+zBzKCSC8V4mcwL
QvcYFPiCpCifDUaS9kup9AsovNvmWTcvuvRUJGJB7VRTZx1SxO58LYLoTGh9PV7Psvyhw/GXYIhF
JDvISBaBJSJVjlUcILTCTmkCjoBMItx+aF9xRFG2iArgLaXNEneJcgd74oB8mw9riQNxobgxBe07
guxW7+d/+aQCuaQ6NUHvuPVb0c4Ul9OTgJnC8g90o6TWRNXhcVhy1uV3XCjrP7u+ONygESY7o3gF
R5Fhbr727zb1baKSM3QvYsCy/DizZbsRzSd/bviG3qX0jXMO4P0Q0YKAF/FhsoxMYxM+KmbliQo3
ejGmH1CVAdMYh/9dRFX1V5LGjr9sCjdmnCjXYZVp1QvIy9746vUkWJXVgNb8azTMwVdfAsQ5EQd+
2MwF3aJ/1MvRxbJFDudfD9tcUQrdwaTScx4n1qa/AHwyZdKUfThMwKXMAoTuQs1XaJf5ReUx7taJ
XDZKHOP2tBBU20euJLSnyTqzsTeWi9HI1dNL2481VbtCTsklLSku9qcLX9B6ZCqCX3bhHNPIdyjq
9Og2VKs8euqb6qrm2/+/DTlvyB/zju2hqL0pV+oFiiTo98W/b2nUL4ehhBlonEJXHBSQuIWmdnxk
sFZfJza0eKujjfXw936GWYF/kgWE8jYgiPpiRZY4iR0LcWauRlnLtGl4uv2vErjdk1GJNdCynVyY
w32LcyP8e/Lz6kpVnkWc46s0j7u4XzLLLz8hFQc8GyHxXxIAS5zGJdRjaFbpu6PFje/786dWaeBk
v7ighrtHMc9HKV8alwuJ8a+sMPRHFDnbT17TKpkSdDciY+1uPRa0YM8pHsZfEykQraVjnEqsQWdS
5a5RidhpK+4cgPd4oDlJvZE+Ylzlt/nS+l4jXBXLXgItpwBOG58xeCywEdgUpailE3KPKZGkxk6o
5ItA1/V3EwDUFUBr8ZfA58j3tXxeNHZC0tOQytStelKwRqe348KfAnByDgXydptDMLnRB23GirFg
uHd12ow/6odJTVjexNMb1FmtUxJegi2X5xAuf9x3UwFAHQJo7kfxqgGkNn4qKybqTp4Lkl+e7w+C
RXG0ZVmwQyGR06oLqAKmW3GUCuwXYRjX9k1D4Ge7hpwW8SCN2wFAfI2f6JO1987WcXmtjR4o16Dw
i5MvvXRHJMmEeRjQR8fGwV4BDCAlcXAhEVbjjDCd+ErT3/Si83QrhVmqMfLtNW79Jpnl3GXwbtZt
dqQhR1GhyW6jyzMGKBbnaXyTBMrPrhWdGabtc+HCuLJEuXGcg71gULthrFT3jtsE+75MlJ135rk+
aqgg2ZyXghZmCNw/rZZFiehSGfHvAkZgVUGgBhEgxF/1rS3EkkI2pNynYeUc98BL5K3TaNl9Iqi8
tryWX5ptjnwyO3humlQ8LpxhtTO8xecaRyOi17pfAqUOXzTp4gquDPz4DD1MCyDr8IvicM6b7XRb
tGUP747jiMU1EHkP93a/yulrvHaFSy+Enky8tDgmfTvNs+2zJ/YF3ppeOSWbIZBSpSdNZTQGiIQY
be5cYpCST5yUZgGowaisnmtztOe3AaJEnj7yru9MzT3K6HE487YLjvBUsLfi5PJIZFT80AXInv+W
sN4rrCy/l1KhyG2keag3XkgJSJFKmC5ZmKICdPrIAWvHgtuTvrdxrATHGHCPfDxRQFVy4CEMSDOr
rMBFxttMgxHzoMXD5c4wRyZNgn6rbqKvWqSTbu3/sLUCEgzu4wiZM3TMspKYyqRWrmG8E4mw5JpL
wAgGfOHRwNfrtZRlmLyV7Y6LGYlgjW/KbxvTPctG2P4ETqY2oivAFX8Tv2U3xBvoZiHZLFJXswpI
b9MIaUcAY7MS7feLLxzD+mjZFzk4fHpFBVbo25wTH+a109t7Rv9jOYzKIzsEMsb+PkR8h/fuREgH
RSN3t1BxUAwgXtoldP53Lk2eldRl7jhlUAJeZcaDVUMdDtRQssg5R+yiAkiUb4wM8uJ7BdypfxM/
W8l2FvzNkwyOqe9pzVgcPbHL72lWJTHJojNOO0unwNfJgsbkuG9gmMK9xDh7eKEsU84ihRmsFsxP
7R9Vu5ra+5/VkLJ0QQEw5ikXsLsBiWsxaZPU5uMQPYqcAONtd5NbEUL+nWJitej6nEfgrVvuwtqM
wi6RMkGBr+JFO74Zwj97RHh9uvPxEMtevwy0U1VmLghiFHrciK+ogFBg5jcYaK33/+94Rf0s8RWk
JMX7ZplizORKgLTo1fohl3kGcBtJA3RLrtO+FQ2o1uNajtvLH/AIJd9AWtCkjkRH9tc/iovgaA2K
Z5e77sebwljaoZ2xy62bBPcg/+F4Wmb4QkYqzDf083uEq31j+QDOKPrWa378RUatogn6M9aGJlti
q6AtXOVOc7yWPFK3ceIAxD26zlXhY0azGQagz1feHaRsp8wmeE6Ug+gurqXPFzsRxNiYfaYWeljW
GAat5m56cUqhLMHjguiqYdUoZDrbGIsUiMxDDlIfTiKPBpwBWNP4fDo+84xt9om92IdjqFcmqIJ4
SkhPj3EQfZGPyNWHvPMT8q2KudD1y5uhlEwaq4pO0dqK7yz9NVOb3URvWhDRPRCQ3qy0IA8uf3B0
67NbQnC0dzGgxI710vwXzl1haPW9cdRLBDqh11vH5MM4HfVTOEp/Bi+ql0TZB4ameS+eU5byRCC2
4AVTUoZBq8RRAeeDfq52SHupmUoZbl0xgHSihUVC0pf0XYHnZGg3m7E4tqIwRcnwNzykBTOfqBsE
iEid9QXjsu8HN2jAa4dDSwrnwpcBGRDIMCXQzOUH8d/Glkjc5hyItg2nJ72gA86YdqHj200P+u9S
/lnRkTjzLWnprPbJCErKOx/tTdCD23Mpw/eS0xuNbZQsHTIj47pULdc77dEqC5AKBD/PLhtVzy8x
807PJnG7OlY3vEe9egk3QZ7WxgfheHsKODqYVXCy6/+Li5pK3wDTjQdKFQHl3Ej+TQ2FmbB2FZtf
zVFxWclNVyhf569xKhfNUf/3PDXInOPWTSGb+1qNWQdXYlRs6ukFEZVk0HKcjqSJ0/GjFEl1YTar
akeGYDB5dWjWP5B/CBXBsZH7a13+eiEqRAgfgyTDVNMN50HLMS/3bDm8wEcJsqt6bf4tzcQUCFC+
zC2+YNbzSwUj/U8/xjz9tZGcchry2Tidh6CXhKhyOGkhISa/U2cccq2IUmGklD6S4g2PWQ8Rml9/
mgiFO+hVoZDak2t3sMEDmu4bxq05f/I+SzAMq7tX0gIJFjKHU6Ry7JztQZJzcA7X6hVISOgRt4n4
KgPhp6UKoJDULBPgnVFGsY8DTgUxcIf40EEmS/fnoPPht7O4skppiSYJtIhYOcdEU/isCVqqvWhU
ZVTVivr7ieLZrhmuEcUOWGhUBACVOYi+TckkVT0K6d8j7RX8FDcBhs2eNU25ynjOrPtJtdyaAjow
aHg0t9ogTRUFECaHvfa+l5bEJPbmEeT3tSxUqMymTcv/vykUFf5UbPhGepN1TidGnHYaCabZynGK
lLI+04qecALbVz1vfM/TwOAjxjhie8I4FVsYzuZzFnBj94tSu+8CL7P8NdJ8qLQeZa8ZfiJCJQn3
B7IVjRnNH9VDR1AmKUWFRU9dgu/yBaEuyenA/333+ebsLlHE2kPOpm0+Z3R3fTju6G0xalb7wa6j
oG0+KbzLtSdAde+tWII5ctyrNK1HGoyLduC7q0dpevVDavpOGqBoqtLX+aCqAOKobNt0p+owm4KT
Ctbh/zSlE8mik5BpedILm7NYBOSolotontlj0gniy0Do7kyflM3GFDeAET2/Kl1hX1d5CzK2TTtB
6HTSCnrf35J0Q5yj3Ojo7dwXq6ZMvAKbHQWsOeVC6XvB4vUjiCX/jb+usNdadXQ96fjxIZ18rKFG
73v/NlpW51iU731Q/90Iqkwp40tnAFbuhV60Ty6/M97BZiGrDjZrMi96jYVFZibR/AK2TKRNxg26
64hUSk4HlmL0CmouQnEyb2K5Jreu8N6Ugk3PXEWLgI5Hyrg7F02mavyssJwYQxeE/pnLeqsjzyHd
dymQcSsTLms+q4uh0iHiD+3nOJMk7YBS3zy5DES6fnXFrBlulnVLoALvx7gQ5PSlALhAxyk5b+15
sS+6Ffz/8btapfcK1tFwtTijXp+h7qW/NknPEP0JTvIwOPJVKbTbhobgOLBGWjXsyQjsa8AAKl9o
XmSd08GgELYB7XJjS/Mkr+UOQ2Y4BBT6h6VHVqPS+pY3VchPkxFNCGtlENh1J26xd7TyTrueNPRW
uOsVVBlHKXXeAF8CHWryHy1AAVai9SK5EORJ4pInxLbC2tlZjh/kpkOOXqglGxhXBpsAXjr5edJv
Nr1ObvJqeOpJXUx4MdyseUwzlGdvl6Jd6z0aj4zI7Ga8FV/ObW/DJqc2FFFAN29YdW58TnTKs8+w
L83jn1YY83phPL/ISOj5d8P+jxjC+U+1FUV47ftebPBrq3+370RZscmhLMmJ46A0i6jfMdq7qx5+
5UrAIr7M++V0fiFDcuBxBDz0V5lr6JehJCBvWZNyVAqwx8r6Q1DAW90rRp2k8kVLUSfDBzrnDtkp
jWn3D13LTQEpj1EvpWL+uu7DbnTH0Sft3rqbPC3OYToIx+NFBNaB2yTmTSwTCRe9f+4gbvgssxdk
JkYg5+1QbqjQz+PJ1JkkLU5euad+tHnf1JxZJLoO+yjQFb4qNhY6T1aDgCefsFUdP501KlH0YixN
zrYiDLhYmFX3D6wNXAxQGj/x/m/tQlQbSqBDobt/N3BRrGD0gPIxSPUepROsy8AHk1dPlvfbqHwF
P+kefB22O01cyYnVvfooEnIHAs+XwyD5WogA95Vpb2l8TdDMmqGALR1ahVReIE20LLDQ+KM0i+FY
qzCvkWon1IaOhLlrQfCqXw0WAk00nIrz5QaGGm4rl6PDhlUodeddJYq/BQROwFSihSvGG3UKjt1n
7hH/qLWziiQsdyPwKUV6Nt2TDCeKc7mvgmf3FC/cBpoTBzcyXjJM4IAB9CkGA6OpHzHoomS4v2TQ
L2VNClodIjN8LwTZgy3Jw+XStZSxHtkZmZUrpbrOS/4CAL9RI0Tni0q+YON69G6UzCkDDZHkTbA8
ZNEvqz3SJ4+cWNei79ckt01BHFZLekdIoLSBdozkoiCq64vI+Pay7Nt/c6L/UbFabCUwVYvXxpDv
RXtp1JYI7CqpFFcmN3q0X/8qrA0ZdqNl1CELosAcqT+f8lTeChbpPrTJWeekngDAaAu9dfNe/IZ8
swGx65zBeSIQJqu2ih4AXRUnKVdf3nHzjVtWZmJCA+hZ3zNXS8n2UGzB5G7YjKs7Z+hdWAkvF7F0
T+Q0ObOUAimseV54nY4SbeNbD1bf+C3t/8J4g19mi3boENW0L2Dg/mV3m4/rvQZ1ImUtg6PWKdP9
zM5FYvnMOpP3odnWSUCEGWcnV7v8I4VYyp8ExY4qrk3nFa2gBR3Wbh6knBNQUMZ/iwSptxDjaIeJ
kNRhrpaqgrfZaDDzAPIJdnFR+0JsT8hq35+e6Q0Mnz/0f7G0q7fCpW6e+Q2MMURSH21zc0z5DlVL
ChAGz90J5UCAjGiPlnfvuF1PpxMhaWlHTVtWePAIemFWLrxv+WXwvqABE9fMaFFHwnXC0quWDxmg
qfqbxmw4193YYYolzCw+52aGpg7OinkBU4NF0Mv785lOfksP1qU19540xaHdICCk4oMkbZpZgMj1
I9LpcjtfqQVGGlVaoQypuT731CMTLOAtXeej+HvtHSKGqqWNMmewfj/zBACSXmyW3UNjfXCqgPi1
6gT3IchIwc3dqwBJyLTjv98zTob0oImZA0GXH0d+iWnntVo8H3NIXG/wehHwE1oYmArJlid9z7Sz
6MREelJf8hP2VyL7SM2Z9SZ6z66xvf81VPiPQyD/L0mVOQfMJk5/h4pzBfi/eaMNebKwlCBC24lt
05iV6VF16RwokFpP5BW9JcCe2+YwdsUGnkG1tVwCau1UF7TNDRsROt/wO2RQob8As529yylwIhWa
dfAR/8at+m6/HRNVA/vMaO8eD3vVz8JDYMuz8gPdWAKnyQ87A8VZXS0J88p9PvGl3h1fEsTUdV8N
Nh3+MQ9WXoLjGEi5k8Sm3L1+/2qnZKdOF2fL2SSeOD2kXCPvlYsQIxFSB1xQLmExQGy1JPN7LqU1
75+CDon036hY7phMd2QOcBCwP1CTam5AMeNkIIniAEIo+aHqDG4+UAYWk1x4haLcQ87qd3fC3vWM
XATESnVSB2gl/skuT0ldcK1456OZoEb2KJKeGOfzGOYeHkLAE1KZhxvdQDXkf35HOSFNLvboodJd
YcG0rsqC6oxIZ4/pfp+fBP1cVkHhDAtzu+xtVyazy/Uy9xqJAmcc9IWhpzq7kJSYeXO3kI2MrN/d
a1Nj8DIR7Mt2P5U4oca/cFTGLF3IsMsGKlqXiVipUbO6hW5pWt6ufwvtl7pUix6jdGOmfG1iXZtZ
D7I+j78Kb3TcREhnT2D8/djslFoE9gvbqO2ubQMlnKto7hEW3EnX6GYOAHkB6yeCTbuaHe1AUM7w
oBBskqkQgs3P2W/VDS/F2pDiSgaZYkb9IyuaApi8y6VzMT4q77Jr6LeMTQcAMa2+kFfWVti5w01D
wSWn/C89mK6Gis3xilyjq71wlZE/GKFZiZ/9GBNqsrjPXW+SjufvmB6eCY2SkGVzWBLT4jMS6uJC
PzYIdBi7Z1fdz3xdlzkLjKDKvxW3GawzCrVTC8ZeVbvU3DbG9H/Mm5oWLLv3REJ14FlVbbCktEEa
a+efT1MhVDo9JSuEEa+thjpVxCQNZey7vtpKsVFb1GvfiCHVcoVt/cf71egyvvRoHgngjPjZ1JuC
meGgInqO1ODCMeUEVpgcR8P+djJxBdSxfpctOiqoRmdMxPgoTS344LTthjr5Ggg8MBtvv2yO4cdU
5dCh1GEEtTEGM29fl8NUHjeuI53OoHhUzbmDrg1ICkPE2YZdrpHjhW+/axLo4fpJeqaiV57EuttN
50Ez5jfaCKSOgXLtHpWRf4wAmk21WlGkRdQBtl3xRC89ydwelko5BPGt3/EYAorqc1vKoeWvdeGE
bs9KuvjSQltrcE6JCdvOqRF3KmfZGV8TXGC5zufETiViECryyzDPj8uuaF9vpGgvoL4G0WxUlYxK
Phpphc6DJtYSyZPxNNFQ0OZKtcEJEHBPbEJOuhEz868bc4G5MMEvT83JAB16xfU5XMFH8YN8fCbQ
a7+Q5znwiteQUcHkXynJNXN/jO8Dw0A543UiP+pvwL/LUlWH9JmIsSwSBG2kj+cK5kFEAymIIINx
zD1Zdt+CcFPI2but92kj/xwwBrWiNyRfcmPd6LO42uv7Hr2Y5hzSHTx8KFnp89x6WPldoyea6F4Y
Lqedzj7YX6Ia2ghNdzGFKMi2NEuFanZfWbOqs8kbVnYXynxlYeNsjDLPbYNEIkx7tgwJgbOPd0a4
6W7LI5usWL3DOmh4FwsEyBrxwewBuDkgMynw5cOnDOKUIdArx6BiA8pTUz5vMZqELMr+ftUGziBH
+0OthLHwag2QmHPRSxvR5FxifLzDVsEbWGaGMKM8o4kN4AWos7TFU0F5KDeUJLYwDlA4JzTOoIFD
oe9aJy/5Qq+YQ+G5I14yNCLhly5JjlsrYs5ZeSSswznOMZ4P577xnru4Xe3nDVGrb+pYipsijYzC
njEmjEBP9VL6OdiWODP3xitKH9nVj7oe230thfaeqYTgkotqAQGoJZU3GsZtjjmlj3vMgeIsUvxS
2av/uz1JhYwqWKUgolNCzkzojE3PJoDElTY51LmlQ0VKLdhPARrtxxZXNVLJkFt73mpeohjEgdLt
qby03A7dEQBVkzJUouZyCkTS3wUtM0Ks5g2RkNUgq1y1TsgEhkLuiSRqPmDmczmaUjpKzzbUU1yS
G8eSGNRpF07iMH/ffwiB+3PpVaJkpFD2wMZUpmcDt3z+zeExf9BSjH4DwRa+Y4LCI2jYR4vr1xGj
IDkxTDlmsBnydIxJ4N6aqAt5+DkARMNilEidj7QSkPJDObrvwEquL1QDgIzwLXUEUb6irCVMWmGp
KInjvc97GF5iB8fbSMPFnXWRGktkHudRiobtGeJt0HuCcCJpPHiBAq/3osn1mL0TA22OsXBC0NMf
OogDPw9NkMsixlY5ApPwCok2UQ/ZLUkkaYJMhKf6VGsfn/+hUN3f3zzJzu9pC2s8AwoDGhSmsEmT
E0OSZNg8Kog8mqT1HtzVIuFz0NGZde8HdOtr94qjA22wHz7xQS6DmN6kgW1vcHj/TGlkfpY3g8Hl
sleMCamNPOcTpJ2Apk5PxZQD7P/zD3LYt1RolehoA2Fuzlfx5u/zd8ebr4MN6fO7sCVIw5T5DdGK
UMVbjsFzB5BO/+zf0+NLx4JWEeeYCHwvOI+Y/M2t2OVs55t/4FfwsY+pooIgC2hxjWw5xnx4Ru6t
Q7ZPSniwxF8YwG2eJEo+wMi+/XFJq4CHgkvcYTJZcWxtIZDAFZYXc2E36cwF8GPYDjvgLr05ncG9
08qNMN/COPWKqALn4uCvQh0FtbNwcTtIySAbZW0Sk8MDxfweA7KXW6EduYGCcNEnBvNJ3G8DYpPs
0LU3p5zKGBOdm2e6Qae+EFqAo/OHdeK4aWiE3g6z7EQpOPcOkEUM3lR+oivYnjrY7eqcFPnTCLYd
BXW62rOo3O9DWGpwggqBDZwv1A9HbSCwB1Czva+DjUOcohxHBeCcG/OTld6u0MP+ZpLL3ZhSPXM5
zLplLCcAsVMpn+ov2gAR1zmsfveb7dTJyVpZuGFUNVQHfy7OPPUXYv1b3pN1eKO+6bEv5XC1dXHy
xlANWw/YeFnzRYAdD0Bg6y2fy8+uj7lnY4hW37qp7t1rCuP64Ytej1MBc2qLm06RTjWKGfHk5jK8
BMGczc5FuhrZ4mynOk4vkYrGcvFwB1GV4ILgxJpGLoo309aSF+Of1zZnQ1HJsmDEHu+OHagG8olu
AdTrAAT0iZ5/wuIswHjRRZZw91kPtLAUZBZhNCcUGDUjxSoGZ4hs0/ldZT/9anpktsxI6kraELik
Fo/r/S7KB0eSPQ8z/0tWLFLSHRfrb/tIBrvsog72x1ZcgTw1qzIAEK752V4hOyFB2tA2RlAzfmQb
HBNxcng8YmCa1eDnOJ5CnGjUiB4HyXOt6PzW+Rt4LgOc9lifaFIYXdWXnvIHuQ4Zm9b1pKUQS8X2
n/RdfnaKO4rAGnDkIGjVhBWmHzuC2MRTBFnl5vZC9Kjm1ruYXUIh45PCd/YwrPmjccu2kMiCmFF2
ZFnHilWM7/52RxQ7BW3+S0i3/flgyrDM9pBrjwbXK39uY77i0hVAOKhJ6nBGORa7V6HMOawPm0dW
VFFYk9eXFhtZca/yFO2NldXMUsyVyMrRjHwhjAwFUYaRiZMkcf6D0azAFtqfkUyxoFgkV4h3VGMN
ptvztGc5aXLP7mGKkJE5N1t8H3A5KqP0lG3qt/2rIi3VMh9gh8CTSkuE6El8ELTetHuTkQLWDW9+
7acDuM3lD98lik/yyhGEPJYgJ9NvYqHwLO24LDS3aCyxd1NkLif0EeaR0YLmLT1+S1vn5f3Duci3
QPZgR4S9W7cHQqdalnvvmnBu+RgDrb6GV9UqiVfdiPa3J01LXEbAGsXgGRlhX3Ka+YGckeFfcbEp
iWOXFu13dW3m/0TgYNAORF8bLM8fKkUffm4Jj5wyNGhjXvaDgbi/iAjgEbfBS8ieIYIrDT45FQg5
Y2jTEPAj/oC1wGlfxvNgaXYvyH4XaUCnARwqGvbpI7/BWK7yk9J17hLFOm5tU1lSqwZx05VeFBL9
AXTKdGjFaBdNB5ERwgufjOySwogcUZFwRWf7ShjE0i5C2Mbn8rpLW/OfQMbuJILPSaibp6zzAf55
etr8E4KUpEjswX3Usfoit7u3EwyEIQrBqpt32R6LwfV5ZP+PlV+z2Tfj1j0X0Gi2rXTuJi1VLdcC
m5Iop9kIqVIULj4MiGtnZzOJxXiLJqJ4ZkvdKEtANjcVvEF96r+YB+whNDXeQmyunk1mJWmmXL7l
LKPO5UoatIgw7SAthT4zJCr5/G2HNqNm96tglq2PH6rn6EckRKFipPaRb4KgncQnYxtA1me/D35D
/qK8ExPlI9JDLlhLJHqZGf8JH1XnyYwiIvSznJ570aDWa+8T+ruo+11UJpO8Qb3Me5V2eosC+ScS
vmz98A6Wu0EifzzLClCxmyOUlfmeC8f0Nk2sRr9QL4Qcmz60kSQExJBSguAw4M90PwF3UZJpDPo9
VOB0LIz8iXKi6ol+HJz2m1infm/sJezKgELXxxIBWTjRxbt1GdngJL6dQeAw5e/jNlcTJoa9asTf
s+iwsHt7eXzJ+N3hUZmjJN4OtV2x6WLZgmaoFQOAiCG7LaVnUUkbFPKOpQvi7+q7KQrkfJjXtKgU
fHWaiI+G5ORQuTr9/c7zkvn1A+IAewdsI+EZDFkfl/ck8Kh55Y+NBgoF2OGG/cmCl4m3/JaxG2bP
hmn2f3vNFQkHEMRhobDB5i7CJSjOjTIWx7AebZEiAxOG/F9bOl7++/K1KXeqiv1T+WhxUL/3dxvx
5Mt3FyeAyItOq11Em1sdZB+7A4uxYwCfEUyoe8y/ildV78467liSnyNTZ3eLpCvW4w7SN6rWAvkF
R9API8ZcKYQpp4Xyzcos6EYJZ81WFQO7iOh3k5AGFH6WE2Eii08AIDJvBgKBpcxJ1wIfzpgm2yY5
7N/QPj9YMgVUBgHlo6ZLIfncXLkeDN28sdx+KWHPmV6A/oLqHObhtReADTQgvhM3TapXoS0FQ42L
cmCIgSL497S9kQXGeqGWSlKYn/R8lRhGbp1YG+/KULTqJYTmgiFUD8eaoiqI01Ujt0LMjIkbPGPa
8E20iwJgmWVhrIwz+XSLHk4vfTmgqVBLZ5OjP2Mx4TedoUghlbTFleU+d9YP3goBnapUMXTTsL5D
F/limRujSMujkv/wDr005ZvDwAF3879LVNVa47Ens4zYeoq6MRu0kNdtec/GdXP0gADmOuNcZj4r
vG32py47YXr8CXAL8YqhFjO4SHeSxylLwLM6gqWo4/5pXgf734I35KbN+7iYJPPPwu/63AF2CHtR
IHFvSuySa4mIF3meOoAp7B1vIxaZWNh7EN2B8GqpCFctgkZaLmHTl7eSwHQYd/iE6LMLLNsnb/1a
2lhykbqVHSENUqmcfjo4lKHNwQprd+BP6OV4mUHEhVjn2JUFUc3NczCB69xhQzV+bLAj0M06HsMI
Jn8zGuoYxTjekmbFvmP0nZh306FX45Vi5qv2VXTBhxqcFp6xaG3rOdnkXJgOc5rBX9kHTQDGr0QM
TfddcA2EmTHhvUQT4uDxZF0rlFmMt+xQ9ZM/Hi9ba19gltBs+uQH2OKrRYrjVheD7YOxf+P/LwEA
NOJdOheWJWgGRPY0Fxv+Rpwr5h+haeq43lK1WAtvu2eGghoUH5I9pgrUcV5zb6CfJ7020sgBqOO6
q+v9nV3ufYotDf2vkrp0xeXLppvbmgUavG/ULGRyD9r3hHAELDX3V2/reGW92ZYnI9+kFzXHuAXE
akov1hpYQaudy18rG6QctyY9VX80jXRKQChTCHb2rOpHGIzoedT10txfVlve4eqcCqDtElEhwseA
WR+DLfxdlRPmiB0ACXXqxMmOcEjX/dh3qoMMJLh9FI7EJ7hqj1Lkjn917wLzTVCVMa9CqfbR3JEe
tqAJwH8+PClred3wWwPKy7yre70Ql9PQ/RqypannYcM5CZaBFXeiJegEQ7XAB+sXZLY3PDBgcRem
TyHoWQdtLLx5MhzjZjdoBVu+X7yJLNCLzsYhhU3l4EYn4QytPtAFcyFF7nKhU/jGbIrrhNO+rA32
pmv28hL+9PC/hSO8y2z/m23oH2X5QiltXquYSB27zIXWYVaXHd4lrk8035NL35BMCx1MRas5Ut4Y
/k53VvMH+7QbmxN9XvO8XyIEr/DlJhBtF1WSuD1+NfC631TNFtKL722wXpTMYUnrNPzqat0xjQhi
wlkNtRS1CuWvArivsUKfkn532WMhOCd55UQytlvjRADSWOeuu+SMFTV1epdSJDaMDelRxIIaVpCo
EZEKAU+PGzx5tJG+ONAyuhwM4O4FDynNUdFs8Yp3Ou1yAmi6k874A/QAB0ssYaQkW2sqzj56Fc8F
NWxmlFlBIsHnuvlylDpqiJ9WGf8vuLquupbTjQTOYfLd9r1AkEvwfyFl3/OU+yjTXTudvUhfBwvr
2E3M++WqFYe8LMhfbPzBv7bDF4BH8M5wnbbQio5EbG4+usrMCBFa1sjkKamZM1js05YQP9D1gGSK
EGm7nSajV7na268g4zxVulDijA/9g3eHxPLvmz9Jk55GnbA3E9+hH+W+02ouwI2k3Duq4pMjxCgu
6ic8M8FNtV4QIoao3WzPDer6SF+hQL/10ih4Khkh7TvS
`protect end_protected
