-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
zfRsfKyVG9WWxdIma2IBCnUJW7jRFvHyEgJCyMOZ+nose0JltQAVM1ElGRA0Hmyd3Ayxk+OSK7by
a1nOiY91h7fE8biqit/AbsSn6iODlVl9yMiz9vFnoVrWD1YmTMKOsmNHmFGitWUrdykTD/nEF+CD
JJHnzc5gEAmV2223oXA7pN9ZlIh5ZBbJ1kMeUrpFSgZpk1WIn0/gz2tooxuJvrlIRMdNOFcjN8Ml
Py10CWQJG1FBpdeUcxlft0MBbcc2Le1UBQ13nlFUNJSUiaccxWgIgbxfq4VWEIhmYWuUhkxLib6K
JWXcaIVHG8rxa/mEJIIrkPbRvoRQTOSaXR4UTg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4672)
`protect data_block
iZV3ldluBRMUGK8DcVQIpxEKul6xqi4Gy0SzdYT4mXTdUs5Myq3v0WQkldvKIEgdPZx/E3QnHZav
xxRc+yLw5FKIR7P1iHTb+eyRFhPsqwEMH+fyq56SHQwry4EtZKjWAPkuf4AAQlpBVLNK98kuy4nj
3JNWteu+dwVWLzlPPVBzGJcn0hB1pVx9mJG/8lA2eErP2kIw8vC8Xn75SpbbVuSsrUhAlY0AFVrq
0Jy7aBoaRCt2SrBPEVq5LbQio0MZUksFYSbVe18bjbRCtyc7I0LCLt9zYSzYNj7a3UenXYJ987ux
/KQ5m0pd1oxKPYYvll4FltF4k7mMuggdgDytN5+b87KXOGmClIJkveBxLezQhN/Vh65xIWnDoNni
7vowQMgDxt000H9tHrVHkD4iEYSRI56TifLGpq4Hw5jcOChT1eyxcDTyRJjRvix5+gHlz93SDmDg
mxkx/ybNejf2Rm+OZqN51okvSUgy3W9xA/8X4tfTw4Sj/tIu3ts5YLkCn/1IGQh6ubc9LML1eNYa
t8jkYSvIPPKjz4EcBRLYIvHno16iT3/30zR9fbTQkCS94W7K3lqkXbewsJarTNx0ckiopRPqubMe
Lvum3GhHb/8fEbUT9/dpq+iGPH5UOT6vexDvrbCqSZpfYmAETifbLjPoTjnheop5HuSYbTF/CONp
9v0BgrnXQLWJ9HRkFhDbPUD+vgrxJCU9iKwG3Xc4DX3aVmoT6EVXGnlQUOuxdlaFNC8hBIaRLDac
s/lPTBPxw6XQzdYSi6RYaCSmA7Vq7P7P0x0/suXx6TpciFy7M3I6luDVUKsPi5VD/fs/oYNaW8W2
+S9R+sFv8AsUyR3Ww/fZi9rafonsBvf6M1lFkcsOB7P4cdTO+/JnkBoFkuAWOAJNluDdTJc+WaDJ
L5YwRbT0d/vFHpwi+Ae0lkWbq77afqX45j6Y1wfdcpZBahErIvu36q65TZv5H6LZoKxoB+0sT4JH
Y1G3x60VtyjCR9YqLrOa9ZOTwjJu5H+Kv5YqXTZxrgwpTARgV2OhVLweWQstcrqiXbc9X6tUJZmo
Z+Ww8xMDQ1JpfqBUOz3/QtyvSTe3+XneOprNKQ2wwgxw7Agy5vp2iZWeU+W2Q0ETWhhdradqA/I2
vTjJXzI/4f+OW5ofoeimgs8TJtESEsRPWQl86+0hvkZVhrDRY6gKp3uwb1vEhhW38rGlYQLNOSU5
SSiNVwd3jFn2uEbaY2jE4g0SGKRcZrbbnmzze/ydqDvDr0kgFsNG8sVn/A+XF1VMkmjAeRU+FwaK
DV8b0fQl/U7PsqdBLJow8vRlxbBUVyRiEUpHWMZnaOzpNIXKJu36zhx2tAyjW4t9LlndT1CiyCKH
DBmdnvn33WUXVuTsarlYNS1FGMTgxxHMpzIv072Ygf52INDDWNArwhc6mBX7K5IuO1rad750J7Hx
XzUoCpibQvzoXel1sr7A/yL2EZ8u2RttTDx3NF680kXOmmbXIxB/b29Affck+at+f7FcPOLlnpv8
Q49g0YYFfztYCSIVGohmY3WtTaK99kKQZd4TbWCnjDJ4tVnw8LeuzJ7Yo0J9qOftMQ6T7rOG9hIM
XKkDPf09hjVrLdodE+ow+Te48bs21bmPGntyf7bP8bTx9dZwpDD8Bss2Wc0fz4mK4LEwAoG4KqP9
/PWCfESqDkbZgofc2kuCoeHsvyMDV252gUqiHysSQHW5s/4aWVGL/3Nmmwa6TyEix3i3ma0kVEf/
BONkOhm1da8SBA2UADEc4z+LTj2bGjPiuXVB6SwSVU9YZG2zdBk+EhReNPMS3023QCSuE6dE41Fd
fwIIx+ql05kHB8y3bvmHELDU+pJITJ9+IrXRg3mOmBomjcA3kxWdlEO0yrpLlKZTCkB3veDapNzb
/U0NQKrXjFgP8TEcgofbBW6rrJ1eTEk1M/Sbk8Kc11pwumm6drzqViGL0HE5eKN7JshnoA2VYOAI
t1yi1N1H9fGOVbnPpeXccVghYVZsHk1hZQPmtfOBnudXye8ufFMdl+/mqlmtH9j8wx+2dqhrV2C+
MsEjkQqmeaHWOP+4rqrnJQgr/pjw/vAvj3CbCTpOu0I83xFmJ3FkBU7w/f/JnZqPws9PC5SvJ789
fz9/enwQ4Gc27qX9MtEMkc3b2FYz11ePysgl0ISCwdiB4/V0JCU6Py/MU3gb1SpShNF6dypqN7+k
9ayRo8TINXZDCtdn0juY3T2QqJ+3TJVolEMY5nmrViXT/b6hwwGoSux0GDoYuUpx9B/rrZ9FUW4t
jZhUNaRl5A2tzCWlQbzEnoWIH49YA79lAw2ffq+5Zsj8tPksh0v/fKy9sarE0YcoGIB6e/haSXaC
reNfJVhrlMi7wV0cQ1qsc4mxDlcE36+iLxILCHWm7WIL5DJpkWkGog+VKRV5n35LmhzP2UiYf+Qe
40/oAgChLB/75LEGdSStIWNyq5OfZiBtN4dqWKtOozn/DL1pZ8DCl/Htgkq3UvgTl7rEbPK2pYAN
iQcSjLgjYyABES3RSui3BtIS+BAzg4gmhamwFqxJbpCOOaF/67/LC1agKPgIzakTCcwNaAVNkN5F
kOvw+aapaCU/XihH/EACeLk6SM4MCOtUZqS0lkCutij8KuguBwtyURc4Dk6apobaWdR+xeodc8YE
2OoMrEUaBr3Kz11h9WqxNjks2ngf2YnUR9tNdkLcHszsDh803tiOexbiwdLKfU4dnTkkrN+jkk10
CvgIvKfU5QGyqSEb0n3XVA9ucVdyO53IXu0O6FC9KpoQCi3LIoUMH/Th+F8UQK1HzArEsZ3+K/NZ
gLSFWiiFGxthJbzqMqRAaq+mQl1erJyKPRvpm0jgnxI5W+fmwajjkePd0AuggWdcZdWnJQiuli2l
u2JnfZO4YUktU5i3BTsgtKi9fLYhl471mAMRa9tcT82sQuKwYNcy35lTqpkW73BX9AuQyYoueVFn
tX+dYhoHsMoRBP9BxUOERgRrzfR6f/DLL3++qQBna2oU1UarMtLbCZsLozwYhWC/OZeSm3RspJti
TWXR9zAXvSeDJm+PY1cIzbzIIT9TaxF9aCBRYqsUF4UJ4Z94EyNpdkaUXBIkzsIlocZDhpw7jKA3
AYS1uyGvhcQ0ItGYOSN74UdjxDx7arW/ezjTnXJwtjHve5o3a7Zw9gIeUo9AzB9vyNGGsL+38oDX
TZcVBZstJrhaViReOiMZ5NjzDxn5gm8+LQVeH3O4YueAD6c07PeRBT3x+Oj7maz3aY8d1Adkx6W6
q2tIrQlY73PQPfwQkE2smZOK7VFvDwjoNEybB4ZK5Wn2DTfk18Qm8fhd3OQRyFW2BNchYQegSVp6
fdIbvB2s4lwn+kU3WaZZPdyDGS23/uZiC7xyZeSWvda6LErHX8BEG1a71nPjatmtvkCbpi2wUvYk
vxK1/YCcEtO2zjfIlXCe7RSfDfBCs8aoAEz3SZwi6p2KWUquVGdj7/hSmb0ehU7Uupo9QsV3lHH0
rMuX1jb9v3dt1NP3stn/aDNL47OBeK6M5JjJcV41dGEUAI0Im8KWRW74Obm2EXjPqJAnShEHEmX2
F0R4y8DJ7d5xnIQfZFKa7FYEaEqtDTpFiM7CeMlIzLz9xlKIZJylcOFsm8JZryDBXvtA47LjQHj/
kordAUXCUrPXsBymIC7LNqHbM4Ie+4snqLaAPt3hBorhrYKj3pYGsGxeAj9ggMLDW3uHA33gc82B
P2YY7zYH/rGtQ8pt5L1oElnhumTIDWHl3PxhUTHH82R1AYLjom6GAdnBadInWQIRf8cfFxNam4gk
zCmrwYgaHLQDLzm4FcorUog6zYPQwfzbbK7GRKy6n37ycfUc8PmUAE3Ty2jBPgPCNV/ISkQG7cz1
qCVPQlXBk9ZCXPypRL/G0M33svjhNJs4K+T+mn1xtII0NCJYwQjZudm7xYj2MNZaD2j4PUuLkkCo
rwz+jUcvO7G8YiZpM0anunzsoPJFdc3B75XJ6vPCXfEqE5Xq91RBIb3GgtcXdlSChEfElRbpgkPC
UCuIm9xMoXh9/Wm9wWaJshEG5sN8laBgsNoS2jI9rHSGqGyK0GTYz+ugpnvMovYJW3XFJVm04NtQ
wVwatSoN3Nhz57b67hzW248VLJ5Y2OwolNPz/pGxDPKY7s+lqfsTzDoe4VGeGKGK6Lngryb/R3pQ
GLzji7qN0aF5aCz5v2dMN37XsWSMWhXlX5+opGbQD02RiwiZNErZV3lRbGhZP5wP7vOi8Cr+CUBo
rp4UqwKv8rjG8p3zxNanbeX/a6e1ENLHKVyuk74RsP9lFkBPd3m7y3NBd9vtehVN7HLb+gOqeopT
/SsIAai4EjCDltep/g8ycuhsBVvC+odMSFnI0BmDU52KD+EtEWvB0lNiR60cvq0svRFRrCZONh6J
D+wyIG2gWJUoMXMB5St+j/2q/ZFByhx29mpA38RZUw5IytcFTkyf+H9tVApk1hyqZPS7h8hWp2Ja
32oXakDTxRl5gxlcr1BEJ/GVmhscG5DfH+Iuj3fjzyplnP10VvsxeBftxmOaiq4gbrNeNSqxbMBV
/fwUXArm4sohqcc/IZBQMzZiYNcKiQESWZL4Kx5nu+LVzOgmEzfYoyOZmE288eXzs0jiPBqA9LKR
NiRHwaTNO4c3b1yXcQse/oVXnHsZwHL15eseZAtqOCnirGtB4XzOj+gA+1YktDZpZELgm8ZtOXy5
/8MlArtIRmL1e7TjTM0/nhcjofsvuIhE4bLo1NALby5WwgHdn1LNKaEBwqqXg/Pr2C8ZQJoEzgwB
0VpUpXTormit4Bi7f/vRi1GxOfVaQe7MEpV5lFaEGh2NqBVmXR9MYicVW6cAJy68BQqlOzvH4I3G
ABvcVkwQ8L+1zyvJEOZ3p/J5Wn03jFfw076rgNKydPO/IsNe+9C18p4bi57Ki5DVcGOfLHLlfyjh
LQ4gB0MxfMqawrybnibrYKe/lK/HPkbtO5KvVGxe6efnQwC2K0pnKDvnY3oB1/dV8KTBITrE6/o9
yj0ZilVhqazXp7lTL7qdUN8fpV4LaSsVidb4fzRSEKTDxZVCV0+PuA5vUOhedPWzgRXn8CTT/Bvl
5NouaqqPagPrJutzw9mSKGKZCgNIbwWPZ6twv5c8Z/Bk8HhdCXaTDkOP8bjs99EAS90+oXuVUBq8
L5Y1GanYLKOa2FoJ4f8/CgXBr1jwwC3CG6pjnv8TlBqG8GOySBDKqmo2BvMzYOgrM3NwAVS2K6U3
WWyTb5rR/QCb1x61Gat89U/bL1jYT+wVHByL/tBo21c/yj2e6fR+o8WLqpP+/YqzTMnFN1xpOgaF
GR4PUhA6wWeDQmHoBxO7Jg2avUPsbJWwoEBAMFojaoFZeGfFThO676PTkV1YzwzJlYsdtmvt4mzw
O0qoF6rnOrrvzdfCQsAs04xG+Wbh1BYi3gXcPR6Re1HLeN3RJWZ0GEvTYnHnbgb5/wS+nsX6EOuA
csCDKWazhgXqzp3CPNS2dbbnmd6x4TUuOMQw4jVlRf+GevD3CF3iZRRDynjPe1nZmsUQPf/Sbv5r
oY/0D727x9HdZKmN2qeqfckNpS5Ll2/pHn9ssEfAWbAnHtGRDXdhbg+Dan561B6cCoQgEUAwUpN/
naxhNte6u20b2E2IeVtWgptuUhAtp1SD9azoxXsQApVeoCKeFTJrhkryXtes4/LTF6Lqm8o3Le6t
8+yAcpKhgfvBqTumRlGUymVVTSZLyO5RpOCfzTmpiaI8N/2yJ8/056s1ylYABckhdIaD8D/2pP5+
OSBAXKNbbuN/w/mUzgxD3tG8nwE/OIBjNv+k0p6fQGC/+KOvquRcFnAYKrL6EGddKjXOO5o0vKJm
+oIDoTcezTbUS3S0a34SCoxgX9x+VvGZFiJi3c9z5X7P9kGmBt74FpbqZ6RTvM2zMmzVBDUO8UHq
JOsdUXhDYDmIQrRWcbmns58Dv9XyyqucTn7kGqzm6kewjCjiJkwx5La3MFlEVDBLlTtFdYtU9MyU
x6pS4OMqVBIhYAH1zuwJCNU6kO7b9TXyNHWK8EClt7I5grtGPbM3H3q3U+vDWA7MIasOjQ6z8CNg
W2cXBa0U4lQAfEHpKmFYgbFdtrYnEXo+PBT2bQH2cXiFYN5tmP4blzRYaPQEtJ6ztqTeO/26/53T
ObbQTM5goHKzQ8tM+blG4ccszbd6xknRJqq7u629F8yHToFVmEG3Ub/3xG9hfa6x2jijJLJZ+A==
`protect end_protected
