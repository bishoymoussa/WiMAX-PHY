-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
qb+0/LDbUBuDsiQL5S5W16jQkWY42SR4olaNK3C/uXhWYGR/qjvOwE8t6cBgFLoNZn2m8Q1MR0bv
qib/XCwY4cMO2O9bpR4yzBiPc0Q8VKhq7FxIER50yKAhd0IMds4XimQIih74XN/+gJLvwkNUksiC
rV7TOkPiNtSGWmDtsdnun967VasHQaGLUpfctJJlRscxVSGk7KJduUyOI4idgWW00NDJ4csksWU5
XEMFRHMecUpK8IAklArwgjfey7/Q4/nTM4eN1YWdKX/tplttcHZ+s9L6iVGfq3zQcrV3BIAVopyR
+6xrsWo6XcH+U4oz8Iy0hCywJ3Hmk4a6g4XFWA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 10592)
`protect data_block
PuyKjmreJ0Uu58H4SU82+Mk3tZHFJErEb7Vi71HcX6BfAU4t0t9qNLREff+Z9WXndrnONuk5Tptv
N7zqYO9N9TC3/NUpTRh/ZO5juS+iTR1sL9ADvURBy1wuGGgp1yIwMQrtv7mX/45yimwV9dLLjZQv
PK6z0IMd7fkX4oM/p+/hLlEfY63cxtrGBYBVRx+q8W9ZkiRZMDh0dzClrDBND5s7B8j7qb+rlhmW
cDLSoHd9/fJ6bMWs5M/eaCj+m9yV6zQPSZlyEbSxC5n/3x6p8SHVIgVUy0p5uj1Ng2ZtBdhgNt+u
SIxwYUBu4t3QMwDQ+9DCcXaKVdeKRPQ0jX1cNKk3Jol3e11YC7Szl/dC48RqoM9L6nfkje+qfthP
jPC+Rsa0xTruNSQYISfkxujZxsZ9nkqxkvuu+7rMfjJq993HI77Y+NRlTQOQfqgVmNjC/qw58U2c
oC2qaCwwl0mc5W14vtrDdQkicem4KXiF1zIDF5pn5VpHXN2dDGROpl4jbqaNYmEGUmKXuxUUplez
KHBCEzZOJX22Z6DykTlG+1iqjzme4mMlsn4MY5XBcMv4vA520qmPtPliPYPC3tc9QRVUvsCUz37w
UbNNwJPkK32VS5gn1icMfgCFRpxlnAPlqnNIxVNu6Rhtg78xj0R6YQqFl2zIYvIE4p7GJuvfqbh1
EhtIKoAbHrh/uFJcbnrzXtgcI5qZ44hERmT39JLdZ5Yp2M/hJMu7frJsPPyZEHLhAXT9j239Dfi2
pb/7N87lhZtvYiAPrKZ5RtVsOrGJdCDeGaM7i73zXktAJOVVjuc5WFmcg6MOcs9SDaOdvfzhmSkP
mszqEBu2cig/yOpb/Wunwom/+xr+TIZH3M8UfbyXqlduP/aBm7XBnMZlyPtUkDuH6joRgq37gOoh
ytEsOgN0I3MuPlYCDvIQqc8NnIbfWdYOYj6I0MrsY+34hJIy8M9vIObyDSXRNmo2Tb4ncUTbP2oX
hAgeWTuz5/IorRP3gWPEzwgNBmL6OdH7entE9GS/I+tD8fu6ct7p4YARqL5AcOYzLChTYtM2yIrw
vF/4xWf7LJat/5Zc4iY+xgi5xV4bLYlrMyx1CzbRB2grm+sBlTl6uQ6W01oLfwXX4X8JEazu1Rz/
SgCM+tWW40Eru5J4yofbr8G/LI+fXMAMq7q4ehTMekGRwvQG+x5XJbSsreXkJlVsaEHuOT2q7d67
uRUPAqP7Tq5f6P0MC3Qx4poUNA0CTEfZrRyljyhLvGBh4O+xa9Yaaydjq7c3Ljv/HWUe/zEEZfD/
Yg0oh/CSsNrpmBQVOXdIg7saedW7l31XbxV8yISg5v2zD/Vs5rYa0rpO0DUXdCD/+oaenw7l3E5d
y4QCywOGkO4rrEhXOa4Fvl5kDsixBhhicgSadesQF0xEC6FbYbt6R5GkGsysXJZGVb1LwqAjvHVh
grYOmYUoH/k1T+kPXhUslvc8JkJQ7192LrDCeU9QwPbZ5v3Qn5fdSP3dzsbB/egv6livyhK/ahRM
vTvYOfOo/3gR5S74kwlVdKZtEX2TmvC9C7lu0FPu+j944T1o9kfpEPlTFihpQYKd0u4ePm8qQYmP
HHbfw6mjk30RbSN74Ow1I1MoEvTPmfGh/QVpDtRVkxhTPuxti9+HLRlwECuU50Lpo54B/y7AbsYD
BAUKrDJeAaWdpOdl5CYXcsec5+F2TJlw/QbK8JIl6+Q6zIAXjYWl3XwrV9lTyq/k3h0Z0HSEzlkX
J3QDGhVoRFadx84vEV4HdRTDgIIW/meJSnR7l+ceCb5FD/ciw3udbNJEskaAWXZNb80pqCnxSM7V
c6JainWx4I6s0X50rwDOHy1fMQhJ+kvxiuHEAJNHJrKID7VU9gGaVRXW0ecNM+PhZJmoMLylfnaw
Zu5FMtOAJdxDGD0hohptca+t3fRX8jTyO8txypSwcpbhQ/Jm7BS5MT+KjctVC0dte3qPrRz0Y/da
shnDq4BCxkqsHM5w9d8gvs5f+A6WMR5NadYTh/G95unzuAzBErBszt8nO2yGhwiKUA4sL6NTxCyl
ecxw+xTnif8GQDvBrsY+bSU9cABMA1ftHsIN9TIub0QruhovLAktq6iyGn54fhvORvDJabVxB1fV
f1z2o9vsanRBjlvg8FIsivwvNyL2gLY6xk0DOrUhw+9ySNH7j80J1AwEFpmRDFs9af9j+GLAn+ix
G1I5MYBELSjZ9Y+KHJUrhVCI/T8lWE4M9Z/cvPMAFDYoMNAVMsdZYasukuNJEQj2PAplJqFnqzDd
9G/qT3GCQQ3Qvtmzi9+HGjt4SZ4yNzX6+zUq67XJx5Sac5x80f1gRqAMFLJjvahfEFsiZ2NgnqF7
CCO4n7LiDiGQQpGFNh7Rw04n3yI76btE1aKKQ0Hi7SGoxZ8IAivtGUCKeSM4zcsdz+6Sy1x0oWiU
q9ZA/Rwm5JQb7EecLUf04WlnhqNJF7iDdd7D+uRvHDf54bOhx9/EMkHlXVYAgtjt81NY4i2/AnzQ
gMqajfJkiYrzm9gxpDn+zU0cYfBJB5ZkQxr8tGbkMpFkwFCMCn/sg/QwtIvLsj5z9hWamzLIizfe
Af4aiYNteBO/L7/FP4PNIjw+8hNFUM+wtM/oIUvK+6GBTbHFiGIUsXBpE+hVB5Z0ZMtN5IQYwd0j
zj5qgjmdKq7gHmHxcAauzfH3MLsNpdWVbrQ4RMW5vGmhkY/uatHaWtNsmTweKe2QITQWF5wF9R8m
vWwl8f1KUOjprPPm/FKKMl0vyz97pU82ve8WakC040bC1EqbQdSoYAclM2ocBvvYWIG+gzChatc9
d8GBk1k/X6LKLA1h4FGwu6vOS2oLJK3KZj7wqCqmNOdOuROdfdak5fhU+GafM9XhOGDtD8dbtDja
QGHJj50j3Ei01B5pAXX3izYn4Uv3KaAj9067WtH9YrUAMsRumfoWWo9vpK9ISGcxfuE0Jja0VRUH
vNbvV7NTTPH9MIfLGrxJ5A/O+NP84HsIfQcMTRz4RxBxyeFjbP+QPA1MU9HBQN6TZS5lt8fWN2vS
ohR49fk3bAKs7tLJStxDBN32Voe/DD0gSaqMtnAQl9tqPPD/sgwI+wzijraXs4XItJeetDLn529i
l6XK/lWz/OhrykckRmAaI3ihIvzo6mq8lNAWZkflGAFoz67JqusjDeVpNjbrZqMUacGF1CrJzyy+
mUeBFLT0kTS/LhgGY+95piVySJOhv2u20LvX4DnUnMeFTb8tmWuncbotLGobhpmJhuSQAcXVAe/M
DoyjWA96hTC4x4VNsqXfIOScLuEVhJgqMeRp6ntVtiwO7NTv8De2B0w1uMG2dk/BDxfFsGY8EWY1
oTalr78Djhxc3MYHw89fwcjVADxsnyeDJTMFK7zrbMky19CImBEtDO5/rKP3EHW2eA/G71Z5SJFJ
9XxgIA/LMq1adVoOIQD70dxls97SJrVf1+WC6WGW+spBwFIp/x96c6Tk1/wI/sFXUrydbX4tETm4
pQcSnnJjI1ZgaodKmHqhTJZHthp9Su9ft3ut+7hodrdWNwZhDhCCr4XWmI7MkZBXw6Msq/UeV5vu
v/4UrqmQ9TddrchFumF0d1AJ6vXgpXPn4mKIl6QZBE6iKv6ROUG84P5ttO0VueIY84KJx45JQTHc
12Nloic5mhHDZhgYYdwczJ8gSeklDXR/iT+IsIGuIVITrmaGxuCl/FpqDM+anv/vUAChLMYMh7Uq
Me3zI1kKnhjTDYMS6dJVc1DM8hRisYJrgL6IReFpDJcLkN3HynvSj0sEYKBWjXGgdwtQK5CQUpq0
ttkZNa74h0yDn7peYui7PXNeLUukS5ZaXyl3LfnGuQ2hGDl9Vekku/D3FL7EQyP00fK18XOJCGEK
JfvkVvnHiU/Zno84dGffuAkbweahyMclN44DCl3//nG5HE7TihKlEtqOjkoAVc03WtCniI2/iZEJ
SvUQromRnPDOGIlTj3lGPgqIA5mPbg+4Fvke7148YGK89meQV9ieFnXfShIaoyLPliG2x4JBY318
M/jD6BefXiZeN7ksflUgAb22YhArwYnnVQHaHpb2ffiIDxPUMIbQxVctLAF2dr3NkNwLtlHAni2P
UR8lQORG3/kcmV+SIGH+2SXkigcwcKn90XDi40sW/PevfyL7PbKcbVnHs/1xr991I+t1KyCxRsiG
AD3AgRKJk0VDkbbwRbiOBchZ0+vGvKKdLQU8Ur/78EsdwIKw36vuMfB5NDrKjKNcQ2zvHOke0vjf
zJd79b0B3+5OqzGm7uQgsK/LrIFj1r2Elavdp7eQf/F6wwViAHk/qgitoGSu0woAOXQ3kms8stNi
MJCjm76Y2pU1DhJxBXe+m2QelURGovZXIci3Exm7b7lJLKyGnB/twFaG4FlOh0B8NRQEZp+yPsiC
ShFiZ/rcZNWaArGg9OEgOieV+HAb6iMW5HTVXqNDnKBlOyqfV+F9bGW/R9dkaYk04qdZ24Go/ENH
wUgVTSTCqPQsssqUIh54LowjV+3t/RroLRDPKUw5zjY3gQNHL6uZIjQQ0jYhq6SUFa2m5B9ecPcz
THg1xEMjcI5q7h8JoFZJYRMGEfapb50OaBdoKlr7c/5KWqwEyboRjP3uOTRFd+6bqwSJGBEb59VW
c1QzRlkr/rKiie/iLQN00vOQUalc9ERavaiYZ1qRE6z9K2v/YqJYtWn8ZPxBpTQA1FaepkgLOCzH
Dz/TYC9eS6+ceHY97XyqyuWZn5rIr6rTgexuPl6NuwxTrfQomzD77dBpNd38zSM5Bu/jicmvidXZ
unbuQjPZIvaO9YCpu4tY38YRUzKG08K7NeZ1gRmI/DBBxwJniKxa8FaxmrDX8hEXtDijzz7zxmo0
yvU6cIqglafSTZGbXIpjF5KgV3Zk9BIf7QR2xtZPVdl55roahqX3QfCqkUE0Yo0Nj2iP75CkQ2GX
mslXkIsuRyEczU7jevaH2FJ5g44jpXksVmTNbiCyJWGItXadeHCUH92MHEYvzjpKFbQXpFFd8afE
sTXGx+R4NpjJO+QCo2IEjkTkGa2UrB3nVwurAaFbZ1vPqQFw88Htao9y7QgV/DQpwnd85yBrKHhj
9YxK3WgZpY+dDS+c/34ogLEAgNqbFHo6d7gIFzJiz6Sljzz1kcotEL7esb5OUw3ga6dwfQ9wUqW+
uceRjkJud6/0i4MR4TswsZupN7tOlvTE9FX8Gb1VaaDEKKBK2z+uRvjYqPJlYi4ZSHUHqcJK0icD
PYqBJdPOg6pBtKFzqbNS43d/putx11s1ve+0wwqyIqfesLx+alIxmp8LxAztyDD1Tj7oRC5IRdJo
rGaI8vYOv1Mo4ylQk8+rlU6xeR8HhYWGJla7D6k8eQGoxmj2CMPUSM2YD0IQrXexIYR4TorBNlwW
JsFYo+MHf87xsPF8tMi4Cz1SVbWcizX8XXPNYkS1vnjeDH0s/OtXL2R6Zr3Oke45LncjWY5fYAHd
rfzUoEP3HRcqtmDX0R7Ocphtw5/BnK9fJEdYO9OUPQo3Xm/mLdUKqJUUYHQLwBtOM6l+BmrQ+2NZ
IXLUUOOfsgmykqJTtNaWCKreCCxJH8q+ImI0aAXQ//2DWagKVVyMn9m2DfdJM6ewydOoWG1tflrZ
syfCzV6PoXYdtINqeheQVClTvsnKKCnnpiAn+VIXjE9Wa85O6KNtWSa0j8M/qR6zBCXFtzqkgQvz
FaM/Tme4Q3wM5umhY91ku+uxJN6yuqtlGdXf4GieQXwghPGb7zNPXJf8yhdEj3nv2hcDdK5zc/rY
1Fed15fGsRKkm2PX+UIjTc0ITfIRZgapWZmtgfuSpOvKhEKoVk1VKzVbaDuHEmqan1/ZxhTsxKdm
2fVzx9t4gQ6n9HTR35BvvhYGXbZMN8DwrgqyumQFt/8IuLpsmsiw1ozAfE2VcDmFm5KpWwuOviU+
q5HFXutmitkSKJvSz6B7ts0Ow5UeF+9MzIKsgvRaphCVerRxgKGCc5OAW9WvTivm0aLFJ/foaHJx
PWrbRanDpVhCrDC/h3QGdFj8IwegBwtWUcFV6suBAhCmgkjBH4ONP98TFiXm4/5ruNOEZoiR7Y4k
RD3DhA8obEkzP/3j1w1dFHkIWY5iRzv+Mw3YwRJeCdw1pdf/j2Nw8oj9EV9lcc7set0UM3onGPP+
dynIKdTRXheMHNKaK793zn8/BL4zShhcjQJffN5qnY/NSV+K1Twf/CUx0ZgSFEedpMlSlTVuqXRu
I6eAi/WINei9uGI6v/o07LZzHYIFJIV5l7vqlngqFvQNZ6d8b9Lly84V5Uzc3FXNxB2hy9dRXfI+
yiQlsQGH9FQKlXBCetP4pkNZ3U83dZhLLCJWJkT53ImT1NuvZ4WhNEPvDFLes3wt+I+UfNKtkoU6
buHKa7TjNqBCVY99DZIENOeDTuPuJr165efnFHmDxe8WAH5OzYyQGkQFmBm0vnhbbt74a9kUgQrT
uChjfoRP3czA8opSH4Vl8LSHlQw/xD/JTlVGUsrX6LPPB+Y4TRZvNWsFammrxAkeihkmbXPUXJtx
aXhbB8lhcotKvmBMHVmKDJlkodPjFNjbCishxf/Wk7/H1HkW1o7Syq6eg94DARAIY0xp+kZSdtXt
C4p9mPYIgfKaOUmCe5i1DjEwPztDn0dI/DODnER3qCbJq5OtA4ok1qbGc62SKE2csURH87ZO2b41
Jmi63DHo6WfeeJ5HCLBK6cEw/j+J9HaF0RMTmYsVWUVwq8ZwQxnRAJcooVF8yeTgI5Q8uIatL6rS
YTqpJfnrwrfpPo0EmvzIJpsPkSAForACqiPH2zi2Ts8UZ7xV0BpheecUstAe0jJk1wy3tDVDePEM
C6ZVxmO3bjmByHuj8P9/OHSOC3qOTmnBY8F1cVX9kO25834K5liDSTuLxyt4FpV/2kP+Ty5bqBL2
wPFkgLMFLihl/Y2QGPEFmMCM8c8foeRDMyi/Fz+6L7fFa/g2p9C1CwdxJhQeKz0Qo1zd8hwq96K0
TU5JLGr9PVi+xasTascs7T++ojphxLQXaJqoKi+uSsgKOjZ0ARdFjAi3n2IsQntjjs6MCWt+us9q
2EtfSg9qGGUQ7+LQaLuPQ6V0hEd65mFWeIwRZkGX0G0ynqPTa5Soq6Lvserh8A06/jKR3Etu51AG
ZnBY2ZKToNo3LrptnX+FYaoHrenfQhQmG5t1ZvAMV4+kfrSu01H5Xq3GNxA4y0ZgptFlhfGI/R4d
zEdHPI0lyKGAiv2ySkl6nu28VyamhEGY0ifb+1XPRI+ggj6v9fi578iMcNCq3lnQ100cUhJEg23F
4qg5abXctHfqFSUSbdivQq/UiaiYguHit0u34VVUh9LOvsZDnFEbyjOCOgKXshpU9OEVL2XyEuTs
5ve+Ye9bj6ef3kNIPWyjpwnXyZde+z4HSRGISMeMl4jxKFVlHCPMyw29Sidrhsb2rwYwQ9lLKcvs
9/V1hDzSEgpWB9WbPA3OcygsAOfob0btR8OroG4F1v9i+xpuTwXNwpo1WRVdev8KnFxZX/sEEQGR
UA9dgka1S+xVVLda3rJyh1d4YDn/a17bLHfpTXnw9Oil/wC2UQTA2FnUVhstxAfk3TRphTPOGVtX
iPaNtMpafKNe0dv0Whitd/++77uqfF12Yu6IqMqhYeTuNNk3cI+ZjEcqw+S1HD9t89mPabFtmx9F
B6QXMrSCzTci3PQO8aQzx+GuPyi9gnYucr11a44eNlCwhdXzeGgmhNycHSUGdkRpEBuUBNMAYPdf
CjntHVDpKO9WopbVQowsEcMFxAB3Galy25N9xdQMKmlf/AEh2I5+G+6KAP4IOMhlgO24WDJJxpBO
Xmx9VIZvLpIeb/G7n8+61K196ScFDmRuWEziMwtEbqWI0lxYL6revl12+Su64exCra2S8vb2L+Tv
xGEDfssawCr2KJhgm6pTjKOzSXnzluHhilY6cKHg3ja7bhHj1UIYCHM1Di2JX+ucfiTKNF5x6e52
JNWjc3TgeCNydyEMBuEZsFMpscdOof04Z3sRET3p6wOlPG73Rfx/dqM6DAsvItuduoNugDspwdhE
eKJoeUzGXPf/1T79zQH2J0YsYRa3CXZSsTqt9P/V9aCa7i30eeQvusOYbjAk/i41vzLFPIi0wRm9
TYAMvPWz/oCH+3SB4lzUz1Wspm80F0/XF14sCZ4YIeaV9iurQ0qHgPAi33b7iuD0bNmWnWMHKLmZ
+v7hc1Jxfx3jzZHKg5rmXPNlNMerHrLLxsJBDkNtaQboE5ipNTwr3Ed/IhFtomPRVJQXm3DzOfK9
qTl/71aB0dpLqcKRtIEnJGiRc7CybYwzqYXTSdw1eN0WTkEdFeKFmJnZRkjCrb0Om5/Y6b0389mV
nPnTx1xWaGP/y5omRC/IRMRx9acVSpdEHVoRsfY1JQQAQJUHFYtDZH6DuujG7YjZhuPJCrWjDN1o
G2b6CnAK9OH8KSzW2cpEMQkD+TXoTE4O806UzrAM9gGiSgq9Z/Nvd6cQ21Y/4NL8wbXlXkLLfFg+
TP2RGuGAI8rqcQO8XkJhGhbaV/aG+66Ggv3j/nOAziuK4UZHmWSzJZqi7zRxYVPMyKPRVPxtO+nB
JM/OnJi7Y67wq8rVQn7hB1GLMkp+HuOZCJfNOaSyW3XvDARTwQGcZyVx6g/MnUl8nqogBOLxnZFA
s61JHm13IFcZoHKcOKHXB1segMvQWCCxzctuehXJgez11mxaWzTRiOVn8eQiiucOuC3OyZFdM2wx
d3d+u3RPwjU6Y5kgTcgCh8cST+IRr+52e03U5wZBOppfC8/voiuKpCwSwvkSXAdw/Y2ZZfcCybJh
ady51kLlOgqOe6EPDsNjlTYC2PZfKzXwzEZ/xNkAblrMFXmMyt2c1X/Jh3Pfamr6WiuKqUAqft4B
jKrH429K6et8Uwdj6BgVBD802IqNdq/8YzfBuDHjIGprfSopzjpH8yozErMVp2Lfjz79owztGN39
ecCC4up8Ww07t1q85wUbBdjgcR4Oj7eRnklUwnbLV1bIMvFRmcelEAatmJSFWLOlFwTmsxPqVsup
kfHHkHZBbOIJuLXa4PbVtRdUpDBcnv6hSmsMXrcE8/JFOxqGW4i/KpBFOTWqjyR+prehPNxdahDo
WgJin88n9BryH0EEUOxmtJ0vp4TH9ORvxRrt29MdMTUalwly5NNd28D3vz0k9Sw0QJDhXnFkf301
4KTmsFlswhOyzjwDO/FjMK/GYQduuEtV2EUfm2mV7U40zi4rMnGK1TatQ0Cx5KMs232AMaToIqqm
HCEx3tlzzKUGHLFAEhrNhkTayilRH/BTKOYyUr7kNA7v9QadPXJPE7bMfFQp0z68NTsiyjx5v+8w
qUhNrsWBB22jVkP+g6W10yi1pZHk6C0BqrF5WvGlUUeQg3V/9ZNbtWD7s8F1vNvFyD7j2MH1Ikqr
Ra4OuaqFB9GlQvUxk2DZRi0CA0ma2eYtIqNxBZUf6M9o1fymjVNw9XIpqUZ4OUFUGzjOtGSwrBgI
juKsqcoyjDJr0swNVDmo3+prRHGiGDZy9U0XjxvJZq3OMPc7Srpxy2H7gfz8sPoNIN4SGsccpsqz
7J9v+sHVYdvY/r5zLJaCgodxe9PuddsxalseynCV/9KbUrwvit+hV+qTaV4DKLYhe3tvgzRk5x7G
tSWMaBy7trUxf2z/88X2UiePWd45t7O5GajuH0uyAt2ZCAcM2KqQeayEPyd1ZAPhd3xKN9tTPtnM
h0NJhlc2ofzfENsYD5G/8DAdMiMn3Rdh7jQPpQGFBSd1ciayw6RgngfH6/zgHwY2zLovcqiIvSYI
2oChG5tKmDLBADorWeS/NkXX7AWR8u+p1PSFwIEfIt39cpvNmf4OYc8IYO6k5KZ0VkLpWI68zKCg
7ti6jUB0wAjJX+57TCauHNyS6sc4kxTfa1v4zvcrwWNHE3cc4d7vedjAtiX8Wx9/ciJlUD0z+lvv
P6psZbIrg3fU3ilOfW1T246+dlV061nRwVjrf+jtzoktSxeWVAmrm9ZbVGOlyPaJEc6+IUoN9oCH
y1PhWFBKhkVUij6cZR0iptQEskkjXarszI09EIWREhEd5M6rP5EWF/F5HPFaB7oNIhtwGVWEJKpz
hIKm/s7ugADo+NilQgcCOzPiNFpkKQNqErD1TqrqbYe7lypgYzNuXBbMlf9GK62A9+kRnuQjEGKj
woLL0W4JsELCTvAXxwFvNqicEEWHbdC2jTRSjlzAbRi9Azr52u2UC9hp8qfioMJ7STk6AO9ynKS3
CCbXOay31Br8nie6Y8ESJOHtVuNwUdYsDAJTfJWcNUMkfqeEmX1jnv/Wvt73Cqbg77FNLtc8H6YQ
KDUbG7q5WCrMaItyIyqfVjPAhcoaoEUL960ulh6UBepE69EsojrpNDgsPCUEvz62Z7i9KB3OM0l8
0kWrRgb2AqWANZhObtp+N/qD23PX3UavKoPd85axHCYYefQ1t4MmELIUQYK3NjAFXbRwAUaL+GLv
CiRGAc5NbUEj+mNjTm2mbzmtO+MwNbxBYwJh5cHG+9Y4gS/Vs2/U6ILQl73Ia/jfaVKRBi7gp449
RwFc7C5ppM/lWB8F7TmNjtvGq2ViW7+Um7wIM/IxNdXc+WOtegcfnihrUn0jkA0HV+4AJmD+7iP1
MmWX2ZLy29xx0vuACs2O5euxhIJrLGSsxGQLaRkZgNJpz2WxRNI1GIZCAhEjS2FPZ6+JNbt7IyCg
RT2fid6psmzu0SAj/ypltXWiB6nRfGB/zRg0JoegwjTmhiU7RNqQLXbZemGZF+/5ic/Ue6na/4TN
NYvPsHrsDS51+AHy17yUUNffPjw3282UG+tNjuQoV+fUmHKVyMsdfqwZ91qTVO3tSAIvhJsdpA5+
Wgv6q7/d+X5myVMyLbcF56pO8RfmY4NVTGhvYX6O6y7Los5Mxl7O4s7SjVM9tnmrRl4a/NkFq1m8
qiWvzsIB+ZCfJM6QWz7uXGtQd1d2y5/Q+Tpx6xxq5k/uw6gn1eKuQil39vmQJVVnfbVJXLoMNFCR
mPqCKXdfiBJ8fZEuEH7qN42iCNnx7WuNFve5xw7tDSge+IlrQwLfX6d8XT/SADu604ZC8AiEtzTM
4HuYGHG/ZK55qYxFhhKq/7wJ6YGgqccTKIHWtPOBrxzbvHoBfnLV1sn2OxIkPYfA2HRMlxciwo28
k/753Pd5YD3/XV0Ny25KEq0uWHpbjjTqFLmpmnDI1JS8cnjgfjxCpR3BWIynuWos1bm0up52zEXg
v6Z5ayyMD+OdScK1RhDsH3LBWlPSt0t9hNmg2gCOgUynOcsdAA5HxSv6w97nyON6PxHuDJQZ/D5D
8YTbk/npj6OevN+5/r/Fr1mcvSPZOSL/V4GI4m9P+sZeygprGQXEoIVf0vsPnEni8wga3rlwe2n0
xXGCxNAXUpHI9R+xmLg0JYpFR6f+/0T3855TeMn+8H5tmW5gPnuF3VJWKT3Z1NFF46aYegswQjxl
Niv5I3gHtV7YrPhJSroAEGutHQ5r/p/6EkLuA4Kqk9142eDTkbrh4AqZ9wlCn+kbdocNthFSlmA6
kHz4dIjFnZOCuh4epFbqsqUhVuO0iv1gMj7jeoDwILLzABQyhKoLBiWxhCaZYFPkEXgy1AN13EDp
BWWbfbCpY5quFMxMeEq0S7pQDdAan0/JZzX2xInvG7xs4O/g+AZZFTEBl2Bbd+CAYMVvnEhXjReW
CkWgpPmJU7jwNBD+J95LA7RioSMpi98Gxhdu/meO6xHJaE99bpfFQAC3d4yss0I3yeKudTGKC00m
X85UA6vD+GsGGu4yZr9edl9eqMIc2Q825oUgAUrTWuiTqunYstG67DXzGaaGn8m7OC9V/dZMLJci
V3zAZcBjg5K+1NcOj+tyABgl8PCZIi83ZCjSh4EgYVcT4N1Ra5736Ry+fJukM2Pt8pp6w5RcGsPE
GftOSR6eNoV5BFoILrvizXgl0hSj61THPhlzHv8qYIvNXqr8Egl6x4qsduaTheyfMX5NlKsmfb6v
M8O1KGDD+r+ZZkQLV/4mvijAtJcH0xgFTqB1C/0VIwhK7Qv66W95bvGq/OIERB89Yk3mHPOnTho1
hs2t+x8Uzgjb8yky4CH7A9N29AZAt5h/97UKkHf6qEh5o63sFq4VWnDThkVjMgzoFxCP7dCvgfu8
Wo6WzItUi+fe1P6beVa1U2oDAYf3dvUElYzUFD/TlsllBeWbTMRwxChxAp2ecnOZQj+eVpGEt2MA
8HJ71r5U4wozUWLTyGTDH8BUDLijey26z41SOsOo0ur8QLF5JvUnmP/PXRGaHT+B/zOFubNNJs0Z
s50Joa4osx833OnMVyrg40UtAfysryBho6xEAodyDDBU0mtCHNcAMFq4kcy1LpPdjK6yXLxrrY8T
iwReQ0f4y230f/M86BSEkR8aeyA+L0tP59J7OGBPbaHUqWkpYK+/FGfv3d1CupGxyovezp7pcaca
ciN+M4KZ3xsz5R9b24nXx8e3EhDMcdiLCBFybkIr+LsnRaRysJ/c0tK79ULtNagIGZViSV1CPX/1
PNeCT+HDEGO3AeNcTTwYGInELXzao/3F//wkcwcSa12oopmGmuS89SC9oFrOz57PR+UbYRyB/a9b
jUqD+01OdFXEJ1NHdeAAMhPG4iHWKUZyNOzFW9ZebYIEhr9SAryGXRHXJ79q3T3ffy/VH14viIML
pvK03YK5J9RhsN+lDlTwg4Y+QrTk2/07i5svm5j578Pe3CIOSQo0RbF9+PiZ8CpTD2yL2IMPPsmQ
5cV3WAZQw83QmdJLXacoq+ji2KoVdeGhFcfHDy6kDRkPrjyxya+akCQBKySMNopbu4NJ+hUHv0ZT
fzZvMcBY3hzRWm31SNEtyQIR1ZH0IanXmel7ZPa+xCDVW1HFkjw/j1CiVIDrzYPkO4Kk1YQvUd0O
VrFQCAOIHJK1mhj4LOtn81E34QZf2Meq/QPmDDPaW2lkDGl6s53bj9xbKHy/MvmGf48hwI67G/ik
rr0fOa72SyKbdQ0eHMuOjtzFFX0SVyK5vZg1Ei5aOrn8PYxfHfQfnyvljWBsk9ff08taJTnmvtCk
dRj9a3OTyDEy3BttY81xStOHcKoRSGVm3tqB5yuiaHeOLnTP2lpfz1ouER2EhyUOpTjlCyegbxMs
Ozozl0d87EzCyAPuqaIvo1C4YGvUj2ZoG4IHcRfIIju1SUgJU2wZ4iZaDDTN0OIWeZkvrg7CSGy6
gKTy0c0JtebjE3wxdUh9rPIRdFUiLkZUGT4ErKZo0+YByHwboUSZ4jbz+Db7slNn6ltq+vHynmXB
ylyhZK/pVREtZGumzKXxerF1CwQg8Q6iyxvpkySnyKZ51OwYnB8p0Fx3/drOY6APgLudf0BpvHwt
UB7o+P1d/dPYTPNFTF0B88cEWqlHEDCJWm+p1+t1JsmXEEtD5RIYmCGH7kxGFqF8JI2E/zDa2qyn
zFqoNGd2+pdmQWRYfmYedbBbogQ+JSqy9S/naDJP4vBUYjK1D2hFU0O9WzNRFiW4Nfri5DWvGtCW
YNrFf2B+1XiuirQfFUS67at2vqSWNxPpgm0j5CaeeoJ+1R8in+or4FdhiG662dOPWm7TR38Ecepy
fDd7uBHiC/qp8DgYGj34J4ljQrndfyFYDiVyPij/SZqdh9JVRW4UNAlgs3n/dx6XolKNOmq6jmlW
O+Kq9Zyma/Rb21mzpmKKT3abzcTp+i4HocyqTlNyxPrmQVdCQh3RTRRbV0a1i7Fo3CynHDHEJNg1
Ynr9u130urlfI3JD9yBoCQ+wkrn12V4r/LAJETsKCXs1l8aPvdbJQHfM48AOJ+WgR9NimD7MpSay
onfKc54+h5jnNbSE10qQLl9TP+6tOpOuNh9X/rq7HztVCdh6xg6m9waFO7SZZ7Ef8+fsfA1zlWCD
My88MFiodLJJg6OBwt3OSY+3+r4TimgpbNxnOMMIpBqy7VwfL6HzjFOvTIwL7oCEeMwymRtkBuLp
yF8pyXXgjaOji4JAumKPhsQYu1ZVMtcHrUn1P+/xdAEt5/mvWzfL+zmuPQKBV68ZAgjce4Sp2zno
yUeNriUTBgHj454VNbs153z1xdkB0Xi1+TL07FOMwKr3rYvRYphD9t/WrU/PrA0=
`protect end_protected
