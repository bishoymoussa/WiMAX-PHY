��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$Rx�y�<��wA�*;�x���@�̦�W�X�fa�M-$u����n~�%���P�$��W��kYَ���P7�?UMfT��q�6�U��k�>����~�\N�(�����X�e���/6U|)�X2pF�]$h���d.���9E�	�IN�f"�\��e�z�y�b�����Oo2�?�qˁ'�͜k-�K�P|����y:����3�l�d���bl��ˢ_�d���kx�rq�mh�MذM�`aS�.�DW�mS�9���Y��+�>��!��!�T�uOB���,��\L�7m�O��W���6����'���j)n_�I����2:��$�K�2�Sʫ��l ��!���{�l����.�j4�	��很�̢=�����N��s���s5���_�R�>����ТP .W;������	�"�מԫ�����]�#7@O+?�⡾�Ԫ���e�O�\A�	�ͼ���ƹ�d�	@�nQ˰��E؁Bf���|D_�%au�-�'���w�*%��"AM$w�*��67������Ic+u�Xaq�<��/$tԵ���.!8(�B���ޱD��6����1_Ǚeȴ@M0��} � ��vS�0��QU�d^����Ȟ��h���s��4��2�E�/�Rl�wd3?���WM`�$×<f�L%p;�]�N���|QkC�	"��޺�	$���F��q��WYB[��]<�u��R�b��S����C��1�)�����*�����Q��F���$��2���I�&�H�ֻ�u�F��շ��md�z1����)���*g:3�������>D%�8qdN�F�ɝ�|�2y�:Sfʘ�Y0����!�rwө%e��
�d����� ���.>h��B�Rn�J��Ij�����L�{��D���K��BwV�0 ?R��XUqHlW����Y�>|0�a!t��wn��:��;���36���Jl'(m�m�{��E����jL �p?p�kw�	|�3&[��]]Ow�����X=����G�;�>�µ��m�%���T���ϟVsDX�^k�|���I+a�4I�tn��m�{	ѥd��T�+�v�vq�MF���a��ǵ~�$��v1�q��/9��|�r
E\:��~�˛<��7g���F����'�AP=�&�[4D]0�~d��H����1��P\o/-2bShE����2������g̻'�p��2-�<�$��_ПE32�:�7�9i�v}@ڳ�4c�uUф���)i�#Oݣh+����!���ܜ�#p1s��I��%P���9�gآ�������U��j_�7��5�p+�X���}�O��\�'�4�-	��VAg+V��,�$X�b7&srˏ� /)�	1}��}��y4_Օ^�/���h�P�,�+U�XR�3F�S��)_��L�J	}*{�F)/�i܍��]��ڊʁ�mc���
#�5�����W�֑�$H�}#.��ed�I���Bg�qF>,��+�M��K,[w1�.Cc����:�,��E���u�ױj������D�i���g=�=�X"�aȘ�W�(qQ�"�sG*�XU�1��v�N�K�ES�ݱR�l���ɴ,����a0#�e�� �����Д��@�7�?��Z2Nj��?HN�Z}CDBf�4���ü��;i@;�H\<�Jd.T��t���HE@J���il�@�A.Їm09X+� _��f�+!�Q��Pi����ã�0�T���y�D��������K$�2k�30���N�T> �B���-��S�[�
��E�8����L�*�Y��/�W{<��A�	Fq47�)⊇�["�����,��n��`���.4:X0��XQהּ�R�{c31��NFF���c��W]V��](m�L��PV~����u�$t9I`�޺�0������$;������_�M�2>Tlpўg�T�z�vC�2so�-)}�E>�O}e��t�z�#���^,��I�;�V���ׯ~ 7������Ι�������X=�WZ�[A��ܻVrފB5�[;pB�=BI2�AL�Y鹬�r�\6?vυCFL�lHAA�sY8���A�\[�1�`���t���/���"{ǩ����I�`n�.��O����+�q�ǆ��r����S�����
���>0�/�gܰ��D��Z��%K�P�LBZV�SG�O9�=�U���>���cȫ��$�n���<8�G�?=e4�'q�T��{/XF����x���`�cp��Ԓ�piy�n�NҾN1*BB\|Q�f�ؙyAm9j�GU�X>C���f�=#��1ѯ�5������V�:�G���vfg��sy��l�ހ���CY�?m���+��.2��ԇi@�h�YmR}��$O���r�b	r`�{��b�DqA��
���n�]�}BL���h��h���ȯskbR��ڡhVMyH���P�~0�l�d�~dϗ�HT���@.�t��<�qB��|W�pfÏ�fQ�/�W�$��������Y�j��&��� ����@9�&6&Ў�m��
"�ft�7gLcd�}�X���ݔ}4v���>��ܔ�
�t�[	����"8����ףߎ�<:�r�&�<��w�t0�3]�g��w���ſ4���}IT{D�P V���o��Rm��gҤ~n�u��B֊�G��*c�6NZf��Ƥ<�?q�,�5-:�%���w��y���O���qN{2���% ����&�k�tY9^Va%�k���!�� ���]�<k���}3���O�k��rY�y���MJ�Hl�}�i�i\ Ynۼ��#�I�Z1��;E��g���5P� ���/zII�ܔ�Ni�b�7�U�� ;�;�+mzQ����\�Ώ~S�M#�o��w���"�/����e�ga��YO�>��{�g	Bwۂ>�'!A%Ws&s�uYz�f�ۺ�VW)��f�H�&ӹF��E�+V���sI@���6�b�F=+/� ��f_h��ݷ�C� c/I���$5C�5����oQ����O���0
*�W�c���iMۭe���!��&��*HE�f���B�H��fKw���������8���f���;s�xH�~�w�=T��Ml[_�VZ]U����o&|M�*�e���Y�oNqh?��!���Dk����I|�,�ؒm�y%s[�:���ؽ�^��s%�:�Ģ�Q~~ߊָҾ�_�yFG(�<L��s��41�u�*9�7xb���@���y�@CT_8�G�Q"Ϙ�*g��"$SNO��_����/���~�����mJ+4��(��7�7Y>�'�ų)��R���⛟��^󾹼��
��x�G_��-����������%ҷ�սRD*�]�nve��7FS��b	7]�mޓ"�jG��5��=-4'gb
�A9�-[�}/�d��f�iTO�$�{C�j�u�4�Tn��R�m��׭��L��3x�MO�L�\'&!~�fNA���ɨ��P��NOz�OA)7��-�3:�����r��0��=��8S"��D
���Z^�.�</�ة�$���9j6)?�h���U'\�7�rW����3b>�S鈗�I�����9DaO����ѢwÅA)k�ޗ
/�}��7�A3Z�E-�J�O��^hc��|�tn�`�h�T���r�w�� o�I�>��*��]��.�7��J���/�_r'��R /�=K�k������EOY���r���(�$0,ܟ�fo�id�4M�t>���}��h�z�c�D�v�1�����aޔ l+Ob����`�-��|e�J����w G<GD�2Y˿]�G5���m�ά���<x3�m<i���C%�����4d��/�6nݠ��d䂅�&&�l
�h',�7�,�y��X+e͇Q��C�mB����`(��=��3�����Mm�y�#�����+� �e��Wu߱�f�����o�n� �4aԽ��c""��$s�ԝ/�A�R̂M���4Eii�j���9qK}G��؊y?'Y��Fi�I$J�L�!���B�͙�&5�j�H�\4�t$z���oٜ����#ݫ�,����y~8�
I�*��@��_���u�C.Ȇ�2��lX����Xk�����8�[���y��tV͗о�+[���$qߏ�à́�2)o�؅�I���+9p,m��0C_ɥ𪸰���ª�l����h9�_�/��)#I�Z���VrI$�!�:��P�T�[K�i	w�n��n^�ď�Y��˴_�{[X�
v0b�r���d:�0�Vg;��lU.�C���#$O�3_~}ƹR�=������佡��?""̱��;�ӂ����N, a�A�`KG%�	W;YE�/�&���ӂ�j6�IOi��1��V���ca� �=�A���~���m-�:��p�c���O��~?g���W���K܆�+�U�%��c��o�1@�M��(�ڪ��IIe���#���d��<���I��̘�G]�O<�A�rox긹� ��f'�q�p��l��c��$�G����Z����ѕ��U��c'9k"��I���DȶW���,7^'U�1?]&"^���V�0�6��>1��l�㈏й����B�Չ{|��|�\����D��7���ٽD("v���087Kݥ�T�7���9�l�����I�D�@��!b�C�L���<�Y���4��ACl����ʴ��P[�������].mw�U�P�`�|`�9��%����Ι6'X�{�e|�e�,s�|%�{��o�0̄���8]v[C�iÓ %��n�uj+�t\�х�&�{�M}��b��}z�e]U;�������3��	�Y�hsRAW ��;���c��U�aw�~��v���7�����yVZ����a;��Ơ�&�Uo(�
��B&d����<TP�M��`d��Wy��(��h�Ѝ�O"��\�z s�i�)���s��^�Jb�,���w'h`����gw˲�)�=�.�|����K�n�3iA�㏽Pg<M+�9O-��a���[�2����q�2&��-�#�d����a7��a2k��dS'wZD��P�8Q!���m;�t�@ �OZh�oԦ�("qi�*
�P�k�h��F'�;H��V��~Z���[r���؞�� >X�͘���n�ߠH�����W�x#�n�Z�N�E(���L��ў^��>�k�P�_�X]G��J}i��W6*'6YP����-���Ə�N�b%O=YRu&��oQ�+ݡ���CSK�%zE�U�{������`v l"��bS"������	����C�wĜV��H�qd��A�x�d�pSA�1���%9�54o���]���Ѯ����G\�����d����=|hE(<�ŝ'�|����{���[���/6��bG1 �? �T\.o�9���㔲��C3�T���G��:�yl�;��eqF��z����!��'df-�Xӥ_^,Zh�9+�yO�.4�"I����f�i�hJ���ݔ�����[p�Ղ��%>[2�����7|�PƉ�W��}uɀ�.�uX�B��>p��]�Uf�5�NQ�� ���X�4��L� �����$\=���$M�y;]TK ��ԓ+��a�#�^L�����<��n���w�O��1oC9�F�O��:�Q]�#�(i-��8��pY����A=����1"ň�����Pd�ӰE������[����4�V����b�x58O�(���ۄ���ڢ��}Y6r�>:?���#��#2'�r���@��%���E�C�BbX4iD�"�H�o���qE/��4h���&��*��M����6���R@R(���1Ơ�k�˶oc*~�� j���#�YG�|D5-� s�I��V4�h�	;p�U"u|M��H����w�F�S4[�
-��>j�_�t`�T7�X��^=�j(�ofً��0�0����@��)Im�3�2�^��'5�R���e��H~�hjl��C0�@�~����l���O�p;Cx�1!�k�F�#���Fg,w�]�������T�m`�7���O���L��=8H���
�V
�}�_�sz%�B�)�s�'T�؄��l���Ҭ��riN��r��֔�S	`D"G�ZH��);�;��=�}8�1j�Ȍ�����Q.{�������(X)�'�ǩ^��Xk�����تUS&̛��H��?*H��3�M|�=@ZοQiJ�]���}���E�`h�2������c1^dp��8cFU~A�a'�#�ڛ�&��wǭ�~�C�����^u !��#������Q�����F���j�Bj����U��u���	�Fk�����y��@ F�g��Ě����+z��O0�X�6���W-��x�
���4�!F�|� �w�$9�W?�􍢅�MyĜ
{fvz닇��4��l��$_i�ؤ�V���̜ttc�w��OH�Rx��S(:r��ٟy��Ԫ�[i�f�+i�0��`>s-�Xc�H��fV����=~��rNu:;�٨��]�O�m��}< �y���/$o�&�J�z���Z�A�0��d-e6�Q�U�ye��~Y������d8D�vV	Q�;���H�6�5Ҵ��(V lE#�J4�'kj.�V��/r�d�V|�Lc��Y��-��m���@@6�Q��'��/��{�cJ����LO��+�
�48��L��l�"&����q���|���f��P�l
zn�����@�l���v0�^lp���˷�E��'#@�b��&�����-?��s䖕�Bn��5�{���I���9"��r�*$�ѐ6���dw��
�c��ɉ�
ۡ�o��:z�pc�R�P��b�5��T�Ȓ��`���m���]|�(�I�5��d� >}[M�xg6P3l�B���B��DzO���=��>����G�K���%���}6��)m"��K.� Ԫ���n������R��V�W@��	kAxPn"�:��V��y�O� ��r	���dM0�އ?�����"�`m�)�=��&��ĕt�nt�Gd���8P�mN�T�X ü��l�SX�d�h�ED71�u�V:�GC��cX'^G�f�w*���lDmEP��Z�jZ5�m&h+|�����]oQ�������:������F@�����J���F�# [��G���P�8]J��Ǖj��j���	/zǤ,an��B@���:�n�qQ���E���Q��/�l\�8��R���a�)��R�`�!ַ��[Q���?�ak���1@���>FxK1�3��~[O�笍g$������0�������G$\�.R��6�X~�4�M���C�I~���q'�4bJ�F��2]T��2Q�bO_��i�2N(<L6;��7q��馭�Ӑ!���]S;��x���=ޮ�.�?y�Rn5-�<��j���1*��z":EHʂk������(=3�rb���1M����TO�9����v:����Xe��6:z���e��	9ٕ�[\*}�W@���I&o���0����8�7��W��-D0þ�%���b6	Q�虧C�<��%4�soV���� E'
L��uh}�}�J�L�@�P�������h�����MM�e��QT�ȸ�SJ�6�z�V��WŨ��=/8�vri4wN)ԛ��Juᲇ�dU���Cu}ݽ�(�Y�\ϛ��l����.�4JU�.�1��(�����'�JA��BT%E˥�1��j�,����Bp_�(���f��۰������yf������K�C9F�@aҪ��.o���1�䝩���SL��7 J��fN���p��h�@������n3�
�P�DE�!*�N��A3�ӯ�!Gt�u�
�~Z-���K }Ȕ�:C�nwΖ�Q��o���[�$��׃�ZV�g,qF+��}}HUz'z(F�T�B�ې�#}����~B?�lZ�#_N\ X�/�\,�Ulo�jP�|�8F�1�e��B�n�pC�y�m���=�>�R%�x'��B~O���6A����q��x���@N&�~�=&�p4��
^V觧��F����eEa-{d�T��hJL���K����'�2�!g�GWt��l&wTX�S���C�7p]����'A4�l��'�����W���w�ܹ��F�5B�+z�0q�kTr�f@?&.k�M���๳���k��A"���Z��{��H�;<��ة����n$��9Q���	Y�>�c��A1� x��BDH�E�����Ay�Tx�IRu���9�P��T�{`{�N�e�)ߨ}�q�	Z��L��Vfc2�߅�3W�|���� �np#1�1@��K�.��F��/��p�ǜ^J�(b������{����rP�g�j�Z���'��0��CJ)5�2Q���a6�tr�i���0�*ܮ���2w{�K�M�5��r%�����*�[�6��]�`�U���h���c�-��w��K!�e0�3�i�Z�.��(�hC���Zϊ�m�����ʡ��1ٙK������ntH��y����y���/-.�8t�����G�@6V]�(��Ԑ�ǁ\*j��SţSB��ŵD��ߧf2�b��#��.��SAg��x�]�
�gf�6��Ω��9&�&�C�,�p2��%U Xg���A��^<�Ҷ��Sm��1�g��a�u)۵l%�NS��8^
2��q�<F#��lC�L�S ����i�dי���������A��P�4r�o?#-�s�T��q�d���n���a"?�CAͿ���\A�\��h7юk�䮤B�ӣ���Q���ðd,��n��R>���������� `�M����$47)On�d	�2|��(�-\:K<hƸU�c���:����躥k�y.΋��^� �֜��p�Y���~�$�&�vs��4v��\Bjƍ	LN�"
��볢jJE�Πb�����^��Ge�p�0���:���g{��궘٣W�wz��N4xm�E9e	զ���������,�6����Y�Hn;$"i��4X�=7L���B*�G��%A��K��^�݁C+�[���|����i�����c��G�s��;m�k�w�5ǹWHZn/�$�Ђ���[P�절��
.�?*	��g�<%�	��4�J�1����&���{��z��[d�A��s	���x U�H�In�C=����').�R��X�c_mh�f�h�"��k"zMh�fD&�_0Ph[A��d⤿��S��"RK�+7%(t�=�!�����@��� O���2!����Ө���{�������Y�+��dAo�!�|�֖���t��h�6�ǈϏ�z>�mE�Y����F |/��~N��(���o �o�:�.4?������*J���&\5�m�Ӏe�y��f�N8����:Z��);V��$��9��8��n]��6��#��x��h4}$�ѩ�~��g��������]`2�
��cp�X%���.���iB��j`B�-k�TP�����9���+UrH�X
���b8��}�g�m�(l�;H�&��_�'��DA��
FSoݘ�ǟe�5h士K=ݪh�)�pÄNLo&���W�k�ㅄ4�p�5K�T����cN�}w7���F3Y���gL��x�����[n�N�N��?�Cc�4��v�Q�/Vp�հ�A�(]�!o	c�mú/!��Gt<=f������3�UG�rJ ��FR��v ౚ/�`��~����A����	-4�C�9��~A�Hճ_&]���vmQ2T��[�����9�&�^\�/v�害aB��[W�53�������F��~ڵ��Rz6�H��5���Ϛ(v���U]4��d�ۀ#�Ub9.��iR���h
�)�t��D*�`����4�,ߴ�]�K�%P��эW��?/�)lGhq!����_�W�	�J�XtJщ��	Q���,��S����q�-���/�D��v?W{7PN�jh2������;#���K�.s��ud��9�J[�U@��y=8T4��M�T�I!� z%j[��H�ٳ�;��$z�E���4a{��cN�	L�������W�[���x!�d_h���3b�A��y!�̲�LW	Y�ߙ��i��]K>R�o�v��A�И�'�m7cg������k����s/���ٖ���;��()�6+l�[��n ���?P���o��2��+d�_y�+�v{��T9�[v;����M|=x���=�+9�&,����ˊ�W�f�hT5{&O�T��<>g���:�s�{Y��<T��ꀨR�sP4�%�D�����sv�?c���^�l�-��	n�I�.Qe�R[A�6V|�/ ���XF��3WO����`� ���C�vT�U@Z�Bo�c5EN�[W�IS�TGs��5E{/��)љc� ���"rSC�!��G�je���kr�F����t�ڃNt=mS}àwg�&�M�n�3��J+��	��
��{��"�5p�"�h-�f_j���p���"�V@@�x=O{��k
2��{�B�ԁ�I��Dk(PY\K3zA�w�㮿���7٩��d��-I�qr��"����ɉ��¤́����x��x4��Ы�`�^�`�"���[IȀr͗�_��_sEc��[�<������[ѿ��7N�=������#�o�DM�?�z�Ӌώ������Gx�>*��3XO
��f��Lȇn!���A򓾷1�����ن�x���\)Qp�o��fon��[�F��;�S���ekx#�97_�7Z���G2<�iNH4��4 �Q����i�zj(u��Ƶr<�WE�S0q�rWiΊ} �Q�� �K;,D���s��#�z��A�+����˓J���-G�d�op��̎w��� zD�[� D�ep�e����H�N��Δ�m�s�y���)*t�!_;��~<<R�N�ڰ`g��=�J�\� �1e�K�7�U�Σ"w6���������F��+���8����'H�h;���!�/Q=TD�@H4�e�ot��J#'[��ҮǾe+:[��{�rC	,����G&�݂�ɫA�: ���4���uV� ��

���4�=r�8��>�?Xl_�t@��;ݠP�~o��	��1��ǲB�2?f]nJ�`���1v�G/A�j�j�p���������r�-Y��Im�!�T��-���Z�n06�_� ��g�*c`�,��JQR�%*���0i�ָĽ�����*��V?�D�sY���E�|�AFc��z�$/E����G�B��&P���e��������C���7��Ւ`�>d�Tq��Q�#�Lal)H R��KQ��g�l�V^{����r��	��
�2�n�����dMnjQJprLK��RW��Q�$C�G��Ay��h���he�5uc�8w�6�+��,��%�Aa�@sD7���=i@�>��b=b�U��{�E�u�-�cI����C��������:L,
�N�ѧĬ���`L0��T�����(��]H���z�h~�ʋ��M�V�1q�h�P4�"���UY&��� ᳏"��<�q7�@	�x�%���ů1X�Šy9e;��W�{�z��\3�8��Mp�D+1qc�9+�G��lD��(x��p26ϒ	Q��j�E0�$��a��Uy#���i��80j1т�D���o�{����6��F�
q�� ���|��|��!�GG�.1�=�N2EI�m�����a�EM-�	�
G0#.��d`�{^KT0Ql�O�G�0�����7 ��m=���%�����e9��U!؁8s�(&�)�����А�d{����lz�#����f}ף��Oc�v!�̀=��><��3�9-ў�����twTXH�#Λ(��$�����X��?Y����� �&@�`�������7�o�KMC*�E�_�Ľt�E<D�ٔ>.o8��d װ,��n+�����(�ߊ[Di�PVQ·�|�-�,��q�SǑ3�t%qK�<��!Ny
���]�^��-ɕ�
m޴X�`25b�����1j�������>�&�G����8����Q��v�Ƥf�&Q�ղx�o,���:â1ҝE���v](ؘ�Q�xQ~��6S�7�>b}/���>��a��zB�e�aV>h�(y�k�h��A0��U�Z� �9J�{z��Bax.�TK�hp�����F�T#��i=Ld�����n�G~��\2�(6�@��G(���Ax�j�uc��0��.Ć�o�Mn�d��1�ʪ�11�u������gF~M�D� �m]D(I1n��"��DP��O)C.ۃ�ZNp|k��S4�cTY��:�"���j�m��%�SŪ�bh}Ye���F�^r�W̄N��а��D&F�L���Z��f�{j����l��'b�����x���=�J"���h��@��q}0>n=��8�bQ�w��<?	��ͻaU� ���'W�%X)(3�$����ʤ�5��m���l������Ǥ�E�!�?��H�?[C�6�˗��X=7��>�dV$g�e�MhʔChn�S*��`�hNJ�g:v2"�p1OH� y�P�c��,CcǢS�c��lٵ���c4_7�z~�̽��~`S�f��6,����1\L��s�
g�G���;�g6[�T�E�EB��N
���}IX�fXL�HT%���^Jh�(&�vGhd%�۷���ܑ��',l=Ȼ��1���\#P�y���H��=�t@�R^������nA�\�E�_�8�V�<�Y��7T�_�ƈOL[(�B1�.،���6	���IZ�'�ىl�n�6K�U	(��>լ10��ֻ��W����%��Y��-U�dM��s��!�[G�j%��0�۔�0��O+~3M��VE���*��*�;<kx[�ڤ��h#z���iwYcS�E\t�'iNf�;N��^�M���KL���;|��{3�Ò��}�9��	��0<l�����!� fS@��; ���)����Ӿ�f�f6]�8i�}��Y(�p�X�ڒ	#5����i��>��9�	�wPD�GaK4�@0�P?D��\�4�����A���&��q���9��^{7� �	���<�v*SLeCi�Y<x����&�6.eB�;732���$�<+�l6��Y�qTn2����b�u�1�F�z��ɜ������=X�RQ�5����yM�ae����}�Lj����dm=#�t���糹yC1㘘.]�P�$d�l�a\�,���=Kw����-X���;��Ŕ�6�Q�[�T$� ��7؃59M���|XX7|[F���mMm�|�`K��u�����5�f�D19b��Ԙr.M?��_v'����2+����D���N���˕�K?J]'�������N�岬�<7�>0��P�iD�и�	�(v��]��[��
��zj<�m��������̐t��H'��&�f�p����{��K7�N�a���2RpR�2��#��F�u��6�MT�sD�N�pK7��dr��Q5�[�CM��Źנ��x{šE�k�el���C��=4�bp�셒��IB��'%�阎�i^lL	�l�����~獧i�Ӭ4M6K`��:6AL�>���ڥ�|2v��1\�\Cp����Zw|�s�X�V�Ra4#H�<�i$���v�.o&�t�H�=i.�`(�V�zFJSALκ`�7�o�*�`��5�re�ҥ4T�����/GS1
8��7�ȁ�\�>B�k�$Ӆ�K7�Fk������{�ܫ���NB������������6 Tڮ�%:���=��1��jt+pJ�ҷ��!ȆCoR3Sc�"�� �Y8���.�א4��b��T���PF��ͭ��{`͌�%]�~�S).�ɠ������!*g��h���Qsfh�o$�C���?�G�X�Xz�㙱����,�F�Vb�:����UC}n�i��\���?�GaI��:}r[f�.�,��VR�CM���W]���i͉�O��ɪG�P=�~�j^2�{����&W�&�G�''�q�C�����b�"W='D�1"��ϐJ�*��d�q�����<����P��aU�8|S5�� ՝�k@�{{ð�����W����o�[ /\�{�NT��+9:Jn<��Q.!�.�<�G�6��+�NM`���!��\�|�]��]L3뚑�a�ʷ��;|H~+)asS\f8�j@�8�1�	XD�t�:���!bdE�({o�:Gޛ �����ԓH�o�E����*����O9�I��̎��3Gc��A�+�X��E�l�����T�>u�k�.�M���Sh���h�Cåh������F��)N��&��;��)GO�G�̭����/ަv�m������m�
�d0���E{�.j{�a��a%"p���A���X����L�z��-P��"��c��h!l�9�5�N������rSe�hG�&�����`" tǂ �4��'����:����작ޥύF�F�EAr�Ky~u���C��K!|��<�I#jT�I�zzƪ��M�y ��e�� ��0�u���BP���,N^���E׸�����s�Q�w��ζ�$@�c|ޙ��m�c�ɞa�"�V�� �٠aT�$�Ka�<�D�����sCa$�I[8��u�ҍvD_�����X��tn��ͷ������L��	}FR�uyδL)�8/K�c�[��T��>@$'Щ���m����Q�	*]AO����.CY������IcO�p��#�w3���4�k"��a�v��{�����\k~�r�
4��\υ�*g��BEg��P�:�Ա��3<y�8A(���+������	����Uy'�d�J� z�ۦ�4"�8A7�\�lFO7���Z=����v��)/�ph��F�4T�Fg�2-�z��ޯ¿������h��k��:�!}b=���WK��8Y��ǎ<;�0��A[[�K���/ �r�ƆŖi��ͳ��Q�V�-����p	�j�G�kkQ5�㡟�4@�lt'�-���W���}cJ����˯c�U@Aa��Ɵ���O���4W?�k߅�o6�u�,�ȏ�D��j!�
�~��!`��퐂�1��tAT��A� ��qe �����$5Js�ҏR�(��=׉�
i�f�).d�+<���|���I� �Tx��qe���I{#П0v-%_o�V��$���ko��U����k}"'��\��w:z�����LC�PjC��*�Gsݶj���£�tZrQ����F�n��)Q��n��`���l�'�@��W�Z�X�u?[૒����*%�6�*���&L$wވ�y���u�I�X&7�N��e۽$nfg�_�ME������vj"�?�E��8�|�s�6R[V�'b����F	SV�{�� �0G8�X/C�8q�P���)�#�J�$�D!<�4�4<3�r�P���0���$lt��9l'���qߖQ�U�B���ٍ�2�T'�UO6���T�o�j��V���i�7)��j��QN*��z}I;���k�:��R�2�} �]��>�随��4!��`��:Y*���a|.Z/����i�����[a!��d��̌���2��zdK|�e���kD�ߧ�+L�I��v��'�nUQM�t��J����a���]g/��+�`p3#����`���4�Rς�
���u���0\�r�G#�gK"�fbՓ�/�m�e�$!��{�⼚CM�1G�s������d�*{{
�%��4���a�
�5	z;�l�	��S?4�!� ����c~&��͝|[�#���PC���Y���+|��vҁR�B,&JƢߦ�J۝�w�C��^@L�9_�/�� ���Mѩ&o�O��u�n12�}
�2��١u����hn߶�{`0�^g*_�Yφ�ч�L�`��yU�P�W�d<�qv���)�4��~�zL��_�\2U�Bx�	>�ۀ�\8�`*���Ca\c`���ҍ}��1���o�V_��C&Q������kk���X.\�)�=����EKK���;P�h^m-zz(�X�3|����u+���m��ē����elB���b�+動�WFV����w(UN�\�'�Y�i;8�.s ����-O�4<�9� ���U|���/�.�I-?���5N������G��
m��yM��˩=�u��AC	��D�>^9I��d;��,
�t� �j]L,��eA'P��O|�*K�L�T'�}:�s�^}��5\���a!$^�� �W�P�l0Ơ'1�Q��q�
���V�~y˔�'��8?Ѷ���I���X�������`3`)���4ij��L6A�R5�N�bp�4����]���O�B@L�3������7Ƴ�^]ͦ�iR�x7�8f��x+!���(S�ҌTB8�|��:m)��|���>�6��QmK��0/C�-�~��L�N�E��q�^��q����,�.LN�)��A �7o5/yfso��H ^?�K�L ��ZNYd��g9<�"$ Q%@�`��4񖇐�q�]���d��`\���yľ��ACZ�����~�n� ����m�n�Ne��h��C&E��,,��"ʿ�9i�JΏ[K̯}�����v��H(�v�)@�)����8������.Ą,�dĎP<�d���c#���W���U��W����Vͣ¿��D�8�>���ON��Hcj��/�)	�y�e	�U�m�w��UN��GC_~7�d�h�EoA"�5sQ�����}��^y!�yRU����A�LIЭ�M��2����&5�4j������ld	����.Ô����k��/�T�
r^{�n&�W��=�/���4>YGy�O2u�:�?ԑN�֕.�-��*	r�a)�튿߆n�0�*��Y�v�TF0j[�?ѿZ���u��k�����替O<p����3��h��N|7M�v	E_�ą�S~��,s`3��\�-���8'��^����|���N���0/��D�$��%�s�n���a�����#q[���d�F�����X8��|!��O��a��F�~;��#mjty�Y�Tl�,?pe���|<N��ܮ`�`3T͔��
<;e���$^�xx7����znΡ�s |Á��`gB��~E�&���B�P�M�u6���k��\j����=U�l��u�4K��iD�(�/3 E�h���
�7kˁ@WcL\n�+�·]�ظ�\�������z?aʻ��e~Ā xB���e����5�Z�'�;
�<�j���0	�Q�aO���Ru8Ɔ���d���f� �;rl���7�nm�B�@��]�#�%��n�r�Եz����ݧ�9��;���?ⵜ=���=z���l�)�r�����
p�У%�B�!J�t��R�P,�#8yp�����_1X��(�.����(36v��t'#�b%'��v�
!�3C�LH@�CM��(�>�����D��;#�� Y��O�ѹ,>~����������;��=�wu�-Q�3�؜�!G�q��[U�#��p7�1c��Re���V	>A	ҟ���	)���]���(߁�i͐�vB�I����P�+�����E�}�o��˚vI>y-�'6s;���)m�b=�+�e�̉��>�.(��qE��(W񿝓Vq���w�z	,_2BY���l�*��S���L��@6���AӚ~��gCV�����^obRZ�~NK=�1����)A�.F#���G���kꝫ�Ib(1����x $������ό��`6��kn;��!�\n��X���eG�˙e��@�8���łLW����0J�>���I/J�Xg���m&�=����<2f[�C�g�@���L��$��.�#��;�"\0��xXh���W3lie�&��^1p>#랬,5Jx�!�|aHL��V��+�JS:N{Nv���I �U�vme��'N�X��|n'�-�V59��k�0t}7�i���~�v�Թ�k�	�u;g��t1�Y���冉��7K0���=��HHʐ�x�P,�7�Q�hZ�T����T��)Cߙ����P�O�fA<������uLs�m�c�U�k�<��w���ux�>��z�9D����J���`�'�qϨG�_�^��G�����N�q��aqH�Ũ�du�u�X��_���5Z�H�[F���ݿQC]"���\6�UI�[�����_�Jxף��܆Ypk26*�0KzG��>��o�P6��ڽ�ZL�
`3֓����P�_�'1#��H[�;�����[[5y#�\>hA��f��J����i+�hfؑ�w_r�؂q+.)���m �`CY[�(�_)�O��A)'}����ܺq"j�q��{���s
A���$a��k��nr���[���rD+s#-��J�@���+֊��7��`6�~K��hE�H��:A�W��DT_[
���	��:���6����� ��I�m��E�Å�����>�֣<cs�`�C�g����x0�4ҟ �S	��D�׻�[�,�e}ȃ�]�B>��0'q¥���o��ŐtF�v��Ly������9{���:�F?���� ����7�h�LP�9�e�dȀt���ަ�GN���'p�N�t3,����������L����czS܂@r�7͒��#b���y4��a� 0���Z�J�F{���I��\h%{�pg~
��cj����$ W�ы���cr�B��F{v���W�߽G�J�i���G���u�����πP�	��<�xXD��n��-C�3����a	���B�֨VT��׶�p2h �tw호�k(��P���&���h����l~�|f�\�&��Vh��F�_ 
ɛ���p�v�t�i C���`��RgT��	U�����XJ��� ��^��S@���;e�nv`h�ʘ �c��I ���I�b����G��­2~�h��G|M���
R���_:�-Dyl������Q�5(�*����n���r(�Hܞ�Õn�ԋ�M�W'�"9���C�G�a���Q��� �LT���` �d�&�l)�L���w��%�-x;��g[�&<�Ci��-�?�N.�7��Z��H9/ZHX��#_�B@;o�yt3�(����HN�4��{�����ehN�mp���60֠O�z�I}¡N7�y"�>�AK�"��-�O�Z+1{j�#��F�$��A�s+��luFen
~ZI�1��Ǿj�+t¿��*�M������v����~�-�ή.b�@mo�/��͜!��^�r"�4r�bp����Fh{�����8]L�Rϓά�QY]�v��q <^�oQ�R��ز=�k��(1��E�O��=���}�<���+4��u��>i2]\�@����ڛQ��)�ի����L��
e���눙�Лs�9ؼ�Vg����;t0�Z�9�8ǜ����"�
C��m��4;�Hc�W�r����V|5DY� %���-�[vv��R߿�y�K�bw1L�1���@��%nbw�N�����T>�е�b ��4�'���Ι���8�5���*���A���z����ۨ�e�г��s�ԑ�	�i�!
���x���' 	��)�'�������Y�X�t�m��pZ�ֽYt�R{$b՝FI�lADQ�mM�D�Ύ�����1�5Ͷ}fOE�_<IB����d41���P5�[�����,���ِ��Ơ�2���B��ڀ;v��5j�Jy{��>x��7��mNs�$T��$���|b��u��m�䠓o��i����3�8�4��x �Z���zuW���"+FFW�!�����C��:_x14�����6q%6� ��Wͨ'�9�u��y�PKw!���P�%�rԣ&��O�]l�|k�츣��"�@�ݝ����ަ�X����f]�o&~��6 �fXH�;�m��Q�E��J&WnLf���.��m�b����e�2D��C�$�)��	�1W��3�x󪄍��v2Fw���pU���Y0Z(��(�)r>$ְ��Ȕ��~��#6U
g��@���ۯ���:��S0&�p��&��t�T.z�-��V�!ibիs���.�ws$�[��E+>�	:ӛf���~z�Wi��a�d�� ����6{ea��$-0�E@4Q���%��nva��ϝ�Zӯoz3�U+o��n@,ة��ͭI�N�$�ח���	���x��M}����8�Tp����	
s9{?ސ
S�2�?��1���|3�S�N��Y�k����¤�y�{���P1I�Y�����lm6߷mi�χ�j�im,Q9��,#��"�Z��,�bj_�qV���'���\�� �q��O���1,m�ұ�#�j;?	EG�j�~���1Y��4
�x�İT�Ñψ�D,m��*�x��I�%�/�s�Sz�9M8�>��뾄����fڀ��Щ��-��ȉ�����1��IݎӁ��s7����1)Wy0-����W�X�40�ٕ����?���ݔK�4ꡀ�!�gڿ�]�g���~v2���eϢP�'�[)N'Ʃme���"QWT�w��s��r>�<������	��\6D��%��
zq���] ���,[�+#R5�0�Lg�+/��T>�����g�5�֕�%K�
$����{ӧy���{9+x��a�:�(V���:T�뀣�'/F�^�J�}L�T6�=β����h���S�!4F5-ǍS�t%?��W�&�B�-�ð�E'�����C, �}�2������zh�w�N��p?�9�[�
}�v�£�/������_a�x<ޫ��J��L�z��,�#$���*�OQSk�9�������cΟ*���T����0�}�*~%�O�)�2tڵ}��7 � 5��>��cٽ����<�L1sŶ���b��}%��N,�V%@��k�W\B��ƘB�4�@1�,�-���0u�ͽjp�9�GS2(b]�O�Z����"z{ ����B�N�ѧ�}G"���xr
D=m@� ʹ�tC\��V�-���m��wZ�?$/h����̤��)�y��ܗ�U�X���5��8��T�_�9We0�V9A�-�N��Q��������-TS\|�ܸ<�W��N-Q�ˌ�h��J͂�Z��=��U�аu�2
�m�G
8:�h�Q�6��R��e�`��3�����/v5�+G�ظ*o���`]7Z��/<��'����mD|׃R뗔Z���#5�� Rnp�@C}-�_����hMH�>�_z�{#�+��cP����Z������L��~,�c5}R9�1�����GWk��g*%#�l�ڟ��>��6��ޅ�]mqv�fM� V Y�/���?�X�� �wm&�$N��l���66v�vrH�X�pr���� �}r���n���l�F�C_�K<Ta��^��sR�:���C�,J!tCq�6�Wҥ�Qq�2ZK���9\L�7�N������2����WCŶ��@���{�/3#�ӌr�u���r\z�5�<��~�b{�(�`��mx̝Ex�ɾݍb����Ϻ"����:�$%1a=�����Sg��O�E�OQN������'���H]�W�7]����SZ�@S�-�|l��ӟ���Z���;�i�/Kި�L+N��b������\��,P�a�@*��s[N�.>�L����u�:"$�,Q�S��Ⱦ)���]7���E�$0�iY�yt$ӯ�u�T�O�~@#�G�n� ��siI���Rgeʚ�HJp�xki��j����~�`��Ci꿍��A�Ӌ���D.?��d ]��FHꍑ�B�1��9�O���Ra*�)+��e5�l������4Zl�ѵ-��,Q/q"=ei�U�`d��BW�5N�4>�XH��	p�P&d)W�Sl��������bv�<�M%��0�+9f���~�އF%4�7gs�&9`�����W>�-�LY�4���-��v!�@'��rR�^�z����&���_ڐC���%\K3��c�@!E����w}�l�.��HA<X�,=�����0I�n����)���6H	�F܎ra�<?3&ݓ�S���)-�i��L�a�j������>Zcұ��2e�^�A�֛0�SF>��J	_�����P��2BD�'�p�n:/�L �\(����z}3AD?D����U�ߥ�|�^1�ػY�q������9��S�sn�?�D��O��W�-��7��j5R!�S�
%�(���AkϗJ!p��!�"+7m��Kx�{�_��_��������G7>b�Yˋ�7���}�6I�l$����k����bj�k]D�YT���V���؝ӷg�`
��v���6>0��xP'����f|�|��3��������ř&�r~������m
c~r��	c��?	(�G�5u�ˁq�'��?u��j�y��Ԛ<�~��8����я�T�
m�Ӣ��r{j�~��w����!,s���j��?D� ���E���ղS�l��j#;���W�n����?��Y�1�H:oL1mJ�a 	��\A/k8p��_d�h��
��\/5u�)|�]�dB:��E�{(�9��H4�EE�{�՟�6��s���;щQSr�Z��B��H�i���`_�O����:������P���#��ׁ\v^҇��`�uZ 8���Z�?0dʼ�0��`�!oy��q�yb؂��;�_>G]%'ք�..,ꛝ�S��h�3nCf��@)�n�{O7��N.y"T1p�^8�F\��I`�i���oe�Yɀ+�ʁѥ��z��a�}Vh<�O{���zA:�C�k�o��L1
]*Ռ'3�9�%%:�E38q�.B���ǋ������8#5(�̮��.T|\���úT�����G_Thp��G/4FȔ���[X�!���f����|`�������`U;��Ņs6&@�0<��oGjnuL�gm�}�޺��W��9����Ҥ#a<�F(9�j�))��E���ZJs��`J���u�3�����MzC],yo�ؾ�a�|Ap,G]�M��oiG�_�`P�'|