-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
fmhCv/a6gkv9rJ3qVxXKAphCLOyyk+VmrRFLI70M7dcJhLzhQ0XbKjjrIg0B9TwWnnEjRR2IRGNZ
LgD/35UTk+AyyVfezg17ifE6I3ZVO6vW5zFpY8PFRZTU2UmCWSMUwrj1d53ZhwkjPyw762MKh6F3
lDjURlw4rEQeYxDMLqz3kPLrnKUkaypp2zUUtHxr9HwNSxarHVv+0wLOXsUBWvN513wq7bdcMqIv
yJIG+v0cjVyD+fusxU028y4OKqQekRYnBKKEJOAb6lfKPuDW6+hUJPwrv7Vq9629pC+5H++wFexB
6QRSJvkY3df1rNKWQZs1U0Q8GBcxY3sQZrz+kw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 30096)
`protect data_block
ZtQUKLBqWg8jP3wUz6wUcF6h7ljcgw/ceptA824K7VF2mcK89Qxp3lOJG82ZclibV5XCusfUgAbf
08h46nYwg9kAHzMhvBbjoAogMUsYS8ykbxuDB+FdRK84V4G9lJtyl12GaFa2801MLW1KfGXpCegN
7v1HnNyWl4o5E3AFBdraHCavCRcz3jb4JltqgoD1POX0FEsU+SBiM1BSB6dXVXbKvVPL0tNAPvBy
K8wWO0upiD0b3W1Gdf4iCYm4M7mowv+1wghHUu6SkzU4C05UdRpxwvNPQ960Q8wkpRJJm2mn7rwS
qk9FGptVa+kRgsC9BrvJdVcnNqPMp0iMrqE4BT26n+B2oVu12BFhsro7mPy+1f9RE4/NTWxfVtsO
BPgQpi1vZzg6QOI8flDY+WMleBc9OCoL/LgW4sW8l7xxZEI6ip+PCbvcRKsxo8W8RIkC/czcW+yc
KPnw19TMnnYcEe+FtOb8f/k5HLAT7Iaa2E0qUooMNNBOStdyfXCjwy9EzD1uLFvgrsOpX7JEtXyd
zTyycCQ+JyUjZvptSGEwH3mC4BKgfxGJN+W1AVtV4qy9iaJl+hznI8ArQwIcQ0LUD4B862PDXeQF
XlUsmOTlZ/62snh1dlOOgys9wuDMu2NS11Rsf+ON1MnxnibHkCizEdRD9SuEC4lGLwKn6EodD3zm
mq5/RNfVt6Yoog24gxr8hgdwkXkk54Jf5kOQYBTkDTULFbYpazu+uv9lhwhMX3twYb0DZT3J5Hpo
vPzt3F73JoGUgyVbb/qOYuHEr3fWAMJQzcneIOJLYs4XHAfw6mXpybmVRMr9HlARJQV7RKZJzxL9
eCFxtRt6C96Zt87Exzs+76SDXBoH517aly+CxjOV9gKF8AI76+7Ns1MjDN7EIvYDU/MehcbrbJ0B
HGHXZF7aQUENt23qzylveER744fOtdOexPijCsv/rMeovqWaD43XtrUARwmOm398x36YgkPIDHk4
wmrYDiMfP1LOwBoFSTt+nol/r2P/kKSgZwV2/XmDRX68uy61eKwg0cYYaYIZu18IUy5UH3FQ8h8o
TW6LDOFzwNZzCkiieOEbn32CD0izhy1N7z/AEb8ena/MMw0t5mJJlH+wnRsT/Li5LiLP8ZXAz+4A
eWHH1/FZmabU7lg2NJ6MfhdS7Pwk3aE0fqOA5C0Zmmmps1X4SVAhZAOwluQIobCKZ4XGc90x4SKh
6UnJU0iSXKpltRpGiI5FkOz04V5oB9Vp7U2Bcq74Tlc4LU9t3XVkz+YXRla92zudwCNSsvcmyW0P
cAlojvvT0fD8Qpo5VnZJgWC3aafjfK7Zl7cHtnCy4IDvms1JoMDWJdWBCD0A8mXZGFL3OH10xjf0
MCK64v27UcRvw1DuJ5hbVuviPcd/RFlybE1yMfZa/xUXGeK8f/HDLhlQ4Ke9VvnZUqrBWW52iJ0L
/LUkIbSgTx0QWBln9A/eFbGX3E7YuLjggFYpF553vRtPVWHTOvk94eNvHuvDqyOSRdmGd1nlDKm4
86Y3dvWWR5jXrrFW34bh5mqp6Kb1o7qUX6HoIAkNDgVUEVz0t6PUIEQmtKi+UV72Rwvd5IzW7fLa
Lz+tGqnfxOZGV+qsNas7ZQ042j/v5EIB8Uag49Kmu8Ly0G+8wq2qXYI+/YgOgzbma4j+79kO/NP4
INfp9cJdD9dI1UcNsD1PbcHkDFLJ0uoHF1YvVTVLcFlfSSIKmGUzwOeo+zx2hkAjO0EX1aayc6PR
qcPt9IZu3kaipxCfbhWsZ8ie9nhi1F+CGik9eHIrdpOx7lco33emHlB4cMWp16t/BfmmqPprjYV9
3Ud3vPMFUTJrU++1LQsYQ8Ahfr5uoF2CxMqPM0U1yRwHL+RA00mv3fnKPCPaQPr7+Jkd8lGSSrPJ
k06DH0gk7jq8oj5hr8mOtFYo5rtJ/6wWEl9NrYZ+YfmpIfKGRnWbmy8Mp3W98qdkTMWFwp4iKqxn
CWOZUln52UmRIRgJhHtyQso44jR78bRbwYGoueZ3gL1mnBZRKNtwY6q1vC5JG76oWzV5oePKPFwD
0i6kVyyRJR6gMDnVqPSJE0Cvp1wKmu63ON8OsT/5bCKjAdtrJ5huGvPdWLpBhWVbIJMopVmEP3oR
6garSs3cM+LIteb4MPoM+O544FESYUkKul1JOJ7Z0xwfqr1Dq+G8ruV25fpKcC3O50J1VRjeKEIa
kir557T2fo03XZaKMEP9jft7oqUWHLleBqVZfdnRimMAXjiF3tsXiXd7rLa4STB5x/N/ul5kdtPv
Yjw7JkQuxA3YLoSPSzoUqcy5iKL7xrnzzznvwC2E4LHRB/Lj2SJUjH/dCl6EoSVXqz+/qaWOylFO
sHxIHEsLh3XjrkXU+66KbMi21HHXMX1k8h7RSb3Dn8zwnR8OTQfFUWvkYURTfUvJsRE9xW1/qopV
oJhCqskzYSAp6QxxfJ2pGlfZZBfnhkwkcaeT1Yg+/MBruWxvcbTZMpMPsxAsrhoCSBjYPw2c1L9O
rQ8eXTANLpt7rAJTiAFnwzozJ/UK6ez+cMG2KklDbUDpxW3QspxDmpDp0wS8CIRA7XGiM32jYMCu
bAnUTgFlEva66iWzL1T64F35TxF6yTYSEsMrp790UvNnoshqBtUr8rjtzQPK3vEDk6o/kiMw5qmm
cFRlSQRwaDh5nkLXT65iY5xh5Hfa7cwfJML5yf66/3A2IOnt/fh9/hmXYQPixThsr8bjayPr9t/X
h2AGgEwIIShOB8u8FuRVqeUBXn13uip3vwhxX04UFNGYllYiwDNOtGHyQ8vSa5iJfomY/N1/4dHu
PYFgTxoQ+yaC5ATZEApLUjyMJW/Ot5OXurRbDEt6CRoOOxZcegUms+jaUfb0N6jFJ2nbBM/BmSfq
7VWar6AmDaltyUvIyYy2d1ScI/8v0srF70T7OvdfRYpFpuOIYJpo3bEdDFkqhTXr1tpa6A7szmyX
Y+LZCKkNvnPEIbfCSpaXgG4h65vBNxd1QiaSSUl1yQV4I7Dmqh3LuacW/OfzINJJ1+6OZlT4E3Cr
CmByuCyEeWl3Q+ORW29gOBgPZygYXjhNRhNEjsVLUSKkGETzOl36dO9eD/snMMY4UvdFc9cnAFSv
rnL/F6WDc2QQ/j6iPTLOTwtJwFvckxD3Ve9OmF47RwHeEzNxbASKAL/1RJzr1VNxpnk5O8dpyTbY
BS3BP7viY9nmFCKQ6R9w0XCoxFrFgwPOdE7EhvFJ5U4jdZV0w5p9/2+kbOhtCekvywBwRhYAzBf5
bE+U4R5XO3iIWwUjovG7SDpo88AZ/dWONoWDRw/4K2xXe8RIZe7qsuBwI+f4hlgpxv39DWSjs2Ac
h12KTJg2Mwfa5foxfDxW53da+fL/KSpU9u+wp8AlNtV/Lt+dQg1lkKvtZ1BePPhop3VuXDmaHl91
ScPbwrqqFg4abUP10Fq+SyCdYDw05cgnbTnrSoDtvkr26kWLDqUev16ibLEFa4kQ7l++/J/rWWGL
S5RMB/kUcHEhFuXjgsLrs+jE2BZ53sEOi36W1whpScNJ/4CZrlK0AfamL51foImXjygFDxI1o44Z
dB2JvB7lsqblbsv25JsNUfYAFi2ay1RZNzIt8HO5CYbfXM9u2hYX0H9PQU71ESHIhhDzoRVbzP+H
KaZij7NNbTz1b1gU4nXFWGF8hHnl6hgEQp8wGyHff14nmH/LrgaxwS5vmLdcnaugZnildMWw8V/R
DoTSMoqoIEo64Dg9cuz9D+1aRBCS4S8fnlbwHophhzno6PLlKEwotJqxduYILkx6Amr7qinXN2Lq
GpzMDEDq/UOJneRwvhxUaEFic/DXXaeIvDAM0cRKaYwI5GI3mRKBVCHporEynb/kuwUsNFLs3ToP
9aYr7/mdX2QKCRr73MRmvXFG24Xb5YG94Jv74kOCtBMwHaEb0BcEkPqdOcRbYNCbGszvvP3L8DvB
CJDqLBotKqFOd80W+vk/nFR2OWbrxK0l22xnka6qrqLd311Yk4OeUaH3/UBnxjMAktJ2P7e++PPX
tl5uBkqHSpZxXSMqTo50T6kFnJJrh6BJdDO0oaiCrTmC9whe+UJsyjy1UiSW4r8FaHCQjK6fYSC/
MNp6q+GVTaDOVK0PLmJUpj15jpwdg95baWiVwrNnsLoYc8bByJ3rV0uPuqhfgbLOqhekBqEYg3jK
mqrf+AErF3jf9JHShXqfAzPoGUPDFQOSfVwyEdRljTDYIjAQejdlAlwVmsTUQlsrfHenOVuW+PFl
hhP79IS0NH2Pb6BZPe6X1jmvs/usB5R8LyU6K8nV4pOgk/a03QWrgzd1TEjRlRn846dswUlTYHNH
bthUAwTndKIDVv1hoj5dxMBfBxq24tdqYRp7gvhtYBwcD+irC2HZCOxPygo++GoekUc2YaK4OAu9
OGN39mMAyWDcgqWDbsuGI1cT3AlmtamsTVBqiXOQUmov4f77yRBdglyrYoByNEjsg9d0luRjX9Bl
sgXTXJCvwcbZGn87tdZfgn/BlTQ0vr2s/wWrjAUpmBTrp9LCaCAVvKV5y2w5HwC/Rs2ESSPVjna/
H5kdHE1YgdTYb8HkRLB3ywbMkc3EoGhgmhXYWHJMGDBqB/TWANJo9dCfID39TZrHMKnbo3z2MXI5
ZqgaCeok+FY723ldbVWPqTDnz8CjmauTPhAKRCNJ44Q6Qnayt+yiUzIX14Yo/+JIPQYUYddwWVzL
oYtWdFmIGWk7IsIML/+n1WAl7XgPgWlFGyzewxthh6DIUGuaa5pWam/QuFUE5p8HU8KRQtA+sorx
508ZHMyESdFIqLL9WO9zmPxZjYylVIh37Ki3wQ+Geh0m5covkuKM0zs43KgupOzDb9fiu4ds7O8x
YzjLpJl7NU1tsYwaST3rObypNYdMA6rI3E6RbQSIzyc0UGgsGdbxazuv3J93oP63m/GNEs+g6p47
HxtDq7UOBgvMlXiLyNL2x2XLL/ihrszr2EHpbncbX5fOFvWbUCLv1vcmHJK/VSdQjYqu7Ga7t2GJ
Exbe00siKbbXgHXwVt+EdpWxPIZjux++T0xaVP/Rn+nctGH0mrOAA3Suf6Uy3uQEZe8byIJNlC5C
8zjJxzkQivApSKnCFgMppjEjMZ3mBBqlbwZkXcP99XXBWUGDUhQtsJEV1wwPDXLJxLLvcAoUt7/v
aR5nIuBQK/LLXhh7U5yl7odi7wvTMvhQ5yiYfPrqgkA7WOMkeegimtCt+NH+t+y04EfjItju69zb
SDZ+iyyjtxtqZ22WXkLFklDfT9EONc4ZLnelNL06wakVSKpOd4JjsfwwtzT/zTeJy1RZoPi/hefP
CYGFtcrGBaVtsSHa0Ik4rH9eFCPLpqfpiOYmyFvGtuwxTwNcAyBmp3adAPotU4y+k6gHtaLSz1oV
6ZZHD0JIi7RAa8KymUAAzrrwJp6aE6b81e4gcQXpyTNSQdAJWTA120gr2s+JJsvmvqFTlm8CF7A8
zsTh/QI8hpkoR50QwqZQQv5TYriEeZ2B2VzMOSvHZhmaMzTA/OXUW39b7z+d+zCfSQa9BmV16EO9
Zjjdxqk4DMIypvp6e0QW7LxUEeeqsKe1Lhf6rdaP5LTt6DM4uM66ZRDtHdCWD9cn5MjAnivfn7+8
tUUWzQBsd0LQrIPwv38vaI5wYvAUoEiCzaMd1NE9jXkosOkc1B1VvwK727g0McHLZrNa2tDbb5v8
4vyvIvEJkOjmxKXHCyHREfXw/yxUEAzvil+wUIlASXqlvCyuAafkdPFJ0W9hjcPq6CE4ZIgSu7QR
EMBJ9CYCDW8Z19cXrIPFKNsb0OLiJNP44dFpmYnXNKtEVodMPIPdBrxN+8mZ0aED1tpWYCI7j24L
7Pj/rSmKe9zvMNyplkzeRlWj1vWQbrcqAVNV/yOjBFVHxgAy+tDbiQpiXb5vbm8kTvhhEvz79C2l
MNLtfXJ6NWNtFKLcVv8xIHVGmJPP/n/0ffi+YLYj7PnFlsLvnsniWU55DxPqowFZC1GgYizOqGyi
LsFyC3y6bpVtskIr51BkiM8UfD7wmVpa3baTGSFOmFX8jBdepkjeZGpfpAUsugHNR50hh6S9YkyK
EuZu61JROqRm1iTM/JhaJvdysUqTcuU+YjGmoI6RRiuBNJ0nI+RuqxSjTfLljQPEq/Lk0TWHRXsK
DTc4T0XQebf6bAtOIGld6WFJfIyDlEvIuNj1y3/rT0N1a8V82yqKBS8Pd96wPTihkjk9M24f1/Ht
pDsT4XtkSd/3iTtrT6bNW2zTshCV9zsUehhZKNCqmfQA9QsNAjIA3Qb3hUHJ9eLcimB/rK/NxAwG
5UJ8QucoCa9VCeYza26IK+P1T+FB+0Z7mByF+rvkRLA56/dNCKmJFVotqPbBX8HRkds7sbAdzSjx
e8seaDoye+DEIyIeKYiPOE9vbfvBbooTGA8FB4jA/mohu1yY+y3dIzR22ZxU+VuxEBJKLJNjtv7+
8+GBKJp2pJckCGYcVSioLLiMrb4j00L20SSXtmNXiFO+drnm+3TeJgQhMebNxZjaw4VtjOFgR0CP
SLDRUjOZS8UDDrqvkxhriSrgjm85J5hBJO5YG1p3N/2xydb1E3tg5gTlkCi93l95S+BKa/eC0jXC
fqlf1Xd/gqv52pr4voPDGhqX8FA9TpRYRROIbEYNYjK09FBeBfJE/hzG4Iwj046DP+Wi+xEABA9U
iTxtveR5D9qQDEF72BaWPo+TbGhhPO+FicNW8peyPiCpGIZOwkWkkOFXLTXiyqTHwW9vJ3eiOhJT
EV4VAcXtEq6TwwNBxy7xc1Gix4v7dPpJ4n4KJk2WLfU7/L1H1aoInJXZfba4kMmHOoOH9qLHSwrV
WtUnH9ymcUMNkywLWWMG/jQeU4kVlSZoVx3GuypiwyFNqz3yyxlp1epVPUFPoa3l4ZKBcJzV+Jfb
jFQObqFDqCUGtD//lA/rzRIc7AVf67IQYXNhswedgPqEwhLQoZyOyY6PMtVEQGDfWvnf75bOryNY
KhYJJTK6M87F1lhs9QR7XnefQw6/V2WGiN6t5EUZ3/53rJNb4UdjZBuMKZRymaI47zvOwcOxnUW/
Sq8del6xLBaw1o0EFzpGRqwX3RHQcfjbPFkkl4kkO7EEGyoog+wn0vjSPWf97AFZMSF3bV23vc6J
+S1FPDs5ORgth9UOxZQV8SYOGZoSgiwPvFd5ZTpgcpqHpll5YadOwjIqLoWBMnpFjz7vEiR2zOor
Vg89lHjLvm6FxbXEFkLJ/I6AOtem3Jr1xsTRJa4D4SaSGqaFhGHnY8ZrJj2B2+V0KIJ2/3QLy/ZK
HzmfzVgaxERFlhMLYJXaqzWs3oie82d0ZOrRiOMnARirTBSrWAdqV0ArPrhqQ2MWRurPpE/ABaJF
iQ5TISSY3Q6OG/tY3ADstgiz9UihzQ6Mw7t6MQaFJY1EerVeE99iYKKtqum91XuxVLuHH/ZbE1Jh
XtnjyXbNUSiCpAjB2ULjxlKHJ9WnKLT67k2S6iUnn3d18i+E+Z1yAo7bQB0Tj+5lyhzxHpdnGKmH
SaqP+cjUrsp/nE+ZVKMjE9R8xThPV+DPzMHo/oRtn3NkODj5EWEf6INCyeLqQeWHdk55DjoQL18+
/LtpQ3KFcr3P6bloz8oPsNb763MGjKwE7Izs1XL96Ix+fnUVPZoMezsIk9Dq38t6LCcTUfNKHZSv
OsdQbD/2vF3+wJdJGEo2+utJVgd3Lkd78261flsvPCAdyGCoPxZ+Y/T3BxAORliY3xo6XUqgp+TP
5O51ZC9n1lCGHPt3Sm/PKmYheohAFdtsg3pEln3bzBTIZIn7RXeSMY3/oHMQuDnNTi+ZJV8cvVCb
xWh8H3lqpKJoT6IofIwpL2znUEqxcx0kbq+iK5pKJu+X3kVsV+620ba+B5QsCxuI19nbtY6Qe3e2
SNnlUJyyQi98/oNn1yoxO079cln/jofBojMLhs4JDhpu5a1cVMFAJlSTF79KyCzEvo8teuHh1KFW
7MvP+4/rj+EZxma6PuXKOfNIXwyHB1JJnlodzfz01PBTGtpT8Dj+SJYCglWsU3hAeSfnrEP6Y/XA
5PDsDwe7CxTpR5HyqOU5aMttywFVDwEV7lcLbiiqMyjPVtXYi6oHWveS3h+vuQvTKCnNC5zCq3Ox
+90mVSCGG53YHOiEWItlFLuLMhsOq7cBJ7iCRntkpJ8BQMOmsT22Z7Tr6tDyofk2sIAzTZVVRuhw
xmXj5gHfCy1d2CaejmmhvIVGUqXLu9beG61GQa/vT5FedlA/WrFYrYIvOvBzMZ37PJZKJwZN8JQr
IzIpSoxdVmckPpWd4csH2bsppUDwdbDNm8tgwK4MUsYbkN0HwK1Cbrb5vtsMxTWrnNWMXpnQYfRl
vZeac6BLhGEqeXEemIxjFZCqXidTdeb+MSpaFqjkgY+K4ApoJRfqbrGyWVkEnamFwIQBP2mUXs16
wDt89w6I9efcZJX4xLvNEMIl14p5JSD9ZdRScQ6SZF3DZ4rLl+7LRpsN8Pb0djVy8Bo4w91OIrAu
yzLCvvLm31RRGMt70XqnBAirYjkQv+RdimGUEu1HDt8NzhgQho6X4hGm+6467LA4XZVXqXPDPGZQ
ZtLZlb/87ThoMUTIrOwjnr/9kAuJKZeCPGloSCsqjCzQEx3tmltcJPYFkdvvi/X/Mxh2nRnzW1Eb
iywqp9LB5GdtM9pijqzkVSCESLXS9FyXRV/JFiJ8+WIHcPIeXPkXgyl8Sklx2vVZB9tbrJrYBUqb
xGTNzbIDmbL8KpiSiCW9TkLx5sIBJ8uVq5+eVIsrV9+9f20GFVkd91IlFi2xqZuJDqk1oGHWvBKK
/2kx5rQjEKFb2fIMYHB0LkgXUWfXFkqH8BXuNHy+YD+O5nidguvbBe3801AaxAOGQU1fRdmP67x4
A4aYG3Q+kwM9mZWGq/H2Z//r8VHUwyu4BCJbvhpW0FerzFftKIF8i5kBG3gRmW+A05uG48FyNYnf
GibjuQRwrlsNzjrActIhsB75CSNI5h7J8wY4B47ULHc/QHKKR4ChtKEmtAAm7epuvCPhGzugr7oy
Tg96uvPybvspKSxOzzry9ppY8m6nOMnqjBTlvkTDSWdtvCbO20mxmFLUO2HV25mG9dyi9GIbe5lj
Hv4dUenmS7gjpx54L1Kj2ZwJRfddMppEvDcOHw8G1NOgHUd4/Ri3t1bOVFQniQ8E6It/GReeXjxX
rwZlggDmUYPv2SRqG0Wv5B4GySaGAU63UjCwBqTlbX0fAjjCfytV17kUBOKSIfHpnOBx6t5IeNTr
tT8IzntS3K9u/7DrDAp1mReByXReaZMt0fxk7a5wCQSk8eU44wSehnnVtuNxw8vK3wx3ueCxdI1s
SqSMSZwbkh7mB3CpfRN5ulnodPkTdk8LsqnYQ/EF23MvaPA64Dr2bElXAJXkde4qX7QksNv9RvvX
gGoK31QiUL9+7Od2+KfoUtEmpGYewE0FRMMgTsnF841hnsTMome3LCyFJmqHElZsx4kV9NJE7Jj+
iZQzwbhtucUiGqyfCyicVDUOs79FmHh61sN+pn9vwZxkr53YayrGSyphMOpwCNgndlXVl+jtqp2r
E/k/Y05ZuGU9U0xKKCY670i1s6ZoXGN0SmevCYzGqFb5wiRthGOjQedykAFI/dPkwXe94tWNaURd
ja59hgJkxr9rWgbWFcYa8oPjfiGNrB+2CJ2+51gnFmIcB+8utoqGW/x2ujsmhVhzenbzTg3KKCxy
jxnB++0xaHjzisoWscKwCVxmnBqEXhqoUQh5h+rAFLtauhJp9OilaE1jMXjJeRm8M1CMxZ4OEUm/
dVlJ49/8FoqEUSaBxXprGs+gKNQJLiRBRFCOgoAXZBRHd4mtqEXx/NIktWamE952nGdGoYBeI4ah
ikYYnAnWC0ETHP1BYuaW+/4lAuKWXt/yvxP2T9xqP1/KGMwWqu+ya2e4aaLS28vLe1KpzmdKEewa
WQHqwyI5SMPOManh6eMqKYPI/Kt+Ya5c34VCUrNqk7sEz9VIDoAw4g5cbTz/v4jaVKm7HRXxXxUK
t1i5Itg3OtximtiiM23vTuUqhcPYuY0BH2uE2e+CmQxvbB6+4lEKYLxR6GJULOYfXcfPMJj/Jsj3
gkZF5CX4/gSE/+B5nZCTCPoWCI3P2M78DfmvupfGnU880e4fUF683YHqfgrbCdn0lafs9SrzZoOO
zhrQCp17zSNyjsevm2OZLpr8X5qVZS21vAp9icO8gKRwZX7rtXoJsYzq+dThfBU+2KRB00g/7ClK
ws/BexOuYQLlFyFvXRTr4O5TF4VckW+lyY8qnSILKMGB5/7+dR6zdHz4njNEmiJ8sZoqAhEUoVSa
J+LsN+1Pt4FVChMVw7hjHw/vrtPNidrEpOYNdXyMPw4zazIHLnzXfYeN3ONqHx/bgNzaCrO+EDBh
T79qjT21P+bKr3BBadm9/GDz2fy8lZOeQ4MkP+614qVTgd8D+FL1lehEwk1S/1AukYxyJRaGt7OI
cPbNwayxyGcGwi05uFyCLmTUvoIDfO5b3QvaN8yCKDoAmU1SD7RoJCEdrbmKGyfUOY/WdDndvUpn
gNptIwW/p99F+uW8eeW0O2RZEQ2+CtLSaEZIz0UNS0WEURIL7xk0R/mlscxpp33LtzYIcQlCVdlE
FhDgT0oedjDbIDhMD3PQu5KaDeb3/i/W7r+2ausgX5xhCc9Pfh0hkzSW3kfyHRmDC31VO5j3di2G
WAuILdwCknTDEl4Zp16GQ3RNy6oeM6XsvS7HHbhrTWjROh7BH1wh60mxThHTqlVRDj+z6agB3GWT
TDCUzZiLvTMf9Iffa151m/RYKL1ZEzBtJrsDgxORAWsum4id1PMwjFhJ04jQiz0xSgpWWouloLXn
LAV/jPgliwwa2eevsL1lvf8XzP3mWvHE4ZCPxpl98dI5eGtkvYRk3vEeeqptSBTvMZY7jbNJ1xjk
mLqtww1DfYXy9bS0S3b2Wx55o8mAAqo39rwf5oQKIjAjWv8MdiJlWjA2gvP5DKkHb9qgsrMy9bYP
PwPY+qdcAawKkIctkqSmpAFeMSLEn23E+BMdaxgk+X4cxzo0itSCn5U4v1OmdPmotdq0OwxpJso4
B9vwfj7w5VwV7834UsvW3Fh/IsjCqaOX3pk51n4beRyAQOVHnr45y9TtRNbpLH4JA7QCpjiLYLiM
lqMg4Tqd6+MqzSTwn1zLedIAXdgpU5j2NKaMzK4clY4W2cKGLr1zbvrbpNk8wSOjT7KDdeP55SR7
MU0Clm7iSsjMwcZ0nPe0thwAZyMkno0hxdA93PVtw/guxaD0ADZ2iJzFtJmA8qxb8hhI4K2Bap7e
TfV1CNQodVJa44a7AaYSm81vF5UFhIq0dQL6l8DAuU7YiN5EzhvVgAen2351o+0YDRrueWLKVNY0
xZWOJ1L2SzhGpwVaL7Z+dn3EbjWieO/x8hXyEcE8D3m1lobipvW2VeZwiLIjOHggcGhY0Z9pvtDl
k4egKimbIle03vv4PwImvrKsjIktKnTPVsnzZD2aakmAL2n7O1syxDP+ymZSU4Ep1zJXyk+TiAL9
HYpZ9xSOPSPGGfz7m9D6FsIERemm948T4z+15ofhQSKwh2b8y7EgzXEfyirtJJy4p6vcgFZEOzho
+GBVz/TrskojUKCDu39HkuDm5bGX7i4+3+kG6vB17GopfnaOhrT30qQ10y5PnWA2xrP236ExJ44b
EV+oJws5fYUMadx+m85hmXTijhE/tOM4dLLgLNr6volyzqBjcWGpzUnbBFZb/vsVvQE0djMvhyn2
wbn4zPJAvHYW5ZhNgf7hF5IUtxlQAUI/95sC3Wm1t8XpqrbBQ1DD+ql5fPI2EuW4fFa8Ta3VKHyG
DudklvU0Po7QhfIlWGCef1kBaG+hzfiyG0i4F/hEX6vuWK94WzxWN9pW4/3d5qDJ6hf3MXMLrIKZ
STvsks/4sIiaHLV86kzH1DxwzanEJRK4c1DNh6UQ3mFKh3X20FTVVdsFx5bqZI8fJLBZc6nGp1py
guQmXIeQAxrFZadJXTZVtVyLA38x5XPrYBmykN5IBSdp1Jg5l1JAq96hCpG22yGz0MZl3lU/uVuC
7SyPSjxGh4xDlFgpwH2ZdWqmjfOaTbYmFzn7d+A4NDfokh2pn1hh2kfqi2QXwArLsRv0GwYKruVa
nqHId//fl+RoY0xGpBBe+ckQUMnB/RrWxSsmUfagv3hlgmMc6sI94LyMmWzNY36Lr/fWC+7sA3Hf
VpWu1u+EBsibOSTsskYkO+ef+xGRQkQatYnYYtUScmmAo3EBN6OsmSNUuxAOfG9pPTNRXBxxQeMj
E31VOL/tyQ703whIpUFbwqg71Sd+eQPBZGDRaCf9cC8atfL0vM5Eh3wtnzw3BAxoYYkOrACSw5i8
++Kj8DFVpG65NCULIumL1sAx/8ASY6eJmY468/SYhv098ZDh+cHxTERNfvNjDGoyUrsWywCyktW0
QHljqr8tzrcRCjOBjKHIabFrKxtkyxB4WUwNWsEQGbSopBbBpQnfL/AtqpwgawOqvS/S32YfsmSM
iwzpyj0dqKOSrELox7sPgToBlSv75gZQvULjHgTFkJipCw/mLcGOghZPlyv+lFpLLZeT/7GqthkB
diSpEl+yMEVsXTYR4Ffqbu3pJ4N/Pu2TErOuLCgutS6ior8awdRBai+BNV/gL8CV2bKRgURBWJVf
fDKQ0+XOYNEgnpAoGfdQK46n5nyB5poEd3gFxsZdOQ1sIJwejrniuGEMOHdH9d6InYGGlKk5fBpQ
d5/gsz1obpn1irRQVuZm6yYlJignY2mX5UO99sfKuAsJPuwq49QLZXeOwp4hA67tmqZr3r0LBMY8
cplD8tT1i1CJDb9AoiGFot8GkRxYPfX51ALUz2zPms3j7uD88jU4Up4kse/nEKuvx5nhluSPPTnk
K525VHpZP+sXJK6Ns8iH4/co869Mm08jcSsmN3VdOZfPuonhgldxuxyXOlDgrFaTSzI8xaR7gf/7
0hTHzUZEhNgjsAaKAFK7hXX2MaRlnu8o+PqqcWZlmbk+JjcsSuhHvrFJRiLqIqS9G4ExVEqjk2Mk
hqRi7UQLoY98zla9Ngdsz3OjNZ/vdUBhVS2SjNAQsgagxRKn4e7MqRYk0WMMHxbMbM4v38+tKf1F
sBfyrQ6s3W8x8kNbcD6Vo68Jh6Gmvxl5U/CTWwyhnjqaKuoF5lMqB65orVoCNsQ5Tk7/36bmALzE
DKLSQcnExCyTUMMJ4kWrpv9ZVoXZVYhy7ekJqSwVJTkDmQjqcMElfuzs9rwUA/U/4XAYze42litQ
Wtf2KZsQ+p5yB9iuiEJFnQXWMOdCZrP2z4KhSOiyN7Uh0VtcOp0WAe7HCNzxkt7ONkp5vwIX3iyZ
TEPpJjiyXTGt5fxosUkwHqguQIHCi0vdNUazDe8Nvn5x1LAz1wEaK9UowOeFWqgSrqWFCCUo7QW0
RWCWIoYBsCBjgdvJL1/aVYmZt8S7nrBm/1c7g8Y3RGwnHFrSu9O9Fxxkh2t7t7kj/Q5I64Zbr8gq
L7SD0WkI71yzDGPl6JRKw8VZqLFW9/7G+KQm+V34EW7Gw20wwN35vmHWMfBsbSrK26mNwSvaGehs
JwZ/6nI3D4TrFqLjQeIJs4wtRHOg0M0XgFJjlC7oyIi1JLSphSyXj6Yvyc6MLqtW9u3zrMQKbBzn
4hEl/aYsWbqJ6vLmeSMSAnI3zvLj/+UCtDtS5ZTjgbcqZIJpu1kkElRx+VOLmiMQHUP4eUUQ2nIY
ZbFuIiHUXtJYBzkfJJ6fH9v2QtsOJLJoRcyLiQwlg++3pXiy+h0d3gQjCqz0TRfx8appjMFsj5fl
5RLGJk3Xcpue6Gs/3K2du3IShGVvRbA2oIu50CIcVmZiGHRGUy8kjm34ylRxY9JaSK+mdOtqEtbA
UlOYJsszWPJ21VM17i5R6JaWSriCGtN+U5LaKDq9ArkQAENqZyGzyaHaD8mVdTgVv6KP0TEnWQoB
sbERgvdGp+V7GpiePkdU3HQLa1YFDpcj6pbZ+kVvA1Pg8FUdwgrA+gA5RoSk61TwgueOUhYxAzfu
jQeR73Xj85QqqUCTHkGNS6LS/jdBUCxljN1GV4o27FPlhS83TQ/L53qsjJr67200m1qw5lhA/pF1
cQg9bUO1pLZMvKonjlKKi0HfqDjZBmWLgHp9KWdtyfT7ldfuTPrQNfr58WF1tv3r6U2j95q3g1bG
nekp8YTrPJ+HnVK/R2pMfyaYDf69/zhb7JprtN3kmuwWnJ6ITs1a6nbU23bYoKEXdfFKftqJKrfd
R4cT3hR639OWrDMrpl1trC0XnMQ/Sve5qrr8g03TNHfsFvgkeibYR1pUjnjd9KLQR3uA88bEJYqk
PdkOWkZM2aOaQeUDUebh7rTRCooHcVei9GE9luQ/Qpr+OegKxqSUiUOQTjeGL5SWAaVJ0qLGXT27
dq2xemhjaxWASEal8unbUx3XlO3P/TF8DmLU/HDappBOa2VZYrg96OqaOuPfnhG9dsmC034LxrS9
yo5Cg8WkaamU89pfSUR3OPrPx7Ey5owYoDjHoxqz/DR6q7xw+PSL0tmpSfadZkAKO6kK7RCnf05j
Z7y1Q5u79wPYcbDkuVZuwDz/S2HenQuuDFfRLztucYtL9QfsafKzCNJFp2qQcno3taQiPwC5r5v3
1A9rhgxg6jdxQ/WH/IbNqnd0tIhut7q6Y8wjgMrJ2VgDosHLSzG4vnmwYgrpyHjRnRLxjDZGZCYX
zxyndwQdfiU3Qv1Fm7vwnoPwrVGzn4b3WWO6u/WjeucIHeEusoVrX5YN6WzgIVR5siWc92YNcPhc
k2qZzedNgop6rvuBnflTHR6JUUeoiMJzaZWL1MB1liYHb1L9936AYzNmtQGj5elcV/bZtB54B/0M
whkjTjd5HuEu9QMCLvyUv6jCE5cnRYzCcpMaQKzueZVW73qT641EitYEF+HPCAmuh+TQgX3lsPBn
+MkwHOL4NHeSwoVjPsUANp8WZKJah/AQms2BxZQaG+fTsx6Cil3ooQIrsXKWawG4ab4nGt44S8Rg
PUiExyn31CnbhNjVwtEKoLwtbwQToczzjLpJzEAq26wdV3dA8EkRtswo1xEhnxrXYDNeKrGYazhk
+iT46qtbUERWjRPCQ6p4j+63RTXLNtvehUqtyotZPz1tyiploCVhKyoRmuhKAv91CU6FQPYbOPyj
QY3qqrReY3RFIUVAG8TPXg7w4/3NrRV3N67fQQHR2Xj2jTWHqIcdKeVqfXxzv8mDbeaqcJE+7p/H
Ual9f0o275OBsRj0g2KhueKWC/VT8SkRwDiCCoM8mQq36poQ9mNSZxiZK1vYTHvo5fUf14katkcv
Sy/q78LYJGZx91O6WCl4ugB/eqlNLMbLMdNCpie/7r82XHLH2a1wyMPHFUWyoCStK1fAA0ihQj4a
SrLC4FkYhP+f3iEaQhcZT2cOEPJomfboDqNtsbJ5X8oFrtBafJpHmULjaIYI2g4Sb/wVa5Y/oOzt
vNEefikOotzfkVg1OCR+x4h5iXHmpmNogfdZEa+FI8VKb2ELjUDEAyvbkV+ZmwbOCbP7RvyFFMhd
8zEzpCOYACisHYZiogEr/W+w3if88o6l/4QEHRmZmVrG5Khk2VFkXf5VCznmCjcs6Is2GZlMhP4p
fw2kceGq5I0j9O6hNDb9lA8Qyllh3zgBYWKoDC44em1arEFpJDbX9iAQCj8l7xnizwKqx7FlEcZS
9yZfWPGSU2f8FeWcMVhgKKrekN9gFOHIzQV5fRT4fyQd39QgnYjKYSvKIB2zH8Bj54Qbh8ysD26n
enRQpcYpCHIG9piJzv46qYpNUWnms0SqmF11nToPpvDvAHTNK5U3+f8mDVByHnO0ppv72wjMzo2i
089PEKLVSP7FmozLe6a/2Uhc3oORGcXnfI7B/VhQHXe4vYJ73TtdIoAxk91+YXBkBWavIRaRh0WF
UOmfeE0YPT+nHxfaRhoEKVE+bp6/Ifr5ynp4pllWtqhTcGpqmCmhi0ma8Gc8kpAY84S9YBZ4DCb4
9zenNTYoQA/p6um21EfaiIxqcDrSIjScfh0Qlw3uHDatgPy7ZHAg1ksej3+A0DRtWKZ+PTQ/Q7Rn
Jgynbfs4XjEc3S44NaT4ACjI02Gf+vjaV5dOOeSr1rNwJcdqxzReauwn4NQEJQhohAXFig63ssbQ
f+vgX+tKKYSLaasgEkQrcFCTx+Ty0gfqPZMrFoFV5SmWvd8MqN3A1ubd+xugivMrOipAqybIZEqy
HjbRoT4VPtZRu7bEWFpujIcTqm+oGHz9AdjJhvSBPDBq4ivnADtXAIdO/YQnpHCmGwLUoblW7151
M1LhMl/J2TM7YT/4CGZkZlCFdKwb0x6bA+E0IrNykeBdr1QlXGc6npubX5MbD+8DYfxmcfXITTzZ
oUU0r3/r3wpvbN+Pe0ObXqsag/cJbWNVn200YWG8qDyTWS73HYi5o7gUhvKgWEHjCDa0YeXH8/N8
8vKBrGuYUZSCHz/1w9yjTywc84GfmONKH9TnNfFSmTdiQrjE6e5H+ehjcANMxcGWX5mOdY27Ntf1
eWpW2WrwBvEOaIlgOH3S/N0Ub3HSnuumiSTkVulwKruyq7X6ATwWHdepFtQ6/2nxA1ozlnCBXDLw
emW28WiThjIc3nLT2RhrVDTlcV8/N1/to2Lm7DrIRXE1IM52OblJfVVVPn4TjbRtvky8Vfe3Ts1Y
rOGf0fcxgEpwUZaIFcIzcF+FlB9TMI0UggVBDqv04UJDTxjq4XK+4jsCmHLnNBxHY0/z/09dVQLG
JSYyEFlVbKrlxRLRGDTe4m8iYDuwm8qlsGBVX6SmXw0hS/0T4KdBYsYM9ueVTBVHE4dE7XXlKESU
OaEELo6anGCfbPhKI4icMApY2id+cVZXnegN1KcuiXZgUMquT5dN58GaAoVM98pAKYKEisSLjqct
rvtj0MGIwQsPtfjsHvvJ8ZN02hKLmH+BaviM2xEX8D9YZ6TikUeZGjGuGGJ09FKgfk95Je44f43U
QDBV2VxIvaPX51K+56FViQncdR4yb5+IAyZ7hlEbFf1dvufF1FvFZwmuRYuEeuEyHv9DSGS1zlsg
TTI+/NwwPTBRJ06l2UJzBSs39HP8M/ggx9I/p6sBfOTc4o0Inersww1hcaDJQjnFpjG+3IZoosZp
W/vuEby+RAvJS1Jk34AUv5YThssQO+2Sr0GqQFL1V04QGuKg8MzVxSXNylmkX2yo3FQXoQ3f6vNS
lghHa4eRoB32ocKRbL+ZQppVurHOeddZG4jWnA6hoWndZQdW/RHa0zLwouwdtbwQVw/7wlxHX5UG
UTHLt35cwuTlToWFHOD8IzHSeccrz77/ethdEMQu52ng3PQ7JJqklUFJpEB591jOA2wniecKHQ07
uZreQynlA1uvKBSctXIA1R6bCIntPOZxMns6RA/JZAU+w3ZDpKFauIjaTyHgPNkDkkldzSkSN9Q6
IljvJFMn4N1/zwK8BIAC8lPUkTgpkRkQSaqjIFEBhyVzJ9EBAfqn4pFAMc67qRItwnx6xqBfNgUz
Ff1gXaJ+NDKtMDq6HMsdMutllXF5D7BmUDm6mXHGOBxLN0IdddXkp0M8i35mfGnOfsA0oPbko48X
41oitKp4He4aU5y0UaCO5ft7T+8lUqW0INRKuQpzGBl0hmCgDVc0N2RsNtOEhkOkZHCp9CSL+Asa
DscH5i+vjtz3KPLpL5sd+qne2jpzSc1zFfgTbJATGzmEmyHdnyQ6BCn4TRKHoVKTN+mQPFiBIFkK
/TCDVU238FHYo+3pOu8XHp8rYdCXLgyUmCtUY3mqTpdRRVEyPCJiEfX6VJI7m3qVokugwVsePe9o
pK0AXsSH8qJ1ATIiec8ZIjTo47Pi+Q+hcaasXm5rjVHavJlL2NbmFZ6qqXlGDGT2Cl04n4tQBwk/
H/McJgP1XSLsIDNhDegR6UHJJ+at1+vaBBvzuOA3ECgApGiWi+byY2aSoSWdpE2GBOCvaHu5nu5f
fMn+V0X3NlNxuyQntk+JRUw0boJlAnbJZuhHEC22nAI1UlGC93OKVEhStuT8e+7KU75vpJz4kECC
2+nQBwMmeJtaeTXOHy4ioWTO6eH+DCHIkKm0+raNZ8N1E/046B6UH7fK0MQBifp8h5f8nSrr0d31
MALBjvlH3PIWsvArufLZThaFSio9whjVoOs1pQIUZkVCrBp5TCyvhyPKRlOgLQ4RN/F47AytFOlg
zdCIuoUFzFgE1bSuc8neaXE+V7m89W5zlFbHl1fhxcKoRsITm+W9VNDul/1flnTSnowB8DwAc5O1
grAmFz7IELQvGTNzXhmZTn1ZxP11a6KphR1fDAp63udvMyArdpucmXsCwzhEBwtZ+xPJqioZjlSZ
NRSTk/IU1m7QTXIhbjdyeXKB7etVGz6G5Swh/aPQs2Olr9QgPfMb3pzOgyL7jSzxnNbPxIZtN8/O
DOHwwqo+DJBTQvRhpMJcbD+3p0tuNYGO5dvL0WVzH8AWpSk6iwwllv7cIDdBLeocsaGXtgDz8UHU
gpIvcpSEbJTY33A8i0g+LhCEw0ccrCG8oao+95NTUZJVregpnzwCEnlXCAK0PRGls+CKwkIltWKy
v2TP2rsrWCzCJmKtE7eRN/oUt5Uq4N1dvlms2kjdevLDiVQ7o1pF72fKj7xyDjkutA2ZBjId4yBi
EaDa6Dxys6ZvDjkHQ79iKQdx3/UiWBeQj8MyiTpDJl0o817bTpiACEA4LHa1mARwDomnP3TCju9r
r0eLc4Qw3duPvdvBOWkVRU64j6pPZPkPP31yXTp7Nwfdcq4iHu8v604pTBGPKsTUdozVV8kskLOQ
+wlpRuRvwop5Pp9jXjlfe7LmEcA50gfSDJQjqs1Ky8edVuNNZ3aF+6hT187xccTvHidks5ekcz/h
IqhSsg5lxbThPBDT0ju9Wd4FAwQ455i9gCnHVnLH96+5awY1M+XBx0FYBgSguR9M0bBR4Iw9z1l0
eeupwJeG/Xmp5W8CKNMthjyDNQBVW718YkYwpuzMilZ82EJbj/zm1xCf0HNctksOGSq8TGwxhcgU
ocF9ROWQUxUK3poZxMRyQvEBtIeUy4pZIyIKDYLfKcO3U/ShaOCo7JM4UmwSkUp3JVQQtTHrVJUg
7mLos9u4pYi7S1kEL8J41hMzFN0uZrhqk0FmH62PgRxtC0s/g/ES78IHyhQj2GcAEpSNMjdGGkEK
QlugyXJjbwXrhNED6mszsmYEwvcUq5M4atIteZY4sH9XsgBAX8yo8Dc7dktAdI/snUaZZHSrPmyw
WN/XiQNw84Pkuev9FRrVc4ZXumlczfPLUhSd/nbb3BTwbXjMiRLYCV3ltToXH2dzmBqQVrHF9qbH
VleJT/pdNF5UELGaSLk+mb6ayhcFciXJefw4jSA2nsIf0ps7cKwVvhfRADShYaTWuOxV2ARe4ttz
fxlgBYN0p3oCp8AclZPGjjYBljm6KO6SOgIJbantc8w+x5aGfglYyqBr+mJ9TbGwpz1/x8gnuKVu
Ql/+PsRtqid1tymEATtJ+suhjQilaa8hkWq6NEJPuTORhfQywbELS8/8OV4+9w0hC78+gZC+yNEU
4xQmPEcIzadtweMdBpixVagZXquh+dk0TY4HynV4lmtQcP1zCm7NQpH36bqY3hKaruvMWaIGY7xp
3mRXqF5YtNG4jzcD6K8m42PIBfdHYFeijUZM2RWRrLK1FkukWZPdEmm0hRuqtlaJwXpTHBHO0Mgy
FjpqMhssgc4r8E8jJY+0SGiZIyIKRAYNqu16p6o05lybTb8OeI0/sBE9ypXF+UYsGLgrz8YUghEA
nWqI79xlbJsPLCply9DH4e2sX2PgRrpPbaYNV40MeAaoElkVpRGJ4VlIi8i6iWKeAMltcObfv0hI
J1GWmg7nksLsh6P1YLQIuYKe8fsKP/CIpwAf6O/YVwgqmqF6qJPco0lCww0XQVwCWXeIUFRaPqBr
c8kR1h9+ahg1XCNDE1qy2oJpDbkoub0cXkVX6TMusr2gQnhAQo/M8h5z5XSne7NrVDqgKP8xU6eX
QGs7pk3GQJDZQI1ua6s9Qs8wfonso89gQDyh4sMkwIDE/ZZJTjV+mTvcnr32OqvxgvY7S7Aly2E2
360VtQEfoddVcAYsKM1vvd/zWcDYxiMUZ9qfGpurWHFF3F+MIwEqRtRkYDxLiqvEsatbE2hOVaX3
eEVYY2TegL0KTBz80i2XZYc/N/jGc9HUf7xDqEVKpSMfXgmFyYpP8cZkIzwr96wzfhhATmeN513X
Uzt/1l7N1bvLZzJcCnwOComEyOd//TSEgHjKpw74x9ka1x/BUHnd7nOy012K9MZt3rtNc0NH7qSM
hW03t32z+ZlKuSy0rpuWpnLlw8gx+YdKHic00aS+mYguBKIcZqWa5NmlLnWSuUgv3huKQXfUaMpW
QZvn0s/Z+FphQgubECTEqqMHawAPlWFiFYJT5tTzIoJElVckUNnC47uydf+ksrg9Axe6kharL1xC
VtpMY17WJ7FZvidP6+WBCIwsd8LOmYakZlTjKkJx2xhzt8m6wLo3kURcNxVMDiVLAZjk59wyBN5/
C/1JSQL3W/rKxkbBDCyVDAt01jliBcTSfrJqk4gjYFg44YsHtShzKJtmrK8Tx0tq2P0X3uSkV30P
gQLYqFq4fHLSs3DJexNoNdtLcwACrmIUXI/7M0GJEXLx7Dzw6IzYCrvB+gyOTFwrmpnLhM5crg4A
vH9iHFni29vy+YkiqlcOdMZEsJVv/nxkrFGE8V39HpWK9mRyv7RIYaEIxz5dJ2p7ppCso8//Lqws
nG+L6X+uKm/mu9M3qggU7DcaLuOpmSKTVO2pHMIo0ENV0REki6Q8i2UiE8DeF82lka6r04ktyiBV
6AZQXIGG4ZXGuDCfw96lfIF6vZfyEXDA6kr1NDxUVvMvYnQMa39JQdz1VeDfzg6yqjBn/PcNQSpE
oHjucm1p4EdSPOmYzcir9U2mnmSA2ol2Kjx79s922g1bOHjE55kwYMEGCJeu9BWIVsSiRYC5BJAe
kPCNN/Yd6xijPlaPibA8kBSDaskmszSgnQWVOyo6Or8WFG+HOUasakLPvBwcIzBpwc6vyGETKgj9
1+B8eBAyRH1DLdn0Efiv1lnVwaTURDeypiokb/d5WE7ioNGmNR+LG4nwA4HWy7tr7yjYC2dseC73
0MoDI2CA06T1DIHxzpaTzUww1PDXUTPA6bxVSGlMw99zNIs83j9t+eGfMekRvMqFBuk0R+90lo+l
h0LVStJSYRhK44TYM2geBDbzR+7AleTQ51ygzpmF5lMc+f04EIFNS8cks9QsPx0eADjBLivdVTUt
MAOqXq8g+B78uVXtIVT3HvKcKP+Q5H220N03rvh332L3dJu1aok0TqGl6powrtq8VeBTZYg+ycM5
a8ONbfks2wOikuZJ+CLttz4xVrHRXU4cvmMJxDFuGRcLtkkp3S/K7fAJtCcuYCcRHJaWPnRxMP7H
Z2nSQJkSHVv7lAbh59mPcflVsVD1s999zcmd00FisaDVrygvmoJ//qagGQ+ftNIiQ7KbyRDX6sh2
cwYGrQg9gep7JTLt8g9HXcpH7aFE+DmiOtDZLUPpD2Y3I5DIuemtXzvI4t1TBms1OQLUfiAhVnMe
96JWZOrlCc+xvGQNkz47MizzoErnOLtgFxPXt9FxafGnKkuxTTx6cHFDfGtMHNBY5bv7OIXZHgr3
1BJBt1oDX+WsFvuoUJO9kBej14puMkMVBc0PVgp7/us5obzsXTn1PkoI1OBkBn/wxrELnYUI6yGt
Z2CjCjti+cgvzZSv7smTTd9qDL0ju6ediAWanvK6uv3GiMPMsu2RoFkg6571cZf+baZdCLpeTkw+
64PRs6lypR6Maa73zholurOlCHEWjXjrHbHZf4wT1PbX4HmiBZKevijdUphdqs1KgUCxzk4kj3gY
zpm+Fuw4cEILfGtCdNxTowFKdBC8i/PHLxpDm6VZ9azQR4gYQ3O3cSa7ZB7NEwIHfvP2nFHs/cwh
YGdGGAAUTI/TJ8lUeWCb3lOrQR+JOFGK6NWMt/jz4eLkObYqyHVEd//WRydI9Xu6XCPoiwBSHOT4
1tZvBG3nP26EsEX7eS7U/IAv/MeI9APCxXj+5QTA56xQCiSnUubBwt3ns2pwY3hSFVzcCKjDfbs9
sYOnO0q43ok5veHM3Q0PwFVLejksUXAXCZhd0I7astZNrdoN77Z/ygm8jX1eWq+he9pyYjpmK2/E
9xsySE/Q39NeSSdGSaJWI6xG0xIuTb94J72ebjbth5ab4X9mKWgbv6aV21j2jIj+RHG5KhBpnCLt
9ZSqcRgT1MQgMvj9gWG3YsLuzU1umNJ/un6aFbvqNktGM7tA2PRyfjMiPlPQly1rOEJdDBpj2JQ3
cgkqMTjLrFBqT8efkiHvIoxS+NhHB0m3XvJ6H16cO3kIZJPYYPhhhbhOghYtjlM+neCvRYoEYCTI
cjsBxUtQtr9nc3kbISCm+rXb5IuI4RKCRBiPd5fzsIx+f1muxl41ZzwLYfHqS80EEGxwWZlacDcR
0nVFgxpx7XtUXZojGT1SfLiw32qECFJCp8CxdMWtNlu5r3g1XqY/NFyOdJlj6l2nGXxvF4Q62D1G
R3kymayJ+kGb3pYiwok59B98+2EzYWRaMleIwRmqbymXW276iJZr52ykoXrMmMehMKUT7qihLITB
UlsdlJLcdRgLZ8JoQyuqxzSv0WgGjteR6Vtivt9babdS0DEoI5GGMAzY3u3TI23QlzFTg3wzlmqh
bGTuouKyE8bwuj4+4HviLDOpGBKjwD2rFkrAV6Paa977/WkOXw4zuB48GK9pCBu7Y49QdcFK0CZz
4J3TDUe16+KCGDjByyp2O/1dg9GvzC09TB2RfgPn6BSCkTtb6RLOqMJIWw0CQWdkcrHIk7lrRh1B
xjXIYcnZdRfGlvEGPVIkvrCChp4iEvW3Ul162jthadcczQKfmIYzp28WL+q82B4O/qGWVmSBd6U2
fkmlslRVicGIRyvjhkhDXHTu8yC34OobgJzSk4z7QyWlM9BcsjhwRuafypAFK7djW96FldIRn1/T
QUrx+Tp+xbJScGfH0Uq7vbLPkPhmlMd3I/V/1/KsyHPUdSjEHfliAmIXEvWPWjo4Vw5b9yZSfZzd
9NNNnysHz1J1lwMHXnzePgR9DhPyJaqpy9xG8KzzLNzXba6Wpf4gxHIrpY1XeV1RqETQf+JU2YxD
Zc8P6E93vOaKz9R23Uk8RMQ5B9mjaTiyaIfPbYkWBn13GHaJf8ev7ch2RWi0IZfIMUS/F4rfNVlp
lwgWiH2UDx1hBqrAVoPrTj2lWYEk0eBorZ0MCpzIfftMU41dJL2YT5N0pjsU9qpzg/kpotdY9DnC
n9h8iqgbdPwun8OwcenI1UK4YtOe8OAs6+T72ngLg9QusDI0NbuFkCibWayXCvfJ1YEN3ozAY6X9
MZg4LAMJzJLCIRbhqFOnQBCMg3/6nFoBj2q7YUZvdsag0YVtPQic9AIOP4BYv7IRKRWLZVkWsCGw
YGCJxx9XNf9Hfzr+1m5KqwKRHAPslVEfpmBW66++lX6+IkGOxaQy01W22W+R47l9ktrgN5FnFD3O
14eRwr3wpA1Nu2pR2cD7hNsEhVnVHx7bOf8jYtrEeOVmEI/mEWQvTgjxe9Hk+jRxi7TX2h+ohr4a
onuGiFA8iL12/vKJt5eX8nUiYUq1zinYr+nU19qaX+NbRVCkZVK4Tvo5jgkc9q6mPGUbr8ypdHz8
qEbyyjnsgjtDmLIgi9t2Te2gUtT/GSBvRGKxbrijwfKYLx0UuMO2mzLn5ESaQPzxhtBfw//yRiXl
JuFkrqKIMtvWxTWSQeqdN60cGMb4THCnOHTByvwkaRQC6+vlDUSBbev/dDXPqbCrCsXYZ5Xo2Ioc
bJ9MTCo19U59wPqV6Zr5u0U8LB+OpQQxb5rXWIiUUwlFZfFhABIRUs0l1hVF21qErLLsEiBu2Xbt
JcaazGnyLKhM7ZmqK8eFnvJyjxNnvzpFeJuxI3q5EX7HHV5xE6P+EjxHK5kiHACDER2jQqoL0iOf
XlfRWqcz1B4vimOJYGF8ZWXqi3UkyzC8K3J15S/LPx5jQZow0s41yKLf0itatk6MQ7KfrOqitXRW
VoUxPsRgLILb3PUDLzMRdIAoQZh6dSVPG1FlLKbSOISm1YhvUD3l204B+dSD8JAA7xs3w6EyYD9Y
mQo1Oy+Htg9iVZyAjNQaotk4QjXOY5vzIHGUp10Kx3ht2CmbsfvHnCE6zlIYzcbJITaf9xrpsNAn
MP2qM8+W/OPxFKvpVqV+/hfkgsSs8Dcx/95nkElF2kxP80cz7ORH66SWMaU50E511VqVvG39pww2
xJpYElMmigmh0Qk6EtvPW9iOc9swXeuMV7Q/gtuQ6QeB28oTH3zAZdcO0xJCzf4WiFibqDfimk0k
59byaiVhdZEqstJPZgpRbicZZ/NRhl3S78YF9cd7P9GOpId0kL+8XCU1GKdqqhqc5kB/MntGI+C4
Xg1eJtLR7jNlhkj0CXeVvU+GYcSfT6fIfg1AX0GXc8H0lp1UpD4qbOp1eZ6al0G9cGVllMjmwpLh
s4oswxYeES+bbrF50xkKwEMRzThWfVIE8twzug9L2gBTdAr8D0CN6qo9I1/NmXv/S5oWA8GQQcjH
Kfdt0qBQjIIfP+A3fPj1mLhVP81bhqN1UFhqR1/2SqHRN6Hz7d2vzvxhoIAzrWrVoF734HKwhji/
wWjysPN81G1PyB8A662vYkg/MDVKaHwXNhuf6JhnmgkjMlp0BPKtUhfOYHxc9UlYi0t+tYQp9AuS
0TkRoYVg9S+4Gykes+Urp1mScivA1SFvKf1o/ERetaeod1R2U6W7tkr1D1R75vcgUQ5XOLZ7b138
RzaDGlDw/i/4NtWpU2384+v/iMdcaKb1yWwmdpY1sws5W18NHDGm+3KGNfl9vKn7TYx116WK7pMx
blX5QsVi4k9z85Oc+Zp8c4y9FwtEn+/78LUuBIi+Mn8bSOvwD97dn3CCLOPQHgrFFeFhUPPJQt9/
CiYU6QtDbH74/uPF+hToi4IzKEDp3bcg9+yStxExKcdTycCcobTqXu91MrIvzh6GfX/Xx8vmBu9C
w8eRAeDnhZGnY4CVJwn19NiD8YIIZ85KmpWcKSzUApGiD8Jb8O8ITYD1Fp+TkyAXHeXw4y1h+8wJ
iM6API1Wn0e4l9tP5AMbaeZRR97cH9eBYj9XgOoKMB+Y0JFXhVw0zlst+qX1ed0lUoyUpxa9wUoQ
tiLvNE4aCNBFZwjLTuQWXk5Eg6OzAro57HmTMNfn6huNhUimNN0C/cx5j+t1ONJhornj6eUhI1e8
ygGcIblAzv1AOKFf1UK4k0wngA2iV7YY3zkkBj1PryaJbFAv4ZyNcY34rM3ZmrxNbAMndMS7wEu/
ncpHIZe+w32bt9YKQo5yJOvmaLKrCtPLUtwRlPSr88BXzhEwR8Pftr54gOI369IUJrJW0U8gDFzn
ezccfGZ0Qdn5QhpRkzIQc+jlp3EDcOTFDowOqxoe4tXcQToQAFfBng0o9k/t6PTLNRWIOH9cIest
BVON+HjLYXHKhLbjrTqPKDcv4SbFJeYjqyoimxYD+y8g7XVzOmzn4yUrnzrtC9tVirHy/pwjX0wa
uHq5vuPqrb+56NWs1XvNWJSswHPv/rmgmtL7/h9ou6ouV65cdzLy8ZTG74/42W3yUThZVlLL2Q27
QadGB+qQYoAKmymfE6R/BolWQLjtyZWhYF3IR0ggC8kG24Kkisk7WDSpIbBe1kTJ8Przo3JyQ6ie
mi/IHGNtdLdZ+w27uKkeUvTfgcBOFC8oukNY4kVdzHvHaqchHe2mS35K1U5H+ofYkKXgoY/0z4xb
WKluRo0rDG2Af+l1iiOYyY5qh+6zGGxoj3PRzlgXvjed+6vGZmdQi7TFQDmBW506Dui88dYfNkKN
7Ld4YODaiFD4rpwIS4V11CRQoXdMMngb4blVl4uaAsbdTPqpUjcA/dyT1s/6dtZlAqTEMzXcP/D8
3LGs4thySQDBAKH+T+n0hPVR8sdJnko0lcb3B5moI4b0hVo/uHDwjqR33pqjVd24hFSK71MaV7BW
/SR1jRtoJ8thQc2SK1jpEDu9iqImVF+1BdD6ko9Y40CoBi2a+1ZHPEjB8fVQnFXM3bR8atecUvVE
S2Bc6Nv/vArgHirxVkgCTY1YuId8gtJQQCpeEqGAfBO0bc8d0LTx5vxLZjwUdfSpZEgs1NfpvA+H
YOBizBkm7tDp8BVb5nFUxn5XwnujrLaqBT0xj1U36mC5cT0VNVPFf2o7AwUENOmkaOq4yOyGSs4M
2imCJamRVSqlpa51m5J21ZpF4I8jIBFe1uizJ3BQuO6FsgJw/XUI0bAmlG1XFsnIe0QN1tEtCjyW
AWvXbiVcEgAyOFb8MV63Ni9tLKq9ben38E+mnIlxUOjsmgu5YB/8kaQF4Nk+vLWJTxnVm1CVVUye
GrF/CvzkRG3ZNy6F/GpEMEQ4bgpVCxMRXm7LlFvGgV4gBTYk2TcJ2abtVeFNvQhs4RGzHvy7sfbf
f66HQ4AwXlUQjh3yb8CrdQNfS/zmmiYsMS1d8ONrMXS5eG5Ci4V8ytyTGf5lMYw+MHKbPiF63KrD
ukVAFyDtZANdpq0xtRuVvnbWR1IyEDxPRCanqLFqqpZr9jF260qlVpzQiQiDOYiD7FDRSAClJZ6W
xd6E9IHvYSHN6lx8UOXIVJ3I9WOh3yGFwqpS5Kh6fooK8V00BsYvhRc9C3/2vBw0LnkLYJS9JjnI
YdeSFIOxzyHBGtKE5yJSSEks4rjwlGBVQQ9ZArVM6iuocNSedpuX0TVFHu9pG1oAHI+jiJqdR3xV
WuqcQMI7tMNEezKxe7VGkYnB9Ub4SELipEKkpAx2WvK7pozTCE60RjOqdoZr1kJr6AhUiYMLb1DD
qSuoitiNMvYB8XoDCxLCHPU9veugzxt6gVDjslbHVkOJClAW8BwQuXhyqa9c59Y15TikNTxWvUkI
lg3rjJ7WdfSTNco6HX0oP0U5rVU2bobN318nlr515U9L01lH/6nSb7RGWUt2wUg1VY/0bMtlNIQp
I/SR+KhQLuQBddcN/9I6YiQS2r2YfuJugkRU0QVizSjp2IrItRbsFASmrs73IACjfhoBRLwIlKJL
nV2xryOY5j17KJDDkpN3qWl48+7qLSz1tkuszD7X4UEUiEPOBamdrjwYO9QtbkmX/qe2VXoimsyw
U9eFKFBNa5QiWiJcbSVsZM0hlxWtJWT74E7zQtFjyOtxoAN5yDvW80NfKg66R/oePjJS2KhaQKO5
XWKhpeCztO/1EyxsSaGx4yEMPAQ18QF5Mg4B4JYjZ56lHEe848y+T1yCcXLLc6H42yUYj8r+Z9d5
z9kfSf1AzSAv1kDnWJFAEA+grRLQ+M9CbwuUJKb/C8QLVoWrykI19Whm+8BzNHJ9Xk4NnbL3EAZu
XIgBlcQUA+ayjmD6Iuk1rS5+EmslW3qBTpOMfbmz0qhn2Xb0csHgCedC1AkPt37Gewx5YV/8rOKW
nxmk0u1a20Lsm3k77Tnv2o1fXRV/p1J0oCbY8JVNZAoOc1laVlSL9NHUfl7PjwXyeZNxvyIlfW+p
JLOw7rd1AEMjklJ7b4wF0nEIlPc1byuMYW/oL77uT1ldyNNK1h3lmUC1EQSLhSk3qaDuWndra/wH
qTi8AmOWaog3gBDHSJlURHCi0oDZ/XW49ieRFyJZLMfmd5NEIKas+RqmzS/15XeZUp2xQtXSj/8T
8niwKduGccEC6m2fFPPQEZkY25oULrRVydqGSvHm6IeU84TwR2AjaKpCJeSGgezr6zsTQKmyhPpj
pTl/yTJhZm0n9OM4LlciyK4gH00pPS1IdCLPdfHsYDJhZEjL/jc8bY5O9ae+rqc46Np5eIn8vLwK
n/IaK2cBD4pUOwWgXEYljHS6rrT/tLdZv/sAqmab09DNQtAFCWKijavxoiwbJrWrO5uyicMpUGAe
ldSb3BLH8juYUOZqKsg6qkWOz0Evb/iGJdkBwRyPMbdfWSYTybV0Pc1yS54pPEVMzM0dJ37AhMWO
/TWR9DIEAzL2EjvyIZ+ndPzuTgJ6okjwdjOuYk8RbyDEFe2iqtAT68Q05eeg8L9Pga35/Xpj9vnF
OqNn0jI0Zg0qAQHajicILPvKHxiNjVMp/X2uPQguwZgzKA3BaP0HJo6mv3Iv7T1C6BRMhXPGjkYf
zXePW4Gx4drY02cgtZcSSusp/Ue4A66Bg+3C53yYYin0QYWaH2hrqdGH89F7cGx0lDFnWVJkmrWu
7FyaiCyL0jMJ0kmoOelQArlRizkuIYwHD1C85fm2S6h6+w1p6vKJKSqXucN8bJsOs0MvbVwnNRqq
RYl0WOjME3bG370G+W/Afe+mfYqBNcUOVVhVeWl46mfYj7zbJXlrtsITU22Da73AcK7VliVRlvqU
AO/Lg+dHI3cgfeY7hHPg3mSbyz2l/prtO3OjZDEYdzq2nNPBiXLpAl15YwpV2Ne/wDZxRucEQj0H
ibGi+nZRi1Rldqs/zulyhq6uBNqrRdymJFyZ9/ijQRjyV0PvVejOElJrk8eLaY3FaocUTWzZt6m4
Xki5jQfhau+pzyYJdDGJqJlU4ZKpVMz0WeYbbRgXogSRoCJhIlPX0QBAqzgCJO8x5TsMqp9uVWoz
JgsNVHaVISl60Z0L5ou1RZ3wmntnLn+8VK/q/VzMlXm+/RCsNbevaBbTVZvP8+WzbX6n72hYB+s4
sr5H/2PU/TUvPPUCfxlyOAD9E004jQ4KEoZypnP6905chseDOp3Dzaj1+ED3oKW44cHyRhfHiJYT
YIzT8TTaVgWELydel4DE9YQUdykBHtFgr5pMzr7IbcVy0FuAXD8A1oR0NaNEohoXSU4PB+6hi8w5
nUeBj9buqCEURLtWJsNEHv8WQ9q86O+b/JwjYme/aoyuWCQDw53cotKO3BDtSV6BNoPcCzp2PafF
Fo2LQ0pwEdh7H2ObImuipvraZzDY5R301gDwBNxeOB68erUyLd2e1+q4S9f15+bnfwGKO+VuqAsq
yBzohIW6HZXgNHNQ8wsYtwZ2n7Yxro0BF8sfg4/DLHzoszcQJ6UqynIk+THBDfb3pEPVr97VJc6z
V+G2riD98orOpUv+Fp3jsQwmQ9ubK3RXCOOkUoroIhR2rcAU7UsndJDuyBsdnpyxUzgMhWf/aFeR
ZELFz82orRuDzHQ02wJc/0+hYCQAP/i9LpPvHI/lkODTqstHAwXr9g5iHWmY2T1GtKR8oW0H9nQh
2S+J4YTnYsuGJS2WV7jMSoTEMTtQu3Oat+/+39GXjmz+s1P6C02pASGOPo96Q7NWRp67hmD+becq
E0rxuJ4+vlAjXw69J1wKbx2E3mpfqvKT++rLa4FK6/XQ0IjKmZ+pqGjh2MnqLclWMATV4M160mZm
DJAkEvQ9a38LQDyTaX+aHt9TXNXNdl4Yi5tnH4+qDT3DEfzrNryYZi126aNNUk1QqKJ+tFh0v0zj
fy50ACwjB7ts8dsT3DiSPtegxMj9de8yobEaHOm9AUXH1o/oCyWAHM2oUhXXfAHsIxFEZn0hS9La
R6PY9D8v2ZGWlLDK559pANba5M2UMU5xg8bWCunRFIfVuvnVk89SWZz+cfQrWum23WVjmKIgyNOH
f1occ8mbqJDtoTSikaxziwVuyiDkF+jLivCU6D6Famun6Ur+pIpIqIANSuHTovWGaekC/nqegACF
AM/M9genXgWd3uGJxQ7Vr7PLfhSV6HhAcAnJETcFzcyshFz7feAEdrcb0xFHV5PPy0J6KVjb2Ned
gnfORirU8ugEW8nx7/KcKDc0NxTOtOBd1hV7f9fbDQwhwubmLAtOU+ch5waRHUwJL1od5tN2Ozw/
Pq+wRNAPZTeU+qDjCiK/ceyVD+Sjomj/1AxjbWebDzvWuE4Jv4Q/Pcj+NljYt2Y+vXjT85+Iv8hr
5ZJDcw3BCu9XclGLG08QFeT6cVrZUR/+G6T3x3jiWzC7GKXJi5iLAudJmfVTf68KkaVaWBxzO+hj
VYDP0dCg+EIhV/fKt5g4UKAC9slmyVKU5TFjZvPqjr7wBLu3GH7NT48lEMucVW1oYJlPOi0l6Fhz
QuFuyCxa2kpd7HAgL/pO+J+AohLpYwggtsgz1ItLdQlylX5fL4DLPW8ejzBVIsM9OkA4+BQYeMRo
Qn4rASRAZ3qZZ+HkfSLIvzIbQbNBC0scLWlrWFhiBL73Rh8q4kUdRCvOm1CMla5Z1mog4EM3SQcG
WqkrAM0gZieluS1p6Jv9i7NQSpHUXQWaf5blklXVU+crnEi1leaIYrcbDXNP/D1FhCOmNRtHbX3Q
4JrXVmeW+a6GEdQEcbc0kPVVV748cZcVxeiXKhC2yQKcelUbISAr4+0kfEng/tjbtEg19SKPHsz5
vhI5s0dvC6pa4xB3iCvpFoS7jpI2T8pMiBGZ6+AlvLv97YDh2OwW5dM8mjk+eKzKS0WFwyUKBMUK
HsJJC3Agba/ik/WGwRnP4NCDVpbcD1iWg0WC9S8hjyJ0MYerl+S6ljD0uZCRtvn5BZ++Kan34V+I
p8GcEc4+HHnemMIIQgiusTcaIymIyfr3w9Fe/vUT72uGbdC8ry7AOzOmXDlSjS+dytsqt45xtzqJ
27oIrCaUMbcCc6oOzQ7nmqHyB6zq3iWIQI1Q1q1fqEWN22xh5nSVeYSVbe2M70ADHsTzpofUcl8P
MPqB42BZBukZ4CnyuCc25Es95ccXStopzI0obHzfTdQ+iy8axc59URBoSXn2unskgvLAOBFX3cus
082uTsjv9RwXaB3zrYWMlErndPZyOm3/nGphEtXlz8ytB7222XtqCu1Jq4WZLsY0vJkZXnymFV+k
/WrCQKZJiaTRZdwrQSC/yWsN8+Q7lJexNWJlMCBQQ9TVsQfV/1He19jbyYVuYfwtPxVJ8SIbb37P
sjUWWz3rbKb091Lens8Vy3/BCAIR/8KCNffBzEJrTKuEOLzjOzEM6jMPYOfd9KEZBIdVSi8oFfDV
T3qBE3Uyk0Al5YEJGVnZB58N3r36Qxspj2ttjIcO/xPPp3Jr89T5LkAwiWjPB4BzmIu5w27bf9yl
4iZe/GiyeACl6XKJCrbcBEXJeUnsvkJ+eLdPltftcI0wjgIqXFJSy+ktYpBzADh/79rUkLtJ64R3
2W78z4VlLlHLSxHyGKI3dJbu/a8+KjJb6nX1eKQ/0+S6Oc1fWs6O4V3++SEIbvjxGcXRP+HDoo7M
Fb/4k+U7kZZVSGAESbKHH9Xe/WdgiZKstlBvqG576+IcOYih2RsOnvqvgiaYVDTZPBNKQ0a8awQf
GxA7WDxUY441CpTUVDD1wYJtF2ByiO96njcWZEiDwe8SG4ZaK7KnqSZlHj85bduzvs/GhjMiJigd
jlSBl4rb3kbvBm1/giGGRj4kapEVC8VGaFeqPX/mmv6lAXx9KY+/L0TyOgPDz8WJg1LoVmlh6TTL
YRAskJpOVsNUHp2x0vgrlojxqUU+dWtax1NT75jp97pbhl8YQUcWtU9hvMVhnvmMLkXMJxE4mDMz
5Fk+GUqHu9OJGOQzUvZgsLhrhsyulyHS3UVKbz2FFeMjuwqVctx/OOjSMr/bkPwALxJDLEAOLzKm
JB9FePnJpxlv8lyU1WDr3L/VnZdaJmk3JRpu+RKzlm+Tj3jpPbRuk3HojQ1iUbRqguPsuZDkmdND
XsaL1ir3dXtHkf/jix/k0SK/UTUx854V8mjPD1y6aZZjzt0EKeKfDq4VniT5vUtCkwk/YYMmyBHG
gsoCSGmPF+6RM5eHUbTi128qO809EI4bipxLqJ4k1mxo3TZdvyH/H04YanMO9GkjugbHTZrkCuT1
yULQkFChCOGubzZ2SbtE8g7sZ33KpgbXP0CKCfXDDrk8me8D2MmqRohK4IjyoTeJeGGD4XrPxriq
XFEVjOgyDwuFgTyyU1og4k7oq6GgjE5+cqiL9OF5nuou1NCLmd6O5HbudNTwnJBoakIEvWlOLB0t
fAao2C5UiruS8K6lhDyLoHxC+AV/QZQNzjpWFCte0unsl0DRUXoPtq4y4UVdtrKnd/2aKKryhhgI
PdUC1g8ggDC+mnksEFWwJzNZ/LGUqL7n/3/2ZZWv+YCXENvHVg4DIaYMu69Y/GxAD4ZBo1NoyUg3
iaU2SNpCAATLCISuSF8O9xaw7Q+9h2xshDiL5tQbiZBvsIWFCDthuaMfJtDQKbopO9ihFcj2d1pj
glLiYZX/jIA3+B5i8JNHlVcD6l9/5lK5AAAY4WX5arrSv4ZbSjxF1LkV8xoDVRr7ZEJKiFEgEAMJ
FH4wEm5b8hWjZ7SRGC+oFK/hUHgWFxH56tW5AHmRaITO44TbHdNAbkPzuEkt6mD49SeWQDmja+WT
c/sVPjG78MDaQnNP6P7FVDYyMNya8cJMLtAGrBJQMB8Q1Fie7iV7VMd0ya89LP5x8qHkS0NNW1OJ
imxe7dhOke6nhjyhfAa6v9UW60fyVsR1TuH6beqtM/8xRzKFH6w37LBdbP0iCQsTulOqLS/x8azG
32gw7je2V5N00DAD9ygG1ZMjWoZPhLOaYtOQtOmEg0dnZaTWBsi040U4jBPddL5sCA3HZlMa0opH
X2y1QlWBITyBVeeXongEW9fJJHtInCAlNXjGKFyGVnp9RlSSjf+hnwbpNYqHS+YW6ipThzijSevi
+qruggIqX8je4Il2Hhg2hkx9UKmlX5CwmbjCWnOr+enclmGuCDC1g2WJ/27+RTg6VKSidXAQ+hwh
lAIf0qz+mSYvLAaGmfmQKRH4D/tSQLQTj4YjhTKnhtxQ9xvYz1zpGGN7Jmlra2Lecv5nmEsMdYK0
3kdV3DaC5U+W7HpVgoFQS1Fue7PgnDtXnep27CAsXJSLys5arH3NKgfdq3SE248tbQ3+bDCAFRx7
/JbDOBM/YFNh4M1xMMdf5dXmFL1RIT5/U5X+7naRqq5nFGGnMZigbVe0/6VkL4VYlU7Dk7B3SFMR
5BJ7oRntamUC0FEyx9YRIAqrPA/AyxDWmms/QcqmXehIGZp5OkhEp7m679SlcKMl+MPLDqXzV519
B4dhimYdZK9SpIyZ5cztCdaoJdNF3ACUQUljK82x20YX85iRLQuj9N78mSF7Nnh6iNlCPSrNEfpY
YPnNtpJe8DducMwEccR4KfTAov9EfuGDsqv+bNsmKckzcH+2q3OQaJX49nOLcbDjzaV2KsI+FQc/
8YL4BHBE5dxLCq5j1wkbmLptvr0KTbIEsFh3ETD5jDmj2nYQfc0rnd5z5sEPOM1+oneDBi+dQHb8
iLHlN4jEyUgSpNy57hhmBq10zIkjfwLxaztCo5RQmJtSjeg0vWHb2b7hOt3vNF1LOB+UXZl3l3k8
ENPWeLNhJLsDml2Ag3D7aSz+0upGx2dtqYGWnNtloHEl4I7AbNKZDHXxMGx5pOvgpEMNYThQNc0E
x3/8tJ6mnneWccFk5+/GGb0GE14NigJ+KEHg53eypFo5/QECHOLm9a9iPfA13TnrVfpVqF+g5W2s
PSPh1ZTl9apLlUnsJ2lW7s7D98XrrSy5m4Poih9UozbIj8zRPXnhs+XkJtVbwJx4nlxsDtEvVL3o
U8MNgt1weiRRaEUefn/rvcOlnV6+QWKKb+dVMtlxn20mXW/yfWzRXkMur+dGI96diach3Rg254ZV
NSpnRYuQDqg0nOqMi5UWRLAUonnnwpummTNXilc7JZCMzzW+KBVYy8elgcbQN2TGrokJPS9Ifoly
AWkcp5Ds4uaJMORGqkOjO/pOivWzhr3y22n4mPDSgFNzxCey6ypgxBywuhrjUm/nlExcxbX8BXyg
qm+NWbskcf2v4XwOWMih36DKMQp3wV0tAdbzY/ucTsxbX51igl5t4bW4NeEMlkIKWx3Ba+X7NgKt
HZp+tTsAogbVUn9fBHyGW4B3o1xgrhAGdIDS1CBpY1+Jt413LbJqnklARfE+m0XgH6+wqS1va48S
2WwQA7GtGILWy/8SYYc4qXmnymxdx6qc3+fI8ppQcy4ejFd6ApoTQNmDFjtmLaxUvkeSNsZAU0bp
XgWokMtzWBZRtbHkg5YM9Q861SF59/+oIudZ0N+VY7ViZClu7/xJ3dhAuoX95JLiJ5KopuSfwhrK
eSkX8Ty5/KCoYmspKwu5Fcrw/RoVfV/iM3sVt32006/cA4eTUQEp/nr5TPo6bOC3wN75ArSx8FuE
DDOIHrLWFfrG6Xy6Lykgz92zNUfVEJL4poA69s12PcowAfZlgHIrPjm52eD84MBdCH1Pg1ppSPEA
lLHc7MIID0OLScsPIp2KS8F7TY98+sQPEN9QVHRBEP1hBn9tEmnR8xaed9bNaRighDPvn20VMFsn
EsfNAVbqz+Lnxh5i2lWrqe1z+78Z3V98+oQ4b3UUWAgKaB5Uwlpc3dQ65eWZ91v0TMY3y0+KrFCx
sxbwomH2AUzbEO3j4qVIehcsxbb9w22u/ZXtyFzc2PSDLTALDIAjiW0M8Hp8TafCOwTSWF58s7xO
qpQfPQeJdq37cW1ntRAMrZCUdQCArSeFRiqttqpRgWZCNkn5SYtKd9On5dqqlgpEyBgEl5Ik2RI7
wI357q0h+BuH8LLfxr8fBiOanpQrcTF1zQjMGYswFYkd179SD0nDlrFTtwtbK8v0HZqC7K3HOyz9
l7xMyxpqvhxaaV6yeV9qtDJl8pl1eu91qLcJaZTn7dwE9gMNd7pFdrrAbe6aoNtzX4GvbDqOfOJ8
/VmOtmgHwCATRVi/OErHFucXBdfvh9+Y7IQwH7Ru8EASnTYrGvzdkwbFCjgRCIQDOdGdDtE61COv
qp3bD0mn+/0vlfHDePmFoXjkikmHqO3k2J3eVKmpRVfTIbxKaaElRDvzyZ30MStUDWNQZtWTK6pb
tMcab9An8yQ+XaTTTGKmcBskyFbEjdjijZtSByCh41YaAclA/KEDkdR3VC9oYLwIxuTTiJLoN7Ln
GOIz0Rp+AIHjFUFjmEA+IcZTs5O42wbwQW7RdCv49dCP4UPLPJXOox7BvLLp24BwWVIAP4sxsnHn
6gnbkwu2x1kZe5EBESo7K7AD5adF2c+xiJRVs07qNYPs5+bayOf1Ij2NuwA2H37u2y3aUMJaCUHH
fzZeqJAYRmO1RNFGW6x6HJkw9V5hLgEqKxUwQVDcOHY93D1uY+0r7cRqTGyrz7HcJM74goUx7dKA
JVB+aM3ILKWiBLSl+HXklxuXF6RddXk6Hfc9MQlxXxITMaH18w6+MV5uH0x5W2+ayF7LmYBTfRzT
ajNeZrpf+jQ/rk4egwu1S9FXb5crAoMW122LWBAjPAXVvaGFMN4hDbQcGe99yrOw/Rkk/FmK1ZZN
otpe+ME32vjb5gaxQk/hj05W0MCygwEUM+UPlJ7P5zqOCWdrrJWxj5icoPBJzcNRfDlVuJr2Jbkp
DWPG/tzwX3RcCveWQa6ESNZsKHt+wHihBeKf7YW00TDCbz2ngQdIzdIDC0mCPcg2p7Rgjli4aONM
L8gSd0MGj6EA8iOyskJpKBBVXXhJfn+el5nWkXmG+HX1ywtYS1xcW3ndmC1SU5rcM7QrsOmU9lkC
/Oh4F0sMd2tlqC2krgUZbKKn6A1+1lT2yN74EXyvSuCmorBLIB7lBuBk8haUnci0xsjLpFOhcDJM
5C/H9tOxLHJNAAMsUkITUh3gSSQpf2XVnEbYJ71tBm+hI3FVx8n2Nfb32P2iOc+HuQrUZkN0VJ1j
dWr7EEE/Ul5FnIqEBImJx2Af0tf2vsSgpar1TVKT9LmG9js8RCUxhQ2WqmBwIswZgXmo9qWCT3AD
OpdUUmeYoifx2dTGyVI4qlXqRW2S9H/frxV7t8M97noMfsTy80CzdppQqN8KBLrPFUiNXWiATW5y
KabMN03FFgFbFyLLA2bZZVjcMrq98vHSD33japNS/FD8ag+UR7SmDjlgxX8MgIX9V/NPlfJVosAi
s7j9o7iQyBe0E0SQfuPvJ1UVUYiFIjaijdPiYtKoiXfT7Ie8TDFzXdNw+dB2WmXARVd/1mr5V2eo
SJ0cBHX8VfaFjsZD8m5eAPR2PskvAVv5az3hqiNi8dAG450PDghXlzGR5+JkEr61hseI5vVSDIGs
zh7at6kM8/eBIVqUUKXftRq+Co/sWgootcb+EhnSo1plmVNusB/mewuolvX3Pmyp/GZIst5Cv+yi
Gn6ofAWgO+o6cj8Pwd1bxQQx3pzUHOy8iTKpGNH/8Pb2PDn7ixBHnqzkvAhoQ34GeNFESkfkka7M
MH05HAFxIyOYKikJbAC/wn4eAfNXuUbhberw25uY1wK34vgAtkmPzOO6fATvfPDzG3Gx+249rQ0h
nAw+rdxAr5jUCC3zKy/R0wThfVnlQTDgQmOGR6yYUD9A6AWT2VecloAOp7kVqftemH/yPoconCjy
VTnJbmnje4T9TUyMv2+ly85OA6KGftnA+ZbncQKbiYQ/V2cEVcfm2SRLEXfrT5EgkofrEKsrYRJA
zqyOKQw+jlP9I8mwnXN6dI6Dfxe1FWEBFMcflnwSQmasAkv9JjXK4Kxz6gOch9Uwk43tTj1N/B8G
fZvX7qoZT6MV3k5HXymM6MP70OPBwq33nbeXvKYrhvZMvfeAf8BuU3mT6MtEnlpGD7hxjAZbgW16
+Fmys7ewFqgziApFh6C6yoiZaFEQgCzYGHbw6jD22yQen+jN2UUA++mso9llH2Vlxru5/9PruETc
jgPnn1IiVdUhItB3C/nFodSe/C09isWtEYrIXn+CuOw2bX+J+MNsH7DwyPeIdZ3hdLF+B8lxYS8P
LzLmQxJeIoE7vN3mzktzA2DxpLmJQD7svp2kSjKoKxxoJsTu/pPxPiZQRl5WXsO5sWHoA01Dspb8
ORyVeI5AwdjIWl6nLUg3xBYy2MyiVYpx5myx3Ebt1xjN2Dan0mzdZ5VkMQXHkmubTi7ebzDPrc+/
xWY5BVO9VehtR8B8py2NPS92lbhlrfHNIIMpU3r7xi7npPmMuNVYWfBNEX4tJS3xeSNxSTMqXPjG
fwWbtu/oJ5cyIDGKYiV4ksEYlU2t5hguqlLJoOJ5hJkihigKPu5GVvjXIIF4sA4GcO1czdAasFBS
rqnX4C52dm2OW/x5MEc5SKavLlk2NnrgW6kZRCtkQX/QwX+te+LWnPH/NhI3/XlLw1a1in5dH0rp
XqDl731KuV6q2E15cz32FE9WKEGqBD1eDtXHtvBGOm1uI3moNRKr9Dsl5n1YVdYbH9j2zY0nG5NO
Gc70r5N4ABRAziWmCj34NlHmawEfAKE6X8dklLCmJKDipDI+eAuHUqkOaUtoDeIhCSx9ptwqa0SQ
hA/2OkhWr4FEOv02wxeVsIeGoHj1PWh9orOUkL/sLGuiYQoN0oMmBK6/rKLnCnE3IfeGA822PNsm
catGXUH8FjO24v655g1LBPsFqaljjaXg+cuXsEHkiRh9TzEQ+31BtrIbwe029b5xNi+iYXOU5epo
s98goKpffmJJudvX6dnbeay868LaDSy0QLXkgQLOgUfW5VU0aEtibFRW0zTeNJUBtmg6ZhJxGkqJ
lHKHlOcxwIA6SHbVWGJg/9ddd+nSNEYc86b7f7R2yKVYoUOjFrahnSZExJEgXf6DyCtKxBPeEWYL
zQ8LVoe2tjGM/Byi7sdzo2MxnW4VYpporwFXMnBkPp81MX/jU8hZ/JmH/hsZMOkrJX+kPMnunxSz
Z5iYv2sftY9lDIpgjP9pEoJeTQwv2wFf9lUKMNNWh0/8voDvtBaHYQiUf32i2A4Nl7bNrbXtMizK
FjIabPuWY48sHlVlU4wVftWerAhXI3dLIEKbuOb/oVUJHJ9aoFEKsx9ntMdLVZjPjc/XiHGEkApb
k12Yl0/394fSA1C2Dy66N6BdlkwIiH43b2meUCCc8CRsLINMLRN8Xz0ga6rRCHJZaGFGs0V+y3p3
4NGqQZHctWNyRtfvURp0yB+JpOJk6gNii3dzrf7VYMUGdlBSIhERLu73ZRC+tbroFnjaEj2VvhNF
glz/d21qrfEbNedhLSakwchibESFRyb3st1zNvJN1XqfFTgZ2B6Ked+199oGXJqfRCIVShCUh7sd
snquJp73QRPDqIo/mRLkeKy0/wvOJK1hfCKpDI/WQAPHg+jchgsivE3SJH9h5ZPC94onqK6wruy9
5XY+yOFF8E7+TRhn8ELTqHXL222U9NVQj5aa2goC7RWh7pVqlEMoAJ9vvFqt0RfK34KMVKq5w+vS
lVAtz3qpsesXW2Cdr0GK/3vIUae5tTntuRYN/knvV3LUS0Cc/5CCfvdA0x+ZtD3dJAsZCUufD6eA
cLXQ9Zri7oBLPF1nNH9c+z2l72kLQXWxdt2PBlulT/sEy9g5QYE/n4VgX4Tn9qu6S67rRR2KOh5o
gzbpxhzJGjfC6MbJxhdx6R8aPHA0rXC68xXyd0Ka+r5FsDpaAw0cgUpExEJNyKcAkp1ee40U0mje
Cf33GGFi79W0j5Ow4iycYNNuIW1TyqSs/+RX6Ovb0ZBsCZu4k06Mx5lB1jINNyc73JM1zd98GIrr
KsZjiwI6Gb4sNOo0FAjLQXseaA9cNoqEHAYD09fsghJPXSMMncenJqmQs/0csNK09WJ3eEwBUpEK
Em7SP1XYmIS83gRmTyCSewPR7V13mGswgFVQQTscNsbRSIL2mhayc9o88D2ym877pkSxfueHyrHL
mou2wpq/25eKw3Xf/0rt+lFvv+5g+3EOkx23HeOWZ/IBjzueHZTllIGbN//yp5o1T9+cz2NlnnRN
oEd0BbzhghU/YQ+W70c1FKJGl8Hem2qCCePVLtM0qs1ON299IKlaWf06UtUWROiAJ5g7WuprDe25
GRc4IqoIouaH4+e0e2yicluZtNu0yZf4aJtIbIiXvZ+Vj6aiVg2Y4jUff9Sg329ZU0JygcjhE+I7
AkWITFOL6+sv55mS4zSVQJ0YH8aiXaRwBd1ZSqKuEYr4UG6EHgvfiti0OYj98jJbB4hlRwcTCgWJ
w774NUnSeQxswCK18MahXrhqjJtDjr+3Rr6BIzso5jyx0POETiR1bk+odrIYFKVJMjdWDzgzDhpl
rAyW8wh27TNwjabrcUpYicOvk2V+Id7QPzIUcQGSrL9uSqbUJf3HynF4zePwsXSChWrXB5T+plHO
IZHNNKqWsoWhrUn5lMKyjvV9cS8D4o5hXKK7waAVfImsGZr9zVAaWI9xhuR7KQl1LldQgVvp6dhx
C6u5RlPdjie3BVZSwI/t+QTLhOPFBar3Y5zCBMuKOLXlrwNg50UzfaVYh51fe3jWILwwxS7vCaAD
rc8hFixDL/5JtchtKGGKynALTvxTxITaUokOUG++nG/4afMqxYT2vGqjFeOkF5YJaTyT3tYgPJhL
MjgGw5IqcVAM4ShtVafmto1PKUPVDYuvcGU3D+bKJTzkRs9pbaX5Cy6eYp/UC/iLXf1k9Ufj1ZIb
SGN/pgJpT8D1Cyxxzjw1mj62p0p28Y3vPhgWNjeALSpSQl+HF/McCEryYvdnGUbmoZYBNb09q3I4
w4LjkQhJynziHnT5ag+4QRSdELs/dV/ZP6ltxo7fpcVc4i6v7tJ7CCCTVwXFUEUB34lHrxYwWQ9/
zUAXZmadoETICgF90yjb2ewMvHJlm5kxiGI/p9JDFNCrvPIce2LMIAcDi/Y09IyS3QDMbcUCEMaX
13lyVFyH68OxvgvyiAj5XiuN8dGqU6ApJHyTlctfSj1mHaFNKpANzGyDtfJAomq1eGAEOS5ea/4E
WVl7+4ASNfPvswOFym+rMBWf4+46q/RENa1ySUksaUcGe3bxww1b7Ahlv+onH2isJ58LCdGDyYpm
uZMGdGTrnBEc+HZ+YnQNKEmwvznlxQzxvdkWlKMgwjs6drRM8OMjFqo0uuZLe3HO1/5xATL7zrzS
NQ90KlyXNHYqNtVPwZd4X9ClenXOKd4YLkbGXTNAxQypnMC7xOrE9y++j/Pw8uciPNtFoUxImujN
oKsNEckneVdYqu1cnJZGKYRynRzk7EVN7QTZ4jGU1Wstp0IQGHg9ajJcia2lcCyKrv39Af52aGif
`protect end_protected
