-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
EDcU4fK5Avb4cTKUQoStOlDeDKt+V9MPBEXAYihKYcOqFQS8Fs9AJQZdsajPAO+tK3cmeZQ4nSJx
muXTKl+FxYJ9qJXb53J87pMitU6D4NBb/xOTjsFgxGP2TX26sItwxOL5jiDS+yiu7LFSXlT3OcND
sN8+2DVew1BXRKrWlR4Bs9R0RpUtH2HPIhN6dZztDrRzDjnLKX4FkI7zrwMbEBs8lcRCi0m2UdhH
cwVXWpr1uiPNRK1F2bl5mcOICSvL1cT05tFKzBjCJk4AA8OBcU5XljzCf/73cx3G88GQp7uuB+d4
jE7K4KucOxr594urdMvmdOZYPgE3qUSUiyTMew==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 13440)
`protect data_block
9nArB1JnVmaBQlh54JalGRRwg+2qdRDvpjak1Z9dfveZBvmBcHGdXzKitibp5Jw1y06TIAZggEJO
od6vKEbGXAnxMcnNQeLwDm+Lsfh+heOAnt01or7SfoRbWKgjKc1TB8z1dpBumrQaXAZEiffrPkyO
qHTd4O7K9G5LqItZ8mqnqLmabQrtkBQjHwnfR47TMg7q4cEXhw7HxAixUX0IWAqsBJ7v7SW/5sxY
NprZxBmSteb11pv4cqt2zfY1l2yjIq0UxZa4WTaqX7/JVZj6o7IKNSL3cUi1uV2+279gOSmQOPxl
Lc+h8Jq6ipyNWV3Jvsn2XrdcZPAOmR1+gXbmx3mLIzVzVF7x3g6lhctkn6GfXg7VTDIpljZvbejT
uat4eYLPQyDmPwqYPnhgNUlPh8+QL756Ya++WZDjVxzsow7vcyKnJQMZ4TKYttoIqRtgnPQRfgbL
TVfQt3BkrshgUSY+YDw6q/Nzs4jig2TDmzJbtwREHHFDoR6RltjhfHPKe9PupmWL5iGE0EQkTtbZ
6xN3QDLMoSNedMi8gG9gV50O5pPiVuoKKen4IAceadHalti9GlBX2TMlo6qvEtuLoRusT5fu1SIj
dWhH3cqWwPCCgOCzth/Nr6IAFFFNiQtEUD9fy5ThvzQh+8eTEaj0/SLAMhfUhn56ehgdrNH+whH1
oPuzVShIYIWKhuwoKBcW/nXzBI47WXg7wOQ9QeEisONPDEK6mROKjnTOYjrANM4TBUHLW1x08DLd
hHRkPIutndf0RfFp8lIvIfv9rUIjapuAZCsvgtPmieUuMY2YgdV/0gyJY9z51wid3GsU7rbiiJ94
I9H3JDVV+jG/7nbDHe2YEzyWIQXi0okRziNM6tmPP7equqDYtIZknnEDB2xpkWIhUypbwmmYDq/h
hJJoJXJhjFABahMsmsaBbivQQJ9bvsjlJuA4QlxrLem6lqyF6xS/+iG5N386/FmuOG4cSJODdenA
dNwxmoIK5rDiMLT1QZ1/PCcT7N73t1Ek9/ObbF1QyyXtDqsLZcXq/paFMfrZBtw8p/HY4yxPBKeT
dO/h3qDd0lOrmATqT+/MAVEXODksv4hoMPkikOwNOwUh8YVzSJVMYVZxG/Vs5zN6j8Kb8Zf2rPv+
NKNEqP6FEgDfhIXnV2UUJQM3uoXiqDZb228090RVn6/bVA8u2nnpoGEvWUImhc3VfKwJlTgPlvj7
e0oJ/Xpx/BNQvG8yph7fQjvcqjU0LnIjKMIgXYUBdF2uB1hUB3DtznYiQm+vpkul+eMgfQp1Oc9u
cuzbXAgl8q30pBT0E0VcxDl60mY5DmyoYXpoR/r1ZHw0B1Phl8qzstu+1x1D8CbsD3XkGLkd7STd
3mpBIGVskg7Iuu6+mkzdDYLQLSGUT4TCMTdtTLrHL7vP0BFcrwvuMifH9OJBxief/Xm48hpT3bIr
a3zUvx1HFuBy1RWJoe3DqslB+kRO0iXGxZVTNC0NEg1zrAOUPG5np8tfa60tmhk3iEbRWe/zdQ4i
8E4i9DP1d9GxgCwqPhJm0/BVZByevAMiq579xOXe4pAnenz+9FvSLdLnBndS9EDUJibn/MVuC6Na
aqJh9fy62jdyLcU5ap92Ueov44Z3qddtPKmPhM5JSrBPpz6v72oJT1ILZdhVSRKkphMuvKEecIi+
6c/guejMlFqmq6vsKLWY9d3mjMyGNa56nag3iaWFxqgUPhCS/n+AoZnU35JkPCR/uv79fJGrYpF9
bApZnWL+7V1FXDxvQKA+NJRKP9fR/Wp6fr52aWyZ6ijMvlVl0s69rH632aJ5IBE7pS3xthQCHMxO
uo+xxB8y3/GFDn07I0qK44/1UUq6wzZ3Oq2+gjo39zwBg4of854wt99V8JCGLKqrfJuZV72WLDIo
jXNwgrMtvRxTnvfjOiZXXVNxi3NMg1kvk7Jq2MZxzmuO6lScYTjSBT3f8R52NoNxJmuFSRaiXSeA
R3YMkp34gM3vXMeGvaP05d4AnYUzdgB/Dm0dWkWgdU0fUOlmOXDTtqOJ3cTxH1a5I8G/ZHDBPGs4
NSyrQoMizvY6uoWGsYCuqdSJ/A8YMbOGz2dODxI2QbAznV3Z5QQK/MuTAIByF88eftHl4gvtKWTm
MQJzqfCWPYsgZT1VahEdrpVPKtql7L2hviQQVDmLv5X5EJBCPw94W2W/NTwMe36+84AkLxlpocLF
0M5YGFipM9IMj+1AfFidzXpY2oSkbTFro0g1AjUBfNlV4WzhR+ux7i7hLuGNfeEHRovUSLcIHJnM
d6B3SV0PIqy9aiqPzs4affIQJFSfShcrETcQ2KrEYsiqy6Edvljdd0xYPb95i0kBY6dsr3kEGlsz
do0pOCDn16hI5slh3pPBEeFp4np/i5qUPiMhifXDpZahoz7cPQK6MmI0O9rRD9NQQRMTfTKBVHEZ
sjVIeBxGxKM16J8a7zPSrgV0T+/zHab0h+zCjVOgzWnl0N+Lh0q4QdkxyN7ZFaIz9vlNnwnygAKp
UDU91J7E9j6qF4c+XX2E9ENTzArPb+b5WALMoBdRwbKjyho8ft7uyt5oYS++mY5K0L7X6Djy0p3D
FTSmCs3v8jptKln/r/c441TqAZZsRY0Gs14CMCPSDQtmINzyI0BAcgss7EpxkMVV+0LYK6ZxgJ87
Da3js0Lu0/vhjugJ6CHFtIEFXxK35X9PNXkQRgVDISDDRzuhG+CbDaGRDnAiaoA8P95LEwR8qNmf
J9m1ldl9dXdLqobkwWC8p0j89BP8qkUZfNFWoc7H4xCyGHxlTKfvykWv2r+hqk7kAYHnfrm/6wzl
LkfI6P5kq/XfN7CTuGoJAeGgW8Sv9nv08fROOjBkGF8PhZhNWs1QkKGrlnd8btT9dZCgswn0h7mx
n27cCZELdcY7SfrJGk6l+sNmqCah60D7wBDVKPpJitf0OZ+H+O2IiefIG0hwMRMbMejVHoBdT9Fw
2fSmsla+zbcjSDPnmQcNNYwq10ILh19HvjF59d6Mh7ZLg13Y9YCmHJxcUss2UFGmtJZtLqouv4HM
ybjGy5D4VBi3T4Pi0HC0Vmv4sgJVP8GjSqqFtnX9qFmqiJz4uNaCZwY4aqbK2BBeictfaRNXiJ62
UuJ9jRrPsuL8mJgZfdly51ab4BpZK/Vs+5FgLc0yBjsoyq+Bw0Bi3SglkoTmCqEfzdnjvRAGPu57
ZbVaSuLkObfCWIRTZFDQ8YkTEc0D+3RVyAnmaAsd5kNHd/cBhdaboIbU1+wxqlX8m8eV5XX8Te9g
fV1qcj/Wpyz3zYuIuAK/piKtbvoBcJXjwCL3KHKHuhQqBc7NLanTo7K1k5/bYtKV5UX/jGmsKYQv
pymwunvlr6jQ7RpUgDRv2ldVAMeIg+7DMabqhKLmCePqzZ3dZ3qC9NP+mZEHWkaq9YwnSefc5Lde
chuW5cj/4Y+4vg0CMQZ7qgUuM2GAfB9b+Z8Gu+RfwrhV7w9uNr0iNdwHLSiozSbqCtwWlyOWDFtn
4//wsMR4sQIOtOS5DVTCMkxYrgpeLJS8INMVhuNJdtVa0lA1vKCbsC/psZWd3oVJd4dnGjIB7ULZ
BrR+c0MveFrloLXwgtZ6T24F5T36KP6w3FZVw6xRi1qbuMIMm1/Y/6H/nERFZVZz0tZTjKccE1CN
ipnQXxW8tWzbyFkraROk4WEYueF+hK3AlGQYx9IilenijvRPvC4N0Z4QpvWVUO+VyKqC4t23xEOK
/zrd9HKTlTdVtcKkTGHmVv+kUp1Z4ITMQN0jA2ijs+glfczVjujIfDGepZghT3Q3n28lXUK3idJ9
x0heIhqLGCYmGoAhBuRgJeByv/EfHflrcUwCW7XWzORqCnhD88eCWwsyA64lCRpc4MR7oIZHXIf8
nDABYsJ+P8ShCBo2UxbpOlk28mDs/0Nm2p+BsLhLrNcqDQU+oiBdGnArjpR/GObVe8Yr2iK3CjOT
jGY816RxtY6poO/JNI5Sp4BKcYfLIMWp6LGn0liZ7XlnY39owjJq1yq7AenqmjETGspyN9R7iqLH
zRR6PqCnB97YKwtUlDmcttqfbOmq7EJKgSwxvpsnwbhw9EVJd1lm2kVqoFxWXj5ZUp5j2zu8B+e2
vKCnYMmzc74kj8SFQm9zXbekoLOPAJUcEfFmLSctP+/Cwxr3+UbCaFKC2YPYy+NP6bz+dGB8OQrI
eEyClLaQaEC6GWHEOtGUxbkz6fahOPpA22rtlyttk6eE6h4jqrbE/hz/8H3vvxROykiqRyivGVuH
PIeSsOR62SqXrAr620TtMkTqNETbLui7ZTdiAxDrx1B9wfNu8OCLk2+WfVVadrPp2d44OPW1XrHt
KG/6yqndHAtmZpJGMKt09xKWK7z535giDC1Na8B/Od+jNN+6N+mDZbrkPyhLtuL9uPf0ZHc9cV/K
ogcH+UPOVLVpxGutcpFCMiUOek1SoCQc8LjOi986BKvxExXvBsFP8+qodt5pv/ah0LNJ6UupKRlI
X8QdsSkjK8iGlRUUSvo7b6f+23I73R4roBPGTmXx/PyvZ0eeX74nEWK0vKx9yvD6AEpEkFVuEMrY
Udtw+7l+IufPcJ/A6EUPAujGufFWw9CRmb3pv9Kni4PIxcPR5X+Dt/5yniI53TcOdTBWAblbqhKF
12btr8jZ1FYL+Mads6o8R61cOyPHf3Sxtg7/qAplu/Wnba2oicMoAv5nR7qYTxVerhKEfBVdIfdM
70FnAl7VnOCv3xNyxYIG8X3IL77d2ZTjJPuI7Hg+rrXemrskbw53kMkDN5jZ71PGQEOgRZpFHNqh
tM+5NF8mr77Ea1idEECESPjdKRoobrvyFKmqBSdZDsV0ZAgUFHiob+c3YRghL3CSsTfaGLdWocIj
a39HQLZsPfT2HbUrEK/hDumTO9ef2jn+1sRna3CkcJt3W3EGTYi7hyO3lxBc7Ktft/G1WduwkQy/
tuy6Gbr6PQN6ZCa2o30W4K8XFzyDGCTteUGXVVJGhurVP7dSndUBMrstdgqMYE3IRIstGcr0jFlp
Sy9esRHwoF+GPHnuErFFZmA37fQRN75JQSao4rR9JCR4W2mBaBPBewJfp3eSUPvyRxcelzkJnzIb
7873HSPllTyAPViHwjWEEMZxTQrDqmMjiOJ323SsfYbrVhaS7xuI23CyjLt5+sDw+KJ70WFpUqgp
cZJb6O7R6VUh3pNY9cYUcKTUD2hsAcJleDM809XB9VBdTaPxWhfxv0zy2eAXycz4euHmYb5wFi02
zh01J7d+yKVfcctXtGho4G/Ai/Bd57vDua9NoplG9kSUDNxyVy3wCex46TWkU9CY9OazA7K7iR4L
rI5Jb/oKivMxF8RJbRuQsXZ1c1Hf4hPTuQ3dBY+ZO9+IsfPyAXvmJ0tftNxc+x4a0WYj3dMJwSoM
hTcOCF2P4ApFiqtnMzsTeLsp4GA115W+y0l4gIKQCBZV3BEpV5nc/kAD3jJyyTc+KmVM2rZxRg+Q
VJYgkL9pWk7vM5Lh8cCBVxH7dzQSErwuwEZ4xJHlk54eCHFhLCoj78E7ZWtL4fij72M2yLp8e3wL
jcbhb189toTVXDOHsFXa9Q3hin8+NGsYAtUXynWoaumpCBATKD0zr4nJ9d2a+9AMP9oSi0jN4vWc
hk5R7IloPXwFgeZdvhhIzmRz/sJ7rLZvV7M/wEbv+xcxGxbOHawrNtOlW7m691cVZh/1VBuCyIc9
rvFkvfp8IGeULn5ZBjURg66aHtnuXAASKgE5B+NIxEz2PRF2MJWw/eA15EdV5pVrWFIB5endUXeX
9hQa8HvEiQwkIqIQ0hiHESeg3VWLjPFW8KoRiVsEdQ1yp8tHTLiMQI3IvClmGD1yskdbx+GL7dmo
rhHB6lS6Z9p3O0ea6wO3LXDbYhoOmWXzSHvJnogVfaaaenxeInp3S/RP2KJ97m0DXCqF4oPm4zgx
qtuYJDzMkn5NIvsFg7FK38QE9gnYekisCCCRkw5ObkaXGM2KsEKh0abT9eDcw4DZqHDz+rTeZR98
+/4mhcxqf5s0s8ZHoFywDtrSiZut216ppwxBhToZLq/9aQePdyn0kQzALcr+ATyiV/pxCZpIs00V
QScGuIMOHwYHStt6YCEnqo/MSSQh86+wFHMhqr6N86K+i4H+RzMsyie7qnfMGnWCIRe5D1ch4glx
AEMfE10KMdL7XJe4df4uizdEdBsqnxhYLN0ZM0jgrvbHR31smDI3juQKYmSVwJ4XplnRDApgExez
I8IfsKgbl/4gBR7JXk+6Epv3fAqy/MswqoRxbdYJH1Z057yNFleVs6l8Nfrrj2gSKPwwniI6+Tyu
2Dtoc/pfjCbYtmGqCQ/toe1gxGW4d9q3Fm1ur/9kMzIVklhspoWWXu6uiV1dA6/Zs8Wp09A/MC+w
1+L1albA48OYw7uZ/EgBkrx+jqoWvvb9rcbqv3sOKdGIHCSxC4LXFPV41Fly+/qsvpvGolJPJx0W
0EL7cnrI1w6KePvkS8ehcADa5UWsU0ojkTzu2MyuapCrMXmt7o5X4wXu0uAOkGcDNqN7lyzqYviD
b0AGwXmJzPONeiQm92QtiJNYCTkxVqD+ipqQZcBGr4zvbAjReKH03GvwoN0tYDCdXSX/L4Bh5K3x
w2yKTJ+mdYJm0VvQnoBs1eczIc7Nk6KEMNjGqJ9b0c6PDeMvIXr0TTC8TiUJ4+fscCfkZzJy/JWv
umUQbo/nR1KvZQ1X5Bw65hy7gh9N8pOi/BQNFJTQBw/BNglV/hyUBrD0peTSRwx1hjxzsxIq5zAZ
MlSIC0sJfzftTwkGoc2DDicg25kwU4TUEGXK9oI/pKz2QSshhIlhYrVtR6TTSVA+H58f+PSUEqFO
PQLcomMXukNs4xFDgnH3Gax59B4uWH90NYPfqWrAcTuopwmg8BuTcmX+4rRfbo+dhsC+dndZlWge
DqwUcRd32VtEY1ZiGq3WHIfLQC444cNI9RfAw541hqmUdozwVoisjqR/oPyySpn6c7wDN4mhSOxH
f0yhc+zIoY3pJtgSTpSoJV8LUe9QBbVZ6AXxXkCCqMnAqdb7VqJjFiTnx0IEz0pH5wsKJZZgl55p
zJp1XtAaQ2VxUwdZ+C5gu4kPtFjQFT02RQ863mtDGVrqO3ZLI/pEGxJLwHr4QVp5Fih6mU5JUYgF
Hvx0jMcQ4h6qaBJRib9oD1qeeGf42yR1iHUBtvAHC9s7b7lb97QLc1ck3S30C8I8NAAgWIAY9HWj
mkZMzB5jTKhZlILtH0s5oq6XbjZHue3FofFW5eOlBGPKFF/OwEjdZCOAIBBSBTQTD0Lu86MPAr2Z
S9ahhW8cNFGyBuQcbtHW6Fri6EujdS6qzMqOXXW5H75EqDwZp9lvOnBLyNFYK6wsT4CKM5eAHOKx
dYs2RwKc4le8SawZMTLT0ExrJ+fql61dhjFhPUf7H6Ev8EcqGO3cf/mqT3AmN7+05GYv2NxgMvuA
TNFinbpd0iZIEgldMYkbLhOzquZjr7/ujtdlVdknJBx69dlPDqVGc27ueaov268iYf+AaH7nJbc6
2QhKcDHw+IuC2vwYXtqyGWwEkBYzs/+5SMU7ABK8myZcQglTP+Y7DW9NMcOLy1kbS51LbG+rEwep
/h+e4yy3ERSnlthpJHpbDi+1R6q8g5sL9i+Ggp+RBUD7viOEiovfjzJXnA8aak/Hj5pZg4Br+bu/
s2vDVGfjICKG3qCZm+pw/UTzgdwVuEBfYXDkCikfTfjz2ydSp61q7IRwr7SEhmWjEmQwz2oCol2c
hHijPsS3mpifA63dw5qSTBaeVA94Y8mFdifi0htkG7YAYq0PMhoV+9LZvn/v40MGxbTNOTYyxO0C
rPbZiQkUUDBqHxCpbBNRR3XJhjDVC43wH/uhn6YmfpqGaCFM5AITrNKWRkcQofpdJN8AIMwSTGMH
cfrmYXq22mqHOhfSOjf+2C3nPB//tenY0E43RmYNj9hcUrBvQvkcflzwlyO8xbB5/wq1D7jDR8Hb
h1YrG3OiZ0wDXNtV6xk3lRajxEtdOCthh3+Ht86TA/7lAj1vLxxB/AmcPd95o1w7Hzs6pv74rQ5m
38gQ9Q55KW2pWM11W98PPrE4jj1M/zx2EyiJ/w5gnq6geYPzArRJzRQV6ROiyfulNPJt4wrYR+Rv
xpL7KnRW9F1oTd8O/Uzz6hBv/7crv9RBl03zOlfA8b+9UaayXmRM8pMv6Cvv25B1DKaTANq8tooc
l/uEyaSl1fz2pMM7We5ht+T9eEqKC8YxXAvFu6xp9B8222yKzI9ztbdy2GS/Wvsz1hKaJtpVcr7H
fq2KYirOVeXDiNj712CuSK0tgvOwhkcpsbN0jcBYrP/G17+W1zss8/tWe0CSmW97EWd88ern2v7l
XCipBVltCpZhQp+LZZKERcd4apTbP2GrDhi6mxeCSbhxAihkPbYV+7rnVE3wEwgVGvXIUFYKohsY
Uw2tPGeag3JwggHTfXrdoCygZIJ/oI/cL84se4ys14XJNJ91C0DtIJbtT3SHV5wu0eyucjtXW2q/
kMvEoaEXYrtnC8IDLcJt9OBoRgYxU1Q2aBufF8PVI6OEBgtJihmo6QXGArSUNV2gBYBgaIDIbSjZ
WGGslKHAQYY22DdHQ7u0y1roJ40/JoQh7VcgnprDDLcM69NptQ+gXhsDzxJPv5KkgutyizPo7VXn
CCsG9CWmPgm+Hi4lj8L+AKvWJj0UrJoM1axXMJIbmtyE7H0H9zHhgWoLM1BP5dmnQKz8KGrmMHsP
9Afv86N92xL/cRR0xhTzLZnvnaYfU9WNYhXasfI8kdkARmrMeq7SSZhQt3fYTJ4GZ4G4cU3t128m
OcL7FahRLPLk8Ljx05QXxlSC9xpHFWtIajkET6swe63pzQVU54WiQqsiKdMjDEEqH+9wmFY7AxTx
Z8oBEBIt3bFOMIg3m3Of05Awn2KPreh4JfEtaiDJWbalM+DMprPRu1nSDQxE36vehruqVTR/NKHZ
hGPmzIQB4sVTnMiQugwkepNj6CZ6lFPDV/SR8WKNUeeO8Zst0FGV0FP5S5ZPAPgbU/K7KlCsk9DA
ZzA0uY5LkUyxMEF4gaClt3DbFW3DpxJYWTrYKKVIJRyFWoPNzpDIjFrilpWWKhqrak3uP2FVHKpA
/bmLhEhlOPU1lLR0XlzEN2gg7k7EldhkVNA2jhjwhjjhjwHoMZKSYKu5kNAfVgaxXd7zimN8Ul4I
qd+ebKZbDEbaizsKJSRbpPrQdadT+uD7QdXIJy3Vybnn4ROk/gXk0JgR5sb/+pS1OMSS8KBW3/Wp
/pZ0jONON9wtmUKbD53cTBTP6bZNpUQNIk3Kjj2oNwOQvHFNcOYvS+C3a/GbHSLxebDBxphXGpq8
CTOh9l9sNJZyglf09Vx1KMmQzyqkDLJDnEMOVMj7KNp5yA+JlgszoP7ngpJ+2R/B7XYR5mNZ9Dvf
qS7NnxxT4DMTAyc/VH/L4SmEqE3FFqAToUFpbMo1K+2sEG9tIHV/8cRE5nqWSHIHdCvxtu4KOm4w
GTwHTeeHH6M72YuZfc8gpl0JosNGBchBOlNB9MSXrlMIvV3w45UCHFriTWR/oiEhbc6yhcJT/MPK
3Zy2oXUb/9VwEqdRVDI7dJAL9w6Pugs8HuS3we/jymWQoJganlZ3ppS1MSQuaFH+7+57HqKtGoV4
ydaeBof/1wu95nr9DiTJ1LcXOfSnO5IyFBJ5Ut3YBkeOxxqeb2/e/AfFq4VoG2e8xKLQnmHJVd8w
o9QVwHwCSDCXNBpjVrJ0+37ElrCjkVcWaqHPzXSC/Ese9r4jZ9svlxtCpZfXJ4eAxXCDObh5KInd
jb3KMRfhVbxH/1A1d8k5sJF/C9PtHYN0bsmqDi7QXorjYGPLHoQdjeKA+YkdOkp7qAOwIXHPzBC5
krCRPX8E8BPcXa+0pPhdgav5R++6rn40RDyHR+ggqXgAMCLuAqlBI6eMSaz0dvD2vkzl9DJrybYH
221soaKkaYltkL05iFqD82rUAW68BSRPyvkOsVml78rlzqBEw44YXT3OBxSrk6VhcJCrGZ9fkx4T
qktyGkeZLU29IKRcWeijMpJW/6W/XXTmQi+oXyzWDXIQ0/LrGAqERhFsjNA2jMALuacTV7khsxZb
igFQz3JuHpZJ5XHLWlQfiac+bB0XYMnjsaHW/3f97Yr0VI1fCfuIppeTIzxXW94lAXLMIYfQLoW1
aTjlyA5nb6SgebUjo0I8uaPlP5esRkHUAns559pfKtr3xqICe2yOKhrA5+kh5gi9Ef+z46PHcTiu
KKi2CzBwTVgP0283vo0F1ZALBqOx7gbApsho2r2qhkK4/RDR0R3KhuD4Ug/jS4XDJwYZrUty3RQi
ryD4B7rwYWh9Xbq3a7LYJ5YP7IhHBZbyqbbNU2SqP3hAsNeTAVZ2ZJVnm2bdUPovdnWXzDt4iP1s
QaTLuUOBsXw71pzk1nZ/vrR1fmnwkCArtUs91/X/udxfnjcWCyu421w6BybTvlpY2AMUt79DjACX
EISs1zzR3eoF0ZKkSmQhWycjWTVqRQubFXSjd2060Iys4su2NhUlbFUdwlFAd1URxRwW1pY8CM/b
xajtZ/LRTXfWAo1EGo/wpba1/W9xi+3F0hY6bm6L6v5jvQ6Tk5HP53qjuvGpn1ErLwK1wRQW/wQn
PlUS7PMmVaKIKYGn5ZgW3T9xt3ioi1UYwkb0B8o37wH3FRcv75VEXTfwG9xsYYF8BX10MizN+Bhg
Nsdg9bjwB7CvGP0U/lqyveORhPVonPKk7mXr1O0f7/Q+UXA3aqM47JbprZSjTiosSGvB+H/wocQp
F5KTxui6QlARvH2YjUK4bixsIci1TCW3UokDJzo1TUnJ+c+arUWUxyuJI/dpF5YFdKqOaZTd9RBA
iX0+nMMAMT9x3sAVbYF+acCetm2WP3G+rq0rSEUkqYJIQMFNl1jDb+W0Tx5c9n/e7Pok8e05yLWL
Ky9nwZzk3fHB51Oprr2rWKKibZ8VCMz8qy8bENG5b5XlHp9kJkCiT8vAW5TzX0pT16dj41fcngWo
vh23G5AD1R1B5Oiy1fM4/mtxXeEfIBCk647ItDpU9V4hGnCYQXGM6uB+yb86hRsFeTZFq43/DB9X
+j50l2I4ekcVi8vOs6NLn6xW4qdtSqntyOMQipQO84cjbwVyEz90Miunz1nzLAbktOPQEutFXBM0
pVUmzsGE3zf7Gd6NA/BPavqjDJWcWKZ4gpLIuRQZwGk94jxHQz5n+yEsjN4iQknaTnEiH7SvCO9M
C9vzhF5LZ3uc/9sV5JMb9aLoXjvJ6XV4DORlqECftG7VOmaKH6J7G8pOcZHaFx1Dn/R68Y2AJ63l
pg+UYyPHu1Zr3+sMBDeuYhNdpHd83yO95+sXUP7F/1QcDtj5lBUASPiuJoCoG8gTDrYlMoIWESFb
caf+0njyoN7pUq0imdaCKTg8qUyBg6bmmXgmSd40W4k90vMHpZr/AqBEWljNS01/PImCYwK1xKV6
39uJcpfyz447YMhbcSEkUsb5IqOK9lze3TSFsMNdyLIP/1qPEHtIFDY+qNGZ8FWo7056/bXh+0x6
3psSZhfZ8IsCXeRiMmucugZaD6Yp6zgKsuWeln5v9uemb3K84EXFoH13tkAQ4hmC4I9Ew+0opmsq
BHPY9ggKB+MMkMD7MFwCRmzobFRfwUyxP9lgqkjwwB+DN0RxYNNGKTKfW7jDiivhsycR+LpjF0mG
FWd/+d30eH+fRR82V7fC7Qjr4Up6ROYozctHUsOFESscgzA3sM37/ZP1e0lYvSJkimaSe+OpG6Mg
7BRJw1ACBiXxArdpmBJYKgIX6X07bym4UvHJS36aoVIXfX+bEuVtgjrRSPj529H5rr4kMGObzHjt
UvxSZI/7vCvYSwl6Y5yTXVhoWXLbakhkMl5i/KQOM3fzNBA1JXyYbXr4nsJ66ze1Hzojm+yts5dr
TUNkBg5s3VF/CWztg+Bvuu2QiWC7qCHi+ckm1fb8kQC/rY10hSHz4Iv6/20l3xF9DMVl51jziL9L
s5sPWQtCO082zf1jzu41RIIpBZLiKTV+LxMB1jqP1xO8Ae6Vw+4XKJAxoL9zDR5yu7Xed2/Yo3Rr
aS+mgaGQ2+SC+ZM2mm6llynAkUJ8mui50a7Zw7XNJHfL8N+P4088t5VWMiEA/fbq69bBFt89JX0g
RmC9X8H7uFVNeo3HJ/QG3NiA/jLqQlU46PY+iHOuXGu/nlU3q1oNrRK59xpDMdyn1Byochir26u2
LbKNgET0FG2SQHNivBNKoWMpZj/IH27g2VsYV/iyiab6VDNUwifOZlLOOdT4z2jZD7skASTe2zRf
NePnfnvKxqz/6FE3k1ETrwZp0p1hRSV8Q1k/xgZjK6aU6j9TsKLLrq09qSFtyajwSYG1aACSAy+R
w0bQV4Qdug+ZAsMaiEqWs9FNPDkOQIsRFkiS8Y7nfw5SEPfM2RjrbeWxNJ48RMl/5djUUPPM2SXc
vMHL2EbSGlGj7vi70iHibVyBbVeOdjb92nBmHZ8gqu6ROqmPsYEZYxIDcrqg+1wSzuaPf4XMuYmP
lWOe+zrXbF/w1zy7KUUfmFvmwlVb5qp61hgt4Ccyt2CwgLDqmnSj3ETYH9AUaqncAZdN3qHCDS/c
D6Rmc9SliDhLspbBLQZzW++qLeHfuWxTrJQZSFdjEO//5Sq5XjfVHgE3iGGiiTVT3L5TE/Sp8jMe
kRTI8JIf7HqTZ+PLfLXlE1TiXO0AXZwEDURMvk8lWCszur+WWD1MclHGswE33hFTNCqUZFhIfjCK
Zmpi6E6SDDOELDJZvnXkRyF7Naj3FH+Ux477C7qMPSKxcKM2L2Xt4jprRqRNRXIboKmpLUguRPlR
usKivTLdpV7doOOqpcvWEWEhjqCwHhl//oG0jI2nUEKxKMKkcH9KarOworzQhK5exsN0U+E/FXjc
Mt+i3FVudI1+PTldAZvbHQcnqvmbwZekSWXlFw787fs6x4tbG4kX/YX0twhbk6p8e3EsgAWAuDtN
xfHPbRblpIfDiuwZEgsI2z/hq7KUVqtOVT+9NXLNPL/5OL3EuDUbx8aHyP71fI/XvUYhG3jTM1m6
+apaf+k1qiPK/tt+t/QqlnofucZW+Lzm16Zxph1EXATM5d4Xh64KpBEsywhAxqTSM4spJVq4GlZl
RC3H7WsS9ZsfiHllX25F2m309cKrtmde5cNONvrO6j3IVQRsQJBZaS9PTf+AIef+n8EFR1ttlTWt
y8SofJYIGwd5bQStYn2ytFNt41VVwD+EpYyuGwOz0ZlJZrA1+EnRTWTq0Dmcsf2cC0gnKnyt9gCG
QWWtXogL7vEHGVTQ78UirebcpznyReCOUzfC31lTV4HBidxe6jFZBnkKbLPRefn1/yPNiPLzRiat
gjxDQzUA/Ne/VgHvk5fWefiJG9r+pPofWYASPeNVRBxFK34I6EB/Byfxw8+dIKzPUCTyRf0ESe0f
lpBtlkt2NFuWMvgZ9wrG8DmgjoxDsMAHNc23Fe1x/HS8gF+MBZdqjDXPhXKPRKcioqXWVvgNhURe
/6J9FAX/2cRnM9BycdB+pUGcR6e9rEclTZN8AV6I+NdJAlmKH6ShbGv1qkJPCvu3LEb69Roy4yGs
PXjN6a6EPiNd0ocRFNAtYdN83b2E+YgIknXL/RRqcfkzDiHqyQ+XN6xy+FfsezGMpbgncXr0dd/b
e26p9hi1/aMQdP4x2uJCFuDo4t3pLaX9rrR0HDRm4A+BzkGTGWgqxUymysfwNBfd4lbHBgY/PuFj
AX/KNVjGqmeyWxQUUJPjiQlLRXDJ17D/a1ltRo09fS5FNWrd22afZAHmHtNBpkPTl4EKom/GxZH5
xYVeITRxvykc/kysFK1BfGBHUtJLb2ffMioQ3Nu5zd5lfyX13A3g4rQtVCyLmeGz22BHGb69O31M
B5F+CzwScw9tYrrbmlZ2bGSmHxFRYv6gtBVNasuDFJl3Ix2olrNpCYWxB108WPfbZL8QZZ4nKCHw
tgANwsJxcxUu1iGRpZ5Zy/eRgFv59xvvHfBREscuDo/EYL+nQdqeCr7XYF44yXYz9+NYM04r152e
Z6Uxz4bMRGZJ6JIx02QjsZqKSMQaygp3s5gTxea+GFLyIIstoONEcxj0oY3tJYuhhXrC/8hNODUh
Lfc/OmfU5W/KuJFsnTt1TTkcGCTihyCK0Kbqa0s3xXsm5Ins+JCsSEXVflVRxGUubPRiGHmE701q
VLdYd/URBb5ok2GZmVJaZ9C+kgRsT/U5mm40plrJPbWDjb9D8ssjp3qR9olgCc9PGbwnZTOOzcjf
jiFnZLoGNknEcwmZEBHpPMkuGTBZrJUoz1ZNiH1p/wRKP9ozYuW3c44ZIrFfXaZFRNLWVoL991hu
Aqd5+9ZwdjG5WIAy1qhVuMTK1gnXdZ6qplcikEtZBGEQzu5wlVwS8Q0h8stclFhqjrdC+eShmsh9
jx0kdSuucafcT1wCV3K7WGKOx1HIfHQlNAya8Eb9HqNPAz1cC4QyVTW/SyRErYkun29jkOyYes9O
y/LUDxSWcTYYSn5WTrE5jfUgjlquhKRCenpHgqOoAJvhpUJ0viUJJtDBH46jK9/SGL+ENHt3dc22
dQovNY5nFuIdCdA4lVt3ff4aiTe+T8TAeAhLa45wJ4pWap34oDJcEOeUumWzcEg/pfThuJj/fDBi
uaz75KNnbnzAIosLu4/x+1i4ZUzYeL9QbnqBWhvj9kxyaKCwa7ftnwbjcdC/AvWcT00kxFZSzXL+
xQi52hW58uG12vC6TcLzaETvgqHRfcvr7Y49vDFhMg2mGxeREPUTJ48Dc5VhrQt3ZuXrk+fblXTU
yB18lc0siahPj7M4M2m34Tsu5U9/6RdQogl+0GyJKwp8d3GQ/5HnCVZRe/fTeeOWtZWJkLf6OAw/
et27AblpSAC7rMHm6iu0Vzdpk0R71CTRDxSDRpK8d2vT5QwOBnH0wbqpINIYCuwpZaCIcAUILORP
sPw5subIRsdUm/gLach5E3NHkhWXCIcsrWWKSRzJWpJpE6T9lx0fBYIHmB3+gBYq5xDQdzQqTLT+
80SdS8cTHCvtxo0RQj+nXHWHE1EwJs1suEA7nAGVPmrTAZNbvYgucFvZWpQa0Pg9+qx4GuaDmPkK
riD/PFDfTcfQni/0jPFT/eqUHMwbH+95o017wrLXhPYavBPmlnWEZWHDyzLoWPqVlnWLWHKLKJIG
MB5HM+IsVis5PPeMA1RhbF7qYM2ZARjOv0Q7J17wRUcs2kiLuyvTAV1/cSme83szB22wEZYkgTw7
cO6az4L56UNij9WmD7TJ9E5Uikg1ZQkank3P72Xykq3sOmRDWeDVHgtGeTkpiBcQg9nl4W4sSbDm
YoT7VPkZmfYMeS0qzzqC+WkLxJ0Vbbu+ynie31padqZGaVBQJzk20st4Tx0vTf6yO1Vb9pIr+BNC
2boic+J81MRRCkoTJE5TcgBLa+RDQwlfapgohJItNXJGxAd4562D0z1Sp1l+n01ro2FWzPUJJx0p
wKafPLd0MGTF8aqVtMpr9rA9TGRyMEruxPAeDXMx39jls06oXPt3v0GMbDjJqfqN83XmsE+ByZ2b
NFX299jcv49Hxe/PiZAU8sUbdHxMNEikOc2iriyAFoyZcxS9ALkuT+6eY9BTXKEqDpCmzpA0JSd3
jFN0apRebuVteqceROFTF4cEuCvteyuccx+gX0sDMWS6F5YlSd4VO4abV2j9NQp4Dg/tN7koj44l
gSRqaHsmghNWB4nF2kvCkeqCK+2i5o4wSeQbUzlq9oMoMH/kAT4Xw7QYBl/n7Od0AQ7xWpdlW4Lv
9vHC2DcnHlL+2BFOnZ3+C4nebTbGAMRjb2DnScgCtfH/yyRlxZU/LW4Kfd+IRigZvh46OEyMmKTR
UTqdQ2j2MkHeq/zxaU/bfi4P+YiDGK7zf6zxUtzLdDdgAL2Hh6qmtfsbUU4k98ZgYWZi/YtXfkin
02CudY7yCzozROgLyfbk/GFw9sGX4rwT0a9xzDl91l+14bT67oTH+67R7Y6bnjHbP+aTFi2cHcPy
LH0K51N6ePMpy1JLbilM8gjlPm/seonApU3G1COcZJ1DRTrDdtmpBUcDUPFUpuTJVqi/CMoT9pQE
gtvrX/HPFD+QJjBfC1iSM5ocHTafK4b6BGYgsD6H2PyvSXRHL1I5VRt+sQNgaDl5JWAs9azF5EO8
rLbGBvWsqq4BIlAHjl0AVfDJ3aksB/BJUwLTcovrRdaTxT5VTa+4xtFhiM+5uSAunw4FxeHZcrJ/
fD8oJ60YEQ5lpUriRYdxoitbMewvvEIwbEyxcJoxWVswvPmNunuhRFd6m8lj11qrBLLp9O8oPSjp
UEVf7nVAA0IRJsK3aX8KsIMNomXANhAGD/oK555jqVcFnzF0t8vi0e7wWlz6CVXOwSIw8bw2KazS
aIWh5GeR47npd4idQ6TCCKeMdWtEA8REwGLKcSRfA00BMpFrG6ec7uaqy5FmiyHsf43fm/SF6AEB
a2lkl1NxW23KG6Uk3QvWTRy+WyghjtR3F3ajbcjHnCRiT5NTOxSzRIM/xzi00m+qebbX2ncWSScQ
ROKeOMWSZjomlG6TJ5NFwEc9JsGKt0o5wHzw4IVswIIe4P7QwmKfMI8GsJrFJoBeUgRFnfqxpfh3
w9qox5/0cLQy1ui3LkjDmXtTVygRpABGl57dWvMhNAhuiCzOza6A8C947A1kHhFsjZCgoAW/ewo0
bHbrD+PPG7nWW21rzwYEWOagPtVtfkdwbpQ8OP+LDfzpzO1/d3eqp/K8mfllzq1Pdu3KLMZjaPfm
n0Jl7anfRPyihHJrtqBAk8vpRTkS/3RwnL/sYE0hZU5NHQxaxjLIrPdTjLj3A/Ifv0frLskds5R1
FIYmugBrGKSNdVI1FBCk9s3cWlKUOJgpYNggTudD0iJGuQS+jugQpvIVsSXeYBij0SmC4gV9J8d7
09aWw1A9PhyHec8aF4Oe9800+OSjMG3i0QfBVrBnpS9IY3geLDXp82f10o/3vm4Bya/Nb6zjYSEH
EMxNhX/b+szGIneDdcVuElb3yPQJwAIHuUSPcupz/3cyGRau+0eiWbBZBWWcEGk71VwQPbsVXdDb
lOkwSlvESioXQLgefgHMyIqv2zV7YXYDP1s/BO9zqrl1mTIx9i+t4VdXJHzIphDd0jIKzLVH25HR
D4a21UVhHTQPrvqEvzDXPQQFcJFIfAANIIuUmeo36aizfFYxShgqVlDEPo8k5GEwmvPNqNdIUwB9
EAc1nWUPcX0iKRfrgMIQ/b00bZSsaBqXwVFmZgCnnbtWhuz75IjafmzTFhMfvCL9JWWTYWi0+5Mp
2pT1xAS4UQ2+AW3nOXci6xfLXptfDoL9pUYf4JeSr1g55EGyCakioNwxxFuyHWq7mGL2kTLha6tY
KhTh8qanPAvHjohRgsk+a516DTS/WBzRGQCCjTav8S57hbK8VmBhFa5VkCoFitjDPxGHTogopm/T
8qqtiDAy/YHeU86DpLdSMdDMtYHAVAVEG+TO2zgR61ZJU8jMkWBSWnQGFUg7AgLfxEx+2nC5hYb9
dz1hs88KPAenGQoVAhZZuR/4UDcwsXvO16YkWCBxTX/vybInUXau9xfz8l5me5OBdLa+9+O/Jv6r
gPRuDR7zd4QBhcCW4gaC7NIUJOVZDH5VjeziOeXRn7dclTQCs0QPyNaJseubB+30+o9HL4QUmfv2
a/yNoYDZy7QgqIdv+Gq2jcNQFVh2Y7MfoBZ+OWTf0gnHjqR6aKqr13pmck1Ez85y+wL7NxUfU3Yx
aDO7Pg5Lm9L7pqkYgQW29maa+i5+c412ASmMueGuTC9+d2b2V3jaBRyIl4xHMOogRg4DcVsdH56e
V4ujUPWG4gkeGzYmXnnVjPPTH3cPW3MlijFaQw+h1Ax5ogWZoCQrwtTwsWB+
`protect end_protected
