-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
MGG0hpVw0pwYJnvHaDUpFdxjqKGdaecQdGLeAMIYU8WCWK5n7NYBxRQCfVvTeWTs2sy8Svjnf2+s
dsKpFaYDy3FIXkyLNXVKaJaUtsKBgU0WL5etRQfqnesjjS/aYbGt+UaTlqOJqW/ZIBNo+cjkxp+U
grGCPywkyhzZjMZkJwNW1jI2S8QmC5DGzjTQByWlBaOtGuiF13prmvG1eDw8kFD/FAiL4klh7FQ6
oRxOwFux4by3oyqLsSBp1A8OdIkoe8cc33/zEQBfQveYrf4MMx1cKefcxOYQ56h5YUO8lHRFtbyq
4S6TCjzJVI4L9gPMttnWfFK23Cyr0eSLd/exQA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 14656)
`protect data_block
poNlD18T0pnSGd/chwr4MZdMJoMALiFjdpS8VqgvYYVXliJHhgHm0WyNnmLO509pd1Roa4Z+4RH7
cZJSi2T1qQ2YScgBc1pp93GJf8d9faJVvmXfwl/z4QGCtODb8loJdavwV7otWAn1QRI5/3lDwVi9
Zq6BJSNvYP9/xGIPBuBHdqNdnAp6A1FlLg5BGQt1rIkSQcPH7469P79YCbZbYF5mz6fduGg+RMRr
/WYb2+Nu1Q7BRhd3DSvd6rwbR4za4NdzK00nVMxb/6ON8R2yVX9Az32vytfGD521qo2Fyl/CQDqm
8Vc8+bpLZX9NKixzl0RjoVt9sXdmQz5lPZ2wg8+sffETFhwsnRSPZRqVw63OhxZlqq5gFLuS9iPK
T/FjQg0dwVvQO17wrqtPUsc5tPCmGJZ+4Zq9a7peT70+9pz6Nd8BE0uk1j4DM8WuRD0PGR/2xfTx
th5ZpiI8m7P/fDWNJEMrZQjVj5qW5MuIuMDG3VXA18gxv8GoWGNE9NzSMbd27u9hLpKc1vt4GnrA
DIFrpjGUAZes9CkYPndECs93aLv2pmNFIoGcPgZt/LnZB8zLrHFCSzRFVK2F2yzUvn1bdOcXoHkh
BGnQVNV5lRHwqLxkMXTD2AkvYgNGw0DtrpbhprTdSXnfntKLC1rkHSMRIXMoSUbL4wcq2wfKk8Pm
0vXk35ykaIceRcrXyOhPPYSV96Wgtc0ssW7UUXT6ob/Nj5BYLpwSguuR6XMEhRK/BmgJgkMe9iAr
it6x8rbl4N9YmakxgDqkstSC3FMMKBC7b1hE7C3K1tQUQgLS1cGtWWU6H9oAKGJSf8cwR0fc4N9y
vgQwR5nhp0sRFga15jZgABE1MKiOpl+uJHqDgSoyFeoweflCPqMC54P4JkyX23oVVy/pPlTv9TbE
0xBq2LDGp9OlCxb+uKdo8ALrTvu+G0ZlMg+1tdzjv+5gFu5y/IVSQAgz7+qH4D31kwpkDXjdD4HQ
ZeR2ZuWX3K8fXS8vekKT4DBgHeoL7qiVX/IMHKhy2C2/3Ee77gFv1rfmdbW2HgPCpq1anMV7IlRS
c+fOcW520kb0vdmuBE4AB/mXmsE6Fn/jEioNP3Y8psBWD/BcJQaIw37v7hzy4Z2ru0GCRaPfD89z
cKy26TZLRqo1p+Bwi5oXO2Q6g7IEpTBNVZg2tNGzKf6OFjeSc9RHnLL/DenV4oF1HgACaTW8jQBl
noZOMa4y2Z4UOUoIoejYBo6q9kzuTEMLKKlOgBiD8U1/VKdM8QPVe+WLI8i7NrTaX0un/Fa+0DdH
rRcWzEU5zVk64PjLCOWLazA/wCtcjm1TacyS/G1HE8pU9u29I3QDr5Py04cy81MIKKdfyHwI1J0E
TJc+hW1UGyBC/2rWIDPb95VaFzDPuzbbGPGxmRW5ZJgAnsj4/DoCqYODDxzo2ktGvv336zOYUkfM
sn+V/nCYOw4mhiNEJSDBMy3PR45CBQVN/Nj2OG44Wyde27OljrrcPrydHdmbgbDrzAC+UfomKSDL
IQmpgaDG8nHaoPA4TP/wv46LP43AWTyU86hUDOgtpwCFQjZjZpXAyPZkembTK+hpiVaqqixmNeew
UgCg6Tl5/YV44nOz5VY+xDCAF7medCoDJt85yZw2ikVOzdAzgQKXiop4G7LdTegSUXdX3ELLpmW1
igOJdmFuyjWQrtdML7DaU/DuVuuPQL5asS4pu3E854s8iuPV0oHqjJ/VY2Av7DQ3nuH+Dd57CBBl
fbXlKjE1qkxf0TN4xGSi+JAr7RNzBbshdvgX9aBcH4pIDQ2sjztDnkzeKCxP+l0hRxhRhi9Yc9sE
YpFmnbm6NFb1Y5zy9o1OrslWbKv+TR2j69ViCLWhozsQgCbHjozVhsTMhnNDO7vy02UKh7Z82jrS
9jzm0cEW/N2W+Awm5Zq4tGMNYEGhDa8qtHmFDznKF7v4A/euczKACCbwqhMy5pmvJKTnPVSCPyUE
pbysZcJatEpnwiDb2/8Gqr8nKni0KSPR8mSW6Zw96krQRhWJ6wW0nTttEC5fk0BggS37VhVoHzrP
Co4niTcRdNKWh2qfoOQUzm6A3W5Paoxwap3T3y5qnhQEkXgXiGTFme5bAiMdhW3zjRrxmoNNiNTP
zVWPZ/60m6ea6miLoV7VxRYiiybRI9ojyIBFwIqziLBviKvOdyTOj2wARTFWt5Vc6hHdQUyHqrdu
ZIuRhuaxHLIq3CfPkZnzSJHcwFbpxMW34VON6Tvv1T2NHZNv2rNQ5mlfpeY/1UM+ESqhUyyn/6p0
ZAmFhYdqbUL3695fFNxkoQPRk8RjMG32QszASDr/lTBG6IbTWPVgM1wjJt5oABxY2LDgUUAiznBP
rPlJOvCY2iUaIhTxVienneGlG405UKuHJcUNRmajwnBy7ihW0CgJby3/fVxpCz/RbY6M3sHAD07Q
GGnbLmWiyrNGyVRD6cwldn6kZJxGyeixuC08Q+V/6Cwis0arSnIQAm51z4myuLl0HHAWERxT61Xk
n/bNoK7wSNqiZy2pQTIywiIgznKWwMUWa6CH/PyX1M9UQFNxCQ/dthcS3OFpS7O1aFc13WcebFRw
5lSfa784tVFC5MKPpOwKAF2VErOLhCSGfZ+yEAfdDPqcIeGYZa3d3NscV1z05CmjUcNbzsAgXAzJ
X8pUT2KtvhMahA6QdZEpR47B7hWvF3Q6JF3VKpw4HJeR7V3A85tXZ9cTRXkjUTkPyxPcjmJNn5qV
LtXm3BYnQnTyYlfVAU2VhIzbOGMauwRFHcUSR83krTxdZ+1gn9FSJPBGThbl7yt9jzZ5iihUaA5Q
UzYlifhG81a3LpgHKbn2Qh4Etqe5kGHq010whaTdQQNHC2F2ONAoGw9EhiWfo9iE1czSeQAhoZMX
Xv+TBbc36Mgqugp03jMgQtYKTyo+dhjKOaNKdWDZ/w2m6EYQjgBxD9IuiI0Ppn5HH8sGepd8DSCR
U/ZlWSNCDwbqmQSYozBqor5AZ9CTXhlyUd5AdDa8szE7eCl4sm7x73MPUX8Z4BtlJIQ29xnK2d2n
VqT5Ie9uJPSHI/OjFbCId8n+/gJJOQh7Lm2Ai+9r2u0DjXk1nKc9W6f5zA8cpm0ponlZWe0kpm0B
YAvQKWp2SrdHEKq7Ii7hfGPUU300UaZjT/RND/CCidHPq5GWvigszrjvLm98a5ykOMTo7u10epnD
16tjpKvnjHnEnHcLJwwL+SW9YPoIMJtlFyNyYJVgY19NFVL5v//mHMXbL6jEijNgDF+dZjwHArD+
fiG0egMDQUaYjk1wzZawIXrUY9K+v3dIP8HrFa+YngrOVX6AwGnKwaEOJXd+vZEZQcKaN8GzvL4L
N5Dde6M+OAaxjA6lZ52nLQ8/hlPzIpEThE8QzjmC+QYn7dkC3dnMRebks2SIfg/QuH3ZoK+hdgBn
dpXH9WUiXjwbRUTjQeTIXVTNPWXp7i2/7OQQ+FU5UjI2TIfFcELdFoGXfWUuG7HYg9kf2Y2igEIj
W0UOhaFhcOOrI50SO7F8DshctQ0huEkltBwlqraYcypQ1xCE8PBv8qHMRzC4NvOs8JtW8//divOZ
pwG7bti4p9gTtQItID21b7cX6GvZRBpm5L8z01lObfLUchvDSYl8+JpWToKgV+UEioq/mj9+uWwX
yVpeqcPOtlY+64E9PVPbaFXNNO5kUI3CEj1VT45uCJtDUh4Haf1zrPL5ibuleWGuV8k5+Uzl5ksQ
XhrabdPk0dfy/eTkxheywTszMpKahaEH2GuAtRfVksOE8JNtxGVz/p6QE6WrKeqSHbbmYY5AyvQn
f2f0p6VqT3NOYESP8kCUPi6jfDXOhOA9rXgzDuyrYF35Qa/7hFYGfSW2Zz4YFQ+0YrLsoo8aC67E
QXe4EILA6blxnrdjvCpUFTpmR4rLsrDNK5/vBHVXLFYzrI4FJzOtHRGNhgM6ewHbLgD58uyvf6ZY
RmcwOIHCEQ1H8CkoSIJFf9uve6AQEuymTWQffj15LZmAwqtvFEnH2FSbIQ2nlrNss8v2Yst9GdEh
BboTpRX/NiFDeIgGdS4QMJ6Y7qjp6T1R8WUFr/PQRV+iEyBJ5q8AGMF25Tg9UIJHyUaLF4Ic4R+u
hutEmCdqPW/ldlWVAyZx/fs5fmTUmk2rkOpgQzpF9jyLiTixPQcd6RDdCYmOB7vPaKoPJYCJjRFu
yX9rfsetFuMd50uWDAdMqgqwQfG7vF4B2DT5XrPo4RfTDXHfM4IUHHTKJiWp9HoktgFE/sRA/gUF
yijB4lR4QuY6WlbkjpC6EizCWEuzf2Pg8A9Tt5NvAt6+BKW8ICvgFaejo3IAY+x7Qzcik4wVRWBh
OVmSs7UUoQmnrVggC2E4zQzDl/l0ST6Uku0Kc0QxiqJ8d/8qNsYZAn7HYF121tAaJ4iWxVhCShw9
NNf0Tw5LoWsy4vg+ph3lMgCaz7yN16xXs5JWlux1V9rIOmpqM4LkC+WgpjDcp3Eku315z2Tc54Df
1WAmvIBQgjkMdv5faRE87emNxrBXASovmZ554T9A+qRFIh0HHbiG/Cj0X/5IkAu3d0/ni1k2jeZ4
enQk89fZlv79WwI/XPlcRmXglqA7+eB6iDF1NtQgHCVQ4Z533e1YOHfC3DWPeQvrgwcx5DP1ibsi
9QpyC0K5ai89mgLvwzWb3v4wqrGtdK5Uv/fJP1tTNR42n5jM1ce28OMmQkGn1+Ic9ZERA8E1ris7
JGNU80UUS5mZArHQQ04YcN2NhiQu0l03/dMJdlak4qd+Vvh8FAodu1egKFhUgpVN5uZktUCz5uuv
3zCThoKFBZ0otRMGCI6XFmBKuEUmTpHv3pyS6mM4LoeB5KFGqM0VW0ecqYU6J9yv/pXTSFb4g4Bb
jNNVrBdRvV1Uja7AL+28Dld9W3HVj28ay4CbqD4fFzNp+/3wBV1qMl59mOWt0Fy371nOkQQ8Zkja
prxNLf0HFBfmUOad8NB2SXlW3CfRloqwE6FGweKMt8OMVFGQp4SP+C14tdWjmwgLTFFcv2GJ+iaI
OmgIihx5p4gdKE8UfP5HuJ+zLp3UrwP1WUXpmaE9h+CAQ5WQBzjRCmfV/uHW+iW1D48gKt6ob9pG
TytWk17lYS8epAvwk3craDkaqqWPM58ers7Nspzbt+GqJ6R0sM+L5zdEeYmyLsa0SJ5EV/HUzHy0
COsh2AKHKidxrS6Hm14OnxGlCkCDxBsuA/krFwXN6k3tBHcIgIhlPJVDFKJxLfI1PcT9C1L4QBj8
06YSN4pxbWn553Mcry3lG+qXOqRPAE9O+B0xCDlgV8df949JAxBXYmHVBsgOyk0Soawl5lE2d2Sn
wooh7wKrHrilC9/6qLv22ut4M513FtnMsXIX84Qs+A2JE0vVYpUwSG7VSJaIW+wUjMCS6EvGCeuw
AUUFkIZ128z+9jZyon5dRbVW9uF3C58iNqHD82S9ZAbtAKJT6+Ybf2JR1t+dRRsUfHzEZ0e0Pvo0
BZADJL2dZMPvl+nWACMsgiaqaFkazvnGcsu6VIkQf9dpvq+sE6r8cHtBvg0Zg1ARvlUgtdL8cWOZ
hfVUiBNmArxTOITSkEy8Acfs4DyzFqO1jghPRvJQYyg6i6Acg8gHImJ5IaO92dTFAFawgGHmg+KD
IHFQAx0zAHQXo9c7fqA6FOwgd2zIwIjwziYaKnJttojxLQkA8IJCAaOCmqQDfZqxmVMl7gDShJ5g
SUKlevPPL6OzZGTJ96KAMF7/cwgVoRL9oODEuNE4cm46dvZEZPwMjpeNmr9wIS6I49yWTxCSNJGR
EyFDtQ4gS48Hh0DYs8e2vhKty+BIWhs2XGnWUnwMnuzw84pg+6xd81+vy5+VqyhMeadmbBc7qTIO
G/lcFPuA0p2lxioV1njnq5j8xuxOQFrYEo9uGDFwan8EVxHEWrNP/LxkAQ5GO9dioqERybdg3QT5
rMrW4koD/dpnPFTtm5PiHQPGQCJT+D81QZUPbhKU26rgqk3hvAql1S1f8GZB/w3787RbgEy72IRg
PG4lrjKx+H5lnH9AVoN019ENeTwL44kYFclI+hW+udLUtK5Zvt5K6JPA6TX0bhvM2/TZHtzFO2RP
mOM1OTydVLWB3vMus22ChiJzeUCseFCrXfAxxspYLH4J9pmWf4RQWIDLiG4FdBI/VgceTHqYQ031
tEpPwUqejKCFVhvZCbjWwRh6vif7JytuSUf3KH6QMfvMGygirTvst+fHWfF1o/YRPVqt/XDVKriE
cULOJV7FcdaQtAAf7OHLtLq1W3Sk23O2NAEZQvYOFGOHkWDRlfKXNZj3nQ5D4qfcx5+u24NSJ20l
KDAxXBu1SNgerTlMC7Cpfrpg/EeR6FJyANPqsXtevE1X6YY1QEiBQzEZTSHeDajVmOcHRaewVDI9
oKurwRTZOCdmpa36GFoq/3Hlypan4fnjg15RfvTwAEh9L1LgQNxV5dA6thRJsr30zgJ/MADuZUEf
zc1qz5r19J5Hm7AHfSuWJn9BUDG/x5U5JHIIIeeaDwa0m8fyj0wd+PthjnEsel9W4b4uUo3Q6Ia7
1PTt62ITQ3cx3jA8uHUQPmK32wYso9Y+EL0TipA/9HqfTHyBmxDtq/Gsoalx3R2sKl4YZKSbmgqt
NK5Pa5gbL38SFimcGbWbMUzuTIHO1gFOcMPymIOliGbtMUf++NNt1f/7LjpTWsLVqt5BsS5hIT/e
M9bxPz33PU+ZmW2WoX2jtv/M3a9kjGz2frI9v52PEKBpuNBXNZq8SsLRNcp7rWtw5G6wc90/vQYg
11F2rA40EXoziM1IDHCgB2kSwwNGmOdB2TIZnz/pNge5AeIjMGF4GLB/V6FvZZYVR7w4va+V/RiW
RqbJ1ikdZKCfhZpJp3bmDFObNtOcOXCg9KB4TKDHP6NqACS+CXRHkyx8pC/HkgxJ9zCBpLxq5qbT
uFtTHrlVngv7m8AvF729QUhJ5+rZ8lvgj9LZcAg0z/Ui4lsPSsxC2Qz7KHZjabmKJnGynNCJzzJy
KP3TSUzYYBrGDxMv+vi61XCs6p6WNeZx6+/VVK46/20QbBJhqJEBvWK+9qkt5ZkGE/SE9yYQz/11
gGbszqVatmU81AHE+gA6aLgSKfs4nzSmCA27P93tVWZxjokzxQG71og4EgcL87xn9yCe/wrdzQ/8
a2JMF+ejRTvP2VgDjSBG2ezvsckJ0QvhTFUb7V8PNwdwo3FOP7ebW5RPuMHPL8TujOll51KMEBJt
APyxe4Oz+7BqyXiQ+CCFCgx8O9FJEW2Khg7a3msYVtvhWHk2SO1dZVuQhhJlKDs3euzh9lqAK1dy
JTvPiuKqM1R0OhZ75PNUnJUwo5UpmhRTM2bN1PugWEalP1wqpI/v+ofmRJ6MgFXYHuzYtOY0No6K
r0V0+vH/4s/gKk73VBn+g+XV6oOOmDmxatxQbAtkw7ph0LWOUR/2EaavrAKDagwfIYdg8+1DD0RT
Mt/sCeFAGMUIgBrCzGndHndo+v5K336cvJUsnuQ/dsaede1cAGZewGopjQ7G1ZWJW6NKWbHHutfF
7uuRc/LiVFwNL85e/3YMJkKrpfPHnubWAi45XZFh4nn+MI1mxTDVtSwyQDr2LGRviolTF1zLlqCU
MsJnvQ04HG9+wQQw9ykct8xChxxzy/meQsSDhrZm7ngplMEyGlGhvtxd9KIUzfFVIfZGvfoGTVOh
7vbE+dSV3pyghr2xiDX3bLIMlaz/QAqNseB+EugrDNBFdta2XazeHRVaVUeTSfbl4vRVgvsTc+e/
QjGF55a9ose6+zMh2yjKC+V/beCO4gW8Vg4CCp9LQu+ExJ4SnL5PSL+bM5UnzbP9YH2UQxIGH8Z6
4mohQfWSy5a3UH4Typw6ob+FhuZAyNJetvZeMeOI0BqTchIkQcvbU7khKfuAqK6uo+jIOdNWJdBb
9RMJGkWpoOtOJ5Y6kmp5/AeDcIsVar4JILWLW2X/G3wB6JUadMaMbsYi/L5Rsv7P2azdkFiEWIAL
5JDM2oiDK1Z/tfIEXQ4drUZ4j6gEfXrUHBS26tNcZZwnuUHPeL7LfQkTeA+8p98SLvfa1/CL0eP5
yom5UtrIqsLoS/R50fDdgCBnm2rBQp+BZBXXGgMyf3LNipAa1w5DGQoKfw61IHtFx0pCPnj1cExJ
qIziMEJ8W2RJAfRz8t/8ihJDtgsw7JGjVFs1dZ0oLEWPUIagTxKDqvLxJ7BoGGfDIKGIdXIPPkrL
6TBbbYYKHhcdis5AznyziAEvJHJFoPEHJ3h8n3PJFmWWoZhcLHK86SJ2j/FQQAfPG205o4gdHKtf
VJ9d8q/eudvvxh8/Sv+P0mQlba4A4MLuGPW46pANfgMPimqA6UTi7vTeiK2NRODn2mlLHTqBG6mV
InOEBeJFMk0XWZj3HW+s9CFz2D2fjQpWHKO2dWgYcLRdAoVlrqcMrHvCpQcnefTYfkhU0W34YLT8
7oA/lXsTWjDKpyMkbUY9zV+0B9SVxWxH/8ax9iYPurDIgq6l1kvZH9hKHCOr3wfleAH5eN9wQSz6
DuKPW6FxzuxOBoXYow7yIb0N4HvRJGFbnuQutHdtcxSH0hXbq2dawP58O9kp6cGVumFBlWh9i/s9
yOjSUmRTvtz39ouwugWJdiJ/Pi0gyiqgzQlqXcN2bYo3QtlKt/XILV5LQAajkDHmR3cder5rbTHy
Xc61Ix21rm386II3YF7cB81kU2qdsfp6tAz0LO+h0recvFPQ6NfVZhkte5eWDDeyRdDRNLgBzfZL
b6gtgAlXkSggPZeg+X6Ypzidti1ClpHWDE3Ke/k5HaTK7o2eRx9y0iSgMrU7Afk638iNzYbPFGLO
/6n/BRRU3VZyquSiV5qkTmhCZMVKL103AAXeBD+rCq+zuqExbQ9CNSMpZP76PYisuIM6ows5VYGZ
t6O4FKDl0l6n1ErB58GY9h2ckaj70TAIDveqP4ExK9jm/nfIAsfCdSdbOMchsKIFvsqn6uYxdfuy
OXYq15WFF2TFk/0mycKyooEI+P1NFqPhjx+k3/QIHbSotwFj/ZpFKJR38Vo7LV5lYtzQDIYLFeG0
JRz9g3Gc4YrJWJ6w81R+FTWj8CiO3Ill8fFrkF9nf68HoCYzfYBP6dhc/diqrFOUZXPLTp5Pe7gQ
cWxoLgFIx5iIKe8wM5EYc+3AmV1ovyRawjdmv8jHLcNSLt3kAdq1e0ntwVqM3RhuyBYLZ2zUg2b5
4RhHNRO9WR9QlsQBcgfX2MwTzzjStYbEMn3fb5eEYzlcwmZoxUWRdc117Wiv75SuIyHrwVjoJTkV
r6U9pHMBMJ4SPbIkm73TBJn73dwuHj3XmYoTPlbUBPM7TWQe6mvGZU2b+3PL4NYk1mPSz2NyAF14
J1W8eJYGMDJu9Cb0+Y1+/DfhmT5gUbM736enFoxSTa1JLc6fsjF4LBU6i9hzoi9pOhx4FZSrubzc
0DyKmA3L7/0virjY47HY+/gv2hZtUdXzmbUdcduoNheH5CekxP/j6VBqg5IS7UM7VMAkTuA1O811
FuAcAC8dF0G7cLzAJmvvmkPXk+4jXG3VbWP/1YGd6pSYryY3J6U2l134m0POIiE6I8hZL+SsIWLg
Yyd3I0FCFjFVhLfHxAezCA0Wv/+AeDTDxPlN0Z58XxG4R2IWuX7rgSl9E89Uk8G4GTjssEsyI2QX
DNtZ1QuShgavA+uK90tuCg0nFxFTviN9JyCB9wFmXO7sqJSL078inznCjnYZm1BOkb4uZ2IUnyha
W3P//XV9aBJn5ELne8blYHoB18GUX1tlDfjDD6syWK/jSlyEeof8Md5GDR2Dxdy+Leza8Fm3DYFE
rDqgTc16epBpSjvYgC0ImuErh8L2vnpcDOoHiV7kJ5lwyTW7knhHcpv09h8XvYZZzDUN2LDmcMTo
oHvP3TcbJa2AzlmliF1oX9bYylWvOeQ9Djw9tGEVi4nZkh+Df9NsaJvHP15FkjkY3a7ih1EltcYM
8Vl3hGeL5ijJ38bLfnqP9GhzMIdH7m0H4ttm1j2/vCt0DlgBidl5L5dbvrVotURhpw8/hMz6akJh
HC0TEteX0iA23tL/OhQxgcCeePHZ/BRQ+JNKZfEa49A8rstrtUHDSgMi9XLq6ucBFhQMmd6rkdID
M1hycc6zg9MOGAGowMGgnj2pwZKkWVoi4K88DM/8LCyFxLJ92cQrc0tq1ugZIZA8wdaiIiPwkYJ9
4gr14Tg1kBBu1B/LdusYyc5HDZBE14Zzr19lHZaXqNlOLYFS1pB9aELsf6j+CsR0dpHg0BoRzCsa
qogqD9+7ieRbUgMklv5D5yilgnZRe9Ci/ACnDQ3pUPbjd3CUpuvjzNMynvwZL1C9oUqhz7qS5LSy
pjtUwWIceTWsj48sY3Cw06/X0t/hpfszubj7QbZQFv9EGu5yZMHS5KOM9sX885LmITf3uQLhXTfn
Hy5jL8s7iWY4zP5xp+ADQMKdpU9xKsF6e/oUx3rah9FUWi+fyi4wnPD7kqTp/jQu7iEk30b+7Etx
sfEjMp5l8Fhtah58kv+COYASrnK55pwaPmGNOj9MaRKnY5s7JKu1dW8PrbDuwdqcRbnyTXpctbm5
5HO8KxeFWtVRRBTO5dchopX9n0RWjKBUTpw4LHpZLPXjlCOC3QPAenfZHuYcZihYhQulo9uxAD2O
lP4nqX4P4Dd/5w4YoWxlDEPyR47yWgDDFtUEi0zg/fbL+M4nxVo5dUVLN9eT+/QcG9CeaqfEDVjx
pE2vSbtuSmC2LckMr8Kathh+2B54wOAaKf6H12QzY5LMFb7ZOBCDa2LL280wWqmBb5e9JDOEOH4r
xhUsYP22KyT8oStDOpVZjjs1C/Fi9tRIwxhos/QUSUW8klkOj1EXky0je6A4yUPy6skRmUygnQPp
KmeHbVhPNbXCNq/TydNIWVkd1pgnjHfTG+GOhrvOjkexBrcUXZNxWzeMpa7U8Zr2aM3E3IvsGMch
vNaNx5qVCreomr77G+NvjblCzzksIPiJoaRQnoIdupms1SoVhgb7ROJuNMctdfeIWwDiNcGfg/kD
MYrG9cs7zJcuGhMzs3Gobo2B/i+daU6XfSFQDNoOtMfskv3QpSmyDHsSIaLeq48BBjjB4a2JlKhg
eRJbsHLLJdCRtfvWZRLiZYtekIxsM/OfDIt3AU7JrY83C1656vohoS5R/P1ighjIAnVItSHPJQ3g
/O00BY2IC8IK4y/uaIwdwI9+WvOh0q9qUZyQBfwOzI44UDaDe1LmMUxYnWnhVXzS69y6jRM3Swid
FA8TxwIndWn9sEY0qqRAttgwOvZmxLdvZwheakzQbt+jzkpSsAD3TO3hn4yO15y9F6veEwe8t5qi
QL8OTebFq1OmDh7jULUtFkzWw6d6jPS+bwUbxffe8qDI/jntNW8QVpy5IS7+5Fp2+A0V+UVF5SfE
pbSuFFmTD85pH4ejQXc5WhPCLztluFIRhywgcvFwVKIuda1n9AI6NWHcJnGMObdZE0A7D9AoTw84
icypb+xqjPWV745JEO/mqS+ubvWzcKeU67MZMYimOcQiM20eo8ev+Y5cUYNxI0N7M9Zknhy5ISCP
WHwpGPAIQjyQocbZvFj3QWJjx3gYVSxBwc0HfLkGlIChBx+qwxjd3uUVdi5ejTO09+CpzYbem9YE
sTqtzBmDmWBLRXqsIb8m/vHKufyAdpQwPVJfbautX5d43ouJWbtN12BEyBKio2i8C/NLd8d7CWkT
4FT5KU3967XDvWj7iEFx5VUUdRLbiIy5iBo7p66KMrhZFHY5NidZNdNoMCwxRmG2fKdLQWxc2Us4
AmKQc/4UfG90O+b9281N5EhyAYyrdkguqJpEBi1Z3zCX5K1YsGgahh0CPoKgNUP/+emoMm6Jh5RB
g/UGz0trtX38DdFYqv62/JjhdlX2KUo6nPUbx2ifWb0+iScKNNdUpw6YmrbF+WMFaZM4GcHw+/9p
XM5ne5leQm5G+RONbbMM20qZiIuUs7RZTLTQCXaij8nmgMVoSKsLUl+y00uBuezH/5Py+gs45lJB
NqexvlO8FhT10G4sCTIKjQAKkba39AOHKYj0xTj5Scv/Fi6WCy2Q3P4NaDlgMhiXHHJT1rNuY9FF
TwuS1+leE5rRZs4nPCdRpnRIvgTlWUDzT3iTdmZ8cE3pu3TjAt1G1G2cNwCNuMEPYJ155P6ZteFr
dOMLfe6uXbeeFlTlxK3rvMQGfcF2W7vqCdrYAvS807NMy1ox9hX9u62E5YY31NTmkU7z7xUU02OT
DkMecA0tV0equ6DtqTah/VnihSr4thj7+sI1QQ2c12RA7VdwXOkGqWWOsOq1kgLOEF6zf7TRj2Q0
oAfM4WBguNQOZz1EoKPM4PHYx+PHztZoUJ6R0sS715DXc0sIvCSFMJT37VCg9n4u+JzkRZVTR3ob
zsvdpEaNiV58QRRoNP+xhzsVnOxij4wAkZ8cYrXi3erNQnOl4y61JGNGFsDB24ExGQELziM8Hss4
+bVr8peAtZq4vmZiMw439oyIKz6EsIfowFrQ5jdbeLmJ6C5bpTWNmnMt+QRsT6oeHLdhbIN9w10V
oekGMeSY1otoEpfSstjrQWtcZuKbuMhf3PfKMbYxfP4EY81Di6uF5/NrIKNWdIjsj7fn4p8BEsLx
aB6bhUT8eMopqXns9rtiYm0tUFjLrPD/lKaJcHH1QUNH2iBlg8X4p4NCmommAFOv1Ly/sKXESmcF
Pop7CPAfdWV5vrZGdirrkSc4io9UfdNQFAWyDzWcTshnrE5DeBTGvlKVIVXnH7meNi0fn+FKc8Sc
Yd48TV2fLC4my/bWu7BdoUaV3SPMhLd1Rq6NQRcuZPDiNn6reJ+r8EBUotqLk0/lqUpNSQZdsmqa
oyalCqncKOfslDGM9s41C/iN5GIFehCKrbK2Kl2AJmuUHnEGjk7Rma80MvVFsYkHkl7anp2gLLO2
tZZ1KSjA/S55BBFyZZhFT2uYudT38yTuftbrgeoXKCdVWourJ9QUm6aBq1FiVz7ulJj8bkmTXPN6
i4l1EGsMegNBBe0a1HrJiURbwAktdSx7RRKnHj7gt5o5aqk6pylyde/3GVVWXQIir6SJrxr7YjV7
Fu8QzZ4rIlmMF1taWb4S4MDo0IXRwlcY5rtVo5ll848kfcbY5tSN5PD5HLwuyo2kVKiVpY/FZMy0
2d9L2rO7G0W0wZbDFIruCnhMpJ9R8OXjFKo+LFuJRuwiSb5J5YlqoPRSjU0maA4dfU2UHVTrFAAK
9v/7Lz8fWGxgwRFPOFX6Apn2Pj4xAAg6h+MFRAs3N8DaF+iGKKEdICEcQO8xktBruDyodZP/qOWo
pHtNlV9Ox4mZZr4pGB01wowJWBU6e7HDe62McLKjMx5CiNG51tcjSrmB7vayVjerb4SBAMk/URE7
A9Q35uu3Y+qO2N165oJUSW4jQqcn+JxqNRDWlqsw4p3FN5LrDsUWqmRojJKjZCYATenWmfErTM7j
484SweoveYatX/0M50Zcf77u1JlEgZR0fULUbShf5w+LmNFEcztzSE8JjkRuJE7GTcq/ZVzFNvLS
4XDJKtBCHhVxrRfcAQHN2c6Nbyl9Sjsi25BnVbnWz+Yg+2Ov3nQfb1yNpbD2UMKOBdZ9zJJ51wA9
p63tZeHcoM6kSzj2zcofQCgcUgzWymfrJJtfJCBT6a9O1ZWQbic+3yt9lT+hNmDobYGGoRnigXOO
vOhRNRUI9TvPl/s4FbunOYhUHFkFfjuGRnIVe8w0fOgGx3msgxSLaN2UX425FBoafcUL5LFnYVGm
MSBmViJAQo9SeuW9/GuU72Kz21I9McUokzty5CNhzUatm1AZXI/v2736CifEndsr2jpmgL/TrbOi
nJMmS829vZ8sS9q4SioucnPgX5bw71RMTBCBICZsv6JRFY6WpX6VNuJbuQevRlJKB64/CPWuPzck
/K5KB7+dKSuUpcEZHlHVl4AYycdgFeiOC4MaSmVKcKExxteN9vn8YzGiU6RF3rPVrP5PCC23D/8m
MUhLl34pI5BG2vishhelgRSg4UXKFkMSNjOz9bVZRFjSsnvtBjlInexK5Zdr3zkuoGp9dfOkKV86
K+oDiav2y+67jyddiQkhhcSex7g7bHnfVDm3CQnZes7LPO9VPj4AX9cLtLKoxn1LE5tZwePorKFV
yKUpgK6IXEVA5idCsgqTkLDEYakqQrb8Tez1EsJPFwtuvZlSIi+hQ14DLdp3NYDwUQOqzxKR9FIw
kCgzvhjIHnKHIrak95PqlVHH9Dl9NbNTYCH2xLhiQWayOgfkS5Hr6OrC2JNHBEQDF3L39ec5167m
qXnSeAwFKKEt5+p7rTqHvr4hhpadvtjqdeVFj/+PLT/DMPFWsY6hlUKljDM2UV6rz0QJUy/RwE/R
kqBFZjntQ+5PfujZx/Om368yJRcSJ0fO40xcFPJud8/dyN16+xcMBXd9QDhI8VvSz4vgNWvJdVmO
gGi19muF4A8uVzQc1Pxqb5Hx3TOH9mRaEq3E45B66T3uv/tYcmhPU60d9J+EyYMhFbmAJJLXlMXr
84jsY1WRV1MpGg88ROUAl3q8Vn/gKoVjbsMprhVw1b50jk4+md/DOn+6IvmTW7sE4X2W9m6B9mk1
GFYiTUehJUwL3ChMgeDOgIzG361BrLgyQPI2I6o8RFkzijqA0Y0X5WWGcm9Ds//bGA1Ab3nlaUai
3pt59bVNoSSv6UPqfbnuzdWw6bv3SyYtXypL6TMi0o3TCXbi5dWysnZppBvIeenRvWGAcxdMljtv
HVcbbzEGWxg6UDoY0JCjK16sfXt87H3e6YC5bpzP9vL0/y7nmpjx2gDHXTkv2Agvb/6jG2kfSKvb
ihnU/W4zaG5Y1jiIfhm4KWksTrfS6QchxUOkdu59Hed+U2+c7sy1e7d0TeLa7yE1Y4vWRn+9m02o
rdHrv57yOwb6cas4vmKaATv3nTAkA1tCNhPvhHSaomOsRe5NexNp4oaPe0jL9Ly4ceApGxNBFNDw
gjh9wOGRF8+xXd8q6Sc1PKRlOA4clo5Muz/MQl6WE3HT2bN5wf1bcctNQpXHbBo59jXFI1ZzjpsD
0dCMtfBqxbE7jTSpGZ8m/ECod/FNOYwwZ9YJt1+TiyAIZdAg/UAI1WaW9f8Zh/YMrl2oL0ZblATe
O1oGRj/0SRZRZzRGuuPMQso7tIJTZfohsNQXyb+wCCxbl3sUFY530vv4lAiA/hbmpz9/oHZy145j
GPSfjGZQC0m7lx0prS6QxXs0gWkGeudmbmG50TBveTp5oItXvURXoY9kw2aq32520zyXTT7RjYQS
cxqFPbUQv3Uw7lOru5oGwNuKV0g3j4b4I2TCZPMfSze0V5U+zO9qbfL09V2oOTHmpfXmixDDw8Qn
I2/kf+UC21yQbXBWCuHpKJxNhmDhpL8MjifTV/WA6YNcmk9uiYXMelIjDLbAJQdV0DQ0nZNx8dlE
LGJdMhM6/HFQyLXFOP8PFDLDRepF2mzYXcKBBgeahLCjEC0wJBwwY1Nxqs+rzwNkoMKHxeTHiEst
vS8FVfyOac6z2uQ9NGHmNCcDxmUoIKXXHdjcVGI59CLVljgITtJy7FGrNgth1OpHetEGitG4EWJ0
qoXTkiJIATHR0EUul+wtoWV+HIe5TCJ+F1iWMp/ouGoYtZAxpkjxnD/CxqjPeS2/6jaae1umV8lN
prn8ctuPt/4lQQZKAq8MIhxDMGbVSsTBM0ENsJcP/jtJ0vkzoKl1+53MnVovgG+mNumQr9jzYAPv
BoMiMQsSgP5YVgyVJkaSmQRObfPFLgNNK7BntU4VdCZn+3MVGJiqAH2J/hTx4emmFnvj4akh3I2d
McfKDq6h7eDCKoVHoCixDPerY3e4FWUyx7bSSikn0ect6hNtNwsmTK3buSYjscQjnS8LyrJhpZL1
0D3AmIlKoRapH5Vml0hGDFjdsGUfMTe4dc36YU3cnavUjNmZwW/Jez3tIyrOxR5JCs9NvVOYZnVW
D9Q2dVk8h04GmCYVIem6WjupXU7MMXIWLpDQmFVQ9lBSwO71mh4MDJUQpl35O1AvtVmw8OfzvKwY
oKTrtjlOS36I+0rBsqgsP49XJpJgb81KejmucXghiBnD65IX2j/TrtFuNTLrTzhx4RQDi7+3l/vq
RCh9mOD60FqkKszynnGYQ38sBVSk4LZJpmQDQxsh0b9M9JXpJWzZGgaPjzKk8En5loTW2RlcJpG9
3GRv4JKMz0TFyMDjNQ411sAF4/nDCRBLPjq0X7tLgXqbBGvF8MaEPChCnInDY+GFbmzf4Ug9xv6N
rGrvx2vY6Ui3J5ROJoSWqa7V1MrsvDRf2gjszdtHVJGMerLw0Xnc/h9ynQL3eEDN48kSvrR3vYd8
QeNv1776rFdYxHWtDbxHVPCfVIXCwiyKH/cVr8mw+hhISWwdPM12kmoJ03+7l22ZXtdSFe9AL+lW
S09TlEYmHKkgr3tjd3nwMJrtRtcH+LyKFcC4SZ8G/HYCKz2xxkcnQvT2NciKT9OvK+xuuK3ZQH0n
CkylqxBZTAFajtYCVx63XqCQzI5EPP5ynZ2R93+BPkQ1xTh41mBiPU7JIilrShDJso1CTQvyiWz7
MwIH7z2m7sfS4Q/WjPhnUN43EwF50trTKildCeVLHlPwXI6uNh8Q6WDkb0jnM4dQ9tkVfJVafCcO
MNPBsPFTJmOddjZv7+CFldasUV1xPdZBYpP0TN55IOCWesDa0FZpj0OD2i3kLw0Wa9rXVu+TS6xC
SbCk+EyFYQPnmxdQn5qUb6MsonXGR9NIPCQU5YN2bqyxh6KPWBkRWEkXtNitVu/Cpb/7rug7+6t3
V/b+cVWrYg/MzM649SpRYeRoZkh+dPckWj+UPmMX3slNtCIYvDeqkWQdOyNFuB/hmbqXUq33XcYY
8Bb/KRqJJ9hfS9TRhoW0Cff2hnHsv0Fh+FagQRQog9pNJkRiKUUmu7fNHbJHTHcolhOdbFR9jHwH
OZy5U2J3DsoWAYH6/LAOPMhBMq91vcaS0f3sbpLyL7xrF1mx2FRKchbcmZeds6ThxHGpeum+15r1
4Ue7hcGtacDGoUj0mSvAIx9qNP4qIq5ZG84JY8Os69khPlTdu2uKdI8XzQmth/lQaJhnlWf6gWP/
ptikPFAU+oE4m2lh+r87Ka6MdO5yUdBoCSaC7KE8KRRG3qf7HbX7esNqal50hFkdh7ZTelfGixUT
WZy672bBCOSqYEXC7EbZ5zdtyRcunVhYbe7jacYQkQH6GJUnyu43lAKgI+ybTt/4GaVxJmoina0R
J8VDBJHxuAAPlZrk1RP6AyX/dLaBqV5Y44RH2cs+z12InEf0sJyGZ25uwJYtpuPJQnDwiW0oLv9W
0+mcUnylP+Bf1SUwsOMkE2+YGQBghFFzSo1fonbgaQQLaeopODBbhWV3jsDceafFFEtXtSgtYLLu
aN2d2mzKEQhMdbaaubZWr7E/DMqeJ3CuV3J8ZhFaKConxeUXgbgbBS3bkQdEaZhmxPQwYxPbxd6K
ntTpOmAPC1lO2jjGPXru29Tpm7oedT/+QJwGEWNd2bloOq1pRsOO9VtfSuleGhpLWR9Jq1d9NWqh
wCNTcZvXN98eyFQDi1/VLcHp6GuFqpi9GoTmw+qj0mP1OMcpZy+hBD//DqY7uZgrDvnhIkzMDCZ1
0YaRGcrZFRUq2Q5ki5xqCGJy6AhOCb+PSXKsbg2WJVpXUk/Xkd9PNa/MowVR/oaqfQoGBz3O2tH9
t7EAHKIQ+HmOAVVu6RwLHI7mntcjxKomsvqOXsnT6ahC936dycKS1r7LAlK9fpTQu2jQy0s4Ti+Q
fwsbPfwg4oPITZi4pYDgTPLGu7bMCsYM9Lht9n41eiEoJw3aFTsmLY9xPRsjkckoRLsEaDslTMOb
BMe8Suj13e2bROdKkHQI52/JpXFAEOm1ch1RGj/8sHQLKIMj1tH+v0g5b22MdWpVz1FFm4Nw68g6
tIdkizvkclf6p2XBiJviWj3rSAwNWyEHA7UqPxSr9pNR8jDwjY1d/4kMYj9j5BEHD6cShNjMc3x/
fMcBejBs15skUHjT6lEpFLT44YrYLtC8M5PXA6cJZHlIo8//LpgN6i/o/X7ODWILOuEkE+QWz01k
rgTYPbzGFCRf1ttfP9RF2mSMfkdnFsm0L0NWe/pEyX4woJ8ckyD4y454U2KStrWcX78scOEFEAql
tUb/aRtmmqRBtybCAAf5yVmwJ546LKwN4vSOYkbv0nbMscXuxBaknJ0UqfDAWg1Wr3bkvxq3FiMQ
ssxKD/lxsi7akAoOcUapWzzF99She4DMaDNEa8GS867zEhKaMgfU/dBlOaCYB4l7sUmHhYn4j+7E
QUBsj50LKP1Re4VRCJOwlpwm7KumpEZnIpLBbgMxhHBrTahuTtWR643B3ZtDknGp7mSSafybqBOk
PcUtSzJrz3NxbgjHUI7pzRj4gLbIH1HQ+Ytkt16GlpoiaUcCuC+368Cv4i+pd+KKqb4Q2KLCJmkX
MLs65yaCRQFloGZ9IiD1oWbfZanOf3rQoNLhIEDdgsG0w2Py4y3enT+ECktX11u3PAdZ6Svy0ozf
7RIGxKfdEvsl64z5/ii+zVHLxNbFgZp4DvyRdfxgXaH3TEBWRrj09nAjU3+X5M1iVk6L8nxdaNUv
dV5VdQXNCpgfvztJCqPbN5I8efI2QhR79PL/ZdqD/w0lHzjtHNV50q72sN4SUIeJ4uKtuZkryrYP
JO2q8Ao4LEewsIbx8y/pQURAo/BfW0tHBFoTGtdFpnyxrpL1jhzFe+3k6m4GBhHI/cf791Je3N1q
pkuM/aD16kmHI9XCL18gQIbFe3s1jSVqfXnq+PNyD0RRWifshBbn4Lz8xXN150qntV0dyzHDXmUX
JpDkoEoB/w3G141s+uWgnBdMJDrDqFSt/TCJHrQDR6ua61YV6WOfWUmsUVWHsehRJwlt9b4qQV/Y
bhY6tylVF5wEsb9iZTHZ8FhvPNlNzwa6ubJyNbJHEo+okyZSI6jem7SrRivpWx6PPpK+87aqgVtD
RVtWlAUpm09lBvMSkE7mGICgApNVxAysc+3NhfsUWDd1WsNWAzFl8ZCn64FSOyNyzOyV+WV7DvfY
mR2616HDsvrli9nvtMBKuVhNZgg/R60JEjRyiKHYujL+FgUBvx0tW0/Zp1QmegqjY3jY8C58vv9A
hCRL6VhPgA7xeWweKwX9WjgbzHYvq12OckaIVmGpxD+Y+3Ebymu9UqOd9IOjooBdSbRWf1DCoaEl
JZRTztQwYF4+Cmjh/OlJBL/raZUlJCr2ix9c182RPa8aZ3VlpI0vDZ/yDeh0kAQOwj4HJ0phqA74
1/geV0o3b0OW9IrW1sTIXYsPVdAjBssMCWpX0daWzxzYMHPoJfJ04sw8E2rr1GqrvUPkuOrB4LsB
p5q6vgR6DHNkgZXraLo50P7tou9W5tgiTdYOh7r50K2zZQfggo9caKc01uBqLPz2R0VScumRwLCu
OqzR+UlZ/EhccZjJ4nqPKCVGKZdQ/WWwtKUZXC5B4r9NkJQEPp3JqnAi32JydcCsGI5F1h6oQDeK
VD1CbIgapQ==
`protect end_protected
