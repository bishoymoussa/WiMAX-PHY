-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
tfx2ZeyKSIo2+kwTAvitKogS8AxiIT5HFWHArCdAfzHLqlMeNvOh7Jar8GPSDxBKwqYaUVn8fwj1
iFuecyvdghoYGhKfb7Qo7JAhnbd9qGIVAT47HFtqN69UlkxAbFAKQAChq5ZAAIcpxMxJdrqXz3Je
FxuZqXNrW05ijfiN5138ddJ2fu2Y+an7SgoBhP5TgOMVhZiMVcv09BjbbyAv4qTP3d284XpuMxyn
q7OjoRpKTpwJspbdKRdKk6Vb39axnkt/XgM9nUD56fpR/DqPDdbO/pW/P0zz4sjCZEcvXWg0KJ5b
ZMnbLyeldhyAmrMh1819RN+RKGr61hrpEWrXuA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5824)
`protect data_block
eH96zI+0BzawVSWF74GcmbHZf3QBxBVGo0fS5cqaEiflqwEVn3ncVbLr4fk8QQJblDRAs/E9o7Ac
o7iXaCDSgfhYXQVOUzqBYSEQkHityCawozMLacilAuGFgu0ZlJoFFydDYGu49h+iRgQAITItI0ep
dqcYNVtcAtiC6y0q1uL3m+ixDs/bhtyFrDVLouGYqZOdroEerwgwqDUK1KkCMBYRrDiKIn3bCCpj
5YiFDrRm/b9raN/f3mq65oi6OK6WFucgYargRdjGb5s/T69O9+OBhb+htGgxzYLC7kqounWPcCw6
3z7/1fLbQ8RH5QOMLazlhuVLR9x5GnEXR3uuHvS4NdeUYyxeicUOwTXkTNqYnj0DGTuXAES/wmN8
/y7oI+Z5GGVVtlXMbL+LdCk4xYAFQWNz0yf2iGg4KVr0Xs+eEyupL+IymlWNNw2TfPpJGxC34tJ3
K0Doctmw/9j1Z4WhLhQTrYdAUjtn3DRjJEKx9YYN68SxyFLPKYd9yP7kSEcCgU30cRHUJXRxciuf
MzQcz9xYGtZ7fNHsCQ33DUZo/yj1bsInGGpih4MGRPm1824oNfz3tb9L9X5/zdamPLuLr0tvxfzI
MAe4QUO9CvvbewORugXvHH4b5sq0BFQnPoDDlX07F0RFv9m95ADw5ZyEnmZl9BeGgTAjvOkgMoIn
4XUKTXr3P8KWYgSOTIzpRldkPu9OHeZlk0Rz0aBDlDDOWCobbOvkwDo7U764zkltfuRWGrO5xN1i
OEYIH+NF44tkVerFM2M4ujg46Aw1gZ8J79bJEi+glUDkQLU/qv4iOk0coYbhZ92fjs25gsfCmasS
Y+IFYLJzqQxpdRuiC1z5bBR/Pmqin+wvQnmNauPEV4W4RyrJmTwBPBJ582rCt9KZ60FsX1QC1768
+Y1801StG1U5T4zRYEjZzjJcNTEupUb1qABbMJDxgE3Qsa0Fn0IHvAyJkzeImNfpS/zii3gzZ4NP
wxGjw23WMqYfeBumPutnYUH+GPAiFhhFsEytGmstJHt774OuUrewWWzcE0mDXuf7goZU2LFJxOke
/HKiodToPWjzvr3jczkBIXrICAaf+d34pbGqfXQuenDJkMksuraI2z4gLV9gWb9KRIR6EEF6ncHC
BoIeA71aaKRzGjeno4TFmP2IDYI6rjwZCVOYgKeHogXxUwDA2ZhFaWw35DyNc4djShKhwl3EmueS
9GvzxU6Bbrw7D5N0sVhBV5VauH3lNIEZCV0jZEBgV3am3mj1ax2zTW1yLOFgO5HQtJNT6ablCdMi
KURkgzTQZgSZfZLKnPz+afmymhIyiF0rc8hsXKND14AyRF3ssJJDykYBRaC2NM6uHPpWehS1hAKp
1mfzSY15HZU5BzUCAWMbO8OsMVRg0//yEXWrcSl5Lbl0Ar9+H5jCmpM8mOd+PH3gZtzwjboA4A/1
SSnW+zSnaTwFuQgQP4he5D1bfCCIj2A47wORdN4dv6jkkbI4C5lb4H71aHEeQv3F7rXNueMFZPRT
wOFniDCuzixvqHrxk8zHbcad+GvxRf8Q9MXm93REFcfuzKVxAYCRJqsX/3Ku5mYJ7gbQKD9/rxSX
afhhLr8Ozop67XEK9MHeCQCOnQsXTbcnGUF5dimelnk7PAHEmsB8pmsdol4PqvrKqeaEZr5ZHr1V
4MaBXDqF5VhdoMogdCtunOJbjHYxzlVGfnDz299ZwOw3nhA3T/3Ykb+nC1Nrusu3hQsRCsXtaFh3
lbqQDMhSEW/V+CbWviHp1G2NmLROw8GdKZX4f83qO/tX/K04PI0uuOlR+OtrveJSDU2HQSrz1xoD
csWgSemJ2qgaR1DMWcqxk99HmNMbzRVrp9l8VyA+STNeMhUtyXM61VN0QiMjeleTt0YABK4yrorW
lFAw7GpHqyiTZfm75w2sal3eDUCw95Hyns+WJ3yio4IsUSWu5WdlYHpADm8vhDAi+yovOMPsBYLZ
7/+1w25t/Wjxv72dm1TtZxEUTiQOe9Oy7ut+icxLPsZumR9WLCPsCztIqF+6ucXO2VxgazA6+Gfn
RDYRUep4FHa488PqKJfoKA7FGDlqPy35Fa1705vQAbtYWO1hmd0EwDz3o1hsN9teBPCNYETU4g2F
F2S2PI2gYgwryV5WllnCZBckkNU7vbqUvSNC6qWq+CqBOa91JD1xZIiWtmJxhR2OhLU9KBfEEEqG
HLGleUDcsz+A79sqpr9feV/TJsXk/epc9fvQuhewYOwX70PK2Klhn8PYVDR5CllBcNTQERwV7Lfr
w5jXzq9JvzhhDtiX4dWERxsGy0c8CCobVRPnxzZcZgIRcAhACWoAwZ8GgGuOsqllJ8yham3zKYSq
cQ11klPgpcRRtaTXuES+6i5D2cZMOapLPlU6nQcSk+ljVy0J6UXlwaYfLNHEVgD/JeeGVtZevAFC
gj6uBzRUhK9JOlTae9xjAOvb8EcmZEuenfxIhwyVdVDrpragpxhfk6QWLPlfNBVArx3lQOUFhPQ2
cj5lcDYavlzZr9Voi24AtAVm9bXh3WJuT2yDFiIMMw3FRogtc9aUmqqI6IdGMJeoihrz1412b2Xo
ie6UUZYVDdMqAGWvnBcmgY7vEYGgcFreLtS/uidoSB6N2VPyDLy5civM9833TYM0vtrHEWYz0inH
KIuPOkomBH9dvMJq+ODXJZfaSps7qv8kSKPgoOPlT7RlqySTgjVkHnFlUmfRNEK3YfLxotaRacuE
hrm4ZNfj+VFW4WRwEX3DnMgug1Ia800KGJurhwR0OkgPQeqKmIuR1nBTdQOXLXoRqljoOFUHWELG
MISk5XWpJVurt3mtzQyYFzlw2Pq5dtS0dLwG4mYh+5Nr3U5a/WrSn/g+/g1ZNr3jjLNyPq+RFuJd
GLKZnrG7Mg2wR/TPkDiIl42r75a7Nt4rosrkZYpnoUx3h0g8C4lD4PM/JmNYQ0jemkBTFTJQw1/W
/YhoCQiH9Y+uCr+e3WOZ+nGYhUn8JE/7e90EfLFRaBhLapPCv3qhjZPEbCfGNO3MryI+AwmVNXzW
/1WXClF4WI1s4cNfTXtD7FKOy3z7IQX9FQKzq+6faTof7usBKighTfjZruSJGddvSv6HK4W3/n9j
XSOLACAGCfD2WyVEg/bA7aZ9yvTU846h40mTyjeKahQtUJij53bNTon7O9+27PLLe7CaUN8t52O3
d6+9GDINadb4QvGnP9CXupqDniPLFFpTaSbwjo9hh9dUriJqrZ5GePeRtfoMtnI5MKZx3WKwzpWD
6r5nudTGGrQJ28tCDi0b4hZzAhHR5HaiC4NmROS1AbXnNuoxw0UDsjeDIQH8ji/RT7HuAoP25SvY
hODEJSnt9XGaCBsiDlW0Iv+30Fa2hr4tBAj1N6HDP8rBGkNm6a33FQ3sThWiBQTwvaXfkzkoLLac
qcPjinLLXqzjCruXQ4jzn7FOjtSe7nLM2xJPGSvNYQ9XOVfety+n8svRl45bSBH3d2N3N7lJfZmw
9wVXDBMIE18KtlRs+0cTDMuefodzFyYEpfWitIZXxEiVaoGq8Ju/I3r99nrQl9/FUxmQuv2ROB2B
YsZXMJVuoiu4VksC9NmLJmoiuA8NFiUS1omEtF11tahCgcsFer1vDPTmndIewvC45qdsUl+vZ+to
hM5zD5CHSewwvWvZg5CguZ0zXadBtwDz2gZul2fCHzWQTUsS2lauvCKcRUDH8t5euT9A4ytKXGB/
dkdfg2RN05PRTLiBZXjSLLRYFWqLG8NQcNtL2Gt7dzYprZDd7vxpJ5tX4kc7M4QnVQVJXjoSIZ7d
0259sP7dQEKbOO8wZMKsv/6J233RvMrkBXKBHCNbOLjI3+2qrTHrakiuqbzKGgfBx9Hi3FDBfe0s
RlxLRdlDWmCoK01rHl9wIm8co8lW2dMqmm5FPCrTkKJBlJDzKlCsTJ3K2wGZcD5Q3GMp7N+i+oPO
SmwvC1A3LLiDIgbDVTq3wb4eN6LgPq6v27iu78ncK2dv69Hc6qA7eLt6aHF7V13DQxB++G8YWuje
0Z94k8Mp9uIE8tgMDpMyVuljqyD9VEx8CJy+Z3s+4oYwNl7AO61Dpx4KQ0kzkLGEZ9UgBtDVF2Cw
q14V9DdTnV4brAdbKQ5uvkWHrCstipE/IvuV20NA2JDuD2opGmbHS43GsjB0x9LBd+aHTOmwm5Mt
IS8qPWwczQqwvrYzxd4F4lH1qmjjTrISNuQVMgvF4/F57hTiGlYJPbcelWO1PkebyF09XLJkBCM3
2MvGGPc37MKmDz6VLwm6fOU01J1g9kxFQqVyjdrQym1NCApa6Fg1WsYCe7XT4n1lkZCwjfymBbMq
GSjKH1ywF7ITMvNkXUhitrUHERcY0JWxcpEYz17zXZxXZ6SdW/smGTdEsu5obm/PQ3SBo+LkySUc
TbB+r6IsoOTtyMKecJ6hBLJMyj3Q1ma5Sq+r7M3QmipB+/6TRvSoxprqA3nCetp0hJUilr10G1uh
KCkDRecQnHieTmR0H7C3/JjOksxYEV7M1YRE7VA1ja6G4dNf8JY3tnISIbyBgPuwEVIbkdS3dnUy
AY25ntMSHoKfxZ1CRQGfBGqkrs5Q89Bs/50bWNqlxd8kMikIacjKZB7P89F+tIW7gYcbLFNX0SFf
5UMpZdIiVFC3WFsGvevc7Om1mry1whFcuiIs4HeGNsmYUCWAXI71trGzaPhcXGVayQ0NNhxVuCes
Ru3XGWFPcfahbZ0uKWkWzdBz55wryh16n+Rdq9oWJIpVrfC+IGWQKKZxY/93ZCIASNd9sj+vTGE+
tMQdxW55UqX7lU4vFOOyixepkXJYHTYh4icK66Wrf9bYFanYxspvxzm5ie/daci/u9NTpuO2EUgX
Fu1Io6pdMitj+qt7vqeSmOCMeemefL0Si70S98vqUs3qFZkLT/5o6mPPLfuEG29V1ZQMrEIkoJCO
fG3o+U8hGpFMNaQ7Scu/zRREJ9Xca62E7Fo1n8jOMfGbptYcEXWBt6EYHOiflrkW/aklW0SDj3uB
husGXr4oJEPNiSBhZif9MIv0MoHarfuuhEYNRolW1n2dkzb61N9rSr+ySLW0RS1FBkxS63YpYxv+
wwM8WYkiyBko80u0L8vel9V7cphXy2zEMjJrXvuV/BXhiSuMKhi/RR6ONKQCmSqpug+y7b+5UvSh
dBSdxpyWb+DkKqo+gDYLOVoiNlFkv41R1iU2ZvB+eEkU8DSyYk1grsWQT9Mp/NKmbH47fdrzIcw1
eWRlNjS0hmyWNmCMshhlB0LZ+Dg9UZiFEbSLRk6Tt2xor3eUxydDyzpIogEeibiVxvKkwS3Hup/9
QNXa8bW4tGXheLtJvFJIRwbRhzCmesGPWa6Jim3VlfmizMn30zZj+IfzGAkQ2lurvm4Mul3Y/GLR
TfTJHaC6YE+TFODXjmijnRMT0WCghvmZQ4Tw1P+RwvV1dQPkRYv6UkZj9frfdPvmWS0oDolevtfY
gNOoXz9K4MPKSt6VR5j7RiDcOOqZGxw2WZ0fhdo/+OwfPmm5LEaCL72Pi30BKhBv4yGw3AZq4EFJ
qtCHyIkcvuHz8d7FsgeDsVa55YriPLB24jLHwZDi+eLxaBq6w8pC0eyJjQxjs0ToMqEZ1akyzPXi
peSx/PqeAMIhgYr7RCAnvKaWHtw310gUtb/zZDXlyLFZtJGKszFFv9c4PLSrdQD7h25a5Ybd7UOW
PlS3HKjL2X2DY4eJ/5sQ0Q+Ce6dhj8RKRTmHli4DpmOgNxvaksg9ouC2wg2kKnqC1H9XbBRi6Ms4
yDsrCT7QnltZxqRf9QFfkqoBCCm/y1NnNG9Yh+tk9npWpO36fE79wl5t468gOD3qe1GkX3OINt5T
kj/SLiY3FO+ENSj4yL6nE7vVdz7YIcECK36IOdb7h401hp4qvmNg2mKhmmXOWG0XuNKZmzpEyEpT
3xXnnY0+GH4WnJhBwYtpVBH0qDoR9evFyqfSz9QN4UHtkrkTzm6XONbPnabhMEjZ0LT/fY2D4q5j
WEKv1rTSt8sWje2M5fkrUiMHgMt9xaetBvcUfvG/wW6QFwOooYCMB4rMJ8JKVnzDncBncMUO30Iv
vDQcVmv1GgNP7pMKJQcpyBBQ3zxg6bYPMJRe969SnXOhIImjqDScrdgBLt2TqFibzYawEt5vWuO4
gcd7MhfCdhMR+6dB1qPB197Yh6eg2DpVZCBVSipYjNXoyH+AgclttEDZMnTnsP2H/ko7oYC5vFgA
Mb0II8vyDtAnw99CeonA9uttJicsZWUVJCV+BSGmtIgucheVpb5xzN9p+u4U3Yks1Qrby+lMfu7c
UmvTQfItvGuwwspL/BA+gqIV2QMozcoy5+9XeeMvSpP0yR5L2rzWze7fDeQWGVfts7TBUJxyWM8m
X9t84GIKr0lv8zjSTEd9ZOVOyYc75zNR/KvESLoNAC4FVJtb32vwtxcCiR/uYdeyjCjwm2rCjDqK
gYiUWLeDyzEN+gnKVIzR7iYen2sXx6BjprY4HJomvHWdxFNQqdb2PY+N99sough9WU5NRF0+l9ow
jDk92Rqoz1+WPKMUEgkfKDqUZUfWNfQjOZHIdDLaODMWwySsrMEAz9pvKgnx13m9cqI2gA6bvwMQ
Yjhc30EL7GoHSpa0c8TX+Acq9q3+OVxEeRQdWXTz6P4wPDXYRhEPUHlvysTevEoTJ/UA+qev0fR6
tudHRvvwwkeGXKSldSS9IIIacnEeyl5cdkESGzWKNOaBidzFlj30NOzl4qm2SyYb9Ddd7HA1Xn6G
vaqua+Vk2VLovuyuTqcfLNH3NDGIZoYAJCueVdzLAlX9Rq8FywX5+E0+j7/zOjLO3wLJj9V6fXvZ
Yi2YfC7XYo3az3x/Bq3il0T+lCxMzeIWEbTNW5PgFtbkCnjM/nrw1wd0A5oQLxPtIZNiqA6rxxR5
ANOj2WgCw65H9dK1Bw08nNyUlppa7XSnCtL0B8RQrCgtWkm9YZmVHWZ4B9Tft49VdMunJbyR59tu
PMYaBLTs9iuhprunI9ozAIWZJZhaKfdck23TKkKByhAYqd8TGAHa6DiedunVuELgzFY3R6fCggQ3
mFL+przFC8YjFcxcmADsWksMxxW4qQLMXI+HYbofubU3JpyBPHRIYLQJD8x6w9UPaGxrxziVGc0Q
2FN9issHOyXqvy+MnhBXux3lDt6jU08k1lZA+cpA4EHoI5XH6B2cjS0B/w2yBcj/WTwGr6MJQ9NI
FuWlsneZx1iSdhUhxwWYvWRMhHSfWwEPIVdMoYEqGzfZPWaP4JSa53SNu8/FVFgSefwK1wGEGQx+
GVNeIZchabnoPhsOTDfP+k50/dlJSxPjo3f/Ci2SBQZCLIFZtaEZe2WGO7dcVEYch1rNej5KM+DM
CfHGp++AtFCMntElBYODnSfY5IBsjhgf8EUMfe+lJ6z1wS1VEQwVwUvkjtrFDSEUQqFV5hFuYpuL
bD7265ALKXpek1Z7zewFfyB/sUzB0XfmHBvTcvaTkjf7OS5snwpEFqr/hzX0LcsIlFhOqWmnbvfN
5+mX/YnODSb2xkijMoS26QTaly4GFLLRXfKnC7J7KjajFK3kqpLfFiGfY068wWsaDXLT/191vHRt
yH+1SqVWMZ3jRpAL0KKmxtUtv1oVuA4zBJJcwzPQjDogd3/UquEDI4rbUIOi88N3gGmry1+isoMm
AZpLcfqI0Br+ADju7SGwqRZLp2+UC9HtuhIsHGAz1cqh9NncX5z20KSiKkPkkYV9Z+0JW7XTJBLA
Pg9Ix7z9fsC5nw==
`protect end_protected
