��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$Rx�y�<��wA�*;�x���@�̦�W�X�fa�M-$u����n~�%���P�$��W��kYَ���P7�?UMfT��q�6�U��k�>����~�\N�(�����X�e���/6U|)�X2pF�]$h���d.���9E��WG��L�X"]�Ad����ľS���8od����e�GT?y	7�������ݵ�^��R�q^]�鍦�����s�ae���h��L��P_���ާ��YЭF���'\��68�b�[����w8�[X��V�F�0͘3����q諵�uW� �h�u\V�?@��_6G�_�*�G���B�絉�f������[�G��U&�����~�F��AׯK1�`c��[<��FY���4I� �#�G��x[X�=�Q1��`��R>(�w����R�O�?����7�,(�H\�#h(W�EH=�������yq��Ѿ��aF����:�U~m<|��.��0=�P/���4ǆ���T(�����3�{r�E[#�
xr�k��'m��S�6�e�4�����L��'��o2���Z�
�@����(��(VQ[���e�S� �	�I`[ؔ���fq�Tv�KV8��f@�tb��o�_1=z��Z�M���mr6�N<
�a��u�9ҷ�%�~.IoK2��rB��[�m�<N���P�� �In�c�6�*JCyǂ�<�{�gb��w��l�m�׹s5�qN���m@��Ϋ��3�߅9�47s�y�z�e��.b&���}��ppy.N��\�4\q������(�=���a��3Ʊ��B��C��b�p�
,u+\ѐ��y���G��|���a!�a�j~�겟�rҒ�'�β�;��e�l�x���S��%O?l�`�#r��*��띭�أ�w`T�im >k~�5��V��r��n���YǸv��AT���2 GR�����ݺ9�
�)��*(V/�׌�	�(�
.��f ��2�Ee�K����kg3`ޅ����g!��ǝ������4�&=�$7�j��<���KV���]�w�dF��^��z�(��޸�a����b�<���6K��W���s%�?�x��^z�H6zI�ܗ�Y+�c�3L���"����i�31�^p�=��?VJ�k�!4X����^���H�eC�.,rg� �,U�g��G�����<�V�.��vc\L��z�W
����8Y �x�ظ��E���v���x/��=��&���`�Z��7G����F{`��9E������E�rR(�3f�5�0>��$��kyϸ�~XY�ۤ���"&�z�y-��Y7(�9�(U��܏���PJ�Bltt �@ן����ՙ1�����U�)f-nZ�D��_����:�x�����=����ֈ���N~OOp�K�{W�'g�L荡��.g�`@c�ʐ谛� ܂�5��x��\e@�"�'�	�ˊ��\n��i��Ia:���r2{��V�s��$�����ܶ���u�IҘ�R�vrKg,E�kZ4aK�/��|��g�X��P��akY��k��[�$��j�N���B;S�['b�ٜG8����A~L7aD� Ƒ��E�˘?�x{6|n��I�>�||���N�����݈+���aᱣQ�|��]2����91�������?@Y�mB�h��?��`�a �xK�
�� ��+����^�cӕ��un�I���(��Ƚ�)\vJ�@%�ʵ�Y�`�t#�3ӳW�,3[����$U���s�ȋ�����w���EC�&��nI/�u�$K����e"ݕ�[0!E�q�bu�RJe��)��͙4�Q��w��O[Ji�R�x'SG%��Ee�ä'���$�������;����X.M8N��>�)�����	�@�W�K���
�A�=]!N��Pk�Z�5�I�h����ľ��!(6���О]X��-��"8���g'7�ep�+�q�����j�_�� #{�)�c�<Ǉ��y(%4ЩNH�6zJ�eV]#�M�OGAUQH�]@�@^+%����
��5?�����ح;�I��m�mBu=�g%��jmwrS�:��k��D:J�ns��p����SZ��O
e�-�/��y�c�.Ґ����T���Js�J�!l=E�(�ؐ �r;����L�Vu�G����`���KtCG�TzFa�J�e@�ܙ�f�p��ľ�<�oִn��U$�!��
c����\�Rְ�|������õ'���y=�ŭ�7�͛����r��Fo��w%5tA���ц��󘁀YN�l���A�xb��HH ��p�pӋ�<g�0vowU�ck\��U�3�0�+z�].JR�P�4��VH�ft_")e\�Hw����!Xo^����Qs��U������/�R�v�2��P��y���w`)�H��GM{�����2��肐��{l�ɖkǒ%9�:6ۮ��T �R�Ɩ�S���
����y(k��L��f�H0a��h8}�����Q�P�zd�K:�S4��x�>��2cL:g���I�I5@K��UX��Fe0�Mm�C�<��JT������F��-B��e��q��t�0�$� ��ץ �l�`p:���~9�h(θ_��#آ���~�����ZN��3����m�5�d���݁ KN$�;������^N3������2�/���G9D��^"p#���PY�F��$����z���ݕTuE�	�:[�:�h�;�3K���}�/r�:`	�u%E-�HO���l3О ����P>�E�;4�˳шM�;�sN��av`�.ӿ8l����x����;,�q�Q�P>� �0^@+6D <O��dv�`�1�w��J�("�~Q�J���*>��	��hRG���S3I}a�pXA��إo�'tD�څ�-��m�	�� a��sK�;,�^�+5$2��/�_lP7������u_ ���/1�6d�)���=XZx��Փ���n���X��>5�_Q#X���7�]�+�!�8�����L'���.�o�A��'2��c*�_r�Z��_m38Cm�ޚ��\I��dCq,;IM�W:��~t��qc,Vj�s��i�4@5���|\��!�]i��rCc�"��P9�\9J�������d��������!֪ �{"n�}0�݈[�Φ���m�W�3A���=Z�X�cY�q���?���?���(x��1z[��/�N�$���<Y����l]i���Y��ٳ�:�Q�>�R̊�@Z�<^XE�5�ݓ�K�M�d��xp�t_/fJ8��m�AmpNm�b}7�����t�U��'7�+��
Q4�E�
�T�I�dX.�{[�m���	�ɏ�:��+.JD���-�O@`IB�~VgZ2
�����Vx�ͩ��v�X���31����[�0���\�W�&�/.��%�iE)�0XM�����W��s~\f�;�=G����h�6�V`�����y�H�M���L�ՄOؓ�C�	�:�sJ��&
=+��n�tmpܟ_��!�o���:�sJ3#��N$o�Xwp{P��x㇒��d��i��#ū�U�c��c����m���R\?��|vhfg��3v� �yf#���s�gJ'm�q�%�;�:�[8��/�>c;�d��Cut0<�p�� �fT���\�]FF��ꥤ;���FU.ajW;���(�l�=�;8]�u���-As���@�5e��#Y����vB������S�L�<`��n)[L"��-��*TIEU~�� c���+o�i���)�@xR��I/s7�w@_��?��-vwv�u-Yؠ�v��R�f�O�6
8�g��J�S��\&de�ںB ��Z�S��Q"u�̒`��#O�::ƹ��>�� o��R��)H�+^q��	��ϱ��h�U����î
�{�.�p�!��?�{:��#�R̴ΰ����'!�����ԭ���LO]S�����߅(�QC��r�����B�J'SB�@��ۤ\�:*J�����W��t*�?���>����)���3T���7��"4�ym����������J��! W�iϯf�S�΂"����ݏ`��
�Ķ8u������0f��^��#ML�cQ'э�ߪ��"��kd���n���1
��;�t��<��ǂ���@5WD΀�E�Eqv��i�m3���w�-O���3���sf2q��=����5ڎ0�������SLHG��H�.z���љ�B�l�G��}�Bf����"�� �^62�H@�����b��nt���ksG ��5�Yk�u�A���}�#�D��1�� +�����B���{fxML,$.b��5*0��	�c;U}.�>֮u3B�1A�T�N%I"�_��
g$q�P��\�T|h���4���(�J���y��4m�[1�(���_��}>���[MO���{�K{�\�2���>J�h��A��b:�[� � �1r|I>(n{�	���	]	��D@�[�٧�?�ڢ�B���a4=��������J�+��
��JJ�'��&F�|�>�{��N�����$����Eأ����J��Z�Y��'ȍu��F���fR�E�S�`�\�T����]��>�z���) �U<4��~����9_8������q��ڏt�+�v_H��3���wO��@������%��Tд��U����q�VעZ��1��u�����}�K����Σ��fRi�������3�7Dߖ�b,�́��W�|�z���,��^��C�.�ڣ�����̆RbU�r�	���+贤�0��`'������۞�i�����U����S+a-���aB�9\�*�y��C4:��?0Phl��'�
u��mRXP4@�'c*��
@II�O�Ͷ$�ۏ��=CAIG04�I�p$�	�c�������,>!.'��O��)�{M�'~��[�zd�L�:�G�	��c����i蕱���T��}9��>H���8�>�&�b���i�2�5WJ�w	�1�P��#e��u)�g��mg�:�_mߊ��r��ȟ�{Ѳ�e��z�d8M�ۏN3��V��~m"�3(H��� P�q�C����EM�0[[�v:��i3���8�o<���v�q�{?f2ad�[��]6��M�^�r/b%����V$�-�V�FSh�㍅r�o �5ᗆg�ǽ�:|-���:�?GOR�㕾�޺�&�c'�?3+�-QR���yd
@d:������Җ�p�.��9�a_ҤSIx/;��хZ��ld"�@i�@��IwuZY��|c$���zٶP�/�e��:�����=�y?��d�'�gN�'Ul:�@�s���0�R�켁�U�t�,�S?�}�O}��ٔ���/}ҋ�q'I.��r5`����h>I�gIM᪤׫.����&�~�f��a<�3
%F�X��n�	xJ����͞D�ҝ�C�6 vu�s��{>w�w
�buE�_���J�����~c=�<Yά�5K�EV�UZ�=1�|�+�S\}���[������*E�j�Ԯ
�P�B�
���+
Lq���(�~ ��'�'�1�c��4�o�}/�J��p�O{�b�aSqd�v��.n꼡Op�����i�%=��9���)rN��ś�[�	 �>T.��� �yԪ�wwv�7���ӄ�E��h]��s:��ƏFt�P�7@�p�0$d��Jal��	��x��B����[pt|���e��W_R9v��-&j�-'��;a��V�GM��C�:Kv��tt'p�k���˄�Pƴ	�p�R	����t��Rp���c;��u��K���J���{���uq�>�����$$��ǀJ׉���vʟ��7�j'��j7�z��V����^�n;�n��d��\�x���PY�3���'�)0��m��.O�w����u/N�۲��D+8�m�/�'Lg���IvX�O���D��;� /σ�0D�5�	��"�k������L<r�g73p3��O�DE�(�K�,O�:�b,B�c�%#��^&�0����6U!-}q��W�u��x��=X�+��j�Y$��1�bJg�m?�
�%!%D���S�1��!��ђ/Ɔ����}�_�yD�.=�B�8�'si�yC/<,�Z�(��|�a�B�e��~����U`��pF��n�Ŷ`]��p�%.�oղ������9U�|�[��JT(1�_�ϑ��u��\�{���&Y�&�:����[%=\ �S2�Fn�{���8�E"�J#��A����C�Y4���@�Nc�7�:CƩ�/E�_m:�]r;<�I�*Ql,*9�� ��RH�#q4 )���j�3��[M?(��n�*':��KKӵ����J���)�.Y�؏���:QbZ�0�P��z�����<i���ld��؛^U�Δ�j�jma��V����j y���\m��w��[�9L�*!��NH����>x�a�"|x�fD�`M�