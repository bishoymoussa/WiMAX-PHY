��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$Rx�y�<��wA�*;�x���@�̦�W�X�fa�M-$u����n~�%���P�$��W��kYَ���P7�?UMfT��q�6�U��k�>����~�\N�(�����X�e���/6U|)�X2pF�]$h���d.���9E��WG��L�X"]�Ad����ľS���8od����e�GT?y	7�������ݵ�^��R�q^]�鍦�����s�ae���h��L��P_���ާ��YЭF���'\��68�b�[����w8�[X��V�F�0͘3����q諵�uW� �h�u\V�?@��_6G�_�*�G���B�絉�f������[�G��U&�����~�F��AׯK1�`c��[<��FY���4I� �#�G��x[X�=�Q1��`��R>(�w����R�O�?����7�,(�H\�#h(W�EH=�������yq��Ѿ��aF����:�U~m<|��.��0=�P/���4ǆ���T(����l:^��$���)�q�R ⾫!�2��s�VX�L
�*g/��-;ɂƊ�_�_�����rS0�t�5� ��u�b��=��*�jD7���rg�QB���+W��;�������G�?Ǔ6���G��+�k�2x����*[��`SE*��s��Q����4�z��_ |��^��-u���vV����%��:��6驩�0�y�5��\^p����2�k�'7� �+y	E��FAE�����T��.��> ��j��(4s�j�6Q5̞��6(;!#������$P�̔\O�� ��;��	�[��*�C*Z�"��R2�%��-�m���V�^�v��������z�Ƶ���fS�m�G���,oﶏ���!�+ĎX���Cz���$�Ё���5�8��B���i�f�^����O�rN	�AԊo�:�C~��z�";� ;��Y��me��xo�1����-*7��{w
���#Q�:�e�~����*v��o��!�oL�t���|Y��/1I���!�Ѓ)����GQ�5^�҄�,�XKӮ�N�����0AX�L���Z2��g9�[
� ��/;����2���hL0���z~,���b^;�oec�'|f���aD���S���e��k�F5�5��%�����&$�gc�N
@�L��48 �(�&����ߢ�f��5?M,��߯]�ʛ�vj��^&��s�/�K+����n�Pȱk��"B]>��S)	dpY�Vy���Z�s#�  ���H.\6�EޏX�)��K�U��0�R��ٿ�r����@bA/�FRb�cğ�/ޣ}��j�
@����D�����9��~���7�c�ߣ��d�*1d��?�[	����\����:h[H�0��A�-��<mi~�m9@���i�RF���V�4�t�ݳ�bN���x��әx*�<����G4iRk�ŕ�u���������W��	�l:j>1�4���d�c���gD�h�ƅ���Ng��F����*���p@皿 �Pb�&�u!��#��H�{��.�����	t����(��,*M�U�@�<�W`�hӟO�h�_+^��{���enA�ۥ�P�5�L�]f}V��w1�b��JC�m�F~g#�6M�}v�h.Fj��M%�6ӣ�j���IEAG�o�2W�W���EG |O�No�PW/���y�98��^@�E����E�6����E-=����2B<."t�A�v�-M��m��1q݇E%��贅�i�� �Z�a�i����J�Z��XZ������e�Z�F(�E�3e�_���%�[�`����a��, �^|�i$��~��z�7C)� v���(�� ������IB���b�8@��¨M�TV����?��)��R,^�׈�������#š����rO|}�$�P ���	N4<�oj\>�6�z�FD�&��,�%�(T�.�l��l��
�[���NJ����Dl��
���E5���&T&�J�j�v�`���p{��]\�P�aWgZ��N}�!aכbk����&ZyUx�yS��[����f�8������� ������ZJ�Z�x�(��4S)ts$<<�����v�@���7/`�lm;�N �$�{������^2��@HK��2��H�2��h���o.��TU�b�����O�C��� �*�_��-��b4	�����F:s��Y�����D�ң=|�/V�g}�����W��y&�����v�Ǻ7�]��J,�r
*��E���Õ�۴hYn�/��ڳ�����bQ�r���\+Z9[0 y��au����p5����<�W)��C=������p4��|ôӘ��U��k�=�jU�{���G���[f�Zх��9��=e��T��F��5/����(�Bo-���[
�r��-d �S�x	U�V��G%4I���[��7N�DI�{�㷵��tE/�<&	~EZ���:n�a��M�ޟm�x���]5m��t>����� ��|������`���Y�No4����q��?q}r�V�0!עP͋j��ҙ�V�s<C;p�=�U�\9y�� ��s^Ư�t=T��X�;��S���������1373��]F�}�y(�B9ɊkC��w�	�D�R�Ծ*��H�q��#>�뼙�1Ϫ��p���%@F tiS;�2�����u9,'��zW��<���e$JK'pab�"	���ڍַ�k�A~%��:%�(�OG&ط�[b���e�2�Pߗ�~�e��"r}_j��(E��hmqi'�s��
*���}A3�h��	�V���oDNHL3_��P3!��lW�b2�u�?O5��C#��+�]�y]��S`e��##D�Է$�H�Eq��-τ�t�l�iu(�H,+��V�ڹR�a�	�GQ�ge�R�,��W��W�6���0_�ae�Y�G�}!�v�=�œ����n�d��i�ԜnkX���3t���u�'�d�;l=
tU�SE'H��Q;F�x���p�4�Ͼ���S5O�#y4R�YTD����f*G����� p�������q����A�O��tL��8̰n��Uo{?����;�/�Rs8��a�hh���Ql��>K����-�����~[��G��v*w~z~���ٽ.[�s����T���Z�fe8JTWF�7�=K��'\�>� �_�;g�Q�U�0�X��^0z/__ťy�\7�W�l@S�qtX�F2L�R4��[��<_9��±�$QaB�c�nٷ�s�Ƽ���Ud��k��yRH���d X:�W�3����SD�a���H�`K��U�Bȭ0���)Hw7)r$U����̃xo�y�q�-�
��n86n��\���%�@a ��ډ��XV:�L�y
/�|/-�Â�DO�`�!�ݖ��n����8�S��۷1j�)���؆c�*P�-��sPR�(�^�j��"X��t�e�Q��]�B�=�������x�k�W_��׮dG�P�Y�V�#c���ׯ-b�3�ǩT=��)�����cR"c�}#����{}l�����+Q�b��zS*�g��b��wF���V��H�*��j���a*�R�;�W$m8�h�����d�3�׋Pi���r���ɬr����e�FrO��C�۟������a�U�Fy�{o�)��bEj��ymn/�U��L�N
�3=L�c���)�߬�VT�n��VF����L�_92�M5f�6����B��2������"�V��+ӵc��-�}haeb㈥Y�z�@�:L�5"�{����Ҵ�e�0��Ą�	�f���@�P���a:����1�A�%/F��W��48]-�&�VʑU�+N��v���2���uz$��o(b��~�t����#�K���7���n��P�7��,bkOΙÊK��ɀ�N����g�i+�Lﶗ�����������M�(HB@��`Oq�9�Z���	�2 Ԥ���c3CZ�7��Q_�ւ�?��`8%�ʆW6'�}�@hME]�Ԣ����)������s�;�(�YO�7J�?jL� �<���9�-^iU���g�����SvL64
u�yxқS)��u���w���n�.Nx��'��c�CR"�c˹`�Ql�\O��.�2�E�ρ��R��AC�����6
y6����1�ԁ��w�3���p�EK:�F����N��Ѣ�D���ۥƝ*v��)�"w��+RJ���pȄ���� 8���a�ؒ�����/�����YvFj1�SKW��!V�-L	�@Pc��+|'���S��H��������S�ln=�W�� �<g�|�̸	v��2%}EM^-V1��Ҹ@}�*����[������c�k����a3��A���?ގiM��j�>��e����-�4�����n���ٶ������ݫ_�s�:	����p��_/s����	�Y�y��;^�����bTYG�m4Ʀ����-�K�v�M�`}���Ak��u�%��fF��GZ�`����G�>��ٞ"� m��A#��b/��� (�l�kz|�!�$֣�k|ۈ˱�#�i>�9w	iݳ��J/g��lT>����M����f���c��.?���f�S����U O�Č_1���?��ZP��W���8H�V�""#n��Z�wO��=��_Kip%�_`�gi�B�b���N����>Dm�x��q���
����G�*���zW�������|YB}�4]J+R�ۦ�c�@c����N:{�Ҧ�P���ȣ�]T�*gdH��Gvf���SԬc�VGi�Z3x����s�f�W}
���:��D�5-��M�3q���JT���,*#P�@*>^���4��i9>�:։�x�'�U��q�C?�7c�VT������?~���%��"zy��G���:�З�h�\���kQR����Z����$*�<��L=v:�gFJ
��~C�B��L&c��ԙXl�q7X.]��v���@�'4n������_�h�o��:>h;��G-e,;��������8��Q�A�ETC��p�'pS����� �?�H.�j�y�P�x��.����e���X&�����b�٤?u8���3���ٓNI���-�hMyokD'�B�֕�?˴ij�&��	"��m&o��9��1R#�f�T��,�q�ܘ�2���W��Rb;�c�Q^�9~>:9��Kt�RKP�s�p6��_����uɇVI�X�[�x��ۑ�<�\�Q�un�!������o!��c�\�85WK!#�_�d�^��LNh,�3�f�@�������2l��=�����4�X ��֊���Ak��ʌ��¨������C^M�~�<�З:��s�;�w�8[# �Y��p���𨊭��S����?�&���(���NC�}��@!6��᧑z���霭�G�|	���TyU�ư|�l��.����ԛ�g9�py1W���֪sv�쵨�~��X2�4.\/�T���qo��U�	�MR���H���0D��(��z�e�Z�z߃.5�y�,� Cͪ��[���<!����Di�l�O�0D�߈6H��2�p���f�[��C�'mdd(尖o=_�t�Y�ifc}1�����P���G�y�@�}�ϯ3�^l� �����u>h�)�2rC X�cy"��rx�72Qf��T�U�6�rYWC�0������	õ��{��f��wʩWt{ l���Ə��R�#:�&���8�2QGSS��'�?:r�7��
G��|�x#.ӫ���"��C~�z-x�#�����`�ͥ~Z�(���6���U#Lhh�&īz�T�vJ��TJ�VK�}S����9\�&�a��I�	^����G�ԉ^�GU�Gl}� �/��N�h]�3�m|;����m����j���Lk�fx�)㬦��[+qX$��-��d2z����x�.��*6�_�y�B�~J�"���$� ��35t4�ICjk�Ӿ��oև�!�v�
��q�&?:F��YUZ�KLVs���$Y��\@j!8��c�p}��g�D
<�����{n��G�&���p�/��Ʊ��'�t����6���z��rƣ�CH ��I�|����l;�x�[�W2PcTM�0����	�:�5Ȋs�*����N�^���w�Yt�kJ(c�F �G'��ɝ�~�6m�!�,�������sW� ��/̐x0�}u~��E��6�7$[gP��5S+�0��U �A!k�}�ڦB-�Y��o>ka�.�1ꔑ���U5���e����,#���e��T-��;>O^�F%���D�2u�j��*T�1���l�g	�{|��aF���gmm��5�Ӌ ���۶߆��?p�o����G��Y��H1�/����芮	��\�<�o`�-�r������mvYI�`�Ti� �쟤"�j��ڧ,�������&�^
�aș�ߥ�\y��GD��ls�h�~��9LW��������kkK�*�6K�f�1]Q�B�����Se�eF��l��B��pb��%�r�s\�?�d!I��V�0t��	��$�n<nڂ<�w��o+6Ë��a�NP����1�`�!^͸����S(�+ �=���o���qĒ;i��uE�R�lP�Y
&�T8г�ڰ�'�.cX*R�������Z�:g\���F��/d�'�2��(��Sq��0��������t��K`T7:#��뒕|�o�a�������?C̼�&O��3ƛJ�� \��'����c'���q�O:T��b,/�����i�z^�<d{b�Y��Bڀ�S&�	*�tq�����$�"G�ueu�ǿ�e�~�r����B��W�,�nK!����G��j�:�����M�g��6��s�� �B{/�g$P�g"���Z�~��V��0u�#�S��D�'�	��WGB*m
���:7�a��4Z�n6�IL���6�"V%��w|ɀ��uvƅ����e�H<�kJyP�I�$q�Nk�z�&���WVx?D�g���h��NLxsՅ��3Q�ܛ�	~ϼ����.�#{�>��o�lx'g���4�8�3���NCcrV娛����kֺ�>�J�ۅ�硽�.?@�y�f�Ƈ��O�	�a<��Ol�e��?��8*K#|�һdj\w�NK븞�Z��e<Nb���`s��z�T��vXbAj5%�b*S�)WM��'�Fv/��>aI^0�Gޕ����pvg͏�7U�ijR���P8Z�3j�̻!3t1ũ�EG6����K���v������ 