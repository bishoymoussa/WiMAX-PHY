-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
K69ULOwQMXwAtBrPH+JaR0zZ/BYFKFsMAIcEVjs/4uM2Uv/8ubc0xQOgZR8vfCf2H0118UQdD4pe
vzQ3OVlwXoRzwa/BuPTwEfDA4OU84yO0fm6teRXTvQbGW1ulVgI5tgjvKWKoIz6VLLP5M1x0HFTb
lAqwEavUkkpvZNOxUg7fYuNMLAsmjmCJreJ3vDM46k7dLLsVehmiQxFfX+OPrvX5UJCGzjP1CeXF
QzOBlL/o9ruBhB7S57A9f1BkTVJa4ujGsB3wqqwFkvwlUFWjc2wNvBMlfW8KDE6XYyuYZGKcQIcc
A2Mn0qCSF0O8oG9Ik+AaOkd52xufAhhq8iCU3w==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 7664)
`protect data_block
ouJAAfEfSui36r+5ENEBZNgJmGw+rXuKxcsCoh2WXaJaxpWVJjntbud4SDf5Pqv3esyXGy+Mq+9f
oD+GKkOzD8xfzltO9VFzVDUyCN4pu97zlCav5unvn2+zRRYwyLDyzgkuUZHhGKRLFNqmVDIZzpbf
jWwMCrDdz1KH8L2iZkPIiThXzveAcfUUtx6i41FKYP732rrXLbnvmE/E2KyO1CwS7p59eGIJKBci
dIJutOB62t2rQQNJ15SEiwAqJeKdZquT/6kaElRN27wmva0A10SnHAvAvPAVI79x+AtooZ3uDnTa
bNRNWGpgH9h4fxJwDzT6/q2MI7lKynTIJdoOa2smDLtiMWX/dSiqOh7IWuHKDKqE5XbL7f4GMuJq
wTay+Fsuo9kop7p388qVOwiJfAo0Q0EwSBwBDKHDTOWdszkDSQcVShg+icHVbhWgDhpBEupuyneD
dAEjNvo0cOg0vnKPjylDe84XBV9qSHOQBTJq3p7MXzzXPaD9s3VbT5kJ2oUJvqSTDdRs/RFgYEDR
7tPGX5mnX6VColxt9+CggtJcMDiLLlY0+0ztyitAx/4KaGLWGhskJGQPsLDGatprnIy37QXT5RGg
GgXF8NF3hDd3LlBVOIJnQHrX2CzMgyMKKDuygcSCy5zzsVuXvvRrokFgmcDC+OtefJZvzWM9dVu9
rjgsAqysbRlLr4eudpwybjAyNYB3qqI5l86L0CWR7Eg+FxsKySBty467SdUGANWlHVhO2+qFk2VN
y9CFc5JjcJRN2SorzCExNz4S6RPXwNwuGjLEDPnxitNK6AzZbvLEalcbJZGu/26vlXlDjiur8Xm9
Q2DezvExL+0stEV0VHeXjAWsU5AL+V8dD0qKCPwHwrRRdYg8/oSXCVVSbshrA9S9yT4DZShQhS+k
QflqQ5qp8SHiYyr1kJ3joZOdSHJFzMt6HFkC6mopKx07xVyuytCma65gOV9ZK4flOmcapyzSfllW
UhpAP3vrz76QO2UHLuHREk84kH4pzzifIAKEYJysebsNsVKidFJsj/4mpKzmMblOgBFWqZ2FjjLj
TMuESWz2+1O8ME5KvMe2kWhER7KhVd4REVr/6be3NrxrwI0nBA05a3BCwNIpZGO7JmULci84hdhd
65LpUuS7JJsLXSh5ULCU3Wa/1RTuxpe0zpoy642p6G49mMU/Do3NoNw2DqLcvYtz4N5SqJpA6NHK
5CYtbFyAWZGtofUVLz27PkfDVzMY0VdsmoyDx26BmA7X33xayNi2YHfiS8PrR0QqVL+dDN1z0DLb
HbaoxPoleNf8x9Hgb7gzODe/J26HCXWnbDLw1KjarEFpvSJQ2LiYSAI5Nx+O1eZYeN6LazOn7+QW
8qDmE82M/Mzm2GdLp5ldM/blbtAaalfPWrFQ98yUFWPKuRJ4hlMcza/VxykKJtNLEHau0N6rM3wL
wmwMw4TptJf+svO4d+Dt2dAsoR4u1HaKzj751Ow/wnqEBzDJ22wzTyhP/FJXiq2gGmAo07ird+Dc
w9EJwYc7qmjtetnQh5laOCJlw4m3wbLybYFEfbcbPGJThk8IY2Bc2ABsUC5bk0aBjl+b7Dh3T8FY
AWiWak2b+QwIALE9zMpMXpiRuVNU3djwlVmGKhFm7EnylXxnCMioIF4PirnIbkvj6pONog8wSB5L
I6fOPl1IiW9GViOie3/qmjqGtNiJKjLWWuliarVn4hhq2JcIOJky6+SyEBtDbjxC9RarfbiWN9i3
tDu98ni3NVnNShIn2LtfR6Qbz3ucti6PL6P7d/vA/iEWjighMw/90EhQhdsaBXVEIrQg1um5eQX5
LEDXTAalaoPu4gjeVa35YzJE8UZqWEnRzBy+5GOICx7X5Mc0h2NKwVVxY+w6gfKZRbEQ1Li3Wz2F
nlqL8FfUr3hhkv6Ye2pjPC4Vi7tRUIkOUBViZpwYhX2PvYGsT81oXhubtXyOfJ+N0gWMh5zwmPJD
0gqbqYGg636ExpmKjCXNET5ugsNSNStI2YUtR0t17u4FOnhe0Coji+QdvGnXRVlsxPzJ+5flz9gq
233aYRdsNeov9LEj7SNq4bCH7mDexkJtao8NYPYg8Lk575rbUyL3Yt9IkFkReVVCqTNJkwR4kgEa
cD7HrjqvW4HhFZ+GlK8R/NcFr/g6U5smDSFa12ZwnadEoGYuyiduyWpF/nJxoAEJJfa+Nxyyz4ui
6dYinWC+7hBWfmbNEkX3/+sMr6Pc887525BkVmK+N8N1MHpE7GEjd/NlMyC/dH8FpHDAXPe7Ejxz
7PDoSFsZ8qLkPr0BAPFM5ZeZl+yyOIzmVL18tls0pVhtzFNyCud5AoB1Gqk8jP2nvy2OJuITg9kB
0p04AbOtX8jNgue6lcKkTmptWZx77Z65ZgkuMUsYIVOzl6qa8nZY2vRC8ApEq/6nOwDBWAMrWG28
k++KFfUcS7GJqVzjMusstWyb6qI1wVGbKX12iPzmuXWbilp8hQZMApS+hSVRAzaKHel+C4imFPeC
mI4gQA94EEQ+fSG0EXyNIJWwADntwhYG2M0QqClIObVZjK8m4IeGiEn7sqeI1SBrcpa5IksjUm9t
TxT5qfFElfnJwHou2mo4eVw4ZqDe2xSx8H78RtSKUXny3NND35D9LPNhVWNTZA5uTz0JpfpSHR9f
yw2UaH09dSzcCF+3EO6qkPzJR7uK8aejTNfyiel6aJIcQw8AakPJ7ixtk3shPZb4JT2AuDxAXpNe
7082mfy1EhWeF3KZxEZLQVPNX8krmu4+nZEuWgW8fETRXnfmPWaTNlE8jN3LUbeiU1O05MBR1wzb
77o5sJOVlRPgVzCNkB7i8zrG/58KOU2+2y78vn2U7bgawk25htR27ImwmvC876+D9Bg556z/5NOn
JvyJIgjMJnYLJBRYY+8PpNE5ZIQm+pBhhPSwiDpV7HnYQjJy8Pvi8zA1kH2osWs5a2oe8jJ/OqBB
g2YG8nwa37zfzABN1e4lGuH5OemVyI94TKqMXuzJAxf8VyjIhTmRgKFu/acU0Z+l8UwC4q44cDB+
sWL5PtMW13F7SvFblljr/9hORygg0aSaxYr3NdH5W4WnlZV6hpWZ3yPEV42fdzX2B6UMbEB6ie4B
3Nt47R1bC9e+5rlkZLf5t7jXeagX5/oX0T11VQRVVEWV5bgI1nFHW+V0zbJCjSdDDx+KDPRO7w4X
h/C+J3IrWlRhCXWl9rJABA7qk8kcSlFTGxuK6QP5L0CP+fNbQXny692VDuJEDj+YimhmpeIdsMJ5
ZTwkDn7kIH6Pxj10mrilW1traB1RIWESDdIErRbQ280GI13RSS/gN1UNdH2aOHvPYF3mRWMSZDoH
wP1WuXvOwQyv1bWl89140FKd5ikIx2Q702Yk7cHyi9Q0Jm2I6nCcCOZwI/mfdB1s9pNOnbqORzXf
QORH1frRHxfLYaO/U5rMP4dd2oxBEhWPqwuPBUwNwNwLosg/wGEfypsWYIrI7dgIqoKbBZhssBSk
YH/uN7fzRsCcUAt9C+iHgBf6IhY9EIXijKcPVJKiBi1x/BpYiSzdmg+4nxmY2/ACxalg2+LvP3nJ
oW52ZwKNXxzV72hDHgY1aSTEN1dlixL/ch2Z9rc48XKkPB9PEEpil7Pfp743L3xOVbR6ckzi5LLt
S3SFA9Ul4Bd7X+DmNjG8WYnECeBFQQvSwuBrGnYFRkzjY/RQTGyi3KvZSvDFAAo0UCoABGiTRGVR
kRhtef4bKdmU/0aUyVapyB+FGtdT3TJIMox47YXC1M3OyUEbSHDPLdP2f194khfeIpRV/8UNl9hG
ckTLO3OZxf9Iw/5g0cu7gi5QuF2GtXscM+jCxppDovjkRyua9S1pBUtb7elq/eA6tdStMTmekyID
r5vuHiqeXCcBuxxhrG1GT7ELD8xRikU8+Copl2Kj5fDZN134t3fPkEe6YrrJHMADpYGsA5ROoNqg
+ITJl+KuC4BMaDtbgRZu/s1961Oxx1ABoCnJwoA4RI+vJDB2shvdc9alhgiWKZFl6wNv3YMy6wHn
8lHl2mc7sLNlfYF0+SrIS9o4iFYvAQj29T5aZk0a2e5U7p3wdYOl54A/D1KBGrI6hrXphpgVYNJ0
7s9dFyo89gWPSVPMHfQiiV+yryuFF2U23h9+a8w6YGpsGIcnaDTnILiwHK40SCtGY3VjeugTF+5K
sFv4VVDhHp9x7JKSj8hY2g/lbDB+QVd4Kj1ORFqGVGAlNhLlRIWiD+wBa50NBCgWkfcgjfgrBEOR
2JxdpRRliPqk4rppCuBn+eYlgd0gsSoI71TscB5UTPCWVVwe1fsMcFzM1reThcYDdF5pi8yMy2o1
IUC1qTzGDS9GvsgCvFvaABwdzPyZ5vJmH2yADZQVNByfwRm99Y2WfdjcSvdmaDcO59CR8atWMR2j
RPZ4Orb4ftj9DyR+b23cJ3+EYxJZ1bal9urMMlNDlI05M92mdmf5og4mKRDcoUat8Isqf2IZ9cgI
cewhGUPLN1FENZEFL5pTeLMI2K1yZvxBAn3tTy60QsLGUT93apuHg8tmpE/4iGXr8CuBKE3PM6dK
XyAV+V1Y47pg4dEui+tEoGfn/SmZVCwraGkA1qCXpqw/GoRsaVm3JVc6pjXedygJyWkqYARMnNfP
Kbj0Ars0ecuP458D7PfCB3+5gl5YopoAr/4Prok3IweNTr+zlp0BtcLFJiE2u/pjBqyy9WKYxes6
eNgFlSQPAiL4zqvyw7wNGo/wgXU4u0wqoyTQBqFFQPwZANDx0yWYtkrWFfra3DyYzwtXnh/9ZLFD
oA+Kykio1lRvMhcRLJzl+9Db4oSM4p2aoGg6ByKHhH+gdmNTEVUHAxHuPYwI5tyunmeQsmmviW3M
HvXE2AyXoGTTl63MHwPYRt6yi7LYE4ZBRvj+d0DA4RKsjBqtAMkUaEEbTQfj9ZNfjLMt1L5zB8M2
LhwhivfRUyK888cB05sug3HERZiWvqTs+St0IJrYyEjF+Aw/CvXYWvmTw6YWFrGPCUleQSY4BxC8
7246jS8hIMeGPN2nUNoZERzPSgQRV2ycyCNNUD9PYwQkiV+1nobIs9gLZ2RASvpt93yK1OFweLzD
F+HLJrCDhbCA9ss3uAgcpvK9zZrbRPvLx+ER4y0QgnUgBusUhHCT9Psw5ta7cg06nfxViRym52ww
RXas/x8vWrLDJPW/Q136yIDs7DNXtA3yB1WHg9Fka66fUTqLF5sc0HR7dDcvgIr86BCJorDsJ/3T
EdtQtfdF0zNt4S3wtUp3ySnsBPJNfR6Jp2VFu+X8iIB8H0SMiXCfkNXit+f4O9eQh72dLzMZ35cX
OFkPpM0VvJTKCDst/P3gySOUhPAP7PQ5bdkZwiCfk5OGKhP4hhQK7g7xGNjq9CszQ69Ib1WIQFh9
FHjIx7zDqaBfsPT6fgZ5QfEMy2h2kfKVldE6byX6ZPS+HptgQXaMv0w3ozsEZMw4sXmK+MlPlsZr
NPCdgqRXZ3UZTSe2HzXxaLl0UM+yP9doLGZDFa+auQjKv2NrQ0bL5lCfdCwoa6R51T+IKMkcEfA7
MWwLVF7xtTPwyN5qh307IJBHrhhRaujBaAQpHB+TPAioK8We6EH1nha+j75TLE+j6nZu4C44Q/ER
6KtDr02/DWo8U7SiVaNymZMndXjwgBPalwnvyDN8GKl4f4/Q53Kwr2xY8nW3mwjNQNyk3Sk4+bxA
rHL+8LWRNCLuif/kC7q9yLRqhS0k1tQU2bCcc5O1jlpPc5bYPNbTeCPs5u5Z3QuxhJyDNdKCZnJT
aPOWHhE+ttR2urx9MjlNUPo7AwManVFqMAM6mxlv12RBysUs4kdDdsUZ30ABFJqicqTyK1l+8E0D
QiCuhDgCph6VkKC+AGMKDUpWKk74wFme2u3K4/WVGd0PBEeevObvGjCckJST8wp0eeJDnYxwRzL4
uW5nwgqMB91OE/ggRonWCEzu/Ja1E8CPB5xvpbXL1WqyRRlitB80uK+l6LPFRxmDPWZ3a284GnBC
8unN3Yo8DU4RGViTthesA4Mzbdz08UdAVApntG3D4XrUrml0/8kBL8KyBVCvsbL2up3I9EGuZULG
g5vhk3nw97CF/PzO4lc791nSPgb9aawEIlgnLnf+c83Tosn05SOP5P2xni+lXJsS4Y0FWlgeVegi
qDzWsMIvWbrFT70a8S6o4zByts7S1N6o6+9aNKLBXiFphJtkMs0iGFEKK3FIjPSXZv9OXFvjWdz/
gEnD75yaQESl6qZLouVs/BY3gBCgZVPdrtRSqhjlrZpceJkES7G1pmiZJglXalIJ2/dJFo+thdJ6
7cWeLO9AXOTJjs1g1HKOoN9KE/yJbjdl9RpCw2dmrPGjtE+ipQ+yRSN0H2TVYLmfXELvQcKY/6hs
6EoLeK+p6ZupOF4q57oOvwy97p7tcSBFdBXPc07NvRjO129yZapa2WZTZDViweSfsogOyoRYTlqu
u52GhS5ichclh/dyFbNj8obaMGlu/ECDxaRhDWba0XzLomz1r5nHsmTxlVFD4nEtXfvlksQVz2aP
mGCLX2sZAfu9gGAHigzbIJKCd3pAru27Rs7d9wIZhT90k6j4Vg2S7JjKMnzKWcuW9W87Phvcj3Or
YSaw5LmpzvGd62S9vlTZYAzxFZ6rRn/gw9gLYsw2VMQ1zri39qELNAS29ZIQ1Y6lGYi9EwJUuSwN
CoDkHbgbtShth3X+4dHfX9BwtWRsCgKiTuS9mPEs4+kSGWnXSPY7SL+vkqsWR1pfE+C5OF5699oZ
yRLchFnbGFg9/zxkD/34bmiC3fw/Ls6n06mSXKXiToKPNOFf8xbeNOWPuqUyk5PecOqyiTrGSixz
prfC+vF4ZrONVoi1kMQscsqbV5jE+ZexAqOz602dHTjbAPTsxatrT3N969f/rs4NyxKnc8fzIp8l
6oh2h73YGYjzR0JW6tOZdt3gFD90/jhcKR0EISBp6T5yxvzSVUkVyM+cofH/ZlkDeRIzZNLurSHa
pFhmV9tk16HXCJPO7edwCFa9VTLmnyWjdqYNrQry5d/TtuLQmW4YQn2MAn25nf5hkq9CjGJAAGnb
owJpr1FFZ1cZtHR2E+2f0mKel6GdB3wsvab4HGZ79Q4AmaOWt/UFtP4/GiwqzpDhemH4MsOF8tnv
wToBnIKFMh5TLYAnnMbhJ8t/R6T3vFdTdEzbEH2782KffG1cdzTD0CrTCRsnYmE3RnYGbLcFG9s5
U2y3Jtr9nbrm6qZiBnqJdRoUYsvYQhIsChsrT3ABpxTiX7N65szC/EXP8uuxQXKxIqR1S8739Dp0
gv6yC26u/OsN10stU/6b/IpexVlgrjilWPaCOIOaXOgnOQvyAqk0/0TkN69c73uRst31/UViucti
iaDqcIgXgcaAmgqAYgzeT0ZXEBNRYjpxOtri6R7dg85mEwWKyGhZFwO341xANZ2jYjVw/n20i3KV
0sOlrsRsACNgg8HSkNWQ7hvW1+Y5V9k0bXcTvcwP/BB8fOGrrg8F4fcLnTuse1yAZm6muJabL28w
xJm1lc+GAt4V8iMxF4zcAXCB3q1JNo0ziae8lkFPBRkd0TRfHNvSoO+X/cXLOoC8mgGI8gMXCOwa
VqPgaTnG9uz0G9kJFI0rgNUPJMx7+grBrTEy0+8ACTKsJOOnGzcmhm+si23YDJeYfElwX7NpUIpE
NiwHpI/s0HlulLfAqyd+XTE+F2U/XyXl8B96LVnxx7wDs5TwO9FYD4O1FyrHMZ8Lxze9HFfzi9rM
akuMkVcFneucwRPCk2M92u0tBSMsZaklBTRwSMG3y47ListoYrFHLPvOy9C82YvP8Z82phIkm+42
zpHCcGleSJJaRvqnky3VmzO4Rhez9VzWfMwTfGVKVHlUnNGlv70X12f6RHJwrhZ7TEJN0QUKZjhh
P+tJoQ6Yl/O0lZvnrU+t8Y6XvhqTnTOkHB5cttHiSTETXA7jT2/eoEp2WvSTIEDZg13AX5r8Putq
eYbhsbbdXOBvBP89yq7EJcLFOQzGQWraPZdR1AF8xl/QuiQZYJ5bwNx3BbFlyz4qCDeHa226CiEM
0694KcUIhIhifiPYUOocZxpFWCdEGuqWdAF8tLhax+v3QMvbpF92w/XdVGhFPGcXRaEZ5LEd7m5h
8VU6jP9f0grKtSg1xdVFtUHsy4OG0IPu8/gtuTp8jsobBA+9fe9qN6Pjup03AbkcfuJFuy8RK4cl
pcfaE9q2uM+R45E58d8po93YbDMr2WDJFTD0iakmyUUcjDg5LafxA4zK6cJjf+4X+50lfby9c/8V
f6QQ+mqnoFfmuBSk5qyda8Kk4SyRvV82FYCqDw7q0xM7Njf8PPQq9ihbJSfqq5MrBs8kCRzU3hBc
sjmc28OIzEYfyc9fYvbWGQJo7RITv959Bnx791pT0Kwqn+12yLG/0HzOFQes0j4SzteYJqtzWd8h
yXfwMNpm79PTqVDJLlB6Qb+h8WFflJr736/3HVo+k6Fg5LcLkGbT+mdscGW2W2YPKqvYVr+6/Flx
JNpm7J+huk8huNZI0wXVIr2t6XG6qbjL10BsoM5rZHm0n/0KrPjVcTgFxVJbog0heF1tj9JhI+9g
wafE/3pPzAre5laMl2q0hIRU+9sug9V0ZytCEhwzAulvDnF+qdKPErXlMbncrH2YGQSRvE2u8Kia
PAC1ZzpQNG/of9nybkEvANr1OaSzk9IkQbqNdcayXuQgaG52phrin06K7bfMMGoncWPTWe4ndzqA
mkRIU+oPAp4tgjezUeYqiybzuKgnGAEHzyOio7b979CP2xoJoB1r+Rc0+s7d/LwOH6oX16c/C5Kw
9i0ATcriCrfnG0azzOEJaiQWKfMBLgKTpeAustomzeMEbHwWe4paDc+hgJFHCmKmrxCNRoLZxqYL
PIy9NtJ3yfkunOUmhzhkMQjveL8FTXqDM7As+sRs4bKf4kRBYac96bJdaRUwjkytl6wzFWNEXXUJ
sqTFNY84KDA0DuPPsXxGqHsOK+VBVRy0NeDbqC6WilBxCfNw3Um/PAzxdy6M9U3ey7uMtUwoI7Vm
P+t/gkz0JuaNZAJsIBSaxWiobWGBlIXPSc6ZS+5AlQvkAqU1bTkYn3Go09kM0z6uj5NzmvT23byO
422XxLGtxsU7EWrmpvZJWL32Zm8ClDXPApxNyNaj6ekxiGZTitc3XW1qeB2MLyfpckRaM+yZhz1Y
yLQ4mABLFIWUnDms1j6Axej+2Gq5egyMFvQUCmOVgZ8RAHcxhJzyIkK4WaE6OoWNJM/RPNKo/U89
/JrXjaZIdqv5SGJtordCKzRYrxxnNPm01N5PGnEyvhz05hvmoFMTogPkgTp9VhxQ/JNNkXNrKm4X
EzwEpELSajyRSsrBI6hlSRTI99mcETiWglpVtSuymB1Zo7CIgIFE6NRZ4bJxSXKgpZQ1mEiuqPEr
1SUlEEaHOYr1lBj+j8Oeajuq6bLYoYLzt1Nr9mdJ0753W9yDWNc1AuL5nr3sATb0D6+IacplgD+G
nNM82RfzROjrvDD8qQ4ODbUvMBQAtDJ8mFgaC7/1Gs2eZi64sxtZtguEOdmzIVo8MOqEfOjOhxPR
7BkGJBXbbJNhDWRFqH4G71p/jNLhuz2h+Q/9djwUHBQWfS9m0gJe8E4oSCMInG6yROeahfwpvZMJ
WID55NF+iGBjLLNJoPPmEC/i+Tfu4yB/Js1ppttQQ7t+c9mIHq2/ofYbwHxRslrW8utZcCznZ4np
exslwspb8xjW41ZXfnzSdL/eab2OPl34FkcCUk3XI38go3Dp73jT6zPkWZI2fKKLT7OoNKolNPX2
MxKYl9nePW6A6XqpYeMSp9oGDpnPvvGjydN+wZ8p5b4fWFeWrPb8rYaewK6yjkbARK8GEt8FtK4t
kBpBUS5IjOxCDh6HtVM2fWsbyB67xp1cIgNASGERNo/hCYpJ4Q9RICDsUzUaRCxKu5Ae9b1QABXX
wnqRAru4zeNMGYJUWffy/zxIvoFueZHqBT2D89TIvsbOxWcY4VkFXd20XANhffWGTXBBUL01AO0Z
gxpgJtNn9/MlzcixGXT6LjFBX8KCwPPRvF0kdOoJW9YsCa2LReUBud6h/nSp2LMYMR9EDkjClgHL
e6HR6r30yQN7usEYcMvs7N75uCf9k8vGVh6Yye6ePzFzvMqadtFb6Zq3NOMLplQWItA0UNqxEpYY
kQ2K8ctpDWztpOQPcsDCpZRZUsFsR31huqA=
`protect end_protected
