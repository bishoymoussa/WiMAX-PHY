��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$Rx�y�<��wA�*;�x���@�̦�W�X�fa�M-$u����n~�%���P�$��W��kYَ���P7�?UMfT��q�6�U��k�>����~�\N�(�����X�e���/6U|)�X2pF�]$h���d.���9E��WG��L�X"]�Ad����ľS���8od����e�GT?y	7�������ݵ�^��R�q^]�鍦�����s�ae���h��L��P_���ާ��YЭF���'\��68�b�[����w8�[X��V�F�0͘3����q諵�uW� �h�u\V�?@��_6G�_�*�G���B�絉�f������[�G��U&�����~�F��AׯK1�`c��[<��FY���4I� �#�G��x[X�=�Q1��`��R>(�w����R�O�?����7�,(�H\�#h(W�EH=�������yq��Ѿ��aF����:�U~m<|��.��0=�P/���4ǆ���T(������v���&P�}<�G�"�H�M�k̟|�@ߩ]�H��%7��� 4c�q�ުX`2��r{PBՇ�t�����6Tp�K��
����U��Lbђ
/xЂ����Jz�����\a$�Pn�[��Nn�\EW7�����[@O�h�ϗ6�$o(Qr�q�������S﫳��E.����(�i���n#����~;8�O�}r�w8t���DU�n�`�Ww��@*��y@0w�=;���v�"�����$eV[�ƌ��_	HS�q�K4;n#��H�pd���\�E�P9�&��f[#��r�]�
�����>�O��Z�ݷ���}����JC����Z�~��v��h�dh���k�/�c�ſ(��Nq� ��Z5�6����`&�n�C�65�<�f<���{%K�$
�HzsQjS�������*'l:� �~�M�%���jW���KD�':�I���4����&p���$K�o��*�Kګ�.���%P�/>?�]~�Uy\��Yv*Z��,����l�@b�!-'}Ī���#R�-���48wv�p�-���0!�#�#y��R����-�;%}��?'x�n/c���UK�t4ӣ��7�Z�hk14�rb�氪��ץb;�bT���je\4/k,cz���z�p)�����@�yw���7���F����3�x?�|~�ɤ� �v���o��H~���,?���6��7�j��p��{f>e t_�I�Ō\�̇�b8otRi�h��T��者^u1V�2܅���M�	��� ����q����������6�	�s��y��5���7���ౝPwb�(�;#&R@48e�(Q�d�mC� bÛ��vl7?}q��Q�xv�I	k���1��d�z�+�?T�T@�NH�g�8\D�/��QwX�����-l��tr��V3f�F]�����Nշ�=u�cWоj6>t�����-�@�[z:{�9�<]��>#�n����c	y4�ܯH���mj7�SĪ@1��ހwa���t]yχ%5.�'T�ץ.�g�|BM0]/���b~*����@���(Q��tZ�HZl�q����8�5~�5қY�y�N��s���4|��"E�d���o�)�Pv�No��܋�5�f��q�mPD�6혵�o��2��	��������v��o�lC�"��g�L�񊃤�V��U��D0ŕ"HT��@�jx�ma���y�aIE� $�ͩ= �1Z�/���|E�<�<f�n��+5��/vz��|�L���q��'������0'��p�^ɿ�>�a�,���l��ӻ���o�{��ET�~�:|�]h^�\'r�d�˝N%Q��Z��I����'��۔>����C��
{UVOh�;�~�����b��)���}�XV���W[;��K��)hT=�g�裭��'�����5/��W�����B������"�*R�E��7*`f�Iv�%G�uM�0��b�鴤.=����}��"�9)��O��
��6��H�#�vG-���_���$2��������"�;�,���sn�_c��;�S�+4����y�8����ZG߷�,B���l�.�U|� �����\��|��_���Vã���E�ŜH;�w��"�*>��ZZbV� :��TFZKCՆ�M�uom��P�_V��3�na(�)"3���^�ZbR�lr\Y�-��+?vwad/��[��VB�H��ɗ&��h-�V�5�>�Xc�Q���l	�9b�V�J��t����~�� _^��'f�����\������K(�5�ӣ+å-ì�U�@gU�{�ۃlo \���w�.)࿹-j�j�کHB���%�U`��	��".�_�� L��pF�v��μ5�
�	q8~�}�|̹}�<�[��ĵ�,$�A�N��HtG?�*8��w�M��^���L2�
��. �FZ�&�Ԍ����(��Յ�q��&ศ�Os�,����_9�N?�8�����-x���/u�Ń�8�@�a��N���N���ؼ���x(N��n:�����W�e����h�EҶVA�ch���&Ơz��1�����b�|bGDrE�H��;�Yhӻm��U\�p�������2}>
0�����N7�cl���n��ɾ?�X�T˖1�I6�hV�b��bd�
�	��$r�;�B�����Dx7��IM=��ي~W�RW���$s���v#E��ܢ�Y/��%),C/���T�n�^�A
6o����n?D�1�s���^��*Ptp�Þ���B�B�ޛ>��'~n���*yc\�%s+��0EFY�:�iU�P�쉲��Ղd�ܖ��u˱��������A�`�x�Z�єr�#gb)��#]����S�ti�Z�GR��\�Rv�{�K�j�.��|@�o�U�T��Xk�7���Yżۉ�@�x&���x����c�*����L.)j�]�6}T+�j��R8����*l�t8F#H`�G�t�+�2s��rc�j���'_�W+c_��������a�vx)���lML�o��^݇z7h[�d�b�����rm���LP��"tS)��2EX�,�`ڗ ���Lg�*�02��>�Sɚ���n�C{�_��I��a*}�^OS}�� q�Y�iR�FT�n\�yb��J���Ѓq��T��b���w�U�ÜP�1MJS=�zfk�03Elxj��<��ٚˀ0��V ք� "��r<���}�:s���H�U�c��g�Y��F��&�J�ᾔ�Š:U\�<�j�x�V���K�/�&BP
����;ezV⇏<�X��7�����g�ln�8P�B+�����m�β�� �%TQ�x<�p�n��(L~e�����
���,�5�v�ó�9�p���:6��B�������|,���ڕ�gL�Q��i}y�h�8��m�;݅�[�mt�g �eo���I�]V+`3���7�� c���:\e4w\�MaaP_b����+G���¾ث}	��;��_�D~�W�q�8{m�K�����d�Zb��{ڊMW�0���`�����#6M�~�p�#5i>�=��<$�x���P��4���<9�vN�%�5������)�z�o2�c#O�Yζ���f�K!S��5������=��Mm���Gx_� ����3���h�piKz�˿�P�B��h���GH���6��	`���S�"`��3����V�� U1�{�����?��"cn�-��\=�#b����n0�pp�]9�	$q���ޏ_�=��(>0���^:�]П�B�c��� q)���eCނ�*�I��9ȥ�,Ɲ�����u��#��Y��K�fn���`A�2�������	��Jk�b#� T�9�|��X�Ih��:�q��'�ldz��\@�Ўi}n!o��|�[�NV�h�[-�@�~��l=�p�� �����o�,B2.]�¹3Y(¼����� ��;�%_�nr���ea�c���}h��"# O��32��t����r۴�" �?#\}O�m�H�6��yz��2��F��
�����"�szi���&zg�bZos���.�̛��A HK��n�gv�0�.OhX%�������퉟xzW��}A��tL-�p����4Ɗ��]�Қ� ��PPW�z*GMb�x�aʿ���+	$Zi�H\c���㤠�>��6���R��y^o��-����X�>��#��t��=@�#��?���A��45{ߕWf�{�v"��uU҇�U;b�i���r����H� ��(󂅦8�I�>��wu��&�A��fCT���o�6�م^�:ejƈ��bլ�[6���j-֦�>�J���6�Zg��F od��M��T]֑��p������r="��gI��������.�n������Y?8��e�1т�T��2��'�	��|�ҵ��E��QD�e(/J�l/�0ϼGy��ݚ���HsaW�?4	������T���ٯ�4��g����A��BpH_Ȯ��&�D	�Tڴ� ��2;d׷�zvx,�\��ЖN^����1,�ɨ9��'���Q<s/���~��+6����v�uc9?��MX�d7PQq��y2�w��^��F6KU��c�FȪT��r$���2(	*�b�B�W��H9Ƨ��n�7ћ-���֎g~��QҘ�i��.�Z��6�
h�6��/uw7��\�$�7�����T�Ǡbi�T�:�N��r`�� �{=>���#ӝ��Kwx�5�ܔ��Y/ ax�>JZn�6�A?����_`�����>�0��1�0��u���Yu�}z
���٥c���g��ܬW�P��7�EW:���z�v�7��v�?�(�p�k����]�(~��x��E�b0�p)��$�F�����H�ܔ�(Nhg`��>v����m�}��4?�Ķ��:�����#j��:�.7.�� J<�����8 ��M1�cTJhN�r`O��LҾZ~j���2�J0�zoMo[�2�C����Ӆ���<݊�q�qnN�x^���K���YvC��!䜰���#A��]��O5�Q�_3E(�i�(+��}U�*��	Pxf��KѦTN@����c�N>�6���J�p�����UC�8yiA��Ȼ��<�fw�	tJǅPw�Ki���9]D}��6����s����;������d�Ƽ#��@ht���lA�$��;�񉠔��]u_�>��EIi�W�b)���_����L1�=s��tC���otQ���L�	V�L�,�\�g�j�F���@Я��s\y�z	A޷߇�@�&�С��|��sa|D��<�KKr,�u%�G'P�y{SU�W��9��S�W��Uz�u�'R�P�&n�U-�CA���p[q)�D��YVp2�֖��v>ſ��F �K�c�RAyV;�������`ܕ���	(�O�3��0Md���ɮŔ��ڬ;i��$�Ow��� ���*�$���u8��R=:U�H�����T�;!��0��ý,��a��)r��4��%��Nyp�*��ڽ����{}JQ��x|W�16�J: �JŐ#�9FMP}E��])�*;�a�s��ѷ�v!{�GB	��+���j�Z�+�2�jp��΂�-�a� U��ۃsj����T��t%U�tbnl��9��2�`�ڪéٱ���,$��;Q@���R])f���M�=��4bt��"�j,�#E� ���3�=�~��o�LR�y��)� %�le(�ez����՗qx���� �	z��HV�aM��45���=L����"0�{,p�xrxQz�@C߾���������_�� ފ��W�~�n`}�͹�3_�%gr ~�ܰ-č��DU.+m+��P�"Ê<'��F|�CH�!�d֪�(~�z�8ȿ� ��s�}�O��4�=8�)M���䆴����":,3������jAank�A� T�Vb�z��:�	�&B�����e�_����?A޳2�w���Ⱦ"ߘ>e&!�դ��C�ۡ��O����a�n��ΊY���كF�a�b;6�/Q+���gR}V��b���� uӎj �ԋ�҆����p�=^��Ƃ��PR8O�IW�.!Y�$O�-K�ǒ� �P��~����,&���[{��3XgcP˙2}҃t72��vV��_c%u�8�,t�̆f�
� s�)�c���F3+�pq��A��W��܅��1���,K^�q����xA4�kN-�����ۉ�A.|����=�g҈��+D���[�Uu|'|�As�-���@Z׿�;���-�i�H=�@\��c+6��^��Ǹ�Fg�D�X���D��!��D2�����/.sϯ"�SD%
Mݜ�X�q �]���i�5�:��[WYr�\}@C�F:�:��v	����A�7_�~ʍq � @��f�0����z�b�.���kG��v��[v�"�)���p�ykR|SB!mr�WO^�K�[��5t�i�!��Fa�R"�_f�3��2 :O6��q�W�UY� bXN"hj)���I#U �A*刌W��/�vD��ٽ@'E�T؀ ^%x��-��Ǿ�O���v��oHO?/��?n<_�o�n��Γ�&!�~&PB��}x�M�����-X��y���C��Ȏ�N��*�?F);޻�$[���+i�%���� �S;e[���6�Qno��!?�p��Lz�7F����~/��'XQp�8Ddxr,�|���ix��-���Uߩ�X���ЛZ�3�$�����PFq�WU�3��]Uq�����o��\�B��7�D rgT�7o���F[4�Z�~�Vu_}߿����@�*���d��*f�z�/��&q��MJ���B�*;uؖ�X߆��t�p
KM��K�Ew�qC��[�U���߆ç��<��p��}`���}oc\w�8-aI��4~cQE���`<�i��:�!y��	"�MVٙxK��:��a����{��l��[,e,��c�T�>)E���ruCJ|�%fuHqs%~�Z,��\��%�F�QzO7�
�XU���/�T�e|S�� ��B�wp�����S'�f��" ,ӷ�8�`؏>F���'P9�޲��q>�J��8ujG���	���~Ch&$���5�4$6[���3oh�d�`��Ҙ2W�����}Q���|������ԭԙT]��Rğ�_��19�cj�M0��9돪�5#�ÿ��l��,S+�dQj�ީ�U������sS�5n��,�W'��q.?����% �'i
u�#�7Q5��$���Z�u���g�fmd�o/-75:�B!����LmY�
����G��X,Ȭd
;�^d��L�x��:IUW�,BH�Bͼػ��8%(0�6��P��B�5�:v����O��޾6<���ݮ�р�f~K��1��?xKOy?��V~�d���W_&�"���"p�oI� 1MQ�
�N�UM�ϟv�)����	f)*0O'!�ޢO<�'�?\x�����Gl0���A�;���_�J�?d:����F�9]���`����z.�� ��ªCҰ�P���V�?�����.II1@�.�k�)%^@�O��3��1Tx�
�x'B�$�����>4[���®�j���N7O_t��dal�P�������e�Vh�f�r���^���	X��4$.�J��+���|�S���N������,�����8Xh'��9ߌ2�<O2#��d�mX�9�B���̱V4��C�����Yܜqcu"�9��<�s�����z�{rO�CT����՟����'�F��������0e���\9��VA��%��"�Y�:.��ݪ��O!��?�������~��ih*"�a�A�����E�0ǖ�cA,l�O.��� �����d�)9��S����4��5���G�&2���b4}J#<����v��M��J��>
�U��p�A���v��`�~Kv%��1F6
�`>��ʙ}��n���i���2e��v��	�2}]	�b�`5��)�~��#�p�־�Xq�9E2ϟ��g�y�'|ۚ>B�7 ]sq.3�ҡV�y��d9�yϤe߃<FCS�����e�/��<�^Lﻟ�*��U�����,��G� cj/s�[��O���j�ʮe�+c���{y��Q���Ѐ^��(C�{8���JZ^�t��]��B�n+������aAK�+nl�#@5��Vb���%�5JT�,<�֓�g���l�ɣ�2d�b/1�_/�`q��o+7�ʀ�
���I�r�ycD[�J�b�b�W�����oڰ
�"D�X/F����<���Z�]���ou7�j35��L\"�g]�����2U=I}�x�<|$
e�Ǽ���J�=�pՓT*Nϵ��8b�N�+�B�����.{.-�H=�;�o%�Z:��+�j<���H��I۞�/^�7���s��%����,*l���+(��F�-�Á��CNQ�6�	��,p���OfȰ�
y0�7K�èk2��8�,�[�@U`�>)~s���Нq�H��a`��"������	Xd�M�@������A^���#���ȁM��߹�:MG�yD�X<r�@�O=݊����b*���m=�p5Ş��;2�}��t���3}n��i�/jy6A�>ZI��G�nl�u$��Ǝ �����v�'�V91z�X�'��^a��<F�@(jy9�3�B��{�s��s�T�ó����ę���1�Kr�|�.U�S��M���r��:�M�$�a����M�g��Y6���Y�=�4�.��W�I��M��)��8�M뮜�y��x�4翼B-jIX�з��e�R�#p</�aЪ%j �ҭ^�"��>D��mxV��+�������#y[!~�� ��y�4p���P[
�>/�v܈n��u�:`R�1^!J���V�Bc�'k�b⚱%�F�#�?�l�-���0	E�J�J�\ס�I��G�g��>�����c�{�v�����!g[����C̷v�BC�e��퍊�*�L�>���'v�*$t���#u�p8XN�,S_d��v�*1�v������}�kN(v���~�:�m=g
���=�Mue�hF���'m�O`��XrEbi{;'���"U0`���"��B]BAbʽBt�V��+|R|�Ʈ		��>�ܗf������z�!`��|!�vi�_snXu��D(�`��C�!nkh�[3�ܖBNw�U��Xo���_-s�U�s��0x��R&r���y3����-�K<A�Va�k��+�.�Kn�X�l3�LB�|���:��<����3���">?���0��2�i�K��͕{�}�������a6�Z��KX/�ݼt��%���3-�c�� s�@����b��{�c�g�m��m0T��t�XDm"��g����՘�Yp&����G��E����	�����*�������nː�ǹ^wdZ&c�:�Z����5���I��"�h����T��%�I���gu}�k�SC�Ե��$0������ �%=H�]Б�8� �c���DD�&_mf�&#z�B�]�vL�6AJ��z����B:�H:�q�!��z￶B�T��
#O�T���0O��2ڻ�I�O#��lh3�V�D��)s�`ps�����kͳ��g��zx�ԶlWE�g妹U�>�O4fD��	o�����)�Ū��&ɵ
��d^�F��3|�؀jm��O��h(צ�wT\�2����ǚ�}�S�$�ϯ/{	��^WίZ<�2��aNmX]c��!�E����]���PƇ3����PY�0��~�?�)+W[�̅��@�#�&2dI-��������xOg)���o�A
���0���J(U��dӭ�t�Y^2%��o� /��5�䍉����G�r�����nuVD�Ki�	�a�$�03≿�n{�
٥��r&���2O��b.y�����ߒg.����K���(����sWk˓OS�~E���:�	;T91.؏u�'N��mWs6��!3��Ɔ�jBSz���!:�K*�^�@�#�;7��E��Nz�T7��
1ҐwY�>�Sx!�-�o����h�.h-���v%��̣|�k�U&�S�$��2�w�����`H7��.PA��n���0����^sꢽ׃���ݮ��O%_*1H�JDos1d/�s�5�M����B��N��~�|)�>U��P�{aJ7Q�H���uy��+�p���Yt�g�2>{�|�9�6�XS��T�&A]|�	8�u����3�94�E��(]t��Vu��G�!�e�~a������a����nQ��7K��<#Fk��������mB��Pr�C�� ���D����=�d&ϒ��W�YZ�������kG=ϩ�W��C��OXN�T��ꢐ63�9�<���3��I���L*n� �q����.�]�#�>��@��I��yDR��� C|[�u���@R�n������V�����v�0Z!�n�l+�r"0��5�w/Տ_I��R��k�%`�Zyn�:D�����'F�I�g�#�����G��|�Ts+ਯ�g��F����_j����]�a�G��,������(�r��	sw�7u�*0���#��}o5����%��D��u���0R�RP�*�?:��Ï�)���� �K@�����0����9E=�Օ��2M�ܪٱ0��\yC�.V�*=X�\��F>PP�����Ry ���B(�I��p΍	���3.���W����
�.�u�ؐ.��8��K��D��q��4r`�q��%1����̥@����]tcX��q$(Lud1�%$J+=���˹���P@Ԑ��|ѭ/8~EUs+���z�u�b�Tg@4��8F�}k�_dx3����\�VΊ�$ �U�`����U�+)��ZK��'W8��k�5��Ou�Nr,���/�5��0[�����O�"s&�g�;炽��������TZ�å�kD�"��kJP�d� \J�����N�]|���_W��y7�'�-�N!�ѓn<ѥ�
�)����W�O��
K���l�ܻ3�5Stɥ��W:��^<��o {u����PW�Q�A,�	Z�� 0��
�@���w\�0�y?�����P�r��"oT"g)�! e���
�cd�]�Bq���  �9�ƖV���|	FX�c����Z~�T�c���c���f��Tf^\9�Ha���
�����`S睲�Kb�E�	�*�j	�ly�9�ӛ�@ ��d�rX��Xv��d���`ј������"���g������B,ҩ�Ct��~��b����
@�v4�>�(ޱ<��c�##�v�x�>�����b�b�8��ϳ��\	!��t]y��̾�Ũ�E� �����0���!w�S���]
RE1�Z�[��7��v��Й�D�(_�o��)gg�����}{�c���B=�;�C����:j*-A�]!Q���2�Ż�HyՐ9gm�����:p~�/x����`G� �\�2���=��@f����p#s�a�3~z�`w�s�	j��L��䐂�rB�ľn
�z�/Hf{A|��WW���%4-��(U��%[߾P;$L�3�����s�z�K��h?b~�	t��]%���AӁ\5G��s�t�%-��`V8`�?&h��Qԗ�J{����[9��-Dsп��������$kv!b��Ȁ�X��p�q��YEg����!�j}"7�`����n��`j#����t����P�ƨ�DY��f�O��g��㲬rc�&ˇf=�~�|朹������b+���#�A�h|��pe1��_h�c.1���;��XeH�(;ma�����lp�Dk2bM�IA&�k������f;�Ǯw�/c�|�E��-ۻuP���&������O�T�3:��>���o$3ƾ5C0d����U�Jg���p/Hꮱ���4���/�	^�fS+ QI!|A�&',�]7��"�B�[�%U/	7H�%a�����h~b)�ݍ@{^s2dq��dF�h���������avlK���n�pzN���X�l`᜗��b�ސ�̂K�k@��)�a����0��Ҏ�F��[�{9�j�j�~�����a5ft��c�FE{Y���k���z��Kǥ�8�Xx����{�%��ܷ��ݰ�^��T�/k��z�K��0Ů�YY�Jn�ebԷe���0ۂ�4�+�H����ŷv쾪��`e��~� �LhR�f.��Ȼɕ3��Ry0����H�W*N�w+��ҵ�i�Y�T0�<@�p�- vn�*Ma�����R���y�@�C> �Y����nfM��w������\K����r�ɧ����HG&g�_3%eĉ�g���Or,�!�V�_h�X����!�)�BHZ��޶@�7���g��J�h�d0�����w�+i<��ƿ��K+⓵(e?�n�(#^d�>����}	WNټ�Y���m��ƿr�RԲ��Ϟ�2	MA�U�]��dB��\�c��=��j^�R���O&*��ʆ����%;r�n��;3W�8���r�BEu{��&[���ĐFR_�����
z��A*�蒽�O$��4=�`�l��]��8�X�	Q�EV/��C���RM"�X}%>#��n6������p���-}��;3���g��D�M}��f����I�h`N�-U@3��'yvG��N)�]�wt˫��h��r�����%��A��I�NǬ
>������鵩�Z[�+w.q�S��"�8i��Mr�="�>��\V^��r(�c��Q�ʪ���=��p���0�4k֭чZV#Fƨ�/:�;��d{�&";?}��6v��������!�b�� 	�e\'��$�ub�����n�s��v���8�϶0	�ɜ"��Z<���0��7���5Ɉ�P3M�%����<q!
٪ ��t1@�3��
9�O���96zp��˦�j��'�{9l�T��l����������pY����D:6���J�	 �A%沕;|D�e�crJ���&n�Z��iq�爢 ށ=_t�z�C̯��	�yz$�/(��qP`ȏ�P���