��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$Rx�y�<��wA�*;�x���@�̦�W�X�fa�M-$u����n~�%���P�$��W��kYَ���P7�?UMfT��q�6�U��k�>����~�\N�(�����X�e���/6U|)�X2pF�]$h���d.���9E��WG��L�X"]�Ad����ľS���8od����e�GT?y	7�������ݵ�^��R�q^]�鍦�����s�ae���h��L��P_���ާ��YЭF���'\��68�b�[����w8�[X��V�F�0͘3����q諵�uW� �h�u\V�?@��_6G�_�*�G���B�絉�f������[�G��U&�����~�F��AׯK1�`c��[<��FY���4I� �#�G��x[X�=�Q1��`��R>(�w����R�O�?����7�,(�H\�#h(W�EH=�������yq��Ѿ��aF����:�U~m<|��.��0=�P/���4ǆ���T(���*�X����	 ���6G�^�w��J�!�nܜ;,�苭z2ƎW4᜞����pT�P�Z��[�`�|����#�MR���7H�&D`�b>����!�k�S����l?_gm�7��\u0�>��(��Q�`�QX��
�WΤ�D>i%�"��YhB�OYs�0yhީ�a�F�M���g}����H�`v� ��?���Y��#!S�1� f����fq�V,���jzć��aJ�@� Dbք��BS�-DLy��O v}Wê��o>��rn�.�d'������?DQH��3l��L��;E��@�����A�����T�ѻ�/,uw�2욘ļ�5���p��:O�S����I��ԑ��HXB�l���H{I+����o���Y���C�*.��o5�#/a��t�@�t��ni����DA��)\~�[������+������j27��?VL�[�4�w����D I�*�X7b.�F@�c*�J����&��)�;�j:�0hi�,�`�}JԎi�y��ٍ��w��`H��=p�C�iv;�1U-�~ϿDPy��jQY��,�7�O����)T@�I�uO ���x�k%h�oC	�����5��%]?QH�S���&�w����G�,zo���*����P��NF��tՓ�*[���y�����hb?"�]f�6����S����X�`���$���Aaӡ�.'���8j������9z i�R(g�7b�j�v��s҂ڸ287^7����$������8���.'��r��v���+��-H�v<G~;�饮7�p	��j�09�(JjX0�	�F���i�_U('����N��.��-�LZ�/A��Z6OT���X#��M������ܾq@�u�46��Ej���V�h~��U�����kV��^,�D�����L��p[�I��)��gh�RZ��R���4f=���}�c�?l(� ���j�����dk�N2\�1�`� 9>�m���*�s�}��ˇY�-:��9��@
r��Bh]��I����}�o�HU=F��@�5ұH�r-���^�~��K'`�R�,�z[Gw�&�e�����qM�vCԉ.�a���w�{�^;۩b�v� ��� ��'�pR����"<L�r����%s��%���ƞkI�ԝƷ�IN�KR�~YlV߀��{�7U�Þ�ܰƈ���|�E����A�U�왑oA/2Dh�L1�j��k&c�9"�-���,�70Y�C�O97��Hu(=~@�Y�m�4R�"�Q1�K^sh��<gXp�S9!y�L0�|��w���TFkRv��`0�g,�:�[{EH�pqhk����l�~���� �-u��k0`����>�d��Oh������_eN�L��	O�����Vo<ЯȍS���禗dTa��?f�" x��S7\x���3&M(-���WֲWǴ��O5���E������ʽ,3V3Q�"F�)����x��PHeP����9b�f�Sq�Ǝ�5~Urg4�c�!�0g4@[���2R9���Y�L�OJxkj4��yJ�X�_]7*��:�/�s��Q����|������� /�#?Пݿ��j��ޱ��b�/��/sCv�P�����˦W�Sͼ�K��2:ɓ����TK������KMǝ�8Ѱ��c���@��	|�	@CJ�5
���AS�@%g�U��Jj0K5ĆX8�Hxs�A�X����Bk/a�u,�B�г���%��cd����S��,�ip{L�C�����S�,�۠��Z���x��M���4M��X�4�&�B<�pI���Ԣ#��Wގ����mX��I�3�$QI$`M��V�U,�ͬ1N�Z�Fj��l85!ٽ[��Q+��3�m�d.P@�־�\H������/V˳`A��� ��>px��-0��6IA�Y)�1!�͸@���B]t0���1RQ�@���ӖǄ����7*�W/w!�GK�Y>b�ut�J"���㤲������f�&~�M1���=f��I�x<Oδ��4R�G�9��(U�"?	 �+'������������Lt*�X����X[O�����Orrt�s��Oae$Z.�3���Z�+TQ|nm��yaގ�1��h\�գ_#ۖiwq�U���A٭�̠wܸ@{��̕���[n�V'
��r���&����V�������W�%�aB�?�p.�P�-�W8u+�����w�`�����B�n�!q {l��e9]jt�X�'I(�,o	�\���D@n;�y��\�a��F_�Zl�O��؊�ß�,��)E�(X�`��� ��.yW��[')X4>����ȏ$��#�ჲ
">ɍ��=�}J���8�h}z$�&`x=O�����Hm��)q�է�I�t������o��pX&��5���g�I}ˠ��`
��_=N	�<�j��*�\^���YĂ��?��2p���u�܅��S~`�$��"G�S^�=I_~�B�{%����	�z	�`�g��/�C�t|		��$�i�� e .`��4DW��T�JS����������]�sQ:O%u�|pv��y b)W�*�HZ81���:�7h=HR�M�����s��Ɯ��L����G���=��#ݒ���dT��k��eT�b��Y�*v���dy*�+����߼��ܨd�r"��ҝ�����De)�|WU0��w��jZX�z�o�d����g�	�	`�N	Ae|zZ1�� $ 
�� N�.b{��.� �o\��w�bx���Y&���Hc5]�gn�C�c*���V���X����<�L��Ү��#p�b��L	{���N3�DJ9��1��r�?�`~I���X�=�y��e��W��Q3���ۇ�x����ػ,�TN\���o�~�\s��\D�*��F��I�2�G�Y��
�%^���.�Ql[
�+��"��0�".���7_�����b�,��L��6w��V�Ÿ�J@���B {]A�-��o�������Q�=ϗ�������x�Wͳ�[�w��$�Nu>���YuP'�;g0����^O�	�h`�Y%��+�����c���5�:�ON�C_dSs9�c,�fA��{� ޜ�Djc8☎9���&���+p��� �#�?���7i�����4�!���^&L�G�$E*��K���Oez���rgv�ݺ��/G���!kM���dVX M����Qg�5M!���E���Bצ\YQC𠓅�e�$�����y��G�Z$��e#˛�o�Ţ�[��=KV|���&+�ҋ�J;��cm�'�;��iD%f���"c��X�v���n0j�ʃ�����ñ3����}O�.���e�&v֊:�0���c�����XU�y��{Ӥ=�Lc�W�f!b/x���B�ɩ���x:w-ErvS��5jx�v��-}
��@>�?,�Q!q�b��~��B���f���H�ԈsBO��z���dV�U��o�c�C��@��p5&��Ϳ��9����ǔ�߫�}&+)��f�+x�$NL�B��ZO�~*��Xj?r�`��/GR��/i����Eb,��P �Y�_~<��{��|## ���|H:gӐ���A^*��o,���F%L"���@`�p�^��<X��K�Xp"�z&5¡��l�ֶ�
ٱ-��-�R]�!1Q���y����0wO������8�>�� ۤI#MG	��A^P�G�b�nU�� ?󠏳����:G����*������V�U8�����8�0I2%5g�:t��3�L���l|._�[�ͮ��(���W���o����`Vw0<�i;��X�=�{[[<��H8����Љ'd��dB���GS�(�����0]����0M����R�T���&(��e�ѡD��7�]���C�ܩ
�^ȸГ�/;	X#�����:��2����J�<E0�p�=��Vw`�-�4��<%�aIgzye��b	4���Vm�&��ӌRk�k���=S��B(0c���n����>&L��d��%���9����Ȳ�\��c��q�GT�ц,x��$��vSxA\��cHj�07��H
�=Ŷ3�d�P��4��x~�t¯��Y0
����](��DD�~b�e� :�ⶦU<�9�nQ�U.�6L�����W�$<n0b4ސ��ߔB�"
�IH=?6԰�]�}n�������-6.a��,�� �m1剷[����,@H�?#�pcau%��*�hSA��Q��,P�
e����%��-�VN�luUO�h��Jb����;������~��%�Y�a�c��"��W����,�\%�aY!k%�
E�r��Q�GR�W�O�@�x���$Y�'��YE�S�(%������F�h���/V����B|�=�c.���H��xh-di����������#�Bv���̱�==�g�G5���-�zЮ	$;QJ2���-�i����c,+<4N�O� ���u:�V��99�&����;�V��LUJa��,�M2����Y�Uxw��s9 ��$k������{-�a���L�~�ꐲ�?c��˙��v�eJ,Λ��� V�J�4����� {~�'�n�pm�:��L���A�o�|�飄}K�7��?c�SaD{f�I��TR �T)�����c�NCF|��uu�[��Y�SJ;��tF�8��
�ji-%P���@�[:�J�	6q���T�$�6	��dJ�{儂J�uTIU\W���C��7�2���6- 볮6���F��a�6��]]��	ħ�;X�	9�m��8
���P�Ἷ`�e�iVD�K>�F��z���5���P9+�|=��,��2o�9P�@���Fm�Ͱ�0&e���
bN�}�B� c$�urd9#��Ubk�	Jy)Sd�h龞�5U�Р�Qcz����Ǆ�ѩ���ݽ�,0���F��B���#�A�T�Ok_t��YfxC�%�$�O���iUK�#����0�Z7=��&`�=�X�kTF��)�z��w�!
� /�F��ف�}���I󂑳�+��6�7���C7�I*t��Sa�&�f�9���>�#ǃ��f����_����y���v�N��4�$�X�@g���McY����΅<wȨh:�l�Y.W���S.lBf9A|���Bp53{�QzfN�U_����a�)�T��>Ć4)�v���x�Px@4_\�ex�A��ʻ���!6�HKm�43��|���2����zM�J1�U�����<�Y��t�Y�Ĵ�A�ɡ�ޞu�q�y�a�f�ċM��G�U(�e��A$&`��R�.^NUc��S ��tZ3F�%�Ģ�uM|������� 5,�0�բk̐��n�଎��H=�����ݱ��"�n�Iؔ�K����)���'�K:�gB6<�=!��1�W���i�0���j�`�eyq�)~��Z�P)��ү��������bb�µә/mX߹c �@;.�U��W�2S�a�fa#��:~�6o����g�?��8�Z�U���A?fw#L��ҡ.�e��Km�?R؀�S��)�0�N��8$р9�}K����s/�"v�:��2ǫ���U�� ����D�Q_�����Y���Ojb��Lf$0ݻ/�	Ǘ<8��"�&�u�4��~�"���r>!��]eAj�l�*D��$���0=��`�	5z_�b$	��2e��T� Q>e-f�n6��˃�U�b��By��hҫ�I}[,CF �����	�P��Q Us�W��<��A^��c�b�k_Q$��T�P2C>J�ŷ�����Q�T[Rw [_�=������)4X�~�o4�N�k�q�vT��P���}(��Ā~
�:wz����^5���wLf'mUL�2_�;�<od�/ʽ�ьjڥ;⣀]/�8��1���EgU�,[��'���X�o#��s!\>��|��o>��D��m
C���_}eA�i�H��?+u��������c�jԯ�F_�%d��(<�R� ��Xb�Hv+�N�W	;أ��$�P/@�Aa�6:b�D�:��Un�k2��_U�/������GX?��E)���TB2[cyʂ��Z��R裀�Q�{�ɋ�4^��L[}\���B�!D:E�.��dC��V)(nFJ��5��b���YNf���OV�3 �e<0�6�4�r���r6SK�"��@�ݛ/����K����*k��D�K@�kz�nx�9b��6n�޳�l�;.ɇl��n�'X��7�f��e�W���`�"O���;��q&�9CPծ+9z&rC�r IzԘa�v�D�����	�U;�Jі8��b�w�bJiѝx�g��^��E
��\��Ѯ_si
x��A��z�"^��μ����_��)Z�]�����q�K��+�"��4�3&����LF�������l3�@�������}�`I��u���iX��1��b�[�E/K�;L�ſTM����Ҩ��TЎbT r��)CQ�N:R�M��,���#V+��7Y!,�~�'���)��UT����V���|EJkF����r,����ަ��F�˧�d;�|�߼!CV�������S6G�<c��c���vǘ�Y���^� �'���'q�������8P��O_!�E@Cq���=]���"��,]�]��Q�f�Ԍy�)P�8��o3��~9�`l���k\��m*U�W����uW� pO�[2�p,o�2*��$w�26�j��n��XL����F������;atuwB�GU~���C�7��)p����UP%�Ϟ��/*3EN�Թ�(��{� �T����s$�zƳ����#�:�9��F)��G�-;  ��w���*�7f� 9�ISa[���\��]wd08a��i-����\]�<��E��w  �;!/�x�V��q)��|��`Kr�1M�pv*�@�ܠw��Ea�e��w���ԕd�@ٗeG�s�)u�Qӏ2�=��{v�>kYm,]�}�Y!_��~|_�����	�q��^ � ���%Iy�7=��0J�����r���^o��,��������k��}5cV�kbao�{X
;`�"c��4�NĔM)ױ�n�����g=8�n<���y;��-BP�&2h�	�m�^1�ި��n��z2 u1�	GKFj�_�m�m��l����O}���AM��q۞���͏��v���@B�D��s�G.@e���s�_��
�J�3�̂K�DC�b� ��-��k�&���ԋu!��)I-4t���;5U�\=n�)Y�f�}�����*��p�?,��xM��X��M��2�����G���u a<Ӓ����|"mB����k�쭯u����Y���?�:��U�D|�ur �?���D�v=}�,��;u�Yl�-Gc���O2�U��C�"7.0aꪷ��q1ҧ5.�*�h'�NRJ��3K:w9�f�b�T��걅*|�T���j�d�q�y}�VD)��n����.�fZ�7�U��8�((��E��8u�n����_�ݝ�|Eu[�c������{Uԝ;!7o�g���;X���5;u��dk��$~,/e)��8Ǒ")���)�v#(��i[ʾ�[���NĨ��h��꣕+5�Ԉ��<���6}z}/��a�MYrAP�6��k�^�!"1�qu�ژ
U�$�Xx���ć���!��l��C��5���v�^��������m��ԙ8�����hkŊ˶�kVJRJ\P�d>[2b�8s%P��un��`
�ɓk�^���~ڇi':�J�@�yr�]Rp]]��f��(�aʚ�Ζ�}@[��8KmMck��.�Nr��&��