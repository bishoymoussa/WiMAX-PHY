-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
AA2TsODRhkXxZq3vIpnim2eihgDHfQlQfuf1z2ahfc7FlgQcLq+vlAy8pycmFXXocq0jrtoKlT9/
OSznExXrgFSn2589YBoDaPdKD3jU8PzEs/hVLuMxJZ9BYpHLIFAC2Avq6lO/Qmpsgx8XAZW+DaFQ
qQWYFegDzzwBHfolzP+YA/F7Q260aP//RT56AGgXSsg5X46mGT8mes7XBv+G7s5yHoHFg1SlXMIh
cJOmCpdxsJu/0RldsmkpbFjsva05wRRkUghRbjP6LFhNDYcGFv4Lbbr17dgu8PrQdm9Shxy22RsB
2kjY1Z9WOsn7K8ue3RpEcuixAIK8L3UDk0nzsA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 72832)
`protect data_block
10l9XYSncneWHSef3xT1GYpEKdW1dBJjgGRGhwzddkWS3/kXPJ26RKWIErFX+YFMMEvXEu9KyXP1
dRtdiO6RSFLLmtd/JZYFkqcFFRhrlmYxawoUbTzX46HGv62LCWrsqQgmlKtrxntSTBODcbjCjkNb
M5E1w/UUT7DIdXBcck0qEYC2istSflSivySSI4FyNgw6HruKEHkM8kW6SyQd42+ZXZDEb4ZnTYzV
y4RMyLC9WGum8ureTfmOPz74r4YspMwX7CYmYo4QYvCz9yp+IbALd0xFW/8WAp8de4F5tMjSvcPk
lwPvIo61hq2tQ5smILmK0hUDRRkzIQTOIHJ3TZCp0d2xjvC8ZH04mnx4ztWPHLqNC1llzxMutPvM
C7F+KUyRDoY3PisNDjAQVaECmTV1p1J/pNbN+p9C2KYTYp+8VSW8qGw2EGU1vOdVDcFh0/YZFMr6
+aezTWn9O9g1FRS7yvEVoeQKeCumtouxMK3QIeukiQZhK2eQH0bMRAxitQEHpMX63lXSMP0Quesi
lOwiHZhvxdV9XMfLCadxbtIwa68sSHOWeUU4KnYtrf0jaOOypJZly9gt4VpXu9V+YlZyMKrAGsye
ATh8a4HGuarn1tijBw0L9HcdC5QhSwXrEmC5QRq5bZatOkf6JDao3quvcom8NgAk+XyCDwFUlH1S
HzaHj6lXLxTGnk17cyFXhL9wAmUySjOU5PVGGgV4TXX9LKVd6g9XEnBtX6zpo0vPSdJOxKDzpJ3o
lzkPbBYGwiBLBtgd8EE724CysP+R3SnGSchqaVJEJK/wOC2NO2bHOftTmp60vefRWPwo8P8Ni2aE
WHzj5m7aOAXPvgSkIUAfuMj0Nszwi8N0iHrEDvjL9pvnQQMnCTONX/fNKr1L5xTy+oQyNKV4xHf5
GQV+9tJwW+YZMEdJuAWd47LY1/aXrkiGy7ll3k+tIe/nC1PimYdszdA9IDEm9/9KiGfDUCaDWbxO
PQ4jo7KaDMjHyMtEgztz4prWEF8tQwqGOg2hbk4dtfxXhrNUbpzFr7IVpDcF0yGm6K/u2PRXV9zd
0OQdx3QLeIZjyv3Dpo19ST0Kya0DCw5+ZjOmkorQ15zkz/cxro7uMKmtEs/2lmk0Ez8+t5NXvDi2
9m+D5YYiwqJb4wLu7LRQ+ilmF1lXnNSBenUFZu201wljsmG6tlI7XSfHrFynysUVIEi4nQe5pG7m
6zUgBv0PEnvrYVLWFCE2ecLOpMECK/UhG5ADNuVGywxOTvAar+Q5usk3UKH96AeKetbykor338uv
m/RuVQpJZTa7FbxBP4kZ/vNO697bFWDT7B1+WnWrYbRJBmzdYfPqj+JvlDEgcpe0xJVpK7i0aio6
KjJD9FTyCxu8TpEfJlaMf2Gs7bapuobuZC1ZQpTezSvH5K6e2PUJY2wV21MJNr03LjrnjxHPWqHO
hwHRfLYaUCBvj9d9xytc3LvllAXvCnTz7IRmMfc/UhuIgkmwv1klzRST1cVDGlBLjE7pQvX1RNZk
5fAZ1Ca3rxlnIAq4/3QPqtmjZKtRr87LhKkLnSFqAyTqoXwc9pLsFp6NfLnQgi9zIRg88DIH2PIl
7j38m7oR1eR+wVU/ITgUP1HAdNt+9rM4Ujc0ZoNEKrkc2TckD0Gn/BqoGuzIKUNIAMFxPNdbdGcl
UICruQU0kY6ehXIMlOOtKzrK8OLiWyikYFQQNeAtMA2jiXinn1ai1RRGOM2TKY1bndaBpZJ15i3p
vHyx1JCYZRsydPxe6gusc1eQ+XnQTHFTdaXOk9YMPN0KapoT4LNof1iLlU9fF/MWxm6qaaDuq5VZ
T+/UT9CpHJLb24FIPjLw3FqP2pDiHbIJL97miUf6T/qXhtJV0PYKm1K+nL7wsUBa+lNxtxPM6VwD
muLFo9sDsRVf97bRFdDy3ZHKm0crHYrmOrVhPCxJcDfuIJ8inOrs78MGF6poWFvYJg55/pgsYCwp
15nyKG0xet3sCK7/WFEaKX1e9xvrNeSAKez/qp1371CI5gzPoDLCIOBuCZLrOL+HkCb4ZGZnetH0
8v1J93UevfrC3EJW+S0kH/reZr+y3642dspN15Sekj6nCoxGj1JJBqDqhyU5RirqJvQ4VFtaPHMi
wEVyZn4mODrlRtWgJCE/qItFrKYe7eSPc+H19gaclMvsd3U14z6YuCYvva+oYfGmgdy4ysrloAcJ
panGDyTXMpohq9bv6R0ezz42ufqbXvuR4zs5JFrBLTw8jLl293n8jgCVkWa6usimfGaOHTnpWQ6X
3wfk12xVPsHLE3+ZCyJ5bA76qQss8HC5omXzDxte1x/7/H+/9zCagKQpkrO09hcKFPlmfOiQmr5p
GK394tPty0HWMvcFwAgjZ/5BwvclXllEJZY4rFOcWDwPSppGcr/BAQXFtOWNA3cqB2uvs7SBgzPD
Qfx6iiCWh+FTZaFN8/gbPLzsTXUyiPFNKLUGDp7kMqmK7EgLTZN395QqRz/8FFoxqoM8m/9AV3j8
4reFiGb+SY/Bu8aawAqaE1a12J+1ise75uM1VXHlJdLi59ULJN/9XAxDvGam/9cbbcNjpMYOw7b+
CXD+gbiHwyDFPBFezgIdCUO9fz7s3L8zTPb71R+jRCREkV+QJdvVXDwpEJq8ujymMUQ0rEHlb3Nm
Cc5I/COdru05KmeV6EaL2sKFIkXmHg5+DxaF1i7Ix93kg8wQBWjbFrQgIqKD7TWhrbloOTIFkf4O
2oy28T0CaU1Zk4WWWZlDYKLBdgldgeMYm7mkRUlUSSqUNuUGrx2STsFuwwZAiguEsBBZDSUjI+ML
P8oBpmAu2cNBQJBCFPzZxebuMsIaBtXIkKWoFiwUAl3A+eUyKYLJuRUizhUGAljPJLDMoC6tEXra
1fqYMPHV17qfpojrII0tLOftcaJsPAKziwXGO1kxMd4YjjCvWReUmP+KIwQ4MBvz1g8YUe6Cj3cs
rIqPjKZHUq1MRxa1sN99qVsvwRa2OqaGNoly/5m5edFL2ufeMjfJojYRg8Lakd9vXR9fnKsSy4Vo
tM1XZTUoqFEy2mgkhL/jmxOMsE+zNwinTnSibsITSZ87+mr15dLxNxZtyzzHkVADDVf2xx9/6DVB
g/CnVzKN1luCVzCIy73kpXSotHWrgp2lITU7CQTUG6j8Hz+e62wxmgBeV/4Bq2QIBj8i6R102eFd
bC8joikp795hk7k7i4lDfCDCPfhCh7ELpmeTDzUl9vjWpFBbtEc2/eEK86iKeCt7mjjaA06+sK2r
hsC4p/asLtzJoGTX7BzOXZMoGUhCr0cZq3yJZhFgg0ksiEMRiWLho2fgVIJp+0rKXVYE0AOlD2cO
IBGd93dFS4iGCLwZzAr0BZYepjoXqyJ9zGdGivjTp84h87VFDoybLB3TvavZnsFmAi52riZ99/vX
yo14AKF6cpIBsRx5ijwUB358cfq6uGCCmtvI3YtlekNNe/v0xJRa1AJc/PqroSgEf1ugfZsglfQW
mf8hi1IYEs5h/EoJ9pVWnVZlRNZudk7bixST6dHELrt517BmWvxE/YNzefpzfe8A48SYvC/IC+Yj
/rM2+RciH1EEwHKnbR1sD6xCtV38pEJYD1Ynn/Z+gJOSe+vGv01f3XieP9tlZv01X3Fa/ea5brSv
VOG24us1eS6eUtUHj/eLxhFr97rRuMmuysibQtPybZTo9/WBgAwa8P9JGxmf7IBEMaD4fW1T+DC9
mmlqwZZkrg6lTCWVAjGWxDsPDeNTrYdqzJDjw95RIR1Imc3PjnnJ3+P5QeAk9iG7jA6in7oPrxPx
Q96qLSRCU7o0E36EBBBG6Y7OMrwigiUMpmL8FJd65fB6Fzdg+6s6u13vcsYI1BbwzP6fDGdK5/BU
DGENGvcqdISmZq4u5/rjlyzjUuu3ip5LO/N59NLT5IItrNZMKyojxOsihverctB0g9zj6W43zydf
VmhcFM/6uF/6nqerzcleWKOYZiq8nXM4wHJ7F7uEOz3N9an8IhFa+75fEfqDFBYhXNmymT74HNYr
nlP9EvMyJfE/oPpEZWqdNgxs6chZJsI7GfnC9ixvRPPxhOkYo58C+pDIV3JZtBaUHRudAEBzPcVl
BB5SVPp6zuRNlVLQ/Xg078WASBL6YR55dbVaEFUV59PhmxgXEoiuv1Nasy5xZD4iVqlRdanhL71J
RDGNw7snVKp+YMW8wjTuOnXuyozjxMGTG9u3zMNgnxqnXvqgcbren1hAOTzC31BpVQyUHwNz1xxv
y5udYMqIma+YMsV3I+C+SotWQkKeV9Ia9ygMbQXVMpSsYnDxZFf2sMqFnplZRlmv2W2/4xQjNBTz
ZyQqX4/Z+L0MQ4Mxx4DTR9z7c+jBRbF8EvA01tq0qf5uiWWVzQwxn2UCtef1UDw6ns8NQhBo9ghu
aa+DFhRnb3MNivU/562LeM9lU4+pOWbUAGubo8HPuHZQkkFl99MwHcQzNTtFonaCCscUwD7d95EK
+kmgeipIuKTdSJnhxV3ZFZo+gnhJqAUqcxBE3D50yVui9g+vse6bg0kszA+PP86Gad5tJWh7JsQ2
r0eibB7yse4niXrCb9ZdOlgg4qjOJ9+ZDiPUGco2kA0pv5aq7bgTk8wb2+k+Wx98PYpECSGaIuqP
4iiXk1FsyYQSUqeqxL/i93W/pV1m3wjSlPqgAIFFd7R9Mbs5GWFuhLelk7/cV6X3RwAJgpuL2Pie
DRcfRg9GlLaqCb18Z7BGAEuSyW40zBPO5FuEXzXyJ9aS4DiSFgLbsN69wUrl4YFG0Cn11wsPiDTc
JhAIdT1wFL8yTkGo1sjTTNvwY2LIV1ktDz2pgue2d31iPymeu+kWSH8qU0ym6VCVYEgSB3Aqu4gQ
Q1M9aZ12iGkF8XAu6JzveP02++u9ehWujAcx3YZMCtzNUX7oem+vVsCiXZcccaGvo6M0aSMQcvR/
p+o/PxsyPyNyK8+FG5knWDLNyQdrqYyuzsXbaCK3NDOmGy9CBFWt+1btQ8miNv98WMYcUtPT3tX5
/Q+j2/ECFxgw4BM62qPHjQ9L53tXsvJ9DWKmHZtd22Ut3MXb1GoZ2rG9ScqNOBqk3VR0MTn7umLF
m+Wi61TjyUHiq2JIXh4SCQj06BykyEojP+gKa0tn2FzWToadKRkGhMN6yMbwQ+wAny1hgNQql90j
rsWUcaMSl2+1lKSNZV0S8z3jiW7Pgib7MhHWvMSg6b5Q0MJp32d5ji+n0aamhRYEwbXYVmnSXmKY
Y4Zj9XY7qn8oqWo5+4L+nNhmst82OtFcIvvlYRtEJjlGxvetvebPYWV5Z14Vv082/EA2p20Hho2S
BgE5AWqQdeIcTl4CvEQPIIkKfU8amlsYEd2gsz0lHiZ1YDr4dvAFZllowmP35PIO9T6UWMLb6w2W
7/hvo+MlyvqE9mszp18UXDxRfMV+pLwIgPwfvovTrg2FYCYUW+7ovK5cjf8jrUFsssBeqB67XIO4
GCJ3+DP87vJRYjnsF0Z6kZlVTwrKriyVc5qz+9Ktz33S5fGYGFM0NyrcBdDNk+GOt0tuHYrXLGCd
e+wNKqKGQjdJwKsYtXvag2ifLWEUMPCbycrwmFHTYSOKrA6AqGSpg/coclmbrlo9lF4k7sXf5gUq
IO2bvvEA8Iy/X66REZG7Q1zOGG7F9Yj0qVoGU0olpLc20JCfRejCjoClmP4uveWxCJs70kdGqEdE
TDT3MHgDOqaui02NiwgYqcPes4O3lhZOU22fGyrUi1gVIZmC1Z4vPvKQoPFY2O8FAaMB5PEwx5gh
tK/pV5vgmr4FVWEWdp/q62TLW5SjrMA5d1QnI2Monxuc72/mG7PWx7e7lZRHjui2gcajsVcUGc3k
pKN6EHy/GGAzxg0kmbIPdAVKDW4pVzVW1JWWYlIwsXlJZp5JgouwEWqC8zgZRmL5NhRNha2sTXWx
PtH3AFFXHbH7mdOyeJkcsuyEqz28MuiLWmzUcBR+HUYiQsE9NwrAzMMkYC9jNeWpwkCLB9GRTcMd
6gwMa8+68rFaa2KNB2IqWqidbRMU+YM6y0NB4yDudaawKkZqxK82/gy6xeMyrF6TmvT1c1aO/vkP
CeH1BpPzvcQNFp6OBw3LtOrRbGFvJfCv0WS5bJTwKp4rk9DaN8LJNO7+G8p0T5fnXLiCcG/d5gXd
cG/MsBKD/7aVhITEptPRhVxH8IWfD5ZN52Dpjx83nMkdW7YWwX/mSThrpMsJqiBYjJltvyEW4cpw
yTKrCIl3e9HkWGNEhwkMyNkm9V2Q8v4UtRu38ITdumlhZVPdMieykIvpQrhyKLtBiibOxeE9miZT
oI1gFkDRlEgw9fAAHsbx73/hg0hx+0pb0R9tvtH5ckETTdk6x0FVxDGRgiSD4MWqhC6BIF/Y3+HP
IExbSHQangTp2Hy7XIhn1q6uZkmxnP4qLpp9ydmhjOKvbw78N8b9EyeSr3iqtKazwrJXqOjb5a9R
hN+Q34m1So3dEZpDdzlf2Fi0ZuO63YOcon6XAVcn55FStt/mlOVIHl9XhMgEFhQd3tjfX0QV89DL
f6td7qx6ERs0pQxH5BBeWPjtMGmsnybpz+DMRZmDPxWSdiQ+r+hNDbYHHqVNwa40MtUk6Eetz7SL
8QsMUfrqLuVls41t1dhLzwKLpcSDd78B9vMYeEnyNPc05JLfO5mTwMrqX2BW8Vz5EtSwqx8mo9jf
RtmjR7lB18hYRtM7Q53Nlh0R/IoWESUITv1S6HltSSU3928IO9C2fn2tYUK8qUkGNExw/YnE0/yp
cSC3lFVZ+62Cs6qSopMiSGTvKU6ZidS2v5xXLp9nvXwB8wraSMZy+Uk1dDBTZc6Dvp/6Oyf2z76b
qFDm1ClVXX1+4fjSSbmJ9Up6urAFnWaOz0lwKAdXXYk7TI9dj0PI1NI3aGWpAZ78Cd8QNk0jqj0t
uZocvgw4q6PzCYl5XqzmiufNyxUCw5eCln5ow6yKEe2WZiovPCjcF2HD+e4r5sYkqLXJchcrqrmY
2hxgQj9eXLYp5ViyUt3DAy+ciWQkhEoCP5Ivl9r4pouPv/FdFN2WjN6qHLfCGDWvRgPIL4tIorU4
KZufxdQHXOK0GsqrWrHKCDWPQ5QNtFC3gxfD/utpXJr6LKP+ItNTlaL9qx2BkHcxgf5NgTLG0vNO
EEsLK73c4Q3MRNMuBvbLZ9uq9GGyBGIV0VPFcKW2TR08PSttOZZg7IGOUHurHDH3+MBRyLHbn4WH
NRkPza3tBfIyj6L0djsEjAhg6ba1hebscwkS/FE5WelX8UDK4HAvAaTskok6Lh+ZxczmKJByMVKG
uEIPg5rXvMxgvq0NmpVBzMcawHm2/8C7GBL1IMdiigqv2xq5LimevNzYET+rTTJT2RWVo+4cioS2
nnehcGneTNx7FoxZFmlfHcNmOa46jEbYPuSXx5EH4UTyD9pogHVgnYN+tZoGZxMT6bVUlQTjBLkZ
1HXkTpX0HtRwVc/u4IYGc6p/h3D8coZtyjxTo6slxaKRbbdk9XCuF+beJBXeRLMUO0c96nBMQ2XT
jQN+wfdltAOd+UJen3+r/w4rjo4kulMR2IFo82vE/ul0WQgtUYosmUB2p+Jq5w1OObzgoYDX0Le4
349VbKocczoH9F2ry1M4CNMQLI+a4xmSotSRUzx9NybbHpLjq1M1Nngjxvf5q1cvqd5TTtnsADY2
Ycwe75NHGxDF1R03jjmVZTGhSZJNCqoqA+4lb8dGrYKInzyj31uZp2npQcvTpeno+KHHCGFoWAJI
LocQn0w9KqBC7U6ULRsg8SIkLhbUoF1JdyxFNUoxkfWGDmOoNtlb0/S3lBC8l23xKu5UlDZuv2VO
gQnLaZ31Z0Hz3WQaetq0LBlJ9UdW5JViAxgu5cPxfxQ7qBwvTEuB+hpx/1u9ZcwbVrM9BLS+rtzS
m0pHLb+14AcBA3oP6K7ari8NWECsC0sR4sNRasMIj840+AOvvg7QRtWWFIKwt0mEaX6ehGM4vbYj
et2qfGZ2rIyTKj+A5PPmDuRXCuhl6gtuNg/dj4GGipb953Po0FqeTggcRN9TDMnFtMlOqhqRh7SV
hzQpTTLEqwlrKPOgY+gdTpltocW8L+gCcG6XJePSL1mIvXrFco5709xdNZ9GBSGdr4K72ovOa8ua
xRL/QBqwuLY16w3EAOJkHTrILzYih222GW04V+Qe3cER1hn0sdbjyUXjG5u+TMFlV9F9rDTPWT6t
ms/iV1W8FCWqyY4JYbC9J0UWHone3Rx3b1t1fVszm+u/94F8e7vqOPe6VKkhCq3TlId/WnFPWwlu
8MH7KGBWqmqrBY0z582KkcIUtXXe4Xz0aV0A40irn+DNlsn0LQu7J13YWh1pN2EPHMQPI9xvUMT2
dQtSeJaOYIPd5MNETsg2BLSbdgjR9Ec9Twnoya3RmWqqyZWcy2UsDvdslXGYtHTwp6VRqWsCn5ah
YWN7nFj1xrc8kr4UPLQeDq7vGhCqyy1edYO+Jco+85hELpcztOluiA3xsRZycoxBfOLJjjgvrZ57
zMU45pmUuYnqduLdsg3nPYZAKqh1BG3t+AvzbdMRwOYLsacQNKaZpi1J6VjE5/nA7SCAmaZE+NwT
I8IYN0RZDvgelV4AcD2iv0AJ0Te6pb5SKsFei65/e6NV5FGCvMktREioj+xk435umPNWQdfwK+Is
Clp5bo7CPNV1spLT9fnyOLOQV5wjOqqcTf2Hx3f4rm/iLmvu69ln9aRNKoqqu+8b7bmq8jfQjXuk
5JlSRnJ6aGavc22kNflAltXJ1v4+QD90yFQINoFrRabou681JTtb+n5dVfSlmAmoGxr3t0SNdqlj
SAxg/xBkUYjI8J25sKhq3HX5m2UYr4mlIumN93yYnt0OE/VcFewX8h1UMJyqalHRNpxHnkzZ2w65
l9gJRiOB0Ronxxea/wHgOHJIT8WfloyzgIcZqpVIGIDMK2lX3VKj5KQyePFYX/+xKus5BUwbcmpX
GQDqEla0A9Pwja8Kg0KX7zA5QXYJ8686o5wJ6HXvsQkcCYGjppoqmYPL1lSJIfVjXrI0gDSGkdQ5
3fBY+TPhsLbfBajbMA6lqFssRNuSgGrI1g4Nw2xMhwv9xOYX4z6e/A3xBixmYovdxbkWQNAH4ViE
KqrJvPiOa57suus1y2EKqPj2WZZpP1G9SXgJC5USWIHJWnL8tYKd33ABnOdDnSds/QbD2BXVNV5j
G2w5igLmSWRC56AFcQbiRiU6TWJ1QKXQEKptiwpwdzgQS4CQD6x7hqQULig6LJrgUsDBNHx+AQDJ
7I9Zjq+qVDy8iZWv1e07nMUVIk7knCzqzDua4o9BdV3hFFt+wuhDXSeIPD5Jov3MNa7Daz71JjHQ
4JkETKpxm/pk684leNSjG5tuC58qEn81wq6wpytQs8N3rtzdZ9id38R3cj21ON5TICOwMbca85bY
cbZC7qomyLVLwoztcXfOoijLWugRJWsSuoV6aFDbignTzCfv2FNUSxiyIdCmtY4rOlqucPnSLwS3
WfVosi4ZqSemWNreycrA6rn2bOmxBmVMmSaJERV2eMNRMCTgyHYxKRwhLrVCKyJXNd8+dv/s4lJV
dU0MfRPy3itIB7UDpLuD9QuK5+sdZTDLduv83/5WSpLCwTxMUIyfyKI0gMbJpq4zIk6hSUihRJSC
dlGn+qPMstfsCQc6IuiCF8RTtztAHejIJ8/nMiR9PKZ9fUd+cRVScsZzMJ55wl6wb+ADqtyngFRP
i9ShEMU1AI/R2StO5bbPRsgifDaegVjbrYE88ZaFLViXfCAxnBe4lE7CvVEF8WOIPJZQoI+yoKnD
qzdk5fw4zeSeXUjUZZZwpHQ4kPQMB0t8y780zzYag65Iy4fq/scVuLANtP3dDoEoTDT06cdj51k/
I2gU+R3njrEmjdALeP8nQoQPGbMl7Ib6TfUVGObfdWsTkrpzKRs5HywpwSr68EkxR4GYgy40MOuJ
IZ6GdYQfff4+j1S9iROvVFRk2aL/Em9u4QSqT/3DfLkJSiXHyqXVCnPwAfHsCdJ2Rzn0K2iyQ8ew
STlo5UdUAyfXXBk++QdRkcqnbBTUw0T/kakFj5+L6HRay3jctpiJ78Vvn4VDY/gS7rvtjIYj4QMl
k+pX0Nah4olqAah7PBcMQJi76AtbhJRv03PXQdBItW8M7qkIKM0Lbt6F9A4MdXyjMQ2tK3FnInT7
WSsXHSQU0SIkwmv8pnv8clLjkP8F+l+v6SRFyeIVCX3x+uPFQrjKFWxZ40vvuFMSLu+y6KuAxBXy
pow6bJfGyiymoHipSoJcVkHdGINOGcqTOTyBr1QKwWPqS2wYGyenEMMZFECjiixAvtezJtKlPtOF
sZrW80qGz3pvh+JmHlRVtiUNEv1HLZWbmkiEe84dI/jOKrlFHkdOkXjak4wViLfGEgPMalXaOzSp
MLmxkLIp4vr30KIiO/M3UWSr9l90xeO0rzpF+cor95m76Pq7N9jjEWTF3Nswx4dNzjSWe2YjEADM
CVt69dSssqwU6QSt9eXSJYO+cgbmObsZrC7qPIZO1AqlVIsM+33lBgtSMGEXKBV45avKrFmK9a/H
ygihga48tPzZ9zYBTd1d553ZI8jkI0UeBWxaXTentL2YHONfsYbj9bVn2W+dJ6ZNjehC2W8LaNF4
DWVKFOlVx0wzMuz4tyETWk0JcB/a9wg8UTCezn/5W2SwXECA5KlPkpIR3FaXxT6UqY257zDQA5bI
WlmZyzCHsysb6CaA5nbO8/gYgpQxAGyXeeu20GDdWqEa8VBWPYy/BE3BDDEt9sLEK5v5jrbSdVVB
m1jQFWDgp0bxzs1EHrc0lu3ONZPAJ+Emke4M0QPOnpx+1M9l9mFrBIHVFm6lkkj66SYJVWN5Mfk2
jO83vdodD0T8Z7kQyLc47NgEe3Lga5ZHDSAvJqLEqjRk5J+peIMKG0K2v0dDa2KCUKrPK7hQwav7
SUDwW+JRsTyhB9oyxT3Xburtawo7kO8MgNLI5Tf6sajsvYl6LV3YHuOlItYyadP3IfOBGgGCZgSb
Amm6KbfvFbnxCWQbwQMzASlw47dYpLyj4fCotxl46itMmMVC+36yF3X8YoHZcYTuo1CgveconPLa
r+RV5dgS59GRGpOMbEmSuQgdz5i2xYEPhId7hdpTxvQdAGD3uvDQCptP293eCc/m9qOCmKRaKPeW
5ghnA0A0E0v9qblydJSwSVwzYWfrx7QAjfKLJAl8Sr4MtQFNd2adcGjzr2LcytJC6wr5vPk3VSaB
kaLZO0zUN+7Ys2nxPbd1Szc2IDEqB2da5sWuDqFUF2iPTfP4o1p/KLfQnl/R0QLuZ8Y8BT52x68r
+dniCgI+hU1hp12Y0HAGHzk7ZlDi0BCBbSk18aPBYkvsud7rCH8tLgxpP0oSf4PGqN42t40eOsIw
et/91PPBNmnXkKcutXhFrpvTpgdR0KLRI0LZly3wOTh4fHDUUGsyJfZgRjDWohFhd0yOyBpXaTxr
irBuIQoRCQVx30XaAv33WecdcHGTQxSE2GVsZrTMQZYsd9/6HiYFS/DNlwz/5zP4NhrjyRLEjoyq
wN6t9Xs33BFCQRDxem/dgGVYd209pofVsDSfqP/4zy6dkCJyRkinJYYYLVVqRGaHSM58ceQxfrH+
tmNeYk8K7gpAYgTXkrNyKSkoCQDeqB9i0ByoVwSuU28H3mymBDA83Ehn7FIxWooUbsEXAJnGqtvX
jLh0gVYdn/ImiYtoduziZej3IMJKO8j+CpbjsKaTeReYYpKHV0rfDSnfWbTb+YE5t2CN2wFlJ7I2
UhvdDkKpHtGqovlJ5ZzgJ+9BMAug91+8LrL6TWperv0jQlttYyq3c2fExIPdkUCBTxLG5f9Qa3HM
pHsYathIiCeg2hdjeIeqQAu8wDsrulRBFedjIwBskZ1m/IRMgirtRGT9xA2TEK48WmgEoMhvqCXA
zb6LtVdpi4apwqiQgPyqhh09D6IPGxbaPheiG1/JveRn/gQWXb2Mr6y+pb5HCPpKs3MV30jJnXFO
bSoaA08RGSMF2AnLzTYH2xM4fs+bpdMFD7iL6tUr61a7eCP2TSKedS3ILTaD+PmKa6Wr920zVnil
YIMmEL0tlzqDTAEahp1qx3mxoIzXcpn6SdNXJSFp30iaJYGkHvgworZqV0qD5aWW6WM/xsYuVtxU
O8KIP+eOPTMUmOqVg0IrshciC7aBbY7RWJDy0j1DGY9RAhabPu7evHjmnmyIwpZ0p1VnApTHnJXV
HGDDcNvhDr0MQ4Za979MWvFjzZz7vJr2Wo/F8NvjDHuDLzX2j5rDzpzqjkix+VERhegmuGj2rQI1
0EoM2H0cKicofoo4uOEP5u5YciCwu5/oYqTr07l2xDkn4Qa3m66eNydcJEOI1p9hDn/0qd6uCYIM
rNVfDEyCApb2FWD5WiH7hi5hPUYtyz4EQ7jHxCHH35uApQDgKkgCMKtZAeDjZYSorunqG60S1PIP
/QFJfHfrQT0pMjTf1zNBdkyDvD54g1DPhySv28PnGMkSowSSGI9XqtA544/A9MwVPx9rPnryiRFN
pKWW1v0oiEzzRWSfNSetde3CVAi0G85fGeSbT4if2yjaTSBKwIjhtYteCrgmI/h3mxQ/5epz2Uu2
w3fYQ2QHmJuzyR2swjppnuemPaA5h9QwJhkAvszAf9wGVBBPLwaWjRxRIrUQTgHEWO09gI5d1vZx
DmSJ+WI2DanSct9LLoWhBQJQ7GRh3dH1nlhOju6zErGHewlTs2ZkBpvhCkQgigelKl2iA6JUQHVo
rp5fcJbxP+5k59wtzTQZHJWc9uZfADKzkYQX0fM9HdVT2uu3r6Mj6ZCGJ2pIc07YVWjZJwhF4h7V
WOM9qt/sAONGzF7s6aKi0rvSDySWr9MJY9XjYYbnaGvfZqM8SrRz+DhrA/Dfs5fuZlE/XgXKZSnV
C6EXo3y+ViCvFcGbvH7DOl/Ihght9sJ+Z3paqAa1qRIedxsmZSikteXlzrNLCpzK5OjQPTTdUX86
hjgFOnJOPBFAKrwGblLoR6eVtXMiU9rVDDRTrvPhziXha7/tCjOH3dqr508hSRzk/8R2fkTzu4fJ
3zbM5fRARvIRYEJsp+WTqQLyJ0dl7QOz8G1PcEcGnnca1aGh41nTv1dgu1k2fRPLKcPzzFMprKng
3UpY1vZFZGyosSyLAoA67hq0zeVk46fA4uDSvbKtB/S01ylVQfUoEKfDN7yAUiTj2KkUVf2+UBUo
l8tJJka/8obMbv/AQqXlmU/6Yla47sghJvr0taN7uH6jBBFwOrq5xPLlXu8apcLjmx3NjLuAHXIV
/xkSvr5dNhwbjYxCpgUlLRtn47vNnzTku2/zJKRnMytouGTj/sMl/nlbU+uwCSETUxSqPHPbuEEt
EYynwp4WKKjsLQKcLS9tU9zeXTnH+7aTgN/JuunzhCMVFBn0oPVkwNq9vsH7ckjk2UjgP31sxmYT
uT+xqykH9DEPZ0iuLjpBWWXCc5s4uRT6W4DKlJOBQLbUOyqhTNiGnOuOOdXmoEm93qpbrxpsIdtf
nD8fZq0dfok5+D948QJJow+Xb/FBJWx+LT0hZecsDjj1jV0STY2U9KA0Arq4ZN/7rDe1Mvakrdi0
nEyuFyH3eEgN8dHCOR608AHJwSaDRR7GfjJb2hs2JfdVRGWvTciGjzvac2zRSNL5LAh/OS93SCOV
0UTnbQoCe7tnmEmGkEweyIhmIVAXH0ljnnZv8ic0DMHcICg6Vc+SWgiG3gAAZ04soSYG2Xwm8X5y
ZYeXXAw7+zgjmLus2SVIslIjHN0Sg/W9u2sCWLaeENOWzNLPPcIJP8KDUJo+Uqm5vplj1EflkWaM
U2d9VUsjZOnXqsk+Ya7HXJT9LqWZFVgxeSkZpIBUStEEBM12yhQYowRZwX5lCD0ZZN++IilQ+yqS
SDCA7q+A5Xv2/BZ9QSQZNA01O2OOryBP1+ggbqjYhDSFgAcUkUdPNuAdSLzVHcJH2s0ueP1pPJEd
ckFcnRo6tAX2K2UVvofx9VGOM4itYOSvQty5kUhRtlHue8iIdOHSEekBdxrB7Kxd7eYgiEKdAIEI
refrFQ3RwChMehA26vvQu/7GirKNhxdezBVoU2jX3V/rIvb2gcKFQUoii51RVqOxcSQ8fINVZGt9
DQa9fGHfh5m8DUQ5L0eITKn6NP2NKiMrolsQGj/IKpmEZ3v3O6EfteDwdUwPDvfaE+cIGU3rHTuF
kEEItecVuQUiUWtnQONNNziVYqEVunhP85cjBctCi3KijS47eCUNmG+f5R0dF+u/jv0bnfZoCI2H
JyOdXMAu/K+rDP56hrY942Pgu/I022fDX9GPbon6w0lro8vt+J3IFGe1vf1mfiLGi3KdgBfzYHg9
qO1eAd7+hjeOOmLotmKHbOBwEcsJpha4zLcaavlheCiekhA/u+y/RB2KGZJCfTftjkYgUgCH+4HG
OeMG9iRhOs1ZuLfN85zWZLVtyAeZVscSBTTOgXOT3W1SrN0ZKjP7vU84tu5kCjqxKf/dniBtOofJ
yKBhpW5aVJ1oi0bLslgQ9NiMZ54L6HZ7Qk4BtTxxqMKvSZBQ3tVvZfoldbCJnDbUboyMYXJ0IVhD
G/MO0/DxV1aFM99cDIm/mGhl73UQ20S9LDRRRD5Hn514GA5mHYhF0TJq5+1zebOO4Slb3i2/aAvY
mTVcvyU0URcwC/pmrv012duJ6sH/xS/+Ylk/FcKD7476umvaOoetl8lMh4Vfcex7BccBdpbxEins
LJ1sVMpvqEhO9XEIbvqOk01eFINsTpy6B9YdYKiilXIGnELvWLOIUzVuiKvYVCmfw48xDYSOFz7M
sbiWI3IQSnf467nY0DvSJi7InxK9l/7wltttve4Ewmt/9+hktnYlxIefYYPZMT6vKS46YQ3vR4xx
YBti+67JJVM2zht0KX982JEdtl2n5VKTV6jI7L/Ad/+TBqzY1yXDyvf6tfjdEIYEhiUhIfE2f1pX
4+9uzsR14q/4SYk7vVk7xcVmL41S5dSKTBUlEw8oqTXm+tsOE/WQtm3QYOwxqb9OFwksR7HfGM/R
HtMfzeOJrGmQlblt2NCu+YcffzEePL2t/iOoLqqtEMPI1VJD+iIFac0Nfdkm3fgsVZK5DxAIa9Cw
5vIVvPpe8KOYS/KSFO0dkNgsSXESXRPzMsanAx09AI9RCShGM795+CYcZQJh4XO8C3ugj1y4sO1x
J96TSoQISr22wzNNmTCw8ePf6z7wccqckP+Y3Pqrs1suybM0RQ0o4WBohf4oBB/JJcZqCJz3ae72
ECYhN+aGkJwLQwgrtSkZulGiX9y2o0YQZTgM56DF8yoxpRfOkTKYCP2uqXtWE/feM8aJRO//nVUT
WdRdOAHNaVUYMWW5QbP4z5pxn4niMZe7QkZTxqxD9nZr+51LapT5jSASIeEvsBXavOz64wYmBQR2
LaQ8YvZx6ODvRJ0lzAbZUR7MIF+RwXFtwrTtlxV/yHczAuuamPHKJP/CMIS3FIQrP6DLsJP4kBex
FHHwwiBtbwruw3fBWObdcvQEgYXOySY3vq88C+8gvY5/PK9t4kJVpdednNy2bGPMMVVjDtRfZALE
luNcceaUZ0QjKnXpF7gdnEOUjKH8DxxJ9w54t5vkW0wF6ERHTSfLzB0G7pNiLPBZuXS7UhKU2nt3
8WILFYI/xt5B3pGWZoqf95056YI+qVorerXLF55XAXRPGqoxyF9NYwnIViwdPwsN/JgnighKKMYz
INz1mdS4mvP60rQ8Su2E/FNj4pRrwzDbkE3GsPMdWc/xynlj4BGCcuE9doPTRlMKlhtZw3i+YGvT
RKE8tsoMUsrjvAiQRVvOQCuLGrZ9ID0hqTVGOo0fjXgFyNZ8UCZWVhAsDDrZpZctPJiXb4ZMHGzj
gcuVTY8s+ChH5IQPhJ9h94DYfBIkpfteCnrvVQnTWhAwS+NdAFRxo9p3vovgMy5bbFLx7SCYWmEt
x5WdJK4KKydj8A4oCdNWRjRCBH9gOSiDqB2HUnQlSGxNAvZhhOjg7tJyivHPUaC7BHKXRNIak6Ko
m8CQxsAV2XTk+s+3sQxfw8egpHHmQaOgnr5ClcqTencyB6UALxxRFv/P/L6kSvqRDgTdV62ZFwNY
0yVGZkXdMw0PYffELUx/IH6iuoCDXnk79QtAjEjwHFsD7UxTrcew44c2h7w8rBRmj9j2OEsZGBlo
RTZaHMIzILJBqoeZ+QCGNZoawUue5XbRMO5uKS3xrGRkDSpKe1wZlGfGX9VuiA6kSrOhX9DJMhrP
bkUDrBvGNEiJnwk9j2epMkF7+4DD71Jtmg2zYo1xwNeoE/5aKfSIQjJWcvqhkP71x3YYU8bAGQ3I
gF6iBRTGUCcCiMMEi+BcEW9aW0Z05LbzGnfviZNdI0hsgBxDjyxWRf7s2b83VETpiPxn4woD8zPu
Am0QVJN079zlLUtrhOZb65FC4U4mvRgLCOWscpwtqYGqUUkbltERG8IQbylpDFrqZKbs1rWwwstT
S/jA2rZSXNX6FStAoMemwW2oOS/lILj06ylC6m79SBaB+WOtMn5PsOcWfeFS8qfsV4yIsOkK3bJn
E1Gz5xOsG48/tevX9DyCy2X7fmPAXodKoeUgrEy9F1EET/r2uCEuLc34n0kt8ynUBluiV2czgz3y
c3Hzw15AS6qCJkl4krnxb9f0iVbeOl5ROow2+F3rVn8iq2TTi6LHlsVLMQ7uSr6Vah9+Ci9zpSCx
yXKH/jwTJkwaZcrayv059cts2tq4HTVYTbo8y08gvtFV14MQOrwk9Cjwzs7WYDbuuZhLJWIT2oRU
u6RUDVZ5KLd/rODLimKKUj790jZW6yPyPWIsi0Z++VfrCCuBUgP/Doo8yFS1sKz4H/R6KaEnD7EA
maBUBbz/6HvvWWYJycAbSnq0799plsi3jjnXqMkbqMW3+hPUsxjU24tJ+mkTlcp5TjwrZqLyzQaS
CTOxdDh87D5SNmrU2i9XYiCsXOd19uTJdZHr0kNKS4a5sAE79IHGR7coQ/7qn2DKXzNdrShp8FMz
SB0Za3TgTeHywihNMQojzszjIRvd7onAfC57GgxyPvvbVDBaSP9XanxphoDGFP1E7o3C8jrSPQDq
mebH+nc2PQdp2HiZYPHwhsJtxGqZsLwys5ONSBXKljFwIYVGV1GrLC+ze0dlHWSTD3MY7aChhhu1
2/Ok69Tg9D2eCPmwn6AbpD+VfjcMr91pbT/0Vc/aXCMlBHAMCFATCfwdlpOjsKOB1tqhtZP+3u3U
Dcxr1I5XfRgaR8FoPFt32Ir3HV5/1r1kzXs4peH3axAaBm4Sz35Xy7COBKErbZIQAA7KGl/JoKDT
kWep0XkNtxRkq2EC6U6uzPLhjICP6ZikAu1SJzp/3z+dmHykO+/QaZ9xU9LZ7eIYSM1Qw2YcJmu3
/qMZve/2Gc0vD9j+R8WXXRN+WLlT2Iwu+ZxxwrMiI1gsZxBW838tB/VMI8UD1lHQ4rr6gr1wef1d
FqBnaHOF0Jgl2Mus0oH5QBdryL/cCk+vdSYFlYHw/r1d/j8AGjRLFbYNdRocXNDFNftYog/Hz+1F
2uU0rZjfRirhT/OUNHJJmDSWAc5xgWhw80Tb2DdwilljC8qd5eSQ/wD4Q2s+xRAsL8q1sn5eaxs4
XCZNxe/wKmjSMsby1hYmzpK7QCYT2ZQ/13MWnt4gb8OWEP1ndco7RSLbGQoKWJEDeZQk6RebWmYV
5vgfSNpmvkwRe3MO6X3TXZHaSvRmwMDyIiKsI5lU7lfu0NZ7T8luI+YQZVYDr4eE8xqaqOQarApU
piK7X/yCdr64nX6ZQNmvXVRaTP+RMtTarlGCvdvaL8z9QyUYEl2jCunKyQES0Lm+P1YW5waLVTt1
BJ0R2o4KIyuOtPDamokjaiFCS2rtqUpfJavWrwM0Q9vywt8hKDcP0uOeusQIYTd3K4hz1QlsTkr4
Erf5KR9f3COY8pzfiI8awh+e8cYVJWOJP2h4OSkwk6HIQzc9TaoeWPyCDCnaIjGPRc6XQx8Jv2Ww
HgCFQV3OViRnRW0GOQZ4G5q5Bj05UlJnF0y8uTqv7jnwZW09Laegj9OdNK5fwvH7JDDL/rr5Y2es
I/1WrZp/9vhWtCILVpS2QNYBJc3Y5fYt7ZbhPgegb76J1vHzKtyQfLSJd8JeAPCVESSHJluF8Dhr
oRa7tLrQJ2VwrJ+6krXxfKukgpA4ChxLtqGsqOJDw8e2W2R5tB4fB6BvMMBN+TfiN+99Clg+nEMl
m19hxLocKkaSatxkk9XIkg5X2yeHUTJRORoloPix6jT79Rrvs7P82N73nZxA5DEs8Rs6qwHZI5rl
CsresqOYdS9r7OMx74ryTo21pVmysZC8dlcQ7OeHljgqT/fDvVju4uHOTY2ACutAcmAKtO1ZBsIY
o/OFiEjItO9vVokif1MRHDPnSXt/PH1TCWmRZvgStBkmUKd9Mr/BcDa5EQ4znfBaZod4hTLcb+48
lSFH/Tl0PU0GbPu0JT8GEE52dI1ogu9QLqa/rhWfATwD7pD7yggfT434oVuNYq1H0LRoiydAnGFZ
qVBtBgydy1TAC4gbviptEGq9uKqVtlS+PADnO8RW1xQu4KtoC84ZNg+rjCMwZA240yadkqGkdW6o
viWkD2APOi9WaTIgOBCvO5Vcku+eDat7XXvPYWLId9/yxP5LBGbxr84RpIBkFkWFMLLbFE3lDtqR
crS6cMmItokMkIlIHfbcREDQvd28383eHiDgDNb+sBIjz5FxgtN2Du9VKGhOzjWvZ2BJDuP/c+Yd
XB0HsjykGmnhVFnPg2LOu+VRo7idU7uMsy7JkKaAAfQ8cA6ufVZoT02YFS6yVAdCkdh1IQFgsdtz
ylHaoiRYG1AtpNhfwxV1dt/Rx+ZWEIJ3EnJXYTV9d66rp6kmxidzElZvhL5cWaY2rcGCBj0eToO6
/3nTdj9sEwkaJ3r2iQDXAFuPh/XzeQ6KKLQVx+tx6mi1X5dsGI2EnT10FjEu9HmJ0kYKjJU9+YwW
7yyaXFcn+ECeEnLcF9jz1/cy0ZG04Ad4ENNk8ZQy95/7+PJncXOnNLr+3hUTf06yjgVZ3/fUS3r4
viWZrPsXjq7mlizQ1ulEYw6tzBuDsOI1ZM0K3wdt2lIgky0HiyV8l34+Fz8x8EzC69v/JA7ySqzr
C8cSfypNBFtRX3guVsMIfuxBN2W+9945f+JcP9CLMkwsyuD3cbm0akCmSRwzR7nXii8OyGZe6upm
INPUCTMCcs8Usc6h+Gmg6sU51TKI1Fkaoj+IwhcgM0Mty9yOmKmMuKPbCFNrFF+uYBF40wKmbD9D
+ufuRfTfp2BZm6U1Oq8Juzyr6huPF+p+uUYzHH/79ZaxR8v6m3wjXvY2XBI7ZZey0Rc37ize8Y+T
G5gw0GHR8OmNCoFaqBa739G02kFyX/rM9rDhOryliITKdTCo03R0TC2hqlKTGQVCw9W8/OPzEak4
WmhPdJcH36qfwb4/B8ozdjf38mrm6uN8yHYdxzORjs58cBVViVFpMmy5cSlZ9hODCPMwkrVPkyN5
PajzIb9l40kljFBcgMlXt/qRX01JD80zRYBN5ztQzBMxCYfotgC49YIzhwbobuadrLQBNQekc5SG
OzzNapcFt5fLo3WRdMDt9otLrt4Blv3iNo20K/CIjL3F88eDDsxPXSfEGOdbh/Nv8MkiU0YBfi36
mg3WhMerFU90DTX3+IdnVkB3MyJTUKriEoHUSBY2F45plaHmQgY2o17n3paOYVTrKlYtcamByOEz
ntAe/HyRSKQFqXZGwONbgGdgkE+n590j5Whi8OCY90NPcDY8+A9sGQ/km47+FCv6fzvFzd7q5pSF
aDUA06WRqpbhzsglbF3D6Jot0v4CW3TJ3pN9JMddXjQn9YEr3s7aAfufItr7bQF7AldDiBh2mAft
Dc4JKKW3OXeW2HjvCE0hxfYrxIRSWCgDct+8lGaO04C1jLV4hWKyhNKm5HyEWUK436gF6vfiOsQv
qo9WLiOCPZn4G9nIIRIuAthGwQfhTBGiZCUzuuWkSmDpUT2xJASVWjQdT6v+Y5WohTgvIeXyzf92
JkUVCCESz7MoJ5vWmuu6wI29rco5IWMesySQxDiBnKV25MBOglxx88ojT9uFPlSnwRKh8ESJcXcT
qz9sfXXdrxSNUMH71wtNuIzP2SMnTFSDm4IgQeSMaWvvp89cxKiUsgiBh0Mtb2hs6PVZ3ceeUoVt
5/rUJjNdCrNf8hWyRdJKzYrZxcJk+Z4GVFWQ73BNmAZV6pPI+3G55oXeJp79DMh5GWY8tvC9q2eS
6vmcqSsVOiCjwJym8k6/t+YQYwF5GduvvhTo+hb0YM/anLAjHJzqYBZ8TiCOXfUUNzZWkA+OrBGM
f8ry8Il7Bsn9tf0fxhWMzuTdzZJoeXE1aX0To0WqRW/JKJST7ZCh43vf9/SR3IDIqY3ChSFXPxnC
twn/IcsiUPM2c3cvsW6/1Uk4map57dmQObDNk+/4VFp1i89pVsuDzjZKkkANae0e4h+ZHdw/v7N0
r1FadpK06rrHMX2Sl1vqtq4+Byn0MghPuhg24UggVOCP4oHwRHv0HbvNI9bdbLBrEXQBNMcilxTg
CgEEfw5C886Kj+lQKJilxNK48nplybG1U/5Z4U5UGBpKDLA2gxqqmYLl/S8YMSPK/EHzfkVySLjG
rRgfgu3RpbsByz0cfiA8Z5n/nN3pigbyKtiVXXUkeZ1jMMi29q++nVY5dXKkKfEnmkZ3XRAihZtG
sWBEA7NB8QAZIygd4kuotG8VNqQMeXjNHsshQx7VYRHkX2wjh3JTq/D4gMWO4eedueLhQ+/4JXK1
xd3xj1bWt33XZSKD0ZrC2psyGKdDzpakmP+DC5uVVUkaEYOSKaVHlKSh/EdzR4HbcL9S3kyjGh68
CCAf9zOk5ctN8lpTpaeCyAwKoA/3U6cnsMO6quEEvC4Tgx5KhD4Aegf7Saj+egcrFCmqKqZiuVrM
NgUxIV+vfC225Co2IT6wVKcAi2EsBlBldouqesGAbAjq5dyPsTlZSjFsveXxs97xXt/8H8/xnUg/
Q36DKTocddt8CgqHG8p3ld1qCTahEJRsAwQBn5F9rLzca5bA+4DKI/HlCGgF1778OltORmib6YGv
XOvS8iwMis7ZsOvbtqwnbMkiULN3xjy/5afC56vZY8GTfUX4QEA4SyYwuNkinBS1cn+ThlF/EQT5
Ub3+8eOVOxWXmg/kZkBiqo3VKLVjd+QlFU4Cy4dNadE379U48hBhR4Hx3XJvnFW5z/AkRJjUM+Mv
1xcnqQNkLohM9gU787JC2EQpR2shMrCS+20ZIOXNVK8naJUQs8UnvozB+UbV0gnlrDlUe3HrjeXx
n4JPF9aIK9UqLXHVeC2TZqgAWIuopkWb430qGhKYg4xRXBVDrZDItbiR75KzWi/zbQzQJEkmnYUo
qn8j84PUXOz3IB95mhkUHHzqqpafNRcm4CfLfhIx/zZiewphAyGG4c0IoOVBv/o4d7p8KwLi1xWZ
Lfr0m3Q/cgbSPha8e/T+JQA5xJuw8HJpqX+aUUHhIg/S6UGKVp4yAafD9FhizEPgJFV/wdxHPqap
TKn6aep9nnV1dMhT2C9RJPHKKbrj/BzuWYXUkA+hd8muWI/mCYA0o54lYzyL5EvgQRmh4ml3onLA
ASdGJeBN9H2cPnzMuDStnPgiEPePuSzIl1TVe1LJTSItkFn3seVCLIYwGmm/sczQXZ886P/FNY1n
eg8YeNRvKL9xeRm0JOdSjfEAaI9hojq/Pg0QO5Sl/uDyWx3hgH765wXqAtWa8HPkHdaymbb9bBBU
nVa7578ZlHKDIXqBrsVTq371gQZbUfOZJdgWPKEN2ZfCyJfTjvbYkFTmmHIM5n6CIK1EhoVdn4up
5svIapH9wSs+qPA2dgyRl/B687k9nbBiVm6hi5kvLyOG4AcPk6pgjDZu2CKSZQOEvxmZgrTRsOFL
oZIfvHk7BZDhA7NQT2Pz8Y+T5WYAld3G6th6Lo1wnpHhmvVOzrJH7u7Gldhd8cRen9cvTNEQRjbb
q/GGjQUUcUr/WHBUhKJKMb3lS6mFHpveQmjGV5ApN/rCcZuL4++QqkXett02yNDS5XY0YFRArTdC
hiiBfBnjL+GKVr5S5AT4tT2MEm5AnLRfdxA1bRw0aI8J+aY1laUQedBJ7yPEQMFIm7NOCJzlj0vm
mfD9RfjZes0jPdtPssbEjfsTbf2ArTnYZUR08+Mne67z/49thYVVWjMdXYa8jR8JN8792pVWI3pa
m3yBI/6Q57+aG1pzq8NR4Wd4D23NhoeYUd0Afv9aR2RSPHukrIhc+/0Aqp+MjGS9SOYTgYwD6qN/
hYYKhEtqD3lZcgAHU/xbHvL/ZZ/J8cdhk0VAW6QdmE2DtEGPby5UiIOfRzGKXVYNYg1dbf2nm4xt
zpzQi1ZcjF2cUoVzCxeYHA7KBqgo1TfcyITG4IbCc9DFUo4XDAUC9UNSAVrAzw2exREDsaMceREn
+eD/w8zi5qnpzmXo1VV5W0S5FPNJ52nqoKjdoZPHP2TffnppgUUP8FGfUp4S/fntqFj463SRmDtK
O4eVp5fJvd+oDiuT7ZxFfzL1YoOfyFab4dVDj/yrSEVk9pBM+MflGSpCnCSiUqdTeNDHuvFRRquD
VuUOK+APo8ZN+TbLZJ935qoMytRUMe15hHqHcB6kLPPlf7U2Xv7u4yxvT11IqMz3GQ7KM6X2rkWq
WdNvRvA3S5LxSlBWwHNH1tAgrWA9C7E2OZB9pGWaRxqA8BJfe4R6DcrWwbf3Y4HijEvU4RyVNe2s
mfE2OH8aqyau5Fg1rmpm5B6E8f1VGGK38ABl7qYKH8ZVU9cD2PGDJbZ67P52o783jou1trl8vAMK
REVu8i32p7SBr6U8pZVNcfbm5vQSyWmPquPf27Y8ejlz1BbdPkEtpH/nEparivZPxbobyApnoimp
gQxw+I847ZmPjKa4pzHYd99W9xkhfWeV1Qr4LQWliI3dw8BV6GuW8nE4J6u7d1+C4C458hMrT56p
7CxQ6kv5PK1ttqGRbO9sFu185VFcC8tzKTYKoox6mjiNsCuugYvcrmETJFG/7Q3CpiBbOLkC15VZ
B7+UaOW7Qt5ash2YB6rfnP2iGOhoJiKcPZkL4k0cFKjKVqPGXROnz/8kKU/W7Qp5RfKd9gUctbHe
VAuXEby/XERA6/3tCLAB9obA3jqaBoyvsSF+F7pN9/iQQu6eqViXhp2q+kZM5GpO+6ZP++AneAgp
e9xahk98DtDxsAFqrNXaoR9kYskvn0No5zUG0PPvybmtyV7LxiQycCQ2WeOgD7AJoTdYVfJ8gLdl
gICH8ldTlImuDqbfh9hgl7jjJ5XQmgmaAxNJyHlWrrAn8aMIPFGLGl7yCHB9q9P1mQEwqOu82nIf
z8/INmbPrLrYfHb7aO48t5JK0yXe28u1JbBMO1ti4GSgGGJMeZcdqbpx2Ha7fKtNAg+BD4azwwoy
IKWLtpTia7hyabiezAwSvCEura/t4cCm4/NvwM8qKWWzQn6rSjuG5vzwhblDBSwjRVx0UhQDyJTQ
+KM9dOaM0wulf8m9ZUPbqYuaOPNTowOZRjHIbjYwZOms9BCduYNxu0g62j4dFJgzBfLirW9E7DHd
JD2jCYdSNHbLLG6gi38+st/4uZaOcSNhoF1+8Ub9aD3Y0S336RmBUoFW0gqKqU8iNZ6s2XfGtxOt
bRsiSiNFxjgVwozP7r8WHvGZhecf6oFTJ/wAPlOiMOQUMaH35L6A3nIiejVEGb1935dUFfiTMhsV
0YYT6rCPB/FcyYSHlH1O5zzrNjqxXpqK0DH9JAjWLlDoWRFDVO/jDagIvqhL8tizKL32vDcyWCl1
t9bvLe69XV4VgWzZ+oi89Dq2fB0QkdSM5OpMuiztVEG5ieBht7niHcXWg9qSs1VuwDv+gWI51HQQ
WMjwES6IOoBTIeE/fz+efiYfPl2MyU2s0CREyegae5yBuEKNnaL75wlqM7Q/o8J4jufkwQXI5P9H
zmI9QHeBaoN8gpwOAPLugSHTooVXKiyAjnjRPVT5wZ18lalIc2YV6DHPV7YqeL8+UIfE670yJ3Tf
yOI7lQLNpcMGkHo/BpOX8ZVAX8b98bzWqeYuxlBzDZRPETJjP9lx2R5mDxWMUxNMU+h4sTNrf/3m
6Ygx3YY0+5z5hZg8oJiIHyfha3PQ0MBLgtfSXRQjBCAAG00F9UKIoDwmsp5a8m7RdYQGI+XHpJpb
FRqH6nGLefGIhrDHl01wC2ZdKezSj4DsCiUt6IDLCShY4HsIa0SIpB+pJ38+I+3mxA5w4hNt/54T
6Ut3iZMUSXzzqc9QqzhIvya8CqeMUx4BfB3r1biW2/5VFuuEbIQ7rh3/qCSGDvXtXR8PKUIb7jya
dMVk8gIak9rcRQKn6JerzzpBME6OGxU81T4rjDHXDbbH0NxgALbYWXeSrTFN7CirMR2aFcd59WTn
K8V+fYN3x9iiTaw80FRGyFk21hK1vOQo71sOJ76SrKPQ7JiSTI3fx/atYnhmpHTgSWUyE9oXQV+n
K8jA9OaPwv/YFlhUqjDBJfKM/l7GV5on6mErpkQYUY37z8R7ywjyShqORRLPtJvTlaQjMQNA702H
J8Ar6PY+XlqYHfVHlwpmfa+qKkMZg8KEtbtEXpDjL3RVw/pkcrVG2N8Jl/7fbGI2AHbWO4gZO4Kr
MipGip2PdQBw//LSGO+fhAg/WSUT2NnlV2+ey9cm7x0z5SpoXSR7aTgR93DTwtV1/mRV60aiqPqD
41ILm4HOmk6IuhKI38TXYEZcFYPGJbYYMFnNOTBLUGK6i733U5uaY57D/1j5aGjb0b5ivWbe5KG/
bGvIAAvtFxATKDLHgXfPb310nOfVbQqbbNqumwqsWLSY+m9BYdQUA3JwPh5UtSHmrYQIvhi6DCDO
BpK1+SMC9q3i/FM58CRkarYoe+EWAB3iRoCFJ2E7OY4kthCq2K9v+3vJhLNE+9TqvUaez2AyeGGR
/bCp7T2YzI2k3Obm+824s19J/Yv/FxUBqHFY9WTqNsSkrxq4+kGcmqlz550M5ukaPU4MIiRJPUKm
td9CvrQaHZC/SDIJbMfO2s7uTOBQb43TjLM62oPFjdiVgi8yOdfUp+nvLH3AXfMMHPuaP9yGKXl2
eib6CERcuXrdKtRoYacE1IsvNkSthYaoAExAP+bAjzhU69v9++avNOm+se9IiTrbJt5VF0j6G9fn
7HI6BlQ2374WpvOuHvEh5FAiBVJZ14HhfwYIbR9mKMG4scmS9jpjt9ITPHHLHji9Rtj8tO0oG2du
kokfZm7qwfe2WVHf9+l11ACPqlBtYwLeHbZXGQYpULfiob7tJu1UTSMIFwErOQqRAeHZWFkKq8Y5
SpL3ti5RtnLtpqCiRUcYrIo0Vzv6vGX3xxKL5tYkIwa2O2qZxafhFrEYUsUXmmlOpHmL1pfZOp39
mF8uKhWcR983wk8BZuCVM+S12W1LXLry3h1V3tlbBQlnUn9uQuCdjSwWMA+hWkt5gOPTUIi9rIn7
z7HFkpFmxENxtCqbTRhPrpAy0MofUuFN0Y5u4jpsOpGpwcsigYJHS9/Jvvd7WQO1Tvo0akAUcpLj
UJdTKQBUr5sNkiuzjq3iZAdwXSqxTWCGg5Y49+peKMnQUfMjsNUL1miNX6ncMxJI1LPcOIvZybdP
neDHuDV/Ql1duZtTtswZG347fisGM6+VNBa+e7QGOj43p9wqceZmCXI3XR7m8sltKMfNXXvVqqRN
rMyVpiPZlXU/VcVtXzXcmsCsguIIO+84uMFttU8qWZ8GR7hy+xUj0HDl8BO/7RVTgh/dUjLUZfIs
h1N9gTMfX+DHk/AYToYz/tUY821Ug03NyfHYRJkpX/Kidz8Xr9vEAOzngEga8hAVA0HcYHZ3amYr
T1oO4e4qVesP8ytKM2ynGzqqcGx+m2GHh9iIKHY3tL+8QS87tG8XoVYLTMHdjNxCR8YMYrQcvurF
69VDqwSFgvgcumZVfxzVqhzu+6fbZ3G5fthPmuORa7YgX/W+o6t8QJaAiWZRRt9AckIPsBYMw5h6
Dss80vQYqqg40dlOhBMZS5JRCyJm0sdXy3tPevQgf//oQuFchO7uA4J/qZKmE6+fDGsU9MHHlxeP
ATjUMHd1th3g7edwS7zUfKSS87qyhs0F9Qo4Wv0fdfJwWp5iRWj/4J2AQWcz/ewMSjZu1lJljCPm
ybF+DBWSEAIYDrJHYR6OfdGc/IhiWePvMIIoDoPmlhhJPKTxYlyBNphADsZzD4J3tjEAJMXDDynq
3/IiQ44FZ1cHz7uE8NazrinHfcbDqgttNt0wu9Q2Gp9KyKWo0TWni+xV9rAKW3uRo1CCnBhPEIS8
AkKRL9G6fQdjirvii6TG3AsRLTm2kwefaquhBKfRMGFMMC4N7YfAGYXeV5dwtl+Ekx7hMm+IjBew
E1lIsN1AT/OBwX4gcKS9pjF+vRwnLHSanp61mVVYkxwiw5tkT25JsliOGbmfE3zX/x60imKILW1g
NVZRfw7LnMFgPsSTgLXfbC+XFxRIiVea4Dv3eijkZimPmdcywnfe0hLcaYrkbzSLmG2SnVBvUOdr
Z3mbn9iwiruB4wFb6o+7f1+xsVBDOHC168nvw6II+aFf07Q9EtiBciX1EHrj222mrmiRNXxlaVW+
c8rwpy4FfyjJn48d13FN5I2t8zRif+B1RUAqg6fMKBAckKVTKJD2t5oBOvAlXgRzEIGGMKVB3t1U
52tpRTV7MIdW015iR9chkb5SHoS8jL3yuAF6CjhDMl69oTxxxndRqF3NEN2LlrwxE5DwRR6PUN0Z
kfaaw+6nA9D/E2SK/3LWxFQ4O12Qy05gWTd/zDfnjSzHrPoMNmwS/TfG31FJcVL/5snrRZPKLdIa
AtrH4HxveVaE9+ke0wxZ6A82I0ek8kccjwy9XC9OcweoNKWzB3y0iKmRt1WaSFO8gWUrcJkX6hAM
lTAkolcxhD+k0HdmJiwbqmboB9mpj3ZLU7HR98G5ESvR8/2zsNHCj/4vTk12BtPUCSrovadqBB2W
cCzu0XM0EoRxmWcBabMtNodoEiJWyBVIL7yBumUf+mkRB8AlYvAI+V3SsSs3SPYHPci/G6gWUDFz
eHZ5lH9r1aY8vPyd8OrNqhpxI1i8DKM6SkIOyXkGcsalxcz5q1y9nwkjq2TMy4XEE5fssDQsdGc8
JZnNkQ/NVmaizV1i3UTAlGpb5Eg5BiG04D/KmPF49eRN9dtjk/YBu86ISg8aRCDcmBHUV60MdUcD
Rz+hvUsxQi0m4p8ao0Ff4kV3jYZXoLcW4vnFyuEQhHQFluNjiq6hf8yJG90GFjwMPJtHgKAqrdKa
YSS4zxAhJoLXAw/Yl3BWRalxQjZV1v+I4y0VCMvUlcrSs5QnVACORblsu/4AEuPMfMuh4nLJOeJ1
oVRiu7iqN+IUZa6XfCMtPznkE/2gHzy3B/4pZHnhAZ4qlirNpMlMQrmnHVdruYsi2HEzoJGyqVkl
REoA2rkNrGcAxPlKycBAzSIpk9TluBGCDwGz7EKnx0NDckukaDdro2Q/sebtcVR6eMrGiBOdFD5z
IpqfQFnahOXp7yIlVzebaZZeosKBao1zUByGcy56vETxvfifE5mHdVMhrrQgyLyVj7yzrMNpD5Tc
EbNQbQ+JhZFmNbvzkSyAwUHloUSwPLf53XCXZixMEdFZld/U0HoJWO8LiN+ogfPjAeeYmdLyQZbJ
JDqFvb+LVgEST1ZBjXr9PQhtuG3NCFJ8MM6jNwVpnDpncdSGJbLKg6Brx63oU8PKZsriVuvSyfNb
2GesIrs+CNtYNXqTiGtU4GfezujqAXy5i8lCc+Zlv59kyfovMY9xYSDvSNKJVjDOlR+zGRSZCasw
bb6oCRFUyjXuFuWdKKj/XQ5mv8KwsngRQGwYDI59hB4rVwjEuge3MdgB+7p6UYU7+pJ+rzaewJA9
EGWWIcbGVx56VZRtof+OpPBx/1Gm4fG43yls/ypxCQq+sYtkznFfka8EHRk6v6wBUuUUzBoF7M+8
rOVuERTbWMT8qy3oGgyh9dg2CetUvmsxQ5ar9lVo4+fqrMeFkaAkjX8Hcw3W5yKGNp6IfRZ+QtJC
2t2TYwnfxwL8cjMMXiVc+YPVg9Dt2PhXTGimOM712eMv+LR6ejTjwp56jRC/hTP7DXYvBzZyQ/I6
WqixRFPs8FXmdy5tCHPFjdOFmO+2AKHG3r+NBZFhz+MS3lEY2gCj0fHyWUypYhYX5fJvgbTdcUNR
hYjm/carAbfuB+dkwxzmmh+Pug2ML6mXYUZJCDcFMHmxISH7dqBJqRfUcrGvAEy4XJBQ3NA/H92z
qzWspNOrswUnL2YgIMkUZU+CDulsORKYr4Tb2pz5D8gAN4qEStZD+gUYAbowhe6rotEguuiQv4Ry
h5Y9QgVZAUE3GO0A5YFCRmq66UQlAFk2VyB86WqnMu4s5pSQQLpDOt9gp44uecBUH2ztRqHmcZ5z
rJdOyIMeNxs9K6aCwGGf/PoiBGVVo9SbUmputaHkRa8CKwMJIshdLRYGB6gbeAhHum8krBlI3MLc
e6WgO2c8KjVlmbbu35+49gaohcuBYKalmhPEmJHQb8P1Jxym1P8XK8H7Dt8A2vA+EXpRxIZaU7TA
YghY/2cYrqOvmQMDoQlDafSZlLpMzcyY89Ylbl/GCiwcvapuBtfoEnNhxV5okMoHm3vkrbZlJvKC
qemubamipV6NB1P/RmCbL+Ztbt6ymRJfg+EM4Igjwy9k1M15lABA+lO0fGHmAy+MrAnqWheI9YUS
vGx5x6INo275KWndIS5ZmTH9ykUGadVwiexjrARQ4AK5leV9yIU8qJaRH4owE0EerA1wz1FB66yt
zSaeZIe3oo1xTsTr9L2IeO8IWRlCG4CSeJhA7rD+aJ2Crs48kwyy6Z1+rnoEh7Dh/+C+A/aAR7P8
OC7OhRB5/S6naimcKvggKZGg/hGUtHIfRg5cNHkCx46Vcl1t7HsJmF/vmfPt9Gbh5FoUafy/ZqDz
4fKc5v6V4OxB3uYixDMl6ssiGz/4ySwuatdsP1fV+hKsM0BmFnT5ys4gF7uWa2nyFgDiS6WaA8m4
NoOEtp6uH8ZjrKtkrb6b/xM5pNR4SnLInX0R20qzm48n6vatHcUrapvb7Rego3HeZZMUQ1NE01qC
LBIuuEKmD81UkYfLcz1g9tMiJOgeqatrlGj3SUW4ozMffDSihq/ZhY0Wta3qAzys7c9fhE8SB8y2
WjMfVIMj7ndLcCr7IDYkkSF4K0Q8k7sXUkLmpC4a0u/pkx38P9XBC2WMjIYw2pT4dMzEBcojwkrF
Zwns1qDqwfTJHoDC+Q9biPt0/DpK0L2sMNWk3VBTZwcy/Ezvq2rkH+K4RzGqPz67rvG+L9HeD79g
3IzdbIXNF4hB7P7o3B+MDbBkyFR8/tusWDPejKEF6QAWtbqA/WPYtMyEFUPpSr+cU4XbLajUfkZM
oTZTnPXmskYxUly7VzhZcfnEQIpO43Ox3715RnTVlaSaBTNL96mHQHfiqVAa0xjx7TFAaIx/He+1
8a4RvIyQBIVHBPr12E8pqeUcFkqs972dRlCgAEYnYt8i7UXdMiZnQjYbqC4hANhnmEwJln/hOvSb
x2jYZZWfDnRD/a1BubLgg/xaI4PCANYToV7hovjJJGV9HDUFexAecN8xQINBLuCzWYIy99XaXpKN
I9eGMdYtE2ZOSD6ggcJwUi5L2YPzPV0nvY0lpwUq0EEVGeQVboB7PuHRZMs7yZpcTGrJWdLppj9p
OErNdEmqpWhrZlyP3C3tyb5GDu7ibcSbFmbt5/beZ4s1dTnZO87IAAWlFUb5Kzn2E9v3ist+CcVf
dKdwAkE1htrELuop50mq2zGfThG8vgFvg14vwu+gDKAdKsuFcAigl1wMFL3Ly+zxnzi+O93QA5gb
f1eVk81g2iJZSOhr411YVjccyY3y7edredZb8J1CFuGNLGvv/H7pt5bqVj+b7fKLZNgUVFP72tgz
PwckEgBpbTbfei+ClEXDIHN9Uc0jx/T68YqQaaBYpxwamDh/pWL8imhx6ouzgV5hPKtq59+E6oyM
CwccSDEGKCFOlQrMSJgKyURrp0hkUy3n30CVatkv9tm8Yyrymx9ESddDiTrXcolQ+lTpDxSukOAx
XGlB8ueKw+UCdOyI6LX8JGesOd5L6FHA7e4gTSCt5fe91fK0kVRhJ8bOAqjfT83I8NX6EaVxiYO0
4RuV4ZomTZBEl+/RmaZw/bJBDnld2YrqIbN5YmkHtpFOFvyjXT2pLATchVDPTmBHPTpokZMj69YH
S56xAVYyNkyOeiVXNIMlfbROCepz8SpvoGJRYHI7OBeG2SRmHa5Oo19LG/YkFR0p68SMc6XeHD9G
XMxTK1upyrCkJYuGig6MlGAN/Lj4rLgOpPrS0GYzulRiyk+dRREToMoV4Qh6Elq/+GycQXsyRH1A
z4xmoDqaSvzqiEi2hQMQ2o2gUDaUsoW5bilns10JKsopBfxr43AXoskIqrbJOw2L9aUfBWZt3X4T
1MMMDRl+OFf6AwScnxEEVP9rkTztTgh5fS1l/3cC06kCwDJtZ62CbxVychDs94gIAK5Co5sXNmNH
Qhzy4enba7+ZL7M+y1lGamfQqvRP6TmzEelLsIkpDiGU1wTfu+Ve0MSd5MVV15xtVZzIhqzHU8LH
v/r7mt7fugaQnPWDDOoXSIykE0k/oYDChm4z3moGh+bZWnuzYRJyjerG/gy35LuBaHtZQl34W3iH
TOoE2MWA6V8zOhP1m5eSWHEy3Io8ksfJ78H+5WHBWg+qDYM0FPp5zvUeMjIGT+0hqYD57j4iilzw
x+biLS711gyeOMVlCo0BRb0tAXIUhYZ7asp8wBEzIGQVN2Esh74ZjYKYOG4l08znpnJXszYo1tbp
gy0SEnQX0WwALYziuzdD47E39HiZSz77Imjf9F42GbjKXf255vjxVytdQWl3wmLVwwpQ9pPY7yGI
xrrg1pydvU6a+RYRErImXpdSlYUIvF38gXR9flTWof7vf+YLCrLKbebRboGdFP6nWC4XuDHxlWUA
2dukMJdyTf7K17d+A7Mbq/Dto5ip+EyM5FVrvkiDoyKQjuGn2hgxB3c/1MAD5axysqcBGLvaep8a
mVQqO3+RhQWfFwIYywDZu4E6iniGlWorC0yv4O2zSpWQJB3n+Ti4xtDEcGRH4dSKLdoOtiuHlVkY
xFy7kXBG9Box0G+OgmgUij3Zh8PRrkESLOL8Tqu8PyyHkRQ1hzGmWduHpoKnSiq6t7Nh2ht4TP3U
hGKmW7JU2XZ8mHdldod4KOOyA56XUPLY4a+ysOVakySIJpTyKx4brGl5lwEf9f7/LBguZJr+l1Tf
tR112LaHZtHq6UAIcDkVLEzNAnUHBPZ60rj3LdHnd+sgYDn4wQFwwkuHXGyHA67xqHq/9XvW3iTC
PipE1Al5mfpJPaWp87CPqc+/ovY1MlSSbZeyIdjQs3HwF/vrkH9dPe3Iiiepr4ZttlBHbYA5W6tm
HRpwO78yr1WEQVmrPGGHg5YhTbz68tBDA9W6Nytw7aOxawseBTMngQnZ/0zo3Fk4HbkHUqo6xonh
/w8mRO26o65EfQYt5GjMag6QEMeWCSA0kyprpnHW4kUdqxHlc8FZ3UeeYbkM4BpXbHvV96oMSIAW
VKbmPieClww5mzEThWw404SwM9jXsmSYa4VSHiZ/6eAdW/q3XYKX8Xwr8QZnDg8K2idi8UtZo810
GgXfYzfpEQ5NtcSGjntwFCDvog1lpK47uKuw4YzWK2/D/EqhACdWyI76QXHCr8B7wEeEG1UrQCto
u+YARarWFbYqpWH+WaHMPT74e6/HCnMY0KLZ9R74BlPDl/TD6XM7sBRBBYI1EoDDshHYI1jR89BJ
jxXrvA/+xndVdpjCJkTSxThjdNd9H1kakN3jo4YyymwQf+F5xtpkH3bxqYa8WV4iiYK4C4qqWfP/
rB06qlBVw8bed9DUVJnajZ++5whPapUdaAhhk9DFSKS4ShLcRtyPgj/VQVoM6QATrw6RdjRinrbG
iFrLdTsm3+E8HAM2fIOm5odVG/0i9/WWe8jOHA7GBxd8eSG3jfqsACfs2heUMuSfegBx3v/Ed1ty
MZ69w8cbtv6ERGdVnqPG9KsZJFdep2v1u8fuIkhfZQ98zYPdyQtpLp+DUAroZENJrhqdzX4mq9fE
EEwDWTcT7IBK/I5GqcJMU50GW//pWj84kQWbcULZwNlR0wIozBiKoRKIJFL9aa6vb6lLYA43WGzx
ZPosfErRXOAbcd21iT/JK/ecTVJX63P5Hwhab/0nSWULWEA0iPrczbQypZCqInkO3cHpDVkNWtb4
6td9d7fspHsQu9vngnsSfMpTT3jWevubLhC8Kopxg4l4DiSSG1vuaWVNn3NcG/a5/NgWPP7WWQMn
pweUuS7eSUJhPp3M6OPujhY+Jpia8LfC2vRARvhKEzjJv9YyrtJFALaREzvxEHxit4KiuevQHsM1
R+ytj+pmPwE3z3ZUAaMLsfpATzibPonTc5JHDpxx0Mh+XFtAU3xFRjw7A6P5E79xBQ+7qepP4LW2
xF2Z1qbpByDct3/mAIUoC60JmpqAMqQBgcrsBet+/QmdFhK+E7/pZrNiUJ+f6j8goEzdi2QZ5qaY
6gdc+7m4Ka/M/bG9GjzW6P6jHoqmZJuuTxTgd+D8IaC/RvXzBqq832KLJCNiii3Zt2gb7SuodZ21
iix6ImSkK8ft+VmJ7Hm5w+RFLejJJYoWP0JemUmsRlsQTDxjCfnSDplUwVjv9VcRSA0hsYCboXuU
qHs0zCipJlOllJ21LZFCcWAt94DWgPlvvvTpQsXXIK92JxIfkIcaZE/T4mFVvYDVm+YXDtJL3KN9
YTzaNbFTP6LWmF27B6sO18fTfnVqsoJ4MoPh0VCp8skobTvWWreoYccfL6v9DiKXAjqHbDRSDb/h
3RT31SA2+QKH55P9fAxQEY87rWgdjKz6KDpjtMO/P6CmYeYCRA8g7jyEbtgGUUp7I5LN24D5xD/4
Mhh0AxT5xfdpSqzguOTC4bCI/PX628rG6QZg7TKMnLmiFmYf+Dlxjm/azGVN+tYRlp/Kb4vQpqwu
k9jTZQYapjc6r831dlvQQXRXxlOF6yE8DwD6+wv0CL5Pf80DJaF1oOa1uHe4BBvvMg+8djhaJVOW
QydlXhqdqAaLclLazod4WKxQBPp+nDLhkL+/EzsptbmrFXVhHjbEIRen4z8XDdCQckAMmYhGPPTK
cmiYy3JUBuDvhhhf7Xbt5WB7U7wDXC8LV/yAmZc7TeHs6D2XC0765i9fR87pQiPFHNJh0hbwF5Jp
qWidDLYGqwwLCDJnLOTkXElnNtfMOh+hsXKoly85M2gi/5lRv47XSVwBe+peNLplTENPdd6x8rW4
9yKNm/93EjkcSPuUIpDaDfo3DYG+LgDhL3BioUuixGj53eofwwrOkk+7a3GC6TlxNSW5qQAglZmB
57WHnUjbpIVcf4gYVHSE7psjY8xMp6DHh0BNOsXDDPokGtsuBo2lulmnzCP1DyhC6WlF6Peixud9
LNWOUus8n0jpCM/cHhS8bz3kNCVVN3d+2C9JcNtCpTI60tMMQEebDvOzyznMIT6om19oLtArwnEj
zoMwXNELSeoHsinTq+tEGXb4qjd3UoztmBfC/MS+2lACw5yc4QcCght5xzC6giZCGpUPQx95cSBK
dgNDdrH5RzrWIR1uHnQbyQwfA2CAMupJtmmgXZmtUOpz1e7CzhfGwG+2vWlZ5s7ED0ivN98glQov
rGLdsGknES6aGqH9G5J3R/5pdn8ppcK2ugJCOcnNHPu/gPbFRtz8mX7eNZU2bAbWAfiVzNULSGq0
yFX5jKuJFIrKpcX5T2fVRuYdZkWZq2bgXlc8Z4AyJwAXy7e+7g2oSeZea9dIRhdIE8/lMb1Uy5QZ
rnRfg2SG9oqU2m9UqgucnEw7EYUs8GLNLxIOpCgej3bmyEX8VWQgQTQO7ChgmN4ceVVzTMHLneVx
idJSZRs1P3757hMCpw2piTAe6mAOhhb7hxvRCgxLUNwL2fy8Nz2KSLkX2AbcZVNbhQJI6J3Uq/Zt
ac3KND8NxLE5znuudhHG0dJA/lYZy1yyycV747QgM3i/U7IqtxIzF6s1FfA2IpUp0k//4ln/WjEu
Bu+oc3n1K7NxVL0SMD6+hR0SIDpBemcAyoVm/FmyRLZAHAW6yPOI8lmrTyy5OY5Ici3I3lemHxh5
ussPeAdzmxqvmZiUZz92D9XqrM9ErMfYP3ki3oeR6YDYf3XQXZxDbRWXgDJl4tSjlGTQpwr5DGli
g04W5W1vd61pL1hKgWj/cM45FkHwJuv4z2aBzebRZFdJCn8lEKU9Mj6kOYWM3hVYjh8uTW21FMCE
gZd01WgFos/rAOgZg79D2WkoC+bSyTkSXik+ALX3ERUOY3pP48371ldZTULxPOyL5eyBuOmF8ZtP
2sYTqJ+RKPrhJcEU45Q5LDGcqt1RqPoDppqgSAlm9f11MIRaZDmgGr2Z0WMEr6eG5JbWo/SDa/3n
EwA8xmznAI1mj1uKJHsI8qnwY3m6cHWvCAiX4b065rnjiFXAe/0W0JvFcaXl3ojKOAYWcHCmhsGc
udjn2SCI1dNNIh1jHSGfAYHBXG+zhQTF6PCAbkUqOz4bAtMcpwrOn+etvR9rvHyVxrzD/yQPOKgl
K/D7vHkU23ndnMA6EMgbzEV4hks2dqXbeq5qk4h95CLr3S3yD/UYULqdrm+wgd3ufDaNIW13xhOa
qvfLAbBEp9cL/bp/KoCkVi4V3t+OVLgZmqWBp9doUIc23KDDwSsv7qgkdnlmMzfwdy40SF5Yp7br
LQOV5m5MhweA48QUTdQ7uJBvXlPmPK/It46t6poRFSaovxFm1FhUGy3ls4ibco5Ay5CYj9vMXKZn
+v9zmvAU/Xum+j9K+yQmdHtScZNrUYApV95frIeAkP9CPBVfrLZg2B7maJJvr8JWxKb8M0ld1ajx
edhwkuZYAheXZWBTqhPntdgMMb1B3V6mFw1+R4DaXfCzHVZ/U/F/x1PCTxcexkf/9+nl23ch8Ky4
cz7CDot98brmuCLdk5puwtZEsrFf+tGad0q9ZH2PP1gXL0i9rowwvWy8bHE1IOkoxFUW7ng91wXQ
XTssLXHSlPocXwEDg4UkWdq+cYk5P97fpv/nq8W83id02eRuNQzoglTVkkIRdDZbkJxm5bT+oPIf
B2F6bnXJuZeQJ9wdXX4uY/nxqmN2lXUBOOHTZ0HOJohbXOLDnncvrYvyekDo+OrOISUd7q0WRik1
aZVv3mTMk4/tOWM7Gq/6TG4hiDrDJzXURVXYXO4ieZp2LV7eezUhjwyhZ7pD4oQm4YmPrg/E5J05
W8C7SUjhvKSeLF7sRlcNq8B4l2IOgTyGMQq+gRBzUB5e6O4FwQ+nqLXM/jGjBDu8Qt4IGNaPgjHI
bCIITizAKoLbpzf0Ts2Mv/2AyskphWk1upg484E44Qvj93YEijxwk2952T0mRwINGLzG1n55dNiK
S+5f950ew442+hBRX7SuPlkAXYYrI5s8vs3yXW5nvSNXz+anpVMdNRPDFOr48cfaZlWsbw53oAuC
Ip7jYK5UcBSVGKfkGKRUGjSI+UUKRIkLU3pRGaBw9r86+fGOY896AsO+EI3DpVp7bZ29dlgGpYGu
p1CGNjnVUjeocmzqQniX4GUa5NO1FlvqySvsEcektzNCYziY1qhgmaaUOtpoNG8CeHx9iTNu/t7H
A4JmUYYkdcrrSC8ok/HXXWg6Gbw9bqcIrk2GHszIiT/07CwMy9viQHHpDD1VYMdiAHJbgIbbh1jy
2J+aGNJjgSMeZ5KCcUONYDpAcyjYoPjk/Tj/8v4eekn6OGcUYJgGcpvjhtTZAndquGmMrf5K5aAl
I8FgS34/cgptpTAF9EaV27bKxLWA7rjrySFvZoC2+Lj/c0iTIPsyLDsmUCyuIZkB9PKDzVYfoNVa
shidzcPH490EPRfZGhaKMCb6EqHFMOvdWK8i1nosSufuX3iSoJXnO5zmDdKliPBRSQA4DmBsRvMU
67RUrBMx49qDflLtDPlYMyiiVGdPDQ7tcIe4EqpHBsrOQ4gW9kkani2i2HH5nsGvd0WL4QUb0VPB
4hQXd4aKpqIY4vTzJIm95gnGBGZJi694VSvLWaYpxUT0FRV6NSz782IcJFdrQP9JZZU4N7R0Ithg
fvlxZos4WN4ncTaIfOtgUTM98611FTOy9ELPVGZrb/kQ6d5uIw4WuCTOrAn8158PCh5CRwhFeR/Q
D8F2R3MMUbgY8sfTShlxe/uWMFSZIGSUjJfIKm1N4b2Pzyfr2x7CdiWOL5jGplLzLEovi25yPSda
kH5EOImBTM0bXyOJaR34XODjK3OML8YXWEvDUR/zTXG6pAsEXR2iCXDS2B40WAJqLYPKuRvBESdt
qSz1DG1WEKa6KHRZZHSU2zF9Xpsh86TkiVGqlgVZ9qoQWP2VOV8I01VHoiQRGcafoDrC2UNj9A5s
hDodin+2Z5MSicFFZTwR6Ft9vRu2pxpFEnQXLhWMImQf9leXY67k86oGRtlG8P2cgsUxbg+YfdAG
xyGyslkQ8N7bNB4B3aok+TDjKFLHfLx44EtN5BWYm/fORpXmYsCGU7gEztMl0k1K/v0LsDfiQ5id
GsJOBVATHlsaB17/9+VhY34OlDRytOQyjZoxwvlZYYpgPOZwR3Wzwq6PNPZ0dimdDKWroWaXhF3i
UzYm3n3l5l1mDBnjCWfDb2b74n7rKzbNGTzg2QB2Z80NRS3ZVzECgYsl4XA8Q9VGA/81Jr/ab8HR
TOxQ6NMN09wuIaSSdBd8PExVaLlELD/7ToAtlttE4+hk66dhpqvxLxyXRX0g/nVa8662galCbyI8
OX2z/v0aT2PLyYZxorqKa9j8ATwrFh9PQUuwqvdk0G+ptXwMZI2kSP7mfb+0z4EwU3jcXdY0FddG
ZvCV6zL7G9g8wMf6JdaSNaolpdtWPTuJcfE3axhgeKrOcMhWuGwFR+epR6ip7rD6w0cNtFXnj1Uw
7qrzZzM6ECmgFthXa6ThqeXl1icoeSv/ki2dsIkXSq+esQKerZs800xeytdOHXCU6n/BujrvW/Wa
BZhnyg5y77tVHhVA/BgPilUEQi63LMeb9q1RHLmwbRrWTaPHPabPNYCNqk+u5hm/C9VRAXtLppEc
OFRg7Nmia0Al/40SSzPr8c8duTuB5TuOKZXhVTYBpD9CbjiKtLo4it6Dgc4BwyDZJYwo9bgGxkMK
txbui2r+LJbRVVilu7fRzJp1Qh7u8ABZbk/ddrU7cUe4n6CkRUNNJShC1UDDKCCYvqgzojI5L+D6
PlCO08r6wlrf5MUUUFTuAPQ222KrJLP3mrjoM7Jwx5Mtm01zUeScsF+Gym8tDu9t81hSHX68o/68
DGA8XecWltMNVSU8QbyH6lCxgLGoY7Fwpa4SW57eMMeXST6iHss74gl1VMhf7Ket0hBMHD+u52PA
/LSopVUQEW2+QntAw7635yaWtSS+ctzSFZiSNPcmgf4tiByqBzw581my+DDecIUKOF+A/TsIRAOm
Cr5w+aY1GzFYcRdW8B8FbfSu5nfkGM7VAWd2ID8tywA3B04wqRfUEquhzz7s90DByqq7NMx1GdQ5
sNurRYWS5ceUcRhVgyOqFGN+8qWdFk1++yPluzwjOeJcyCL943MxGSPGYBPyGOp+BOTFe4QF6+Lb
VAyG35YTEYTz6Kq8nh7lsMj+GBHWCBC5M86TIO9u5AJ7asTraId0oNF6j1pF2viOWLh1n/Y2mFn8
NqlEdclapWor1Z4RvR/j4ii3URdP2w9sIrIkpuwJRMR4B8ZlhLARfdDB/GdJdUyxblJawpesMTnN
zoGOMhQJO6EQSRX4azAw63fUFCY/iEgDrC/cRRoQZzCb1qt3ruIYvgpsi0JJb9VQeDYnk3e7wUl2
IIMyn4jpVq0xydwlAVrDQKft2Iop6rXd9vSyK0tlze4fckNsFaSUnRfikXZSr+/tDgtDwqXPLLMc
0+SSzCdNHO226l9ZByyvOcAlc6/penhdhpihrSoWN9JwcQk7HSiGO3UA5YujXHpjry4C9jy8JvQG
MCDeNYK6TiFnV/2I5bvOmUUdDTFRVWrGi8r/PFVcL4ZXZzS/Ey6xPLfyW+b2FrX740Qv2uYM1BYg
sNEdm2WosZaiXoMcq7eYyqSpLktoyhD6nWWO5a2HZv4XnWeVdxRnSKgTF04bC0mQ95Zgss2zrOo3
B3GqwTmnH17yZx6/8lNzWTtWka3RqyUzPvdRkLovott9zKKGAPe0iKXOPQz5kiCYtdHyJ848jHpe
+jD2T3ShFjt82KLbaw43RGRnfyqSmWldXiV64IX/1LanTebNMcCB5M3w5YQWGGZIbyt4FHC+2wg3
fj6xBztwMUqcBzPdG9p/YiBH7BmDt7F/NqtUJATCgrAh2wpzW/nGBP+2btdVsN9JX+UaDLjBLZuW
KKfyLUlxXv86hpCRWLSsAuYCmnGznWSzZ0jusf+gj0obNw7YkiHnviN5Lvig0QF7NgEvSzvKR4As
luisHUijFiK9nWqiXYFcrg3ugONCbtd/HcfQgD98VuFvleQlS4fL6FBVWSHx0aifnnuN3l6MBcT9
7tzlKTn9m78ckT/WCNGqFGoAK0hyHaZJGP+m4HlHDcncx/2s2HNpqtkjD73IyNBWYKVXJMVZ4mfb
7uuTHuv3wwPaBy9IDwTxazkPqwZlmNkLW12SKEGIL2UVSmNaJe+7UFqUOsebGGuN95gX9Jcdm/HG
7jciCB6pfwk2rh0aQuZKYSvG9sn8HPYZnLsKR++teAqjs5oITA42MD58H0NOoEjrbGaxtZN9IYA4
au89tJQngaM1MRmNGHalATtXF86UZavp1yPqJxWKbPxAlFI6+Qq0s+5HXNNp1gVGPzl7zIB5IZ2g
C1Ot5Dv16e3ShokZwh3YCEHuMncqNC2LrzkTzLMYAx9s0843XVwJfqoW3VmIrpG3Tgcqk0N74pbe
EHpTa6zoSI4e2abPVXAwkhBnsqiTSwHooFUMXEj3eJe8LaXN6LKWkrg2WeyjvRg3q4i1RKopjCX5
UwaWXV8F/ZgYF+rfx6FHBCTf3LOjWcy9JexSTa3nUKDbzI3dcOe2fbIdXfVAqVxLf5JCkEtlt3iM
gNxt+j8725uYM+tvYLwe0phEsG11tHnqThXPfnqYiCn3Eruu6cdsMXEckDBmqGCHW+TA4G52HSdK
2ecYRX38hhc5+bWtybCFvTD7t9Ru/bRdyi0w5S9eD/s23EhVFmH7mBcI5GWC0fDrxwtfQ90V47Rc
6z0X20mrXozZ7pvIryKkTN5j5k6AWkYfuCoWj83tsDxmsN7wFNs3o/rTGImo8I4XjoV7iaRMv5bz
YpkymJ47XeyF84Lsmijv2kar3p56XebVeQFiho5PjgoQXzI9zFDNE8jvTqnUhE1XPGRaNmoWGYVl
nd21q0tWdCCXLX+9bPlbbQOOHz4t7zqetlS141AdNaA9UdTYD//CRum3lKvo7HSUsX4Kpkh7Biuo
sWrf4DupbNzRsL9xN7nVdwK4KP41LZZBqfg7F+mB0ZF6hskAtH2UtjszAscrddbhVnhCVrnV9E4L
bXna5IgUHzShuknE/LNDBZJ2/Ex36Q9n31yZN/N7JiY6h/8iZ94zH/QDc+fENfVcMIYU3tHwfIqE
BAl6l7ivG7RdnD43v+oopeSLxVt10MRLlyTWCzHCp/rzCQ0d6TgxoB9PoLpa39P565JD2Esw0Ekx
wpna7w5uNG56A6NpDlylHzX2Wcm58G7AlpbqPg0N7tW+J5pdpJOMXIOUKtUFk2pYkixEVHNiFqgi
Co9u+1bPWoXG+dz0iTg7vTaR2OBzG35tn1JcYakaQOtQqwqiWOeZcZ1jJxQjHBGe9yjIWA+z33Ws
x2Zx0m7W2qwbOTPEx9tmRmXCVcYdqc5JXP5wrfiUl0vyti38ZU7c2LehKcUHkwAhQDlg4R53CTgz
wVqk1hsYMx878ozeyRt4zPXsvzr3gvT5e6O2VpvZEGHf4kfvbragIlsw7BgG3W/KK5VTaHJHtSF/
Ltz3CrFGJQVhuvZZOicNKpLmDpPjMS6Gz+gBPY9P9cxCFKMFK8xXLHskkdBs3q8HO7XDW1Z3bnvn
OfYcUaCgFR+5Po3igQOxjEfqJTwu8XNg1fVhkqIfi2jP+6iTBLUZdvuXCmQV9t7jw3TqeV/rQdJl
2a1ZljeR206EkFXmRKuA6ilc2PxFM5o1UPr2QxecANgYp4wso6Jjak1v8gJoDF0iFqrzNqHzTID3
nHU4ipYL4xnLMJTvEtFez8CryggVY8YDqstJ0m87yWzg3k3W4LU8B+QNV6KcJGQXtGnerqVS72kK
dopNRXIBQxKZeEO2rYt+KXsueuAFV8QGnx+DV0fylwz0HV1LPjOXTbGgR9l/br/34LJpN2GdNOLL
f7MVEkbrOUbkHvwpDlZBa4C9gTLIywoG4Z69jYnmtO+7mdP9U1kRKJFc2ZZuv8BT+gwcieLJoCTc
NlGc0X8VxtU9Ji1SJhB595TeCyzl+fXqePPX7spGISZEAWs4C6Y3OQlk0/6LWC05wrZTtXkxgN56
pjxHnK/nO8M12PGbzUXXppA2pnrNQ0S32G1lX81BazS/NHec0BeI/N2jE9CCvdCQ5/g5W89FOZzk
ZpduiDgE58MXBYhmwTk/AchugGufI/RdO9wYnSJiIBPSXjZPxlt/TQLUknIHtYyLPTTmluYwx/su
ImWTnjwdScsVIcuNcJncRL1AJBIloISCf6yCORkx1jtFkHuDX/Wr+OwkKsNWa8tDYWqdvUoqQoAj
W9r5KAA1iJ8XrJDGfsonQqffMH80dX8w95/R3lGVWNJX8Aa43Iequ1UJQzI+/5mSoJbXrywnS1Hi
B8moLfRwYHTcdmUDJLJE1Klu+Q9zGTKjtjKGHUSppUxGByFuzkCLOE9U0L7sHMdSdx1vF6ImhqZv
+CnbCy0ucjJCHjHYZ7sxRQ//N45DHclZdPMj8RR87Z0maqP7iZcWDa4TrxUtd6b68iqn2ip1O7CH
9ZVgPNfDOINm7nbAo3Ud4rKGg7xyQr3MSGviIJHXjiKolyjVcn8GYymZVlZxSMK/LL2lgbTVb6NO
vgGHb3DFwzNmsXoA6tGUpY2vR4WCJw4+a4UpZt+Usgn8a/BgVnXSUuVVq/kQw2PGU3xuv+G6ALrD
5MFDqW9D0Fe2r4dyqRyCQEj+yz2sYkZWr20iIK6GQdLcbxu8d6bXbLKzlJqq8obSYAhVWu7NSulH
zjwxIZBshs4REWSDSzxvSq3OrP9Qf1sKIaniwRNPxU8Hycca3veql1VF0i61FBDl/kTs5tqdjQC9
QPaZye195Q3qbP62FRqv84frkTkKBGfvG9kh2ixeVmSZ1t9EgKrZSELGrvM7A2GgWEyv3UaIHl/L
D9Zc3e6s2M4w5YiW1ZnyTuCLRLzCMFMPJCQyGML538vRE9ho9J3MZM9Lq0U50phBcDLPF6Nq9SG0
xqFrseRhujNaQLMBAHuQpB6dKFm6zacQ6CuRjlGgY0LpURejJOWlQkGg5kwO938c5Nz+FAYkFq9G
eg3UfMPW0+Yxhck8qKFAsvXJHPo0C19TqrLaYXGc5rrF0fJ6w/ekSAoX+/ekK02TESO8ElblIm+H
q2gSsC854u07X6By3780KklMUOL92SFVEZZCwOYqJ2KDLetr0daz0uX9EbOcYdJBoSfTrF6OhADj
vdCCPoVe+eWuwpv5bWV1KoAPtomSbpEhnvoI/wootK1uHoMn2oaBNnEc7AE/ycUx4uhrQLHQL/yA
nkIt56Nn/9fqTosA6e6PyNVX5ayQB7cXdelw6IpUdiE9VV8Kn4GxRXcoCbpG5Kd8jqET2bd86hJB
PySogYOM8v7PeY9ScBgppoEksS6fhwd2VaYG6s1MpckD88rC43TNZxwLdcYJ55Sos9MjQ5HFTdkg
/ngAW02hY0Tx3z391wYC90A6yoNrmIdSiQBPBZSbS8zRS3TZLhOIBm0mQRD4w9v120pEdZoFXFKs
sgfCyZl3JgH7EOKRcLpLKtcRMyqg7FBVebcKibbOe72vO58Xqx6OpSIGbQVVRUEtnuiQyR67PGCO
ycmhGeYcp/oKo6nj/YOTICetJGBR5Ap3gvAfw7ry2wrybFdR3GsBAADVR1pVj8d0rmu92zbUNyTz
Wcx10Hz2Cj9CQvDsgxaBwa+hQQ4zj0EvlKnAGZZVZSWNpkR1DGUpq8t+C9LmP8WzbBA0WS47AVwh
E6daIhPq7OYVuTK83xmSDLWaL5V9fzS+ZNRjuvVFUHfJiFLLqNVBzc8VRqs1S3FFhUNyI1ZgIxhd
/0tJmIwpOTVPBCXNT0J9Aa7oIDvLV2ri78DLq3LCQNLlviOpkWFZQYrHtHAW/FavpEx//NRiKHGz
fzlcwfvfjubJSXT8wUE4LWoxNRFBOx27oADTL3h4KWax8uHhN8k+JrivTEj1CeTg+mg0pKRLS0Hy
if4ZDjONs+WR5AyHJND3Pl8crCR8bMjgW3q7kCOqOuJuRbtINniC2zO5KsU6705Q5q5Rin9VU5/7
gSakai19FN7lXOiFZbkd4V6epuBmec1Pa3496RyCYYVWlusXZwOif6NJzGaAwrJVrN7Bq1VjuMkT
V6V9yWTUKNPULhcaTToxeCMiAlfdZH1iNCL3wx7+xXxpd4UEp0YG9my8e8FijvDf2WEoe2ePvmVc
jZ4wE7M0L0LDzfZJQRXsUd9UqmZOQ7AXq0zuEg7GpuOEJnXL9hBNB2w744W0Wy4m4D0jPib91Aqv
PSNGSCUOxC3kp+IOVdT1kHVPLGZSiqGELlzo6BqUrXHm1cx3Pl2R+YUcfN+T6TSgh63/23azLEJc
bz2QXTYMavhUo3oBmKNazT8S4+xv/eierZNksuiNuYqpW4Z3ydKGAf+itaJmeadSJjrFkUR9YrOS
0Jq6FknvbsOT+6gZCkaRZFQ+E4qO/UhpRCO/WM6e4pgRqND/QXv3yhK6H0cajpueKQwuWtsT4ZLz
cJYro7YblXuJqZk4bT3JGxEZGjfgtNd1BSyDwadbb10ib5H8Yq8SHjJLjAhmtZ7KIK995S/VPjgS
7NyCCGPFaoD+2sMfr71GBCPLwgC3E5OGHTPKNb3zmSZXE6MRiRd4WApc99GzeZEZxxWWzhkPhUP5
Hwei/IcQdAo5KZRWrFgLjskrxDmLyTC06N36AGZDqlPEJDjAS91RFEonKGAyJZzFdb2ZxqQxicsh
JTGaqmBMx1toTzNdwBHGsfW+xaN64VkQH3yJBp7GTzUnO7SSDzYx5tBjeJhskDNMvjWSn4p5hCqa
IBw7HfmP6aX38AZPkJ6H3/xw4e/vLW9XRCw8QW6nDnlr0Ky0sakX/J71228hMstb3zLjTodZwq50
fgRW7SXUafmX8BlA0kavhiKFz25ZBYjB7cNARuUbNyfbimHI5TxF25dT44RSZk/2qXyjCxA+cjq4
NELbhfBHkFWBvxjyjKZkmM+mlLnsJi6yb4K9ccAJ+S2we48KSds3bacR1zDi9Qt3BJQxHYpEF1Fy
FGj5XZP9bfoA2TQPcdQ+SYfrgzGUUShR3DRlY6v5fon23CprM8l1FzHALwRyoTueO5mtoAR2kozX
XjjGuBQXTWQXiRvExQBNL5bgy3XMkbMHxi5nRoYzI22Ejz+rIM5hLFN8KO0Kv2Io23tkomjWM+8y
13cmFWHiUKTpid2W11iqY+YPhqvy3Zggq0z3Mp3zh+JWODIztvD6cgAlCbH15xqIj+iIIg6Amqs6
fcR863GuaCkMQTWBl0CUf8+nopoRYh3Yo82rGGplXN+Dw/R/LtoSG3IazSTbnE3lTxNXIM4X457b
oWdfoMr+O+HxwKZ25V5pfkWpOk3cihRX+yP5Ug33IPXqoXmU+yFg+dTmoqjbKy5pgO59BGRGikq8
EGSe0+KWC1bBi7AL7BOLiBKTDPSk6d4IjvWR1guHI+JKe7dYZq7PbfwiKtzkSw0+0NU22vqt7+1U
130wheecmriy1DbeJlr4Qx85CBdxf/M5M9l4UvwLSFhTJ5xgfa1LKToP9eqZAszfl0cOi5+LufgJ
/NTK17NR0+/+wwpwY3kXh5rI93Gvf2PLN6tQfJ1DTbFdLmgnG0Nqibrj6XMSf0SRIvVdMdAIh59Z
DeRWWUJyM+hAtzrlNP8Pjv7wiA2vU11TTJFFX9ZSAb//evQlLnquliY1ssSbVSXybz235W8erNCa
HcPnsh2xTv5tjGahSGm/DMHQCvKH2FVI1yT5ft5I9w0CBVV9hJ6/XKLzxzP+qWzOZJO2ZpOXo8v+
6lcZas3eBCRb2SB6tM6nzh+J7Iu3ufjFBtg3haPIBF+XhmKtCpPNftKtdxtPEd6WkZYj2sGYmBoz
45IBVmmE0WRZgmtscn3BIuKiWH3P7CLFPOAQ4n4SpReg3PNvVrJNgcmG5qe4slOWai5572Cxyrhg
d0afTY9M6EOqPCeWuRl57PgO8U369+n+jOg3GeK9ux3A8CxQ66Rzsq8nQ1+oLYWeqAw4yHkgNMpu
pfe5sEmt/9eFZFG+kkRAG8kV/F2g+kOFTKnG2deIdZJ+fmdxwLY7KW+LG0nbwvE9vekFCFxielAv
rbhl54oMu6b3jmDxtbq/9O8mRZBxin6O2aV28JZ4RD9jjGi1yTIN1jEouv0ahgqqmvUjYtvW4L5f
srKqjSUGDxR384dSfoc9XheNmVD+kuteSIKb8ky3IR0t8ss+pTduddtEYH464nRgwSPzu/rWYaBg
tYkYKeq1oDY+LHLS+N7S1LYMoL3se6GlX2IjHpoPcbcVRJtXNYlHHxdKZWu7uTuSxL7Bi1hAtCAl
kcyXBRYR8SLgoWDRKJqcu1OepfqLRYIfvYrQwsqryp/cuCxng+sdczEbpTBBljfeM+cXSjlqfzSY
4/cYzS8L1HeGkil+qNHGl8yHtstW81H7wo594s9ndbZuiamSzJ0nMrMote9zFoFy8Wm9COTRDdO+
yhJnJojUQxgo7bg/3FYpnrXC/+XB5JCVBPLrFs9v+oY0AuajmAhRP/g44aSUBlBkcnUjfLWoexbD
bFO2AZBXVuqEYhi2/cEsKyPteosNtbxu2+6qyICalz6VrHZjinO1PeNEz/S0OFKH04Hh6seQfBwT
t9QolsinG+FGHKqHjK1wwBOSwAalLFcktzE1c77rv14bKEOEffiABOhQZOhiJ79eCtIkznlJWjzg
W9+fmSkPzPZ59tF5xzPlzpbXnK4LNKggVO/o4+RZp1o0nQhGgbf5Br+uRv+Lxhq4kxocvFQ1TYLB
mYVEml8EstuCGUJiZEp8am4XNDwnYr4u9fMWoCdjZNg2NCjdjulBkPpyRzJ4eqDNyH1tox52TlU0
puKJ0sYHqIbPdWcSE7qRCJcIQp07EkWSrgf3oGYiPTQ+k9mDNGrUWYbln497dIzVmoj5Z3ICN7Ja
ztxInE7jO+JO48lgj6ViosaDgdp8vOEVKkW6u+fol7soLWFXKE8y4goghGfkdtH0t/G4vYrc/SEb
d2l5KZwoZ7+1z5rfUGdY7Paf45kVVSdavjaw04mzwZ6ezJpipLNv9eI1cBnq+/jqSfzvarEleC5a
PNTeEn0VRktjnhOXtW5dyDRFNHmMbBCeIaRx3IBDJwioikU5ns+WNZ17iIyxyqKsXM4ZgxPcNALJ
YA1XGAnBF5iNadnaa0udKQPrUn8N4+8ppf0zKBCPQ6vGC+od3rNCr6Uz0tVyVx/YKT4689hc3it4
Ic06DeTvpsmdnpgNgHJ2jnndscJSg1QGNSMgb18P2SsrWvN67dOWj7tvJcLDVvX9S2cimbbQ3yua
9RRFvmK1Lr6K37T680CyI0MS+sTvPM5s/A1luTtndT8qaS68z+Ge3cdgxZgx1kGTW2aqHMYhQiCV
1XcJnhIgNIrw7G8QRkCYSUFt9y/ciivBdBNFSBEvONuy0q5lxaIZVHGrntmS8lz8ep9iuP826QUE
gPEZ72aVF2Ew6VlpRYNd1L8jfiERYrDr0TXTTdtdhFAbjw/vwD/0vmpEXZCCNC9YAM5o/k70ocrR
ssx67O5nw6g/KzhPrm0aGI4HTimOB7G6+HJpvMVNL2tWsQj4FNFqBockLZgauNC25a9Yv3ybpROn
GcsZm91su1WbA5UqEsC9qXEDWEcqApcQS3w6rFwA1s0fZzVVyYve3j0bLQ2VmIzYcWkpY/75G/uR
w40j8zV4MFhFGqBBi0NR2tY9TuTozcc8ge9Fr7DxQMYi0AvKsN7rEzorjsZNz6xpFdrCMaOi6fAg
Qw3p4DJlrMW+XU8ob0qvER2tIjtCR/CAeZx39CA/RkUmdoTEFVEQ86XoxYYp3PDxgVHLenelM4ZT
snyejRdK/OYUDVQk8EIqIFijx3hS8uRxMkmik69bj9FN3raVX9r+2FvAqzlpaa4L6mAhthBptZlS
hc1MblaNVaGrP14RA80Zukb4u+YbtEjQ7VA2agsuhd1NmAqRoytcFUMwkjun8OVxKTIeuf9ia41v
Dq8ilP94CyMS2EIduWNyFxWzTHmgrxaQbNs0HpfYk04qD2+LLEoymWbHbHFlcsPW5BsyQzwknZdD
WZ5euEy2oWkUbdlK2iPHygvc+1NlVaeSNCpm3kewv7JQhVnKH0o/bTrb1FYwtS/1pQQN0lr7UQjS
OKAy1mMFC351XvGnBOb9DS8Vv8CvwbdCsmbgQIFMeDqzhztdrRyDsswyBgk9fBY/BsoFYxuwwfbp
5aaAVtLEmumr0wzIsTjZ02pqDQltF37DYQTnosG/Msn/KfWsjQxA6mRt9WEZfcWBz33eTExAj4Pu
Rl3uSG6qnEc8Im3OZqPr9SzKEPTqjOeOinZL7C69WWxHws5KT13fSaXK4vzgopBlzKFFWxzo4ebC
PwAFjwe9X2TcwLBrdheMzP0CphBxRaft6ili6/h7H762/0ThdP68faoh3ZU2vP5UUd1Bcdz2C61E
vUpkEV3IFLIBDza3WXE9kQABBkIg5O+shZRbNc+aKvTvcn9SP62N6BwpOCmogSoPFSO2RtosnSEm
c6wsdvMRZr7Cfb6nccTVY6CiaofjW0V4rBAJRhfO/fy7B1jh6gID/bZR0T56kyjO+BF5MeF9xsdo
oglTv3edg2B4QTJ6l9mmMftvD40jKMgOP9HeIWhQC8v79synU0ileu3bb8TgiQDPGaksfacfXoW8
GB/ViMnQGxQXF9XJ2JhpNTGJeTIm3ElxpDQQ9OQ6nKXACDLourWw5dAw6GZBUzqLcRvNCPzwfxHC
LyOrXbCG6mmRBusmLDGcZdGk8by5W1n4CD4HzZNEJOElvAd+sM03fYX463AqpBG7QpRZXXf/8YSs
lirtpaqKTeFrZ/suiebazH3O53hKoBn5CVyz0lZP9aZIIvDQB6Qj4DcyJjwTyKGOPyitneWQUVPG
m4T80vRDsodGSp+jdHNhUvTqZ3VYT8hTYB+nUPCoF1NiM9WkwDA6iSqPCrEGUqLrRh1UnzFNhMpJ
7kvCdEmfjTvs1umgz4lcFZE6ds/M4vBPO01fqqJa8ba8B4PjlPvq5UnmXyVYDy/2Ec9CZL5+YeZb
TbK7I5qpHHSkpVdD2nGLMpj+i72DOmEbIultJzlAzKAqFXafUbsIXPlcmekyQQKNyqVyQazJMGs8
JPNNh2kWGOxgimdmYy3Gt6BUNREessrfcG+k2YuQEUf6qdkfuEsbozEzID5aYcHStdQk4OUf4dog
em1113L7/FB8Ai4F8xrPaah2eDp5F8O3AnhrVoCYUx1FJK6ftjG6jPWfiiQCPwbSIfo48BsPG87q
U4ypbxRG+kKGex2fWiP5+KhQlB4pYMETFS4eWW4yvH8SXSBY9oFvuIdFOpjg83pMelE6KnPoyo6f
Jb+ZfAX61/DTFfzCY7181HHz9PBXPFOjOPboSN3O37g4ATwg2HL0qjYfqLnqoOhQlZBAE0rZCdMc
1L+b5Sl5JBkyEDG9o+mD2+ESXRa24HTeHiJVvW4YzTWKQ0dJcYgtXhDP6S1zVHVaJp/81hJPlvv7
vFgXCq/5ykrLxygl1roRb3cbnD5VLPpJEXHPWqtagS0BzUzPgpz/qwPxonph3mlzm9E4p4IE3Mv+
+9E0v/vUQM346gr5ArcDWKdkeBZVJEe1+6cRmGe/J4CauwUxsgcCdceBmIKAyYk47u7VpEmd5KgP
y9+1W0jrMGFGXrt6+2vMLgqvE4AAmTBCN0/ivgX5YPM2Y+7xa14Rj0GCc2vMAMmOpx4zgAnS6OMB
h7CXVnimpVpYHMqWtEuT4q7ksxWzYyBzyCEBQzB7m10SiyDO5psKPZ1ETEPHNpT0copVgH5ryrIl
m2KOJYafAfUtVzHNC3FP3nhexfX0XkljsL3uI3833X4KrHnQXmhW35g0YApzjNqZkWTD0g4qdTIk
j0EW0GzrVpXoqSM8ax5H6uym4iiyCf/299MdqMr1E5abf7blH5ybCRzzbcsYypXNRi12VSVhfPLH
ovTrXUrcllAOP0JNciPd8YPhvpIF2nIgjzaRJLCE+xFbBooRXCDRLduCNmWcuRAzKtuXuX/SCtWH
rY39c3a4RvY9pKlmCOqI6dUZs60xUj/D2sIL29LeHe7MxWtRiY7FrXG5IvK8bGnL4XOd7COl9JMi
4XAULQV1EdoQ7q4u404FhopEGuvhCxyjl35WmMSWANG9aiFzyma+1PlrgWHGNGN/Wbkuemnk7lUh
symLVaosfy5XkeyEDfozb1aWwTwYA60Q6dlYBQbjcHYpFqLtecSIhtmPyf0DL6uNw9QXAwXLTlzb
Mx0oIf1xuBo8M2ns0p8NN5AwIWScKkc/lnCpGCT6quvMEL4p5GzXD08yr4FrzuDdFSvqtRtya9yi
6CdyAI1+udab4nO1uR3wxshIN+V01uRdbltrn+ga6JtWXMAqldoVlLrVLVmgQTueJzAw8zhB/ltT
R6j3lmWZhfol6OCxUpQspSRUpSCizUjM7P7thRWIQeky0FByfZwFuQ9z/BUvTrK7gAD+y+4kpf3I
S4w83hMV7qmIl/JS8wvxZGGmima9fIfm+HGu50+GVuLZshQNQe51VPYECzmTTQXQ3U9wmcVFnVdx
XEpNaPldFb9eG3Rrukz0YuAm+r6tIkCFNhNeBN53kxEA4RudTs2P//Q27c8bvgwnneQN+9+Hynnq
LmNcylou2JXtMfj0IBT/j21JsqLVF/ls0u8dx10AT5544O300dNWgGIrmMKR9wANv4rwIC75DOaZ
M0dGW5fjGSkgn0TH2QjTK9Fo8L/YM9Rlgv7Ro5GQzWaazxfGT/FIYHns9M93eIqKq1zIxjlPRx+6
VOkBBHa1a4pc21aZ/55PyebwEPIZPBOtRDkHVXn0My+qZNC7Bh0XH4eGBFOMbHMB6uwAHK+W6EJQ
F9cREzWg+nmRDYVvmocF4WpwiRnMLG+DhSpnasuQzxkg+Ndwj6mSRlVaNFN8SA6GUehAdT9zQmca
8+dCTCGkADDNhwPimgFNrXVvP5KFSFgtTdQMSQBkYRUGHX7grBY3BK7lvhqexUnMk5YuxBLbVB0F
52RuAZi1/80YELf9gs1+swR10SAYiPs3Zdjeq8LXbLxx441Ycv/pxRlCA0M0EJZqm0XqN251B6tH
TD6t4rAy1AHu3ApuqNRnLw+rw1UNDFaIv5bQd/aMwV0k0BB14KQp1D/4S8Dv1SqoHg5Koucw6dRW
wlzbnSI+xPT2YGgHAf68rq6CBudmpaogn4y701vaAvsbcijeDvhEYLjgsmxJSp4bobzxvvNZoEIZ
vNjFUS9dh/XDJ7GkbC9upuLAc9acZCFEAYB68mTp+LFxyTePHOVrB3OUuzYS1FlvI7MuSEsg5ylj
opZojbIh93CesQv839dQPxyharM0OmKWdHRHw9zTpwG9DHPuilCMEM4ZCkAM/kSCMsxhJX7vG5IY
+Kk3l2N/zUzJzz8S1T6jPIdB4Y19nCTSjJ/oLk4Q45fQTX17zO4UrbN37f1GSmRwO5vG457BKOFq
beVvLwe3YTqwM85n9gZkSjZ1YS8gNMzeXuCdB8jp9jmLz47Kig/HpvG6XcNUU+GzfHDCfXVk5XIt
z+ZaU916bwgvS881L8B8hNR20DW/1YEnABejTrxrZtfZlG+rs0u0gljXvS7mXvJg68JtBqKEejv5
4r6jgFDc8181pqXho5mSrDgIMZnkLrrUon44rGlGmwOL7XkIPqNECR8z0id17CgxncCw5zGT3mrV
tCJfnlP+2UbfSJhuLih7GWsa7sFzPh1MADwXx2NyARcgNvztyFLQQoi1sm6AUW4L7PJD40SFbAN3
OHn1/GYTNJa1rbnq5oE02nhELRvtFRo+FAR44zDzY3kEx99VZPBIppET+8CO6zIWEFWiZ5lICnSJ
02PDLP6wWHMCCI732m3ekUZUi5WdlBCYRiEkNrBA1AZz6S1y4MNtNwSumD2tuHut/ewwBJyPCgzU
fPSCrzNlcfHM6vKbn8KsC7NcUhZS05E7VXyGbe0/bFb08Pz/+VrTq2QCi4WsNqdp8uAWpOrIDAnH
jP4Mn8Hf9M1tQAoQIv5dwdVu8xE3W1LNi5yiWOu6meDdnLDzn9eYD/1+rM+BwwloNXSzYdiYZqcP
b5coMkED4M/oGnx8sZmcnPOHrdZbsWtKUlAkvGYEMuSk6sTvtWl/Q4vHUTt0QRtafwu9qmgYFZAk
uNZKYqoWjLgxc1WghvrMynBQxPI3t4hJU8db60Anp4jw+oP6g4L+mz0o6m16C2dImkV0LYB47uKV
veQdq4hb+Vo/mdU9UIJHx0NZJmUTBEGDZ8UC8HOZEh6reytcuJ6whtkP+iq9FmmtCULLnz34zFC9
DndrZv6Yz9Dg3HNO5lKRyVxdnbtN4xcjDnTTqu2Os6V2scFenMVhzD4xMA1XXKxOukLvVnphJD5x
Ln8pxYnBZ5xvgHOftrBynvxHLtE3CtqFkoGJ6R73Au8iZVYu5ypQ00iKIBAfCTAZ9dU/D6tWgaaX
JTCEOqbi3BtbznPOz+szfDzXoOqNxor50MEn1eEdvp2+LZtdtzB8vR2pofDpZZoIf4fTiiuqKQXB
FndZCjoJNKyGint5h4GkdGq61OaaYSN5O1RBUSFLhwRCY7wSRE7YEA0YscCQwYaeSNzQzxvfjM5M
WexyEMqtz5Zg16O2Kpxk9G4Yq9TGNHTX/nsTdjgkwUJ2xta8pUx4c87zw1ShiPVSX0KcAEYXV343
b1ETk2cZZhZrk/MEF/dY8QShE8vR3xIueWpWEI7uZnEKUuJDLKSMYaioXZvnaF7bGx4/cwmik54Z
Fk/Z2XzhYNo8SiZkDX1bicmrQm5gCg1rlcy7p2Hj0dTxVoYqf9B8S9EdluMr67bJzBB4EquB7ANd
teaXZ0o4fv94uPEUSSgylf6eI6HG5C+He5dsBcjZEV1OiFz5LRVecG1mnZmQAOj4P0/XzAgdbmVK
tO+eSPGOma8CXjUjVwcgSaYTQOi4gZyUiCT6f+UQT2TaaxJddUQ6F2HFNCRKjLJwr6LiEZfjpp4L
Mgxm0rgPWvEUrCu+HGnukrjDswt9LwCtfXMVUZm84qsFKdrubTRVNDwozNNNWytai3cuFAdUG1CT
/X9ygTmeUpFpnTGcpJ1NdwPWPlqgzs4RMqqIX2OiBU00hUY2LyI83z8g6MK23yorQC2zkbIvprN3
HI3FZmTEbQK4ygGs3aR9tbm7/dIh9W3wWhmuLabZayPdY2wjR7BUtf9jYIUk6qI6PER+J4799oPh
kxtYrWpkE5LEvVM0lrADNND0XPiIhfrxqDaZSu2GwZmmS6IWAiiNJh79VdYyBaFJlFj53iHimo33
smWs9Jb/qKxQ+zUibyHFJLNgX9DWoeiWuyHJUG+NCap8cMRcUEcSwMphSwKrAPbkH6P+MKGsy6Cx
0NXA17saxlcCBDCsmhf9yXXlyQhsgK/fL30H3Z/cM79GHq2KlDtYgLuZVb3A+rafvYeBgqOvV6d6
6TIfgtCp62AKfEd/SnCIQecz++Pw/RI5rekUet1QbAI02iPF2etmUtOxer1JUFxMXgn6+HQn52y/
3A9Ikn8H/hxT+j4/OvrINNVaFYaWHkuA4FbzTmqhDfxQR2baOBBWU6Fw3SzZTqyCqaI2cGp/vYqt
KLj1gz3rn7+8vkHosTLfz+t7wDCze8Xtt6agdeZ/2ItnpYF9nWIjT6dik0xAHnUH3eHZMs644QuD
f9O4gjdzxEi1IKOz8x33ZWCSAhJhRvr1cxemLjWYH8OOkAi59m+F/SXuX3MLrLCixL/TCHPO2BGm
AjLgLu4nLJYFigqBzBU2ofoqSMQigDWPQYSDacqufV/1Mo0WTc1fllCEzBovxIldNHHbAsfEVwf5
2U7ma+WLOLKofOEXVxhQd77iregaP114Gne2/Ii2DuVG8ng73h4KhaTReOJ4pkalYzylWEmW3hfd
ZsgiXs/swpyWFxAUweNuj38bbaE7aaz5jzWCZhFs9BSeO95g7/Vjr41D/XO60AU6Kr5C+KAZ4WCg
/Rll1qtDf/R+sUL7pzsyeCiXEeiXvLqh2bIlpstQDAJumXA7RxaofQZXMmOSqhcEIZK2zad6uKrh
CX3pv1sL/AdA+koO2bPJqx/UwENrcUMR+1XHqG2ySg233G4oW2dhWTRmTSQGugZUpvtMOK2budle
2oA5cGgUwFDQ4RLoBCeOHYYEejeGZ6SyupFv+UEtjc6cZtnn0JpvafGoIlf1T/vZMVKE8fdtAanb
zQFPsSGRb/FwJFIN2+bKtZBfFXDG7UrPL/g4cu9chtTcOxt/ef1CklaGHK/B3+6Xf6k1x+1kW6Kz
GXXmGmMVw0Yo0OxIKkoTx5DuLnmlFpBg069VedPITjPNMgfeYuxOHdYb/DXmZaussZSiAv62ohiI
J9eCWZkMbZ5EqEPDsE+Mi7gqQan1/jj7zAg9FrMK4DbsoiPISriVJESt/cnhkNI3Qd5sRnizLHG3
O6WF5vW5b62T6ZGXgbprKGZgSgxEewi5PDOtyTN1U0Lo2H/5pCZas1yo3ZCZEG/wlY89g1DH5Ca+
CFYiN7GsLQhqxEHOA02zQJF6ZvqsxcVugKGEXS90rjZLQPc//9CSm+xp52Wv9d/EVKq2iR8fr6yA
TJ4zhRPMquWduRh2hcz2GuxNqr7mkYy+wS8mlL+eW/LU+5W7fY8WQsekEEj17M+XyV6Deg/u/nLe
r0zCWMbok+5kk6D/O5oAcXlvOutYeZphzxiaSAJ2UnRQIKIhK+MsuJmHzlyJCytQfA/8YOOGv6t/
zxHYFxhci+NCjJds38pj85IK7pCS7oeMS9SbRZKzfhf3zSHh9KUpAAFoG/YtDjYgwmV3TB9pSXD/
3C5jw9gqs8z8p5eFjDfdd1vZ/mrisYCJfC5YeOP+elE5mcaDEkSQ7PlzTQg9pTEQdsfx4igDyv99
K2xrzINYSwlHRQ3AacMkc0PkUz/cylUyoxCxYVZfwLU8CUBdp7YMSQu0v4H2akecnKOPUozq5Bc9
QbDzzKorpET895xLx0DbFPRtGdJfHOdkeFVKIjY676pLyXXQ8UJ6L3drxFEJPp4K9Pp68u3+Xxwo
EQaC3bvGwfcr21niWbtNy6WGxPwWsLR+9whonw0Eou/1zNa6LclBqsW1Cj7RJY7KHReCdOvvcQz3
mh6b2sQO/fq4aYdX0I1HKXHK6AWXEMjiLv7Xw+jH93C/FFoA87vK1QBvAIZuaQQ7Ft8VOpvjVTE+
5l7iTO2+DUuVTHhGJBWs2rx7folXkmCpMvkRArTJXts9BB8OI9kFyl/TH1srG+BGi6cMvxzssCqj
1Oa1VgedMLEahB3sApdWuuOwub2Uq5bOzi1d70MRAyMUi4YLLjlXxquzndPLlUxiincfAbo70IZN
hlPrhDbbppOVgaWC9GcHGePuK38hHl2E1TM5fpZ0kUbfC6MbGlT12sT60tgrbhzC/t1l3xU/qTJl
OlTfXEmN94JEeL5qMJoJ3LwhdDYRzheSrixChIkBCPpiTimZXEOmJ49mhpU6RGaoAMMsypPBQItP
WeLeotjaWSbL4tMU+cXxf2ANEWaSwRHGgzm57h+LKMWaGLCVk93g5h3LFCMK8vFBchLA0mGtZasH
HYuBDUJmqmeWWPpFTQWOncc8C04PyMD7SPdatVj+GUtDuCdTlClB78D8T4TI7ptKgfHXnLQ4LaO3
jUZtAhAgHHzBxnIjr+k337xrAwOoMhDoFALBNS3M+n03+jy5ZgTlgLD5oS8GCYci/Na2PoDX+tIB
PkKOr2u79b5lQvpE7AUi/lJahKEH8uPBz3vYpvcGe1ojYWpDrA2kCpMtU7CL0QQqWIE8rkpb+p/A
CD1I5n1MJEuzHPxrA1/Mjtn+RV9ILs2UKTVf1qM6ZzK/x4ZfjsEOktHNKx1oux25NxLgLyfz8EHb
ZocDLSEc3BQG1HBh1dzOvkEzs6gFJX/QnFJRTzP7OXqcZMIpO57REBFQ7RBHBtG90SIKyR2+hEK1
Uu2mbrmaPclmURDQe/QStK5vkHktaLalt5A09KGY9L7vkzDRLkV62nfBfCBwMvEVcTUAi5nzNFcN
yxXLGY/LmX/09ZDvuinUsvcY32pWEbxCtRjTei2fFhERctVlsswQOWUbZ2aEdpAM1ELZxHRcFosf
SAmOrgFG68be37CA9oYHsm4YAiGi6JO8mLXjmA+nRslrp0iHQz0k9ImCeJib7xtwFSI1quHh4PeR
9HVj1seUqHLrmD8tosz15F17JTjAskgnfUnS69Y59x8E4h8hWZPg91VkyJnP6Hsw/nw0UijfGXg1
VmVIYINNi+nhJZMgVmX3u+zl0mOempRZUlhB1UyFcSwSMVmZFM3/jJmC+gDlFWrLy+2e133CkrVc
y0jOz7Pzh0fAuoH2e/X3xPX9VcFlmZE20Z5Sprlp9GzhmEqKPPsJ3bBFUHsGtEGCYCxIPytFD6UJ
ibEik7fwCJOGTp2cg7R5g1MnGwHLnlmG1Vvh/BXhtb+Va0sps3bcQv2LGLAiSOZ/aHq4X/MqOo3e
HSUDCzWMVZZLL5oL74Bj/PBiKffbY/gWTZajcwbdv/eHjCFjIro+S0wpsN2FX4DzXnk+l3rkS+DG
rdoQdiTymWECC0vZRJwljW94coPayga5zmthMsUX56Bk25JzCkabkZazzq9bpYYxZXbwlegnzwMo
xIEA8J/XvF8cdP4oVmK4MMlQSU2U2lXNVBtf4WWHmKqjdir90xnSGWh5UOIPxHU5POVuuD9pZCbh
+lp52fwb2R45nZ67Yq5flHXVGynLOw+wCp8VMx9qyfcNSoFCLc4S2PgWo/iABKN7fh+ptUMBI0bN
vJBogP0GygxSJ6hBpO2oh22iNjkwu3ijjnMWgSI0UCPCKEdvzzWZqtvHQLqWWSNE05GkQz5QspU7
LQ9U1G8pifYBES0eeEgYgz86/mkVMAtgM6rA3BKlxqW6PgY//H+cCycAkap5FQ7QE7zipeAYttVe
FmFnQbKnGTtvfNwxB6OXjUpLVQMmv/9XqTLofScpUbsRBSPmZ1Qi8W8amjM1B94h+98X4HUcCGw1
5+nguMPtt514M2yrz5Rzx6azBcVAx7IrJD8Cq77hbTWAJsK1Lk/pp1efbQwiONVLkscLse/LZMHQ
YKMpJ6z5awKQY9AA1M1MpOw++NTpdSOvpZeiDl0FTU6RVHkKA32+60ueNkMlZ3ziMbLh5/RECqWR
3qlW130Suy9bTE7Mehj1XPY4uDsmz9WZklDEk7S9zGapMMWYR4ExYLZLRHFRZFPyOHX/z320NxUx
MvYXlQJUpwBmQues7+MrzHzfzcmY71uxYt7DVvR8BvZrqtisuepHU6pd6oPJBf1LQGmeZI1kEd00
nSMBBsv6ZVSxSYIDDcZYG5cer4Fn35cjDGERJLb2GSC5K8k2xpIgi/JMt5lePQrCW8ZfcVqSc+I/
CsRCeCRnMFtJFYR2DbzEPwcYjIqKZOaesv4XLnkxOnCZJddMRqG6PfktTFc52DC3aULJzLGuKcAM
cerAi9GjExSfcArRSvTsRfrpIv6f5/nbF62kC3DU525T5c/g1ZUQMI2sU8NhG2Dqgpw79hPjO60w
UrqbrLpXoJKLn8KZOkpFCrtXqgr9V3t0O4e/JuzU2L5yLzMlYs195SI5MzBxha67mXoxwZRUP2DV
9l4xSYV+yIB1z+QGiBHu+FiWcmPEtADRIRGqwIQA90FWe7gLPeQQk0Lm4DDZQv+t9LB+FDL7WGJa
jjON02dxv5CCcyXJnJMOCbhrA16vRezURZ/u3A9nOAazA7OFrWo9oyxOWZhjOCsLS3CcpFV5PiUf
N8ydtFX+v7sjYX054/QTtaGB66Ta/IuAKU3X7av1u0lY/N4x4kdB9VkLMnbES49YvpC3WBvp9ouR
ER4WWjrnn5aae31f03cPrbRJo3yYfTOSuwwaXBn4bZpCbfV8DnLpOXFBedeyQYlR/GLNpXkjCv2H
1yr60FprAkBvQzzSV2mhQaD9Uyb6qpUGMoxgugTeyxDO+qy54Xr51hb4VnI1SnsqC6VOl5B4TK/h
SqFPIGN9Peu7bYMcYQzXqiT2TQgLdp4gUWoVRKdrcFDJr5MvH8mOvMvtTvMlEH8vfXf1+SPXpE2F
vmM1xub13jr4QtU1XUeTrVUbX81LKsWoQBlJv6ihNXYhNpkVB8Xz7VQy21aeS1yOjXSCP1TjLsRJ
FvmmG7L8dzLQ3xJwPFOQujee+jecntTdn8xtw+etXxPiu1Lrirnv5YvUO/y65bkS9n5KmfMXCe9a
ahu0jyna9M+/zWBWvjXZiGAAO9lp2aWn19UrIkbzBC2cysHq0K8lYsUaXkPOieKdPaurYUiMqA6e
K1/c+jXJg5oVeCvsF1SRhSjTDj4dhGb1VmiK47Ost8iF7uylf0GIT2WHjH9W2CodVErEi7wjd/Zq
qN9fW1Zv3rRaKU2DZhIvDWVQHESYdVAJZkzjjiQr8nvs4QYGK84TOnCelc3aS0JCaipJLuGNgRFf
a4FJfLohiDnwHYntHJkUEVYShcII4eZkWj7pDy3bckPfI7y+br6BOusW3NLV4ca5rGUvqyGdw5Ei
RSS0EqMDOlMlujeY5CfLp0s1zazLvdKq75vD+aKJo0Z9aLnRvXcvULLLc3tYg5ipGwoJfYscpfbd
LAzf4l6brUR2GcvFRS8r/k595yi6MHMBMDuE5RDkYLPDqu5fjdad9mklmreeKBoYqYgxTL3zUG6R
jvUMQKhNZKkuBlL3ThPBVQOZlis2TNqbatxgasy/1+q8ouenGJDUuzI9wHt5k8UY1FUIjHj4z6EE
p2jv1W0UAtE53+FAmmWrzaRcjfkVcVXSnLeiiHallFMXG4GjoSmkkjzZnHo7MT3tbtcTutPpIUPx
c43oJ3aUr3JDJfdU0AH/ETU87WDCDMjdNP73ePxp50BvswI4ehP9RrYgmp1Dr14bze+qgrlfwLme
dKnwe96U7xfFOxjXiOTrwKU4telD3ZtajZ7fTEfPCeyvHWtK/9LH5RDA9VBqpT4EMvytmloswVNu
unCOZ8tu43Ue1MPvKHSHFMMMkLCz57x5a8bvJe0C+6DQtywgAMLeV2RQQwOy3ItHIoxhbwf4OAPn
O7/92YtDTTLTIDNo+4ITIjfCikWU74a8EKBCX832XxG2aLCh9dPc8iiKC2OaaZBpBa5PYCr6I4C+
CG5Ami8Eew1SqzQNyw6JknCLgrSrmXY/bogdyPdEkJNcQlvrLfdQq8sHg4621iJzj61Mjhv9h144
1zeqmXcQwp06ZGkG+ezb4KhL5IAtCQHFMNRC2Wp8PkDbBQVxcsZixm5ZuG+w7UsR1ia+bVonAc40
RV+ZnOZoa/m5p/LQVo0DYoEg1DGLlSRA+HpireJhbrCmZ37l6y/366Ps991cksY935g9tSmaIfN+
h8p3EoyD3gm1kT5Q9svQwFcRJIotVgAiPkUh3c1sRNpSWcr5fe0q6bfqOMV3gDpeLGHqSivDw5h8
Rbw2b4REEJeEURfXnTZAUtzLep7tJX5ARm/Qb5yqWLKapNrkbAcpmAlJ0KjHYHn9SdIJVU2rkNA8
32NwlIxiDl1xwQoRrphOACltJvjcA2ejSBxbEF4JzW8rpBDCfXMMp+Q2FwWOJLGBjdFH71F7TpgO
tcREXqa0OVkNPqcLfOhbuJyjmdRUyzMYl0mPyd2SvuNRDi7578bG3dz8mLJ2UEelk6EQcnDmsroM
fvZmtEOKmXO42ul3bgCwM9HFj2f8Q9x2XFnv6e+jsRvT2DWcnhkXxhrIgPLl6zLN141rSrA6AKIh
Bcx687Fuc92leIEFYu3BPKE3y2GnJs8YquKGNpuoGj/4ooSA85LjAmYwuBC1XKv1medYtxa56uXg
+fOXa0ynHAz81fpHkdwp5kIHqOok1/tGae3++c6REfbyHDPB+y8Pgji6TFzH/MULhkbyEoHfQupk
78w+lb6uhKqwCT+hZ5cEVRbcQvIWzM5VyDy1gCo401pM8IwC6P4rYbEnyaHaRy89HE4qHFlU5L7q
++Ca2d2RQeT1woby3TxDS2r7W8AsAOuzRg7vn5GeUITYHK+JDlu2ldYNS1ip9Xy/LFTwBq9bDXrU
rD3M2gG6bm/ugqnEAlVojwdTc/gAibra4BzSUxFidVYOo7LMy3CfYeMO1H9+QIRiQ4C8UqkmbCqW
ZL077WxK86rZrlulVV49Nu0nNjjQUV1wDPCnQR/gTdD5mz25NVmN1YibkwuSJiFoLtSb5pyzDHJf
JJTB0N+l8Lxbr+qXc8ISdwbH9wxMxKtTLGsge2Gh7DE8gyleRF3fFOjwm2inf+Txsq9YOA4Q7jmk
PlkdBEZ0zA0AOM0lAxDU8wgcOgQbRbxP/9YHfmc2DcGj9mGBjl+Nj8+u/kxrowXYVX/JvN6W/8ue
pP7ef1+35BGXErW9Lk9A/tK+tkFHIqiQPutEi8Fup6OXIkBuVsbzLN6Ka9aRviDwH3jb23VipCmg
fHKblKwDitgm7zmdNRgu8Z5bEWLFsKHWkjytf/YSl7SgI5Qkb0PUo9Le8MVzS7qrgjQb71C+pHzw
gCJRrSbjNHxBBC/Zxn1a9gAvjRGLAdNAjp7Gdhi61e/l5lup2Q1XbfH9/f451VRi+W1oVhSL/Nwt
ygRvqmCLYp1e/lDmIsAPxsVSb8cNhi/QP5v90Se5KY+xYitrUKh6saS+3h0x84tYxCwBMk9Mxlxg
kcinTvaXz7cfx5TQ2GEwiEzOcuv3Vs81OKuU45ieNsSztEq1Ga0fsW04Iv6kA/TcI6O4BnT0bcW2
x7Pq220hYSOCxvDg0LoIg9L9zAwduEPVPdo02OpKEPD7xqM9pDenA/WwdFdUBcytJ+voCgP+Byc1
l6y3dKkkWr8CEBfZhKljVNEN30SiwKngvQUorJ/kZ1r33gtpBRGDON8+uihLcjoLQGxjThWlVDZx
lPpLViptIvFjfz5yzurRQ+LMG25uFYsZjkXoi7t4FU778M9Z5ExEng4wG7LV4OIwFgekNHUZ+x3V
RI3HJ/18k7V3MSkZWOJT6LY8KrnwdxIHw3pAQJ6B/814+JjSlbSKK8b7fvVBqEom1ilRUvFbLDlL
A9ryMovIKGlIsLl3cOGg1494ZO4ZpgYECyF42xCZmlG25icukJmYeSC0yFj2x8gXIr9edACAPBBY
agTJRsRuP1P6i5kPTpMY0Rq4ZxaVGRd24dYsFzYtFcxh7gEcdZUQPVfZbAP+KWWF8/pSR8qFTX5T
xeIN/2YijclWR+dJidi+ZMYgWsoslb5MwTBuWAzJbzMK2uBdeJkJSKnQ9SwQemn8a3g3OrwYfN1l
d97WlF4Z9jHNc6fuSxc+A06Ri0L7RzDnXotzMv6viSrRGOrmQGg1MZ0A1I3Pl/VzHDHUQYN0rRsP
LsMUVfP7AoEwHwBk5n9o8pk16x6XtK4sTyaVo3dUNF2b10WWuxvOagCScCJusPyroTFXyQ5mGIJF
yA7Jq3ejb/Guuy7RqjqfGatLXQUJ+hMUudyjfhjn8guu1GoBi+T/ktwAVjxJX3D4yJSdGLgcSLyu
CYmFdwmftmxBjc8xgr8UzlXzAfMuzsXUZuY8YvAdp1yjXAYypvjqqRlfkvedEuO+iswPtQyumm18
rsG2ZFMfMtOH/zHr8dH55wl9OBgwSqIDbqfVAMTdvE6E/63iw+jpKKRNUg1KaBkAird3AZA+01eG
32Srzj+YEzsMAIEzaI0qjZirp5U7uIunJ/SSw84y0U6cvD94qxxPnNEAgz7rIKEHHKIv6//W7SNo
TJPbR/7bq+UtVXkok1tas9Kf4mf5O+HJlAqAyIGjlw4B3WrwSGe5dmsqceXFN7oBtd30EvBFfskG
nnUwLcYnnC2Xxd4/LseSPO2hOZBf2Nk3CD+BEEDTZcWkKu836SIVVnxkIfeq3lIvXZykjZWjzTD+
W/87YMoZZXpaAKLRFbYinMgJfHucY58LiZBDNZqpyemSCmSCdUb9IFJiB4720TaVyt4CsRw7x4xs
WWi7Yv/FeDc6jwdtDs2bS2aBc0jHRMpzZ3mh0WMT/tBYS8VAgEg4CTiIb2ZkGYC29KyIZfa8Irpu
gPzYJ7tzdTkR/nfBdl2Xi66f/6KUj/jZ7EdSeRmKG2QSAZwKbmgijMhxrRl0RezTv2wZ5cORwQf2
fD/VNrumhSBkfXWpPy6v4QTadD427HRML9wi5HCr50byFpDEB3Rdb+VD+9V+/RAWD2moTLcbroAu
RPVqn8OId0u2UJKgWatpw5Xl29cjLAp89W3R5wGRJjgtYvXkqXUFLwCXj/3e3mpCtrLw4KR/dBl4
GvieV2Oi5vrOPg15RoWlX6BCxaPmsaPeLITUAFzY1siK1vsgCxK2ZVKyZs+SyaucLnXfKfzt9Yxq
C4Qzt2f/VKs5f+0jjM3SGsdFnINYjXhOYjC7dF7vMJGWiQFNKDwmmzvl2xQbmIYTUDmJCtQaeF1p
QF/Hu5HHtKfKM0Si48xf/dYTJNV60pbzRBUX18djbnx/vWcrm6igdckv5TNqUUOk3c+BFLtBHwtu
WK5Jjn9+p4AvzO3re6PeuFScZFr7o0s8PhvFXGrLgGY3iHHPpC6AHwUoP9BOhppmpKp0LoXjbRFn
a2AASZk7AFyvrKV3ST7nZrMUehCUwhikMl0Z7MeThJtBK4jfS1uYnVsH6Qp3zW8Bz+tHt2wIyrbw
lY/kc8Fcj+uuOAI5UE3h1fFPNOQ3lPPZZWpfCsOHen1xD5gDyLoFYoTyGaiNDGgtPDxvHDoCd4rh
79MG8lh8v5xIJ0mxJszSw3twTRJ/L/eHa/2OFfj52HeLJBHumVtVu1tz+DjXJAOdZGIGzFfpDonM
DCFLPPnUinLKYOcJeLhqgtHVvGmd1whLh4Hb+vvvdKhySuPN7jMib05pf3H8chPZh9FuL/aJlxwg
zu4EWoBenTWmzchdK2RTn8UtxN40tztBtRT0aJgt1m9SG6XhOYtmLK8hcbA2mgORf0rZCF7eZWBb
celEWWjDpMdJ1TnqerK18LlNoPaUG52FG3uR5u0iiVGRfG8LqRU76faeKdVeSbvRBhhjq3/ocwmm
D9aZ/coXxYnmx5zP67j/dxWhs+XrEnEFi0Z/Fz2NaCNTy4R4g/b9B1kjbJPCvPXeSwG8sgM/65j7
IIgEw0jRBEGKN38XFEQOQfYWZCmIJlS286Sv/Y2DPMXBJuyxLq0NWb24Y4f2VaOI7d2+GdBApuYm
6kKs+NSKK5U4kanK4ETThdvl0no0DXfsZ2i7eDj4pHxawZTIndegrvvEM3Q1yfAW2ansqAiehRps
hhOv60eKhBcp0Q577nhGKPhO8Q50HKIULfhCWZcuL9PtGp+mfTKlJgE9PCxv+E7zdIoMvY+E4zo5
Ls4quBXceQJcaenUhiOrRF+HyRRIikkaWnkKGPH9ImCN40cU8hz1LEUhKKNOWxGpJ+5xhFyKAUl1
wh432cp7RebdS5mRu3VWFjjzIqwaIriqor7ak8S29kNXbrcrYRhuLm7/BKUxp46PVKs9LdgdFWTs
ODqHwQ4bUDA4oZLuUtmrl6JgLq9yVq2MgeVdReptJResCEDXFpu2Qf03rQxQ8JkRWclR3qZ1mhJc
lYkiR+NnFzY+ry3ILi5S61rnPzDQSmwb+/YpgHIulC4I/fcmmKnx+TeyH7BJC9urkEX5PR/pXLoc
PrSCGlAa4WvZMsVPkt6UhMflb4OI/ppFDj9elh/HiuFYz0dEn0ebJl1bgd5y0Og2Dn2P1sYb+qYH
sClCzmNbeZcpmbikIgYPgpQ3lrbMq1pwjcFpN0+IquoWjppjCvdAAJsWliwVuqU0shqekY3YtZJf
rWZYcWMgaG+5Kyag4MgpWY0L5i7ARk35O8o10sI3ijnIxBF+StEvk5Dsl4bn9WKN3SCr1JugYq0r
M4Q0jy5fdLxAso034MwirVQfPdYVadfwyfEHoR4nnt6X9cIEEXRjKDcnC5zQRyQ/N7b1Nbbyf+ia
8aBVsyWmwD9Bl3IDq3gXteuctopvswvxfqeGF6OuemWWxSKXCk14Of4CK3tQ1pWkSmQ7Dhsy5Hio
Vi9F6qvArjdJM11zkDrRRH9owTBriytBRZtO10+vWdkWhgVyjzZGoWd9O1Ae5Tzxb1TnqhLgqzNR
7hbyS2s7+fDuVTYIpJ9UmKJtawEv7yGlBw/StUPg37yi7Cn3stcw/oWx6tlQx7DM6CD63/lDtXJ3
HYttQ12juAAFEFwktKlODP1zWXJID1H9gDYKwKAOzsxSQW+mjIEPrbhBDM7oFk2cvq/ptoi+W7rG
rtNwnME66RuhuzBsDlcy93PLBzIAVfQJwfx5t+sUWYnwA5z20Us7trGEiVgg87uRsnmJncabo0n3
FouLFjMMc1c70xF4PkEDOEvDbTySHToV7wsszrruqIo/pwqSSsH6Vkz1zXr/XtqgvkSGAf1F1xhB
1Tx7run0X6TioQ7Hxoo6KxV3uti5cmsL0Y0zHCAhtyNfNIdRS+LLRD8WH68vXcsc+vwn+8vMeS9H
tQddNLJG/PXbK0+Y5VuBTr//wC4uM2mLK4jNFHH8vjQv5e/EVpDwVwfN1ghLbC2lmmta8QBFZoUG
ZBTKG2Q9Yz5eFe56RqGdlqmpncMC0ZcVkzuEyFLfqoTIznbgMXDpN/DrPS407/C4k3KESHjv1lyG
Me37HzE1i33L3pqH5c+o7+gMf4hi7Mo4qcDy9p+JHK02AB8K07/D0+al2hJgeqWnp5lynEqlmh8k
Q3pT6FbeZ3G1fx+Hm4TdquUUS+Spy+v1Rb0uKWKto4NbYY3zoggyxQ713t5MUY6d/Bw5UCPipbCr
oSUf2p6ncQwoimTq7E1FbV1FU4swRe7Z3PIGCTCZOovhj6Uymct9bykNauh/jF/3iXiu4P1AdfGG
FHlDNZrjk93hb9UL+L8+XS8h0otI1JwX7sBrrJ1KqURrAvwTvyHxKFuFqtT5s2rA6M83nzsngeJH
ND4IiXGf6ANqLDG7Ul48TzyOwWnv9oLswDx9vYEuTFr8D93nF5JATQjOwDZCY+RhKYzQ77qIsa/F
lWKwtCJpJ3TrZqXJuV6ifBCiuoi0DUrWgPmnl3J4cXlm2DhEf4m0pFyEvUUancW3syQn8bfL7rpf
7PmMHPKBsi3zX3UqpjJIz6bRUloT/WVToTV3ZfWcWfyumDmPBoiWimY9iU74iKLzZY43B8ofpF0a
zPR708ODVaMVEpBU4cw/t3U4vOzPkdVdvvZg8kkBFyIjsANLX5AH0EmBKz8Y/Yt0uVaYdPN4W6IL
eUqwVX4BPFdg7ohhz73IygYkqH98AAVC5LG6UFU7/frw6BEkdGMAYa9HtqkqGvUuNwJbbKRWZG7d
jsiQgFdpDuR/gzIbX85ElLROXmYj05QnqD3vyQ2jqJf5C5JVlycae+shvV2B7fEcz0D58HgXlsvE
pRkLauVfDoK7e0gSTHPTiTmXysjK/LpLKB4gjFXH0WY2zdK46LMtF+dxZ7kPUt1VFjpHc6Ff/vTB
5pbeMTLEv1uZ02NzL684/MNc5131DOkWKO+qpN14Pwcxdti7PLRG39nSOARbroM0DVSrwUnQU8ph
NtoffefTpqJoydRWvPRFIh0kUoTyrx/qUfbs4c21D0LbF7n05yMvp3Tyk9gLz3btwETkJO9rRlKX
f8x/b47LSlvck1uOC2o7a4mFnW1BVyGzXONxgb75lDbHzGD3aDMZuTcN0MpJjEH58ZGoPbDkh1rW
53nsmXazjMlrw348XML4YFNkUWuInnkEEI2aHoxGnMNo8f/gHl9fqcaV1JET17YarrLF7Jt5/FKv
DKFLIepwws4dg4Qn0y4NOxxr0TktN1CM9MHV3RMwrOtU3JE9mAvE8jAfWw5Gp/m/Zk9MlT3VAWRZ
sSY9QLLzkgc6RkMp8t3xN84HwHz5umvM6VH5m1jFE4gKn2swbdVYba0a/wLTvQlmTy50Ux3yFLi+
pLSfCIQ/oNQKrDtcsCJcUZz47unDo5Rwq4ZTzRlHZaeFAJgpPxIRb5IORfmvEZ1mz/14e/fEtu9X
RTz9fu050uUmHadxUmCugRXCdMXzQZavr3JIc/Ss6SxTDq9z/csObgzW7J4SATcR6Y3RUmklbg9f
/Gx5x6QyDUiD2eIsLhYtjgy92AfpCxkXgRVARQgGiNaK2hh0LdspGitEw9X5GP1eQobdYH1Qyu6f
c6A02Q/Y/LuyA77rGAr43e3qhC1Oc/D9N8aZ/bqwklvNKpIG2QqLZxteHubKeTfs4jWuyMal4yF7
mb41jAtg+Bd+Rrh3538TsnSsF03VXr8TaoaHt2faqNZjtXw+0upaSnV7eQhlcV0MZM+FEpb1MzlY
2hT0h/6Zo6HSincJqpJ1hNylQhXhU7W/MtmdxAcatkcWJRqpgnJ76s2cQHfoveaFEj6JYFmBJGf4
XThwyan/8JdyxYhAozpfluLy+IAr+T3BK11TYwD1EYstv6maEmvBfQ/KT3nB9g+/vnxJCYXHi6ty
A0rPuey5z24D+Yb1X/2c+2VEPYSQrKsbSc2aUqWD3qCb1SESYgV6Nkvj+vV/puxZS2ETKwoKjCqm
OparRDHlvGcXewmPCeNIwWa3wksG3H8+ULIgtw+L5Tab2ZI5LGj6V/mW3yLCsZ5lmDG1heOGcFug
7h5RJlXcg3N2wpsiUFnVq3kHDmPGL/tT7Kof6lSI1j/LyoC2q0WpPGWPtgksjFLHJpDiXmP78N7R
j8ZX7kNuZN8DUdXdJZoYmi66eLzzRyZmOBBbL0vScmhdh8+tssBVdCnkVEkM1G2pI2M+DO2PnWZL
z6lmKqIdHNlLRoG1rMYK1/y4Y2BP3Iw1WQdemh/qp4sJm02b0Yk3f3Qz9fnfujjRQyQWyvFa/VWV
HjGKhDyLZBMWzCiLRuha+kPxIuzah8MCUgVOGF3kP2HjGo5jXCIcqxJ8PrERcIJlYYnpfB5eit4p
pyEV28go3s0tHNnS+IR5rcQQkXAI/q0AjfsD+NvCivGOTTjURcjk02+/Y46rQgtUu6Sv+z4o+7Nk
F5hnfnJ/bnlSWIUeD5dLm0Rlacla4dwcygt/KNcCaIQch9EMeI5HnH53LkYGsCqGzFTtwA22SdKV
M0RB3/BXNbLhD2nb66WG5HYH6QnRSGlZh5D6sIJwOtT6WXbmUgzRbedNimtFdKIYn3iqwM/P9++c
YMINqI2L+vRm/h/w5Z4XmA/VgmGfgm2M68ajyhB8zULnScuKcWhmnIFiHhNROybuW9X+avzsOM5a
vKpfkOlGkyON1qV0r7QhioEHCN0Y20tVnOvRbgqhXraTMM6DIa9qM/WMWGp1wfj8WHzse4CHMOyx
fQAkRF5ByWL1AWSYVrHv9lweoEcU7Dnpi7N458pQQYR7im4BwBSGqVvGeDhSeD7XnNzVbN2n6f7M
hr18Vf5iCvqz4/j7cmLbRjIAQu1lpsUTiwDxVm1bAn862PlN1O2fKRYbE1dSlqiPoQLxllyQzFXx
QZ8KUN/+JjBa+Do3MJQRHenIn91e2JoQS4Q7xNuIH4YT6ZXs1Qx7IREY4avqfCYNEBf+m2YXly47
MwDDSZDfqbuiouWgCECvb2sZHiu2scJudTI3obxag3o5aW2YXB0t5NSnWtj7QSdG+GXCGl9Z/x7L
X9oZ2HM0m2rz7uby+u0nSMtcyKEsyx2uXFxa58pjYgfOCpzxB9xygOYOTSrFY9ZvUUZWqeODRFRX
rvJ5ulHYdEThWSIubAYxVLvWmszwof7wgK+C+qZ0t0+w9vuSa98hFv+Owe/zjO0DmR3RfPPY9Lm9
rALoJbWc7Ppf9+Pxugda9BXLMrly9Yq2AOAB+E9TGZdb1Ni8L6yhGHusZF8h8pihVlW91bpmpQWN
iWiidxMCdd84Hwne9GfSdgKLjunCXBge61v91Pz2pjuzlFErZWe6VCJQX3yIsfg55zfYrYZi5/wA
hWzR1KhJH2k/w0P40uTZc1vo6Ya7Xnl2uxlVnO95HTOO0+Pgalokj5bfWIn+5HjER+FcihtkKlR8
HuPhxGArB0TdmGvK/Mglt9Daw4NCFYlXAPFgjWZp6NfIiITbTBl3CuPR9mf/Ow6kscvXtxQEfdih
JNrlQv1a/vAbP/KiOD3SV6/J5ARjQJBrn1r3jsjEsYAyIn4GZdxJtsLaKwdyvTJJn/OeR5Vaj2Z9
8rNqdfSHCuQxgy8fKyKAHQCMPu7Cbp3NQVjCBf2SL18oy/GJMo2BhAc43J4Du86dVCkIuAUblSBG
CQLRF8Felwowms3/e+iQzhgjVFp4oLzITGLTNDcIGYvxnblinzs920w8Ub+g2qQSIq1RyEeI1nYi
IbbT85YPyyFar34GviMK6ft52n7NOd4sSSN8L3tlcNWewRk9gccDRG1xpiUTq7OvioBUsULUFqt1
69rKdkqMqLPXJJuYGchQTYR9f+5IZSjQof5PsDOMDixrfk7Kwe+q7Savx6QrbFbLM9abmcD3cfi/
pzJKN/vYXWakpka3Q/wxT+Rh5rEfJmr77xuhC0wM0yHLqbzk4Edpw2h6s8S7JAgEBp1/u7JYkXiO
ZmcpYFDNWfrxySUv+dTA1NA2Jy7iPvgr9f1HbItVYlurc1fOcfarqjTcPzgh+jhFjY7cR16qQ/1J
rZXYxpBo/5cByLjfyDYwBh9jLmJ3siFeSbrjKspnILZEvULGqYETy6P48vWFjDsZP1DDcoKHeS6C
qn4qQlYqmtbazUegaXpRVB5zBp6OZTV5zSegM07GsXNJSzxOkTZSLoM6V7Td0xygcrDbpagDk2ig
ipjx+IbYT0JpMCCO/ZuUfUwut446/SEU0zIXXkr4T6xf9uFq4CrdPU3PnXbGzx+lk3mh+XC+JkQr
NyJFr8XYEKHrrl2OCJ1KM08iRYqwDEngGLv0AHdkK2Y/62fgC4VAdE9IuIrXvTWu6jnYFYHRklmW
Ab2MErr+LTxR5tq1+WAMQAlZZwwa51vV4y1NEiA85tGSuLUPwqDJ15ufsA67v/fOZbks0m3wkbAh
Pql+bu6OBaRU9Ij3xHkQvG1IZfzOXgTVq6uVUy7M0ZNv3YXKoP/TRGKYV1Z3sFNPxGEB5TsrGbDP
aCsXrVXrX+j2UagX+cMEXBIbub9tvDiQIFAFT2quDskxAHqyDxEvre4twdLeKn5CfRwXDoOFrLHW
xvKhZJKe9OpXa0XTr3obCeIGsaHWK/C/VlNoebH/Xy8jLSbaLJsBq0gLCchRp5+J8RWf1u54l3/g
33fSkGNAJUu116YeH3jTgB7kx4YYvef/rs7yLVHGIZf8nEVilcf29PY0kHFLOeh+U8pupfNYf8/+
/tsQ0BT/RJkXhtEudX3/lcYe1H1rE0Wc7pxr+M8BFIcxTKTe97ufQHVu/UUxDuEk+dLSqzLJRUrY
DEUHduSuQYteLuOfq1F+6T24I16cl4mcbcyBKzqNrxpHN3lAQmt4X+oPBushrgBVHw/NEFl4bPPo
gTm6HzUhMerf62zwlAfHQ8sVLzjDTq2Jrnyb93KWX8W11oVvP6r+tIh2Jh0IRTB+xdFX9zNzLXGB
OUfyeSM3v1Km1JoDVlqiL0mnbCms5Xh2+/z+p6OgiZY3Kv84KnDwMqk1/b580BD1dwC6PVi7Xn8v
n4f49lfTnH1h6yp2oRynkAHQNYT5OLkNgC5ie2wIfqARULNNKtRj6zO1FOwXhOwjiOBv0tg7JrdR
i0BiuT+Gyag9tKx+GJvlDb+jzVBRGeFpPO0qtDLSjkZ1egUOnl99OnHjrSuwLGvI7kvAV+snCYcz
oyaPOY6aZXhL+mI+9JezmzuVvJfYTpSgPj+Iw7PfenzQKbI80K9dmBlaJ0iPytt1oIRibUVdcsho
RfW0cw+fk0esr0uJkF0d63rdeL0fA/29x5CY5mWyhjSxabEcPveJJpsPgPR6digS6ayVFQklioYB
SXq4VYLmBIBuZONsT/WdlaenqNDDi0t58P26okAcbfhUMlz6z/nHp7YkBb27OyuHzL9cQuUQQqf+
iYNn9DBrqAVMGZahL/Zek3Y3vPnXNy3k+uuNqXJO+vkXJcrgFb0lPhuH8ms2WIcqkrufEMkaOsGt
Qvdd6zB+ZE2iUCRz93/5nPHLpPjk552opkIJ0uVTS+ynka5igYn/GScamw/LevbmIF+q8V4X2Nxe
KSwxNjtne2JeOklCbUwXvbxnJT0JCoJCF4jPzq2xC9OgJatQZoEFKNTKgUpVZqT0ppd5z6Bpc8Rx
Qi7Dp62n9MpHv3gPkTYzn+/kAjeH/DXhdwMaggB1cRZsynUdUE1KcbYXx2SBvQ4skGAR+0mLB4gt
n5Yy8Kjx7zIKOJhCflOeKxvft/VyKXvX3LS68fJtQI8hm1uYwu4YeV/oVTiSCTEzp4jEBLdnSfm6
9mgwCoTB37/znfMe60RkRhbl2vRHLnLc800Lqgi5kRy01uKCoFB3EC3CUP1uT2fvMheLPpP8/J/h
sv/3DU35cdBMpiMF+mBs1pULoXVrIKhey6Uc/FmWK4IUX2zavQ5QCWsZ/auOBalBt8oM4XozmDI0
LFUFWEanU7xSrT88//nbaIJMQHa6s2wCKd2UMXCDNIlSV0NsiXoP9zdBEibCI0z/5NYQTKfhn208
5c1jH4jhN6dSSZHdM8Lpg6H1GA09D8y2uFMaKso8VcUQ8aVsfMjFjAjq4tWHv1bLX/turrX9xbmA
fFc14QUyVvo2jsm2hBaI6gfgF0nGKqceraXqKWft6aRCukbCBcnug8OaguH9jBP0k0N3qgv0p+ai
JLD2g5ynUeYH7Kxnva4gNG4c9xQrtPTL0ysLx68fzO/8zSntELPeEI6OA4zYWhn8/9PvAwhyE9Qo
sIFMMPYsCi21nVD7Fvz2w2E2URZoT8i9TV3QstZFLcrFzxyAhuDPjZxC5rHW8zMKjEzA0vIAMEJR
SWkJnAJdQF5dHedeQVWK/Tia3mComSO4vpoYUx339ABY0udyJ5vbxDjNm0WgrT3FFPjh7eTIt+yi
RuANCV9CfqTqbWtoYIelT740XnaqLC5KvyMWPlAXtNbpXK53Hywq75ZsdRlAIERXipr1fygM+HVy
G9eIJ8m4dSJoPoxGJ2vn+HNFBgqGgynEvwG7NB7zJeYaS+V4+DgWNLYt+4+lF2p5R7NJT27tHhPq
NdcW9UI+pj4DDHM+pd/FqGqNLOH667LDmbbCnw8YZA0duv3bDmeFhcEIeoxP3w0pMeYX7pdQoiPY
Z/TseSFt91vUCfgs5IZk7X0hvFPYgrRYPLeoNRyRctrrovG4CGNQjy5zHCdUjDDkGPuplvb8gtE/
7kYYYuHjYiir8hF3PPKEg5k/R8JmkZZHq2tHRS69CbEgepd8mqn6LQrWWkNBFx8F2N+ZVJEBWIWK
w/DKyhpjJLd8yhvHs/Y9Pfzku33AptYKjNxGJUdj5npJVQ1Za+nPexDXwFGcdxyIppRGsICKTVOJ
zPlKBaFzxxyAzfoyMe7KBHoXLJ0gdhtbt42kjZjDV0P+lDAKaUXJL2DQDDJ1DWeTXUUcVFkaiXu6
ZqP7G2ihC1oBMAC31LsUXpAZO8qz6hu0urcun2woKBqiS4sZeDfUHSs+5iXxAbwQ8fxaGD5tf0Ou
vVXpvxOkGodfSx10IG5naLG0w2/fbP0Mwpkncoe+X6vA75bQ5UcmHqlqpVzyS4U/OemBMlKdC99H
KXQ18NUILepPVNBbYoU8dGc34TWAgQpnSUTA6f/W+0/Hr0HG+qDKqQ/AxPRClw4rMcvALrReIA4l
t8tFpsoNMSyTGd/+Wk3gQkQP/hMw4dFCrbZ/+oMmz06PUgp9QD3RVsF/6AhQMJOHby6rER9ECbV4
ydGgUayw/VFYrUvrB4imZ21WeNC3GTo438r1iPUcayP0+FL6GO8rSY+QpAm4nMCjMuG+kiZtvyb1
FLljdnYk07ZRRU/VkfDWj69CyeCdKI7Vq0nOzfRzcjbAcOWt9fdRmWa2FADp04p41+57PQYaA1Td
vIVKlC9P4g1e1HnR8WMD550JrcwTCdIgh5mV1mAzwOIC5uEx3MwE2EaF9tLukF1+Vb84FEu/Bbnx
0VHYI8ODJtMXI/ZZjJ5Dfbd+697ttJBISMVBdfh25qQIH1Bi50MnbZVgllz3AsI2RRZZh13oSENr
LEdyb4lev0xIpl9MOG0nKOKsBAgISzv5Zdh4R8y6xRCW/lrSjZFSYUFlly9nSmKcGwM1aTSEPVGT
SBHGjaEPwaDaFTL3WEvHnyTVDXMNzaIrt7+mdSMcweeX4rg/lQL2WcK3uxRWQ5DGslOcs1PGaF/E
ej4LvT2hOFONtW8HxY5qTMruHpBVcubjBuGNM5JIkKmCQHh3YiV09m3biYqJTU8VNyqve9z/iRMm
7U5BIe3xniGOtcuW4hAaOr7Q/L7IeIQDYcb5e6DuRnloQDG6KU6K3h4hXxznwpbBtLynmPipWvKl
U03bmM+hpmVYyaW37mV/A+EjyHccXYTblYWDcYTqmFErYtOvdPez9gIpaNPO34NHhjlc4IspR8Pg
tYdq51zpFRGYDv22TkBv2eKjcx5eOUaa52V/BvlMn9Lr6vvLJNswTIcfCYy/y+yFb7gKfwUpAxck
Wm9nm8dIOWpiwslg+Ik1DKUxJAjS427fnQGlKUHZ404SfW+NQyFFKxI/PHNvWMM2O8572NRPREZZ
0Z7xaizSTEuE8L29yrnLdiMBO+Jwxauf1s1ud/kRh1M85JU4tTsx9hxoceEQL65zjbL7516Xu+i1
RusKCdwvv6RCYO4VW+jrd29tt5nn/Q8UBnyP/xTgQVtj+t/3Rt7BuqZs8udDQNhYSeP2FKbGC6Gx
tznYEyaHQHgUgyCZW9/rPXDF5ACot09yehI/574xu2TPiFxAPMAakiZvf7JkJOqybQvAGawgl9bQ
IyqoqGwm4LQDiBekY3k9NIe5ZikrPX1RE+W5uXZjRGR7ZIStyiGowHARLoLLhZINAyopAi1cnOWC
tMUJTo8UB23ySB4Icx+2o+Wbyu61F0zoWiBVAheKgpZNQ2R1yVWeEI3dTXTo+IEk6kZ7mfEL3kyq
Z6ODg0JzLu9Zh9YObDZJlpr03CFBDGQpEtmV6trMuHO4oqNIv/STgbhZsMdS/5ZoyivSR9iLRpK0
qLiZ897FPolvQDLvEktNfy4N+Pn2uQ3SKaVauE5qnCRQsMXgpqJFLwJSR6J1CAfIJMVRL56D2NAX
RJMmSzdSdAj8fH/o3M1YxwJdYXJyRfZnfDQutNqxBlMHJhq3lVhNy8JemoF5we4X8pIkIQXhnUK9
l17PLfR6WlnxwbISOD+dU08Xlqz+GOZZE3xuXOngiYTiLTzH4akbW9Ph3LQ2ABpaxrdSx/+vKYIe
OzE4AB7pCIXVcHl11JznOxR3LzkCzpppf4oqk61FAmZdWhwYSYSiMU9Lu0+Shtw14+NNF2ch+Kd5
dTWiPApdbuZmPkEbWk1/ljah+4VnoQuBcWExGVs0jZ/hkP8YhAA7gMsYvHOjP/evzYuBmYPePhBv
1x8wtrfUFCbuI5kPnsFa9Ren1ShFS1yO0nFmfmdY8ZXsk7NSkPVBSnrigw4B5CZrd8pc34a5+Fpw
/tWqwj6Ss54KgVNxQByNZ3On8nS9dK5u1IJcm7wBec12VAFARz6Pn8FVxfZMm96arZx08/J/PKT1
WnFYNr/oU5bTRcuOEc74R69m5O5WGCON1QcuA5QS0tMqWWHaTko0gp4Azft6tGhBVvSr6FABzac6
b02r5Cutf/sbOfPZHHpyx9/bIcXKLuxG6/XeVf/SUhf2R7UrrBnKN0HF8NLRbJchLlqEsKYunNZB
74gYSIvk+W0yRiD1hu9Jij+HXfMFeBxxP6kbprh1iziWGPSzemplkkP1SAhdC1NZOQmTU/+0tkkW
i4Fm+S7a/Yh3RNmYetWkk2BwalnQliBCSJ5FY/jpt4S2IrtGNBpfX34j9Za+I0S+/Is0U34LIL3D
/hNkUWFReli2H2VqU+d+MZSF9sXQPqsgvDE7nsEUeLBNiJiAl+++V9Rrjuw4dugULTxDI+7j2PZm
DBpYRRexIPpZnuiWr/YCYqokK3bkJdhG9epGITDO4Y/zfMYOGH89OfNv6Ogv5ODkJ0yU6Cf8jbrv
Bp1I7qaXM0+XNJuA6XV8JN0nxdWTLqdMsuq6sHedgjmE7/El3oCdQMTX+uT/ymKDcKo2Cz3N5T1z
fYcKunrmdY/uFqJSwGiQKLFISHmE3PPYL9o1zCM77GWgMTnEpI7OOmz5TwnU9otiaiQfD5Y6vEho
jp29LDJhHGxjDIWn8x9wFV36nNzFGtIXj260MqqmyX3YuzZGexqKvQhIl7iMnLiFZm0u7RRGvzNV
78dHt1R/aHk0u2uGzHKdZr4xU0uRMAXROiJOKtyGblPRr0aW3gncEvCZGd+4P7KKYdMlC9hFqSKf
ivZ5+oGDwen2m7VIQNNdQQFWocXaxCsR+X5oeRHwEtB2SI8W2pmLsg3IoVYj+0y+h/fbzJAej2ed
Og099FYCnLafclCQG2HVFxf1qo0p2pWbdTOOj03xZ9Wu+MakMPY/d2mHHr5MktnKsq9BBwWwXrcV
5BvLP1AV6rb1/ra9L5QDYflDWpXC84tbc1+bOF535OKnpBQgUe2GbV6SCKHxnZQPrT+BqP6UuiX2
ilPXMbVQRv06hT2Yr4/7c06lYrToMPwDeYHB99+d57dBQoKmglpkRE09rheFX0SNjRbcEdNRu0yf
1eUYFbf/GWQ52QBqKSZeoRUcBJOMzr6kZMspVvpHHmlhMSQHH8CPa3Qc2r55BNnV64a2HF5JPbgy
23nJqAB1eXDYPWaNDdSe+7WX0cp1j6a5lO0B2Nj/HCfjwhnkYpXpsIQK2QR2Ks3ODDJ9IxS5w9kp
E7XyaevReacih3jvL0ELm5EhN/W8epJ0/jSbsMnGH9885nvq3UAR/Uy7fzhgnqSAzveLFqkK49EM
QzLk4mz90rN2kBc/yjckMUbdgTtk69lgvp8s9DCyJDNQ+ZvAp8U3rahIsRNvY2/NFiMmhTgNswll
wNYc5jX/Lg1yjLC6lnKt0Gg0r407rQRhbeTXGJIeQUvQ+1JHqgJrBfFurnXSYcfb8SdpuQi8efXa
lHMEch++xiO4zR6Ssk/4FZZyFvdNim1rVeR015TC7yVOXIqnaaXSaOEN09W3Xh+ldjweq9j9uOKi
cJehLBR+At/UntxWKsSeGc6ZnTcWgmRm/UnrI2kOhKTgp1ZwpBq/+LRBV7vZRkAV+U8cP1eELYGg
PHGpPCwVz+1tcm/LzMQikmoc7UX6eCzyOghzfMzloU/+R2VZMOaofmPFRpu9s5LkD/vwKJs1uBeM
R7XTj4bS2JG+BPNhF/XaTOZTWAJIXj8EDJ22z1tGyxACRCKXUSXuTylSmExycBqBLAQliOXrmQJ3
kRpY2Mpgu73zuTxZciW+YCCweC5NNZGL2WFre3jbkdCfFMMRaHw4h8mGRpD2CeDvd25ZFT8mquM3
CzL4NbXXYaYwlch/CDuBjN3WIMJMQX6scTI3s+/wZG4j1QaPSQyhb/8hrS4URCX4oNM3e4pes2+c
F7dOSvFeAXrfFlR/Rvgvgpoc/DM8sotsMgmzeiGNXIls/L04T0XeZ4sEBDomdSQdoPQk8P8klpzY
P1CcSv3h+22qi07vAIpGlafuQFF3gen3VAOTA32a6wtAhrA7JAvlC3cvdivq1eYB9DdvZnX70fFa
JsDB7UXyRzE3yuM/Np/au4EwP/Wer4qf98UP0+9QvH45tv7PSJ7+2bF++YTf6F1wvEZchfQ/ZaZc
XKNDIcwi4fi1sV5G220+8rsQ4sIx4doaRSk3S0cj7Er6MKTnJ+MjAt5YQZFU2AzzLmqisto/9KxW
FJIZYHB/x0FKrKua4ezmHspdlcObqzI+gupY0HAmr5JbW15u0e/Vej9yoV5F0x7vxSZdJo5yPGNR
H5RH9CFDpwsQmasgPAeyhHynbMR8QQfUJPeAKQ4YRGGPbN8s5XubZ4NSY/+BHCQuWYkvdiEXw2+Q
rMdyi7aMJmzMR5vwNA4PJqIgjES9/DttwNNXkXVe/EHZ5i/hSLFcdeR0IqeluldbKpNnFrU5SHTc
sQAEHN8FFxAtDFmja81oJiFQiS+wT/W2iomuVYvTSCBW4SYRJqwLEiKYXgz3IepteQ+JTomcOnHq
RSaEcr13X4eBWb1ypo4SqA5z6thfoIO01iP3qRYndPIX2aS2N2d7tf90S9XaPuJ9kKYa3KYQBKtZ
QjpkvadRxiF4006WK097OKG05VHh7VVEVOmfJPbkdIw4HpdXLIYRZtbnmCCq7Pd6C6S67LYUEbfO
6dEDabheLerbCCwHm+h98ak1o2qLhMsFiod1Abj1W+Lgzplzj/9bS2g7MvpaOEIrDvrjLwdu+ndl
V76/CmeFjZVJ3U7BGFBkrJH5bOFUk1KgZV66vEvVNHTxDbpo7DWZO3m3JuPJZt24xAmRTxVafk3X
XzCv+a2woB+tsLWRJl553STStGXxv41r+RGbCx5qhdcEBg6yxnBE+hy/YIkHVRvYLGYqoJVxiiHR
P04S6MinYa2Z01gG274jUJpq2obL09Cjzc+sl5qNkAUojW1dcKBBg8LWEXpe5vjo4uYsfCloWHMj
4zAYxsm39g1gotFapKgh+764mWHU9X5aMaSnxjDPEC87uxu7jcOsmfpHy8/bv6Oq28rNQqRwrrrY
5arnAm8jL8p2C66Uk6KEKcmFUmvNTrZFACpBy0jJp1rlRDp6ZPfRg25kPrufc56bHgJ/pT3wt0O/
Ugvd32WvCLzB+gesL/OetnUYrMUhGLmZBKkx4ahAfERX2QtjAuK5Sy9+YmGs7STgBehyjos9/hYX
8aFl1HdLn060oY03molRvV6xDvsvguLXDnuLMNOnTb2pwmkhL6oGYSHgA3x7sbrLEF4M2XVS5h0+
bcpqBROHwgYEPSK+tuty7rqhB+BiG5ThSesUS31AwBXP0Oo/12hMI0kdaytTHJj9h90ezV8EboO0
fZN59Ssa5QyAgYv2DYgcKqVrg7HW85tXQJfcGaw/q8oJ6Lf0N7EtyidMPMd+Q8ZS5+2C5hjZQJzc
ctDRLo29ezbn3Z/v/HsvFh+aq6ox9lh2h+efUOCktwMmvMDfade2M1hJpxPWIRYuC8LEhyfdlV2Q
kNS8oEqS2Qt/n9NsR8TZZSnfAp+kxabHsEBg5KGP478Yc+ncywRL3s+uK/J8sRz//RaNkmuDnMG5
uG0yH0pSaoMgLFunRpbBdk5djiYyFrWJwWO5nBOlyP89BduiKysJFO8XWJhDuPXP+Iy+zxfhKlHI
Iwtp0fXYmkSRp+hL2jCCD0BV0d4E8SRhK8AeHaDgcXN1k9cgfmVwvvdshGHR2Bhf9MCcNuUmhyho
f9G7JH1dxminHCEwYvukcFMVQJfnJj/crnYU+RvK3AgeyamIk+mjSjD/SckkTaePeb40BIV6WzGB
Ki+gkWFP2Woir8URqcG5YnT8y+S9R9t4uvI2kfpCkrJdWnZFGa4tnD5nOScBrJ7IC9YZCimdwCdd
BkOlLftMAJPTWbUqbCsyBr0mX+NRhFKW+aRd3CAZyj7QeHjzUeagI5r6Pg0F1kECOSqHXPKVVTNf
D/O4kBNbJDX4RWwdhNap01+iY3jWSMDcS0QAbAtI/TPMqyk2wd+XnvnpywlQC8oORLdXrrl7A/Xe
z/DDdNkQaqbcwUdzsKvDu0KujpjaOG5dp+4btcJmiSi7X9kdxpQnqaBkEhKj+rcvowKGhJFzQILl
ea0Hc7ol1PJiuC8if6jR5Fl8NnQE3pOzYbT2/ZNt/AkNTAaS2Q0reHgF4me7L2P65s3EnkWsLb/k
G41AgXhRNhaxZHvoXKUAnPtGfAarC8T53rKhhLUJA7tNjN+NeSbSNERR+e/Z/sTR4clCp3hK1dd7
JXZ2lw1hV4a7kl2AmGe5VJ1RztTLbLYSkfSossFabAtnpoo6P3oSxJwnvq1IihegHY1+b+sDhPN1
v456jKnn71LWkZi+CcKBzDJl5HSYLt51Z0P64+jPYZ6o4MXMHAIIemYr8CoePS6KFG+nugn6S8Pn
Ueifz4D5g/vK2Bba1n744s/7Q/ZaKSMapUaWGhci3pAoKxaRVsJ/CyJwez0eRiye0vv8VRK1xzlp
5ziyEssi5Ba/9U/a1daRFZ9ilUztQoKylg+rpKU2pF1wiDwh/6C+0hoeO57vjdkvfsxv1UH280bK
n94GKaVREYhThIcobwVwBSn+tPTUiD2hZFmjGM4NeY5RiDl9aceA2rgQaRki484biiayV1N5UEMn
NXDfZzfQStu9ApuUwilM7qrPxL2uBXcaYkisl+D2tOZP10sSbiHuTLY1obOHlRs9BWTCmzntPRrr
zbnkpdecIr22Pffq4hG42eipHl2v1JvJ9jBG4+PIwqRwgAdWnLdk0u26Wc0+NyWp77qG6L/fIteW
+BNAGYJcnARO6lFH4NuWtmMZrP+/mWYJf2cTLSZT8Ln8YVogXwpGpCaLb3QmUTbYse5lq2r4jyRl
LCDLHTUyQRbfCIyjxrS1c9lmhXXD2/xIHkaJiXGednbn8fypOEOyfFaoKwJe5nuTiSJd7IaRFe8W
yrlZzzR8K4WLfiKB5ixUMWl0Pav1NPBBZvo9MBHLlFZAldKiYYAYb8phYw0HAp376PqQY0i1a5WZ
J0yoz+PuLHqWPeWppkrLFMuAB2FCb+NLE+CQ+tJpILsBzCLYCy7sDTRt9DM38Nw6VfdSldfXVr1z
TnAH8L0RNp+WqRGz1CHAm2NgeytGew3eH1QDQ6fEByiElOKzznXly64Bhb1qjgOythFosx05ETge
4SAnNSF98w85KS10FJE0yBR5bABFkZikwoEsB0nIkS3TQddIseSWfdt5Bv4hQpgkiuxZTOV4N4N0
Zyp0A/7JGQUz5N7ExIRCWA1/3CE09tySuY1h1GCSeCiPNxiGGnjZT+nR1TA2Rjq9UYuoII7uIO+T
B9jrpIi9avTDsqOosTK7wY8QBdefrD7hugAn83ZVuF07Hpk4Y/FhNLNHUm6fZxTJFAgPUmlf58YI
vBXVYrrxyqFtSyAEtaj98m9FpaM1+N7chw0y85vIvM8htSQlJ20XTBDF/9YmORYRO+HVO2/d0m67
GnomYbxvpmZ8E+Vd/ZPa5jqnKdWveTVeKdfIerKbGu1fi6BzZtPvHxe1jwWV8S9mzqQDaHMNLIoK
31haTKWXi/KmbZOCn+whdLf/Ua9AmrCNbaqLM/OQVr4incGzIzuf1WUOmxQHxAssHqD0q+XJIy7W
nqDbeewkHyaOuQNh8UrDvzgUtTgHRQZkxq8hhsAHtgx2lNwxn2fmMDqtY+UzeUBm9pBGZCPzzyZf
GQ2a65EzBbMZqJdne6JBjChOPNZPm1uyDVTTKYa4VJ2aIXnI8gs9DTjTASDUa8NZhkuIBVVzy1/Z
EttlK7LyuOt/t0tk/HuuRLu7m9QfyrJ9sl/SykQFI8yhzT/H8AuzJW/+dUanZqyRhMD8HgLjIzFA
0ZqFmsSYmmIrhiNu7MIa0DXrDn+uZdG5X/4jxUgz2Wxuh5+qLHS3Tq86TL00yBI9/PxUm4XdJ2q3
JBirx/qRjUvjh18KY61yTmMYMr5SwmKbXhgz2k+Sb9PnOhK80A1kAPtLpSsG3iQnLUYrwrSw+Eti
Y/72LhWzH2m/WpvDgugbfT44Zru6BRlwHC0tmiHrlnhAGehgHjl27u7tlzf6P39zyh0WEyRO7sqO
YX//iHo/XV8f01wpfYrPbXE7WYdwRr5GHeoHmvAtW4GLYz60CzV6dIZP6SSJm166Mz4tL+kfi0yT
3U2pxPJRnFKBimB345To4OwDGtFrf7UmwCNRkJ/j4LR2L7Uy/rgVSj8zkHlB2Rxzgw+cj1IUlxND
MxG807vjFcGZBnvAJ4AkxSxo0wTJobVvJ37W3kR2QsdCfkFbaYvXd1fLsALdiDGzFFeHybWPjJkR
mv3nxKypK2qHtiOZGGFRD6JmP7ZIGJvacNNvjomGyHQJv60bajr1dgE1KLOsgA9/tOJiBr8iWqr+
DYgQ+q09gZv8G/fNXKsMk1uZzL8S0BFnRJDfj/+onNxC8Pr4VCcHz+Hk8p/aYLMu1shf80uE9fTF
Lo7UHcWdrA8Y/2jJ9iCic8JeIzHA1LJ33eo1F6sXCxroskXsO6HEcvl4nu20GkR95Bu+1dlYDoGX
2orChJ5+B1hjf/M6VQt51x+Hx5vFrYEFpt0sjkuQ4U/6uR7ikGB2D7dmO2hkwQ0lWDZvTkLUe2O8
oloGbQc9CpIFiZx27ye4q0ueBDuaF55bTjXW+PVlF+3VEt3JH/7aidxk4FRvHU+qmwIcguFYbkRh
QX54MJvJRicZqvXmNxIXMXfc33/OcY0lsc44rzY2tpLC0pMW+bk1AFp9aylkhzShkcO15C1MzvR8
rfJ63XqFLK6uj62VOSaOAOCIAueTfbS91DAvY4Rlfb3ieHdBFv1dysSh0PKn+3+iNSc/dBNQXMlb
Y8yk/8xcaPfpveaC80gBbfSXkXee60al3cDpFRFbUthcXl+JYRyl4sbN4l3DgJz8Ddw52yBFleKs
xoygzEgItYLv58GX/NgnZCG5HAtCzQakBoYl4VrLgreKuv9bm3/i394OeGNex1/hQCpZQHZAkEvv
lLt5qFzHZm4zhx4eNGZv1dojCrNQjPs5DB+12H8oKwRFaoaXzg/GtsjluMMTVdaTryQCIpYu+za+
DLQ3ubq+L18KEB7UGz5Yrbrt8sDFZ+B4tlT6IGwRSR869WSRVhrmfhL5eLstFFnKVgkIyvpcgIPR
zF/qOWaq75tYlY+rKi4QeMkYrT9+A0zfOE/UFDMzsV/wAku3FBNK7FpeX+Y3nVEjUsB6X6pNKdrT
TSJBpPnt/mL3R6temrat/caix+t5l243wXLyY6axNLZp5/HiQOiUGCPu6Yyc+c5WqZ+pSXHblxfn
Kd3LxsjFXI8HjT9PnYuFx9fWRCS73+LJAHs/eHZfS0A0cGkwCos+bmNI3tZ3tntNM8j5dqimJLS3
RIu6m1plHEndtXdR4ChJZ4t4jxdxup7sCFXxyCrSNMDJchuUk9ebk4L4VJAz5FQKRPcZfXhcpl9h
dChP/+J3kCGyCGBooZWVgt9RGsYfzQkD2+Q6f0l9Df676UKzs7QuMBCvnLmhvpjc92s2MHrpGS8+
+soQmSipaw10Nyg9qnb5PlSvvwdoadRS4nnJlj5/rmG0sr/ElRhC23VnvPTixi6ajidm+1EnsUzn
n7l31gPy1sm6kgEcODB/R/+0MuYtZPgtBULlyW5/kdxjwQprnET3MjSNpdqV/Etq2XbWhBJ17bYB
yiVkXNisJ0aIv9yd+TS3Cj8nbdUALThMPyBDirPDCA5/NnH0PjGMMlaziAhCaOSgiYkdr1wbJgoi
2+C8KEKZHjPvB5PLBVXqVKKvMksTdXqkR8Cn1VjUNB4Tjmt06kygsupCA6MTm1PSuGMwF5IPkwBC
6ZmMtaomHq9sebWfWfrg3VT8Kcd4ISabNRtpl6byhTxQsdqZcxPBlBogblJIJWklRsTnw031xiCC
hla+r7S5melev6tM8POnojM+ZT676ey3xqRhq2tcDtD/vWYpS6/PECF+G2GZFMQQv/jrAoMOalkZ
hraHhYaI4aI+OQ+NMTo27CLLSlfvHGl5Ff1lyQnBMBEYfh1FHZgL+KQpWOTxe5sWfUh0sjvnEDxS
s0zurx/WFnhVvwkJ3AoQxdzHNFEIkOPjuZOOyNhRQOWWj9lHzO4HOUjxyqzq7+Ky60WTQe8lYJRv
P4XTeLiLnnDoJSlUpZs/26zjsUiKTrc5dgTpWM5vUMJ+YTNlcI7ptjLXypiXbiz0Dezst6GA3cd8
vFqyKMg7k5udycQ9bVqnIkEFVx4jyo2xOHUd7RNk0mKcAbnKoObaFFqhXltqgdF2KJEhHVvDyw3b
r6yk+jmeY2mUUAvB9NTxSNbVegIX4irl5H9j2o5dymQ2ZXcrY9I0xh/bhVr8+BjqKgvhW+Et9Mhg
FVmueQPLKiIsEvbegucbc0Ta8tsc5amsclFoseNkHZldWg2atinquNcarlTzyuWFE4lzqQ0S4VVW
XLxxr9XFOVdASvrLKHjyRX9R1eNs4chueIaqz8DNh9/8wQToIJ2SEGLlBhe31dGdNi54y7e/Ftos
gTTC11wMcs0MVkIcHXjo5opnqATdOEjARi578RQrYVaovfEWd4QBRaWSMatLL/thOD2e5ROyEY2F
l2ENN947qKUC53PpgLpf7nH0/UhDEX5dShbN9nuVPCiL99HYyWAc4EswlHaYmJxpHsiSTgSx2Gk7
Mfj23fqEwyl08PiGjupvvMK2iQGQraTks07Bt6PpDWbxAxw853icbXNrp4yAbkfw4b4JRwBNApPB
PGlBpd2/DGj7cc5Z5GEKB6U77ruCmEImti5y3fpqY9qZZeQojmWryuknfrtenDlanXp5sNaJKu9Y
6U2q7dKHt033Xzd+PulXXzQIIi3PXlANxZPxP+6qEoX4oK77WTtW9KeLKJ/zWELyqFi9wPtz6hfS
BCCdYQAnX9dmJPQ7K5tKvbauzAjZ5WzdGggga2jyyF2K277YHTE0gKkW/A+qkcmsxSUgwXgvo/vO
S1kqUG8uhjga6KBV/a1TLN7YDafezYLxtZRMQyORGnetH4QqI6O7CfTQLZ7w/gwwkVvMesQWy5GV
LAFplXPGmZMCj1ATV4Ai/Q+aj8JVuIn5WKP1JZok+gOeM/m2XM3Hn/TMtNRMh3NGnr0Nr7cSUZa4
g3BSMKfdNQhxH3Pz4sioHbigEUH42mJbkv/Jm8ltee4lYvZrN6hInofK4bCUd337BaUmWOiAXXB2
Ez7h1v+aGi/TWVh/zSyYYWR7FrC6vYCpQyAq3uxq9FHogp1ywFyhIsnc/fr0bz155D04hQH+UYLX
KK9yYEt0Hs+UowPqF38BPKnbysExwqqUz+HqFI5dc/dcJx8P084aKSGoFpJOpJNqVTAFktfiaOUT
EJp19mcp0aPszPw/RBU3GbJ30CvIbYj/Gqb2xDLUbI4z2ezsqff1OA5O/psMAp6UhZtZ1FS4yDlc
qDsViIL5NJh7atgfTQ6eesUKTUnM6BOOsTtCzdOtSbKwozO6wk5eeoXVC0Xl5ncFZsitl7B9YpDm
BIcqczyIDBJVFBkH1KQyA+TZRoX70Tg/GngZLOLtNj41CdG3+YoCC/2fJrjzRK1IpdhTuTmQBZQY
R4r3khjkXUyM/LSiJ+uXmFdLSZJLqvag7DOqko8jsKamXHhxyJzah6EVv7+BOnACjGvYDiutTj4x
bUbOx/PIFV4MlA4HbKIUJGAIzV+NzB+rnlUJAUsh+GLn27Tn3hHfbHuIDk4S+QZDM/Jz7XPeCxyw
JAPhhzc9GiZufj2d1A0OT+RH6pixRjKz7dn//X8xUNrbhl3g//x//fVWcHTIOqxkODJYSCnPDEYj
fLHv9MenVizMWUle/+Zfy2WNDTJLRphm9ivOETgUZCx/WN4L7T5d/F0xlemkomKem2TCJFNtGDbK
5kPMsXemP0c4AMnOrJHZN6ifWqxnSxoqOZGIgVCpgtW9Zv1RiaNmE0k5NdWIlf6WjXgGqTZYqOVa
yNUwYeraQ5FTabGF3yx8H+7gCtvjquc7nziyKkCzT55MZkC4fJ+xezzVkZBgsrqbatPSUe5LX8dX
CtA8h0HN+2UnukVjhSG9MpbpWLSj8MNakBGBU2b9C4ezQIdEAMVjxK0mUn39RCAYH9L2vHvU0iOi
fXLcWF1zUr47fGvnsHrQ1Icjyy/CoXxT2FjkiXuDZZzw875r+gUXcyl6khQyE8jwDut5MKp03QhI
gRrbdL59cskccJLD6z9H9sJpAPONUM6V1NPB9OC8CuNKQCzubBOaZy1uM6lCnJIdRtpJWmlY98dx
OOpHwcf0f8n2l0tG+170UdVIYl/X5SypSJyLBoS+I+wMOl0Y+uCZZOjRy3+z1Eybh0+qsx7mPHYv
XCvAqyzFpFISd68ZG7b89P50Q64u1KtdGrLZYa8a2bOuGmm1HWNR1Ix+gonun72+rS77RFj+2HsZ
VasIRXxIWW5L62PUkOi9P01W9ZgPF+FwA5PWo3Sq8RHm49jdqE6NTTkfOnjOUA6ZHJWNB6V54q2V
zEI6GXw2gE3dpNvj8SzUEtQ3/DWhZB3DeeZXF0E0mqgwEprwMpfJCopaf4c1PXNhmxBRzhc3E4o5
zzc0FSqmkHEEXkgd3DDS+ftc8b9JmJ92XgfokMqAHkLTtZMCa4QaG2hk+JhCc5kN2/MiFMq4h3cX
3askwLC3O5PhfX9plNroMQWxkqb+ltzRGYKbwvzT0/hsM/MrK0ZqJrbBk773mS0+C5AEFYPIaUi/
NZ5Wi36YWz49M4eQ9hLKPCVUpnm7UcsLkneC0XcFGKf80C83ukAlvf6pnX/yyESV+fLXms+GEKcN
uPeQEXojOjowXKUBKVdACzbYPB1lB9qaGzue/b8VJYhezZXZy5+GRqMUC039HAVSh/XQIWju+U6S
lmCYq0SJitchXFV1nbdcTA3jUwR73TdBYx5X2WvJPGPyR0lV/3IM4uPWPhSWToTsYaCGD1yLOpIC
bThBlrrVr0R6ZIntzS5349TT1cNQx+ViplrUIZQu0W5KJ/SJlyjxIAwY2DYe8NjAg893Ql8RkmXR
64GVmZy2/iluB5VWoqMxR8pdBJXzE7qNYAHFGEc7opBvhpUvLvJcQ7r+wZo9Gi+KS9gOQIqhbxF5
nKyHKB6LjVKJqj28d+Iev4/HLCWwQpcWUx1ri7cPXKS6lB1P5/h9tnOaFq+xyMvSK97MM660FUwN
Et6HmeHqCHdimQEdiiczrAnI1p4SG9efCwY9uGyY7aI6HOJ5P6gHLX9JzNB+QXhe4ZkDja4HDGR8
pJ6zCOOMXLu+k7t8vhv4vMTxtL2+7QXjrZpgXhNy540Xvr6Jf5kGd+WAHmRk/fd2m/3iWx67xIWC
1guteUcreBewP+5orilvKI0b9c6Yd7UcfVHkrbzGJ4hK87gLfxG2/790RZdiSrrSyIJHzWuPS3VU
Ap4h9RhNJxRi+nc7nCdT0EiImTMSOTtLwslsYfuiixdRQofuJSq/wz8RYuCtvb4Dqm3NCaKArxkw
ChoS1OegeqTS7jg1U0GjrlAmFxFAycAxCAX/rFP41JRTHv96D1CkgU5buux5AVFEUGP5577k8gL/
9zIH8hALtwwwzbmaQPjvZdDLMnBNlUYwwaX/L6i1UzfOGGt9qxx7zxnqx6VQsO34/L37ecJxsv5g
QlBI5+QgdDPiOGpJ5wloeYTS5V/fX7Z78F4WbcClgpV/F6klW5S9KG9whnMjr6RKiTPsmQoK9n7q
uAWIB/4ws9PBVqpno/OErVVlsFZRlov9Ikg0/yL9Ai/BxFHtKBQ50a1gMxJEyT0WDPRmjv0mG3x1
xCXgsddT9Bjzxub0SPgK24eF5Vdu7SQrsll4K7d2pvnvvUtOrXKhL2MunOClaD+DOJxHNnz1g0Vn
M4t0+pkAYs94D1HLw115BxeLocmuDRD/fpMSiAXy1ZW0IArbKSs+hU1dapRF2JOoU9cJNAu/4XEV
t5/pC9gMnBqaJOYsXW3d1449KNuJsfXOnek31z/5Rjce+KtqN6EssZjk8HMt3weQveyGg53zUqq+
ChEeSV14sopFgg/Pi+0Ni/wrvOnzU9ZCFU5SYwkCLo/uhABp5Rt6Bw7lGIUPDk15+pC49DC1KXK0
ZkEfYXEPx0x+4RdL7jR/0pwLkxqQu94Rg0MYNbki96XdLCgA2k4r5r4R/ilonEnUecZpRiELVhWg
DMACIwYrR18KitDr3U15eLQ006ocZR5OgNTTuNR2ktxd3+OTiEIVTcyrbSxiQiAjbAtvkUKqJdPZ
/D75Um1bnmk3M4ThPb/kq5uTIqpKAdwahvQW/17enRTX6iHOR04Tgad8aOwEewyTN/UFVQevnIgA
Bh70S1JRkS4Uyfy/X+TLit4c8Wz3D2pXB90XL5Fme9HG5m3UxoyLbY0GS9MKg9QiPiZu1FLdF22Z
QuAuzJm1Eazu3K23wV5dG/rCPN3ldb4MdbASlGO7NJQHJ26Ohy8jvaEw6mHCkDGO+3dwq7CiS6aR
F+wLAzckPwoY25kht9aqs7Cn8Jkil3iRn5j+0U+XfFU0Np4EPYVvLUyHDpNjnA1gq1JK0WlLAs/h
tBK0mwVQMIy/xI6UUdKGJl2v2t45AY/Sj83q8c2zUw3xkWnwKf9kEdubK69nZtB5c+ilWIU1A7/5
lzxOxhwHTraP3eVcM3OdyVZCukKT4LVJiSIakCR6wuI8yIQ9f5FSH82sarTJ1Tq2o0xbMKK9DSB3
vRXjJSdkzFC4ZZiDvpJxwEZjuqk2GkKs5xgCMrJVY8gdFW0Hl6EQ/7dtYzxyDkpekKd587NJOCu8
5jFmTCBFoAudsMc0ejYY4BfctTy3FWAAs94YsKVI8g0R3Nc+YBgivnM2gDgx89s+8vGMjzSG3ePx
ayvzLMpzlJPWgluPi+L29G3XJxCBwfS24S6LYDli6XOvTh9zfzyJ/Mt6XlDyTc/ja1tGRU+ndhx2
ExsG4e9qxzDGQ6UYvoSStocvhHvBsW6a3wnlHKDACtfCj6VfCTBsnW7Mmv1eAsqvbhPyXAsrLswj
gaWn5O6g1nteNEjBkttCoaxMcCPDE9h7uvYPhADcZRjBcSUIY0fmhJZ8BlCjYbcJmSMpS51P4MZp
OkucjU4Jzk2wjv0n+82UjBLlA1rqv5O7PWO4DIvI+h0BJ0NFS2vQMO6O2m0n5S7gSzdoJLu1RmAx
o1iGlfSU+Mcu/I05ftQD/qIkl65FViriejVXE85Q20dOcPhq5ygT7UtJV7TAFF7v45KDuHDbjyiD
+TpD7NYtJYBa3ZJiD4EroJOsFdnimN8AWg4r+TGp3P176cmEYpGFrSN0vL55iRk3hUBE0WRSShaX
lU2AnEbZkAIzj9fLg2y5d8j9SKm1nlGdJ8Exwik+SOj6EOZ9veMBcp3MgfOGIOMP7v+Kc4ZXbG9b
XigAbEoDUwNZqc4iu8RJc79zU+imchfrvcL+hreDPxtkzCuZPefQNN9O8eEJrKfF++6oIDHNe2ui
dMamJMU1oArsg2+Q8zfIQ6TAj7ikNSW+xfwEXm8EFd9WH7R3+U4NUQ3ISQ/vW365upIVTkw23G6s
w+e/jWiZXIZcY78gH3k/PzNIjxTmRnHJ7lOAsX8aRQQbDsWxXALJVe6czK+IaHHHz1AanQg+oKRq
+pvIl2kLCorLFXjSTcRO+9E4Gig7bP/UvZMOUeTwKea+LpeQNAr7uGMOBHRKtDFhe2/Zo6TBVLsu
xw2i/zE4ilo0jp1L+cJ4psi0HPP70RF/ac/iJw1eu4GKBfPshkqMamfx0EzKFJzJh6Zc0Pvty4Ry
so8NnAP/Oq2AK/IpSXGNUk5zxtwTII+32tQxlpRgfWLrb9saqyrN8c4XSbaeuViVwwgySLgSCE6o
6++xg8LNmloeNe3E5/9NdR9y2twXUgb5ZzFSi/azbOaKW04ZIzu5EOx6tq+wiEnvllvCumZouwGx
PacXdYitm5I9po21gTGMl422EA+zLem9woNHexaKQcBCnmKE7zQY+H3gPbYiI6GALeWYPR5AtbHp
eX2RLnOQseafV4odulAc6Nxa233bj8Wr7Xr5DZMxvnNm9j38lpB327k5eZOiS8LYo+Q6VqOgFjwQ
Ej2JNpdRpOAZGd7vGKadZhtjHGty7w4xkdpyakbU06dTUZwRQZOmtOkYTU1h6gUIyxaAbhsQs4Vf
N5lzGBqwKAndL0LLs/4TdlW1R0fle2dGdFNqG0Xqqedbw+cCMaZxNz48petW0s6VyBkdVfsVpPps
uGtq9nXMlZJmFMzr9Sy1XJFy0tjVP7FIogldFqw/pW0LAil0TQmV2BElajW4K2MpzEXInrRvt9xz
KP++OPDq7QMrOqsJcpWCJXeJCxNr4knyqufQDZNzo0bqlJduaW4BhquMN+rxU43WnCALXCl8+1lb
LEMk/xjcaKBKj1l5cp29B/eYRa9DsF/5G6U+Gdxpwi6/EJ5C5Q0wSZr33ZDEYoFbf5j8ZP1dxjEp
Zjow/u+pEEpn5cG/Jch/MxRDNaURaV0/hAau72a0wyUIO7Y76rswlj1HSpk5Tbg1VD4EOO1VzC1K
Hs2Ia1FHz6/tl+foqDbUzhrvxDAbTBj89OzMKcd54WsiPqW01iLgUiTBFQFrNeL1FTahP2GAYq2U
kqQYxnyefB9AYnIFQlpDlE+oDwfhJkza6P4UplKcGz/Nu1+7YOinPDyo5YHwW36548i5iDM6Lj4D
sUP6HE56i/w1IpVhXDjyUEhs4Rj/Nc0fkR3RlDCZaa4+C1wJ/CgWCuFSF45Z4GrfxG9tZEWmw8U8
sk4rBr7vqr7xrF0F3qTnPu4RJ7KY/A1+Iax2wOlq9vRLUkJYgYLkKbdlV8Hj1WGMOeOInDK2l6gE
jmYg1srCUB6ZjRDbhrYm1qrsUhlO59w1O+lSJF+Jdu29GxlGyvZhUB3/Pb5KgYfK3vk0crWNsKvQ
r7NMAvyhKxbWcgzNDXCwpOMoEWEELHD0Erjp4G+Teow5Id94xHX8Y6INmDb/mjDYYm9j+XMJxUK1
ZDR7jsqU4rDvytTd7PXnAsXZk/C7/UYC5oZbQW1VIikwGV1Fw3z+AJQpC0aD8wqbvDzqQG1VmA+u
+/HH82cXyeCfQYq4vXoNL8UYftK2ifx/V1zbcWfwc4yR/g/JQPA3wvbqJYUw83CnsmZ5jmVJjyXv
aTtGQMKKmBzwioSDtI5IPM0K7UDPVfP+XEILKYkz0UFkBwfI+1ZXGmLkCa0/SnpGSA0MIihhqbFg
NkcMp1uT3FdKvARxFIyyYfu3CdRij+L5XnZjApZEDa4YePQCnR7sXTXemMm062Ka0OLpxGXE/CZK
pReSnfRFD/uYRxQZgqlxOQTu+zmwwTNlyTYQx8E3gqfxMFp/ZPiEWihCRSdKxwVPqqhU3HtUqI+8
6E+nMGDlXiJ6rr01oaannqYYRsL9VM/wqM+JxvLphYTx1pvFHmyZrm/B9k3pUcPPy6I8XUXIXr7j
9oiv/wSbvRx+/Zyhsj8IrTJkvDCKE3g0F5R30RFmmg6j7M1uE5yxYk8Pz9N2JtA4X+aIiosfyXKt
utIm/xWSlPXvq4Fv1pTN9yQ+wgcgQfL98nZrbyt7WRbf9Q2E5KAF35kX4eB58tXQTrPQAoYuBJOI
GMF4XZxcjI+/MAP+5/F6QQPjtj59PMHhhtNPi01fnzg2FUL9DGQXGRuc0nGsCo4EHtIyUgitE3eU
ZUsNkGu/uT0vXrC6bTPj+G5vc+LvUX7iVon81cr455LzMSHwK6DHFi5ONV37WjK1xec5WsbhdECv
rMLvlK1RDWxxd/5zC688X2YdBspwE6HUcr+UD4EE47i5QYFuwFrej0xehdlfI4xJBTeccoEn1+HL
yFBk5R7r5wn69ppLaHCWYRkiyX0O1t5ZtT7+EuP3xAFermkAkOG4cSa6MBWky/oFsxFNEoHxreFa
npv0lkBDjSk74pbpaPyFkTC5S5j/WsIqjg2PEwJE22lLSFvWsCCDReUCqf6ry4zr8IiclPZmwBSr
Regv6h9psTnbh/q7klj4kEoc6xCOsHLEs6BmRpgjHbMUezYHV7i0koyDGupLVDDzQtTXGRy4J4lk
ZPukiHgCkoZ3KfoP6E/tpOGjJspRI+hiiZHoge/Cb8waZOxyWaDEAhaALsaeH8/C9/a/gA82CJvu
Nyqwr3ycSOEjeMSZYu02vMo6ZATAoJ5AzyBR7X5OFMyX3akxhXhjWixc7tlxV6aHEE8HQhWakSDQ
CI2uoTLdL50eRRRMiXtJv94vuP8y9IfoCojVPVkIU6LZXHFJR1/5y7TW6Qzb+kAnCLtOkkf5JAq7
Pid+cp1ipnc9pDSe5HeOFpaNwaOvrnF3Z74X1uPBPgIaSpIkppoC7A1arJnuAsXtdoumt0FbWGV0
UG9y+UwGS3dr1OmLcpXRULTaceArpeGwS/SgS7s8O+PFrKHkJqiTjiTQrSWGJ3Ud9c5qWt5qC8O6
5yVpMhmC07BICyPPGBuuR4JYahRE191UlG2pf8Qd22shfGsKTHRnrRLQAUikmBTTjxsby15PUQsQ
nxDavUWFoJ0x1fCpzDKZoXiKABMlEb8nfvfTx28Fke2NPP0bhiLe65MpQWlhAin2Onv871g8HoiG
J2xrRjfBQ/3VVrKFYa4lw69uvWUK4wxUhPnuGZp7pu7MI2v8Q4DNcYYrcbD4OvBZr3tCZ0udOc1x
konyZQIV1pbOw3g8SbQQy21YVETM1CiIP4RO2D7Ny8O2viqTbJ7H00NB6/qjAyKDBcS0VbEmayPN
dQv68ZrkuN8eRCCnkpNR2XZWmtNZg7VllcOAB5m+fgsph5DkVITcDHVNNrxlF7a73E1bjK7/38Z+
G2CmhyVbyO7Tkg9Uqpur896dliTHGrsAUaYtLo249hQjZO6qqlf9se2dWH1Q3Hy1eViwBjuEmFPx
PDtJdWBEZDcegQfGIBrW4Bd/OtqIfsV7NPTcJql1sXKWjIgWXmDIdOv7WovHnPzgNRICPkNA6LxV
2pBLHaIgkQsqW81afTjGciddxvaz+Y1kxHsogQpREe0F22zZOdB05g4MX1Ml5Gmuq4OS0DGvf9Ke
J/uWf5bhq95HA0SHlkF3amTbjYijvCG6sboanEMPCRbKb0OgJnH8Vm4I0YIovpZ47ftMUoI6k+L3
dxNQ9aCDBgskOHjtspUAnGLVBNUhK05hQWx2nlewFqVLuq8JhfEm+W4H290Rbak/Ud9/okqKpftp
ggSEQw1bGhStVC93UNK//63Rb3VdZoLRnQ+NznhxJCMPeCvVC/qBLU/vii7jxS4dPjk6wnKS8hzo
KF9e3HHuTSm/VePMko31T90MclqNWBZ+yWGXec4FOc3s8maLhTisWjRUhNeGBh6R6ox0RimykgFp
plMlHspVT3EzDOHch2UduXdyJIn/KNMl4ASqnDapSJftwHroqaoozLlbhl6nCgnbrBzkvlh4Ah/w
UUIftRGY7CPvrFKz459zdWFi4QDzNJ12SFTeJQ1ap3h1px/KkK14FEe7StmVaEvsa0BGwqbTnpd/
7sZFZ1+Z4F7gqGRfiOk4QzplE7thwtOqW9F3//dCWkE2y5iuDXbGt3XmH5ZvyU4wrNLp6zikgPkb
u9GAnazYWcy4Q8cO5/j03zjhvIGvTViTTBci5BdXoWm43Ec5IUFHELvRhToVEDEQRylV65XmkQp4
CJ/xNMLU35ppxvTk4VwJrKLtee6OnXl+fJIn7kcFcg1TRyv6gYrDo5B7iZA+wy7ryYAi3E+qVHFO
E1HBlwdfjOBAIOKrEF1YGxAL1pHy2zxaE6XaoWFGHl1TxC4v87jIJUC77a7GQqQ6QZdbs9+u8xUE
3JAQ1kE03ggoNVgdPU1u2i8bopGkuVxs2L+GX9MmfFVl1KmEOlrR/2ZrmUaZf4a1gzfGeUBq3bdx
2d16tWygbMsDxkDjZZi3Z8psCBtVajyZhSx/OnZnRITOVepUiB0lj29svqc/mb0UlH96yGIKPII1
AQL/jwbF6Mz08+5KeiqBX4ITfsNLNvyxSCalTPgUCsZiNHmYJKX/IEIYpUWsXXozMuSMy6UZkS0q
nmxpDe8/+RHlud+7bgxrpHCJPd2IJcoJXoTkpmb4J78BNPf4XFzv/OAtPrlZ4euULDe8oTZOr4N1
cliLegUM4XM9b8CGXBC8NEZLGDjUl8s5nSkTBjnDsd/iTt/cCgb3k4N3BQjze5Nw6UIQw28LyxM8
T7bLv2FpvKFP/3fLnV79SIzx7WJVX3kVsVckNwAc0NqsgmbqjRIopGl+/FDFRT5fO7ICRYyAzCAl
kyS15vgPYIDIwDz/w0ZH7p5Bpz54E2GqyeZc/XlvrTwM2Qw7upD19XhUwmzcbov/FBUIxIcQSQ3m
UQzC+J+mYXGXPBBuplS8pPZMatMP5/j8ABRbSxmxV69OgKpar8wvenTUAlXWwgEbiNT2BiwiXQ1r
BCf0gUsv6uW5sZevnR2WlBVdY42cNgFyZd5X3R7z2xF+H+jnD15+9yLuApEfvXeDP9bO+MBwEKlf
OrP9p0kxqz4qLbulkIaQvjpdo+8yr66BkP2L4EWoHxcErSL1diy9YLb+OQIrhhz6A4nBycn6hUee
T7CMf7pOAh4gsjPYWZBXat+nYUnmvbW+YJBVANxf6a1pmtq2N+rMJLGH22/v4rvqEN6MunY30IAC
VKoWtBtBiw5Bo1DMUAONNqQ1K30Wst9M+FajOnWeTTyKzS6OjihcXOnaysMO8hO60ljX1rO6X25n
AhTL6DTacz1NupXsgL3qEcTsXdlYKZbw/QkJaHeTsuZ0n44/CptvyvCQV25OWTwlic+Z90SuigSR
NkuLyVpuSetWvlYgFMX449DzN7YTHnxJf/dsGY5t9avHN5ZYuvjKHm2eXDuEfFg6zKUPHAqT1fqv
ZpPyN3DvcoNyo11sI/3VXbwf228wMMI0amLRu6JlIrl1zCA7v6qJXUPGWxjECzth95bIZcuvGzjF
AdmFn+toO1mIff/gxa7OxsIi68n+P2oQOTbKbWS9MyDbzByYtW4d3QpgSMtrvHxuHiRzABunm26E
bbnMbNPAt1WRd5URmmsRgAePYDiq/Hh9kZFBkmpE0gH7XSVgI87jOXr/Ih/yJHK/Ix9DO6YxR0Ez
ZFg1lMgL0BOvu2eAKyis03sW7adaJk4uKak9oqOVm/OJ8SX+Mey5EeIZH3KZ9nHPi1xCsNvUNssz
d6jOUNUP0tPGxwLebFj78mMmufKttbXk/fH6gDijHRHE0U3AsLnL5cz1AlRKK3LCP7btt0GPggVG
pxXIXFUS1836S7+zeFpCgKo6tygl/cumB5Xg6O+LJoX7/Fk3UNiGLFlkeGeudeAYxlpcw3n+NsBS
ImkzRPgfQzdA8iWnCMLvvhV8eYUVORmp6CYHhYUPGpPv3uh3INYmobaIoMMqJbOadnLPILY1YQ1X
FRWiwUOM2AnOkH5z6cgCdqpssPwJVk9d3yBpXbJ9jyFyMWPKuZ9LqF0eCZfqdq7It6WGYoTrBtHG
A5YTuWxSRrhaVuO9XlPQwNl61ToFMYdnxpSQN4n6NXZOJ6QpOZ5WQdVsCV85llZ6pgQiPf8E0swF
YoSzO6tLNChuOGVUECn/UhR8WX3x9LAqaarU9ATEOP49cd4B9YessQZYqoSlmpy/rYwlqYcz8Q6C
LlZIvXfeI85282syntFPErRwgUys8xRMa6T578i1MoymDEQTgnRjkDKTZJ6aGj/oL7CQM+3hqaAw
rhmdS2nDYrflbWNooFLpW2KyBa4zsW9ESLcVtyZFawBRwDjylXFthgRzthe9w151UgvapM1GiS4b
y71Vj9FRagY5ItkQV/4bCHGqDfuBIqVGgNMzTnQ98kPSpddrIziGGqXI/B84cZWIXXtP+ZUNN0aR
kjoC48SMl4bWBxEt745+u1ZHQ/BTCaepgvv82g95TQ4AhNfA4p3TzEBVvd5/bQG7JCZH1UkqKBNY
GG1vG/d0F1Z4z8l1uuDqwLGvPV+uYHsWPDlNKUBqSWTqggzTGflFzWGbieSFKSNfDE6ZM/wzkAdB
8TummIQ9D5/pInoLejcC4OOHaf5vDgmceEmX5sQ5BPdo1Hsdscbye2zCn/mTEF9jQCnITYc4Kpz0
cRCd/1uev5wLP1rS3lucSSAXdlgitBAPLtSrSL5Qvu9nuMO0zvnAjXUZA54iEA4vt81Hy9UT2gvk
2tf1MFDlvlW8JM69KiDj16iuVjp1IQXuhkMOb3+BHWsrUmsZoZZZ9PlE3nJUHkmQLlqxYj2rU15n
Y2uH6REtXVpf0fb76Fx1KQc0GdYjGa5AVNJqaQAddjkKNLHVfYrBm0tfhdtq3Rfa7Jf1VXKDDJEA
XTtTFDy6FItFsfgVDkJaF53+eiKAxQYUTyAHbKozA5fvyZyb5KGNR9Ya2sB3vWWJtzBtKsBuIFzP
VOnvtr1NK3wM0v5x7zAHHacS79eRPHbpjUYxxtI4ku2rWNtTwVoFbIqfo5+BeoU9I10n6UCXXizi
HrJ5RrevSy7fAOHhnVqbI6/XQmRSjeM7+8mckhUnvIRUz9Jv8LLCeJstMACVPmVF7dbfyq/GE1P6
88ZAMQ2YTsXODZgGgEMfrRaEj5q2mGSHzTqxlPd0lCOmbN8o1W2cQwml5BcGVgF43GWNGfz8zSje
dPmnX9m1kvfOQWknkarhKK/VHLJmscCnbh88DmlZYYzGmsvm5fU/KujXKsGbxhwTu21T0+9kV6VV
qFnZ7YyjuowNFnB8v7mvCsGkVYN1McfG0GvBLHHxU+Yg2lmtcNpy1BmCce38NvkPk/L52dnqrqJy
TmI+OMYHP/Q+/3WrPlbttuZSis5i1QmA+SVEBNcnGNAUWPXxBEXYTzM+PNthCxgDHfhKQ3rhQ7qX
N2avMouy/gEqirtNM0F38Mum3bi2S2Fafgkbvhnnxmalb9f0sf3uvBYIg4SEiZjr4RO0C/LBX30a
vB3wt+7FVJNUjVuuhQRCUCj6LLG4Xad4NTsK0oANDoa/DZJ9QBC4tW8aj2sRZoWAGPIpULt9fffQ
BJLyX5PRw1GGo5XUo4GeTGd2PZYTxkhT0/kUJ3G+BAsFdcHlb0eFfzvBOR/ELFMYh4XhsjvX4KlD
WBwqs8dQ4MgIBWLortN1swUPRDiaYedynPzsXLyB6BVyuVtkVkzhVGdrIe12v1kptUDgv38n80Am
Pr45OA+zAT3/afjn4oHm9Fo/nPtllwcSScaDwWqmRXOFrbYePABmvObNfr4MOd8jkusLgo21XTit
9UF1h+AWJZA+FacSk1ePd6wgCpswbAA5t6gwspjU1nRSUVUX6kq06ZFZKOvEFCurlhmgTy1qs3uq
lfqaKy7ktGCZxRRUYVlXocj6Wg4FCGa1Kfmu1Bbb1HmThJksU0AXd60+REPRxQim/hZkqH68RnoR
AF1fgUQAC5fgNOuc/DJD+7fk5zydoqEi0nI+2daYt2bDy5M0TYxO3Zxj4QgJGmVORZI0OhG7Ey/l
IestsrNUI2Y7tFUlrw7y9Ae2Td9u2apkVV+mbdMIJFF0llAb5BkP7MLVGrQrc75s6IWChgS2BxFO
8JHWMhLWGI+y9BnKtm2TqHURI6d3u7yCBJBtjH21ryzInIoV+YtPjkr9eDHf8kUOKIuYj1+P3hjg
ojDYu0fJhB84urOks0aX4yIfZa9LjOkalvF9sR7vh8+5VotJm4yk6ypaGtMKnH3PspkR5NUNuEx9
NUElle0cUDR31jGCspqXsK18LzZV6WzcfVWZ0kHCjJ0hbjqn6ygbxFaO3f0diTVqpLw2sA8qH3Xo
BLPdHEdQ/rNyWuY1aiVuQFZ7HCheH+XIGDLtZZEjdRHYoXaYJoyQTMf2icttNWJTNhfREBvm0X6H
mobti2EfhUX7W/zTElNeVRenHPpDxnBqtntcc5VCMX1z1BPAJim/ipzapBBbM2PSflYQdZlecrQF
ciWQdPgo5Vzo8ppqQEHi3bsOVPJgQP6kpgJsTR8t0NXb0GLZMZaay+vTPFPpr4SLWMtuf96dUpiv
i3CkNx+9sAeWKnwvqrM70z+SbnU0r6+fjzrEnCH+I6M0S25ddFTqbkXPq6RniziNK089WmfKMGOT
qcK8PA/fDT3Z/pDoVw1mAfofmUqWRx6piH7rAdrpLC13229/3bFXRWOV+wCKRTgQjWzD9AFl33En
RszP4AHBLz/LJRCf79UkaBBV0CAQerhNJ5hGkCTbWgjau1Kw006f7mrUBFB6c24JySVjuAFH2Bxg
9LmIoLaGyG5sa409JnIUWqeLXiNmEWEYBei8XF+pBLboa7DKw3sDw2UFZcgq3+mbxH2p/AhIB9WQ
t045K9E0rC5aeUfE4+8ZU4zU2I3mpGaTHlPErUFbsrlvLS+Sqmi0fDSTeVT+52pa4NGf3Ln05cMU
ZTL3KorFUvZo8DIxazZ5MRmRlVWNsY7x3VKDTG6iDrnQoqx0OmU3gmd1HyUUhaRaIp+NcsagHH1I
ew4csRsaE6SeyWCQaa7mIp8IW69u2GVQnFTEiZ1wFJ7goWx/BekNK703ajxSO1S36DneiwRGaKtW
I+7vaS75F2URj4kdpaNkMWU9/rtPgVy+A5T9Te7YcFlwxCEWVB3M9k19VMkeDpW3E5gfmIkbctRd
4OXkMzo6nKD5x2CUBeGPFMni4N5kZG3cJOq/apSXkMT5f2cHqm8uIgHv+01N8Ngx0tXyQ4pGuUZM
BuWxYjO3blu+QqKqQIOnQX637KP9bWyJxjH3IWhVFMEdM0dfKw8OaPTDTpOJfsgg6bdO3FQqfJGw
we0YBcF+xxTuv+/7tY3+1sp5UVbNtjVE6J1+fbwGY+rhj/uhTxdmqsBYcoJRJdocfmzhU9tW5CHi
26o0CDiVa5DIO5g53s/9pqnNREnRCu4CNvKlm1vUaGilbCS1TCYBra9y/snTDji+tQNAX3+Lzlw/
3ofXkX4+xA8MPGeVwEWYGFDANu6ask9a8rvIT9VG6qxYsQV/U/jrHJMzKSHscp4bhwXZpTzVQXKV
dKSOCE98iUI/RO7ValJY8if7j6GyX3VvASOP9CEyR/kYJHkIp+/sWeVyD9wJS8+5wM2wtPPxYdAA
T6Ve+8bE3Q+Rp35i2KiD8QkUNM5cbRoxydev3kyoEt5u24VeZqU8lQSF4YxyrTc2jNJnj/Eu/yHS
Wh7CuU5gyIvOvpwkBFflZlkCfmw8FTpK7VI0PG1pJWrDGnNWgdx4dAM6nWe/Ro4imURFoq0ZiUsq
DHL27O3RPW/OGALoi6BsZhFFrDMgke+W309eLVlACVEOWyyZkyD80lLRIWwk4spM+dYipiBOxV+o
FyN8ReZJoMwLRVyKpWul23KuuroMQjB+ik1tW8+91WYTgXcywCQUmbLynFq7ij59VNvg6ypybSez
CKVoubMuP9CWE6X84hALZ//9TU7YzSwgz1g6T+qZfHpip49CSYVpSnVIWAaPiYF7653qug5VIC0z
4jrD/Ab+pi4uyNhwi/DOoqCE6gO92ca54O55AMbnG0xfOKPj4T3fAfl93KD8nMSoAHPWZVmsgWh1
Or0FLOxZxhS6hJJvn6ZUrnePCT1xXO9fJPoE16szW5x9jcmuFu1tZQGZytShFIRA38vAjgPWZ3Dn
xPYNXhUC15E1nHDiwRrQ3nDwoEUt4ZKRn1luo5U5ejcycotOtReKc+bhzWnIETrPmgbC/nvin9JH
2X8FR0P2AVFUQx51o/mZbfbpIwfBWVAiEJgpYWK1RgTSzLmr0d2YGs8GE83wzUmGWh0uRns4I3QA
YJrAze4iiJcbKZ7WeGUcWZcMkY+eLrh44tKDUY/t4qHgw1KiJjCdzXgy7/b78hYl+n0/FlLMJmVL
FkDgW95ZZCBKdeCPmikiOB1KXYhDjU9XA2rN1hBcql7eH93lndN/2Ig+tIBdhDm2ntbdYV+SMZfG
SbZAvfS1vjFbGdwt4wMIiJM+YPJvfph38u1EXl/VbgeDsuxIBCotcomFSMA8ljKrnPdTz2BjPWB/
Glx95sXEMrM7VqzJ2YRhgtGoMc/ikZ/lbxcSqjbh1CdpO2ql48Fyo6zxYr0XHMwmDbM5Y9ksePI8
DJwU3Kq7FxJrvyLcbABobKSgTBCFEdcAU3UREBEVndkCR9p/jExaRIdVQ9t9WZWrrTeTzypANkek
y9WHJSv4PvaF4tDqGIa/LgSqwJvSy6/PhVAmUSlKf/L/etWlsEE3Q1MlTh9GIdzEH64Q6QlDNrrV
qRxSZjgUHyFEoB73nS0JOfSIpL240U0szJuFaabWBmiS9wmPbgjtGsOQUWxjjYGsAIDtDJEsqaTs
yc1xWPqn4AKgHBZiq8HoxftfkH1YmEML+Kh/LYFIsatasW1CQ9xahrdIS/kWdvJvvHuldnH8s4u9
WWvgDXKwGLGImJ4g+c0QuvFAxgA62Kp7yM/byc5oC4a4lfoiYEK+FjB5H9KKKIsZFsTP2BoMFZV7
zCBFTL1AgKSTTHBCG0CgAyNH0bmNoJr60Xuy+tWs6CP7HNpb18kRdKccMT19gW7ju0CCiFH+cWGS
tIRFSmLh/NQEuVtOVkNROG6VRzNxRNxKYTRL6QS77cnB3IeXm7R76sVtxYokNWlGFzNA1qFuitka
uCgwZLXqH/jKy1oxa8gfmoCojg4k1anLkc1YXeo0WA7wWzIB9L7G8Va4IJefok2D8lNuGNIZLAVW
NKugg8BQ5G19ihbzZ3iaJ84D7K821TYG9QrPLbqq3+opxHz6FsZJY9GOzRinvOLwX4OPi+a5in0f
bMNG/N/amcnESPavwEEoCbVXfbY76YmUI9yQwO+nrSNOorfxCO5bC3bIqa0QvlOU+8CkRb/jY5Li
rZYUSDcaYAiIUGvxB1Spn+wDzWhint0NMZkW7094kmmSO/k6Fha6ThPms6+AaEc4BS+wWekjRax+
LfL3qB8zVYvAI8M7CVrQZiWsNi7CGsr2kpCE3IJYXC3JlrFiygdOkIOzCw==
`protect end_protected
