-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
soRiy7+m8Lr0R2RDgxxTj27EqI/MM3dv4SgSZ0ORv+7NSHn4SdFJSCjYjVD1xbQvRuDfH7pqKiLC
uTRvCer5Oa6LUnbO4I28BECmCTDviUKW0gOUdgrhlk+DzMYsMeQMUFUZJYJPE7bkPRShv+Bw9H+p
tD/CUquJn/nNAmkaY3nlBRQ6UnYAmNK0YKdVgAwZx3NS4p6cjgl90SVPGNgT6noHt9j1eesNt8n2
t911HEHE7NaE1OahdJRiR+HLFOOqLrmRgmokY3KRg/+KS+dDV+EY9BTKEjOiqiJoOiPC2RXuPfJj
lvow6tzqs7uSFFLnWYXCjy2kH3L206o9UKmpsw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 56272)
`protect data_block
k+NDNfc9E5AtivQdK1De1nsrULcvjo0lKqNT+wC/zALKXddsWrthIu6suDGZHGeDpjxsbh7w81B1
YpGWMzoFaUyOmr6oWx9H48k3yLrMyUZ1cz7B+/mD7vBha3tM2ZsKaxufj0dBNr2RpxTsi4Mg5adQ
4+S9aF4Dymecz20swYELogyVplrSbPdaY4y3OOpsE8Mv5QhrnrgQRCQyoZ1WLAB3v9qwbzYlz/Mm
LLWTQyKWRI4vHYE16Hj/0E33qJkoZNTCLpVHx24ctUzeCESKRXi3pyf73Lpg4EKXXVCzx9zmpyu+
keAogsuW1UlZxTDzRxQoTsiC+DBWtA6C1FE6Nm9LjBrZKUMgIll64gJZkcePyaJ5wSISJw6hdqwi
iOZLAQ1WFUFPazP2cX0c5U7U7jY1o+RAGAzxukPUPE1a63O9vWSSO1qRMcXQV+7LFJq+Ki6dUaEX
rkVF7Gy3oGjDe9RizGVM+hMG+1Bx3g/PTjSzVEnwetOhK0tXdLM+hyMPIaxTMFJDwoqluHry8F17
muLwQ/AQGlQ0DvBEAk8r7W19rJg3zL/z26urx7nGlFXmn5mruF4qF4ka7Ivg2kTyz+kcOzp5OA51
lZhzp2pZz9yOHNw/5ovNeO65FF8/irpZiEB83n5SNQeu9mVPCVIJNd/NQIjIHyOBf03wC4XWSK4F
cK8OqLVy+aVK7+OFzIr8hULIwph7mjphPIki4JrhegVmPjfm4aREVSbyxVYbfnnwFzIzuYQ7PdEo
/pVXIl45mvUWdrZ7Ieim4kPnAIcIhaKZmECJams4DfVKxa1Bsp523XWKxmkTI5GttVmMl1OL7uGb
kZHpBWeaCInzLbVQw3HMVuD0SqrfkaP9fcr36Sp3RIOxIEYHZbFpHQ9qj3kByP8KX/TcOBVolc5X
IYCPur4PC9stU0UZXUO3gA3zVYxn6yID84cfhxmNswUBHp20WU9/0MAeYDkFUYg+lARH29Z4QndY
QKmAj6AVdVaihhvNmD/7zqgZl5pl4MYOQP4BbF3bK663t03Q+UtNJfl3eBQPMJTqpaZExfedHTQK
zQH41Np+5EpqCrwXcchuvMeF0Jeu7gCt0vc1zpWiTgrY7dtDfFA2qeDt4QrbbhGEhWvxVqF96Etv
lqVV+9wfwqcq3p4LxwUmxlAKfWcJgAYpdcWVImRPyGjRPsxeYy5UH0MjPaCB7qfw8084jCumc/ci
iNZEtET4cX7dNuPU4O63wpB2aFniaxXPX+8JkQ/FeR48IacerzH0Ofvdb0alDtGjXkm9oZu70pUE
jstR9oyhiY5wCR3JOapbS+xXK9hxpTKdq4hNcLxdj+KReaKvKVha0PzgdeYHHYvpuVY/E06iDlfn
eIH4zBJxqxa9WpqpJNUyGMr+tuscbVczofXQepYhPfhuKCD/p9EiWhwMdbRRDGbdzfiimh/DWOsP
Ry6yO2L6RHXDxRVPDz212uIDHRLIFiDkgtSkfSA5np2nbuaVYKM3E75pvvFGRFLLYEpAc2HZVvOi
BSV4WfJKtDEvwBTIyn4jDnQ4vVApOsOYmiQg/DaNFasCdz51+8qPoqT6BOH4PtpE2nvk4Li3gop2
GgtQgBBpP+DuGjiff/nuFP3uBlvgcRUbVzlfjd9H6x3/EKTOns0TMDfB4LgI+SzN+M3I8ZevphAC
ul+jXbqDiPRjGzXTBwHnho/c5Y4JBxy8PVPydMLOeJNZ7X0l6b9u9F8mVGDoGaNtZO3cTjbedbcg
3+Q2k41oDjqC/3u0QSMyyr4umTSQGIyT5RyW/JIdt3kC+hOyAr0S8akEHHgoA31opiwtKCbvInmj
3j1PintOGaQa7utfBOOvYnIVmhoauhs41JOkAYgIQLTsXYtmKL9nQfIWRP9+Xva/oJ63htbe3CWS
R2/qCEckY7C632QAdhMHa+HkQV5b9rPC2qVViFY7tLnvbbSwv7K92Vf2xh+sbp7+QxB+2ubh3YLi
Z2TiX2uYEF19lLfkENVHXFek41RkmbWuqPcZM3TnRLS3JKsg4hHU+aKdiUJ4iCyAO3tR7J4IhbU0
AbGIfyT/ecbYFddA3vrC1nWHC1O532OKUhLpbKFk8gmwSUHxwIXKfKUJdn12e+GQStY+TE+yn/WC
9Q7SOtj9chColIkFjhjIPgGzj4zLYvMr2zCnlfVyEVu/dtWjSs9xOR+9XyLevQKj9zSJkS5+kJUT
lv6dSp9kgjBttSK4ts+WPUcvxPl9j6gviHoX22MLetJItPD+OWadMXzi88f9G2WXB8DJZquYBROP
NFn5rSC60B3dWWMoFK2NwgAQZoozmuJcxQnmYLOzG1QST40Qpx40sU2JUWGJxKxwdkwdBaoDxCJx
BQmD/Vg1wze6j/Y4epe9T2q/Gy+8z61Zg+ky2J8ao2LSAHEIropbuM30Reid/tT9NvpeNdRzU8wf
N5EuDkER+jLE3SkBVYGJV/NkqPAJjsez24x3qUBz9dEB17G+q3A9HsctV7LV/sphJgIzjqsnZAU3
M3kalKAYsMu87h1dXpOPEoQ5Oaw2Xn8Wp/Usuznl4CHGkYMcdWTDvglXEnht8EI9wpMiHDkZpQuk
2vZs/HvDUaJv5MleardxK6qmcSEQXU/QArUsfomJ6lZLMoHbnbQaNtTp2esSP6Mxet0TJEdVrB6Q
Lv69jkXE5zAkD18WZk9wIZaCbHQns2RYrLgqJqb8QT5GwoiNfFuUS8vI0+koNmrtVJt/53XuXoyL
uNb5ia/CLcxjgiD9mk7kNpxj8zxEgXRXIEd1pFsBnepfrD/njjCoPOx9oeCY/OxJlbHJQ9QUAdHq
KKslcXQHYzN0Uu7vovy/gja7lScyl+s1Bz9qXErGrjAAaTpwFFsX9/OTWKzZ5vq/WYYRdSXqkh3f
7Exm+mSONHf8h46u29xYDSKWcjSbOfoDnawe2Z+G1WoM3weC2SeDloRWtWw8UHOl0iCv3Ulwptal
pHHTzXs8/9BObadmFDNWhiQ0KdeBPZeuoRMULIZCLtGU5S9M+4v3pz4YBhJ5YyjJnaCfgTrIzWdj
DxSf1bE8ordoff7s+Hn5XHgNoWP0Qv55LIg5cVPJ6HX1s/cLeEIO87OBFGGgn5HRXtL0d7sMXM8v
rrAD9LJ8Lkm1DBxff0jCjX2smVaq4bYiyvJ76rbK8QQJl0RtqYNZeG+A71RAphzEQI7VIZak8vdK
LNWRo4NER6ChJ/3+4yuyQ/6T1PPb48WtAf/l4BOm6H+g8TW4jhzXM1LetgwnTzQ93dn5E2iUtG3G
8WOV++3emgBtHv3pNH109d+VQK0bG0MDRGCoHqjTItj5jf3A6/Fn2yKpDnx67Kz1WcZppwiiDRt5
NWIP2CbASejGv/vHuo1uFbx/YnXgdVTBmpHR2fNGsboafNHOI3yC5JquZ2bvMAi2Nn/+hyio91n4
7roBPkpHsesWnD7N5l35vdCJI985gdc0Db+/+/LbszHU2ZIdmle9LTmuu7JHi1oHzUB1Lbh0MEWF
nkLKnb8/GRf/TzKmCFrOO15afEzrunXDwqh2ol8w0knixpMyhjtUmymbnWl6mSxL6aiKiPixkSca
DAA+YSOJgz0XlG38tyq82ew8MvlnfkrCS+C/MJ/vhp0upxsMqGmBK2mSEbLEtIjsXgBcmHCvtdFq
BU1jDjJlXcQMdDsd2lYgWxGE1eVUaIrxwDNLggGvmKWw1Tf/ADPOlmAdwz0ANxhCkN3MLEOfpCcY
LmTZgExunRR+h7MQuRs1WKByzjz8Zk7QxYtthxfXmG9SfNDkrS4s7DvWRZenrblPnpF6vPWzJZjX
+pvM5VW0f7XGUBZ+ERppoDjOKkPzYzzx4tRuuBWF36hsEbh/GwAsNGQk9IauroS0OuqpEeTkOt7c
e4k4uMVa4Fb+zZFsN740AnjB5f3a3E8jXUU/TSWXP6FhpcxGqT85W8MzgLfzwiV1HZGAXwO2l5Wg
va7VZmN5UUAvsfpvDCdOWQ3BlOlmtw1xCaQkG3cDGNhvzYDUUverz51LKm6gR0Gq9j+TojDXsER1
2YwT5ozOYSglJNZwcpA1U39PSiJ+0WXpUBiUe15ld5aJCxj0S9WrZlibX/NOBVaqtaVvXo26JTmG
rSEcrdQBbPkIwbTDRNpJiN1shCplqKsCn7+Jv6KFQhotnBK1ym3Q0/cJIOydMDhjchDp3AVfMqd3
ackuxyh4uAWeTBuJPUeyTVnmOCDCkZQtEYkDNc9UtMoO7rudTzNnHktnFhoH0pA6D/Bj+mCLE8OP
epZbeTnVFGxCYJuib/Do8PKVFYodWjFWWmLdwr+/qPOd+ViK/FvUjMNwBUOVXH/FMC59auBbbTPm
40Pa3Dj28sokQ5r9QgxT9NmdtQCyxwnMulobTRkrsl1+tSVKUqtuANn79yP01Cj43VgIhLg94T4C
KiAJ86oJwXGydTThpr1YgSGsDLg0AaxuTuZN1zz6LvCg5We1tJKbkOO2mZYOwFEF+iBYceU6xKiG
xYHG0BDddhoMoZ8uIMIjMseerFEnq7ze871qO4lxPq46evMpCebQuZoIrvv8lx0VBTcRIxLcgO6r
Od8845SBB3U4PZMN3v6+hH2wG5dRSTXCbsyITJnM7kjxCPTs3riqB6m6KXoHeyn/CEO/4/ruorBn
2cjlKGDH5ofd32wp8vArp4/3FI5KSdH4wuyCeIxKUQBYvIxxHlqKJm78UvjVPzo4dkj7fLvy+eeP
8yOduEmJqQmHF80FRfNr67VaVqor1a6TaSBCUp/gJMNCR9K7Dmh87Kx7+NBvyqIhwoRi8gQWgpt4
d6YHULnPIzwu2mqFG1h2LUHQaw2EHa2dC2e07MFVFXM4d4fJcGkDmu2Q8YG4KtCSiDyOrRrU7Usp
epexuTj9TaOKElwh9vFYv24qI0/RC4BpSvhte2FMQNmu4uonaLO3rfTNCOB/mJF0mzEUse1M6oHX
DoKLdYu29KFjKhj9UzGm/pwoDRHB/6BM747Ns22omNUSyAkY0+TczXHg1Yg/GNgEBpno0FxmBUzE
WbRkpJoihyC3v3QtO3xvGs0TlT5d4EpgHdy+ZqbAnJwl9OXLPYNyeZy2QXxbHVwLqM0qOKXB0J1t
d4ztXv2MItGwYaRGIpi4OCHDKYPi9MjNj17f6SLafWKHZsrW7dounJWtJxs0FLBhBASTqiwtQjm9
u4irOOgW9CAMTfnH11SSGkolemoRSXO5976Yd+77KBzU31uRy39zV9LQiLs9afRajV1hO+8Hro9Q
ZidflMRiavbcrg2wxXzWJ5PGQNsPts9J+GI+ls16Zvv87v0EswS2Kd5sykyS/DGT34YEV4GCrqEG
wZoPHpaVmJqgkczZTjKoAugewnMjF9zxeFiUg54QAolDtqBJMGeO0WXKZJW5O8n7+OCo/H+lH/t4
oxWgiuT9IUjcpB6zXcNABeq6RdTDdfy8cvt0UQsfyCORfa2Sz1/dQCErP9Kju5MU3MFAKZIieQuI
TxW9+WBKjZU3Bvh3E/euWgLFyGCbc2eMzQZsB4S+xuI6GKAehzCEjrW+OpfWuLG8hbgRQTAWRAL2
Nals515Y+fA8i6T328+TiKip7dYPEW0drM4NQkNtZBvBcjIaTSUc0fZQZvMI45e7tA0nUBycVoLL
QsHlA7prQsAW1oAySQxlMXKTHOq6Hikie83y0F64hxkXITaDH1I2hzhFgfyFQnV57jOAg7axaB1g
jKHpRIirEv0lU6cJ3JMOKssJSZ7j+1hEgueazgHeLCoSJM/WwqaEPT/eyl9jLbugmpbc671H9jVp
KRcDFUFCBpby79p785G/iQXnRRP6NY4lFRY/ZNcyePL4KIAtj87p6OIztYYWniIN6gWciuUfi+8e
MFsF0uekMY9u88zWGRAgQbd8pLGWc33y7aN13/i+OkBui4ib4SwQBf5Vrt7iC4VKNC0rQxUt0cGA
+ejLSmPgehJCrvjUtVZeZBqltl2+qwsgPjisI8zRLucvAjYF1Y+GDX0eJ6IgFQef/WhjyyE/pk3g
ScClLyRxZW6itnIgj+lka4039hoRg/xTtTedLfkN1lPC5YtOAlX9sLdYOyHirXw6Yx2zFZNz6vC2
azNUcu3BsLBMUV9yu6YCMIo+IAWKmow6qblvRHUf5hfRvymRk4WYLRdzXUQCr1lGxRj8qIB7qZkX
2k26y1InqQCVPnIYe1dCaFPsZVT6TAvuVnu/0GewVGAeHGGyIPBhyVqAUBrvDxBnw9EwscBaOtjZ
A1hKGcciCJmDGxP03CIJ5AEWAdRlOC8QLKEZtkMlwkkIGjmCRFso6mR3O6SZpML0rJNnoxOZ71+8
v+NYPX3TlCvYjgPDK3+6vDbgI8ClIc/t9VnJX09ITqbLpYIzyiF/xdT0oU/WBe9O0yUu0PxN/3e2
sSvM6AzX55T/2ctCDWwoY9xpjvVZrbfBsx6KJ0MxH0T+OfMWeEUoGgoSOzA3/WpXYaz8UPRL1/1g
kX/a72hr1fbYErluXq2hz7kRiXq9mVX53pqiQxqIojO5vLSbNlkuc265xBLV14rR1tblVGtJLBdF
Trx5eeWacaZcdlxNlMfeVJkLuTStzkDDHnV/0ygQtUqXlEj8Ckqa97niVzBK/zCD7LpAPoqkYH1v
mjLCImz/Lxuy4LPQaK9nWEY4RoxBSxhpH3TMdCtRHUREtaVSTVOo4SYyu27PXuXHCW0HKIubjQWe
RWL4goo0veFyLlJHOpe1udKfOTWdKyr5zF+dZ/FkIlqxELNfhhN/7g7Y7HJXSjb+7sQmTmvqWRki
ZaN+1leNoYamnLR9f8thpMqMr2NSfKtSclhvAgJxhxHcv4wHsHYRhTovqI65ZhaBMLivYBg+mP6R
qanto6VolndfiVPjjWiWjhKLGV7CPhBpGwxqHlF5OwAQNTT/c0NsljLiNorYVGSRhYgiQGQDfn3B
0XRRI4TO9rIe0Bmg5Sl/QFj4H4w4Zee4QOd4A4VZGLK0Vtx1k1uVdbY1miiy5fu9ngZS/191uGbf
XE5tokLaBw32RviY0vLJnLIu/rkXjI1c/u11bGy9Aj4XGgfPwiroq94eRpixQf8+Ur4KpWkbfKv2
97owXYoLdiuBNxJ1vnmLifaPG3K5KGRIdKWJY5HPlkBtctyzcJQOhOQngE5segKQ+qpj1ectMLNr
RPH6NLmbTkLj999o2MtHkryYllKALHoi0/oTsufGMjXouFUTO8FG6+i7ta2SwXObAcsgTuuPsyit
nsHaaQDEJiInJqmjLAKzo6keb+64tZpWhQHUbyP46AfRejV468oaEeIZQ1omzEwlMJoijalFKwgL
Z5pf3JDEzJ8mV9dmaKY+THs1vmhYkr6yHxD1jQsHmUwhJQUXpIsg1ZdfqOIDgkCJ0fCAFBMtPH+0
483laFDHTdUXANILgspXxrcVFlLMUompCVvfFxZWQgXvYoQAfY62uVaG/kjpVrOSp91/HFMCAtsX
KELzf9wABmcLQmSYPAOdJZoS15wqB6YBIWs7x1GuoIfSZdx4JhjCOuaBHj4XH/9kCPM+DPw10sZT
NK9+OmG6e1azo92Z3iaC1vFRVmX/x+GuupWJFiyf1u55efRd9Mg6/YWLQo/X6Nx34WeccsEyLvbR
szR35Xi0CUlyZN57FzTDceUCeUTbeFUihDkCn80psBphjl8G3xFnVkaJOv0RCqieYgwXJRjuKOoo
CVnfxcVGZ21uDuigp9sW/TGiFEiq3VE02tVMKDcOnZM46WjDfNeqziUG5mD+vbWUMCOhWQXX9PF/
pGq6JfjVQaN9CsUQbl0bnk8UlBnBcrwk4N7muRxm3ZaBsH8NnrzQwvert8mUGc7owH1rs/gYNp45
tD5MWx5VKpUOSJGE3p8Rbt27V+kFJv5jSBECNG3oCORzFdiOaI40UxJZWyTFVhUuZ7n+XZXuBCiC
wlxUPamqzLyqF2flRXu4MdXQNr+vUgIBdpolIcR8uhpko9O47wcfcc1MmiKbMnvsCFxlddzKXJ3d
OGJX6YczjUotR0HVaTRzWaa+Hpol3UhRQCNksaVfSf+KM4p7nkYJwgXZ177l6E8ZUlY35s62mUsj
opt2nYJ15h4CkBg6PTSOBhEvW1EzvG086KlQZser52+H6WWgtGAU0Nf5BPUw57D6a0o8DhCFn/QP
oIUWj5fao71xzjWZ096wAFrqhjobrjwIkaKgweVwTOIl06bPdZMV6d4zy4QCHhC9XCCBAJHwvWRc
o2pREDiXXx3mySD7hq1hU6dSmBe325bHHOC/WdzunMdoVzuNCOW6KO8efvJl0pVo34y3+cvwq+fI
WvjAeDW0LJ+CYu0mkCOjlUwv0ul1/b29bFqa9AeFs9+tPEXlfUztAixxCaqUk3bkxBPUXP8qrHd7
f1/YeMGjWt1QyMe8B9qXt4KcRuiuO9dvp/vXPul2RyZuDuqITtoTfgWPUs4qF3lROLxvjqEkwPdo
ULVAILmE5SZ/uTCpYosa8RoLDUpu0PIBaNV0MwixdcVR2LZ7INO2YFwOJpgSwwzb7tBvwV5RA0iL
szVd9JKItw9ov9SRFilJV21+ANumsHqBeXy0w5IZQ/jSsXa47BkvRokATCNc32Lf0lUZ3Ra0PFMX
B9EG2QLBTXe6k6RSkCnwqSYytNeWVJRQsDklyb5sdtdQp71KCH424s1Ojud4MctAKmInqB33IrsO
txLVdWHHw+DrFdPKCyKFrGRPCfwlbVbAQ+orAu+gcdD7FHkTAl4Kk51BaU7d/lRYVX35oyb7dTHA
J9IYZMn62GyJIPnTmUYX8TlxSr1+FLz+sbS6aUwsGaNJ7ZTC9xbghWau2VTByMcrB6kjeVzfOSBm
OYppIlXHqJJzclT9wLP7I25zc7PLTl+EosPKqfKnZBB6J4PvC04nBL7pIlOxLAAvjjBB58tgeU9s
s+yW9Mo7E7ZMzgEiRGESv0P7+PZGi66iIIhpgIXpPsRl04eC1oN2YsR7Mwz8DcH8YImphhgWZX7Y
TGykUN884U0O8W99/Yu3rEszxoWDh0HfLVn/VVaIsnju//NJd3ZTgRgnTI4wuHJpP9Ix0cn0OyFy
yEhCgU8cjRmyuKaH/f0h0N/EGGh4KS4sTCfEms+NebrYan44Ak+MQAg4It/Sk/bYO1kPDOtnms9Q
BmvLCBXVcBSDQVmcjxUo5hwTzkh288z+Xa1Lx+jTlzd6+d7vmPX56Tk9BXNu9gs0hNT30PPvJ22T
Xfz2r6cb/ry55bKYT31c6Nrj1xiPEtbAkSiiKOKdYD9rlhXA5oo3aCZHZSyK5eaZBjzeFR6Pl1o4
eY5uroU1Z9LjNoMGUsxhAm7Rxarsre0Gml1qUDUaY9B4Or546YrKHAKMZECrZnC9DDySPwwvjjlh
JCjAyxA8/mLXnJEJXt+1jmK+T/6POuGqDzOBPU00XNZf3JY+agnmp3AAu+gI6fEHQmRM4nZZBmTt
CjhiUyVUYG0CAzd0hntm32L3xAuX0kbqXLJUhco3Q41y2jvUrNvoTawulOVZ5wC2E6AC36eX2bJZ
HYCyiA9TIvow89af182cU1xLU65IhgWlyaKHIYFyMPG5mIAU/GCq/rHudy+cte4keypr/D2ZxCkr
Xv41MqfcOAY93j5PWujXBjmV8pN4kQ3mnN8aZbiudod2HKUyK7mUNSo5OwjekCWAIX282hOCC8Az
kbZiqeJUOR6Z5uf25Y7EvwXO4m5i0rnMy+Lnw7OQd3KT0TteVqfFNnggiFjUszJaqNnXYQFiKBqi
IoJkQFFBmxBOjSGUVlC9Pn8Y8iDD6j74BdyHJxiFMmUb+vMbY7HuEYOMHFqSPCKrz2NqE1jPBDwU
Btg7Z0Ys6VLuXYS8p0i8Pg7ncHFmszLWgrE3aUKGO+XUrmEgH9/wG2VWIivVDEwb7CRwczgr7kkx
O0B2x+1/TQM8UY0ljuqGoROvkJ7ebnNFS4exG8VJY3MrNCD0b+TIrz4bjgTwTJkE8JnX1tDxFMGn
aCUwJpkOcFmUqq6mJMlKslQ8ouPI6GlK647FHk7NRR/+EsR/y+3LPySkOw20tz978F2ERPOL1nWn
EjqA9JjMI6ZSpWzNfVyQd9xr1k90UDBg+A4Kf2VXhwJpAkxnIYT6NlX3fdWODW5hogEKdzgXQiQR
1h3sdDMWukB7w3iBIZbFkBmIWwCh/TWDeD6/O+lWXGGfqnB0AIWzyaA9o2k9CMiSn0iW2zSLEjqx
qJnLJcUNPHoFpjRfeY3AXTaRBRtGeJOigyExdrOl44uooJlDN1mG8YE3gsFu5XMj62/o3NT0Zgee
mxMDwMg0IO/c9KCbNUFsPYmsxoy+AIVtCf5gAw4fEe06kwLE9l0A6PeZHU9f0M6Ky5sdW+QPQgTj
XsBgqJzlDzYK/Z2nHrGO49U7Ki1IGsQViL8DNe65rI6sgEfF9/iBbsicg/SbWcpMzuY7UwdNVyXN
ofFDXnrn7NSso0zxSGY0x0jXga08Ip99n0WWuJOTh+kAVNzRUld7ZyiBrYWVJ29c8LLa7grBbPPw
cx1FRAXme04cEF53yf4YSoO/U0cRm8lf4Pacs4Q+ag3A6KfDh9LQdyGO8aO9qxQoeNUmAkjojcBJ
mwuNs6nSHlhlMCgR3URio6LgtkXhx2pIX7GfxMMVkjW0QvgQS7roAN0ll2tVxgh1rDh6TXWntB9A
ocSjL78M+N0KDvJBKDxBVSglJmUhpoyteFxH7kP+518TRsmGvbgpuIZZ0JlGxw5s2dOn0tYF2bmi
ATmewKdYlc+dUBNCloEQ63yYIrDS5TwT2Cs9hf/7IDhxeHCLU9wagwKOfWdKfByASkN1hMXklKDE
6o0dCtlv8LNMMtDmbwRzsroY7YFQMH2hFa136qWZ/BuqOcIUgHbzMqk2jMYwdGKdE0f1b2CTepJp
vQ6H+oAhsn4oQ58ZfW2oueklFC1z+GZI0Hxy6wsj1apsbEYDUwFGzVKkJXdByrIZzD+L/iyEL46k
RlqwF//4r/XBMvFp6mjDg3PBuP436wm3wQkfWTWLGk8YHS5UQlCALR52EqWBc/XKFDF1R8BcLRkN
E1TqNqX1pdyBTkgGEoOuSxjkXBatiZQQyr9KnzpJ5tAsvJVtAJTQdOdBgJlnpgs/CZe2vCAr38JJ
3E8AUMvb/fCVew+cFgkqSgoooOiIzJ//m6mVSH0m5vwMuEuKiAQ9Dqh3LUNR+lRzfeHYKV+N5y65
M1mTV5LdiTIbm9Snv7I7EgucuHi7LXXnkGAxFfMwIqURlnHwOii07CtcQnvNSKhRBEZXEt7laAXV
a3UiQ5J7r+PisRmFtEeg/Bh5DUVY3AOgWQ8zub+1HKdTOSPZweu6dKp8FLm6u5SfpcAL63AnoqX6
k/bRZ2UfQAkgNwbSsW5cC0CIMY8RaappEQO2+M0Gx0gum1itPODgAMSPrsMKI0KrqGQJOoaRX/cU
lNLgelBrPXFqrE/UxA8OzHtvMmNpoaf2uPCaM+4RlWezTy1U4t1p2YTnElEhlCzi9aBEpm28PrbR
OCPXpU7oa3clZ9ZyZcbxyg+Mlr0Ewq8hMbaZUKaVcl15Wm4wHZwDOCWgqaBB5qwFd6fiYXfUvfSS
J6tDHrjX/Nr3xLWsFilKec9GLDREoLZcoJjlbCxkM3HffPlGQ4dW73oz0sJzU4jcHlimsMyn5HhE
Mm4K6tb19aq05KQVn9n+ZoyrGAFKI27eWgob/uF53P4KYm2riqBsotRn3WlpSgwUtdxCGx8rcMds
bfrW01awQ3mrb+6tpfCppZb9/MQaIE05/x4Tl3Lp85ARYTMlWtvU+6g800GILo6Yu/By/1FN5lVs
RhBlYPsiExa0x3OFMY2sMyvjMxvB/lBqavc/Wiuq8KtTYJZI8ibOadf2hFIQPBABJ17aFo3e4+fq
OF7VefYLuocWSV8RBwKl4YodUuMImobcoZDiUGrY6B7xmD/6kuWqH0/6tAW1va1/fNSn3jai4h2l
SmSubkppcRvEwFnoHjazDTHrhAkho52DQGUHbZdqkvwARokh/gN8hlc7/TwMpiFLcbwQ0p/y57AA
B/GyCz2SAzLklkVY/upu7fZF+VheHjjjWwNTdTAri8BkRmmmRhpyH7CTJ5LohtQkSf8eE8L3alWF
Z8xisVFYEYcMf/RusVyx08hq3fxdWW69KCTvYQecTDonxnKyeUdlYtdhlfrp9SQ5NL22psyBkNq2
jhn6OPDKJM/rC8A3gL0AG2C2ZG/2L+kEgeFHYHDvJcS5VcKZhxPpCRF8z55IfnoTtBtK4xrx42rl
K7KbFu8T/08ivKJ57PjzPXm64A0Z3kRR/LUTNq2lk6WhqO5rBo+XHZZs0XLu6xbxqgFWH++WH/L5
AwTTk9YQGxOZu/3o0LebbUmuVsIh0Xcg7g2tlzSG+gtahI4VmH2ZYLlm+pEQsnP2e3otnaxDZACW
zbGBJNkqZ9sBiiVdkSWdma5dF/q9QVQlq/WzmmzIKkzXnpKEoh1+Fw5grsJwW9WwTUkh9LmrIHza
mqoXQvJIO3YC+B/hAH8zrhZZ183pv5GhxsvT3Xw/lkPexc4uTigKsJyWbDJpCcPTYlXQY4WtRKlv
5cfmoDYUloFcZu9CyguJeH0xL6oGa0kvdAASQBED2QdsPrD00QN2micxQtpUVtA+9sYJ3Hwrsou1
5A+qoXJEjPBB8HDa/9kWNcj7GigKw9XDjP9Zti89v63TWhxreOXjoK0asdffD8bH2yLhtvwOp1E4
mW4wuzMalJmzCEI2buWixjEOCsVF8dEOYSnGTtZqFB6cER5Azyd+rjZqe11asuAWvGrQjdxNYfH5
02GlJe8osIJXrQdyDJ5rDaYH/yFfC1sLltIcflb2yNnYdMQ4tNcEBSXEit686sZqYq9lGyyZT7g4
a9JJDZrLa6hWF78PZpq/yhPiTtpxNcWAFTMrltcXHFjt5I+lq/dK95+qPWAdK38d1O9BsHE0VK2t
I067/+wuBaarQCabm2CtnNzlWqT3o5BPF4dOyJTxp5BsW3TndI6Yt8/N94W0Nur2w46OTuIM6Hl2
0iLIr3Jg42LnGqEcepjDMOCA8HDs820iadba/S7RVsJoSr4kLCfQG04jFCD5pkHxPp2AP4Kmois9
HzSg899xQ1zC1Nvc6hfMiUgYb8aV54Vc8CkSyLyey174vzjhzzEUZTI80pQRtFHtlykfv8AEmXP6
uUFVtwovAzfL8zs0Fev+ZVNCi+njBEGFM0nN0VscVkH9jZaNH9pqDzqLDc2YHX7NWvZLxOWGvtcK
pYnnTD4MdzzvU1ZxYKhtKl8Xk/XxTziP/DZr80dtQr00pqbHE0IcAX5IwAaUOjMaW5mHBmzGxKVq
6pX8hQQvT7/hVxXaME3kEnsEHD8dRpdN3uMGkDNggd0ghDxoloJMFv82eXwfwjajPp5bCTV4bO9Y
YM11ZbpOsnLQoxiB1YSV28k7v+hBnqo0WPIuqeO+Y3h6CzJbdxOQqdpY4R2ewGHLSvG4JbiTVYoV
OtNJbjqU2LcA0GEXW5fS5FRXMak73LKem0QkX6ZFCwNkhf1R8o2SRImvejTmDijjXS6hXFCJOZIG
Xvj4T6IbWhFYBdO7Uw8q6nygdDPMVCgKWRhqD8FFU4x4+s0vJmuwtzgXdOG4uGsfPndixUf/zKzf
p8qZHQntFqgTd9uE5gTLQJ0lS9dnscWNnoPJ9dZqCASu66D1ecE+ZTIeCsYfWSIfWe8iePLFMEm1
0Ec4+hMq1odvuHXXseLIPHsKQs6uDZy2qRprSmkXx68yJrkM0B3PIKEmCiAaMwPPB+r0vDTy3szB
d1uIVyo8W2BoZmo2I/L7qo23Na4v3JCpuuxyx9I2KoR6RNNcH13WZs8QoyPBLhFIHysACw7QWMgw
07lM1xZzqFubRthlzWyOtie6Rvz47ryZfIj2Itg7qeyczPMJBY2Hh2vdpulgyqLwk5C1I/tIQa0b
EfSk4Z7CVgnL+U7TIBDR4TSCD4bb89J8KA72wn2hhTMa+/ku6qcQF+0GcY+tDG2sMgxO7O+f1SHu
KK9oCD4EFa+upmIB1ewWAlu+RRX0xFtIIleFtv5APBaIvSXvkm4SS9Edv9fRw6dnr0Iut4VhPkKe
xio+3/FaNKgEfK6u3da8DYLz0AF77e6UwW3JuWw7TKEpqG0+lErivsOK32cUSMnL6tlkXHlh8Pvs
eTrf11PRaFamCHP3QDMWuyimcYHi5GcSJ4ecn6O43oRGaRvyrUZIzsHQT+X70mT2g4Nx5EmwzAm7
VbaUo+B1ljypkahcDM061dLEpiWsLt9sH3Di25SHQ6MqDVGYTOWD0buJASY2FnbOHuPZX1akkZ/S
Xbc5QHe84lcqlYfuTy5ZKFd44ttBvu0bgq/Ub364HxSv7PiE3dIY3oDqlfQDrveZeBlOQCXyQGM5
MaWETjcJAhckkH0bw9o2SQ6RmAGqa5M9SjORllOnBrgxVmvbhFgyAgPwaOhpVFCJm2l2YN4mmlW0
Tt+r2d96uW8JbM7YsPhs9Yf8y6NxZiBzegKKJ/pH1BYtVRw8oxlBtMHR6rgcC/RNU30/KMpGKFMV
piaRR2mpxZucEFHprhGZQL9qOEKPx1MfHIsFPiByyJxWugWrjb2629/3z1Onxoa3B5huCk4Uy/5L
45W43Lk/xO+rj1eAYuJInMpwvCN7rKOpFmOlJoDw7jjOLglL/jMZdkhPM3XnMCryZwxeCK+Ozor6
5jFrfp1RdwxyLVnQY62gvjFG2GwOYjOVvbj31Y3hTJNTIa8mKzvSQnNar/K+9PHfPilPkBj/y9to
14w0A3a4a9mJf3uiNTe+X5aEcR3g1TajKGGVC34OnPLixQ2YV/PFi9ZwIASaP4IHwSkHE1r35lkj
4pHaytYuTVpyz9v5V5QNaAf3nJh8CJtkT82rK9Sniht5jkYZ50xzIoqPFpmKIdIxub+Xigp9dAjo
l+0mR0fL61R9h6Bicuf+xnzVB0fzmD9+kCSx4SEOYLk5OJBZ2HazeOc4ELtjdaozICQirrYUxuzw
BdV4xMEicpRbqryPZHHlTwBk4Ki2LMul8/yLXAIkrozod/SYd5+3ZjUY0LTZO7abzN8NbgM8vwdj
lt4rrf9tVIJavcR6ebRz+tqTgsyH3j8nu3ZOlx7e8cdLXiSYDWJwgkfxCpcJRMseRyr/HigqwfVo
xUv8j7ff/gTVIV/GGg6Rwni8AVY6iAX1R0+5xBHXg13zdp2Y4ksSbJ0OEU9Fv0F2pfL8qiaZVP32
dKVXg3cIPwBfWBmkYbkAO54Un4FWhGiSIL5IV8T9VtwcdBNdQ7U5JJCU6jFabxjoYFRkl/iQDpqD
PyaegAlkxhr3EhI4eo/3bgM1ZwFIxBw+mZltKFYZYvuos4ln3SOekjYae3hkKHFpvAy9CWzGPSlJ
fG6nDYIWcTaO3aAA+wGKAOUQP/jDPubzoIBxvBlMdZs+V+fzBAQmBChOkhU4gP6cOjLkPJVj27xX
+t1w4cy+DTRk4jVC2FrRcTRIRuOcPHdDmwDjM/GftwuktToHnYlKrvvNEx+s19/Hy0w9z9fU/FLa
tyHtvDKN/G4KX7n1EnXHiE51cU5vtTHEMkKXJPhDogF3TGy3xlHM1oeRZMzhOPQTtyILkXdW/lyh
0Z41sZH+DBJLAp7NaD1fXQ3VViUGOLxYvQu2uIfUWIGeAW7loGtulG7X1IWDdq/bBm/ba7rxiTVR
eRe1B/HGxGKvrDQ3MMmHehUY3vqx+V8JuJeQuKP1AfcttYf78mdI1p1meA4D/1fGFhdHhay1Hdb2
s9Mm55HJUbnqSRvJGN6hwNIvTYEiA1/2FpY540nneG0UmPDG4QpykIOl+S0K4ksZAdm55CiM6AYt
5/MJ50uNb0HNRGPYVsLCTpAFNRnB4I7mnMTpV5pfo4wEtfjrL6+bjCzsonWjKZh9rWKZps2MUUxb
rhSG+mN9MWOyKdK56Zvl2HIgKRo6vdFcm66ZNCMMp60oISb0ik7DvtkCEnQoEnS6t9QXgD3u/79N
YqHp4KFT4JrA1mGGTFUFqdAJ3uFiKMxWQbOkyK5J5gl/ZYRVZa9e6492c0d56gtGohByWyM1GGjd
xbfTspEU+ugzFZuvQ+sD5Pp9GvnUZpOsFDZU/PuIpCt+UyPLd327lIcQPbvEGLbTTEQByq8F5xGN
yHQHKI+RZJ62CJpn8WvQifI9aBIfTNe7/uGzpJ81lERg4WbKmx3IvXjDxGF4fGStrVo1btzsuD8I
QUAU4AdH+FoIe2mdQTVQYrnpsNZ4G/5jxZpMheErxFvSKKFPePnp9L+/hbmyPAa7EjjMqB6L8YUI
Q9JXkdrEn0ZaZ7rZIYet2pVQY/NkOV25mRalIz+6IiqlcsDiK+lNXH6IE8DarU7GDB5b3OVdRLlp
bWTmTtTBXMwTaIY9d+K5Ff4pMOi8/CKyw1a+C6NZiAL0+cYwvUlVmFz8AN53bpJO2F9sdzfyUEnA
I6eZPTzBBedkWDoFC1mGRPT/XRZeFiMmeGlF/ABAkV7lkYM/kpOizv5DX/hU1vj0yJLjzKmeInY8
YTxBSSE1h0uLUnNZRGB6RZxiBQh75kYKqZQZXqAkg6TSh2XO4J6ZRjKKpzkThdtkEnVbpRIm0NTF
tm/l5z+VRFQ70/+XeosQyediCOsO7zunJmzi9z1kNcsxliIW7GO7VZJDGmHCoNPEYY4YZAOKUE+m
yZWwBnvTm85CwDrnQWgtHwx3Xn2jSZUzpW7t5/QqgDyKSRcp5Sa1i4z3oh30+r+t3LzkLFj8bwRf
EMnA+di/PVyulUr3ouMSgoOXkcRrsAm0QCxeuXDkDDuzO/kCMN1K/waH96ziryIfEiqUQJvVBKc6
ZWpLPPQvGviun6NxG3U/V2TXZC+yAr9Ft1+OAjHFK8eqURLHWzuKAzDn6OjY7AaLHpNZkAd//HqA
TarjcjdAI4W/YdcyjxnR451Q5kCvhjutwtMl4weznfZgmE7HDsw87M3JIQLFGJfglma/pbJVMK8h
qrAugsyCcEouppXBQOxP5bUMxqhms/ArQN8v6RnJDetpXlmIdZdWgjTYryNWxg2HDuhBwJ+9jNWz
q+VJ76hBCGYrISQVzgm7KnKxwGZ0bC08AhKKAvjxFwpQzKmQjYtdFHpyVjaW2wAIQn/hHem7RS+F
FZCsdUVs7Hv+ivsxzmO7uo2QNFi6vah//YBQima6TI1PaQBgbo0dfEuDHKsrkq4P0azPEtFFCoke
zXYJQkIWWwIG//Ibd9EBorL/P5i8TCNNnbFHRcSusNaPuNPBwlLAm+zK6LldwJ2bNb0VUGHMxE4/
FiTzvgNLuB4bA/DjsH9MnZnCnKMbBnIOaSn/hz3TZv4ya7FEU6in0cUKtgOoNXkbRjfH0UotURlL
1WZI/qZhMKhF2rNWJkWulDydWvj40/sd0sJnfTsLhCQRPTj/s2YIUUh1tWQ0Bz7zs1P9LriY++jw
FL/PEvmgQzIHmhp0XdmNrwsoEmsObzxcARD9Xyu6nY2nzULrmqvSjEMbcuLSNRy2XLjd5xx+Al0n
IvSchlaNTByJcdc1X+zyqaZgMoqtX3hEMt7zGn9bCa21KxXzzrNZ7/AxDVx2urvPQCb6KNLqvoU/
PGAmyQydkaqtAy4R2yIYiNm8i9RPll4L5LIbUW1ucnRcEIIsJBdboZzUPKRD7sP7IxLlMwSJyyrc
Z2lUhZ6dWxA19cXPoggKHx0Ecsm4sK9ozFlRVmNGUNwTDh0y+1PGpi000VkwCfUwFNJ5A9/kaut6
nQxXsBwSx4gNVo7KUYI6xYdEIEovkknBstj9cWv33jYp5Cprbp+UiPl5NfH1Mx29YsEjPF8OJ2JY
aNfpJGhBcwPeRseM7DbtZkA1R97M3zCsmphQvKzfWZSVrC6zLfEWV570ZfzdbA4H30AcMjjdr+LK
55N0j00Z+RVtHFmbBlDdP//buQLcQXdLmjYGiFrEByPYL+H7DI3i7DFyAJYa2SoIDVYAaaUJUKLY
K42fCbrMiHn2zRCW6RRjcaV4IYehJuS9woDYqIL+3KHq1+QVEQw0eTKD8nQsjyE9XS77VwPRKytB
9HSBBxnB++Dw7hAbxrlx2gb0w4FfJ4wiw/01G4eYTuz4YnPcsdFngl16fS2mIOM5vXIBerXPBdsF
Lz3/Ab+3WHPAwpmAL/RkAIVgrrAH/+Wzvln8XY+TSOaIwI71CI++b8Ma4VZSt9zTiN92gwqiB1Tp
TKsCXY3whmPwRqOQz3c4KZmiHHZciXZy+OgLRq0y3LFSZ1CeAzoTmqY3RA6Q4X6OaJkuTCJIDY/V
X73nrnjZPauydTe5qy5qr4WS6j620EgS9GJH2XqlTVsZnvgKd34gJMQRrGKsOH7tOvaozJyxDRh3
Zkj+wmr+UdsMNQ10z4KPZiYcfhbm+rrBeQqgtXNtjoU+ori6nawrd3UZpVasCI9aY/VIW3Tb6Krx
5H3409fbNsUuiS3ulS3KBOJw7LTjUzfl5HRu+kR8rdfzRCVkv0x/K9UkBpQIu76ROCK2nK79ePuO
Ar7xVvKo030mTh4gg1vTR+Kj4f+a/afZAX1wc6pNHvosezoQseilpYDHnhiPVQ4+ZQaLeJmKw84q
2I4DyFSs54AUP5xd9P5+8tJWW/pLRm9tIR7Hh6jXJgI8xaMWl+FI7qlmdU8iHEgHKET8Bc8yph8n
dF2pMbePuZabvBFjRBclnxuehCNY0PWxhFYygBbv2T6Cgy9C3qbE+CWP5Dfe6uyzbYzH+y6Gdori
N5mGOSUgjqSPLOyE7C/t38l6Defyp5h7LdwEJyD3INV/Hndz3dWmLYHD0Z76TOFTt35EQMpt8VSX
I4IRbhjutp19EkppxtljqKBn7Kx/9VBbj9KSGwq1oby5OKWPZUhg9UIwcSV/XkUVXKyFC0o+f9X/
4+CwJVuGyaUg/S87h8dr7FYTAnWVFLS79j1lcPAY+xODOh03KVz9p2AAzICdLyZXAU8i2VbMr42z
4a03JH44oaCitc/jFETHFZXvcm38U+rZl66bcFcPbSMvPtgvhBaVTjUTMysqpkoNjlBwTBX1erK8
zI5T7I+cnl/3ffwS6uG6TfmnghfQt/pwXpe12AElk+/mnDelEJa0+bd06vPEhbsazyrsLvn/VUqc
wZJhSEoKr0kvweoWAzookrhnnNqY+ARcvEdA9+L602r8/TxSbLDLP0tJlhPTfoEqktiT1f56noqJ
MRapvx8+9exZYDV3HaIy+QqDEvzVppRmMaNvMtPWESJiI74ApVwDHaQQhtKjt1v2UpuQynXObub3
pIBtimMrYBdtsnJCxh0Ihax014bD2uzd/3TpIUQXU5MSYjw22XYnZbsbY4SLp7xemRkLsCqpFR+H
5tAKfdlLvF8++zIh6sy5elJlq9jf6ft+tWzutCz4nEtSroPsHW34ssuCUPuVeHZtiioeTXWE1v6O
QxLXX3uvYiKSJISyBNm9WV5gCiGMCZ33GfSoTVKZGYkTiZtXyI6LPMni5yKipynAAWsIAQyALC3y
8MA8CnfE7J6Bkl3i7/zNwNYPKjCvojmp6OP85ojwYccY0RxeHgFrrd7PW4O9P/YZ7lWBdBptCBAR
wKtzhllMhTbOKxq18wtKbokLNmNA1MTGsd2cF+XSIVIdkS/WtOBd/ZYuRilYINm8WaBJIO3JVZjN
G1Z7dLmmdXe91fLlnEM3u/vQ/BvsNXrC8Of/8yR6x25JKFhg54Cf2QEfhTf17IafGZET7o783yLM
m5Q8kxwOPDgbd4uXcrdAvnXMvfBnkDCju7adgpZHheipTo+B24mhMpkaIzD1epNKTBJ4wv+1M4DW
bkkbN9q85sMEeaWF4g/umIkDpV2Gdbb9G5Vgcf3d6XD+g0hLGpFKti/Lvh4u2Nx08DrYwwNsqcp6
JAx2vnfM1+fdYIw6dta6OeXDdUreLATS5xR4u1resKnhUwVsI7DvX8R1Y7k8faTnM+giabfvc4jG
+gaJ6VED4a5NgAgwoAdMO3Nq1SILe/62VD5LzqKsgmX0TgRvgzVLh3cOR4jkL1C8Ns552YQLhmG6
Gd530ay/Js4izSgYmVyXzeWuGrTFoSaAmIw6Ep5tApERjyxGasVMuELyNEU9D5ngKlsgkDU7yY/n
rYGXtVUs3SZ6vwnEb5TkIGvaOejqICV3ht3nh3F1HKcCvBz2HLSmx3e3nwKi9VuxXwXSgJO+ZRnH
3DrAjGlj/GLH/Wg9/8oM6CYk+kBuE72g5k6XEfN5wZzaGvRR/k2g0dzq0N9ftNfcoPTC/uk7B5Wq
Iyd5rReFSVp1BgZKHxyeCQY5qOG2HQg56W5oxT4JOVhNm/SiZ6nmSMVGGjuZrB2wS6FpS91f8IQ1
ntdveyxwcqj6yAl7k1HIKj7GHT4ps7t/fxMZdnCT4msZhaDwzHbH6gQt6E/EP/C+MrPGCB7DSvIm
BxZaE+5qvAm6gjZ6Fr6gptMStp1ZfvXcHOmvHACkvFLyt8pOb8Z55rl7YFS4JXEp1e/CCulvCl4I
ZGC21nmJRCNdSbr1KWxQ7QNyV4SywVwMQhgdxS6jt+oEih7U1ScMfZYOGzixEwAxao9zpc4atnZ9
cGbvTDYJn1hXJXHJ23MQ8PCXcaFvGrwH4nXUWGsA6eIiUxtWtH+B3EuONsBk7RQlCHbsrxtiRx+w
25dWPPpVdoP0MsxTlvYOJUIOIcS4uuAKvP1vGKtv9vaTn5VoYSbZyBdJaLVJDL7ULsxtWQ6HgJwK
/+OJPYEiGtmez0HW1Ik7aOFUOVNemjn9NQJNSNAj4mpH1RwlHX0gp+M0TlFntDEBm5NcFGFwZLtZ
7iLM8jo0v/q8pefxNArzyt20znlysleY30iKJjVZLF2EV7Hytb/zEPyLOEGyZ2zeCpSqZw4fXGZu
gwXJmiSLoOjx+2pIybXbZnpIWK0nrbmb+tH5sjted6bNlimlj6IaqWKwTHjserFL2uRN5h2xgmoN
JmaKCApdeO+PNbY7B6gapwLSV0sTlMswkhWAd2vnkQ0LvDD69ekLv56De0eG6sSJOL5Wqc92rrtA
FBVJpByOhX660cOy8+KLkADmf0HfT9Es4Vf5NcfE/DfgLCP7ml0bQKPvmh7QuQnWjf6edW+qdEdf
HRhOIC/gVZimCObX7JEKiA6PezdyqItSIjEQdiVwD5G/h7iE9u/Tow73Vqcs2hjcqtppb/TR8Q7V
gAJpwy6JBxf94edZLUoi7pIXumAiNU/i466BRluRpziA5ricKdI0Y+XPl6K/nk6MSUPqpzEhgO7p
YXL66TJE2lk2cYcx7WfovQN7Oml4knwfIIn8FJtw5XWb5nhfeXTzSwHn9rpTZ7J+0s6bv2PXifby
IuHqTs8WW6eXHSAj6W8HqNl438Fge3LYH5dhV0V5mABxX3dKqubSP53bn8B1Zu7+lBalnG9CXZy4
BCbDKpxqvT5wQXMPDD0TnOezGxCat6Xl3F7gaJvYBYwlG4TmSrW4P9GtnPcH5NcWl7owXTU+xIgR
GVKwLbNsxc/jEVR47OZTOBhX86T3Y+dxAHjggrksnyfK9oiC3wu3ERotex+F2t6ODPacWGZMltgk
KPlk7qkau61gD5bEBNVNVeYB0wz2TYuflzTFr8GrpF2txIhglQkqyGQtL0nzYJEWg9A5nWVIYwBY
lpzGmO1fPH2O7J7rxQ4ko0M2uHVzK8ze/Eg6uoZ9jyVRwX+zCwgqSJf0+dSRjC/J9SPTRNpsMSad
uiAy99pLiFUvxhvLSlpjTHOzRYHBz6QRIHwizIWizMO3jPzc/MJIPmCpXDT4YpHXDjOrshhpfSAO
VhWTDOvBn4cNtRIXgvy0lm4jyQzy8yvx+ckNfSh9HpE70keW+iLG9ZOlPZuSWzlND4lsBA7gKxhY
LHc4BCOQnmj4zO6QcStyLOLqkhCygGEcuBwna2MWIZkBGRk91cAm8SM+acXEmeUdNgNCEd/I/Z8g
xzTt1Wrsu9GxFkKrrA5YVH8amC6xUGf8F4tgmtwH8YL96DNDNeWFFpJM8gObuPk9DIyeVIiXH8TH
PgzOns/wO7eZkpVgSHJ1v7NwZRrMbFGVmBVr6bnzD3l7iVktBtLjokACeynf/KNjMCfVYanEHE/9
e0/QeZKr+xSDlKgSavQwOjJ9ZvbqpkzOpJ/Gs9bRMVQ/X3jweVWaxIZUgH0uP2VIgOC0YY8w40m0
IQa0fzVDMb9kaWNPf0OvEXVILxNKdxiMuZyHgpcIYXxWid1r2Ei3Mi5nQzgoZOzmAkHKSRIV7kH5
Hefr5lqsdMf56v9D9cPhPN0Buz2j65KfbO5uYqHVU+jZgUDr2fDIaIT04FWCASrapTb6bMJ+OOld
wDxbvuTV9+rgwbLFbWWtj9oRpKFH+sAP2qVI9qkzIdogP5h0RnERZ32m0+AOyGN4gdlyDchWHL/t
ZVCPR/egl9aRMbjdiBuFITNLme4XM0kZtS9V8Y3u41RH8YWHyVnH4f/c3pGx6WPpQXMeg1QbBKyq
doohj7EmgfinU6DwoZ9s85Jyz9WIttkFmibCVRhvDxnu9Jk7gHP1t9HHuTGKmMNfA7nkvn6FAy88
c5e8I77Vn+BgZ9gZkDO3XjLuvms1+0hdrxAMAcloKYsM4NYGjUP3/MyWM3R8ddOlLrev/66DfUI+
wSM2pu/McdwQtoIaucu2n8LE86RxX8evT86KPxknbPdyQlClpna+AJB1Oofcm1oIIaRWc3icg8qB
UKRO6t/JhES327idibMoHRvX9toW4BGOu0ZX1dadskSAcHK7qxXx1gLw0aN4PMJBLhxUWJ9QK6AP
kpzLpAOc3TUqf4aMOFo+zj8LBPruvlf2asIP5Ut3B5N4G29dwA3vrBHSUzsPPPuxTI2UcHH0UzBh
oRSz2p481fIXwJbs8ExlEjpLBx/TAtjcubunxKjJffXJQpB7KX/SaSPeowCYjuy2ZC3OimdffHET
kkobMoLRBP07LUXx9YTLNGAK/DTGlciSwKTkWh0r1HQOKERkw5PQXigtPuw0a0YjU9Bz9+bM7CSm
yUpt5f6o9SBVnsRJL8kEtpsYte72gFqu5Prb//Wy23KPNLLZeSEj29VwaqbhT/4bCTNFKLRjYyDV
wJ1TdVQX2dPRt8de9ZCOAeoDtmUUxnG8OBEzD7dVEPKBDh8EEI0yJb6toniMlUg8kRJaR5J6QRPw
POg6EEJmG/Vczz6eFRj9iW+7BvYMbDiniZ/uF2b1eschVv8t/G/qrOpkWUzLe9TXTzWEfx9mOA/C
tKXiIhcn3FIhcr6tcamWhT6KVrP8PncAwi1E2GfAMy3AN7vkcamFWmrpmmvgQzMTG8Wzf/aqYdkf
ALgx4YYyUxrt9TYqwmzN2SR+bwVBQj+fbsqNfpIKp5nadUxUD/WaJmf/fqk4U5BPGllNSGSijCGN
mmZ5yj4C33dUV/hJZw0LEmhETdmL2gQXWI6BKZ8sutD4Ldy4/vf1Y3yZGwVlx6s+IQSFT+STccHD
kXuDIUrYWxeyGwrP3Rbgh904cj8LGlDNZsK342gKCVX9TPxkDeWA/KCBewKVox/LswHk75Qy9wcl
uAWyeSU15+FtyR9sCgZYtM9CdHhikrg80iY0srOIK25W2XJ93QJomBuhreSHcKdgEtuUl8Y1XEmK
q0e7xKTrvUdiaWiK0tXqxTdYy1YvG9+ySMO+9XIbYuebNL5iaqi6Jd6ZM5xmSRle0+8vRA4wwv7i
6vXacwsNXI/SwZoJN0ji5ypbGNoT61zlKILrS+8Oykc2eCnM1pPehC9IXylEgeEfaYJNUEjLigkw
ofYqPtG705mieK+4w8Y/zIAF5UDzztRNYdt3y6bZgzT1iDBIhMbizmhzQlCurGcYRCcNjEzEDaM1
m19p2dcnZ0ISupT3ASGjB1Kwb48e/wng0NDjqVLIokREpeHr8afVm/UsuK8ySRtYCx4i7tZEPvJA
NIDFoO2abkJVZ8SwR+WpwmDPmActh62T/1KgxcU67MqmFJJHAJYUC6LRcVEeIXaSMrr5msAaN8Lq
A53qDvdVyI/v53ENGaN/SamI39MUmFHc6cMOswE/7DnQ51Zj+IiUIb1xO7JvnF5t0nn1Egd3SJL0
RONstmc/g0GFPKtyOJf74ybqua8Ev3YmOkNNrqyrZoVKERGTseL51engygBMJJBAukBSq+B5mGLi
R74Sg1np99Ik2R2ftTaXfQQmnqGOwRGZi/dI85zz6hlQvLLr3i79nGDcnPkbsKysfoFtH0SX8Bxe
Za2cDMXjyt2ddmERvEcNvm0zgmynNNAOGgksPglCRWDGfIfLCb7S1aL3LKwcarBovb7ZZTFvOQQV
rFMlHf62mXdHp5xJQ0aRVKU2Pe2kcl1XmQuJzH0ZLq0NzwDuIZwTDLxyA5x2o2mNP9czLG+HiuTs
E5IcwtYrTnVJOvaat6M9iFqTkUZpgrPFxyDPuS3FHtvMJGAId4FuhQkEMwFI77X/vrtQkfalGkVj
r82pUqztrlhADH2ggqRCNuSbbWYHzTyvXRplUCcoxh4TsycZht7mcC+vjy69XB0uqa9741c1P9mx
lkaEJVnfeCkuBVLNt8ADfAK6r9m16yYo/cIDBZdqpzENM2l8Dau3d0e2ufZYiUFp+WTCKcjyGEVv
VA3ZBgEMjL4DZefYTrpRfCm9mGP7zuZrR8wbU2wkRFZphxrkxvZCqh/QyDGx6PTikdgeG/v+Oj0X
GAphZE8Ah3Vd0+jkJoj8sFi//jWVkaIEsluBjet7GWZeIC+AJDiZrHAxqJcpn7vXffksSsRnuxxb
sy1N6Is+rm8kW3COpWz9LKPU5WgixMS+y7YNhPq2BWOEzB122YmsWgfQB6GWVJs5njgvC9YpX83B
9glliKmydAnfI4FrvSSyFcM819E3aJ2g7w8BYybd37u4sztdx6LrRYiLv9iHjYA7muH+nd/JBhKD
Gagx05cpPq+ZQt5heig/r9pw5+kudaYT4LQSRqgNOOU+juDyACvuwDe2yYKLcVH+6xwtaFFgOxcZ
k7jl0JJvLgu08cqf+zO/YbOg1PqXaVEWzEtTG4PNC0THoqYn76azzcf28yIJGfB7zW9Vh8/+6hDZ
vh6rofptnnQiMh7rx3rQ7MdNKBy2V0wLrAn2/mgYOPZ5LZxAA+cepq2AXp0g0aEnz1oeZtFz1YAr
yg4hbDkMA/Omq8LA7UVwU5wcc0pt8ALHeG6iRBoahzgY2KL+jH6QX6c3WcSqI6E2joAvYxsePV87
HCtc+/EIzrrXWJ9X8sgfEM4NU0Km6xHl6XFGfwSpaS7GdXmPy9KS9B32ZWpgP6PYSiyvdT6reEYB
DIkHzbu92wGFRy2YD6j020H4dRoVLvUzYKezP1Wq0xraAeS/qZpvpo/axr9MsHazLHF++vThFYOK
J38pd3vTjtCOwHYtx5ltqkqsYz15Udvoq+r60ImHXCSj59HqtUTfiifMcAQ2ZQkIYuJLgwg4D4Vc
v7dNnCJhKqFyxFMJqao86Q8IUaVY0XwbWPW1z3UgTeUmpUoxBJrWAEc020RuK+LJype0ZOAUzBTu
KNs2ELkVXHldRvUIGsRrzS2aX8fkv3hETWFT0xc7G/Wz/pGBSkkSgJ80rkPhu7x3kF018tQGGHrT
73HU/i5lNapda4AKFdxBtMqIW0ORjgpafm64TmzlrpQoZxYoonDpBYPjFZN3Q6597JZ3MhgoMInA
Kcw4dxB0+T2Q9rc5H/Pg5f+BbVIqYh/ds6xWMMQdcuRDMEpf2UKfyu1lboQHJrP/sN2IWTkQM9Q9
cBzNDFccYXUUs1mSZfi9eCk7XjpjS6nol++NRq5eYWbsa/XAx8+X0CpMPvtFlepmfP21zfBu/BHE
jNVVqy+GiBrByJEIzAHistPN/oT3E2foVvsJcv8LZEw1IC6lvfxOBTblowmIDCp4962oEa5UdWll
NjZDyx5Wn3keBHL5bXaNuji4sfL/BRVC/TIpFapMP4sDI8Z/QI9hMD5rfoFeSLWKhbHJFiSeiNO+
M7AwTAXJbAwj4PnV3rerJamuCDTHBB2L+LTpLjXMZi7C1iwB5j3qwnCLF3j+JsJz444Xgff8DYaS
8xAoN49th/I0JjjOhnts2rcTfr6z79OwKcdgi4CBxPraPeINW0BHitYuaH4AXPrRlojUGELhlol4
OyRkrsln+64pTig2r2WW6XcRhLgPsXfOdKe37ZAyXnWN3eI8I0mv/ZXfzhZ7CzO4eGtrHYO6ckWg
iVQFF2VdvGWKld8Kf7rASTkGPB+WOomiNyBNUOMcCTeM3NfyUGj8wlXywB3rgx6+J1KYfzp8VEDk
zocb7izgj/dx7Ul5PAzxpy/KBzdSKoQX3sYmyjKD9iJiYEjoSkUNDMsrATKNsR/ikWYmqzb0wHy+
gRigulyNScSQKJ5lnWBjvhuY/aFKW37/0fYFuliCV4r0M91DU6HO6d5zALCmyi5S2S4Hp8WbQ0Rj
PEhKvxf+TjNlB+QX1utUOHfP4WKyiuZ//s69KM/hz/LuHSYuEQ/bIWOBxReu2GYyv4l++FMmh8aB
eED6/Q4MtohYUg7JNZ1zFTvOyZIEpscO0W9ZWBsHxkPR6vYjzhh7uzp0WQlCInyZhckl+A1oXhLa
SYUnE6EIMvxsF5CsFVxtOqjMRf9Eyz3X+atWQI147ede5bhctUwSKDVA3BVWaKNpzXnSDLnuLo2T
QBwiuIlU27sbqCDKMzlrqxKzVCmelfcGo8pdoQ//txNdHbqu5yEU4xKRurtpVSkJ6vXWR8ldg2E4
Bf02EbmOAz6ABSOUtd8fxmK9YWYZibMZnCDNtuAuIY8qNIc0Gn/34E6wSiBUm9AmKvV5QqGz1+nl
qjAWQGTsHMgYAyz48Evwjz9cTLiDKLFVU92m8EG1j+DQd6Ysv7C3WWbsLI+TQas8PVV3ZZZDj36k
KtGzV8z0AMoMIhRwdn8q54GvakjFkqyJwdVw8wT2kTHmxxia5gTvbWz0F3S1+XiYgDcowxrgXTRM
VQ+b95eybVFUMuybK9rEkWgoWvDevCR4WH2xR+J2eUWLpCFXs8kq2Ovh9t/PukW+E7xa4GoVnfK1
pUWImcDTQfuaCVWWEEwSgmL058CxMFhL/R2xrAOs46CFVNHkT0NensNysoOUCpK6FMu9mAFNO67H
ayfvt808OPM8HFAcO7Gn3dUKKyX4gMzICOQv48pKHvmWag3whCcOnBINVk0dYr/EqPl9FkC3GkIF
EFlynGe5jbmOdJj/U4Ov/e45JSkTEmrJDxlHcR62gjEmuGM8dn4UU2XNuoskPYREMVwvwPZs7pxT
SyZ3Rl/uP8AhBQwySUc0y0jSdLeDpeyvy1lVm5BbBTypHUWr/8hMLL4tkockdsjsulG6Z0115ZvY
piDtdI0NjDWkl44YSmmQcxJz7zyoJ48stPMKFUnKRZ1JrakpBvc2MCaPsLHsBhJgyBWnveZusi4m
wMLWNVN/iJMij33msC9bUreKKQqHwjj5rYh2frkt+2Pi/+spnddbddjkRHTyEoEkUcmyrvqREYeo
oDRXemsUhUzUEIWVhd/c5F8hS6Q+HeC13OuvA3vXnmCjg9jSC9LB4aE8XW+hZ55eLT6+VyPJUW28
tK1A2RuuudF0SDxagY7qTsLbhOXzM1ILQL3+3+C0/nhmEdioW+v5EWEJkkb/832HDzoYvzxYi41c
e+j+MKl2LxWHC22JovEpqUy29k6gV47uYLLg8POxpGDe4FaGUYdu2Qxi1uA2+Odd0cknXS7gjEPh
wlPgPmQdkQNbMw+0BIRlpBeyLmCt32yUnKXzLzsdYBRj/P0aE6g5H9Ze2o+73os7SMpf9cgy7DJD
SyylJYmqb6z9kdptftCGCJ7y/qHxtjo96EIvXFAzTYNCEtlak0fDuMlfKOh2Uc1Ez1umcgi1PBPO
tKm7b5krb9WKE19w2pSyJWIrefnVxBVFXk7ayVdnCgEn7CKg4p1hJAoPGcPON+mtselG5dSxdXXx
Qf+27eCPicHRS/5l5SWQAchqTAP2Cl8f4T5cU9X0WXeumxf8VyrMmWBIUA/9bOIhUP/+f0kMEbtx
bAyEEBnVsnCeIncR7yuTpIM6grS1SN0b4Y4zq7xaaS3TJNfdcUtT9vRRaD12Eh6nIjfa59ZsATdU
GjwTLZwfgioWr7Pq4Z+EK/Lkujdqxu97DO/dVb9Up9ZLavKxllQYBN0RLex5wbHSzfEvdck2mZkB
4xDhTM5Y0NK3LdMnxxvmK4MbQak896wCCpcNVmrRbtzb5qvR6PgEjCtr8Gak4Q3musDmxC84Yfgc
HuBFzab9FzMjfUZw8VPpJUoeJO49JNedYdEWC3LNjpmBxcqTX7NXjMJZYn5sgZYuXB9Qof6qrGSY
1WiB4C+qSd+ZF85C4or+Lh7Dd9Myx5x9SZkME/sR291UIMf3hm9AKj37DVHbsII9tQVoNHPYlmiM
XS900dtqVQjzkBtCETeJS/JtthhUEOriGtHhuhmz2dthjfKf0A2NZA2Ij8aeQEpguNxEuQs8YVYI
3RqLH+XWO0Hj++GIAGnqyqcNaQioDg19x1kGVc3o2pLQESkmChOzL5ky+LN+tbzsA3CxHvP0m1A7
obydLHk791ueR2fU/MMwhfer1jZkCYBlfdsQmwA+0VWmSZ/zytyV+q+Lck1ZfBsY7W0l768F77tU
DWGG4r8s5nVZMXsdIx7xAVISijjzR+Azs7vP4iPIkNLBQKlNll9orhllnKBYrRXFTsCyFjjFCqEW
Kol9eTszjvgVwxCzqceQcY26RxdQkcrpz05kB1X9pO2vcjFjJ32Zd6ai51a2Z8wQVm/IbfXM4Zq0
SQqeX0HfA+hDeDhtGIPVb8zilJqTCWXCb8BHJYEMP+ajcUNd7JunLbmXLi10rRxXwCNUJwLH1RNl
myZibD3JCFQ/RGW5svfGrG+1K6f9UF00zb168FvZbuKqtnlQ4KyPfvO8OZMdjGhJNgiHnHOu388h
qptcwO49rtAgELPyJXEYbN6NC6/t8JI0NRGc3VBpEdIOwJytD4N6QV42lwVWd4M+XSkDwp4bLusg
SL7QyVm28FE8GnVdZAI2VYedzmcdUeR/rjDmcc1cOp0jfrQWiFHzrjdWVIrfmYnzVT/9YXu1rwNG
Un2fuYsqymf9WrFfqFAu+Yhp58bTx/VLuJhq+cmj8cjsFdmcJ1HGUfsKrcq2RaqM3a0gyg5PwA2R
nTiMvwXeBv37sLSCz/we4eVt5Z/0TEzjSLJJbY5xmiVT02hX8XJZ+wFafP8IvH3LkicnhGNdft9W
hSLoy28KCGhfeeP9857G0S62NwMWcib3VGpRDW4SyvTCMBN1tN4yqVNPFE50+NHymSwYms+qsPOd
shyUUEd4cYBTK+zOXPbdlgUPN7VOUQdGxOtVbUreywOZ2Nl3QpAZK8yujCGDscsFjtOCj7MpoRQ+
21KrBJlu91mQIumsuwtFGcdJVp35HTzrVqm+9wsKSnW8EYncYi5+J741BUxdBPRDoUmEYq1vXmcG
/tOc7sRvCPSquAHzL68MixHqsG8LlUKNJSOuTwdJJohSKWQ1cEFV9IkOdITtFQxEWH82DGsuB/xc
Q1gRcUXUWU6raLCCxdyJbCFXgAR4IYsS/2/nv3hbAIt9j0PRtaf1JQfbk/Knzfk8w+GJEZsqEgqH
hOpqULF8iTx3a531A0YuRvWooBnbUmY13LxOVvNUh7cJqNtGFJIYpi6zpcSxVNZjj4rFPlRRSCIb
kHD8ZLRPak7HuanCfbZVJ88SNQxhCY5YTAxQKAMvhYpUDo7laRi5NghZ8WUyorzpZfEXIojmDhl6
IoMAhHgBd1cCKlzgYs0Klk6u/mdIjVNco5B5y3wi0mUQcYWwk/zm9Nh4IMqDGTOXo6+ZQbEaSDEk
3dy+P7Ca6RAprHFaqnu3kpge8nc2lCevtjONskGYJMsaMvgzdVk8HYurR9+rZ7VKv40Og2y6s6Cd
ZQUcD+1QhizXqIoH/3OA1ETh7y2sQMT++PbaZ7tk3yPS+FCwv3b49MVl+s1VeTgW2Nn7FEjN4QX4
Lm5Avrlv/ItEwEGprCPckrsfu3N9kQoGKeAovNHpDlQIAO3oRaU6+3mF/tpXx8H1FJ6M+qHhRfyW
hZJ0CB/A8HaBukvojIOqtBJKHwfK3OZ0c8eNeyWJeb/ae/wq7uU+GF2X6cPhEROL4NlvfuGl94ko
XR6Wstchz0kwXJoFRPgwhaE5A/rKCsmA5srK0KxhxGjOuwRTGjAQcwvdvoe1Ft/MksSitGzcww8L
Ltv+i9FXbZXPbzkIi3tah/4oAyt8vmu3MeM7v5ReiN+F7LqIOGrcTxRW6bkji3OccRD5JUrgAy5G
hAJIY+vvBqVlVxRKCgCIMv1Vs19+OpOT8iXCJLKrgqtnSB6HN+t822szfmwGRCNXwoQSL8/dL9S4
79zdPPk5EoV9xye42ZYQDHzNILxexrlBTsMOwu9FG4/JgGPtpT4EE4Xc3yWiGcUsfGB8RFopGZyD
sO/8TetbfjNzVCSEh9FE+SxZwV3gEKKWFHUs8seRvDwzJid391/g2/utDJoPD0gOpJRR/Jv769zc
I0z8J+mQllRY75/ztbp46KfCV9EMXmOAQxv5DAVyruclEREn6f8Qf7HH1tMBmYNDG2cY0Nzn99ar
58gu6J4n5LNjYlZfdVE8Q20PvfVBq10PLvj1zESiHBAjJAuBquYpXUlUs4hMc5fuwmUIPLaQGVMo
H82LgCq0eb7YaavqNxBDmFBhlSiK3DPGbeX3DOZF3TpadTqqtOfrswRhdkaLVqUNZlpB3IpXE7Sv
GSjh3l3m4CzSpI5DMKx+NA7q2tvQSr28AtPvfpBUQdnLNn/uxlsUncmIWM0VXWaTPo0FZELcX+4p
TKyYP15Kb9BDirG84+GjT8cJCTUMrAJ4k/JWdLlInXaxFlpfGWgh8L6FUoB34wWQM0J7YcNc12kB
1pq/UF0GOkdCgzYjzzQ4qDlqhvMasJVcsfrISAKEIVFy2AVa3GpxPraLa3dalPy2LedOO+Ax+4Z/
PvxlzNFRBqk3vS8MHA0J/o9jeRVYCsSoTEJDFXekgtWu/qiFUSsAqFWkny3Z5S5gk6Mxie0q8v2B
kUt8BTSJ+guincGB3lZXo/m1YmL0v3ZY7a4mGcvXU4/ZxVFN+i7IVdNJDAp7FlON9KD8Fi/fIVfm
9k0xvFKpWa+u2CxqnBhjbO0M3uD9IwLvLX2xVm387hMp122pW4gVWrPbrqWf8G2wxA2JpMoovYNa
/sHe6wE2BP1cGesZlwWNv/oUK9KZqSibvLXvDSjaJEVUzrP1qqaQ3Ht044VxDYdRVJTovjw7IjPl
7PFZPnCYxwvjFswu3fUi+DsJf6pwA5ZGAo8fE78El3OmWQXf6FDn0cjw6me8A1RoV5kvrR3fYUp6
PJRE5/5SVLmwc8ZqO060JVtXRW/uzi+/ft1aLC9p2kp6BM+Rt7cbq1cjlV6qjyfbSvl3hNSWforK
Gf5Kb4vHIg8y50WDQ/k608ttRV/g7HCF2D7d/88q5ZKO6hhM5tgou+FBc/Rfc+wNimPN1e+e016Z
eniukiZ8bT+4Uv6nQ7PvGHDoeebd6RQetAgVqqc6+CCw5uIOHD5+yD1x+U5lglEjb+HXg05MpLB6
hw1W6k8pBqoabBimPGdZ1/OPnYRy2ZS5XzG0a9uXjDg4q+obdi+fzhRqffqTI5INr9bReDOa+Evd
lhrVwBqWpjARG6f0WKhOcktuVwH7SBVrxK9Ixqkd99/EdlQA2qp1zB3mhYF05tjCA6Ge1qfTi6V0
W2MSr30PA0FYxYu5aeSbajD6EfZdxZe7nVe7CcnanS+kqAFbW9GX6/ysT8hX430yufndFnv1Lsf1
v3lSxecIzp6XBlyOi7a9g5Zqj+sD5By0ZMd2Zf+XBpXJ29vqHqRz02I3CkXaTPxB1HJCE/iscWjr
+x5VgYSKDMFtVKbpVdY8BXduT9YV4yVW9lMryAtCCIp9BY/iDQZYyBW8cf7dKtwAbvjy5R+1fou8
Y784+IBkBaYWLhIc/ShEXlr7lJ+2pv278y0LlPzhH344ACVow31EFHGDRynZSHbJ5CporZCm6cFr
KBe7hAwYVJFbyoJ64fABJlEzZy4BVc9L3y+2XfWIGT9FROo/k3pAU/Fkb8Z+45UJXVVaeTXgzOIS
etWzf4zh2Dzz6Sflal0xYo8hy4AG2/ZGQt3pj7EocIKKeTB2ZrLw1Apl8Q549JKWb5CYjapbFnsP
k/V8r2sEToF4kbd1TtI2D+9mDbi/YcUlerCfOeaDL9iKKCUCuEnufGDUDncB2i1TVmAsQmi5WeJ4
H5XlK6BzfObieArZMcfkNr85mo9GREgGypnLnVC3thT2gHpYUXc2yBHiNh0CyWSyVADRMjQqU0GK
Qt+ZNffE4YQ3AI0wr+PyribGGkmnx1E3TxZOENZkBl6rbHUU0O2JEeiTN2s9uuiJ/aUYBE+lQ7nn
4u12vonBPiNbd7+13Gsmjot2ysjH7JYzEOXsScgYp2HutvIt/maUuDJjnDfuDaXT5JdxnXANopGb
/bgb9HapJfgqeKOgm9BG1w9TKvBd+dR9A15jfoJjm4KMeAVelOCMHRW9F7iyqI6T6CNNR1Z6gOzY
oeFpYzsyyxyUxaAKvLdKP5zDYQH1odXqW3R1cNqgWYOIsM7JOTIOyqWyTMqsqzETv8V4qLvP5LVg
LXSEeq/0cOIZ6pec7ZiZo0Zy/qdiQw+QVlWeKZmlVVn8HDrhLJeAw6qCh0DikW4b1Tqwl9KrQfZJ
GOqXXdA0YWlC0JVILcs3blrs4ORZDqthz391oBpEoGx031PfPe2HaB/bnFbVsULMeTt6BS4hMhVF
tg8lhvakakHp2lA67zzrOPiE7Gpx/yV49iaSdVOYKx7i+fImqha82STtEpYli+8bJEv7HUVMBC1l
7dDo2oezJwxmyMxuOHw/kw0N20ZDa+a/EJENccACM7oUJL7TqG5v79h/LVDbzAojTNr9qhbUz2cA
FQBn183OasrK3xICB0jUHXqrl/o21aobBn+zGI5f0JDBMFp6ejJr2WBXJAdtBzis023fUEH2orvE
Qvvyal4d4/fD4/OA3ORnvhnYW0/nMo+fguWIPODsKjW0mC762QpBuQPUJIpUN+5x0+CxVrFxQn7q
RvzCwsDvfE6PpeDW82EFG1BdmaSCUnCni/TEnQpoSNh25verm8cUunRoPeLEZLdTsTVbJ0/eey0T
0RWakoO2K0xPUgG/Q3DZz5qsUANfuMlU4sbaCPcNXkMNTVr92Nq3/DU2fRS5gPfrP63bKZaYKvsB
MmJn4ebhkJ3m0HHkrGQFuSOTrwQuOnRyQqaDY77xCxVyMBcTsguUVYCM1YmZTORsnHf4R2fWTaXN
VXSTOdvjxSnk2BaLxxupgIu3c8gohMaDw8dYcMj5gTKzcRAtLLBDXrd8Oc/LIPqBYkkdCU8vYZlZ
tyAbKsXZEFrp/nveTH+nOGa/VTJiFua6PhRSkXE8+POBKEmQi0Wnye9mAm3k6R0CCUUPQOUvfjYn
7fcZguBtvzrU+/hobucHp4bGeiCWJuPBP7or1QkYO14Ui4+BIPZnvRqJvUsBN+OUH7HwdYCTcOmg
tjY4rTrZ6tk845Rd90uXX9c/Bo3tnmkwVlWoUiUcepvH0sarK840j/yUIduVI+KF5otA+2UkFee9
Hw5lm131lES776mwEl1ck2nZayu9IrQ6vhYBDxbYRhEqdjb0EYxjUp5kfC1aoAxhlaWtr0VlrRbq
VLuJDLICsJ68n1WELWNRzvMqD0RKln4qWTIuhe1Bbszr5iOpX/i34M7FFd9LT7KUGEgeleKaFYtm
+5hLWTDuElIJZamUrRbtlR+ZvwLW0EFDq9C0TF6WeUBbGo7E/AJ39Nwz7+cibPwgWdsK7WoSQ5OD
90a8UP5qhpjAYY0Svzbsg/CfWfLP3T8osI4cYzcA1ATw3vvMmHZKOKkfUgszdij9GPr7kmwtRtQ4
7mvvXXiXKZRh2wvVTkPvHQbq2KO2m03VfGoBI24j9Qlp4tb5plhYfn3jFl3YFV1SAtkfidom6HaU
h8Z/qwb/3p2IRKONCP0VV4paxEdo5CGprpLblra0nXMXxXvlNXGujmCUWLfrq3WtqJ2CyZnDnwi2
TEL8rxntrXVCuBoXvMwz9aAMQQYreAvh+78GSKOEPcuFhF93IsLG+05jjdGNL+/Fn+7VnwNZQtqB
qlRp4U49HcjL+wrvuH2iYz9SYw3fP8bipDuEEv9XS3ljxfVm75ORblmoefhOPDtx3Zzi00chh4Zl
j+yAo753yXg4cql2uqDzBZQwaae7QmM/wRarq93J4w0j05F/ucQWKgLaQnIPG94a63Cob8X2PNRQ
5G75oiPc37yBxkmVrg+MMt1AKK6h2O77pkQFAzZBaYRZ2ErOuqAH3uIrtsTZyA6F6yl5haikXBkP
ikKG98vmHtpjBk3gn43GBbiEdFIFvuxgSnCBjvXG+MCkAQmfU8Dfkf1M6jGmgybGOyap3zME5pgC
8+fNp7Nz+1/uUrRvY8SvDbGrK5vkUhK7wOOGozQ+0UvHZ0M0Y1Ps1Y7nWuSeAaQlV7l+78O0MYxr
wP9tMSe3Tox/LHN9JK0NjhujNaTVILN81jqfYhnaHw+gohvCAOC1p1v5CSQPQgW8Y8f30hrTRI/g
19uxyd2SkZJTBD9dIm6yUqTk9xft4evWtGCht+8Jbci4t8yaaJoWpmDFQq+RMoJtxa7XZHogc/5M
XaHTyPTmfpKLI5OVWyx/p9igIbgR6dtIGoVptU4n4jpfnJSNKvbhntTL+wudVbhxL21E2RaYZNo3
uvLO/KZ9vX3DwSIi2BWfx2v9NQ49mcOLpg74+iJQOgFMD/54oXaPyMWwcEAPXhniKl+xqASLxgBB
SgFKu6TYRjWGAh2wWE/UvXPDH1dQm6jPQgNCCz9tQ61e/r0UI9volTbgUVgK+UOVeO4S9nf90jFo
aBJSkvNcUEJqBoStYPe6IDTHQ7bJi6x+VsKDPhTi5526CKYgpTA9O6clzPPMDgYZToFzurTd8fKv
aTv4SuPAKXkp+AoCUzSVXSIM/JY3mNT+IjEYCbKEm4w2AmI9iXhJG0pBf8FYBIHokFMKaRij5q0Y
QBlJMh4ykgriLhAfoi7yW2s9zoQZS8RNd1ZB2vKHVtqoQyCDg/yEujVpUpOrB/nVAJPDMX0lGF34
wKdIA47li2uROq5xL3NvegEoieCAudNJbAQ6LsYxw8zCbagaD2vKkadrOBz8b1QV7UKnAQulPFmO
ONC4/T+oVmIfpmlWjy07i+66uqPrzDU0rVpTPKcYCZM8is0DMMLE81xHeV3QbcRmyuy5SfNApmC1
bNy//VDYW5A3tlNe6+UiElv664BpkDYr+Yi5iFyTwY2D6ss3rRT4PnXhOnVSUdAUysHuf2g7w68E
AzaqoTQlkQWu2vbNXLBQH3XPLN4ns8jQfySl5+xF76xcSqVCKbAgwb1IJEcqqARH6BFah7ORWKBk
y7rNFGMRaB1rwaQ0X913Q7E5w5wOOSal7rBIU2GyDPXMbF7za7eWNEeUOegDv609x31hUzSAmU/s
zAyFCYzN2lJOz2ZsoKdmEEEjiDhNfuwoSX3Be4Y933eFXCVGQARcjr2hsMd52CN40O4zUcDWCmTm
YoJNUejpFliYfgeJ1ENCKNYhxZ0iNhk4bReUK10BUvtMf7O4gplHyCwJIkK0tM+XrzXVfFxPMvTa
iNuIUzAbmOpbz78jkhQIhmHhW6YbHE+m5O/jUlbeS3mRFC1xzdpH/FD2cbQl38as/i2mLgtAnNXJ
6w7zbxQjc0m2qPa99Mm2degPGAvdtRXzjMKeMjyFj7+u0Z+CGyGIrsUwxZ4k7+aLHZ8z2HoaPxNK
BocrDJLKIKTCP+ICUoMrXO4k1QIxDnBAAhU3yhHhr175Yv/SsGYcvSk82fVeU9nHUGHoWS88sqi2
hJm+iVkGAgH5QAiele7X0FR0jXHf2JutqnYT/+/MzKBBAs/z2nKBL2ZCU/tkUhQlZywu2qf01aa5
WRaqjhEeLqG1FwfpkkOvboyjWL4P+pcsWX4T+7CowtENx66hfLUIfaiqOu14tnGIRVp7urhdDIk9
vdtXoiYGsjea+YUOPizvNB/m9p2aWsVj8yjLfIpS5X6vZsHG+tdoIUPhnYQjhQuoIoIPXq0wc7yE
YVj86aHzy9g58bWBc5bcSK9M2EVeY5184fYVzV73UQuOjCdcJDZqDhMww7Ln0vdoVP1hi/yYU1RI
1linZIm93SpI27PQQ5YB+F2czVly3vq6XRbDP3nnzYAhQH9HRZF6Yz7rd6R26YRzLkrxXp9jBd1Q
d9nWd8w/V7vB2cSfm8jsfWJYWxpSmIXXDPcysBLh00JxitT58jHzQgPgVI4+WZgFMZUUuS9oPCNV
rBf6Q6yT8otXnddSViBvsIVAQonURCYLr3w9XlBom90YcNUkyaguhpYHIgaCLKSs/1GevwZkwtUi
rOZHfhxjYGw2O+25MPzjOAOB1tEsPC66jMVQwym6yVYLwZ5iZjeO9+XBSzmWhxWOBFUfbbDv9XTW
Qfuw3BEk0+tlEHfa5o74o0wuvPXxjg76e/z/8DJ9O+PKCfCgLMIVcGqZBUyRVa7hILc7/pBELRQ2
D0yGkxXU53F9xwq3pJ4PcSPSMbuQA78kjYFEeCv15VAajc2LpBEdAgG49HRP2tpbrPG7t0d3ynv0
A2gK6Wpd3UQYCN++sdE6qFDiUae53kBBxHJ2L4xcG0EORm9rhgFGLemhPxLnuIfpByBr1eoD8Ws/
XAFlScVJS5ZVWvxEfjxQeG9bchsF/kmX8MgYjvN+WVDvSe/jrsKxTDUD25pimbhVaNXErIBWIRMA
AgsvDKeWj9R4qg8vgaDZVvCFP8VwhJ4UP0oNMA3h9BFv7vqnXq7eLIPM/857tOOqMI5MDIbB2uQA
4sxK+OLU3vw3KEFAYc9wkTH6dDB7Mvq3ns1aXNNa/ynriHFRmoBeLVozeGCdAvz9sPzM5gNMNrkR
EekSZXYYQykV796kt87DJ9q5Vwgnt3cr9qZT8jusum9tChJonBYrp/fkFGIfiJgCBRbWh7I3eRR6
eueN5IxZmKOE6rmww3zmX9tk6TI7oWWkgczvhiFoJ9P3sQSr69bIoZ86yKyhnCwTCfLCYnQqEZRd
ajOikNlG33q14GEdSSR8J8kGebUQQpOzOTjU19wIG0fv+woOK1iH4htJIsOy4mf0CVXEFw/9ZSie
Sm2lglVB2hvQ9TksR95hLBHi7A9mk0NV39LjzuDScTpYGUYIZTlkrDEHaGk4hn52YDkGjwwmYoy2
pM1pyv9a6ye0r/Kg9dwF+9JLCy4QYBZYre4ZYpVtNc7Fe5yDFZA/5Dw5r1yERV7I5kmblPKnUdrc
onVOF+qcn/MTxDctnCGtKONDmgNlvxv416A93rIc5kWUB/oznoOAljmhlaSp71MsPlGgzbfOiiD5
xVaGomUiFTaO0ff/9cReV4RhA8MyQztDZ4wWo/IDa9bU644dFnb6m0w6fzeoecpniKazRApp+EME
90+/DQ/Zla15OJ8sGzt1Q6sPsM5F+IHOj0HYEYMLklcw1S8rXiSzGde5Ed/KRpQEP1A7UhSCZXS1
IB51vqY6r8ydoiD+7SVHf6/QmntP334Vt0K63SWWs32YgBYcmVNh3Kbhf+oiPPpEPw/xk12SodsO
YKzJ1+oa+hW/eFyi7oSZ8MGw9BDDhWQ9tyB9JwHdMEquueONZsoGSHXy9HSjK3LrxSwfhJYUgRy+
LlI+2O0/PU1IuKLTJELD6Po6CsL+PLz9Z3vVR0LnruUDw+5VqT0vXd8J+HjlQvC4duS6cH4y22V5
G2PYH430RcvR3BPmSRiPTChQsh+8hYWMg653eiP8UhvC8bN7blpAMDyOQpFJBAx1TzN306zPxpGO
VbKiG8Jsgn+mN0uALRHJQ3CLsL6aaKxuypl1JjQeDh0R+BGn35kW1zivWZKslmnf0CnxElhMTysh
cTU5o6CpABC0w0XCbV8geU/lI+yNEUMPzp1vvzZxR/O5e8F7xdK8HRP/Yw/Lm9jVb223NpMtu5JK
mNmdy6Eh8kywICcZRUdAC0Z6Df3gs3l4lr0KkRZrjtTM8m0HjWzRxuy2Nyq2ZCQxkJOxlzhiL9jR
lpQzQlCJeV41fvvYRfmc3X31OQr0ATLhVueDKepWVPYbTjpMgFwFnuiAHtFq71Jw7oOqqgiR489j
oPuB3Pejy5cS2hLHHSR39syN+0uq8A39QpmU1CWIsiDNf3vYr2lD9jQsKBSS+iJb7j/jgXDiCvdm
E0IugqQTegh4J3Q6tL6O4JdPzA7bG/cdWO8wlQa8BSMaNykd0SBHQZSvvlib0r4+4lY4OV3p+vib
RPZeRZBf5qHkGXlXEwgM/hPXG29IrT/D6FLcobO25UaFMoYLdqRWjrn4s+bBHVF2QjVQmrlgIYeL
qXngDr1CMJqRWtqPEOT/uviDdCEggtI/WLyhoXA++zWIlgSnWOQjmD8UWF1V5BEQsopr4Y0JzzTv
C9379P9UEg+4ugoGmJlFV9S1xjXAxXchyJdCuaBj0xNc0hihzV/Pn7WUOyBPVUUvagxgEQ/nSN7F
MO5SbP+sC8z8QjSS85IUh9QmUj7WfTl3GgUZIVI5dC1boYUhOdpdyuaR3LLga6onkZ9RxayI9/Fp
hj8AkMTHYqMEEAvKj9GYKPPxxPFVKdJEOkaGz/IGYQubWRBEB9FjXLwoy3s9uuPR+JjKBHo/tZMl
tzGXRjvdsw5HFSffUvYGqF442Gc3kCsEdIYJj9wZgmbh6cnDepgaAUECiWLa4rGTuReWxDNmyDLJ
LfyoHPBWa1A/585IRFptLE2McFkyCL4f5ESM/kNpky68knjuqlXaVmzdAZGvxiToWvHcDEWuW3SL
Akto6xNyPaKBrjDGH5PwIZT4oYVqQgNZqA7xSDZPb6TSNThFrvLJYIwYpazAPQdQeLkmzfzji8wa
NVCBXzwcEt984903Uuzh7QH0xfo3p8glwxBGLXkXCcgjTFUCuSpHn2pesbeFJdiDui9imqKwGftJ
S2X60KFIO7vj6x8Roip+8Cc9Vi9bhiDEk+mT2DFGAKwK+8r3SNg4mr0b2JMyKice/sSnDfxxgEzQ
EOOKW8sAXMWs41hC3+t1W3+uImFK/R5q3U4l2XqGfnuC8WlGoBduX1GKHh6FwtxDxkO8q6DO/BCq
V7NIuviXjIhHnQ0njiiPyrueN62LtNLJ8bNAG5RlEWGU+ucMnSWR+JXHQoBW3gtbuBpeScKoDMQq
gQTNnU71rrOb7/yT+UhUxjCYyXKAcZQEluRyk/5LFovR7sc2IrLVWNGkgxypEEQqJeHWjuA0ytsH
jQF2FCSZHcsuREk+lNTgCEcY8oOEpZI03/2ZKKRy1XEa1IIy7fyph5GIZNDe4Jqgl3kvv35CHxb4
AIlj1diMuIknz/IStTH95NA1yZG+7lEBJ78i4d6Vl2aFXl/gDDxVBmJTxLRIOYS0sRVi8ohLpLQE
61r31sTznOa7cnkL/QTMI1874xl+vQBe/cEXu2vRr7Tzr21UYbLKpHsaOFODlQ8AT2Q+EBP0hSuP
iRfZeoidLtqzt45PgbXL6SIO7jXzGk3+8+9P5oM39LAMuz/ZNYg1UJ0xnGUkaWheosVZCLVdyGBg
rWCfBGagQg8sxqNV6W964T9Ocz8jbgGhxvVLCC3koVqFXjMwIl+SWWqzknZi76u+Oe+ixgk5DpbJ
8Qw1UeKqk/YrBZ4al+DpxIf592M4ACzxjBcr/lQMfJrTfYGgP6aEsc77/HvG5UNLvNnGgmJLixiC
w6tS8fB3WomWn6al7wBqe0fVvSl9E3V3aVxfuKpdpvIEPokuFm8MM0Ut1vNawNYfHoiZFC8YgqxH
G8dgA/pmiIVWoEDYpt9PhFgAQfdxwvCyW0kyT5a5XH8DEcug5EnxIV5yUOQwQ9mCvM7dhTZ/2XM5
tHi278TluqYYc4PAmNshxr3vfEl6ebtoUezC6l1el9JdFjCFDCAfw9MHjzoXS9VAvvGGVce8CZNO
87J65vrYK6QHbdCObLPYad0kh0m3DkxxJJ/Ba074P0DFsVNCoK3hjc0hvzi/2AsvgrlLTHGNnKob
p5UeLJGBzj2YQOv4uW8xLpPhPIDL7L2lXG1rcJDnwWlD7/JTfHVYTglLQMeMveTpczj+tb50koQg
ljCloSuNjJ17zPDfghNd0gUmI5kpGaHRCZpMFOtBpBnWxaGEMuX7xTOKkiLednlIAKy2mSTRsZid
Wh1pECtbNbIIPrr3KP0/12X3eaVW3Ko2ro9Ce03K+9uEx45kLU67eaaeIvy86ZnMM/xL/piTNJG1
OMSbjJiEH0c/m6Xw1YA2rpj6+uY1/++pRoTMStqlMq8Wbvn4V7IwAGFNYFdekBFF6y47tXttl3bi
fTu/E0j4bsCVzuZCRzucvqWG906JNbDdsc4DBWO5XgD0ldSeoSL9sGe0/sYVsdcdATEsFeOUpCjv
w/QkSNNSqxy7aHvT4nI5+PGySmn3OkPV7OyUM+NR3Ni8he9eHZr4XwJrfNdEDxSgAmrdXecz9ipM
Ni6pv+CCBjNZAnapxm2i/30RRRWD+7lAOjRws/4Yv1BxC4AuB4eOsudcSn0aRqfQ3T6qeN4/douX
dpSnR1u9XmqyN+W6b3cmql97gtJC6KoHop/2qUXAV2IR+t6msVKt541eCb1bakaCrNYN+QuRttqC
skLFnXJ3tEIjlWN2emdRbzsihhyk8NupHWRY0fVEZTGl6qAs0nK6rxNAj0DbTkb5YduGRDVAJTPJ
FLMYOxQ0n4WE9OvYdf6Vqf2fJx3t2QgEWL1YUpHx6zpJkHSJp7iXoluE9VdYVfh8qKc4p9HJFW15
TtZ41DRKwHZBRsqGFwKaGR2WhInyFAwwTL+UKJgxxCMpJHFNqgEA8VIP8xJBU1/dfWHk44dkIquj
8Jv1KUQ8kLaWpJUt48zMT8xol24hGDmWYXMJ/DnGORPvjQUzbMDSEn+oOjnWOzJk5sVhNwgac5f4
dGJFP1GZ0rTQmz2Cn62JK7nhaFqnQBd6BkpG11I12Zh/WfsVQnlmGucbnuP8Bln/A20SR9iALMyg
GFu4ZtEZJP7y+g+nLGXPWOqQxpCgTvh9CXgjhduIBuBPDPSeBnZ15CI2SymaZBnmtG+Bn3askMRG
Rh6UHXOLuiSZton5i1XAPDTGNS3c89AFTgVlEnV1EM6so/kYwaFs83/owEfD9FE2T6L0M6PSfv3t
zpu4n2B+5EWu18MTjkDgRC0idRI0zfpW75D2H5TWYuB12sS52w8CgYa3W8hXWOQeeHXF/o5dimIs
gpcnFW+p8DU+6ybkJ75ocy9IsHzMBTaMFpnnbrLHVNd65ykpMfoxEAOEITBGaliZxtL+ttqC3fQx
zU+J2Hmxu8LHrUDHv3IMVMiSw1pdN8hnvvTu0dBHe/fZA4Z8m92ZDogJ64KTNy2D/g1xTXljtOMe
4yQoVj00slI7/Z9gbnKn+YintBmzJe1ojtznzpScogjdMm4IRKUgy+iF791j6uzSsYrzVSM9bnFj
/ThWQv9BNCO8UBLrkl5OL4E8hO0PVlXLNK3NKSjrorEqc0k3JrfVVAFJoggCdSrfqqfeFPGTw9Iy
sYLT7hMNn7513acjp6MNJz385JaoL+2OxzaEAMuvXad54oDL5Ax0Xhc3WvDvQpMvT/wupv6jibn1
jHaEucdaGWwiAJNvux3tefp5uMDN9QLXGSBa1RgSEfga92/SKhZISARYFwtexJ3FaFdnM/BKxW2V
y2s+22RMeIc5rPBaOy1Gz+jbLFHW5CRsUPuWD+gD6CNoDxPwwINjXl+jFEBkBhgi6m40leyoBUDb
TE0/+Q0yqfzB8lmmcmq+uEqDHBn7YV5Basr9Ioid+Q8nY2GTpf0RW4ZQRukoquAyvltrg6IqgLtM
f4kYkv2M4k3UsHNeIQO4L7Jig9kJVa7VWvikLf/Mgaw2fuhc1O0y/JOhudAMf4NE5QDHmjycg79Q
gOYZ274kOysbIMo+wK5uHPUwOSslbIGRg3LOwdPzkb+4VR1qTJh0NfqyfU6VohoW65g6iHOMw9WI
9Tu5yK4jqPQV24t6bA+THFsygVaHvy61NtpmJeyKFr+K0GJCGTr7TDdyGKVEyyyLUbcA8j4+mpDL
6yzDR1TN0i6JfJa1fWom8cjmSjckbK5q4zdrOp00h0OyMRljwpE7GCepS8Q/H4a+kN2NRIwR0/gN
pn2fS3A6qTKPMbwJWzGDBjJInHs7LMK/fAnlvhnrDzcARAw7aP2ORdGnhYLmgQVKpOvqpVzn6sNL
vgkjAzHW9/pSbPfNBUFrUwKK5HukE5Py6c5Ll/VsVV6WZ950MSihVwMOi2PlwVGrwOaoB/SmxQb0
iBQULuuPOQ61tAc8tnUCoUPs+1gKzQklveoyHnQziyjS3kB6HFwCSevmVrfgEjnK6Ln1I53ABXd+
f02DmFSM/daSsWAeGhAfiCS1FMhhd/9PN6V+Of1ykh3uqZNIz1Z5XlAR8CTXU0hn6kvUcAa7zWZC
/0+Ftr5mzblS2TM5sumD7qrK3HwPE7OHWvYN61pIle9fSaPMkJUcmb3grjBGw9FTDnI1IdSTk6NQ
sQqfmdJ5OZidsvtQOhGKn2GIy3rVLKeWgNG6PtrsPxUI3UWTnobsH2U6wUfzAD4zNtyWJ8bH3SaK
/mq5j+eVhbwQAX8Q44BsmIVZXSQHmKArPymfDUIRhhJ/uk97l7b4AEvmTOJfV7IPhk9JKMfruO7/
ERJL4gXI1Uj/OjI1MFfq3SeJ6R7NOliKjzexCYUGgKtYyAZz9iWGk0SjQeR4VZldXQeSFOY4VdfW
20fXMTKfIe+Wx9t4D7NUa9WLnPIHq94aB3pb4iTGhTymQCKNPdUCDEvxohYEBc5wYRQjS89zuxKL
3NQx8EqujdbnpXpcQQDgo99HMZ8MEt5A83HFkLftPSDgn+HBJ/qcPB+BBVgwgG++vEMCRL4Yqkps
+eRJPrCuz59WdpPOYM8cCadJRUUOIrRrxy8FmmIHa2SKHg7jEooW34d6LxqekxSGOrFJpwnV+QNi
HooxtAT06wkJGqSrIiC1ouM6THiSQZhiv5dDh+xJlUuH31A91OvjD+MGeE0cak+HPzVgB2Cwoz4z
ELYNK7d9TXB/4Mxx+XlOKVnOmMpYiqbHS2m20In0gE1RJ0MooRw3Ps/69asZ3MLXuRYgw1Ga4TEc
sONDqcsrwN3A+TxC96cqt691UzxAOB867UHLJCaeyAQLC1qmGeCK+ioXQody0HnyTbzQL8ypOEWQ
VlEaP0hlrnGa5bBNWd4mqJBK6JoYD6rOuTnpkfLQowby4yl6DhDiIeRzyCF/z/UiBWgQz6EIKNEQ
Rl8iPxmPiutOpRTGatkdmZwUjp45pMzPuweCkr4bP2Bi2e7voNCK24EUzXNRgvE9nRBnXrFma3Xk
cDS0cnyyZRbSWEyNR9qfyUvqLxd6w2yIKrgN8tZsWzjnjqU0NCxNavEXHJlW2ZrTJEcZ13KLtHH/
vQ4xUAXo1FonHKRlS689GnJ2LziIUyx9aUf9hZLyBEeijt3kX9+JkcXoFQsnnzWsIF64W08bx7V5
nzp9s/JN4QiQxOeik6V7CcvIodttx1XLg9Ed7UeDwKJgYCwO0KHvl/Gw07aeIWuQiDg6IoZ0gbnA
1hFK8WaCvDfD710wwyJfU/a2FJQdzyVuUL09GbDJWwQYyxiY9v40Ex4AUjKHd3M+zeMabAGeIVYT
WOWuKXw5VBGm+pZ1kIUaKi3O/oswzTr2L0LJCLC9SrljgAgCBkzXBLPQBVlTjJMaJAfDZ6qC7fWy
9Co4a1jcG/pll4RTk805pVuG73i0N/lwhNsz9050AWCqq7uScO6ZrC7A8qWbaMOml6heP3Jh6XDk
AV0F4ci2O1jRJJRKDlSq8LUOr+7/iqeHh3tMTQtnMBMKVgBu0tFuQ7Z8kmArcTjC2f/64wOMCM0S
Wn9TRfExKmvv/mp6Nx1D09lSfns2MUoMyDf227ye6eeO5eqinPwpTMnmYs/kzFjflwXc0BfnoDlv
0IU7slb3u2402QCzFtWB7MytepWaYwIlTAwK1Kk6vVdsyPgbeB5bUziSgyJCPzku7HM93ciZOQ7Z
UxjtwutW6XxbSfhMb043i5voS6d3UJTXYWdBWBzSAlZletu156aeThCFyDst3PC0/w6LO1YTm3b8
EGC9C6KIQSgIYU1y9IyQ+Lk4fnyeranv4kYCtRCkKuHVrjLC3+r6jVXQ3cLdjVFUUS7R39kzE6sT
3CZtRyYjikKdkRph+FJhKO9NuK63yUg1PIOG02i9iXRbfHRJbvI++e6hx6Ig36jRsL35upd73VMS
hIYr+YHrhzyku1O60Oh1sz+aM37fuxhQmoqm//Thhq5lsvc8hWT8OAyMj+wh5Z4rQ17/falb0AjG
HaU3xAWew8vXp/ryQUbPXtTuemg/Y4HZzeTMDsAdO7YB/jI8aV2CEb1LvaoeSXA0EG+p5puCKUO5
1WAbsVwnRQyq15aPhGEGBNFmEG/EmXhrI7OHi3nKGPRgucRHnzei0Yr/mpGTxBWa9VJyZHgL7Nwy
+BIKOBfapZ/+jimwtUMRHdc01qWTeV4Bqyq1ZD8cnlB9ngX8EBHZckDmHQE1ezoxeHf69KAE2qWs
w3vhfcEAQEFchgEvasSFk89x64gybej/noY8R2rfGdSrof4TAeGFBK+Agdtau44SFcnyfl9V0mF5
9cEmQhd1S/xURG7IFPRV8I3R3SiEkhtXkuyomXmvLT4uwq6/kCpm0nUfMEAmudJrRuEMUW/xwXZx
hQTKKP06rFAnTg1OlKDNksQkcER5+MT/1Qobhj3KvrC1MZAY6W9ELozqLdzRXsNToeyojZBsRydr
FYpzAfwgxIlkm5c5wzzrrBKYI+A1U05+xjvDHAB4KoBDx5PbdBLdSkrtYxXqB/01825HyWB62d8Q
QzHAYO0KyQfsjCzbBr1nE9cqmfEtkX5+U5wL3kCUIlB0oLYvKkeaKKUFrUqeLLTj6eJ82ghe9c4T
Hfing0qlB3yIZam4IYTmhJ4McLrZBOlXGoDx8lf7NX77DK7nM/QomoYHecQSMlAjuZgl1ftQMhDL
oS2Zy+tYgSmkjgJqZ/a14SAs1RH6VJL9GtmAMffS+Y/qXvqpIAuOCC9OQXz4bJpSbBtoQNXgHEdd
DHUEhycDZsi3JXWqH+MjfkyASbdh+5wAMB7mvZG9rguOmgbaIC9qY8u2//geZiPVD+jzsCN9ttmY
0M25jm3ebYmBTRTz1vx9i//tHIfOdDRtcCw1Mn3WxJCgDAjVrApNc9Uxikge45x4zXxYBFCyooy5
TasZ9JqA4JWA/67cy/sHwjaTTcrWZDRBWw2D4Dd3/o5G9Qso+ztqs1DJ2qtYdV2rXutTOAueb0XJ
tzIH9UlpJyjSVbXyypm0/Hy47ht52e7tQSFDEvbz/toNJTnioLVFONPkb1OhhH3njnGWkoLznf2m
DybVY6qxVbZeMtJkKLFs3xSbIpxFiNXhcJl/N40hJEda6boib9YVTkMVFjiZb2GigRfoJQd+Kj7v
60/sMlG7tiiaX5RMKtsLOrECRNXDd7vN7EFD1DSJ26WIj58jTWTUsAPs4IQLgqFxTc64nmaLwnhD
vUr8i35p9mMkQ7ZWgnYOfgNga2t0QyQFvcGwG6EuyY6uj3kNvvUtkNJ1UmGf9+D46jjY2fXubK7N
z6Ntti8oEdBF3zDarNs7+5SUWetoSrYMX5koFSoJCYn7z+SfGofksS8wjhfJ9FLLgyyKVis5NFor
LYRvxC6BXMWoXSRORO4/gYcDo0w/Zj4Gb7zYc4Qc6y0Eke3u5QCnfYqw52hj1B5fJWTgW6YSgda/
8atp4wRqUtQjPXPqLg4lPnDL+BgjpV7pTIDwpZREGhxCq8q3riLFeg2/5CHDAaa1OYbdpoWZfyVE
QkuJUSPgUDPCaXhfcjDpravYwr1eDyzZMCMedOmV3HFinuhNjhJaBQxkt1UCzbzG4abqoPjtSHoY
40XNr9+OOyrbpA8LNj+lY5o4h1+mnMCBlR3F1xYYwd8eu1iTJxDQM2zerDMYyB45pWugpae8o8He
JxEphT0Ut5DE+E3z9gIy9R4l5S9mpgZRjMvtzMxmhxz52YANTOJnN8Ax6BGgkqBLAenZ5du7mbhV
0HFTj/4R1VSmYhJoPctrIHMhf54jQ5sUMEG534CwAt8znomcSxxZJAe4pUeTLxSehBBfCdUBWU6r
WhVPEW5uT7AtzvvkIVsR4JPhsIRxOaSUI6808a34mM9urw88l9NLYyoIE03ckm5XNdevfsgP6bQS
3VxrgbP/2+gpAD1nR0WkVuaRocESfSHb0ey96GdbZjtjLr7hl5n8WS1nH8RsnhcAsbTE0fmp4KK8
N30h0CsQUvZ95wc6xH//484hWMNP1EFnckGWj4sPvttG/1cahSCmKII2dmsNNF501VLQnrdKWguG
jcbzmrH1GKaZMwrqSXwVsXbMgPiQHx4oCkLcaLSRz7SYmkMErYqJC2zvMmBB/dHSuy3fFFParuMz
Xq0Bwh2dGl577X8Cg+ZzC87p0ZE4Fe+HUv3qIqIRbfxqpcRzOo5m0EfFOCnmvS0tXqYF8+MEXatE
FsYopdyHm6pTLWNsUh3ndFpFONfLbtthbu9yy2y57izLgf2Pt6LI2C/18NW2yKRCGEGLFkrQr9zH
S3+NoPl5emo6VPnXIXWzqdOn9KFnGbuYeoF8lsAGxSKNp7xJ9eywLOPn8BfZXG6TRq4j1NUX9FwU
5DJQ/CiaFcQYf4gxlg0fA2M0bLsIqlNisinz3QZXGLPXh/sKfZSppWrG2/MTlob0aRiwFbr3WAlP
dS0iRTUobRJ/TTHKWTomXPirFAVPNzbVIbtJSkx1CQCgNtU3JOewf1TiHmIp0rvlm98vRSwqTxRC
xgAm0xCZxlurHxV6tgFcvH1O3zWrZajcbBjjTTW2PTgG4W70Gc0ws0rpMBWZ97Oxay41uB/tmE97
Hu+knQ/NIs2EnX/xSnMYKwAadoDaD4h8bqPolpC07dk3cfyNxPbexd83EUEABBxGguTE1M8B2oYX
RuMZcCQbpviNye38NIdbjpuNffkcxhU8pFrQySAYqv1wA0fZ5auKIDqTjGVSHx17s+gkPFGg8Gxq
ryjTUI/hu5iHbD3jX0FJRdV13/yQgnk86Ipx7fQsQEyVbQgvYFf23eAQ/j5T0tGPIz2njqwlXaXd
tgRzKGj87QTHS7AkFWVGfHnlLmkACwbCh8XMoEIeFL5U8FHL1a8JgIFeNqlHVdyizl0De7f3CgpH
l1OKav+1J+ZHQN+qKUGGinWByG+fjzufKtGkgbQjQ/OWEBuR/d/UZTf/mV5MhzrN7gFeSUStggCu
8L/vpuBv3frJD/haB0+6I2j4oEBRZ1b2mNNLDQqY5fyfD7rKzIFlKrU0P04DeeKby7iD++5gp/Vl
OmqWA3ImblgasKCFXB/ZGx2iKnWAhxacJ90YhFSpj9Q5YiyK/k3bkSve+rcaNscWRQVzHSFvvJsY
flqAFENUDnBQa7RSWBYLd2aWE0oVxLQZgSCFjqvntRHlqjmYfJnH71swW7KJ7gcI4TfjM68zTsJL
4daGAusXfVinwlkSfQ5VEXriTS4VRM2+OKDZD6+0+4fq8zLr8W7gX/wbcbhOVLd+UD2zBbu0Bttm
FMUH5GSKK9PApCf7o5dmO84cfNl7lj0uEwBJCNr4fixm6OkJgv3LR6rApVHNt1KIL7nDzg9qZaI1
iz0WbW37c2gIrDlsLcDcnYb2whbTBNNfj6RoFV8L9rq6e2GURRwkZb3LFudWt4fSC6pIJpGJ0Ddr
R172hktpxWLwQD9naMxhN/W+JI4D/2PRtQISLNFXb9R3vs4DQbLmJSmVjs6ZCwwMMnVG4K+oBXI6
lVOB8c1ceWJ+AJQ+g1QAwi0tEoW/W58yFQnD6jZ18fQg84ediYIH/MDufz7DOmCOWABeKdQlV6PJ
7cwrDFDoks2/a9sMJaxQv6kdPutLV+119IyPilbgWyWLsBbI1meTQ+MVkf+rF89Q1Ed4f54Nq8DI
GbabnOMeHDg+ZjRbdbdU2179G5gXzbp9HVH/vSF3UWFlZO3EfpMbfzSyJ4avwe+EgBu/HlGqd4l+
TR17S0MNRB5NqxaCx/DOFcCrx9XWrccjtC0OSRNlxfQXbvbKF3npq5CUFIh8w3Ekl0ldwkGA0BJ+
wbHhRPXscZzVWxfGkzRsgEw94vwXIOUtIMsdGjM7V1Te5sWLQSJxfq5MucoUNj5QoBQ2uD2lr5rW
pF1ZxirPJO6mkLL+kzx1ifJ2Ed/JOLEzd81HPpbcLISF0Q9nrcBEA5eXG3wDUsDjEyVJbMPhKvoU
/5m0Y9EUw6lZsYo/5kKxSU+XjSdLTeXY50OiDhuhmB9ZrncdVGcPcSVmHES3fASsfA2YGtE1r4O2
u/mciee3ZweXq7cZTC/WWSEiJMxfye2Owjf9o838njRe2PwqHDXuv3EFedsmKZZ6WrIgKRlWYZS3
4VAqAwZKXPCCZAXFKWlunRl2AXrSLOCESTiZI/V0dPLnxUHNfReV9xR9IDPYRskrMWNMh2qM64OI
37JWNrgeGn8NdqRO0YTj/PdlJnu9Lw47olSff3iccxN/ZS6/1e201EN2UNs6DzGLcYhG9AkxU/Bk
0M04bYLr4UObADGg4L9HJu/Z//7pso4/q/4ZK6jYngM/iBV4Qmkin1TRJXkwW7x92W4/BRTMzsDm
c8J5U/2qlcBHAmrbjSi6sLuQOlVin6nM2D2a1ZBCpNS+2+2vLUAz/BwiJAwyk4X3VnhAkB/b0b6e
SUmdCBLnYYWNtHTkf6NmCSXSfjl2ab3RPUQyHsCjLhatCcWo/RAuZVJ/DxtuhrjHcurYh+R0iEdo
tfDIhMFaatJpFKf8xcInpwvOjaWl0SlnCbXQvj6tMy8yJMLI4CdBRjnO1TnR2OvkdTVOtEadfzCZ
a71BtVzElGkKxKf35lt81y3vRexBqHhLyZraE75Eu6F6ppwwDQtoITX95V11z5Rr1Obe9/Gkf+PE
ZIPcwUqqx/6yJ8zWXT0a7r6VdpbHJaF1xSfRY7HD6KkocFjxXwbyjpH7/LG4y+C51t/fqqOazdtk
6Mm7xGe+PJbD65t7KsqkAibg4c6kCV4Ps809xdxHkWfyfamSdpEA+4UidwbOj9qMrirvQDkZeZHi
7wdCNigMPoZck1ZMP1ya1iuGp8saDXLqRKsjWk5bb44kqEJ2lKE6um1bWYvDkYhtqksmnhdwb7qX
ohBZ7cvygimo1HUcXmIoIzcdLf/lQOfs7vIbpjcDzFr3R4jR0JsWF4ObXVXvzm+vqURDGWzbX5NU
W9ecZShQZGg7fmyGxw4ZbUBKHzvdyROimqSZkrbprqlDMfHThzFd6FPubPWtZ1Cc1pGB9YBm2T54
HZz9XMFd0rHEvKGaQvUBnXgEPKFactQhbxjbT1/+GGC2FC8xXGVryXZFj1/vVV8ojBqe/THbFD0r
OUSRKlO7U2zo7oulGm7Le6DOVetS7P267eA078c7A6X4Ux2qPhQVDDOXMaX9q0+vczy2VE2kZdpa
0S/FaeETPZaXww5YDehdQD3JZz+acDCace/wtqiyNX/kmCei8W+zi5AcoSaeI2ZehYgzfBHD7gxT
4+869xysqtugzCZFbb8co0yCD8kNv5tWbnzGXPPPRDSCvIVgVVD9pjT+gqfW8jf9goy4fG7ODfQO
286F+fWZYXNzMVUP285iqGNIbNCB83JyUwWqkM3T+FTXn2VbtMLTOqeJknMDtf/aAbn9VSFHiRmo
QoPfgPHdxoSTt+1MNa/Sn2Xs2fuBx5rVcSRvTXWApitiaZzJEuTZvNXQdlp34IyBnQWZQ+NhPn0n
SKPg15y+r/LaGpIJqCJxrDpGKwHvt6T73m+3CEicC8XuEce15mz+bFHcoEw/hQ2F6/6q/lb5eqXD
grwvH7mpMz0yeMAviRFjd8B4Yz3jBXUw4Fh57nYXNF+iMr8LHGsO9ro0StYX1ywI67gCuBtMI+zh
bVR83QpBvs8kyO277xZP8FnRRZKWRn7sGk3r7PL02XRSUvrdqLVaahttOkbMjsJ7pN7uPub70uT4
M181lP8ub71REAdysCfCDhUGCMJdEf0A1Umnw2pydZ+7pIzJR809btQQfeW1aXBD7c7c4rBF+A/N
aJLhLvoLTZX7rfFLL+cFD/t5AqOMJladX275R6WXTfdU8PhZnsQeryp6LakuieuO/Xy5MM+F+eMJ
XAGooBzUUi9KVQcuKQedx8jw1naKgCrVQ3pWsulg30CXnDJ+tXZwkA1WjyDYTYRlVC+OE980r5w7
GrDS76VhB0hEUBfH6eNKMkbwKhhcnqmcJSkZ8yUAWJllA7Ege2b+Rm3iHP4muE7DACU6bvJP5AIM
OYbDYhmHlk9/8KBNY0g9FwQcZoI8MAepzQ4UMegP/CA8XEsHCPYwaulnRNp9xD0OBDN+Z044zPHx
pO79UbM8q6oL0Lvd2Ged0VHXfSsf/gimi2tAchSfxyRGmN/PR2Te2OlSyoXElDP0Ads6t19ZAZ9c
sDAsWreyi7n6fhjTpQEz77Kvm5DIjswan4gJ6WaYwFW7SoHRr30PD9Se1MwT2+hQgaTnXbSU/Z26
SA5QbpsHV0ewd8IxONj0MwRt7pinWSOzynislhsNXWu7FcTi++L6sdj+eBZcelw4iKX4IeeDv+ML
ULcwhK7nITY85FGYa/ntYdVCE8Pi2E/tX9nEYq9dWDcW2l6QG+WBlA7k13bT/Pm/Hj2YTdQdMRfK
7Y5WlWBN53+JbUuVe6wIUcUtDy3gA/9qbFZiTK3gMFsFJLQuDaM4CNziZ2Z7Ie1NLdc9owc6Hv4+
+1K2oYwWdVU9FWBDvFUn/+ZAoqHqYMBPr+K/pQkjpOz2HIcgLKA06qRlLfCKZx7nfgrD37/+jiLk
MPGCFnATodqWvMaoxLuuFgHOVeaWDp0sopx5KBNuEZx/Z5OhiSNUlvc+fnOG66Xp/HS5ZJ/hjdsD
7boJG16GFN298olvsebydkqWzMBiX+Qe2IHDq6GhxAvuRdwPfnoiKMuebBaKQlFTE+PhdcQixxTA
W5KNNstbgqKVgLsW7XAOCn1bzLj8KehsDDeKonBwWPA73UNltE8pKz6JXq88G3q+8oVWy+Huvk0L
s11knJKDynRxTkVgyPfWFQ+F8FPUn1mjLLT1u5dxd3RlImJnTB2JIprzhFryNjW6LDCGXePXQbl9
P989KSaI8dTLyLcQMgfBK1mhxEnx6BfyNI3OuoqOt1H+uU2dgPjzfdI+r+KAhygvY0Gz/2XusAdb
Pc47FQMj4nchy6bfzTqUPJqZHpeT4CZ5A+nWJBd/+xSB5oi4D5kjvGh98nHlOUEWVpi48atwnQ90
OalmODP9EnwGdw0M+DOkZp5CO6m33TtlTakO3tAyCPVKVIHHV5lHaF2aqxECpLCw4fbfMnB10jNV
Hb+BdbYfciccdAru0KwkAiTPLR/fWx4VI8i0A5mr2dlVY84pwcLgI5ZNXNobPztL/z5qEaiGwlcF
WWAqbL3Z3NrZdL4YafgT3NUoolab5gTaw6uLCXrxr+EqyArXdKLrl4X7etMP6n8F1Fbvt33Z3o93
wCb8DNCcMyD8AHfFzzPTlogy80SIvB4wbkHTxscQ9VJXPrk6/lBqWmZXR2UyFUBXM+DnDkSF3D1y
eOyVNugpO20LIygGQ/mY5WQiQVkXqPpVwWXxMLjFEXRMQklMl/IQ+j7VsoFs87e4ny9wu6pG7k4v
VjhFeWXwrqN0xtHEeBUGzyeM5PR/OkvEUyZfeMJklOlOywHeuS+sDOzHy2EyYRMppNwzfpUxGPRr
xAEqzrzenrclM590ZZf5mW/zAcvM7B+ODDO4edq6EgFRmfwqb/Ww3938WyTbFS1wAKtY7X30RZH4
3x7BATbsPSjiudPdnoUr0BqRb0CRE2uoJOH0ZjBaFxkkeXWp8/i5Qsk6P0ZXpHS8qNKDsiMZtoYW
7Ynfomq4b/bzup1HuTUes3DWayfZkMB8AsmnONWw+RpkhXhwsv5px+qBPLrbdYt9fioRWXOsQXah
80sCr5KKvFmE1S0djlDsEQ+pO6iQHTb+haHOZF5yN7uN5/7nhxx6V9UnxWiqOiMKyc0L6TcBnO0m
KReULnGcGp5d5PG0zFbgJeL4Ll4vDI33tN2ztsQRhCX6tpweFubFpHEyHdin96dQKFYCIqUymLMT
Aa0rcoaW71ouPwWSdqo1ox+zys7jwvvLG2fyBxIkuNwoZqFb/kBR5pbFT0ETq1J2IdZ4gosdkt6b
pw6/un8ioQSQLDKDeQFpmYkl6M47tEDrate2bpY+PGL3DDNYekwV1WsRAwfYZTa53FcL2bFrnv9z
38tZq4+/vOMJ5b5OZ7qlOUZB3od8hqkipVmo9C7fIrzwu79dp6vvNkrD4OxOjIUWb2eGbU7OxNHN
JwQmR5V+rE0kyBL4JeHXkwQ3eMIvI9HzX9bOFCS6MCW7/mhHGlIXcWg+6qvOyiaOtyThaauW8JQU
vK6M+hNQMUQmsUybylbz0s6zaVhm3HL8PEa4SSul9vIRCTJ0IXNtDPFiZ1LOSttLCB+NJ8q8l7bI
xLjshEzhGRs9L9eIhVB+CaVcNmvW3nc0qqIZ+EM6cJSfXa7+02fAcbZWNPZV95dpTlQqnTbRZq1e
4c8kvInenQYlJoCQ/p220DBjjNbgql+Vw5ydAQOrmJpbDDD3sAsWtD4Yoo4SYFHMZMvUJHmwDHDu
dTcoBcFnZPncpb+hXrT9kX85aklu34eyPf9/Ybur34Aq+erUoPl7iMWUdXOOweeMUuFt39rgKVIf
652G49FwYgY7BDyqE1qZsRe5OAVEOh7Ed12YAHno90fImQCW3WyNQGS4FY7rGF1L/Lh1dn8RdN/h
SBOhrIOItk/Pz/VsG2A42YDCQgvhJvt8jzuRpwkJ8qvxDZgt13b2n5EzKsv3zWTPZ7AXq/rH50gr
R30YC2xXBkZqPaRj+bIybKffDrOHBshzhc/RfCHg4JyzwGKCppjLTprMnLKs6zbLpys5kr50TjTs
7rqS9nk4eKb/s/GvtJiOvc7xqssO//umplCGbhgyrEXpx94qXGEmT+g2DAeb3dH54bMxbP5UMJ5Y
aww7HwKPRo/cyzwvEFVhbAHPQ8CKWDX5rva85XC6B3FCHwmU5IIsVzyUBOaYA/9o0kjLQoNYdK43
ObJf0qsbA9gDUUcfcQmE4qzTcgZk0DsIIwmOVh/9Zj0CmfwtSXO7dVeNtoCu6DriIWls1EZmsKKE
KDakw1rgbgxu0ifwM7JUgxJzFEHuUCgEv3jC+qvql0bVJTRDI+dvnmwNrqLZTQeU+C6ZkiB17uys
eP4TGyiFxOyw9kkfQYV2zvNJ7ixgqA9mStjRU6UcTvnJtMvKth9YFN7BhMmeEvc4JQ40MJqjEgy0
Xm19R1bqXiLYCV5kljvHjsRuNxU97uFWwk8Z6Nn9CSyWUt/rANC7DkTiCiMXM6Mr3wdlIUDiS9h7
NY0DMJKAeCUQhWqIHXD0CMy5kal8rEBR3DzgLgjYCenmW3acze8i83nXLpZjrb1jIY/WmUIhZv/H
wXALu/nrTneUOqaMnGOe8HRz6w6c1F8NOmK0fRKQ1y81eou21NkO7T3WrytP5kI0vFQfGwx9J/Ir
yuZykKSbCNyVlJjcHcvyeFULawBrDCPEK6xL03RWTtk98JNVCPk2EFjnCvHzZvO0mp6iyyMG31XV
+ONtjLcIJh8rm+45ElsurDGYNFDX5vKe9v4ZT7jIH63FzjVlbu2REVVpO5vK0YRvvyLgdMXldQU8
71w8Ppr1uK+E3Dgr1iFhgWiG8cgRtBdZM+ypaco73scGdfupfXotLTC+D7eJqXX6zg5kESRbJUwL
SxK6MBQnDUH2X8nNMrhyTtC8CI7RXNCJFneeoQprp1mWO8Ofvymueb1bKcQZurCEpzEdlukwzQGH
8/dcGuobQAirk8ByJeGlsu2ZEXwJ6qjm+Nnt+Er3P4Knd2edSc4DKjz14ta5myjVeQEvlVb3flWE
4GJlzRReVTehteCjg/gcbJKz72fNSdPdmd8V9o1CRJpVhO2ONPMP6vEbmNxGnHhDpjB1prs/j3nr
QDUqo2OneBhPBFRYie2psGIHXDcPFb1wuO2p4qYDv0omH1vKLY8E9WiRpOSDwX0UyvW8QwJ1gxFZ
nzfzdADKvVVr/GiCU/r+2RAcq+QGHzo5w71sEAknSUY48UyAHYhldCh4ERJfAvYavncEa5xkGhqB
UJJa/+X6h/Zet+/bHFxTDLMd34wTJ93rqxeGNy33JJrIHu6YDwNBBjqZTV5XPL8eQkTbdIFx1kN7
N1EzdCsB/+kGes7JAvKLqze2L7QXkxldmvV2fOZIGso291Zi/Xk++jqDM+sdZcZv96BszFWP9Ikf
DflvSxpLs5hnnDAGpPiP/gV8SR1dkJS16lN0ETW3WljsaloxYb7QCQIRHyz/nuZIVKjpqOuayTVm
jYUFb/KiV+oulS1SZ7DrNbwIIrXZfTiSP3ovvDBBpIPsGQVQSQS95GA3fc4nbnQ6AG16WBpZd50O
37nsV1Kp30RK7nxuyg6pPH+vMMgoFCeQVPQacV+4XwiDs0H1saQb95BeDGHcyT4sKMgFh+nDGDKe
xHo/UKbEilRBpCDcbLDxRhjoQtUdHfVxT/iICnfPLjcCOvdk93C1VyEXc3Ap+OKXYcLOcaRQ09zf
wdPyhLWic8PzaxuV47/C6Y1F8crtCVf/ND8S7WbyGt155fhjVLyDBhWDeEH8Mqcu4yB/CEKHypzQ
x4xv+CyEPLd7sA015YHRd7koKdx8av2puVhaWeTuVQ4O0bgsgHtrn5iTZXltdfWQOazl+My45T/b
2FhplL3asKwpGiHeLMRDQn6e3HBC9Bj1ZHJSLa/Je7mXZWpix37iLbf7sPpLdCLJ7Y2HZRs26Fpg
zFiGmuD//6aqnt/gqYG06sVinbNUrP+3t9Q31g23JMVpj4Lw8mLGTmyssZfrWwl41R7bRTGQFV4u
q+RcKc+EimekJjR8PnML68/vn3KQKHlX2H7mdxDCjhY/SxfCFJ/BtyOjXHCRh0zf33OxMoV5L25V
zf/yBcWI4Us4TF2pvBNmL+ncRGsH45F6o08OQcwpWxvSBhnc3PfgpQ3rIAVFgrTPwQyWbskS/XR5
TMRD2GMzIEQfiprikyPlpoxBqC6IaFupN+adkFhLFYv/bjtD3c6yogqOGulPkavQaxeuqjazy+OF
YiH/4X4JFnCvELeZHvzqcdQ+ObXzmVY8zms1mQA4z3y2Rl3mCu6yhE1xYsWIv+Uo/XHHUZ0wKMci
c8U66h/DI5KRf+wduHceUk/l4HkC/exOhkHymOZduxdA2obNCEwgQszsOxR4jfG3Y+qXAs2hKNka
5CvOxljsAl3uQ9gbEVersN5emAKoD/XN6wbYH4h/LdF4bErEywcbuDN1QH8/WGnArR6oYpxLVHGf
a16BJLP+GWbHTPs/ybA8x2hl0XiVf4nx67k1PTbF1PnCGhSwUvl7t7eFKhWk9ZHvZiJfc71RPb+I
xXjbwxDqcs1dPJ8F7jY75ijqcpC5Va1JLStWmDLHA8x8WEFKn+7w8z+3ZCvFQVNEg6j0CvPLAIQK
ayQ0mLCkJ02RfgryltNNO8G+RYUMRsVWxo4Ge651A9OInf5uVyyIlDBnjEZBIYIqzDAd6E0rFIox
If/nsgYKi5NA1FovmRTFF+3yUyKaZmNz6X1Zw8kpfi9XgkZo4BA5iXF49LF1MApdgytd8uXBeH8P
AOR54FjM9q0/Zz0FtYKTLOv3nlPH6IuKVli+gWF0km2kfn4emo3rv1YZna+yjLLUu9PAHvaUt6TK
F8yz6HLPrrWh2lPZPQl+d0Isi/lZ/nTpp2VI8ycOjA9IiA8VdeHys8sBHOodmsrjc/nq5c+En61Z
cDviYQbvWdxmQVpDiLDvYszT+3BYqA3nsl4+SOShIHPY8TqmuMVmW8HdT1fZSMH0oI1Mhrg1mcG7
puizFaO2CMpgXRgsgDMPFD9TnWrEHnxx2JNrqS2gGNnsSnmTxbMkIk7YVp4smMHeG070MU8azL0H
/KOz6erniQAVb2yu0Xvdpwtl4+On4pmIBlI+DqvlI+J9JxN/V6CT+d8dx9KhSq9xmhVaTwiHa9B3
9zWHX7WjY2WU+6cD4nsZ7u3tUTt8bSTiBFjdmwObk4hFZQzRmkHP0jRVQK4CcksADRVJSnBN7AeV
sxj3cf2QwX8DlJmsLAQ9cp2uFO6bTgKdOQnzNf3aXML9LN5wDwgpNzBw1DlOKKuBH7eN6VjqNV65
uNMLzl3nPxkDo1gkdBdYa3pbqjXb7+q1XidBT7zYTH+NNaFidU8xQ/DRgPItOoZK8DYL6bv6I1OS
RgNkmaqHUyjFbfIyxCsc6mn6GaqOnTIk5KBXHBnCXG6nuuogY3Mha7MhXr/G4UGAhwrfJo8TPGrB
CSuEVLMu1rwBkKfzwaoViWBhAB+T0H2Oz4KLBHL6ZLy5jAjOFd3ffbfMp/WGfs0hLlLXRoTPuKp5
put3PUtBcP+hmYy7lO+CylceYmXUVGwDyjQ6Ykxic0omn/n/3JwAVuRsXNhabwnZNamxNCllLGK8
pXaevc6/ih+0nixWDuHGcB8G4f5teKLjKHpvYhY/6vjIe0QA2c/r42mKdFCEz/jm71bPa1rD3oXi
zRK1D/xVwgEuP3K4d+zzFt53mWNsrGLeIKYgIKcQQkV1kE1xHQ7C1e2oila1eiQxIMr4DN10L2zE
9HlqkSR5OIhYe2+9LB7CbdBZe1OShrn7Y3P8gVOkDt/tOrwlElUFL3IiLBNYSZBmReSMZqDqCyl2
6kTjXX5Vz4tmKCtOmcC03idWtyVQYh2jNDIevPPvaoIpSMot2bMd1TvD0/T28A84E2rnXm73EWk/
0bn+SsJFJFHFU+gYHzUsLBFXFY2J/p+cQflG0/FeWOZFCiiA3u+YlVkAe9OnWpkfETru8WJNOYvW
8hePwBi7rS86VPB8V2GSwYyYZ9wlFUWLtKvXnrU7WltJgdUP98So1xyaxjm53Px6EWslWfKyW7+d
QF96kCboub97dDZLM55X/edbDvIzhU1ABWwIgfKSgz6ma0/9i9PF2m/kktntfotw51+lcMjGbbgE
+NWnuAuNvuU8huLECuU10kjIQgej5xTdnJ9EFQxUZQomzWHoCnuDgwli4lHvGGl5jncSvWksMFSV
3D40xl3w1R7B25/DbytRQYzwo/EucEi9c/5bVPCZJyAS9Xo+BHbbKcjBYtQuAglXqWGxamRiK2uH
t8OXWnKW8/wOgveL2nypRl0AqKRys10HUKAGIQnIv7pNT5uQqzSDygpRbdPsWkGPxM6ZZ5uv7VmG
FA6Awc+S6fhHPPP5GLgLQR0q96bYEypEUji3aK7hvt6x43BoVqYmIKwEugmzcs5X7gcA8NoldsSp
8OKXGUla9dOwg+AbWqux6hv4pnC0/exaPF+cTiEfC/1K6gGLm3DGU8wsf1S0ONmTq5JY2JhR1GLw
9+KKXmYSLRB3K1+2fMTsmx5IOmB5IK/3z1RTRRbnFmv23KVxq6wVk6HcXLhQ6/tGVKo2eWWRDtew
W6iQjv3mUALpAe3D6yc5N6IdXxUYOeStHG4U8Sj3WuJHAc0fbB9FZCAEi/tQN0sNJh7NAAF8dFdr
tfOx1zYUofHNDuZwmDOazpt7FKiyF5oFkJApRqo/CO3jHHkX+BGT0tR4YK4jvkHYz414Z+YJZOxT
EyF/splA0/HDI5q8LKJTcVZGQ401IclA3+S1NSslrlva11uBxrrK8M40PzVR50YH9EU1SJFdZpGI
OYf3br214Fqg+OI+aR1NTyT0X35B+915McJ89JTBBieacaE6BI3qrCy0M57gNBprqX27TqhkLss8
7HjHvZEqOfORC7pK5MNcsCftAx0y6Nql3kg223AgLPzBAVdNulc38UMM29FscpXv2m8YKzdDJMfk
OrBc0qN+4Y4kMQJgF8zAPry0ZjwmcZCjm6YEtoPtZTXu0eCog8Tt0gU+a9SiCfs2EXBSoiUB8Yzf
hp2ByqwJ9PhVZzqTpMFxUKuyIQ2Zf5oKg29OAbLSHy7G7WsV929p58c2QQXdeXkpw6huzuVHpeH7
vETx7axObDWhn+J1ioCgxXpqVBIWrXsrmxBQtl67ULO+lv38R9lrBUS2CBD256NYcjWIX7qSnxMa
NUF7wv1LUXQwTb7Z1jNujZUVkDHqHxywVScgwGOCuhBtN0dZjoI65pTBz0+VrGp0YdeCHWKI8fV2
Cwn2CmXTzjdaMesxhMTBQYH6cVFAZ5XgbBsLROOR65aeOS/bDdD9ea+asfUhWT0rWS1o9Yw1bdg1
pXUhdyT6D7EbCHygW58FvuikMGEh7laDetIjij1ug42PDDGo73955koaakwrxBaErS/16c46LRzd
CV2Br4o/6BRUJ2oZ5shchDU/xaqQdPGbGq+u9QS9W/ybpAUEhV//A7T0k99fwv6BDSYSmiAB3peg
YX05fb5Wex0VWwSRlp6uN3PrVtSUwBmehIOpIoIN/4o5SWMue2xbk7jiC/Flh39e/fWCnyqmSpGg
pDVk+fA66hA69LC21z6ZWEzLwxlAntN4VavppOtH0Sh36VggFlsAteu0OVhR0yFRplQlmXOWBhdN
CqRJSHIRjJ5XIs68SVSTSXIgCeT9vuohjjtEpqaKHWr1CTfniuVgX+56Y3ngQQqsF0qczOUFeryP
poo7jBduwhoxTiN1EfgynZwa58PiY+WoMm/ult3+irlcOQwDx3dQn0AhX0vAhl9zhW9Rh3czroYt
NIysIreGLHpQycUL9amtU4EymN7/PCql/ybmme+4TBleki6L4gBlFRVGYXvwtpwjefAI5lNPt5Xz
vQ0vYCjlVMamaO3o/A5zN8+ogKFTHAN4RgTwAB12rxRJBej1ZKJCp9qHrpDAGrth2NcwqVvv//fh
HOrHWChmba2KE35bbs203ihlQsFKwmEWUBftUZcVtxySkIoEIsKJsL18gj1ZIg3/iHzgEksZXeqq
8grLAC0BtVAsGvEcZh2cnd6r3re8TnaESrQ9OnkV0EJ0WUNbPM+AP1n43t3gPdgvUqK6TBEs109x
TmJL79hQq+l7rPG22kqK7IDrlExnvOvl0+XSfHzFjA57uJZbNyRqEhaHp+9z/I4epQhp6xQ3l74r
+r7JhjpF93EPccBjvHJNew4V+q2IV+jm2XxayRg6+akdDTxjhjzG7r0E2d6onxqKWtUej+uEPjY/
gFG4mkvI3Ddj+Ulkmymwy2TBGw/XzHSPg/cqgNsUT+4eOAmS3iTOFjCItm2oW3+E/XyHCUeAB3CZ
JQcjDUD7RCR95J65pZk/JSZeYuLJO6NiVwgelzXcZ/4ahaSRJLhgioM86BQFFFzHGjwljrPE7UyY
MBM3VdICvEw18c+gg79yWPNM1wCTl8MLNf1Al3zhCgCSC6AOlsTJ+3ZaUr0/xgWFHz5z1XJJLlOm
COSMaCHjA9I4+EdofbTCyPmBu41TvIqIZPhEgMhwXjlSEtQmwrb3KZpX9e6te+R34ATiGybC+FKt
tmOEip/98YgzcZ200475oJUCXowVVhl01TB3dEe++epd/B7OiEAIHQtgCoi7brVKRQgSjAqncMhV
m0/vyfKL4jZXS8fb1dZSny3HQ8iK2mKvd9tv+Nt9fU787hpUE/xZM/p6W9Kdk5fXD9L2Ad9gVsno
QBTxG7fLJuHcbAOvO2xVyyGN98pxJueohRs+VzbkmBYtY+uMJ2O8gkBjN5O9vcVub3vpXyQIuLQu
d3q3TLmXKyO4kikVq87uEJq8AWsOpMIFqWUFJMOo+2C0nTJnjMv5e4UGUumyvyYjLX7cEq/lmIuK
uKW/pr8sGObJbBFIaMQRTeQOzsp8dhPi5ekM9J50xY6ZTf1K6610Xa8/e373tPOcUTfL9bLGm8IT
td69MCLU11SsgmMHB7Kp7ADZmqarISTlm72oS1UVs2mqtJg1w8OzYihv5DGwBaRTJHANo6xzhIdX
F1I6aAgZ/Iu49PXQFQoOMxADEb4ScCpl2um4JoRC0yoZ6XsUfkj/3w/hPP8BakNoQ+e+nGeFe3lU
gI548r+PIyG4r3ris8H0fIwM6gQSJs9ERPMBvwrG1mhwOmApYPbipQQNy0WvOzkNW63drUEovro1
ml5mff4bWQU82FTuHXKVgKbG+98A48nFVEHq1/2GMfq9pa+1WSpzz1i7Z72t2M6lI4nAzauXR2dR
lCYhDAwbQdHdQZp7aCk2WbYMXQx9NlJqduibfTujcUWDooul3ACfsebkpoAl35Ng1mjM68us+5NB
VAqQPcGZATk1wqaFdN/4LBQvIpE5Houv+zcw8lKZqYNWh87iyx82c5fRBHzWzBJiVsqcYnHocuad
7Ear6HTz75BubxOg3BQoP0WVG9blCRg+wj5NBlHgYPJZEh0yH7aBmtHycu5horR1APzf8F1nfTe4
F12sF5q+F2R6S3d/Mf4ILGQFxg6BhrqJOUN5YlZxZyaX8C597f8APquIUF6RuUqjUhaBtbRrJQEl
A6t5KPA8HF/eF7kca82YW3XizvwgUjmJIMRBILlGSUcjREDAtL5Ry5UN1dGOWF9H6Sy+9u7qJW+F
6Uo3+Ty40woUiHJ9nwWX0MCTk1Jemm2og75/cwnZB7DfX8XY0wtsK5wqgV3ghKy4yukJX1VrhPqY
TvBW8elBngwEBswUN5VtRhnR+xYj+52exkmHLljY1n5oh0kh2MhBWgX61cs+iCsPJEGlAqwdrgBX
q9y62fsXBzoSOk6DvjUDMk+93aG58DfvIaXwV6sOnB/Ld340rzWXHwqk4+I86AeGW+IyksNCaDvK
wTDOSrbRuNpczUc2K0hzTAy5mh10lfvCmgME2WnqfOHEsndjyMb4qyYmREhnYUxlCLGN3Cp2iktE
eKSOCJ1r7NOleuDhedgev6tbozqa8kE4/BlJYcsiiwXymzZkpICF/x2CLrjxDCoSmzfgtdnb+6o7
MztGODAVJmLxEGf0qV6WW2PpVfFW54LqGh5AYixr8VyrRBXBr4/E1nPGighNb4MOKoVxhe2966/v
ktx12vRHCOTLFLGpQ4UIQM7xCCzOT3oXQpIa5rw3VNg2Qt6nYUNtCi6fwP7XDBKT0Ae02pljcYL3
cGb1NZfUAzO4RVRQkpqu2w1bRATFZ/kHMzytjvDr9TCURCpv8O6bJuQuhJ8kzwCES3K98eXXy58i
Nrj4KoOBHIBu+A5WoEpZUvm2OH1qcSKjwarTieHUsvu0SknXXaoe1MoT4d27R6Sg/q7n2bhmWhmm
PEfPKHAX/1oG5lXdp7JzgyFtSEYdfY8g5MRJV7+C5A6M1/KILwfmAwBfOhzx9Sedjgz/zBS8E+sP
yADpTG0++G/SQk0Pv/AsuOOy3Ua5LKjJOdL5QPitV4p9FOmdRM8Sme/tf9df5s6lDOmJKVCm/NfD
5EQmGikFkyukcPik6uS6vp56DIRp4wVHSTXmE5BLfV+p1jUyRw968SzOdOxmxp3UjDHoH+6cnX8S
kgeUsi3y0XTz8bXS8ja/0eNrgruvQ89jvMvKCHq91Nvks77MuFPhbAP14quQkHX2vmisI9lCrsn2
PmQ+gQ7AsgDxo1yjtYDeOFGw3HYBZQy4ccLTVapxChnZAduj6pxrkX7lDfqM3s5eoG6jsHghf+nw
Mlys70FFXlRJgAJOyzReAwNj1ZRrVV4Q3lfetR4ZWHKAR58Gd3c1itMDKzwMiOLCRWuTw1xWYqtY
e54GFIpl0sUsPxPw8mLDJMcMwTjWVvElFM3nYMesl6tRwB1fQuSMIKBJY8Qs7DdFUZ9l8V00LGmL
qursCFfQfoRdDRAVXbnBfEhc5J98CJ1ocIPeDZC1X4Rmt4SZoqTfJqf0yW7oJfc1N3thGh0rkGdM
y2/2YUwUMG7bfqbxgzNjKqFc5Y3I1Dre+X5isrEGFViYxswrvqxpL9zU8t1GUbo6sFT8o8+QGLJ/
5oW6Qb+6yQnngqNKYQNPT5s/4JlCyP8dCeLEWRHs0JPU9qMevTvNrwXZ3PpBUfDy2nir6oli6yLy
49Z1OMujEmGlrVdVsIn+sZ0QFQ4rOl7QYyxSmqQHTNdhmZiUdaXvpJqsgL2yt3jxl4/l17V4rJOY
Ud2rQce+CIRBtngPZMrfWE8B8T/qoKFKdBVVTvL5BcYa31GUmoGWlbEq5jFE1GSDdXa8C7diE4LO
oQDrQDDfNxVQNqOxhvuI5d0ZQyuJDtdAKufmtiLtJp7QmD0VPPT6urE1/TgT+kqCmrNo+R8ZXIV3
kVIOedCI57KnRnHw50qGPuamFj1WFdKL78XjlP1F2Z77A2CofnouWjzjl6HIv4K1JBn27vLr6LQ/
vQ0nk5uqcKOcv3dvl16BLrmaYi0BEG9IDSeFH5mzsBZmqlXbs9JGyaPgTtbDTqgrZiyeDDEhBFeP
DJOvb+24daCTvsUrc+6pb2U6kZBqNhxQAuPRd59BBGjy8gu6ylh90CCqwGc0/SpfRfdY125vK6HS
bQGtq3Rg1chmlx2QX3jaIpQGrV0nQcxThqm2I3nL8+f+pom+A39vykDx36cNRnfwTWZi76cK5Mcx
qNizLdr+cZFmVQCsVkusvZqzyjr/ctMoQhcTdxiYjYpjfWK8JDVhDZ6KjKSJjn4I2GwZVCE2xs1B
zyuIgPxxb5O2EhUhnspjCHCcu0uZKIsBxq92VBlll0gVzNzQGBqQ/xkamyV7q/ZqkijhXY0OWYOa
NmN7AnInQa5dQLxWVMXLYd3rHO78fvfVbWlD7ZiqHAm3/yMNgaMzjOFEma9EnflAPvc/3gYb/iZY
8VFoLt0nIgXvsD6HGk2PxBBJU0L597DjHzDWTgL0LQcwbKQ72/ybmHCixvvnYdjhKulbI1nM4wqw
9vaNQeNrW2AYO/pSEtf28VUgDkEQ9f3ZcPAIMpnJqCXOOmqBE81CJvMJoITQizLfYe1OwZ9GP+t/
vDC6OCds4hzOvo9Eiunu2KaAVAwwgQkNnPU6Pk85OeBlR43CwmeSr20qcCUIQF4YXtkDld0KY51V
ByVVz+mtiSKlo1oY+v8ijGBd/RvEUpQh9088tXYLrzXrnuZxkufvQbj4UuMVN9CAlLtiMBpUH2QF
DSWsPDjHJQyOINqdzN/XvfIEzh6ETQbC5JSiRU3T3US0hFnJyZ9QEBd6JbSKcoYVbJJ4j+LF2sLM
q67vQZRI4d3jMmbN9bvMbn9iV4opP8x12bg7KnXZ8Z1TMqk6aBT3gWQxPlSIrqSpbUqjcSLoRGyW
bpseZu6bOPlPRm8zum5NF5LjmYXR5TGJO0e3lwx/+MMdW0TC41TxDmxSeTwrW/4jceeDa3TIUy7f
5AHSHAy8l4u9iq6tFp9GoLOza6BKrbJQWETlvDtSS4q5jx/zw5ZeT8TcC4XVWNCTTTJKkVtfjDmt
x3GK2JwOLWvuJTLXmJS/CPMUo1A/uh5Aoh9pQywr/DoDOf70D6OKm8xT5F4ugNXKg3wIcvgMnnDF
vnJzlQRoOIyqrR6zRfeQ9+25fmSNz4OOaS/FWZAjDp3AmgVQCBQdnOeV3fcVtlKWcoOKSW6RXLq8
MNwqeGbYk7YD0n7aSX6c4MKgnWueiV6ynHTNfVVyUX4R3IAaLE+6MiS+jug8VEJB1sH2DuKoADam
v8ENW+KMykjfnkcls3DomFfN7dsEkSuF1MJ2KNbYcHcNM2KplTPNymMwTTvS7fdKwYpLvNLxt1iD
6GPd+mSDBNYdbF41vc6UZmvJOQ390bbMajblPJkVa6CLHHVCzO2r1NPK+b4xJsVoul6b+xuUQ5P5
uwKJQ1XOBWIUrkE7GkVgDdMlm53Xvv068+fgorjJq8bkGGxYq/SA1uxcihQ72ODnudnMUC2Wk8gI
24+U5HSlIm+V4/Bq5MwI6CxOERt7Y4qS86Bo8dVhTjJLXVG3423zZ2WsMuAxRojEiVJUuVEOaB0B
vSnYOwA5kCTRmF8Z7GQ2GFbg85SbSJ686Hxb1Ta9c/I3zMb8zgiVu8MjWtDFxBHPmpjydwN8IlsL
Jc8+kfzqZ9uu3Wke87kzAWOWXzPxqEgBmYIJ7hwyqVdjPoXRP8mpIbLno9JUZZuAjuX5ywPTGb5Y
q0Uc0PuJbX/E7liP7swmo74k0f3a+r2UVzQaT1wCv99Aq9Jtu0tbWlaMQ/M8jD/l2ZRAHX2DNh1I
9heYZWf8b5v1foW5a2kQO9iVw4J9M3S/ZsvzK6NLwHHmpsgbAi6l/rJRfoM5epILfg3zI4mX/F/R
on6iYRRbgoonp5r8tn8CGCq9mYbSfEO9Y8tP+9Pl7cTQYTYp96o/GVRsYG1ipi015+x1e+SS+5gk
LInYDPULYKVGoru1CUfARwi0BjhX5gBGRdg7/QbseTqhTYt2KaBpwV6vbX3c9GFjaaIhalpLpbAs
M9zeJJ2CbbJldO48jDR1uj2j2JHsiyyYMag97nsVgMdWrRE/Bx8jtESYzCq6BLDvBMTLD5OVamhB
pVACIw1N+nDFCCf6kglWNtFqHfEkOzQik1Tg4K9gSR91ZysWt4eHY+LLjypMZQ/Q1az6R6z2gEJO
ZTjnWqJcUaxDnTVqjXljh3iKIKfzlJh30Gm1TUf6tF3nDNAwEVjvaeEPTKMDPxmHqgrcRqGn7kWQ
FkNgBxt6fqOOH1jk84DwGv3cDhhtWLL9JfwdWakn4TNMqZDrOfycng8TG6wHYvoWaREus9GDJdpu
MveEMUW0AV+dQjr/ZaxBzRflrNNPg+6O5JfsW1FeWmfpbH6sZ2oQy6YhX8lrWKO+p3zUpy9NuocY
cmQrlTVymgk7n5un3hMLMkJ5ASkcxyk7lavspx3/bY3EVTTR3HifrryBR20cfq9w8OOBwy1uC9iI
SJM7uyKLkRvk9lPmeEzuCWkKzgIW/hrJFgY66H5li71Y29hwxuMJCIn6QR3QRcevVr3kU0Uj+Ub7
ObC+JeHQMXwNBv5VUJT9I8AQ50hZKopwTTItjm+1Ab5SIzXugljzI9jfx+GxVGDxanp9zRokByqy
wP8OVleu0awR+44ywQDsKgM1YBcTdyS9HmaFNUWisako5wpxVv4jgHfi+tl8laQJ5kVOb4s5QuTK
UkISNTcdbiwvKXRec1TkCwDI6C8x0DiUy47debUb1HAgbvBmxDbUtcD18wNIglrbwwHxu19GdkAN
hvNy0mxl6b7C5rc0THEHBR7DHcmbV8iM/VSVAfGCvHfql12pj+W4LBgxPd5zhUwuNIM9+sFZGe6s
kaqXZ8TTe9gosWLRmPAuyjpTKZMAqNTZ4oF9eWsZD7hO/gvlgSlMXI08GXSperxG5dq2F2QymYOd
eVF1kLjJt/hxVqFIVYNpRvsJTQs+B2IDS86IQ+MUYLNJa8yIdFxqACepxkvz9d9gpgMYpKDxFxHL
H4wPgC/1JWeeOeTcCIhpaJtvvQTvIxAJG+5i0hvCBT7OsKXP9HJShZG5+LDiLIYxxSuU3ClxD6Dl
KA9t/OTbS7CTH6BVqmJ67bmU3RVQrRcch1bGC3EPvCkSRrk7THWWRoMX/JSVIEPy/AXp82szngAF
3DWwGPrBM5Qncho43RCdos0z5C0XAymRw4r/TESuvwJZotc/q18o8aZpxNax9fd+QlRA1VzBvRIo
tRTMZTWGuP7T+3Il/s2Sp1cEjpP0CDjjleXx2Lqt+x9+ZqqXX0wBvr7HZUtm2bbK0xI+RrLWYV5L
Up0SM0nw4XZkEmd9HxvyZ6YlQOSLIQSFmihIjQaYXPADAztNcRcJ+ZdC+5f3KzIOMw2w98oNM4aJ
D5K36uXG+Or0eHghjw3lg4rIFe0LiViQqKrf8k7jvPT7CDn7IXHAKrucnc3odrdmfQ0c1WYNytc/
ixez9qSkmtfilYdBfjSeBXNDvDip2ICT2IbN9qe61wqh8iQMl9c/4BXGq+IwmBaumlUmG09F/LV7
RhyH0B1zLXvJ02Ek+UmkYhTozbVY2tukcPoQS6EXo6C7wI1oTiDFUPy1xl+c/bQr/vvyc/yBzkDW
VqoW+zgFKPJfNp6DilR9tZEyZamHIICsMRFdYRCSFSSdcgUZgSyvK8GF9OUGf70qUmQvAAFyALLp
1UJ3D4felEQ4xxp9CjN0gjA/HYuj3sNJzHldFQuukxv1YOwJ6nfRhrbj7bXNdUMYLvlIaSldB6/L
12F4j1N2x0kmLYSEVV9emNTWo5vZOsV0xTs7TNm0OJ0CnAGWzRW6zC0YrfLbuEmdbBORenfso0E5
xF7jZjOaa45OP6lAw8ppCyUSOQ5cCiwY1NR5ZWKTf0Rm2Dv3eB50jtPE1kJnbw8SLCuPvVX71ixT
PBdPssYDXJfIUAr7ypf28k/YreuxEXt71e9tomV4CUXiIBXIHgrvZFCASSY2Pi3/QXdAIN6H9tta
wg8qPs+4KWjr8kOjQCyPNN2t4/aEhy+p8MxsFOVt8oTm3xO/Fhfne6q8Z9FAE/MDvWrIFHY4mwXA
oTw/9/PgXk0RIvH6EKD3YM42/3dEosgejlSwFVbXySMG1RdE8DaLo52l2LkJiv03phogOkNYJJRX
QxL77J86NhvUGODsChalQDtDes2byXcZXgz/dsdROjSERBeCvHp08wnWwCxaX0l8AYbN0Ae3xOsG
6ZYCci+h4bd87FxNwpGlzy70GtEWPXL4fVFrGBPzr+IvLh+ImqpjgMHt5tBYReRSAA6rXV42zXnZ
PYL+0fPpVv6l3q3/UVwh5F9h+SWl28sv39tQQQ4D0p792EPzlZzFvjBsJ53RA85Dqqe/JixBIUhT
8eqxAtXZEkxpry/HXaF5huAKSb/hHzy5thOgR+Jly9nroF2SooGTofucFBsNB/pj73j2D10quAki
uvx7AppIKaItAI2yrWeP3XIX4fWFKdMubOD+ALdyGcHHEhaCyGmoyJ39EfK6Ks7zakfjHTU6JN4x
4yqCfqEqmZ0TxHiHokjXaP7ds1SfU/SpyaNmiw1pWFBAut0EF5P1oxoC0w/wnly6H2OMJlGQaGEo
xLfzh+/DXxZ0JM66peFtma9m2oC2EhoSJJQjYSd1iYmcFMPpupp8OIIWP2TvViM5XgrBTXHzoV6B
7x03fGjWbPAQE5IM0w3FSe56LBvrsWGXx0CXkV1lnHKl5OOUrwEfVzAC+z8l1/8PCvGeVQzEcqWE
D+CAqHviFrErOkrNtG78HHMxWNxzVRfgRZyiXFzWbG1q0fc7gtxfMnzqNP1AZRUwXb5DoEuJsOuh
ikROmwFDC7vowikmNwqHGQXgRyyvWzrBVZnBVpruPcodxiOyO/skM3rxdKQ6Hk+9rkYIXqOrzZYr
OP/aNTcib9tjptHYQENNsbbX0pyCG9TgMEFf95jEm2mq8BOOb5vzqfwIe6U36uKRSahQ4JOJn82P
mZVvKZPpGw83hwEZfMPPQTlHRHkZol4F+JU7EYQnXuPCcTxiUD5T14qtO6tT339P1nTXItiumyaq
2B7wqaEGe8PF6fnSDe/L8n5vJFEHNKJiQSqwsZOtGjD7kBshUa/0rOTBMQbZOUNinfjIv5D7DdNU
lhMVHtbNJaV8Rz7qyy2/UfpN+TXGe39DPpzVjbjXd+LCJh3VcO2n5d/1QkEIooIaY7yD3zzawtPe
R6RShptjIU6ZaJ7oGqjWxmVTip/EzCdXJ6je3BCXDc25WV5uRHZjTuKTJGstb2okz+wYG27J0SPk
NUDDNVbrn2pUpGcM6SC2cqwG94Dcwo/9GABF1TLJHdPDHmpklYuB3nTJyjEa9bFw2oHm81ZoyjCp
sjkPy3Z2QukdCJe2lU8TSFj31BeHAiUhlFfs+N7gA48G98G8wL/FDH/NWJL6LJoUYj0GNlgdamjw
6GvAne2Tws8EJhlNVtlbfNa1PZmXpKXBwu2glxRKtPla1wiVzz3WVTeIL30Fb8QpwUNeig42OF4t
WT4is1kC3fHekFdCL8z4ZWVckjpLMd8LYWrNOL8wtvB9pJ6nXdUScIMz2CPHHNUCFJ5GhZW/u7Dr
Hx+cLK2Mp2+cBMqgizHAgYYcR7AgiLmPre3cP8I+zo5+zaEwj4zTRnT/zsOCjJHOvud4l4+ca+36
bdy1iorhrq2GMJJhoBlXX3fponojDD+uoVuAMQiLhDlf33GhFyax0oTUhH/dRxWGIsNvBHWoyG9b
RYundLpA+bevJjLeV429lqR1mz3j59qIz9sXW4yyOrCJ4yemW0+nrQKZT4aZWbp9GNFuxQAs4TKw
cR5GIj8/QrtaPv+oMi3prBgLeEyFYY/DNH5NF/AF1TFKv5yT7hVU2Zp7RtPrk7WR3IHmb0fUhNEF
LWw2cmMx0vp7XtkqiweglaeWviiIpKAbyC7sQUY/Hzq8VoTJrJ3frMb41Vln2n9S+AcXfLJ9LySL
Btv6yFy9XXymn9dBBbAVWy/u/9GQ64wyQSXdlw0rl5pKA9onVMLejE+wLSMTTQgtxr2iWGnOkVeU
Raw00CbRJ0P7T8Y8RYb8lWdgIxXSexz7fvnuMZbsNee7xh08I5HRJa81AmyvJBIbriXuYAu9lNJ7
BYVEyWiwccdgs1iagvL37CF5wTtGYshZoUF5UAa7F8haP8LJKgSUfNBCk1VCEUZaiLbu8rcj1Na7
yZ/6g9Owgo6RZ9VpIbD7uPwZPEFz1WzjwnFRe2brPK86a3jzVt3/up8q0j9vlspjbtqLPnrswyFR
WCGXq4HcVQRDLk8O5r8gyC/RKMgLwrrO4NbSp9Z02ykvdL1XELiJvlwOESCjN6TXyfbWl8JCbkrR
03uqjNY2ghQD+BgonHDxHa6Az3RXcFq+6/Fs60guogdwbC6c5sojImFs0Cnh5mUGdkz3AKIwuT3+
rWEyKng396VPT5D4a6vDfccqflrMjZCsCFFMzoCPUrNGK9Z/xyfc6J0OAHuHXjXvyiBb/622EmPY
pVUMRYBxJl14A8zZM2TRZgbhU00PlHCqGd5m3zWqec+6NtTtKXFBhs0mSYbJQuPGE1PXQ+8DNS86
jiX2e0iL95JwuR2oq/zjXqgYvGo2yszJJtbdav0SbltaHFZxLpFNNHvB03Z2t/cDldozWVVYOKnl
GH7IBxTCaLVDEym+j6I/LzwKOVEEDY06E0O5W/kzHhkDvv03cf68x2vl0r84XoQdY9YaFZx3FrQM
wz8khIPvO35CEbKF0uaYDDdrIwmkCdQODYe7NnGJd8X75cnl9+rh0NtMtm+dmwdrgz5s8t5qRHzF
CEa379xQhW+QgoebnyUD4v/VVEI46dlY1dh6O1mbBwbbX3RJ1GY6rN1zYBl3/6zpRETOQH3lWhT4
sqeEEwYvC+7fWCduRtr29IJLNcDpCdF2M16cR5TNZSfHQ36AwVE7WZIV95+KRARWCKbYrUcRkKVF
fT8zzgyoVaey9NQ0FfpWUn3685bguzUMrfZtNg+nfkDpxVSDI05Ej1vyRgit4J/a81sS8tOkmkZh
walPAVrIcrZpV005evFWk4g5FloLcF25P877wjSiT3uHMDsCm45y/X5Yq/d4wciegdh40bwcRvKI
s03Z5/NXffJHjcQW3kxDezR4WZJhNOA1NY6F2Lzz59iw4V2NogC5IEkPMZ3OjqzHIBJ1+3YFpcXF
AvG09EQA10k2Snjp35uotAC/sJDCK6sEcMoI4Iv/lfKiZxccTKNrfQ1mbqjgD95Pa5YXsOU4ZTRI
9wFN+Zk/O8xc5VIGBWlHp0idUQWs7hMBzJU5kUK5bbK2W7YHYcJMA/NuGNdmIGF7EfmTkfNUqxDr
VVqE9HqvLz/jNwj/18NOQ9EQvMhcq+dmNENU4Kk6hFJbjY7xN+/4PEebrCeKr4vMKocxBT6cdKAx
xMsDgwMIFph3G5aGzKPmiKPlDt6+24TlEQaBVwgo5FdN+QwykcX04n3Sc6WA7gq1xsSqDndGVByl
fzACHlSaO6nwWT+NJnkRizsVGzGJezdYWTscqpaxFBNnYBTvaYq8y/KDW7yjiwirJMTU6zWX0b+f
rpuunjH0G+FmNEXmW2qe+qfwKnIu05QfPhR9yfXjKCPigtvfqHOThd0hxQW3354myKk8gUcoZonV
fvW1c3LmqkUEDGjZ871Eu75/+ir+spPhPsDCjXlG2fJkVlW+zRyrV0XaVIh1dxiiI6THlbn+FigL
wIoIHdVnqUakOzPnL87EFialOuZmsWEvoozeyIGYZo2kTMQKLXlsCUYVwD+JB1ZpmfGG7o+8NCSO
3S2RDymjC/LcupUUA2nldN2tNo5C5sV1XYnvau8qYzRMED1FoSFfdERbA5CtMoEZsWoNecQG26dG
3QAima8mrhpfoLDXzTW0qkyf/wL+9QGhQlu10hPHJU5oG12jHWLFjX+eHI3q271cY3Ii/nH/YlQb
bMPLkuxq8tJE5TOZDnsmQxt1lM2XR9Oiv+Eehng070EFgl9K0LXevPSI6C9CA0hPEn+m5Tebum0V
Egar/btqiDXsTEEOwkV2IKQtaCGnuuA/Tc1Uzdx4LBD5JguSi3MTT4bSvGbsMvL0khZkL8N3tW2q
OagjcFjlneOsqcCWAqJ6XYVMExR3/hr3tua8dssiB1jSnhGd1miWVf96AgK3/H3kOL/ZIF+YNU1D
qR5NWCeKqnX5JcV/vs1c9aEHyiifHBXM82LyALIei/VIRLef9uD2foPg7Z+DN1qB+hrI6T9T1N5y
ccTnXSDzsjGrV2l64n5H8TjjaLxfqIrUx6/ZAb91bahXPTGoaQUNAvORZXBHzsARKs7q7Jv4dCb5
+n86Treq4aRuJeKbbFPwaQxhfcDLtFZPHMn3s9BbVoUYytkr0Q+jRbOCGVWuhtNRs6Rwqs2p9xqL
1FEykW+jDBjK7uY80AscC5QQXQrQsof62StxA4sGLdb442arVxbWAMwlp0b9p++8z62biB8c4+aB
THYtKl1bixGKsNYEdpliTZSm5EXS67jqvtSTt0j7Ozj7XAA2OL2/9hA9GJaVj9tWVNUFDdr9pUtP
eCmMVHen3mN77hwFzH+s9hAD+VjSyFUBbSJaqc7Y0IuWsMN1HQhDu9NBdpq0GRF0DfgaY7N0mwlk
c3OPgv6eWRBKfMRZgcmZk652P69sZYRwupwU0/jylhbWWW3O3dIqqrOmJ2pumsZ9w4hZbgWuVBkO
FENZR1n9icW3Ct7pscFlHhZ2tkV5suQcCE7Lpx6IhvglnIplvZhLgbYfGNJHNH9tT/Odl+P4mjoO
LH9WPosq7yaXhCeVFFKvOqx5BFfKBhyBD892fepsqODdsX30/iDqPsjsIetG1CTtYUBmDlGFl+Aq
JBrEPlHboqDKWCbVFxPDC9p1zb2TyTmK0qWhg35vX+nYq+Xg9/mxainmcRnxVJh3jK1a5rbRnSOU
vDMlafhAEpVbtit8jc4Y0T811Ai7Mj1T8/lZWB/8JEveZIK9HtRV8OUuYZ49fo8zQtjt55WSo58A
+79Jy3JV1QpUBHslcoVnUHB5L74BOqJs9HKkNg14/NiOQrdZqAAV6HrHJdG4Q7EFF7R9rt+GKkAv
IXlDM0qK0SpiIp49fZK4YccwVjOBiMiWrw34IgCFDtnFRINCMm7HYBa69ElF6awLvcAqWVlVZr2C
+AJMXPj970aIWly8k+i8d566jeysT6+BvEOuUC/aomFkMC3pOYDcpGGi7eJlPBRkHdIO9UmVFUeT
nlR+WVF2t3PGaHpu9y5xjT67vxR4fHSWUPIJkSsZcmZ0PSoMEr0X/Uvzzue/xkHEZoXuu9pABQyU
8lmsV4OGqTKtm9Srp3wTHLZylDMSiJmUJQlWETMnOZMLV8lI5we/2mDycubKSfDQdoZNigzZnCi/
NJDCvUzCuma8EAf8ngcPYCf+V5yDRrnpt7Gr487ilHshPKRZA1WqVMouMZKVrdX6t334DGoQ9ZSH
0X+v7BJaB+kEyGso0eTniqzmDTgGzG//Hg/BmYjVr2FXA/CgCW1hNy00gDXe7dhSK9YBM2M8lwHD
AvjP4tSVFAGAuTTaOSDZHtnwX532px4awPHNL/dpbs7pW7keuCpEXJP2r6qLbkMGSjEh6kAd7FtC
LgRm1LNPNxkpThPDLJ4PPUyqQumXyq3oHyFGdNrQw0QF084loB6XaiFIe1FKa6hq21yN+82BbCJ3
4C1/HKWYSsKMFLwdFujkAsOQqxkn/F9nhqR8xO2JXw0uw0tXc9w0OAB/vc8dmZv9zc21+pWx1T1H
tZpx006VgQdv0eYgb1Hff7lwWDO9tpFzOVEz8L8wVtmwwsc4w3TRwum0bJiG4B5cbheRqEhETHOh
gIlIiqBS+GICv51KeKoCLaWDa+tnjQ1q6Zo6wA3F0+IfIDFBwVgdiXN7LoP9jxxh22lVpv0educb
lsA9Zz6upEdgD3KpUGjF7/TwjVSbctw8uv9VG2C6YoCj9U8l+OgEyd7lxUAmaiNvDkoae8HRbn2d
eQD3Whfhic+YrTWolhI6JQB3FFuEX3Is7aps7a8dFuuB2aHc6oqLcjwVtnvE3X4P1tCfDSc37FFz
0YtQWSNx3aqgREsZ6KzPq8puLxNm4VArSo9kpw0LXV8WfBwZxcJlch2GiCsVaTWD6C3DZN6PYsLe
UhlwKahOHlhGRGdYVwJSauEJodK/JrMoa6mfkrcVLBLfUN38a1x60tDriB6KL3Z2VKDe4n4R9UoA
X6KmL0sArLbyDDLIUiQgRCY1BzWqH9AQLfjBx7+gJqWoVyV73leFkFgmalfSEORHthKmlHK1avrb
m6jan+UqVSNpc1rzKiOY2PXLLWIb7wDZ1Q9NMT4yjyaQN4RwJEqRw85SinSYKuq+kcsuERQFjZwf
yY4LmbcLnK6mql/omdNdR+rdsSYMuO+KEMDL1FJhwFy/0Ck9E/ykzbKE3zFdvf8ooOPRQS6Gcn80
1oACTf2XXtSuza0VbK2cX344YgaiBnQiJbr0jJsOO5tB3WwSM+Q6pMpLGHf0dbhAzw7MajhiRqGy
Rd7u8jsftAFiRDMiOdEBcapJaLPptxmJFlEurMw96KZlqj3f8mvwEyZGA9gMcdehppHKTNTftRGl
kn0kD3Cf1p3eNiD5dyW0vNvnU5TpwdtbnwFvY0K4usixJhHKraREluKKj35ft/p9IYkMEZR3ugyk
e3KLyhLq7RW/vM5/ErnkNNz8CzpNzJplk/CjDq1NwxrxQW1c79w4rNwUhwGCvx+yCenOGdEFUU7B
SQQNWN25C0MMCXcgSZ+5D20tDkNbvhcIP0gNGDGo6ODWWBeC+5uYXWpCuhYf7iEbnvgZw9Ca5EHx
kyo07knKpM80kgRwRTb9E1bUcBziibyNd8Q682I1+urkUNUMqXo4t9Ob6m0u4/YSkCxfEokioF0a
rn8Sm4+NovSX9eyG6RAQ3Q/kB6f8Re4vUKmqqsnhTIWO9RVzw0s35Mk57tMhFexE5nlD3TzdS3IB
JuHY/IF3hsx5wof/qM5XnKdt/0on5qk5AoZwYuesr/7ZZVAcc14et78AUFLNKDI1+d4PaUM83a4H
btVUaze4WOPZYxVTBY0dLBO0PJNshJhDVjqUPZicKQfdNWcN/YSVh3XGCdIFZs1hy0iZgOdrcqLM
oXXFDdN83IL3w5btQZ/ItmOXrpZd75vvCOGPl5G8eMCxrfJh5uaLLU3GghIwt6lvhfQrnJiJm3EF
BL1A8KWUvo2GAy0tflduJ5ApV7eXYCp+0zzl/ZZq4K1hRopv8f9ESChdgZRRr2FdcAkVaymla7Di
L4WSyIXh0qwLyq2I8Z5tpHAsDalhxAHSWsxJTZ3el7dudnqkLGo1RGl2QGX34EIolHpZMbO/D92H
Ij4uqyz+v814eX2Bfi1KgZPQgh3Ow+h/QSpdmzYyygT7NiHZVYLlFhFDp8o0qal6M3sV0t3fD8JY
M5RWKzZDFura1xK9IUBBdvZMBZoxGE03HsEMBf7kDXzP6BylroIJEWeqlQ3UGZrjgGgQh4hwECGR
LwjOFkUJeu9YGZOIkqNbwjU+Yp9Hx95XEygqMhIPmriNiUn0ETsbQLxqQ9Hph+inuzrfwHrDUCDT
kU7MdPIP1h45ig3PWj1mgRv2F9dKVQy5A/19fhtW3pOL/9A2Q8Fb0ooalWEuypgyjQC2AfLNxkF9
HbyXRxGuaEkLXZT0RMGL+ylvJ/qqurJohdIPkzAiU/RzmFF0E+qu7l21n5YlwFkssUwJKbf2K3TQ
cAmSHQKTxnJBeTwwz73/wE+VDnbNJhnZo1W++/FrBoGXWYikJj8iVcozM+YfpIc4gvOW7k/Yl5pH
DEMtYiRrLpCd29rJN7Ukw5thcfH4qo+VCMRoIHI7sLoglwusFazWRv74Hy/k8XelnOPs6WYWfyAg
YJlTeSSGZKYDJbgpxOFeuIo5Komtuwu4+qdx7702NEVUYhxVZwWFB3RIC/tQkQ8NBbIYtLDsow9/
SjyxzHmaNWlCULl7VkIcHPQ1u9gtJsrmChhpF/FuAMSpRWEuOSSRTuGMm8s1e6skTy2JiR4+DeFO
dFRGDQRRTnGfH57Vy6O1qSMU+qYDBxyWwOob8fBXwqtJ2+HLZ6BJHLdqHfx4eXByl7dFKJNyHGh7
VbVqQYQY27xuxhW/RP19qkjTLsVXAGhqGP/NqMylJOOzOAVyoq12m67ga4csoYfWz2eiwQ5VuIaJ
1vxNZp+j8/3hKqk7IVSIPi1R+MHQG4K/lz+Hdbqs5OVWPu5YGeHkIVkVHxea+v7U4sm63NxJrHjp
Xyncnqdu1n2TkUQpRpW/u94Spl222717gfZ+ry8+rxcuU4xCQx0WbqRXIQ+2/3jmhMaSZ7vQWotA
qR/KPERuAIqthZSyxXLpAxsaKS4vfWTD1VJeQr09yLWrvuDRxTweWmJuBQ5w3mACscZa95colx6a
4Yjc8pqPSP2h/UwhrgP4E0qUthjjE6awIXYUcuahFt4LCuAZNzdHRIZxvv0qcq2aK10cUXa3otFN
N3ipFE8qAAwXD7ZAubItkRIiRWTTFEdARyEuAIRJ3lwgGc+aR1T7QuaKsZf2xNY9FMHK7XfAYD+2
F0KMQNzu39nW+Nx1aA==
`protect end_protected
