��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$Rx�y�<��wA�*;�x���@�̦�W�X�fa�M-$u����n~�%���P�$��W��kYَ���P7�?UMfT��q�6�U��k�>����~�\N�(�����X�e���/6U|)�X2pF�]$h���d.���9E�	�IN�f"�\��e�z�y�b�����Oo2�?�qˁ'�͜k-�K�P|����y:����3�l�d���bl��ˢ_�d���kx�rq�mh�MذM�`aS�.�DW�mS�9���Y��+�>��!��!�T�uOB���,��\L�7m�O��W���6����'���j)n_�I����2:��$�K�2�Sʫ��l ��!���{�l����.�j4�	��很�̢=�����N��s���s5���_�R�>����ТP .W;������	�"�מԫ�����]�#7@O+?�⡾�Ԫ���e�O�\A�	�ͼ���ƹ�d�	@�nQ˰��E؁Bf���|D_�%au�-�'���w�*%��"AM$w�*V�[S�Q<1�Ɔ9Fz��>cTt���Y�2�)_�D��#�V�,kN.�Tq�_CZk ��AA������a����8P�|�����,o�9ܗ.��`8��ݾ��0�)@W��`�1H��MJ��$�H��hPa��_��"��x�8'٥�gK����j��&m�+���8x��8ic-n����[� |���Ar�͑h� AmȅE@��:�:� :+��嶶�I�uPh{�A%�»����Ϸ	uof!�9۸uQ���1{D�
+��`;C��F�� Ҁ�É���E����B 
�{��k�i?��%���EU����};�&8��j��nUja��`�h��f���=q���MUJe��[ti���&��GI�"�������h��$�����$�p��-�b�n� 	חj5~�؟���1Q�7R�?qk�B�x�*��R~-���O�����E�G8ܾnb�#��^3���@[M+q�s�K�%M?�ʶ5*#�.��V�%�����L�;�-�}s߄e�I%g#�0=�i�G:��e�\��ח�����e�
hE�^�k��?�+�K~N��J?�����3�;�㈄m��k�0��P��0�߿��,���kSI?���;�}��R���P�Ց�����0DB��;�KbL�omS>O;|=v&����[��l���É�Nws&��F��[��R�������ftc�� ��.Wn���>T����7-�f��RUJr,�m0�6�ܷ7,��}����.auNTbÛv~��T&3��D�STCP�yk�d��YJV��*���;� ^�O�W�c䈵�,�8�_�΢[���yt♎	�Z�Ӗ.=#����de��Ʌ���K7��Ҧ5&k2���ޗ�{�?��=�_	��uu����f��p�E�k��#�\ڟɰ���nΧ1~�ϝ��L=صXVy�Pg+�@�	���_�� ٕ}i�f�Ļ9�bg5Ό-�-����xb��ջ�[Vӂ"]� @4������B$7�S���!~���t�-7S���r�g1t�5�|D�nH��q��P�k�U|E o ��y�>L����I?�hIvW 63��^#I�v�웶��H�_�"�`��Ur����!7
X�S�&�M��Q�a�{4 �g�ӵ�4FuΗ�q&uɰ}��qJ;|u��� �k������&�G9Gr<�ǒ�M��;bkaP�A6r3�J�k	#zW��R�e��W���o�&�~}��N-GB�eJ��~�����k�>����1�gV_�K{Ro�2�>�YPM^6�>�'t}K\	V��1�N�����l�W��M�k�.��'���9��S7"8����!��q-���\˫��� ���zU\u/| ���I��V������K@e���:^�ҋɅ_��?�bp�{����@�Cv��l(�xz>��W  a䠾h�i��Mu�	xW�bu�R%����P���W�"U��#�ɾO�~�0�(��K�Q�҆{��θ�#.ن�,56��;�]���t�A�Z������[Y�?�`�E<D=>��@�N<"�J ��l{1�!�R�����%�,�q��#�f�4Ee������q�����MD��^M�����F$툑�^�|my���<��#0#�MB�˅�J9b�A.2F�c�0f�e��%���mad�>�X�*���HQR����Z�`�3g��|*��&��'��$|zb.��j�n'�r]�;g�t�|[��y�߉f<<�{k^>�"+3
�DU^�lĲ�����&�v5��ݝ���U��*�����jT*똕ZM�~�S�&n�]Ar=#'b�G�<b˯���W8�23�HM>9�3�0�xϖ�<p��M�X��T�?�}ݪBF#�C�YA[F���-«!}���6f@�᱑`�Ug��~�)�\�Txnuz1eD�� {���i�4�g!�d��K�.	`f�c�a#�(���{��a�ԋ�pS�5':]��� 0�8��*���lLvosGiy������Vf�h���H�}s +�D�w��ʴ��B_:)�Y���QR�N����R��7J^^����n'P���)�X�NҴ� ;��S\�DhNlŸ�g�ChR%/� D]ޢ>�b�x��7d�v�~�[(����zi�Xg+\�l����c��Fئ��GI���̦N�f��7�=�ϲɼ��RC;��l>4���I\>���c���w�'�Y�4�-~�#�1p�6ת���X	��ܶ��Ы/���t���,qx���階���7�L&�w��,��?�X
p��~�Q����y�俘�)��ʶS'ۙ��ët/*;3���3����_���P�-J�̽{r�|�O�h�.�n�&�������ݽ%ԓ5�� �C��6���f�ڽ�seo�#�Ve�^Y���>�S��q5�pJ=�0~��$lC==Oy��8�I:4�I��7��s�����in�T��Gi��KyI���8��q|��bw�����v��'��:�Ό��3�#>�A>D[�Vq�X��'�Z�b��y	6�|��[*Gg��Qm���zR�k�"=���a���^^<6+�����l��/�Ѹ#^Iᙡ���� �Eu��d�>)�4�ԡ�b��>:�-'�Y�5�ϲ�9��j4"�Mkۊ��@(����#/�����⾷x��������V���8��1S� :rx�m�D�+���Ou�wHF[�?���}��[���K�20Ua<64P��P�+s�,,z�~|$�r��q�M&�������$𼵳]��_�k���P��]�����ώ�W�V���1����&Yerω%��l^��[�f�Y�tK	��VK��Ȼ��.d�3�Uo�/�r�v�@@Β@NN�S��*�Ao�p���S�<P��E_��QwЊN�aϖ5�_�s������e6�ڰ���R}Eg�"�\_G���G��-���[��i�P`�pF��Įޚ�)��0o5� <n�\f�i����E��}��o��ڧN�Ժs�R[�%Pc3'<��i���W;��e�jz|�J�\������f�oqj������ൿ�$����#p[�gp�� �X�&��[7��r��݋l��kB �"��;)�S]�+ΥE�M/t+�b8!���X��&l�9�R�W�\B_��X�о��WX}V�"n��=LU�x�y��~<���&��e5�WfMҠoJ.�P�V{)�H���s>�������T����ar�}=̓'����!O�L9�sA��ic�O_	(��K��������ӧOcd�b��y�˥�$@i�ЌR���ǆu4&z�NY+Vջ�L(L?��rۭ6N'
�
)�e�}�g$BQ��&�ܐ�{�H�.��{������x�	�R}�OR�����;\���� �!���\tDRO���_��Sg�k�^>U����u�	��d��A�8Z�E���V*9M�]���&����S���>J���#A�����A�<���T�*L���(!�ߙ�t���x���|Ƌ�o�� ���_���	Ra��}�[��24����E������6�yx�A:_�KJJ�,5�0n+8�.>35.,�ERV�\�o)��r��R�B
�?KF����GC��(�Y�i�w�J��l�Q/�E:� ӳ{"V�]7h�83)67�h(K��"��}��n�s�vp�i	��Uw~��{	��W�oZ�fd����ǉ�z�h�*}+��;
c��2L\��J%�\���?Mc��ٽ��L[�<��S��C��īn��ʳ|)�vῑVߩC�8s_�[y���/Wf\Zӱez����t�[��5����XL����]Lil��j\q)C�)]����#�ܯ��S��� �>���lxAce�� R�,nE'��C��=�2+�+r�S�O�-͊�ǘ3g#�g��ផm7�8<�2��z(�xBL�(8���ƈ�Ί�ťV��_P�O��_�CYO�Ih)6�I���_�8��ʕ�{��$ϝ�9�����*�:�g#�b)�Ǆ��w�b�7j
��.@S�M;r�j�pyr�Bh�a`�\�g��7m�b42\�ԐX��O��(��� e;`z�G"����'�E�X��4fb��������IN�4��t��|VQ�}Ò�J�!�wxHTZD}�o�%�C��A�p�!H�V�Lq���j����<Z��Tif���Ҭ����0F��cGI�s$� �k��x���)~gsӐifBNѵ?� ���HfbY3��<�JRi��++��#(�������A��M�"9��>("1�Q�Qן��n�~���v�*Q6<�A]����U��ɟ��Q$7}�,�I#3��^�'�'�=]��4�zӡ7ļr�A-5�6��Ci$Q��չ�QDc�5}��F^*(��}!��z&�5�"A���]Mb�����+�^�+oLƶ֭�Ή'������2e�v�?8���ٽx�܀j�Gc:,�?s�N��`)0��N�b?��J�Ʊ�&�Y��\��-�$}�<�#d��B�������F���~��ڰ�"x�'mt��lI3F�r#I�NN\�7|�b
�C;���fd?����&��{�t����K9sz���Q�{gx�퍶]��3���dx.Lnb�/�Pf���x�ޒ'4�}܎P���aP�FȊ��ޔȌ�@y���콚��Fz�����#�q���Q�s��*�k��{e{<wgz���i��Q�jF��[�H�!��M�E���Cf�� {�6$<��n�ϵ#����g�1t�]�x$�)w/�ܤ��_���Fz�x�Lgc��⭌�L���OLb���~���q^�M���10VMf �K.�|��˾UҲѡN>h���W�Q�a��՟Υ����i��rW{���<�W����#�x<�Β��#���+�hF	��M�Q1v��&	�"y��Z�\����hŢ����H��=���o_�GGR�%#�%:�����n���=F��)�8�ȓ����1�7���]�?��'y���Ŷ��zRAq�q�k�T%��a�ˊi�(���0�hw�J���y��{[�*R��z�T6NH�+{oa�����S[��`��<�,�!٠��gܪ�������ņQax����v,���� U����A�e��'���3�=y2��y���^4�v:��g���f� ���F�8�F�Dd� �<�,��Y�EV�k�2�e��}1�.�}�"w?Q�m�����3)�1΀q��k:�s��i;��94�,�VY{~��<�mG��M�I�ٛ�Q-GJ?5w�r)���jS��]�y�"f��u�`" ������m>�i|Tr�-�1��\� ��v�/S�˙�"�gZ+9�C<n�k�[TN�{��2W��=-��\�Х��	M�O"x*ȢK����#��g���m�/S`���ꙣk��ʞ�G�Lٯ�A7w#�b�W�_:�,�I�p��B��P�Y�;�z�c^Boq��b\D�&�W�W�2 �4���w�>}��E2��i�uC\�9N/Jb���(z̓Q��q�]�y�b�Nb�~�j����.\a�ͬRr�1Вq����IxO���;X�02�L�Dta���b�	)�0����"���[�pM�m:3�����U�RBL�{�k�9�G귅�d�R[���=���c5#,����JT�zi<r0v���Q,3��޲��������x<l��131��M���*����,����[���=�CՕ��9 ���x�K����8��U t��5�4e��<A��B���Z+�?�_�*OSؼ�9\cL��s�aHxJԪ���7��$;o���ԝ@�~[��8̩b��gsȨCr�6���m3<b�����~��#[�6�1���c���d���听�:�vcxeL�jm�~ɉ��n��%�p}h&��b(J��~K(��v�'	% ������!�9Z��FH�����hz�p�sĒ��0Al�$R*g�w�U�E��