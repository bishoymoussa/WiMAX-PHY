-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
p/22kqq6F5/qHi14IPZlrq0ba4xqR8QGK77W+wPlgSP9YmgPe9ppNjb3BC8mpPZMGXwNe5ixww2x
Gr2ErF/c4EK1WNxtN+Pm7lAErOQY4odOE5nG25gGlxDkzZRMfPXg3M/oGBBGVNzb1tI9IiTSzr24
/+FEB85ZvwLrLqXEu5C0udjtefQmLU8lUYy2vblyzOWpTqy6QqWh1BrAKFLhlGcZpKQT+hJN3QLq
WoK9pSbfT7XTXASi/7f55xbZ5xHW/t5p1X0D5e6E0RxBrX0W4tUUhOBqlrHHkX4dzxPXNj6OVN1k
w3oF+ntLb3p6ZdkkqP5T/Js+UoRtGbo4YrGn1w==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 25136)
`protect data_block
Rc2JBDIwzP6L/iC2fmqKAKHfLalkbR+0pI2V6K0zGOu/P3WxSm0a/Mq955d7+YTTiy333THQOiCU
EZHkYSXFW3utuTSmgAfkHzz0aBIcf+Wh9A/LjedFcC3TigyXD4wk7eC2eoha7CnjdELlz86PRbns
p76dzY3wFlgfub5NDLEmrSuCI2fVGn/MdJyURQMmNA740Y+SASWh/iMD78kTu/csLp5ijyAKOeIS
iCzAodaeIvfBtUHd/hJdgkHewTrXH29OvcqXVvLUAQh865nRuuGJHq6XBQJ1KGfAqxLeYxH0Yk/v
xkPD2gWf3mOfvNUmhFqRPO3pNp+YXN72NqzjCMDgXdDFCKP5qsNIqAfB3Ujh3MLaoi1QVw7Gg8dr
y/SPmTT236P+Ryd1MkaQ8pq/hSusUvp08vpkvYkiiu/QKiOk4R1ldHZV6IGy2KR4BoK5Eup7x/Yp
nMFK44lVBBKkRh6VhYahJBJkBot+KzLiSelyLb8gbcYpEp6728QQiQi9DYPboy3mCozabhSAHhHY
yXg7UsRFZ9ocJMQwEF3ThgojBLNyAchXj/6tYZ9dC6fTgO1q9dqzU3P4nRrU4be0acmnwPe1cj/8
mCXSCnw+27EEO45GPUSUp8Vt2v1QNkV+acRUkh9RwZC2DpKz9EDji3MB2mG0Nfkqh54WQa2huAGf
XjQ7a9gVI+kUgmzptBecOwQdykXv2rQVrwuKbKCvJE4zIrc1vxpdRKu47KWGE5sVg1bNfMcMoJdc
vEMubZuKbuPIuwfZxFBb88rlm1xLtNWwmwo1r6EXI8+4GmWN4Z0zn7r7aLChP1lsC5Nis288NdPA
ElpvQzMfz1IYw4BdDSx3TntDrFFI8NI9W0XcxhsZ22y4Zwkrn97g4JEjBQf9xN1SZ7C5JAn26wBE
cJHRjdj8VBBRsPN1kDNk17nyrT0bJhCitYZBBILst6qVQRl2pmXl9lGyIc6CwkFe7IYNf0a7YhNE
PnuQwENsRxLZ7m94/XHIGvX0SEHQflmK3xk+aVHl7JNYObjQMh/Bd+j/kmoXPsu80OWMmneHBQWR
JcF7fNO3cqQdkNKYNUlW1ZjYbiEIpflRCoXjWUM4Z3s5pjBRF/EH6Q0JOgVRy0TIWYm5TW9Fq9OM
gF1ljc2+vpk/nXbLkxMyeWzDThAqXHez007qy5NAA0Uxm797lzMRIF9eYwDPliGJN6D4gab5+/d3
S71H00uNJJ+xQKNaIxIciaCHteUGeXxqDYzMftly/VtWMXhGXCuo8ug4Mct5cTmgWH/L5ZQEVVI1
ZKvKgRJISNy2dzz42PZypB2gF1KP0NvEqHZmp5pO+MukobtB7i/QeFQn4qrTL1ZhLfpNOsXJp6ni
y8oLcJO7TUvhx/RX00kJ+YI6lEM3y6fys5tKykpZuUJ1clpfrqbZc6oR/5ztokshUaANHmvzl4vO
PzLyJow0pOVqVs557pIe6Kg1dR7qHqAY3fAHi9eSbpcM/9eCnVrbvPigXLQwukdXrRWz5mF8l8Ns
MdI/58fVCqlpARm5wREK5CsIQI/W3YI8n7m9gxcvKi7zNwRaclzL0nfkK7L0bPSyiuTJhRMwA/8f
rFr1LolKDOzlKXnP/Rj7Y2KYtd+ci0SNTqaN7EfuJdaLES1CjPKoyTdT6aq15DK7oSHTtl6J/puu
1uwdpuyPm0UQMVfsLFs9ZoslsBZl0qagD6Q+wPYyIx880SrQYOI3XPvJ3w5iwTUAVwrB/XxH5FSD
Ze6Uzo9tPpYnK1mFSBjx8lLE0Ybqxrd+Q+1F9iS4a1/hV98l5/S7BFGpzRCb2K6oXE7LAm5D9qiH
MPWaVZV1oZrsegOTZznRp0iIYF4tuTFamzLovAPZDVHX3wD7AZEpEPyfllC1NOzy02693Luy/Z7V
6uU0ybUGmAolEP22dqlG+N1xpugQ3NFdsW8Xa2H4tGyXBc9gb0qIgW2+MTtYo+TX4Sb3xKPQK/57
3mu3ao8nIgnnm+XRdkrdppD/q8YBRBDt3lFthH1ajLiZ+X7HTcTWQBiATM7uxcOZfXg7nt2Ib9Pc
o4yLIqbwRdMP06IKM4ipiToTQ0hEw5J64PSGVXpSi4gXdgsptA++ko0ABZX5SpYeiUU7aB9EBV8a
C1Dc3pBqQKF9VMMN2OLRCO5mUALovN2aUYET7R7nMb9Dl6RGjLvXgxR05d+Cs14P53sYXpce1X4M
w8upXtxsbLhYfO9CyUfg0Tx25R5D5XAIMIPAKQSl9IopcR0xc4oi0FChrHGYUKCTF65FQk4qqlVW
fdvgERRouKZeIqrUh/1k7I0llN6j/0x6zV3GEjW1RYprYe+HitQxRkMVcAuKyokQudcFwnmrxXtm
2/jhIJVai5aDPBF4+BT7mz8aKh/dU1ct6g19LTV+AJCubRaNA2sch+/MA4NJDr46d0tIaCDfAkZ/
gsZRgywaMadHWrCJCXv+5YFjYL7LGjBcpfFuqNMcwqN051uulcAbRtbdbupO89BWYsXEeam/OBfq
OhvJl+NfXihK+nCv1BSgoGALRidmGweQOVifFuZTMmAuEoFiKU2YILtQp3AcFVJ0HtypezICVsWM
lQF+ARqumWJNyvt1+olK0bptQsgG/QZCHQikBGe3zdfJ3oh96YbycEDoM5EI97WK+il6XmezfJX5
SbiYXRZD7tYpWPpTUFUMWtbuFpWe+mp/w9maKH6EgoJ1UEmOgoN9tfp8v1/+hidlHtKLTq/1InQs
BxMTNAnE+ppSgoz214UWfoVH0A9bDGrJJoXuq8it64Bzsg4q3BVL9wKk3YYrjbfno2Y5GWtGhRfn
iqzrXIQqASkNpYbOlB2NwxVk4+Lt9ub42rk/NxwUOtQgqYocvdKc5n9wKiiPUfTAma11Yvbbo7+Q
bLEwO2XnzCl4kCP0kHJ6Kr3lf+WnRF8t+LmjOioGdQpTyRYsu5On9SjUBxTmXeN8cAIFhzRng909
5ofoaraScz59pv7rzdYcrwKTSFBaeCgKQQwD6L5GdI2hPxEJB6S0Dwsa4erMimfxlzoId69sr0i+
ocxztmUJzFeRfODyvvg9pgOPebt3GhPS22t+B3dX/NONqqqHFITtEkWmI3QlprXR2HXq2xa53wDo
ZFM9UibVid/OZddZ9g3H4KHfefuRKvB6KnHotvXGR2Qmdds/a4xn+sZrQvRMMtpNVWw2J1T34llX
AtFySNyxIrsIquddEOtohW8UHEA39EAi/Dkd2SwI6oElhKHMWjDQJmWEkfn5wraD3EhuJF2jS5b6
65DVGrawD5OVhvDk5EJpWIwAT2XfdFQ7z+Q5UttthenFG0J5MkxXqalMrVXbieGkkTFenAMi22Lc
P0tcwZTtdf7T4cBMCz6K8Xj4MWRxIAb6+6PBQHBkudA57N3CiOlzLZrcTZQgMlvT0hGKeOhNO2yS
3a5QIJbMvLCQcAY/okg3liqj3MgKxapFjEgXTU6lvM2WCOOwwNOkUooWLCtGeSnEyC8WHZEz+14o
JaoJ7T5le56Mc/sj8y2oE8Kd2xj7cUIPoCGRjpvbKlwAb5A4/vF/hurxItjNM9cWcyb2Q+zrDYrm
jz6TWlb8R/heuRU/FiM9j7cZTBGEepAwK5lm5CFCdTWAIK0qeCzof5nNtcSClDbEX1fFH4HmI11/
xDDUCON6r4JhM7LenuuzvinNP3LA3CO2b93fEzmRPlq8H2TF5HQQvYfVUsuz5enEUx93zzOtaNNZ
5OS/u94gq+CpxjtfO8gJ66OCyQJh7RZBFZRLTjPKEWw30CAgalNMBHoCRbKA6mb2tbHexZArsjbh
sn2IBnkCVBBCRf8A924UA0XrEwXSGolpqP9t8p9mLZGWlk9ioH2PlzSSLu+BRoM0BIYIPkP9wTSY
RaTotjVXufH0g5ZCJvjLQIQd6VwYCLhTdUlNdCsASIkrbhYquWlHFjEtyxKgIRUw4kGb/oQqVd0C
uG7i4F0Y+RNQSEHtG2S5hA4oiL4/U/V4Gu4sh4khTM1i2xQwG0Q7IZKEIxN3z9UGyHXvHb1x57+s
yQDK9O7PvToUB+DkkX5XUGy97sbFVHZItIOaCTTEqJNy+nAXQU8rVRjvQcXdxV4QkRyPwb+f3JAL
6ondL37RBAHHhlUrF6uTjHGT6IWE58Un8uWEUXp09DsH5urUybktFtLYnx2RWNwBCb5FX+5FUObE
riPdvo4bK7tlPgvvU+9lBrdqwGZOPCBxbOpeZEz5uIAPGN9JUJ7g7dB8kVOyMvF4jQZXoATjh9o0
1Pq0nll7UKK43uxdincmecnRGWat8dRErfOHQw6x2GTmbcq0ePLZUac0+4ffL3/udV+Rw8VUK7EG
qZ1+Rz5YjjWcgGeD8KS5H8sfXNmfGtj9uDLXQwtTz3Rk/fXV33U4QFF/bASO0tFiMCQuBiqGzZ5E
KfrFy6E9I5/zXsBaeV8gCP4BBFSeDIJsAu7z2SEiZlDm5sSnNUub1E90LPOV4M1BuHpKW8ZRoYQE
wPbI/xNmrKSppYONyUkLSJSOKJuHZDygFJizXjJby2KQBuUbH4Aonhsx03enxmZ6CduZoMAqhS7e
UDqkpvFuT3c4vOB9ULqGoMu9qFkECHpUyZBGR/7uoovqSqohr8fFY9AIrNaOOGFHZSiU6EhBiRme
SdlwLedWnF+qzKy3B+mLHRnKrDqd/hjq5mNB4eVnv0Yy02suX3pITnnuQvd4+cKWXKD9qbJLHK5j
qC75rOH21WMGGYn8fO1MOEQsU7UR8GW0jL3fqOf9BG94Uck83ar02bXBSCb2JebdzFa+LyBIX7K8
s8oxJhzBddRcaci3Lb+tIh7JEF9tCqw6N2e1G4ezqT/VNkaWhH4eSant31Aq7V8ZQORtb1SegxMF
Tdkac7JJmPGwrQo5Fxqi3AZuiylza9nb4n8vdrxXIi3Q1+tY6yKdTK/4qeXjXGrOn/C8EyrvRa5T
xHa7kWYd2nIE0PI7xWWywI0ROg/t5486O3ZRHZrP8GWArRC2gFVU4BWpO7LqKV27y4lV7v9NUm4p
d5KaC04aiZPToKR1Oymh64JwDb57aWdcvHc/8cYB+OEg0NVkcc+OeSLiTPm9sDutjgYgroerOhng
MfTNp/oLMteCtWYS15f0Dc3BVDeyfjffFS3gCkZpYip1TNXrum2HxKfeO7BerxTDLYmzvYbtn7/H
nwcld9lxlkzI5fN8XukMY1N5UX12uDMk38rJHhirzYfbQARkyjF3j10zt7WoK5g0s53e6AwiFDjb
0huH3xmGsIynTzrvENU4ZmTNjlgExbxYnSc4K1DqaUwXI2/AUhqIAgH7ZNyv5HbU4GWDgv6eKjS7
4EulkykExzmzTTYQ0gwpQKWtgoi3jNKaU9u9spX5GvSrBMWelh90yO07RIhQ0ntEP72TY/lujQrP
j71Y9G3fRYzD+zLixE1vC14/FLFbihqiUl3P80Obk5bb6TmCiASz+XO6DecuYOJVkOQrK7Hsv9p0
EKDexQtejowWZm2Z4wq+SlYu0ZK2LAUtJv8Tt8048LF6RUQ0Br9YqV4Vx743oxWy+2+p3ZggtwGi
LtGxmcUpmGv0wJlbxMXjMujtezIrUHPrhSEANSYLDWXQ31phvqDQ3NihE+1inlVjPi3KTWo4ikSf
4ppQcjBP9vGFzDv7+EQL+uLUjxglfhytgLhtew8zJ8fv8vMKauNHYNdsf2iEUfL+0bmjvKlRQ2Mu
gtDjYe+KTdHwQCdVlQ7Ekr9sBBS2KiHj8rs+eGyCXshzywK8b40W0875/UxdrUnDEg2b9ATo6q/J
gpuqAYfxY54bCsyq+Spii9dLaaxPuWickwJ2XZS7zPaKYruNEhdjtem/vZ44SD8r1yzLWwr87vp0
y7i86mM4n5As0iuPKD4l4e9voCOk7C93q2C1yW5fLgwoz6oU4hWth3CIwiRJ8wbw49haRf6+UQAa
iPxNCUD3EXxFLiY14kYnIOKkrOx9f7K991ztS6y9/gRS3tSvJZ4/wYKx5d4f3CJiPzneKRDqZweg
mOlKAWAbFjFEClYExKxTEmo2qZawwV79OlVcnsbzHXX8ONF/IhiAmnrwTYZgaMUgiyTZ5/Il7cSv
rAXLdAVj9lGFj9dQHDrohnEznRCC4flBBuYsAOfGNguETqAgPvxI27I/0BEksrKurKX0xNcKuSLw
ONGheOdNfdYSDyaECyiKUDJmtAB0ndoM2N1TcAF3GHHows7EgFhuCeG9Ji21MZMvPnfXEwbHbJq7
lTTdI2LgK6xSajFKZVImwYDvnW8gkP8ft6FftGn+SQmSBeFzqz7W21j/hXe+v3Nx3xC0RYQv3Unq
5kxdJF1ND6r+mPaxx2K7ckvNTWy+RhtTDpf5aQ3EOceZV/FdhKPivvbK4AZ86rk3qirxDPuIjRfU
ICwu40BMXwiWzYFjk9T4Q1g+dQb9RLlhOUGkpCoPGOGDLInjTCCYEKISGk1odLPcWdwYJFdT/ha+
ZJBpbrVGTr2bfuCyBR+20bv+D/r8KLgl+2HjDPVqbPpwjDKlJe1NLZfBctNRcwDivatiXbSZkFTy
a4f4mchKDUd8Vn8N2TWjDQPxCZYw4152B5kSSJmW+C++Q1PYaXH3LohFA1NfDn9soYgsJs6MFvfK
RG18kShorcdaG4jsHHjSUn7GTxO1d6TfQMVXwiLZT7DF2NgRpOuk3BLh7dXMniy5HfYJyIJKaxyH
V68gbtHDfke0hq1PA6ohJXiappmLPjcdjeAt39mj0ImtPK3vLrLOBP8bcsRl201bRBSyu55HlWpd
MQG0+kNZNUZ1tMn0y5xOAdWBdW4R6pmq6/QxtCdIJh2c7RaAzC9tTtbQco8ELmKBs/8qFwGvrnCB
pqCGMx6jw6NIuW2IAIs9jHpgzp5k2rheclk71kBVYmIxZU8/gutohRlxZ01DnCWSv7MvTgeYBWzl
tcxslgXWjsECtvaejTxAmt5vLsdY5E8acedCJtqwUxPj0gFNob6zC+Yzw9SWOxnyF+xX8TpNGEWy
Kz4fRI9VSBlQnj4tHT16q2lSnssWVEhWjmzDCN5dDDOFS82u/bYqbnhdH/gYs7a8kwyx3/XuTUgr
w4aM+Lrt5dWNQMj+M/GZm9hxyU8m01oWl0uxOcLP61OJ5cI/WLOGcPKoACQll7KXlHqblmMxN2Rd
VGw28bNh05uITOSkLcokFnQDX7bZd3Q+wHmmSjokD4ua5q4Em1WLnJWIUYsAJ6aceBQgx//JwA5g
SbtrYZQ6zfA70Y8WMm56PV1BspkvIe01DCNLI/IQWJdjuAyuKWcL06cj8trS0k6Ar/Vpu9X4FbOV
58AoRy7VOn8CE6AnN09cIyN95aBnAWI4Zjch1zxI5b50QsFkGU1R1F/IzGtLviCKuHuoeaVKtnlr
QtSTlLCRhxWmK2lDGrvO5ZfRMuWJ/pDvPWuI/BwW0KkvC884KDJHa5wU8Vj5Q4MKNCMh0HVrwyAM
DZ42+kTCMXQkkxOL+rtR3GKwIbTpnVpSMP0adF3t4DaQvyE7QEwwghWBqXVM14TetFyqxm7RK4M1
k4PSvawQldpnp8osTSUAEpBdc9g8kPCMf2Z3niCAy9398ZoTLP7g3BKsPhKSUIKvmWwTUKD2xiLE
VEzbHhVIgcH1tTgievCx2aCgMBWUPL3YogP+ke6slrpz5EMKhyfC8K6GlO/R1FymvulxJXIvRcu1
lCelyabAldEX0tnA4TB9o6k3DZrKhVPomccJuI4yRDTF04YGxdetFn2eFZV8DUdVprnOgXyE77vD
ZsXQZUlOIU+NcrGXDzLa8vOdipmoRnT1OYyNu+DXNSJ5mYYdLK40kvBESyxz112ysODzIGo7kJWP
TEXc2/LwFajvkcCbBeZqZkVpdrVOnCneTnAQ/AZzabrYujgzIZft84eEw5DVbboxhzuG6VjWRJ6z
K+SM2gjdZooWORseP8mfxpWtnj2LRnypRmOuk7PKBJiaFVzT3YXMf5f5brnYedUqTazRbre0zNTj
7QASbxLTLaSWgL0GnJ5sJi1L9BhQEGBsC33R4O/0zKkx+Xbkcu2fpEAW6/jKiLJsIcyBDj5Dk22r
bxFVuCxXf0DF4twpSwIYdfj2x/kiOEXvsuH2PBATBv/jajsQxylEzAGkRbO5+PjowCV0C9krY3NC
GBsnit3zFKnzNFdE0w88LoqA3XjQJ5YbzqLkoOLSxuolHMcaAu23Vc5bxCNAFh+SeoJxBS4W9AI1
sS4bnqOHoPRtdirV4BF0tj/wwAzoAscaED74xvS+mwF6NKx2qOoOb2rI903uSehMWw2S6cHO0165
TUBSFzNkjhANjSdjWtQLEFrOqOUR7eNoDZguVmWAFibtyOwkyQN1GG8I2p8okYvQbL/nyLSvR4v+
m/nzUvy3Yi6vP7SXAFEIJLInZ57AZhGLoKVQSIxRiTUZOjr895/hkmgR8RD2DRvQVbdqkPDZU9YH
LDZKovv7YoyHwRP0vkB+1EVnQP0dbhuwwkVKiywBqpDJnhozKfJUuSlha2TPXEzxbdNWB/fOc2ei
9qDsuZxYdDxcQ4FQKZHvgwSsHwCgKwdg6bjFMkdslnUEDOTXbr4YeJY5VDHP3oPe9gZiGqy43s/q
+y+fKcbdXsOZ+gRaAjHNzsZrn/YHy+ubDbhh4eRkVyZZspviPROKxtsOfK2zW2hB5Jkc3xBgfitv
68kf99v4L3EyPcKPW8KClTT/c7WU9oXNmGPf5V6R341BR+r/kxoJpyBxuTdHoisFmctrxVORwbK1
w5FMAlvVcbBevzBTERAsPSuYKkhrN0UnRf4vx4in/cfzru7P1w7NxSKw1TwCJy7J7HBjqzpzIA6c
smFoJ+mwVgiwccU3tAZaBqfjQpybHkHkFgCicH9muMZIJ1/RhG2UgGRqYEQkQS2KY8i7xU3ocJeh
B4ypHivD/ComRWTF87UjmIFnWwzEDKAyw3Hs0E5kwzfvrVMIJuVRLo6sdd/hkMybY/Ao2bylT3aD
jkFP7yre2qlTBBfxYoOrVQmS91wOr/RI6dzkvbUt1seRo7dTQooBrnfuMMrsiauoMnh66cTmwVzr
QhTrG5UVAiQCEHJN/9trLAnsCjrSajkGcS5j/sSxAt3SIP0mBr1pg5p5wvD1cZTUpuYzdNDe4Vpg
ORPUwSOujvljv7/z6Ao0lYaRBHa/gs8wL2rQuaYeYpIuvPbAqR9bDBeg2QAt4JX+LJDQ9BBc97Fv
pt9TKmexFJGvww/0jAM578aGaU+7CnEl9T/rbaYrCT6am6J8lHBK74xNzlpBB1ftPBEouucE4Iim
9T7X8EreVUKOI8+MWnTIE+K3RAPzw54231PuCO3tH+GhWWYNhQfNJqlXzIbMf1SM4E6ehz8SeWCc
qhMJGXpPEQAUSiB1earaOSTleoAxHr4G9wx3Eu0V8iANYIoWZ8fannIRQ0sT8KRXWmirDQVh3TlI
cd5NSDZAuPP9UqPgydo3s2GTPQJPaWTENxJCSA6/nUAaAdCVxR70/q7mZI2pkAL4Tr9VwEYT7hqz
kasT+os/UYJutw0702grv1NwKtsJpzB+NnI4cNBoVtXYmIKyweBBfMDq/fgmF8tTnTYaczceNWBe
ak8a1RpsOe9lp/gcbaDEXBvJpW1In9g0rj+x7GnvzUZslEY4NB3TU3p6AAoMO16WeqO/x7tN1VEZ
6H7KxlpRyHB2yhESNy3/gktL3wjxacjQ3qS31YmsbrygRPtcun0bPoXxZtYFMEP1pvdob9qOTV1M
7RJfGhmSG1tp/ZjGoqxY38bnyl2exR9mrAtMbvjrmEtZkqF+2WdijNilhl1j8UWueV5tAY+WhAMH
m39MAmB8fV/kSZXeTSwyeIkzARDo3QqqE2I8wLqePPxi/wBarRky8sQKus6wiDznKAnNsyKkRhl7
Sq+mlQcNGLNNCunRXHJVwuxBplyvrpayFhVxXdWzC7h57iROyCxXXloOHMq0Vr7uEd7wMZrsg5bv
aDKBgR3565Xcwhe8/zQoacgPc6CG6cQFUvJ+D3OCkZOt9C35qQVL7DOO0bz+U3ssYMYMcqUCtctF
6K7Ehb2UQF7vnF874JRJs1S7AI+4XdQNpDBjW9dzH7w3Ju4+WRLTPrvckvUyNKTj5lc/4xcUYyO1
f+V0JDRaPvDuQtVlJA3of2VIxp+oAa6NpKslF41JbGfq+ewLN/DCft5VmVYnLAe79hs6NLxoTBMC
ffC+gIxYPc4oKomnFZ7oEux5fY7SElUNV9x1w1AKQeMpoc84/C7ImsuXIkhhdrSyuoJtNKNM4UJ5
m+I2hr0eKi2Edm4/ZsboDCIOzvsK4u9FYWyYXXP1xstbLDNESUjY2ETEKXCl0HQ229+vYd8BinZq
0yszsxOVhXLz1x4P6G932wf+6irRYu6hHG60aiEYtVyG/0D1PQpc2xx2UQdKo8RYpR/oi29y+6P4
P0vXzFH9hAIoyAcBkw8eSH6s9CYDziYdmLIo5nGxnphDS47AI1CZPHxPebIYmoWFy2unjORRea5W
RJ+/ySEQD0a/F2bhptWhiclUoNc0IQ9lblO+FDh94CPu1mRBBO/lQbZMeHRX6wG9TXYVJmsGo3Rp
VPBL0hKZ1vxwlA8CCEc9iWz5jIT4RHCLkiELVABszsUIoWvqTlFkCj6cr9yxlLmSXqN+qHgqxOQ2
ZDdwLGhKxm9tI0cF8Xsc6WIZeecbSWwEU69wa4eV6moAwHAPVgX/rBTlYXm9Vs00ZazRq7yMn8bv
f4aM4MFKlBp458Ta93szBotECfATXIwrLSdCDaHoio7fa4q/f/xhPKjbwodTVY4uiZiBDfHXdSVC
C580FvZGkl0auexqaK9p7Z0Eo5AeHRzJ50vJq+V+ZqXQS70qP3NKDQAk5HGNpi/m8wwezN1N/OMX
aAPnQXS+4gJ77rnLus9z9rmU0qOr/67EJ6G9o+xaDD5BxuRmfTgD7Dxy0pDgscBeY7BXS4Ts3D8k
u9f4Qj15TpeqmfM/MK0WIyrLNRBcltvFWvPGglau5/6bpQKsoXP0GN5DkMJGO7l0g36K66gFKPQ5
0/UpNOX/rIdzMiYlIwFFP75wDjWSuBUWyPSBklxkYaqMyG2/qUR0/eAefODmyEkzENFlPiIvPrUS
qcJEL3CVNfKLqAHKblMj1djh5nPpZykWTdoZdhTLSd1z7xji9wpW9IPl0uQjK46Q2XbDvWHCufRR
Z/txzc0jHvu7B+FaMOzggFStKN7pCoWCyzwO9h+J6XAe9xMZnfqTkDNkVPZkE9luQcQ8jUeiOu4d
9wcNXeL18g28/3DilUd24v3fhQvxsN+DBAEfKjlUiNh27HLdxhMUcFfdd41jihv4iuKRyTQGvgCy
zLhfT5J+dXJU0du+SXpRi4OODVA9hjJEh/mhnrZBd0UGa5rDlplvHcBOxulxZTjdscJmlU68UXdI
zYjRpxOxT5Te91rrWw3ur4tIM9TRlvAz/VPlCTumy/EaKpwXLOawQdqctUc0sNvi552kjel2bNTr
4+f6CiyZT4BiSb71CHeozzqwUwIssXhBjcCxU9z9rtKIfw1Id4Zkcgb/KlGUn/z8Q+jfRaIde+9S
YyApPCAfNt6z63kK1iEd6eVz0NxHbCxFkJKNFz/RxZjtx7cRw+utcsoIczZy2LNUhSZbOj/ZJp7L
bRQtPLAA6rAwYLR33SIBALhJTtPWkNCQyj1Vac3xOLg7W/gNG/Jp1QKmw/PzQ4tGWxuGeiLTnIot
Ekb0FlrBZIxqOZgazOuBRjt9BdvSeHUiDbdWrik5hRoJ3YuvEt4mWkk5XFECUCINrKSv0xk0LZHI
z7icLyQgeY2OzQG7TRvxuU9wGik1M4KNUnBohlOEf4XcNlojYSTc6js3m1zoc8Lsq5QQ13qgiu3X
uT2oQiP86GdtFqSTpSuVwocVyexTYHhw3RVRYx19igVzf4nR42nrFTDN/hXvv4z74cg5V2QJ/1K9
o3Mi3M6JMKbXnd7gg72FEzmpfqpTgza+Sd1foCafXTZZ5h5Fh27jr7qMuSkTnR1n8mtBniunKm1R
pl86dvnbBCKTcEe9o2LXv1wd2EkkDvcOv5W5eb5IRC/GfcuTLjFtQBona7AXyES6zIk6YJ6ytJGd
qetG8pA0MwLuzet3A1U/H+ccpToWHggGFkyCh4+Nna7SWodRkEgt4K9cZACs3jXvBLNN2b4WKrow
c//nq/eH71u+ofyAoVEuN/jEAWZ8Kq6ZRsgM6zjjf0DJkWeEEru2qHv3sxXFp1JMGKw/pWNkdNCo
/6hR3lNECT4ff4cPrTTfEbEzCA4rbL+DnwE+VUbcxWxsTOBWih3XKnzU+oKDAMpk3MiXr7bzNaCr
jpvVkLDSJESAb6voVJxYb6uuLR902FdOxZY221u0HYY71WLRg9D72iWv+HtaHHwkph6TBsCAc+E7
Gs0QqCWWJCj782QTyya0ahh7lMTuo7e9+sqXxOQQbK0WGFqgRqdTPa30D0Vefpq3rsJ14J7nDR1f
HDms9N7eYF/BE03WOSj5XIZnEoMVz8W8sW8BpBIXeTziLdA5yoAqQpLj/v0RUMoQ6E4gdixlPahy
Aj2L+7O1l5bFpETVobh7tfZlC9AMH7tITQFjLT/Cc2chiP7flCK9WeF4v+cPwX6D/tSq8j6aaJfB
Bf8KDxxlNDUfLZTAmb/A6Of5qD//T1BsBhNWRErW2wy9gSg7jBdadchIQoiOF7QmujD0WVUyIaXd
h3jM4/scx0E65t1VY2PgMlCg+B5ad6aGzJJrPJKdYtgtTyNKTQOlWCxh6bskjEYjfl9jmFq+SreA
7271o7cWM98GXWQOReOawZ4lMmyN9XqU7A6l7PZo3P8SWdLHXIDdubXlLyXVL/CyIRpsqPekM2PZ
oIp3J+JkMjeEnxt1oa8XEhAhMyif9o/PIwEcUpc3YZtxYzbrKvnYuaDAt2p4q30C7Af86saV/2/R
iZzkTEoKmN/hj0epIOiytAg+rQ/ogOZDX2PABTuJyKuVNvfIaKLqxgBxS4q5tH6szQPMQq+SofuO
zhIDpvcjsWpjHoQGPtA1H8xalfofDFmBxBDy/an0oU5RraKQD4mL8maA8v8iAfJlDMiZ8NBRcl5U
ANIRKQa7+08FddH2n/QLJVo+G94UYaHplAJ+xHHo3L5BxoCrJT6YWteojVN+/Gtwf6+xwSPmrqSB
+2n3GkUM+niGRL14AMHFPQ7RKJxza4iWOdgcIF29/VsHXNzYh2GsUoCXwC8gvtrSg2EoxaquPiMF
4CGE0Ud5VWg5bJRDko5a5S+rYZwKUbKdHnTRN9LFReGEG3U047P27vfSg2rQisqWvJ35+YxhEZ4p
eI0Zjb6oS76KM5pxpPl2n5C8qAMA+yO11JvV5t9ROLmANwsK823B7FKFM+YtfCECMyOZUOjJhLUA
fO/cNdj27yG81qc4sbnziN5nrDCF3Cbirr7V5cZiughagCE1UHxFgaru8c9N39b/zsUrKssJ71iS
V0qykHBjxsaUhiS9jVsA61yc2tE9BDZO/1zq+fzhNxdMVSkHKPU1RDbvEwDKryOLNXrhTbwy1C1a
aLDlwdYqK8EsixgZ0x+m6j7Im2TTLFqe5D2vIQQ27GDwkcqIbZaEKysuTKew1rWbruwPiRHLkejQ
Icp3Xt0F5oq3WUl/M1wVP759s6ybpGc5QDFAxjgb0vLfkJYriUk58j5TK4MeRObqrhYK7413wBA8
4fEv2w9iLrUAxUyHdYjSmGWq0k8rlcZyG+o2CCKh/ZD/TDeFd6TCdlUMM1wI0hBCofLocSzjLpGS
G0ibq5CqbspLFx8y6BCEG+/ZGvloIfWXmZ79g6bkXFfXmKLkqUmU5Vzz0BX5d+xaRARvfiXRUxfV
9izUs/Vqo0moHzcSZtW09NaxRlwLnqQB2m8lYkoSXTsqjgwX2p8XexYwlEnkwv8/GHrQDBEXL3a2
xWoYWLRlDwtd3kxa7fJuF40MBAfB34CyApAuA8823K62r+MuZEDQXLeV6SNBEPYfpD9M5WKK0TO3
srtnu2BxAjK4PyXtF4GVB7m7BnPVT51neFEIYBW8wDn1FuH9yanLtAwvNIbNiQ7JuABf/vYN+F31
M/UjnArDfDvR0v6Err/4TBjKyhHLM9pUjBA9xunsYpkfKm9zPR4ZFZIcEoHF+cpuaZ39SxwMpy1f
dIDd3Eg0JGEdDlZ7bZsNwo1ffKd1htBfipk7E7aFRtH76hWFNR/LB+pvt7/AHwthqAZzPVLAF3qO
fI5jYx/zrg45nq+WPs3NpmfzEh/Xj6nbujqTpUEnh1ecEL3wbpPxHS9j8IV0GOI++KZyQu8bgoUi
0O4tAeV6JzBYQMFYa41f9DK7SbhvmlFUi2morw+Ku0kMpEKNHJyY12gcmOlLB3odCvb9kXB5zONX
KTVPOVnvKv2DLB/GdNNT75xa6leZZYdXfVUokJCUjfUweJ7XPDqMyFsm8BjBTYFeOajeQ7iLO5dI
KUN0WnPomJYjfiNdg7V9XfOJCQSbqjfXBTWeHMqs4ZVSVPxtylY6z9f5sp97nzYgPFlpPcX3NgI7
/zwcX352vE2yaMwgbhzLMFSEr35BqIXBAdRpFLZR/GFi/PgI3uX1t3PBMJHhxZQZ/KZc/O1XKw3b
1k38DEYF/Dk+juJmvYYcDcQUxwASYks3IvwR60LiEcl3sikcQUvoqubkldZYu5cVdrkDWcOvamns
rRQbJJt+CBg43luFvC0LT/bD6T5DhKh1TINfxWxwI8unNk1lYMO76Nb6WT3h1JcDh8U1aC1TqbtE
p2xmkGOTXCXkdoOJ0KF+aOfQnQ26WTjYAbXD2/mSzPwuK88RWkrxAYnNyKmcMQI56bgkBg8scIVh
MvRMLiRQeIvVg5ZJAJQkLZFaS9h52XeH6I6Ixc/i2LGDR0TIMjP1dSXYA0MxIvZP1OcCxEodbqSs
DtLMi0ISDNPv96ycWcMO8nd4neekKlP1veQ/g8MchfCAb7qiJ3HwNs7u3BbRF6QPIwrFG3cx77oR
eFFPktXi8JDWCxbyy8m1wk7GlbjQV/p+f+R/JnpLC1Ijn2qw/ZL/kVIUtYvg2qXmYcanWNx80ZAn
NCCM+s8s66GiL4vZPbsQsMNTbVOLnDH3HZHDrzteeL8MvPrSRjG4MEMI8eP8/bK0E4UWgBtdmdF/
oNUxUMaZWbpwf3GbeEmyPpjYtkSrgUx7Jf7+UUWcJnExLsLmJFRr/xeGmK/3ENM5ML8R0cIO30JG
iXCcP4e9wqSmdhwU6QeFv5uKlj3PpFYsdJ/CPORPOYrCKhitJ4S9ES1QvCkwZHg3+7MIgQ1mwzb5
PbifgmsQOiKhOzcAEpFETM5YvFPOgO1e0xKHoOR2mFOks1wB9Bq2WJijz5QAbzETeWvMeY9yUIDI
hiJsUrRulzBGEDWdnYWHtE5iqel+0n3kaPUCsgUVtM4KABNjylleAx84RBhf+zF0uMqJBkk2wveG
LEaYg4eSttMoUdSiR6RXHJFITpnRpq6EtnBRWbupu+Yu6tDsYjXfbzI/X54gpLXtCISEGFtFg1Wj
+a1kpq2fGuYlxfAInprXON5o4F/KhnsOefWxr8XN5sXUqH3nclRa5jGCDmzIRuubVrkaaCPxuC1N
zLGjQ31D4b6hW5MbN20hv6MVVQjydbERwOlVdP99X8/gGy/Lz/1hCO9+aMfV/A7I6cgHJlax4nY6
h0i0nHRhJZzqFRqam7Qpx4YkU+ejQ7zeDBXWafosyMnrmiWXINcW39PgezxOQhGpe/i17K5q59UD
SmtUQxXq44TsENYaZJqXDqD5+ecShMRsVeMwZKFH+uevSvPuhN6BkXAWsNDQMDCGfTl9/zCyhKX6
wkSuu5EBi6f7Awid8eSIi7IKw5FN8VL3VXH9kPKmvgdFcmt6i4chaJErpvkqWctCG0msHPiCdWZA
bh7JMiiqNbhPmPbSBYb2bhXXdOiqfIc2iPM8S0DcQE5y+3X2L1hEoKgN9b+II0ppk0yIm7Mrn06y
EssyOODCWBR+PZWqvuIoFaRQKBLJSvydfCjHj/oqakNn+rDMBL+Imlt5c3GQLURXGZ362dJH3Iua
zBX8H5JXHuX1Eq8efqSwzPurSeNGuq6oLdkP+9Zs7/Fm6ZrUm0xECpROWNSVVIkFGoGdxX/jdxUx
RbFYYZoo9oOZVtcs7gKyBVHVTFFGVCJaj6NaT49u/yjKZ2DlU4jZegl4OGOs3Jl97jaUswcvkWH1
BNrYDCt4A7lZMW1v7ZPkejU+DT4I7rjMlqUVi0XcUlbKg8SI/Vji1TvTHE0i5MATT60msSNXinR5
Qg3XrYJW2imdlSf+vmkMYY7JmqeuSTgWp/UawK0WoNLObZVDQPHuryHhZIgX547MU26xSSSPE+Fg
2f28unk4yjr51JDUhmw59F4UQdRhTcKuKjGIcgew9BxsoRNtU+003nzbkTyevV5lACTc1jJodRzJ
UQw5mTBViAly4j2rA9tDXMwYIM+TVf53wxjRRmegXaElHty0Q/eBeqYLQG9M87oPqTb+A5V3AILM
NaSsP/Pf8r2AqotacGyScXnucoq5QgBNJknA3yCsgzrqTKKNZMwmx8THRiT4cIRCqseLnf5m2GbT
8q8RPxcennmWWeHRcjdv6MXo3CauwrhccyyNR1qgi+jQAi9GLVDZkG7aAnE+nj3tLYOGAqnOtHu/
YkfE3uPqrXL6OTlAfeTcCTVIjZSEQo+HklVuEacAr4AdwjleRpj4OvlzAB3tx5S0dCZyYIVXUjQY
p+ZtxYtrwKQXx5bjl44nsoLy5qI2kpLW7PXnpJ44f63KVvId4dcGBUmnNL+1XQ0MNO7+S9AX6Ldq
kTiX9BBGryOq+48mW7kS5LoNet62T8Ww6h+wP7DxoHB6AEsqzSiKYc1WQCeHVLaLg2sbQ29Q2CC0
H4DYK7CaX/wCdu4+RxDC3k7g0/ZKfMaItauzgi8g+/jplJN29ND8u8eSBReVH/ssXO0t5Y/z+vKD
Qr7fvADL+n0UYzP8F8OpdG+rqR3thqAKXk/LDIVGUoSm6/0TQTMWV4emU11TqnWbO72Hko98oeLl
iEILewGDPJScg5vsdXJKJJ0YqB3YHHll26sJ8SYIEXEgU6j3PcUD0X85zpFVfFVMZiPGvVpZtcI1
3eBpWrHdb81bfKo6iwj0DU2PKKdHbM7ofGW3DwLgNVNRM+t8OKJw6RMYOX0QG2R0eq3o10ef7XK8
i0dB4prAzV1dobYSYGd8kRdGtqHopr5Wg2Ll2RRIEKcZuNctM0kTq6vnkrSYl1k+FQmbT5Gz/DWI
ZRcHXhlYiGMmG+65D6eUlcTzh1odvKHwQxmtJ7//37gBEUqVpmGnCPm/5S9bg0TN39yplMTbVpJU
RtQ8xG6o3XFkSP2VVX8RvGWj95lVE7r7/zKTuiVflwyy8dxc1nAcBACTILA6Ld5zTl7Z+EaiktsB
ocdy44EsP4MAKZEOX4xtdU0ZGEoXAXD1PuV/4I42BUSMtwUD5e2Q0NR0T2P3uzMFkBFP02GKYmag
XrzGCYsKiu785T/DtFvRnXmb/UbIekJz+fbRViHbjoYj5nxdEH0zy5E2cJHrWMRxQC6qLqJIOLra
GCqb0kwVM9xfV65O3ToE72uMmUP9Kod0NraP74oppUXgrAf204BAbCkZIt3EWhrunZ9q+z6ZM4dg
xO3p9nE+Z305HD1R8GRiWWRinBAlAFhG6ow2DpwXIAR8kMMeVOPC/jE0qc+7OcppXwriw1qttCEw
X0b5F8vTOMDSy5ouXw6+HrwjkW6pRGe2fYnBUAEydCZNiMCKvC0ihy324tSMOUKUcMYWHRa4LEkF
NY0ozxR8eteEdvQFji7WUhkNJ57XXK+RRJIvsbamYkuC7+9GtrxXTqAVWiV37jHuRrvrdNG1Iq+7
wJ9OMDqNtNm5QWH83D5QeZ/W8b7lULdR1VUXZFzyP5Bx9iaI84spfa/1tZppzjgZgY7vtrm/6Elg
6B0DgajOM1iXDuKVUUwsofFhop3DESelKmZcs5ji4kLg4d2sdSQ5/PgDvddd9VP3Xtanc93hs2Hh
RI7/pHqZksbUsbjIBNAbTMWxswzmn2Qo9R34l0ronNepfbFXdXaafo7s2EFPqUETT3r+9DS0WeQb
ZZkDefcHPuzuD7/uizJXxvxrlYirwgoiX/5lvcVrCGfCOPVdgxLklQV0CaCxnOZzCH9tUA1ieoNZ
evsfoP0F1TK7LBSw9oj9Bl91j8t74eALzUVdcj+AFYMdexP9xMZHhizf53CjvMbhWQ3woyhG/z3B
ENwMwM75VkWSx2YUEC7ntbAwj1taO1NJ6jKSs2xRZgNwFkmqpoDgFLWA9+eAfY5u139/zvLjx2n/
n836lnsK4RvBXR8/bcjlpPwlgy6zM+BG/sbxYMOnqJn9ry9gOfWbZlkrXMVOiOICz1k39FHfHdsh
GEFf2Hd6Vd/4nxCMmsD3oFVEZrQfMiqWoxqhsht8s8QuWXTRiYGZxDWQCXHU3Ip/P1g/6TCuEb3W
mggkGqyq3D/ULWpseK/6nsT8Q1QEgcnhgq3+MaYhV3zstmp/8iVye+Iz538devP2wBY/M85ZjtAQ
JyK8B6busrICNAmH8GcMxqbYe0Yn3f7Djms2fVUoajh+JXFhVhPNHvWwUIC+AFq2gNmME3MBCn0r
P6quWOg4wdTX/kEnkLcFPeLPCcutk0YAS2wLCfg77msZq8TEouKQDEyxnuE5SmvdRxP27vKH4YoO
pWJFLeyRUZrxVroSYNGa3Lptvs011lAV70u6RG8euyPRw0GcBxLlf5oSi8mEwpIoUWXHSeifKS18
AjXH+5H8YYRsrk+UzU1lKNu6M8+YLXm2dktG2/Yxa2MDcCokUacyd8UwQJxzc73K4sr6/357S5l8
DgNJ9CWFllkrAHnmdRlNMpYnfXBpo8WWvvfqcbeaDBTpvgwSW8ouYV7HIYIUtX+52AYeco1DVAMO
l+5WPKa/9NGYmqrCzYWM/1IBrudZEG4E7IiPL4cAfcmOamNKhk8qH+oEE85SC+Bi7ZiCihRKScu+
JYgC8qEwQHvdf8PLIhkfPpxCDw2ugI8HWSDIm1GokVnncUn8JIsJGVbfLwI0WAo1cNxNem7UkwQL
TMYR0lvEI7YyiiRWaqe2FWmrUEWS6m6GPyXug08zOSdOncssqA+TAsWfzbqylwb04DcCc2YGAWPy
SkiI7/deZXpoF6Yi5gl6MaWVePRbctnqv90vH0RR1+AKIJ6KpLUe3Qb6mpPoZErE87YWR1XOlpwE
m0mloFrnmAvBsV1U/0wj26gmWp3ugJ9LoEWYqRDsaApkdAaC3LZWFXSx6qW3ENh6bbadQ7Ms+zaK
bB3wG5e1l2vpaul8/LJgYEWxBxosOe+8Z1ILj65CVn7gVpPeVF6SbheM+0it53S2RMQ8Q9VMhMAY
XFPc76y0cGXvXKCoJP21edwkrw3dvlv71lfXzX0WH57ZpgCkD3L/dg0JCtXE84yeYy2RA5Atwn3f
KqGEEDHHqJhwI+g4/FgV8qLkbwNY2nFdZ0dOfLOD/N7dKQhxgd8n24tZupHJf83pBJ6yjR/fTBv+
m4n2TaQISlgUrfsZhGlHxKGRPRGVY29MuSxMU6XEtnVUKNoBmDQMp+kYHL46Sp+vkXvunc98dpge
4zcAXnRk97QUaHM22FpE+D3AjfFOJ+b02pjxwi6MajbMuw0ne60wDziZYQ6WZsIQUbaamN2DSPmO
cryrE3FvdwqQtbdflOkb1+/sl2a/KjfK7wyPGk5T5An3ugpZh6ruFtYhshvQ6LX8iNMRD+eW/w4h
sdqibjGr/TjiuDUSAzcNmTbj4LBp9ML4GA6vt3RCj1NzaLEHO0vAjG8kUWpPlDHFMw/73yZwoQLG
Sr9suctbLyPB8SWFY0WFYy6+2TRMB9750W4OGLRCLJtGZzj8XRWcSXWzb6pYkZhazs6VhSwOCyy/
gO4+EBKgZLqhiyDddYUTiJpzqQEHgY1qK6utzEIpXQzA/Z6P51jhSkayxvQDEG9lWkDYh30O27kO
sLqTWHxnqq7p3yYRNY0EvFa/Ke/U7Q+vSD0y3hq0fdzYQs/xh+h46vH8L9hGuN/FARQgq0soMCg3
p78P/aj4Lp8HLuTZrjmHsnV9myNDlKX90vubdsHEIHuGBoQaWL803ovGtT9ewdKBigBEHpTw+jJB
66og7fj43SA1uh1NWYtXPdwdkxvWTRzOIVm36P9dt7TYZENND9Vj/3aSS2+5iJt/tHW7mxT7cIwo
WDae+/6EXk7+fhzJshoVl4hbIJ0jv1iUjXEvWEDt2SFMQMOLArv1L9VJLDZFhn9TD8AjrpKK9kYR
6IRJby4HrQcBxI6esbPs7jwTLLSCJ9PFsJzdn7Dn48phA2pOpTcYUCcB4CqDZ+RhLknfISH09lVc
aUFstblwncY/4WsbQoeiKBuhsSnBvNlGMIoxVQVBB8LeGzqkS2/vt9VkhKTxmvY9Uxo667CKA0i3
4OrzwTIiRHTgvRpDTR1UeI0MBzq0GD41KByt1lhvsSfLz6LpCkPQGVdITbPyo/nPpyWEd6JysadL
AUhDg5NE+YEiAJ6CZQQAvCneftKUstohwKfAy30XxTNU1TI6hnk/lDriss9191Wvt0Ylf6cTS0Ri
qbQQLeXsY3u88uaa2dO7ZMTI/+CykRIsuRRIt/VjC3NTiPoqhc7sq0FyN0zwHg67Hxs/GHmuDLS6
EipHg/L2hGv8KmRRkwx4gg36N97oMhQ8VpNRGGimAF9a3Tadp12gBxcCWCqKN/OGZa9HZYanXj2u
Uow5+2n1zzsBGgZunZyAyuQGs1WjT8F91ZTtJSsZTlxk7z3J6+MsX+SsJTe+XmYI1U5My+/D3+ld
zMcZ+gIfOGO/O2lOhdbza3TLzeXJiKu6nhsb9wVnI/+Ds+4MCnvCHf6rclvmC9R4YO39lWxrs3Vu
ID4IQK9vBIPu/GGGR7s8BO20CgDfuNBP8YUvPwF4IsE1IlvFIDlgheTIPZANwviJY8BetAIEHwCU
U/U90GZk/wQSoH4WBw3rQYPYwYxnrpJeDiJUyMJq32Z9O5OOxVx14t0SqJBcGeyAdnxDZM+8PbPT
7NOMbmIc7znWrH7TVKgnGAqszCNhvPvvN28KeuUAsYoOFC1rc77sQoVfNJ9Bj10drtfQ90At1rDs
IpCGaPBb7nSnKQ2Y4VrIrDtlOVgCtEle0AiDyllyUy8eJ2CKtCtvuaj1GMLUYwX824+jXsj3/YDe
f3uPPJRMEB9Q4SKBe8oO4XnJu5Hk0zhMZ6dbBHiKF1nDb+3AuXdGqC1+CHf+9fgiFieVs3/uilIy
2fqjIQBGIu0gWGmhsmgJdiknczA9KFZngH3l52DQFaib03pBk3A0krb1DCMDOBgJ7pl+GDCR0rAm
i0fBFZn/IdfVyuRmf8/PHV1ZxJoeHCyZnYdN9E8vTJAwR4LHexqIzuEH9EFXfPHpgXz/49UZPwU7
VcILrCSH2fyZ97nOJC9kr4debTK5apYSqcD2qIU3Ho0Dk1jA8cRYNdsLfgm6s7opt+z6HJvMFuB1
DxjHCraU+e3jE15u2KA3zKJQprngpRYKFy/b3nJKw8upmzEPbN9o3cgLF2rs0fKMoNNB17gUwG3/
VigC4//U1RdOLFVn3ZbZLB0uVNl/Q6UpFYABuGlUqckY0wZn1VOe7UP48UPhF+hHjqNP0rt1QTAU
lwFYIvst8Bf2JEza4r82Py6jcRyDx12PzA0nwIY9PbBsqwoG+ll3F/jsevJB+iubvYM9scgdgZ88
fgOk+rWDYUy9LNl4bYZTAcwIYc6PpUW6LkVb3/7porb+vc8Ahmj8DEF0zCARjiK4BrnZRk7Ss5on
f7ujCkiGdCNcZvL0CM55MQVTIomWhywrr7WALQtFaElodG6SYZoGqneylc7zp7X9cejch7gSdXUv
MxdYvDlbNieMe1YuSiss5vQSPHIc5k1VrWmduinJyySBLNFdd/CXqLYe28eXDWGsgY64U/xmyAIL
ENLwePl/CFn5aPW5xzPjUW9gIBJMqSPkuR0VBN4Qiut/yud7xftxVWf/06vnfkndGKyZv1v3akFz
++HZdCyaP8evdMpI6wqwYQW4p8KH69CWgR0sZM3G4hvd8u4FROXHdPxBakeGHhTVE0z0qlLkAwlf
2OijngHuz/6XCb9HrbIXlg/slJ2hTIusUN6i79pUpq6tTu+ljP2zstfSG8d28O1bANYXXkq3ulbi
0cWwmMn8pnfDrAtikqYM8XZ1zsIxZ11M+X58quSzxN0JJgPnxCwD6llojrw84+rA/YSFb3r8wAy7
MhdwUftJNcuMoisiFTMKlAjk3GS+LqKyzuCJtLFe6U5jW7Rlm0kDuT6e524eFSl1deupQC+T6+oP
7vrofjOuuw1jLI4YnD9gUz/IMvEeiXNxzg+SaMhHcwt1smBjGhSSl/nMAE0+7yWQuVkBPdm9wN+t
IIsHyAN6HPSQ30e8gIxTdFZ3yvVcbCdQu1BMWb44hrXAf4Dknp+ZER4A0D4zS7wL3l3AAj+jv3ah
G+iW8CuH3caqgrkZiw4jnSWzrqS/xZBXEm3eGVpjcCImMDHiW43D5pql2KUN1AK6doCZIre0CneP
yUEN86Yv0R+BTTbO4uwj9OkVc93vm8GVKkpb4VC092LHfCTJvPlxLM1ao1AaWVHV0ZeBSn4S86kj
+SkiBL7mOraqTj30cslApLZae/zEk6FjtkPYLTvFlJgvBBKBqBAap9boqeXCzESSOeu2XuyO+1N7
ZZDAIF++6Dz61QiP+35KRCTc0EsHdjmnDX4wqODsseGyVWCeQk2HkTdXYZ8cJSEq2sIVnTknHIIX
6wE0OusW+gQl8rDdfIbpTGZqV3HjSyr7pSZucvUcvsp//NkEy8zsoHQTYoewsyoH1hLa10jByVZC
1exgZILqtsznPjP+j0yrF2j9j6wzW/nQSI6MLH9j058OuF/WAEv4Mc/IqyRP28Zd4qMBI7AnUpd7
+mN42oKX+dpQVimHy3D8knLrn4V5dlovGL5P9f/klo4+OA6EYXWnu33ST650JliR4whXiocwYBo7
FeSYPWX6pZXTrOMHy8wHYbvXH2dH6MC/qk5okIG1ojt6qlO2E7gIEPZiAds033yoGn8DN2u9ZWsT
ff/n8BXs+gJNXQpcyvrmG4by1YFcqp+k1be1TWQT3tJErg2CaswYcpkDmskN2pJZHUx0HvzIaaJP
xpsFxAFE7tkCmajcKCo9vFJBdDSrVwNhcR262RUmLGDaPrVm78rk2fTlcUWj9c0gOROpWdMyrO9h
6mKPVmjkeWSvF/pKNwxwg8d80KPNY15rKmUTexxSvmwKbnV2KiQ0UH/4xZ3Ie4cM/9u6C4yg67AU
GE8X0cWTBMAh0Bl4dPn52vomV73cA+0gORwLkKLSOkNEVOsYhqjDxQ+TI5qzSZS+LE/hsWxx8piG
oTmxm3m5kTWOmDtYHOXlyZuNit7gsfcSHfCxTuhhR5oJe4GGvVovuoeQYuzfRECIwlBinPY/aHZD
3AegwyENDOnAUFrODE3NfmYyc4SLjFQpIIGavQ+eOrXaffk7QHg+NcxF8mt6W48fRIvYIIG6UZxL
o68MQ5vU49yuv5oIgOgeiTHTV2FgiAFYrMXSSfPD/H3fkxVX6eS1EV2J01namsb26akx6IrzUdR6
JELhjTtBa65+9JTVmYY3/JfCwyFr133XGP0QczHSq9u1qciS2PqO8TAPWVwGsnRZx5WKCHm5kR0D
a7386BnwLQkStAF1zZ90FuxwvNcEtJuT0ZcprM0Ko5mQVHvYppDDkImdqOh3abpOGcexEEp24Flj
vVC945t9ARwovw1VBYSvN3SINfTknVHhebGjBmCCvI9Bvrs5wLNXVOLmCnEo2tIFfrfgIUHJmkOH
QY6bzQycfenGR8c+OTp43tg8BSJNMypWMX7SHD5dzcqQU6NSi07w0H46IJ7qXcXhNJ0wWjfCuWFN
LnLTLX6i1qbeL2TEWZh8yR6ZxKwMwn6h0kwWzDKThjYDheN+ZPWI7EUHq5eWQ7E1DNw7i1GuA3q3
Eb2fCuFB+G1badO/m6Fp1STbqIY9MTmfrC39EN/C33NIZOZNTOGp0bnKOJTUl0Hv0J8HuoCK48Cq
12rKIj9+irxt5/cTxxDgWizce4Zz2XTogO79hlpcy8AXqWReFmA96/yVlT0YFRQB/3j8wCyKbldB
2HjHgIAnMHOP5C3q/xrrvPBbYVdQaMWNCrdgTHSN4eJT6890bBi/4jM0tdX/PiEEDjwUHO2y3EUR
uvY472NR4w9sZ1mxE7pR8sZxfMJ8Lni79WV8WMMiKMbO4SNK4xPd+i+wWI4RFIQiov/gsrdpVsjw
sa5mGvSktdqYPgejpUd834mm4FHXO2iDtOGfD6J7C+PdgrwxeYbBOjDjqeafYnGkDyXHOcTWA9oE
5dc6tTVuLd5Nd+Up8dAf0Kt5kv758KqUNpxPfRJtESh1h3eP9imgcCeHa3PHPSLbhh5YYIvnHZqo
cBPt08Y08bdSobxXpXnXIN8EEuIkB0qmpBiNEMYfJSi3gTYkOGVCV4BYaOhcbrIe8PUB/Bls6ZyI
/TLqEKbK5mSI/T38Uq+WSTmvTXtEDcXyz6ldJfY03NrknY8UDymnUhw2b9zM6hS8JlcL8fDARtNA
JOCY+Urq90DctU5e+Oe5l4r61ETcRDAYCRgdZp4im0KpbWnUhuxNDsbdI168nKlRZLH9qpilEkQJ
O4m3z3TnkHLERCQShn3wyD7Mo13y5IyW8NjVxQPY2XMwxqRXv2K1focaqZU9iaLYGU/FTzgHgBmy
X1f1x7P+4++7ojxXu8J57oUPpvEvgotBLcMw1lDuL/cBQoNua9Vjjk3H4zy1uno8tzuHffFfunUz
uJaUa9kOHktm1oWxDxa4V/k+Thn6zQpTE2OEYI2zWcwNvZXtR3Y8xTa7ej76ZQbSZEWi/Tj3EHPO
kVQxvdy2Hi6xgZebLco8MTd1RE5tGQN19hPJre4lMiBx2uoesPM9P4MWmxF5/D92klmoSKsOMGKU
TLmuKOXNI7K2LZGKIaXBTLd1a0/g/l5Q+iEjYsGtkvscVZUZnq3KB6UO74xFODwMy7segdcats09
Q5CuEd6ppMjwvAjK5olYi2+5ww4HiCidnpHdGrOkdw7I55zApXmla1dkG4Wi0bvEqbmAkQczmw3R
map4lHnSs9bWoplwSRs7ECbIPpMtWNaR8r5OX/2/kHx/9z7jRMPjzlKK3K5kjEFbAPHCJ0EZTi+i
sDaxOTV18fAq537Jed6zESVGeZ/euko59PDyQzN9xu5srxQTvK2HBZwJNXkzx49oJTxM2ume3W1A
TvneG6LKRYS9RD5rUqbDF4e0IOuSUzNpwu8MjQzZ97WBe+8/0q2Yu3R7lbstE6ofdBw5OG+sgNYt
S5OMs9U8OBe4/bXhSDkhvEcn9iVEMNgDdEXqigh1KkJwLHqOS3PXgbGfL05iJAw4dvzhEMZiNPNk
BkO9IjO6D/5Q+XAhJOGv4He5XCthSSKMcqrd28l0111PmpjD+ZFHYijUylap3QXWNT/e3oN5NCBN
U2OpG8FOFFpi8CyP4RCyqfrNYe2WnDYKeGLK68DW5UtWk0o6gwwg1ra+CfGYWVUgsINe+Kc80i6C
Nl1rea9EEd9hLQmAD4tatsy+ZrDSSx6XaCE1I/L81p+gHSQBEQbaA4TwiVoWdhtLkV1zTLOzO/ku
8MTFH3/hsezC70/oz1dK/eMTfT9NihLdpLhTpQQAK2RUQZurh6pHUDxMI7O2wL74vtB7nllBUEQw
UmDsXrCrFJD6RPjX2AB11Xbqmqs7ezAUzYCWg/6k75D24N3wimM7jMht6/mK464MZWSpW66jaSmb
Oc1tpbxOuty3CnfWEuToCh4BA/tpOzMRiHv4KGVEYlnxG+jWr27DIRrNydHp3/x45g4Nwugau02b
Q0lujweZmQA3mEgmLsodzMC50UQWk4EufxCiIhq8R7T3JNDQ3smrgapQx4LDJy9NIukJJ4a8o+WR
5XdSOedlxzcYNsR6w82w54BjT7nvkWoJM4gR26oSHQK9wLJXl6wLPw3mCXTM88rIER86+nPWXeOS
oJUn7T3bDw1qXAuTW85DgC0yiZgC8bcswWH3hh85Mqtr96DITfXMjL6cJzTN/EV6jTzRqNOnjJN0
K2xYHs2GbEI8PcmqFXGdKYs9C4CbS5jz8SXSKpDjTOYpnuwAGuNqbaVo0+8XI3/9UBSSUmInuv9i
IsnRp53JIz9wwpd+h7HoJaprmk+gq6CrFrUysKOI0+BJO8+yvz3pXsQm5Hgt2QHL4pFpEiyKC8wi
0fj2j/PTxz1XsZdPndv03mOk7QUhaBpCA01DJNz31/vVMM61s+ucM1Lykiph9Y3+CzYAtVvSgKZh
+DormoppyYtDveBDJ6SZvb6mWO2SOwvjgqKdjteFZ8+LCw6P+SkazQq2SJoRs1JeeQjupFHJs6co
4PF38p4bREwp3s2b4cZ/hXpwfsscfXTg3Y5HlsWzv13NO+YqzjrYa5+cYXqfmp+XpYjnthXQZGwY
FnKzUOtDTGkEvHGLSlwL+mC+Kml9/Wmj45RS0ZReAjrhsYZp8qnQxZfOwk+CK8KwQF+m+7huRR2/
SjUUB/jP0sTKOfdIkwf7uucqyOANHMea2fbSS8uJrKn3meVZk5MuOL7ZHRe9J1LY/at/2eqdAzXF
V5LX22tvAYy/AIvlZqYk1Pkp16Xhphe/Ocv4GkW7ltfLq88a3cxtp3Uhi9lxfQ24zHGG5x3snuvI
wnJLUzsD/eTSioo5bgCMLyKC+NFruRzz0XqtLLDMXVrJoUOUINVjcH00f00rNPIGO8rilAGLGq8w
apcvQ693CWuioAyDVFGKSTpx4wHCtW5te5jmn6TunlQNGtM+Jsk/+5F8LaTWvoKSx7POOJ1diV5/
atUWKO2FdwJA81L+qRcMPVnl3GHjyHxJ+q4mE20yPOY2rwGYpsXd8e6OQD1/c354/FrgnXU2EPM5
mp5exftrb11tZzEX2CWNg76a2puY5JlQB0wIc2nHPslPIwbowUZcZeYoejUu3Jr+U1m8oJSwz3Gz
S43FB8CkIVpobeiSW+ekCAVX+QENsisIlDUQfVzHjH32v/Zy6+sqE9LTAf5EoZxFZVOqt+46QJca
zm/AzyouO+ZIjiz6sIP0HIn6+a9nLis8yrp0qQeLRXIvCsBd1K9tImfiHg21IWfQpAIwwyAoRvfy
0ql4Npn7keVkCStBcl7MtwBwUtHy64O9LFhJ+pCnBasvFUKxI2dx6RWNVO5LzvmGrg10uRB4PZhR
e6yddsVWGBhSCl2Trenx9ak4bZIUYBVcMWz6JfCpM+kfwZD6hK4Ml6gE6oTWj1MIuLoeXkzAGaXx
4Svk435BRMnIntJ4C5yW3+V0Y1fZcb4bBdWGBVqVnqL1rO6PCDTihPYJwaXw6vkW6BO2ajzqwRK/
INVdsxnQu1vOvrKlnZwsIm+Gf8wFXrzjGFZPXgQ7acpzNLGu8cvMyNdwp+tLUl8ZPWNjjUKrE4zn
hcIwmNtPiGWaTOYUv0DpMdHE/tVp5tF+nfwIvQiDW6Ory297Y+Nh7VnkmN03sW1HusaZZCuh/iob
dqM9aitIq4e1mAAuYwQ6nN3LZeElxdn58RCPsmSjIztH0ulZnALkY89+IOlN9NbtOQon/U/+udnr
M+Ay/Z+VHt0SLHW8f/634x++UA2Gudf8+ShNH1F8nu1xeQx6nZNYxMvWCsLLahBv4n8yZoGpXafa
asa7CAWEx5TNQQw/Woq4vBmRXz1OUi0GDFRR32OopUomAxDWNULyQW1CYGKThPGcawnR5ics/NLT
/3IRUFCQ25jxcdrca4Tmhlev7Py/5h543+Q7QbkxMc+tZvcQbZ/GLF6FlAmFwlCWNilmhzn3edxL
BjHBhXT5Lla+9I6tPB5i4+nm1u2soUHGd7HaXRb6Zrt1zebAwAqULFVdcR1n6Ptvfo4bcaWkkZUh
l7qyRSRw+SwTig3vLCaTqcIuHi7J04xDhaYkpPVMQ2Imxjro1sya/slDnbW0tc2rw5MRUgujUnX8
FeINDeqiPzgp8LnAJ8t7kK5/C4UL16rZj/VyeAofQ+xz2+hRRpqgIhHINbQhd7+gdbrev/gZ2EvX
hEq86YndcFUmbc7srQomaav8Utp5Wydb0FyDDRd2I3e6wjW1nioN4APfQeuVJ406FFe7qJ/8xEPQ
rXDiZptlndFHpH/BYOM4GTJAg/gX8FeZtn/hGcPW9QXPi363bZJ8FSqI1UDkynJBRja4bXA/tpUi
6Qm6uXnGGXGKO78NImrpR3csVkaD5AEjxRwQXu06dWNSRnFWZ6XjfsgJMr170lPViLpsHzPhTDya
f8bMvZBd7fLgwN/Qjrqy6dgkdm+YI8JBLgVVa2dXK+RVfg9K+2kQy3oIUd3ekZGpD+pklQqNwT9C
3QPzrOynplrBjZaVdw3r8GRlfKHBCEAyO/FVxEfct2wbK6HkPpL2Jkw4T8ol52lVywl5VlrIPFuP
Uh+fH7vqsAslvzUUqSLrlUY5Y3m0ZSg3dg7eY5PRSHtWaQS4zp1dTToondvTdsprqHnYd/b+Dz8N
r1M1TVFsv6CMfVxvdp99qlGY2I6EymsKcAS+u4PruNt9E/nhWGpkB8nstlMXdm84Uak/1U7YBQa2
Pdqboc1lRVFPgIDWPdXm+bgEDljDNC5NGKOZJ+/LprLq2KeYFI+S6P8bbtbkb9yIP9wFhAwdd2s5
V7TtF4B0nlD/LSI59Zyp22wMTQ7tPMz6ya877yXsJp0zrbvaG/dyZkHsB1ihm7V8I9Qc6GjitoH5
JNttrFFywRl2h4eVkkkGPSLd4uSGD8pbnJRMyF7zYfzaq0L8AFzouY2M8922KTLrFef6Lp2/41Ea
6/ww1cEHg/9RsDcbUB5aHyoC0FSVkHf+s2zafy78jt1gRC+K0RKCc1NrRYltOvhdFpZHTWXiF72y
Izr3OLUHyimSnm0OELTwJYefgT2yevNF1XOtGvFguB469lff8+WbziSI4lhAJJopEkzGoCv/stqe
Fwnq7Ihkz31UhUUSzuy4oFHeI41Axe5R8SW2Xx3i/GkP6cB4I/RiYW6AXZqWXWMOnY0cWT/8Qj9I
mL0ekmpi9riix2JgaPQRQsUnC+t9yDTqattFDiUZrECxPCKywW8PU9JQ88aHN9GsVoc0gLJUif/y
wHS745pnV4d2vQTLdWSTT/QboM11hI9N5v1P1QPPw0slXbyIRDy9hskHMusfpkoc14q5jAKmFZiy
HjmKe0yklYD7XH9tRsgiANEHlPXRID6pX+efEBKhoF3BNYYAu/Ojlg72zQ4V0UrOdthQfIgVLyci
2T94483wC2Yuq1LdWBjb44bXhm0afmmg5m7KlJgAV+Ces5q2tBdU+YyKzr8R4/bOO3dJ7shXQsNj
TfWzZybacxNCRJM26sD7vz3cjM/70OlTAhg1GAgNT+IYzY3uU88N7sFWJtCg93XQaBTys14qjs3r
Suqh+kyvJ/dnUvLu+B2udiF0pyOPPMw+IxM07KtHanDgRf3lcmLCovIkGX3EKGrAk0fCINWjlnZn
/AAJ/Nwl5AVoABdGwRYL6rar1GxsHTxkDkg57/66V98dOaPzIc7P1aU2Dd/5GbB9iesoMvtqIlkY
lzSrlo360OApBjJr1laF+zbf4mGoI/hjGTRzkwqDd2LKtZqfeBePaWEMP7zjZVQD9PQ9WWSxFS9T
Xonu9+CdpkiTS9cKL+W99sIt1IPMuDcnzG/7ut6K40ulHTt8+es4OgI/Q9PMLDU8+wGCzmIHu/fU
ql3XULM8GYmh3L2tmrZacxzW1HxdQ5s0s1TJIQBRzq0np6YfnkSaXpI4FzsbC6Am1+Mt32K7qplq
agn7Jj2RB4N6FYl7GUf5yZ3dEqPqb1SW62qwZmshXHalPnfdaM2YlGOmep6jLsvFWP2x8hvxveLq
78IPVYFQnuoDoGZfmcMaMnSMPxiTW9VjVg4Nt1Z6d47q5qFpNang+jo8CRxgZRc+O84mX6xJzwqq
QjD4MgDoR5T8spnTTygos+leuo44cAwr4Cz9NtW9LZpSXEpsTxHyLXtrgP3+GZtx/inMQoFB7qUL
83O+KmvSoA13vuWnOQ3jIJ4b2eSM5Vb8EfdUUbdQBEl+cwNgR03v/v3OTOPsfcFYH7gfKp3q+v6b
ehhHtJlKs73Av/TWV8HDQ/1DHAPV4bKQctrrp1VblumxOkOBbxpKVRSJ9q6m0L3heownvkmu6ScK
7i2wnlXhVTtgTSc/1JfPdMoO0Bea5Q1sCj+ezOnQSgmLH3wq7q790MNyFeOaqOh29CN4YvNRvkX0
ZrXJiM/M2TJobtMpgpFQlTs0Xy1CpTa1lsdESPcpb3RJZm9mTMv2MDrL9Zq8aftuEE6cL4lT3Gbt
jl3XiM5WAGjuKfLimW7e7AGri0DeY6kdstFTyacRI8SPta8FxyUnGMH3ySVM3DDdRIvs+jGEWKAK
9r+67jVwdQSH3TVoOI3O8ZeNefDoXOS0RyeggZKoVaA1uPsHzSA/gcM9mZZUrf0fjeKIoPDlIA9T
RJpClVX4NC3nkYmCQ7AHy1TUInMQI7FciNpa2PKGM60jSL2VeQdWapjcYih1m6nFIimF7Gfs25Zh
ZG5/Te9qDqCioTJIcHuJbdIrUHFqJwO5fVW47o2Xbboo/bPf3TlFA+jWxaKQZ+OiT7dEaX7/WBYb
Epbxx+kVuOzvY/QdDMnSFJkZMPRlAyvCj8LJT6Vmok2dehICI4asstksoRb5EpWrAyDe5e1cyO5F
pRNWG2DErst1E6BtImmtQk4IpuzfjXQXloQP8Al0THUSVhEH4OTj+b1EWSAsi/y1RCXVw17YjdNF
77gY6mKgMrqBXHwtsy5G0Iy7vpqMJryVNXnAURjLSBQbc8JlqOmLUkvge820HQaiffhSXA9Orfg3
ydmGrGiSTODLPbGhTk/PKXQ+QgxpJnTq76ZR9g+tPEGcP3hr81mRfv6sisAgtRMtJhviI/mSKtkr
4WJwEVK+g+YV1UqvFkmj33tcSJtjaubgupju1r3mOQIJY+mfpYZHm5YB7I0C9luQgyiWUi9n1YWG
nLW3L+zN54kO0BXekDrEOo2PfKT7Gpx6iZHk5vB30bogNfyTQkW10zY8mreJ6n+C8/PZGhlQT1YO
KJGt8ve3MtTVi88HY/2S8a9WoFpp4Sy3BvDDDWLDs3U3i7+r6up6VRsafmE4AxdgXdpWixY9u48p
4DgtgDUB1q5R7hQ7Z1Zor4iTd37++f7PP8s+0gB0eGg8nls/aJ0K7rj1aG1PRE1k+zFWLZza73JB
isHndnPr4ClSsKYidV+ndZuYX7Big9b15XuQ0N4A9dNdYadawjAL6qAm+mlODIePvPJL3yHB2+0f
XlC4/FBOLhDfxVLsSxoGQxd2DzrkQKnrze+7uBJHr8QvKiEWVhN3B0Y8TMj32L9wW1nQ4gTQa8pR
WgoEu2CltlhIim9MNxW7phNNutIxmxAf5L6XJQxHLB+ojZFs6c6TRWlj6/1PmgDxMf2cwlGy6FRS
0OV/dNElyjQ0IMzYx4kqi4Ey6+umDuxSuigOxxRp6KJ7LUHTdTIh5Mw2YuxR+9vmYqzPNqC68d9K
v+/oYLG/IQfhN3Tib31aXQHLr1K5lAZFWGqSN5cuRGhqjY8YOFyPi/kQdtfj6Dwkh9KMO4gA/wnV
Jh81MlDumE7wGcJBvQiIUSiF1xQUujuf61zpbLBC65BSZnY/3ppVKGPBrK/vVujDEzW71dZpvc62
UtUUqm/x9sgJ3Z5T7XjDdlWgmKmDgQ6gBmnezYxbP5XvhF8+MWbCkZRiaSfgiBVECYFs7ItjaaxG
qFfmAQbP+QKWcM8tj37y7+wCd8vA3v9d0ZA/XKTa91crlIPGoVnvjjRjJQOS11hVYEsbZoawIQ8I
WWcvHUxBSUYqblrNZ0RnSLTtM3E6D3eZrOcqj9i26MY+P1lT7DcSPT379MFkSz1D8aThPeZV6BDs
vAUg0JAKVvmOLwHonWxKb/e4t4WDlM9RQNMhTC72VueODRdLDIBPry/umivEmDrV3Yje77P9t391
7nf7eys5NIgnTrnpxrArT3IuVbWjPnKKc8B4J287l8i03fmdVesiP+ffFV0qRwXXTAuffyy+zP8p
6HSze9/TbupTfIScG5uS+KnnDl0k47VN9Ety4xDvjNoiN3qShxNVS7HZiVKVz206LnA1XN1GK8eA
fUeyCbtDPhUWvgRwnQeGIw+u27terEZiDf5jKGbQdjYAThcXT9jfhfcrwJiW98IGsb4ofAm41fVb
qPThHwsufQLuGDfT7sdyUyYddWjBl1+CH0h5n68W4j+Rpxri74rKlIYrAdGRpKtupfikLUTdRaop
eprs0RZXM+/XgSV03bxfifqTG0jjET1YCzmx9cepcFviBC37KuLaHFOmPsbYBYuWwhl9Nmbxqzs5
3b5IKve1pB9ycptHkTwVq/WetJf3V+KLqJSu0VY2EYsgs/gz1Kw4dqAnWFs+R+InbNFpyDbpW60P
jCVsUqN1wrTZQ4q8q3hjQC9IdhJ/OGgBUi2WUh94yF6x58Nf4bp81uSSCLhYqPWA+eyOdKuNX6s5
h8FYzHkWUlN9cCs9QJfts+b4oiZvPnvByqRzC+gqQ7OmZ+xH9dy0gptpR5I+Dk0LB462kjEOSqQK
s1o0SRdEQ7oQHyZcW7q8Xh4jpWUQbFlRteZL/lDRK48+G1G/wHUJFteq7tXfOHDlqt0YFBBJqZag
RpQRh+ZD3nxrCGUb2BacIF4u9CcntrMp9fuE306p2cjLw2Hqm3GYdfkCr9f4tG82a4JWh2+zEDux
ckT4/g2AgWHp5CaY1leC9zJ/tQJybs8aUYh67DYHQHBLoMOaDp0Qk3St91Ky9m6EhuCRGF6SJyOJ
/R86WDzQCvAMgg77a/dsIk+JhqnjtrLMkD/89kxjB3PsYF+UHbMngn9UhgUcEEKCWw6/VxfI4NJR
s6CewxfBvu/Mc7gtIeRpfTkCWcNPEIdKdyVjO+EPJ7kBZr1zAPNQ1DQi3lWc2DVlOZ7GQtT7WVN4
3kiUCemofR0AXWfPJr92DuOkxXzTM3aXZKmpZLqTC8q6KdeRM9UkITZqs1Um38Q/g2O/dMFFlDLH
iQLwnHPVr7hcwaZH3iCqN1dX3N8wi1Bvu8wZ+sg7r7hRjvJPOO+Q8q+hIyNjDAEQo+buDzdtae3C
gEnRu2/8QY7XezhmaovGl5QkbxglsqigN46oDB/8fEKRL9Ivh7FHGOaEm3KMVBowUaZYh2Bv1vcJ
wmViwDAyg7FbCYdBSjUbCyAuZBu98y5dxRK4+BEDkWhWaUF1qrJYl0vCZTZpKNDL1PVe+kf824z0
zQtRZQA/j6F67p6vjxqPitgL7l54NSjynrL+T2i0rUy5/f56yKoxK6zlyZ+AI1rgQUMgdqYeu0Bt
4AzFi+nW5x+zsV/WQJQspLsj3yO8U45NEGK2jBJn9F1+waBKiSI4fK4BQbG7Tv8IrZoV7rWPJqg=
`protect end_protected
