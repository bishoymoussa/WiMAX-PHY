-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
o/si62S9miYlEYEVbCV6RoE5UUhQB4FXSGdvAGyYwLTBspJ3FgvIDYp/s7bEkyS+yDuzzjZMsX6R
onoQO5Y1uefCrdS2AsAVRek06U+nVcL2xB03M1ZX0SvToleMcQpUeHVjZWXMFYIwI9NUZLNTCqd0
PpR760IOZFsJjRgFkBDdGvtH7bnvQrqM6ApgtSKRrBorASSWj+8cFcrmcqgTaRFxmZ8Hd6xAx3tD
wW/jFHjlWCUwGZ4PwaAOgfyKWHOOigvlXEOk567/AOjI27hkhaTY4ofOhbghV3paLMyaa2cp/Rl4
i3iYVVNekHdN4DeexL2fhqc6f+XRuAU8ZC8eLQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 21168)
`protect data_block
gqMitRV0IRuJ1kX4dGn+eu6fCIcR/1riW4zF2NnFDhIoonGk7FKiLH89sY5mowUZL+SZn04Gl0K6
ntZS5fI4rpN6nwG0rK+prYfsGvcihtAcOelobKlvWu4vGLG7u1GzFpQA4Qnm3orMaUEHBCnyC8Ep
lzSy3WR462IUC8UQ64kahoUqdjNN/f+Rr27r8+t1v8sB+L6xIG5Dvr2h7RJWk6LAn8FBf48sfhSp
0cDoFd/Oc28kelsBKRIDEOzwtRGHQoqOXjNnO9P5uAN47K3jpBxpwjxGSypR8We4sHjYkAC5iJ5e
+onvdEoxnMzZ3GsylCTX/l4T2syZb2vjLgi1xSNSD/Awv05efjeOiNey5Zh44Bi/3iR2+9pCkM5H
4WpLaClpKQNOXcnbTWSCuO62/a5GuCyvlQ25Yje6MqbMa0eg263hB5mQocbcMYCuNNfXpOUe3rV6
TFNeo3SXw5DTk9m96HUOQyJ5/EapiuBf/juiC4NXZd0Xbcla5OT/C4i+Ok33LJHQUdSGvP46WJaE
hPcmnSJRQ1VJg62qZ3H5WhswVknXahVdf4yP8hND+78aQoaU5/NxfI0F8TmGKWgZmynzTTpG+GuK
p2WKUYeQlOwlLAFhaI5SP66F7JCUhKDtyfAkwxdubziGwBA2a2E+4x0X7wbq7s+hsGZU0dEojniL
nosInnw/px4JOCtWc3Z/mJ50e2i7NYQYr0PuAyRryqA0jGm9gr0/AAmfMVf+QQThMTfl0pYZXWh2
NsVJi4IsOwX8BO4f7je7tbkufZsTCifB+TnghrLl6+Of5Ci4ou+4eYlY+FQRKacn8wYVpw5ZeHZ6
vYgPjsMSykYD8uJrG6wnxB2JrpJw++WLSdm3mdq979euWFs8+GlBIjORUwUmCZbPWk7VrrBmnbYR
shH5w1ZrntuCYUjrIOoXRH/5+hJYTcHzx9DveP70CKrUBfEZF1rHUdLyZbLRpY7I6wOCNBVWGNBa
CnTQnP8I2HhSm+0Z7njUVebl5hgPdZqTjuRAapbug7s78DXzIZ1WC45FUQTUPdQ7qeti1HpcYp2S
MCtYNL/+Pg6Oa75LcNbiLKDCWbVFhLGoUjeleCk91SFq0GTwUCDVQUl9sD8+oppgvGsSHiaPHT8R
Uk35a6oH1exM5KfTYqXjGw651cqiZTLqr8GVVRSSi2cDDi/fGiSb+BOTZv8ZKJmfsULt5MTvl9eR
jBFg5BhlPOGPHPVvZBi+LF8QsTQ1XZrKJSsJuXjcQbeQGOYxQ27gk/BFjgzbgXNr0G0lsw1gnAWT
dvJ5aF4K6/EUxcii/bS+iWvd6Pc3ai/s7x/DIcofS77OjNE5V9NIc0bwrjHuc7nQxbOT+pJNMmsT
fh7KEaBm9oKDHxDxLyD+/MGDCuj6mN62jEkmc07bqzHmPcdRdI5a4QJq5Uckg9veqaGy2T0WJRfB
iLllgNDJX4xMIqJiyrk1g8Ne6efl1y0RT1K7IkQUje35dMOG5NFsTrt+y7eZQXZjRWHZVJn3vAnH
IA1rwRX1zSs5z+RH/xqoSmuq0ICNQgxmY5P2IcUrG6/r1+QS7pcO+sH6lniHdWme/9urvPHfVLne
qduRlWr8vpqm1hGDPWvHV9kr9Vksjb9UNKsXxPzqa8SD3WxwGAG3lSwYuiCa2w1w1Oatd5ms8Dh7
2M8IyeFl9aCrZlg1G2XBjun6+ZRV0wXpin0/nEigQTki2crQrY7RU7U2/NM5AjLAIizxVZn4VDgE
6cOTq2OHEtPrwF41jz/9EsWxzakhBNLHagnAs9AS1Cb5YtdhYWm9PKcfKnGWDOdzSfDt3f6mw2Su
8jkJldKCYNPDUd+QTZTKBq57lZ+uYK4oLBZbWbcpWW3rQOZwhsjyZwFd5MyE1/APCDKi7T44clvb
+ljIBwh+EFvMoDEzuWVfCZE/5rmgmfqQBO7EfKGgbEeT/hN0TVAP+mN4967YyVl1KyQQBr7y00VE
fp6j63GMJF3zvmjjwgRdl8fTVgswthmtT+x2Lz6KiSAMA4Jcl2ybXedRXAma9o9EUYd/+b5C1f1j
+gk3YX56VdJOxt1+lXCsO8iGO18aCfhT+ol1nrfinerotu+a9aIFyfHBDO9Eyg/JXXkr0OUa3/ni
OS6il1s9pfkwwPJEKZxwIFtF98kMRyUhGfqAM0OuTuaf+3lzpXk3/Q1/g2HBNCkoFOR859tY/Nq5
fZoIA5WJPMfrnnHCPq3C5booBrnc3+bt3ZJtdGAuu2XrcoPqE7PQ7RK4R3eGwBqAQEpGXrGuAIPp
gM6+40wWCnt8CCE1wL17BmkwFSrlhbW7S2/2pzFMHzIzX4j20r0qzt3mytfwitb+sLj3vRZUmhNR
4QwORI+qtYfQ1D+jf3XPyLVSFODf28stH3uya9W1CQ/aTpAluBXQirN3K1fjqxzgzW11H1OJaME/
q72VbBjsVOKULjxO7m+8Yaz2iu3M9pmj3bsgWf7fSW1CTwcfOS4xRHJhquXiRifswZETwJc381Kn
Tx2ik8zJg122hmNjNsOYh8S3721XMVJZIATkVBXLbAXAIqlaj/H1bX3CWlvCcGKLgFitGmlTHWZL
0+gV+bSEZvNQLnVFK5/ndVu/AKQngVXuxo8XPkTYpHERkNvdLbOLYF+WlMkak/DAJEucqreAMKwx
gT8y/i0AOl8tDrvDt+vgzyMZUiJe30wSaSn6VtZvBm+a32A9YmasASPA3sTmr/cLaxQtJojX6Lw1
2/yMg96HN73Ab/R63nrnpAusplr/f3adQDcqctJv7VCOKtOaIt9W4WGwtlIAfVSzMB6dL2OvXyW4
cXlid84rYtHepvsUVKv2l1dhUcbsJBw3wnQJgZHpkqehFYwiTtgh18KEA5QBp9M785ozxA5dxJN+
Aqm1if2gV69w4PW64VdDNL4Kb5fhjtHkmcSeHNU9fNSIAefBHnO6hes0L5Zd6zkVnO4luL+ajs5e
QHxTgtBvZJ9yf6fszGKi2HEoYOqNy3EVzbFQ0uA9x6X/63e2xcs1pGmf9N9AuQC1Y6ZbrRI3oxtU
miH5w2Pp6al3yzUf+FYrGL0NoY++Gyh2nd9KrRzGTZD9F04LKlu2DMiVxv5UETQ4jUW275j13md+
fEWeTjIUJiCkv3lAPdI+AfhhR/f4xmope+PuLdeAhj/oxM27WQQ7x1daCrw+qTkE22MMYZcTEF2+
3cA7Z58G9HEWEqYqWvlcBkZtt38mY0+48x9KEmMSum4TIIwTNRaUzegjhPHCelhM7aCicZ8xa5Kr
2Uyztz0QAHtya6r05AZHR+NfRR5BfYaViiLIUrOJ73RvarKUq3Xzzs659b265FJtvQPu6OsfXLmf
LG2qj7UmzfhnsXQMxczTKEcmbdy4hsZ0ozdIuiyKmSQ/30ea30pD5r16+z58ibX/K9OhEpdRSlI6
71kCFEsmdZhz0/lE687eQh7KcXIOgSHjlOLazWmcsgSX3Gpxbgx1hIaC3I5uIej0BgiFmsIQ65qk
emjGeZ6kBT1/hP6gzHjL2JuHNr+D7GFwcNS2ETJAKj5NXqKT0Ewx8l1FeeL0j0Na8xUo0M2s9c44
pfHxVrCRqmv7s+KyXLH3Eh4kDzeyVNeJCDkEUisylw62cXWjngGvXYWABOnOcsIHEs15bhlbl1lf
IytF7Z4xQIk+aCJSj+Wo+VuI/mlp92JMCgHHw4BMmd6Y++yLaVgLXH09oXFPh3TQlnGMkVwc6oSp
K7bK5pwAOKyH3YwXiUX9OakRJ2O2ihqdePPLy/kJOWZ+ihoKJNXm6pW+g6+YOoCkd47SQ4CvN5nz
164IfE1fDaqEbjg07mKf+BkI9Lf5DOZwVFeAJ8gC9EBxECQwUAZHNjURD557PsmUg5eBOpDamXeA
ul8DMJp26d2/gFR3bQURRLkdu4Jugw6L4czoBwA46Znq/kqDgo6sgV6EMSucVp6/4Z9II9quFnOo
1M7RmVjCzzVTGcRNS1kNvhr3frNtuMIcNhLQeb1+EFe/NYPi+DrjS68fYCZ1x9vtmI848CKm1vJX
Y2slX4NyRh1F0kC8evraURElkVkSddPGDQUV34voF6FvR4tNXCay2IBS1Gfcw/IK07CsLKAorHFm
b/1x8mUE++BdYMgqo2La4OE9PCCj0ts9jZk12Z1a+SVmuXAgwsU0a/xeVaZzR6ui6EmY95l+ZO7X
BwJJLjTCR99vI6eaFfS2a7pd4zT1hlqdF3JgEZWjTIHVOPg29ACS0wU70avqQUr9oDVvn3Et869h
HhOvQAPdbu+6I/uzmaT9YUcdpRKEXIvUUOrCBHOaMDVJop9sVHvgFdCJuyJhqcM+bmgIUsVxAExk
4VeCilw5XjMLLoaGJrVXKvpcgYVmaG+5qiPY0pZcrYAPdb8pS2c30dV6gQIJXcpotKRb94X3O1hw
dtb9fILkXVvzLAe2jljZpSryZ8nA4AsdMJwocPJP7kYMdD0n2A4wkqunrubpCw1H7EuYsdliAx6f
NcwSPbKqLqZe8XJxK1VzLlDPlmDbvztNEtkH35hDCk6IAJE26o+LL6/a/ypRXofXfTJz7c/7QTUg
cjTjiEJpANC2elAO+V7oCikGCpUKhFpsqEAYOv7P2hbqmuCvW40Xk2Fp7FR1WB0LGgyyQK+h7DZ6
4iJlJYy0D+DouZ5VAsAb0wUpPT2dzk9aPig/1IlvenLQuLswxKMTqk2Fqnd6xJXQAz7BdKrWdu9B
HqtotVpvc4UNfmBgqUG0H6cGGrVxsgi7QWO0+d8RrI43yxvBNQsCLingMhsE2mvaYN4Ahn6jwPkP
dV8wcLpt0CAja/0ipQ4bpFhGrkME6SYpuq67OYMU612FBwqjH1stPiRfYnvY0gb8sN7oWDV97En7
4WRwCzmstf8QfuWKX5nobGtFCM1Wxb8RiaooHIYA89ubFIsEKPY6ltxi0GyCdx0Rii6kDTd5KLuj
Luk1Yjs3tN+QqJsKfClpYOus1kNBFfdp6e9BrUPS5Cq71pMGwTiy+qPf/kYIJWPzvg7iYluB7vvP
N5P8l4kkiH4icaMbYaa9bj9ChZwXCJsJscdV17pcrsmOxFeBSQeAy9x1LP0ARS+QhhaSxzz6E+/n
mcWli1f0ArbtD3Mw2CuiSwm+icCMeIsqBa7138IoSO/g6XkcibGgwz4knYTNx688Gm4b/YUtJzij
RUQVgXLEuAi34kTxqfs9p+gImKoJpVZjv80NhMy/2UfuDdlpWB8DF0ZtCyK52ffMSn14TUiVFbtW
KQda17xU7nJ3lwKi6xZW32R0GPlpdq4N5mwnVKgwWIzI0wP078P8WFMGggJVQ6BPp2lrrIVE0b5O
O6ZhJuv8Nq65xJwHfUZJBqlcNuw6Gt31EJONOMzlKDL4gc01rUHjyIIAsW2JC9ayVzhNr3cabePH
CTtoWNqpCuQMErRS0SUQKRAuqfj71FOER4/zJb1Zx+L5LOrmhCmOp7pNvRGdGL+GPnqmkf6QfL0b
VaRCWhZtx8AG1CehMKqN4XhXKorSSiS1GEoACe8pxH/h+Rlko7iTX1ZvcUEBiPpJC7bXIf5X2IfE
VIpuoPyFsRqrUauaD7TDv3q+7HZFp1mi+jd2XU1Z05YskplN9czafoOpLmJuXxqEaoLTlw4F7pkU
+/pNsdsceNPfY1ZsnoRrhqb1G+fcZsuKrEGP/oNULVvSfk9NhAkZKysrPTTB/2q3xWjxxeeknpHH
Zo535dIfKw94TIRfD5BkgK4rC0oWSUEDZlAdvWq44RlncivA/D7b1VDDO8OIA3J1EFo0Rqkagki0
L4xwzYVSJKk8orDDglP01mNJDP+zSwPtIyPdx6ZR5JatOuaLIwXnAnY2W6YL1nqijMmYCJhdnLKx
BTA9KVzEaquwf2bntjccXDA/1b80ALwrPD+6QdvnjbERl50e1mQ2Y0+Ohj5/YUqSYhvNctm4O9mn
zKZec8XiHVwNVbMTeloICggyxQdVPLULeYCsJYlJQTs7MDFw3R62y+buged8aYT7z3onD3lEcc6f
lbPlZL17CtxYgtYsDMS5VfX39IVlyIfsZUvMnp9kESCrCXQDgY0W7q6Xh465cq6Mwp7NeEchDwrz
qkTdCwROodCrbGcJIDpisvvVPnxU96D8Mp71seqAzcRK+wiMtDVXfXSY1gCbe0FD3fFCMWAqZ319
DpGZmC8aLlqjuKd6JzCD0HTpzTFf9ntuY1cTbbNl43P2x723vhLPCzbQ6aNV5ebikzWMem51jM7r
cwFQxkXm5bYSHRERLA6z0mU8qi9cWti6PUM+yEu5ckyIMz4zJpjT5CBQeqw26NMh+6/hgsebEOih
EbHi0zo47i5aKTcgTAWGABMOWDj2g8AUOco5EHOBz7m0RUZkcP8kQktTitjDXsfJC3+xW64qaWIl
9ykX3FzHwNS2Y+VnZR1pFmbX4sz2oEIGggeV0ZDReI1UgeGrSn2dQGl0ajwWqaQo1seXtCQ/gKyQ
jPtSEr04XsxgFAGIfblSW8PG30uj19tmHy8z1E2r9BbwrZk7Ox0waoMaESEi5M2vnXN9dab4nyGy
EXezdQ+1wIa7IiRlKfzpZt2WoDGqMo3t/yM2Ow5AVy98FzBbiUS9LmXfVU8O11eKaOjeyBeYKrjO
nUBx9Q90q75h/Auf8rb0LVuM6MS/7xebQqPYlVPpFu0NpaU/eEPTgJlh5UDgb4FwMxaRgnGeCpD5
KDLN0B8IhpN5HZyxByhixnT0lZDShwOhHtRQ1ksNBKhKQo+3TUIBhsTIfBGy1Pchd29yv5XO6py7
MW5xM6h2CMIjHIaIoCsr5xV4MCwJvNaa9U01CEMz4kPZzJaV0NdHL3hy1hONhZIBXj6asS+nSNnl
e/rpdvWG/z7qfPCnqRcq04ly3TDM6UUi5BGQbJhLEN3vtk/1D9SRS3Q6yaDwRdjNai58yax1aUk5
w01f/+oBhiZk1A+19CImb/2u8fdA3fnhZ6zy+cEM/Ngb9HBIe/yNgYF6w1hS+Nh8H679RZ9pkyyk
7kNwbq2h4p2Nxr1dj6bDHr+8GOpK/kZXvFjSh0JO9n2gK/5v5sWLe0IJV4vgz7TkmfDibB84z5XE
29n71fhPJwRmMCNnCBgjXesTBrV55cXFwusomjxJOMIYkZOSiyGK6SW6+tX4QKqT+OCh/aG8PZHi
u5oR7a+1+BO5397P/uzoM+u1lFDP/TQB56yG2JXyR2xjY49f5MEzGIgvCaddNSP3+XIXBgYcXtcy
fT6i2khxqRzqaTS/Rc0eVMKh67JeV1FdTA665RoH++pvVYwA77fnhWgRzZO+nYj+YJI0VKQdMugl
iUVfFHo8adrkGfknWIqHff8a3jqmO93oPxUkeC0AbLaLaU4InHBZAYaczrPmmk33r2BM17cEfKtv
+F3sD8KxO6emPQyUjiiGawETbioNqIWJ1iIo9N/zgOsBgbLevGBNXRHi2Y5dvd6VayyQ7uRlf49o
w+/WQM2jUEpDwFPOEIehOz9Hm3GpWuw/Bdsi2q5BPqsWvBwdoNruCNcS/eA7JP0NHymtveaNTlu4
LIqeRN6Z+5CuP7aYFzMTfmgj1/l3aW+bPjHmEIpreMnk6BRe7YpVfQ7x4+/3TIr90g7UQ3Axl4DW
zzkyL9eT1JhA2oFqTl8WMfKOJLms6ki5TdAY+9rhjOcIT5m5FlrUzxKaLgha5n7jQZbzpCvRtw8D
nEToaijiegrJ7Z1x+u7HqKjpdrcEUiyfE7AO+V1Bi1LHCNpP1ebjALhO+BnD9Uw+0SuvQYMZ0SwW
MOCj3ergQBy5wxAauPdq07uU3kiphniGYVVoBEms1K7aVWCdRQ+E4NUSlzB+aZ3DAeQFz9+Kg2fX
QRKFveXSysIrAcsyXpQlRV/sLNvRRobM+M/y6fz3POYTY0qX4P6Sd/xAC/iHrRpv1uzD/7FkVDjS
OOG52dSHPhAunx/HeVioyKCT9fRxCw1a9TSdqzA1zRhcRPHNwdSUeWy/aZwD4lMAtZ5K5qDU0fDV
m71ypk0nlOml8BpMNzGsQxgeVGGuLnPnlBzzHsqTjZ2NkyoO6JZ2bcbPiDDD/YGYHNZA6pF4xYYC
BK8XA+7/LGbFVLGrnWYPrcqOFQwBUaOwNXLsrNFZSopxaw/+Z/06RoLDW2fX7THrhsWqUwqqh//9
2f2/532VcQ6yFSmVFBH60Rsa5sVD0DrXr5LkyyYXgwC6eo0kYmPbQqZ8ZDNH3JcbkE81IYvop7nY
k6iGT/9ZXbOzWS5VtHuEOiJgj41Kr29NXMRcXA9RaUOCaDpgZNo5CYQGz1xSn9UwGwAJc1Vj/Qy3
RW0RxyO2G7PkITsfTE4hxDDhrtyM0kePvdiT2qRs3h0s34FVbbE+EGgh+2pSPs76PtfYv6hNRey0
bMaCzEE9GD9ztwC9ZC6fI6bKSuNVoPlJBuZOEppvl0cFu1GXaEm7MWkGYu6REhqb8tKjdYiIAbQZ
6LQtltniMl5N4wvXu1kID0DoFfBi9KDpGmLHS5biwy9XP6OT0W6JgczqHc++R3iSCei5rNH57Y0g
S1GeBgELn8JqQVrlPVhpUAzMYrrMgEidWaQaZiw4lr3+9wrAl+DhBfADh9yJccWZUDGMnxkB9wO0
UAtoaEVgvXer50U5YKhzv6XhANAw405xjSLUWBRsuC4hhfBHxKNEXjVkHYLPYxwGRoGPLT6CbUTi
o3CLoq6eAqZUMO37HPXWP302WjZxQ/iHEU2tavVr1oN7I6TdY1Pm1HiuUvScP+fHOCLm84DJFQ3f
OVa3y/yAgis5YO+HeNEzimQA8G7BtzY+0XdAUW4x01yfx4gx1JaFTRo0U7EOs4fSKvvEDxWDO6i5
LBdfKzM9eXYCIGhNBPo0jpG75hUE/4T4isbGWEoQ3RoGJ4Pg8sFqw2kT5yCVYl7evGuDNnYR1meB
BXAbxyMrw3/G/m1hbLHQ1oDAHgIXKdpisR45YUzW1CZpnBjCC0wg+goDVlh23/Pz3vjNmmWosR+h
yMDT7V0HCMmGwwPE38KBvlC0ST888URa4hAA1pk6rWglWvlR3TfkZ56pty6xjmZjYhu4CbL461RO
Msv8woQIc+SjQY3IrV/8ol8428Y8WMSpF5U9si7uXPUmSU+WfSb4KskmaLUOk5kiJFQgxgNdJjxw
sFcDgR9kjvtN4H4GP/0bsv+ok7vpg/6alG0XYAiCpHkCYIZnE1syBypvwDB4FhfN/6tP13oJunTL
ugMfavcekjYg0tZeW0IuLrQ38P1bg3dq8dzpRHxreYJ1aK+18cwZVsE4gAaiw/wXTjye6unXv6j3
+FDuhKDOw6JpGnY65LGvJpApflD+5jleAn0G+ZaBCESENFb2bdUiqJWGF80s/Mz6+0TdkL4uK/tc
36cITA+B0m8ic+fCEXK/ziB2/+tyiXxhtUDJxCOfep1pRG/VaxsC5REG9uSX3Mvs0xJvr+dYHLHf
n5PEOgrz0v/dHjvbwOFyM1Rp/vCzu02AqCmjZ0nSnV5PNYaQYf37ytI34c5Cv2ihLn4Wao9WSTf4
s7sTWQXaKiGfP8I9FhJmJ+PJPffAe428Ad1H6LbDNQxaDR2A5HmxqHByjiMNTZj0OV6NnF/wSGtQ
BHgH6ORXIxAg2mVT7WtCDp773XERaJN9ZjNyQARvDN2ezuHtR9mD2TTUlwVeJi7FeCIN2+Kizo+w
Q+xsH1q6T/gHRJZNd1XQtFsUdL860UeuDuU5hIsj8xfSLhPpppZWO/8WNQK9xFhcaybKhZuQJGVx
e7M3OuJD5KP1M1fIBYYWjgYomJB8pihHtFDO4jsRfylldXtveAeyew5hzpuh+GLKHHQLxhDb36W3
FJhW6jKTZWQduwCP/bZlIEVVSPv6hZPxjaEfI1hUN0f+N9lpPL6Wfjk51kLUUi6rn1CxMIs3DWQ8
LK0XvpExLDpnFW7+yPcA5YgQ1OtQj9fqrFWM8I30Dm5JVQdj0B6CuU83CZ+TudGlJ3yofHppvqYi
I+H3CNSCikt1gvtzflcULjKI4MLz8HSZOmQFxXPpVOVcvoBN4e/Ri85fy2LUkn05hL4JDZzLyqUx
SlcKb066dzyS3mRwtZ9CXsUFb5dtdPdOpe4IevvaQnVl2JHiPmDoOIpmuwx9aK9Fd5Vy66eEQowp
WZH5eZB3IeDSDiUXpPER/yehbk8iHUsJSmSJhZYRmKVfWyQIABWJ8aSws68X//ZfBTu72ZzGXGJR
ssrzaTUDWvC1kJTNuSm7E2W8yYc3YHWv9icVlrKfpjniJXbpr6Qwr0wJT394MOMQIHxL7XVXeFT2
FgMK/nVZAu08gfDHJu1la6rkVocu0UJy7rN2wAItx/wMWVck2QoXlnxbiBxEko/S9qwWn1sAcVMr
sKZmEZie/4/EEpk4j5pOEApNRZNFsme1v4HPmx1sPWXThksLB6EN4GKBPqtZvdLTjXxMfcEuMH4l
BCNzxejJ/0a2K2pOBjyKaIZk6SZ1JROQhFZvjqDMJ3Nzo4eoDHcUdeFlE1U2hTYxDp3EslQz2eNS
awuDtCR1w/efOD3IvCFAC1tPAegglNSryF0s/XjGUSk7ag2uQ9o87GAPoydNd4ranLXvwc4Aztsg
0MOzASd0ulTXQ39VhS1DdUQlTLfm1o6chbHAqoXjuv0qjX0kM5LE/FTj0r+PiGIKKMX7g7lgYCuw
VLHC03OA7v/gxUAfI1d9IZQY4+SwAdZHp8VbtPAgIxqgWgaZgO8/DQubp5/eeM8p+lF2nbts3UtB
1Ri8UfvDlyjbpDCp46qy9LHaU7IITdZFsP1FS9fUVHuKLDbzQT0f2flU0YFfnI4OqOIOP5Ckd4Bx
74eXWyVpPwVmeHaJazqk0QtzPcXP70ECicW0qczjyjkFe17eGb9a3d4DOrlXclhEGeRKgGYCB6+X
IXeZKIcz84xnPZJ9SWmRdQVnbHjkHatLE2scomxuI0y0mozkUrRLFtNsD2IU/aKEd6S0kssO69Ia
U6qu8eM5IjnSLs/YM/0chs/qOYzuunaTH5a5WGF/LsWh1VvI8X4W2vKm15Sq9qp0e64HhTx2hZJE
g+SzW1MfbRfUx7SjYYvqT/v1UB+aXDTPoXlTH5v9KRD/aZJprqDV8GEEKCuVx82BkfUAToS3HYBk
iCB52VP9e0z/UzJ6TAp9IEDJo4EHsjWmPjSq7dXjDctwsaw4QVeJZoi8wtQjlD8vN6n5qBzqA0rd
8Uql8FeLo80gEoy2DnqKIIOQSSNACeN4KsqRBnb293QdzftWQj4ckE2RLGbkSUeBV43TPe/oyuXc
JbJImQdMlQtrdOEKw1lwiih7FFtMsds74ZNEhpOX+ZhNRjP6dR2GcpIzeZy+re0LhPH93uNQxbkn
oVTEvCcHLpeqD8zMS2S6FQ43oBze+EnVWytoNU80ZxwMq1skq5jiPZIuc7KVZ+6lTdRUzTwveKwj
yCZIw1gQNfxtRdeHEjvjVKPkYf9QIcDBdUuM5F2F6woSaJyRg9Lm1kgk9RRpf38NBhwKAY9z2FOz
XMXlDcBCiJt9uE9D2UnFI6Y8dsuLbXedrtnb9V8jmx/ugwWhk5J4lXP/jBHHpL8jB2AQE3XjDR6H
vqGybS/G9nI7ZU18ugSurIbdXd//7bMDlAoe2CNRNAfStry7o3IEtsXCbna3SAjP1NcpenbyZMxE
hSWYwQz8XSczSPpnu7mUiipbPzDAZ1UzIglDXmu9IEUoVZrGeRGr7hfPTnziFa5jZrkTKG+mQxRd
LYNUIJHjGD7UPxvI3C6IPxNR08sbD2HuI+Ot5qAGSCbQo07vCs4fZP1i2KqrLaX2ROofOk+K+MGe
GnopTYyHuT6PSGYXo8RWklI5hsB9w3s4P8E3QD6Ogump7lcUp8qAkidYpXyYB8OG7XnZfYWKXrQW
Q8+FfmG/XD08yaFs235BTWmsP6YgQH7JdrNO8R3oJL27NdsVg+oIJu485euRdnUafrWUyn/B0Hm9
LWTG48gVD7zSXtbCwncrobKhGTx7DJu8MY0z2U7U6+xAaSFiev0KmjuYDKyR2ceEG/YbCUOl4QgP
h4mt/PaTvv6TfLsfDbm0AO8CgzEv7xvOGrO1nPjAdLrkkDmSdItEY/NxV1XsvaPqzS95IYgjaV8h
uHHi5OgXR9lnM1Kpfh8LEkVziWltiQcEDai28ATp55200zv2RjsQ4+irmhRidDfYtLZbVRse42ab
L4Of9rO+kd0AO/Z+LYy+xctS43aO5XtTRHEWQoQZLHgFoei0291qydUhHcCrvpnOFyPVFObgsb6A
HfsfVsYRG2AQLCwEYp20udGorcmfBnGdIUKgJj0tx6kiddFaB9rWCSmdJaU2dz6o6RqVTdVitdTy
uTCWh4I/CyqjjIpGhDt4yjqqsu0NkSujAF/v8KtRVSRbq6r67yn5TAp3eelvabnQ7xKvSiiC0X66
iZP9kwgeSOfmYPb243DbUt7gz0jq2CDJ8ZVduIUQ1ekezvUqMzo/Bbq5ZXSyLxb0jl7CXvTkg3LG
DmOAPKUEMqanGLv2W4zqVI9bLBw8jBqCOhE8aVVf1HZAD4ZkDhl1IvMLKE4bkbbIqMY5voDv6sLu
gLtJAEFTHA/d5IweLRvUDuu3jGvrAdPXzD9QLbZh/NL9PGlUspu6QkPOChhZlTPHXbn2yIw+mQu+
qOWzYZJe5RlamGfwm7cjwxhj2j1XjNO0Ux+Eav0rI+WeJSVFsnPkdwzzF759cctJOrNPRcgu8ole
zwJs+VadVigiynahLTJGua08pqQJVSiW+/fc7a/CU7WY8HO2r/28q8QHbmsJPbspYoh9DZlJQtXi
lbmSD+aA2/vhaqgeqeL/f5ZJB+RDdBWJEKh6Tz7TimiVoqcqBcwDZj/kbXWKsZVKXNFmrud644qB
7U8JD4wiERA+4O7auutrriR2NuSInzCHasLG1ycUGzETXJ4okIBAJ0AOvOJg3LWXJSrn2/iIUmao
V2WY495QGK8RdnLi3O2GqWnFLKTtRI3gVjlXx4K+tbRv4LX8+nl+H2164wWP8hyzqh8/Ur7zQ/Ga
b3x9LxupYXaeS8EPNr5Nfp1aBydkPPQWviyBoLhv0k73qFGRE+TKSUXWswURY7H1wLbws6rRJvu9
cEKGvy0OX5Tk7a3X8/dnzvH+3rzOc/U8+xsDDRqHSJ+5ZHkWardFF+W0h/SoG37DIVwFej5qnYDx
ywfIZlOwEmOirET5chqaF0kvrwdHj16cGJHmFabBWKCL4yGfBhrtsmvamzvxIWjdyanLIXffs3M4
dN6pkBqJXD1fAHehlrhy3RzusOPiPBCzhaUZMl4C1e+nIsHxstu+IylTGADt7IW91ZEQmEQ9QWWG
ta0l2pB6dfMTgo5dfxHb73gmWTPh0Ao8ViK5cA1LUqZ1Xiq/n1To7ZN6kmZGABREj6258J7ZdAs7
rpN6KN/G/M7LKORBWiPe4wSA7ZJf22UIkpZwapBjr8EG12TsPHiubudJiv0A4GSKyGRsfzJFJpuF
l7VJe72yu1P7xQlUtmQmVo4DYMNH+PZR/Q9s0izESRZ4WpROtVb92xRJdf3aZel757U7r+3gmRRP
o93RRIdu5qnf9BaFJr78Zv3dDE8EwyydtpVC6VcC52TRPaA36tW8Yw8ywwWHV33Ue554PKpUvjBz
St08XVeRzF1DEmmZA+vIeBzfK7JPRXDryUfauD+Jqj5qbej594uQOTCoHZmQBlA87kppaWUGTcB8
nDwZJKCZ45T8RRmR0uMa7PZQfR/JmdShLLEg01iS890n0FC8niqzxrBDPhXNbqeDDzzMdyPqkZ4J
oL8fLBjlQ+8zOCDNmCJuI7igX7SdYrYuLfXByHm3qQAXAJQrA73L023gjYTXp/AXTBOpeKob0fqq
EbPFjtQEOnTL7erQtrsDc1G3NbhO16Ezc8gxozR/B/0WsIGy+72lRgmEusSwZP8rRpLj8H+6MHu5
3FGVcGGt4Qx7aU6lLgbko8aOCqtyJLYXYLhFGgDfnemVQ/iNCaM2LDghju9BUbPbYgpASROjHuTu
nDYpToiFpJNAJW/+fl81OtnLpgBmjuLOvSv0cAbBe2dFaMtCVZ8PSyPVxDMNqEHAWfRnsnqhcEYZ
8lE3d+tSlj1AZ26Sv6BMQvt0bdHSTEqY6a4bJCjrxJCiX9ndOK/VPaIhcOnNtDPckSH2z86gbeYu
AunNQ9mlAWqk2LuzMbQGwkXRm9bikllrAgklBHsew6K+vzL5wpBbB1uZEiBHEpr0IPqYD16h8NEM
lGxMXEm2KQz8CC8fPNuOUoVGU8cTOZtQjg+octVl0ulHxVDe1G5xBuDwIEdtyKQtP8QEfQ0GNvyP
OK/BtSnxNNgrdLeKo6ljTMa3xTwG2gtOCjUKKlyi/f//QlxjGwi2XNxJ4Tta5NjuyWvQNXl3P8hd
fNtmB7Yq9wbUxYnlWT3QwgFeWc0EDldnBC9o15MnDx+TLV6aPKknLG5AA2JYMVWKO8LOjdd4B+iF
waNNzjhjYre/lVc4KXLOrAE4sz+YFtK0IKezwsxi50CcQ0gnQlHHCRX3fgv+kSSwvF04hlOn6eJQ
+cb6BzuMwYKcy7Xovgc2rkG0n2m7jmvpWgwSrLGc1ug3s/zjQd5aaTulioFue0FD9ioGNXzHs5UY
bUYm/l9/yKTCYNyyweU1V6C9DZQHS1xMq2B7ZPSchUosx4agp9+6rGKP1u1sneSR2fViGtuqVw9p
0MZraOKQv4Q+0nBVeExnt8wN+TPhdyXALJXR6rJkk+CWVDZMDUYXzyLglc2IKsylZymhPxm2sfQu
4ADezeCBfqOd63Yp37ukz4E8QYV6e5bET3XnkwgG+15O3yfB2F3ewNjbRIqg0RVZoNIF21lQtVNS
SWYJhDhyoY2MXgsQIbHW7PRoEwR0NzkZB8bEI0qb0TCTLcS6NgudnI/phKPIN7nfftPkNiV2sCAM
fkVMmjCKKBM4hnebfRCVNHIDXTFw8McR2OdzFvM628DMw90ouRDCmFW93KnBvKltAF4UMsimkfHL
R8k6g7tj8UJ524m474ITrE7vef4CyyFnqrUpAyzH7m1u51opQKZrucRHzVqtRih+Pw8+JbEA5I6V
ZbJQVZPqPF0jeZ02QO9jbH4hsnj0ET7TJGWzzIowl0OUdiW6IQruLw3DIzNYcvqKsekfk6YJM55j
Rd/pzlmZysLPjyrKPkr0fZ2WxtyDR9Voi1svQgMzdZTL04qwh4PrAg7y+MsOl/xOjgXc2I7Q/k+2
0ySfpCmqqwOChzBOZMBnfHArITgNumaqTxNpzRVW3ONJlnOyzUYs76zzv/UMaEKQlNsQUSrzhoYg
36T2ETjVKe24nyRkeXSsp12YZJU8wn0ZG+BS2RX/4QwbD1CdDdTiwkheH2RiUoBx1HpsrUvrHheq
eXJsjepJgBmNRF9EuQE+NuHaN8wBjnh60YYaszFywYezCluSmIEyAnSEMKQY4tE7UffWA0l/RsEn
GcQ5VXw9G8/l/h1rITzg6CTOAfYKgqx9JSRBLqOE6YDrikzveDWbIgWsnFx1/nyZijFKWiflN7AT
LFU6xr7N9v2pOF6ZpkewwQLcLL1IOPS/o72mXv4mDfmd+N7/PthY6QQYap6cAwUCoMH4FAXl9T47
nccAebRWHFE2EBwnCkxrQ4vyGF7Hh/RDbmOFglo6bMwIQMDw15YmnpoUmDED4ef+c57XPSaXM+dp
2VxRI25ZlrXp80tcR9A/qPf/EgT7JdEcVA4v5wpso4stOOshMQlE/ZngVv4VJQfLeRI3aSWTsHJR
0ZmGiAmuWsQ8NZXyQKMAQXhl38aHMyGSllVyX9NynkUzdcEq35V2LCtxpa0WA6FXwikE51skD0Pu
X7Rqq2vPWyWRdnRJYdm34dCJnm4Gf2w+iVfjZWOiLbcPKPeqkaeg88NtY4z4NsFbfw9xEN7o3WYU
GdXYxHRCT8f3yyrStFRgHP2bGrMRuCgPEO/mCZhjqI7fJhQW2G9eRg1MALEoilhogxan98M4fi7B
SzIzn7adQk3j2VKrqcQRYKM3ZOYPegYE/vnrb6u8h6AwtUxao6Ngh6tB+C9Am0hDA/EwNi6q9rXt
L3SYUpTjnI/V9wLjfQJFOmbiDY+rCBxkz2BqIdQyoAVqcqIC8dwB9xZnCJmkrtaaZZTC/pLXP2DT
7jw3OvqObFfU1XO+nKedgWd7TYZ5Fd3q/l7eOucyceTQHmh4w4AY5hnNldDAtP8jqDzVLGNrwf3p
6HXnh3nnQ9/46zptcPD7THyvlpAIvD/AkLuD/A6AJPoZ9JX8EAkGb18FrkdoVh7jvYOIR7R+TYzu
S1MZhpoiZqrqDe0W6Kp3qPk1WQD+UcDBFYkAjmVXPG9iR0QcmasKJJXV/pUNxYyDjfd+2ngu/dD9
b+96LsQTJIZ8Xmq9kGhD0LeNDM+ZDbPo73ALRY6SEmE53PJiu7BN9aopwze6xlirLvI7YdOTahpc
+673vARcL9C86PODRtM9Vap6fq7ZqX0SYUIvNkyC7d4x83j5tPzE+WfVoPmjwUSvIaGmw7S0STAV
jXiVljEBYN9K4ptgQ3f9M/xCX8BmDTnOUb/BBbMr2mRuq8aaHFTkEFOGC4nZO8GgGa7KsAGGOgV0
TYN8uIk1Xx0jKRcuKSg+e+i2L9L0G/A1GFL15x+x+CnD0cdf3yAtnEIvvvg727tYaI4lKF/eqIIp
ZqKRzMNTFQUbnL2KzJV1xUz+KC1SxjpjBobFncSm24PZ/R6F6CLiKxiyE2G+ikT9f2jS/MFxH1ko
3JkKbt0/qkD0ajjhOFJEJqn+6KGwtWuyBJrQxoDk3xFUB2XHXQTlqMGiSEcY8wfeR4XBFGL2GPum
jrdUje6t2gd5GKbeo/uG/ubv9+v1ykAszkthAPXQrkYBUM8o9wq3jebkwF5kdoyHeBEx6I470G6+
W0v43clzyR1zXGeTRsY/U/iZUng0r5uFsZJILe3xtUoW7q0zrmqTJ057qXtFrp4swHLcnRsSdnBf
0zbm5jrnnUILAtKxUeGZtpS7rUmdK2H5nbSRBGMixPDlVFnpxDXdSVATXXyHqodYRMv3hiOcgMGY
PSAW02SLe7o64jQpAaStFbKsdob+mOGQ49Wx4ZkvWR7iQBD2maFvPnZfVnhrP2aVxlFb6Y4IogQN
x1J9bAYKa2kcKJQ0f7wKlYGAY9jGOGSCaScL+oWTqTx+CFKY7PWueWD6wHteNl65Q1EzH8Z60POQ
Bp1GJSPV7P3A0z9VjR9qacIgEJu/5LF9Cv0OZ3CTdBMCQagPMALDVzO0DT7m/EAmxIWH7O8sBdkd
5rAHX7crggOSKYOK3iN/M4BoBqWsIVarFOsGCKo0nw4v+JgthBDwtBZQHMNSvDYG9ifaFeVQuSKm
ThGC/z+NJWi7UggMS7xWEYxj9iDsRFVKn7Po41VTAUr42Sa0YoCucNUkHKPLJHLIHfRiacjO8F21
aqBCCP6fTreMEutF5cjnDmIAm/Z5zSRUz6Ryy0mGwavqfp4ai9IqcxJ0MdGbXoFzD5gLzOO170ZY
HCz1rauN3GDuuXC7Iq0XvLGmAZyoF8SEDMfjlqfogPwzk4ulU2szc747R1Fu6Zj0YxaawCtfnJIG
1rVBTq4ueot+W32S/3WSHZtdb9ERsCDuZzRhHuo3sVyTMpv69oZp6mCiGF/KMp//4vHlFGKnlIG9
DHRMjzKnR9woF/WQYg/nUDr3iV1To/PlPsm1QyCz8Vknynnt1BxYr9t/Ts27VN1plVSLIQz7pN8m
LW8zzQtor4INTODY4nj4HQDvJA1VpwDtgoJ/PfBl3kaC95DzRR9vU5WpwdjErm/v1xBjQvtGBmnx
Rh2uyaEVo13C2ZjBHBv3m5g9wwoIyU9kXg97SIEqnUXuX13uoT4GXoNLvPuRiEVcLET19t62wcDN
3DMgUIBrhJrLlxcmvYvFg7YTLvBL/pDSrlpLpwaC9wQvgEZZsRZHuOKbnXAh1nBQZ+QQIRo3obRS
hV+mMznMkfoc/ftbf9dnmM3qltp08GQESVS+UxA333rcSRp1eh6smEIDjJ/alR5MOTGj7ENMttDB
NW93n9ij+gw2ZFysBTkYsoI1PxDk0CvYfZYi4XA+aepPy/2U50MMzw+S3+Dosuv8QBIzOm5+t2rD
1a/XR78o+hX8Gdifl2w8mxuDdbp6JFLrUc5+wct+RjE/JbaoV0X5fEmElBY6rISSZQY87SQ5L6ki
ELYhBLwm79p9GcgtoNJUSPFJekUjKN6WqcQ9eQsh2DNhAAu+8jRhdyykkno9bA2fbbUxgvM4Xysg
llMqWDlxz310TmgYhbbmRrD4yJ2Tl89+1+1ocDfhnQOArDCNmQhzM0GvdD6rdz6jf6qPKttfjJNk
mOvOzqQ5aT2SfBrCMbv1bGAfqaaaV1k3iJmxYUc477V0C2Av/2lZUvwUrhe18ODn3MQ+JCMz4P8t
d2JcHgzQ3OnWBJfUAqHkxOfb3quHzcQa08TKE9X0Ufw9i7w8gMgnE5VFrR7dZFzyQbD/ck0x0Gyn
cIt15EwjNx0JklA/+LPqnXd/YsbuvBkZUaklu2BfeCeKjrHfUwiflRV2sFXQebasi5QX9kyfwHNa
oKD8cMbBrAAP4Qnl857DkNrqA0qq2dyK6q1Gz2W6f7brdUNYaSf3OPaaOTpmgvofh/7k3tKoTc4V
ZdAFuPKH+cJPyFMurxmftProOXIHNsJnlBsMshR6yoloLM2p+iSiRhFZJvua8ZoT/i1jp+gpK893
67oikwi7LNlaXLRRZxQQGAi0IiwmEcVrR+aGXila6rMyyZQk7MYzMJmlYMLKIbL1WhMggbl6bN3l
lR5TugqF1yh682kyomw/+udd2Rg2NZrIqJ90icZP+LphpAaHZPDRcdCD7SwnZXa+3sz6y4479Elu
lsLgdYPyfdKSpbsEK0m/gR4Yz99Depg7gjtjxEt1wGzH8GyQbRz4wWZwIkYP3MLPp9Ed3BtyoMSn
h2VL8c0zmWl1kkFeqR8PlF/K4BjHX9VRIG7bcVbfKLbvWQRc15HIXbr/lMoQz51XsahaNQYj2RLw
C0PgRbGbKMyed0BGld82uydGnzym51artTnevDDM9v0xG8UrnbWos9IxFR43jQEuL6IYH8vwGVar
klWyRdpciWWdj2bz5fxqESl29XIR4L2dGWRUcb9U6USf/HLmieWV5Y8rddTTDpnPeNhZMFnACjb0
Jo9EBRS/C2EkO8ycf7lPbQlrdsm4XvaOFK7lXwpqxQFtDcuDe63sMbP51Wx0icT5wCWhcrBXTket
dPHbVVcRYMPq1uYIintwuCeXv1FskXYUzfQA1RkrsnALv2a05AKI0xVkSnrMv0PPOqJUfDcY96KB
9LzASP8sec/gdWxfgZ9WmYmEFN4hIUUsFt1n5BdwIyQ+BJN0YFTCQstSqSpyWP5bGal9wDWJImFd
YovlbEg2NSP6qfEj3z6MZw+zWt5Y9MU5s7TYJyc94IfEpaAh3tWPrT3m31gMc5EuTNJ7KzknyPqm
sbjkK33qoduoTHHKNRBrsJR2SMh52bZY+8I2SiDtyYjMuqe4jFbXG4AFxGVdNvSxFCRRFCrKHVBx
MVOJ/Kgd/ZF5/3vBkpbauGRN6FgUWE0hlgUWfVMbL/i2tBllywvQ5XFwsSM72sku/TP1jW0Tplza
G7s4A2oNdV9QMfCD5bUlIdVzYoTLaDndefO4CDJG1hEuD98Fyrj1sJ8mK4phpk2udDceUiQbs6/F
nkvlinuvkIPb5PQC0br33dUpc2cRoJMhkqKvjRWPZbWVUoj1lhEBQqSXkgzBc01W3NGyvT3T6M2N
Kxh3LY9hEXAzUNQ+5hVwUmFdeCB51xwlSCCxdpCwhePz269yrNvFjD+MWDQy8qlDfHnmUKFw8vnM
8t0d4MHnt9BbgEQxrvJO5f6i/LH2vRKey+qOagoKDWwD5mNK8MhrN9eYloFjGGL2L2uJFlunQ6WJ
jyVulh8PmV1JMFh0VsPJXpz+0HjbWMf1hZlGC8FC0CBXO45b5RZRzrz6sUeFlTiRdVy+6CO8+kCw
aXcqjyoWsaND1dhuzk8yrhTbKvTHxe2ZJO67xtMSF2zQ4W7VchI7/RybDf+gzAbzwcV4EPkTppPu
b9x4BA88h9J4ix7GTva6qBSWCrJ765UNstpxY8zuwwiyZBMpDbrTx2/ywtla47fPDm+n3D0O0v6F
/w9Xgf8uR9L3n2E9JYNrR3iYVqY4bXJ5dtn71LV7BT2Frcsb8zjkpXRKMM0wWF0VPSk7/clA+Kd3
Fc+XIDUL4s6Tj98xI/pfJmVYoPGCTq2jjC2xg8HzbJCjbheRRuKzwH0J/t+fMouVHy95CdW+N3uZ
jwR/A1G+Yz647K5tbEdqVHlvH9x4azV+vf4+zSIe6z17BHIq5ZbLL828obpYrqVKc9HBTiNVvC6P
UmBiLc9YA4Mgoj1n6Q37A45ZZBEWkh7N3rZ9RMdTZPdNuc718JWggTWTlj97LZWEZ1TQSit0khMU
ZPu/mgvXZxlLqYuChMVrDeGo89obe2y8I/1T5/2BVUrdmO+XyNpYB5sp3cMzy7Vcn9rjkhwnaxqu
BKgV++0wNy5N5ibwrldflQwxfkdpeUS/41pCXlCmSmEW4VSKJnojt7DhAEthE9pFBTKwEemMJP8b
L17qsi1uamzQQsjfPL+SFBHdJY6CM/af0OGYv4CZmfncL9EwqmaQhVLFngty7VrgblD/ZnsTVGz3
+tWLK7N+BswNYEal+h0dY1j0/AHHRa5/7rvI9+Ov8azDdoDPyFxJaPc8aI0ai+w4TkCn79ip/3Aw
HuN4MptRgImVU+KnHRlDwDH8sn/hRM1DTkTMtMOFYLDgqA36yONIHyCqWBeXut9ZSMIjQO2O1yIR
4JnDbYhoPqDBq8R5GxAsy4+nbuFcmk4DIhlHCzonEJlApMqypxlhpCwdfNN5/hbQWaXRKoa0Ni/r
hk6db6koJWr8kr9mVvzViKa65NQqqixgBBRmwV2juHz9RdOVPOFxUxiRrF5pVdA8mnQSAqUtYrKC
WYr5ehTqnU9QMS1ysWvcp1C1CC5Q01HMSZ5P59kyfBfcJVVz9E6SG6tYNTXg3NxDsnZkxLr3kOJ2
AqekY0inmimNKjPyesxSTLZ5Xs9tIuxV4Jo6VWFhz1zkZQXL+a1NA8FZmw60QKn8y7gCd2VGWHrf
CcRAxJu/sqgKC9/xvmuhFyxWKBnoqG7tOpPWHmQJT0avDKmbdnSiLXV+lgEdyxzUCrWuAMKb7/Pg
OYTdlAjAJU4BZ3svzzEksFn96oPoG7oGn0yXZlbuI2hKHKFzdXZUmwaAzRfjFEZ0BUsp1/kyc/UG
iHo8V7fYMPZOQU0YszEOeZQPIfMDHLXtycQ0xJmgWV9hjeD6gJ1FgXJ6unAdz82YTtiizsS8/Ki5
UnUPS7OLodUjdNezlgE5KnY+Sjwi6Wdbg78N2lAIXxe7FPogSsabH6NUBMQDD4BR4VEdf3F7JOne
9VY9uEU/s1SR6JbseuKtP9uhjTEaShGEBhf0l1roSL/VMZh63A0uqEhQcHFzaU0XnrtN4/xq/zWy
9Ucx8o18Q3gzFbNORRBc0gVe8h9xC4bVvjcgKr6oELf2SqdjGN90mUsFjnAZxDBqo2ILHSAV3kM4
SL3dBvmFPcjnwOxj9qccIbpqN7adHgjFeydX+homjzmoYlNWL0+EDwTgST94WIqCjZknSDMreBwo
qTldizO6a1fJLeVx6u9rG/XUwn7XjytW4HlfnYXuMn5G3smWqBY5V2LhdovQZYMRv/uxi0EQfqmQ
43+mVNTCj3tSh7rSx294ZI3bAO30sWc6X7qTenWcEYfVafMZxTxA73GSNOJ38zAAYvq112F2FgVz
6pMUT1Av5Vs18o01KBHs/YOIL9BYjZ6jVxa9Kz9HPncnjwKzbVUrmeHOydLyVBqOVvg1jGmKCA1A
HrwtNnDFvpJ1hwDuwFSohJBj3owOS5uMjtFUKgWuhpmkvxEhs+LtU9KQjzYysL0JJLom5iBGuBMR
ROFAaURqrBPh8m2wuU1qef3agpg8cd+AS6FWYWxOucr2/0Qy8cv+NnmfL5mc6GsOpctA/MKxl57v
iYdmJGcwxV0T0Moxv6VXhJklkAub9Eyhn6hiyiF1TLh3wpQbFgClG3dlTqL7qW+TMz2Axl/gHtI+
anVUls/+JuxDjVZS9Yz9B4jcabzloPj6JtHML8XADihppiL9vPRSSZepDxgP+NEHY7O/KrHBYdq1
DkPPTXPFTxtraiHvItcrUO4F/NNY5PlOs1HFNx1WC/3H+UWSuuXSUAZ8bUjEtXPFAdTLTArBp48n
D4qd7oiR/CWfLZ6J+cWL5zpipMAfEbQFhqsDjbcrfXBdBgztosMYScH5mfcvRBjhbZP+WCLI6a1I
68FrhNk5RePZY0DsFOIHzsi5uGrVIhDUtSDX9glAr0CxC2rigHMKNtK5FCcrEjS4szX1GpJ8/59V
GwFhAHG+sR0asIUpAQq8/W67xFxDG29cIgXuMWW2A6yH0q8BrNEmdZ8+r0i1gd+Zr+rUDfMTfl2C
22dDSOj7KHKeiHZ+Qt+wSVclRvuk5Cr3KNPh/foq+WJlBQwIJpE+Re/5TmdBc/tJMysNkyXQ2nLZ
eCeqcNCucBgaKOCRmJHXDchiDuivqpi8FA0sLqgYP4aj/U/Bhs8W2WQ4SG+/FkVF3FHJllZYNGuz
+2FPdvVHd8HrluQ3RAMBMHc0eb3ofGaA60jVlsbj7q08HwguVLNP5vCIwaPsqGB2sx/f0KeoMyNH
0Q9kPAynue7TAyHMf8eXe4akendQwyPxKfdXGvy+Jz0gpAiFQYoHpKMR3U5OnboVBAX2gY2Hp3e/
XggehMZb/uKlX0/Uz2PMMDNUHz8mAS0CRh4tgITBiG/R2UP71kWxI6hPBoDYPGDsO51+T46vGwvJ
HEmtZXQ6kl4MTQ0Pn87g0WXlK+pE6mqtUwQQ1krO0UVSBLORrsDm9PByI6PLil39KYIJnd+JVigb
CRzlpNIq7oIihLgWH5IH8FjBS6lj4nPMtZb8iMB9Ce5lfPFBURXKRMtyjJh1bkB1wO8arzm4RmSQ
RXTBlX3Pz87jKhXAoHS+2Jx0/XGZsaaxx+0oYphqtJPDiCJ/znJKqZE2Iszu+sMm2MY5vyucNhKL
o/DZBsCjvljzyqZtHukg3bZmqKdhTAKWHe7MteEQd72OOc1J9n8UVvXw1xVVUKEQR0E+Wa4Qt//B
Kmuw3lmsY66XSezKtR84VxD7TBno/vxqoCviANJELLqisS+uG3AOnKF/E2vLo4yN/iCzVz+Lb1I/
GXrouMAvKxMcbnsPBZ++AeWNoFkK3w1PRRT1QK5a88dtVyxt2jFLFYw240dB8ia5/zO7tGm8rOG5
uC+7FAmKfO2Cuzv6RqyFRUcz59emIdIiMNouPC/jy3MNlLBMJnQdh+TIBRixhh18IzxKXglwG/ug
ejaplLadnTvp95SKcLbP4MfU/lq00LiN95jJVYvfLmwMGDlD/yNnZZetIlOyxnEaaKN55ev4tvP8
e1XFDcEvwP9A/Bfyk4/3iw9Z3Qqgf267V+1eDd25XayPGBEIqg9ghD76nVYdx+uvdabn/OlpNj9Y
JcpZuxye2MYJvU126rQh+0nTbIafsV4ODUimb1NzimJkGOHu3YtyWuXd0U2422En3IYhhsJcHXdB
SwN2+HmIqXSi5emSUSKjr4ptEYbuRlXPKAOPks8zzbnmd6M+YE8wEQO6h5UKGXrtU7+BlCkkLbvE
0eVQUpGrsEyVB+f/FnUwnWeMECsLpXL01n8D7tdIcPFsKLm7ywaO2ArxmRCq7Z2oaDy+v6/EzwxO
8o8e98WVGiwk9OlU1xqdA8RCWltSF29MzvcOqIYZSJJUqVDTICVh0c6KoS32WxtVeQDDqAf5opB8
j55xC0ivjmVi8k50ld9+l7D563alw5z7f/3y9q8zaisDn8vG1ybdxHBnoyaHPKyGIyzmy/fQ8TA0
aBiZc2kBoXFH3VMjArZepmeK4TaPeQee4TqWiOMtYTCFDKj+6ivLQ/aFj3jF8HFa1Fl/wopI2tr0
hOlEuXLKEe3VeIGp+fke8BlFjsZ4cWVVYr2/DrQt2yXZGMq80TtiQ3GUVjiG3Q1lxsqytkVU70Tf
8fiqwN5iN9ZtNIBg2zdm8Czx5LBfcjGfp8wBTSaSa3MHByFqC4dYFPNAaBHeDj0msK3Kgz0nzVPV
rOrSOyh86ZgUQmG+wqrwP+BBYiRO6P1nG38xX0edWAggj5PjmiSP6Ujo97qopJ1OlTOTfjot+DOy
FD1WUAyv29i/AUavbEFjS1WvFG3QN9FAyN6xAclstxbIoA06NHbeT0J7qwaMXM/txW3wDyxV3oVF
j9+ryRIU01SBCiWNZ8o7Tvskl4yoZMvX4WkncY9gQz2uJGH+tikB32Sebz4mgvAx3xcjiGZVpWWp
w4LdfAMRQkfq0qPz0v4lQvLbX1I3qDerUarLAEC+HiwtLnE2M68Ibkz/rYKl27hHNzeO6LqwHT8R
r1fsy5fFnez/RjAWhjgflnkB/ZZulacLRI3vhkRm58I+PeXv5qGtKxae65Yda47sRKhoxRJ19FRx
V49e6Q3iavyBRVVwk/vSBBl/DS3zk356TnZ623tahSz2HxCgbU+JUIgIQBmIGMscamyOop8XkgQ9
TXZupnwMfyauqtjxXJhayz5gJZSdAF27FhY4f3eehNGvcLHzJD7VbdtdyARl6t0p1KrN+BDptHIx
H6PshdI7j5/pzucMWA8HD7yTD13edPDEQ3pOX5tppON96dfWkJulXC5OJxRh26a4urocEWVwb5U+
ufDoNMN4BPJC5hQ4iviVpGyBA8ZZybC4OM0ug211D35FXvMwtZT+PC4vw5XvjUPbRiSLM5QQrNS0
7J1luK+Ldbb0ipwJTowVYKPoq/24Vg/rccy6zP0WnK3RvsBR8nnqPdhU/WW3lUYkeia6acojoBlX
eefDSR0F0UzoJD2VJwo43j3lmwLm0kJ+B957Kw6ezplUIECOCCGV/737RBejni2Ekn44mrn9/IR8
JdT05eBkP+kQ3TAkcZ/VmSjKeu2CF3w1EEFP9mDt3Psfp1FHHwQYJnyANLOpbiMQ0KNT77H37QDW
svvd+IW/F9t0mTQ08vPo3lzmsBhFAL9Jt7xnr2QeiO2hWzbMxD7kbHQfvEK6KGmbtDHpjK6ZaweV
22qi8td4n9iMEK0cqEEyebVNviAlKvyI18m0qpAhB2iDVqGCoRTETRei68E5X9yzqJ/flvuuuGSy
0EXdpCiBvYv+KluyKxTZlILAmWOgEo/XkyHqHxDwAkuU+shA/gP4ykyQ1HujToS+K7gw+wAFKiJD
W/u6tcLM/TpA3UyiMo4okzyqDV1Fnz4cRLt4aQdsGRj9B+fowJduHI127cSgS8piOljTTDCmWZ5M
CSR5PbTN1XwMJiyMe7Vf+wJGTnGC/tuMjBr9ULnM1q3wauu7Pp7MlNWi1+v6/6AgNqNhAv2Xzm7h
YcLXppLJGmOvcpHp9X/RXmO3CQr4km0d0FV3VBMfxj3RsvXT85CE9p5Sd3m1BDwPJqwwWMxYMZsF
pijoclQ92FsCDp1cvTJmS9lofMpEpTBjylgZc37VGKFX/qUtSRsc5SdAMgezlK1w0JDZVcFF00H1
kWr2Iep/brtqz4Iw93D630KBUaR111WBXUw+FoEEm75wEe5exqD5BdE90BuiJmXL9NCxFSqVVWvS
XgWNolc2wgpjJKPjxDolmON2o7caeRaZpHntVn7gqiE1GtOg88y4KRBmBXQmWeX2WHnZPWIQi3TR
CVosHJ+MN0WsB3fBLPGGfwiWaZ/ngib339JpXI1nLWiVJxoBTXSf2UdTwsyMUgWmZHevEiWflVH3
Xalq7BRBDcnPbyfNmyQTS3UgupHbEsFzOFK53NdQepnGT36SiDBSeShyVmtryEmRgCSXD5AjvDZP
h5Xoei8i78OdwVuAKNNi5ug3DNnnYpqR1ebGb9U7R1eTnv1q5thEPJPJk4bPWba5UZEua+0ZUlPA
0iTnaR1zuk3A/cvkLVGpg+GomTBYEuN0iXlPBWm2Jf2VyrojDP7lESKbsx2R38F/KaIXmsioOj+1
vu54IZz9JHrEysjdk1u4CPdmIA4B01/k2N2tmR6WF6BnLYGjUxoZV4FiNjeGVkSvTsbpVF8H65ot
lUt4dD0hKzirHbgYzjrBM/OZcWfzJTvpgP9IG+xK9Le40UfxEImjbUu+o/n9LSoRIrYv74eaKvys
kf2+RX30LXDySW3yDmrrbeo7z5MdHJc5t05s36KeHVXpCpRyb3iKn+GrLNzPQwEt/8Qs+g1z0Y0B
wR2V1gUQfOZ3F5oPOu6TgV0HMciXZB7xWvn0CV0MApKCtdbXAAfRchuu+bJpqE0bYuyDCXmTjeWV
zY6ieWPhL8txEzK4c98gDFYc+Kk0kajWzRwbry7KCzwi3eoyh2HrkjJ9rMerkAlxQv+zcpZQaxyi
eU86FVHe9mdlVz/CXfRImU0ArF4dqAiZ2Usw79LdFJRUuwvZ/2Erf0ivc2qDT13nIbFFDiSxgzfd
Ay8evpHur0hX2+Z3EbpLG8P/jxflcDV5LL4Iz/L6hzU2mtHhfrepw8DChe4qnc3NiEGQ2B1QBj/0
6bVnbxvi4KR3pb5jq1lK+Ki3b+SYcICZNojbcrdyFzkkFXGglK8J4X1wCzJy8I/DI692PNQ2vIPk
yj4R3JzPQZTq2QtTjEw5VUHqwkcqm8baQbcX5iVJjIlwXTJXA2hfVBW1qrgPcvR5t45aocy3VZAw
XUausz5JoF1nnTSyb1ile143Avd+hGl0IRxeGmLyPFbkPdeJtvq9NBZxMXK4YLtAMtlpszJAKkLg
VP69lm8OlVMIvytfoqE1DugxL1comDBDKIkLg2twqMNRpF10ywQXkZavQU1yerCLrFozA8xIf/Tb
lQhFe5du/LjgcUXUiGYeoGullxZwxFmNIiybob+V6whfemgn8mPKONB0LlGFPnaEKmhf4nKtrDgu
UzYfX/TkJy8NcAH4pT4btWlCFDp8EvPu+ZeKdLIigt2JR6/aaEQKllYl5FDNgtq2gXrBCB+C6MOU
HETqEedzxTEGaOg0xQiuulBlQTNAhRaA578344GWfRljBHehVceOd5wqjpih6U/Td9t9lwBNRIdL
VPwnnzacfstcV3WcpLqC9Lg3K1wRUppMTtgYR4REuXbnqFg5r8eg0R11ovoEsnUbysJ/V5ja9RDY
4UdYyLL2tUGMyPkLO+C0ZRQCR94L3dLVlN2g8fQ9hjlac/H/gzDpxcmtvFtfL1z3JZ48cu6fvIFO
YNr3jqK+1OK0k6a8z+LRoRsC1kWanfty5uKmQkuSNbtShe6ej2uQ3yEHKK3BxOE3gl/Se/ok3WKG
DGNiEkBk/rWQ7NB28IoOrNXC0S31NJpg9ekGXsuPypcNAU5yrqKoPJAOurmCQT5jnt9GJYk+TsBj
fMZ2d7uwsDjVlwpM1sgM0IOjbTAQd26MFS5Wlkik1kxR3Ql0lRIkTKPBUfl+T4hAYtlENuVJXPu8
3OuOY8AWT1WY1Y6abiucAE0E6AjBDZao4x5IoBqCKQo65HgZcp3yEKZ+MjOD35Kj4iaorKfoCbRp
1BGkpRcdsA3lC7wa7f53tfE833b4UzsFBbXcwzaXVQbxT1eEnu7JpqNvpPNzQCbeuS4KEWUihJ4H
lDiZPxfAMTnn6SFQHZtB9cKse0UZgESJtB/1C9bxukmKYRfhVBKsPt2AFiW5WuqsWsIRXFoA+moH
w13UGvNuSbcF95NogBNuAnSBEOpaQNQ/XGPYu+gzPgCzkFhf1HhbpnM0OKiIZP0UzPsO/iFIQBB9
ZtLGKzP9MQbocLil0Jul5QlNi7oiW3swXpYM1N8xcNjxB57BHeMJ0yqLxfSNBm76N/zsF/BD3KrZ
AibCkchvRG42v9cHEJW+YXm0FsEMIQVf1wILPsBKoHXKFDQCrwm3jJIH4gqSpBKjvTE+M11e3GdF
MLK5sTKP98b4byydiHlxd0AZU/4bOEnPaoHe5TlQ4VI3uWsvuk6w8oi62R9qH+2IHFOpUfObQNnY
+UdIuIybjZg9smXtcuFZP55VeZ4WI8FoAivoogioSCpaCuGU4j655rSn08uF6dCR00Z0epNL04IJ
FGWYEwOGQdNkB66MO9ovYsIP2AeMh2AAtKog4M+cafEgShleJqRLy+a+trJKDvqDDT/gaCVCGKLh
JDxM4sc2d+DLCSJpuCMVmb7I3a5y
`protect end_protected
