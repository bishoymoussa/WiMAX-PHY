-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
iDIIQZ3DRuBbIVvkvtGSi+5/C1DRFAYLOeSTLCIb1hAYMoL/gkY2sY6alA6UV3ZOqkdrYMlRMIPq
D9xzhUmWeEuaOpimMZVyaAuoSoYM5nks/hleQq4SEIu2hdZblonWKWOzOb+p/JpLxC/goWeiD2k0
BlbR4ahOYzh8vkLikRBo3MZhnsMlO1ZtprpPPMNJjzqCBzzMzBAYTX3vyyhc4Iqvcm4ijA7UqTld
F1YE1OFYYEcxbHAurHyRID9rCnQmmw7N9oX2Sy2r/JYgEUhiNBJ52Kfb8TtcS3NnD5WNs8k0Rlr6
GpcjMm+U2luGoSBLouztZB3YC6O7YUWyGsRsZg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 194096)
`protect data_block
8G7ePG4LO67qmjY/O85yHrcP9yAAoDd1t9Tz9MvNaTY1aZB/K+Av9vNo6Uo5tDXJxtUduoDjJWPd
EdNWlxwEwAW/ZKhupBAmWVZkDLleHFe7myh9AgaGypTFCbcKwOCilY0IKmBjUCCGy+r0SGD15x+g
T1Dz+AQ7oxnng5OKBUwtZjiJWQD4qP54LY8xuw+ByEQzjciFO4hOqoJGlwl70N/GacDW9EvB415K
C/9/YBsv4gUBnTCt0jH8elCK0swhq3v1JJjsfjLVbj06q6jvIdY5g2hF2CRXFRHwj0pco4uXFrU2
o17TYnraGsKU9pBzQPsgP5YN+2KxGftsYXNGbTAf9oGGDhWzw8sChEYHEK5oQW8tHVRs0MlXU80o
8sgEgP9V7gdqK0Hl8w80d6ulgwDXj1bXtvZ5rWAfor4DpmN8++DPpqyn+2nehDlEQrEOA3CWN1G/
pvxxM5IwwfbUAib6ZIMCdyBv8QmAEz9bUNXonnn8/wQAx0/m1AprWKI9cUsd8OqRb/QC0KXk/S59
sE3GAvJ2ug9dg+5bycyWtdyGY07jHUisbB1QD4S6whqhXh29T8QHcNAV5ZfvqRPp4SOn8VMhFk5S
dC7p9QzMpKUWQTzh+C0F7tlHg3nXP++buj7byV9a+Xll5TiZX0+g8kp9wuFMXo+4rO1E4gRQ6j9H
2wa/7d5qPVHUo899X5CrlW3ymOhNRNrMSMqO4kdxDJZqjZh/l0RnlJiyInGPNnuogIN4We9repPV
soFJZ+JRvJZMNXPBVneD1s3HAYIF/W8oUa0RJyYQcvG5dqqthfpwS+JHMC0Y7EbIlhzTUsTIoQxv
2c9CYNWwmMQseZofPKz9444PJqIZShUJdauXFzRrQVForIsaK/7gNfe2HySZc6xETR0Z9fcIwHAW
WmGVFtQ80BsUjq+NTFTMNnh3D68X3P/ZqPygK/krNVEiJRUCpY30jp3uVPHRTxM2JqzdtDe/fKte
rqtOcmuQImZlPiQeIdmg1+8aVP3EHB48EplN4z/cKtfCpNhVeU9/RiNPBV+t8F1BFamb/q99njKJ
c61I3wSje0MvkDfQUO4992amU3e5coBT4zS1/3tai/FrXq53VAqo340ZsPlbzFhPofSIuqwFbqzR
/G59gKeHvCj2JGm7RkVGh/VDfrk+GS6r8CUUv4ImJ++8HD0HPTx3wRLuAiVMnkvhH/78qrugi+VS
8lPlxIhePdXUb4Ng5i+XWEIQwTxp90CtNhHyFMzFWoHPwNCp5gT6DraNMsG0bt25WaoIT/pNfJW8
4rzqghVIU7IXblvvVFzujcvlGpZqvyeOc6W6hjeTsiKaE8SlQgM9aGjjSSOfc09K1A4vxAu5uGEj
ZhgtDVHtfSj1bEo7yviTuiycCVibaWdq9JzVktXeV9E5ZSD0xBP70TbLACIqFP0U6ghoRD6ZmoFx
P8/PeOlTNf1lLXxNbgWVB4XvUkH5aWSR22S+BZLDw22RkYNXqCLx8eMHs6dTfHXV4RtuFQPQedvK
s0RGbv2WGX0P0baeyjprrM168nKdfoMQmTPtuimV4svH8UvxLSXP179bJ6HglgQhyglBrxfv3INS
//2zMJY7fd38zH7T88waP5uDX6E3HOpI/2dQAUPNA82bGHFIhsNmHrQRxtx9KKpsAHOz09BCygpU
jebki/axa0wUQvGdsJ4iCnA+Purbbht6VwgGIoFRwlZ8I2Q01KqeAOWzXNkDEZkCVoJD/4cKUU6U
PpPTFOhzoU4CGpQe7D45tNwZsSRLzI9546QIndcLTCSsEo4w+7FPfzSkUUbyFi6+gHvWLsgtQPoz
TIXj/CAvKPl7rJj+QjkXmpVr8qvIVDs3YymUya2loUNYjda+hC0o9lkvXovBvN1tg93nRPp++hna
GkUQQOr+o65Y3on+tshJfC0wa1ui91oI7k7SrqBGRccsSZJawPCyzC/eJx7DO1r/f+oef2B2egS1
TUp32Fwwodd5XL5QBADRErJDUoDG+G2MATNKTq5pEIRzUU+Hb+N/aMmiGmBOOWjOh9x1Awmu/vpP
r15tq+wtsTuX6UiGYS12wncWXkbj6dvryi3gjnwl/ddheSeYhNCGtFOA8ECG7rB/yeiLlnYn1o0Z
NqyX4HqL8a86fz7i7vLuvX0aYWn/pkntJFrGSl64B9JY6A6qMqeRlU1AgO1j/XydW9MCbZPHWgOq
sdZeHfFBZ82vdVTDbiNFGRkV9sshHiJwBWKuKNc6av/FlGJt1v5lgarePPLflEMeI2xD2xRypkFn
uzmVO6KOHwAALCPwtFx9mUFj8YysSFjNdBTKhFw6GcpJvMT7GE2OSgILMO3kUyYZA/Oa5iraFLBa
tBp9E6mT7z3tsx/NHwVx8q+iA2XDP72KNOGZAlMcTXPh/jyO1k83U9F/3hm4tM3ZoeBYySIwRXka
amfdSCEZxz5EWDYrVVPQwPztXZTi3G4iwMrs2TyzPuMIB40FGSIuHQopfkc78fVsY10IUcNqczIb
d5Tv2so7mPj91xfXb/ayyL+v7mfBHp55qO3uaCdX6275XP8FA1pe1RMIYu2Eq4+snWrCNmM8IfaA
WhRN9p2LN1OGiGYg1BLsHWYDRlwNsBVuKD2YxAXABEaItC7KnSAwY6wTVpbJmmHPyaQM7cW7y71Y
B5Boo34zPGeSSOgDGwbYthBuftubjWa87zo3d5DBmj/+17A6WtFyV3mqLemKO/tDC3BnOLymHyA2
3MaBxn35CNit0wni8yFiK5erqumgOL9vfb31fPKLjk6kbIoJlQjsYldKjSLb1xoWO2i48iscQSd8
HNQAV2aQ5Q1+dukNFMjgzmo3QYRnRCatf4W7hSjHmLPd2g8bPzyvj6wEG7898iL1t/ChYDTJA5vQ
O7MiM8fK6SlyV+0jw/ncw68AHof6kXAeR0dWoQXN4p6lDVtEsEcbjuxpBKgHxJTHCjg4aVThJFM1
VZYJ6n6KHLtAwAwFji2q5+hCxQrcwq3rrdL3FqSy3bs88OGkTlRSHPUuwPWUbZFXlSOTCNeRzkq5
xhnnhpW8KhEecwUYs3QUqsGV3Gx4jTlbRhMmS0S3dYCKWK2P5D/BtzrYSfN57RBYBlQjZNRVATv3
IgnAbpq/yO02SY1W4ehSYvgMvJ6Pa/NVwZ8AqK5VVo6KS/LAlVcvNgbxPz5ZZPiDaKLSuriHznwW
oQA3TinTXWfOW/s54uJvb0upQTBSzA3nivW9i1WwU1iD94CVy7zUA3aL8m0w+chqwLBsV/TiMrtT
ClMHosy8CjzVa6CRh67EjXT1vEjJScVTx+37YKlbkJiNfCbD06ZR/vLKla1HYlWF3GWhUz5BzpaE
EqRgTTYzkAxjoaDkB1JAn7WFMzUUYVe3d38aS3RwET8H1eY51wDS8n5nWEFFsUYM0f+I4RGDIwDT
xMa0n51S7GqTry53HqcqoLCPI/r9+Z5xmXh119L2Qbg/n8oLcvyVEAyZyKmtYMzvb6nz/I52THTV
XXwXKdQkXwREPa1G3JL0QnG5GQwiQmlsnUdHbgqDqpzi8K7rKqY5aeR6qTYfNgr+NJwn9LGR5dSp
/ugKtCqAnx9oNIBgmvj9TZ3BsYjnRmFDnpWvtHinroDg6mi6X8hHBkc4SX9GG+VFpjSlzdr1v1BQ
Wm27qER63SOzCFYgAQhOrdkVjeY6YOsCCNK06JUw5zh9RRFijoz8/easxxPZT6EyHr8vMvK0Uh/0
AxwzMcNZH7unjwHjOUqf8NHWIdcfLJQt0/QGwqxLPauqCXq1mwa/zkRZqoQmm9mzyxY5aTHNJhIp
ZBLwyffHbh4XUxag9SkPtVinrMwDOHhTsHDsiFE1ZTJwGMZGEWmBuxhufP2n94iS4Scrq09hpFLk
qPwl6sV9Gpd3YK7NU3Ob3Q2HN9+zMtqZ/r0w7i0Rme9yx8cjrMowoIFbK3LpllORykZXAAH1nKzo
ugvrA9rP7Il1yxrufBaZJHK4A1kVPfJDsl4sJ1ZWYUuo9sNkq+yB0wWlKvv989u0ULjWhey4xB5n
bEbYX/rBmbjq71UIrUBCM4p+NxkhPpr6fqVm8R56/qPULGcu09drkCWk0HwaPgzztcGZ5SBPhcxg
bmQaen0PYITnCpkoO+jYSw4tB6bn4yZEEm8VXwu9Bsv/p++tCPuu0b94tQOVyx+XzhwAb6M8qqpA
Ql0n3qP3jZ7n6clw/1nIMPH/W+i0cjq2o/LYXNrnJSmljGgbtFHF9tdbVbnGPADghMYKTvjJMBNA
czcmv4bitpch8elxmx9BoBbmniQK7bRdZgtINCZ7ZE/arcL7SETl1CoPo/SXIdH/tY/dvkWhFeSD
U2yNifdygkxyumU6RSU9k9UI53kAFI//5orIuArLz46dK+nA+KXLkE2X0nsqcWORYi0D0HziwmkQ
9G+HmNJjBZE+adO6jVsVEtsDth5TOmo9nIznvNN5C7vHR6hYlrIQW66GytUKS6N1JVRDILRkXTq1
x1yD71ldxc0wiawyn+Z2wZAHuQiIELPzftSKcd/FQU8ekDduKtK31KXmVRhBgMdGlb9nwTtmlJdR
Hvh3ilHRtbuyoIY8vKwhg5Sl0kU4uEiFO6+GovCoWRlXjMdeDtDdx4bGJ5g0hHdHKE/sAMeXwNf1
hS4jZ/NyPPCOzIwNfKLMqAbpi9cQQNu5FBxqMCaYnxC9Qp/ZT/iQmFhT8o6D6pe+rZDsnr70hSpZ
ZUO8ixDVGK8Rg2+9sXngpvOu4gklWwO1RL+mBxsW1jD5fkoRNGweYk5VbtM6F/NnJbnmgbi0vyLN
KvJN/lIlavUw574WFtvWfFGABH+52bcAJqykrhmX6yynSnjkD18ZkXYkyLZ7PI9SliMBoTCnzNlR
yVd1fDm7V2lFngkPDQ5yah6e7qi2lk3ujsLqD1D10ZdcKOWiU55l9sEamVm8phlgYVf6+/bgSIDJ
NjTiBvK2Q4AjoS0P0q1prz7CG8KGldrR7jUHyWXpEWzWBwyNnTHhYl4/vQOaRWqMej2lRbvbh3oQ
9QvQaeKI622hE3Z2teLbxch/zXuSGZcq6AvGS3TcIr5QKcVTfHppu/z4R0c3xcwfEH3Xre+IVe/u
+q44d8HGXFYCx0+y2tNf4FiFnlVEyqLcE4JL6pzt4OzNuUayvsPCRDE7RdeYMsNXEGTMoXey+z/m
YMLNnEFa9SJUZxvbAvxlvFSLSNoP2SqGg77+wWcQUkxKvM9KeXcjMFY6WpNbokeh/wz005t1R9PP
R8FySM5q9SJD1w/goy52CDsEiQKmsg2P1Uy6cGUWpHUdSNNVh5vUJo4MpK45HZerZ0kLnD1H3LBr
u4SgYlpwOgNqRCrpQXAzt/wcZ9nElYgM+rj6zF0rrb2krz0nScjUqeB0agl0GBqvh8ERNiO+aPmO
2GTc/XJrKpQv0jYkfY0q9FfD4XloCdr0HFio/R7kYAi33tpU47GIchvX+IGxot7go+XQUiBgbR9s
VnPEI+sL3+gdyxeJoo6zk2gOKqLx1z8XX6Hpyn5oVy4JQJv768QxDbncu8LLjc0khGsMObHFKX9Q
JKJc2g7zaja9Rj2h8w483txG/XG+0YZDi2HQB2W/BT5lfu7ACoEzpo+3oufzXjrSolh8ytc3bUdq
FaaZnQhCl68OawJvpymvFbdATo3c4D5+Il7rCrPfuMffBXrpAyIzLilORrBpOK8WxwhabO9TRH06
pxA6CH77B+EJuSVUqp2cIK7l4dpWsAmVoDU6hCBl7PAFju7ut6eTC9/yGK8NootOnPsOHGuSW6bv
rIFU1+7L6gmvvUI90DhOiO06+XXwjxzmauojSJe+rnn+IPcbyg4Iom8Dzfw9g2JP3M+V+Eol/UBb
ZgBzz/MsgUAoKF5a0JMYGfFlWfCnaHTl7TTFJ623Bde51JoJiAERtdC57m9+wo9HDq5S605bPECp
crD3luiOJus+TxR4o7iPzNPjDECnWuIAYgl6wjIS9RUxaNr+KcTPD0XxdJur2//bdyApqS7bvGlE
oz09Bbx4QUwHQ7VtD9h9DpUIvId+Lo7qmjFxcp1nwIhhPnDam+YcZp4Kf8dQWqIRNpj8kILRqpvA
DfvapA+azjcuRrCczM1Q9wmDepZ+QxmIyvWr2xMYe6aNUvoBBMcZrCDiQc1Ok9Lj/xSFQ9irMW7Z
S3UjnqNQ95SNg+86v97C8n/C18GzNNABb+dU67i9j7o5gmWy7Hi6Zbk5t0HXpaz5dLFx89CNHAkg
boO9Sb4G5plVrwoiPfIUb8TpTeMqmoyTSdGXovjS6gACh3+BTCJ4vUrpfTqySTXoAlPqvw9FTAnV
E2iuY3stv83rfcMx/tt6VOdCSPkvZHhL+EzaaKn73Nx15EIAeBPEMMg8qP3gTCGj0Hi4ihLNG7jU
E6q136E+Kijxu4hGRX6H/a0kOvMESJFg6fFsSEe0VTK1tzv4Bbt105neOQn1wsGV2ooXf5Ujz8iq
RC48LqOurQXbxHPutFR9R9ykjdVpFT1ljP8CCT32U138TiJFTqn0bEIQF/AjrkN5lzFCrhw87/8X
8RR+Bl7gwQv2PxlJWCgTwGSzP8+2iFfrnLcHwTHCW+ftV1JVvxAFHsX08hkaijna49fCrf6BhHKg
oVAIYJyPpWcqqphXeVuNWypsrj6AMBjfJskuGJN2xM5meYLLZeQBPuigmMbUIctLSaVng7dsEfUL
0eVMHpmLnSvNSK/ygiHRYEnCxwnetpPl7AQLnLRG02qBjnhpw24cjGlp697W1NUm3Er2k7S5Po3t
BF9HPzKrqGHaC4CLYqL18SvlW3QzVTf/9LcaC7Jet6pBMp3j75tPtTnaS+JcAIG7MLGyQz7rHLnm
jEZ8Bmsi6rdEdt4Vawql6q90fQG+k23lrP+gPNov12nrjcNVRE4RFGSkNw4Z0iPE9W+qV80a+wc+
jqDKyDfLc5BJ0wit/5fWVWNHCN9wZvfQJJ27T79qxxKMC0VfsYG3ikrDiaHbvHAcazNwG3PN4Zox
QQ5b4IN1/plvfU/jNjmlGGLHCAzNrQ7gCpPOWw3tGjTRfAaO5WMmNmyXJEJPhc98PiIjbC8FInkc
ePW2ApxHrTSRQz5Fieff9wDQxNXByPXZPXbEFhk3+pR+99VoGGKQTgu4FtIC0QsXxQFaaalTxdXM
6PTXubpGWjmDZ/9MoS3hZWKIJxyZCyx3SJM9qDLreokpw8tQFDPSyUxNGZEJOWuxPwySJMUtCuJ1
fNt4huu7YxBCdAtbI7VSiQ5IPWSmAOBDC4VZyBOmZmH/l+Tke7FlZhvD4jbQYz+DzvmNvEHePFMt
hr48B1rJU4uVV6nkJ6eK1yu9rkJKl1c4EQWorkfHVKI23hrI3gHAhGMJ1bwL7BCXHk+Oay7SBE4b
Eeju9xoYGRmfNS0OwmkLpSCJVBFnSyimxuhUhq+R0PcrnccTbqyOwM5XcwsgnGXuOghxlfVhvr60
Tf30pHxTVWe5EhpiTzjnMZRQ6Hxn6A3pvx7X5itl1dnWjgIUeZekBLpR48k0lHktU8WSDdoU9ryv
O41A5k9Aug6zwXBZZvv7B7U2Tc5QDDimuvMusSvdcQ8TK9sfwgxwIHpRXcpVIQUAV2tE4D7rJmzl
lHq7SaW3E3u8LZzgEex29L6RDwElmKgzKx9/4KEXeZyPV4b4agUeJ0XvVo67bR+ZoWVq+UhvtZOU
zFFHT1XPZln1PLFxhhEi1ZyDMAUceUgxPGHg6PPXu+zEcbPii++avR6K/TiUHtHzWJU1YvWSZgX+
+5PdggvS3qQIcDmdKtahGLGG7fZUKlPZanY3DHz+TsHbXSBiDG+3lBA64f+Zo5qyiHmQj6kbN1YB
K8i18ay9rghQo90Zyj3dwu/TyKcY+nodvaBjsWQaNn2+sLYbt+/9M/t1y6gVUMYdxPKOldGgCpo8
lY1e9a4sZE2VZ6/RRCoKInbni9ki2wuP+FNEYGsuVOLH7kxih/gYf32VCcf3hu0yfJYjgTN7loTj
fABvzRs9zYeRpfIRLpTHl/nt3GhULJzYVfiKdONncbt0r1IUuB0c7w4tCD1wkWpoTDTMo+veNTsO
QYWXhpgQf6ZQT5CGIkDbZyC1b6I+HBpw8FS3DF39nhN4GG8H3c7jrJhOxfV8VJZ0x8qVNwxrqMuU
bNbn5LYimyupTDvYzudj2WiJKMUO5nfO9BJpJdUUKF3dUKT5G3l5lfpFPb4XpF1u9lz1i8fEG2al
Xws+1hnW97YQ8+FCif5jpQ+Ob6DD8MTITWdaiJoVNsPsEfVXkQcG9PSGJALWHbJQH9Lmvc6IKwCt
gXOWTeDYB6u+IaED6pDeK1QY3Dufk4DvN0zKRFapeBYJgeYX62DCSD6Ysks/uRUkD2VeFS5+h/ms
ARtkQJ/pILlM8kj6WLtGcyrcN3PaPHUhGk9tboEsE9/TyCR1yqq563sizjQAqzFPNlUl6TvEMOrB
v/1mBUNuwpJn6YwDI01xz9WTpqyQra4YQ5zN24R7XZuEYM/aq9JfFdvSPyLufVXedBukpPw9ws9I
KSJ+UrTFh7zQLnq/6u2pL7j1gsq9C9+VFm8vosL0Efsg10Psh4G2wQKVQ0ufC4ia2/JfjVxvEd1x
Wo6d28Hw4Gcc1MGRQX4NQp1Pdxm5jwggNjjkXZUZw0tOwK0OKqPNIDIU+8s7iuAZgURETdtW5/Bo
KQBsPCRwC2QUNQ9ezNyNya8DOtoVTU5GJ8dx2zq4+PiOLs7qNyAomojjL6Lo3MMD4ycTAj6CCGdq
gD+GSeIeU0RLAk0vGC5fLtKYlpB0zldxtJfUDuLio+1FP8FaGDVtTCt+7436ZLmz9N/B2JIpVr3k
PhFZx++eEeXlNNULCIhrVF9AytXFHbn6CNmiXuUGNqJGi1ckRjx/kNrwhVPJ600EdZm8WMsDAuQ7
331D1krr1iAODaGET9hTK+zHgwGislf5BJh9oC0H22aYo4YTCCkDTO9ol2C0ArlyIDCDfyK/igNu
wNEMgz5vPL9QR5oWuNXH2KcXX5NRgE38n5RaH+u7MrMy5p9Qi48fK7YpHtGKsetC69ZPrBG3IH9D
AV1WWohPdfzqpwODx5egWJE2lzW0XePZoMUpUwxU9EUlAYFdaYNWewjEENOfvFHLnSkdpomuhuhr
It2JSuhQBaXEUREhmhmYfmPJ7RrWkmUje+CwQ5W+JF47aemr/03n8uuawVDLdBK4ZadQ6zRhu+fl
8eO7r365mjCce/ZDh5BhPgP3JmTcGKeon4i2U9zZOUkJMaanKBLK/6Tv7y+Z+Ksch5l+hmtevxFr
gV4TkZm/31sR1CeE2NKM+RuXbHcIn8/daXn16Rh9+iV/wFsa1KuhuHRvZDjhm+h6SJMVmCVMpKB/
bn76bn+dKLbebRj95L66QqZhzS8SXlP1rhqh3sbTcTXuVk3QciXGDmQQ3np0j60H2iRIdlx1/6Jb
jC2y0l6t4mTqgVToQLYz6VN/ncG3RjsnWGIsXcA0OJSXmwtrgHpp/nIu3194+FlZq5WgjNgdOlNz
3U93NcoEx9lN63XexFNUSL6FL70GLzlLST7whdyh+qg0fkQI69rHCJoTS2HEkTSmL9A5fY8t7GoY
PUaPZYVVL1u7EWk5T4ZOyjfKwgGnAYC8/mpd8IP+tNQ2vQgTVeDMBnXt7aWoezmQBpSuEDTJgab2
FM/KzoXOscvUAX76FvEK+1Izj2zLnvGHCdrBL4L42+ZqqFyQtu8flZexKbuPlNjGdNOI0BbGRcw2
eqKuJby4WpAmvWq9x4AiTaMFXBMd80kC4ZMmdHe3xspklFhyL/H88C10osthfswuEoreg7HdFLbp
9sTKZQoZ/6IQwePWD+cb/UdQcwTN8yeHoaXeFGya7IGAdzuiO6p0LkwbooHK17YXNosUBwsDJEkN
ui/siWrBm/kNw/PhQwzlfS8hcEs0jp4zL1zV/aV0btsxen2/x3R+Pb+d7eIoOYcA9yaRpH++mpg9
DkPVgcmEw/VYcfo7EOZ1Ays5fdh3p+3q3RorOcqgxOJukvCEKbhYPpJbWaMfi+TsDgpode/LYhGX
XekVwlHwZ7dTFvYLBM0+AJdT4aG5fXGA3D9xpbWZ7zNieNAABfaIJTIVrrwKrlcqusngD2ASlmfc
zq9esV7ChnF1lGuyWc1fc+71os+e4UNhRN78Z/9sEu0kOfUf16fBSXVDWvVfxSchR1VJw99KIRmR
sqAgXR5Zlo7Y7O1/P9IaHZ6TTLJeFWHb9/R3PuwPNltT/WnxwAHhoCJvQDbzuCRLWCc+jrtJIjf9
z/FPBXIQ21OecLVc2hxwQBh65HvkI3D6vC4XX0cTsrdaPx/ddnXdgt2XLJ5KJVPb1QuZA8Qunr66
kiKtue6wQooWbu9gtQaTvdp9wyVBkRKPrOHDm0IUvP7cia3MdfvTPZc+kB8BltO6i7JVVZX8ZzSV
uOE+DTPQbuCLYAP2sIk15gkyjVb7KuTUJ8yLq+MUs2abLBKRaaf91x41tr8jYwvcETnsWW5STyxB
8662gD/uGuVPKRR4TUG6FsDUUm4E/nF5QrWNFfo9cGPO9k7kySFLFm53Un4aThIYk//EVNZZY85J
aaOs93/E6dT2/EdxeijfwwXV/m/YmJ0HTaYEvN+Y7rrFzEpvGi4VZfOWKpOs8mQpDhqbVtx3kY2Z
3F6KBBbC9lLcvapujRZGnRY9QERdeKsN6M6QsX5slhKe9C03TBvqm+t57gy8yCv9DaEq7JnwiiU9
7UZhwRFQDpFWQ158xb7+N9oohpkqE3y6t7G7kNBtIF9lZpH55mpuU3Ub9Z+zRmpLMpDX+A/2Srkb
mOTqLXHwwLedGBTK8298RwSfwN8YCBKrXAcamv8cxJE9BK52hcEmExVnotBBi0njptHbrOepZYXf
WC/P31rJaX75HNVEQN4HJlkl1TwyLwJ3ucGEn/Q1SydJ6uFvJMAiAGPzocSO3yqljtRsAHrwJE6Y
k10rzDjLBhclVJAykbqYI/NiiYvjZnEbqm9rFwONxV6fR8Xajf1E3eqlmvuAxTdnbMxCclnaITol
BmXkjGjGvgcGdeZRDVF0M1WWS1ptXxHcucw4+xKoPtzW8HgJojikiTYZw1RNaeYSsfEbOCJLxnOQ
VMk9rlI7bUOAHdnn2HfDEnmTQOQDoCTMH9XPqFf9FShmFBA7jm/zlLuU0k2DzlP8lZYfBn3Tpgw/
zmmiPKZcr7sXeRZ68WHZ7Qfeflg7Jg368wqTH1TJ7XrULtYRwQj8Ko/cpMOWlyoKjAVnA8MDTItl
XqdyO1gkpl1Qs1/b3hDwpYwm7G27OLdH6+oEIBh3Y5KWlpd9tb7kn2NMnnUgtwLpoRR1s8Q8x002
MKo5L+RSlXyKDnhQXa1lzurgjJzn+eaKyN4y4+yLDGM9m2OaQprztLsg0WsD4H/sIyPJpwyAor4a
1ty4HDdNhxfdkSPRbeH62ECbv2QxqMiK8Ow3J4Ym54M9CmtjIGvSG9kWOAhd4DtQE7WGoCUVMZWU
nEj0DNv8NzU3iD39TgXy8K4PZw62yke2hb32NIlSBjJjT5ua3p/iv46H0xFWRaJmd9a5ZtO02Eb3
ifbfUAPidhfwq0pntGdhWRSvb61f+ljbqMj6yfOAyACeMMNRy6kw7Am5p/gOSdL3f5REpVyfJM6/
p6u+E/NTHMc2JGL7fD2KVqcJ7NhCsrAplB0zpudUUW5Tu8Wp1ZBl5kROcITLCyacctAY9UJIUq6L
yQRyrB2ZbcdU6FbrinIR4q5ABlHK5qArxxNSR3OSNstYo06skAI2QtpYMOw6ra7Q8FW22nOGKsyZ
Lm2JeVkCjeDdp3MXBjGty9HmnIG8GRygMSmTUu8Ft1tlGCs/EEE4x54nurX4o4bDUNZuAzmfvxBO
Be4KhZ18sKyg62rXVtMX8TkJdMUQZaXp0g0J25L0uJQKyyM1MXyWrMt3/8PRTiEv8uyIRNlUACkc
h6mlt7bbFOZMreOqbH5NrMQTC0GtVYe/eWVyfho4KKQ82XOAWPJSh/+HnbdlU4jbUkG7zefhv/P9
aEQPSXpUWquZyPI2IiV7RHvizQi750OOvlphS/rS8fzl/HoXZgLsAqGQbjfyuzjXBlEzB77cQnlA
i3LciPlD9O4lj1HElmGQruUnb7z02fJHiK1O3cjQ7CRdTR+hTZmjScykNwGblbEdsawloj/nafaT
2wzH27K2nuxZDoqh4OZ7/cAK+0BOq5KVtHOhBePOQhGq+4m/Nw0uVH4MfycS4q3GCgduxyy9SsKO
R5r/8tcA+sRKCeabmuQ8Q4H8VNV/MUajeEwPK407gsJNiPb19IonsD1C0lRf+ssqpMZinaXa6XSc
9hAxz9duvr/hgitcrUcXGWiplBOyOa4oYD+Uwg6iAPOhoDuweRYQrDSTi4WvoBuGwm+5Inu7MnNe
5+lKyhwHP4CbgyygAwObS+m/Lh/Scv8B5ojnVqpr0eV0ZCflMM331EiEHRe3RHAJmJ+o2wnpVozc
J6dy13hT163BeOA5JKpf/GqD7yXcsP5XtgZTaLPtLIZ1X4EpheAYGCrZkf5inXML9HsvKNo5hMHv
tFpBjt4ZBhyBy0tkOoF+7rDmEI0UwmMDijIEaBE4UyXeuLExuo4U9MhROhA7wijPPeMOCr4ur0eB
1xuss/fpDWuU3K1igk/zEwbTvBe1TJ+f4CE187FYWjJrgz5xOvmEGO6sOVvqtY6x0wJFQzih89ue
Fx7zolOZ118azPtd+dnGYARd2TP2ADXDYOt5rN0C36ei7Q7N3ntBQy9/GhmkJF5/t0Lt/x0gZTa8
3LGgXw3rpS1o70ps8c+zcJaiJ1PL9rdp1B/Akh80HRmwEw/hlpvL1VtJ+ACyplwgRo129o2/gQjE
h14PSe9bEEOfV9secraJ14y9jWA1T4jk4S/dm1nKRKqaivC5FiEbqZwbcCRH8x1atvAxEBovWMRl
Utc2xPDbfKamtb6B2vZnijpN+gZbAlg8p0WwCjxCShjCw7aTmr0J3RDFmVcBX4SAm6TmcWamM2FI
6eucD2qXU040nJybPMMnauU8oMEeijNjP5mA8595F9oYMtzJXXR7sHemsVu9FXGTZmQXadS1WvuC
aGaIBWdIEhMFk4Be1iXV/7UqnhpJ/1yRJPbj42Vooi+jSNBttlGXsmPh3SMZNK3cW7psEXEeW0/D
UNb9f20O5SpTDo8ZD27GGELvwchDoOxJyeBu2vSTZrYt+sduD96AiiqgjrfyEK/2zMWcyTNr0O8Z
rjHVg6SaT5PV2jDC8kWI6YfzWuu+nmW0I9KLdOAlKMeikYIpAaKToHh11ZSi1nwFCYMg6TJ8gXEL
u1oIe5glEd5dX3kLqOBuEshoXNnRylHxPSx2KDRF5Tv15EyYFZk5P1oLvpBfMr7FhS7UAtbmLC+3
BZ2UTz62P5gpP/1CtsP7uh6L/ICnV3iJl1fplg7NPMRhnFWRx162fzU1ThwHTYV1RfNJAmT7OGjz
Ds/neaz5IucNqWBcTXzMAWm462xLZ9L6kk++QHtEyvPL3RxHPAbjHgTpuOT93z5o53rpDtQxEK9r
CBGp6MZv7IO4tmWlkw1cwYxVVNaRApAqD9a67gp9zDPyQ75EvOiO5x2bS2zqfJRexgzEeleVCC2j
st/f9/jdlFjrecee3k0r8ItmexkZM1SV8MOsh6FgcK1DpbumHkG2zpN2c6MiNRbqSNtr+kTeOjqT
nMpO5aU1erjxqHV+weRL26C5IxjbixFDt/zuvcaNESjDBXGAijm0H5PMOmZmyPa6184pOx+WycxC
OzQdHF3noeuitDGNXklcYE9ltVIkryNGFb1fc01ACq5HWQ0t24x7hNDFibqRzbrt1GH0wrX66sKG
YNkr7u+88sO1+bwS9HXJBrH2tsvlJzPbsMMGy1MD9cGe/1ZLsilZL9G9iN24hL/0SHtpD4tbtoui
94f6EsCDa4/BULPxrMMBZED9htIgGMXKxKgfz/DWgShttVYIGC0HKPh+Tc4fuxyDHcSKJZbVR58o
0QA7IFrQbiI/xN8SaZt/jX6+X8+xqiiYRqv9nkyxvWdjHg4GLvAkBYqZblJGvdqk2Bo4lF/ceWzk
ugmAkLcoKq+0SninrWpkzBK6ZnW5vbfxSZxW1bcwtY3fMkLCn1GAUMkATwdoJmppbWOsiWjIeJqo
9lHopfg+eOfg7/3ZYLcFozqJlXv8XHKkstFvE3OuUqLu3sm+piXiAPRennsPpzCUlT5HJEYj2Olv
hp28PYRJxstdFYBn14t1de85AQGsLCQYxd1M4uT4Y61Ew4dc/kVhTow7c9CKyX9/keyn9OHzUrFT
GInlpZ0Bvem7iglU/evRkpN61NRwHeh2ghL8+DbMndiCnCZjvlPzRQ3Kwpiune22Kdjq1XTQhpHf
kzRlhE9wbEZ+iOZvqSbbHR7xtSQ7zWHlNJS3X/HQYTyUxgs/bvvg/ZQV5pl9yvbpVcW9zN72SyY5
kCU6IaxbWgcNdgOzzQ/ks8aU39zDqN0EmIont34aF46XQbU1rYTL+bnT6uxxqfQgOo7b1fO6fdTY
ZqT5bREOe9HKpOpcpnDb56dmZ2fdrc1p6PBwDt5w8kHOBmXQRkks5tps4rJOZpRvBebXLB0hdUHz
1bECtcSpH0ENaSwjYifAF5MD6OfwddU/U2eBGTU0ozSXTLLCuJiabX+uhgk7YcmqY4zC9S10rB0A
Ake9BMdOaJKNEZnJbuIGLuhEMPYuf9w5WwSeIyv8Hi0R5Etn/Gex0O9Q2TiH7Hqow8grZlltjhjH
LoWTHogTJYIaxSx5iQoehy7XcrlCxHUC7gk+MNNAzwZmviFMXv2vbPFjgTrW0gVnAXHdQ8C9T7qh
cbYI1y5oyikAtmS8Rnw8nzco/JnBau4AM2vCUVB470sgaKUcu8MFjT3AgFk1eT7TV4q+DMjclqPI
7WGRk58DJp8jlj+94fgDMGobYHCl4HpVSEYjIGemYhynFmseOgp90hmGBsZiMXRYcIpl87K8c91Z
TvfmCaW1DVn/KN0eWbICC6/qKEzB826/MwMQvCC2AHocDJFS6H//03089GpmGuBdP++7o5IYGxLI
t8UUbzkTwkrkSnBHmOVTn9KJVgbGZ3ImKd+hqO0LgArDxiWMsb/IBCa4unfrGBZ9FJa7YxkJVCoi
1DuIn2RlGyqXdFS91zFkvJMMWmn1tyoPVo2RLkAZ+vFJSFuKRGN4zILN249jj2uMLmxtO+Twes6/
2O/AbDKip6ivI5iYtohO5tu79otAfcX9PDqE8WkPkpZIiXgmVUribHhnIhlwqzQTfPV9NbW6OyOq
fwpNFEM1tazScDNUfWz2rxD1Y7bfYt3kDgrqiLMJvUBgmhjAdNebjWoH0Qu5/mt/JNXo0DT1zn6a
fghNOr7YrEZeRVmIjmMBPI8GSIQna0JOmejWS2bkeMHj2PL1oylE4iypJbeN1Ho4fed/Ld3i4OgZ
xfzLc6cixh9iRCJo0qO0NyaEF81YZNVl5+Wrp6CDuey1SphTMwCxL3RMSvn8ysM6nv8tPqu4wpsZ
1nbgggj5hoHphpRCrp6rECsZibfonRuRBv7LQ+u+qR72JOl0wWQSKyDOBQUmqd6FYBQVu60oaMLQ
F4+cA6NkPq9qPAl0iYoo02HWq54cdub7sXxo570OYQgF88rx5U/CUBbaFXrSXeQhv9J0c/gTOfSy
HeBNQz9lHBiCtr6Z91Gq7V++a/q3WjwcjWu1RhIAZEqRKW9nMd4QugkjTBxSndwUlXmOcl5P9YTc
+lWTN4aPQpwG8gMIADR8VrqCox50s8oMIoF0HmR0A4KPNQLoOcNDwYVAVdaC89RYPCIxbE5Xzboi
mKvDiTVHsGSioyEMR3k7f2PQI2CYOmVT3KIJ5lcldAVqZ2fr+25XOt3zwLqb9mQSx9QGlMj21UBB
hdXqjaC3PGDxRV0OL7bWb8BZH99hxAPaFwcDNZEKxn6rfdpUcgQV1paMVivhyDasPE6N4Q8cap0M
hTGxW16qwAL+XTgUbjTnV3CLSHOKBBcPP3Mv+mUCymsG5KY2lWItr2WutVjeMvg3AqnrWtfGia2m
oQtkwopi4fLixDiWOTMHkrognpWaVd7jBVDl1lh2UycTuloJzqcClxNN02V5zHaU5IHzVesOuWVg
V3v8Pr3HKV1g2DkGppMdmZzHW+NF3JndEy0F8pEOwAD+EzS4VckFUCq5exQfKClpRRql7hhh7V4V
g2EwLGmZGmOdsXXwOAPPTBVEA1laC/fvP6KJUqmHBUJwxUCJri2a3E0sftmzQRlmHuoBcMWS0Cex
HTwDoPctL40/fFXjrjdsfXjNEWCd8h8eeV8K7T+AuQKTLzknFoGtJH5jTbAqvgT0djy2lXnlT9BO
VBNLv7124+qUERXhl3HQzaxFKUhRwa7+JBv1aiW0ig1H+87Vw6retk8jmjGrxrScoLmvYi/3Uxy9
YJGadoqmfh1x1eAdgL5LsXEOw+yiH3e53mjCryY5T+fHRt6QKIL51jVzjSE/pbCuVP17CXwCUR5c
8Wrg5o37oL+sd7EvQLUDwArdAhy42RHcYLvLukimERBdS8Lu/MPgDom0/D0CYPDLD759Y/maFglj
lVDMw0eLcwkYmQN0QclIpcaJFf8F9eW8+3l7Rt+eKeBECNIU/0m1EQ/8yCeZf8cLLxoFOV0THpKA
R8OFj109gLXPUJ6IsNGHgNmGCfBK91dxlMmfHfDxJbb2DaDpC+S3j32vcEc/KkmNV2Xk2XL1Hm8C
dh1u7JybgX6FLpNCdg0ODzfa3mtqodkM8pnqcnatp+SRwgqsQVdBCp3yCitqGTuLPZPuVg9eH8XU
Ql76+O3ZCJhvWJfXI7dl1phQIYtfssnjSa8S6bPzo7czfGtBU4QBPHDZE9e6ChMz+262+56osfDX
QWKZdTdB7FufmsgXa9w8RrksrV3Au+5wymsF/62QovM/DNRmmC4nKbk/1EpcH3eLfcl5HX2eUy3R
p4wKESRlZPzSrchshAQ8SSLZ7BgL4aaXifHv359kErBH/IpKXZz2gzvsz8ykAr0EE6TIeBCIoBgo
/NQunCek7oWmw2m/PuthjLPCWujjzN6X62XjkbROj0IqazNVM3JLI4Gx5CNGvcrvngHylsfn+146
dTKNufZ1dE/6oTIrzzEYfuxKf50PmKMYOQYMCY+5wLep347bmzEVD8Fc702cKf9V7iXfaKA/CWkX
WYQpPbHUMal5q6qj38PI5ivrU0BAzuRl1nSJT7MfuH+Weic21rmnf1XMx+dIDLvfaqQ7C9d+amKl
8DwI2lJPDI4YmUlqsg80WbzAuLS0wD1tafeUMIhq6CHJuOH7Q2qUF871AnrKDw0mN2/w375vdN6I
clvlVeU7oeSfXn5QZBlGRLCfbmgDYQo3Pi8oNj553IKV6xjFQ7QRVwbDpvT28Omd96jHtSHFzc2Q
XKfCHgxQytZd8p29NtVTzj0AGtE2X6fLyPdyNu27G8QLJcrEJO9va1o8A/+NtLow08tMNk8VQBnI
uqhy3+2XmTUA4Z9Tnzbxjt1LpyMfzQOKVogOhy0QIRxJNi7orMGFvv1JKkQjIflcxo8ZWdG37vH6
I21usq3U0Tj+5gK+6TVkb10LgvRHh5KmIveCiW+0ronBH6IHOGF+XwCF/o8piYmgyIAa8NeFn7yK
7fLlwnGY1BevBYtR9g9+LVcSxR0Fz36e8ffcc3c1IA7KqX6oB7jZ+dzkrFEvnanAAtY8/xtxvglL
yOZNcsYJpb7Ni1fiLQH3wLJiTjYj7mFQgeS9nqj/E0WZAvqcC2D4/4RqRRvI/H1SIbQEz9MTEagJ
YMMW/+yy+RGpJBPXntm4/QLn/9LzfIyddj9cXP4uBh5Se/fgZCwFxOU+7Kq1gN6zUWNCUuXaPa5E
BFrPiArtdt7fxodJXzJo4Iodet99Jzk78QGd3nVppBl6oRvTP21myrle/fy8TGM6CHyKm594xDop
2qhZ4XFW8wmqc875uaQIc/ftu0I17UceviAernJilf8wQ3kG9ZZYRCq9mNtkPccgqajXGwq8m21J
lxo3mWe+vPOV0BE8+sR1I3icxGwldlQjHLyW9XVR2Tt6sENqnMqTkYAIoAXPaCAiHLBvSuesx4Mb
uAsEByzXQ5DDrweUH9WsP1xnvNbOtmQCqSOIgSyjQnsrV7EAc1MUCUELgLZUzsG5Yqs80jW1pCIw
7Xn1dT/u9tpMgJGHwYwbNiP5zk05wrnl1CfUnOFCUTn+opC4wQpMSwZjntBiiVfdBH1Wlr1/fwTB
CRliNR22ufZR6G6/hjvD2x4PfuvbloJ/6p+a8IU+2292z7O89Q9yfMGWFYqfKOACdHSGBg/po+aH
r5jh1Kt2Tv6yayGslQQBgN37D4AO66rKOHitR7GIUDGmaDJcS4Cw687ixnp752dj83o7nOWa/r/d
3hnRYmEErymPwrVJXEp0wG64GCKTQY8X4SNi90tleekz2rJh4kQceA8C1U/k1fH+Y/IzCrz8h/42
jE9AGYOJPAV5cMf8TzQezmOIrKieko0NlOh3wNDX66SYVYo7Y3N3++w5ALWBXDg3h9jameEwsZ6Z
cEzPzB735rZZd1UVX0kMGAaP5BmiO4EQdche7Z37/3/EmYcnyO7VbPgEEvekunDyxrqmQfbRBRpG
itkq5zxCZBi5zGRYQYdPEKCu/XFIMDH6SGlJBOLx2a1FondRWyWMt1FJk/+FgM4EnX7ovNmDCdh7
r1Pyf+qqUxik6lnfjovTg435h8rgRIin2/L/55qYdIsqe9n+yFKBxxs33EaFVfiOivL5EwidUeb4
RtuZN0dzwisG07jzSnYznfveu7KCpAEe5XaxZpsXagmCb/bGQE/uW1h8rKNAzRgK7b0rfQhh6ec8
KmNviGBpFrng1BqDFaza6agq8R0pXtcradRsIHNN3Ke3aWtljNuPWTE0eLqoEjTGd6/c+MzQhBXP
gqUGAJyQK4yxrmCC43kM5+2a1zeqgRekn9sXIIczhUuP0hDiWU5F8/sfVOeuI3j/Cff70qT7yHun
PeTSwfaFcrNYGEJyMgaxExoxLUywhfppxYkVHgOgo7eI6hVOLyO6p/KH09Z1h7dFnbRGCjxgsjF/
A3g4RV9lQkwf1WmxuoO0IdhQJriSOilkT4TW7st7KfpoOZQ2ubY8F0zyxJbJ79iSXisZPfGGSjnk
ikZrxSMq5xyiXxq4z1bn2K5AwfA1MAMKF4r53PNe5fwDn/va7E/T6YJDj3r7FNORvDf4C4onupje
//K+KtmzN9TvJ3Nt0hudwZjYlob8jvWpUO5ZK9nG7w6RJyzDELN3ZOv79mQ76yxBcgSAAxyvw5q3
4zWM0W2IXdlQY+10nuY5VIPmjvnwqoViDlDFBIxDKT2NGhZTTLhJOoRUFy2Ni6xXbL94wBLfHlsb
x3tlbeYECxeyugFYkGLrHPlZm4XFopHm6lruF+uQGKVVn0PLfhunN4EQ1+bHsKWOtESphzXCvFOp
tmIb7moc8xNh770JXLm8MqiiUux6TxNbQJQxO76bo58AgXObunk7wpw/qgMzEctBRMvRNzv+uHUv
O/nk5gcguu2JXjrsz9JwbZXBaw4WhYApE+EtMzJ5m0EsDVbRfX//Ps2/e6R1dLmhXRGbXnnty4NL
gGDhoT1/QHKNcVAp0OqgqyjEob9FFtgCZATPieY9Sxf2gg4Hi9TAscb+jLS25NE5pr9uKf+V7u3e
Ev1MX7JZ4dXBa3AlR4NPZV2z2wY+8QEt6dylLpXIaCYYddPdhNe9M0lwhS2OoF7Yrl4q3/55vmth
4xOefWkEwWjds4RY6zkEuy+s1Mu4fqVkcomgfg5sYBY+3XWMnudgZ7RVMoGNN3EUZPsM35VBrQ6y
4ZB4fFzuOBOhOEVH6tIOS7le2OFwlB/leExWRB/qfOKrn4PyJ+WjvxfwxQHsgGVNnR+/G7/nRBNy
RjyctdwqAm/G0RoztWBAjY6kBkEcUiksAyRDdXy67JC4kgmOW0QPfTFwbx2YJP30aV1NVEmDuubq
uKWLp2xyu6NULL+fYsu5l0Ccr/C85TcZ7m/y7XRtuAh05dR8gH6b/3cDCOmlJu3+EIgibJnlFeJ8
KpCR51uYW+EsfVPKe3kZNJPBX9oLwRlnXzedKqDdiGeE+jn11vogPxk2CoBXP4EI0sG1IC14gyJm
ZYJBv6NaLIRSr7ZiVPDibFnD6MuEosqBfJpmOOQbDIs1kvMIkfo+j7rveXbjgPkPIatHzfMHC2NP
Ti+9ghaI8jcBkpSMXoZWel1U0LmVdVMugkAEKhsrTyCTSeAQPIkIyJDiUU+X0HFuBVN/Orx+T/JM
RiM8zdrAuvQrs54FQSKd0B2ercINtO46wInedBdR8XSTjzO2i4gpqGSv0LtRgChTyqXC8zgqUBRD
BZn5Gd2gXiLohJUmryut8juYS5j3vf4dOlhStGOfq2NY474QycHzBiEWf1eQtgWVpKYpcjHM41Mv
zEc8RBZaguy6mXGodXFgc7ew2MbaUfje2V0RLY/uPujJWqk6qaHcKNGcK+FgnAlvd+D3qSIdjXlb
UGsMe+G/d7aPNdZ4Ab6ktHWuXtqtqx/N5yUqQs86Ja07thFtsn/4jcip07X9YfzTE2mNrhLK4bf4
PD2COX8IeExdDDkTHW9hUg6a67mdLhtc+6LrNw/ZUoBhQca6BMJloTrV2DLiq2Xa6Ro5v2kmubwI
YICu65CFMz+temxhN87YxXrYbMX9u49KyjXuTW0m1xOZcl35pkyKEN9K1T+vTpCf6hu+O7el8RPV
mJ3SryqYLhnjJIjZDw7p0CdeODmLjkQug3KI1gsim31I6T9oN1GKwePcXMnhnKNaPqmvrmMs7lxt
T1Vhdo4bKGyqPgRNX/M+uxKWQdqp/EPVU+OA0DMIOFOP0WNFAUBx/XxKc/e32RFgA03xq44TCcDd
Y+w/CAFqIYrLMhE9QFQHp4UfE/O0i1pPGUYYrEBGZ8c5NnmRVVD1gvUghArZjedDWdBpIhJnqVK8
ZVWllXtAVTUXAyMVLsN6MDb58M+UYzu+0QWdWmNN3kpP47yTCUDCjBdOygZ5glRjggLDGPqZObZi
P9al1Ld2R3YtlDTms9pWOb4j8bsuVBuQ7aG5eBljD+zozXJykPwxNzHXSUilE7iHcHRpVraWXxEL
Sa++oBtsP+5O6r2LvJcJkIyR1iS1Yc2UM9ahkdZiC2LLJpDU3jvjtFd4HxBWW0yTsWGQNZyi+Y4R
h9khPr9ieUyr/mDsFiZja/23dXLZN0NFvQIUZRgJrWcH11ukbVGAAkhoHtQzn7aGt6+PzoAZzvbq
Pef9G4coN3P8ZUNfcOvgpNjpbKKqOmAGF8enWRVZ3LnlsQ38BADWP+ht4zRIbQoqs4xE7iHKX4Xf
iZEOQSg8lhDhpTtcrhtb67/jldvsvFYKWDIlXcrvvx7ChggSPAuFiMThfaKC64QYrVDW3gKHaxWA
MJ3ssdu677r/u+kvaX3IdnQ+hwp3yCOot9uWfAHtPvbOFsiYml7+uuYFSrHQgCQh8Pm1de3TWKga
MB1JFMYRM8geJYnjpZHR8a9kYMjUJl7ZQ3tFFNRDHS39QrySeWZJuBV9uSQF7PYw5B1AoHPDlUZx
bn7kPzz/kHC8g0yQUyEzB6raZhvAajZe/CAEYFU3DZwGOI6F8z172zcKCYRSaWAQAxq5kIKu4e7P
3/fJjnHKQur0VgC8lUhXn1Ycir+3Z79gs3T/1zOIN93IVS+CdKK9wuy/XCnOBU9o/zgMJkHkhSmv
5oY6FHwo0OjcKIUZE7Rnuf2lKpjFu0C44bQyO2Kt1W3w/URaQ+SN63J1ZDUNONYyaWh/ayuxBbev
qfo1AdXz4Hh7eJsK/bAkg7g9778rbnESVDcAthF5mMhSC4kQK5tsTqG6ZYXrQeHp9T85X2eUGU7V
fswtKfixkgGOci05qApfsO6o4PlMWiJ/R4Kvx9vTh8P/E0DznwL+6kPq02Kp377/P1cgeAds/N+X
7te69u2RWyjiHbfOgvoJcAYhbWaTwlpzl3zOD33ldi2/g/+0sN1MandwU74+380jcNLUtFdbCAK4
v7FEJywni+szYKZNAqttW1rUzfb/qyQBksxCDxudkpG/xP1ocFyXofjELXeooMBnuuhuzE+KauSa
E09bmgeDCQND7M3AuLlIQ9wBWIue9IvgIij+PoS3npVwxey3Vf7QnSeEOSVZ4mG4LsCgDQPaRWsL
aMJOn1jSZHNQXfmd1PEZIcmtwKgKwm58hNO3NQn/zVT2bUZGBqOXSvtkvmy85/JBq+u2vgayNAYZ
c/dFrRaA9tH7SrWfgr1pJfAJnpVYiwQ8pA+h55BsetEYs6WDfiIyagS/QFiGIY2HgozcWjKv65hG
l2XW3YWKH1E73+vBV2C1/ES2m+BPQEVd6c73PXzJTlQsRno79w23eo4G1KZHYuD6lQgXpcbC9lO9
IDVx7Oo6s6K2b0zQpwPY8Ld4JcEJ8L8P7GTCOePmh0+SCrMO8vbYouWIwheCMc1BQ5QFhhbWT48J
i+6k593zRqgHYa0OKSMczZIOqQ0lKIwyT9WI0uSGR0BSzrvhzEPy/yvKioxgEj/MZuDroop8VeJM
o8aCK8fCxnVjs9iTcQwJq6z7Lue6bzltdpJYJlHcqmrFO1NIojfb9BY5pLFyPXqYL8isIk+nxd+2
d3GHKLrHb62D02kWQWUkY8xsMCIHgb9kEGZA7gfBYtE+ffq+U9ciUfea3oSTbJoGBk4C8dJ2d6Qn
+guUaekC+9BF2/V3AsJKAnvfQl/YJC1RTflxVCC19NZQAGp/fKyqAdpjK/N2OyojeyEp49ztaVJN
w50dCSGOOuAQ2+MUV1JG+EIW1VtMVV3frfm0JOx34NrLKsSko4hoqRG2uO1zByIE6vQ4FUS4fL/Z
x49THuV7/xW9OZGXFJOo03t4qVZhciUSow3yjcj6xKT088L4rFNRpd0GLkeX2DkU1DMZGVIxOW1z
hLVRzC9GbHr3I3jfV1Cn8H/ddLGhvPNs/6fA26eTfrAZEu0EgWDcSgF2ByxH6YYmun7hvAlvbm+b
VuyAEIBzN5YNCdQ4GFYu6T6T0l5ulcrAmHXL+uh6Z9NWsRo84ygfWHVhbUqurhKzy1ZDDOuN0Gcg
lAx4QcNfYkzkhw85KaAldokbV+l+dCNl2FLUFYPVUXtqdOY5CW7MAdg5EX9/8wUvJ0B0lguOBBGq
XZ4UvpdA0qhiLYnBPe7jQGYeN9U1wf8KgQG0Ey6DcHApUmISFBr+S1FjSICOzWZZd/XEilsV8YcH
lWg3At62VJHG9ZsQyxWAWy3SsIqRH5bkrq1izPMjVObNMiinjO48PcZQldF/rowYjE85pT4pUEjb
UerG5NQr8qQ7USenpE1oAgVbdHwGaXvzJkTfs1Bx4iN8MylxMZPDn9wpcbvqhBZUKHBeV130feKn
ShTqrsyDkmTThWUrVFohdpFI/N4Lq78X5qzxn3DJSzT+1D1nWMw9konimVTjIM5VURC45ZWnyxlW
eyYEW99ZVpKCUz4VORGmEbN0wS7Ng/HMrPd5HIDNd7VwYp72T/Dumxn3mHTDKl9f3oaI8Zdnsh/e
/v32qsxj3ci8hM87vlja+GSTG4+pXeh9Pm31UtaQ3XJaYRl8aSbV8CHBgl6o+kvl51YbKla6QVFb
QgtXLoJVAx0leDS7NVTxWqbTDJjrnrqzFbWZUfGFQhUEPcwO0C6pl+sWdJcNWBNrUe8IONIccv+T
Kjr4d3g7ABsggXsk6dks8l6+Uy4muNddvwZ1ViAHysF8l4BnNTHICJxZ5kTd8gTJRbATz6gT/FwF
wzHErHxQL9qFx0efkDHA45cSXoi2Qd7wHIyF8rGbVN5G3YKhYYqTclLGRTO76dJvVuLlIgy19onj
/cCJvKlxPBSy2ReB8HM9POVkPL7Jpe2QFZ72p+lwyiIQ+7HaXFKOzq6W6/OL2LnioD6S6SkBQaZz
sOBQotrV+soHhCWNKwkegbojnB55aiU1Kndztljb6YKK+/0UBPBZZ1AFWHOKW5aUDbZx0RAFIWdP
gxUBHUbel7CTfk99LncP0TvXIamed0Q/gjzJRaesuSMKy9qlJru0NzG8gKiSpBPYlX7JQ21G1Ywt
6eaB0kT2EUJk+snRRPDQ1rJg3itTUoKrWGnNHgAWATT3wGC5CioMk8CnxwlHrjn9sPzQ95M0XBWG
nz830TnDjEah5tnkdgbOCbuXl4/2SEdD8OWyGfs4m7BheGgcPnczRYuGpX08tNFxfZs9N4wZZU3P
fGvfnGdm59aMx51gPysg3e0LZXJG8ljijmVFgaZGrAO3/yuPDi2NpOsM1UH1SIjXVRIrJZeMJY0Z
A+Bgmk6eRJczpn5cUmrEMSSxtvMXUpHM0tUWf7Yr1B/z9wiPKl3sTsEgBklkz0TtX1HEzZCJXXG3
oV0DNoY4onzzdGveAIsJK8XPArqYkIX7jTXh29Jn7aXEvE+o8rsZCGM3M9qjjMBPZDcOEgGu4oBL
PVcwcpag7pb5DNWBFX1ZkK/02QZtcPX+Hi08+bW7ih6p5FB8x7/CCKNncIpmC8bb4k6UgUe2ekMY
DdCnize16eR77aP2gjcBQP/9PnQL4TVvqBhfU7klbNmQVfZeCeBLAu6ZUt8Sb/J5QH+4QY3r/oNt
2GjEBoRI8f5xXyx3LUNaoijEZFzVAA1m8yALtoJfyhmh0AAhSx+qDcifuQQP21XsCQQlAdd+Ioxx
7CY9TMbM5TNh583atL8Nd8ivXFTcQcgKt+8OmFfmLLmyFIEKoKl/RoWMeyshFL+AeR2bb7ukIR38
BS7+HFMMM6i3pxeKczUxeCCEygJ4oRs696Fu2jvvPKbZDvsp6KXdLdnvV++rSdauoNiSkce0S4gg
39oBL7gakcw+pgcQ1KFb9jf8ummnkI6IxK5oO1XOEffnPWeq0F0qNRE72yjGZT6J3r41hQ2WIh7w
IhiA3oxl+Dy3OCDG7fLO8z8i3UsomRB2EAJRZjHFli/wnUuqWodLVirkjViohxpeLM39z9zv8tIx
VyFc95CnTbmq/u68qn2SJE+Xp6GoXNsEgtSxkuNhtfHcT5BRlL1v+3Keqsoq12T2NGpfua/Zx+Br
Rbq+3zqU2yroxvcwIw2unfEOO/EjKcr03GszcxduhYT+8GLXegORMq4VECE9b+ntDPLjM03dpXy2
5Gz0l0+Jwg6LOxoymo0qsj6Dut2fG3swXlp5TzhQPkXsdKxNesnZgzlAqqZJHUNIhNj9Gm25FYTD
MYHHWLPjqETn2Yh2jSJVAaBIqA9ML3JJkmydPTLLZ0WgMmGZrithyx6ZSC3vXh+j3Sm2ktm8BmW0
eDSpNwZgxLgECdp9c/8bGrubjKhJ5zY5EIZndNWl0Zj4fD+Ua1u4giyUgj924tiWhI+7j6YkhNl8
t/XDD128qSj5EUd8e5IBKttvbieHEDNLmwvBWgVdFhvpt54hv4g3pU3cWvcuJ643jF0vMZmnCZQn
rS4HGZwo87lWGITffhUGB0Rj4js1FGs5GP+7GlltvEdaQmdJoun08nZGK91lLcKS7fomPR3Ulkc4
2cR5b509lKbc9BnWOsEP5A25bAdEdVCNM7ZBZzjYmqvxLppubL5g7tW190FFGmSOHsooYofCFzIk
xuHXLxqDALrneo/ZysUcu9bAtxkcAJM3QHbixg79jPv8ZlBjhniMClWhhXCcJA6qelqtiDzEBlUU
UVgFYrIMdkexBmYlNlo1nZmyaQa/+RVWrxfmJR/9Qb5s/FQAT0NxBcqyT2EOdtW08+RymNqbHL2I
2D69hRsCChu//OMAKkWCcmICQ5DnHaFpBwyyZ2sudReWIiOqz1s2c0fKx3bqeSzjNbCGfpfZoVtb
r5HjAtpx7UOVy7Qkrq07J0QQyH9MrWfx2HEPwH44mb9pl0ggcjMdhvf1AQ2QUmYFG+HNcMK2RDBQ
a/HoQDsREPEJTz55zoOgQLV5DlHW8CCDRUgenc6XEnR2GWEnn7D6tPZ5xf54Ze7/DsIWw4jb0/UZ
FoK56eHI+cUKa4+gEpdX24bh7JRsmlUxQGxmZcTjj4N0I4aJALaKoFJPnmir1q0QJw+kKZD6Uvp3
tiekV857q0fcxxq6WDhhtAWUxgSXZTZXmCf/B0c7GL04+Nlj0+3ND2frV6MYF3IvZUsotSmDASP3
3/ou6JRu9Qyr/GyOH2Q6+2KeYnuKLD3zewNowrVX4WPu+VxZX4MB2gikMxwLRWtKAfMxCKmx0JMu
RWshlfxKQoxEaK0ZqP42owyRFohImavp2EWXgvjJtKI5jrl4GqtWnxL6+HkZ6DNWv2fHQNYJ+vc9
Kv++Kr5LR/KB+BTBT1DvU/owY+3VoVvj3wb9N+hqcpeedJvNvlaXkiGgm1Dy6SmWhQ/EIylqBLgZ
1A6ENh6+xBTpsBOjxA0U9eshVlieBo9ArDfyu9zByYpIqcUMKexu0chHQ4BTYwApKXB9NAgeCmE9
DzlndzCKiFmaBM6ds9eymnAe/1K2AAdXhHG1WgbnF/n63/hYxcvo5S0O8ojbRuaSJiqAVVbaP3BE
EAOcJQNnMtAK4HQ8OdpIQ8iCLLMRUBeZeh8V95C/bVAu87SstheFQ1NQzBQ+01WfDyrcul25arbq
RD63ie74CmkgadOGoAiITspvOxxkB2sjlcxkZjCz7qrO4YM2Pq1W+LuRvO1unJYmnu9Q0rqMFcZP
S9dkGmI/Bq0+YLrZUZnzXWDTVwIaFshFHfn9M9h4+7W2QTGi5QRayx9TaAFBqrmL8TQQUkbNYUrn
Cm38KUWY8c0PT7sEzwFKxsH2Ivqo4tMWcB8Y92Ws+GosSn+f+KqI4f9ZUioiYmFQjatvhibs7xim
NigDWmjCNeXunA1JlbzAAtwR9qHozhC/YfO0+toVgcwxv/RYcuBUHpMdYPEBk5EwVoJ/WCOI3gGv
2Pnq9r43AZjM2NpcYq5E9BMq+/HcvutX+r6RhA2qS5QKC/P9wCOvLiQZmS9Ywby6wagoGPnrU5BU
+nSbKFEQ5fwYMGB3wEw24PQI28CBDF8/LJK2HrDoLLHJckjV4fLLWxwY0i7Q1WqBP75aavEg8kyC
NFbRss/ZG4jU9nhqOq4y0F3i5O8yuBC0gDqkRNw0fyw97tYovhptGCE6Y7rKDg/nEYsv+2DJxT/q
pyA89eVlVOdVbZ1jLtTA/YO1XNbXskNsnIo0syYcvGDedn7bPFt5U5dy054a7MCXp86JAhxEc1mB
+PePBje1E44bl4Rl2hOvkjodHUQodGoAxbuFMlQxeSzcU/YR+MS6LJpThXtNnMCJEp3tRl7WVqSv
IRinqQiT4yVHukSBy2VwxkSaZiaC/9R9covIzJWdwPOtRVunihZsm4cjnBsOWK3qDH5DtWhyvGbk
dgG1yjmjYk2ToovmOXRDf28COPSQBkDNqer4/VLt270UzpBy/oc8d8I5q+jt/1Dqaasuwmh9++Sl
at1FGlUqLA9k7H2WczQJccKs2ZTkKZE7ijUHVC2fMVQRPlJhqpLnCzyQU6+7Jl/vgT1GAzsNvV/6
1rnXqc2lI8CIlG6SwFPWnrwj1Ca6e6BtlhJ5HlOJn82Sxlm/hHhbdTYQmC9C+nsS081x0JN80nH+
n3oqzd0+L0m9Gl2h59UhsyLOmA/SylPHpaBH6xzsTpwqSkybuw51WiuVf3iRGvpdjG5hCqGTT2UW
aBs+8XMD/spQoE+Rxxa1bK4Q5zA/9sVm9L2T1ntzUKbosG2NoBvLQRPMwEEatcIJMrsenIIkFtJM
17uqNiLP1kVcm0cTxsMjhVWUeGDSOA+ZReyI/5my3tnvlefidivM34wI75S0Kk6L7IGphOIz7FK1
hfS9oiFkpZT/SLipmXsHW2PPQdB0TC2fI3pX7ZQvLmBiCO/S3BXOrwPrSQzEG+IcqKgAqRLswB7p
zN6HE27cXekUF/FduCmhC/ePNAR4tknCFNjtMBQYkGx3kqs+MjabBYNqMRJB5CIh8GVPZIlP9koa
ExM8geTKXnzb0I77+Jw/guyqVyBhCW+pqDNPaXFJsnQ0t426LTke566dVbqnpVwFxsoEKLCQzitI
fRMNUvcvncBM+ePf5Dlm7Nja/7CIJ++svg7b7Vt6aeKoGxjXhKfIckmQun4AKc4ueiqyqHP9xBCR
1ybN/slxsZeN0NaeaJxYfhfS2tAcD6omYfHujhyNENNSr/lUsJK7NG6aZw4IDqABR0G6PIaN/KiX
snKD0J8vLl1aEZzqEG4gPDcEzsmRkj/H0AkHflzfSL3MlVUhObZcvMcJeYuIuVpf5MTbqgumr7a7
BMg34bSN7ELEjOgg/uh+0n20euJO5m/lapOXmAEepg8PpC4H7rwCpCppgf4T6mFncB2iEf3PUULZ
cA4yFp6cMwXcOU7TLZ0nFTpXZdEoGgVSrBHRi3zDJnxj9LuFNPDB8XErRehMSSnuS0nrnW0JHrQi
zEzAC06cBwK/uLIz3zBVPqthU47VGLwJWJlxcEgzlQaQwq0yhJLM2WG+2pUTyMUlmC7KZJ7r8oZH
rlKpdYH/jx99ucaiOdHxvMD11ro9Xr+i8eUrYIS/MICpwnv8l76sMB5+AshRYEZBgD9bM++ADtQY
BxHGYQeSjBoGC6hK/nJM+jP7/Ipz3uzDpW1kfF1KwUVqbueSK9ERF6gTJg03yja+oPgqB56js2oa
jbkH/e46Ab5tSn+OvTjh3c4Hpi0V5rFP8sL/F+aYzwUJ7Jx9spPiQ4hW+NClLnLKYQzoCWslUbkd
woFp5/DbNoe55jPbqJHnRmm2O2Cg3lEXbyY0zVxO+/WDSIR79Kb4Z39zAMgpmr78zux3QgVNXbkg
c2gSATN9RUbaO1Y2CSMmPyiWd0WFWePV/FozJ+me/xP1uIMcvfl5R9fLQAM4mcgVJz1ycCMHH5nm
36oREwZSFwI6NmJIxcoq4B3O5HpL8E0r7snf2kdtYKTp2R9B3u6YftupdFWsOOy4DNv+dvgVsJRQ
Bc/odAbYZS1NmzQj3wfqtk+0U/8/R5mItLzmz8icN7kMdEcqTIsFJRoe649iJbDIpDCvmK6R4/Of
YXQq62lYFWjfVBlwhj2GcSBeuydoqmGD/dSJTr5f3tgKwEgON/25U9oqO6WNEbCbwDX39wQNPzvH
PdjwxC1y9QNPNAW5zYGD/yOohz3hjGrPiUj15WTEHJDYnHScJ0NEEJmQVyQCUwwzSvp/Swr68FfB
wNDeUDrgd+1CD44fiTlNyAc1lapMK68aNhxrdZOmMb3H/K1VLIJP3UqKc9GclKVMkWx9bTscISSB
LG/3Qo1B/TVlT5gAVEv1s5ueEKRbtp35mTXPa73/LX1ZoKkwYNnElAqCvwEpkYQdMpUuYgpbuC/P
6xrrzjvsQWUHeWlMNlVs2AOR3s6DRG5FBfMvMb3sUL22XEu9zQa73zvQA5MbgN4ZRCO5hcz83PGT
BmPcpyGlG/cr9KpYvD0+VHW6KUJynD6GuOdv2ST0jrSGLE5rBc2UkNuppKC5OGduqIZaQZy2Upei
BYDtn1R3sAsKhdAxyOowHxRpf+RBssYxJ2TI5jXPOr9JHBqI6giJbFtBYNwXG2EcGsZB3dnneqD2
ptNYIbOkdy1HedA089Sq5iFCN2mqRFiT0ayxfOrPlBr/4txvPbQ+sdX1GeQh6rZ+dULEq7iTZ1Sc
yqp76P2hIARfXQylKuwfDJi2kxp4ldlHIeLRia0uTzIG1rNXCT+8Fea4Mf7mWm2MwF96ntgcPz/F
9Xj4Df29ZdwRX7Kze97jf9mZQc+A+r9n6dnslFNQjQQH0u2E7PUIMFfMMu9Qg5ahwdlpeEJwX5Y/
AopbXNW8/cRysTB7iCnw9bJLs5lGhzzGaygcIGlWyDuaIxNNWJirz6DXkGjW9HDsZwlzKc8x2E+a
N2QmmqMrAazKHBZ1aOFHdymUGWANc/sKuO7lQvcw5MHsVoYxJ1fnE+wd6nCXzcqP5ZRY4UNpsvu6
Ed8lNyaAyLfGjpkLsj9tmaD9d/K/ExedOunzSaxLyflvH0XI3H4St8TYVJglJrmyAp2RWtdIVD8c
7bZujS8PaH9spcTFCX81guK4LDs9T3CrXH6PyMOyOj+XqmActWXwM+9FLI6q7qbFBAuCBkYlVS8S
xWl3E5FP6d4GsUwP54YBazfmLAsP596TrGwgAyshhl7I+1tZPg1pJRZ6ZWD7Tk+kmt8PzJL0bjEG
99+4L8lIopqvwLM8YhrhYfROCTQJEIuu6tVunefkqn2o5Ufwtsw0FsF6u6nJ5CSLD+Qe9IeI/9hJ
Dw5VCoflm40y0MACJIL3ng8771/qkSS6NHHKlqT3k+4JE3nrnDMYUWnoT4bQM9BbJkQFKK9G5DrN
BrdHJf1yF2ZRsEGXxn6cUCAFV1IFk8vn/zXoLAMhvqO70VfxB3lq1IaxtznSEnFFyh8zCzSAqSEE
yIftYz1uY4VR31emRLi2jmLM7MiW/pWGey67lm65ZfLMFyNDURh7pdPmc6HrpA5shNjTY4zgm5Sf
JQpXj0rtD68fWGHMozZA1oQIvrnN+EWIauQCOdG104qdofMGN6GNYQJBZKJ5Ap+EYeXPgk3viWlH
BtRhDejklCtPjZbuIzqYsag7rXQYlTsEr4AKnKitU0hCVRyjlx1HJDTY131t+2lCLnaDJgH2w8F1
YieAyOLj7j7d9VSw7ZsqGOEoR5x2HlpS+r9czh6zXenuKjTvjpcOjE6tmqBhs/2vmpMzA/Y0/4we
cXkNxGXo/C0H7HxRsli3QKs8XwJWlERz6/CIWbVC8iIB4q1VY25alBrikOY+FXFQ03Fsld+k1rWb
H1P0gR4XodhJYSewKOwbtM7khIFUA01iW65fT5jqWjd1fY4ha0kAkdiLqslaOP1SYi5T9UfY6V62
7zq4C0rxdECNyjUpR6LIosU7uUZS2TknB2pMPgv2KiuZfgmN4CI0+6vilrSC3UbhWLS6NP/n7FNy
dFTENwaJHTC4WutccQiN9TVSLLOXzewYVKpP9o3rpD6XJwA2dcYdN7GTwfUXRb1oRfOPQWi4SGw9
lcPhaAQynEvH7eHpCW7rf4GMpVrQwcfbPQu1GX2cmVBdeS0PX4bldg4J6726D4c5AsLI2jDuJY37
oawlA7/qNvlu26q2maoLpllQ/+/SI63rp3swWk/aH/ugLTxl9lU8AYZr2aJ2BfXIYKOzQiHnvc4b
bFB0aCxCn31AaJa+AB5SYaqZMBIgFIG0E6Jk6WGOKTFBDO431jkjSP5h8ohq/+qM4PEQf4Y+2xC/
fgUXBOBThHMIPinrx3V5T5SFpaZ9jy8N9hIpnWEok92obDnbb5Sv0bHcDRCWHKz0R9Hpnp7tSosu
wrjtg9BKLurdP4NcIbv7wlCDRKrkt6H/fVIfAJv3Lmn4asjvGQKwUPMSHeLC2Xkyp1qCiA9xvDAU
d72OmYWYuGVc6Rx353opLndspePz3oI8vQvsGNS8tlmAhLiyOon1BCEOMFlYdoQNLg32oLC5gBB/
dQ8Ys7gHhk7n+/288ys/z85tV/32u6vmEQ0WZ073wNAihKTXZQd9vvncQUG9sYY8CKXKEcNI11Hc
3si5321eIXhT1wTxkH+XVH0KdPGF3kO7c3fTmarya7oKhVhQqmgzhhJo3wA4qKauV4Drbm7rxUxi
/6CmAN1F8CLYnbI+mJprb0OVaAklhzhcHuZHooi2YMvgymEyW63FeDkFLFtb3h79kNWcfzPh8TBq
/nYYETwBluGT1ncoth2D5Maa8AC2J8Wx1UMyAORPKkUx7uNZmfPXgAfShjI4hilX+SIrrad8siOJ
oFM0VF41cr9TynEDzFtwoZQ2CptseEUmmr3kyuQqxvo+BLuxES6GolH4oLYXoJji1wXvyX9asduk
dLpps2y4bkWiPg3iAvwQPf/VkKfXJXzME8Ago6q3tZkPp3FQIM44lYBo25dudYxk6HblkH523DB0
ifjKobCeFW4HT8uiSRVRN9rohAputBM9VEkWi2p3hRHoJGCpnRPCbeUv3K4w25Myr4DPnnDpIpok
Ilq3qKKfYx6xXcnNz1mYoAm/2hVbvEgmvJpL+wElpI+/2PwVyo7PU3qwAEMQQBXH8XiubUQUKCRA
dKh9nIosFiqPRBQ7uGD99J4xOw9LbG+f1JznhxwmcW1b/IltYYgIHd9wHt+XpHVmYnELUa61xvU5
ya2nr+0VMZs1qpbI9C10cl8MTfI1lymQexMWA7hLKCgELsSJxxxek3HsrwOxbKneiARLahkfGcPq
xcJA0Ing3BEydlYpaxwiH/Axk/y/nT5SckqR6UgnoxRWLYFQOiSdN+Z6ImMfRletuxWhLMr77CQq
7pJ+Zh3MFq4FzrM4spQ8zH0iBwXeLkwENgryEh+VRc/vcE6AkAqgaGJsBALMU0TGdDpf9tzCZ4ho
mWEj4dhznnJ6dOogCydqy/BuUDjnJI7RS2UMe4JDAHyxAVdYi96zNZ6O+zGim2TFz/yaGJmHdovL
J3BnFYdvkmqkzGID6HB21NKE1JrKLroz1f7IQgJ+HYdVjQazHZN74hur5bnSvzpio10limf1bYXF
IhtwmjVqH02Rx2nys6AiJ50N1mm8mv0dzA8yljQ5/OWoAVVQGQxNF4bb3mb7jcd4MWXh4oSekbAf
7Mupc4P3IY4sTbPnoxsuGH3lYgzCdFVmJ4ujZHd3EPGMfAgYNpX7Et/aMxEL7i6m5nWV26UZVBUE
Fwk9NgKkmLNN4USeOiudd2Eonn4lGsVB7ojqezQLxJupwKI20VvIxbQfq4fg1uo0/VWCb+Cq3isp
eGokHBcoqIe3PExX9tHwa29/ZUygLZSTEzXDVxDRp4PPBdIIpWN4QZyYMstZ0ka2awhu0iQHfqb7
cCYKfDjHUNm5pW6NFTwhzbMDJRiEtRO12U6uPJz4X4PPMeaDbpAmLkfjt6ekBMdjW4+3KM1tBcSN
9mvVNu801z0RiegtZKQGeDwBmw4PAcEc86FLbNw9zREe7ow9UqX22YRBtYrv0NlAKwI/LXzXtUaj
fJXsaLBtKaLFryVtoxqyhoUw8fYBe497HCypO8tCSLiU2/YsLALq0zCK3nWyK9pwcCxcdaSQ7w34
Vo7aqQUR96awmX+uom6T6kOyIp/iNE0m6Iq5MMwqpjEPz79O9bOFl83R2oSyxd61onxD+NYdg31Y
EukdbRByk+zfc1ojwJIV7mZ5NsBK0mshWcwFwmPMJR3TEkR0+dRCDeBh8XBAkn2eGenkoWDPlznP
hlrWAfoRm5CJG+jb6rQSGhzQ9WZUytmDWdmjd0IK92RYFW9c+pF3QGvXB7B6aF7sT8HU2zbQ1L3s
i4aEtuFRzkU4F1bKiYJG/z/AR2/m1p6R6B6KDGTsVAdjXX59snIpmqFDTa5fpJEVIu/q8U2zbErp
Lp4K2bnNKQ6zqKiiArZQJQGh/xq0r/glSWKTXuj+e/Rp7tl+GqBb+2/IuQlVvvcV3gs487q026DG
4eq4rOJUcHpMOJG9ik6zd4QC+TGMYl/4UwiAncZFUruA1gd4JxwnaoNjJ1Gi/etthYEZkAmcGY4x
4DVUzLkLMeIDQ3DjonWVGM5uyXvnf+S0R9eVlMKrgA19a22f1ai0zvke3I58zPpn6zfH5gUF1NDh
nXhe9Bi76LKfpPLqB+ozBH4hogTL/UB8DClYAX+Qo6PmSZ2bVzBObDM9Np/k+MILjx7ucG2OOmN/
eNXmwnAoQNbMXC+wGh5qiWqNSiSp6+Ioj+Q++UI+FtXOS0MlaK5itHpNkkUlsy/P3pklou1k+fxJ
jS+NGOp9xBc3Z2FR0Txz2ynXlyKTjCpDtFjoN/m2sckSE/IoRHWoEMdfaFU4kqEgVe7b1A8jZEr4
gFotnZPNGX1t2fDgx7T4E27gRZ9Gf/gegy0QsRJWoRlz75Pd+JmSZuSnrwzB/+4TC0W72u8BxhHM
HHuA9v7eJNnjsLpfXEYNaJmCuxkRKmaE0l8TAJE9q6nPTMF3oagKQNAlHK65n6Aod3FSrDGBG//r
ftDCkJ9lAH9ZPCEy4nd/b3zhO7L1EWidmlyK8J8Aqm+yJNGkziSW03YG3ouXq339QALSy2ev804s
DVp5ZTgryWflaw6YEsg6wwdGINR/OPWL4DVn0KVt+flXDiceqRNSZTqlTpD+y4yXQRqDmAS16InH
0VuWqLfpOPlz38aS6tFp+iaX0YRcUf8G3uSdw8CAPngTMv1z9uVNJHJXVCcrKVw/AgNJoHN+SY+U
n3gJqqdV5QFFQ1sKmfjbLmP1v02hjD/I8ap73N2W5ZmQx6HhDnNi256Nex4rROVJm3oSFD6uKjTS
jyOD41/k/N/jpys9Atc4OWAselV9m98d/Q56JCAPIyOSCGUmm1uOK+5crhYoSCZyJxAuRGx4chSS
EofOvosb+0Jw8sbmCqQwqMPQqkuSM33FhGo/Mbwv4Qk5XD28sosyO4aToCYesYh5T400zS5kDt/B
f36Zqo+UzhnH9ZPcN29IcEXrd9ZMST4GJODQQHsTsnkvaD1C1GwEoBNpItYDNgcgTGakDpWp06rd
gwkYuKbvpsSlxQQJDGHWeZqdIXhdcg7ggNgtiqXb4PpEkrLugtJxbGPIbZc9LiFTLvG4jMUAYoS9
VHGVJVpYrUuUb2lSvQ7IuYI/zL9WA3D8mjlzUeJSlBC/N3IqfgjHQSaiVL0JO4NyDWE+MpGb1O2E
Ai6vcpdtLtVsDbiBl1iFJbQYxD2uw/oRvyLh9Mp5Qcbn7QEEeAMChr0mZ8+KpWUF4DrpHLhb2UEk
MvgQ9mpR2JsXQT+vQhZ8Ki150WqdhfdsGv1xS8s41xQ2wyrsiQfTzLLaor0BYlYSHGjMjhoevy16
NKsiNKp8rIqBikZU6JKxPEA0IvYm2Fn1eB3D7O3qd2fTNnDSpfvWRPBAuEaMqGDV1LaFfJYmP4Kl
dEIOqzgk9Q1WMhZvEg6kCigHK+KS6/HpZXorT2l9jOHdy9gnrPizLDLvUMRBqkJC7jEoYwTu7r9S
f7PE7LsJ+ziUuDvSmg8ajspz/xfqe65/syYZxtMECZFIjYDBUivbgksSbFKVhuThtaN+JfSRZuNu
AfSSWlMxw1TU17TI7kItW/MYegtPbFJMR3iwmoPTFkrGgO7mKJKByf1ewOZmRn/+X5iwI83d+Qyn
IRTqkMcJFyfKWXDW2hziSKG5t+PvWLgmqSeioNay1ygbJTB+U/+QKk+mgvUDhGkDLDmA6TdmQ7ug
egcKOh6AWwVxoEgX8R0FXvaF0803gq7J+8JwMV7lGmfJem+TMrKxnZzXx6T/JSqAr0WrXorJrxcV
MY6HBpfgrvax1mncYKf9cfYGyjIf9VSM7wXnmNu7kPdWmR9i3onmx93Pi1lyP1Y8eaJ9MRZb7eey
f8yfxaBpJojQkgVhJ8q7APr3wJoTXNCADzaiA+uRggRpxuAvpqtFLW828VgO91R5h3JzEM9uf3V7
60RmezKUPfJTxzgxtrxS1v6NTECqx9K2Lbs0CULsQS5ZJbM2f+MAuzV+An5ORJvCjR8OEovIjy3N
OH336cK03kEypAKcN6qeVKv5HyZ2iea5FxrwCZPbYNHXuTI+0/RBhQzoBxVLa152u3OsMnV04Qfy
vnFIjEs+YLoD3j9tB2k4DLyOLF+adkI1IysI0tqPEenlijv/WEM1oSWq9kTWYaXP2dm++jwazmm6
QyUevVHVS3oKeRUxzh5FTMT+4aJL4zZA3TiQw6dCLH4vmm3Q9hOavzIpeYFyRTxg6nlTNvaFKgDT
ICQJw72VcsIO3ZAQcgUaA2JEzbmQMDjW29B/qgBEdbiy8fYjEKrCuO0Ah0nYk+C5RJV50ep65BBj
FvK1N7oc3Ro+Wk3fD29ZZICRco1PRMNwfNvg8KZvWgQ68gekmh7DWquhsZ54Tn0vbi9HQmVkol41
LSy4wmQn9cmbxojAuR6iiLa9GYgo6ZHRh9GZ+yvuve7DGrI7QFtJIxHsOTF0FF+RRsF5Qw3GChvd
eGOxrSW03fdpx1VGs1cU6m/GjUsFyrwyxLYA4DcN1Hl96QwxKj4dlL/kjVl9iGyGHxsVP8Jq/W0i
ADgAdvaWOC0mhNBYZtpnMOT6h00cDbBuWamN/MljL/VHEeE3avQJvC18kQmsblmYn9mUQPFpUmLF
aAi7A3Cch1NSW/pxfrCczwlp88M827nekRz2q4qPVFnbXvZZuJlvyIayrEVi/u9foU45ZV8nI1xk
JQAhtPIto253ZJll7xmyOtXXK4rmr8LPrVVtOpJuOPdkfvLrmi3MUiKw72xArLUrW9vSO4L3DPtI
T+2RvtCcNu6sBCBY5FAso9qTpE3BYxIFwaSKYhOaZgPPwPW2mdbVNENo2Ti200Vxr8zDt24GUXzk
4qFZ+w9yUeAtek9VXvTL4JCxC48LuuIVzuL5Vg3Upri0WgzZF68KlaInEWAsaUVvdEvvHbMZr7IW
XF/5shfovqUqrbzcbeaqowistO7JAY0VSAnLCg5AjW73ZNjHnEsyCY8QTQBmzwPMQRfrrATRGWk7
luqUVHORy3J40B5HDQbJleWHqHWArbfqJXrAgNa/fcP6OgNLr9TeDM8hjGXJZjSdV0cck3PYaiP9
IKhOY1iIPTvib1rlgjXxCtD7k02XHeIHgESqQ1Zf75sHJSO2pRXvzxUrab2hEroqcgYjSFbiPA2Y
4XdDME04DkKSeujNEq0z6I+WQ79mctUUEXGkZ1XgRJQsecWSMolxm50/ayAPLJwtinlirc1pmYqW
+sLrsdfejTGCApR+hatrwtJShsnUOuyAvjX8tipGoqh8tq/ZHeGyqHW4+kJpAq7HT2KgpHQ81VXU
NX+JtKdJK211HkP/5/gC5x5HcgfPvi5HSbIWCXdJqxZCPrbrJvalqHnBc4m+35C8TKb4Loe8zHhi
PAbawg8qxSdfT+RqoWTC4R6SNnR/f9lyUGsPQxbI8JsYh6/EYUirl1YzKE6lHwVrspO4Xc/+WFb5
AjnaxhfEg/3lJyDu2DEIzGRrtx/60Mkd+F3BFSHWPCYlJhfZY2aeESmIqiNn8XSffcUi8VCSujwM
XKwuvAjZ3hWuKOucC9YM9rx5FtTlU9X6hBUEHwINyBnkdt9jg6FpRxtGP+D8Wj0FFOJfamsA8YO7
iupMLdN1UDr2huxVShVTu5uVKb0l9oHuyil++0jC93teCikZqpRSZI4o7CR/KQjo9uLAlG8DKQGq
PTbE6E36/ki2NNvwBfsUmdFwjs8Qj3bNLSqFwK0r4ByZfi+bj9CUgWYvQ6URH+4ejqBY3Lf1irvj
r1M1eNFSm6I+U9nyYPMmaoJksei8EDtyM2U0Ya1ScTG5AXEKPIhNb1lSSpTJqO/sTTIn7GaLFA+j
l43YRMcW9q7sJ7E49wOBA2LMjkRMIVouJsRuaRavRwQkrGktx4VXkjZ1UNpFGdbDcXg/HXvh7hSX
hDtvdtHRfqeeaz4PGEApBpbNutkOsTLY3xvLEY5KFxWVOwMhyTv92Gm017wn3ndIZ5Dtx2VQeyvG
Vs2CFy2oxgMVC2HSYVYeH0W5yOJS3iZLLfbzL+6t+Bkd9udSrDIxrLoFVn7oSfFbtcmaTLP88ZLL
Fj/waZdq/zt8B/vvWj9W8v2zscmjQS1qsaJk1l2CV1aVJ0h7JnFf70nxZZMIhW81jfniHnE4WzFK
RjmUFqAbToqUc3QkM0HQwcn61mxSKiExAb5PoS5RbZpF2rqQPz+sYhfceqn4EPE7HWT44JDH7e6r
8zwfNvPbfusLsJjuSLq2wSDr3B91iU48n1C6Qnj6R6qc7Lan9cutw3Diy7KJRM1sZkgxs/Q6aWvL
lniEP0DiXRNjTguAOKa+CiW+uF0v1c59SvdAhgJhH7EMiBG0IvwSFj4KkS2hu3/S+f/YZckwhi/T
Ut1a2XiupACl9W0ucghscwhBMkVUMdxAIn8mos/s16vAfKCFSc+IcamzCzq1Cp8U9ixtP+HKiZ/q
PA3cRABF0cNXkfBzPd+fEU/C9lIjkpyym8fZ9P4/hw8hmxw6+iNjr0tfhsDhX+lfhjFnRNpg7DwE
y6NBqpj/grLD2POqXFsXr3LeBNc1zqIloD9ZdbB8coZCLlosgwSP3dUBUxnWT+DYtDsWGuzykRua
EhPod2bSmX+85PP78fp7K9/sTq8jOwab9rkhhnbdM0jvfzj+XyICANvD/SU+htHujoQhRXuj47Wy
8BjoahejiyUrpSMOr4RjqfEXmPNiNteA6RJAJgEZS/udsQjV5sF5EQGfTkmyJKioljvdCDXWAegQ
8ySlyQEIk3qCL8Ugf56ybYN/nhwb1wsPTLLCGsURDQs4iZYgEHeIIvo1mx2Fu4P+74gzom7so+bU
+o/lFUclmaXPnKQ0bT3nU6rdDYzsE9R/v/PS/VPt0kzRqsm6IYLab8slCTET3YtYtxeMx2PUdNy2
fR7GqWvRjDpYHTJ/Yqb15jlvjQz/OG8TVu9Qeh9rM+q5uHYNg543R/eUNzsn98n4X1+21Eqo39IO
IKT0Iee1k5VcR5l6M0vGygj5/WrHs2gmO244peniBpv1yK6zcxFB4lhBXNJBEeB1tz/Y3tNqEt7/
gHBEnIfLm5M2juXIQtehUsT8HES9V88mS/P71CtVaPoTbt4vmDGf6Yd4VISr1HeEqnN4kjkwuqVk
T+fIdQqXNs1Zw5zCLIuWZNhaJeJPsYWqJxTo+MDGQHaEroiNVmvPqlCTg/GnnyTk0Qj5a/ltwZJq
boN63xBuianknZmR9Gd5H+D5xRn/UcYVo0DJ0mjx2QFmmYJLEk0AcqyMwDp/EkTvwElatoX7oM2j
OSlcCyJs41i5pXsq+8qsIfgz93+1qxfRS6gzOdYbVIE/A3CVfb8VAj1oS7iG1KC1d86L8+ASnD35
KzFfwyy7zHKKqqzQlA6PjzmmqMH92Tyxx/B7LLH4lHisETNnV1f94OldKr1027nJPX1e4AoztL7o
xyKpPQZSjryTvpc3ptFzAirT5eVr2gMyRQWpWDcx4fL6TI0SX8zVNWXEqzXHjfnpiueQlweAlIQb
3ac6QXqeAKVUMmW78ob+zggFz+EdcNTlkCzCv71DnCrgU5s/UqhZPIcx5hDE0Ttje8kt/5tdh6oR
+tYPz+uzMwxu7uTotdXQ+cOsgDK/8V5KEz12/xntjauLtbsbvOgBTB66n5bhgfD0oiPCkXQxbsJ0
cNzQIaaA1/N8wQdXjBbdpXipVjLRHBMlIfWaprBUvYxTU9k85YEZeGItp3XBbJFI+YNY0CpN5XlK
wxrjHUxCcID+vhHouCVGhxmjbivPhc6IbLgH10TM8fhgvR94+2vO7G8xoU6xi9DsEijge+vzBQdg
4lKfP8F2SEvSIerv3LPhoNYPNa1T62ZERGKnBVCKMLZC3AoRV9P9LZFqUd7CddoLXDM5drdhYPVD
7pecV1foCyHFllqRkmTyXcY2Iif9SdIBkJrx/GEP0nl2JFLPpScynOFXAukv3pFTu6UelX21P4GJ
G9pr2osy3vZXTFZYc8uipY2o+yW9eT2SNvmqsQX3FSgAl9fEY/Akc8ukTqqnjKgJG1gfE9uMAFbh
tAKCBNy1SUqqMwdufX3YmIXTvQkz/N7XB46i9C0BVeq7bwMzIv2m6jFDikhi9gtRt9X3BvIJO3EM
mPDkT46/KnEq411amXsn507Ktz8sIOv/Sgghi3nVmtz6tecHVtuhMPM3dI0OpysmtyLkH3L5LIDB
l/kXbO2ZZ7/vzMR5Bye7zFkonGEk2SSgsvQyAqHQfRhre8HJDjwJelhaqA0utxe+YHdhZHFUiKbk
K/zOpysCICrSLUEgH6OR4m1DtpUjiTCV26YJrCgp70kNW+rSN0idy0pl6L6dSvVrTHbRSEbBInS5
ACVQ3wHDOcs+S/Kh7Au8g9jlgqsfhHYuHOrxWoTYhCikurRHW4IGgHGLPSVwUboyN+L6gzPi/eci
GDtCozYcrKP++GZk6+5CYcyYYs1jDbFEvGvEEnlLenuK/+ifz4s1bBKilQmrguRMtkHH6GDYOGYj
0Cie6WUiJoAJ26To4GhZJqqvaV9/e6u/cAZdhsU3a4dhbJvw2mACbfHiWf2k5rI4bl4nrSW4dF6S
36bGy2SQKAM6Xk/I1qvrbJd8NR/luWqjeemNLXRZSrW0vkXxygvH1QOPfLf9ktBOIiXUAET16e4O
iWEajKGu2a++VnnMv93VHnnbxZ42Wq6equ/KDzdt0Ubn2IASy+wIRxXYeHrvoOBFehjEAt4aMTu0
6Uz1Pgf05T6vIt5DLLaGXIs+MIGLVdjX3AXVPCg77OLy+f5vhhhuqqqIOpUoHQxJfAY9VkzY5pBr
MQW0DNG/74v35Wu76GWuJ3FlWBtGEtSiTyqS74M19IbH/oEkbIhajEs7g0jnMOIRZn20ZtkZXbJf
GxRPfT3KTT4yc7+8elHamZJcKt72SSVd5yYV/R5TXzx6PDapAVr6FOlpn0Ooar5QN63FVxZ10W0U
zoGiEPljmnRbM7NvqS9QEmqU5uOV7Nb0yd8fTJfec22jCVEFe/+rXDTbqO3+GfpKKiOGQYiK2Nsi
6ut7UCSJ5+swmqJNY16xKChgei9IBulE3/u8h0T9+riCYw8CjFEXfZExi+DE2m0dd/y5jfJlLFS/
z9xtgFniPo0sURfeuPPptcFifxzoIcDhrIfwBvGmQ/pqbAtLsPKTxsPgCgSuQFvgdmBeUd208Ql6
AQ9feQSsIT1mz9TnJ46EaENTobSq5rB+L3Ra2vF8AEw53Ja+xb1vK4NSdNFuYIUFkm65073O2zgx
Hs4iQxI3NsjqLpaLFsqq4miY0Gaht+uTIySIWGQcFxF+B0+NYucGl3f89YuXErXT69Mo41VgS5NN
P0L27QPNi13xuebftJ/Ji7r1Ope8joLX/EASwVI1ym1c2mFZepK/sLNPnfRKJadgaMdQX+pC3vaS
2QSua84JPbstEMHGo/H+Gryp5T2CUY1Bt6lmKjcxg8BmIzR1Lt0Rqkk4LQq1XPPeByTDzAdq27lL
4vc/oB7q4ELom6BngQRAtE44FUTN3YRVPyyTed37AQbaWI2bHVP8R0yU2N3LCSFEQJLiOySvAJFR
vqr1DgLvKzfGMJyLd4ERp3TQaZeYO6N0EL7UJmF3Szlq+pQpgJetSvn4Jw+rpGrq3cyqMO2r4u/T
icWRUaKuv7Er6nhy5A6hvQcK95trN4AK6RvmDI7LrxlW300NuRH0+2uNtoefiWCTrnx0H1Pyru37
7cPuR1oIvG0Sx8vwjqDjpLaz17juDKr2uyLqiBrxOHKWnFC59vwAhPqARv1qdkBa9hf5E8Ngv9VI
GAEv/9T0FV1H1uDc7wuz9vWxSw1XQnLjnD/gtmGTvVzywFUJaFLmUF0gSG4j/KEjJoBsbw7sx/k9
U74w1QZTMc2f+rZhFviQfFzlvoL4c3wO3pFBQEok/lDcRXwr6Asy9cFy9w4ckLjFfY7CzGZ7soZG
Z8f8ypUG4NPjiOCGsz77VLFSKSU18vQTL/uRIxKPOKn3DwNTZ4D4WpEmbAKspLuvBZlMHKdHHrAN
oJgJila3OYZAtvdE/Lf5c+9hypyaxd2z8z6lBDs0VhffuWocapT2fHZRFEKdvMvbiG91hdhnhOD5
OKFWtUZayznpWo5qzsz6MQWsdoe+Re9NOPq+4eImCckVYKXd+ATNN4tT612W8VWGS67ItnfaBIYH
0DZMcE5IIZLV1UQ3n0rrD67OmN4t5Yx2HxBnjzC1XCy2PHncyxTUlqkBSu6xRQC3+uP06h0taKmh
fYK4TBNIHSKNLpbfaZhF9orf9LjRIEXVvcxrG00d2uOmbritAx+0ut+dZB0l4KU9h+fWAnyoPUs2
Ze6uZd7OcYvOmYHVKxtLTbXser5J6orzf3SHU9kP+snyZlKALYSxEsH3Z9hIIliocBxP7gLaRiwf
+lBkKyPMQanF9zebd58C8Q9e7ZO7uzJvMLWL3eNN+KcW2hBjlyhIhztptFZuibH6Ug5pG7advgjF
LK+C6tK1CHHV23x7abPunJlKFoDSfMIY9gTR6uElqMqjyMIBcWIlkNf5a4pcb54oBrTRrXXm/4lB
+stPzPhMuPyVPjihG3rrwy2247Eotwg66lk+Vd6LOyDie9SouQIG4auQE9F+1JsfSlKSECOdQ4vv
zTiHAO0ItFDmJrqJINmitoGZpY7tDBPYYYK8LN3Bhun/ssiwzyzpcjYJAKvN0PtyGmqa9MDihTGV
teRhR2aSwPRdYM2qbtO3LwxaHH2j2T5ZDgUSM1DFkm9Mw7VoqzkgdTCa2Nzuju4naijebUd10q8T
vgWzipymetnl6zPge/8WySze9DJj8CQxlMYUZ7xKISY6FuVmwP2JtxZuK+bIJ2huPMHZuwNG0VHn
93Nj9PcAdPa7rqqINCZdi82AgoMQJ90PSjll2zl8y1IS+RmdHsYvZkb2S2jr+eQcHXbdx1RRddBE
sxbr1TD19nvphLqk74GlxinGqF+Gk7IBGJNPOAJuRgoAOZfQuIinePbark6H7zjB46RvfDPgS6QC
WU4ybMyu2wZc69YhEXnGj12a7oglsZXxnN0fUkl13a9KGZA2SScr6ZJw09JLQ1Cw6zRymP9qS2Ao
DheoHenhneoGR9mOpHDneKc19/7aFb97TfO73WXCaRT5qghuSX5bu9MTL2QSj0rXz3h1IfwFcGLH
bl6wXLmCe4mdjmcoIrSGHY50vlCEWtVadaESHWKgs8Me9Ig6/Jc5Zww9PswY5EKPwSudBdKRCCaZ
n66BN0Y7gTpeZl6p11uOegCXq9WEYVNtVYoirc3el4+tDWcfpizhPuTYW2NHojC+v8PVvzD+iKg0
3NED21YPwp8A8RMy+BuhAJltCWaScQ5Sm6qBhQqrF9jAKxwPmpsMShxsX9BZHztXO7OezZjTb9w5
qco0rdzcsG15dm0eALNoEPiDvCmLihy8gZ5gDUeOqgcPmedRZYKx1rF0rzs6hYEUGFACa8ZlTcwc
b5Vc/x0tgczmIJmu4W92nuKLfnIyAfnhzCOrO/WPum1j+JqepyAhKn2CRSoFo8L/GG9/pvk9kX40
RIrna8S2Sp+b/4VJ+k6EgazyanlCqJm+jVC1CZMcT2vH/5qhGorWcuJc+rWlvdN+SOzJvXunYz8L
P9RIAbbE/EUtD8TMg2XWzhjvzqUiba5AJafQn+w5M2OH8NB0PlGnjcmyNcJ/KvxzpjdWsn/YpNj4
lZ4JT1+TR0mSZkfEW8x/TK3iH7XXb3CLnUjRtBFfCpRVzdc/EWpWCSsg52MtOrkwXmPCTKRNBt1Q
0r3lW55dqOoaHtDALttSLSGv86L2lhEhihR33yp1p7XAiB+uoJS1NgA7MhlJ60d7VcskssMaKYGr
WntEvegjPHaFAph+Phz7KdiMKar0bSU2j4R3k2xKeMuUnizF7HppuwTFUElqnhbEYthQ/AAYOOzk
ycR1nSRdraSBh+/I9rAX/2AnBg5JWW7XerFO/I4rKx6+0ASjO80pKlI9JNYIisTp7p0p1IJqRB5H
+bYGlqG9myfItO3+mTmqTw5+Jt7m4zscGUahCiHP4jfiw+PBm42dYBRiqGNNan0DVoNAXqbz97dN
tQQmTAD+an0on5pDcG/r6InROTGJXJikX4f0m6ISOg5ur1npPALkBb4lSZXP4QuZvvU44Tzg8dpw
UyqfexpKfsmzBdfdtwNHBfj/9/iGh0HAfluphoinD78LV0CqAwnhGhvfsX+5gsaVYjkPNFSqTKHf
D2JrqsahmbmQPR0PK2z4GWcCe5wGMLiGaniBFyGty/iHhR85K3Rb4oOL1ik+LhCt/tv2ZYSnDT+R
1xEQjAAsrdI+kl/Tajl13vxX007qiIhUbhoNzJzLSy+wunZyvndrxtQIOKbJPmj8UCFR7fS84C1B
YfFVpviPs+2yF10HkLBWOTHGYIrTA/6DJkOoooT2Z4+Zsh/+azf/aGGzAlEd3/vQd+V19dgQgdiF
eJy3VQxFSr+6gSqqHI6311lA/9Uj1GxasNzbeqMktClTKSP86NZHSIvuhtSaX106VJPZIM3KZLHp
FICimDJS3jcVw2+ukVRjYCqxzJjsl2W4wHELyHf/8GagNh9hB/eyzHtQnoO0ISoB7TgDv3lCmlTj
6fvCtSLFqbN56l54UXKbxWgb/gMJZSsBdT1eV1syw3wIt2yDUtayJpBqDq9N/whid0iVcrMLQIjF
eIA8rsORWW6pr/rXm5dCx4+79YnzG2ziqUFRyHO5ctdTvel7WbKGSCUQoCnYa9dfhslglXvprzVn
0v/OcAK+mmMyQP6qk4tsJAeUgw7fhSRFTZRsb4PXiJXiG2fsVYbVZf35txtsDoryJAJtfSrKMNEK
svoL+DkdvV+ZeNlEpd262dG9BBIh7Fg6MQor2MxnW5DZXZyBmzDXKlIbSC+yh+usxN4uwp8JhAwt
QeIGfYbpUTKq2U5sRQtMoZvjtnTX8gtn0Ix3EWEZahfQOdP7z3vNL9CUmBGGMTOxNjtaZM9RtAgQ
Q8u+eOjYgX3M9qQO1IzCoafeCLvLLwwCPXXw3l29qv/u1AMdr1NSqk/uHd0vci4NetmnCxOuRnX2
IKH6w5O7t6gmyd6bJ38R2o+UdpF+NTA4xstaXudBIcQ96IQI/amT+9XVrKNBhVJmWkxK4woJIcuL
unuSD9/J2m3jVsj5zs5HLJrLJz1TBPhfG35KQC0uNXsfY+Sw1hUKmZTWDWMDvw+K5InmwcpPDP8e
GFyApI+trI2PW8/wZQSAU8ZSdSUS28+v6qtEViEflAj8V5GK6YuRyjDHDGPNYSg7+14leCOnpapY
/Z3q2GKD4gDZA0u8OwItW+4QPEXQIs/9vQjaqRLZYQX+5RhRa5LCpZkhonAr4ZUKDI9KpXnfSOzR
/4MsZGRyS/IdIE38Fg4gjh7oK6rBNzC1fmuoiayLQ6ryXqh7D7Xe6C2++2Th/QuMswgtNxilyPt/
1PjosmlqSYqNo4xCj9cJuHDVdYVDZOxwIoiSNpiM0azvFETg0bl/MwXn8SpIaxgFn6AfGUp81cvW
AbFqagr1d1gUoqAGmNIP/IcElISQss18dQa1Ehd5JhpC5GmOna7LJJpXs28oQ7JUvALrZe47A0rd
VbZiYQH18U/9uy5Dyz/4Gccy9kzFYMjN4vDFKCwbSJ0/54MhmcvsBJviaP1juPg15SNzwK7xSvQ7
qkxliTxXjL1gAeEHhmoxcKPVGSC4CSUdxYCT1x2QLGU+CNOfkQQsWySylvc867IOg4shiABe6sla
I0KqQfxnh2V02uLLBS3ZTCjWcVEivlvXRcs01JWCx4VAXBVLS4f3ZM/SRVThbgsWk9lhYgDKOZfR
CHTGWakQZZfXbqOA3bSc7fsvB/vICHhLb47sow6YxMy4EdOYMsDlQ1WZAHUJsP1SFMjh1kn1x4zi
kKhK5gwGLLcF22vbDYjPJTPVK2xbzBOEiTnKdxmeNv2yx6Ell+D6cRYNnn66um7DSy75J8pJWoII
XHotU+tV4X4I3qQth2uRUv3vonb9epARjQ4qlKhReYAZxnB2YHplaS4/6zC2aCNpUYBkORhMma07
UiylCLpxJlYiCilHzTUSBWrKo0oU0ITw5W9DGbJeek9UUNhJOC5Tn2o+1t3w+/lNdz8Kf1zmRE/p
ruf8elwWBRRWaaH4D9OfScKshiEzyksKoeQy/G1ssF5vidOW0bE6Hm8JMoFszfH62HervZwn0Hbo
n6crfbXcHuPW+27OOSSh1Y6l9LXBXZ7NDmd5oEn1uZcFcr4V6pmwRFnrbK3n9MHdFPIpgwm/LkhF
fkY0EfutgjPVNFww65d9vI2vx86tnJJ2CCS7kpUPp2C2V4hjq351+ssUatXuqO87YLAZI0rxZ+n8
ypFFub6IvhNnav6yIfUcj9G1g9aUP2Nsnj3Ne0sPBFW1xFwYQmHJslXTl+MP+vZUExoI4Mgjqmmd
bR0ZxlwbLwyED/1cr8jLCUeZT5wgSr05GL+QjJvYlidqdFvWde6ejSU/kYx/58rtgj87lMv1Allv
q5258efHHh4typuuOI9LoY0eIByBZI7a4mSH+b1wzGcm9ebrvQS/kIr0YOBsM2n7PS0dBTunn/kN
2FDJMk7n9mr1vOpGt9kChrFI3Jlqy/PT3ppy7nOp0vD4RoVVe55Ok8QpWhknQCdRwWEzv60GYrYX
R2AuAQ7/m8ZyRzttlbAb2/gPPWXNahAKcY/PumcN/ckYBWwduNugImhjynlsy+ft7zNphDxmci2K
O4auuElDy5EWkyu8QlOCnoasfPMFCZUzRmxGf691SYVdKd9NICERauvQrpNfpsPBc271HNbUanC0
r/cXiIEsMxbl8/YjYbNqCPSJotTilN9v5iCeh+uOxEPwvXVkMqUnG8VrIxmcloqVBPXflb2y7Oc4
U+BBF+wyMHqDgu7mca1VDbLu8GTIXLs5W640AG25xmDzlJ1bRTugG14z1a15NB+kAbELaMH2UcnJ
TtVaTrBR5gF/rknrsu2p3xZIlx+k0+pr0IFAv6X8iH5BPG8V2luoFi+CBYuPdJEpi+MCSd9xDzpZ
jntTL7uF39OrbbuC5BRxoq+UXTUeGbzR3w2v/4IeIJPu7/CE5y7AT7/r7eCVTQdlwESiBOZC1shk
QYqBqOTgaZUy1LP7MoI4dmuKCm1gizFXzaCJFagbFw9iZyusAMrIroQ2/uV7M0DZhk9zBxAbAmZc
0YJwp94i2CD3LH+LegXGhwDcbvaiDjIFIM9cYZ2OAI739XEbNvQb7WAtAss7r+X3GO/3k0ogOCUz
fVnLAV8+h2WZsQQX0w3Yj27hxjUy9PZguG9FKnyTYEs4v4+PXtBdzwSES9fFuASuJ0VKfS6iTTks
bRgy0DCRYMSp/x9eFiDntAYW63ZO/PnQuvm08wIgp+UG44trtZ0IPC7u6A1hy6FXtTdiK/ytX5EB
Y5H8BVaISlZv9bmF8PqIOukEr5padwVdsYi/dRUbpZ5ZSjNdb47BtUfU6oTPph3ih/Mr/kRmTIjg
jcEAgosor1J2XHPs3krn6J3U263XHCQXSyXu6W4k6UQhrN4sbO93bAKdoLKpg5gZ3t8tRCVRW40O
zCnHGkx0r5S/f56WTZzyddF8fgz50DTJ3Bv/kzlj8QtWoTYBAXFpRtXSEBiN1MB6yoM4QXEKe0T4
JCnKv5iYZYpR0NfX0BcqV2ua43SHhdH+MDqbhorrK0SqX6il5jxg55ljdiyjXY4Z8Sih58gEha7d
z+ipfO7ZTsyz8G/MYjzAw+7EGjZYMAiLT07Y91UHGsdIVwmIxaZ/v4wtV0ms5GLjkGEVnN0vUiig
JhI6BC6u4sZ3D72muRVexA0PKRQUsnKopUTmG81qtxdwLJfF0mEcFAZzuTQAVYBJRR/EVPfXsRph
FUsSChhwGl5+xP9lvsjTI8+2RGN2rEKnHCT474lAr7E7YYSJr+KpayBwRgAoL9o2/WUK2a8T09Qp
nxVxtmkBj6+4lfRJFac6WjiZqQaOcQwYRnWfA9hGtR+ILFCfAKa/rhEYvwR4BD1HKKN55/dxTA17
eu0l2kPINJ9USPzVS0paq+SwfzsgH3zrxvGLmxVhfBFaWO+OIysR3EIGKhccBGkTJQt7k5czOIbX
C0oeqChT+9MtCVCqdW7PD/wwflT96m07V64bU7OLhQgoLqGRCfKttwoplpbzZGcP3nKkq23Vdq7T
iheTRYf7R5tdoRw/nkjO63iwsiHMpK+QPPnvKP37L1C28ynrrUouSfCALeTOKZZYieFyYui+e9Dd
2no447eC3jlOWAHe/49V8Qrnvw9U2bDdlBaVr5JpyUSLMID8WbCdN0APL/fZ7HcOYITyu39MG0Vi
y33syHD2fh+sTjUhbKA9HncS6/9V3+dCbZSMUFcsVUsaknXYBg8i1lgZmRsCRqrIGy4Ni05oW5P7
XHUwKn+QMmEOM5qKu0/9pFZfmuA4SoJ+DtmG1yKRqSZ0r8/G2J9DZBWRK+MbR12jq1TYRmpSt3ZH
w2p+sXaqtQ00KHQpLUN4ZAnZXEKCC23z7l6sUTur4CPnDUtlXr8TYKcgZ2J4z+Srf4/5eI2tNNzI
HxPpULm0iUgixTMGJn/wzEVSWLEyeZUFCvRd2d3dPAI88M9qUxCkVL5w5MxAO1edlu/CRhJviC8B
J7vTuqm4Bg23BAVKixnpPHQ+J83O6VCPrXCqmLud/zdfqJg7eVgwyE51rjRHuWqm9M0uRzh+Xsm6
JuHZ9RglW7SIxqmdT9Jkz7ipFOQtSgtYw9wimzZ28taPe+qyd8di3UqiUU+KyUOnw6MzuLtB3/ND
7iIdaGXGg/FoThUjsTdw6ojWclzFhMBQTKLfelvbfcnnRZx50TS5to6GzBzxV9Nfrba6ttPkTxYp
xVK+W6norsctsWyj3ATiCT4uhAW6xv/ZxX73gWyisBeLON+yLBcZbAw2Yor87QGjUsS1+e6/ZqUC
TRduHtlrKY2DmTW4pn8e/d/05Pnm0BKs4yurzerH6bDWOgXFfZ5PWd8/BYU2v+FcUP+w+9IyGXeq
W7bdvTxV9OBcFO7UicCpge0reY35bYbILtkJPMWgnfPM3JbvE+x1TFdKESm6NLVz9GJSiF4bENA7
0HLCV21uNnmWVA6hVQqlMPBJErFZ8d3dMzVpBJeJeXo8zMAkXuU5e5I2Xbqr1RD1yFSD83y/kbnB
kIJmkqFqThjJMAgAHkXHP17GL1frdSZy/NkClHb3tFB9S4rTEqdMtDEtAoA0KG2OSaEu38Yb0Zn1
FWgQ22yExtjvmoVB8QAUbkaAKutqLiAJ+dtPSQb7cvvNXKHN+5r6ShH3NfAT7qmG/N1N1Z9C3dMe
i6lrAEakru9kvxm2QFRVT+2vquaf7wiGFrLHz7HRE/V/I19UolZ8MB5tdW0EcvZ+CRxkQUYDHI2F
HBOhIbcJVDu+aE2NPkSMiDSs/b2rVt6sF4hjmnZGg56n9dqM1sc4WC5jbxq+ljWLA9NMde281w3J
7lZQrosTkKkSmS5guaO4Iuv9Elcmf7hBZZg2hDoUD56NGShOfNNa0iLCP89/ZlQqd0UEp9YOuE6B
GTqjiEfFBRaRY+EXHuoqDOQWM/tn/sFS+Isk4dcQbKqGJFEugr57HmKdLmDT6h9XyExNPrVPNILu
B85fRoHmOtIi/jhRVYThg3WNyD3Ia0w+8arrsE83p02SOFAGLLBn4imLL43fT1vp88UgiAjwAbXi
a28a/kj5wgwQtG7mLCcljfLJ/W9I8Qb/oyn4yPThK6pz2G07iTBZ5BCzuLmxn6E4+lSiyhTDhlDu
P4+dq6NPYmsVpG18ook4RohUsoxRKd/dQPsegAPX3IghqHMLxeOrV/Y3IxkZR8movb90SD67XCQI
/MqbCiRDZFayZJNiQcBoV9Sm+92k50OjpFnaLbgQ9/9sWSe3ziQ6DunwGEA3aAVo1sipyAxlrT37
3U0CI1NJ1G9k62Q7a4HxBuBBWRunzwVuoOKJLidIiRdFlGtUm8EORrwxuMfpCUwWx3fGW7jB+xuZ
UbrDWcwIj9AZmD3x28TXAxvltEIeWdt4PAr+B3x92XATbMu5GV/ge7e+7qo8SPXiLKa0dkgwyUcY
8RKO3+uduVhzBj0cgtGKCYFv5Com+b1mfFD0OL+9A+dDPQB51cf8wedgs9bpkDwthYNGiftXrgzQ
Zd7CwaopMzUwjbnWcLMzw7rF9RWQwxty130W596x0KKEJDhWkQulJnemrmHrN+BILrEaQKSdHC+i
JtTQeH+GtYj/Srub28aPL+im/PUoGL/uphlKQu62rqdSVRSZZpz/FbkZ3rjNy476l9w+BDDdfkr/
7dD0xEuInPMeDfhunxMxnba6okHhbJEcAmLVfueOaj53kVYv/8Hla4im3PhIQ2VCw9+HiZ50U39n
l+SfGpcpSefVKS/JMFnSMCq08kTaokZDBBC5KV6esAeoyGjFZdOE6VsaKxkd58bcdKlWB3+zUh9n
pEzyxuAKzyQcbeFL/2hoRwNMsKF9HJkJArseRplljE7hdjhzQpxsDgJdBfaVWttnyubkU+CCKUdL
6nXOODyqGDbohM1iw4o7q4TTzTYDFFVA10M1mu1fAkOIYZzRyjqUprz1rZXky6HfvX2lXJLiSb1b
8WM9YKeBYbNyceomAdRIUYTxdLDb0pqa/zyheqY6kESiLHv6oWWMEN9+btNzo0KxgZ5ww+dHiMdY
yp8eEwPdVbgSzavoWysjvx7a1c35ZN6WarwRQgt8xFaKWzziR22rbaoZapiDEX6rxWAaAcTGrHYS
UcBcajwsV7hUJr0NMn3UbB5Q1l8dYEHXJWWZqjmJ8TLPFxAzz/6MLgOpivPQNA6jP5D9r2l65nGc
NQPK4oi/Vs8YnGy35JSogcRCjH6FCDwJz8BVGVtS/6IRgBI6+/ELSXPk6CPadtWeV0RqyCyuYrNW
v/oV4adiJQZ/aogYh+2h4grt4Em72jYwOltzC54cF6P1iFUGxyo9mt+z7kmA1wKUng8Q0KBL83fU
IJgbkGYPNjganr6Kkx+byOpJPVNK0aMICVvQPQIWTmPUcoepIWoxlcRs0S6zKpGV5JXnRmFPp6TM
D+zHHWM8phYhN5GFd9daHMwB2KgbB7u+R/5GcyW3/yHgs253JfvMjndAMo2R30rCQPnzKg/iNRXX
8yfJYGADE3o6IOC7dieG2ni8O2uGR+MxDUCdx7xFophpEgm7NvUXVELolfKxjrtdi/6yBt8N2cJY
d73t3nBGekTXYMJsDOehnJvlOI9u9ZwZGgU+zel3Vo5auOi8z0vbkjtFYaUdG7iBhu/GKIisLHBa
xD9+VNSoQFEMJIUI49cNXbs3DEo6XQl6GrOCYiDOzbhmtS8tcZM4q8hfzjaOAGn2ncNV/8Lun4/C
GpntA/JYOdyf/Kq2ISipZcsS1zb2yX/GoCf/W/xrqvVU+MCtxFFBxqiahpbTNeIqQJn+DdJQyvgw
w21RHd7FTEfXjZ+pJyk+AKGkkxCPOA9iFQYJru0hQiY0/IL0inou4jsO0uaEyWBLp+BAot7rQZz0
vBZ3pKpu8Xhek9rn5xYq4BTRGAgiiYlbrGaaUY4nza6u5BhOCklZfJAfmKJCJnjzUuA6qLVSxFSY
293oFiUPCXzsDFbpYZ8RDPnGEUdYRCi5KdBvXvmJWlsU9dCIo/EAh5iNN1XvKJISS+UwfXmz3KRX
JhJ6u8HyuUGhfd7+VrffRUi9sqWQrVLNUKsXq7/krRLReNhUUAKbowBBJYHdHOuVgrEtznECGs5I
nL7Wce+WMKp1MogSd3gNuWsFRSHgwM7V9Skj0kciGWXLPpDLzZ5a2A2d9a1T7T+vM5Nu46sDfUJo
mMb3KDpZuIO5zr3xLD+HKpiJMDeDuzyNIfWbhPXp7/iCwNn4Qf/g0+SRq/8d4vMpTZBMeZAsUwk7
y0Eiu+f8N+fEOym4NIoDDf94A28uJAvyTKUwVvmqSBFCXgPq/ek0uK3tjC1Aw504I8C0YLtM22DF
PAlWaQlkSvzqn2z6CvTWgwcfjzOYfo9bT+l2zW+kMHuE2rEnekMd+p4l4SRwUInhNmhZqOJV+ydA
hAS+NFQPE19h3K1PulCxaU5II3a/vmtkav58POyUZmVRPFnaVwBLODQqM5HS7dkjMXq3kldYUKbD
4i0QwsM2n9Jlh6VD4B/DBcjloLRryqRnXqQJRfWWyWgZ05ZLVGMcpl1oGnbIMsb2f2uc0nhCbpV7
zkAwCPiwXCRXg4wasZ/viC2Mv+90b2UnH+D5z1xEKaa+DFrSzxlF4BSd+8KIZD33MLfApDwXTl06
4zRrqbN+VUnNspXW45bAfzH7vbtF3kF2DAq4F9VYYpnzxA7rsuAKNENh1qAsVjLGgmCZopmW+dzl
D1vEbQ/Pg6r65n2iHNRk8/it/ZZNjF81umRqdbEcxsvdDX47bSUHiuZ6jsp5ePbm6ESKRqImW/8O
Xt7POPyvS2EWfThqtxJ0m5wRilaNOurrojC1o8ONi66uyStML3oqf7LUOk/7vV6cIGNzAIEO8VIe
P9brI1Vccy1WoITpkh54YgIpT+riIbafJ/DAHbQ1sfdZzHTwMU+sJKUul3D+fEgNwP574ZQpTP8l
TRJ5kZ955eEDenYoAkLWCKOAbPLY/6V8M8qd18OOG4tLea5YcqhU4bdDlbxWXhgvBkDUA5sak96m
9smmFFQE6z5DPlb+fz5Ib7pubnsRscoMPBTJRgP+krOEmijsKjoSbGgNj1xw/vztbqn83hhI57Ba
4vbVtLxQpPdip7f8vLbFnG5/m4LAcXNZ42HWlMFn4AE93mAOFwLNCp2i7WuZl7/A3MUM86wcL2Q6
KsvXvx9DbVRrfDuovmiBKtJ33Fw+pu6d05NQakNPhMP/qGe6u0ZuHwSdkQQmikK3r1r8Of1kxsAw
7rMxqcoEfkA0f9sC685cCZ5+Yfmsr+jSRIvRgLMSi0lzNf3SVf1pATzQbM/GcVQAyt+93nKwLZcO
kTDOgCVP7onqhC8pFGE5oql6bZW4+9zvzvD962Qm6ZeGABpSz40n69AJ61Ts5j07G39b3gfQ5n7D
RWs1XwmgevLL7h7d2zbouMrw07dx+8VxkpFKq2gw9cTnm+OAB7+ZF/brNhsRrtsUBBaEV/sYttPK
AnvdFMkstaroXz/viFzgkOFCriynVJ4cGWkkSxeKqe94SdrVMDUAYuSEVy5eZuBJz0ewuk9aVtUa
2OoR6IrswKgyqcB34JPGiEII5IPoVBgk3wBqa/k6Y14jYd7Mb0+raE8zBMsd3ltrZv2a1ODcybQ7
BjlkppSXhE1pPdWtVSOBO9g5Qba0wfvv5E0gr++LqEBlKpZPErJ3XW/rIC7BVdV5HcNvTbY5J9Tt
HNuC7h65ZR9UFS9knzBrfMXf6aVDZzvb7o9qxj7EUtCDjKBYd6XZFMAqPJbSwhi82VKwrIge2xPV
0xpNnYZs6IfyaJ6W9CjLtt7m+CIHpIeQlr/rDLxZtWcyLKJaq4AtWM9PUBGRz3JBnce52U6yXXi9
Fv1nEVKoOhiDc8DDqE8Ctrx8R8Cdqc/+tnL5V+mJbVcTNgp7diPQXNXGgRgGBJqnEz9mZpBHcWQ6
4cwbONRsuD24dH6d9eWakAFmmclTToDU5HQoG3NMjNWeT2h5JRizs0IAevdzRddFuFABEVQ0+SM4
I1vbHr2vs8l/PQ583blkRY78AZKL/CoqwLQ6Pmq0AsU189ztwre/ZLaSOLyuU731XGLRJQnu0Z1o
C8YDc786jwgcdmA+K4VUZk28Xh4Dsn4UsVgkd30OcHzyD8hN30mZZeRDKpo6viLNY34/w4r7l9T2
MtiIHoH6mxtm0nnviL7TrlaYPPR0MamA7G2VSStl1Z1BH3Xl5n4ecl38U0YxSzg/jjULDy/x0nDz
hsjUoh74AGihfb6iZF3vwZ1GQtWGnK+5VVcmDAApdy+GEkKYCKJyAEqrI/Jgn0jdIQoohPeTd/qE
ZREvsAuHiUS26W2qv574myH2RSSiBThl9quimmMhiCUoCdQgUiACOMUoHm34zcBUuaTxpo9qz4Dt
PvxA/u+3wd2hea/RCuJxGlJJyF3VVY77r2mgB/cIz0NGtTkOjCRdDJshFz5qg4HWLB1AgkI68Ju7
Dj3DzJogo7jknuNOBxb03BwAjxi1ExId3922bOnrqa374N6908nTDHagZz55jJGZB3npE/stDfRg
GsLkCkRM88jMVh6x2EbC2dNJm0LVwyNIOnC5jiiGpdHm9Cg62tmOW0Y4rQ7p9K27uEHFU5UcKAJQ
nbmHHkbsWfdpRbIwKiBuSy8HCv7+mvAoaRvacORqaCrfm3XvB0S6du8G7ppG2UWqDORXpDWMJIVc
bTjTnAZCaYMtIwl4BPN7uIV33IFeJpnLpk5ZN3kiBIX4NE7w020HSv++uJaV6D/l2yKtYLHhag1q
aoYnls9lPF33Htq+JwkIX9arEGARYQbNE4fHR5cnqEXhZ4voxWlBS1T5cz3Yrff5SOSCsyBnG5k7
tmsatnR+ha2fwRyt8JPwpd7WoM0j8lZ9LKxVfQVvdqzxjzUIeMieE0bn1ocW+A7bJrGDbuTsIQta
QcrK/ichBy+CygOpl7e66RmScZsgCk+WtG0m5Y5SgXLmCj5yzDepBmy7ALpxza9aDSqIEbbyfa9r
uV+PKtC7a305FUAiQHYn6H9CjaXhkubU6mHQC/wYAwCdfNCmKPSysh9HjNIWi2/eTlKGFtDVXiaq
EwLmKEfBtSIReKnM1Qxm6WeDB8PS4zN2VFALow6s2vyRWnRoHtFD8FxXHRAHMbDVDRVdCiWoNQJn
sFtzAdnyfALhFeHK5GY7u6er93oNReLGLWZ83c8G5ez8/WZaI2JtZgo/TXfiKPZfezjcflvW9om9
Wud4obP9YoEBpv1ZthQ6KNsUCSiS8PdYK0PWu+U65NthhRgX3aAGBJ6IztK5eexsMdNHTuD/fIil
MsilaE7zwNbB80t/PXVUeUc+wNwiiuxbY9CrcLPQ1rO+HOMpIyhczsRlok7PxMqZh6O5xzW33MQF
O60Px26E5zkdSOSty5CI1PO+wL/AgJ8Fi76FSWqBNdPk5PmSLqlzJlOZezdZQJNZLF8BbXLUV8SX
UoVygIFvKWExFFdFiwMPZm/M+tpjUA+k+phJD57ki7BB1mCnSxawNHSdjN2+DQa4yMN5CUhl5NAr
yy+YQiRrplbRfTSKWUn6pUMf63bxFj2P9SuruKZhdb6Do+kuAt4GPGDpjpyJDwagt6aI7G7L+MCM
0M7/ZuDwHfBvLliy2ysAz4a4VKGH24RhiZs+kRIS8SUSWBo4Y6j/rQLIqDag96SGYU4dDxIiehtC
iS9cigXx4e18YotESq/CphwAGU8Fu/1TPc98Y0Tg7vjQAA1aLXxEVLMAdTy3uPw4NWZB8EAjcwQZ
BoB10yytMbW4tVBYD9T+JeDd7KlvoM1QU2dPd0UWiDBuo+OjUksyXXEh5fqMbg2F/ydkkZv4q7WE
+6BVbZBW2c9e3WMDo3l16xwjTPJabL5oN+BbW24fx+fCwfdHynFhbj1osD5tWzWf4nqQAhiwNWZ3
+l5DDkr2RqkTcYjfwn9pd2qVdhggrFW5eTPEPgY/wfd4+5iXDSldZ+dtpzZb2QrirRd75+7/z9gw
oRGrwk2y33P7KPjNx62Y2oLHUMitBY5NdpRkgQGkg/0eDrMhRQ4aozheLNiWahPbZ8xwwCGe9Lbs
q1x7w8/a+XFZnDWrmUX59HcXmcYXuvoX7GwMA9kr2YCM2X9yZpG1UOf4Uj5m+N6UGMDrRJEVJSHs
rjkFyw8N2XKZmK3meeg47cqTR66x/IvFSHOzy5WEO9d4id1GxUv+/ysx7d+sNDf4vT20Z9PXStUT
HcLFoZ0SMJopsVySUXyIRgw8WkxPukQS2Q24B4Xt524VvZGx4+aG7+czR9hbnGhoeACNYNF70dlU
oTlirsRDMpu+ULi7IdeXCvVkfoeBPgrdFwHKMkC311U3lezT4sHepGHrSqKVKoVlFRyfLhTZmOrs
OXttVM6RoHCXuzyvJV+CaRMUJpo5Yar6BQQ3Wx5sg4LQxT693nD7wjl8OiA1wZYjsFTqwlA7jTF4
4fmvH0EZTZdaB3pFGFAE+Hv/YhKa0hetmHAfQAQufcP4BT0qSlTy1T0Vxu8/mzj2qb/7g+I2Jejr
LrbmovUlARfOD0sxRN259F/LhLySUZTbc4ZOh4B3KUfSb7jIGkHpto2Bk+G+HROsUzRWdCv19Yo1
B1xu5B53avGvgzgYycEHQbZcM0BduXNc3oYzVlmaFhj73nFx9OXpOANWfkRjLm/t2LHBgpZ00We1
mg0PNXmiAqDz+KtV2en/klPqenM13WhbOR4Y4CbyIuRycMnZjcC1DYYg0t2t3SgpkYOkQQ0H+yZF
uE9FOxMnYiIm2Rlb+0dHMgj4pXoQLue+I/OMhZphTeX3RQNfrEKDDkPAAa71lCmlKExd+y5k5AQT
Z6mX8Kd4k4zTlF/X9NtC8CmGF1YAIR8aNDNkMJ3+acAqGeTwEa3Gnl3UWSBkMia6zhACw/DFry3C
58T7fqhY268XT7ZeNdznn8bITIKYVquDl4LEFhUJ0YIgQwo/vpJDrirJE1RW4MZt1I0O6k61xVv/
OY08x/UzcQoZCUzJosacXllJJ48K4lLMdhDtPNZQrx3s2sA9bcODUVSNlwIUdpIG/JHxQR+7dVJC
iELODpgB2l++uulp1i4MpnN6Bj6acgg1ViQibfEP5gsCRcuV8qSmW2so2EMP3AGyXm0L06rkATxo
BwX6kwExR3ZVuxAqQ+rIuOkdvaRZJTVfzdUL40dG0iZLcSIZ5NEslYiHnkg2fZA1HarVW0BQb9AF
uHrhcxkhTPIBIHgIXdEYgDfaecqnWsYnn8IVhKlG8HwiPaDR4QIO02QA5GZaZ/cDvqLjQceRDda+
6waec8fGtbGVMB4Sezka2o016KYaS8bc/WgfM5hf2DOjrRoZd831eMWUuNYiG6azKRgvuvoZGMcu
QSj7oj2DFUks9MPGoATI7yDMBxfU22yUyU4Bl0/K7yEoFkOFk8/hZc5aLD9uPpKMef5P4QbWn7Q6
Z7vhnL4GZKHViIyTdgZzmFf2zv9n+wZs6XGd17WXQGaMFU7dkaG5vGyQjvmvG7PZSifuR+cPVaLz
HvXdjEIzrQseRQ2NyPju0diIcFQ+iUbPCbDNgkqK6Hi15PJGJq1CPZy296gWStqmgFCrTnD/6ZEm
Cycn8AaZoQFr7o8IQWdhCc2/CC28x+G+Fu0/CCTAvUAqfC5ZzrIrMEo1zVRq2+gIgiDQYLM2PLUX
f7lML+ZQeEUbZXtx1pzmBAp170LAj1P7eZD0lbHvbfDFpDxeTNtCGous8GjL2kfPfmJ24N7Z3SsC
frf6uq7xUgoMgG4/+UC1miN7SMKkvhQLySJJ8hi4fghRYu3N8lttABCMNUEFSeNnyKFT36pqK3eN
VNkC0p1hC0bI4+Bxtpx0Kh3ILw6XKnUyo6MZ7IdVCuP1KH6ZpTMbn8i9c56oI8OL294h5+El6qn0
Z0VB/tuSp04EuWkWvX7F9z6IusnKvtmLNzFMP3H8uERbV4Z+BhbpxAmiO4JJI4MKy87neh4Pzedo
T2QOSbdMY68r89FxM/npa+JTimV9q8/jpHayVJmbrcEPwuSnsVg3Qh+2yYhB6TWuJuRVUyLc8EHM
g+3ao+NUu7GXg69bHvZCiIaEMeHZfr/yP0wNBJ7cksyEKF9tl0MfG66q+5ibJ1Y5N6bjuBdhFibr
H8OEx5VZ1VFV1CcbHbKDLXQEfNN0N/q79phAfyJryuDP2qs1sBHH7TkpsenvP8s4obhHa4Gsu8ci
1EkjMy624hxF+nzgZ5sqGbnisJQdjMofekRnY86Wq2jkm0QYYYVketyr4idfPlan5IabuMi3k8JT
nnGTS8M+C6oe2D7x+iWJjDPVu8ziNIGaIhM+SU8G9+SayZKyjdB5wTPWwYbQFEqTm6K+BPFDuI13
spRdYlDZfgcHZBjYdp8dkh5RKASwmcEs32nB9qNik3vAywECiVJpWPpj/JbZBAmQy4FfCq3F6ts9
ynjtQeuJu8EP6QG7jh9SIvLrDNTaWPo9ZwlqKcU1Oys/qKa4OowOaZIVSIWdYmpeKhYfY2Ku/alL
ZH+jrNsfPrPPzUdSJZ48kvoYM8mCj1gHBl5TI8WKjA2OdQRqQ6+mMup6DfE2msL1N+QVjA46R/9c
bVnSaQbWX1pcKu7W1K+s0qpgq8xYtDwRZ627I0uLBrI4y8xCWAkTrDk+IHgS5hYA8BMxuzzvIVIH
/RYTR4g0Vu0oDzuh9sOQc5m+Elmji/isrzqaidXa9Jyw74GibeNLEesvs9daJ3mKil+D5zu0gUCa
PtSVSaSsAYW/U1tWZzk8nsiF/Kk6ItbP6ZkENqNZtRkMmdHouPC8RElrxaqDcbriUAF6DHRh7crC
ZDe/wYq7rFiYE8NmmdDaXBIW2O69h7JgvARHZ+j3MDoPLJ9SkMA0t9MeoDCHGgfK//GMobju6xoa
7I7K14R0UcWY5KNTYHYgHYdAo8BLyC1Ln/XVrpg9ZnbE9TX4ihAGYjz6BaUHYwCHgJVJZ7S8VfZU
IHA7pD+/rGt+kR+hTyaooLiFQ0dFvChtVUcwRDE6TFZTqFS4hz9mg9/Pagn1FnVaAfVyp6qHEMYh
y+34y/fa5qjOtOed+z+oYya9HGPErzOjzmuVxQjtz0x93FPGq5gx5TyRkAJ30jrcPl91PL0L3QND
6sJYhyVXrdQ5VhmnNRcDsL5dGi11Db3bgzShc6CSGWHUO0CagZ3DZRreTpXPJi7UdTG4ZNFTMjfP
ERJPWhdRgQZtTS637WsmuSra7vbeBjRwRYXerGivmRoLtR67g70H+wlHySdSfcvOb0OzFxy+HcFb
y9SpkOXlRkGFOuKodDGrBRqhcvtbG+G/O8wX+g6FUv+aT1xdC1F0YC5IHNOHMhDty2aUO9kdpY62
Rm4FXETPDYPuoeR852+5bcGUvF3KrFqgGN21XqqABBFMMtHPYafZVS7ySRi4pcB5oJ4OczwaVNKU
uw+nnS9Wq+2i3ztcNpCFsdGAPqbjS2Mj4jj8KCRWO3IDDCcpe1+/E9G5q3eHHMTcCOGqEOtrI1Ki
tPAs1KKS4nEZm9FoAvJKdNsmt8R8r7vZzCVNGPttxpH8uUBNvnKzh28XFynPfuoXJ8Gls//2pf9U
wsccB48qU3WROFjWMchTlXmW8MZWrkD6SxfiQaCgEj24fXs8V+H/fGJiCQv2fxqEjJsE3KPCs2G/
hoCVHhcSSsgk+zVWzNbw5IFWk2FAzqtNNw4Z+WAjaXEcNQICEiEOsIfEe5k+4+CLGUjl/JXxW1CX
Ep9UCGB6T4CwV5aoro9WhhvQpz2fMbPcEXd3zql6eE1/CvzgVnWoWVjnTT3MkE8dMd3tCl+FwnSs
ifO2sIzPraPnIP2HdSSTQnHsHLvnjaGobUsHgS2QJ+210Xo2EDgP2YR9Jf4ZPgCsmZJOwSkHUfh0
AEVm16r27fczczb0Rj9s/NdvkIGfrF2g6QDe+6hdEkw3Y2NNZ53D20cpOJvUgZ3z2YOjm+s54H2H
LZ7xsh9EnvLunA2KCUC2dUCDF/2hNU9dOwbURiMMnaCYHJnPE/aWs9NyMGBw2x5E2oM0tVkUZHlY
PZnLs0csRzGIv+o8lCd4w/KIrfEkIZ777sVHozKTIUYoPSVehZgGA5HfTPKWpD2VnEvvkITBhLct
38TYUToK5VwjhauCIN1q7zMsuDKryZN03lLi2wJ5pK9w3yMMbt6+Ayh2UVv8Kn0Mx9/4FpqRVZcB
pTaD4eZtQzpqHHeq931+ohomWFf9nBaMqwAKF/KtbrcQow+s+MQokHy2LZXEidaykjOsL+w36uCE
oHoFTi5It7PpH5/XSE/rEQxA/Ic659OInoz0tdq5QlIFWdWWPg7kD617qcdyOot+ODzyMsY2SLwr
h879EqSVAGobyXxSuCH1hDXPw+f4MgPc84MMLwtrIkiQIpEvpmVtndungM+hEoSkY3P8YlE07GtH
iSLfywXqIj89iHVT45DWdXTTRebXWkDjzQ59n+yOO3O1YPph3vCaYZafDAY+R9PCOw7mlNYRb0nW
76wUcMFXal0UfdJJ414bruPLa4KQqKCuRf6SkXITpM8Kr6gdugurzmk6p/qn9AC+UyLGivI+X8T6
Tv9oQfHVOgl7cUGtd/8y30CI6uGC5PrWJx/TjulBeYgUwTmG8Fri2iXuR6copRWi00w4MrD9DpCc
cel8wIWSMnq5WssEFuOjECSz+EycVBkorptTfQgSjLZLbn+OIb4N/AyGVu626f82VDakRpGlT/Dw
fsSMLUsQnTTJrl8QSft/meEJvIlrTJY4bqjwSRoaSxWYArkPcAPB9+YbldHBp2fmBCbmcdgCqdDC
Qw4GYkp+3xuBGCtIvqg1TDsmkNak8uU94KFoQymzLbuK/1GamH+NJ92YM7c6k1G51+92dDWMAjay
9XU3TXci5U3weZ/+1tzilSgPyD97/R5NOK7sHsO/miFD1SM316UM8RoCh2HXcIZ1dpodanAebtaJ
iX6vwcRuJhuYBz/6YfRRTv+lx1YD5j8Z3U9YWOzbAcOwV0JEZW7Ce5o4mdLotpWNn3EKQRSH5kby
JKcrq2zRV/cRgXl8//tLYCFeAReGkdIb01BJw4WmAzI2lxMBVHAywt3YBrYR5InvhU7gGzqilK+f
udGmZcZ4Oy+tjAGqMOqsq9BU55qtue4+ePdcn6snwSrwFNLVr6b7TVz5C+A7W6NBOvC2BLKBfiR/
w9ipYKTtD/zmWiOaz60YRD9byku4MMAR18cu64bubrWQasOzNQWcIYsgmmO4REmUl8SS7uZNSj25
QNw4N7lRpVMW4/p44UFxfvsET4CJxVVLDzv0wBUZY18zisNvvg0CPbZgGcZ3mhd1tJcruC8ciWpf
N84bsL2/2C9pfNJM7fVLVAKo0aViqorOsMEkV+OOdPhE3jtVYePftNVQKaVhhCl2js0/hSfuXW0c
/LI3u3UVVyu5c/ueH7+F+RxqOod/BmcMb6dqvn4WHSVds4x4s3lMr9uP3HfS2pozePE2/t0Q16qt
0Um3FaxZP11DOQFOIK43SQsTdVbQvUtSAh0T1JaHzgTCTK46iwuRaBwbLrX5N4hSuSFAegdNO8QN
otC0riH8Tu9mE1uLDO9FiOdQUNBUwOaqlueaAfOhdqIavkIX+7W7ya9rmwjaeM1rznld9hAXlBeE
lk8iB7KzhD8DZRbQ0XuYMSdbzreR6pPBPv34hpzHoZCCPtKb9n7obGaDKUk9MW1iIOIGSCVhWX3g
xqGI9Ks8i1mw0VTmZWnwEmADBt+A+PnLFyBA7NHWyBBydYpovU7qM03wGzMtINxpRcijuNQIuAph
iEXPofbHyYbjNBzt+JoELRGogsXJp9UdaVvIGM1MxbQCs8duAaAH58VPWsYh1re/WmUb1bqxPW3x
uZHJmy+7S2Q6iOKxQPHpr3yhW7wfJwKTmLOAeqkQoB3+pr0l7OUDZzmh2dMp0Mg4503kdGtLPP6n
0uhx6AtJwh7eivmoPm+J58o2w5J7w52k0Hq5cqPmE7AGTpKDCaoEbJ7kjbUJFEeZkCg2AhsnJZrn
qPbiJ3q2QzTNMnetkxMsP7etJNEqAeJydaYp4JBTIBrQmVJvnQve2L2W97/Ca9ANUw7DZWGQ9PUy
MveZz8p2Jj2lbxwGxwt3hEnyFKb+7WDwodjnmcnEVCP2RDpbgVGQnTa974yAhgrcmSc9nOPq8Ipd
srB58jnonzyo5YCeiqHeJNtUIwXIeDr+dR1OCGsL+wgREE5H0uyeE6YdkeEf0SYxAqFvaTkd/bag
xUdMUixNhwEiFWMglWKHV74CNTXLQ/Jg0zBsMoSVVKQsqKmbChqWX8aaVmn59uZIJBDdXXHgUn90
XTceJttT5SQiDotWfWCZ5lhV7w3DzxfjFPTxCzXVvKmIcfLO8iDzHDkuFN4AJFSNkFf4uhfAS8Sj
h/BP6plsJEVuS7aYkqUzNflZT4oM1yZU7ZXWZ+vzOX93x3FiJL7M2pKmSQlBwcw9OpoQjmEi/nC0
MUOxuwVY6JKTcquByo2y2c8f5h+Xad2a/1IvS9a2xdzCBj1OIINyZ8ahGf60qjJQpR7W4KZzecYT
38NtlQKnr3w9fdlqfMJLhYdrS2k2vBD74iKz7ThjJqGYzl1kDvH/cU9L9PRgVAEC390mzrS1Rkgt
xIh8XZrCJGjrUg/zUIbc/kh/s4qmf8z94LBd5DAara6nK+ymYq+qfvhTfv9ASqjdA4pNxj+SdNOy
mwDtbv1ScVcMP8VF8iW023iZOLJcaOHLSTAjcsEDtnslIgp1LkoxgITrG5L7o3iCfq7B/1cLAyL7
pYciAQh9mChcV20zgKyMUYVbafzBoL5ZB/1xRQdP2f1exTtVftDTmA1RVHeDkG0efFzvbsEY5Ezj
JA+rpMxjdE9S89FXfS1UucVWJLT4kBcwDN/mAIFZ8grY4XNg7TeGw1JmRRdMAA3xUpwDjoGic2f6
QhwfRnS1kNu3tsBjUrCML06J9uIjkwi8/NAOyNp2j3RBHQYQUp7D88j6CUD1fxysNHCJrXU40G5G
EKYMZzHMbNTpFrmkECNBt7i0NJdK/ajEC8zxUCmj6k9NnPAcKl6xw49b9h/EfO0skMVfPqCU6stD
lhGL2io6MEbSsRD/w/DPSYSjERI5LYUp5wdlWipr/4TQQrWI/umXrXtqhgtRzIX2L4Yxt0RaneX3
luSPFLqS/Wrb1y/xa3c3uzY7wAb3SjEiLbUFXPeaFR0fL2iahc02i1LjEgMm0NPhoY9zANJkKgwZ
0384BBGsB5iUKjJNiO7PLWnZtC8FgiDe187AcXtIwGloxtePkRiCsKR1FIqVuM4sZKrsA1LdDY7j
ucQc7CLL80zeHsExP21TVOJLZzASpivTD38UEZ6yEIUuUaLO/6r+CFcZCkkBhCPn1VqgQkKgr6/T
JFZiUFnnr8hO3MJbcJ1WFE4UsfegkjF+K/RQHAsAsQ9QKC8jnCfV/CRPO6Dvb0dIfYCX88d9n6+R
NMx8KySnQAUdUNNgh1Gi+pfKodVj8A+ApsiaUjcluDagwZ3NIQazKmtFxTDPsfx2rit2+17nMdJs
g4aGwnlnyEPBOxNnj9xLTQAtqAWe0ZAlRbYSfdaWuwAM9PNlVI5RZCqvDIF6sGC2OblIACo1ANlR
Li5uZ08m7i8+pPld6sY2d+WPfYNBXJRKKGzPhV6ij695xipmlI8LlWTCxbhagV/oHzCL7RNUA5ki
EjGbkalMY6uAXO4pY06xcer98PGE3F9b9B0KynbCdZ1oH9OJImw+gGQUx3b8K/zOWoT0qmzqd7Vv
qs5yGSI37R+/XJcy/R+1p7LFxWYHEsygZrpNWwDgz4rSN/JCyvtDSWRqnvm/CZI0MH/gew7b0p2s
p1dSj4r/KERlQKVMyjJXoCkD5Y7OJduZlIKDm8wOL7TcRXYcdcSUc0vJanVb0mefzfyGvfVlAhvO
GkbBOFbT9fO850hu2fXnC6I/F4BgsFkQshqWOmZUe714KGjRh39T7gMSusRU7Y61eCmi0840/r91
W9i2z8eRiHt6sqaDgQLMg+gQzTbSkxBaiYxuEpd83E5Zx2UF81j9uUPlZKgGU2UWjJ5e0/5K0xZ/
Dnos9LsJ41hXNVGupNZ5jc6Yu0uu8Yxv9JrvMvKqOSTl1F9KjjpGkyq+YX0wyWg7KbswiN3dlbxJ
B/X9DitX8I5PWli5ZFoAYGpUCAin/UTZ5mfXt/sOgu8kiML8hz4/DbijMObSKcbgBHiVEe3DRXmD
6evSb3KxzZ//t6D3+Fj+e3JwAYefCbNG9JneWG8aRegmMr8ctvj5smfCsOiopbmTiYhV8SoqygMs
+5n++IOMTXy2bIYx8UpJDDtJx4A9aF9kCzdTxmXSNn8wKkRoCQ+DVXcwS6DYezV7bBHnF02Ghif+
mthT11a8//JVTtt36+7m/g5HsbCElgWhE80n01ypduNu7UH0BuFQk5URJy8XUxI5Q7HbrH4wP2M1
2idBygBN5yGsVR3AFlieDgg90co/dM668cGeXqNjnNRfMYgAuGuc9mt8wwTjHvETmCVLkzpmJSIy
1c+1w5urGg8KHm/7Y0JBRspZzLKlTxI7Dy6/gd2XlPcJl0KXDvVSIrftBkIAyLC2/uuHmAX7Y4BV
O7wUXXKpDErl5vnbB2GqOtzpqUPPV6503y7fQ+bIqI4/ZxNeI42gKTivopRtyQ767pBLTGdI5MRq
wW2ckuelz6p4s2fWmfeNyBsTGx+0V6TFWfZ/5yFxH2coxPbyC9dUTSIHrs66oKRv9DG6TH7enIjA
AnCS/8W2Qnl/Z4WHgV+FW1Nwj+ytZn9q750fY/63lRP63ZJfIp44zixtmt8ugNb37YjtP4rEL2qB
hEkQlBWxPWzzvpcOjwZmTkv1GXU+lhYH99ImJVFHftDju191B73UozFFi392qf//oi941Rxrj1rG
y+5Yz0nj0TYBAEU8g5eLtuptbqqwSD1Wd3hZJ8F0Xr6f2fE3wnmIsTocZhceMRVcm1665q51hYax
LXYGluKoWMRMl5WOYIg8N6v0NzoaL4ETRn8DEIsSaI3c3OTXyWmD8msAr09LvejRWyV0Ry5r22uG
TXoqIRj2/LEmgmJEkzi1LXcRIsQWhGfncmOjOoRlXnkQK+3dzizAOh+JBfQgEQK6W9xcau9SXMYj
dTs8MTjmDFOPEQpJBSAeOkmI4qTmP95Nfz1oT7Acu2fGR45g17qQmKTLKXwkcoO2AQkbG58Gau1J
lxxUKelORHQgaERMhetUinm36O5lUW6E4Xmkwy1pM48zR5MXJjVqBykChxoTYXTYa3v+rlNVIIGd
b/mIOH+VcRbSlXP0occdJeuVDI117avtoOmHColxmxAeuN1nMn/oYaMB/Hww1RTpTx0q11lJrI7M
lC+vYaNv/5cdeHg6H186gSdqSd/Q16ByYRLOK9kFroPmCVaqgPEsRqyLawU/98XJYQ/+rkDQLkhQ
MjQlFBO7P5uHxSDd0PVXHIyA6pYAbm9Wcd1fdr5orIFEYSqRsu75JGjFCF6omj8ALOUzW0BUXlFl
J2jKgXfXgjRfBDhiXnR3j/1LY/TjLeEGmyJdYfLmJ7aa8drrMSwsjm6Uq9kJFWbuogXeCR1mLlQ5
ntOaP6ZDDVsqfIKWi0Ra6bWRetxR0WuanWIv/hv9KIZLZ0tcXgM2VnBjjnsZV12oZHwjW8nFi3/G
ewNZZrqJeKa6WgNm9aqbPFICrONmsd5tlfsmInB3sRWDHdzLpbY8gTGg1dVI4vuJVQi/ePNWHaBk
cCfhJqofwNctEJd+95N4GpAn4OnJ06bbyk1DurEsO2APbIejUtQHhLe16EzG9EXYwdOm6UXgG7tk
N2Zlz/NHuQEtRm+OXgE1QgTzwgj3izlg4OtRKKH3y1e8aVsML9kd3shgLklAxpDF4oWEJTXc9q/U
eloCF0vNpiVJFMjr71LEf5201jvo/qF2QkYFh6eaGfjAq+OTRV3RcR/lm3cLYvnDITXTaKeYkjgA
dfE577BEwsH0dS796GZaQXsLxwLCmcvriv36hcMzKW9smuIN3j0IxbO1hqCWWJcW36PqG0Ftq+5h
Vnv6V18zWDASh4GkZlta7wzlVP6047qjQEQ7BukrwURlH5TOqHI6nP1uz5+quX4mukVNJw4HZQED
/rCwUkbL1EEJ8hPA+MzqfgjzjqnQxCX4JEwiO100JY6WcvvOJPRF0FXdmeM/YUPfY83XFycuw6fI
SVOzkjce/JLa9YAldI3x9w2nfZievddRSEoUvCC6WDiKoJwvjSzhy6Ro2aDNJ6L8Q9rFVi/HdUlW
AeFdqc7N57LDs4DuydUGaJKN4y7+M++Pfnq3sx1axOwtCH6RmDw9ImJmYkEsTUgpnBQFD8Rb+EAH
6j39xVRAoJcy8D1JJIZmff3VVvdT+TLB2OPeWHdYNzupONNIIqx5dIdkVQxMezCQvwYUuPSbJcmB
vCAWK/LqPFqqyG/qpqLsUeRzaLp+gLE9raS6+vNT8bOVOTi2TaBYzFNSC7sMSPhkMub7Vt9n9ffp
sYa4Y/yIXLiMyIe/4mhvZaEi9Olji6FfS36o15bM/XD7wnVmBV2fT4hybvIknbdvUTJHxNJ40hQ2
LceUegejGJ/91KcgxyGYJ5qINH2tYwKIM/rFPS/Si16AdfyxH4HCU6jeox+1tHAjP4NwTGT9oYkg
Xk9XgLOxa99RXPJMYY2ycImTVQEwwyYYpwaNV8c8KWlzvu5SrZI6GUictE5OfMYD7DygYOvothTg
U//Xc4/pS+AGJuAl/IHVQOPywTwNzVt9NcUUulcW2AauPrm0NSIooM2XQ6QyqfrgbY7Vt6LIbKwK
VZwj+fqzl+KHmjcCnpYJ2EdeCRekuENgtItwWvcxVf+pVvdRa5zcpNxwZ4YIFJ6ywluBulgIBUdl
6MnrmJqDbh9cotC/jzlygkD87Bilb6rlhDl8BuHcGIo74FW3adFlNq79ykw6EZeNODdTQ/Ge96ia
fVQQyz1DUs/pKNv0VJs48rf9yP6s+0f5N7oeeYJT4rvapqY9CtZHhRZLBmG1QAm1ycplYi5dXvIf
LHCHN4l2bSGLOnomQUInC6vBmDmrjJ6ZZVoCzMRjGPd5xU42etgmSGF3fsz8ZjK41AZ+8EDu7vtx
A/QNJ105mvivASbzqYq9/QlfzefDgxcF3Jj0WDzGSeZbEI3szgVBvJauwuzlFIsVVfh4NK1LJUfN
67W6PgsL5tN6Wx9mdFiaOgMTrQHrezz0e8UHAnYvXYcPSxCrX/0KcExOLCE5c5VIrubocdoRisiR
JEcsnfGDqm5WJc/u2tRF4ga5/CjSG4RofDmXbH41s1JFhMTwkU0vCBvqpwyx8zXlZmJlvZCa346w
9Abtgk0KOGGuLv0BoEwZ2u77oOY8DTq73Sm4yU15p/uQONmHHjJ19o/KTeNZ0HEBSTMAZp12/tQr
mUl+ARnPFG4XyexcqfxL/n94U8wTYTeUwJDwE6xuGpHITdQ+8P1JcJSkvP5BCl46raI0rO+RQi6W
4ky4192kxyNzpV6cZrC+0JE1vPseSpUbo2EBF9w8fOg/c1hEjD/1VisMaJrv4BDhEZj2gPaktNzb
O8pM95oNcWznZLqBkt5nb+lzBtEQubYEMBLiKoJVQnh3xudwERACWWoIH8yxlGKto+KJWE+28FLO
uqCcyXR5+vqVLi4XwTHe5ZT9fboGCZOvpEroyEFOpZV7BruLSRyXXVXtwLgLa6cHmrRDmgpibaxo
z8eaMzX39qHoSD54s4H4S0W111etWFaDyUAKqc0lODyqCKH6tE7li838SMPkc2oGB1IGrb7xwmNp
5jESdxRXSy2dgQL1OP6n2/1U5zUOfVv8jqbglSGniBp0W/1ajnZDjJp6Oxq1sEG8FKhsewY5oUX3
lY6QRAq1kbLxErU2Cv3Q+yoU4AxToC+vQTO6JhKO5cqSecfm0xUIgWDFhMj+b1sZrupwH/WHGQxA
6hgXMObWYZ4NnjY9s5AUPykA8Z3M/l8mAHzhGjfZSU6VNCuXfYnksPB4CnwBxn/pLQYvXkMcwo9l
pa/jXi2WPp5FkWsddX4vtfCpwvKaNh1SAKK6MHfCk/seow2XSo7YZsE0V1j2oNquKAw8k8eJ8jWn
vX6KGMeg++nuMTjochVkW225Uisd2HMyuen1BMGjerXX6J8jFxZNmzQnUNFNS3zm5MZ68YURItu+
6fzx+dWOggLfQI4qGsuJc5/pxcu+Zx6HmKFUj4DuEeaZ1+V8SfnrpP3XOQFnWEI88Df6snPAG6Hf
hhrvWylnVKvQ7W2kwtJ3R4LdHJhBwrrgRkRZ4Qm/kOkVKzRzn8XIVU9Gs6yUP7HVln9YAzhrBdjz
2dafjI4ZK37GdIEDJcS7COSkj02UNAAdxRm7k1QRxKpXnK7De/Na6XrHeoEuVOMMqk12KxqY/cCA
UAq8W2RIKRHydn4epEM8wzJk3ZMfMlSNEX7KCpzIZNMfEDv2RFP2O6ft9jkd314iZzJ2PlioBd3g
QTxLuz1MbODlVEbH/0Lh6JU3WkObdnjIVWWFsGEPaKdeJlsO0tfU9crRDPkb4oJjzPQrqNxEKouL
vTZSMle4MW/+Yt8f1JDevaLGf2Mjf1ICPO7EJDzNIjVGiucl47jwmHYmasVKTb9FvE387sEYrVEN
lGcN9IqzTLcwBxb1dXQQwm/oWMQDwgeOxCOwUsyoIL9M+/0Q+/Xg0l4pjrlJExSbyyxDvXnQ13l6
OqIugF580PFot5JtE14wzTCJE9wqHuVBnZKthhWFAgsFUxl5HUc4QuedIJRuPbKJ7fcXP+XJ3YKC
n6cB2Lgnwp6ILi7cf5VJFPXvrN0R95cAa6IrgCpFp4wDW0w7zdMEu+FkL9YNzmjdMWcSlB+gyTJ7
oElKOtyG73Eaafsk1WC2BxqJBBPPOy7fmIRKn90NMljx8CRHuKkDfTa5nvff4tw5ff/C9kT+YdgP
Q36zWERmYcSJ0dMnIcS7YLxSI5Yq04vZY0PHiJ3X0jpuEiJumy2nCABWCDW0uzyOQOb6VyjVr8/V
WwHjMSB4vr4J+6E7E/p6EE8L11SBKQ9731bhDOlroRsqbJtR41CnEOP6LPbicaabgsVt/A0+mFii
Y5no+eudb5R3R2rXBfEDii+rFcvzCw68d1yk6hujrcqfgyTo9QOmjc2kdDjZSrUF3vb2EJhnvUpI
5tMA9rEAPtMArM72rau1agaGl83crMGrizc4terlh6B4jODXaX2Vd9yGHPaq9A1F5E8/xhaGS9p4
Emf+iOYZDDQ5NQSqDAa3egnUmyWGdN4uqOfZiRoyfkP5/yV1zAP9goOruKL4FirPHROdrkJqDew1
MVEQQ1LFIjpzFA+4w0q9JHOROffd3kBDqaMGMPf98PejBrgPLWjXzyywdbTUJrrWYUZp0NWUY82c
qLyl0GK7CLoo9paAk7AZ+5zQmoQ+krO3CLrnZye206ZK8Jz5UF1BgPR1VM/Bt03/AAAcN5DiUpj4
7lYcdS5ooKhmcK0sxYABK1aoyhyNgB8DnG12uLmXPSw1JNof61HSjnhp5KBWD9lTUyw+Lu1IzXh0
mYRcltqDAdMDyGV1bzyc2nUHt6/1CfXFtCG5J2joelSc0MRKrsMkDPSEnyZV52ZOQEihRTt1pyRr
r92J6GM+ucink0Ha/iZQDSRVA4u/B6ZH7VExQ82RDLP02JIjxN50BCfl9hlnSTEZjCV5EEIBmFGs
+6Hnq7DSjwIEFOSyBSTFQgAmA8f7okfn0NTOZCWaBMhx1UCXNVfbLMnG1Fm2tXiUjsK4DaEma/wb
T0lguA8/SA5hrPV230BJkuuFs8sI8TswLd6LpvGK4CvRUSlLx9TLG2uM8xibISlXkutOclPd0UAI
NVe6catJQbcRuYhUabeKMlVrLTMF8jzQFrYFQStRTIP4HikjYnFN1EDCl2ezUqO2lgAOrOKsIiDv
wLliotTCiwSNKRLkNpnVSFY/P3nWrM+0TZtKzYURBgUD9wVfPybP0LsDn15NYSymfYtSOWR2gp7y
Lws6P8cwSRpAvAOVGKxks1Vwj2FmYx8O9R48uUUFfOooD+aD49U96v8AAaqBaGjc3bIuSvJvtb7S
ejlErnnbr3s6U5mWUR7uwEJRnadqfvZi7dz1NP1ZlDKq4QNpgHo8GoJ+Bv+UrDIjUb72yRibN5QQ
Yv+JkF0l8uMMApDOBJGSaIpmdNk3Ewkb2Qy5B685BeJLKFYZQpDHL1wGL6BNO3WYlV4e6vvAtRZw
yjkVO5X+d9d3R4K6oTru2IW1NqFfu7YBc1DYAuzl1QZN0Nd2zwbQCgVS5RPEeF+Y+cYZHAF0kNs5
sVIyRIprTyXuwyegy7ZS9UtrM7v8LzB+R9YPhtGU8lxl/j7Nl6CqahMwled3mVVj/o4Gry39cTN/
2JM+AlwgREsbFKs8X9kVxtOurm3KVRpSvYB7QnXBVwEX06FHCQeWrS8nSjIlrLOyJolHQK9vU6JR
mZxSp2rN32QNjsKY+ot4QSh3kWGHJt8BxIiZQTWLE+aM/Kw5oYywvdQPoNXp2Obcp2R5EItQqXAU
VasYnr9oVjIIKidY3Ao4VAcemfxZmik0k4qWzqriPJEkRpqJlEYR7Me09R9ExdgPkeCdbwg6cBAz
BtECHtK3ZIsDhYW5xOXeh8c1+dvMS6FjpCwpBaGqTnj9k8BffovuwXkfD/BciGnB5BxtZLSgQzHK
YLOwIvXulqU2h3aMgq/i95j8a0kHtSWYs81MNH5HX8qXqVc9b52VPkCc/tJ9nhbLEzJ5cR3jZp1X
Wt9dIDSXAWSNtkky38B+m9yEKpzdTWmg1WSDKOKSOw5PcV4oo8Y78rWcbwAqAxIQnBR4I98KXpV1
utxBh0Kme+8+6t8o1DmOuYGALH4+j8WZxdptCzrAssQLdKGbzdnIR4X38ebfvuYcoUJEevIDZXVa
n+jLLZlmaFK47qV0K7Hy1zf0GUMSKTRvbr/nPkNM1M+u2Z3I0wQvuixUljsXF/0HVxfVLeCXwA2H
/cDvRMB5a9sZJv5QGxFl9tljlimh62x4rmIIWBDRwM5fVId6TO+YYU8AkPxQ9KSNwzW7m6EkIgud
ZdcEYxjjA93rip2bDqJRrH4mDIe2/nThMCA7wTkBDiMcjW68UetcJo/YLSXYLjj8aVM8j4mrSdSi
dMz1bgXtibNjXDiiCgXl2Iquyh+ChsI3cue8uNpZ6YJbsAj1t3SgQSfWHQ8DY7qa1gIUIykE6zK9
62j9dJrNfh6wGBNdqelN2+61y/74Rkz1hvAfqCa6aop53MDsh4S7/T9mdQC0QRK56JfqAiACCFLu
nUdu7XL8A/RRQATH1Go/skXOIGWYsHTfnHpDvGSWsyFVrCFTZIsJUtFEH+1qQDfimsUvQH3jBmkt
qNCDtBdnkyU/agDperXyUoUNnLaIp8ASLHDVLO/tJUuG2McqPxHvMCHLMJwW5MAMOL6ntImao3Q7
RvVChemway8k5Tpi2a3BroEyvGYA2elt3H1aFn/sHpO1DoDErKl6NOXw++ylcMt73i7X9d2gWhjl
lUsJ71UAA+/82LvbrT8BdM+0kaqAR4Bx1iV9du9oxh8HknK6qe+aWplQ+gLeBPtLjS+mNJzpShDI
zasPmSgwQ+nzGTHlUTY7+87Q0OruiYMC+q9bEqQB53s+Cfq9e/3dDcH7e/ByfCz8yuCJz935hUCB
Lul4ADfDrSAn0lFHkeMnr0/sm7A/oidrFFsRiJdDt1zcRJ1DiP5qTjEp2Bxx4NDExJoj3vCE+T+S
bDdwfgDqzNZ0o3ntOn7F0oNKbMy0HsH/1wjMot2v2acx+sr9ZcIfD3S0oVmf+Q2n41mn+Fes3DL0
LjG7hvzTUj1+30uG+N2jIEUvlVO/7r1/WGF4i32w35qTjbASS8nP7Tx8e8yiW8Xxlq4/MS017PEr
kd8tvtr6OHOSyY+yVIlyCQjIDhNYFcBgX+sZ5zmhR+OP4nZSrbvh44HnHWSuC49q/E7pbe38bBO9
E9gWkkIoxkWwSm+uEAs1bsg34tsRkZq0RSksDlKHCXlE4XIDx5TBs5qzyGQmJIfvZPkDcBSkOtaS
btCWbFj53AJ5oN3aj1h2o7nAA1JMXK4M1fUBoc89HF5SgTqNH7iAtV3EjM49WMoAeTRLxD8MB/IL
9JkgqWV1Asz89Uw5QCtksjd6BqyI0grWi8nAe68QGT4ts96NNZ7uFx86+e5GIrddjWizT6y5+ixT
GWBH5129AaqCH1vZLFpwp4Jy/8ulU13PLeeXioFTNvKQ2zNwqg7KXlQsBBSMGRt1cRhpBScy78JF
aOWtazl096L17Qy5tZiL6gtNR1aY5x7sf+zvwDvaqFUp/SWi1JYbBTfBo/XlD8eLM8dF2XrB/BR8
uyoEtZ9v/DHQKd9Jhz7/ZqyFj3EUVANq/u/DRpuaIUAzXtjg/GZ2sUmNN41dPUclvf3Hd8bF23us
VzoLTaxMSrnLeAMqGi9CKA/nMkN/KhywOg9AHVHEcphkgs3gFu1ckomcqjeYIzk9t9J3jIS/NWYs
wUwvEsfYY3egLFBwcZzJSfZ1sMUfDhwJvPp/HeRFAxrCmWmkWFtTT52GOOuWVsAcs+p/l6Pnd7uF
5IGV6OV6M3NNkNK8ok4hrTAMwvapD7Im4R6Su6NS5xV3ETeZNrVmJwtSu8nfmvs7RuscnKLPOyxz
SaPzcZTtqDER+s+GK0e+S9MdilqZvzNQHrP+FxhJNv9OfMlGzNOdF5W09JZg1fV6iHDo6CynLUSk
POJq29ar4QtISmUFO27NTqxGiMA1pBSTd3eZyQTKZAxfhq8f5AQUQFlbLpAGozhyeF9Kf+PfYTEN
loCsARfJipnUVIBQN5WILE9lK8G1+UmBd8Gu/Lg81y0B/mF3hcX3elm+yUTomaDTxEQTLayr7Sic
ZXXnjLtYSS9qyP72vzkIXQa2DGN42uOo9+tKdtcPFKnZGfosSUxlDaLNguywf+KZCSlpICAwBW9t
Qdf2YBXoPjqloJWanpXnS3O9dgUpQ1WGLJDcUe2mLVdUQnFBADtwoeCQ1ZLCAL+Xpj23IO2LoCfe
7LFC9evdfBEWvWpusYDiTngb3HXKgwgGS9XCwhKYn/PcbndYXJspSa3uykOQfFo3XwHHbH4x+sNC
7pYGpTfYSN/UxJSNPIC8e6rhGVYsyrP8pV+59EHqsBulaiI7+uiCOtjeiKGC3W64OgU/x4bqsW/1
n8naSUa1g3hmIshMRFOwJYjixQkZdjXCm2mDrWKiJVqMd/t6YDXD8BYVmnrOhigw5bzt7kzWf1zI
o01SFLQCf1AgDO1zHjic3RmUU433qE2qiE/oB8NcHPrgsvkknf7D2xbrjt5myJs2T/+lCw+7ZvQ6
Rh25Ws5NAmwNlMnLlgRxQwIl3aEB53Z5ZMwS/P3oyY0OjIDuwL1Ddt2noTYSLMmVYgPesUP8MmVC
daoLodpDLNE5Jt/aqqxXRXem9UzquVRfmuJulTJQcm+4+nc9PfdlLfivnRfAkvsNuEu+CPLMEZ92
5mp5uRGqmAckFrqggk96q/p12Xmcyc3d/NDNkqWYLON+VDuAyhufV22HgX6CTeM0PxyNqkDC6FPs
H+cnTjaHbD8+AFguE/EGMAr+Eiw1IB1MMbUZDGKuykS+lLM0PRcuuUaG+Nf5odbleOG7sd8Wuy4+
PBWA41QXF8A+Yt4ibaSt8qNmROQ/7zAr8O0o7YBNNQzpuiHxtIkY63v9FDQ8CKSIjzu/qyi4GAJ4
M5kSnnqo0sRNpAgY+yz+mdnaUN9n3R+Q638yVM25dbWHkq9s+KyhLzsrbUtWQvdrlFDWPVReduGg
458flNuoHJH8TIE3rf38lupvyNywY3OoPQlxymA/JzzB4RdLifnaSkoyOop9H8HAxbHuQ7cIpiUR
OfYkxyhdxJ61LTFsHEnhs7QfWcIJu2vptF5PeRmV9Vo/FDAtFUIA/5FTiFURhvc9kwzCs4uS3SCa
fWnfKRrJ9BgAPewUQNdhF7bI/eOhXpu9OGHiF6yzbWj72WcNA22UUN92HZabZwAzAX6PUTcD0VJZ
4Fs356bNFu6NFv2pSU6BNKtwd0qM6X5epIXa0eNP/xJZOzE6mYGGgmt5HYc5tOqMUHtG7oCOtGZK
rb9blSw+Lg9HbvLG0KjslDC4RIJ5HS6RRcx9/DDH1SG+dGjFIKsg2YEnGTuaW7NXBb28dWZSJwNA
odss7SHxTgFfEGLjIwOTLVuyUgazKSDUgfJuynNtW/+KnSjjbl1UXw2Po79fPWYxe0NSrRCWhCGi
NX2b/mCZa8uxrGAEU3AsGPTJQMDvTEt+3wS2lnAfkJ0owvs8/17AY8TqqaQXNwTnDMevD8GOzlZx
dgHX911RaRUyeYnAVS3ZcLXn1IkzyYCLBP1qQ5tCQMfka4MM8tTnlUP9A9mVKRQg8SYoPMiwSacd
UnvhDsekFx+6HbkFukn6y19dI3bgKDCMH3gI+vPBoYnupyShoV0ukeGp4K1p4Kws1VTmhqJ7ZwGT
o1yFh3hCU20qF1hZ4bEdY7FxKG8uXL8OVQGW7ZQd91qzQFLBRT9YUtMxnkbFqdrVADNnj2gc7PUE
br1Kc1GfzVuIGT6eTDGleOMqHoOBvkkrqNPRCO30paFaubSRdqjGy8khS5lVBTRz9vzZS6rDyqw3
IQsVUK1GJhZSOCtgL1wVl6OhOk9HjOSvuvcQ6HSPlh2L449mJ0GSzuNeJXFHY72YxrwlCNfQr61k
/F0HVwX1/XyKjaF3xoy+0+5ifHIC5RJn7MJVUeoVmCijbVnUlJVdKXJCRcXQZXFIXkBKxVZZwSm7
7qSfWNZCcMLv2w1xlMRpnP9uLNmUahfCgOCMu9NsYU7vyJV8y58nSZzvkhSeHEYsJUWR73G0eW8B
48hKPquOvV1n3nkU0X1+Z4FRusyQsY6/gZK+m5VmRg0Z5c1+t07b+9AP36nYJS5Ugg42z/j+M1It
HialZq650GZs7t5NzerZZnumiwm1+RK0nWx+IdaqeSLc2WlaWAqpO5gVVQA0BHZIACoo122fvRa5
QxpL7w8rbl0eX6B6tKJEJOzNGQzt3Qew+LpeFzKuMNaeWyAlWUrjqsl3ni3E0hc0biJz3q3cCu5m
t+h0Nnq3wCejMZc62LDs+baCC6Mgx7DFOE/6+mbKMhjI5q7kZL9ioXELJXMiiXwOKL1KXJ7KaKem
kFV4Y6VPsTk9UbEEFwhMx3T76YVcfjWAQhht6QXTiRQijFEI0AT9q+dk6T/0JFDL6w7SHlj6jfp/
6pQcfOGW35+XAtxB96/4CFam7b5g6Bg47svJZIUlLzPpvRaiZbhW2CkJznFw0Jq78ulLF4ZtFbob
VMLEYerEMCBB8FQ6EUm5g2S1KU6XYSdwf3Hgf2YLGF3Go2JObItzRft7dDE8zX4h8KhT02zjC6Oz
IHFbvEitQGYs0BOVJvjxc/XO4F72vW5OCa7PlwoyvjIYW5rF8ksSVp+0SATiJjI+Hk6xRD9pxlCx
wIX5dc6pTSYK1+9QYt5hVRRzrry6otOTnb5AZpmWrdp5H3JOMSI9DhG0HIdGqX057cG50W026Ug3
bCQo/WXolcUAHLnyr62horGiB99uopeNMNtjI9X/nZ7Ir2W2AokxF7HG55r6/wVdnK0tZ3pUtxPX
g0zOBGcD5QNd3DvIc++uoZg4m/BTqSeuyz43je/KZVgbBunbtzH4swd17iGFiJa/K+PUp/xWT8G0
8MN7qshz954X7XmAjP4LcuccuXdhPLqzGZqch809D/6x1sTPDwI5yUOUdPOiTbJmixIrbQ/TuvIn
oIoJ8MT+wP81Qeszb0/T6TpVB7RpqWTL2Op7EN1AaAYtaeT+/Dn/PEm/7FKvjKV7eI+56XmTNWcQ
mR7o1BmI/f/4txno0lFLkGIdjLW2dSzZyv8/xka0sJqdAnWKxon0vpQHLy2d9hGbuH5eC8yP9/Pb
++gQhf960HOD83aS+ufsUaVGqgE+TXS/IyPaGUy/jwteVVgNcoO7VlFM7yDaxWvLK/tTifb/Uyq2
EbAPCrL/eM2iJhTta1qwHCmzGQexcrk3/i0QrmeCUgwgRjvzh7SgXfQ6ipfJSsSuFnEgLq/i7Big
qrm+k6uionuIHGGYmaqfJNqemqzR//hACS3+cp7SHxvJNEerEZQrdfMJiQipDxa/k13GBkDH9iZ7
Ya3kCRPF9ZRmuPGsdPxJCgWrpeepU3hFRgkTFU93gqoKFOoFZUv+OisJhL9SMDbiOWQRkvrIOWY3
vGup6uMqdQszITkvtHKZBa45H9ni6+yqLdDLlaTcNIvdtq6T5rAcpx8J1ws9R8R84lEa3hifmfL8
cadzDppwS8cPzkqtS2eugPPL2oX2v4w867mactQeXTpJ/4394eF1FcrwmKCaPSIyAsNAfhpRUh98
pj6KJ1c6Nq2kuYuqyHtghiDSHXialzXsSO3JWrwqVbrXzRLalUSTcJfh+p/j7Cw/0WboVTk0tBZD
nk9C5veegrU4l2Y/JULWo22CzAwjZdQ0T0yR3aFfoA2fEbsvgMhdLpyvxuvC+MNiggV4yDKaQl8z
dg2KHpR6Wblsr1ANPcFYaqDn+34XFBS3KBrqzyL+Bwe9JK2OfaRUiqDXJvMckb35KbjNauXQKJkr
HXGZMLRX51oQGkjqG878mRivGo0k9tDGMWHJR83ncQ62N5ZKnQ2EnSahN/XOKsQwU3kPND0AmUgT
HuraLpJ0fjiGKbhBx2yCgLjG+TGUPjIVx06bf9i4zija6LaJDkjIuh6iINFm1SvCm41r9ivzQi6G
LWwM/RUfMLzaIwjEYUig1Igm/UA/UvAsXcfj1FnoPB9QOtDCUc2TQk8FHP9Y26p/7Rp0CB7pLDlZ
rOCvDmmaeBpJjFa7ua72i22ZuDQapptShk0yUBG1VeRbTW6Tu/5ueyl2vcle6pp4wC2HB97Jq6GQ
HdsOMUCKIegOejmNALIBpl0rr9ENdfoI3XKgJo4zRuuQkSUb+/dLusUuwKNz5fYr6k3RHgLawU+G
JwLHcVBgZazAXRV3LzwX2znRlQ6MqGshZbWNQPxuvimQkUTBwDR4Xo8SSREk6qYu9VStfP5kxsac
LROeIs7LEfrk9P788q+Y3971qUrjuakt1VifV0HODQeqOu83+BveN3RI6WgVXeSlsZMXO47Q5dnA
Q76RFoQHtfVEN5ylA2ugtCoHakxfgRAnkwzRqwkzzXY4xvQMf8+8iOa2tvxvnzaiNnxrQ/h9fq3z
kJQNINR39pDKmF/jQodC12u4oWNt7tzPuAnY/iiAEdmtMUhtRp9JTM98kjvT3DrfEI/DM9uKxKVj
cdzGmpDs6Bn/NRZRgoRRefMjEzI+5Ge79l+1JhqmFQM+oDuJYt0Wd7NFbbwKafkNAUkTiQcMxM63
EGU99FBLxrpfBnHFVnGihOzr8zjNW6S7RP7stMRLlSuKZXPjoaYyfmPCvjW1/hWUVwqswg/ZjOhz
wTMcIFhwOmos0vRDl0eoGI1uM2EGuN46E8il/oszeoIn+ztj/bx0V3dAFwK2Yg6J1zpnCqXUa1kV
U0WaHzIxtU1GWGiGt6EUKQz4y2MEF0hKmSuLv3rl2fKKYJakxqvO7zqVzv5yIcGsgpq7YuF1XzVl
VI1VF6z1wSn/PYVLQqoNUN0ZXPq0+ANlA6nT8dHKI6kjpFca1FfkUFBSiFAMclDANf1KCaCHZxUq
MeodXwqkZNPWLFJEWw/W7fc2l/gLgtaeoUqUgnSoUQ0OdMAH6VSnI1mCSbjL+5ti5hCHkqAedyHI
Mk5xAf035NCclIXG6pnUMCI7DLDsiTelqayocux9kqFwO2MNTzeS9+zzlUVrKjUXJYFVgxklW8h3
Y/UhAJUVwnCV8z9vEvMDDSyMcp4kGGOuZKg2F0tNcp1yMb3ziYAjLPMNmRbs6IzWt852iWFM1dSZ
js74Cbq1DUxV7y6RghZTXx7bt3CpYp31CYa3e/qYyToUEScvoZi406wkllxnLDlN1D9CgQglYIFB
xNPD73u+iAa5VlLkxQ2dkI3e/CAxpHVXSOtf67zQILDEE8K8ZcJdNpddIHxx2+3tJspiyQFfqBxV
GjmNiIKi7a7YA1jXYocLbII/pQbT/rXM/uwziYB8dKoWfBnHb8QD128InuqYzRGeQs4JG9JOWMPR
DQVno9e8TIbwIapy81/mvk30f7Tl4CelthPft+2SRMIEhfsSBU9ngYD9gIpRJQWltjM44v+bj+8f
srdhHsNFTboSoHfvrFyA6P46HbSIuzw+SFZx6ZgO1QDBgfXNv/iKlA40UxA9X0T7XGE6N07NORc3
7AZ6fYyZIH9HMGLJgNRV3rg4+utvrRen8QWxVSnhYgsdKMHccK2IlIOG1o9FKxQieybjJJZDHd2s
c1yUcMUGgD27A54g2Xw1medYWYPimUh/g367i/rPSbRGxzmOhfM/yjhabd/TeJb9zgVZBC0DV14q
ZsJig5/dy7Q9kLXwefZm8ghwFAiHlJnd3ShU6rvBbWjbt6jMa5lp/m88Rru/dUT2zbXCOBeG5328
vTz0wnRfspodLmZyrhkeAnMY6ihGMD3uz3nXokdPyUv8QYxQmEc+c3ICdgcJzQW9kcmkBSpzZx9K
2K1+eiAfzgtK2t01XUgK3pVXE1UzUzgA77fgzul3YCv4RTI+RNa3bfXrUtOo41d64F93CygcDL+b
JhenvRqBMWqQ3u0iSAw1TilSTZwDq9neYfnxYj1wQJh4l4ZC+WJzgDDlo+NXC3GN7Nr8gh13Za/U
/rFgxVOCss6XyYGHOywB+NIrczqFrl3yr9QQJoKhVwGbFbMJi3+tOl2KQKsUEL/nZMLnYxn+G4mH
v6135bThi8uEcQSLcNI88Vc/wVtFxgeYlctj7NkF3N1gslP+BtmHYs5kO17yFniysAaxtV8ByvXV
/gesQz1GX4GYh1ORH1DOAxDZDVVPhOwWiqhTTJYvmtDuuPKUAuD93xrM8ZNpLsStX/5wBFmDzCK+
YF1MShuH118Z4zHRxZg83RpJ5FD5iVhyaIpOnvRj6Se0phqfRlmvBZuwATNBnDxhbVB+DUi4VWfL
812beZIO4LFFQx1VcmLJUGk7UiqOgpG+9lnZ2P1or8qU1JQ1l9iHI1pXdcawisToLdrIxY8G2v4w
DQxeg/cZu70TrPSfiuULiWbA3rauQpsfB42ob8Ix/L27/i+zd98HHgyNcuJlFEV2oUTMmjYJu0nW
oxBQnB822Z3pLZ6K0RPwLL62YP4g5QyqsWVMusLNs1FQDBxxM2YpefDbx3ru9ubA8caIOnbEZ2Fg
LDM2ry+gjxgS1z3Zhmcxqb5qtU5Fb05dSz8Sr9ZDWwL2CVA32riIUwxp79sj4ySsIbPWpmR+1PX9
WslbsNCEl7EPWMolTZUYJlruhe4pUoQytFcQ3jUZwqlgU0NZs8MtT7wUXJr1zxc9GZKW3bWlPp+z
LMnGZnl/Hanjcz2Z34B5ate9cy1o/gg3aabGlnJWdY64auvuSIQwbzElIDjvJ3dr3SrRN7OCC/Cq
jO6bk99QsFuhfSaNIt9bUTV/C6KiQvPupYImutyKI/mGgZDFi6tPKWnVmKNoraONMIvIdLuRMK7u
3+FWznPJEQDIPOCCXsYFHcVDFIc/ie9nc4yj4E9NWVRZWCnkUhNPLD2pQp+vDGYKpJADzdACZJYO
N8CGNJx8ThzgAfW3bfS7O41YAqqZnoiJ/xySQIrmQDWynFMQ0bTJftpXicUVg5buBUryDG1ofOzP
fBKUATSOYP4Sh1wnANHfoJPxGa1xMyOVj0AIw7FCkFXcqLs5QF/ok/m9rl/Sw1KMuh39oleIISL5
kmmWBqj+B1TkuNMLzzc+F8ami4keX7DbDcMF/rYPHoN5VJM9vI7RC1Qo6GRfZ8Vewf45sOdp3xm4
7dtBqyMzkjAJHZBcDNnxZzbIh0qrfyc3b9CctWDUXS9vKEMkOK9a7V+SZQvjGFUpUEDJqqNjauQQ
JOsZRnmmYuMazrbMDeCHBF+98xlICiBzzb7z95r/rPsGN29YnhOM7Z0F2W7BdPz3VCQPu5VGbrhz
crzyRfocJPVs35A8oW+adhFX/VkEpSzCSOKLzsDVQyOut24bwKLFD5YYrQI9Ji2lBXyz81qQzyYq
eKC9r1XaJ6Pq4DpZxwcXFfQDikjwMO7hzIBr2x8AXzct7wlE+CTyziLKTNGiXTLsmMGLx7NwdTK0
ZQ/L0jO0UGViORKLfaSyraZ4uDWBIDkLhm0bzREl5NuoHV1HmlyYTFPERHlIOLe+9tZaOsEyUclL
LMTmN/3W/OlBZTF+Ee+Vf8JXFefA6FEf1gvJtzMhLVxdSGTA2ZTH6TUVZWl+6aaX42RRhTOlbHX4
KM5wOnVzZvM++cnz64II0yMgRa/FYvdQI5AVLKw6UhpArgv6Rg4g0xo1hKuMQVLTR5nDTA0ICUi1
n0b0toAbDwoVYML93g6HS2Y3L7jAOClUr7iquPRucXlvqQDT+5V6713YW/X51YYMOfnOpjyEApNc
dhEc0u2lZ90LlAMSaAz7BxFnpvKyuzjVZ9uwt5Mm9GhucJk7nQQO8KkuXn5UECoMzGRLatmP+Jio
8uPmp2z5LmuzQWc8Mrth7NjApGPVNdbdBJZHlFkmilm/74hiJmP89sR0RNG+rW8QjcUvF3qsGB8l
FJ/yGIoFtNJ/cf9NNjx2Ys2CJC1vOjfw6e/iyONSdjgl+ZmJSKvKmm/BNpOeiGQRCluxkAwbmeu/
dRMULSooPBGqsVdY6gWNrYGhs+6hs5i5fNFdlWdrZXLwvg7ybk0+fHetE6/PlFboJD8UU3X3kljM
CxG/LYEICqaJYT11VsM+Xrkg/RDkl4bWR5QzMQx5Fk2K0HJoVfJqkQsic5vxoAJLIbAsUBW1YnyP
rI/cmlb/oZgUYXjDtRnBm+KxDh2acHI3Ou6/NYeEX1MSEA3no4qPBmoqu04C8q4gjUX3LkRlUlrw
5swtgVpkobdQv6OCyPFSbcjVwVMPmNbCmZTnRzDH5uXhTkdDuwD0MjFekL0mTXUWN/Da+5Iy9g8/
pTwIgC3CdN+NfxJyNHrlR3NEdocPEXWH6eCThmBLNHX4mtiTjFyE4A5zfBfuySqRcoy5Fm3FVHUH
6pOMuuMZmGsnw8KsHmwH2x7RqD2LP3dO6eQqDLJiaTlBUrmbv7AytcSDl2HrHh7PQPghg+5RKhsx
2T0TEj8gTXmgvUdQcLxMW9N5gFGtUjFqDJMYBrc3MG52jbExnIRknkiDkllcr9iYQ0Cdf3ORw5+t
++zjGmMbJ4a67dkrLpm4ULUTk3zO/dVjNot/gRhyEhIQezGLb2U0RuZwvRtwGOqhGy2bhWv0Sv4z
MWAMgQqUy00YpW6FEwMstfmHGAqXCFJCEoMhPIsDZmtJMMR0zSJpGNsi5tt0FR5E/e/M1WBlOyDC
WxKu5IfdHz1Z24jO6SDUoL7jJDyQn94NA+PKblrjkSPk0e9TNe47U7UxUilTv5chZV6AlK9ZIT72
6zkitmBfBwfgDUfhgPovJtcwUAOXOdOLmwEVWRXYOZt15x9XcTXm2WCn01WaFnoJt7GQwnTBAjTl
4yxXuyhHV2k0M5XJb1STUFujIsJl7f/blw3UI9ETDO28LeQXwHra7fi5nNuZKlI3cxdeavid6Fpz
oC++OMDP+CF7oAookR4AsMoKhdZ6MzyZnxBhnt2CrlTS62mrUUKlekEc705OUcUcN43FaGV8f9E3
7hiDRU7F0O7z48pVlnXiyIzhmEIpNU+dsY1DKHcWnNdNxryhoJ4t9ZBQARVU8KvG1gvxVGA8Iybk
YVF6IgZVf0sbxYYNCF+7g2SsYFgdjFwJ3GhGCae/4AE1KewDtC81fwprX3NWhkxlBYfreXpvI+xY
ax3ZhzRYF1fBLxgodoTWfSIPf24j9uOw+AUigQ6T1U81treIaxozHnZsvFKng15IJ5/1cNp1ngcG
8ROnQHY5P+aONzIK6bwXYMtNpOfS06lXYGT7Ctj81Gh0sniNQ8n5YHgEyz6YCDB/mSpdnqBbabV/
Du32VrOJb/V6fbi+edTV//7Z8rVv4caVFD0padEOoLgyNoPB1CAcL8UE59ZZ3IharcOL0bLnQr9A
cmO9fwlT9FQzu+wsihzDPCSSUvl1LiME9b5kkx89cf5SlGdOA6pyGMdrX6zGwvJxfUG568W+lUuq
4is0Mdzzt4e+T2KnHObU47yrTO+8xCfep/IT5R3w8dRl+125pcTPkG4cf3uLceS3cMwqru21RX2G
zYJaVBuLMzTMqiBZoDfIQDRnOKK3GZ7xwhgkCFCBhj2flkMF5Oq8A+PY/SAVwzudhx1ar3KcVV/H
hpxsU+Wv8qVm2OHng9bYDq3oc5vCJcybo92dZ2OWoAVcOhUVuNrOpBprETHIvc7IFYb/9QoV+aXV
yahgBxq22Pt4CzyhM3EPGUHiGsu9WR725OUw7gzEBmp/DnMtpLcn6Tbok58+u0WNIpGSbyMCpBBb
ces9TmJSA/MGNwOCJe7C4GkPYjX7cqaNNngtR3lqed9OmkOo38Imac3E5S1H6U+dNP0KDSw7U/xL
3TibDSDII+UjOGwiV3XO2cFDX6JH6zCgguo39uOAHmRftJkMQ5KpzPykC1OApgYgtR1xuXfEPdZ+
KQ08nWiy4iQAEWFbKqOktm9FywxxRvnP5A66gm/FtOKEUzTlWpm9hwS3Xh4REkktQzZUn0WOd3V9
AsPyHOwBU5xIqoPPkLwwAcnNqIVbneauym+PiQkycdZY+AdGvsbJ9YQjdrwKDZPpjitW9uZolwxY
7837+iuojNhNvrCh6qnfUW3dL2oWFlxELsdtsTfrgdNumI0jf3XImKQuI5IL3RGYdrAq1PJgUkQD
Hro/MLeg/gYwb7OmBzG03fugWoeeYpAONHTX5Y9tHprhrefGr9hyJCtRTdoHLuPOMBsEWa9WBUb1
y1//WJEpS+dxT7LM3j4wHo/CaM5RhK+rL+PMY8dEHfk8VsxsokRaa15cMet2Lft5YA6hDcI2a1vE
Y4gxg7c7d/PoRgPXfUuD6sAHePWwwNDAYTyFtD898Z2D/MHUizwtzcdCbxTa3fpJ/SDn/NAvxXxG
5Vh8y07xtgwEOyBw+MIwoi9L5V4UwRdc+zTCAEZXj/ukT+p9qTjyDGDbvbjwSlcbB17V3upw+5pb
3Tg+hg3b874pTHC10y+ge7IRInjYDU5/Ff1K2H6SUeYlv7WkKQWfpN0/psW8k6PmDcehxHD7przF
XA5wUavb/AgtcMlwtxzLu0cJ9HazMMsjVRvIOkL4L/jrBYTqjjs87/fMjYxPbSNu3HcyrWxBBUlK
QZegAJFBiviaVbWmOHP5GO3V2Iit906xYiwjdP6E/6iGIqEdiD6HhwrKdyhBifbN2Sn2IKSDU064
ZoxwB2hKdPByC7sp4FM0LNc0khfW/g4GE1yfuLvqyPoNIlt62P0bPHZpT+6UOUkwWOT9q6S/jLfv
BB1S9FoqnoeJba3tDqc8I24WGPcfuevAlAVrbS+BsvjU1GUgTcloxVJBgRdOgF/RnEnxwxGUncRP
cSeehQ0wa1Qx3ioriOIhV6A5h70/ZKbY/FuAEqEqkrXjV9D1fFsMj0vGGac+/yZvfcNEdjpLU/p0
b9xKHa333wZjdtnW4H8ACyqmx80/P5oBvH/aVFZcoqysb8XgsbB5imBc9DNiPsCnhMPYZfY0DQVw
sdRlwuzsU44s2Zz3/X7ik2+5b3ne4ya+0TJeQFR9CD5mTy9oAd6odwfBC5q6AxFaQ/z8rdNHIFQk
ab6j8P16L2hem98WdOnVHLBRrs117zLfEjd6hSE496mjKGSVX0QVwtpvZJB5JHFmYkNkdwtMH5Kl
b1suxQCzXduoncHmw1wiz2jlMXnRedIsWd3kc082MQQP2Q+ZQoK+TSG2CsPQpb0s95ze3bEk0ugB
5l8qAK/Y659zWW8baOJOypcFP26Bpwya2euyyDEEFaZw77tFZB9O0jjL97hnP1kohpXznyIuM13K
n00s98CUL0DZHGNh9X8ykDTRJLzcE5i6jCn8kw3wlklXxT5Y0MidcCSktbc7zIZws0V/bAIivhjO
p25gtmMllodgEofwFAIbYUjXgXzcXwDEMMShQnJ73lL22BUQ/2wTvM7ygTn3RhsdyktZMjW+bDl9
/JsY/lJfKk06urWlyGpcY3m7Y31hXkR05YdJPW49uQoZOW5yzm++P3Qmdw5YDGzTHm1Po77XRZyF
sP2JLs3Pj8XV8SQmX1fbnx0Ff8D3HSZYygNJiuBPhalJqWtZwPEuG/e5M4CDcRmBdtOUIR1DU2nm
Tlr3V/TLPBjcb13Mv87zadyelZNI1U8a9xgRr5/dDKYa0W75lJmcJrLrTjQjXD80d8jqwH1oyel1
gFiy0XUEg4DDdDOj3as9YPMOy91LR6i7ItoTgqzoRfDGhI6qvtV7M5dmdtci0V0CP01n4smQ62HB
MvRWzFpgUdonMQw6Xjb5Ym9jfQl1EbxMnVvXSYn6/iXa2U4MVVppP/EHM2FDUgCQoiSaw2IwWjo1
vyWd6ly8qnbL9Jph314kcOK6haOPZw7O4UWX0q3fQ0z+5cLpcCsk8WLS3q+xHCRPflSAofVI7kB5
Vo7xKBa8yUBlRcQiM9V8PoJd2HVEPT2QnpWIPWYif63ZFjR4WBYiOpdSTFMwsH+Jx2a5+O6CE9Jv
cK5vKOONYWvVWN4F0wQ7NxZsWs3rKrux4Z0Xm1Ay6L7fHj8wcz/vwCFgtW3FB81P3Y4XmfiNooyV
g7+O+aHNtMZaYUsAFSnrkPGgtPQ8HuVw1nGJH4nzPBGAABAZhhIbeSNhhO3OlOLoMj4BQicwQ/KD
8nwN5pFTo/PsT9tdCEAEXmQNOhGS8Db1X31Au+H6MMoM9dEYgzN4xiTmnqfFQxQj8zI+7PtDGmU0
ju7uPF4sMnpRXjfwTydK+kvE8MyapkBLl+GEu1HYOKHUE7YrDnisKErmjqZgwPik81XTsr3W1KJT
wDcNJG7i6sqeMvFNq5kW9JNR/QhGSekUIgpvL/xUg6MmZCBiFEZWV9t+Gfvto3SY96634G8yqvyu
QBQhJFdvlmBGtc9OjQKmNKK/JFOfQ4ivJqGSdu61BXEnl2iGn6qPDZTw3kfiMyyG/u76rm3aS/pF
IVuAmclpMC0ZWSzYRAO9qeWZbq8uLZk6khNX4Csjy5lAvo/JeiNPFka3W15E85Z+2fU+GxwLLVQ2
e1ndOHkTcNRXec4TfinBCOrlmC09lcmSpP2hAZuMA1bJz8Dw2o7Q2OlHeRV9EolTGX0yZSZ6Dd45
C+yKQP9vDtNRREscK1nCY4kPwpQai291MepkQ1S4mPaE4MY0peMCBr5zLgmFXXyY4KJAfPIv4NQ9
i52FGDNIRp6U+OYsVoNiboezMI2NpZY224Ua4J+vgqBe/nUiMiwxwvREJNh924MpwTxRy/W7wiiA
rK3r3p4JJ+p6Jx8e/nrxP5r4yWqaVGbhNHn9I5ptjcmzMI51dyFjr5CAzq7G2amqlKjQwA/cVNeq
mo/jeacIz2KeKmih4VWKAPNzAyJjJMRgtDIl3YGKcVbm6QEKy6S6S5Q3Otwjwu57/iMThg6TxCO1
twfYN1SOXBJ9+eZaPVRghjgKZ7UCFMHnbE0gxxyyPNVPa/SqzOV2XxJHEJr1DXPkkTIRYB1g7PRE
iXwftGMAFdIPAK35KjmKZJoNYdhWjYz5gNvSLAcV55S0It8AxGIHalXjc+SADXidP0cL90ielM8c
aoB6HC+QamnoY6rQMS/059ckUQpyg4O8hd8TeiBbcqjtXBvo/0E7V9A8YJ9gTOutcfFdZGHSh3bF
uvtg0ZL8qzTsLnIA5YlG4PFBfqU6uRd5PLugcF/saFoOkSkwzs3Lm1rxoSEn3YWPU8Sf6uOLAPXm
Gt6uxUev3bE/S1H9dW6PtxMLDryFMhm2LTCSiV3OZ9XuS8AzB2cQmmqx7qIJyV1+co77UJgcw1TL
BWvz78mcYQHKlAXbxGK6pbyuCWyOIseGWuOobFuWWTrbPHWh1gBvKk+XAEDzSISxyQccPY4Ypbb5
rwGXY9KwOS4QsbIPrvX1UmkxMg5phW9qjWBI6hnXUMAs2YevWlwJ1dh3BYHj/B64cEeSn5Rp7tLq
DNQhAL9IJO+RTosQn7UxX/pzrq9uhFmDMWjieWc/CfDCogPcRTWlDGjBYbhnO4DC/qSifH8bE02Y
WSyjaghNMeNrQVPDfI7a3yN7LZogUM9lALZOP1aYa22YN7ukQH8aH3X3cM4sECCJce6cRZI+fRzu
XDzJHf4pAwGBA2tVFgqPbYYnG9qDdrd1jdDcPWBz+yClSklKb+N0/2JT3mC5naqeXv4rDZIxSQ9b
MmOeUEyh72z/xbOMz72YlbeAX0qUw3MLXf5G6Bzkb1wYnvek6EphdZkWyYJ/aW+0uLoWiQVgk7am
ObsO1s2l18eyUPOIif7GFqDGFNCv1pWcOFq0vBir0UjP6GN2Ze+7Smu4WzX07W9EK5ziwdOYcZgp
7cHGm+BvNBui2LmUweOc1jp7xgIX1RNqtulytChq5/bH5zl7oblqIrCoI+e2cIxuzWdNx0UuyDBQ
uo3odpKxPWc5/X+cKRtKw6nFb7VMwHg58LePef17RJNGodTXMNK1r00Y7HouV6IxEMF43oFjRD6C
mrc7rdnJ/54tMuAWSOHXBISImECJKdAHosId+DUvAC6joGO3ng9p54RXMRzmB9MWlQl1paExELCA
g8Dys4F3O5dp42DEqRPVkoaGUzC9gcDavkohYhwUfPh+zngGAXFSy9lFw2/bT2/v2l9IK8Z4HwTe
pBF5FWg+iLVqqe2pNsGZYhigqyfuRYN59UyBSiaX6VQzZ9T7CREDoikNHhESxAnx0pkjgtbjvOgA
ij56BygcL5CIwdP1FukoxoQf5+diCdn0tPyOH5SX/Y4vLfv1WFQS7cSOtT+JgfTQ6IH4UVNwdhLG
AIdTBVqfXqtWna9PtXfaKA0AdnyqO47gCzoBsZbeWZJjBCMISWD+SOfLKrja/lD/ZlS8DIJJQ4YZ
MJq1b0tluvdHbp9l8c8LUmqT249GgtXHoOu+KV4mRxvXT0ZfkZTUh7pT7u4+aL2WCc13EsulDows
f8GWDYo32bnKSXlGC/xh+v0H8qknfpl630yhNN7E6r65dheTR2E2q5pL9T4LN6jb21pmk/FkGwR5
Wo6/p5Oga6TI97BvLjN1qE7eECXiKE5E0ABkl8hpwRroi1HnQtg63zrs07dsrWLDzC65H8VyP/hV
UCcNX0nXuy/ADmvJrnIMWyt+VI1rH0zm6GDFemWMHmNmE8PiaPH91h79NKwgi3qdghVCzjevLAeW
838HNMZ0oKrIKYzEqiq7tE17kBtjo9hgyKzVI33wo60rrEFqlDku7zLWdGOuXzC1PKEdV00FCCr+
UYgTmnZZ8Kpi7o8UEGnZfoP8gf7v0qCjws1Ol3X/pvG1ii9m3W0Kb7jGhKf2/MyydMKLrPFl2SSh
91CcIU0rSgTlsY4c5Y32eDn+QIHOzd/PBfpjM1YBMruuBLz3TPWHVMmKNbQq2k1v0nHB5YENVraE
51SFvZp1IMOecrJzCJ3XeuN0RKQ90J5VcnGp5CXl0pwfMad1oTkBuc7Qf2QJqXSQoF5FKTb0fCLl
AzWP1VJFZhHVZ9A5BVQTqRUKOi1NzlA9y+z+UYqcYI5rmH1uPV0m5cFoqz4+rK07hmt/tDqHEqwg
82yyNpwO1MwMoEChjd7W46HC4WGSDsmXqcXP+bTtSDOdtehLZfTTgVuHL/ANh729P1WoSix6mpVm
21dBZZo+3UHvUo1f5PG3F9vJYptReXtu7LEdK6Dur8HkYwVWeh2P9wRkTLGNKfXBaCiSmNmk4k+M
jG82DcCN+akziLBJT/w5e81O28pCbzqYDTBBjqA8V5Ln0S78Bf/4+iJCuY4tLery3A5HvMeHbP0j
ZdjeSzAvJI5FhXqjLuFEb7gv0ZcYXNCE9DLn2eg2kappbZhCPnvVxkkMw3hz0WMeiEQch390+c9C
gCrrGQ8L1o/kNWVbisKcdS1tLoXj1+yrqU0tDhVo7uMY50ggyiy+kUOnPNuGEWyNYGeNdh3DvmDO
qDIZdv6CrtwwNQlDSQpADl5BHt4skSuCmUdkmFWdnI573ZF7YE4nEBRvSgju+XpXm2uimycJ58wh
D3Jluu7y5OYBvQv+AjV3QKbGItKcWQtylGSr/SovKUdMIPL7wpKH5ufWWpbFVA0IN1DIlHDv5ZzG
IxWeRrP2UnFEOdIz+qrb/qBCcYcprAz5CHAvkp+MV23S4IClASAfFA5ihhevixhEKv79+E6Y3+US
EvOWecEJ+byEj7gf2UuVWBvXE/ALMiGVMwqiWguCZcyUe/J0I8NijFowEnbYomA7MZSaQi0rXALb
Se3seYqQ9Cp6OXM17EcK6AwKY7OHJ7EujKmEZp6gPI+hiKfqM9b/CMmfEGf4SEJAMsSYVLGn8k7t
9kGcLQNX2Ivq+QMUZPAFDaNuyozuDfidAT2hIi9osxSdQ3+Wme9LSbT50P5nZjnHix+7LNdSZJXJ
ClTpgI8EH67Ojk/Qcybrrfho7mGyANX6jGBlaaWKUjSodSy7+MONqfhNBr544yDgdNLzajX+HWPN
hZT57ZRtY/wZX7e61VOkp8Kh+NoHTS0qkUVBVX4IXyD+JSJrRdVhJ+SupLnXODfS8SA4QoRR8SHQ
dd6rbrnLHHh8frTZGBZAxUz90Fg98fiq73/5bt2FCuN2v7q3+M6OcSnCuopXmOeNN8+pBPWFiKQh
1ICZGskAScFjYOHiGowtaJB5PZsUeWfEagop7JOpimDOGQKCjVarj8xktWItfJzMgWMTVjr+dtB0
XLzwAau/qpV8xGDxcvzTbG6nHEp1QsjKedFWHZnU9rOTWfZHlOcmMwCpKnDHFVCUBLir+2CmhnSH
/TrDlRWy7mybItSemZcuXRym6M0TX/BkOkYvuHVH7/gMZk7D5XKdCuLmFUXi4NQYMenCohOOC0+y
bmzAsnQ4ddlI+J6ekty8Mailp6PTNRFmLUV7xRJ8USuPB04NXns2AgSDA007omky3XrMZvjLoEQY
U9AEsXLRaSSvE5mtLoSogE78ndrf2OZPVIFaFqmWOgvAcGuf/nEhx0XBMSMIqZUFECK/mWEjoD5r
yHBuXkNqqfIN5OOW+UWZOXIrFUB1qRyxEDjBlQsC0rse1NpyoTBcm65Pp3NhHjQMSHTTOIeL8ZXr
nwwK3AqQEpEY1GMrnrNlbmQj9DHDjd2devwT8Hv/jfhLHjQIubG8wmAqLIifqeehN7Rctau7hF3H
NCgTlT7tNTLtOV0WOyV91CqhyWjO1CrOveNJOiMaib/HQ+rHmAGuqWo+BvgyDxBYqEj4960DTidA
LbM9qhoy0Gw7Tm5qPmyteTVa9vGNDu6Za51FkPOZ3/30EqcAt1f0Ez9gL+EPCYBT0yoxb66jduvL
3bbbUHP6yolbvQpDwSeS2kFhjT7GjcVspuFVPCuDPo7b/9XKRv6tTzy+Qcis4dgTUs1SL1yRpcQ0
DLExqeeI7BW2bBrArhry4VqRby+FGlaJ+oq6PrCVZ73vdDdqoZKkyLpFD5udUJZtv1u/kpXtrT/x
AWbN1nsK7IRRLC8qJokvm/SEGktqDMXstP98s5dvmPFynTy3shgAdyPOBaRPwYkHvUihhsgMMvf/
JdMu+1IMow48ZJ7nAZ64amFRK9YaleV8W/vEs0i5f35ilsXmKTP/GWN+PhODzXTQQCbDmyA0yrEs
K1rIjVhV+U9oyveMN0j7QFefROc/swAywhFFIDGnkJBCjMwYtP5qf/Nb9IVOuTD6N8yQ51AO0K7A
LO8CFd5Sw3ZaSKOEZL2oG/dCfMPbymKP4kKehjCws+Iembq9vG56SByRC/+r5uwylgV8Zm5eLtB2
lEgIwKbe8A0VA5GFk+PcRS1JsL5fBBGiNCIZOJczD8IEmeWPAobq5c4moh/UHUbpc/0uOhVxqPT+
Q2lp9/OkXcP1v6R48n5uVpSg/t70oST6/Qqk64+bP3DcLBVyBmr54PmJzdwLCVmiel2NND01rGGg
j33iirmXszFj9BVQsBUZQfE+Oc7VNhjp/GEMTsSt0VG7bDHKijbqr0Dt4TJQ0YvRgG9QYeN2mnwA
Oe98300K24mb1544pE9d4Yb6zV5dP0SE35FOMcn68JZmBRFYmBybHlANBm5d6zfkbD0HQCZX4ZEJ
CsGpIgTTWLtkMIhG3heXSCp6QAFZgXeO0b+fZzVQ1aG6odRC9cMDSOB7BvHGIN5YGkSsgMA6NWyq
pl4eFqnsfOSIY4kN5UQaY9k63t8YVjjSbdvsiZNxkbJUX9Ngs62udX/PFyG9NpbzAiVJX3Z5FUH+
fcMtlLmd4Vwf7s3O+joqTOOjfZUvTq7PUL1seo3S3eprDBzMy0ayvwuHZLXEdEXk81tl4+Mun2Rm
s2GPVxnt5h56lE7MXO7/BGkCIHqXZpOsrmDcjzdPrsuFqhreM6yeg2NUJ0QjmNxNtRc1k+Ufx0qd
Of2bP16W5s5DTHP/0fniQk990NvdtM/HsYV7IQRf6SjENCb/tkuRER43DbBrW2yLHG2CK9PCk8p5
zPVCYsEDeTNWlfLPA55aKRutUjYX0oeqW2W0mB+o+UZ07kARIowEVUf0GpEHXZg+sKtiv1jfCfGh
nxn3z17q61nmRnGFeeZ1rzbQH8VzN0LxgNRdoAwQXuIC1dcUNtg39+tbvbTVklHxuNiEJhPvKlfM
O82zFI2CGn20w2PSUbLfGemVuC6DaCxdEDUvmpzLTpcMLJOB62e0cb+yEc9njB1r51J8Q40iJ3e7
llf5Cq5TMNczVYciQ+c0v2f3Yq15JtT9+AYFDkGh84PgmMx/0GLow7qlBS3Bwqp5mH/IB1hPV/WW
qYd4xBGDHcumnKUkbjQolUtkkxqKsIoJ0EuBmD5uS0MFUoi8d5wFgU5yLGcHzfG6FluJsckbdsKl
1No2E6GRFX+HtliSQ5fNpcMyY/VgQ+dfmNkPgYTQNuxBrWQgpi433j/+Fgt5qQgWrGlETCE5UYyo
EIhs/Asi6cIG0BHN5+h+gCywoLkWaAoSRy+Al+tq4QL6ymi7L6Ui01CZek8VAV/z1JJf54QyX01V
t1awO7tDfePRzUYYP08Sa4UXQbRpB7sVV4dbYoPxrHmm+gBOZooeJZEhAyQS3RsOG9kwQ7ePVuy1
Ht0IGdhzaa9hJ0r/H7hCysR1FRs0TZvsTGlgFE5IQZVNTBDzAeFRQ4VaxcMlf2/1ieJ+/4yopw7U
bKw5IAVCLf0kmCf9oGk6wlhYKSKEyCF6iCVzahGyPrO9m2f9rpTpM/oiy2B/qYpE2WvdE60eOSfm
/ZjJ5TukbmcHWBythC0xq9vwPp0CGrliC4ZTnj9k9RJw9x3xgNjrUL/YXK+yNtNKxyjHkc3Q98Em
IoS5k6cs6ZhbDpshEJS0ArKuIzX3xV0sxF6OMlLC2JwXU+01mszfk3YzjsjhKoeMBtke9mX5UjW3
4dL0PYfSkHXFJUfNRpz7ogyHe8zyYpo0f4mmXzVhzHF9rRxmLqnV+dy3vlD4Zv38lmawN5NBA0mT
aiTZEGlMh1lh8wEkEf/VXV4tjVrX39EnugV7mwoxdcFl1vBS+/eMVGmWCv15LqOnOc8itNQeiOLA
A17MUGWMmJ+iz2nwyIv+VPhxr9oMyCg5xL3bBKMBKbDC4pkjefFriBRrLVDnhAs0TkM8yS9Bwn+T
1mu5Z8yZQoYwkxJ1iETW4AZVs4oy40zuP2avCWqQbbSlEKXs7kp0nqpd5q8lYIL8Co0sqPCO/jex
xQRIIX0QUbGdCVHOWgq0/VgrH9BPh249lQ2CKwqfg1h8PM2pgd3bvrO1oQkN2QlLbeqTrTTCCNk/
94u1gRcMaloN2qt+VYsFigN4TVluIYY6atpn5jEjwrpcsRWNegLP0aSbYjA/wEYgcNubEGXVNNx+
69PuSp5xfmKhEilI/jyc7a1FWmhR8r4sYKetjZ2h1gAMfTEGpxL0GRgebqtfEKjr2zIQF2eKqyMC
gLkFPNvhHEWD7KXRu2TbdmNFXubZvD3QSmc2QrAsFzpHNKNNszfuBEsKSBQoNu3TPCy0SqoIgEAC
e0+lUs4E3gabfVI8gmTW8+rz57DXW2OHecF+nZJBj9xFRTCfYijredUz9fvhIez9kUV+FiCvsDF4
el4sks1Lf79GcwjMvM/p9N8l6LrhHd20S/p5AcSOugYjbwP0FZt6L11imxYSmwW59icO3o2EckYL
JS3R0kB/Ngndg0iazo7uUVR8I/OtQxiOvDPO+Nx2zsvZ85+p6AyoZR9AVOV7rxNl5tkLI0mmbtyt
BMIgYNnSWl4Sr8y2q2ttkJtUxoqafApy6H4a1usiMg0/JYzg9zCJq9NaY1zNVAp0TMEw5A/+7bJU
UFGc8iz/WURtOItshpId8bVOh+dBn22nOGdufZYbLhJSEFab4i184jEuTZv9B/k4anrp2UIe1L33
RtnPXWg82EQw6/RjoXyIWnPHtx3DIyhca5OPbzAqO8AQAGjt+P9Cnd5t8nnDASsRWLuJOxWE0MjJ
AKECrQyQscRyh7+UKtMPLaDmCpRZ3mvx+3oQyX9jYLQUNj3HBX+4dyQOWW9DRsY/ClTYchLjo7g+
lmZHls51SjzwIZOPuc4QIXTTz35A9ySNpOOjJfIKWB+PNWFnywhh/FDCU+teARa4RZmnDkaN3geY
LJa6VjcrqrHgH8z9/Tzt73Xw19CsDhw5VZYbHQx3EKV7FJP1Re9oWUuZ3M1Od7EE5IhJTmOeItCe
Znlk5p2hegupRq7tVwlASI5qY5tui8EhirbymgVp7rIeOJN004dOkQ/vtULgAXpi2AJfsdv07Lia
yp/Xa2kLXe6j28DORrE0+Cof+ZYVJgykpO/ALITlWIAUkDavdeKGuAPk9/AOdLDPf1M1U/NCVr51
A1Df43xhmRovabVEIMdmlaChWmrGTRGHg/ONdhMj0pl96p7xq86ZRspxeGny0MmYwJItz2HbiqqW
1OgFeou2e9+r+BQ8QIIlAb7hbs11/tdWkQvJY2BP/SpXpASKCcP0V8VcDrguXB/vRhalS3FMnmez
vvqVzRXBDiAvo1WaAdMDtV1Cho3IC+euJeXJGDJpBrPYU2jQvZRTYWbBbTUd+pDdUYF/YhhkU0Oj
5fGqvPv/j08CMkDgdWUSzFDdGSzjWxn4ndp2ica0fUQLgMtVC2mFLIrOSJ8yQ/OpaRhNy/zaKU3I
j53UAnIhNyCvDWbarRt1hjm73k48u1q06S/UAKCZuIf76cmRjwD9h0CVRQbKw5U8qTodYV9Hrf9I
JaAxZ+/oipokpSm2Z7kNRJq6HHvnwT0pw/7nFgJd1o7jcgIu8748q7Va5/1PU22wygEw6fzVouCZ
sTIXRTXpYhCG9Zp17SLPLa9ph4k40867GAVO/E4S6DK2QHPkY9iRytp4y0ErXpcnU9H3goSIBpc3
i+I2pOuhf1e439pKOX45jp9AQJ86GOzjgp5EutdUg2qMhDXRb68iGsBP1uakHh/wWIbnp+JIRnGO
Cl7tW4kRVc3Cw7fUiqYdU9DgoGG4RqoOxRGgGmGkPy0a+pkLfWjUkoI+rrCeUvCUifvIDz60Lla7
BHOpSoG1/FRfaRCV2U8N+/rmEkyyjI0ssgw2ofEI2kbtCVTUQDwXP7lhv3kXyXjfrQ0w3Ydu7q8Z
Hkmgu+WXn0l/VAXBLmgm2m3YTroE5aPEcQZxlcyHfNmyBgnHmSEHlg4q044zvlKR2ZSFEaCQ+XRk
k+rQv8Xg/4dDGaYrc01MM36IzxfIb1C2BziLraD88uPY7WVFW4TRfsnLaXZ8NuhLYLEgQB59lrCl
66eIhs1m+tp9K5oxakRv/rSanh+bY5D6REmQhu98yYS2o1VmAfDidThOd7EPo4VE6vE9O9GC3ahE
xYct9+2ALj9ayZF4L+OEPBQuxlLHyOrLIeIwU6+2sACRa1mdgOivsIAlsJG/8E0puEl6FRYBviHe
XOjcCLkhQLdwPCkoMBLS8ILWSg9oCavw6YoLEj63e2A7OrnszaeQZYSvQI5rsDsZRz5BDq5UZ0pI
9Q458DMwhdSBzC+qs8jq5vhcVKJiZXhTtfWLgM3kV0K8D+igTJ7oHJBNOpXKvc9qQYFR5XD4KU35
mJkxfVeRHh46WqTDc7sve6fGwRUp5lKyegIZuxxduttCFBSy2A/PFCl4d/rEYn/rDZPkuubHGpWR
xkCzOdGnlP3dTefn55a9Qiy7TvQ99HMvIAT8vZsNrH7/YOEUbYKSY+XpI0PPu8cHsyqj/AWv0DCe
qA0yupOLg2vNV92RVPESPFuruuXC5+t/MmGN52s+euQa4MjfC7S2C6qtSc4v++RSh59XEXXkL5qW
sQjNzO4iGiyPoy3n14oPwWLPJOXgGi2PXRvHLicC+edsr4mQlCTSytmR+CG+pT0YJJUkrecHwZR8
FnMJI3U2GaF1NOAVj3AfNDh7g7lX3o1gCwZh8keKhzLI6UWOSR8QXaiorpvRJCln/R9SQnbBZ4yR
OlJHqMFgEWunnEWAnodQO25C6CYTfSV9rAWNhkhUUZK5kV3ym3UCuSJ0pGeTFe8JwTZV0jkDgJ2N
IWb4pYsISHju9JLqXzbj8stHL/cPfpfsdsC4AJrgwyOhEON3wzw1fbkFFKgVzUxRq7dTrDwkyukK
M7qh26Eo18mR3Mugax194bAPMfFO88CFgWp440bg3wUvZoZFcExjUNkI6jAwY4Yae/3hGrSzp97Y
6cZdlTNErRqoQvpeFm6Cmwhhp+UKPF/wBkdXb7atMF0kOxaIxWuHhixb3Qj9f4fVdpL5UvKYHIOV
6GhS4Vo8pXOBCvlBrshZW6cIFn/2T5Tz+QPX6SzItv0N7iYToKn4vQAImIgIZ+4PURmyKiqregrK
Ph3Q3+98t+j39bzR9NzYyKtmnlXV+/2Nv7W3hdrVrpvdfYBBb5c0GSl1mDw8/e9fFh8+Oi8PntKM
AGafrHrkkoHIDFuIiJtlULOAE4mxBJKCEUYXlUaifuvzlthTVkBUAsDrEcqciA8Z+WboAajZRTB4
h4JsZk3Awoqr1YGpuuLu+qW979e4IRP9ULe8PrFQntGf4p8Ew4tdcCWPoIJ8abqRJtbjPDUlYD+/
4BrfwsbkxtvTAfRey737vX+T8DDvgKpwrg8MYCflw8lVVtby/NzMfiAPgPvw3jXztxGhx8Ji+lf3
nVlws5Bqnv3HkgCIdjPRV7GIYbfnL5snBjfcpM5lKQCzx0fiZkLZvqVgozS/QqvdUZMfOyi6F1U9
Fy3OACN5rXgjIsVFtGTvFqlVGB9IclcczI1ON4wk6tECnjZJFxoriLep9ufXOpmwKFaUP/8Pz2+3
i8FzjSrRXADWzimaQ4v0d7VOvkpc1sdt29RQQpYgq0IVO8VXWoOSHasySbB7NHVVfvWlFAwmycrr
wWgQZKb1EqXIYMSChab+JpFFIlxp2Ly2shxLpPskKhjKHrU4ytvS3CIy2cIpu5ZrRw2RIwqhK+Z3
7L7pFjOCKrlYUh2CM4esgF1H4X+9Fdm4ypQ4jWXweYRaQp+8XJoxh4uKXMbq3SQixOVeoUpM2GbL
3h8AOD/T/BctucpOFKo0ba4Gu/BQEfsQy6t2/T9NFxjai3LdMFWEf8NkbO6pHqhlLO34tIi0PvIB
PX9WKPzBFxSgoHUJet9I8JL0R16CTiR/poBwT5sD9w1Og12avsRaxyExQssWu0do+MQ1rGAPYmu6
PIxuMJOnOww7onJwEVaWRzRUnZ90vpkXbpPGzO14S0EIfDB+6LNdkeVyS7zd48f7QvMHlLeW/001
/FvsLjykV1o81BjuWNYqt6p3DZFnNQioNyDVhaNj3bp6742bTHLTLB7VYYGWuTkVv/4ZpHfnZfYZ
SsxudKWiJuO68cLIm8IR2eagLXlJlSF7wUciwL542WWBwuQAJTMuHTpAsPEWNM2A2kFp20iMCEGg
575OCB8LazctZ9AZnnW71qUnc4GaLJn2gFCsqGa/Pnr9oL3YMyevnZOx29uJ4mUUBDokHH8aPkaL
1PlMrs+zeVeJl1JdJjKibryk2pLICYWD16JVv2dGwIDMww8RJnMTA/gOU/cpfwJDMXBAgbFsE0/u
m73TJBc/3k5nyPQwKpyccELlc0nDrTS3kypm+gpSQLp1IV001agJnce8aliVUmCu1kX95RW/KeaS
DVrhPzqjGt6L+nDkr3YF18+MH4AzwCtOFO1FM/2dPexwkIQ04MzENTCz/ae5ztUapLO5nTNnAJ6B
kcb0zdqWrR1ydSL+65enLjhAzWC0IA7heeHxerJlMoWbJcaw/TOubK2nk1rfOSd7hiRmG9q+WFDv
HUIE5j6reFFKK3v67wQqY5aEGUwYWKySmkB69p8eghxuL2+jNo6pA6rz4a+ACrs85TV1pFh/C1Jn
65uIEzVYknkBqVcRO+fyO47N6JgFR+1/GIpV6yjBJ9LwMrK6L4T51e20m3Qvk2V2Z0h8PU4zH0OK
XVYVxOMCWGnYMYzAhw9pwuXpSrETOOwvWw4Qxzl2hVKAwjsHajScKe1X7YIDRLwJ5Fdi6PFZ8Epa
mhZOESgei+edJl3PpfUtXJ3Vae5cjgjMn2jIy8LERjWC9t1o55lOYXc/6D9Q5juR0pOWDGa9BYjf
ZEwmK/L9db3r6teFf5XaRTkyuiBjAs9BzJR2grAvdmaIzA020SJWVJzLHlkeXLn+KNi0bm+LQIBC
5c8n6K5PwhqJKQ6rocc4ZiiInXFEV5L1GF+NcQH1ZCBt+UaDdMAazQ9skkPyy6aUXKPLc5Gnlo0C
tjeOBw6riK+14AiRW0I3E3z3Bu3I1oFTnQd2DERTa+vQub7eyLstZfeyCXOFaq0fPRQe9v3IOTj1
QO7xZurzRzLn5yNQtv8hymUABt5x/YQu2ewFGWbm/yarGFcg8lPemuzZsJXjtp0HWEsAhACg7EZ2
JdfaZ5/OyP0AGEyObHTLSAylo5PR9eFLLx8Bvch2nvpHMZ9INSzv1aLLv9IFOuZbftLDNwsn3YPn
Uhw5FTr9MdDPQv92qEJwwKveb+CLUQWj4nOgk9Aw0nEJbi+GOajeptpRvqQNT6sD4hEWSkCuZOzw
2k0WmLMhdh6XKDDVR3vacLtSmYXE4i8ftq6sq+plLWxZ2ZheIiA2+cK+D9ACOBjkk4u4HINFFDoE
F3IgZz3vs/SfNz0ZD6AkQVWqgsfgsmcdH45ycYpOXUxXZd+wcTptYH6oFBEettf2RKP0Qya+3hMz
YJSnz+QyhtiIxaxxapk8pRF3ccGwRrhO/q5U4fQTXK11hg1I7ZrZ2kHutdZRhmVXPsvATOKStzhL
Zhl+hpa9fYUEk5E6I9lWVovHusSZn4JKeNGD428wrcWdhYGR7F06pfGnGl+WzPIb3974GGwJ3H+a
rwrY1D5ycLwnq6t8KkuT2OUdB4xK0ka6oAdFrPRmxZGATeGibjw0Qp1ii196joIbTklNLGD6EoRr
e+Z08bSKaI8Tklx9zXAPaT3QFV7DqjDNeaYfxnbq23nBiKOxNOs95vxz6dbgjtIYIpWe7t2bvVAP
lQhQQ4V8477HORNChvKtOuuAUM5VgIz9AX0nxYCQCKF0nnLurtPqSpXBbACLuhLXsN8FRF6ynidQ
9O0TUqkUqADFGenVHSfV43gJKMGRt2OzfoLgxQXgGlo5cFxmXyedUu8vfHzhZe9yzSh5/LlFycvE
ceR42nLFOB5eyHLseC8E6aaEhugp/HgSZQ7QVpC6M7tgBEc7smeK4gscBZRLxnhdJAXNSeLljz+h
5LbOsfieNAuXqrNRsj1eEHIJb/qdphxZhKtL+LNVz5VfTxFTYbkZ92sTAB9uyw5rwswIwTY9fnWO
U+0z185A7IVXpFYDRiZL2FuCcJUOyl53tze6l6dHWncpTP39WiwSsgtrTWHLYSLjBiIKWDi+fgZi
RarSOUw6Jmo16bljmfB574ANfWHh+OVsg05V7aE52CBoeBoqPqz6MZOWFxnCbjgA7Uf1VdtWoVFN
UHjGzqkTgMsYa/VFJxFT/SDxRyjQFNkbrZGvGpdISq3nC2t0IPdzDrnmvDXfErk03XyAqf119LWM
QU49BA7fSYJ44xrAR8XWGUrxQWNDXU4R8pS2HWScOZXrmdN5IsBpy8YkJT8UTlwR5eBeQcQL5460
bAovxMit8aigBJv2013RpXKe/qfQGHqs0yBi4IZtvzXjThNLkje6ikHXmGjZ2YKD1mzaV0V8JJ3d
4AeypjOte/opKVAzWYxml8U/lNIZO6Ht1x/6rQ2Pk/KcbVylKz4LWX0Efw1J3RCdfeQfwEYQiXbe
GapR0eEs6iwo1FGldMsqOdbZdQCxJ7SbQI6twsP1as3r+9dVhrPDGQJKA89AnDgKaZDxi/rpwNEQ
pDk9TPMWlulo/LA+8aEetBoVuC0S9rzx29KtB2N4k7wEUFWZfkA/TAvHLX/MhGj78qR5ELhaogKh
Yp64Mw8w87O6FpoMJB0Qgbk/E/v1vnu6xEbJI9BnFbfeEfVnrkHFkcu04jy9krfXDC1Bl1FfV/gi
QvUpfs7q/zqGtcSt8lkrKLBvKrrNwAGlPKj9T2eas+QjLU8PtDG5upqxms1kL6fIOTKagi6ruTEd
plsFQZsz9xWk10qAFkvD2GjTy78+LllP00o+SxESGuYYILtvlbIk/cM8a/+2wa7xnPXFvq1kYFBf
Zllaz5Vr6plaMAvkbuQ0leT/7KcfuZKaZ5g8JopDW8BCJiUow3bbf+3xOdqZ6jLwQ/n2YbMoPoHF
67T6M7Z8omqu73mu4F3PutY0BXDtt0uchjBQHg2mjmwJCnxDE3wN478gLYBlcvOqo1W2Exw46ZXk
K+v5ooVtamTKvMHXmjHDWQAHzcYR9Seup64jB9qwlMKRynY3CB/OpBWSXtK/c29Aue1M8Hxw7B89
quzwdtxgVG1+f2DpafrcXLYodirn+DAtV60/uXQNg/iUA36NDoEE5SBHgg4KFlkBIhocboF0cAwB
PILf8bWCcj1IO+x5BFBxvqA5Hj8S1VnA5pi6fJV4tysbJNcFwBPT2lYN7T9EKMGIOr4Ji6L9BekE
06eaMo8cPIAsjxT8/vxRYoQLuolfiIH8el4cs8VZW3p36KUzkhyOkp52NlAccIX5xD9P5lpR1c+b
FG7X1ySQLsMWIFE8HAj59GnysRGKFw+AYIYgrsxMEZ9MxtxPiFiP8AJXBwOS/hXIIr0v76TTGlQQ
wHm7DAmIe4YnQHCCkwuiTIRHw1t+nWiU1/hnALfC6doY78LlGnL8ZFbSCRdaZxGDy6WrXZWTR7ot
HZZ9HJya12yTuP9xMjhMnNMQKk6zC3JDi+vadkwbJnTg0ehaOLYoyyC+VMMTYuM7X5B0zV8P8s9R
g9WK1JCn+m3UAwbqTs/NMRSE68HO1YbMuiFYYNCBAJY1aHjkCchhiQN6Lu+mIJQfZK329GQUYxXf
NaGSuRs7PveF24iddUvXcUHJyAywmMr4WrToGtqnB03XPl33Qm4GTW5DkrlWaRfrwkMvTVYPQmBD
Pysl0bmuhfISHUEEpbcTYalt/vGpY96XL6UxqKLb8Hgm4IPDP273gIPorftHjf+3b40qFccyMgU+
P/BghKt36//ecEQgGe/0piFxqmZANuXps6lnuAx7cs0U9YD5VlG7CwXXr9bymYegcb2a2EvaW2ID
qLNwGqb1QDAzlEIupkUsHPMoeaTg7Ek97Bnk0yG4IgUDFFch5YZ4oEM/lRGgCRLvrZGMD9M0p/PB
EMW2UFLEynBfXt09fauy273c5372T7MT/F6tx5YayCvrttwyDOfEq7ZSA9L8UJQbGUHPZTW5+PzR
/Ahu5bj0FMx9WKMe4Wsb6Tt6G3j59SyPB3N8kfLdLLBT3WX2fCnYT/69MAasWXF+MZJffGbzTEXq
7b8CBo2g+SR7an+7TxcJcNaDBVJ7/Mj5n4X+skdnOtybjFWnd0AKXvyO9YJqa3QN2kaggpRjsEIs
CryGLwQuiJvmIA9mwPQs1PYeZgOVc2a8A+szIIol/r+eGa3eWxtyuy6bJnfyU+6yWK4VgAeXBGcn
2UcZGto1AURgcLsnSaRV/P8L4NvXFniNGQOMHZewScUme+qUa5FJOMr/aHTVHGKCCdneFJO1UQ28
MQlnLL4skcCy9OaqaYn/erx+Jd67s6sjfPEc14BKa7Vm0Wxnuk4fZK1lM9rNGiTowvvkieJWhZud
o81PMGyg2ZhPhk90WUKRVBU9PGk+evhY4S9l7SEMzbYMpEU+kjdLXp/w+sT2mDveuDCAxrge4UI5
D3SyDIcfsACjjerU9BsNxEXrvXZUFnzw1sYF2lPMji0Tsrfqb6YEGYarajSiSwWs/xtXM5BDRTCi
m0d7AY9D3MrJz5dbWrUTf28BgtIJzlWrfq8ta+mPv719wBRfQ/N003Hv+WxfvfxGvtP8Ln2eqnG8
U9CkeBSQMjif9w+ii3410It2XtfdNXWsykFbHNq0M88o7NE7Z02+w9YfrsrUG1nlG2sdbCKQKHfj
Q8Jz62lrrp7vruGkcdw5EanhPE6V/njfsg95jiyiI84MZGawY9awX66Hw+YNxHBnAD2dcz+GGzvW
5/qC8o7crSO5Kd4HUQ4lxCCqBKgBn0kksPNsziWLLlgRumHaq+/l/Kxk3SGl66TQ3rVfIA7w0EkE
zLmMLRmgX1D4qvUDmX8By1+ySgXqVV9v2gHdh3CSd1g7Bs9HxjtyKIJYLBqKsm1gy0uCJ1mK3loc
nxjPQTKcTNVffrYrX3RqhbT7O3Nx7iAZAWOps+HBEF7AhoO7noCMO17b+RxTlxbR363Od/R9yRGF
aKiMS6bwnTFO7f/7eYrKUJfD/kreDWzMI2Nfu1c5/CDXhXDoJ0nL2Z4ds8MNClyDm3m9neqgyfK2
rt5qtSrICyHd9iHiz/YVg3RehyY5GDtj9Qnlo7Ghvo0NkHdU8OQY5TOefMJ3h8gDUYBSKw+Vb0py
cofr68Q7rLAFp4EHNtV+uvybvEwRMnoZK1XthVMJlDqR+/+mWDErJZQmnWrkJ/8GE60TiB1ygMOE
5mo+vJ2VoMmoOgHdJUQPCzbUZoSY/fjRN+OaW7n5ofxcRdk6lOsnuKHZTyh47IELTg+YpXZFDpmT
bbAfozaseayyygRXSy64cMYGxqeUqwt5eiAblk3/oDlV+WX8oUEDQxXPzFISLi6ZBacZsmlxY9DM
rwzBlSXcjud38C9E6YitnaHhjUHoC4VxqC4KpVLx1+KkkrFTUg1RUa/DgPQHgWH4lK1aMfkpyRKw
Y53fFVlk7Z05zV7X2fHKq06IREcoweXjlK+nO9zepgFQtRyX0ndaOceQMme6sBkWApRwap7OMOgd
UbUHc0PyJLrNezyeSXsYx6BNIFyfh+tZ/hVIN8IDA6+pdF+16yAOriz7dv5GT0HDE9/QAFTV2GK9
PUS+IS0VstJBiiOKc3w7pSMf+aMeuXSTZS5MDIMolsD4dwvHxFXZu+Gx/EetJNahfbDQ6A1KYuh3
XP4swayZBfYfN0159fD64WlppPwYDZ2XEHJ88Iyt55sYwPB6OTZxrs4IUoHMk00osoi6yvz2Cwtb
qp25jfFpM+EYvmqw7f+pLeMKEXD8zSC1YazPyaiGIT+W+VSMZZxWAhLvQwFrWXYItdPtLMmpCtQK
GBrBX9mzcf8IWutN3y2htrVq/S+gPm6xT4ip5l35brAAsFoRCnsiUgoZzuAzKbJmLJKsRVUuW7fO
ecxBLi2TrjLqFjsDH7U3I4L/V3spPe0VaYFhU75gCFEXviu1tegCmnNb/7eW0RRintYQH+YfT7sh
7FAkDNzthij5iIWCfmtLcZS/g4dcuGcrGJ/GOh2nt2VijmXZLILQPR0cjTwVfO39fPb45UyKM3Wv
EbqtwcAEBBYSnR6u1Qa6hoIbtuHOJjckD57f+bu3zU04dw0HKt/DVZWyrCGTNJDXwpdLXiN817mi
4VPUaAGfcqdE/ZsJMs3CeckNEi4C9gn9yAN8836EsseIOR4QLMSZxQFdCN0UiTa/H+dzKldQocP+
65MqozUaEFEUrIap0pzbBBpMECcNx60Zqy7mIm/cSkYjw323PyHZjTKoNUD9jTJbNldGrQ4jwBKX
fliZbA1tgnP+0k4MfwNZdDHjUO1KTXx//Kr+B1XyeCOCOXcknQTPnYCYfXsFBL/xEQKZz5M+WxJz
bwqmC0QpONG36rj/9aT29VCc5keG3xO7Er8GOOm9yOx0abCi9gffDTfrCgvpPgADAFGvJK8ey2CM
mc1hv7RJzBS3mmN94PjpGtsZNY7YLLoSQ0WViTDRA9545iQ5ajX56q7lGkOVoqxmlo+FOn04wjcW
Fwk8HGwRkvgJeqIt/hECXA/4M/rDgEnHVpSuBuxNv9Q85GfZR46ENbnOWdiRbRJgE+kKVwfpZIex
8w8uhh/0RGJ3DGa2rVmbzrAzn1VrbTZ6Bd9qEcaK5tPsJAn7xQcdKBU+2ITwZTmaV9wR3iYQVT3C
ACxO+sDjzd31YaGAcGpALzUwT0eUPxuGEplTTpN0dqQZE3+ounS5hz7bYV9cLHqFspN8pVY8sXYN
FtBSqhALPJqlu1l2mfFaInjkvFfuWcC97nnqIq73YyUJPp/uGryBnzjhD/7yuQO25FqUkftn7E/o
dLZ7++T4AFiocMxWp9Q1z5yytDH9qcN8IWW7zWmWikXdnh65x91duNUVZS8GzSYA4cAoLBtOXP1T
UHDO3CmYk8ZywR3nn0R5jVyEbTLLQFRa92bHOi4wlmuw1Vtv+Dxv0/orfOomhexAlkH6KqMDqWe7
FyADijH+hUfbNi+XdPvnJ7uNe6/kGJzmm2FZCzYBqW2nakYPnB+2F/NfH7Qua96Dcz3OA/S9guOE
1a8W0K2Hs7nCgqGBzZX+yuQdxs9de2KXo6+4romFto+sNciB8dYpRqWJ6ZlNvYvBgn060o5torUq
ejYh0HYcgxLRM35hR3hbvv7wP6H+glIBEhuQ9KqNHCKoCPoqMm3wLiCb3fGSabq51KMiHuzBA1SL
t6M+3ShS5m3IiyCoxIXLCEu+TJoh0PglzN61l0BaiXOE9dQ+fS0MAH+x4zU1Mq5yyBF12lJJbyn0
r1OrHILiA7Z2h2gOIb7r8lu1MWGNWTWUf7ZdPT7JUIBKlljGr3rJPVUn2PB3gtD3gUO+CwZVpZdz
30r/Mk2VT6vm1m+ctzanZtCxNnB93Ok/mrzgGAiWXiu8WZmAJ/I2n3+2d+m9tXlK9DHIdGwO2sXs
+V2O5vrGq144xAERl2eDbjAHvR1Qw59gWgWFrP2Bck07lCfWDg/XDp88YkL1KYWdo+E06Mdp8wCZ
ONILP0BLv+lrwFTphuSpwNsfIvDBiw7qY2fO80CqplbHQCXPBjvSpopl3oxsrGfCUw3xHSt5MNMG
EmoyAgVDjlgK9zF/of8gSZ9bnP1/kXIaWJPsrWaQ5Jk487O2AhgLwWKSEatqi4Ea7q+SojhEdVDy
YVFqdVQ1aJsg6L/gS4JQq7B+0tSI485YSYuZlBrMlGapu16ObtfM1NOhx8k+AuUe5vqOZ9AdiHux
ZEXo3MC5DhvbqWrU5MHQJ9dKBg/bd4R7iApvPQo2zyzB5GeDqPTuN8d0fpcAJRsLCMp5xGAgvgfB
Jp9KdOXKWONcCT9upYbQCNeCMI/KfSSH0D3LKax6Z/tavAEI2jaXt4E+MoED51spLHo9FQ1REVrW
YzqeWRKAQH93i+B/HxBGzntcSrNKlK5R0+CeRUyj1OFygOjDH6CsQjFbeJueo1KIGBGPDOSw/pPk
hwiBmsKW/Ot8NRZG0q19V0K9oaede+K92FIcKNl/Jc5SkhAVSQSWNmiHNONI9bHJg2ztnhr7b1+v
BTJPpnUzOiOjJ/VPYvJyPquU9f3KjpSuDizmbN8H7suu1x2S/HQPfl2EgldQOAd7vNQgUFoZpoSV
TG4GasbfdVxBzZuqGpyKVDeHaWFJo4t8B8mXfBdlM/bqEn7AIFqs3lrhO1zfAS+2Dr5jPOUmZ517
k/Lx/3xA9oxSn99HgFytgX3kk7VpD4Lvp8SJK0vUopT/vpMFCKffCuR+elFk4lEqIt41Eg1vZFRA
3wrK3ADzbt9WWo7Zx5Kc7c+1rIaMtlryUD4azLS9+gfr3D6Yqf5gl+pynKy5bfAAesLKEBWSi5EW
062/R4ebJVsyeh/tYH9OM1RSxOSLcI3l/r/iDfSouaKF31oHbgReBXGlRnkeCNv8ukiQT2z9VoPa
3jsRE+JdfaWgKNljsNPLXEXpaRhQ7wbULsgAzZ0XoaiIunN2khCAouRf/xxM9MXtoLMoTFmDtZLN
1whniXjTrm85UnQDzzslqTOj5soC00q53Uq83zPxTmMRNv9r5mPHz+xPgQ18hgdHIvCgPOhaZ2y+
yjHdF11jyOG/Ow2PtOfvkHLHBowEkjp4fcP8c77RWNKkgcwGAWEdvHLEzhB/unUZgEEHwrUZriAf
UpH0ApA8LP2XHp35+ECfLcnS82hJCEJ6bQ1NLwLMZazA7Mov32d7ZTgqiCvJmPuiQYG21TAv83aJ
jXoiNblPDPh1bIQUHXIUuZnlNLo1Vfk2JntS7k2DrfvUnys4gpHnvaR61n4+GA0pWy9youncUrQi
pJLdt6HtC8IzfCodCXOYni7R4iJdRPrBByUD3FlHGZnMVcgZIBooX0RccbWEP9hChdoAxqrPdf0/
M40zhpXbOvPIf7gFquTO2EQGG/l/fnoVFV07ge96d2c9KLrLYK0zFPbVn9Js+0YWcjhby/nEeSEl
JXZvGesNEo3FGGWBmVevyMVnfui38NJwD3wakGOFE9QZ7mnouJe+4kuqKq0lBlJBxZ1dsWdC9tCu
/haP945sKtIWRLrqfQN5zf8tlfrGwYxbOgCJaTHwm/bbgHyAh/VkesFolBVUsJOiMdA2kIt8C97c
ZBoplHSI0//rW/BRlfMRTNLHlEu8iwmlt2BbfN4fp/DjzHGMg4jX+sm+JcdqhxQvETBI5STM87gn
XQBXLHnAjRAE/OI0YZ73LGTxmhaAm7OLnkRv9Y+Q3IrWaSyHGbAtnf5NFMNA6UuFNjH7vb0xLDEL
vnED++zyB8jfdLsRi2BC3xxxfOChhsdWiOea6wSRh1eqyFMVEhhReCipNKkBEluGJ29DQkAZtJni
j+GUY99XCNDPPprXvc1t4Qp6tBHEPDUowe8uiQ5oCDJbtUE0ziOhBxaG1j2SMmlYMTUiiwBkkQME
y01WE6FN0osMYzRmgOe5YdqcS+tI4rW7L0aDLFIsgJOod+2gvSbsimQOoICofTXAsmgiRKMlyX3m
Xasu2L/vlMUTc7NdI5V2vHZd0B6ZpP/7LMF60busXsr7lsS5cEgC/OaYW7iCbt6lg86+tBON08WR
MZeMRFcO4XfrTMneSrheYeFXbF6LBND9GajBbyu8umKsEpG0GGKDDTXNBh7aoIyll3xV6EiJiTlp
QrTePyCeSnaEEslzTxzsGgpscZdiNQakk9mQOnRj2RNfmzlMyGUvtn61tQ3n/XeQ5ZVog684hMBP
lUcAiN7w5ZUZfLIKNrL3Mew/han0w2HK90rsOOmuEjCyz/8ejC35gWW8xzoUiAoGOTwVs7l+/+0Z
p1ghKWOPEmx+fzXEej17823ab04ko6YBxgo/mlNMP/PTp/rmFOKtf+jSuFm6P5bpSUwPhPhEpcht
qnuWgIykTmejg7xFMZbO0LTroOnDcPBIuUdFuwjpwLiX8XFR9yHywSESfJzGhgUajD+qnlGhwYu6
kaKDDgcaBYGjJO0iKUn7wyklCm68nCH4ZwWpJ3nUUzUHAZ8AaeVf2YxywekLZfeU4+NvmKR3EwFS
GT0uAM2CHfnlHmhSu/nFE0j5Hqkz3Kz8FKdoEIZeKnV/y3uUVXZ0vFKMl3aojUxS8hAKzJbHaBQE
J03EC95WbRL9DPyU9YOm+d/i42HTKXM8CzexqU/hZOGJ/GUBnrZRvU01lc/tds4PNl43R19a2Z5e
wQacUCykxYdllAZvm+5oCz/rQn4idWYqhAP8unKBL2hToWxFvSNeTZkucG+/5303hPEldFz0+ELe
Qm/wdbxZ/QeSk5l2Ah3m/+B6RgWi8hEsZn8IZzbGLwSShTwPOVcoKjIVulJEu9NsIvhcCTOAmssX
FE8E6pgGZM3dT16USIQJ3TMwsAVJYcVn9+hV9G9Vk7p9Qkyfx/uaKkWR53RqleC3NhOhLfQ8YEe9
VGH0Ev612pnFhhJqcHxfUdjr/51zcHqBzE8TykJXPaOcUNVL6AWMdyx2wk/C+sNo+fA5goG5APSe
QKMWMqWGblJNk/SgFR2GO4HqgcMV2a82kP1STFJeLR/9UDfD7OkVZYzzekK1CqrrpccNpEec4GC7
4d3RFrVRVHjura7JrFxythZXugY2oJqEHZ/BGVTnxz4ysQc5udPVzuwgLJtKJ9iPqoOR+GvGMGgH
TUz4V/lmnew++RasaCj4GdW3+uuafag64ENhN6sBeLU0Bnug80i/yulRCeTC+pgCzPKIYJMXYf9t
jdzDMKbDi4mmw75qT4idRzcdp+7BCAk9vLOlc3Ufq+30iJhghLLdosBl9pXaWjU2cQ5KCfZOtg/3
aicrG03iGzRaJxveisIgTlFPRaJDGQE4xMq9DP2r2RvloWKiUBsmgTDNkyYDK8+0iwmjv8B2NHey
PMlkpt/O2shepm7RIhBHPLWGr/GjaS06mM9wUPJovvVi7sAp4BAjEnvYwt2Ehl882x2JMBn5vTh0
Az6X1JZ34unV8M7TzZvvd4fSEEE0YYpyxYucM1jZOIK7ceE3brSt5FBjtRkth07m80ZWH46jXYj1
mlyjzLijqK7VLpbEEt6ubqlVhBzi2nq9Zds5vWl3Ku+l1GZ9rU5pS6WmPNU5goyQRogg0qflzgtt
uBrgZ0TV7mCCKXEM7SPoWWQCwgGD5e+1RaAKA1HeFpuGx2IM97HlHJ1ueZVvyH9LDHW6ZwATGQ7B
VMc4VDLcyWwwyk8JqjC60Ff9YF1ceniJpdxL2tQse9R0LXn8kc0QbsonRudMnZdhqEDgelGbEW0O
xqLqidPK1Ts8XOSF98KO1KdBS7eP1uS24GivuzFyOL/pO2XxwVUlkLd7kD6qbA+YTR/pon7EWC5X
p2pmbZ8EzY7F0GYGQqh6VyNUleLaZL99wl7dyGHSVdgds0M7fMPfr+KvDmJGVX0YFNu0uDYTZ/l0
PWMBGw1IDs4W20FJvKq5G0ywioIyu1+yOMMbbndyzgnI/X2Rg+iGw8iJ1F5y+FcQ26Z84SZBKagD
bHMZzCMhp6/R1lvPwNNVi/3WCahWXcLAFEtTGQkOmvyZvtvVCR3daBzj//ONkBUQfZWNV0CCmFwQ
xzmmts/bM7rS5Go6Rr4K8hIfter+rQrstRrRVaeAvgHduZNe0ylb3IL1I7RFHiSAQnTHkyQZemfk
VUldpqxDcFRGG7jrNwEN+irx8AspvBEIC32Fi3aFplEzi4O9A1ZqJrO6GAybDLBZZ0yTMcc/sBgC
ETLNz+YIfrRKC9CeavSgOLrJQbK0KABKeHQUjYHMODGrx1Hg+0GgqvKDOtwoDDUQnDk+vjWhlfX5
yutS8u9daIvCWpkIxdmOM0hTPXiqvrloGdcyBwubdsWNN2NGIUEguQEX6TQ9y5k8fssNkGni4/dV
KAEN3jif7MsC3DriykkBX2Fg8cqAJ69CN1oKvQErb59UvVRrzU+/0/s1coc/AoGJR4qV+C6ZLuJH
5XdGDN6AMF/5Dcl5rdWPXwJ6iKexcJySKE6EuIxY3jwh270RBwKQgTPScjLxZkKBOZ8PTWEkJngE
MAmT5SoeUL0yidzx+JMcwl6PD3px9Zdfs+w5z6u8aeoT4zEprpwKxe5wBRWRch5ssIgIwtkA7d0c
h05HzeI8QdzH2XxN8DGDYuOcIA4nBPoipUgZr87n/uIijLZUI2hFplp08ADwNGjzqYo+RcoaNnjy
2VQ0UI/m4cy8yit8T0V6RkWGmBRSgVcHqfy7V0Tou3ApnxMtyeea4wuCBCJ4T6OS/2OGGfxGjKS4
6UgYSV9N+NZkaBE2F4hP2HFZjTJBwryjZiUeRwpl1jVi6leStT2lqW0cp+i5Np88Olm8oDPWd2ZM
5i9xQqWDe/esn5kL17zq+RDna0ZRgzw1a+IyuCytWHQJpcmsG1JV4ev5mrr2WtwGdTF1gWFIG+kW
tDJEO8qq0EK2d7x2nPJlKvu1nZ0WLzVTP3dQUdMXEdgDlobrH07NmnFuG9kBFLyrEgm0+Zt6cPAY
X8IRqI/oXfFWGmirGMn+Rme+cILAT0VTppq8VytgbYwXKkO9ovKrca2SptCdGm709+upWxh9dw9Z
7CQAaPX6EbD8K1f6Q+qz9tPQqCvHeCkWaaAYAd6uUHnNbIjaddP7RNLoBxNTUnlvwGw0xUFp8aTZ
sjhqZXROmuBM7I2rr7oCa9xLiNfLRDiD78N+zgd+lupHZrCQoGcDUpDuu/8HrqlR1abGB4iEkbog
vuY/jWStYEGGeLKETXC5Hy6ptpceeRM48WxdsKNKhP2QjHPi8jBmp9RFrLYzsWrEz9ez4spLbhx3
2uRlDzBVdE0O86XrIYbNm/NK6SORJwc1pRVxIjNgE16TEVFNKv634M/WtWroF1EKwGpFo54KsmHQ
48rRl/MM+JMoMcJWgxoEOnASISAbZ8+4InAohh4iaq+cDQpOxV2K7zcER7VOrFqQYhD1r1n0GmG9
SjAJG/tNImapAsvl2Qgghh65lMteg9EHAlcgVxcUTRj0FxOAL/N3zuhWJ2V6uyTfv0WLAqTikLlY
bLEn4Xp+OWIllKXt3gJWaBcyqNtMLzjZyru2002jT72B7xPgJehGTsNebsFjM8vsC20jkPvHNGcs
aKGvJYSmOXY5OcJ9V2YoK87sezwtnFV0SPJ/QtnSdX+ib50U0yfeqPyZo7rlkAa0lYvMfG+3s/5k
bKwOeeUdI00hWT06vSExXGSMt9RVUxGmffO0UjDHPgaZhVGcyV3QV4XKo1tRupyjSGq4ijAQsQau
gnIBuJms/y4ekw7mBrL+SkBvK6dOKdJDWxl2YvO05cTx+ucNT05xx12i93fI1HDdRVDIBr+NNKhq
OICds3/8ukKTMdA42GrrTQLE+aSCMICx9+wwz1QlXLsJpOpRqOn52y6rz9+k26TO6RVNVR62Ib5z
snwgHtqt4TXKXHE8OxFi+weevQUs3904QSCfnsKMxMHFx3xyhEw4RNiM3evtPvGE4u2iPWw+8aUv
Y7LFl9OwyFkxc22Nn0aXaWqytVma8Kge9u5M/XWouu/x8KNHoCorYBK6MX0RQeljK8K7cSGA/3Ys
7Imzhpibr7D/31h8vJn+d4p+6CO55Kz19JoBBAVbIUnYTTA2iIY9amJqOKE7wtt4atZRLCNRz7MR
YFIz0baCVijcwUHtAu2HIL+xfzn5o2BfHWoUHQzKRUqoMct3vSQyJlUSqIrTlAuHsZmgdFtFhPSx
3pWFka+AGqy7kFKOOUzJaZwbKTfG+qD9suvWDCW2+xm0HC7zhPUIpYd0rEbz2j6OTECzHbVy25i/
JkOZ98Xhd5Lm4kRDUM8TDIprA+EuGCbvJgLZP99yvsU3Lmqznz96pP54UlY9BEOTS8TPwxB/gG2d
EYKH8dUsiOoDzKBIyFH18eSVNZEgIU7nMc7ym7Kikba9sSz0gKdRH5ezW1hCVOiUkbkeqeRdxYBX
Yd6a2vxFKEnERGvg20v2hbFm9XVLBX3gLFH2/y1X/wXpJMRG48X+ha19FQhx/uaSOMlbHUMCrP9I
ZBrgqtbrz2OVpw54MXVRh5/kFfwtQzMg74I/Eiane3w6m0KDba+Z/zESrIptPwy4QwtQderTvcTz
AfBv/SS0lQp5XoiNmfmNSqOcIQMzQut3s1OOr8Y95qnDK7zf6tBhg4DDMaf1OFk9yC4k1Qx4bxpF
LC4nW0tIHqNA1LYPwLPUy/cLXuTLQKsb/j2RLDcT/iREnQTrhy/EfnDO/QQFtdAve2l4txUHq90W
zDlxtdoJmaoPwT9Fw8Dj40rbXxGHM7/0QWiLxyHX+UKutG3aFqw/K0PEazbD5MKvIrzD1lYotMwN
JDDTwfU6ppWjmRBPLOwN4uxXtNlfDjJCR77Nk1LIAMEphdVWiOHG4yptCvOblkF+cKqh5EizDTVY
q+dULSypAivfrY2ilmD93NgPwSpetWANOcc1/k1Q06BN0PEiAukY3EoCeLBk0nTM+THaGHjm6PO/
isfsZY2540cZTkacfr9PCQv1X4P2u6Moous11qaUtxyoUEECJBgnMYJ2xsPCEuQMFybSnZhCYBjy
UmPVv3l+oOnUUGMvztT0xMQYIqVNYHHwVtNiuvW1qnET9+dGVthFZh0UgplAWjdBqcmr3VxyqZK7
twq8RoxfJ3MghAYASbWeOGzS9LJttRP90ZrNdk9ui2b4NBvyiw93UBUoonlYwNPhKN77Ag+2lLf3
VfB2BrLrZikkwK1rZ6TgS6oksFXvfnfWucmi/56go0HkveLkJYzxYFg9WMRevUGl5HhfzHCcZGHA
uetDMJ5Lya+tyQF0TcJgYE26fyrX1vvCh6lGxlG8SZtUUapoy3dICdgST6oGApVHCh5j8zt1+8bE
y3E7eXYEVjRbp2b1QuiH0DEJu3iHo/fKAXPETDxx09kfdVYdRlvdQs/aulBMeSwlnPhAJD4TzJMH
mPfQnH0nDGBL5zn6Nl71yKKOiMDF5ulvww3AaTfLuShDcNl45l3bPQzZyZixL2iEUSpQc8Wyn3ln
Hjx/hPPrneAPCi50OTqlpoEHgkY+6Vodq98W9SKtNeEKUY9RNjvxXr6yA8ylBrEytZtQAQirsH+1
nFGWNO1geMzhbPqSCkPed6SwdqM19A1mb0aacCGQ2UfJxcNA7YtHQsAfPo3dnSVypH7WR7L8xQBf
yk16NFz259zx/i8cMtbU8akBSx9eFlgVXBcDWMT9HLz9IxUiAy6n5v4T/0Ya3rv23CCQyIxWCr5H
/ijk5U7M6cD8wC7q01+hpTp5sVdO11em73sUSalFBbaI14qTa8AOeqztfJZY8w9fv96vrlf47x8R
3xDFcELiDvMd9sgWqixorqWCtrDYr2+SsmPulYPbb1Ob+IxmxmhStigBr6xNDga0AAABMAX8H9qi
tMHGeEaP5p1KQ4qUxFEoxRfj2yrmQ3pRJwGCr2oGRysiXMPpWxELQj+JAdCAa50m+qk/ubAIZHs+
jVZ59c96We3l/A939N9/UclhT66n5ehI3MqxqOkrZc97u0PPYellmHdozQDZomDg4JQkSp3lA4HO
nvC/0TL+XtoBguKZvFNdXGGTQw9Osiqt/qH3RSblT/qoOUU7LsmLBmcHyRgr45wh398AH1xugSxt
2kBQUad0Va7faNJq46tfA/0ImArZsNNoxUoRWfTuTsqVaejTJWX9DMiewv1C3MxuivlJ0LHzg86P
gi+qXtm5wnK6UouBSxOdpX0hoJ9uvJOBjr7ptuDCQALuEO0I0RjeMQloCejg6PpAT9dEG3DFncp0
I2huc3fKCltDpeanEXuzOSL7QUPUN1D/YdzgAonSmJNFMXXgCFeHBam199aobmyCMCqozYsSAY3/
ba7drlDleS1vTt0b2eTbVNTiyhvwxpgJMwsQZrTTeUO7reOgoSn4CgmPNxt51ZNxD+usOa8wZErG
2yrjkP2OFKNHdRoMYu0YlNmZlccfyt/DtHJYC2z+Zq3YUe4v65aZR+80sSk+EnrW3W9jUn25CuNI
1CmNtS2ZsZ4i6+mGqLgoM1J/oCyyWLjBjHqdZBssJ8f1kRZn/BLLxveNqQ58GQqQqEL3lR/qgThv
EhAnADRQjFHwcQ/7uFkiku3EuumuCYwOPaUHKH1GdFJNXixWvJDrXbk7AwXlTYk23mW9rRxTaFi4
inOSPV3MIC7Hs1ZuFhe8o0SSJz5rF0Qeap1iabe02CHnT5Z+q5agJxx2LPF7+ND+xoDzqvA5l1RF
x1Gcb+W225vXsCdXhVj+W7opqOu8co8ZproeXoEitABarv7TN7Dq/LlgQsdqp/dOevyTPUf9lMg5
TSQnXwzSenJYEnS/DaPRz5/C5OUm2RxcMlyiuZaJP3zyoCsCaC6XRiKqSqYZSUa8qqO6IpdiFwSj
yAmpqvdEAYOgYyV6nTkuLtANoL0A0+V+xaSuJ4f4gh7Su0cx0/qejyc++Esj7Yyjyb+53HUVcSpV
FHmlFxbCRqm6eG/DIIFFFFBMZ5XmL7/xPuFNymVQbniU5eXirJrhdn7zx/dxpAlDoB1Mu4OdDWWn
Lt/LRxP9E2qP8iXY538w3yupeAJEkQyAm7cN0ecB67lB1d3YBaFAUWG/S9PoGl+urGN5//lI1HL5
l+bl/jwDaohPQanDY7QA1EMsArV4fi2ZYTTo+63YvQ/w7zHTfbjtJ389OKP87nOI1zN5J+82S7Qw
0lcAheTQ23/t+kjQqwkGqdZUTVD6elP6gmVxksD2fc4AvkvHYOFyqmpGRjL9Uyx/eV17m1CdWgWS
la6FofDQ6y6thra5Azn4BErghaxL8LKBQnkoxDqJyR8HTj8Y3DTRHF/sosP1YkCEdO3kj0D/dVfM
+LGHiDYgxNlk/GKhxFaKnYUhMn3ojxAX2u1GDRQ1Qd3Qp4qDzXFKknbCGs6ob3LpGEOQpYkyt5Y8
pyhj9qttGA24xE+tUC5ZbJqvaU4SU/xul+3NqE8ovYzrukQdnyOEpLUY471ioHJaQ32hQ304/Yh6
YPO3SVEmlxZwaIri+dkEXpVG8tSsKUjX2QXin1bUGm+mBaix41BNGQZhv4tjMDZHBFws9gyDJxI+
mbrhGld2raaHL74uUEGpFjjSCF2ysn/ojQADVcUlqFy2JaZVXOOK2jZrS3RKkNp5Ke72ZhnNDAhk
guvacoBLYtFdqwgy6tAuO+Q9paSm89KJX0XV9ysRR9ltJB6oSfNu+Ru1FhVazlrI/Cm2q8scsXmM
wr59mgGMQHJ8GoetiazUP7l3QxDuQiSn4d77L65H3ZvtmNN1dvhhBrc4oSPdvMiawdd8UvXHZpZh
6C7p7wK++8n2iv4iUP1jJ43pe9zastmJhGCox7Gt42Y0Vs8QXaiZHn/XtoIc7bvPvn871at0+jJh
2SAdrYP3Orfr6fds/9N+Kx+zkR44hN6GIyZc9Vqi13qaHURnyzrK1bcvTZAV07NuaZua4XQD8iju
ENcy1lqKeAJGZzqAwuceYaLt2mHw+vWaAqx4HgM5wotrblAGdwnrqR83AH7BsMokvQ57PujrPV5b
Ydhh3LMPkbrMNxS0Lpn9SRW4dY1V7k16cFFaI0u3g6O1aQDwvFskzQ7jLCm1KSTVGPVuAxK/lYKY
oeK7ROiEBT4giQFqOOsWZAX/0zeEy8Vfxo+LsWWaoPDK2O+ZgjQRQN88+g3/iewgWclY6clKkFCC
jbUbfxOPP2F79XkYzp2BcRvhGL3lUYmN1CBYJEFqOtd12S2XxIwlzW+9atUFeGSRmLPqeR5QmSwJ
N9DaajqWwFQmCtCbPuWaOBkLTBQhZ6k6itNqwV7hVYuMur1ckX3ix+HuKclrGdEXMKu8JGYc5bga
1r/6vV/nRdXqLLX/ithBcSbwAlERzdK54pilDNb1ptYcw4s06puWenMSsBEI+XvNA3tURPLih5mr
NFvytfvAs0oi6WWYpmBKJfXRaViDM165PnH1eLeBSSEXt0UI23yFaNEhaKsBufn4F4Q+DYvY4Is0
tItZNeTbe8alSLMq3TYT/lcASONcNQ4M+FaksubgGTxfqa02F/dfmPDPeylNaNXzGWrEpKIfC22k
see2OfqHByXmYtR9WeuLOdirg286RN7oVgz+0vMbk4mTsMQZYojkIMMUDfOs2nkosGr6oBlBp3r4
lZCXN2kgTXvUEE0Wk4YWbQ1vhqTgV4zM4YmQd5jL9ThHE8C35GEZOdDfixhIz0my49663vNhJACH
rzaF4+wNndrCP04cl1Avibhi0JzcIwIVDnb7CLMKKIIMjlgiruyJDt+8Wbf2MncNcMU6zBw1bB8j
gcxGHIPt6Ju25xNBBpzhj8yfkm0D6/aJz3z9RcvCr4pLe3Zjm2pip0YcMCaYDbgW1HTjot2jB1K2
QdH7Wp00vqvHcVe6iQfJdwg3vztugU4+C+ywnkwcDEHNa4FoYuOjozWOtg+DLe3ui7z6Pdb4cPIc
C/qUSvm8ANFJhvoTrgjavEFA837/Vq1WeX5jVHCtXVlf85WRMQB7h0YdSPVQb2qV+QLaLfXPM/08
9YL26aoXsyVLgcYWHtgMI2YXLDD/A1wWKJ1uR+KvVsQ0mSV9qp8ot6wvZx2u3Ihanh2KmS+W4jnN
cgPUtshXi4OmBXtr2pWAA6zZS1BGSSPh1y0Nz0q0BqbdfezHbgU7EQVGUaMahL+MWTE9rHoqIHfm
6hFW7SW4mHXysxqIZaNFELhZFB/IIoYDRc3IuJy/gjyI9g9/5erHNg1GSTDjxJgEs5MN3NW2guvy
pu8ybWsBt/t389r5eVAf9XqtjHY2C+ATG2WOziUVl6JqMwMNL0DGsb/vcTNIOfljsC3nIKickgnw
2jWe5ete+0FkLcAcum/JyzO6tWlRzK3SiCcSS61YlPppS1baxRdsKBHde1zIAcaBQvaujGfMZlkF
GSU+S2byE/f0+g18G9YxdlQGpnmqh5Shax9w3rFJkL6/A/9uHJV+Egz4411oUNcbVQ7FV2MsFVvL
3MXJMsjqvf3G/rBk9hCzqWwlXV0XwiNcDaAtSKWmaFU2IeOiFRaVIXEDWMhGPSQDwUG/n+Q37anr
i0x7yOa8LmL6ldZ7GiazcYr5/FbeyD96bJkHO6/KwJaC50HLTCE1qRMiJ0U6NPpVNYizZYbpqjOk
zPd+n3i0DM2fpnmhJlbGAIJn67njXiZDhtQkcDarKBZ1IY7VvbOlqLa/mkheOSv1b6UeYXzt8imK
bFeN8g+yWSJbTSC4xbOiGNbV5q/YVgenlTZPVDQlQfxIWuhahUPJhPKuyAOaTTTOQA5eCa6sMfy+
NrtBM0K7NBeRPOo0WOqnVsGqrlDfQ22KZPQJoVmh9XElQTTkTt8syPx2kbpVCHot83ZkSX92iQFh
nC584ls9q8IWKEGUOJWt/vrRL5nqXmYA5oB01eKXvGOVMrqOK6L8O5t35RSdOp8s7otqoQn4D+5D
OZG+48HUJUXT3j/3H9Sm4Dw83eUoIuXohh0cw2eJnUodea391xpBFIWxJroa2adNsxAwhv234Nmk
10JoIqV5Lsi8YbcfD/3lyZ6DwpQGldGca14SPPY7B6J15saIGgmM+U8ONZWswkQ73TbyRPFzsj2/
ILO5KCF7JBr6A34J4V9g352sENxxX7+Nvi4QEsBbGTh22E4qmEf3qK+8+GOHmuiBdqa0BVmL52oJ
ztdG4IOYb19gyX9qNvowZ+2OD/eoHXdvHVALB+f5GPpVofjTvKeLy9XOYxW8WPAo13G2cqJMeNd/
p8fyx9y746g1X7d4ig3C2bi9oePf7pUIctgGrXH5dC5yhpyB9Y34uDXkhekkmsL6UStsuP68aW1p
482oLrmTBQhf7H52VUwAQ9GQSH5kuaD8wFHhiT95aHpw6vdHGDQFT5nKIck/lPeXUY41e+hFrhi9
GQlh60dZuNSkaYJcWmPFKDMIpi+gV8/+lk4qanP8FPL3/ZMMLkoUQjkP/j4UtLhcka92olfVYexu
urJ2Xi2dC4dWOFR1Jvc3geGAcRDkF6tTVmNR3vEHdtZCO/13Chi5eEAXNT0TF58oezVveM9/N5e+
PN3SCtdExtVTdwJxMmxSKcWXjRXCyqEf5N/zsgHQIrjDRBB6jcukGHyAeubefmaOqYjFLqxyvF8T
vTPwH3LZRmimPTixyfMBQ6TDAErZAAOX6IaIqnV4S+wdjOasJZkzPlVgxl1rqjONsn8G4qru7Dng
DNmsXGYH7qBtMmZSNDPW0xq63Ojsx8a8Mqhka2D0qQJcg1pnfPbhIki+KktIpAJE57ss6AK6WYRu
MCkTOSV3G/4so5BgzT3hFYqO9jatE7Aba9mrxqQV6z6/s5caRHSWq3IICtVSVlEcGIXoZMlvQ/F/
WQ/IUh1BGNDM6+VU+3UzvA7E0h772a2AnC3XINqItiiXD1IdTUNESnArwvLXB4x6GChcdANoVqif
gDqLVrkCfvLGDVImNJT3GyRnoC02gH2RA+YVvIQJGrFzpNKkDuC/qZSZ1DGE6RRg2gtRyDeyk3p6
o0mkz5PE2EKrJq2RB9Tw/oxNIs0/mk6Ed10M6htNn9+UiVQMrEkRhz88k8NosfzMjG9v1H3i5hR9
i5wP1tKNtbkA7yZY0wQL6yJfvOCoUzasJv/2LCpfi3UwTWNyvbWRAECfj0zcwD1QSNQp6taVewVn
bLieI0il2qji2uu2B9tLej80iLwqAacOYjbZaoerHEa6CBsBFJQW8gcZCDTvjj2oThsOVc/wTmso
9wmtq7MbWMeTPkG1savLM4HqRCQQ2uqEbbDQOl2OOyCg/569QAIJ9TPF0PaDPjIgesXA47LXZ6Sk
K/ymtL2G/Xd+Dff+eHvL4czcdbmrdiTXVsVbp153gNInuBnCqm9Q7GyMi7idFPeOwqifB4sPDaaT
c3iZ1kRx9t9ieeD7LvZlSEOy3AHr8y6uXZJepbPwsIFHZzrD4dchpKSEoZVCgEm7pLqbqDhIN9Ar
1SrwIWf7gMOYATSe/1vzj44L2lm0o5LQyV4PtLwMAKUrosuU11bwrHPXZd3RhYr4snXZhXsZiA8s
0elhjeDjyVqXr1AeLZzCrcJ6u+lCFYhv/YjV6tB9BTCDyb7lSCihPQm2v9UgaBc7vdpTjq45b38j
2vDr3hiQ9v8l9fmLDZ208GQDr/kSiIUolaLPPOjENu1wnIyYuJMqZNWc7jbeZXBbm8hnDILnlkSB
tvVvlczOTBPw3rZfqSX7gfEK94RIcLBlPxzZJbtmR/J9Xv3DizB5Yihs/foHkae1+5/GVi3Lgm5i
aM8lMcerzyT68RV4Bnfs86PrtN34dVgAL2XJ/9qWSg7QKcPZ4wG8+garbfa620ZcDDt45p/W+VWN
DHcdabGZhAnXkoZk6yga24jkqZdfQFSO2/4MXvt3wYmuav2z8ABY2AHdznAgll0+r72+RPB93RJd
mFETUhK/1Ld/vbaCvBqnSk8ajyEcsoVyuLwBI3YipeQQ+FdCln9EEyXU2YJ+FRDrW2RUtXcRiwRS
EP17V34NWgd39FCVYVRkgmAPWG14hgxtc8ki9z3yocY1QbMJDEStUk0nQr99lTe1S5GlH2javfUz
31ArAaYcCb2UF/v3VYuzXxh8XgCqUHTxZb/PZ5SmI+5VDWgrp9QoE7Lt+IUFYJggIPQ7err5BBuu
jKYH1UYs2hUiUShoDcXNsJUNY+bfzlA5UZ37W5J4QyRu/6MB6+04dWsbwk8oa3DPk6fMrgdo3W8Y
/fvACPq2/gcqqiFml87Uh5Imb377RvDvgNFAHlkvT1KvEuhgeB+YhCWTlAzVzy8p2C5afU3PmURu
nghulfVs9GjUxiaRK8ycXMYnQp2xx7ouwxklYQ7AbexvcQWVbUJwbEFLB4cf6RQP8M8P/BuwncuM
OMvAnmCldSzzwJFJ6mOrfgkDTDu07oiz7+FE1tjSA8L3Tyzhm6eNXWZpu0smN84I1Ij7Plbkeobd
tmzrt+uLJs2zYqZWyMXVcNF6VyUr7/wmJ0nEnLOeojyZKYXYrHuvZNwloubP+8rm+NHsV3oFLlHF
EG2FoKZECcNfh/F/HbgERo5HPvRNmOpf/fd00vW2E2lLxX9z+4hBqT3x9Z5Trr300mmW28NERMl2
CXuTMU3S1BTszLugpB0rdEmPGh0eHME6R1gGs0a4cAuB3ZKEa/ENN58kQ92oow/fE1oxwET9jTMq
sOaHLsMXVj3NFAlUWF9jVUZVocPbYZv5bPWyfjYX6WSAjZ/kSb0I6duze6dectkx3g4C7ozjlkth
EKsMh/9QsWH9NLR6HPhjVOpv+Kxjceo63/Ge1cEYgwzXQco7oUslPCUoNt1ggNdZCxoQ33IbYbyL
R3diTtcnZ3zEJl1QveRCHSc46Tj8z3R/D7whrPBpKcGvryFxDkoqmgt/siqKKUbtzh7kVNI8LmKD
ClWHbru9h9rClW0amJiBp9ofuGuYBTmKFgeH0ZRp/eZkV7xpNQgCe4otwrUjXREv9HbBiw+QXmmn
Gzv6wA3Rsg9ZwaPDCveGVHb7pC5ac6aa/BmK/ZqrMFCvZECZ6AnwW+L2N/fbZ37bJ4C5Z4PP7yIw
+1A+EElsH5zOdyvjwkkh5qOSLg6wrpvtZF+xxypul0RrZe7DL8oUxIgniH167rrQrSKRr+UokIlw
zI89YUKmMYHJdHB3dz4mJi/9qwJMwCYGHRr2aARmUu48oqz0cjDGsCHovIEo9mk7jj4Mh7K/sX1f
mERatSOUiBSSf91xkX2E9ssCbOCydmN2ue64bJZ18GvmKTWviHnnG6wcjHx2dYuDhVfOIgYMHcLN
vZ/LuYcEc7pV4JAs57J8vkgDE80j0pYENWtn8U/mSEdH8pehkkb68t7I4eaT28k/beb1/i1lExWc
Wo5EYUYwN2c/uChiseTLX7UpTO3qfNhIgdPIIhASOKtcryTBA8/846kep+B3Yq10UeQ245Q+3qXd
AyKgQjmjukrP3RtBQKXLJqyZ6lTB06jUx5TxSJKxcX4kxjzlHChZAREyKAIj6ylCDGGOUzMAHQ3w
oh6UbTdamXx/2LUiHbZEPKEA9zX6g1XqClfz7O9BmyY5rWNsZVvMHu4trMP6sEFITvDyor7C+R2g
zTOBYlgWR6YCRQudNRmtnx6+ewniEqcKYDTStQne/8NBFoRl8tTbM9sOLGlLgXpdsV8WbQyE8Ga3
mPds/O6N0QtIiAXNwtB/gu5r55zHZ1j2ODcOdr3GE4O9dSssXDXG//u3bDYApjlSOsYwZxZsoFBf
Tyaz+V+U6RGVizzBJVeaX7Cp1JJAZYWArXlYzmriRCJGQjeaij8w+asj/zG1z/CyeuedRW0+K+F5
AKDd+nsUhpRzicVHGHmJ+s5CS37B3Tmn6BZC2N2LYu6aSPzOEz8d4gviG/STHJaaT5H3puJAx2MY
5HUOEOn971ggUpkoi6w+UvjScJ59H+5kubij5yHInSdqiKeVg33xU8i8LA+LL1TtQvwu3l44qxKv
rZ5l0YUiL7a9CmnIddkdQpdwh2nZgnQrf7ZNn45hnwm1Po05F3bXtHiS+11swvd+UIx77HXjwzO2
6KTocTaGkkuNr9ezvyuqKKDCLvEHcbq/8M+YoOfyQmvwBWsLQiqlAiZmj9HhGFatX8wPR7WVuzvn
jk+cnRTEwe1w42ge543tWevBCLzaOeua/aZdoxSU60CU1N5lmORedyOSnSUTtblHIZ0TiJmCKVQV
lF1sjo3zUqqoQltSHoa4cubzMjoGB8BdAYSGXsuSPvrYOqSCVAaVunTsnNpHqSGwSaiot1md1f1V
+VthpjlgZYEJhLoOhlMoxXTsoyGgm8v7biKDKi8/f4xdR7tRVaAdrhM/zW7QrCZOZLfX3VQIxlig
XZx5iiVa6lgIR9LQjwAzcVZ+2mBxUWsTpRxpI8hnkP0uEd72eUkDhmuhLKAb0D4HRITIgHE4uLgM
n3MjXHk2TAFV4O/Mf30csxC70vVIJmTUfwp/Sg3waPWFxTCP3hMO2Axzd8RaXGVonsas/+a3mpPT
tORs1aCpXbPm/9WMNHFUASGg+M18OlqGITUSGO7jdkGrtcc7GmCtcmolU1G/OX05DL0n04NPgUCd
r2B55jSoCqccyF5s/DGcwkUz+tLouiI8xAZZv5amSNnYuZO0qCRZ33JCr6UaUAq5rmzcMts43cQX
ruWzpFI+HXy/Ppww2JiMU+/wgtD8iw50rtxLnd4nBZJPWIVNcg8AA097OJcPQUtUTmuWb0MfF/a6
6ZbjKi6pFt9l9W9A1db1U4UpGBrrcxZnzl+Ne3F9YbuibgGOqRpv64XajfoXAVLA96A61VuWtwBT
nSvhROkhxQYa2jO6tEAb4I5NtnBtcyHTGM25ebd1AAeqIi1dwX1WhUUdKoCWOBDVi3nxadmc6qRn
8VvyFjEyMU7XU6Dy8cndPSognPGQCVQVgfxp0/6H5o1UJ9RuqO8RdWW0vwC+rtIeFmeVd2C3lGps
GiD1igm6dZWoWha+VmLz0FyCBwLRekC+UxZnSofHw5iDBQuFRquwl3uYZ7wAR6l7p90aOLJxKKpd
4VasP0XzScgxn7qAC6LatrTJeR+H9gKYe8UHEU1AURGeOad3uI/zHmsbPhhexdkEhMUZmhEPekwI
d6rfT1a7x30Mvr/kQaXlXhuo2Pex9ILC9KUaiwYB8wm+YVVq3iJByyXi3ayVabncEQ7avHXHbpCg
zUSrIQ00P9CxdCdczHAiKGXMJ739L77Av18UQa+uAxzDzWE9TyiY9GDSd0HJsoh06RZEwXIbiqFE
Tk6BefyQGfV+YWblv/F8iofIa370xvb21xklaUIPDmLrMGs2vLAnooIRziNhSLsIDC7naggA7vv6
GV8RzWzyfUqR/qFWSNVzVQbOESZIeo7YjSCL4kFCKh8PUmg+m9JHwvBG+N4oaxQOmTvF7ge0D0GH
Rn47Yu+2vqfIJKjq/PTiBn/BQyKb0P2f5/0Yo9HU1l67kWFMpaaUQk11H+0IEBC3sSXb4iD9vAT3
M9+UiskyHy7cM/99vccs+0ky1f46GSZToPL2tlUn4OutODIrVLwyb/tTha63T3M3USYqXsC9BGAK
HZKiQptdcGGHyqnuQ2k8ThYfRBruaRGjBvtvWsQgN5JWhmYv8+oqJcLeXCpfO2CyrcXAHf7ovGSx
u6HJtC/2GoxfzLiztmbQnw9F7R/bNqFubRp0+rzxwCQvsl6wG4ur3NtosrbAngVR74XxCTYREOjd
KmMbNT8QHSMgYifQJQmjfbNxKDqwtnE4rsOz8us75E18BzXsb/J9phB6YPQwAO9PKBA/QIcemW7r
73xTJOENmLrqHjZNaAw596e2P53tfOA1xR6QoxycYqkvQycy92buNr1i5efBIvNZW1zADhSYweo2
TvRfbQ5elW6UdEJBZ7fvF6T8ZZdw/anMOS8NS1LystE531LbPGxWTNGBuiMPWFtOQT4c7lDFQGih
Wpt0TbLliS0XAw0Vlr97/gZhtlBZQMbQa9kDX/qPQ376DFaKWFTue3Zu1QBorgJOOfQ9zaAKqPmD
X2LGgY07VmHEPWqUcxul3vS39YXEgvzjjsMqsFdf/okTmZhV2eGP97Y3jGzd/y2XedHB9hqTkQ6k
LsbVy+MMV72RBVOowC42M/RTxHt+JX7AiT1+Wy6t9CcrQheowIkAU3J82JfwcCygj7iLG/PyErfB
UMV1YKRMlrSUX68v4Bbw1OUuKJWjH8XnySAw/zsB7tRzR/AV6Hve4kYLeVg8mvjXl5vGq36cNR4w
fCQeG1Wu5MDAGLK6MNetlUFY2H//nfAD/RWwKhtEd8QuS8dptObgqBNowGf5zNxp4Meo0gSwFgAb
uSriCT03uWG5uyWaV27+aMQFmRg6rZQmhw06V/8n1nAki5UC7R0Zn2Mdi2nNsUmPMQZNJ8Pi77sV
bBpdOns8N1XVIyWJv6ATRx0IMOQmeP7njR6DAWeQrnzlXfxLHE5nfuozk/3WAC4HRB3CfR8zV+EU
DeczL5E1alTQ5sDIDmocpgsb14XpZX7E/8g57bVFIYj4KK73rQwO3WJ7IMS5rb+wc1013wcR6CVm
SmvPkwx3eFHJGyQoXGl+wson7vpZvLdNyNuEJpulgU7CPcHntgEr+8FgyjFikZeyeX4P6X6eds1Q
MJ9T0/REneiXB1q+47e01TFVHdg40Em+DEveroAQk3JYCm/BxLOATh4Ijf+kDt8bgw2dNtEgDd1f
LXbXT4QTDRYhATYxWJMc9Nm0729sH9OH5e5zYAL9saUwAhGFq9Bu1+SHKvVH6i6U5/nNIjccwHjP
7BqegR8LD0ucAFDB7FBDBRI4fIZw/8NPkV5nTuvMX4uvXtecuMy8Cn61+hMKw58UsZr+9OgiCr4r
5L2yxqDksZltmNBrTWACpX67fXhGUVWNc64hxU+5o0IGDF18D3QR3Q46GnuIhqhT6c8FRFhhq+wW
2ca17Gm1GZUTfH0CLl9IjpneIxf/9MAVH9DqSiK6u0g6tX6YAjazRjrvOqaao8sXzgFtJKnRlsnd
lTfnIDUi5P7kowk0WQ7RwMZarj19uWO3g6iMrJMvLMx3ij6GDtD8DYJ0IvzGpUTfW2mYx7J76Thq
IebdmoDteLV9EzhX9RpB4u8jp9mlV8lG69xScv7vu6CkeiYX27jhdmKcI/udFswtbkcqThMhTkgH
Ti/ai9Q+/nRZswX6HluPdLI6VIRUq67vhF0BqTi8hWvUgGSO4bzkcMkNl/WF4VWTd/uOxvCeN83/
3rSr58ILyCyIyY2/R7mkG0AiLun49hwirygefEVUoxNg32pTqsJ7HY3Xe3Y0KbE5AIiv98BwwjPo
C1p5PMrhx98sBiS9nkdLNm5gItnzJwJg0eQDpIBtdQpQoPWoZNc+vnjgvsO1iRy6AMGH305E2TGu
D06ICkN9NB/Bv8I3EzaUwX9ZwFGhSNDRlLTjuuH8+THdl0d2IaQ+1YzSjrwWBIEc1RDbP+SYhu20
3Z+gsZ1PmR/4vwRQSKEhZij+gtqS5BR3NpDhEP9+DNcPllXFZuzzaYcVyoRAulHVl6yPSK/K6hZL
2SatSRSnBtMVQ9V63pl2C586CQS3Mtyw/jsB0c2N78XO3WR09Ck4PSEGdGCAp+MRwv8UBholhcbt
VNiVaeV4Eoh/7KLc5tXGU79IrPI2Cw4tJFlZW5Ft0aq+nsnoV9UdCO8jR25xh9QXjNFmy2dQWGSx
XvSiKJxp2PGoFFUdhVbTnV/iRfvq7ZMTSRXu9kSUvYWU9Coa2fuJGJniSH45JEN8kw0RbpAPM+9V
GFLHh9iuV5gmQNkwL4aqpwigdpf0lxBL+331BEmiPyRUx020dhMwmWFeBn023Ts2yS6jjYiLq5nT
WcIZMbAlb7hMGwnqtV+8+O/GnozP7ki2EX5wkU/KIB6F1LvIssNlxrU+oVoxHivYES+/qhG/2EzS
aVmnOc9B0+NeTo2pZJbDu9uwE2JKF02i5gBYDzSs3vuYVoM7pJgL2XuOib+HUJU2QapUc6kXI3ca
j26doVz9iOChCJBgrN+aUx5rkVOOJmRZwuv4jAkGvqPS30agcwt0FHBF+DFyOmrGR+NRmXTaNEBY
LuLhHZdGg+ZMDQTkeT7kdQlJXI/yv21JDOBWZr0ZlAuwYaGiVFD2gl71uDNFYmjaqyHsL4L9LVhJ
r2PjsayXAlAYY9NdNrhNFkHN7WQooNurjVYX02+U7N2227adQsSdKDGTuUsaovFn+u9MoetSfpuh
7ZRBtrDDHDFkzF/Pee3QqDDsjzDYTdfNAdEXYhpy+ffw4tZIeNDiDRVvLHXY7MX2IABk+2EKlSbg
/Hd4C/MtSqn9R4zocp6HcJk/vyUUS+LvbjvCj15S48190o0mWsjOGvzquIH3m5le5La/E7X8rrzv
RFLm38XIg5GVxQDZrNLSmAzajNvVaiTGm5qnzcOBN9h2+/5GDQbBgvOrFjh96sEGeXbbhs6tJ8CK
od1GO2s83PD3ZfVyTNgmYssgd6AUGi9X3pViH2DVb32llWXRvt+0coXM+SrK6xdLqjBvBR8nEyI3
87mQ6GNg67yrVyIz/72ta9XwOprSWA2i4cmdYJxRe7Zqtr4BPkXUFDqInHSUrBdYCVH4sX37kBhV
v7w6Tj98GE90xPW6o3TSRixUWPXRFVZzcoJR2vsXbfVmg9Jj3lVexWIHHa/nsgVM+s00hM2NNrg5
iNCBazfdKxL0Ps1jtKAqMgeE7BaytT9EMoxuy+/ckWpte3Bm2EcAAtC7BerRFBkyKtkgXZU52upK
jpq2+5vBooj2n6ysVPI0sDLOXRJEqIK7a+Ns1p8kv9TvHQoWRkoZzGlBV+OO0WEWfyb26mroLXUy
poXxUUBswzKuLboAewpYAXfxIqtg1mQXd4yuaJZWj5oKIntuF8bN2qolKJ4avPZPBL8fChZIX2FC
T+mXAt9OAAwIdXI49W0573HLFGKNntA4AtD/nBqSFq8pf6VP8ksLQ2i2MRxVWpzEiAnxzSr+459o
w0UWM/+M18WBS9NYm4559OKVSC6bzkO7KTo2oMtdNMA+Qj5n5aUzYvtxFgFopaXareWA7odxKrVb
G097z8PGY7h+F4SyAEd3fVQghIxj/YnV2S52OejhLa+pcgGc3mxZbyy2G1bWKgi99rB3peHQsxpG
mPSX4SZWfZJGCzjTq7G5oDqCcLlwt3IA7edYT6Roate9uhouwUXIIF+aUxK3FfSd+pj8NgVF6YUG
4jS/p5JUGoNGLvQ3vKFBid5x+jtgJmXXAQxXFEcXyghk8A3I6AiH9iVcC5rvoKL0jHoWimUNJdVv
FWDnyEXF+/VnJngZ3uVHkOys6uxVrZVPWjSI2FfkX0cPFGDGeqvUlaXhMveW7Xs9apMDXCzGRNFU
sNg0klcTHKNY0Y0fWfkltn+VZJj/Id3OtKhliGopFqF2HaiKJlbjQcDnZ1wzwS2rl/1OOaC70z6l
rtVgr/zB0lfLTKNleMOHz0zKPWc+IJe7AkOEW2c7OtJ0S1i1NmUkJqxdvEX28oTd58BDJ49yNTqf
EcMGpm7+Xg+CNzj8XROrFB/pJ9N7WsPOhlnZLpIcSMY8S2gu1aWSPEsGhww94MvN4sJZjcZMXVZV
Lu03WeAhVehKnK3X8H3njnQaKLxG7iOvVxOjxXT/3lkgEpGpoYvIohGfB+wrA9WMnWf33Mq4S6+6
o93EBPB34IWXdNjM3TP77YqEskimhadEhLvgL6+Inc6mmKihyO4uIJwUr1bMT7K3TjTZQQAqDyUI
TGoRDhOPEdbGsGcUNM71uQOOAPCASP7bw+Mux9/fjOqJHK5+/qrO4tCUf1LF5tyMGO6cnRm3SbCq
WLpcjDhBwm5WESzQ5eV3XoYiHpKkVsm8B3utJ5ebNHC2BeQQOhfBM41xUqKBoL8qOF4H0UHCK2Tp
lRZnZ/CyXxP3xx04BXE7Xy3TOzEwkFWu3uQxPUFnMVekHR4yNnSRGh2R9dBR4MX9gTnlgSo7tQqp
Y6VMJkMgox3MC0hM9ezfb6wwD2XdbLPA4LLZ3voENb5Ft72bhZ80Mpi+fJQDLYcv+Lqfo9a5zrtz
a/FfQh6lm+WAwWTli1jWp1gOnyv6E5asVJ43f54/UIo4BdAU9mDORhO0/7UpBulSmcrzTpyy4quF
ag9LzCmYPW8R8kX1/je4SCkJdNOyIwjIZJJP1MYWS/hoLfbSB4j1oWFb6bRA3qqbV97KigXtcu/v
9Tc8W7ICJdduEW1gDOKbX4iiyBiEswozYF+wKwzVRapb0sqsK76B+1prs77/pd6D1lBOMoiF9grv
hxHWqzuzebZyJfGHWX5RZd+PcGO/s1OrwCszGI4V0HwttCEvwo13XIg4/VhzpyuVC6LhjWk34Nyb
d0MlXeDSe9fAM/TKpoz7V4xcADiQqC1QSALWgSTspCFX2pXi+d8Jjiv/SZLQ8+/l3LmF8hOQb515
DheODcD6ZKp3/FOB27yD8xvQpAnwxCZFgrakomKaxym20prW5AS17LCn/AHewY1FT16PYk+VmFCq
5xWvKLhj9/EHDZQBeSdTDzrRfZ8ReiqW2/Xt9+v8FUuiQbrQK3uDmjGlfLxKkWvGaJ9jXzvZfrrd
EMo2M/PutkaNCFknUowRaQxLCWQKdFsGrOVbtcY90RPSfES1yM90OujUIYVbcZndSpKRgyJim0E1
HoJ+mj2/aSzKhp4dFiBWdMBm9JuyIHnogDvDobyQ/rLen7XGohoh8vP/pwJGHWtfEKqC9ATJ+zaW
KpKdNAfoWFTx7JrWJnYuC/I351S5/oP45oMNN9ij1xjCAQdJdoJaeQZXC79b3lu9kwD4rgSXChiH
KLXwQPq5WokEIFvfwRu2cqPSXF2onAHRSzIoi9gQuSZ5PIZqUbX1/+kBa9bWip6vhukHyiw1u/5l
Idz4wY1VgJFKdBafXzeHMQ6Vo8NIqSUmSvoKzi9zoMmRD6KclW6sig0abPl3FW4TAOTVtwR5U/gg
KlxHmxqrcZjPRGtk/MqxOgewGVOiG4UR84TexlDIM1tV4mxdLSVpcjNCGLvey0NNZCwaBhPeqVc6
xaXfJpeLRYEI5G2xoAA37y6yNwKFlwzo3jard/LnojVpEUUbAnK6MrUqTEZmnQtUOxoDqKejV8yt
qJnSIZTdBRjGctpcw7DXxh7hSpCuAkfBxdIO1MpuhRUszbOCgNOK6cH92pcaTaNzA+2sz60P0PEg
ROfDHWmOkL0AuwYu6xWQdvseLh3XR+lwtlgAheHa7maFFVvR8Y1Sy8hP8T85gi1RfxA7rY2k8TNe
FTnEzyFe/m38VJAISeVT24uJ/icLitko27Jdbh5e/cWv+RqHizK1SCXOdsQV7P9WqvLG7TniUQwp
qPV4pwa3kzrRvJ5pPKRkKCBsEemXgHkTyZc/41VU7vbgtBu3TFcwIYlYTjdCdbt4HmWIyoP+TAHY
emUmWsUryCZO1o5okEDXHpo1pYKf+KKpkVDSTb7Cb1t3bD0Wh9e0jjYdh66CnKx4WNq4Jqk4ckQ/
7XBDEDm3t3c+0hKwBGV4ZiYKCxyjXr34wJdPHXn5bB6hpRutX20S7i8baUAOCUy+fJRKKrdlo8rI
sC1oEneVuSuUQtp7orO6wq+HwP3PB7dUCc6ycH4r4Jkz11+xrcemR5uuoIBaKS8gn9OZ4qI5xEr7
zQFVJahScCMLK8SLzigz1MouJfpMTW3YOpXwZ6BL7ZckSpdRTLEY6GM1z/YSP1D3TgO4alpxgW6I
1o3sHRWcx2szRaNHIxlqkUI4vN1XlRecDRNRK1OA2kemt4U4XfIL+TO31cqlWKH6O2RwxICyqQXm
OF2z7MJ46lrzfHyHiXvMm11BRHT1XY1olBmJkRXMj334oQXirJuiQtUyO8q96gNU5uaDXF/ueBvC
H36Wf0MTaM4EQCzpYa5yM2VE3VsmkN2dIB/xXi8inQFXD7+VBTEkXRptJoyPjOW297g7XWjE5JMT
sUGlNOFF3cU+Y5/zZzjrrZlZgwYdiZVpcwR5ueHLN21pcUiIBO6T7p5bA7IRkf5SECornga7GRrL
mnFg7djdCuJfZZoq1noDvyPTKQWgWSyTe4NHLYNWsdbwDwvYMb3amkX73P9i/Yvi+Nr7H5h3wMkC
a3oIUGp5WP4Dw0rUBbNtyIuE297fB1wF/9BAeK9StJynlBek3+o7cS5B8q+eUBnkQ9NBBMjQ9+Wh
gt07IJ3L3ualVm0dsYxXtDIdsT+6wGOGRI5jQYhn8GRamK/BSFKYg7MRwYsAdW0A5sVEiGbS3yxA
36+igqRaabFpGLNLXtGuqmgltxDIiVCu22g1Fmm/lSN7pdwieyVulGr3pjlAbEJiS2i3eys35OJr
DX78bM0slYDuN6+GOntKlo87xqJYZrDBz11q9tfwspxUqrX0vGFbYdJqbmPH1S5uP80TlLwR5/Fk
3ETh+yU7vRScX9Wm/8hEC53fqchIn9YKAlHAK/fYwXk9ifB15vnTZfBCRhwjOoQ3qhf1mmd5Lsba
Ol9YrCW/LsDvT230HfHl85qtRNdUP7jUtB9sGNCNgtnAG9kEdt8nm/5B9oxFXCiGb0SsSEbxpaUn
Sv7vDvWc60Rf4HNEDOkC8kHzzn+Ur2yYfzu1wNS3Rxd54BYf9QCJ8o/slzHS7/s4p/RSMYARf79w
GdbKn8HN5RKUxLzjSa/XSBZgpP8DUJpKAwU9xmH3BKlTMgRVbkOVdaSWp27nAQcKXxNVl1wHUrYQ
CqBDHo3/ooIkOAmbsim7cjsiOviCWBrLAEWs7qOSiOQlLxtx6tqtHOJDuoqHs2W/HqP4aP6d1ELO
L7HniLrepMjgSFu4bQXi973O6Vvvkjd/pC+wqEeRDm4HMe12qIBcuTPfwpaDTGc2Hb8CwPtpjL0v
vc0FkgJp0Cr2N7mJnuKzaizhzRfNfMuVgzyyCHps7eHk4PaBXYhHlBk7FouCyhhWAAUa1BM2CcWC
ekM2V3Hm4Nu7BvdVd6vNAkh6GkzfQiOrnlNAkMxIToYWWP7sXj8dSUrjA6ljGVTIppUPLc6bYqwA
eN8oZMwhB4EvwvM7HT1wQxAp/5buYQ6X7NKIAbWPAGX6FDYPxWkLazSzNVpR9uoKLB+LyQrb6xEm
C4/85NGzp0qaiguGKAYYepzN1DCFI4fhGvsEHi/B4TJ8FWFdspYJVr5e/lfJ41rVExDuRPhZ+Owx
S5ijXgzQNKqBPx7yLqOfXwtsSA7hhBVjUHhkh3xZCUsHQkgCWoLA8cvwQ0xJRcyesU2a+19B/LOp
UCHFVaARL39JAx80/iaTFuEtJdCMZ8bhhMKxUYHvkvu7oH75OTmver5gOtbHOkaSDr45DmZYLgx3
gJQMRtsCBCJi3+5rGp2Rfb0obzm4VJRUeymTRCGVcY+vZZOfaElLFjM5NEyudivr50RIC4b85x9A
1hLTyzNgjR9MLAgPhywLqfOIlgahHQoXhPv7c/OP5Pas1OjCHXHITtXPfIfgKdTh2wP0tcaaAeoL
zn5LUgc9p/p+rsEWznFakaL76AYqORM7qJdxs/dQnzk209mSq25M5BCFyWbWxwKwe3uFOzZLTpy4
Ds0eV5EXDtJeBG5NUnLkGz/5iMmC6R53mxOueqasHmnPimin87jnUY2zC+D5eEJZc+BMLw19tqy6
abbQR8vrx+S0gii8Di4aCdafEm5wG9xyOLtLjZX81dqSqLEn04OwWQTYzh9TY8euYHnZH54mS5ox
CzVPPmxRAaXh8LKAjJiv1c1WUyTXHnGb1kSjDr7QExEr+tnWeTyL2oRLN92X4usJ+LK12oE6tAxA
C7A9uqB3f0XW3fgeEqq6WuNp2xBkNWcmO4jBbdF6ysirbZZUc7denxKSwKH6r3h1+BnzrTj/VJ60
t2hv6n213ZIo5v95fiDz8fqKcmxFg42zG0KYtDif7PTgSZgSPesamd6w5pEIdf+4MLrxWNffBZbN
Vo9D7b9yt/9ncRoPdmtqdk88ijYVj1G0bVTulxENLm0RSG6rv93ez3m6e0IwmymecKU1Cy7c+tL6
70BJs1tgj6IsA1O2XaeTkCFEQnuxG1dZqHZwwAvx5UzcdTSTAeZO3be+qfeEM7+uD2l1aWAuWzOl
65nhtnqAugKt8bpLhtrwtTarZVNUi3kbmKUrQF/9asYY51Y0rBKCHc98DCr6xOJUgwKuSrh4aJGe
1uB0dCo6MX+Di2lhL6EYinOz+FKRi9fDdnVZJCEo3bzU0KNrP1VPf+DxzypyHcv/s2GUbOARMDvJ
/SEVVZVqjrRBdGFAN2oAK3Nr13/zmdTbFuo8CM070SreFf60dBxyXHOBe/2LW27Z+Kez2+heKSJ7
OySQmmNAIAwbR4H+9T1V64CP8FA4wsbtXDcERrr6LT5nYEt/9UPGz7o5gwtHkOPXXoLrsb5eXrbU
gsYGE3jYN6PexV8Ym8OamoLv45ZVFl///BX6yqPoqj4EODnQz8kPnrYYgboThocLvi7xrF7JTiaM
C5soWqgwCR6/dJNftBLR43QK1hljb4BMeocgB4NpdYehgLFnrMc26YBTZVfJ/4RuNojDdpzsuDLd
LNUCEDOeuLAUyNGD/cAMsqf0w+DnSTVba5VfjqYi/6uu1SGk2fMXXhzqx6cXSRDHCOtJVfn5EYmT
aiWyOmm2XSIBNqyxW5lANSur1Qy8caW5d2436WVq6pMCwyOGeGOsMq33MRZPALp6+Wta08iJGFQc
tF8x7i6KsSMZA0UHTGBFXvI8/5ssB785Ixy2N7iOd7qJAm6WRutkVGBYvM8ahlDn4chXpQM9EOda
vc8lXQG28w+049vKZVSYxSlRN45a0MuvHAeAMmfaKyIo+Yqn230LSmiSi9WlOua42alD/9Jgs6lC
4Hx25vAn2Hd2B7oh5jahzNggkw9iHNJkZwsnVKW1z9pT7FpXa9/ysldXAg1kbvfIsNrjsx9fmGkr
rHx1opFPdlg/S6p6HHl93HYinPiPdifQ2i7qTU35vBevXouw2ES1ZqopFKVfnlBevFaIwOjVs01H
7O/hecBCL1WjIr2JihXS9Pm1WQaUMuirk4M4+cbmvoYzWlfqcczmkXxL7N8u4C6VpSipWBL2bVQI
2gZbgo3+OBrR2DVodh4TP4m9rtZJs8EtBwG4VnGwVPrXtC808O1zNcgvHMYbMwN5jddxABg9Iz2X
0wgUR5T/ZsTkupdD4sFK+zAQQqHhQ5CAWGpi/g67uzhBQt36zRZT7Z12CsoG2qkL98bjn0JckAq2
w3EA9rzfAN2Tm3y04uc53rL1YlXNuzLutuFTOvFxOwkgIM/sIfjeI93LjW+lSIY9e8mGMcDKtxyb
wbPiUrhkCLVdv3em1lpCzuneKOr67SaswYrPnc2EHT7dxWfLXrsOWcpIimRRJcgi2YHhZJBU9scU
dHZlxn98bssEW7Pnpj9DRcBrOJlIkUsSnDS/OYPdMJ1CoE7UI5dxNjlrplaRgzGGsLiaYbSDBbUs
UdwI8MEMX4Q4pQsgoBBohSaE2MDXwAtZ3TkDLnJ4dFRV5sYNaR1vr1b49sBfE9RXPjhJOp0hSfUq
KkyaUab9ATyzmwLSyrcP7lm/ec0YPs1BFNTBvofkdY4qe6m9pjOMM9kMSLByhyNtBAApMIMlN1F2
h5gVGB78nmBx8uf8ElNhOrK/vhwqwLuI299g0c7rznFqzI8qttkGBYgTue2AHfcybs0JMsqUYsWc
pHktKdCRAyol8gMtqiioNNld1vLJYZfFrkAdv/c1adlDK7BzTlqil1l0mKcjotRS3Vm/UAVzJID3
P3zt/ZctN9i4/NMb2ULJ6QltQ3bzz/ulenTAzRUuWE13fwWvlSvniscUvTi75JsswbsvbkvUUwS5
62QbbWijPHA9hJ00DpApyVPUJJjpE18sOTsBkhoczWoHZ71tSHrOuXVEuOET9UOYiN+Wogw6Xw+V
vfYrGSMUzWUy+75knJPxkYDGxBYQBZ7NsOkAUHzEHafoy17yQI9BXgLr1zi89J/HWswuFl4W94Fn
9HHDKZ1pDauV1J1qmLoOpKGJc//qdG4MX97RzK8Wy6c5vh2S8DSVKfkpOpBEr5ha+q93bPDx/IZW
SKFnxs7sBJFfCC4NkobIiaYpqh9jb19MSF6RXSDw1zs0/6dQotDCSrdLXYXOmt+f3DKyidaPoGuV
66/872Ry/tRfaQCh8F/0N64PfzfLfKSJIjXZjBQPbshUiBSq1A81BR9ClXAHYN+2NsIR5OI0Pikq
6frTjlUDFJz9zBO+LH1h6IpqFIoUyBFJbRK1HR3z70g+MSXiVWoKlvArsZK1I1dodk5O3tTN3qZM
W1az1uImMxy1ommZa9riOdfJTK4GXTfi9n/m5j+l0+c9J4aAcQ4acgjQb37U/UHbhDBglUho4CP5
+goIKLWvRV7ENw++Lu3ig2/ss+g607BegG5JBzHWW0HDkwLeOBSMfdrXaSToeFeZWSUdsXfKd38z
kSritVtjpRP5F8zt+ZxNEVabF9i2G0bDZazNRHjbrXrcYqKQqDD1sTra682qy9vwcMUEdqS/eYTx
msLuz5I+sV04588KzazCstvDe/V2R1ATO6ACn6o/GcihSrNW/Fv+SnIlNqowhy3nK9gwCj/Hofar
RjtvCKU3s1oEbQNIrkNt+jwCt/BFfpZch4m7rKrAaUVTo1xY/dHpdK8ExnwH7JG2QwVAobbAzhXC
v7kZhhPk+Pvkkj4GroHdVcO/40MQyllz9DP9YXFvNCxPJzREDOAJ3uE+byP3QMLJnr0t8+g9ehRj
pCUwQxxubjxIxhs0otf1PwxXUSm79SRc81AW1100vLBsszQni2jrWdxArxDJNNllE19friq+Q31x
s9BOowt3kMmr8km6g7oULBHo5RtTfg6gGWTfiL/j3b/AswNihgeh0dtmxmxgdmx2WA+VdbrW00lI
rRfW7Upjwl/4X0WKziXABtoquNueqvusMLpwfod+l7vThpHcQZnQ3exh9/zvwxLX83WCKmDyUjPs
rTVEAd3uQa63KOX0z1qTpSBpG6Pxlz1I5KyDjBcGsMMecYlgQQqZ4wlGnXSuQeKyTzvjmJsTIAPz
YyC+Ssp8v5G3hSdJfxK9zDXsTjQaUvC0HSjCH2IN8Kh033CmrAaJmCduJs7SiglxHAY97WXpS0jb
LqHFdRLwDLcOozhowZfGOoVQP2wRwUK/9XWPHo/JpnRIx/5a9vfnSDkzCStEp5DdcEl2tvB0Sows
GVum3K5vitB8wItvkOIbQOgcHOYEbv/T8BxrqLtUqEMkJjhMs73rV+Ss/eV82LbAeyCtzm8AKpEQ
rvu84PRP80YIbr84l6azNRd11U2/4r7nR4jljTjSnnVL9hlDWjqR7vWj3dBksuKWc4E8hvOgTTdL
0RU1oXhjcAaf0wzdnBKBfP9C3ixeM3o9sUKgaYxobotfALQNGUs8Ig2MDAC83Q82ItWXpOaLt2k0
Vu1vPQWeZH5JfooONE0acq6QbOZOeSK6+3leUnmyBhiNkz6DYa4dwXGDVJKQDujyptvZD43fqgYH
PNK506TOlNlPxaf3UdGZI4121wULyGNEOeEM7XDTmJzfD+GryyAQmq6KHxvbP+WxzLRkOQWLyaua
AGvZtF17FI1clNSWbXuzZtMvLhbnXb9Dag8rODWydl8rT1oqIbE9e6najbdM5LW41dzwr9Ml9D53
vl6AKzLpGtXJJjT6j2GtV6xqb0+7wdkQq3DE7AP9Ch5938Eh1/WJifG7qAsAJVItENQtebqqJC4k
xTorVgN/rNuwMK6lL29yKszP0xgEAZkKmmriLYzfWFO8i60qDWXcNhH65CXy0XOAquko5ciIp9AJ
C5pJQVYHO6mSPePlAZm4TZcQrfgKDRm6Zb+ADbECzHygmiqTODSGQXm2BkWIio/nykKsGiSJdQ2B
9m8hwxGrT5i1Jv7qBzmHT5OFjsfrLByB3VSwtm7Sj0cWyzMyjw6XbKBl9R2fbhZrYHANNrlS0RKo
n/gkdx0STvL8uT3rVrYrn6+JdB+zJigX28y4wl3niLJbbBsD6SYlbfs5MAM2aZ4PEZkLYCk7Z8im
rXRU7COeZSwBb6b7zblya6eiNFZSoSNM+J99Rn1Y4SK1GOfMO7EzC2Pf4oWUvZAB89z/Apt9SwRQ
jgs3dETqILG62kT586edoLcZP+vesSFwwqfZTiHREBRfHmReqYwhP7z5HVWj2mbWR3vt6oCKtC9L
7SZfARoNTrpGucmQnHl/wX95hRgClmhU8VcOi/DohQbHzL5zOsYgEPvr76nK+hz5HpUOlGFIl2uf
i50KEmDFo7TqOx29tc6j2cZcZSAVd/HqVg59YSvSu/O5Xbuj2aJp4ZcDhWv2D0BlYtNBJ9zMpseY
fzqvUSUmzsU0wN3BbBmUcqzb2iXHAWgA2SkQsjN5lxQ+aRHD7C8JmEqAk8urlwcWbp+06joukWv2
u2iQpo0JjmQxfVGB3z8cjMqkPct3DTTHyFn+/y5spjhWKZuHAuLVl+MgDsUWaEnkoUF5DFA+TrTU
kAezQ3tdgW0CPjZBthjU8krlX//fKKrOKotPKwe//TjHSOaA4+owjsx1LK9v9Mf0fbfzL/63kWdd
oQnPUY3LERyMYTc4RMxkjTmpKRmueYrLVTklyqCcUk+MU1gQRf443PYlIr7x2VgWeoSsoNAIDYvV
2Z1dCrhOwTrCq6O0cIxJYqXQ/gatsOBmZkkLed1smIosyAOV/AjhTiGomFGC7vzAkLDtqazEVTn7
4DduvQidEeA7Wt9iremUVgOg3R14MXInYNxfZQhgUc5FRO3Xro/utxOMip/xsgkladuSboLX+j3l
AhKVKSDYZyQ5DcCJi3bNJPR65bkVLT0TAy6D+FNkmPvANnKuoxnozp7jM9fyS4AsaeWh92NJoBcr
Vu2/kXrZi4i+X0A3RnQLDHU5SSVwR4eZE8H0pQj2zCDLlmvYUvosUNYyPkRDaNcItMYSoyXGsO39
2qFOokLXwuZVfz+R//TpTkFX2lldcCqxJayc3I2RHjPTdA1hGmc+LeBIW3ZRQCAc9PQdRAeZaN7w
OY7CNjZYc4Bz7pJy6xY62tartHP8Cwg1DYWa/nh76GiLJ3lf2XZ0f6/w/TeImCSO3zDkoJ9L2++y
W0FKJJq1hvxF3RxuRESMPw+Zc1O8mDVdPAGMN7Ykb/pfrY1nnSkhIvmUYUDh94e1BWQsYGE1XmoY
yoRkMAlQwL1sEGWwKihLYflbIX+su4D+zLf09H3wfalv4sm6bHz5ad7qJJEB/u+E7S27bOhJxztl
YI+jrFmgCKmDxJjHFHEob1L9FWu58QTgFWoAVr6N3rD1gfTEFV/xJEzlvaTm6+9qgdZTAgQwoVo0
j+KPcL2fNz/UktjxLzT1N+bEHO/MR/ES7FtRAwjgG/XAJ2NAinTAOyotTnulkpLL3Nv7p8icLrQa
vwqNPOkdbJ154T39GB4/uef7zUemcxWu2WJsDoRD8pgqQGpypPGxZscd6bqYipDX4ROvllS8vA6Z
u5a9vsq23dw3XM3Y38pGyWNFMBG+wS2sgxRC7J8v9aM/FQBngDKjsX2FP5banM15EAI9XRRl+xlS
D3vYNu82QjHskVJ3tIIFdZ5R8bq4MTfTneFM1SapylU5l43TkpYJ1ac8UBIrOJ66huFrgkBILMcQ
MDxblkVdfaW3BwOyvd3I9NQsDNADT58o+f0qwSZ5Lt4vNadI6js2gFxtmdY8FvC8nGcyD/EvKf38
kVOKkKQa82WCq6RZeW4+GLWp5ZZ/cqX0c3OXPZK1F/DaUB8gYZuwGPVlAUmZAXJeOnM3XwmAMIM7
v1LKn8q/0axTKYsHw2rzgPfXXHkPVhD/2G+5/7PDzihy4BjWOVWLxEokFUwG59EXBHEL0RzmCv+L
CbCllg09a8O3o1DhWuzr9RN2fBazqtjZF1vRWf+HhQ8/bnacZkUKdRLkwk++zrTkZIncH+jCa82Y
ACWgQkZ6HtMxwmYB0RRJqVV5hUZspnMVfbQw3n82Sq0JaqU65FmRTbWOhX3MZniiCJ4DTg7qgVgw
U1Czbj+N2bYg+51pkhpuZPYE+SPVlITpo8erfxxaXSZDki/uHVjfBd3kb2DRY0J1xPT2SDhERzRX
XahKuccQW3ecEqMva+PXmrFMGF4bZay63gkoIXOG0SsmWLQiA5czTTQa/ruMY/1IHxqOZzWdSVjI
8V37k5I1p85NCz4G5fRk9lFBQ4ROr+SiQr7cZEvqHnCT9xxqnjwrLT0nGZpW9eW8I0nSvxb+aitn
NJOMWPYbNt8jhdh0ZRy+UjSCcPYg/Is+DZPrmiQXTi3Ur/dAd7k/KV0Cv19CVioEG+L+ZEHrLP5B
RWcss2kAsFBS5qVwiDc0m0B9f+x/GluTKliCWRRtvql0BOkC2b8u0aDUj6pJbTSqVBgl+T61z8Yg
CW/5IWlh/42NtI4y3Nte0bAj8es+XJkBQ3iZX2f4uZldI9M0D6+B7fAA8bxw3U1UCKDk9Fuq1a/G
ig2YF6OyEgpa0RG1x8Zm6uAKUOCoDBXKpu2Vyc/tmo5rnwc3A6bwkp4wAnBPvO5XmLfypErVR/Zb
z8t0h6R3J8Fv6VzArFESQ+SPHqTROr0VWmaHGvhC8tF4UwDAsGF6jPG8IV5AbMtHFD5ByYG79VjI
cX/9aXUlkGJQxaec/2OJsbjbERJL42o5KdrRhR0lXGVandPliPJKryxQeARZKQ6XeVtLR2geyAMe
qLa2m8b+GmDBltU4wCfaxzLW623ByygXO+2rQN5ffOKB9s/tQzdfNsdN78rgzLm9zabWlE7SgxWs
b8Jm51+6KZZVORQ3sWc2sVApWWqmCcaR92payDHh5tFeQf4Tr0PfO4L0DjtWV4e+MwQXWbGgVVRd
Sa9BTEjPHAWq6+Ed9U1KpRwD217H+OzWFBVj2xSGMVD+c3Ht1i1Cgq3k0sv/bZgCAvC51CxDqMCB
31xVYmpQoACS2SLvTpRT26z853kLYjp6Ox2Ij7Bux/tJSc7HukziLpkjbUCYpUmBwLSp7Ge00Gxi
+iZh3SzMXhQEV7Y/PVA6CviRY/kSW9W2tZYpSV5l2N3KTAOzJZmWjpQXt6I1VrIeFoZZPvFIeOvv
tU1b1pdraBtiYcEnLCWnl+iUS3g5MxAsiOlYlVYVS6YSf5yZQ2sPlt2rRBjl1Gz4Xlrf2VXo0l5s
5e9Ul/uMIMqcjhWL1/950ABd9+cUPDgJj84exmVMdXtD201tlfSnUsNhRcu1LVve7WGQfST+sE8X
Dqn65dqXpThzJ9bIijbVQQCgHE7mwhezF9eALHXD0BBnBvdDUaFweYPws0P8GOoA9hf4Lv72RvYi
1eDdxaQbBW1wqDUxkNNuE9ZRMXcspiObQh9UGTBp+l+Cpp1ykXWes5TEvTZ9H3GCdmNjh9IKvaMb
Moli1BipM6X5/ehq4fgwwCSzDygSLvnx2r6bMrnh1WOdhPFvPFssWgs1NOQw/uDjk+Ca3YIUkXiN
wmvF1ui6x65bevWOK/J6XAVyBTC+P8pqn5ktSN7Xu+ShZcjmXHmdNzqtS1GENDpo19nlm4/fF0Xs
OCI46SDWibybiAprV6DSW0ghGUfCw0VuvHum7t250JKNZzEH+x43r+ZcMDNMr43mb418la2agGuZ
an2x/inAnPWF3HijLfyg26x1s8lK7E07OJWSg/35fZVn5F2y+cS7cC7ShkW/lZ3tj1HG9Tg7Ribh
GD3CV7N0YLBSr8fvbI4kTJBJY+xAMY9MIai+F5XgY2krrqlwf08XUxeyjYOt0AibcxBPxCQsSI1G
9ntrYVNUzqOIy0ju/4nWrAnaI9at+/BqY9jiUERV4KzQRCJll34ntB5PVRiWCobUqv4K0ftIQTyi
D/ys14woQfBdi7HVtQGskaIw0p2e7Nm7d3wooSOshOwMgO156J5z87NrgUu4KkatQLiB4XnqIw/i
p3O/8mas1V7/1gJsg/TL7vPI0rT+7R5lxgeMEUPSxfIMMDj7tHMCGPpcTUE8QvN1aSk1ttjbIhbg
C5hGv0tZ1Wdbty3GE5n1mbC0gxANTDSaWclbk9/iVB8O+onRmkMqsXtT1T3exHuVu+H+cK9BXRjr
zvmQoUjxiSwnHeZkjLqrU7jMGKVl7c97Xh1HYuZ1ZxFmtSZc5zCGJkK7vIAhn33EUGaBvX3nAj8I
RaeTtVtsm1dMv0tij9ndzMmEAUoHdANOST56ojEoUAkBwtH81yYbDFmTUlRH93k+ku44U/wB3Zdy
o+Oyad55H493Eakc9g10vkuG4OeAx0/33ljJiF78IajG+WRME7MbQZ/Mma1Gb1ThT/2GEBEui5/d
wXzfF3VIXFa5jxopM/MLwFs/2Xz1fBjJX0Drky+0v6Wiy7UEMb4cAzoBXupaUD3zyzOj5ZH9D8ZZ
+yShkqs1dEWX1azWPhfYxzlrOFoVfhlktp1/b0J5NAGERfTiZn51BFGjrjIQhWtAqhf85qiV4kPg
+LGof4mSvUd6cjVHUDB94bERV86d2Ii+BZb/zMqq6ULilScR3+Su1CchzFUSLTCwmFJMAMjSGWE+
Qp/5Vl9v2uWgmzZL0ZA2PL+50QH3gHRnPVOEH7wNnNDEryEMhXQRjWJW/xhL9tgATUj3Mv1Na5GH
LdW8ek2CFxuVPCqTz7kxYhN34DlDZ2a+43k/jt9XIfGqJJ5uxv82F/72pnXin5OW9eBG4aqFSkDO
R/KZAWFJOnd7fLEjw/E4N47XYq2THd2WbJWUxLXWYWduTSzs0v2ULIc/Oe3jO5q1DikMH1JX4jV6
aTvTwI6KYzZQLyW2A/VrNxONbU56tZ+4lvAfxBTeqLfGrdYV+kfVV8GrT9BXosTCKpX5fkgAfjRc
nm6eMRkvSBOL6itt785zEvymo3nVjbIDQwqMPh+7oX+HPq+N5cToxZlynzHw7lHiVoRnkA83C/ON
6urS0T7ULmYqXeOxOM/VzrJ+95nWItUt0JfBhD2wL355mn6Ln1DeieznoyyzLY6hiO2OQH1CGdU4
vsqTL7rEG+9AmtTcnw+VenPxzJ0Q3zKbY/Fuu8WK7fx7mvkucztSRbM5RGUHqsWThLzTebuuDjiu
vMHQ6cRzH4EGUa0YtjECC8nCyON/e77GUNZiuPDKXdYj/a/DnhNQfcDm9ub1phONsA1JFJhyiWjJ
4ky54qiJIyjXzz/Mqn+RhvVobM10UhE4GAE+cg6mTA9ViPXunS2av4KFDw93Kc3Clp7PonARFm49
nm1SJgIodSOQhJOAg/AAUB623vEdjX/xq9ROThROUwe33inrLVjm5JKh3T6+qHYYTqyUYynP2GVN
6Hpt2ExOTPDWRFJw7auN7jFrmlJjcSf2g6kEWvad+fuuuzRUpYxQPl+c0sOfHGhZ4qLLG55OFbvM
OxVNm5DWtAfEKA30C6tEgE+vY8niVFOfaXQtQRPz7XR/aGwxeFZUkKw96GdHGFraueH+mdyLUhgY
9ciFqUYxWEt7aX3CsTYM66kuRq4vdnphChJkqbMkHi6R6nTaehJGdj8Bo+vGhMKT9XBJPUN0p1xK
GZIuqinfT/5zDeEEqVQ8nVftNegtCkN4FP8fj2M8H/t4b65jAGik7nTfF5b77ipXzVVWFp2+QeBx
zMquWxnw4ljI39kwDh2NNH+VwaQeGgmCo+ZBbFFM4fgU8uh0SBqLQm+QpGt6myN0LVgs+rmFNgNR
PBEEbzb3Y1/82dT5V+Id7EpLDeeUFqNsb0MRJ35FGHolH3JwXdG5sc4asneP0veESs5nce1tjOvg
MsDgo9Xji4ShXwbOhIiLSwqN/XqdN45Ik//xkTU5Q5y/NcB0SI2WrPAmxi9tOn4ZD6bD8tBIPmiM
o8bVzrrdhj7Kug4eUMy9yJl/TfvSJuBpO0NWFfIc6XKC8EdwjrV1yPaz5pV9Ncy1vDoreZDYjMHM
DtNP3sgJ1i8TrHCwxsaMpmVYNcTSuZwo6d8OvlRqSMpKImal5qOfe9HpYLXM3h2tOZu2EzXOJ+GW
ABR93BMYfqSs1yd65IqnMvcim85DIwmRDKqCPm3bOH8jSu0ctjT2Dc9hySGa0wHbYeVkQg/czMw+
7MXTNSljOS6YoK0pHu5ZlhCxQoQi8KoaeqTaxEEDDx6315SQrsw71eII6x66z3caCy/RWCZUePdx
lRBqE5R7y/Y/L/7ZFbGQBjcWFvh1ZYlyHOUjYlzlxFy2H67fTQUzouC1bmjMjAi9VSdjrDv/pBs/
XhLF6RuZqybAc+9r7HusvhNxCGz3JZzHA5zjHQ/mV9AoR1L72GFInohiRBtX9DG0wXiHRHY8rLG7
08uGzDwGaIAu1gNN6mgzMO85ZuAZ3+LgsAtiuyAkbWkJU1SxuWtT04tqaRTBqOjITyZmsPkQVhnj
jZwnuRJzERcRsFP3uX0WG87HZWucJP0mNWbZt65BZaOH60SWlyDKQvLfj1XjY0dMSYyxLIYrUdQN
Xnf1dlsUEUx48LBVAyGGbkeHbggBOtptqNVjUSBG9A7g6znU29IRqf3VsORIkvksnpJGTBDB4Qxc
GdmARM1SwYU9o4bdeXFXfL3QGXQPYhUjzBnFbcCC16mzsNszos8XnoiDz39dsoqhdYZcFh+mIELE
wtgoT0amVy4QrKztM2j0K5xTrNB7QGx0Sja1WJj4Z7MrEAXK5cy+FFeNl+3TzIUsykfoFEmi6k4K
8ezn6eudAgbdv8WpfXEu4Uo1OhLY6HbKh1LmesPADIAWMmJS1Gp4Ucl0pp71hROzGmVXfxoRiXCf
NjNrZqFo53/P/b27yeoB71UOeTL+ZjIeER9hxYXtYwk1wwJy6eM++X6AqbDU7nFoCVvOdgpSjvmR
pQs+VzpC1b1Ns2HAUDgzB65kb50w2KaU4ubcYtN31gOHSuHD4kKI6D1b1RlPZpvdccKvXK8SukT1
iRxTfSOgtE4aGFGg/MImcmQtP4v6qbc73XU/3RLB4Lg3DqH/QNSkcQeZT9ba80Va/EkHhEQbaoxa
g1YpDvJDStFlJ7VarWylLXapl/JhmJrGZkcGVsp3FCGeVNeSn4Kv1PZaJms+SjACKvWKndSF6q2p
sfD26npnLNeyo+zVR5J85CPvzb7sIQweNe1cRD0c6Rf9yrUPeYJAzotaXg5rkpoWipZvaGxTGVeX
VCTV4TmNXHoFRVFpw879DTnb5S1F6QyR0YZQ3Yfou+SvCjeFDo301NpSzUN3xrAueIXiw93uZbau
AfI0HSGo0eCMAKWGICIF9RsLq/ZI12nsuaAZvNogqwpc9ZwD0j0fpqttjtX8JA+NRC99Ou4agKSD
gSz5AyXifmZL0Tio04mJY+Wo8rQddmJzQ9KV1/WfYeoPj4+a2SVaWUtA+OVdZE9oeFkr3rrMuAyY
wUM8jvDfRXqTyyJqoOCjR62sYWvzP7Kn7xlqQHlo6vyynWthGHmeoJuG2vrm4dIV3hgC2vWQaCIM
wWsaV1Tu13F5tLjkCwBbe7bgEo0c/8y8z6juRlqF54mIj8ztgOGNZYDo1XXN7unGvQsxobY63cIp
OwTWKP5u5h9Y392kPUxq+CWslfngEfE3KHXbPSO0rkTRxe5/uo+C/CoNKkOL20CBp4xZYDebnYSE
oKktVCjdNGfu99Sq/fBYJlkkuOAQJeM0YxLEb//ZbNEnZMg0GrmIr2bwx42vwM2fzB82HzwGbPi9
4S2VzT7Yppq99pz7NIoydl5AkyXunF4DwvKC26b8bGijOa5ovAgSf2FscQC4GOyIJiY9/PuNgz5u
1ffSc3ETB5ug7djMhMwGuhahVYQg+MFoEEOo7u0nTuDhUTuwqU4Tjgm2HN2Xex1u+YF4B5jfjdn4
CqSjT1pqXQxepJCY9SzRJ+hMUXk06e3xJRg7GWArKFOEf6hhFj+gGUTWyVndmyDT+0HH02TgeXGp
N4CQmhzvOI8eoOIl6tGGm0c75zyyCwzZwVRmNyHOkWo/AadcrtZvXT+HPWjeHGflxN5qAF1X5hJL
BAQOv1toRFV2MznwREYG0wFmaGlERpbem89NevzffWApiTxyh+6zoIGFXsk1d2aFCaBb1WvNLqWK
LUybRInBg2EZgWE5Mip7czgocgqxQYj26ArNmBwZI9m15henBMQtdBDuKrkSpn0nXPSNnv4RPbyh
kyGwzo8fvKLfz9P6fMQbdRk/FOIB5UDVFjpFDSaLNdXSNbSKn7TsPAOK21fzI0vv/A2wUj1zL1Pu
0gGxrfNV6MfqRRD9mIfHgFW5OLPOY8ZA7wF7UVgwDkPGZFN8Px3J3WWVjzE3VZTseXyLwEE9m2Hz
KX9I4I3KbVy183Bnxho0pv5tyGBwvWHHaARouLL4JC/pMn3b3aNqvAOUWJvAiRQAHQHarNXg5hnw
Wp/m/M6DykQfb4VWRaKp11OaiJ3aMOWzOs7+qqwFFQLx/KHJA5UfAzk4i0xW/SpQtTdqS9JkyQli
5yDChkQWJ7Ckyf2M2ILXkFU5qtBFxcHvLCCibOPvdsmr/orKF13W8Rs7RcDlDfqJnS01v9jDcAer
D7yzs9AQpeiTebsXn8OvSJeAu29tV45DqrSgoVZMVJlNsSBL0zK5FXIjZfOvp3lRuj9wbNJDBO3c
9hUUb0To5oIvoGdLgJ9HrjtAQ9BNyZ8hNP+z12J6BGYKbj7/mQ4f2cHnjHrBU2vNVrzoUwDooTjW
Nw/bz1EPYBmkV9XFn5Mh8nllmWStFSM4XDwMHvS7xWnxzvcR6fXVxuyU61AfvGPY5/jH0K2wlKY/
6C4wcnefhsTkPHSMUChxVsYH3jULenkI8M782PLD0HViHI6n7vsNchbu7/PzgLFtLnzQNNymswoV
yuvHIy3zct1o3jeyvUsIUcXTkp4yZH5SWB0qiMWnsDNNur/gRfn3Ne9M0AvxNr3RG12OoFNydGjR
z4A7iNH9AgY82pfzg7oj711QplmtT9RCyNcfWVPMt9wYDBXu/iKTeBgqtGwFN/blRZmBTW1mQX8J
g/by1nFtAFigPQCg37VCH1lwAu4elt72uToK4gGWPnjLjhEp6nQJV7tSkNlb3NbzXs7Z2jeaRy+q
E5anSi8wjAmHncNttAAkRUEweQ5q2ig9KkHDOLvedJzNprjhVultDt+2PLS3gO22TtZc9hY6dTOt
G89xePXwGcmB2gEA6+8r4+Y7a7wlPldlNf2CK6GLJkADElk9wSdhB3bVNrma6xuS48BXUhw6e+z/
yrtzhTcIuDxBdTgSmXnK8SkhQXhpzwZaNCQfXxRKq3e9j0JAhBRz4u6XT32su/pWqRjTT+KmNmEv
HjDMFKNQfQxscN3N5qMENa0YXWCMVwdxupQ0yKSusI65LUlrIvKtj7IyzcXYhmGnZ/AvzWPQM5qF
Fp1LqI+I4OcIm2TF8B2zSQ0ex8Rrtf/ltQW2sg9jDqC8lP185kI0/tOjItaZI+8sX8kIHTup8QYP
tKnmV32jRGHmYtrObDmJcmhEWGlwYldUMZfK9n0Len0k+isKVt834IEyhZM38Q5o7EFwO7yfHVvg
JiIVGoiQIY94G+nMQZpVRDeSdzdGYZc6S9hTZfzH0vQqf3KACq4FoxVOGm4x617vEPu72jXoIYDN
6kJdhMsS6rTZfz2t8g6rqwULrd/A3Zd2MVJMzDvDcZCKaPmA8oh4CI8qtvhH5/Q+JAggnuq0rI3k
l9HD7KB+fm8bXqda9VC+JylE2Yjhp6XqDBUiI0dcr8ssqmrx7/UuDm5eYwZQzT7Pg7ZorGYcdMRr
HK5qC4KHR/Y5Ixku3jfrzTt9cHyaeJqSCv5lpqNdAe/6zkPNlrTF5U5E4/NmDGSjcMvvA8a5Ymo8
ZsMBcxngfmhpREQtpTSI9wkwMA+xoh9ANzelVbbfhRuFtekHfQRb+lQxRvdzaySq1L0ZHPAlzRcE
2x/jxyjjeyoh0Fe01a6NMS39zLdAc2gLocJR0KOuc7zLm3H2TjgLRjB4RAYvZWuX5RAYHeNusvM0
OZY3w3m2AHPbuRcEm7ag9HaRkspc9rPMEvxVLpE+ZlnQacaQux5UL9w1Fl/g9jkTj4OYSBelrPsf
dC7lNa9T4T2aqeiY4ERPDfxr+euRGCluKKqaqJWQ0yuJpeYJo56RDtci7G9eOnIeRP7QnGMEelKw
nTCEIt7l7uKO+wAcwyFVOHEe2spoN9FXAl+92Z/UVeog4A5YbCai6oG+sHBzNF7MBXmdQ+FHMSl2
kwInZ7Ta+ieKt6fSBKStyeLR2lFiuQQK80P8AcQEwHnpfIXs8r1RjIHhkeMN147scD8I3aIS/1/J
dxweNzwBh8iTbksgfB6IV/560n2sWozU/OKe7GwkL2B5c8+Lsb4MY7IeVnf+krkbdnvJC4yCbGvj
0fzmnQHBnsn+F4VKUVD/BadWQnLuwk8GLs8cDY02cy4d3b2VMPIkp93Z2dDXOP1vGrWbvo5glMcP
HTXMgdfIYq9EzcqLKE5m6klPm4AIvKfbfnEsDH4Y5Bc1lSKvikbi5Ww0VDo2kvER1lNRcZQ8lbPC
mRL/FDnq0G9R3jXIIKLJRNpBgrSKEgaBEPmZ+SjubtzMvCCwxw0CRTrDRBrgTpfuGTaNdtWYK2UH
JblbhMvlIZcLTK5UEEBpE23aMyTr/AXe6Q5fFFrJI7TyHSlncZp4L2KZddamQ+Yiig/cnna65hhA
kilDLcGXYpx1g99dpTF8Oi0VxKBmUynT5uJzbhMgYP0seCJ6D6rPP26K104kQwBAOieic11qafd1
0RQK5JNanjpex6O/gH7vz3dQJR+zotMvpCnIV9KIUpqowM78Uj6ADpwyl55SqcZ8zEYYihd8Nxcs
ULnqv/zqNQiF8kvVWrhl0IxvarcWXO5G65E5fXhZs5RTxK1ux1+fIIPBgkFuM+hW2HrYJpbgxl0o
ThRbFZNU+kQ/Vj8FEIDJ7RQpnINO3LfFouAfm+O2QU1yyHAfqGmdFiDHk4akcDmdOxyU/wJXWHWm
T3dSjjvKT9BQiVUB8x51TZbNlrOdG6JBGmgmZT1IAUaE2+M+2sUvE3s3MyKS/WADAvGIlRYd4bJn
ittgTIagU98yzPNtif9QSUAeKGCWj9RmpvXmLOAYDHx1q7AfZghZkRJ358thUBcHtxyhDONBb54e
jtRvrbTeeloP8J4DleQPpXbrtDsk+lV6KwX46bDOmFHa/ngcKflubR+AsL3Iun1xbBverHYFGO0m
bRiVDHWaeugv4dAh0+pASWRXoC82jKurEktKqmD9/J1cNS4kd43UPL3C5tjtI3PH60HLDyA9qEC7
ZWNEBfn/IP0oa/T8tzF+OSkil/ewDychZAZIzldBNWQXqyQwUyxJOUGefv/paR9fKuVTRi3TsPuZ
+h0Kko6HCA3bN5xnJ+xf2x4msfnjke6oFH4hkPrueFiYE3tE0Ewh2/N1nVDGkNEoUWNqKCjhsAYI
bxCu9O6nOsBj0RUEe+FRaw+2AMubr4jNOhOx/Apmmbv75duQSenFCDWX4nlb6tsJuI43dvSrDRZu
G61zf7cewMVQRwb9tHNH3hC7SADMspP6TS5TqEO+WSqllea+0pakgiVKjSplxco0LxczMxYT08VE
PrHb5714CyEklBR31hQ9LvbBZcEehnuAC/hnQGwblLb/d6wvqLX73SGBu4wJT2sk8AGPdzIvBL3s
dOWN6X+U0np/5jdbwrtH8XiyZN5Q5w4clXFYokD3gITEhhykic0yRz/FdB0Kxua2+UDzwNoAzG31
rg9NKXjmUSz71K7bok6wsa6u03jteBTqKgQJ/C603fum3710odjypQowSrssy5wgGKDU9NNlyrWg
B5TpAyId3H8dMmgKgiZbymlBfB+A2ndA1HEUkG8D1cYj9JG/rDb6A15let6Fw2+WzPAOx7IOAJwR
r6O+ULbrBrFgBKtQutoh3t+graTEekfam1ILd6L8zm51q7YvzNgTsGJFpb+r+PlrNHJDZJOOd5Ie
XKJbFe01Y8nbUL4xWkn+DtcGGL9zg3flZNMAfR/tKfeuFWZv5DVN+n1Bt3aF4x6cdx//hWDdcSNZ
lUGcldSytxO66/grp4SCDpXBpU6QWZ3zs3MIdtG3A8MfMC2gQWIiMHgBKVkOvRvAaVKjzferjNAe
qoUrDT9MzYWKCh56JvH+eY/j3zAJvCAzYIDFTB2CcjllKoIpewTt1v6PbpAkRas7EfGzIWgp+KcQ
Eau4xFjpKdgEJN3fQsBgbgOhWDfD4JLAIRWTGVW+aO/gt7LONZex2v604RvmKwh+jgTqVr/2kAGU
F95k8H4Q9YVg5ovprJb6zhgXM2na2ylaf0PTRjtc6npNQ0hiInxAyBOGpHjlPR2PpbmWT0KN4r2D
F1SCcw7tRBZQtiN8PJJxGSy7gPBzRJEGfX15Oxv/pMwIddTtWu47zqmLpQ/tuUYV6TJouRxWr3M/
mGSjzqXHNh4SXWWVWfq6uTEkGjDi9910QBrSPgVBOETpoT6QSqtMBsQ+T89PO0RvXQxnJprSJJyA
GDj1c61Ubposhrcx4ch4VdHZMBt7rj4GnpIC9g03WzidfbreA2cO7n5X19JMeaSVHEptqUgXxTXr
OmZEEFc+rzLFpzf/GQEAbQXx6lSfLKeGD1/jH7JLIHlGZqWjTIYHEqTPJlkpqGVxnEHgq4zD5v1g
+T3qfNy+lxcCyfS8Tsy6hsuO0XTb5Dqjkpi4wc+9t3SY92m9x1Zu/tSa+uMUG2hVIgoPxM0XBSNv
i7EkZ8pAVhNBGnsixeTsumfQlK0nQk/Y9CuGBE3ZifCFQYHKkGySM55jscO6w5zmcHbifiPnYAb5
RLsvEmvSn9jHefbkIbrlq9i87tE/El8A3693ijHd+xXJxPepiS2kSUHBprvOqTy7pGwHIf+doOFM
G78OdxAGtyke/k17QlOzhgIlLYcq4eV/gPwwR5p0kVX8UWMlcXfWrAhu779q7+/ppmhBx6eeX4PP
j17HTOaxGSUhnpzFBJoymSXbna3EzpVTMOH0ChbmyEVOjQB4ozgeR1m2vQulaFnNS7Dyh6iiOuf3
Uc4mzCqvGB1PHkZl0m8hjTvcyNo6zwBO8kRYXV6kLZtEX/x/htAJbOc4OOt8CEuQNN1E/rfHJTwc
4R1CGWMqSElk91/3wzOG2tQrkaIabAhp9vNcGXsPoYEiaGnPZqb87igxPtq02nXqXtsB7LVYqilB
MxM7naVKMoOPT12fJ2LLkErhKI0ChGHQUJ6bN321168XKzaJ5lEdxgOpaAlgVmnnqx8hSoHHfJhw
F8uUW98/1T2XFTCulamiHpZKqK61pPW+PSGn15LVumzfj54Jeb7qOu1q9JQ1r2DP6lNzNgbs8vst
94iZ7JA755+0D56w8JvjxGj1D4FzmXnBAeeAtLOybb7v3yeV7Pek78Bnc1yJHTGbcUsuvPU5aqfO
lwxwM1yJfdH9HTO+Xd60FV0yzrLWodUg4LoGqukvN1386kNVRo0GoGbaY5vfurNqPvZyJWwQzU8E
MurYYyg4VYFy/CFsAOCRU6tWn7Bf38edLQliKuGkl0oMA7O4IThNAUgySQ/zYCzVGg3olIOFzqMK
ZTq/ycv9HoSNV/QxnlgRiat3n40zGjp/oQ/51mJpcHicNoLYtvKNCROuaxxDDsSw0hzrtDPYUEIX
QdSKM4XBfPhf67guCJji5NyGxwSD0yAjGs6nyyXXs7ewuQ9CgN81DEYaQdWVXZlhgQZFTEC1+WY/
rQKAokzmsviaxV74kNxZjO1D83kEhSSerO7RmwVeNklt72T7bSDz7G/bNhGMzEela4ILqa5Z3IKO
Eh04puHT8BTndxyAzqOuXU9LAc+oxhaoF9Kyo89DOCLm8JxZN778zsVbUUdlXvafbJP83M6L/DLP
wtrAVu8ryyl/5yGVlRglFleXW0DC4Dm/QnTCDiLFOaT9+yhvFK4vsH5F7ZOBBX1h4ovTGHY0WKzw
4v7e4TlrYAjjhXKUlZ6W0idWzVBwQ7ZfIIMAjmlgduD7D8BJdm2iP2J2DmeihjjKsvSRPcL0sm5X
V3iDNTYkg3szXKYRC/+GPI1MuErMdJzngmnOzu0rgPfvRmZ40iz1gtOhdbXTEThe5XUGmWoQjcCu
CQRJdd7l0uAbXUGNLklKwc3gvmVAZSJKyAgsCrhgD7rQ48jYuILFuY+RTVTmJCG8xr6YQfmrFCzw
vEltEC8fUCUzNF+hbh0pgi5UzciCV1TaUT7mdBCmtfRkcFypSAC4aYE/LdoFYSz4e55t8kCfmD/q
q9y0ofcQFgEl0og+rVKurvkuaywlSYG+kDn9R2oQlYV+nzyXy6YKjW6A9jE1KkuwmltbVuxU66sY
d+ufQzoML2D/twC0Es9NMUk5GRRrMfpnWYdPsNiHoK6lKGI0HC5WlA16v7aULK1qHOfb6aAWkQT4
J1jhsGm09Y0wU5Nb1X6SYbsG2xR6YAqHaQwY4gG4bEw3GBxi62AoIFLpheabjJF+cqIBzanuPxSv
doSqZv6VsDCxMi2l0B913WTxXvR9pPgK9F4/vkgb+tqBL1SQeFwrOFLsvBtNh51yJv+lhwtrqwkJ
qAosZDddayYd/5X6sgJUfUn96QoKc45vv2qLusFLScTZDDue8KfzN4j9KfW997e5+X9KomgJCkbQ
WQbE/G4tUVPpm9pYjAvp2pYKxX28/a8/SaHGXAq1KsJ3AEBNSwUJVmDDoSv9Q0AkRA9dJl97xFLX
CFX0bLpJbcKeyHrCub3YMetQ8dxkc/M7VOjGZ0/7++LBlJLtVaNc83outJBxjGrosp9wBTIcM+93
LUqYQhwUrXE2RF7b4j8frAyjDp8S/4fO7KBtCehAJDlpRIFhRTTpvEftnu9cIEK2QiUdGBke0KA/
WlRMZcEaaYdJb/LCMxDpwEHDDsVaCGicRavyiXvCaS8CwykQQtZVSAFz++80a0dC3WcW47qO9Rfh
r6w4giVJAzPyQ3XILMuga0YD1AbIes12xDYXf1RsqI54qWU/3MgHUu2eK8GNkWOnTAefxOFlw1M7
PSw24iWHmfqVJ6EFMuC2DuSPZ5Ra6mXdYY2zHpKtYATlbWW7zTXqhifxoqS2pDf9N0zT6W/JThnv
pY/8PQNtn/pFFFQZzknubYGxwQdgcPbP9k9QipgwUiMh57NnO4ILtYE4pEnJbzVpog8oaw5a8EkE
lLE+v0wn+KtAlLk5CkfMB5vdcfYMEYG2QZJjHePafAsNjzLkfWkjCgizAFr688XKAPKbNVlWBxbO
B3hx5L05uhurw6JbTmKk75iwNSKql2dY4gMGs7qBQw1eWDBdeEAIaFLFsoR9M+/AUA2tJlQ8KuUq
gGMDfJOKsvdBSycjOO95SQpdbS6H0xFNzWq1N090Ikeau8866TwsHrxzquXJxl+TCfY4lrjZ+A62
vNsip9dgCjBBPQ5N5ACLYLXyVB2qFTYZJh0tXiEemzrSQ2yL+fiCtY1bBZvJmPzLT29caHgwd+A1
SfZNIuPEooMJ3C5rqa3U40w+efMK7SGQz80cuXGyVgg905l9HgKXGvgS0RgNBM2H6Tvhp+KpCIMA
To0dQ5AEOOWn3F0ud6FtlvR/tMTZ42ZkIBsuLs9p0UJoCe/my+oFB1c1IrYQZrPO84ukA0Nv/VLP
7ZiqjZNwPybcRfi2s2TxKOHODylxHyyke2ymAo/QA5eAX83td0syPZWERWyJWpKAeLgG2OjzMY75
3AS2ACcguEMZihDB3tmUF/da50qvVBqxVDPuVcc7ygheCxCsmn2aVFpY1Z+FNC2dEnrB58z3krWY
lRYmGJ78ikHIyPgFUjjspzn860jml7dw5mpAhoc/lU0fKYnZnJn2LHWPmqdbvPPmrXF8rL2eV2rA
M72AAuW7aY0nXYLSR+7P8K1DRjO/J7X7aSUjMsjThWCLzfUEd/y8Dg4ogsy5aQvkRkyhxNopctS2
3o35rhlNtf1Kt+IDUgWHw75B4EXKbDKhh1YBBzf7ZmsmZq4uXZ6BV4kvEaSV379b7UbRFrrkR1hi
i/1Lt+U47tvjEKYj3GMiiBQsKrdml4unw/vPL+NC4Q9yqVQeOYyaTkwFzPH+657XywJ6dU5k2nJQ
vWVeVesK8SJLGu/EAW+0jvSjI896EAtClYdJWK90pukWhTPu0yUmcLm2eRqKyx1c15OSAyWsjfN9
GjYWwkS6V1IOhXYr7CqyUBV4uPnr3SmW0ik/ZuaIv5SwXO5dEYPR1FkearlISJJHhRFP+rcFN5nm
4IXbqw6DPT02hhCrUdQlJlZs6+lVa9BN7bnajI0dXIAZMcylYwciT4M4p00u0ppfNWQHyH76bQVV
vHJDsxCXFLdKD7g7OiLcU7YQDo+XISn62hON6gxd0fzEkIApsvevX7+Gut7+sw4r84y9QunanOrv
9WmFP3KJJgEcp7Sq+qyu9+1zYrlS8WsYegwByuigB+9oqRjZ3ZivXUWOridRB/l1FiuhPVEkjd7b
eC+UeD3veJ62z4JBrU2Bh617iAQgJ+efIoMsU5qNXlo2Yu9LHxJMBqfgo85Mj7odpYRuacgBJN2b
BNCzx8zKfDJS7dyOf5lRmP6fLLACKnXO6Zo0peigKUEykJCbwVj0ovPNLbUHn5qJ8gQ3BxmdmG4B
SGNDwsnhttUffjU5j0RuThC54r1VIugf59emVuB3V3C2eiOH6zYTigwRa6iTjLH31t1ZWMzrVQnX
A2K2Z7WB+9qZt8WXLonxW9O7yHCStKdrh/Vl1YXMDBdltdnApVJ7Fsngn1FaOkJUh4RbR9vZk0ET
yxAz6DP25VAETLEq1CuPJ5Ku0AsFQAA7UWn4CoGV62YXXWhL2+z5uoSRX5Y91zIMVVlRgTC84Vl0
8AzEA5FWY39ySRojuBUQAtZ01emEjUDYwv7XDAMaD5fVaeZSG2gJo6XGAKlxVHr1de8W2JVm6OPd
9HknzH7Ug9X/AxM9HvgfPirYXTP7qtTyP3eilsKvMZ/PagIftxBy1ALUPfOLcKiXRjfnQEHwqFzh
vWrNr2wa0dD6ZJJIPaRyHeckY0fr8pvIFEGPvENMnPncl8uh0Q49Fsot+2uzzsjPYIsKJoIX+zBr
P00YemaPbWVCWuCQKdxSi0yYh3JtEGdMsMd+YsH2hJ8BY+PCpsbo/yZQF05HICQ2bpi5TL14U3RC
V6oHfzU8TJzMakWZigXanubXj/Ckwx/hRKsH9WCj19Kl1NXMi3V7nJRbdipxB692xgPN71McxQ6Y
io+r5t70zPi0v1HGZgoCg3yOOunM1x+GNHtFcvsy8kNCpiDvhrkdFoCazLFIRx8CissSxm8k74ax
7v46kAMf5LV2LFKRroB8cDKt39bZ3i2NUqPvfevUPR38GZbTGjACGVXrKSfcjjVRCg6OKNoi0H2h
smmQQm3eazBlC6VD6qlREEqzQ909l8PfHtKuCqhfAvYJNNODQmsyWoBlLuo4qoCyDObaEW6TG8sU
wIa/bNBq4JdBON/HcDaBpXulDHpVBnYvWkJRZGq4n/Eg18WmlWP0punMQwFSol5F5x04fixhXUcS
cNg5YKKe3jEY8QW9P+jI/exIewpOcJs/qEwRj77uPrUDe+9oipaDM1nMv40N3SNMmqwODYCHA5HD
n+z3ROUhalV9lzUpP+/+tXyLfthfJrTgzHkIjAjdhwA72+inea75HCwbmhqstQIVs/xBe2MoKu64
c/8N40FsLjrfZnKEi1wquTqdQ4v/E8b0JY91NB6zumZuPcicRxBfUm1QrzcxufRZSpP5UuJvO6lq
6l2zegPNpp17SIntMw0I1DPJWZwFCwv/vSqiie1cMKDF1L5Wms7zgWlBIqZWH2VDVCrBOFvTRnG6
GkOjDvYOd7+7Jgd6UUyGT4qbglaF6lwJFueREtHTCZ/doZ8xWsYk0vVzhjg9ZmeJMsceBVsmRqlI
+lIVXbce0FpbzuDSE3ALUzFfviTYpgdqBRdnroRtdghMEHx+Rsg3G1osLnD7aZJQZYxabLYD7nkp
h8oW9oLP2VduSpXm4mYfIsqW2ty1euyVTlxT/4twmV+mVoIVEeJhHbqQYyPy1mHjDefueyXb1w38
DiBg3ZHp5Q6PXVkC/Xo34HI7kaqgSPn/Dit1LMwoY95ffBfiMeqSNcyjJgW/rBfMOEoedKT1Qnea
oTt0Nol0SXLfS52w8lWt5LkCh7t3JJvRpg3iZC0NbpzuJEceNebTBebyjv/3i64ZBChdMXcotmaN
JHsS10wwMXnte4ohaYEZSOeNiy2+F+0QD1DOwrJuBuyrGTKxxFAN/ZDBKuMzLk1Y4b7rI9N8MeqO
+U4uPsoIUOPm2Sj3jX/n+rrpCc68nYoaKIOvvUq3Cc+MEoDePQtTgpPN/oGnwmycX8Cb0LYrRRcn
trQF88eeXszMjQqc9Gd7eK3dnEu4ESNphMzKvxOuX6zExY5Jirhj+fKMk4LMwaWkX2AcDzrGW4Wy
C4M2NmKxTroH5Gn9YMSoMRz0X9hFZGVIoU+hXwWJdRFqEw67yRdjgEZg/AWDziu6LUdyBi1UlL19
vrsOdZ9UxFVehr2TGPwLpaCyHI2eUi4ECuaEb1gueaALCM8vIS2DhWQbaaHeni68arMiXUE50dpV
bu6KmsrxJ+vaQ5LPNSWvpYbZaR90cQknHGIhGfOu4Al6YcTiRH6mA/Z4ZE9AURTYBvzNjnjioE1Y
nTj43//90MzhEE/kxsoKiL+kYCPjPEDAhEWtBokuV3io7XTrVfjWBzvhIzIUr3hgG+bcq60GoJ/5
MY1FZ0ewqt3t6gNZQvj+3c7g4gyELfjOVZPBmZdFks8e/hPsyAjLsm9zeYKNAYzdCWghToYWJO1D
yME0nqj7R7nowIgl4BBTIKu3zVVzx5YsJ0WAQv3tSkLxYpH2nMKEFlOHlt/ewHBXqlM2rR/gqVAS
qohDiYsuODgK0lCqA5naOcw3+N1J9dGmdoiA3Z5UVcpAdG6jlXg6P7+yRxuSCBQOnBU1Hl/Do7d3
GADt9KKwhelGFG1ixct8JS2MwcBHYLYcDPNE7xeU7NCky3ks+jex2ZsQ/PXq8W3bIRuUYt2gT8X3
1XWBR58setWfR2KWGQl4q9lvgpnLYw1hUOqD9exFp1Jnydg9WSYNpiZFdMZVHX7vCIGwlihTpEud
9p9jddfoHwIE9T5wahgaib13M0+eL3QjvFgoZeQ7pmzE82SIytgTqNe8kzY74OPIuBn9S1JPi42v
mTByTd8iIewlpnowxzUHDr4Ej6FeKIUn9ANoQN9L8m9GBSv1Ycu92pnCAKy8vU6mDyjSkMqIFrzR
UdZZNfLig4NPFzHRvEi+xibNYsvqb2+D2+re2wqQMbHprUX5FoBOhgqtGqu7L5GuOIQY6RX66G9T
BoffhdiQeP5tKPzXfltuJCcH88k2m4X7rIO4KKWc0p/g4eZeE4gxNhiZxUBQ89DJnZYKjWSNytfV
0TYYL3yFp7OrUVIGbCUSveqi5hEVC4g1feKDAHaSE6WcqwddJ3OmwNmt0raZxCxpfYDlalRjjjfa
tYlXaSbsPPkavVE/8spnmYx5F3Zud9InJgwin5AZA0CiMZWSTkkDSHDu9y32D7bIN2pGdDZtC74b
quxVMbTIPUprAArv7V2A3bJgDTB0sT839Jececl1cLhyG4DW04wDh0b+xI18pVmZ6Kc5UygCks1q
j1AOPgpib/S/UrRqHC/+BGfz5QV4vkFiHpZ5DFQx6XYYeJ6XHRJd6+1E7y3H1iJDdCdnOcfohi83
RAVB74aCtul6HgjU1jadN1tF3Qds7dHSqF6MkIho6iH8i6Nyb5HdibSf+jX1Lt/sfQaBr+HFpT5r
esp72Mty33bFgCSxPlh0iPel8l/I396Ls0rSHTRXrCxUPzesMz1TAlAQ46/rz5n/58kWKfAigxqt
+9I5VDO6oleQaoEhm2flWdeGfBqaOGxBeXk2zonODQwvWKK6RcSOBRm2UbwZqp79MjKa/PqMQ9pI
c8ci1P3da7ejmUwljIgBbHb3AidhIS8qjKdUr4T08Opo2ZztWQtuLgGV8lo7vvpwqOPI7dGb9ZRE
UnV2KNZijusbX4nIYjp+xpp7gL7OTGQjcqrknzhl+os0UQPmlm7eVmrmCu/u+NVpgbhnLcJ3k3a7
jgX0pw0o4QjI4bqQGCWnJFzzac4z11yvS90TjFfqEsCqKLYKSVVQmmeojWgkzbS83baNyGk45eWY
wODI0DDVWirDY+ZbfND74ltOL9U4dxL2/fdvA7LIxdwMYP3qF6GpM+9i5OCJiVosxjubOC7sAYPT
n6hWUojtlOmsyEZTgDY+DY2JlvV93aUWtDIRnABhrI9Ow66pblI3zBNXl5WDxMVoA8jrZG2IbgI6
ToJcenuyES2m8/6k0Q0/k8gWpZ1s8b38M2ys67QvcdvICDezWYsI+4gDllfjDvg1OMZnUzhbvQm9
7aUqP+8OWGcvE9RrSyrzquQaDHurQ/pHv90hazT8aQCsdkSJaTXpceyThcIE4d6/g+OgsyzxsObF
GE/NFoMSJYb9Ga8ITfyhdwe5acVxh78nKFxTrGWOxIWxNG7Q/dez3KDlWEgpQso2C69EtUqDvW/y
2IMn7sW5RwFa2OMYI/+2ReV0uIsMpW1QQPcPiu/mTegksQ8ujAuVvGmfgT14TJZS8Tjjo60Ljast
RKSMg3llDLtSanwSZTywlEfuJy5bco3o96Ry2bDsJXYA/X5Haj93RCnYkKdM3xlD2LRoKw6956R4
o8y5rnU41wyhEKzqTSb1xb4p38v5dQNCebsuYWSXdAN+dzWtTimimzAV9jUWRly+oPzZOVvceJSp
qW7qZDuZcOVtTh4DlllJ65b5qHV6FxwZI7TWRd51a6KutAvyCCpQQqpWH1Mf9Buu3kfGE1Bpld36
4mJCs75Fn8+RfhT1zjquBGkwa8OVO+a6EL+abEmgPbGWJX6CB9vSC11P/YPZperfRUpRXSBjGjCR
pULnRbkeaaVIgij/uHH4hJKkMHBiHne94svzVVMPMBLg4wWVQtIKQGmPthNnXXEwQazjjcSILH7c
xZOzAI607mvjoGhrvWh5M8Zmb5tAfE2io1HIlY3pufIAw0BbxWYu+NjuCHtrALSj7zk9BrvQYqL1
pvIVafUGNcmcF6kCyq67PyIVJbCd706LbFyrGCVtiYxAHuwJrRZkfBlOOLNTUYv6tUDXPkDeeB/P
m7qvcpRCGahsRqOUXRF0/jdLrTTqB3XRq1wu0rAPavjQsd1xMa7h0an6/eetChakAV6EUHXlgoQd
Sy1og9Ni+Y51wypEpIfxGqpyMvJxZZiFj/QKDM+8rMMrT6/d6DShSY3Sphv6OUfxVo1tHlQI141d
8tyUVT83fxqyqoUhFhze20/yVLb9rSVqTQ51ZZRImQKN2K9OZjyfaFzl3glu/uWqkDbye7ALf0BQ
xPpWC3kTYjjkLjZR+iJnE5KKj//t53G0lMFSKxuwJVT2UNbIbQqemKwygIx+7wtGa8qJSwccx+Pr
0fnUDWrFtKP13UqFaP3vBJt8XSWe7pAURHPZQOTORBWUu7O46RIOyU//lbE5CDHJSZtXA3yjLibl
bhscpI9DxFmQpHygyu/w0supfFXz4uUjN+we6F3RDP1GVtW5ldp1H3rpVrj1ASfsZqYgNdf+Id8G
7MZuA+IHnPLH8b47Yj7vcAsNY1dB9CCId5jd/Q7iZ+6cudMI/fAJfP7AOiNwqA1SE4VPVvYj094b
NKuz14kLdFS894IQY0Uh7x4GmM7DIMCr74YYHtPxuFSl8xkoeQjYMIQx92FPs4hHQbiP2bRuTzVR
/CriDIgvxFUNQP39i5hg9mphtL8E6lItq6bC94OtkLqO0er7ajruzJWDiBhFB0CdsNhd9A7S3mB1
AwJzkPsKljlIxCXSMdEf+BrgCkGHH+97twq8zvDL3rjgknX49mG8J3AcU1eBJn3Z8fLW8saSpOOQ
XXjuvG3RfHYa3+lxxOOsNK8C7xSk1dc3NoMmKWUbEY0mHKQ0x16w0JsyWoZ39FQ6LC/lWWjwCxGJ
9X49xHgb85qTgRaudIlj0pNOBXXZITOE8t1I6ArITahkyN1JcMXGUUhnpjkzngsZMcZQcrfrEGb0
B3x58DPQ+cuEWMBig24QWQ728UA+oKGTlpBKtXUtkh+NCqcxwsAMBZsOe/dZH43eZbonzwzBOnHS
tC5XFQ6B/n1jeD9fnzxtrWkQlLljpIR7KzLYJP9GApGH3PYEnDmhyL+QC72wEIxAZso4aeAO067v
FzSymkSxjDbvpR/t+in9RUZu63AECpy1bMeH7l+RtJxFjJa6T4UGTj1yy4Bl1MqrjkJ4E77/xcOx
ZVhyw54f2Vr3SaY6l4xQbUySYBj7fVepFQDn6I00TQ2DD4BNFqATju9+zFClaVVYu9rqM6OJO+gE
deX23K+nTLCktOasl13+vik9u/BH61YOhowbnKyvv64rNN5rPbCy/DAkFZ0FI/z/KNCXfCKzuBzn
rHv8JkKMisH3oUPbwiGtUTBc1/DA00m/JARGOzgZbDxnp009RsXwjZrWWgR5ZvIT7C1aeRTxOHak
CCw2ucafQZ8wMM7JoC8qXtXxA69rek32bXOeY5dMrghmIEyfXhWxM2V7FXoPuZcWS9fjNlXLoAU8
byymANXahm2cmq3hvVKE0N80eybWCt+5KxhIe1bMTaUgUODTkxJLQ+UVOAsSJ9myFXqQ5LGt8K07
XgMiTPDvt8Cowi4ACWF8dASCtzPs/r5OOllT5p2xY4MPaWD/je/ZL9WacHXi72K2p+WLCoXyrFI+
efvJQfXL0BZmdfWN+bSDHciTza/M5hJUGgqsNdEAnonz2ebkrrz1WS6uo09LrnsWuZ5yn3t/4aWf
JuVA4h5N4I61/QY/jUAxsvyHL0GjdkS07peaCW2dw/3vyYstQRYDXuWTk0hW0zvbS3vkRVGI+40E
bKDoeRI33LFRC02yhfegZwydREfh5APDPDFIKo1npHTKMV8XqDC3IO+G9iUPrRB613EiKj5EiVtR
i+sCZjGr58AhxGmZRJeAfv7q8kxH5I9jyWguIo2CwZqTApopswHRjw0D5+dUZNKkiKj1KhU527i4
YHlsaVnPsLHCIPv5tj3Unh0/wr0lrDm1S07rHevgSH804JS5dM6kOZruSFkRv8PM8htR+hX7P/yy
6lQG4dF933nsnRMiNvrmNo6wfqfOsqb1aQsB3B97ellRKGkKVSQNWgCjyqN8QOaRVH3jBiJhBbJz
Cyl9Ed2J/SMwDEITqcBXxY/iBgE9xr01yVsdU8KwSuy5ei+4zOFfkSRS1Q2o/UaxJde8m0qDe9xB
e3yG9iAigmkETU4SCMsZQHub5HN8X9ln2GGSaz6Bl2QT1IDgbmLGTwPT69lQyQqjlroY8GiYVtis
IM/caaETeCfrjjSZJiPrDa2mgGBWdfZdMdnzreXVLHIRrz4J2kel+nlRwQmTjdrXn73rAyc3SDhJ
SeZzN7YTeBibdMPD4vJmYWElHKfie3enUfoYR74HHkh09NlU+fLlWBzZ8azeFrlOzeHSMVx2vh7R
BSP1VKUX4IHpOGZW9TFJH7ykLonCuaNGI4Fv2NAxkol+y7v1/9jufvPk6zNenWfQdqdaVXou/ZqK
QOiLSj+K9ZNRkDSP3FueSR2YrWUjO9uqa4gcyXYQ1U1u0PCcwQKCsQDz1y6PqX0039vCZpIYH77/
yVkdQn1pcQVbD5HKc/2ZGfmLKJ234QJM3P+0UbYl99TMNzmzrkUf2RIM9IigR4h/s9pH6zFlVAiD
qz34N3biN5i4XFf9QxaXDb9JEPi/lHFfxlxW6r6BlSo3SsU4hiGbP3lb3Q5bvIKFTQx+B7l6CccJ
DvaA0EZjpzWJn5WU/2OW/gfQP0dmxIa8NcW+Lvaba7RN3fz32BsxImLNCgiNCe+GF/RM7zD9bc5p
vylO5h/okNYVeXv8bdkz0CLYavrr1aqA78KJbm8ahaoAyn8vLYCKXoj+SyiZVLWHHEjIx9RMouZ+
qKp8/HyBGpdmLlSzeVzpk72lZycFrH7BNE5oS0f8DtCvMOmMmnELH0O8yIjSkjqOEs4OFZeXA22r
PiK0q0la/xKUOooneLqBKEW6Ea12KHufk1akLErV5TW0s0114Ye9FgG8J227XhwXH7QRY8KwbNcg
LgIKjysJbtwxKP0Yca5ErzaWmflTNFoHDond3dOZnpPbRjk1hXNly1pfhgOqibBcV/Oq2E3GzAOX
DTCO3G+MUW2BqpoDc3r1ysx2KTNSaHHTghFkIP7uM9Gq3YLQH5jZUaTFBSCzlK0xGXLMaUQTwa0A
IFABVWatFEIsMjbx3w2lUebsfPGzER6MY3SXI3RYUH5IH7jggRvPLNBYg1IVhnO5OTM63fLDh0tI
fnB2tQzht2pF+0kPvk53EKJ0+P+l8n6rVFiqYpQkyf8an8bfRt0C430u+V/oRTDIppb8oTYT2iPh
BtEtyGsVzY5bKT5/ny2a0B82aD15DGX/FnsCktY/gcFYKSRVewwc8dioiAGX73dKpjwx3yhSsikw
2quMbUhv2UGauCfGK+0UlWQ+oy0ishVtC6Tnn8x3qbud214jWF1ToXliT8v7gcWhu/KHOFfOEFF4
kEQFannDwXo1xgmC95d4OyoFe5SuTePmtSbNH1LiT64Y4aS0izHmtm3dVVRvtGbnKroI9rX70zVJ
5/SoU9NKtH/Wq8nURo6liGeliBYH4xDufPxLDp1cHxziCD2E9ZD74f8M3WK8QhTQCeWN/ti0gCiW
ZIxu8Og/d29gT9BOHnmGICakpw4sf2fHsXZrSpGDxOmtXxEvDcwm6EpFtcVJ3+Fmv1ID8Ia+j0nX
8uqaTk36+MjifAf15MM9CWnrtFkx0rCuRub2V22DEkAoSI8UnI62MHL1cb1q0WUFDvrrhD6fToeQ
rxAzG3ZHyeuheGZCuv2/zp253okiPiqV4ozxZ4HUqH2QKU8Fkn4L19N8z8u/ye49tXJ8IXdu9Nlz
BtA/Hzwn1rQCYvJ+ax0cqeP2L+Pgp0CWFMRsrHTr4GdHSbB/TsVwwhRs7c+DLUBK/37FbZHxCT4F
u/0zrj7fPY9U954osW0P1+QQPm3+xGYaxxPkNhDVIhoMVfjLlR+9FfcURLphRSvjeCICB9PgZhM/
0TuqCtu67/I4QelSeMfv6HEFre4p96Viyfx0Z0AkOU1wtR428nrTV4P9NhByyInkGgRGUlv0vlzs
Buu1qoI+vzTseVUi9hJ4lM0kOae6KC9J21NeKV7kUnqNYXFoodEtXYDLOETOli+GeykSK1lsYLzo
BQwpUOwVLCSPaDp7NVf+XpuUUXOWvcrUHnmOGWVZIf03B7neflH+/BSbiXmpdTlcvVvR4Vi0P4dp
AWN7rVaBSUXgnN09Kn+MbQR8sIGxIuYHGD7HELJyixb160F1PGYJLr8Kzs4ZtyyTPx8/D2Advg2m
m0X6/J3h3Hzt0Ba5DSS7NL+MxBkKXcNkzp4ua0j1SrWHImswf22OlDD/B6Vl69n0pvyckfW1BAvf
E+xGp8RABK0w1ZusOCzaU5BIX9cy61MKsiV+v6yutW/9ByMBXp1QG5ZPxjExfaqOmFirX72grwuN
t2wbDfNIBK67OVu+8ovZk5QkvLZJj/2hRO5C7/sbAbKbBhP0i5vt8pj9K7xMjTzfJssRtRSV4EC8
0OK8lS9F6byQjVjYKYxgiSPhVS7snPV5c5yyb65hA1w/s/le4Tgz3oZx5sJqHGvgx+eOAfqNxam1
oLRg3p7YIKq5QYnOKbf6Fl7b38WbDmB+a85AqjZI7KXkpmYzoWdWSrm4orHXLFJZSx5sovMCKu45
vS7o+82iOGN9E9XDOHXTltQQnubpG8deih4GQGVL8vsODHLZGn5YhUHJEp7ueusgvPZR7Tf2Xoga
ZpUgCP1aodWtFR5momPRWxU3M1YDFKW6s9kuxb/bfBpltR6ufEzeRgYplGA6kbAN39rbQQuW+KnP
z55IMme50sscwM+o7/f+2vn9OxSMzbLHlZuuiK02uvzka5Qrw4Al6cxTf1wT5RTFlQgwhpXP+z8s
i19eRSUE8pNvABQpHcNP/kQwsn1JkTcgxO8siWxT8Sa96T/fkZijVBXrwtZL9d59e8Xi7wJZAngn
LdwZdoiwnFG0l5ZHCMkBQJAYWpF5Flrkt7bshJlZWEj7zSql/GJjpkcxO33xZwRYuBRiedD0bRmG
rTJS72Zn5Ouc+3UUCteNwVIFigiyMCQ/5NkIjMq2dE2WO607LTwwXbkzFZuDvLLYSOPd8NF6GroF
NXyxBWdOgnL0YFC7nOoPhX+tvuUjDYLQ7KxSUAR4lExaN+2XAfGqBAKrA/b+QMnsjhKWqpeuUlnb
WYhooMNayqw82cx2W+cJjMoAw6BEhPviuVKwj6O7K2SnEU8+Bhaq7tibvXggSUmdpfk8whBVZyPj
eDqXmZpHzTbRufeJN68URjz2OnsRRg5cZZO0fhAdTZPvoU2u1FfM8koehV6kDHMojL/5tNEXtgvl
F4mO/KPMoqLT/axmiJ3ExpN8/YpKAKIPGjLKXKMYeTYYlC5AQCOa8Fh2nONFg8L3IkCW79zP4x6g
rlunXjLPrjCjHBz7blN3FtvxOjwkBiR1sFkyn+vgep58mCb/kAwIb7rwVvbSDCQu7T6aNrIciMfu
jmNJ7K/aDsTu5D6hxkiCkHIBBsnhhwdnJjzqfCapBSdyDjddqOg+sHlNFZ4rafYP8c72pQrGfz2T
/hc4/lmYVNhthJmFTmY+hhksSflj81heKfxKxsiN3mUH3z2bfiiE1g6YnriiT5m5qpdT987Go2sV
0dO3izajsKwltIvlybSJLBOYWeu6EgrYoYQi1qDYcRP8vUOs8koTLOSI/VoPKongH+XdHy3dR6Ln
s/4HGDtVRYyLEzHZypGg6i7S9ESgU0PNLmZyVXBjti1J0Qu/DkQhPLUHQ48cnQNmoIRPUZpCXZRl
ydAwuXsdWf6WqsB1LrY4tObbRcrugmy+GWWqt/jPWfWLCQ3qaMndjn3oy+ebG/H4+IjkkdTQ2STh
8UfKBeM0ysAEd+WI8xD18x4Z4sTu4Colce5foDc+QK2RguvZukBe/Ki0o1Y2RerU3+4txsch8AcE
bFiwq1RDH2wjL/uPz4sa+bfs85Gr7EXB6xdFKS21ULlh3FnaHn0yKS42Kbvyk7TkJOePpGKRsbnZ
XrBhb5+2NWyC7uaTWNXSQdkBLWbA0BntBTRapRdg0Hn3N7nHGaoUia96uvKJVghhB+g+GLR4igte
BXyTxyiR/t7g3/LaJT9e51UVX/zhaCQ247Y6TzFf8tabOELr5xy0GEtXlXq2Yb2xaWA+iuhCxwJV
kChupmP3ftNvQCdTPGcLy9yajvUPfCAEMKVKv93SABP//iu7a0o/9HodbJTrF81dK/VobBwb8bBf
Y2Uv7pazEE30wqUXrvHObyYwDlFwN/s62TtoaC2wUSxjTw7eP0f1XvKixeP2c2wWZCXjM5hyxHOM
TpG+L31EFwoQ0HIKEvslfwrUYMt7MyN9sifygXmKF5SlCvOXKgsANjHA2LyR+884y7yDvmVc4GaP
X/CLNiGCt7YBBXx1I1Scl5TDGDsVbcZMwTOGPX3MhRuek5ydw/9jVpCWSfdhyjMmrUjTFghig6os
Shd/y3EnOtrbJBOgOew/xMA+qLFU0XIT2OTo0ItEevS/rUbK7+qfiyXMWMDucCrcJ01zfvnTeeTg
wK6dxf+N5aHEddyqDWqRorxtTyJKv+FkUmmvq+EWDaqSK4wN3Ck1FfzpJHyA+H25P09BbQbD8mEW
XbQhuLQNew1WoGKV1srKy69It52BO0gDlXtygVfwyCmUWclp4onZIiiTXkj/fLAesuIC9ZVE6Vmu
7Fns8mjK94kttPsrkTrGehikrsFERBGCsp1crsJGh8ePwrlNlakOwPGSIZaaUeooxSP7jXNDgy6q
P7nI5nKKb06VGgNJM4MOfpaubGH/zNaGLjPaN73gUBkan4XuoqJjy6zkrASQqu6UuHuxGX0iTGpm
bB5wo9X/qQr4d4EEV9hd2mD2FwwZQ/Y6KvqAXymlT32wLIyZ2tF3DT2E/ECHuLeJj8k7BOCOclE+
Tsj+VmxSWDb2LC4Il2ME4D6XidGwpRyC3YxU+pP8qJsCpq0tYb2NLblpZDed6sPS0xYT1VFOVQjq
H+Mmbwj148iyn/z+WcDfdSkrKPZ5Z1SYX3UQ8usAPv/5rKWq5vaJtfBK8/OVrTUo19oP9i8/xQQI
dIAJlNHhVh6NHySB0pY1YR+pEU7KUABfFD9QfGy8yzWbKmD4EF3tseLdfrVrh33HYw/chKKV7737
X8kCt44hMDQXl0SZYzVzqOBLKN+bC3zvrSXBTcKJeRXyI0Bhg6X5NsFQmwAi8/ZWUpS9PYxbeY7s
HLZHn/FoMqcRbcmpCxRSF62anMbqF46e8/beiJkh2FdXo5SgUszcJvM7CGbNA+60EV/80pR4kRBj
i22Me/KiruTPMq/bnOUpmkFGYdDD9IFltHGLDxH1+YS+cKd7g7R8fKqozuwnu5UNOps/WF6KD676
iuf2841QhRKBJJ9h6wR2rabDtlrjnYdzDXLJUcSLrIo6u5xRJMRRP4Hy7R4PX7dxKuAtEb2UhpPC
bImENkY48SlAKkryMUZBh7YEv9j2A/kqkQBvyNPS7X/vhpIqDFrqS06SiNaj3KeWWXkG0AHIW2ad
EBPSM61oDbEKLWn3WhQB0wSpzIiStQROQsqB+U35f5HMRe6ln1Ej9wl/gHj1Fjsc4IKnAMdkJ1pt
ezMYVVfTJOMjvaanIYigHoNz3liuPcWUfV6ayyyPZWWa6RL75k7cSJxqstpCuPmqP8yqwL+/34Z/
sCbUUoaROaSS5/007gptxPfWDNq0zX7U8+ADE75m6ZGl2insBBfFta9Fz4fzAQDhaptMjS1cPOAO
aifxAzomv9RJaA6lb2XpCB73IS4fAiOaw1GwMbu1LrdvSQwKWUhdhgAiWlJ4322UH7UQeVkdb6df
3n0KJjGxLotZUws88XKLb2G0Rgsn6ujgutp6FQZGKDQiVX19+VXEAnECDnuDS4PRKlM9wiCC9ZK5
qqDQep3pL4R3q8kGcsBP4k6ltMObJJDw251VGHFZbLsfmwZhtWNbjeL9mX4IH701rS6D7n2PjlaN
BnQHC1bXu2MoVjwMQNnjrZt1yCuUlWWTDThfJrhiWrduBGQNzKrwc/NGkOvt5VrVDuw1Wmyx0X1w
rQH9pIOmgnvGJI7YkE0gE4b1HErI2eBKpvAKeEe3jwNAPo8a6KE2Q1FIFipIHf4Ls/Cvy3g4FCAi
I9mp9imjgstPWkGjd3nm3qxFBRYuJXqPEwglg3esoakcatU4mfmDJ59HwY/QJTv7ZHmF8HF/7NzG
fEQ8crQeVFV2w2TXo5blR7lcLOBR5msrrEEwytaFj5R7IFm2rVQj1tVPGnjokXxWYKz4J0AuuDWj
OtjTc88mvdm+NbRlBJW1RqhlocyodzRKk2THtaaCWSXCPXzlkeiLdmxCadeagDCNWmPY0If0lmaR
RS3nzbOgWx/4PW4bkkuT4IFGjf5Cm9IVemwJCB7ZysRqNdYVdjOdxltm+7GonRP8URHAT0/QNai/
9rJTwI9KGqJZ+FW+VejIxoY183fdyyLKMIU/PNvwwtUq+5LZB9M2ey1SrV2wgCcnHqkZfqYOzXfa
eavmCUsMAQgija6Vkm9zgQU1mpwDAq1giePnzjYPTPPrWCKVRpPl5oIST6gylB3ceurOJffeiEUQ
/CpcI2Xs/GjRgt4lNypVvhjPUspBuIyr8i/Omru4UXqGabaUZdScysvtWLxpm6IJZgcUg3YbGVon
V6IdfTsSRCo2jEJlwjfULZoHO1AgTjkpRsXMFQtEvFGDSOuvbuFQkT5PR5fUwW5zhY2lizmQ53vf
Tl7Ua5Ceb9J6g5v869aPxCD25D0qgtpl4hJ6RJz7QMGwplG8EDceC/wTWoShqrOL4JEowfEYqm3y
zU87rzBvWr/yEDmhO8/GrGp5YLfryEp/jckTkUPfL+P/qRWbJyUT+oRxBdkDY6/fP+fg+AGAPOtM
5whx3NhFT6pHthfm9ZgkxsAgOr2oWhe+VNubnyBpWs85jzqYX41V1LTIrkw7zsPeR0j8OF9RBowz
vjr+1VggkHr8zEMenrWr2/X5VscNz3UrOmcEgEPmd1fVz8oZK24jdGAqLw1qUtQ5HbMzIOUK0grp
p2aynyMyPu2wNUCVN7IRpWv5Ww7XTjl0j99Q41l7jqH5QmvRG9dXApaKFYa7t9rbamXiTVSrAzSm
/HcJptjtuLs/jtg/xip/ZG/8L4DNqbIypu4pOVoUYQcXY9hHEm9jQkRSSldQoX1sArtWYwJoxGbl
lQoBege94NI45w45MzC+5zQcd2X1caX9y0aQ/M0j3yyYhWwMAmU0CPuyhbRUmSo9K5T/TCnIA7Oa
9DW3ewzZO2oUnBkKIeeuOTS2gbOULy0jB/xX1SvZo8OVb0BivmlKSnSgHYehxFpjCHQwkcIRyiAB
nMDx6vphmE7mcJf+vwh5YC7WL0pVMZAQc143f5njROmjzE6lo2fjsKPraF6Dqx17EWl9qq4kGpCZ
BfGrMlhwnsqltZcXz6NgwMD/5K/q4OX/hkpm7OF+YNq67tBWZUL6e3bQXNCncpOLblFdFqYJEF+S
7STB9idofQUU9JHbBvBb2O3aqvohEp36g/Yygi4uCt42fCAVFLHiW/G0CdjyLiqueG6Zl1c7KwyP
a4zItJxud3q+DRk7ekw7eS/pkK/aWw0baOrSSufzVqVIJTUG+2wb/m9DsitQ+xCJV/0yUSBM/Z+D
szhnqRJV3LAurg/8eDEa0KLDAd5IJ1P3GAuvUFQaLa64GcCweSD8yVU/Q9NdwhnMFvyPtl8h0c50
XkE2gsEsiqx2vuof/g54XHGflx0siFH3yvL22uH5xm4qUZ9/CxOA1c4VE/yBv4zWxZVQlj8cDZpj
yheXrxaWysFokhyN6bqNvtd3cutqp1OEOmpE3gHrn/4+pYy7UwEFk6xCTBuwmanABMLVkcB6p3uS
WQKwEj9EcKS9YawKY+wJfdvpRGhB/6E6pPV8WRVr9nKI5bfZkGqfoxh9OPHiDqu4syu0N7eKJduL
tI/GyA3VXWJ12OhNOpj7A4l2C90jf8MqmgGy+jhbGaVbc/0Cpcb0dAomSGXdXJBnyo1VUQi0dKHI
EdIOAKa6UQ+gPBw6CiP57tToB8v8rqj2yBsQpxYawhU3X3XT+5rtc187nxek93vK5Qj6vaQn2Fsz
D+vfimympziDGDF5fxKumCoC/t7U+lm8V8nF/aHoVSiCiJTaa/03/6pDSQRvqJvh7/Bp1LqL+Gvp
+NHWoc3MOWXUQxTPeuzRcSd9KpUFtuvvtL/accHRpTJuk7efv2wyq0RRv+QdSBq0CwJQbqBZEUDl
3P1zcqnvWz1DSIsQXXuC8ZaCKoZVzUyBf/+OVgFlgLrr/cJHYH/+n5bT2/7Of00nEhmG2b6tiUmi
W2KQbK1rUPevhQs1XWVqowUi7xr5w9oSDvJMgCS7UR4zBzpWEVvc+kwJQnB/kaxjtbL+mrcUumQ6
R9TnEuw+f1Ewfx8IRF5U0R6hzymrEAzJf9ROZpxzomQTYeuSOMnpZUzqmHcTn+Gs1CZxlloQawcG
67877zqD5MF03RG/XapRBkG7S93mxDnEKTVZU1Wl0cyUVFIpPPQABqh+4z74EYBu8MeBeaCkzLgY
tsTrXgBHzLQG2uEvRE4KE4eK48GRD9ukiCF6a2lb+flKQzlbwbFQBNwufNL3oHhB+iufoOKG43Z+
MjqYK0iazqwLda19VXkHT4XCp4OOGaNjOwpGTyfskfDJ5M9CfY6UzFO8jrjS0mCtbx80ymR1vBCI
UxfxV+e+X7hdY1IqWpCP0DhqJ32Y1KtQOfqhrovUFUDJbjK2dUy3KeON1oLM2IJ2HXcHKG/CMi4O
fpfrPzVZh5j+MM44rH2LkUv43FTU+TRK0rN9sX6u2lh5D1C4oX+69i6wJGDbqqNdHfKGxGHRmV+B
trlBV+fJJOQrY4z1kLPaCtC9Q/XifogmAv00ThP+BI5UUdGFLjri0O/vO7eoP3xqd69MbdPLLhEf
Zd3DD4tF1SuI49/bc2Ev/nxuscQ/m5dnP2L0ksuCzOxrl3Ry4Q5iCWT8eHJi5lKog414I8A7w0rb
q8qbVgpdIxTmqniS2jOOK2+FmfTQiX3ngVcT1Fk163lhSQWiGdB2IrQ20Wek3BpWn57ualuVP6cO
OV2Os8fRwyK0IKYodbN5Sa/Efd5e3IYu9SsJEKAoC1hR023ZEUcJzPW7IDEZvC+no7HLK2N13Wfe
3czkXLCTRolKJ8pfUz9prpCPMvjZnskX9oQ+OGhwSbJ39Qk/BeuUXMrpaMKYISJBoMazVLfSVL/v
VFNTkeSc4Yqwexb/V9EJLjKytOTpjjHPoR1oQr+hOTEqmOIUalWvD03OVK5wNi8yAP12CEDylnKB
nG0fEQOslgvWESOLCVlAxFaW4mb7xQOW2Q5DRutJYQlkJZDSjprXN5NzDiJwbiac5lhznwcDjQjR
3OCAG2RVjfzsTVJSI1Bfu+msfgthnC3bWmVhcvRp8D53ELQBzHLEyjdSMFdVht5lPAmXmxXLu9XW
LjgUFEE2SAIOfX04X4JFX4I/frOZBwA7FqYb4+8HSv1hJNRy764WAxNagmwI+Q3w4vf7jgApjlyr
q26uQazqVyU24dkLHzE8kacmnS3ho8pV7QQasP+96Vws6QKAerLp793rETlOiPgHtTuoAZoPE9uE
WMy5xDyqYQWw7QHXqE41XDHP1GOgaH/IJftBWoQOMo3x/7L6X3jLW+eHHKFeLgBdtDcu2ePrmN4w
VPZldCl4EvT228cz2KIb2tXsvtTjIXN52Xk4g1Y0bOxE0H9zAnfeJ4y9ydHLZpZRsYnelKh4X3vC
O3xHBRGSXOxooUnWwCvRBuVWVVZzb21UlP3jf7uvjQvtgvMks/P0p1iuE4bIzAHskameudfKf8M+
So8SmRC/q2o90aO4TVJSJUWluPn47dMPr0+1xkw8A/+WIZuFn4pRU9fKchyMyzzWhVbVlFvwi5W5
ky13xDHh99xSWsG0njLU1EDhzbdUXhXVHysdr0N7FuthHKrM2lAOhqLaz5OfFkGYO023n475EaXL
Iyc1igTG6bbwlEO/KTGvzR4ihCyg06vgxPTS4BM+vOZ4oSSnCphTIpmKzKSd5T2GB0RWU7lePRqa
GdB8vALfDQScA86J9DNdc2qoJRo75djoMdBNMhUr3sIet62WYbp8MALYISbQm0A/Zh+R1ijC2dDM
wBb0LtxbYU3q8PZCLB/fnTSgzipL6dDGspUPXxAGm+zeKmQp2kLSmWqkGvPusZb1F9fUz0Ym6JWQ
XCwL8e+6/PuKX3i3FQH87NnQPLqCM78w/SeNMF4gqN30e7mEJJPnhhs3XBTJaVoZ0qZ3FSnhg4G4
1jwsNELL9m3Zq/E4tGQlrctsJGLiOY5cspgb3EG4bnbIZkU2vNWBgWyvL4ihjSo+J9ytzqa2HWwW
q/PvNuwxuvxBHIsLl3bx/RZbfzI05GaOnTrC75QohBy44dVFTsSkfagkYAsNeyx+VULa/wJ+oX/J
2F7zDt1DEDF6YnKuzmjcdB5Sle9te6nNTI3EAEE63RJMUJQJ//3W8NUkJx3kAHRR/j+xD7XVaIrR
GMPEhovAnl8AZcB7FMoAFXaVZTYHHePoG4lihD/tQt98nfDxXVL1fp8hHppIEsnQCbGTWpyyKARO
TGK+LVrpE41g+SOZTx9BZqVv2iZAD7uVE8Zi2s92FfaKF3VX7T2S7ta/cW+iNDlL0h3zLZgQOw+L
H1f+GkQwH0ubG2bg0W83voBUfkXYqIBbz7qrlu3Hzal/aRCW7csGhyCo0mH1u19eP3hcvumkhcsZ
uL26X6KRG1y88LwEpQD/NKIaJors1zk2yTT1CUUq+n7zCRYvAn6/tukmrpKMfdAWW4OqAUi2+dRh
RVS+oNAHJ04cPApyiX3/UNxpKrINW246F+ZeKgWSGSSHkijD4prWqk1UEkUt2V0G37mDGTNjhjsn
WOHMLJY/P9V/KvM68SvfL4hWNYT8621cwMf15oFFt48GMuLosz5CuELQnDKdm77O+4D1ujJb0Q45
hGYg8pQvapq7HuEHXBtnjlXMcAEFP0BKsl4gSdH+hmYqvq5ikPFQuYRziJVWveLiBaFXcZWn9rdZ
w7xT4M8E6zIYIh/oDTCnP1nz9cOs6+0zQpLbeX9BDwxt98hoJ+tJRdN6mkxhuH+CHdJaxI4WRwAH
4r0HpEqHORzJ0/uceBMFFGru7IIATxZbMSFGewIKu1T0oHz+zkBtAEqGdutRX3pJTabg6T1lv6z8
L3CLCaTP41xERhYq9s3j3VHCkK76x0spWbFIClycf8ggjmQgR5loNJ7CpuzR6MRIeCqc1LfG3H37
G0mfD09HndK6soZdyuuL/E4DAYoR9ocYi6X0u1+8jUkkbIhNRIofl/dd4X9irvAVmjsq4pGFa8d8
JEbH9Ga0liVYyiWR6ohjXithWXJSHsWAbuKLmqo3ybnyvnxyoAIoKApYQgb6CQcuK9c7TsN3Q4jg
VxII7TMqzBJohDnVcQl1Mh4sybn7Qv+HFeYXn6ukjYrqdVyqLmVE8MdxDeLanEi93fYlrH2963PT
v4nODA+WtA87RZyNe6lZb0NI3WURR2WlWVfsfa4tNF5neI5KVOCsMGRxJS6IpMHjvwyWttaZapjd
GAIjmhf87ys6C4MUQJdg/cJk2nyRLpF4rqRQfiLjEdJWSxD+t6e9D+axmjOz4J+xXZx4VE2Ywxpf
9yhkROogPh45SujHt5mBJ4eO77agwtUV/gbIx23KUhcyMFh8bBp42Kv289hZReEpNyK6ZSFw1Ecw
tKzQf5wvoUN/vBqF25TPLpPBG7Rb6HmM9PIGqCedmEt5jo/MfuadfqJDzXLBCD3ad57hljx3cfIz
p3Vk/+Gdg5x0NKpO0dbhkEVSs5b74U5SdFdL4j0xDUW+WvbQ0VzMRplRdf9kxnGJhRDp+S/RN5ps
sOIrSqfFPVB63/kUTFxRpAG56u/gHl8Uk1tbwtvLCZ6UIkeZ196m/DhaWolEkG1prfcuA7PziqkP
tmA7f+X0TfUWD1yl46mt5wr5w4JDW5I3tQhtK3sR+lKDs2y2k9RFOuqFMiJ7xwkN8rfsqo4B2tx0
TFeVDUKXC8HXFugyxPzv/GTxP/7v+8Slq8TMJDjo9vjJVq1zvuSJWNBh0CXjuNhW7sUwOpiJbBbS
S/7oGvf8YGzu5TCN3qTBn5LGJb9dD3Jhv2dDZ/UcWodz7kuLGVNE6FG98FFzRsfphQUxV9qytfG+
WV0XE9JZjep5oqVHPaAJm6fK05vnR4SClvzTpM2H5gSrsXRqyAQNJQ4Lx/7TPNLv0UxztkxvEFlp
TSi4N7N07XJncPfyyJ6uTZylcCzSGe7VdSAFaI6yFXWQtLsr8h1Xw3c+9qieIxGUFHzp3E7MkDlq
laHvlcj20TafNf8QRcCbFKC0hUIkqzRHmF1AuTmqAP9/rLa1+OEWH6bzpbPaqbAOxTSRpCM/r0EX
upc1ucgfi2Mmk4iP3S0fEobt1v55A1s44jBLqOd9cbFRinsoj02eoJB0DiQb9GP+X6YzD9My75jA
MUGpKgF22uDscx5q5VThWsZIRO6nEZvTLrawS6NjGi1r7ADZYhKSCelnujwjM68feVjt+HgLRAGU
/S10slCTXnhltWrHw2ybzIye27prVlST7M5wLX0fwOvZQ6GBgQJZxl1l8+ToOIM6w1NbMmATp6MS
cpL5BrACz+s21oP465llQPf77R0uJPaZZxHijcnZfOsC5g9Y51FQP+dx2Mf5dgZdOSVPScXdF4Xl
MtfeJC+x19gQw1c+vOeD7WGfrJt3V/B5t2gWk/WdAPDj0PoSwRHNNQfzqsLzhVckBMtyJk0lVy+o
KZ9vcSPDHCEda2ReNxi5THlVR+NiG6vsKiyAFEHJyq06A2uKYRt4DHqSWZm/3IwaCKntW5vOmsp6
B9ldbvYi12s40+eBv4yVSo/LebgOYLG0nKVHDGVqKgv9X5YA55UEYYb2yxKRxsOEUcLQlAWYlRY3
F4C/c5kWBZRUJ3hNCbQPt2X3UybipEyj7ziAb1VYiTqREpFu8futLqhciudWWtwgstVj3a4k/bXx
FaZyp14YkuwdJKNFIT+C1AkvFJ2YwVXVN7dMggP4De+ty7E8HyekeDhvy/jayji5GvtICEEbsgmO
JSAx9sFF1xIasmhML/g/YxcKft+ZfcOW7leZffu+gNI/voBx14BU25XSn0hviiR/4G8+25LB6VlS
1oc5ea37LI6xWkrH2SVnl4GBmcManTRuWiQjmrtmWuP1G0n7ZFEvCz7jwL45Hzy7nsHSgvtgLMZW
O/vTTYPZjwaUoQ3tpZVvuwugpgdKtSDxCjq1RJ2sjUoETuvMhIAMRyKXZr1945Cv5K5F7WSvnnqY
Viz1GwGRiDVMN2FS7aLNVEXlFXrjLm1gyDYbhi78Df48fZ2wYpY0QkjljJBeF+wvsI/aaPWRH6Hc
ihylbEaMOLuLl/Ukaovzv1oqFPlT9F10p5ipDVJE4GQMhFwpJw63yQfjRvLqhkVEpaX/kKAgSbWg
zQ2Rs+2bGhEcTElw+DCkaE7O9Zdy7njsqZHNjy1cKfyMXyBnMJz10kxMzc1V0bLY/zmnLe1btJ7b
TyzXJZrAUvdjswbPP+L/lHsqivbAP69dKoA8nf7f5KLMuSPl8kwvD1VNSXS8gMi5U6mqROY5dWiz
Fo/kBKTHDHI/SsMvALr0+w4xH7cwLo4qydjEy2TxdmPLFqIdCqUmTCsEjhfza5aerQVjWt3CWqxX
GxZxw0iow1UNyHZL0vuJkjRjiU8+1txmMhU2UmWdXOv+nv7PQWjDZnJbLoe+GVYOyNpk2I5PMDXh
xkpXfK3xjRW2G9I2qQ5gdOd0pTa+LntnCjLNG15FFwr3eSdGyG7HALVE/aVoTxxiYhmSf3QMKKuS
L+78KOl2tfSyN7B/JaZgQ8FUW3ymP5uM7KCbnDOnNZKNQXAuk/QJe6ZqJgH5m8EQMR6HJ5Tx0io8
77iAgANGh3Nj1iJeANscQhNMIXF41x0ItQSaWHEFiYNMP7w5rgl2Ypj0ftrTgxhzU5DC6c13+tEy
UwF+lr3YqXBFoCE0JvYy0xAIFhejJwOS4BClb7HaapNBZSEceuOjEMCRoZ8/dbNashcOtLFd2d8h
qCNOoG7GP6LdpWeMIXk2AsgyIjGf9BBf0RaiuLJompGBN0nWYdFb3aP5M3/ZHIIJUNS3YNNduDmA
3ErKYqUQbHugdOQpFvQK+8VEtVuquDQRUDiR9LjOtwR5+TzO3i0M4+zNGJvxol5dXzjFmNI44cbc
vm4c/FZpFKJRAkAKhsTJwAPThgP/AtjR6PgW++1qWGGw8KpJUz4oc5AeNiufshac+edyAkGWMY1n
Xp6fAoAXFzi/4Y10+Lh74hMhJOFPV5lcZEjW5k2Zyhm+kmQWRTPUXN7WOhRORqFIEybknasEuNfF
Fd+bytAiCK1+gFYa9wDs2ZM92ff9I+ZzxN6pqUrUq4BGZgqYfPd9nsi3N7SF/1+bf6THt6bGgCOh
pwpucmnuv11SxC8O89ob1J3E3BPkk+dDKhI6WnDUfgVVR+iCuucdXtuDSdW8izyAEqy17CuciFEX
oqzqo0Iur65udYxITCgXSSwdnXJrTgoFzK2F0uBc7KEBmxHPL+f31wgndcHzrayfmavdHu0yVgfQ
udn5QKgP81rEgHJGluiiupLmkWX0/NKrsyQNVCEIHuh0vLydNgiHJ03ue2jH6Uck0PM+5YwUB65H
laz223b7w7qcTQOxJsJNdA2dnupa3ZK3xFMFlRqGGG5JWNjAS12zCwP4Ea7O4G5xRy5OeluJ6UK/
saElpshRV4CYWxec0YQm3gYrGK9Gqwx3f9oZ8B15iVYvsYNZrsj/zgyYhm28baRfRRY/CRFLgz9g
OKlWwhezd7vRoAIE8pQjFH/eRogeS9DVnt04UC3Q4AWxU8f8aO7D1LQ5urj72GMP2u58IrOnCczQ
er+Xy6FgvJVz6JCEviGHFIcaZLcIz6jl6vHN9BhheHCpzKupmszavkYJ9SOwnNJRWh22MFUxWGzS
MqkgpwoUd7zSd16r9S09QRRKHBIwKKkNHMMhaKooVRBYyoI/oy3x3y/2Ofita9EiXuZduUmNMs4O
uwRK11n2VtjpVe81FPdt9GWjdbOCmNX/F7FwoqGRNXQqRj4+J8ZIeGzS3xUM5mLslUSy+EfVn03o
yHJOnQuVgOp7pEMhnmv+d5Nhy9wW8+FbMOBsv8Mkj5ATy27g4kiQmLAWd/cXdXfVI98m10aFIP3c
u1u1JAT+WA21ZdfFxL8Ai1EY8YiKUQVb+mhQvpLVnf7o+ijpUipJcowM65m26nZYn9tlTFw4hqlz
5F11ekF6Q5DbGycGsaOpSXc4kspyoi/SH+8EPrpmlEjhMcrismimMnzAFHhbUaqfzW78PujHV2lW
mcz6/ZS0VxAB+5WIgDfjqAEPrVNFKz5tNB49a7vZccbtDomjJ+hQhQiEYgMOZqBpiNZmWgFtZd7S
KNZCcXGZJXkphxff3L/forvdGwygDXL1wZdXv0tSeitjzkzN6P9/+y1UT/z7QLjXjdnJtRnQiqdn
VMwHhcc0q72YQb/PEmV8dHt96oF+wwAVpPjgqV7KAtVK9ZgcQjxE+pweznU5bcad4RVN/BnGaI/o
HB+hxVKQVd83op1ZFcIAdJAs6cwgsWX6enBKAOtO1PZJ6zoRaVRe+ulFg7qCRz8YjQk/mbodzOwj
dzs8N/J1Nm8aiK2zAybGNzklxd1tFB/pgNVaItFQHZ0Br/KPis5quSGEkXeAnp+uYQBnWiYuEhXN
wJ0ISOq73uQNsiFpuDaSawFxfXfXKyUmRBBotW+Z86MT83u3gpxEuor3/V/qKZKtXbwqj9zvRTV9
4wawZHZuXWQSklsjzrScdxqqo8PBgJVXlTgED/BmOtY3C6pJ+Ncobxh3if2MXlpCiHF88HOAiFdw
qe562po/vbRGLwHZ5fyt/1qS5AwgcrVdLsThdLbY6aKTHhFT7FZs7wML9FNltkm9sfFLOOQJ5Brn
uGFDtxTnCFQZ2CyyVzVEZTBoqChmu3esjJ43Mu5XXxvp1fOn4eEnSYllS9ygwlnjXfC1StMKLzsE
DYECv3yTYRG2ghul7yQtrmQNlo22+5RMg95dI4CyviMJd9GcV18AlDQjwTqfdJE96ZRSM1/R0lBJ
eP/Lri8x2L3AM2mitnjMzRDbxmW30hhDCOTXu7z8hc0t+sKw+nInRk/h4+nOD/Jc6QgXJ2dYJMXd
ZZiUYSVUSQO9/loA7OzOlYdnTknWQNqbWV+LzP4DWIx/DmmsLAG/7Md3ZxUQGWMbJ626X3kq0R7J
R4CDVoPsGQPMCHLFCUANbELZe/AD+RBD+s1SLRmcMrGFUrodoOJHKvUuTCYunYrMctUgBH1SP4Yi
7EDNbaMe9cN9NpHka1moVS8wcZN/xetM5H0J3fW+di2EqWYFU5riiDaNPCiFCeqPB9iD1ncd1XuI
pH365CUe2FHP1aF2UNDVAYXYzaNpx1RkIQdNpHHXAACbTDgLXJiSeEmQC/6FGQ0s6lCEAvLZwDD6
Pq7TAwLKq+5jhtdx47G8+teN16+E2OQ466n3YqC1l6RpgL6Nq9C0GRUVAv3ke6/euHL8VK43BlZs
NMEvH1dIASZFYNh646x6wWpjbbc91bHltIgbeSOYyrqempEjvE0lbaquyrIH7z7WGjcki0Zn4WSH
17W+Vvd5rXop/B3m2IDsGLaWb+0SRB+G/XdwGX1oOwdKdTH0ni0vh+r2uuMndkNCEjKbFbTDgsp5
3pLiQJTAmsEGcEK5CUoKW27XTM12he+sEBQETlKtKybhSkAsQNNEbQTm8kM9EsLwGER92IwTc0Xs
eBp6zpGzpJ3W6mNZNojCN/mCa2OgMAEompTBn1uWq8/bZJR5AktxaXviVry2PWdT6lwn5lP+cQSn
S21R7BMlwAC/a3/0R8EH1GrOeGTTieKY+aVZ5PsbYy4MBZ0vqeuzPihE8FYQwGOzDr8BX6x/Snn3
HlvrGXMx3RSwcbPGMtW0oSK37sbTuORYeoTd4QTgx3gDOtp2yalhuFeCB+FHIlcrdZc2goFvFNH5
8h/3o6xfQBAYbkOYKL9Zbu4aYpxkltVJ5pmZpauWNQh25aoAKiyHJ1oiUX8rXKr/EvhcuN9xHl0L
jecl6yp/qv7AU6i7sF9nq8weXED3fLsIpxpHsQMyHJ1ac/80t5oJdNkykDDQUHeRMY7ya/NpwWX+
z70yJY2wtQzdIpKwj+0MzACRG4PU9EUWSXq5tr4LN+Rhm3PjmJhkQw/GbOCj5K4yYqjiKtwStoYv
7KFjRW9+R/ui4hseyeWVI0oivfvtbhtwkK8TjWt8ftOrtSvNQtrtB+rlQMOEr9lCuwkr85mhXj+R
DdaZLu1TkpSX47p5DCZjrDrDrtUXHwz5CQML1ifCMO8eMMlLFd7y2fwXDGqTeduEF3z8wizRaA2d
qrdqHTIYiRTqDEQr3TQxwGwrfurExoH5Rq+/5abVV8/GyudPeHqGkGWl+QrUkSkVnSWJ3j9H6Bug
wqjXEtjIZe0Se0402ab+tS6zxsAX+IBVhAgSsYNsWE4VHnVZR6s30NqHPc0wqbD946BUepF2WtDM
OaLfJjDiYQx414dJaFZxv16hudDl+lC/W/dotUXZDlVp7lpJ1Aeam/fIJiYZTfXp8bdS4WFDlMX6
/w+A7z1bu68PvdsTR2ePpPwVKO3b83XSkCfe6uXiKkJU9iXqiOBmznjvMNOq0DA4RVnf3ny6Jf7g
RdDqJeRdr3fMmq5TWdQ7WTJMnzHpkgtU0o+DU9rdjdcbgh4WJD8kn4X1AyM9JCoa2zBmTpic06Fj
UaqejpXL03iBbqM6kpUp4MMKikoGfYraJb4IDgToH0suKNiorzQDwVlDf4Y7iieOwNqamTDQMymj
fGUBcEt61U+ldFDw/1NdInhxSK+hDvNcg+b8zbxrwWJAWwwSfAp9GTCocuQymqMkpri/cX1V8W+T
A7xXhYks1R7bf5ZrY6MsCIp8mL+hswOF9sR8bePO/DIV0a2tA5v2rTtw9+R/509Paw5w9/2Wwj1c
zN09xUP3leOWq1fjwBFlaGHtP1nQGoreiOw6nv7aWu0AOLGRl+bKzcB5pq7yAJPDSojW6v+bQfJL
yk+ILOhDkrEKwoN9SmR9Sl3KsM8si7qxNM6gSt2RTwyC2B/1ENWa7OH8xm64WBVLX8VVtXfzhRQB
iFyCJ1mfcEJHYMbEAH6QJkxNLEChl3UW8t5eScyDZO8OCeSYXNjLh/5CDWqYvc4sgGXf2+fEAb0B
CSwJNRkc+IRxZJ78snSY73jkBR82g0WA+6e45W2M0Rw6t/BR9BlT3sGI6N5LcFmbdVu0Q0AYvrX7
0unK+d2U8pWfonGIPBKVynhdROdDSU8mvE/mdjxNh8luiyF5lw4NrYOcL+lTD1Gu0RlsuCnBlRd+
h4VgkV3tnZzyKXqCiF42VcAzTTe/xi1Ck6iyFBIijDZ5KCTvQKQ9jQP3vo9Vp5NLczA211baFnmF
ksMjtFArYW0EHLbjfyUV7MnTFZNZDvM4Fqe4l1NfmqwMzoyxXQQCqQA+R54sDkLhsUKAXUiLUzfK
B3Hfxzh05JgPfsoz4A1nMdxFOeZWAmmjw8ERLngpt8Fx4LMVWZzAAQaDSgvpvE/jtn/ULonxFPRd
bKuL/v4BpYoRiC8S4cUhqKdiUmznhQ23tht0Hot93Y++hcHrKt8RmWB5OxsQ3BkTZkXkjfT/bwcD
D3Yd66A8JJIKAYKtRNbK0IT7NE+IhFvKpWaYftaC7ROg4ZI06OirMFz9lQPFgi+a2shjtKXgMd5y
eoCV+XCdrQMeuxA/8j0RrotX1uMAGPLSFfSAjH3ImAAm8XCY1EDDDfJ9HytJFcueJRVXgEgvcyW5
XcKY8+tvGwi+1CmaWtZ/eQTn3JFBVfZXVw5ETFWDIoTsiecvJ3p4wwZeeZNZ+Xzu2MBR9jcxY6qO
EA58KZ5cJyooKy2cLFcjw6EiITk+8JI/Uv01/QsDQ42taqQhyoBLjiVErJJXk2h16FCgGo5/rDmW
iyCwEP70sfZT/oU115ZCW+mcZk7Jw24SaVAQwDTKOF830gtiDO2kUpa+UKB+eY6i7pmQzy3E6OdC
QOobzVYAzR92IHuofOEK8cxt9pOWx1aLQ1+Pi6+GDPhR8IqhsTAq6Yo5237fJaEfsEeTFM/KS3jB
Wl9GI0w7z/b0ddtE74d2uX+3AYapVvVmyLmhbmZHIIHQKs3yQcJ//ntCsLOM7VmcmIBme4H8h5I4
633x5x0iMq2HZi8xMkcU7aCtK4xIJiZEQQXhdBj9I7dPVAoBtTuVG0c7IhkZdPEtgzEl51xqo7co
vAlO5bmtU72aQ3P/vGxZABTxjF0ZjWekcI45v4XbdkBxFtRnDN5OpZF9kRxSRWGzP1MaCHrIf9Ib
cBrglHIqVvcCN77pG8hBT1kvLroPjq5bJwemP0jvXCoqcRrx9wabosSNdj9GS11SgdvVRuAeTZuk
ubND7tjqDnmJ8/tXPvTze5tuA2azKnpIV0f3z/KWnGn1tdq3iBql+AWzztGbCXCGdRhOT5nrMfaO
LhlRm9Y4kSMHEUEZ0KW8ie49Aww8CqvOLj/4JtMA9mLPDKiSaGWA7hiuaCpNNJDQWNio7cnPkizu
zbG4j+5tUmyW38y9lk3yjrKC5LCZdd1mKZi9Sm3RDH1/IVVF3jP54586MpuRsrxBqqFtiZUm8enV
fjU47f57pV4E4n0VdUPT1Fg5A6ic4D9Cx7pRYFaygjh3Zyy0IGe6iQCKED3AfA2Bx5T0UpW6e6Ly
4xsmZ0KRmorcZcQDEoNwOq5kS2TgzT/zGmB//gA92zakYpkT6m3I5bk6dm2VAWGEOAL8kA+mF0d7
0cLQBC2Ic+o4ByI5Bmb04qBSky7IH8cQI8whHRrro1Y75X5vpT5TZfrZUXx4k4l40M6qxKz631ss
1VQOAtu9hIBhZBEQ4e7kXFS9yShPXMzp5SEiCYf7O6fWpfO1nuNXk/2si+BQ7RZQZaoydB2oW6jr
LrF2BRU8xEIxw5z1G1mqVzNendPhFtxZoNstLKS42faxNfPbrFh7rA3pCJfPnEJ7jw3R1ohZ24K+
1JL+Eu65X/RzMdZ/I9DISwKZOLbRpRyrXnoQtgU1KUXUS7me0qfiyDTjbvmaPreUPh1RMgDHqnxS
eAE/XOtOhwUhtDrOZ/hjYo1EZgG2xQvv82Yg1uWBcL63rcEzQUXVfbk3T66ltoVj8VdoVnteztS0
er3WNWdzgpJypoeeHKCFswWMsJzDg1sfOiQLPwG75ucGPmLUcU/SI/09ck4QbwCbiLeH2Ut4q6Bz
2kZKvWk1vXWns0sMthOg6jVVb9ckAiL+cMXSI78VZd0SP7lEc3x+LmIb4lHGL193Rc6aTrx21/x0
mp0joTisvI4zXSWQ7+zBSTpIiekjOfkcHz3udB1BagKEo6ZorZMUvgCk9Dkk2yy2Of5RcNAPbrlx
2gXXLNmWKWUo9nb+PLBp4jeHAmqp294RbKpY6YNQKb4Emg7QBHyFKR/Zee8ul7+FLL0siqIHFP4C
SFPg+VuhSNOL+PZqnei1pIYS70aIx9Z/CpyUjcxUyAq8FSdKzfsjI6jzCCC9puQgq7lqyfy+IayQ
8p8sxGGoHAYwVDj55gwPZnTncpo23q7cvG8xzst0BE8GaiVRtg2Oiggv3D0nd5nW4AVePOe65hTE
xEUd/SfMcJYt6C5S8zcoc49NANQ3tvaE7MXUGOR32r3tek+0k7skxY521Cocngpl9Rz3zM+XmFZ0
6FCf5w7asrB3uaPNtQwJnBKPWGwGmdwbAdKI5PWoE1EZKbrZUsR1y+NTmicnesauqMZvkg29lbul
aMEL89FNdN6HdUKZQ5F+lKqf1i7I1VMFVcxlPOtGGDeBb2CJiB3sfUr9SQxuF5SoWY7hSaF9381A
lLfWtnweGyqRf4q5DQfVRVpPEJQeNB26Ckhk2jwmgzikp7OQSE7wCEUekzxgRErolCdNDA3y16dQ
gHOox7WWHj9lqkL1jUNNyuUM6OR1hyVZC0JhS4zdFOpb/r6cNGbTJASEJQRiHT1Ad00EXh/0uMtA
ZUGsOlbjzWh9ywKYsFzd+AS/iLszAZw+PtTi8msKp0ia6b2nlFZiVPq+UU5jCcq7FaCpfKn3ozsw
W8wbwUxrq82SyrUDrcxa+PTDlpJClZuI8/5Q5Ap5PHsGw5vEoKPVrMI5FnHNj0AxH2ilYkDxMq8K
XrlY60tFRC836fqdlM5mBzdEz+iFnOcfOCJHdanBUaM/j0acRahhwpKT7ufGMeCFN7qpD4U7aZwM
BnjX2Coh4rjsgc+BfjeRS3PvlVHL+oItZv/knBcGqz0+Ss18tmxaHqFQOOTT2IbdY3/wnyBpNDpW
gDhooc26fli48GIY26HxMC2peRIIkZVfTJKsIcc0Jp+FuqhAJ9syLDgTabPNc3I8k6xNGiW/Gjjb
z7+jQWiS1kGRed2SroXTq0xoedKIoT9encgjl9K+3k1xIdF0jvpsQSuBxTK8LE82zr09iEUeSPgc
FOadZQyKGC3h7xxzNpQ9/Yi0AsrpIZIDafLGWbhOc6JeFJQtSk5DtPU3C3griCNiSyBtV4fUo8S3
V49DyVTmUX2Qt72MgUYy2r6VhZHZFPTekVX8Xffgb63Y3TvAoAHDPkSkz99ArbsL3WqdHcITr4DQ
iRiCk6gXPXxLYpRQmBf6EQueAlWTPaFb52f9keg9K2iHW0kxlgqeNJCIwfKmbKu/3xwWxVMjjKIH
QvC28fNJ1xn+COHzQ8B2VmTYfZJMtnIj4J3PFVEHEwiA0Y3xSnorjlv2r6zGcZkg63xqhI/10D1Z
Hf/Ta5Z2BIOUIxwK2TScOyTeXC6FwMUKWwwX5rKw+aiui9AgWedct4RpZ8k8DfLqEocuBdmysdHF
dMjwIojvH8+oVOuM6zDWt2A7gd64aRfADvXLA2l7A30tUWIJyf5z7m+sLIXyqq1aDr7eMxo46+At
AE638JNWIyp2C/97dezYLbWSm+RwbM2fGQ3mMbYFBWSwBIMdZ8NxweY3Fltz0XArtFrxE+stE1HY
P2df219E+nR+CnW4AGzpTfPabNFYlN9SLOGOtgwLYOjhVeDD83FeH/pRaZvJPIRqu7Uv7Ib1WwrR
e0/rUS1xwryJ2WcEQjYaZC0f5E+NlaoR2IQhxauDKzzDrOSb2c3hr/1Xt+qIEI+4YwRES18eww5a
/rIorS7hODZAPa2aoqSgL9HkaDE+ZP1lek6BSthB4fyRwLnnfeDpDZpdcGMHfIHBKJMUEveg01gZ
93UiqG9nf6a3kFnRcp+rEfx9Gx8fuqqg6igkjpuNXRyEq2nMTC0BMOnfdFd4obM5Bu0HxtrMZxAv
G9eIst12mFfoxOCx6cf73vJgBCk9l3YRSHqfOj2QiqulNxVbO5q1PlPGSvj6pV11bTH64QIDUjP+
207FbmsEKda18CAH7jL1w44ooOCTEi5hcZzSz7N+WVoPn2ZA7GE6Bj/U/aimjihPPCsjCBNQCIne
Xa0VrTXsPvT1hIkTbo+2VAmRoQSLo1iCNB3lk9ndV5ODKRRoVjjJnZi0mNhOaFgEBw6WFfNU221U
Zf2xsk4xb+b/v4TSGhBszr3kF2lKmuA2KW4NcNQZstj1E+S+83WBIXSz3+LaVgVMsExIjn/vHVT2
0UL+dO6hRJT+F3fLeEZshPWiZKj96GIawUq8L2H3jSjfC4/MDOOu5bDQ6i6lzUONeQnsi++2SITs
4UX1r9CF/3Wg2r0RmaMB3NTfEmUDr8rIOCMmIfleBdTRPd/JkZENc3+VSukEh+un+8l+8CZn052e
epyly9UKnzu2l4DXNxJx1BSRE614XJ/i5yZze/1Yb/LBG8cLXUstJJNiuEkd0h1BYOtMJCapRhN2
oDguMdvpWJRZDXewZTNjgkIn1gsgPLwr2gPFt+7sVutZiAizgwhE8MxS+YRUfiRo3H0JihDGrJz9
HR0l69egagU4ABdGyIXvSLUPwYP+/nQ2ObFlrQTI2N/55JXW8dxJydY+IiuedXU8gSi8Mjf1wBwz
PMQuwg4JsGwEn18Pwm/eMQBR3Nmv4wNmstJgi30kmo90eeE9AZfPFYYPK5S+FbS36mZLW/rJoCbT
PKUnf2AnOTNmodTZ/IHybGCy/18QAlF6nrOmOzDU66G3/1QvFwRU8/lFOFjI6XRVGAPAmrbgNpEb
HPkYRWz5ujF264DiTiD+/U0efkvq2Fyn5vOeGrAmf0ZE5YYLhHZ3sqGX3ST8xtDqnLEvirte4l6L
MExmNdndXhIeY1XgXCTPzsWxEJYt95FGPRUKvbpWzbxvSs1cVsBxEenQFfbz4ZzUYi++S/QMQJ9Y
/lrgdoWv3B9vLTew0Cq4529bZC6aAKAIpWglQh6Mpy0i+9CtMhBKKs3pfhI98HfBQN/ml1qoPZfI
aU5PvR3ufl+O9WS8j0exOKcyHh/zVqfq6nVjib+JMSRDYKzQF4i4BoI4m3y0000pPUqaY8lbliVC
uGsPYGckw9D34ROfYE8wdQS2E47GaNxCsoGu8UmLQQlRdAn9e/CBaQWQR5KztSNEOaD49o+aFrEx
al6MVko3537lus2KEe78Byry+1KOxw/QFCKSjZNaU34KvlB6d48APgjRht1vCG+hpSyiwBbEkBrP
2Y3XchjtuGJx76541ehkpNe2A7Ps+u4DVMBKK+PUlsxbvm140Ewq2GWg4t/3aSau2qYMz0p9uml9
ldujIY9JYgkaWQ7+Die6/2u6QhyaWbdMTw8IbWlrPVtuTZbmA3Fyl3izJmlyhS5ZX8i9xR3BTDl7
EVzLZY/zRDuJa5fcMI+lUWw0MD3KfoL+C7jIEER1bw1071/OKfVboumlADM+6bg9K5RdDssWV9zp
iXYO7mlfmPQhS1YfaNTJkIigfO3FIasF+NRgFajLQJ1K5e0U2dusbiWNMBZ5lCJE73c2jXzI5p6a
j/FpcbroBbP4CswiYP1lJhkEXAHN7LH2uM5JkBJRN+xt3uX07tez8CgfBDM514RXJylUU8X5UUDy
xD4iJQMq9U2mkJiZVXepTT589RQb14S7J1QJ02D51+aKZPjlHgxf64tK7sPsOKxHWcmcyFFUbBGU
qU4nY9WG7yBBVCPnAjoZqFjkMQBRlKEBhuGaSE46yjM8W+GzZMmP+ZUQMtlCGr0wS1iFDqyGA9fl
wXC4fv8R7SIA4X32sYZDQuC1pBTe/3DSg78r5m7fdLZn1shv8SLPPf4fLf92/IQn3xhocRAa8yIf
LaJ7RQRXCUfVjvdoa9ibBciRAOEL/lrv65SrufYw4zllrZ03ucJk91G116lLfr2JzmVq/SHogBJs
QReDWsZoZmX/FmOySKlNk6BfA71w53LAkP8uwtAwTuk78pibKGuzeyJ5f+J6JAK5tKDamUU6Auun
JPVQ874KCvSEczBFR7y0zkuMaCnzmsO2wyRntCrpRxao6ZWsmD547FLLCE7i9vmewCWf7jD0wuRn
AD8hr7YrTSZTm+ipYatFJpY5Ra0lNOUVdGEvTtQKnSrTVplmnX8cor9ZmWFItmEqmvDqsndugen9
42cK50CKJ9U3Rq97G16TzXSwF8OKLYQsstj4blzq4dsFyvQIIQuqDK6uPhYNz5qYSPpqR8lZUjJy
bDxsxmwR0iOn43NU8TdaTj3sDz/+chHZofTD7ybntyQJ7xsvQJH8QR2WBIPNPod8Rb4tegsTvcOT
9uLW3GBi8UwNW799KR9HaH1zbt7rjcLGAZbk1HoBYVT5/Xu71AZ9MDnR/gmMKUD4bbQLDaDc2qwo
iI/P1KMYUGPClr4Z/2JDpL/XP61HTGvZn8f1rvgsomkCkAQCtK1ICw3mUFJ0Iqw7lQgYdT52g1Hn
2ZxBWb5Eovv6UpCbOK/LbKvprWmYps+hjvIIx3YWvrdI8yaEAPsm73TDrLp2bSY+8kHBjkna9w0B
1XJxD3iA/NYZW+9oY9ThpDW5hcW3DLQQknMhpsQf5+8nH35+fpDVJ+Af29AcPKyWpgNWJlk1I1yY
h4Odn16hw368EjqTfHeLxU2iLxFZc3doIJYvCp7Bct07L9eV7gWzM1fK3Q0T9ca6iZ/OILREpvs4
lRTTvJrl40zRTbQS5f97RzKUcar18PpBLK79Z/kWV7fPH37Rwdqm5Ot2ILp/ycQlq8Et8E2STIJl
0FwXpJfLXI/Z8I6poqjwxZbwZio+5qIfV8dfmp+d60MxI9CED46Ybe3SneG4YIZpfWWQSckQ4Pip
/srhrYBrJ3AWpkuDpkvxR+idtbm5xAqQzjpK6foz0V637//wEGulj+AqoKrSTWXiO5wKyqJACIOd
4CDjC4Vmjdzca8pfhl2VxVbkhi33N7r3VMlNjrDQP4G4nOdNdwUBMYHWNb/7CNAHfboGtjFpfO6Y
5qD3BuVU22aSd72zHJlSAeDYz7q5i+uckEDkpNQeIewBMu9pyw9L9QE1MZdt7xOkLzAlhftOu960
Yz85SgxWuL2+E5U6Dss5eHnX6M0WUNdWWErOVLnGHDAEIDHtlbqfXx5/aNl/0VOGm90574aly9ck
8N4FgNPMZL6odeD21cyCVMNsUpQ/Tss6N3s/lNxnwOUekJmZLUGKUqjuJ8UzrqymUSTMVzSSsaD4
Xa5Aetkq+Wg1kFcRXFxRwvrPDRZTRt5uhr8+tqQL8gslnRHmsDT8cHOtn19HoiOZwi/F9iThRdmR
3WEyuE8xg9QovCiGVCjijgsnZuSI3NdFTDQStRPLIG9FHjEzhaE/ApC0Fbt5Ugyqzx+kf/PPpoYi
OI2KGtBTY2G1vShYQ0CwAy7/Vh223f6w/iHdC/8l/7nEL2VOkafXXnFO75gJIJoS7R8805eaSBRm
HcXMYnhrzX1lJN6lVXIKIV2pDpZlizqhkqmuJuz+pvDtGYel5p+9I2ayV8BW31QyuOf6SVS1Vciq
MYKCXqD4YxryTWlgGKuNd7dVaS4bj9gftl/cJ+CawsgUEIEeTCpDZ501JxPopoRhWh6tXQ8Ezcf2
YXzcfwURZJFhctYxtWYJJBO++ERqle2tcr/fCdSfjIck1F1fsObEgIZO8PNotQ/HeOSekh0GeVQN
He5ubtfOJEEe7iKpCXGSA2nC7SUWOJoxbBPL0R5SPriLOiHifo6OtRFrmtDyTjM5VaBNIUfn18Pe
Y26R0u2RHLK2bzQMXAQHwOb40HjC27BJ0BdOBRl/W4aLQlsMHuohFSVYTvEL9XXJUH7C0cTxx4jF
O2M9lCte6hBFJhdiM6sHFCBxIay4OPtg2fYXHhg/XX6EZiWSs5uuTVBYAXPU37cldPgv5M4tmL1Y
gKWyNLsrDIb5SN3OLImg3KP+q1NEyVS4EpGHF0EF2xlVz9vL0eA0g3sksqOkoaNBBlos5uv/T+Zu
vhOdoXB2RCDpGYbOj46t04Ue5NH99jzRtgEBf9iq4/00xL7egz5W+Yox+H8dd5dKnQLtei8gzGku
QwxPp68xOMlQnhXrgbzFizpi/GWxJINwdNTbF5d6y9gRf1nBeMuVRKzGmGXILw5IXw+cuYJrlO4+
3GTJ/NCDvE6WewwoWSIPERwPWlB7MxgKYgZXgG7HyXqOUEYvv20gMJVhJrwX2qbOmdXZ5RU8EgWL
zFPjbLL0nj+iHjyFuL2RwP5FU7TmZF/xPG5d1AsgV1jU6nXI4/paKwQ6jKruGThAga8ukSrk3ojM
r4g09UtkxxjD14xuHPil9TOSp96+1aMwp+EqfXWm9FFIQo/YrbO2vR2TO1mtOeNkrR7akLJsZkDY
/DXRnzlsEQBC8hFloVAsQX3EhyEQE3XJRUKoLU3Iu2pVp8s3x8k6m1qksqoOY0fpcAML5uzpZtef
EJfX2tw2GM1atU3HrterK+UFTme3nXzoh/HmZckw+hn4jLnCQg/4//z15PKv20BPFw94JYNl6y+1
tgQU7DQpbjkq9AA4pI9sLSpVFXmVMnEZykQkXGuiebgV6l8Dv6lSicQgjbRYluNOz2/30BpubeWl
x/48wZBqWLzObAG1tP1D85PWiTc0YyPNfCZV6SG4kv4TzCg8XG+g495AOsYFHS1aLN8RWPzy8Stc
S3BJTS5jyvRQbqyXcXv3mUgjAl9P+IYSOHDyReHz+xUDehQQSNHO3xqkLhhBzqNht3wHhxv4l044
C26wn11EmRSEu4z3NJFhp377vdA9BhdVKe+WBGzyKcAlL4CX9OYTLOqPzLMJl+FHxbQRsBtJsqhv
NpfJY/SdBCo8Tx0kmXICDQbjnspV7S9A1++hD9UPFx0cbn+zFiBIsRpwF32LaOk7NChKb3LUYN5g
sA9iOZkGMuNpLwJOtmChoWBJ/r/Yh2W8wVXEXOlQ+NM+OQv9lGHLs0RjTxFUll61hf2y1JRdq96I
loc4svk9xrZ9YdEcIs82AqOnKYOUzLd76EBWv3p5hP8gPsUHEqaklf/X1a1y+ZSwOSIpfsDCsLiF
E8d+JAIvCgdkwXFdHY3JgoLsxQ8zO/PoUUgi9HMurcAhMp5QtogiRSzhnXP6ljs3TCOzfb/Xn6bt
HkGC1vxI8S/xj/KhdewyXNeqW0jieb5ZAnu8qa2g17UJMs9BwZQNbDcUMNfnRTU3M7RDvbwdXerb
XlxhYp3v89motWKEhYtmbzT0Uw+rAxmsOCay4llqD/l4h1qdWKvAowiPGip3PCu9LUwnh+1mJQ0P
WSeDNRYYJBFnC6tPnE+aQg57ndihq188oGMWDQuMgn4e+Z1rYEHFIK2XgNZzaYy5dKez8grM7Q8b
RrJoat6yI/ETKhRLe+WlEfZneBCRaZ99erhM+U0gsDvVmCRxKvxXG+XvQSgJ10VxbtSeh758vvTX
3XO2mZ9+SGLpPFvJMXHS0kxJrNCV2vz98emygVVo3KBJHEy/FyXhmuDyBoQXKSmHgj4cOeOK2hD1
bvyx1ZuAF9w5DdIzQ4QgKBr4crBpLsmQ2tx+ku2f5K6uLvE0S9quo1OTXwtE2cRw64Ay/KIEqhT4
s+oYLB5OwfAU+z3TcxltGgAjsaJGboEmmrxC+ktLPN2OJGEIqQ/hbZRrJIpwcHLep5QuxRIdr9jF
NtSXnBqVE4F/iHjvHwBk4L1pblRmUC0VRrA003IGM6ALyu1s3XwC9DkkVPqHtxaLSRRyiPKs/EEz
A9YXUhDrYnuID9try6LR5x1VCh0nOhiswNsY7OZbn3l2v64q0Y9UlZRpksec2Opxv/i+Q9G1oIc3
FJVXdjutczJbK7txiOCZU7e9UAKTy6leAYDYBVD5cF9rMMxevc1x1I/TPKfmFq+VhnyD370+gkGt
ty4eXigSaQjjdJ8cISVIxHme5Z4rEnxv9veNnahMze7Sg7zZCucX9PpnIFdB5MIgV038loO7Mj+T
0V8PgyPhPxnk9uc4yndzUoD6UGGKAM/Qfkkf01CCAhA8uy7CBxLJS+CUoLDnHLMqiReIljWK/lwi
CM4AJBfebuz/9s1IDoAmxugXao/z/qu/GS4HyOyegPanpeDUGur/3USG7mgdm515oA9JcM1uMGT3
xmktT8Rx9YkZs2orZb0HOmtdGPDzIBNJ+volYqsSOS9omnyrtpr8Vun9ro/AJAvPYu2gv8JCXxlT
WeOs5rsyaylC6COEjSOXVWhFBHlHs+YROK3STWMV2ZgJPe314Lx/8jfS/Z9NLKNPRDfRbQ5rhN26
6k6yeN6koQeo8wO+BgxmrqulRglnw5JW0i0cQh4ce4C4JfDvEqPYRf45rDSMBJPMWDeZSun8ELxx
Pzk/cFn8c2jvA7mEaJ26VG6HxzeRcD7S/eKWdpkkTUyYp5+YWf/dfsRMIsAiPbdu86XYrOL7+WT8
rPg4z59krXvbCndKPnS3p5doaYZA8F8ewMbVcALVXLmwxOaq06VkySmGo2UojxkgzpXZqkTwLbaf
lokPG0yF5JZeSLHyoR2NqNPw9DO9hFyrNrsGiYo/HMc4nuI/JjTV7uR6NCopigWLo0ruKTsqB+fB
MWkycp0ULqIML/o513UOyBrMC6yf97wHaVA4LQ2o8PRCsa0FLZsly4iu1pMB9NDKXUAl7L5p/T5p
FgiFuKJ7Vw+91zqihuuq00A+cMsAQrUgZiDUOnxgaRntU5K9T9sjkMhJjC8rz8FtQRDbrAH8K36a
aYdzk8ZIF01APuP1Wb5uyikwZxv533Tz5rvKTJXRQMk0X9vKASqE3jm5n+ANAdZU+Ll++VXfLPRn
mLE7J7laLFilXKABl7AbTNzbxs0qzHRvNe39LIbHOFIT0pS2Ou3LBamLJxHxj3nSTJL1IM0aRQ8N
rMc7fvTcvVCj8/p98s6uUThxXF2hMR3M55w6CKNNPcr4MS1QzkLcHU3elcebMPCmlsJMICO5WJSu
ZerIpA3TPE7IjTnrwc/U1wa41pJYkJ66wwCnn0gVgdi5cNmTS5JQ5YLiv9n+qE71S+R8FN16HzP5
CAcLjaQWHcMFP45QMLJqavjfC/W7OgF/W9TtKbcB1qY1CYVzw+0pi3Kh4Brei1nFuIWxjaUgAubC
U+NGwgbrujljpH8gzIGStrK85j4YJtAfceorTwMSGO8QBkgKMAyv1ozOGz83EKzsh/+svZ1oxp/h
ogZwnfd/9pFYqAD7YwPfG2af7ewhXgQMpd/qlfMn+Hby/AAEUzapN3U5lYGMYSddJdYXGP/ZdIQh
V2NzNdfy48KP8LbvY8sxb19ggXJtOLoBtxyC36qV1R732iDdRkKNtjulLIfTLfPiRQ6T/UtfP6j9
NkQKbPS7C6GRAg2ZKZs7nVxwrGeE/ktCwExv5smd4lGLNDnFEOG4DugUln7i/DrpdntfSUTkYcYW
u+totVNLjI81uvTza5QlnrkEczgATAV372t0mLFZRzHXI1+a+Lc1Wb7qBjhUIxcDvtghyXHgFB3s
VxSXzsCwAFp5lCZqir7Suv5n7kQT8Dg6Zl9ZU+CKJ3IigFLlDrnU7O1eP6AkHyOn3u7Atr28BbqY
4Y67C/pCqeKN+vO416maA7r7V/FAchXml1s7ljJJ8pGwnByS66MVn0jOZppONkjJ3/XXx8ENdsjw
2Iz5OplRHzzAzTO5CBPJS7Qd7epDBd/Z3hzokTsCiwuT7gCM9eXg4hp81YBnOJApl5IPFgeNcwWV
j9mcVcpOmVZW4CJMHo8htxohQ3Ofaf3R39pkMmDT2Xqd15zzXgnDaVM9G05vOOx6dk6ZA/jZLzGt
AyEWC0PgckuQ6+nGp2+FAnekipJCv7qYU3rS3U5BX2yGuD5DrN7HkYOxLqAjcPgK1o0tUdoAU3qu
ACPvTiQpMcMqSfbK/wreJHz149oPE5RL8ukmNckRUiHU1xJvZ3+UZmMVdHcQpGWksQNYciJ+wltY
Sf+fQg/l6FEW4qME6TqlHHDhsaTBvXWBNlu3EVDWWRzkzopptPzJa0tExj7L8QZ4UKM/iGiREGFT
ZLt1Wq4EA79a78r/+UZ8f5muYe8YmdwlnTXCMSn4xTkNQOeo7IbVcTG/9hBjg+xhflZVZJivJCLH
mviPGAPh4aMdC3JIbQtjfmbl77lYWRcQubkM98R+aOU7ZjYSSEh5wcSRjCkMmB1wbkNF90f7yG0f
COQy75ntLOjYYaJQGoUnWqFKLHSeOc9Brf5v0Qkj1U18kVq+YEnbV1KvFBiPOuDAyDdu1ojovaT7
ah/8rtmp6b9D2Sd0g4QwMSTphHGYLZscgLRHqXsbaLeC3JZyp7du+V2kOJ0p+oG3C0+PPWTDR9cM
N20/0G1MYz2MZzyiLGAG0AVnmcO/mEDLvQk87Jqmj7g7x043LJlvc2ZXUr1V+8FlVkSoMWvjc2iL
FbogknKtjIUtM3LJhSNbG4wHg990Fqbf+4qAW/wZJ9CvF8USpkitB29uL94XXee52hvCR0DzJFEF
pzPXd3IZLIf0NQFLgB7NU363g/tUGAw048L6c0/JkXxOIdtwTlFTKay5VdZOyytHQXEldX4MVhDx
rL1X5VtQAhl0HLliZ3IMcea4gQKUvX276ipInkCbVnVOQFkTgLCCxLRphstmR3p4hL0FQIwPGcvN
qWBJ3n2Sd04OE+gmT5EUeW051FkAjGefceTmYz/PPiEadns+q4PhpJYLqTv8i4/Yy7jYDqeVW4rM
9K4EeNjYtafxU/QL91VQ2CZEpMVh+S837KqNrUKNvI6CJDTbu9l7WPKsTuYwUSiocpw/hQV0haiO
B3Kz63i5Shxe/l+6odQnu7aTKuFWcP45Rd2U8thlcKzrxNgTmtgnNTCbbJ9g0GjWJPnCWdkXwqxX
9TKkn7uEbSQG68M052MvUX/13UO8mjWz2F2c/kds2J0Z3Vq0lVAP8pPD7goqSmrlj543gV2b7znd
ufl7kOrGdPRl605ojo/6d0XCdzqLqVj3sfU2jui35DGq0dF7raZM6m7Kiqp5Cu9ke3vLiZErhcsE
V2a4FjbVrFDQhXSCwwLr5Y1IEmqpJTqY6q1cGZkK9wuxC3Ee5j5YNizAPAQhlwytJ/jxvaZFH4xe
XILhBU+WDR2P6QiukbAW5uivx8dVrIrMDlEtJuxVDOyoNK4TINXWyNmTHGyeNd0e7PkBLxpjoA4t
824TTDvQi4WWAoWthS8yWzE5kyLAHRwVg2BlTmyomdLeR+Q7G/NBOFGncwyoLl6geXYqPYKzBYXI
fcY7bI+KWfdv3qVOhnY62pQkJI0gPFhr3/yLW4LV2mRTERIA+FFVW274bqktmPlGSryX2AmDkT3D
Fo0ls1dtPzX/upnY9B0HB25NVW6JScOF8BcCK+bXrEPVBmYopp+mPgZFt4NG8qPA6iGSTxE9o7gv
w6Cj7dJOlXwiFY9HnebxVaW0vwwE7Lejk2v+GVhM6pjPMh89Nh9MCkpYsfqkZl6bu4KtvsdB4Oag
d/RHlRzL/+dXkSyW+6Ja+j/+KBIs+UADcG73sGkjFB72wla7Q8JbPcmfvRS8RFvnQGCSBTXJVwhQ
zwHzD2uYngKNm/X4f3DnBiOzZS+fED2OJ0J4J8wyndG9msBNKEEu4iB8GG3Oq7s05JGubo0i3b1Y
6nP/Ln8utjAf3LYbXV8rSLnHTK5/4Tozid5iGnHOR8S3INbdQxkzJLPrRWViggTmBsN4vDDapupk
XgYGXIHH81us+ujMJ3YuPrMsbLLWAoDYSBAhRNbeFMHJDdr9BdMqvFkFhYm/KJAXBVk19o4XUlLR
Ax3ftMJzO9/MaFEO7FpB9bEiI3TIO+GgbINNEOKy2pHUzcLQHByTvw+ZM5gBZzr4buF7QJxJjmAT
JdEu5hHgUCB+bzg9/IgraTnHnEPK7ke+iGGLNktLqfy5AM5exB9SUZOc1F5IlGpEv20Mg1ZoE+UI
OiOkxAPH38UuPKhqpd8vSa/0pFV+xPd5m+6T8O5oQp4WrZbwJK1j4KQnTyMSFldiAk2DPCyeBFEU
1wentGZNLA+Q454JlcqxGJvbLppqk2jlgb35ZRxvGOi6qStbRmEcKNye4578ybSaFt6/RJ5RiuRH
uSI8Un8sivSZTWriEFf4GRPtVqBwH7y1tUVCVdd8G9MLmp4f4F7s6lj6ZnCa+ssvb/KgkeBiLwQ0
C3eUb60ncqaLdpUDtMkumCY8LRHTOnTklirIX8kw7x3j93PcOZbQSaDlEQXCT03Jb52IVlqNGgEL
um0O/M1a+1y3GF9qT/gRk2mhFvXqgdhhIiZ9BkBeWZTTljlys74ccOQJjU35EQiF4SxwQhUFFym5
sjMTCt773iy74CoAm+Y7yQEAqBqQLDh6Oy8l97KlBdlUADfwHz10khKvd7qobpU46tHXneyZuvnP
y1z+qY1RJIIRRlrt8K1QwCHYo5EI0qf2GKhY4Ebk8ukliHnDX66aEsUgywd+mfYrrWs041EoEOYo
bJkITrDD684o9leHBnGrwm8mYaIFufILKkSQY2AWzK0EqGHjwKS4a8dO0bbrhCnTmiSLUZuVcjaV
ptG6YDzX8CLZ6b3n51A+kLFH3RXC2qbflbM2WriyCJ/c78Q1lkrJT+H69rrtufsC3RiICetBZ08s
8nXOlN/JV6LJ/5QPsmvGTsrtxHf/b2t3kqhtd1kmJGHSSJ9oR4p+foGYlMJS7yYLj7C2ACZ1yfbl
im9uzgCknRXZlHv8lOzbfQpUbQBLy2shfPFDtESLdASPQvTy25gyjtUvVG88q+mHen+Saf+7ItuS
jB6YkAOA+cRIpVVCnhbazKnaJHWRonZsGmY4vSA1BCE6KIMFOjGEq/KTIlc06Q+rQJRVGq2ZXhDd
iq3ZhhEQDjAmr76U0I4vUBYF1AiTWHy8/wf11rqcKjFhGMbYaJVD4JnrVVnlP+lqe7DWeCRaPlCh
HAIIDg9p7TCPo2ijNwoowPMxBYF+zDj3ePXD9ypGB8BFyU5qeVT8YZCJT/gq1qasnw3lmpbbBH+I
Q0UfSySjcUiil+alFbsQcY3ayWvtEsxBGx3LmIO+VgYWbIKZIfd5CJFO2y7RKtTmJkV6LcJml6xY
uAPqnDhfd634uGnoXC6edGSz370HmZAg8r/VrG9P1Vn3tGBoIbCWWMRraOJk4tf96iM3sHFVJurx
9X25ck4EVgh4YwTIt9I69fATFV4LmfWD82ginBuGafI6+C/6rzPagQZZOwEmxz3GQJ1zuBjVIjPJ
8CmVKl/eHg3q4UDdggqZz3YzcCpqQt3P5jBz9B/RFAfIU1lM4eDj+q66q+W7TRNcpfW3naW8t/dD
tBYQgGmOoUG7EPo34pioEGDMaNlfpMMmVPGaioBhhgK/ZQGPIIt2/aEiCu/Fb9aqFcLP9wrBOE+E
H/CunYjzHQbY7K3BY78AAMwhKIPSDoNRQAfpFshE2X3OC/ZF0+iA9kHvOBV2rrliQc8o2IxvSRPr
t6Ql5VrJBx1hv+xwYLsdz1hO2VhtPhuLliZX13f5KPlw1unKPCPYjeMVmontrfWWfWsGlkgcN/gY
n4fgubTocYc6l0xwJoXDj2UryZjiD/G6FggjYnSdyBjJTozphkMF/MbLJwAabQok5jlhICGrRLDT
p9CvhProiWssgqcdazggqaQPz8ZEHa5otSMS+B4ORYDVfAL1zN8YBWQSBa4ImN+J2a8nW16w/t0f
vonUNkuYU2WIp7ftAA3iTG+FfqDx0wJWoXACeSsqz3eX1KlukTaD/EhbzLw/zlZBKVAUXNVu30UU
4+FSV9bx5e4Mb6FxP4pAoUgAFtfkEp8P49KIzSEmA3ncJduMO2jvYCwSuFD2EPTW2eTvPFC9Y+xg
zfB6JK3Mrt/A5YMw0V8p61gTYMyg+nT9Q28+Ec/ynN+zLPs9WkOAPC8Vds6KKGnSXkxwbqnBh68E
yGQx61RNGV01d4caD6s0ATW3DaUUHv/uwsEKFQRKWVN9nqzGWZcJvMi7UtnQEfh1wdW5mOq6nw+B
26c0FVVoIEmcAT+AEWSj/m5IAxddCciGAawk920yhGm16eqTNuvowaU6rHo2npsFrOZx/nzKqEZC
PN24MSOzkXYPWqbOeFDiaTaxZWziYQLx/RGZ9SMbISOEKz1XykdyErMuO5HjTgFpE+XKsGxPbkTx
BiSYn1bRiTG4WkaNRvwOFDS46FBY1TZ57omvz1262yY0MwNLizh3BHXit5CX6Uh+WCyvrQzfIrZV
mRVTLuJadbbp13yi5cOoKULyGp3knL/Gzpz8CyrklA1SwnUmVovtWhDJrIQVMQORVAIMxxq7oqWm
TJfEQNMvXN/srjvDw4mwL2drpEJKfDcz9SyCe5w8ya56dxTtDeiz+QsnvGn+Fr2FlMlL7gjtpoga
XuONxb7c2hopP8TfVpeYarzHASSh1ohAXOLarotuLSvhdwZ0GGq8dHAEAacjHDPAZKNYCoH+10up
xeZAR21S+g2S7P6pfJcXrmtor0GqneSXB/rMyEJ7rVZfSZYNUAx4Esgl+5UWr8ONjVrwEeaPCdDi
yAThRDyvPritNAMZInKawZkwIGORWykllhB+Uctvd80vR5JN2fklViDMb76Q1yscXoqfQ4d+00zS
G20Y+4hPTJ1XNWi1G2fzkKuxL9Qw08aHoL3eEJ+JBvneFOz6M3xoP1NYnIamsl7fsUs+53tbZKxW
5PCAL/Gh2ic9I9CwzTMJvzBeXvQd4IyMbEcbPdzdhRSjRaBAXo5vZa3fnH9xuK53OedIsohywN1e
x4FKYhh3i/OSM+c19CRanvFu8ZWR97aqwYYmis9aIm11lLEvHWeKzCU5Fk5oeSNPAC2td7tgQkyJ
rPJUX3iQ7cYs7TiZajxCcEzFD42CvY+opcRjJof5BL6FdH9RFiqrt4ftlE4Ti+KdrjBSmlVXNA/C
JLWOqlR9dp4cpwhD8DTSSr+jg1Obb/oR0OQt/wFgTTKhV0TRV0ROrejyxhNs9i6NMTVZpIb+uMfu
F46p8WU1xs761zWMonpcFjbbJK/lF2NGh9gCy7XHOde0ozR5VlzbWGXzxxRHPXMi415CauVPGhDW
9NdDaX+MIITaIJIuwx0BwEf9LSPdg28pAkGfXBiep111zM2BeHdqUSzlMesdqKrBg35ExQwdf3ed
lqiGUXPro8K3Zq/Xzf9uFFNpqd+y7Cs7cJNWWqDnRRE7F32zpDEipYsgJ1rWd2nnAQ4K3qt/w4VS
MG29CNbykRmEuIoMjoUQ575KL09KaCE01xT2/D51FJBFlieWdfFAdknb3DJSJYBlwzPIkISUAOlN
6pkXM+Z9TJsYraZhTxDDs9HDO5AfFljlTghkZWLVD3bll0hVEBtMES8DhnMHb8lBFpi5Ixpq0AQh
eoSejCU5EVubd4BuhmgtaximeC/4ZNE7XcrEkzVLgAlOK2OeCJ6OPlK3CDL0jfXVv5rG0Xe7oU5g
Uv8omsGJVQWkHSUGI31TbPwQu9wgC47G5TNhk5BHK9eUiDllnREBWRQFkelszAauo9rMjqDYidXF
way4ThA7974+QCysMKtJdVQjrxRwfg+8yiL4LSsbSvOux7W7zllNDlb97JT1B21hk62YO/RwxDSx
0NurDG80PEgo/XhdFW/65H54RzVEFp4ztmpHnLL8mZ24yYghHXm7ey9ooRdeS1DYAFXQKK3EaK97
O3pMAXkqws+B/hxIvq0NtAIK95UxLEBxOMVYfsM0+JvACG1cyRHvulKoj86N4j22w9nEPPT6daJM
XJXz2+4GdlQ8rPyjCR+2FFf/R2GXKGWCSCZGNgliZY+0xoLdCDZlVhPpJ/gi2KT1AZ14C+qV35n9
ce56fqovjRxlqmIO8yyZXBl2EpJRHvzRJX9zByHyPM3yYEXM4wJM+Ahd96G9MeI3t3IkLFmXptA3
FlFRiv0ioArgPrGkYjE2AOXi6hwKfVSjLpaMBbWnk7eBm6BAXzPPa+U4FiKmB1uPQG3BuCLaeSC2
9ohxjuXqkZNt0yQTdjO/5gjUGeCW/QMnQGyrReKrpx5n8cXN4XS5OOTCF75uEZWOCRjONGGTgWrr
1ozkEGAdy7AEEIKcm/7kOC3KZKMdWxlIKhCX2+PLhBJMNZoTCfeS5K7WYHekhHeoAX3vqw9hDiu5
kIXWLhpdvSwizi4MfsUn5aUmw1rZx2NIZYfdfw5pLy93EB5Rtwoidicf2G/ZSthPuR00/xXZ9huE
x6YY0nZINgbddXTiU/RlCSGH3g6MTD0Rdhxm7LPbxdg6U3qSUKA28g5Z38nrllKieMK9P9/HwEjx
uqWWvQ0y/R+7VbIFPOfXTm9x2JAhOpWAgAE+miEeHQ2d7BrS4EEOANki7NoVkvFN5DQi+5tjH2Fz
2IAJFte+tkiqEgb7zevtaChytc8M8Z+ofyDTNxlIdzhxASw79DE98zy1LZts8vjT2TVrmDlSeHBx
66iPRWlH1er9w6uZqe4i1Z962cQe3juvnxIL8nNlcBDI2Fef2BFcEjga+p9BiQ4EQNlGltNQ9pqn
oMYmPC6c2Vaih6CJwUzHHWMt9fHCgInTg1KBN+T6C7fgQ+wgHUXXEX9fvwX/TqZinOXkI/Sbyt7h
CtFHFNS4u5Nqe8MbriAvNTdheL4d9eCBNFbqnkZ25wQicU92sA9/bJsQ15Zd2Jhmey+GaCUBDOxr
G206Toml4KieSn0U8KxptUvk3usrJvauUXzchUwvI4z1zhhkIAO+fjZZwGAjAk53rfvNGSLns7Ff
qt1CcHMf6F5OfqDn6XIvCvOJ8TlSiWp1YvazBvBsjI5KMAxUM5r5qiI8fJBXgLRZ7+Reuyve+ufT
ldm/Ob2+wP9U3wACUIHwx92oFvY9OeSYDbXNu065HzuSI/fYJlMLdpM/8L1bY+xErS+jxcrF0ICV
TZD2Un+dIa6RbjsYsLaff3ZDshtoXi9EaYhyppPKVoW887bgMSiIEUgYfIrW8Zt0mojJwoFvgG3R
hyBaHpVAL5Bz4kSbwI4S2m0W7TqS8mWubaXtiXjGqccvZ+ZZ0CnEdNpMiNgmmPt9iKbWv7huTYUo
Ryj6YIYMyvIf2UH9amoJUcv6PhawDF0jsg+3af291srKxnoCO+kVW9nOeBEF8/9Shno6LHX4eUGl
YX0/yRbvCQzucCWLRpfQBuBSP0SVFd6DKIQ8esx1y0yuVX0CdwGktS4sRfnfiAXTIheSPXNOe/Mh
5IJZGNuzp4qblv3VIB0uJUdOLbIXKs6/M81+SZL0ZYNBriykFlpcRvkSCYhMx895XV9cOhZtE2Ob
IBqc6VL7da7GKK8aRmxPa+Gmb4BhmuUHxiviu6+0H+FAn8TAay9/Os0h3s8LsG63SLUMeuQ4WLK6
DPvfg8UiddBBhngKVL7+MdRYvMZpuA2cNqP05yXl8gEeMh/H2tyliHAVPM+u/Rixnq5g0vaoh0Qk
rx0RgK9jv6UTcqeKXm+Uqje+3q6QhjuPny8kaCSKEBMa2NZjRhd/Roh9LYm1s/friReyEVPFhHRk
KvB73XenUbdBVhWXAz5L5wVuSxqgy2XrItS4k7ePfJLzLH9gZyzIecUlkY9AAROFnKXG5DCBQHSB
4aXiNZn8Nx3t1qoumIZMvoX4rXkDY0TA95s4ICBBQ7yPYRUZOCfmhHHHckWP0+MrWt9MxBYCvz1N
ewprJ+Bqz4qyLFXXtW1VrFLimLO+JbWQgiQjnlCs1xcAxVLPq6BTYeVN4lOUe/HEMKiUD3ig/uyt
jD5l/ftxQgacMH7TNo/yfffFtaCTsDd2VUMg9C7OiTLxUtWG8SpJgwIQ8tJHKCrie+A617z5ijm9
qwQQYm/4dRLMDL77fHnvt90NQTv70F25hItXcYvSNFiz884X085s27JLzhixek1crGDQGF4w3HXg
LNixn0j08HD6kZkDfFlVbJBceHeLvMf2keWgPqCzrcr0AEEziO2NFWWtWpTcc9e0t8w3j7AImsVw
vMoFzQFxZQHn6GQksNOXBrHQ2iKkQGivGZsegoXYVLlZ7hk44eV6Lie8A+Hbp8p08Nqdr4vZYN1D
Uq/yISVPtsvkeNZXJj3YBq5XyfPGshJTMplUWQPdtGxLGB7WzIQ5tzm61xPQd7ATLXpJCsENx19M
ZfXBurJ5Hwr+4QrKz2r+CZgz0V5TzwrFhiHqjkZiYMl1P3wgBm9WmavP3PwoXv6sn4Ajdo027ebW
CCk0ejGTf8sYt2No62ygVcbxO5OWbvq1trLH1ZT2zVfJNooJog/gLsat42hE9EhaVEjtUqGX594s
mu6LMRPf+LbdFoW5wFC+TIFpBvwCPl4Edjw3/l6ZH+z+kByTTfNKba9NjFGHXDxtuy40kGOXkz0f
7PNr/q2/UB8+UkMhwnf6Y+hbwqqE62soRQ3HkSWx5XxQlm3M0M2r3f4/ENrxSt+QVd4yWEYk0g4C
o1s4168IjXuazYyfwLEuNt9nSQIpAAKgcyRuL3/UK1G+23cjrI+4R+n4fspJ4GP3w0YYU7GYCJJs
+Wa7MP3k0M8ZHRI1gLkHK2C6EZyl7aAUrXLSY0IomJW9O7X6Ax4FjEe3dx55WVIbFMVbMnF9N/GZ
meral5woR/JVJCXg6URgc2T3q7vEahamH45n/o4FzBRCc5+V/Nvz1XHYkDmNQVMeEALm0E+9pR6d
PzhLluu10oVbe+raj6rHeNKi+NqCoqBVFSd/pJAix0oLQZh578rSTyD0ooneIwBkHsodCYPZnjZw
KxHow2VI5oZXcBI1rVtE42xNn+fCHSQExcm4jwEfLx8SiuugsvVNZ0qe/aHzKBhLSeWOOlOz0N0M
Xzbm7qxAwMTRBHgPDQJqT7chvIivh7dTw/es/EkV5ICdnxV+9q4fpXv7hNerv7DPZFnc6+to1jZg
Zh5ttM1cXeoQEqlZ8gR23iz3F6JAb92wFO6ugzsAm68Tf+UtaN49iivfoQ/OSe1q1xKml6kUkNO4
ixg02VUiWl4JrBDyBNN2uXPRPx/wOXHrTRVaZWFk4OeWL2ykckhVkLUYDMArD5Cd+VxFsbqyVVrO
LKFPI7kXT4PyK/uKCY2JE02K2nsGFw739KNblh0eJsU4fMwwnHnwYw8m8R4rFYD6bwR5FDaCXfn0
O9YmHZ1/5IDUQjEI4AtbqWn1m6oDUatktbl8dbpbnIZ01u8SaZRBtsAm3Xl6S67bWvlvKK+0uIIx
qt9QAkyJ1UwKtLqa0rSg5YR6J9dlcB5SR70888r0zJznvrWq+oLO9+chxYrmUKyDSGdiRGFAQHQf
MsuIlea/kIugj+A1w+bgYukSYxTjXolljM57mHbdtD94aAUIZhW39g1a2Irn+W2gERbkvMFPP112
g4F9i3UFE3FVU5Lsi+kOL5+igR7o6J5t+v8Cbj0ktYzUNDMCZo4weK1fykQSbS+Ro8Mw1a+nCm3A
8fYyskWUZvvane9PVASierYZdbzSMHZPJJipXcEzquxxU1NBqotPw1Fain6RwYknWde8BDuCviSt
jbZ8gi1PkadU5kKniE5tVTqp2teQ5rRPgruxtAcDoRiL3pvxZTVJEX2MIh8eiaZnzc2LGLXG7GgE
M/13nlTMzf4lOWAkRzCHZLHmxvQzn7p9QSUIpmmE9XHBFZuCz0guB0TH3TznywdkBRszMB/odmtG
uOMe6x4Vo7MGg7+xx5Yda0PHpqHIyJI5vHattzU1PsNGKeEnU15sPif6sGCEzwBYOtfxIw/HMoiX
eZnmghBnrMezs7SZ0LzlYCdC6d7RlyR3EllloOEw2RpLlFMlb4XM+KnN2fWok5CZ41RqkJnGzzqq
emQ5H63OchOk19sgHXuFHMVmXnVOETI5IUA2IDpXhzjdJYKWf2PTgOMFeRzwRBxqUs8tFtXZN8gZ
RMPIeQks4ryopY66oU18/TFzpVjiPN9m6UsDoxTVW8w7+MXOhBnsTmMgL7PCWV41oL+SRWJgkQgZ
nuce2ngKuVOumXuTpsS5gUrn5Z8G58O69JGGMnO8TI5xmCvJMXkC6hPY7peE7LirZYK/YXOcPbjV
UPkmoY1tN05pYdcYZ87E2eAJ4grkRwmZmZLLVLYBPjnKyU2Aq1m5aA51+FmguG07lRHxSxzNEG14
4npKa+JUjYb6kPTY0CDjGM+qQLMZm5fc18LGEO9qE2bNWmKma45Jj8QPAS+2ez0CR24xHOlmoT7d
BIADvhAGUbvzqIks01BIcPNdfwwq2p8PizYMp84r9vB5Y0tBYo8kvTWq44m+NnhmkJKHDU8RNhkK
HwB/PIkyEG2ttY5GIFA+9fJktTTUgDc8+Vgi5J9eK3RvFAr/OWAeB6DKuYWCVZxHavPyXyPjcb5z
kLALvxAFPu8qaI2i2o+/ge7hjNMiB0HKGF16axS9cT6ky6Q0ds8XijRXYlIGAUR22p5jAk4xnr5p
9sd27uEmqldFQ4AG5YcwK6p2bZY56snLto89LxHDTK2DIS7T/l9hcF3S8YIWrvzGXn9sFxNBcOCH
3U4g7Tx/2QhzNzCCQv6esltkmOOg7gwDAFbiLplqXGaSvVCh/KaLSqvAI3gESrQ4vZI0Jpj1HKBj
nvRwQCbpnxGAA6/TBr/9uVV4llr6xetj6ZRIKl10t/AfJI3ZXQ87gTGK33d88CLPRv6zO3H8qSZv
rMG+E+sz1aazVQGty2efxTyZ2xTKagWZGyplYlIZRd5hiyYDC2mpvbmPBmD9/j+oX5aE5n/KP8bk
E2vRDj9scC6HXn5ZXlULN1+y3iGRG2CBGTOzm3zyPy23lsLamiVKPDhzt1ouMOG4BXQvxpF56bvc
vPE8x8tYyb4e76kGY5hJz/LDoBg4+JE1xsOn7B2mYH5jDyv3KRh2TDbyxLZ1p3MD3A9Ierf9ye4I
Q5OdCTDNrXUpwzkypDk40mA5rhG20RyizdZ0uEMbgLP7BBg/r7+YZTb+g6ig7GB7+aBe4Rekx5UA
0c7c+1jYX/05jxTGLuueoxVo/kmfceHI1A2WpV/y4SW0uYTa5wslQquEL1Y1uAW4iblDoaGbIi67
XTdSnu8uaRPbH32ZJ/jrRpn6AskB5HbV0ib1mJRld2lly1nn8T7+sGouKsq/+Ss8xfYhcZBgy09g
KiN3jEyqsG1v1/M0pDQ06fEB9d+6EaMn26VnUkj8+OIo2o06Lz4zTuO3bts+hc/u+AteLfdsshoE
w6uL9ym1urs0Hxm6HppqZfCitvhMYGir5aTqooYhAeTcQuGwEVwuXjI+NbNmlega/rv8pMg3DXRQ
uu4bzdg1J9/gWXJv2rrhwcASFqx5tNVq4nEbcIGE/Zqc9kZTOWTN5w8WfKjTVKJvksHj1ElrfS+u
1DSMfJRXKfUGwse+AkqbTdjhX1sD8HpJWggZcy2NipFpoobk4ZaVaTnDAytalCKJ5RocPjw2cQ5+
NC2Cj3mRNDeeWbv2rkFHAWH1iKwHS47rGdABsfU3Hw+A2hG54zm07sKv2rL8/33NHu8F7dSLzvVN
x7fMQc48bmukhw35y8HmKfmakO6Kx2cAOlh5csxnxS6JXqOJIeLyIGze11gC5USip0VYKic6y0Gt
iRrU0pWew68wamc4lHqQ05a6u9lCK89Zo4ATQKCquviJkb0FS3V9k7bVbPk5kBzD5wS7QYGcaL3G
r64nLypYgzy9z+8thWik0xnsWrA5N/as7uZpg143FNltxGPRkSKrhTwmWe/Dm5vn4hFUWFNFv+Bu
IE4zflmfSq67iqu0BOxLOB18H+qUoqaBg3Uya+oXD0C1LHbWc2NVBOmfZ+maWWb9ySaTh5zCgLx1
H45nHVyMKU+OcMmlFuPWQhx6a4tSIqRCWw5JojSEJbFcUM8an5kc2quGrqCfRmMxHtQDxmPQKmXz
9YTWMccrxaQGQdiGYAJcVKhc3VubNRxuO9FelpKBiFc6N0pt+psE1csulWzUo9myGuWgQ8HHv32l
CPlZ2JiyYjWsIg4x7doLFXrOtuBuLDC59GFVjhdSdThimFVgrOnD4LtQAItB+aCYHL6A8Tn+impE
S5niAtQFs85SyitRdLt5eSnx8BDS9x98ODNGIbghrVyr/7in6jtgpAURhjV/ANtY2wDej3XIDhWd
yZrTQOViyT3sCJhseOXZhN8OOxkxcxaXGVtwoY/azOh9RNqpfZtEyghtR4j1YsdqY43BSNMUsWn5
ts0OwrN9e4c2Q0xlz5GDztSBGcLoi6N+tW78HMxWBN/u7M018my91cNcd1AwztzrMzFcM15byLvg
RwX0bCZzPb7Ui+oMDEsEUo2DvkM9NWlGG60z616dimoZpDx3/6Y/pIjKgDbPCm/FNQqxv9eVV5j4
hLAzUAnNlY2gW8cNDv7Pz7qf9toL42OlNEQmNZZ2J0yp2DY/VufCVsMk2AgZleFpvrKPzqbA2GX0
s/j+skBSogMjK7PpVJ7gcT2ptgd1fbPuRX9413mKEjQeH4XKuK7/Q4iUy1SmY1z9BFEy9HKDhUc7
N9f6BZY4sIAJpIlB1C6F1R/Rxf0HecXjROOL4yhwfHSOpNKyHF9ialxDnOiT/9zTS7UoyuJt1t0X
184wtGRbbMmdhAKPgB5vYKqX9wr1si+NHlVmdeX+kP+KxOHQXFRwvkAIyN7Xnxb0zn728Ufl4t4g
pyRUIcUmK2p1mpQFGanxo4wPreOAQ8UGbd6oWAl3cXr7qR3ArhBhUGYnMsQv9jtpmG0u3HwdJ1ce
HC2T4z3pjgmFJI5Csqh5givdxfHEXkoz/VqCgEQa89Qv7jO/UFQVAmCGYnZd1gFBxlQyMxR9S69E
nTCmg/9FVr2parTlRTSQ+qtF6kGLjCRhhmKw6XkSzKzuz2mvUS+tFPG4Se3ebpHunZsX0qtDwafl
K15ZfBY2AO3LbrA+7ShBWuXBonjotjTA665v7+VPA9h/Y1Q7lgQ9bPbcYSYR/PCxZaASDvH3cU6U
Yag+9QONOLb2mIFXQma3BJmxy3PTT5CgFeQoC1kBgWcVZK1cjQMzxyzkLamQ8KBOk2Qlww9/rXoT
TFaqo7dOVrPAZG1LZeYNK5iwCvrDsjwNNMM1Rw1ys145l6XF87s0Ya3d4hFQG2ErUizPIUh6nfzH
Ru9mEgfFSU3xwEmcc6LAgNn2deSvbeQq2OlIWeYGzRAW4bjMlONzM2/M3+2JUUrMnQg5P/r0+oU7
O8K+x4qMeZDZXUkgDdB4Exglw8+lmkFaHfhyeVHY8L/p/JkG/TBSQxcBGxxPXkCkXgRPLvBU6So2
zZutqCEoBFv7rNH1TSPZS06lQzPXDTzIICpvatiksUo1e7c+HZB4Vj37gxZyYEL2OzzU4QsIJZXh
KBIGZTnWMB1wT1Mly55yVCVFxAQztzu+/8wA8t3C7qBitTZMguuZyt5FgoAkp7k36d13nQlPdX2b
+xbhmbtmc4MaTZ1zMpTCUQQ0gKjXIHMRco3iv46cb5LejsKyYet+lyz/O32l0iCxT6BiNWjaZ/Mk
UM6c9brDy7LGlZV8/O1JrDXTcL0C5e+acAY3A6SOie1Qv+MNxmcRPbN8oTZUJUYQOKioF6sQ9RIp
KlsVmoPIcse019jPa3uZB/0AZsdh8x7yiLwi7VriYicAVWSaAsSjQuxd/8jJze01ZCi7M3Pm5ZlP
dHyF73OgekphFRzLXibfrlrAuKxM3MsjZMebPp/fL9oM0Lp8wXUfX18NhdM4Weg07wKvfEQg0A1o
0IJBHUrYHX/idJvqyZaD658DrWTuVKOXSQThmZ8CJlb3h6N2eM0kOsQe+NK+8nhAgr2dkrDyqIxX
NRI9vye2dAKLNHZQU1bOqIX0WvTddVoHybOsUhHKWcfbESkKUswNeecGP1K/oTrKC6wl2/SyuwaI
qeNBsKeFdHm4m+mJX8NS6Qe2BixGgy3liTZsacqxcZZ7fJ8eO+Ghi2dHnCgQUHmZTl6ky2luCemP
rlqX1Bd0pMB2MOjQjnr/ikXMoHrEPEVkDBV8iAgF2CKGeS+Oy5CXLn1ilaIBTl1sclqjAgeaa+Hf
e5j0CfzYBvbcGs+NhZhGqFSD2QBhouke+T1zA91lYCsm0BCd86MYPcQ6XPCpZHT6M09+xDdTan1z
65TRKTBsKwkkNt+JOZeSkKhEu+nTzruGnHm8JspKy/8BKPI5x9BJ7LOwcI9OS+HIPdUfDCF4agwk
Wq9SoaLAyFsKqo6UMh9VQ7b5KoYvb9+a+Q/CNqQQIlOiGVqvuSBNcpyYlyt6L8ob/5UbnYRr3fHF
of5SGHhtIaXohYqMkI/7AkuuzWCTN8Qs0yu8jMIl6b5zhFuksd6rpKVPsqquYYW/ky8Ham9Zm+QW
H7YQcnKG8F4haR5UDbRMGhS3Srf3iq6KyScgLYw6cAvynWkG9SN/l6WjQaTEwpgEGqjz05MkcwtL
o+D/t0xxPQZFygBtKd5/WrJn8s1rpmSaaJFhCDqqecQw6Q9wChB1IFPHa784n27ZPg6zBNRaFjLr
Wqk3HNtzMOD+ogMmoUZnpv2Rj0/ZWqNXQivsgWos5fVATKVSQQOB75Sj1ZH5Ge9zJOXb44o/weTN
XFmC41/Z55XU9YH8IRmhk1iTFT+CnGmqLUOhlOvMSN4wBP6mA1Ef07a3Fk+t16uWIGV83yUFJ4Q6
NCR9QqKVhCPcU/Kqi4pi9iWMBzZyfxKjbbVQRYp/+twovc8nM1lZb4DyfM+BRuUmYGdaxezZHn7U
p5Qzp/b/MlW/jcG7GiavKbyUFDgg7QjtD/hDOnJAclU2RrWugOR6nc7j3qcj7AvnTO0lxwCPGtQr
S9O/JxZ+bUB6ywIKYPr+RMg1PVMyiFc2RmbEM3eudJ7rk254C44pwr1kl9CcuDyM3qMS234XWyLm
bMNHClnk5KpSTGXxMOpUCSzHVs3LQ3xitkJUS3Uqv/YtNlHGY5TZ5lnzNBvL48rL3nYequERlI+T
z8OjZdlIRpBIARD9OEuJhIGwkTyaYKwLby6hngejH7+X/ZGFOBdQBZUcxQs1449Y0dUtisUZrmwM
X7xR2DtjZsDZokj0phza/+DgfX5VVdbh0AFFpyo1rYzAkal+RnGTIjbTPx2h3DkU7rN+fmm23v91
uQOknuAgZPMNuFO5qLLtW1S3Kust8+C6w++7QtMni+RZSr9R8IjVop5RtGK8eXayvgYR65hTC1hI
XuaDxaDz+m91K+3hiCiqWOwqDL8Dn1HTKDvan+SrWQFr+dJ/4ReASTc2ve7zqOQTUI8H4RnrMcUD
N5xkTi6OThrhS+Og6tXDfcEvQT83gvJYHjZ5ix/aRKa/ohI2y3M2eD97qITk1giHxwCVGDCzrXtN
P+8ODQ0SjAC+1BFi1xSadi4H69JUJqlfMovs7si80cdNOaYYH6MEhvBBbxwJdwYJAJMntGqQyIpR
uE4UiqB88exUu6ocy01oNFgkr79LZCQA7EJtPTz88915hHed5pJMBbW8uJ35Hs5mFthgXqH6iPiJ
Ca5+KmBhgU3NjGOzMzNvQF0d1dmBRXu2FSyPCls2Xx/ZbmmzZ8TKruk+MM43CC3+yJUQjLwwLYLu
WqqfNBPkLDj7kqdU8r7ul1yXZz2REC/zpO9Mi9mWspIA8BIQ5R0pTC90I3y4rUiSiMqxNqS9KRwP
zVbpCXydf0IvQ/ldvMYNCRHmE1BoNPLfgp9g/gDsIgclAlQdj2T9O/bxn4kvTJQEqpqQFChKchLU
VkjicFu2P/UQR2Ktx13nBcDRzlQtnXZyG+nyRd6dbFMOYYKpQVlIC6OE3QnKIxtBcQsu9t6lf5Ae
VlV69Fk9LaLceZfQ4416K2QmNHXZqeCIjyUW0dGCqJNGD/C/2CtltVkQom5BPnQ6D5bBYJysAIF0
PSknA9UjTGKuA8tuzITjqhHGio0rd+UgfLeiVlSJ88FOVoR6nfsucXR1S2r26rPzgkZVLZd3nqhH
WNj9bi718WuiLkAcfUvl0fLq/5BQ3+yKRzXYn8BadKMhP1wRhEzFXNR3wQygOqxvd+WT1CEfEzT5
m82PUuHXCnvpand9vjoz6aySTa1d8tK/oV7xJtknS3oVNkYGsEQKQOSYlD/YLzBAaVAKTKe0xqGM
W/Cn9gDR8Tgy8LJ3nmkQpk7jAphxmbjrlLgfG6IwHPUzGLhCR+vxnbn/9PSxX0tIVq426b1p9jzY
WlkaaP57xlGrvGK/Xu4sZkOexHLFbiC1BAMJQ6R4abgNJ8GX4hsdWdl3ibH+uUAUbZkhT4ZJHjRr
bhlGp0NX3ytjOtTs9RcSl8fUHbozyJcnaakl1pNC/Bac87Dr3r4iBNcMrkp5FfGbg4CvCJwBuZ6q
mLy8cstrFkBJJdJ1FALYIUeKIG+tT0pjOgEMHWmc6QiKUi7DTUrdRgqwRED931KV8xVgBNpQ3fJl
sn773Ot+Xu7jRpnc5QRV4aUcYH4aM91bZrS2UZ2gQUvwdU2W7lV5KxxrE0t6Aix3oA+dKTZyabAJ
nb1niKgKeBYq0Gwhgo3GeLtz2tBmgLe+DNroT7Og6IBd4JPxRZwHmXvtJ79iituqVlp0RPW9AiPD
eEr9Qj0WDJCqAUgdvkqqQwXXYvAvwSEQdKjaB+2j0uDU5xpJmoIyEB2lUHVKbWTfPiF/cgshXQzV
CadLxOUlEDONxAqXyAXoAuGSQjt8QH0Nfyz8RL3iThBGF3GAE8BSY13BNiR45y+dkIHa8CowD6Xl
Xh6SBwHi6/2TxTWZzfnWO1NNxz03VBYkvz4kAtOKLZNcD3VSdjUrUY6BeRw4SR6+92TQMtPoNFOp
yttOg4+uB40W+68QJyvXBgwyvL9v982k328i99SnTRvyLvM6FbqeggQL2wrbCqas3Iy87nhcJswB
CCDnzUdpZOEExa4bpGj4auNZSPM/ueiQI2DMdMPQdYojGHRzHyhwHtBV614qsp59xOSJzW+VMrpD
Avpbc2Xzv5+Vms/euN84TvVZmkrx/x27jRD1fiaVUIxlM/iICR3hRxRrZ2fljxXc7JxbwMrvBqxj
Bfx06qgIzS8Izu/RMceINRQk9rMoAhOcNd5r70XBcV2fwyx5gyZrcayVuqDIoQaNI5Sk8b6MRrqD
EbyeETY+6usZc44bmjMYd3oxOTPZEamElbisEViu2oUcbmTn4tqlf0ZimqdzCAgyOXw89STp8zZr
nVj0UQSq2AEBzwQ6XE5lntkdApURvflk8xMRiaDcHE5fPyrIp4ow9KXadvMYHJmsv4H+h2CeNfDm
CtanZUhDuWcwpaPl/Wp1lIdq3Oq9HjIVHU7QEWcYIc0qu+J4u192tWWvA+UtUmoDu1l9S/QDz1Re
ezWYzl9Peff9DxuNBzRJnKZ/VZYjMbrz4iZbty3frSX80l8jNGko1xibMCdRpepxZVBb0OT4t3+X
2cx2k147/jN7ca4GIQmClx5uqsOicwXiV9J918vY+qRw4EiiVg72IslNB+9umKYJYwyyEZDaZLgy
j5IKQjKO9gyVBOaVhlEqxbYWwFHpJOYz9x/VjaZzqZkTheXWALmxkOjrCGNH6Xvezw217lQL/azZ
RAQCgRkCzwiiwoS4iTotrk8XvkH5nDjScG4hoHg9QzMtFQARwvlWIVv5AEtC5TnaoortLbLsCPs0
nE/OZWPmxVgxJMSXfUiYfSmsM06IJxLC6NgI13bqHTBPqG9vOlPJqvI2qm7lo9YSrICOgjZu6d3N
02d3DW4SM+Fq0w3S8pSEahfIm2kEZFOj5Xz7ytm59VrH3mAZBQGlT2kw7ZeYCcTEiVBIbnra6Qxp
gwhm8qbn2yC9sRCwowSZfPVN/bM0Q8+s+7oQ0nWqIkpTPssDosGGJkrXaOEA7WvXNqruDSvwa9OP
73oNrAoFqc519LBoLunz2q49azgIiiCL7kP91UD/3h4Ai6cqbT7ohG6IXbM5FbSOwmnsnwSsUfN+
ZGa9HdgICFl+/1Sbu/s8OCMAzfzxWMGd8hsCsVh20uhJF0Ldn9lHlLt6YG4EsyTrFXJqtAfV1aVb
PZ/J8E/gj1cC1NKWnXzB8ul7xd3u+fuenrMUCRvUhQk+x5s/zfszkZ0ExSv/Go8HhKi+bWgWPwpf
r6gAxk4OGBUolhzt89Y1URpGzomWGBWFh4Jdnp3PdIc/8KTbDfEaYNRfISlJxWWzIKd4lSnEu5o7
sPJkfmp/Oi288tZbi6kU8fyM2rjtJ+6BZWBw8eW/RsS161ykPNkEmrlNNTnx4bGEM832AXqiFV8/
1kzLcfbZiMP8Hz1YgIT7AaXX+Yc98xBV1kyRj6CiYdSWGkr9UKK8GUYJuJMmWAKNY19LCw/FRolh
byEvMuS8Y2Ez9j0mmRMw/j69/H3lhj9Td/Zku1oX3b3MIiFaDmLB3gf24uBEkeMhi1RNtdsKVXF1
B4uwhPgz6799ZgLQofFcRqUWbnuK5OWSKvT/RbjU/tGVsW5jEKgHC0AoOKXOW+AYjmVQAfn/DR7I
cePGWX0RPsE1adHG7vmeNNLTLB2959K4ZE3fidtN6rT7RtxOBgJwIgkIoQiBfGQF6OU0BNyinJ+3
KdDxxDGppTLbIhjoD1wp0lybaiHT8S+BrsQJQhbNOOYKVVdoN3AxnXOZ0nrV6r3YewEv5O9CHW5q
C7aAR4m6gNM+iIe6MPGp4D5L2jUY6WR9uTwTLJPY9mn1VOid6CC9HW4OwAROEYTn+5LHQnI6s8Ma
QMwYC5ZVF4LdrlmEhkDp1qu/S4YvFiSYX/caL4FZos9WFs95f6/N8laOcg+ojJZYDFq4aKoKjaPg
KwVclJNnRsoVtI9OAsnrXLLbtVmGuSbXe4vZWzx1M/aikiABg0BsVJwFxSRy3qldQkVRV1R9vN2+
W4MjgsqRjepA38ozpJI+GzBqcbES4Y5MkjkjQkVT1Nrb/GiDSXWYAwM+ln/kJWKHQLAvphzX3yWh
p9cwTQdBUYrfANCtKiq/BTE6E6HhQBhvK0I0OAMTRSoCSsTHu3fl+vsJhp4Ius1wsfpWdJw/Z7/I
l1ZVHT6fDezEAmHgrLoXUqfmhY1/VBYiaVvp4sbnniHizfb5l6Nw5RLaprmoHhlMTka9giVrA+dX
ufyrp4D4vZdJ+umge3L6CLX7aaGGN//OwVr4wyB0Ug2gDf5Imk0TVJJHnKpGurYF1ZMv0Q9Hrpcd
X020cOhWvum8uLsRcU0HeHBHwoOYqm0glya0qKXfzBKH7YNe4fRojMLhu6rT8F4tDcxnpXbOeQyj
m6aBBAwGOL5ttXzccQZTnSLilnf8vMJK+V8Uyfv45PKmiSx8AFTPzsdo0LF6e0GkbqAsenTfunMd
E2c6kQoQZbCvQWg45hdJEwbpFztJJ3vCdBk7f4uAC+/o24YCtO3wYwXhhZi9tGh5aESNAwvMumFg
DlvZ4ZjKtlxALNwCs8J4JPn/1d0QM8o/1tS2QAxJ/bg2p6xIkEPEwpnSyvGini4WFi/UxsTw7IVv
0dcLv5KXPsGZOHm+6T70w5qXhjxA8qqCIPjfZUumRBONPlfDnIRS1Fg58Q//snO0C77/myQcs488
f530UOjmKRGZ2ZbYt50X7s305YRkyz1vYb85+XNlw24uimap7e+gdnWK/o56NIf7u9HMgJwh2kAg
i3vbADsP4XAqOhgi5iuTX8FyrXergqpFMzZPvZHpRCAI6LPz2Zuw/8MeKVpgnK27hGL+uKSHrq85
rJg3FukdyT+b4nIlv3+p80taesbmNSCZz+q1fXrHPIs0auAFfxZbMxFaJcweBFLMXvnHHni6aHx4
aYed3n3lAuFEnfmviELLYvBxwJYhDnAfGCmmqIoL6zC4kV3ZnaE7EvDjp2DtUMyOD9iv8FBQ4V1d
MxREqX7qUaDRzGIbcnIJC113Z9YLIFUa3iSaQqUun+4iTtV12u23aYZ5CaLB/rGz8fYmFAzNiVIp
dmMV0XtTyVuXUSGchcwSxMjuhHfGTpyb6mBPIjcbcSvAyOHjMORBnE8XdE2fp7HP37GZ+t77/fZq
1CInrwXJNCwcipCFmw6dQhhSEuWw1cRxP9oampPNYcWhpiijUhRsz9gWW/MDIdMEsFfMPiIqB1ps
5V9rKOIxvGAvtVtTa6pXh9k2Q3geHZ23xaNfVmpA/bfM+8Yn9T/DxcqAgBtFP97fS5tdTPry0fuv
flSrnL7DRq0Xz6Lq911zzHO3CtreIWK7cx3bmhcIc2DRsV1i3P6wUPsrl+3xZds46/kYA6yFYWEE
RPuZpMmuOTXsyU5kUXsbdaPOWyc2+91dbkeOM3POsD7UMnyHr1Y1LLi8PRrMmIkHgwyJkPiMgScG
ldNeRVa1pV+H72AQKhWeM6mkMapsggal1MCqWINZYs7kGzpWCTdc6S+tVTwrv3PpvwUBEDNtM9+I
cyn00MSL9HLXC+bOie7+Arri1afCRQ5gnfS3AMAy2G/9/spFKz+we3Uf9VkN7I8Z+bdFDXwNfqpp
0xCg6AhV7p7fVo2QMJZ0ErEkS6RzIYnZHwFOfpATppV3y4aJP8xNAI0lE+KWZSI7cfQg04jPhqM2
JBF2i4PS9O4nZ8NZLZ5KR94cC8YLxt8MVLO08fwSSodxSxzvMt0b1gWlrMHw8hALxpYY+cCOXbSD
4GpQFC+wN/5zs4r0urP41Mj05wPy+9M4rqsWqN9mnGvUnzbIZCPitFDzpVEouMDHhfS2D5Z+HDhC
xrFHBAxg/ByuLlEA8W3wJjZfAYj83Ew3IvOsKFpx+CZo1Pt/vGbdNIsF+KgQiVWZ+vZ3p9BSD/ne
rgSAWawSQfVPrIPHZvBD9NHGYfxBw3hAORNTKxRKg9N3kBSfNjqQtGbulUATpj0wjo6fQeRzqLdQ
3d9//DOmdg32qcAlEOpfKXsLof0ICNHZzeXggZw+uizCAvk+jgeF4PRz7VRYIGf/LiVJhQZ/PriG
d/7rjnBMFskmWukQhV7RDVjNHU6BrErLhkLaO20Jw25LGXVyrp7p4WtiQlEPXCpTW/lB9KNOCUxb
5Hlt4BbFA6f4Ow4c0ltu7B9RBgksa/BHUJ+rlOqfWr+bU2o6nyelR25wNvK5hte+/1D2NHkHtPcB
5mTw4oerDHnJONah6APHqChZs7gPoWDDeIoP5ZZufml50oHTMLFNUKJ/xHGUTorwfUh/Mj4gdKo2
n2kPm4sjHEotMRXaepHaThfIF00EJR7tPPdF0sBuRrVgCDDt9eQN/JX0STHZfnmpwKg5RYbdhFWo
9xfBaNdVJqMW5DNXQgCG1aXnQoaNvKz2AcQpteSTOGYBp2O9GrBv6bJIsQthBdsOZH+9fnvPVdrS
w6muon4boJfJ7E0vO/IC75SLHLO8v9ke3fwECI/EMeBoCSTZHmZHUQRxmUC6/d/x0rvY9tDjmFtW
VfP04BJDdlemwqJLA7lIqzndK/PbZnNThb3LHjoKNmM/z5Ph/YgoNjcpfFHy/rHSC3lA49PLsLxd
ttH0hhcbdJRjG/sUgFBUiJbwHoGA6b3uznalaUZju73bhM+OfCai08d8YGa9FTbr0DlPIcDPnvZb
EkRvnMnRJ2+mnJcNYg/nJEGCj88awEySTwzkZrw3HAvPKbb19Y5A0wCd18rVjZqBKqA0r/e1jGoh
cYMJ+fP1vIYXDsUlQwX+DJFUYMESMEga5UEO0Sz6fT3svkqu1gf0bi5BqUWY5g0KMxKEhcqlSFYL
WekwuBvbtkOhu4/tJ5snfFEdPzCAuJ/TiLD4hRiX4jirDrAAZm8zy2kHp3eHtbfoBUylrFm1JXL+
zwYzkLDNvfdEqcZR6pDrlqWXCO76R0XwqfuClNKTQ3uAgcd8RAWtwvFUIuOORFMj1Dzm51voa6IF
yuxkEyWyX/R0vJGZgDHcbG+flvDBIbwU4a1eIrgxFkvjvf5pHqdu7q4WlpurSxDqySxDtYi7PuyQ
amZcnPYtS/sjxRJ1FbTYpdBOEA0RcW0GnoPEmrru4R5vpdgNUC3l377NHgfv7uT4+2MRGbfXfK58
FqRSDarA3rCNLESX6jXCz+OAqUhLUxtXOYMZZajhfAbUXL2wI4X0dECCmiY2pRBHQKg+Gs76G5Su
QfQ8dk+dCMbLl6MXBbSTixp0dPAoeyHbbYjOXISKGx6YkNwE9Ni/6QOyvixXDLa3srVbsbzPqGHR
jic/gINshEo4Ea0PlZGOua9xbfafSLI+Rjh0NaiTW7RY2fBVnpW23jySFozZ91gDp4yjrbOg4Qcc
EWYP4pTXUV5zXRviY2hIC8ysGNmLfBDtBoAGoazYZZPjYdI57HkLOA5MscrwfmmqiEhj5R4t91xM
udm47gdfsSIlMeikicwGn40ohJfwr5hD0MhjrUXA+TRqJkJu4K/9ImbNSodHAbyIHWa+kjIQLs3q
llnGYB1eV65YqegCm7eMJpJ2NqFosFFuzebUur2dKM0WA/Rp1bwl/UxbZhdNvWjAxrk/VBkuTfxF
tcfWoi6uRPFS0Wb78Uu/I9FXgxH96IcVmBfDvkXNrjE3UOOTampluguZ80nDUDdEmlmRQTnXVRIl
kvhZYLSbDmklYs4BX4os89t0hLP99E1PSU5QlTVK5OQ3jydSfT5VwyoIQt+gO2f+82X4himHsXB/
0AcOYXVqNXbhutRx8dgrS6uc6qr4u6hRnNgbU6xzR6JwnppucDtKXYfRc/obcq2gEaw+CwcnoHpA
SFQZH6hVCI/AMt1xDk0vykYlKpwWDtB/NvLfzNtQh5gMcpgW/ARe395GuMp65OSvNn8ip3CkjtnG
dOXWr/PcjQmDS/IgQcMjkPEsZSbFqscY+5q15+y1i0Y45cjwN6I1Ji3hS6pgIOF9iYpzVoRqK3r8
lFY/2uYM/KhIlYN1Br6xr2f+Jk/3XIdzVnODOfQM/pY6XQ2I1Zk7SRposUFOtH0ethR/3lUQVN8R
2IS7ip++ZznB9LtbrGFc0YX7ZI/oGCEnz3izr2qHnmCxU6V6PPY+acAyWa1Ppo1mIR4zj3Ifo1OL
NHzELeXlLY6okP627p+x3WSYa8krnrSY18yjDlf3KGlg3qzXrymeRs3rdoU13FXgV3uGnpwgbpJT
oJphu8kOoex4UFWAbagKXxRJOKPa21mW0KUQ1QhYMCKQVFhvoPtOzX7utmMkBgyzTuh7QU0HEnLQ
hW8xyO7mG+6nnmcpZFIb8YbnK2ii0qCktjKugaf995QklBa5zh5Oqwf8IJDMkQzkMh79ZRKf/lID
NKrzqZhekn9dPtFux+1gMEvWIjMX3pEx/1PcwhGbvq9pMCq+p/IgtYhqBPkurO0+5uBi+zN8Peik
AgprYSftXzbo1u3lR25j/5t59COKzchpixCPPVk7HRhVS1IzC2Kpfn2kRu50WpXwPUxRxs+/FpdZ
Qbxl0qvhpEmLAcSCSNNQAQEk8Xw4A/Snuy6jZbL6kL7AhFW9w9LWiphhzerBDO2kuTz+WjZE3ui9
bi1jfNYL8NnTiTgoxO4Fmn5k10cTvJ4KjofHb7Ho9iPN7IlWv2qc2XawdquJ7vjYt5LuZnx68XqF
yQ0RRdBqXi4zUwUrePFXYP0nQ/2/i1Xu+5pO6PE7yr+sj/tiYAmYONYD/UxyDzmtPbTnVAJtjaSn
eXaybHqlWhg8+axm/+/HyKdZMXxRn9i24/tw0eS1hFqqaW5GBjzdFWC62Lk4Axy0PjVHdouvyWEH
aIEqvqQvDThAql6mfOxB0jcsm8dDo4hmzqLcx1S91jNLjmWqDQeJp+9fgVDqtlQ73RvhECXZ7ews
xniozeUvWkJacdDDhRB93PAXAq46LvHZUcDxVy40i+TzDP193RjvzNosmV3uPbq3XBcf59iSKpcX
5ho4Kx8aq1F/npieq49ky22jhzcQ8mWt266CCf7Ai5QJkPmcwmA69SOunvwAUf46gvfQeGyOTk3x
FHYwuudDyosbhnCMpukPpd/xw9wydc4VErY+1EEVf1mFYSgvIdCE2VjXqiI+mxy3YJSweQ2re1LG
70aQjQCcvzE305NWxq/0IdUH86LdMrTCckqfDlOJ445y+Y2/HWEzl2CQ/y6nvN8Ae1p7fhXZth9a
5LxhI9zE3JN5yQbLA+sudOdzlnKUNDJufh4mWtgNJve1hrPTnsDwUUNagrRmV1QebVl4/KcPgxKK
BAB0jnz8zg1HO2eDkXDsSLUlh9kuKdvCJn2B1J8sb4m4D+3o+AZ42ECceFSUz6Mb/X+LDCknW1Re
XlQaYvEJxVsZeCju3kXZGPEDXHOvBMqbxVu36DyTNvXsoUxUYgdEesuK/rstS7eIeUpZ1JBiZWFj
Ch/O0kVtiEwv+Ifeylaqv0vSc9dHksvD16l8JbZkIirjrzFXehHrDzH7ApMfI3wU7vyctz/iZpdU
xqrWBdMPtO9x6pJqxal6DtkNMFfantRWQmPqmg1firw7OUe5w2n2hP4TD0NK2vC0B3rWCEuKJDRL
bCQ2cFgLx2FilbVMwbzmXlhsfRRKu7aDxrWFqveKGjwCdUlJB3VETa1lP63LG5R9lOh3KzH7aoSF
6fI+O/FPBMzgYE4YyXjopqyvUcgCy8pTxiDP7ncbp3Ujhx4o+jLfA9OVdTyh8OqP3gdkSy1X/9m0
DFlV/mJYZ4EcGWr9E056GY7ws4eBKD0/OsFTpjSLzHSiDJA1ZDFgSJ1yXfFi+XKUNQFLaFBAiA3i
TrU+uDfzsW/LO96YdAUF0QjsEQIP/cfH9NB4Kc8N/UvAgvnjeS5BUUU3gvEW7xVD6H+BqlywH99x
O7uMR5a18XH1yI4DE3paMuW6EErYJ81e1e1wiNg/lq2TwNr+wCPJ0Spx4FwP41zj2M3pr6Q8rY6T
wKIKRazsg46aE+1xoavatqUlPDA7pD3LIs8A+4kwvkOy00dBW56UENnb5hNnaSHAZFBM4vDKZdtj
9HrUjzIefUv0mcLfTOYnFxtBIKY1TAgP9AU/LTvzpbofqdDL3DXGwdEmn9W7UWL1LHKq3+RjsPW4
lfFJ9bSSlrp53rnWOPI5/cX5/rC58/fd86LhXFmUkYKJCwZV8+VhPlYYwGtJeDUH43Q6lGir611E
dWBVxPTX4EQfTkWOY6Jqd6ynLZGsc6wpPqE/fuC8u/a5fKBlF14hdkXN757Y66j8gTmXDOwx8mXq
UVYV34F6I9amvLzGhbCBOv7NdFi54njMDS8ZXHIGC1rZ2/tFjtjbetgyMEMz/rjE/b6lKiyjmqBI
vSecwn/P3N8xMRgc2NVR6lU7KZtj+eZdrjwKzD6B8kuKOzgiSh9RLL253H5y7MjsNpkq2XPA34+v
Pq+L7RtxQos8GnMdHXFa1a3VGoKQ+yxkhEmpTj1L5aV94GwMTIYHB4nGKjEgFTIGoMFrJLU6MoPS
gCiR7l5rRdoAZJ2jzzqSA/XuVR7FwaENBc+B/ysvWUt3nszzb0kUwGmBWbtI3vHlJp+kPFnN/qw8
at/z7YTOzIPweuiaA/AZiPQfa2kx+eTcvjV19RrQ1ZuC6UM9WfuJyMuUz9zwr5MKggBljpEuXKrs
9Zg91VnD33ksK0Vn35fU99nGtU0LkUWve66Xg0yzJQd6LiW/2wYEQ7kAjY7M56Ot4Y/6ajrieSPy
TOpLoMxElOrfeErQ6OsCWE4wmSoY89aaRcJU5yDInJmK6q8Vdmt3yKeNLCfjJFb7Wdj7D6MzgY1C
7ZudmzE8bZEBq2bQ65G0WQMThmAM3PyS+B+k4Vr/T0mohrZSWzM04gkUMvx0HDyAvHZuWK9pPkRw
BIxg00gjvJlVaEQtveBclYZTQgNVZXmmakQG4wRxcsk+AEVKryaIoS4f3qskv8ha6pOOdvf+CcZM
f3gpgX0hYBoPhCBLXimrvGP8VXPMgtXKMef+7juUyp2CP2+clbd5bPD7lodH6LztKCJxt1OYpma5
Wj56kshWrKI/Uq+Hgd5EaMttjjkL1PFcObOG1THAqZgERQnK7FsbHiPa1AA6Mpw2RJj/iQyQHwY0
0GHF7nkdud+2CR3RBoU5hbfeYEmbajtcJ8Y3mfpW1wGwj4klolnkPQaYVxznpDG5jZ0SsdPxDm2G
pWXVckZC4c2HSQ3A+y5XVtyRLcvGLC2iuDZQ7z0GjM6QIxAL+x0Iy3/Pb/Q9ETuHV8uOWqC925t3
0pjQ5ffgNRA4ZuxhLy5tLYvl5856zwSrQo7NdHNgEq9+T/E5rzzkZrYKR7izqop9riSpFSQbMdsj
9qQZVTbJljM7xYrux4qF7WtRNb9ITAKeBB3WVzpbzN+a52GdhdFJ/QE57iWH8ic4vutTgT6S7hqe
m/IQtjxxaaj9WehWgl1vFskGdkOflGW/O8+ggEfE99jjBK6Ka4KXOm0fi07rPLpKlAX28PocyUaD
sK24iGPs9K8FwCP4IRCsqJ98HxQ/hVRIsSUuGKsz7iyZ4IDOqfpyUDukK6bt9sdmoQKP7T1DtozW
C3jfnq+ii0OXVTkvhLa8HgOEz68GUR8FPqrJM9MZenCVgsqXu1nm3S0d1TxLk10qVYIoMuf8WaQF
ScsLlL5PdWPYbyx8Vp7ZoLSxvz2uSkeTs59ppLb9y3Vu8NEQAUVwo35K7ryj/zal0BUwhA30OsMP
75Yw7dnf8iO9PVTZuMd6oA5KazKmWHHyRGUzkxQ4Tv9WGxTJckJjdtUGf6ShcBOLFWuh+eB/f6Rp
VBGcLYCKu+6HVBiQTfE4+ADmvZKgL51LLfiZAkmZyc9J0aRWuAlC5zUB1FuOQmEOLKwZT3l3QCjh
rIFS60LlLd2rYV2epSij9PiI3hfAHnO1q9nNcXjN5B/gNvvpIJvFdDCUyVxDtjJtzW5jZqbsHGZO
DnaT3RZpN9SzsVmalFlDKipn6LsRQahsasJE2bZIhsn1GuaCy8WtuoCKZhGnylbQIY7KXxb1XqCs
xYwitlpxZJab/EB8wt8GpeD58TN+NV645kh9Q9v119gJ4TSoYjeYS2+D4wL14EEmp+xXWMuIX8Pb
BeY3kPFddPFEG72O4TpZjc7AWFBx36MhVzVevQBpzUm2fbfMHZH7iwq58/YLUappf2VGoCQijQLY
elJQMdr8UPMdFpQ5bbmjV1CZYZf1wfXPYKJ2Xvf4ZGruCo5PL4qrQz0EoY1Djo6KjQCYkjJL8l3b
xOSZnKVnZufUV6Vtk3XLdURmcFdHD48E8A2bN94Qk0NXprw5raPDSNz0N28QTvb+mXVmkAqprjWi
cxXu2iL4NAbV80xEmBZ053kdXC2ZYFKzi/7yO+ZDstcHshW9uI0c3yrA2DhhjCYIF2GbKSwq8jrf
whMwxEFH/QWWLUYH++eTUlRyp+gKyIn4+pI5uZaP5v+Rs7TSQvoDiEksd1j2kzz/JI+qn60o557C
xp78I2krYXy+JiDmdxhwfva1R0dNqEa7dNv1AvRvick1ab5yUyxQMCAKOzUQfH2yu75CREujmBs6
Z8kG6lOT0b6NLX7ERjPGlfb/J/dziijy2V59B31i1E1viz1VMi3Ux/brecfNKVNzARHtb4mbvh4h
GTRz6UNKyC/1J8BDPdEBOUgBedEpVrb9U/IJlx8w30VqYY5P1PZ5Al3ixNukf/YnAh5oLVdI8sWZ
5xzUDpFt8FPOGf+9COKz0Z0dIAUOM9HzGeTYuYvhyzoHqU0Yb16JbBbsukLxE3httDgTI0r/DxJ1
5UvBnac/UlaEGkUzwfElQFvel2kjrfu2r1lnyFJCMNLxjt2D6k3qnW7caIJw0WeRKgQLhk4LcmCV
bfw7t8gD4EQl+YtolK6DI1lx4UhqGCWEUXFpjVNmjtfoxWsIo1cw02yhKrk+bD8R0S6KD/IJW7jB
FpL4Pjol2PMc+/wfqoAFIn6LAbsU8xBG3ghx8DOWP1BDy+nd0H5/k2t3k6rOcEWtBpJDzwmZweLZ
o8DNTEMK7ncG3fTEMm/CmE7Vd2sxTX3Rou00Dv6cyli1St5CVKZSxJXyHM/ACMjx5P0TINOqswfB
7Vr0OWy1ny67nZpcF11aTbpT98gLIUKysyVWqQe+JlhC5jeqAMHb/lcLw8e+vA4ZZ6sZTW06ii1f
JsvVwAgtNr3T6VFHhuYDhtj/rw/heeq1kEFcet8x04a785JVl+W1c56M5d50zs5It7+gizfazrwT
4y/wFF7NRZwfvCBsbZ2aXFkTAaGyrRSYJBzPrO2ALW679Ymu/2063dQTxp6aQ2qGOSsB9kVooRWb
OfLaWmS5mEJFIS5HYhBcvEw8TBDQIjZEUft52emZN699MyqXFywrMXgZ/9Yp2YaOfILjcL9Df6bN
HkrMuactV3CxSlg/7o9+haLo9nanMOsa4yIYG9+EkTkhLcL3w75O3gWeEwCCUGU552rix3e3M0X9
IkZZy/guz0xO1fwAnE+/QHMfDqdlWatn8TQfMEZ4DPDas6+epJmt0uy+HSNSRDx7Vnl0iluNjOhE
s/NMHItw+hqnGCqOFZ5qUVlDWlmCdeyZWpEmXE+Xf8F3j63RODsl/7teCDmftxexHLwv8e/1EcW8
byTTv3nCPByUWOSJBNFPU2rbH/1EEDJyv/ly9kdvE7E/zVVpErF4+qvLEM7ZLgqn0J3pjIaLNDbQ
hByQcFWX2eiMELqzunJXyG+qqCpTqEaMaNKNslwdQ0blIBFSeM0/Gmm76fvnRwoQyFFV+lXsqTMC
LEOeN4QRXUoU36by1+Ek3bpYtOvvo6lzgdloex45Bl/bB+EUqqIsMmSDFKKTXjqJHiYVzef0iTpa
mnpMym0ajyG4B0J4WtkO8X9f+8DVLNk3PfJHQfI4DfUb0jikIhxvLeN3hUAaOlwrw73bvMFK08fm
JfQBYdccxnU3TufP/gEG8XQ2gnXOfyQpufmW75S7txkEeG+P8PxJYgbkFIQdieHOhQyYM5K6nCQe
ecEedpuR5G0E6rvavMEoOM7T3+p2ZLF4LknK1brwzdXa/pnN4vIOCpZEgco7X49Xvo47E/c9Sm3B
j5AsGl8owYlpZaNJDi4fqhsJKgSWFVRw4EGIg+dkpsVNd7s9kK121axTLnxktwSqiwVjhtf9u49r
dKJwAFMLKjxAEUmGFTcje+TgYyxnJEY9js3qMD1ACTNnYJHxPfH5ymAjVwRRQhqSO1jmXB+9Ldlw
RVQa9rKiu9h3qtELRkgXTXfca/rmyvccG6hO6mRpvQxUB9GUfc/2X8PE864AJ9dJhAEwgQAG3/U4
RvS35CdMoBlgLLQZGJpe2KSzlHyJPBp1axkI6Z1bg6THphlphMlaBaEzYZUbdS0jzyytvnBlbPtE
OGGyKQ0XT+mtdUSCX5vOqLdVPJplhd5oQxhBU0/cCp3BekE9H+84QA1GsdhL50ufCuJMTUq2ZfVc
3zJk5JFTVHDRzx+kPg1W8lpoBfxMRlKxKJ14S+Ajz2kdFtCheDwvmSUkMFQpcOiLmxTRuj1GHSBE
0loj4j2SfTZGcGN9IXcXx4eSIq5gBvNOwOTWtzIqdkyrEDoIAdB4XDOotmCd1Z76MwWrRbEj3g/D
YFe/7rSjgxIl7Pfz39EuAS0v98SPrQfPmH/J0T6VUFRuh03kgQlNfAfjcJFmypylJAk0RiGJ9hh7
ed4UK8w5HW8UmT54N/E6xL8BxD48S3LW993J3KqNaSbxqZ4oZPpdunQiAgCSMHg3kApcQAACcn/G
SIS1UH6oFU2IvWiYDuGQ3zqd5yJ/T6CETQb9N2TZnV2dc6xmF4Y7l6+I5nZGtEEXKp5IU4YyIWfz
++TglP7XIILq+aDmEaWHI8W5GgI6NxVg+iFqIaSOacp6/fzhXlFQkMh/L/acd3IHrAE0zG/rt/bf
82gGRk/Y1afNcw/sjQm9MVv//6KSR2ngfvfofD8h12AwxCjrdO+4PdQ1+jGZWkskXJid+vE8yL+O
EveZZ/9KRJGaNrwDjG4ts1scPz+RJ1n5m3ISqoWnnmt6ui3TYwAy6bBG3MwH+iE/jrJ0Hugp/ryH
kd7cTCmu72x7WazZyWbZJ3BBrMqx5hiJ+HDZHTfafY+DkilPEqBR9m+vXMCqd0DWioLNQ1GBF/+c
SHfpVQ1BYndfFa1+xBDhNtCIjZ2RA9ryz1Tx14m07fzgM/N2wJVXhP1HAeGBbbdZo12yItI0ruCH
zzAuaUOnmRQio3Rd3M9dIuIRseeVUfnEJvGDrYXWn5PM/aGP5PXZPi+uYZ+dwT8BgLiMipogd+VA
W993HVnQPVIAhc9iRb5Rgt88d4L1jRT+Q7F3zgLpzu7a5XeHL/7CpBIt36HDHWPCEdbL+DR3oOcI
nnwE8Cw0V1TbehbwtahK/znM9SaZ8iM60cJnW5AOhQ0Ily3k+QxRpxhJZ53qfeLTQLBdLSmfrCXd
5b3HSiLMO7R+RsPgHXB4XRJwy3M+IK+8JQLH0zFJx1U4mal5le4gi7X3Z70F7gk2r2pP/bT0Bwte
de5X57dPJ+5qIyiGVOQrM5D7xslvCVxKtL7Om1YJtSGRGoum5BC3xZvkqkWYPkJjr+kWgXQJTEVI
aIrbw+S4BQodfdGtrgNLl7/yvWQlHtaZPdjsS8TlfJAk++/6PBYzl/sC5iEaHrPGAPaKuc5jcYjB
IhuEoj/Ve0J3qji0SLXZnIlyeEQcNDJDzXJOBitiLa9ix5Of7v1d3qZESSznFIBf3ItnjG5a24pY
uAG0ZeF7dOMenb/TSEdRiI81ynBaYeQfIFD9iyskJVR9YLB7Y3XoE4zi3AXQ+WfB2mRfNBgvMI1o
KZr/KzuPl2Msi3O1VlNvMOxYkpZgVJ01ero0EJE0xnsxcW4IM/lYQH1F79clGeoGXlMBVcPZ1mxr
cuydsrO3wi8OtlhirocQxzxv5XO4RTelWvVoXW9jEtzN9krrOvQqJoDgTnGqomJx+BO9Qiu6vb4z
cyAuEnxRwubPMdWgH7a31ubVYFS3qm+K08uxHmghImDIzyooJ9xauaS4MAeU7MvkmfTFrml+w9mO
PsnJd3kqHTXeq7dH8WsGKmnm+bIwzb9mtIsIpa/ODHS1G6QCVhKOe5Th9aWkk2we7R6zP2dKiBjw
yREfXXRLqd3bljACkm5drKO+CRVYt7zMKLR2ttxpdpZ3tsKTRH48HG5IkxAIIuy5Otza4opPURtN
qJwZ+Bg6kkinOz/T8AKF5RnE706MVJ5mZ8Qv0wzbWunCrGQW9yueLMB3VAbitszWTBwPNsTur39T
nMfYRDwBt8o4HtVen/Y+8IgjZg5ztiYyeowe2M5JHPBXIH2OJ+fsvAnaCfSk9fia3QOgKSdEq1+G
Bek8/yxrqofsXOFT+YBdaxbmXks5DKVFsOLiaVNMGoCb/ivJC+wK6+ebs3BnN0ICYdsgMUengpoc
Okwb6bhflQivrvddm/EFXnjQCGC58dDKfTMAnO0dXtgPi6sg5z0Aa37EesieXDV0VZ0URQci+iAC
7Ah9fUezrSAncTXGtw03hF9/IKCHUA987vRyHelcFTuuzPBRKTaqzgLKaSjnBazlDn54ykHiEfTF
WIJAWjsgjJl+InNiYvo27hqCmEAAkyg0XUi+8zGDqhx4RTR6V/OwhWtPMpQH7zLO1duDbaDaIjKU
amc0HDifxSdfIJUoLY4wwxa20dJEO+OMUZAbccPW4ThU3XK5LjcQC0RVPUM9i70yoehmyZqqbGMK
N/F7ndGT/elwmlEATtmm2cXCZOnH1r+ww37wjaiOP+kRMnh+YxN2W8q1Y6G02c+YGwiZj91QbCdc
/urBMccdP03v+bksRiDQo1FGt047cOXM6cWYs+2f29JQKGOCmU1QiiNjxTqSllgXhwrc0G04DbJ7
69BTeRkiNt453znP+cLO4djhaZvN8uGmiSpnP+OnQheh1X898I9gpU3OPoTVzhiu/YpGBENuisQ7
S/jbJEqkic/AQ5/UsfLebb+DGM5wEQVDn3vZc2oByDBmawk4ntMJPWN9jD0NLFl35CpZa6kO/Z3I
3TQ7ZGRCm3t9G9iAxCFDjVjSNPprWX6aSzfeJTnH+X7fb8/1HLjdIHIOyeIGrl1QYtdeTQtT/WAo
XlNnwYMg0Xox8gpPESCjFg/mPDR4fCPaqt5G6J4TCV9plEk7S1ERJU2V29yQDj+lzD+569AewRsA
y856LsE9jnfZPIwW5inhhmgcUXeTg0UQ5JOw1H5TgLKrTAKwgSH730MArXS9yw/H6liDz5g5IGS1
9fo6qaZZfEYWKy5IKctvQtrX1VY/UfcozmeMmQpX/E8/SGp7zgqypxcg0oJyQwGCj737IrKyCW0k
jWpdO6sQJ96ySdCaaEZWH0s52zGcBc+8J18jKdyZsiphwHap6aqCbHp6BNhmDU+dZ2FFXoP9NaJR
KaUbHuS/+U1dDOeW2Ob9FF+rW7/ZS1N1gN8UTvsZ4JrAQJZ9vpO79YXani6RohykHXbAM0TnOA9d
SZ8JD7t/20o5B3UYx0Jr62YvU0WUSWjmzLjtNfXLQJIxHhPopuv7gsR+yTgYBiAC5d7jLi//1mqt
uMfr35prEIc8XE5XMvqBSBujBTZ0f7NszKkBq8VoR/IWaQNRZjBop7pDRaas6R6iHGvuJJN0MV3f
h3bK+FTzt13v7uMguIaDPlEadMRr5Ywev4zFTSocENgl99cruc61IccHT7bM/b48gIyFi5izVkuN
3M0qflZ77i5jM//GRfzzo+9tnEzztOQfaoivbcdim7Zr8O7foEPGDMByvmQNku7L5xFty6QfjM1N
0y/oifAVOJl43uYz1fzdesrFb0vBsqXy2ewsvuOMRpZ9yfjipI036tF+m+10Az3puu1vYCEKcHgf
lCwW/zAb72M46jhMb2/5e0S9IhQqz/7FrA0qojv8cLVlExhx5sYrF4N4WcEq+FQUQg0hBVdpybJQ
fVGxLN2jEqDIqCxLms0L9xWK4Z4QqqmGOwr4UfUiSXT6B1cvXUSXgOpy53mje+WfavsW0oTB1NA5
7DSfPahcMwUTtYigj2M1fYjYI99/4xVa3vb+9XzZtlhYkZtymvUI6CiOI6FbRow/sfm6bLJRiC8A
uWnPmhTS9583Ii0e1LNRsM4dnf0x6jwId6FOrL1v+A+mllPDGU3wCDcGlY2aY49v0r/t9/RMIbQM
6XZtCYkenXCZfLDdfm0nnNYu8hOuZCVMNJhbH2BhiYw1vBTVMDxZD8MpRWxoPQmI5cVWNYVDGiNF
q6b1BYd9452txL+HOxzOH+l/vj7E/pIzyOu4/R5c8Ry8mFMjYUUZmgvw5pfkT89DLupIHuLFSrjE
lAXLEanvYtMxgzctuzJTqG2rng75ESqAwj7R/v7EpgqIypp+DiMRVAoqvRCTDD3b7k6oj6atl612
Vfix2KmOWBjQQBFhXVV0JyEjJiATSMhhiXNSCmGwdaaXKNpOwfMMKL96/rGHNoWkK7wxsGLh5xkb
QbAlFc2f/Fy4s7F0BH91KZPsxknAz9iIsPFYRtW+uPe7+ImzDnXnY4uchcZbXmnCKEgr77ZZwA1V
6HWPkXdbfgmELOeHb9VoIvSGbLGcBoBD43DCCcsWsD8rqJwuy4GN9vuf76V5ojAB4hAzy7ITTDdX
mXkQVu9llr0g/T/3vn40u0TWIdwUPY2B70aYA7nsdzt0+kllBnRVS+ijse7Z7TVtx9n/96OnXLoW
DFqRW2yl9rBD3a2/L3aW/J17NGEivgBw7EKnkqV6KRqOPWvzFRE5g45TGpUOvwN8h0MZS4dx+mjD
MXc8A7NGt5iKIKAF7iPKeEJCDrxa8XOOp3qxT27HktZt8SfvxZhNKc5Q0BT51co3lLpiYxQJdt7v
9pGtJBefi/sjzXYbIA/3pKqfpP6LHmOcQNaiCXFbR6m348UD2GHn0XbRgw/POfeUOIBCX+bUkIce
LWDyqW/HEqa+CV3lwffogWvhhsP151OB8EnFTQh9a7LU73gSeWNokpinBTeldrdJsljimH/VWHhX
4MyHSmZPuGz/87wT/s5YJDQ5F5IuzQwLwQ/1PwkShQeATG1aV+tdevhnYyy+MwaXCSRaUh83Fb04
cYLvjPGdS4Z7HPMt7pJ0WiP50yPgzRvzaaPPeP9NYvbldCON7J0S9fMtuQDoz0DPz+f2irBuXJRf
aooGmdYphUo1RqV3xUFFV5r46OnDg3dPQ1bAJsim7WW1B0P592sy5ffrmV9zQ4O8h++ELax8EbNT
K6TUzfP2I4fStrI3F2PphlpsNVSTMJZCFl9noMWhvKUTZ2nGinZYsrsCr8ngCESZYkT5D1SX6d1z
Ct4SYV2SQVnAzustwq/gxqcUTw7EpUPb1uBxHdITP3ud8tkRMDLtJUQMMoNAgZD2vPkwlCHzKko4
brJG5+q0mvt8+1NAOVMrGEuO7hGedv0FRv/6CWXsFNxxGisBXbOevyD/cM/Q3SsmRX4MP0FoqVUt
bfpJfRDO6W/UWKEokPZR1/6oNCl/13n21XHqw4+tyzpWHpq/t+c72NIGQdSB1SUZtc8MndhQ7uk6
f1NxGj8972YQI9wuxmt9fGRhappZkCPMXWmfur5lp8Uz+KBFfpwolGNr2r4CQzMiiGxNK7CZNIo2
jLBCb9oz6I7svvDpbLCvJJkCxctuYRO4guL8JSqWT1xiQqXJ2GiqXFtDudnldjb7zcZu7PCfDsPh
6oURBiyxfNMlyB1wxqJIn0vFaKQEpVbvjgprYKqtkNsGW/e6z5v1ic4fZJ1Qq5LIM9mY1CEUVxxV
04YoTc67SMLcfolWAd9ptua6JELYxGppm/KRE826b18vZW1Q3c5Jj5nqHNPo0d/h1dW2toopUI05
F0IYQDvt0Lbzl9wjYSpkZ00m4Nm/vgRjVEnfsebjlhgpzoNS/esG1e+6YII0BF1y3aLZLFIyjfLF
GXxGTlYDLD9Mjdtg205GMsdVt/Zb90sxmqGGBYGICxlqbcjP7j5hF/ogGl8eXIn0zwQp52tVeh4U
Vh64LgU0Ama/rujUtVRA1pnGkpyh0qQWfLCIqltlQkqmXFyJESynckRGOqxCRj8RV3nJ1CozOVOX
P+i+BneGsh+1spVaEzR5aXJ+ilD37tCwskAvBes0w/n5pEKD7FUmJ0Pg7dx4AMXB+3lDiSKaflKD
yUZTg4+AytTfxxPhhEtACS/rOqh8V1YSOD3YbnXLwEq55l/LOKanCJomNckqtBNGX8uJ5KWbYMzT
F66lTzn5AYThTtaIxejepFZMCIrMjdBcIx2FkXMQhEaaG2gGzV190tdq1Y99oLPL5UBmUebQozfY
9NyyPHDiROVVYyqUQZQc8tGy345feN/Vqo/ntsQwLyFRslCIVvcd0+Hto7cvZViG1A+labPdcCj2
GmHPHi6s31+k6pkg6olvpTwi5ouGJgrVN1NSlK0GhyUh8nRWxc1B0w5r58mz5m5SmVLKJUrIS8rl
Z9y8CrzXtPHaxrtFuAxO+uNgNZHQ/D0RNsmr3E0lnA7IeHpqmN0Nz+fgrUZ3FDBYKseESuVJX8pN
2lI9BTi7v/wBX8upTQAjgQttgId7em6/r/0jQFj4VFD8vFpnpGH9mErrzLlSrjtjct7EKHWN/M7Q
440d4XOQDM+tBTVDEVllqzpA9oO6TyjTRQ9Nnhj8qMTV6yw6murdo9wQaBOD46hYwMWDl5W0MvxL
CnJSytKou61ysJeQt57SGKcq4UXjyP65ixKAuqO4BxDvyY53cQ2mi3A1cvvsTGYebUJpUwjoLcww
riptSRsQLdOy0QiHUf+2yvXETez8t1VJgpV2raJYcCi6nW7TElZa/lTsQ/rmPVq83NrFUMwfhqsH
E0/SGbiH765Jp2cOrTU2Mtyu1UsEdNzP7Jj6opi/R5jwofGC6bkCvkoaoWN8z7yh0cYMsdnLVtS3
Fz5eKmStXrk49vX2swS5PaFyEge06NS2HwxnmFSIM9aukPiwY+nh+GosAsApGC2HbtI626l5gmP3
NB5DLoMUe2JkQNv8T+nGkecn9ZgLy3OwbVaFo1ewZlMaVOLAmb/Vrw3+uKgfKi0V2twPhH8I0J41
D1jgxYKappXvFkSHAMeu/CFe4oozy964IIvYQ5fDWyNhxe8tI7wpyebkuxTMQQIK+EgdeUdRRoAs
UOx53vWuyZSp/WUIyRW0NDkfC9u5nrO5JiiM0FvY7txzT4NggsCK/yYPSK/xF5oj//O4EjjbK9W9
Ib9gJTCuVQuge/Dt+vCJXbUtiY/yHzlRctzpQMCVWslWXUzMNuJwDUzbVk4gE99WTL4mX/USUyqY
u0dZYLLG8xEWm1j/K/shHn/nAb9UBxAXHYsOBDS3BsjNyyizMjxN4ERbKcvsIiSaMSudZCtWp0Uf
eB8awo8k0s5Mou1q7EyNI4BADw1PSOcnQBVO/z9Qa1F7m7DaiaR5gS2CwkcfQi7zwnmvY69QQ3/B
cGAFg1TZC0js2UQK6RqmvfiS8zBv1cMbPJyDKomMmo0cDmBGD7swUc5o/bKDQhf9rbvTNsghvXG/
x0ErMd1AnCt+XkWk9sJQJvvTf87aarYIhhELkeOf2p9fgZ5bkVNANXTh83WmCUGLZbc3Lf8dGTRm
8CGUSaA7OUWKglpQNIRVSv6HD6QUlAzI201tOu9fgP5Olq1E8Y0VVBv3NBuIUxtcHVCBRKRgLF9+
6s83lMjVgITvIXwD0D4MU0uGUrg6g4V3D1DlC66fYCzxgNWfAasBJM5ewYuWWHZ0VXL6gbFuNEiG
V8fyPeU/HIY8aY/r39VzhHMS7Qi6OEs27yU3NjcSAZ/RyqRlr+1jsy8bjyhmRivLzYI79wcqs0x+
M8Tn9YDYvdpcCf5KFNOCShgH7CDyS0XF2xZU4aSra8A2cyzxWHk2pMTb1By4FUp/xOjMBGPhLkdO
ocX6x8niswuytV8EQSto7zK7RisOI7SXGAAyAcs4jNjh92KbGkjVF814ZQk+sy6DFffq7JcqqqPu
uzlZDpmAqjbRxhJbT8Ucd6i6QF+9M6WmhpeBxeGncVFkbwP5Q7mk45DRw12GWQQQQEIQtrvk0Pvp
ycr5+bjFbVVtpQVXMMTH6v5JAeZAdzSHmf4uCIodQYbUGPfAQsk5/kjSjoO9xFRuqT2d5Dhg/P2X
CoE0O5GkZX8zzSocNb+3x3mql2DexUFrasR2lOj5c9IdDrIbZjP33WbnrcwqixUH4bBrhFHCB7ns
jPVsDiGlij0dIbMTIZY3VJcAX5gF7tJNDivO/AgHgUT+LkcJFMnMnGzzmdAWRUuQeixfeDCDd/18
RcfE+cCRY4umHphWWqNRulyZ4y/XmfpdEPewYwxPnsq08rPdOLSQBIeIr+ke4Ip9yHArkrmGLv0j
DlSTxciMGSNhK2GU7xx/XTGWVfr4ssWYjCp5Y1z/CBkaG1rVL1wxHA/lUs8y5veoLwYkgipSXbaf
8D1uSfeebUkDWCGZpKkwi+AukUPnPq/3Bh7oZKy54XnRNfVeutmeHsdXOwRGUaldy8RdHdxVaEzn
we95nlBvW3Tg1IhKixhUFcZC9zJYlLS0MMslKTAJ2gCd8PHM1+Lg5kgeFUA7s33rFySf8JsFApoj
oUh0btI/iRMen6EpNyYT5COiJtf/g1Nt0wBv1kS79UZ8+UrO2hCqyUc4bNoaIhkwy+Ot27wHw+Jg
PMWv6cMGBZXzdKvq66NTPWB96XEQ76rX4PnV0/lb/uL6dfS1rG6LzGjVi0ALpgCDwbt/5wwKc9cM
qmsMsOnkMJyFws6IDnm56B8Y9MmXpfpwpDQD/ikS/GV21uKicDKakurFj5XQsT8kJ1/HQj/V5tFM
guaqLMhxNDqR+PFVEZIdiVTNx46N7OlqzZK/o1HG/9lIpsGw4Jo2wIEUZ+tzv26Zy98KFa3KGd+e
Me3FxWFpcfJo/o+Kv/rwwdqllaMMCy6QEVBNxiVYQMK0KwCzOpsjA6SR9dAestQAQ6eozzKRfsVx
mPXRG5y3pCxvOAQDX2WJWmHpaLhDdSyU/16mx1rWsoImNbBxuFUEygR6iUiQf40o1MOTisJ99uSY
3/b8C9vozJxNA+SOX/laSGCOCBaJkzIPHD1V0nDdcwvxemlqYBcqOzYi6xWgjWTS9Wp+CFjsBkYy
IWCnJDr6XM3XyXSRrrQi2qAVPxtCzY+Ezh/eH8u7wMmS0p5zsyrItq1ldbcp3TaxDX2ujb8ejx/I
f9/ME+ADqi/27geSO5C6e6/rEaaLgx97Gbx0ZZtRxq7Lv7qWSjMsLGEJt8Jjq7CqcCUWCHwkqzMf
vktgrdT0KBNBGYAwfbxFfZMxaqOcHNRAbS26vhnWRc2u0G6PbgfU3YwFEfVt3pPyoZK1TX1tOwe4
qssLuhFmocoNBgwqwDUAQgMMEUtu4RsM3mqRgRxXiTtZNTeZrehsnCHNGGB3zM9nZl2tZXUl6pw9
QoHmB0ehDoAsdbSZf7B11BNkw9ZIYQkpRkieNENiLuex9Ao0rmxVNOkDC338ZTCLSdT8xmwmxpey
vPPhl+9VnTV70I/ztbykRQaGm6snHz2BuZ/BFLCTd4zgKS5qcDc/7dwAMZWQHpfmq77hyTspdIRf
zoMg4i4FPbe99I45lxF0qyoOW4ieRKYzsxWESIxqwZmoZ8uSvTA5Jx/0JVLxv4ZlWohwbXmiD/BE
3RQm85cIQPiax/zj9XxVJf3fTp6gYTsqwoxwBL5nyUA/mQgqbb+yy6eQEJ6sFhjLXR770unD2WbP
F/IEKVW8JGy/2JWrlUwIwETQhNQf6iBVisQ6L8ZuX5RqfIZmJVxTQIMcz+4MmaPwELLCyBmJbAaO
kHnv2rhxOK1omd8+Y0T2RjM++Rjne6WRLQ5SZPyNK2YcpH20YjQDLWVtO6xPOqXW6SV4+vr8GleF
poEztOU8qXWpyDFpiBnHhdj4Jh+8K8c0PCJe01xpM9L+e7rLhFY1lDMuIIZgiwcUnBK2SspyJ1hv
JQKZIdI5zwiCGwyRpq+o+t5T8wCWKy6unAfIgKhjrmJw1AcS/GSPqA5VMdX7HP/y1bRLUV2zAbdo
Cinh8skZ9oSOY85A4deOjsSQkxe45S5Ql2NR1hIVY7ELGK37n5xx1Ds+rUFWqKmXHUeJIhg/Sg+z
fQ31/R4gm/9xQt1BeW+zNgaHCaLblD17K1IRuBUXp4tvvxD7KR8LBWAARU5nkxzx0x4A3mk+IOk0
pNFG5NoYP5qdqhqoyjrSRFmWPWEdu/l+wZLVJm4/1FBy4rjTOYPwz7Pkyav1S9P9657qCghOwbIJ
JfDeAoDUvlBSiq2mUSnUJBbvEs1b5P7PTJMAaRvcStBBvK548/Z4SO/LdO2xf+9f9CSduWzJ5J1K
ee8ffHXG+v/0CIOKaxm5fzi/8yqGaQi+Ppw9dkCHBjcPBsK8lsVObmZT4xQNGJQuO+OfYVX+4P24
Nvt/7EZCIZPfDkLFGVqLxfjzFfGjE6wjBgBkGmJfgINK2x+uRFv+xjxhoGhCJ18dTu9qRlbb3Wha
MhZ+2pydfwHNaqAjz/z3TwOAjK9JWJP7cNZw+WqSbWpugCs/XeufxH02zlnYMpZ/jsUNRQWhufwJ
DAXXFpuW3eZzsK6SZFaC/xuzU2TMR4X1qRrKt1yF8QW+kjNz9W8vwyE/lYmCXrxtnWTV3s1S1iGB
V5R3o1fM9PiTKXA4qMBq6H/OXQvMJdwhOwJhWK3jeBaKnoebTVJVUu6VhjzFxU4JjggH0+jA0gR0
txjQRyJlsy1YyrbTbZnn6YddxWJ/tKV2OSks387CtYbgi98vd21n5EUeCCpR0aLeHqM5dFAlIxV7
CsEDLb2y4iZuq3lyi6e2YKdZ9ZN2dHCzdroQHz+1VmrH37PbrUciloO6yLmysgkVPUtMyhFwJ6+H
fhNU7Mtx8SLevmGuHNGGgoDzZYcoOUmB75govPyC98FScM22xljAmLeNivp9ttyzUDY59zzD0b7C
lMz1E4w1KKYZRKHY9964ov+o/r7sBnrXoiT9/T6bm8CV1qvR5ZMiZ838vyzmE13jKdMDYGoC95eF
eT9XjAqU+sb+gSB1c7d2nW/DyBGY+WkGvXaifCNB0KGC7vUq0bquPWilPwRcO37u9EwatbTGtWQY
vLGkOwlh372mHNium4jPy8hlAeF7xOENzvAmEN1jy5iWEmLYUi2Ed1Vwz+sEnalYYXBDh2RkmQeV
C68opYlvMXdTMN7N/Qa5Xp3U3KS1SG2onOpO6kTaNNs3uZLncj/yAGc7UUXoJNXhP4fECmdNLdVq
g20fHiOZTMuewUbYs+3d91S5x20PL/lkv7H+uvg5a50+uCTM0qmyWJSG25y6kanDhXFwTW17rsOY
Q1vgiLq4qaCsI//lxdaDD+08ZytAI3UapEBQOuEMP52B8VC6L03D0SDKGRZuiY24b7IZ/6zvMuTO
6zDLLBibNY36gKycPYAdNdrLpb4tUmvyvn9Rr7tTJqY6g3zWog8YKb3NmXGS3Zdegcj3wM+jJPpV
iY6H4AKsBGpGuVICCK7WaRjhdO4hA3TbtdM/a+JQ79FOkOF6Is8TYJLF5bCNbLifgS4YLZD+5JbK
kF+JWxF5OnwZO66WKwILJj/u+zJ7Z81NeRORJHgfCDC5cqjcPJN9XbfqCRoM8R61eu7bBJi0TLlE
AFP7yI7+u7U2jIglq5VhQ20PliF7J7i0ArXVE8yZ1+42MX5m3JPUB46P6TaHJX/P5xiJUSYqWyZi
OvnNbmb4DQoCVbYe7sGdYd2BlzFk9ZEKIYJVIk/z4h9tOSCjHw8NzZssPkw12AIPK5h8cLN46da8
s3YOntzBJXk5XYIVUeaZmV6EQKy6zmbGei01uFihbAsvFuZvb/lAMmbYMDTsUrmgSJgQ49YxI348
eEQyPjiiCVpKw47YuPfB1ja5xeTftNYMPohAxqDvJoxdy20n/nuTmsVXbm/sK9FrLgq/5YtvNg1D
HezXVljxGN1uAUQOYV06+ePjMJI3Tcl5xVNov7Wpq9J/fE0YevPSxmw2Ed0ufrlumy1IiFsOpzKy
LAJvTKkJPPk6Z9RLcuieqTtyv4vSEylifSpkTGROy6NqPDImKV25vTIbSk5GR8QjHeMCIu8FEaut
wrsAQg7yGwMACPtMAGSm7JYBZfvfXTmU4IQ4lsCjGO9DaPPaMIw1Hd+ZyzMtDrs5zhrISGD/QaL/
Amnrzt8STNUgXWw/pPao2vDFwzc27aNEpuHlTqVca1Jeof1EOWTax/YchASqWFiEOJVdjY/JfM28
sPMCCZf2GH5bwKMd3CfOwZ7n46+1wvBq30fodBWkwG3pryJCM2qN9xztY3zHO5jK1Izu4DZDOs7H
ix2Qy+clKnzuAZXWJNBoWhcPTjjW35ZHmdtiH7OWTYSnXgeSiODpaeoInCZjgKdCyaTTu03provn
0whgijsKb+w8FgibXJ5gh19opk0je1AxEgZ92ZII1hKrrppRw+tWDXokZG5jGURVJjS3lxkjs8Lg
fpyzzrBpzMLFP45hSOeHNSpXydk9YyHXb46sEUM8+SapEBb8LIFMYESMO7HU2P/thmA28xVShlie
t7l8WJX4b03Nb5EPJlBukADZChuPNVoiDEdoQ9kYozAKqMOXFjrMQK+UjGyuv9rD5rNlsOadRtDw
G4xYKWtarqjNXwOBqnX13+lH7uIqjlYLWeulQsUcBgoLGsMyFpgpcVir+ShswuWo5KN0TTWlDXR4
azva3vGdaF0v2SJLTFV0rYutibgVMmI6PfuWyTAN5Qih8wzPxN2gr/fyHl5koPU/WjoWKQbXkD+4
I+yS10zw/oj9ZfUfahDdK5SD1H+rjpaPxMnp4oa8GvVuhsiBQ5NSfccCbpRrplxzChZi9DNipOl9
aN9WlQu9Gmg45uffnr9trX1ujofsiqd/fhWEH5lMGM7W2QAQlYQdwwp0FXpyuszIrPsBZUIPVuXJ
K2qfU8Ua46RqwubQhBhP/hRY9so84ZNal+RcvJtsuBeGz9oBBn0NJ3R0gKlHYXKLDUE2kL6rK689
bUQPK0th5IhAfALwspo/nYNaTbihIhutBuZnyUoZx02efjTeTrojxCLGnSxt8xOKzMw9YHyfSTtl
CFgONMyKm4NZY5uYVENXiU9RVUJPZtndh1Qzy8h9Zq1BjJSPGgGNQGkE0zAPmgLqfYGuFl1BU4F0
ehW4yIfbd29oZXs1YEi8AgpvTEYpn6CprmN4+DRVtDsFndm4EU5UxEm6IGYAv8aWaRQVwGwKzTMN
YovkFs3/QDEEcVUJiHvMKLXGTwrQ5C6Hu6YfH5X1qaJRt/lhbwTAES9xvv1G8WsUSrTYzPW5Inqm
E9gvPZU4ZSxKMYLZIRepG/Klb2UaNrdUw92Ofd2sHSoxhkprt9Mq+W2ruYeWW4aNvHtu20xBPMqy
OsgS9u09/EAV8mp1HcfLtJLymu6gC7rXuZrC+PJlcG5e1TcXFgJKsv03QZm8zy9lKlT/3ivXvdK2
byrvO0IDHZnGq4ZDV8YmYiJtYjb3qrnaebhK8Q1IpIHJtYoRoa0x0rLQuMZwypLJajDQ2rHE5plZ
ntQd2RL7sIOyfI7LsbFO5WGOXueZz6lneiKKCckZgnLmZduO2fFIRdchne811AFQCQq5lvRnmj/r
Bsihs1cTzdQKepLsoIwEtGT2e7/u79qbmjJe8Gx3Kz2G6eYp7BsgEPK6hmB2q3QUwTrbjF2PtY2r
/Elnjzp/O2ZRmAqfbpPVsO5pY1HYU/vq9sdKFUX1Fvb18ac6WxCSS+G7rvAcFXSbF/dJ7I8eYzB4
4xt449G1OybJQI3qGtQmlRW8iFRjZ+dfOGcrw57dzG7HZpnWocOZJNfVB3CT3W29/8sJGrr2VmwW
zir3SEcL9tVpfwuiXZqeOoa5BQOGcW+wYKoSqBG7SK1pO0Hz/0f5H1sUeeXlKX0rLHT2Ja9mjVzu
JbYReGTqIQ9U27QQLEJwucdFfwDAbQKmHZLa0I/Nv2wyFAOqroAPedHyHp9eErC2BC5EJrQIMxe6
r8WrxzlHHlmXF5E74+4HEAK+RLbUatHpb/z0XxZ5gBkHBLIK0G5ABTBzny39hkgyKUVHlLQaNSw0
BoEXJlOrbLHzg4T3xTws2rJkfPdY5YKOcEFKf1BYog+fCyegtGPIuBD/ZYJGXyBvSd8k3TJjvxyV
UTNKOBu9FJMVxrHL3j6K6e6FG85gGqExqW+R1WnJiS1B1TRMEmPInuR5f/7O7vsbVve6EVMGbamk
lpW3q+7xcOq7DUae/bhfIRU5IK5+SBay7eiowPnSy1akDCS4C+gjNBug8afR1xjDlyzSE6GeLCnW
7iuxlrF5kAeMaGcDJPOIZfIHrbjEQ1Im+GhoOerQVDQYGihliXFKujUzoG8vyxT24spjOGBGwp1n
0VM88YY8Xl90nTDlmZd8IyQLImXWK0CeEnpXP9iUjnJK2jHaQHZqLmQJWaVyampE5I6W01H/NTp9
h5HmS0cZCMr3sTptbZ+usn9ktYIG0LjyHDWX6+NuORryFcRLt9iJP2jB5usWMbJ8H4eSahLoNIHB
E9eVok86VesFTjiO6Kl/zgjLT5K4T/XPCazGxwawzeNffIBUmKO18ptaocjSHja0jZyIXWBSZLyO
J1PruAmwmdCyuoRWkOWey6gYch6/ecFPL386U20QaITaNTXsy7J1AeUnxgGRnFJB0jIHQxgEK+zN
gB1bI8kofZazBA0k3yj8gofjJibgTOfcGJrjZsak3rwkHv30SMXm1DpfdYlRQ0YI02oGu0TI6y2R
DUs6l2rTgbvDozaTqROaQlLNBuxoic41UA+rjlUylWQjXTiWpU/k2sPAJBzs0uMIvQe6CZy5Vkxz
9PBeCMgDLwp9F1XsywRERmw8O5YFQSJZkTS5XOuy9mKAiYmaAjsP938Bo4wGBuRCcc2iKrcstC30
sESYeFPVrn2ZMQKhTFWuKO/58O5gYun411nXaXs9OiVxoyHBHdL6Na9BTCQ8fNKJRPFCNfQB3u5G
vp3nYLjAFAf4gqKzU0HNtVtUVtBkAzlcRiC0sTGJFdXTTzlz+28d/5god0QyRlmf1F2CCG6ZePcU
LyafI5CA1wtijEvhvmrO8mQRhN+DWck5gm9n5XGpTNe991iXiqf1AJX1mKN68IPYcFlCY4Fesjy7
5zJKK7C4wMrdAYUow0syQrbLJsBWqL4wmfPhFbp7kggv/+bTuUU2/uNp+j0dAOaFRycECA1CA9jQ
vU4LV6kMJpf3unjDRg8XeHvoJGeTycM5+z9ztPjuSjZzfzEr9nC7ZY3jR+UX2wbr+Mt3ssbj5K5E
mrd/gpxKU97MAvO6QtTiXg/qgyZeypZ+afpCPe8/X+Y9CA49Xo5sJ/a7i8ZFeIhu0TDCqLt71tfq
2NH0mnC8nol9Y9tAPiadzL4yoNc+n5StZRf8RbHHw2/JlrZjUZhrHpG3UXmxOw3I+/tdbRQWWCdQ
rG/myvgjwCnThPKwfLwS4IY9vRsWlSe4D4iVPF/q+IzlWr00oA+QvuiR2NTsvds2vLvrX78Hp51v
MpWU9jLvUJ/1k/y4aB7kzrOAyU3AL69Z7MV7sRM4UiLIZcf6uuf2WhASwz1M8kvxJw4Lr5Ojv4xV
qRUc1Pf4NjcddfBig+6zL5kFVVEuNUWwxMLvOhwmLdcOFPGZeWx82I+HZ6piuS38qeS93MFNUe8l
H8mF5TGtaQUraD1cNQPHSEk5r3uQy1Hn1XWDdlhE8jKa/uQ2fngqxsfWNsfOQNBthHbDwMm3XJ8C
flJ2WQYaVKl7crq9I9RCMBlghz2cV48p0SBL1cVQkQ3lOqsg4IGFlgeIis7Q0P2bCHPphKJiGL2A
f+aur5gx7cfxJsUw5ebCsgRrQCwKIMWYAnkfHT7xkzGumiTXH16Ve7WCwwkVuxDBrrBGi7ItVb3P
EPSz/VzrY4l2iGFTkXXbwSSOux64jz9I7Y5zkswRYbnJSo9Dzz2QS+tz40oXfbvQawqjuTzG1YJE
F+Ab+wKJF5gqOnMimpaVeBiFSdyK8qT5FY0N3OYrm/MM8YqGC3GPE+iAOTIyOXcIDrCBx2/nvCNj
UA6HvcI4cTpXOyQogsv+jW1IofoYYeicKrREPTmSpcvi9ncQN1grbutHTSliQlTU+f6dslH/mt+p
VS4qzT7+6mXXyM5bItienjcu+X+ZIR/HTFPSYxfvVY/oQ+ARtxjGTE+tQLzNeJA+22krLWhth1Ob
GDyPkX8acRpMCJR/wJqTJzGPJyHdFUvk7xa6OPLYvG4Kco0FHx+peefWLlGYublF2JIeGydFRc6O
zN+woSOyX6JD7qeVv0TeNo89xPQoetgD3MvTfoXutsWNd+PJ/7YpKtPB+Mefqw3uGH1heVdCn0G1
QSR5qmqT2mXcYWuvlkMvMVJZ//zGtPZy4KfY3W8qrcl/RrQx2XLFc68vbKWYOLxgFp+/2y/JtAHC
pA9EzPFWGhWu3orcqPiHD1mPzHUl5gt3GAqXBm+r+Fmuye2LEQvqqQSOyFnZCOFSABJlGnoFlD9Q
IjOJXFcxVPZs4wwc7//q9coNo78ATHN7GumTdOyRxgcJGY6fjzf+Nlv4BUSyCYygRWNogbz1Jz7e
zoUwWDdiAisbFBWeXkGkgjYN/jRNqYzey++GfTpbaadffjJ65VRtZ1KEQv8uiOsyj9Xbhe/A8WXe
Qv04F9l13Ozreijvu7RSudZmnvF7IONfk4+Nby3u6rsinn8i4FYScNDLJJBwI279rr9PwdPZRrvh
tGH9sYhgcIwXIH6uMImz6QMN/l7AYOdS2OZy0NyQfwkhPyMuQRwqNhrQsbB/3IVZuCFKa2/PEPgZ
I8j+iz0L/uPv3fqns0LxcQI8qvASZufeNEPfaipsM87atoCXdZAysBuTKlDwiEKWEcvS7/kzyoxo
vg3PTmeS22poKyyv1+oIFHItkAUdHxfote02EG2jiVYcUICGAvKF87qm9LT9+Z8VKOllNf8QS+rn
Zun6/ZCbZBAIUYu9wzoffrpnkCOo3F5hX0pHLJP7p8Exq8O1fTGM6Sqde1cvW12c/R7T35FpTMxW
8acl3s9dyJ18u23j13EFN2rFNyrG3DeU3YkfzQDNi7uLJaXUAeMiYwvMNg6MPm03hlQH48THeUGh
0wr7hMZGQVCNIDzsUIQiZjhgX4PF9i4+wT26O9ppV9gRyCFQVYN4mb1QgFWMQdABsdvmE/4/TDwu
11az5EKthmEBpJz0YbmtkOOUdKojMi1cwojH7hAFlFxVsqkaTf0gwgYdPPvtWVTF8BLyjIwv+tgf
2jYSxf9hu541eLqDfz5Tw1ywbrzJHc8sXN6hxsJmrsVV3ols+EhEM2nQQOo5ffQ9M1H7TQu355pb
cHNhpuQLSzf4bMGYbNKdYabGY1WA0pwKVfioJZfVvV0PrMbvpX/gZp1dwMjcqnb7Ew/pmZVyf8wh
l14vn1Qoer2gfJluNyQWfdxlZxXYFYT2IAUnYqmjHwvZUfvJVGdh/qK/HXfLorfBEOBWj4WUab2D
nm1RsIRbeRcaXHLwEKKhV4i9kZemSuxKO4wf4PUMi9+ptC8agLnWFk/shNtGKBtYGWH4rKR1ds28
sKuYq2wzTD8W+C/mqZEhLOV7AIVoWx/B9kNKsJi5OgHu0rOdh8s/7QR5Li7L/mXd6UZf4X6b6NKM
XrkL3L6Yaykt3DqXQg5Re/5U/uBw4MLhtsCK5+dsX5tMvCf8qtxCyFItlzefb8eBSU1Pqvhd3K4R
3pA8sd6dzwpw39gmm2YcWHU0c4G3zZskvT/0/RDXFnWP4i7N83m1P0cX20d729nteGBX+1Jw2jrR
adTg2bO/xA8Esg7Mqlaf67uyR/mlDKcFrvdgJYw7Dag6DgA6ToIVJFjuFviw3IiErMDr2geXVJfL
/svTnWx4DQzaqRc32zz7xTRRKUII+7H5MWSZM3NTjRE7XkQN8Wy5CiqlI3FJuCa9CKSSlTycJe2t
LjHpFGqVOApV9DYlnnqAJrNj1/CfD/OZ6pMOKWUxg1fwiaNZINSWqojgNJXas8YWtLmnZOXyEW9W
hsKV758b7C8FzMkhSX5CNntpWVZjSAThla60fsxcjlN22kVgUybZjGY572ReSan7EIUlkMhh2Ppb
S6f1Skh/koaQ82Y9epeTSCO714T+CULHbSCjoMX2q+NcqNyowLdsceZX6SaytWVpfXcX1ygbKLYT
8pAkf5ARfi0O2BUTMK4G4/W8Nb+IuYF2ZuhxFcVzjky5qWpXwVljx6ZItUP6/5FSgTgz8ny2KpJl
zA3D4OKMY/D+lnc6DJ7lCVaRuhYyDwcxnu2aS5tkJ93aTY90COtwPJjZiAjr0maqny3ag+jchZWb
U8jRnxXOCah4UucJSx68ciUJg8n8v3SbVxX67fQJIA+ZEt7GC9Bbuqdz1cy1KzANl9iurMzmz7i0
GJKnKIqTaw9vuCOQPrEPecsdEnSjjM/Fvpgv+A5v86cSmUqvcQbhgRjUkqkGNsP3qAlp8n3nmjaj
LJ7YvAobLCEgwLuh2D5F+Z7Va8Ja1WvArA8hmF035F7t0+RTo9U6mZs9+9tmx6XLi0xE6O16/fJp
gvi0A5UJyo0aBAsD1307iO6ONoM+nZhohr3/O4jFJ6ScuD0XEkNLmigoT7NBjxeaDOpHEu6TlRHA
4M+b8M8FNUUr/yj0qSZ95Zzo9/HtCzXCNA0HOb562geuQAp7sE0E7gDBXQ7UWPNIJw2dCFwn0tk/
hXREuT8V6ipR/gxJTHl95bzrNkMc4lxyeyiv9ZR5T8ht4in7pajNRCKA4YVrXjwlX6sC5Pl4hWRF
9yoVRVr6QnY7rO0JP9y+7mjmoYHdJkkiMluGiQoc7sP2iObz5RSfXedEmPokhWgeVjsmjSzI/vev
rfk3G8nVEAmzIgsFHNaRQ8rfkF22Ew5rNh7/bMnbiiDBE7KHTxh1YrrMyEPiIdwSPD8t21cxJoZv
46jLlzJ4A/pakDKHyTVVdUXyKTGbZ/dRUI2A8SMRktDi4f3BbXQukxQVFw+JMapjPqPyqmgP8KCS
wJHPv1vL5Uv+3WfrdzPR5yHYIVECuFLfjA3iLBVMmIpvTDXWc/nj/5WbrUWRJVCDc4lJev1e4aZc
mn6rzOx9UJm5PBCPlWxC8NZyABev4uWjtRdWmunI4XKTE3mRmu05dvSUhP6VVpaOBZXIctqhbKvk
9dimVQmPkjC0pmiHRsSZ/Wr8aQ5SeHkF9Om0K5wjIE/k01u0vVld63tDGfR5P0I5h3cQMsDGHx+s
cJQGGWJORUjzL/DeHEzuHS51Prc+pCAUL3/RN1WWQm1k2ptP5L/F1jFDiEs5IZK5uumGt/YfUyqR
6rxIMZ95bM3Q0PzIO6OeZkuUxq2mqbeNWWUil0F3my3UY2S3JmrS1WOdtg6pIG57LnpOkhmOGWAw
3xZ60IRAvmo/9R2k3xzADbLYZ/O9LgokJTc4+ElaFyyxA1L+uDzNfR2N/6lPKO3uWA+2lvUnn9Os
RRm/nhnTrE/ba7o7UzdVvyVnjF3pFukt7D1kETUMXwmoehQr17uMNJoecXz+WrV5I9LBwmZWLDNm
rBh0IhnOa7YRezuUPj+F7ULXVmx05n5/1TxyLjn3dCbXLdFaS/+WX6poNFod2yxtYsa0AQI+7YQF
Y4pfR2ABFaGNpc3aAmG4kgGTRvw0i6kYJOtSZjiwzFq6jXnwp5xby6HjNLowiHU2o0Ipq73bx928
lonGSNsjCNDBJSaqfFOvBcPKu6pF23pB1oBQbllC3bzlpBXRRinzmtuLT99c2cZRw8DOIkR4cD9Y
zfhu+2eszv1Z0066KgZEt+jT+aQMBbUXpp7jv+aiifgSSh0hh4dTHHEMDP3efhQdWHc0qz3LrfGH
2sxIPHzJrH3VGe/RlFqs/Xs6P4dG6MUwMh0mJ5NUUbFMrKO9tj5U8cEi2z1S965ZeXJN4nwM+cWe
4nH2KnAPwS+K8X/ksgMXkvOEiHmvksA+hpAn5XojX1P+j94+xGv+wz/NPSZGRq/LTKugaah6gfrL
BmaThzVrA0Vz2bpEWg6089Y0EWcbRebn7ZiEnFy/z9hU1RjgCfYKIgjk/JvR5RtOXp/SHuvvkmTo
SmUnQIhNH+EZYKe2kpoWCPDqjL85BH+W0mcPZCPUX5pANsoXWk2A4WXp6jlUs3fvGWa0dbjIjhSV
GQ5onSlJdSsed5rg08fwaezDr8WXK1GGWwdqJI5+57o2823q6n8i87clrg1chNB8P/Wjudwjbhee
g2wniVZmS9EVv7p8bR+fpq1NBhbYqvmP4yiHWKlTWiKZPG5xZE272j34BiiPVKheZZRnc10pElnM
OsBy8vQcYQ3S0UYR3nyQD04lEw7YZp7lUUsnTmH52kWbd0BCTOHUvTh8GydlKlQEIqz2cKh2pcFu
UGdB0jPeo3bMi6+NFNP/3hpCLtF/ykojWRVjSYCVnoh1M/M+rHpDHD0iVbqM43LfTrh/BSGYPFnO
jD2wBu7BNqNSWyCMjFruqMT814/Y+OIc3l4/VYTNyIYYVdMmGoP5pbbdlA52w6ryMFJWVFoivx00
UCvePMx+f98cEStIoTkZsw6p7LzRVQUyjTtKuh3BfzXgqx+Cmt51Av+frgjPmv9iieTm2GHIoZw4
FrcBvWnCWx5n9slvO1Krioewls1g+CAxAwPyVh0gjzfjhUtb7BaPH5rxqV5kZzDp36fyTAdrRpdM
PsDpL8MAzwLXmtLvfKApn3tWs5AfiNJ9fDIWYXehgYdygHRTBSXbvo90wvr12PVi0a6jUbUXqkqf
WQNw9IRJzY96IHVmC9cVMwDsNWz3CX4V24x5CvK/YIwmCEoiY7kJgdP3ZIxqLjc8OO3eswPavl95
ptH9Aw9u9RzbE1NPuCxuS0hEeu+RVOJ7zwDvQHsyErCVYMHPiDwAK6DFsc3wlDr83ky1K+9r+ng2
kqRdrCf2RMYn3DaHY/4MVi1Lcc43ht4QpmVWR7RKOA4L7NyrxVFV+RN3oTX+9WgXyv5b2fgNhlC1
4J1/kdtI51XkQm66nZUZBaGC8kYprgMOUyW0fR33hwaJ9HE1AZC3zZ4lJEzAuxP/e/F14+SACEri
FqRjBIQ78vMQVG16BF8aheukeOXqTbUzTY5tnrZ7sTMCNp9Mjd6rOaKsROwaa/YDbS3hIlXbs9WV
9ghtnmhw55ldyKmUL5evFg9irymAtPCBDWmH0uGewmtqbkPtjKYuXS2AXeIPngpT6Ti4PfE58gwG
lFBITi/+tpvEAa6vxuLBpE0qimhxyMngwPgUSkHGBEE3i6UZIJupBvmC4NXimMPBNRrR8brersNT
t52DVuGMczUXb+NPmijFwdgBZNsaf7nWEYx0FALcPprOGdRfkYHP3x9kFFzjso4VzeXdHnryZGf5
xuFjxL+0KachJGKADnj6KOTAbSQxnsbK1YV+eSWHuJQDZ7pOKdzMt5wk/Js/zVSkztciwA2BV5TM
dWzeRaF955/qQ4n08V+TFrDHoXh3uwbMjAmqzoZnmuKUQXdxJENshXgGiUSzSucol3r4lU5hyMRq
fT/a6poP8FfQ6cceIB27owmoKBgP1ecNY0mHXGHD2SZIFp/58HyHKw/ottrp6COKvYACYC4Ds6dL
YzGPmOa5TyBGWaLy/jo6cvZv+Jk4hfnKNkvKlblXP9+vDt2Y4YE6ZSQb4iNF9xtk8Dn8073o6f4z
TcXVTJjkKXxnEgDXcfFxhpDPR+taMLixMhNmKSmU/td1mGSPkJyvpg22D/x+QrEtR5yTPOQFVsrC
R1I4tVMt6NRCyq00Bas8sL+lzg3X2D6l62cZWTe+00aOtiUiPDZaUm49bHqhU7TfWXj08Eusn2lz
GoNUi2lahilfyGuvWGwDuOdOgseI088lBZTw2OAKzaxV2r0B2QVH2bPqJFLK101wtxqhZLESCmx5
l2BAI1NRZIZmziF6btsj326ZIwfq7eyqBqJSsug9yuPml7uBAK6AZHWRIdzKUrqgpHEiODZh9v+2
8lwtuBE9tT3HsBasen05+5OouC0P2sy4G8NdvxvNGNZT6n4ir4RBoHkVsCpsGV1jpTmnPxNs5Sr2
IxnHINCpHczzXe6a8WgJ68DTGhtq40odTehtjRP0RhsH1BaOYHN5KQPi5b7ZtJC5PEsInMUWMFnm
6M0MX/s/nQemD2HlDGg8gLIvLuFdCTdo5DSt9ZwW0YTwHXQgHdJaqPQhzcOsHWhXWMGA3Etlzfqw
7Tj6B6UB4z+hGOT9doaq3gDin4OIGoOmwyYcXPKn2EEwvVBZ9vsvNGi3iF5ylwSsnXTdGHXAi1S2
93FtfzCpRz8mGVdgiV2QTno0UTkJruPcEwOiFTILTA9wWAP9vzAI1YlwfFWY+v9muYQ3+TpAwJxP
4YeD3bApHtqQAiLKbi1nWsgPbtoexg+WnR3RVcA2QygorXT2n9bTCSWNr9lN8GKvC5XB8PFln+dX
PkWvWEdYM1ZF6IMBF/1C5PFnuJNbZh8RSyUwwM5dPO5e8SYLv5XjVSguYCs/61MCbCBU0UV2Gs7v
xA/PuFGtrAQesvkuNfUmbmpl0lt+24c1futFzyU97qVj/utDYpca/7z8iuU59TK1cVmTNSCm1PWo
s8vob4D74S7ftDyeT2EIE1haQM6vGaZT5R97w51B13nHbknlG44coCk4YydfpF/8uGVcT4tGxF0H
C+f70mQDFyqLDof9GEIYeOAr7WE0MBGkFbDLEgaehn3v1gRK9k/O10SBmn7vQYdZxVOtP1QX6rn/
ztcUe6cQCtSm06JeIuQTj2eB6IZMV9WybA4eeBNeFZ1RYhlziaoKLcQZ8tII0l+IDZjsthXZ8u6o
gNAvFWziLMK5Y5HeilygWEntOc7We3GA1F06v0/ydAS9adIloxLrU2TuzJ+21TxaXTgxd55audn+
9swImYKYUIuSSBRMHj2ikZhenjNOgyZr1/+JgmW0htjGmAqum/ZE1oIHC3HYu/MQx00Jfl2Vm4mJ
1z6HVOu/8M7d/lolem/v/NQK+hZ3TI0Y5ORgRF76d8XQN5gsO+plvVlIwOseopNE5zeQw16C9Oug
Fd8JdOFSPLCAZDVqgGisYo+dJ/0/6ADx2/QqN9i9Ll6np2dCCsRKtQH34+ewzNhfyMFfrGiomCyJ
2qO5osEV1VTb3YCFMIJC0HWmnWvX5ySsYzWlul3qdIxwHtgfBrUIh/qZC2t53FlOrmhtZ0bEtgTz
nrd0KzQbhZyhlAnVHUlsAxwly62xyaDpVpu8eaFEgspOAnnHGJh3odY4btjdk/161nUU7ECwHyr3
IELJUGGDhgBoYkRqWdmi5mYMIxSxXJdEW31IvuFjShnWmBaTjxI2fVmRfQR05hSsFJfFPKyHvDJ8
80i/kL+J8VTsxxirQKtSn3aaD/37C7z2z3/AFLePcgpIft/zUKhdRP9JUVDfBHHeqP3zMmDtFnGh
oiZfXVrP+gqgt0A4CBIi7syUUqs9+1wl44+5K5+HQAkjYbxc2CsAjfylxiSmDzYTx226kpsmAfZc
qi3cKvFZ5jlY6i4QvSNOIfAmyuW3qy+WaEtou9N6/vGVgDwnmvMbV9dBW38NHqyRbrKbMQbStXOM
vNbsQI4I7wbGSJf1ulLqOEVtwp4DJoAJFRk+mKeQRUvUJJr0AXo90PDMkG4/7kgaenGf8rCmD01E
juo/ia1k4uH+2FN0d1tx/s2jCmFMt437IapzBOqEBczGc6H+Zv7jX2niy6hcFWjv7ffa6uIOPWGm
FEsy3XkZD5J76X2iStMQQrH5PGBv2GrKDgEe9rjrKna5g7azCcFdI1O/rIMMeh2IZQrON9YR27h/
QimTb6nMSM3yCBH9P95KT2d4FOPPNBDcpK7zplbb2hL7Ka1bec2DSeK15LAxwmW8QcedE7y5z7G6
F7AjOy6KOrfYBRUrmx8piqKt7SJzLgd1pWgjo39yBo39zEHKY9LtxEoE40wuXucKQgYvNydI26k1
vg98JulTwc/+Mm61AdeO82lu8CFonq8Xu/aEbqTxjiqxMTwsrnNh5QflEAUh6HI2iJbQKYMyT6kQ
1zw8T3vWNY3ES1EEQozH5yQbv2Pez/I/Jc0t+LpPuDlkMAEOu1YoYe6iOok8gJPrSCjT3S+p3IuS
1uzEugUHHA0qheLiZ0a72sBZBJSHridlBaz0Wwm+tozvsbBp9tIQuCWZXu3PWp9T7ppPtktseU29
luEDMpMuvhPdhb9OlcUCN7nZWcqx+I/8c4MJLjXAHT4Vn8mTDjG5z66REm5FjxdWCzGfZn+s3a5I
Ik7Sxl4/2IEsxK7vQo4FlT+4Tu4Anl7OGy4tlsSNcuLJ7Y1UQKpovf1XmDeUglHx4RnAZV5zNsJg
SdBZFzMZrpVAN8/uWULTx6BGO7WOZylmr8xHDbk4ng3hJmOwlXzvXZjNjyWvpTQTh/CCghu9KPmA
HcBILKJok0i/e2fVFzdq9Up2n5NL1g3c8Cmb1yKog0o6UMCTbNw9eL00f4Yr99pprdXniYyfT63v
LS12itUnyhiqpJoqhaurG9I4unwTWVCBahrNMe74sCZwq05Vv/hOj4Zu9zVPp2TTdmaZ6fCS9WsS
/RDOJT3rvq9RIRQwwPm5r3vSNJzhuHxKvVPUJmvQyzOTjm8BiqzpdTTjlOzHGyhSxLXGjsLmK1KA
c+GEx4CKuvhMFQ/fE6UxtNm8DgR5yUOfa66kiSEjyDPVno6Jq/Mu3GHLnaq8K41qz9IDGZONgmsy
dwBRLQRgNG0S64GoWaeJbIpM6mJoc//y6+sVuWa26hBSiYwv4yknxCKPZCDVAQ493XuLr6cGc9L3
Wjflx716oUxsyejBLmIiuqlR/jtKyxKK4jz6hdRpyx9fY768xHtlZ5kN057ka1Au4ysUr2f9pLFY
0gi1LNitERYE3GydQ2fphZ6TizvWO7Ks3ACoMpH7N0+wOQ+zuQkhNGdSecbcvfTDCVa4lwrzNJ9I
dL2IwI9sfNXp5Gq4z29dBATs0Z5gpCZ+WiIAzSy5P4WxkAgpU3o92T/K3LItJ75n5XUnoRMIQqgr
ReP+7JMciUSpqRhZ8jms/21Jrh6kBkmTib1LQrf9/cnffQk3rN75f9bYrYs/yjtl5wImrkpMARcK
VeXrGsWxp7Sqb+OWh0JAIbBNHJkQ+t5mOcV8qLA8swP1Nzo7OzQxJ5vfvATJjeDylIF/QA5SuYmY
OIua8HrGrIaGF+xlljvjRhofBlq7HIU7YYaYOCGqT7BzqJW+xEvCsMiT6fUwKtNXakEfF2ECBwX3
adLYoiBFkr77CvMV+3rmQV33giwB3lJsHtHmq4qwEiMCWj2/vaGLcN7v2qUgT2W5GoXurLr+rujF
k+E0VgGzbibuVQs+fpNaG4qLhpAzfq9DdiGin+SMILeb0Fle2MHXn+67leFvqm7GxmUdvtFsqrrK
HdLgVwa4jgbkWpkfOeI86sbbCvBUvi3zhuY+R9ysarm2YLl4xFLf1rKlgl3maKT+0IpMOg1GtkJi
BcF+5GYJ/aqblDAh3NLilfFX675t2GWk+iFbLpORilHFuoyqjup4Rw2aE5kpgni3fc1H3cmZoEsJ
7Ck1sxxyJ0XLL+TDfRhlqFmDEXLGMk/Yc4KU4bUICDEdeZzlp76pk0n1Ey2ILCgnxitsVERg4gVq
boaKQbye0Ar9cCUWZbZWeYX1tGDlZOQ/jvt3tVqGiLsnCfVtZQxnHK427FdpUQVKph0ENqXF5yGD
j09vqa8CIPrQGw74Nr0pzJxtlgWP64mXjTJpl2WuP/gwRSKz3ReYLSTm8N7JDeUbWnb7OJByiKaW
pE6XQN02I7FroN3+SQO/63ihmHIfRXKxXPWq3wPxciHyh8zkjcTYfcHt8FE8/oW4UQ64h1HaOFe3
9P5Lf2U6AQpr2sLftkTZNJl7SDHX5g7ZI6XVGg/DTLPqBA3TmsmkyS00srhKQrkod7olrMqaUieG
nI563IAklAwhAkGxiNkBUZCV8767jbbBW0ml+o87/iMojPLw7CotltFEPLb6H17EDPUZ49w5zI5Y
YfbJ3PXllms15FWXzTqgsOTCoLy/8zqd2jxp14Uepb2yV+S2vNSE4x10YFd8Jt5ziENH2GT41n4P
F7Hr96KnXhMhmXA7gAjG4/11QFNEwJfExmnz4XFlhY9JIiT1SUHVVM8cagpDcHP6Fn5P2/b1ao+5
Xw1m+xVS3G/5W5nb1RSnjRqgo51jEkoyqqG8woDfeJC4Ysp29X9L3N5AWnC5Ui/NponX+jaTFBAu
mQsP0qxGOiycZUEHng4SvQ32hhXKirfuu9abH3sjLMtNcHG3ncl9mUWCmfLNb1fONUPGqIeUb+uX
7ZIT2n5mBbKc2NILJkUWl5b5UoxM4xyJqjARt6piFq509b2jqbGDd3PYNHFmxuSxH9HGxxv2lHAI
iP5EyTzJQONErcTyx/ciij9vgrgzwzwjP/aMM4KRXjvsU52V2n1WXXCwpGiFw2zEA0v6m3L3u8dI
LjjFj0OtCEFuP8ZZiEA4QJ/YvQwlITNUVj2VngNTKb4/NzRSUhOyQrSAYssp/aF5ukxJoxLmkuVC
TLf4v5+D9Equof6A9uDPBqsri5yBweqqIrT1O9uwCVXD+tnGqrle5VC/osIRWex5zHZIBUBJMoEn
N7WYf1D0ysuW+HGUxe+BWo8gfSyjXadOc+AwYg5U2Iht3GRYMFCmZ/eSXf+9cNl1LYRMW442fQ0O
puI1GmUfT9jw/fqeCFsNY2Ew4BLt5ZlMInUhOiSNHjIsge+MQsbbuLumGOa/qq047IR0Iha/vnQJ
g83FISOe7Zq2a0PjWXk6koL62SWjP9TR/PdQOoB9jpvFdX1emzoKzW4pJ8OjJS/dcUhnrUtclf5r
9fpzETrxyJHI9ngjAIVxLVNOn45a2wWn/33WNxuvWGjCQwONfL727SnFLOrnMybglv7mfJ+5qn/P
2C9rM9Dexumf88RrRaVUR3fWncsg2qRryT/tztzAkb89VmNJqVn0JHsKHjFIkLvC9kaiFJLCGTCa
PM/Rpo8d2o50WaxdgsqPINXNh26xfjxWvkXzpOoUuDqKqvQsKum1LHq63gz+uUuxHhFbTkW91pEd
3WvO0vtLkC/qNppNjBARhzK4pZOAMHWnAxKLBGVxkHa03cLRITovuXW8q+z9UMwnqX0Q/bju3rRk
mk9YR3a6vnGhaBCwh8jMtzOs5+3KpVj+DEYEtq0x/XbLvh/Nax91sPowyGwKPPDPClvDMA1QTke7
NQlV9/7Ti7fOBLTOTD7mJwzXmtnPg75+zo6LLkg34x9rH7f7tCt5V39hYhmXurkqMwBwzO88x831
130ERlC/6i1JkwnuHFmehd3f48maGVCyoQk3dZt85qPh2JnjlSfumerYjtOfzeFoPvzVtRPbSJsQ
BRoMdcpoeNbbLXcbq+NuaQF/2Gv1gkMNW6Itd+XDWUbuXaJH7JZEHS8Zg8qqy+9WSg/IsdK/NHTc
c695lb++uzwy6E9zJR/W/EZg1ztOSzQLe9m9QOGOiSlYHRso+hW9nByK98KBNd8P5oYR8Okk4N9P
SgoDheY+7FBKjfVAZBrub18Qapc7oDKq2FIesl07ApO371/r1g+nk3Ny7saysHnuVbcYa2y0xMyM
r+WB9eZ5HlH6Iifa/5ttUHnuJ+tMs0kKPmT86no0Qh3bwWjKvIULINbkHUpxZUlkn4N0doJiPsV6
gJ4oQ08rEtbHQHjVjRVlXysgCuKgF0Oo30I9pZkf+Hr328J1TrtJvtrzSuOb367IeJcNnne/N/9K
hJy+Vv9QnM/1131mwaVgDvTO1GDECIKGYczxbN3ia/ZxVb9O8jDvjOuElxDahjxRc2PAWt+hRggI
8GfcYt2+lvLJBOtlirvff+nudzQmurC0inBIbx3/hCMuH8sZ9+vke17AI1DdlOR2YB+mLnTQVhFz
PNbEyKtdJKB4ddIU3cA0qNjLm/6rDKtEIhJS6N5Ob+vKejkSJE4e9fgMRqsDmYIa+phFaumM69wE
/dHra17xg85q6V69nkbN8WupDJh909Ka/oonVYHEgzxl/xjdotHvim8b3aCfPULGfzeuUZlZ0gok
8ZLGHBEaNaLxPMQWESefGs2UrbbnLh2IIvSvKVz96efdc62+IYCS696kkHISIvytc/Yo17duzNXW
E9Dx+k6hY7K8ubHs970FaPCmhRN2gG2wTXsQLNc2HF1Q3sRiJ4bJFRrek3avtfUPAI41EkpVbgiH
sj2IbH5IN1bnhnuRpsUhtjoEH4V5reL3Zk22ovRuW4Z4SFjXeo9P/2x+aw+LtMRMLdn8iPZATrQv
8GrMlBtjYNWKgs/jSqlVXjiRohyLtAkPIOhrywMcxPOVnj3ixMorlmneg5cI1xibIAxR0vBRBbEd
G1iYT2bdnn6gU7ltdikzwJvZxG9zLnBXj8+TiUqKDksTjJmwS0BzJwdMQMciA8PYeYKOddX3gD2Y
9is592NfIJtp0cs4X5PvKAoEXHjF3Ct3mQLi0RA4hvgvNPEfslEJlgV97TAif6xE1LOjxJxJfM71
J7D0nL+1Zl20tQeSB8SftvBCvy/KOIzkg40APg6rKbXAWz9hJcixvVRUAcJkPuRIr7c8CRv/m1Mb
25gUkKetgviPINluWWp2ZYQniA1uhdTkMRWwWvYCMTitRERHIthwrfiH0wQ1KcnbEaovWjo6kydu
slpUY8IQNyq24fXk4zD9cqVGa6cy/NpSwrT9S3903Sa5XDr5sf0HS5nq9aSQcAL3dYpAeiknS2LL
B2+lcTjPDhN7Xqwxw6BsxhoJxyo7hydevpRijpmo5t/uvRUFzBeK649QKlfy3cCcv4cSZ8qmnMEZ
C70vSiEdl2xtyqq5N6/ljUyEHf4QKCNBfTj1FJnNt+p4ilOH70k3nJgF4TiwO6BDCHOhhsALSZBL
qhlS/axU6qZuzOYxUSm2q7xJd/7VhlK2O4ja8Da2eO32LZbTmb01yjg5heUeJ11KP8XPXQgsbl4p
oBfDQpTqebAus4V1l+x1LIZ0+d9sSPGcvwwCGNU2Dex7blxVrkeoco79TwH632TkVkLEMTkuiLQz
yP57URCZ8I+2DMXbfDqYfP1eklblucDEKasftukE1JsPjrWmPlJ7O9JWzhkWe98hA0R+MNWg1YBI
w+TPRwYtf6TwEvXU95g4vJOGMQDRbDzfG6IyQQct6yKumybh4jRCmlN6gCx1L6NMhWJg3KDxvRLV
CcrQjtU7bKyzFHyzkw7cwR99qbuxoYwyicqtfFjYTdljFXIZvs/HkUzqWSSG//eQHlfGsZuNCD67
9QHZ2k+khJrd6L+RfPp0JVDyL416OI7w22tl3cA5V2ExwD0pDOvjjoh/8aCnyhbfX1uIhsqdswlf
O0tkmR6miDoWlGn6BWfaRmzS/ICQQIiWD9TjVXttEb11MO0DHEsQExpTF0uPgu/7xBF7TuwKhghN
75impvxNBjA5XwVSLjjPjX+0EHBNDSnfqwNv9dpAb/w6lRBx5RIPjSiozPazZww2PoI/0poLdKzP
LEaocNj410HZejS+21feMAKXbq0p3g4ZyIPIU0a7YNb6bADyHq7n6BQme7b4vMfLaLDNUQoN/AbA
z+6ymPXnLV1+PUHnTrHBx442ZSADJOMObADKIjcB/SjjNy2ODqG9E0h0bh7qnEUYUR2xDjNxu8sZ
AWskv0DYfQIh1pnDOOLn4k+vdETRrj1Y2wzGPOo4fCfsfgmo1fikihCF4/XWhdSJ59WhJovQjmDq
ZQUtW5uDaZ1gkbTj3QDeYJe68jI97AxrtwuJimyqKQY4LJ22jY/fMJT+f1k4a0SUW71R/HUO/r8o
QWdwSopw1aH5oFDO8kYLmpzQBtTgllcJsPMzJeR7hfsMldWqimGcpCVtQIxkDaC2Go70qLmDjZU+
e5BHdX+b5ZHloJzvFCfNb5uTHgZ17fI6ndzf3ZB7IMSlr/xvsK16rUK/oKnT4fLQ4g/QoQQ7JCYo
LExdE03GXIizn6WKfJtrbio/CdvOAaLyfuFzPSwey1fq9kmRcAZJSLLsS6NL3yI8GN6aUufQy9VB
0vryakNsBG4L8zNQoWDwiZ9nVjDseRA38a1r08zE0tGW+W6OV3qbX5i3EUwGCwlr2bF6XStfD3p8
PvKrSFgrzIR4c0SSFaIv5VHYIDx/idQpw60iNv6XQVryu5a5Qvwfkme79hgS9XrJnzmdoiV1tl3I
i3YCF/vF3zLGJbNYU5GCy3ZqKjD1g3+zrzbtUf7ia/zubAP64O01IHzr4GhHtIl82v7LGOS+EIDS
r6Hm4A8OoB2rMVOLX5PHYuwGCLbJfewPVcTciShCJFgu4QcLs+9GqDC9X2rQ0iFEE42O3ciBEe5v
Co0OM7HcDTTglZTlVMpb7qdRW3bmA3gOFzYS1BRmnwGU6sC5ssfHy7IXiLeA/7VSfFWLBhYULlQI
bz0UB5ltm96HQ1sszLo5+4EE40EzPI8pn7e56yWtclux880PVx5fMAWxF1H5jktHj9dYRYxQomid
Z8KKcxC7FrkKO+diur31aREZJ2vGjOcYRbyA+VlzePEDc0cUPozi5spUlwqEUKSWrpOQA2eN9iJc
fUf83NJvDsuPPBzicbrv5R7n8WxFIGTs5TMvzplyct398tK5pWp6TJK+HCsAfb+CeOzsn6UAsacc
DC6Vb57mk3V7EXKivC1FPOi3jOGCq60Z/oQnrAnI/3BNpXlyFJcXuqZUcTGOJWsR1ktHF6tpOf6Z
lixDxP+dZxRuiCzKAnXzig+ow3Mk9AKwwHGkiqGBwTAdqLeH2on1MfMAddHpZw47UnRqIdVhW43u
ZNBvMYqhpSJFeDj+LwKCf0/YDn2+PrUSLCjb+2eYmu3jYZmJiyLOKKNOwIB67p5+Vy9sRPAmxVGq
RR8xPl4PgZQSsY+ytxUnkmc20XzBUHycIUH7EfUnetYBTcfijynfLKmkHSCvs4W3ou1NCAFk6qRZ
6yuaMxZ41jHReui+OUI8pczmHIxoWWmmFIN3QpfI/f1naDUrrNKjfxTkbZV5spqLUA21si3nCKEg
OjS5k3lxNb1YDE+tK44me0+HpDm+jORJIcC5p2fp6l8PmSKSI/M1twtTAHGlO3qqGpJx3QnB6hBx
2XVPY0Bi6+OMX5okQhRv1uwxRqt0EYOCuWFjtlyALIQ9fMv+SnuE9fSFFD+HUqbzZvrHGj3kIfDA
M9uj87JEQXvXHzaPjTU2THOLrzhv1PrsvR8F4q3mJiLKdAPVGnQCn2mqye09/XklMvhw+tF+gQBw
8SRfhYbvezBkKoH2O9K0Fy1CwgJx4DRakzkLl2xY0lSAAo7LBxWnc3dF2JkqDmEo9uiowfTE0a64
QlAh4yeZjZiabAkDIvSWEu2c5b4q1NqdoThpeumQlwZcuqcGl1bJy1RZoBgrHWPhPJKKe5lE+dw0
1nx8tE5pcS/+vUbjM+4qAhvG7ZlsyFdfrkH7iYnsyPEVgsBeci2IDLiNo314lhM+T9fIB//k2k8o
BQKuRdtA2kSY4+rDeYzs1KQlIrvzN+y5h0V+0Z1nqK/aPffjUmYbGdb87UikepEdL548rp9KEp9T
bmCXnRXe+jBP3WL7YKi8XO9Mo3Ffht1bhz0dS/e3w2bRyVpteERr8PLHkCHjalyHeCTT3+9/9UAd
gTAH4C/n05weV+auv82XNiXiJwzKztof/oTZdi+NlBWS4XBDIhcuxU9SGa+5tSkhtUVSAlePkIQ5
MdKfxnwtnxGDyYWzgBbShqk/Rl2tOHTi40+l4ja+n4rMfVf8LsxWTqZHrRi/L7Jz8FtNgWcdEGtD
wJK4K3GkQHCO6infZlf667qtn97mJojeDYTCJO00ZaRqGibLNvUvJeIaHjLsgDC9dL++OZvQE4lp
p+ugux+owBdkTI1M+TkhYj39VHg33IdfM/t3hwpLQQ3mUnSXppPq9dONlN3ZT+gq3CxamIMSv+Jb
5EFqhHEMcoXPeO5QpNBwyXqm+GGT/9SKYal51FJO+RXxPfcuRMzdhnbo9ch9dTPjSSZgAJRv6VUb
FbHKEVkoO+BZzRmeI6IArJHvI8OiNHs7AE1Sl15LhuCMGKjBELBbdGhHXBb4xIHv96eJyaxLrXoS
I/uNCDKZfI9WArsElznMakO0klSIBDISaMpJK7CUXyD1MmdIbwoI9MNtENaWLcDKZIHuoKBBulm+
fQCqVB2XnFY5SbSjR1Q4dnagDUj9eAi/NAtoz2zILhdPNt5yL1ZoJCMZl+VAtJml4HXSUTnX+B/6
XmwE4OMgCnfO/46xfZ5F/sTnvWbEO5tqdaosjIOucbg2sp+VZmoEEde9BdTpVNLeqouW/eXqPzQh
PwqCcu482AdKWqskJmCx5UIbUPZtwd0+8Qx8ArDVs9mHjYBY+jW3aemqmI7zezcNgVEWcu2R2ixN
bh6hYXD1oHAY+kbDHJSuC1wRPuXiBhss5mdKSHwW1YlSj1o6QZbj7dZcYPfNIwulotYoTe3KZVN7
lzjMU2B5CuQR6G9AqBNNYMFfUbqBbMul4/4peQj2PDvdNpNVu4b2BL2CKbAlwWsksDpFKmxgaoU0
Xm48/xxR0EbxlanNY6PTDu34Io9FMUHqeOOk5yLlcD3nk4+KSHWCzNpGX9Db35Vgq6gFWBj/4DEH
JQqtncBCuAYOprnkYGaysodJS2uT8c6pYOhggLZvwrIW1mTkJxfTD/0b0NXO60Pjdv1CPxRM9qF7
Z2SLk7fXhWktjc0F/1o7OTpPw+jEe8+/eWyN2fIrMWuw/xB02wOthR2bjMbMqpf4kO1SeX5Wh8Gd
SLN6xftnB3d7EdPUticg/0pGnQ7kqv9dEkTkuJquZ6Bg+FUDI/5xNsL7ppTf/NJrJUtVUnfGE9rW
76XFc5ofEFKR94EutPw3xHTUfbb48EBBkG2twKRqzHXcA+pG/dpcB3bQgpYqp3/hqT0GuCB70m/U
YLsSwXvQzYEq089XZWziWht1+Q2f2a2l29/Te2lRaZSGAUxqhEnrHsJA89cNzn4YLruxD3I/wJBu
smyziIbEJknLFtKeLBhNw7iw8pIEQnit5CuS28RPH7fMZaNds+MGW0A1fjmkmJ2X+9HSUKfuc2oa
9OJ3g9IJmfk8I/wYYZM4ZaGbLJNAdu8TaNNAMlGoJ+QrN/hgHr1aobEvRFpJfaesiGg4QU02KuEC
P4WrP8hxKiH1Yn2Q+V2vS9XScLM5jNiwZk07RLBSBbPll76T8ZeM2ln0zeLhmnkH6ONoSXjmhIiq
U33byDSkEurHk2BfEYAasW5A+ic3ZpNb7ko0Q1zL6q7eZogStCIGsV09JrEwdvWWUlrHQN0FpsqN
iNPvqmEqIdvBGM7hllf5atigplnwvQJBNvojwa0nYhgYGXyCi7gE7bp5ZC00XaIGDkQGXc1fWkPT
NjtVg/VfftkGVDJ8nr6nThbOmNALffkzlg+aJsv6h+PERXtol/y1tpW/vNpSOpc9M5/qhGNy5YY4
B4hAGNaMAB7z+f74+mTULLvqQYieNUlQYewM+Vb/s36gA/KbQ0CxPC4FXFhoTuAcObKRyqkDC3WS
ue2DDpgbGBxRUKCqiFTn67vo8/rAZ/tUoSJFhkifkzyGz/wy5vBW5g8SdgrgZYkeQxa2vffilKil
Ry/iMCoUhg4nEhX9hoLH2JV/7tfu9nQQeypf1H9vStjYLexUH2HUHjvHxOJg7o+cQSQp90gzuXCq
0C7OUD9TM/8vpt519taTbJUXSiMw/bBG2OBW6/HsRRdLdROIDhlZx3TfSntt5K0a8XXTMEQoGskF
/+zj5OSr56d9IzWzuv0TJkuP5gY1XJ2dFI8nuV0iqss0nu8hGZvd3KJ8/12lDJcSWO9j6tSYH4o4
b/LbNB0r+3xj0GdVThQutLzUi780AAmKneAQ7+mVSqVl5CUWAHXsbhOu+WBmQC0x7IGpTtJ+FdAC
bBv+L/uykeH27yUpgURek20VwVkmXsOOPBLAI1P6fydKP6nSF3p7M0Mx4hLxJspYOI9wiHw+5pGE
ZlKplGUkgAQWw4CtDc8wUJh6HzXZ56GFAgdJEn46RwxhinPZf07//XK/f4Cl5KXRwamx2z1kt6kG
c6b7wfxkUC2EQ5q4BFFH1wHm3YKFeX2+MZFr6ptgMseNn7iQFtVsugguWGC1ugNC1a0kp2/NPop5
A5F7cdMjtOL/swR3RmuQCiUZzf9/JVfyPMsaXzCcy+fm/37FesO9B/sq9e5V9FrQHvtQ4E501O3O
qeym7w7IKcVwh4UWj7bRHV2dAkjOhErsr+B5HasCXb4lAat2g/w8CCKHqiGYs3dBjNsk2wakmMfF
z1wowke9e58xWPS01xUicEcv2dDe00ALbVNyT8mKxxqPAdTQKRf/W1Gnw8c5BxhtQwxsrLzNp63f
Pssw2O3yczVjwK3KO5IOqRz1VcMxDmNVy2JF5Dt1StSV6jfrGdVlAIuB/6C8eCfD19JnxmzGeTjx
rp85LRs+vE+LZe1et14WSwa5QsDO89OQ1IihzCTkFeJgmsj06lKxeg3cr9Ngl2CoMNMtuNha4tbC
x7SUVyQZD5707anF+L1GrEaPM2XFf+931vmu6AdhSspJlv9H3Hv/Af5WwpMzYu6lCdvqqW+bGAwm
RVxUeIY/NZSVVsrEnWQaAoSq8bbC0cJzLMhbf30uNV11Ewzl7Jj4EGqNjWZxdhDfXfi612RDYX+X
D4jhMq14BITvuSKpnZP6f0is48/KN4kby6q8NbgWrKUjXtkxU4K/zYB3VAdHv1s2/ap+X2ud+hp3
mlSDm+Q7wuInG7EDakyYsfgZaHZsGekY9i6LkUrOy/Cw2bQn6KW3QQkQb6qxtxPao7fZ/Pvb3+on
q6izjuGl02IhQ06QtEKqyYsy6jUnzki6YpM3gXiUvZojn+9maJdctSj2vtD3jCauQr19HsRrVR5B
rsYh2+xexyPxJLBnebzoHeFnG9HgaPzVejJcdKEsbUc87/WLQOZzPg48F1JnZS8T4tHFmohp47QY
2oS/Z7WWVo/SerEKXnkXCWXpXduedYvBLY4cBe4E1YaCbRsiinMrKQEFbEieSyEPaEwzK+iGaUir
3HtrQEAEzdJCLXhyey33E4gmnXuskG4vWdTxTqGvLEmmkp+nhKZUKzf7BjvMhMWRvw850xwTJFZA
nVkm0YWG8P8A/JkkrLn4xeX0WDj8IAUZIA0RbFmPfDAqNJoZK3JoWdAAlCdTOhzMOnIRTaQj36vY
FezamzN4STOQutOESSwAnLcozzb7yvnT85qQq8X34sbi4Ws2IUkhiddhY63DotKkFZbDTXDBj5lD
KNI8vfwBcfQchTgOlH+So7MtNIIHmmpHAGCIdbN69ndwz2l1bqKJfBdVux1NHamRjRfCk0eP3Onn
53f92mPUFKqWl4IWWF+RnF6B9ChOc/tHXE0gbyVc4nvmrYxypZER6Z9Icx24fQ/BReweII4sWPZf
Vv3PelPDmno3zZ9Fe/KXQ2+/o85ZOgjrDnMVbn06Cm166cCzNsM6bPQ4XE4vUQDOerZR5Nx0FdtR
MicYXrxq3zegkBJCYJy8iKTWf8XvFobGU+LTo7x3otm6rVZNBg9PPawdC84EBvZalInpI7pGbgXu
n8KVFQrKARjDu33wTaVLCuwwsgWQuUhSp2EHNdpRbzZEPOOhOZwlZZ24FP/jMC0j5LED7vCtewOD
fhVizgPqFpWP9dp/f1qt9JjZMROYZPBZ9H2k0D1hGwixsjfOfjb4eYA25pS2jQtoxmIc+ryBkubo
LZ3MVV83F5yabJyNegidNaYimfCCMErzYrEpDxX3mVmAD+Tg/HDaDE9llsOV/VMLeFIWzOwQyECK
kraxbFAsMlQplorIGGvSlm/zzPgzbFGdwJu0A3Xkvpw+sEILSJBNjVlJ+aezkCwFSBYFoptvbtSU
nFTJL6MdILOi0mgoVL5VFH1QnBo24flI3W1irMfOGbDm90zJ85BZ3URaLiineo8sVMV5NymGZ1Ia
7dr/5XdqC7BF0UWR60VEQM4sypFPGnv8ZnzyZ+bTNbZ0fnchHH64IReqt/kdglPniuRRFP+BUGFT
SKaMU34+vW3lNlw26VAm4IEwo58ExmdgNqN98P4VgueIGN3TvjwIngOgSQD5oHVFP0W5/MEfi8C8
Ara6LLCRLerigJH5Mroy0+LDJghTfFEu6AKLaB6LrLRzwNMav2tbgx6eTqjFQPubCOlzX4ke9gpa
QkGBrH5c/hZohDoXZ4EWuXlU5Axh80+K+9TP5LNYZ+wsXEvIk8M90JpfUf2WR4Oh/9i4gc4nKAhb
98/P5ZIGYJ57x6VUq8WCwdeqd9Y1GtZLhQn3IbBx3TvH/Idn2MB7wKrfZn67f3NVuJi3+guOBNoT
RwzSYVpat0ELyeuJOoBXWYjKUq364QTwtujYQ5lkKXkVIQhnNOI1gzgZhI2Q8LygDOjqIzAWvNCJ
GzZy4B/p8AVH0ghu2rltEqFpLIirVSI1RofeI76A07ITN8Foh2RSBt0H2S7sByInPFLGmaa6kXcE
zbEGd0s52rI03OESIK+9CinG/Q0H3s6iXCik3zeWFkbi/8jJ2AZqw00FyloDrcpco8EhvIQPDzxp
jc7cogPo7OP94PZN8lu3UJYpxcnZqqIvOTKd4/FgJGRaqnyAtuwFo4W1W2edX7SVSuWAPx/SAS03
uPekIYxKnyOU+O6JmX1D236tL8D3UOmKnb8NDWBvKAsuD9NX7Q++rX7FADJZuARyx2lrt/1X1ZWV
hXSe43P2eXRhMn7gzkhep8TF8f62ai7RIPrXLg0Wf1nYP/IFike3l1OsulQiE8yP4x5lL2B4LwNH
voFgugmXzasVooSf/yZaIEju7jH/STTo7swjlSO5yJ7KkgL7Ry3cr5ZWvtRCA4jxN2RRt13JmrAm
ktpbUACBiY+Hpe6vHzJ4XWqNeFawpip8LLutCAaBvDbtpv2RqGrGOE+31JgNJnFKQznF6Lk59gqX
JF4gDFFyqWbcFB9gJEqf0UmXZvz9VdeyZn1WYak9cLIZLB2lXgZ6N7C8PzWcBVR5zXv5qetvJhm0
LAi09X6pZmVp4+3GzTjF9pgDzhW2BAhdJu9ixtXPpbNWPQT7yIbQ7wx0PP4RSh1CfB5dCJ704t+v
yINPvXMA2U9gupw3NrQEsoWq9hJLdZXBKDMogTWjxeK0dZAA8xI4s9uqKhrG8GIcUa/UfjX3ffA5
XScOzQ8Ssegt9PtY6uQKQbQ4c9YdzO9YYAHZJSI+AUSgEhY33zqwmPENhOKMa/BLTI2ML4gJotxC
HKw+XUgMSQd0heDNxVQ4jJQJmPMGBgwLEvgSqi+5ZFCTNsitt3a3EJ9Vz2bLn5CROpC+A9Kazw9z
B4lRFgMZThzlQW+Y0odG5ciKWMoSHQHcgNXkd7dDBlfQ7ea7ZNzmAit5nrG+eMfQpWy9SyUEvtFR
+fpfzYZKNn5P6KtyCskmueKQxuUUaYqcdArFNeOSkK+ZVj7rKkwzfVk7Sk03hTttKDjjzLcYRiCa
XcSKm8eqOMXXKlDbbcM3o3nlnYxFlZSmP/SVBnQ/zjpZiSeSsVUzaMrkjvDbIWmL8rEWNNCoL3rn
KBMu67kW+vZIv6bfamxD/kOzk1PWFVBRitQvb9P5w27PpZZ9Szjndkj4L/WmkmvMOkuGmOa6NbWq
zBdgGdZ+k4+20Jtgbkit+X6/sz7I9H0loHGJT4wzT9TgXjSOwphrhrGsJNNQ10RH/3GiaKpMMKqk
5oXFlAGhuWib4cm2CDRBhUuC0z5KOc5pKviyAZ6YAjehkXzhaCrPGjkSyNAT2C+RBHMGx3Jt5fYQ
jn2n8UnW3JWQPfj2PxfoD4kAWmDso9Z02N81Xk1QzHS3Ajw290ZOwGaO1n9LuDqXxZsNvTefHk5N
llHUtS49zAYdswtapD0WyqpDJD33PaKuwfYbNXk8i5Di0POvfDMChg/SbXPrizLS/6B00cCxQJ3g
KH1/EIOsKYcbr3/FnrYudyxIEFZyttADrmuzwS3UlRBDwgNz7GlGy6xItWMELsRm2w+HGTfdUsxo
YsE/b0kH+UZkwgRNuFOejoWovA0ZsKJ/6Y29ivoCl3oQo5lXV9bG9BC7v+hjhk0tqYwJJ4kKOK0I
SV/qokbLAwmkZnCleWS05u8KLpJ62I/bs5xD536gO48uIVs+Q4WTc91SVhlFnzfV7DL+kgL/QY4s
3RXf/VwnF09nDj/9UNTPkKalOwhuNv429HmKue5KCFNxr23I/0DxIBOo/uX49Uq29cZQg64Y41lz
npqOB8gX0iL9KxDJCU6vPemYw2i1bv2ZE0TTqYnNx5qFhcTVLBIctUdAFJiWfzFxs/mKW5YysvFo
QCNytkAqIBpiPxZQgwjgx/6RgGMcRU6R5TAAAXLU5IH+BGxSEyLJCSoc+mwiQoSOksdW73Ko5m5C
pSORT7SA41nDL6xrECSUqA/2I+ACUzDoxKgGym85Qau791bZi0moPXdX7jtFEo1GzPtUrBwSr2nh
jymV1UOuWZbvTYlJyV4L4JJBTAKj+l3+G3KaqcNaoPQ6XLLtr3XTiUZEit6T/k3rM7FhuDKPlLOF
ZGSutOOj+A1Sqemfx0eXVPqp5bv9UuA3pf8tUwBk/kBQsqhhFNCKBFK6THOQajzCY6x4IkN9ikDY
5+yoqVfytRk7ulppZAvxql0/1LYeGvBfeL2X5BWUw/fsDbs2Tf4FB4FQejL9DfoOh5miWSS3JV5d
eHLTc/mWFSQcUYQTX/2A5kwK54UFTiYwFVXBGauqkulrirm9nX2mDhcxlLIbd5kXbD7wtCmtnC8o
DMKcl8SUxCz/cKWYR82Pj0G48iBwrhqM/BaWPVWhCe6YhcLnY10+8YsnHG6YzSrlwibdcD4r2pyS
Fx8VWZ0Ic9g/qfgAXeMJqTFBgT0FvlUs6pBRM7BW42h5rTGmAo6bIVWwSXUKGCBVpTjbPBmc8CqA
hENMW0GkTeL94dEUJ20Mgmd0g44WNtTUSF6N7G8djcgyHOCuEb4nr/RVE2kwKSocv96lBCK0ZOyS
wiHngWBMEf2UOOTo3nF38g4N1jU+wsFGKKmS0SyDK+ZhTY47luK1nuLpC6ZoPx7V8qdE3WP6bZwe
SejPi6YTspDVRY/hvucFtSQnJ5eER+3HWUXTIJCqtVMTV2tc+/rmbbOWdeDvXCROxy0Lme1LqK8f
MZGMomcssVAAjfD48g54GaXYDOHzCpWnws9SzMD1Ny4SWrLmof66NuUnRi68v0UeMkTrkzTRoK+w
+Wx6w+4qXdyvzzQirme2momDaqdV7HYh/5MSAbGD8y2W5NyLqmucRq09mBM8m3BEeGYoQH9oM5Ty
GC1fFxWvooLUkSqineexZjrX63XlDCT0SxTni2kCvt3cbiqU9hmE4RynHaFWzsgoJqiJtROdjG5V
kZ9VFCXrqjatdd9TIfI491xl48qXCkjIDcQwnHYZo2tb+NFft/JfAkcGb1hlykED7gf8ftrxBbFV
+bP7Vty7TUK4llNkUgW2diCvAs4OCtspsWOyI+iNyz1Ricxo06kxXXFRON0TWVCIwPxIOoNh3Kxu
l6UGDBENcFXL+PqZrK4pcdIUmLh4d5Npp9O5Dtw8+jL+6en9puK+mk//gq0oVDuFoUXbOksyJbTC
tExRF/nrY0Uq6eNhI6Ca59BUD4CJ5a4knxQ3BlayB+54CymBAcnQ9KKoIuT/aWMiGEbFGT/8mX5o
+9ykKfzlnW/UfhmbApahgJCALafswt+hxF4VgU0vUpyAO576felhD0YPUcBvyDfjOB6dPHA8E15D
t9m1nrVlkbSKzpUxHOGjhjEZFnyiIn+phzooxGcTxm8QMVyISTmg42fj1h+g/ArIP01Wuo9U7cIf
mjPsBacHx0JbjovrjMZPCo0cms/FPlfImcE5gEQksEKSyEycDsc7hb8RBowG/a1kjM4sOEmtBTt9
0qXNnHHWr39o3lp0WRTI7AMVVVjc1nL+3woHcdJmYBaP1qfGyAjAfOJU76ULx8Xbrt8BqNhjW9Du
nR3xlDKxXMOIoe/IMcfOP1BRnvPLHeSZlDKktCotwZepNmNamcJ8AgJYHACI/t0KVDakewGq14hu
MASfeuWm2vmFQ+RmgMIlT8oKxLsMuClicOcZdwkQSAyjFIpY5NX8lYHEcY7NCHwgJgHQnTfIbxEC
X5qSGiXDuOsVKT/BVZjstBI8SrC1Sc7X3VXDSZs4pFKsSEHq5M+fb3xWLo4OmFkURZsyX5K8lNY/
xIAU94rMXnVfOt135HZs9Ib8MCdXs5nPIgyzHtnI9FMhReQk5QnfKJjTriLy9oMNtHXjOeXAmqM+
74tIbgZDI1ajy1fz0Jewqxx7tqKsjjUxEwdl1xEpIFHagBlJufMOFe/G1aP0z7R/iUeQUtABK92g
a2Ht19OckhHrNkFtZMsRFEQ+9oJczFHJ0Lrc6Cpw+nKCMh+f+Zq6ABgRGBzeY0vOhWdrRr8rGwN5
N4bgjVoLDpgdMXUeyUuDchE8KKP61A+CZRZb5tzWu6NDULUwZ+rDePO0n7AU01cPcPFY0dn9YHAo
a6hu7hXytFhTgG3/awHq6z8Ryt6pYhEcP8ADZsF50K8+FazUhOOutoDKGtygkKE/+OjEcCJUkhxg
Eo8jCJV7GafN0YQ114RWtydeQI1zdO1c5wDW3UK3eyDvDi7Lr2X+cnmun0jN/MlWJcqcHmvL/won
EZKtc6KrCLV1kgZSBXvfnBN3yw33F+C2qWO00s//8yfqAEBIl6ICM/FSFmMFC8oR2cr2GiC0UiSw
cnZi5aKVc/vGT9zlRAB+6OpDtWG2OPSMMzBYJV6uh1eMxkq8vzggvex9JLVkbKd9hIeuJXI+oQxJ
V0Un13WoIZkThUGhyaTXRWz1N+4Ux4RxHJ3zX2e0In+hP/ViW8ICWQHlXDUI4o6bgECrdxctwO04
rgENOZDma/tqXaIKne8WaltNjJFyxgQehW7a+SzZcm/ChvHLCXZzbFhtymkJwJe3cuYE1pACYHg9
1CB0OrMwTWmImLJ9Ih0FujBEBI+h1T3OIjydvmPiDjDUDthtt/ZY1iwBORLDABvVHsGtsNfrU9JH
SJl79F7aYSr2LZsmgt8xBdtTGMrEXp6k6xBAym+iPP+EVV9LdgwzbC0EGhhfRp6m5Kyy4/+BtQRl
pzKfM2U0Hk+cX+bOOa5bq1MUTTp4ydReyoBL8v8VsT/TXo9Qer6r+lyjZU8TB9FRDNDu/znTjmhB
kTKNKBEif1yzhBs9wCQcR/SbQZ6T5C3TX7WL5Oo7ReX4VCsmddXpqmFmve+GBesR3bhD5A5ViL4Q
XJtTh5UmRPchCqIL2xZjAn+i8iccN3+V8CaRrmrcsKmKN/yaPDtCb+vf3MMX6hK+gZapLFh7AyQn
uDooOdAw9kRQPn7haVH/BI5cGmxCk+w4J3AMZnsDLuXfgsFGZCeH/xZmXX6YeZJwuiYf7EU1U7Vk
yDOQosb23cqsFXmcu9cHktr7Q4qUbI1kNq8EnfK7wP9G2hmE2e2dXkvT0neJhzNmrN9bIXWr//UM
YpY0XGXD6mSpLbyLS9VLSpb6CtsnTu+KeNfGVRq3ItkKWtL85JZ26sND2NTvl17NODN2EuEYvjx5
e4ArWOeJfYyuzzDUYfYjJxLKWSKQqaof1nV+EryZUcQ29z5xHM6P5JHLg4ewhTFmlYIN8X8M6lvP
OEHxj4YVuZ98eTPJmX/IbQBTcQmCyk7o/Wuq9oonDQotOfDw89n6gUUJbSsPvk3cxQiuoSxyHJ/i
e4al5cebjc8kRVA4ge7oWJlAferjISbSdj/Xzs84aDWVMzkyYgjaAS7ZDXXrUT+xZ57N+q2UUOOX
SEW93VLZjx80bJcrMHdExvfWyjIo51XenGhDcY+fDwXVv5/IN7LtB+phV3Je0el1viNQXu83LFb4
PQRpKRB/+CW6sHVeq9/9qdcwQBg3YLy+PWKFgv2gZKKlnpRlPymGByNqA3S2mBth2DW5wwF++ZJD
ygYIe01lChjpqmpqI+GMzbXtUzQBKbu6M3Q1AKBnVqBjKvfR1tR7EeMdUdqWh7vQtgbieXSONJUw
fUOnXpU3ZKRk7cXZKmD8oETiovND85Y3v/I2iLjE/nR2/amFvv5PVaSLuZm8nCml3Y1Kye9VU/AV
aNJrqBZUw4eMtQpPuNmSBkr6uLB9GtHveDcIxgpxEgCU+0YvCK7byek+RjhWUfbs0cU8bw8dEixs
syR2MSOZgbK0W/ddrTgZGmBGZw0HqpaJHKrD1bdMy+dsmua44TdbfXt/xfZUPDv7hDXyCLMKkToZ
AVTz0gf0wSZXJE6r3VXk/RqhigyatQgb5/FoSqLjayuWgiUxX+tqiEVsHR+wf0aEKcVxo8G+JSLG
i6LttPg2hjNqMHNj6JLCZyhkUN57n3c7Rx6iCxB86BL1zW7hrwP/9laoIzQnjEq3gx5oQ6KsSKmd
UCFTvfkXvvCPZ4ZPtIsIiEwboSaXs+XKdin8V++KZYj8jkqEmWkT/HjCrJoR8UWF1uLbzhIkqbkb
XkjN7tm/K1PD3nYOBVpIgeLH1ZLN83T2Ozoq7MwSfJDGp5xgd8gc9HzIWxFS1Wd5NhtXZ1aqEdde
xw7odtC9LLuj9cOS1wRG1DPZJA7ajcd0wwg4fKixIo0iBMoWHUu0OOBT4ZP91jbhWKKo7iPAUn/y
XcxVOQohp7ah7a5rqCXS/dlQrB0MsJVJPMRVTdm3yxQegPYVewQgpOsPVDzek1/HAwe/8ZbfC1E1
6T3o+qcB2jecHzRaADr3pQYFIsGXWjuc9RWsFIvKEDhxgAPMZC2TBrduCQi2XbzsO8daJPngwopt
wXW2SJQAgLJ9N+e0nnI3CWGaWSS9wt9p4XD/YCulLgCFn7coeiqUsTO5yonzZayA4os4r4zZlR8y
ubYDu4tXAQjMedQvdwfCf/8pyFLSFubWm24392tYS0lHFRmZWX4oO8LDIQf8ZsLmXVja5B/yvpKR
KwWf0LFXLR2nwyEpfdIKCwyIWJQ/Bp8jGIqF+OibugkDT3Zk+APfFKxdsqXzzl/A4GO6awrzgiuV
eYbfdvpdvhPEsWK09jxSxTqPq/2i4I8wCPla6tHBSXfLgMyjSN+pyMnq39UZWzZWmnSF4pCgA+jY
/dv5uYHwZO8rlkeUsGU4wHj5ACPLUCyx0GgNb2ckGjaiQgrNG4KJ3NFLfvnq30woszGai7NMK9dt
UWN1aG0Fg6MfuNLvQ3CU/pPN9TnU5nmx4TK6C/lsDYHK2H5K9UsQhwSGuLp7GOjLWmGkbgGtaVCU
bckoChdMEBi5ENIo+1LT9In+FhRGe90QTzV2310YbtM2LQB47BsMcTA4moMQb3rijxKZ6ntpTDew
wbvDVBnaMYM1Vu86W9azwiS6u0wzUVFX8X3awibpJGfFPLnY44ZWQwI1MiqEV1TY/Z6DM7giptoN
uLsIKnC8aCP+WoInH76bvm+IRVJN+6BSId/6hn6MiRziZ03i8RIekfaZwrALBh+Ju5Hp4jvP9EFl
O5Xlsv/2zSJBwlejpH4ebtvz6s3b0UrTfjKUx4MBZwFTbSMGCmAyEynNRdN7EUPQZGOy27U0cExT
d73LbtU1xZxAZY7uKYhmgTcNmGqL7mKiYhxT06QtuYPu+Q/quJDdna/Ikaod4FPbXMwKzgAMhNdg
GsDsWMKu3f5fVu76wDm8nJNyzVxyxY/Nbu2zGf4GBQnHklL5ut6daWDk45agTrtOa9G7B+i5YS8j
IsVpkeZauyDcQSA/iWZ4CPdht0mP3ce1ouDhMZHafrsMlC+5oBvakCGoRjl6uFZBr6S8U/9wEzO7
TGqgXkJQ8kxQPqtF0hB5llw4+csB72MeIStocd0gcJnyiCP0jSy6HkbmTKwQ4Mly0yVneNjB6GVq
vY96DVnRtWSd/mMv2cBAKd/4h7PyliC2KUmoIiEXkiWg22O/7EsF+//AfLnHy/XE5+EMafDVkvBm
kzRBu6w3lPRFVYFofgUpbrJJpobGJMSs/9JuvzsU/hgR4O7FxqT5H0VrOjwrCtyYiWD0oILzmp1s
Ql1OYU1cv6qdTrPdJUSc+WKhAWVOFpeJvkWV/kQgq1BEx2uz1RoIdSaNE6YSpjc4Y3+vmXkmJQNj
bnzjvSnc5YC/jNV7pRx+1vFokodHTPT4K4hmXAJZ2QfmBfU8cixunLs9J983HUZCJ6fr33gTt0AB
Q2I2N1nH1lwkiTBIjDNtcClo8cVv9Wp0caTtTD2HVzj83QFr+iVVnTsKHJiDGAsr+jEUoORG5hdk
GUaokwfNzzdKoN4=
`protect end_protected
