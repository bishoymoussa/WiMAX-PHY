-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
pNSDl163x5gzL7GwSv1T5BKF6/J0J9BnVgRn3rlucGF3UY8zi/JPMXV6JxeLVM+KxHFarjFD3RYT
O8rTW/pe4bR8Dvu9qev7uBdtqts/95DiUleJFu2mimsI4v3j7f84AONRtFXu1Lhz8FqhPg0n6/VD
T/Tcbrs13xXnbbAxlnqyffY6JV+jbXWdFBR2u9AYhaDnXSQdrxWHvStsJDEFiBg+Q02itXQcG8TM
rEmtXcEk3zjwg7druxThpeLfR4TbGvQmzsYNsZ0qyTRZU74xTzz3vqLtwxmmFbfPbOVBRn/BMif4
UdKqaCloaKauo9aynQYri9vfTM4RN9Qjus+ZSg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 8880)
`protect data_block
N1mhJMvbarsv8b/SqnL6fRn+1rRsWLYnOKSrHBXpjOo68KuYeR/WCw2/fU2RKdytSzssusswHrB8
iO+w1AVgiOgUywLlCIK4k32xZKe/LstH9+xLD3fvrUqC7bMGIs/PpPQdY1OiEKhEGtpdkbiYtZlz
3d5ss91VUzroQJmzbHnnfls5MZ9R0O/Qvs8klOXPl9hkHzMeQdpVaU9KD89lZFrS4ZaHNsccW4dX
To1uQXpKG1l6+J4/5JGPiigmVMhGi2t8kRc8QUg/5P8U31Y3WqJKiJ3Ws8tKgDQu8plJortupdCr
VJ2OZqNzMtJ8JoF15qod1qVlcMZ3smuWDkQDutY/vTDwCfk4asfgCEjXhozpzK0+E4afrEnNPDJZ
31eiEC+GwJooEiWiYHaz4S0GRfGmWGzIseeODsbxLeOFfaqM7fM3peoYU3IJyupp/LaL4qzKI91M
9v4oWwEwU5qMpaIPrfeiUC5sPyXHpdSuNFXjmYebsskHwwNRVK4OJIx2bFSyQiwXzgWmGY7faBI1
yl/xj4C5EROZjZE8D6OSIkKgSonmJR6zBiNAA1HxTtw6+k6gGe2MHoS2t79nAyn+TAqJ5vQcl57h
xCL4QJUeKSQOn2OYnkOxwf27WKlGLW3O3xxvvcCY3ohJa5HBxa1qTdNKVTd+zC6+BfUGqTNWeQ+L
EqauoSnmDDGV2icjiNC0jxuXCJAzMDOFPjw98TMYLUViszlFURGGFUoM2k9UhI3QCKLpGn7FgrVm
Hu6z59NUGWZCV9JIa9RFJ8h+M/r3SPFhZBAguM+QlRdfi0Pk6rfrX/YtCqriHiZ3G3OSUSwXrnAS
i18gOxkwcH4WbUt9zshzLe63gMqN+6gX0i9BPuc9f0AOF7ikybEjbtQYjQMcnExMCQq0Drt3HLd0
compPuy0iIbsfzY3zgv47QFdLvDVqvwnbciQCkHQJ9aV6oKSboYSP0wJx0KDILMYbghDnsz9qz0a
5F99Ks4/BePbwuHNlD5iUtC0duxC9JuglYtm/WVy2xN2ZOVPKSxw2f2AdWeV676SDFrQ91DSa5wf
CLnkIKfzLiqLWperh2X+OYjrZhuPq9Z2zG2LTBtA8FUtjs9FdIL+6+bColnj5WpuKVnk8jwSVlLS
jYJXo1oFrX34CPHSWTl/D6e+IJFsiIK+gAiL8S23RPS7MU/5gaDTR4H2rIad6A6y+j2uQxbuScXy
8rQe53sDO9PtIbRESQ3CvODU70rqqHBvzL8siAeV7hBSzyyZl4gT0D/QkQ2HKb1veOqKZia0y33y
8DMeZLOBopgN05tkDprONs5fAyJqwc89oxSBsOVQTSTHZD3/3Q1cQlYpYtQy5JbfJh+lGk9UPgGQ
jZh7yNRHvy4TFgJx/Gn8bsrPO5iHChrqp1c5sIccrpG5pFqOqm3Xxo7QScziZ7zGaeSdpJ5T/mh3
vxWwnxsDo2UdN2OYMCwVNKiOXF+ACV4v+VMWyElJ/rLtSB+B70sMiom94waLAvFgkHpam/3UFXCc
4k46bmwyTgk9iXrR9gxdEeXQ56GpOAgu9jYy8FlSwaSUCnDOfxII6O+xfXl/XrmciCIaCmnHhnWM
UW79rbAHAk9iovL2YLkFrh4zTm0aZSqqBhYqitgCJDCosV8dkvAfBRYYOJjL146ukF6JPuKsjVQ1
iiOyi8KSMZiKlek5uYw7M+Gq99DdBVlu1eSxjjDDdlPRDUxAA+/cGfjlwvJzNh2DcETCKJoFnVE3
Owm9//HjS/k25hI3vePsVWPoGlTIu17E4wxznvqaIkJqmindUz7AVlsKCHKr8fUmdexlacIV4pXb
d7KsLmmw3/9wciCmdFta7aZ1fMHA6MrgVS3xnJo+g6V3HYI/XYZC6NnZN6BF6vS4ay7I0J/VbFSI
D6iDZygcMzrcwJSCtoBXPcU0ZCgZM5060hmNQra8NMnaapcCyUZGI2cE947/tCy1FUIDPleZ0IFQ
QjoWoRSUM00lf9FpaNoj+q9ZnvWxyFuKalY69FApwQVynBb3anXSlwWMN3kENk+pgFNg4I/qnvy5
5z0u6OZ3AwtC9gARZp9ZP09vZyhStIJ6rNCulQDIV3bZnSF9uRD8COZTTxge3AnmX4Gn84mIfuG4
+bu2iKLBx5NsYijWI90iL0nMGUPFYx5teQ1+K7H5QDnUiZpbQG0xx8t6kQsZvwZhg2leYGts2FdO
foWmsqVvAMJVfpygziDNWbNuGzrierY8WRx3PZIxvmJU263wzl/NtaqXLlZ8gNN9XAJSXLjLSVen
QfoMGpJ37m/gyEpPrMHeUxeUUDQNl8vjR4j/GOcbipwqczYo3iQnyPGIJqjGauARz+i28QNqe3XG
2Tv/e9zeNMC3gQ/D15uDb+fh752HcN7rYy56KkQ1yC/9C0Nnl8609iVd2jHRr9qyPIlZ+Ps5s8t3
F3DwGSmqy8eaC1NL5Nd07TUqiBRQR9lELNhLbgtnpctUt7j2zToverdW+1Sz9SlHFm7ndxwTuPNz
fjcMvbk3ctUiKCYFq6RN73P/hZV4nwMuTBsmvPqV9w/173eQmDJ375zwtfNnxBLn2lH+SuSkquBI
a3vKC4Sa2Pm10v8Oz4deJPmNYoFGtiPBsE0SBrXDkb6uCQC0LN0zVctOXBEQEFIpaTxMUnCPjaSa
Mw6CBHrLZp2gi0KJUcbzehwctUafaqm9sF3yR604ys6i6F8ZYDJ4b0jxG4IO2tyPmYcGplj0/jqo
/2moTeyHKIkbm+5BTMiVkA3qIN9Sofdh+RsY87IMp+OZUsaaW2R9+0DqblCpgK4XSyGWH6WI/oHu
va/jEMbfz6abpTqI2Gr1liUWcJqE7PtzVgUcXQRNyXK1Ibma26FLrLDGiEJJR3Hil++MvStCgmNd
LxF1CgDpNPr3bnpValOjLX9/Wxp4sAKWMFtoJd/a3MldK5K0HJPrRfNqYll4Z0LSfHCSyT8AZLM8
HCmp1MJVISnKSvBTDrZZR+4icuSCsesqkL8XC4rqCjI6zDo4TgpdWE20sTwaEsETnvmoGeZIcdgE
zfTMen/nOQ6I4MYvIgll7smvcB2ZPhSKFpLeX+4rY/poDasBVJhDxZQmOJGL3oVEzC2IhbywOvxj
jUEh7EcJm6+Nl/CLzqPUf49VhEDrukklaYnPpJ8JzmCtEAgjs2oiAUzAm6IXRCi+Lu1QOMM5kcc3
rN6C743Z0E2xgim14dIzI4z3fbceXiJ6Tqu3aJHA7Krim2Mi0D2LJ4VmuQGOSgJWV+UN6ODxSC/S
kLzqfjEQHw9/bN1IVmp3qAy3kXVYdv8/gbJy+EDvPt6nTq7Y3e6KCMhWcUUcFVgJ0W1kZSUjHSE5
bk2A+pN227Hupnve0pwQtlWsDvjESyDGjWo8GKRTBRg6TRUM9tE/rgVRZNeUd92A2ZI0VG+S2zt1
YPcRLv5K6fb2ENyD/wuNq6W6TdFkr2BA62HKKV1n1P2VSAh/8rAUkiid4pnrABg3izRt+nPkrJgO
uT23ZxcGvpJ6KaGjtg/xQoSr3NdWM0lGi6Zam6iLAkhb37ZJm9rNrlsM9vic7rLLTrP9MhhCI3pu
ahM7g39GFOCEiJmzXYQBbKZVfCCtn2RfupImI47ySs4ptOA/pm7e/TzTsfqEuTfpfJ28rDzKcalN
JipSlcN3iFuXbHgS4PT8TZ3tTaRucqOZLaGnCg94S75HPZybRSkJ3nMiqXW7X2Gym6srxW1M9TDP
Nc76W7LqIqh5ReFIt/9+0J59kb8eMHRDpbHThfHBzXGLxEhTQ3cKUPt3tFWwKcImp2N3Xex03tLb
49QF7ahVchf6/bSMcQzmB+cSne1VhfryV4+dLY090+fbKZBlS5CdIyizDsveALNgY8R2h1GuAs95
FO0KZ1RjySKrXE0Pe4dJ3S9gcb3StVvzS/NWCjtSaeSqS6kGnIRYZegXhayfgwADkfePU5yH7Wk0
YmIWaTHeWxkRqPcikrueEKBA54cUe6+PBoplI1Rf3jstv3pdXUSbFflP8UgTPK+HovsX/hegAbIz
81xvIbYA6nOxhVdtOuay2cK8O6xu+H5dprYrMUX9SgJCizku7QG95o/f45ykHLImhu+f9bEx+7wW
D3jQIZlLYp4I28ZUMP2eXn12lb1LU0iLFwZ3Nok/kswRaj8qiLhjKPnwVFhY60LhA0UKjL6VTwws
ng2OSlvqrmOjRkXp96WHenzQ6AIiUvjJWbpcJxmfB3Ge7EDm2AdVhM0oqulDNKYc7im7/N1Fc9OB
3clcVv45Jab4w2Mj9jhK9qCwI1E7jF/eqfx1fFs79f/+4zPjn1Av14VNyFJ7+EUYRQV3KABC9BcJ
iS8jkN2OnJU0haPH+eEbsdLHLjkzTherjvm2VZ1SqwjaeB+vt07K8Ge5oQQrDaGoK48i4k8lIAou
YcXR+JZzIc81QTCwGz4y30PgGGZhadggbYoFMNzjgNMJW8KtUY0d82TiJoxhGGXvODN5PIFDAws9
2u1qORbi3p4SPqWVHmYKT1cIxGzdcKUo0KJ9WjU3eOAU8L/zhSzKMxr5BYBhhIYBPL5THy4t+6u6
Iml79aJNCVvbQ10iJzrydXJZzL4AfxRlUpb2G/2C+xtYwpLKSMscNLQPgyTuzoU7DebhePjhEox+
3/rDuWlR8gcq14dnHLRhMC/78xxKV8RwcCLEJMPwr23GLCMYyGJO3+6A9qRhXQoKfBcy+0VlKB4G
xgBp4MYxJsoZ/D5mmgY4G1EsAiWHjNJiKQa6u9rxp042phwRVsMq8oMEEMJsQMmH1T4SWZwAjg6N
sc/Po52JGsbSISjg3LL6JetPIRJmFFMyxeaUhfL0opaOPLa9kSiMqeSi15xTV1gJ3JSna9jLdoCM
rDnqhL7/CRgtOuCwz4eriSiVJhQ5m5xIZuRKZO7salwQeh0V7Vjuu+mYSHRNYdl866pNfL4SH3r8
8izvtcpMKe9l9rGklnq3BoUG6/ObN0HtjsEFSLSnw/Jqbs0XY0k9iDH2rgTF84MhVXpIqJBA6usB
6CU/a8NvShEG+P6ZTsWlxgYvFkoLSAMPouRztgdQYFKzh5rcaMEnZ5MMbGxWiKOpSKpnYJKRkp8Q
9vfDyis5Yd8/MGJ+HvgQuIPeokwuEA3ck3VVA0vWqXWkebTbJfsUK5jXnijmPOychBlGuug3ECJp
k/EQNXwwVWF/aCmHKUmAbMCsRLUE3RrFWA9wjlHM187FXZWfWDdthNOmCXdMo5UyJ7tiX1h1jLu6
LlqWCr8ghw79P2z8r6Jjk2GSzH09ANZ4nAPIYuwKQUIrMXrw29KfsOXjq8CPkG2VXd/BoYLu7IVQ
JpOK5lH/cT3W++SHXwoO+ihNYix6lxlAIGWrasEHu9GXatXUt/ozPhbRneWLKNXe/RegnNyGeXBG
rFjmvy3IyDfUZ3SWlZhg+COo/R3zWP4wmPjiQAokMYFA7F20g6S49xeype+XpEyaTMwxKEsCjlV2
7v2kknHjTxMGXgTlGaxzRypYA/VEtTc8eMoFvcU32yTpBJmfcCSSd0vlSGhXkTP2dEH//qpsGt6A
aMwEi+KrSinHXDH7Ev6XPluxB4H+VB27ppXSLLEtx5sO1O1JNZDJJdo5dBrjOfz+LMqltLFOjsqc
butahNqYbupYbChZ6IQT6eyvIRgfEYx2A9l5s5FZyOx0CFELoNuMuTLZNU6Xr8K/gr/mg49XmB+R
Vyv54Ol3HMsa6EYiSHAexQ9+A8YW0s+yR8m+DBQ8cT+vCIM8DebB8m4C1qrgxOoQ5+7tRhW5bd8f
u+hg0tJ5oNk9vGa8Tc4U5dK/4z3l6n4eQrLK9BuSgDrCfWxIH+eUScjOL0NWDDcYbJxFDjvf8WNd
E7z4x9QEghsB5EaHyexzpW4td8nmqrLy72Ir0gplAPxyurJVsSJ3SlWw+317tsk+7uoX8JsRMmEn
HTGaVw7k2V6lc0rL4Cm1uenlg66kYafWIm3jIgNY5iwqaFhOP1yRxeHcOvgY/i8siPxzmzRw/iU0
3SvLWjmHg7SIk6gCs6IHnqamM75n9ebg4Sg+Pb7NH0TYNGg56WvXIGJbQCc5Ad8jizlAN76eVlmp
DEr9XQ+4bUQUTkKib5FFdKOmVpdrxXwY0xOiYJM8w+vdkBHUVG7D9nQyHr2MCEDNe43qC6LK/htO
sqr0QlVeerYY6RuAaWYCiOjXfsXz0fofg97/je0hrVNmGA9z0FP7WP/fBPXwNdsEnPxgcK6Ie+oN
ccnkTsgE7F8VnyLTVP4c2emqWhfkOPWzw5rA6UvnsPv8NJMhx0d2Tiiv27xBgiUgjwoVyf1GaBxz
wJ4AkkyXOafe5L8apno2b01f7MTEpuVZtNBVMqg7871b+wEr7xEre9a2SfKijJrDJX2bem8IKhWc
ibDcxB0FOx8HAi/PzC97lUtIxYHru1kDrhjevWiDFgVJCY5LB/QUJLX2XQWTGs0hMyTZZIkPzbxr
qcOx8JdoemRhtyzgo/K3spkstfZG0cS5gb9HzVJQuPYwf3Ko6nmyigQkM08g6klEcjYOS+TDozUE
uSxy15nyjH/yxo8vpxQDdq8yY9bXF+NNr4d8zOYRF8hQ/fEj57Hbj2uvgERxYOaLmPlRsyeDfAos
/JWS8+x+11OQO/Rzr+F2at0YkavoAh3HDLdst4fLfDSJBTtkaKTL2tpuvN/2iDVq52/hcDdlB1yi
m2dyIkWXaGIxRf6shY9rUg+Bu7KqR6AQULU9gm3JUVEHPKi013PbVRS2CpAsF82W8Io69Vmve6ii
q5qikjcv40BLulNJ8zhxNbLPARGthBTz2/peo6ZdmBGtQzsVdvPoIAwTn7NaHKpZ0kGUMB8gzdyQ
XLo/OxmLbJkxCiSH79M4tVwLFv9WLJwkuKrvWzDQ8+b7ovb6KgFE3DOYbs9Fn9wwa15Omt0yp9Fs
Lpo8pHN9gfAkjiyNRdOKGRW7BYiWMonTlWHBR5A9uHGheQk0ljtVj/7mi6pOgyrOG3N42iWycXfn
RoKhpF8D7f8qelifBSc2dPaHp8TPuCgunC2nABwQn9Ae0OVkUXoMc+SzNTupBrp7ErAYJHlTbiw9
7gFWR4e2PdLLjc8unqQS4AEnH1AO6PnunDSY9eBH13ECYp+3o3nGzUeada+PWOMMlD+QhvsPHjM6
LdNAs4rK5fnDn6z3T/aahJ2+/oED+EQE7DFLOdIjqsdfnw7/vxVPC+dRmH3QexYOBO+HSJcSfWCT
mYBGDytLJaNdLC6vESkJ2bhXy0E8jRuwJ5OAy+2Cxz0uDL2LkprhQjuDmXmgQewW6Z2dlkNupHOq
ktf18OWeq3Hf6txtE8gbFUpcoGdyj1TvzVoFRHPtr6Kp6BWgio5N1a3Hw+poAFwm9lFXj3HEZPxL
4yGO13MQlTFF8phS8CkO7vpb7cv5qcevDMJOK5U9bxphL9DYC6mB6F4SUAMLowuYNsENuy2T9rgj
3y68vJ397yZbrxX2BNsZFW9zbTa4OAT/x+DOg7pnVUz/NBZaudmEuF92AF6d2qfqDFx0J9+HbYpa
bCZvA3MBJbuonH0w6IAnKPHA2wK5FuBXwiMUmJvJmWdkKh2dtNXlwkj8X/kwFbc+2eFh7845oP5o
mOe6ZNi5zunkI3Yh2rdh25e4DQGqk4m56SPm00eva4RwVG2UdKklaJiOcmvXuiQsbkPMb3IHc8or
NUTn3VOMUYrlcnFYP23Fpg/aWWlGdVDZJJWef9w7UfVGzUIk2bxCxjYaww7v+ZRH39dG7w/CPtsm
eZYvnoVBbNQDzdPBDTUyBUJaEMQWnxL8NgGsCKxoThBYU1aTw2M8pBHYBIqVGexu+b/aJPNn5CJ2
jE0GWjGyknLttfszRNKCz2RCc+OYVl+HalBru2SM5UALjJJ4rVANheIcWVX2l4sptXkD5WpeC+PR
fesiF2re39BZeQHE4SFs37Lt+AvFMw5h/MW689Z0pJsD0rkchO8uqwHAq4/eaDgNLbAQIhvw+5oO
xRH0M+zEn3V++D5u1+ej/3/2B2QitL3j1kjO9cChQjS7MAYp1mXCI3TLFAFVx/bNXKoBId7Bm6FQ
LnJcQ2+kFWNuYAb/yBavQwJ4P6RVktX6hbnhzO9/MuijR//9fAjWxlE7xr4nyESsBaOTlDF3OJls
0nemUDKjZx5yTll2hK9PeEGz2RcM3ojwmwYepKy/7LF5TK9LxqST8w+/E/H8ttadpm25Lgv+Ft28
7vSa3ubdsVApbYs1NQqxLR0vnVHGcsEjAISYwpmU4LS4aPEnBnK3ehqlqeW6EGKX/MU53/vQcc9y
Senh8GeNOB/+5KliG44xPsPvIQErqxar4f7UhZkEWqWwrujzv9aWC4Sb5DDaBEMymD0yTpFLUJg6
JKEJIRu1yc5kVPzLGs5FcCqInzo/CNRkafxHkEOVs6fs86Byui6PT5t6kG3hHoWPBi7B3xo5fVgl
nCuUNuHpr3Ub0gZVN/Un1IxHbWtPeCFV9lCYU+pKemNfp9jmaTCL6fGAkMizGZekdqcOrgBIf3N2
1/6iXd64BZ7SwMAQUtDm7Hbvq6adGw31uDI/3iw9uk4dm/XaeeBtEUa32zMGz5tNxBzv/whFUyv/
LymBiY8+OJETKbl0Y5Dm36eN3clGoRIRAdfZMtGWQ9SWitoCrHqRMKBahQN8x2/kys2sPZJkw+nz
WegMHaaYvZQhZZiHvr/GUXXQQI30JA/p00IXz/1yd1b9+ttKIsP4zPniIhXYPlTPvf2ZLd0P0fFA
s+krQLtMUYNvxEAh5CmawjY1r6ZxZHipL/xEXud8o5g5/NgLnNo222JlO7EacbXzQ+Aj7GGeofzE
2+A1+ydtqznMK7aI29RAGdGwFjFP+FHWmW/F6ihASW4kPTBIGTdJMFICHVZSi/hYfsALSj1++Y2C
SzsOijMvwPNsE/NNnN9yQl9dIDCuX20gIFSO4OTz54vjI+ZCvxfEMD0G8EQvi/rho/OLLjjTX0qF
hV4oV+gWE93qbVmaqSB4KTu0EvyR+ZyeQU0O2eB/DcLVNrZaXfCozO4pmgcsWbRnTvasxM6GAs9p
jumWH9LHd25hpQt1gbhpOKuhwx17qGqrTRa5y9SkjDkjU7QDggf4wexEHlPSWFneLUSwAs7qAPHF
eTEeGTmIxrvy0sEKfmamB66KFrYG6Zs/kpeQCiofYBRouVwrFvgUr8QnFCds5LY+V+sVS6BJJrK7
wTuT0vJdwrlhMBChDPuq9bWazr6yC03XZLlmxhsoSpqiIMRhiOXBAt8hDlZmA7OO/GwmALhl1w/b
rMVmpJPOnSxiaZM4ayARG9updtjw1gyQGZ1RNIqCYtewPVOJq4/nr18oomzO+SQEF+9IpiDpQ0od
Y+eaaw6BQACEX5OPvLo+AtaPRl99k4OjsqslFiDWnyTYkYOKgVbnUZWFZWlCR9xpdo7keUaFIcHO
MnTUV0bGjq15M9vcdsrHbX4zmHXQHYNMaX6rTmFZaLmfCBMJuzWu+nRZlRjad1mocTYf9Xps9WSi
Anb/F22gjQAj/lmYKL5xCHsv2lD2TwLr84uu+dku8T380fUKBhUHHCznJ85HhS3L++xFHCbdlksr
667r+l8wwXQhyg82HRZgPCcgMvCpMkymqGq5g41GxeD0idkZXyDqBbZ5WxBXlvgQlgUX/Lh0DS7o
38Og5fsXZXNvKdcsS8Ro9ao8KTEPYpGo+mEFSNEGYVxxwkntCauCtmEo+PvTehWd/VX9QW+cOaOb
JJAYmdD5IJ0kDomQbiaZ1+AL/kj4FaBoDLC41e7D2MQ4ccAUMU8VJBLym98n+iMOB2orKhsRQXpK
Ye9Kn6uMzRDqBnsQjnRsRUGwv1Vcc5ildbAPIrCI8zJLQFksSwGaDZZp6y6IzgQKYbs71RmYFbl/
0MbbVwdQTS/BimeFjLwnM7Dw1IYGT0NTVRdi+mF0I9GbTLpfuttc2/ew1n0Dw14+1OM3SwwzGGL5
ftV+zK2smllGMRNE5Dl36hJjWfAYieWN4Dq1kXhi7eHDzivT5uY9jMXe/0Q4FTJj1oTtDjORFLlJ
+eH9N5bw9zQDgJ8yHjz0cq9aeX+rs6K9fHM0VbiJ+o46JwG+D0uBDJVrqORTm0qVDsI4VPgqvRb/
uhvEVZojr6JGFS51rWDbcxKd6xoET0hxH5PABa9hwDtM2eneX1/g05m4na4IEvfQ+4XkI8ewZLJL
h5Atdaghs5T7SYIcdPfz8jkFrdZF6IxXkuAEuvIm8yN2Z7W92RF9umK1W37gkfEMwPKmWH9LcnwT
8+v4AAYOzScqMZ3J46FYRwm3QNs23pVEwhPHV7v4rQeOf/OmWMexElo1CuPPO1aLNKBx8KpBG10U
QBcQRG0wZF9R5lMHzJYP7//iComkWosBSiGNaefCc1wRX0q7Une8Ryu1mFRoOLySJygo2f85bjQZ
EZtQVrazup5JXxSccSXJ0Xi/OV4MBqkPTwIsx8UCX4S2sgF7pZ2c4HaBpDqro4rUnFw83tkHuexc
D8eryTYiZXv4zyfnwdp1rm2SKgz0e5ENG4AsKhUlK6MeOedhu/kZL/K4ROtuLQyX6Ism8Dd62oqV
T3QDg2u84wGSqI+bkWjWqyCpvpOgqIP+0jdbcRfqogiUhcVp1X2LUXAUM+ziYE0ifXSL+Dt7y2BG
jbQ5+JIZ2UR8txlDgZgT4ZGbgYRgZpgDxP1CU9yFk67jrhZDqGGFR1h4oUuZXzKby1esjaxUk6b1
wDGJDlwu7OBnHgIORaN3VeCoIscj4vkPTI+uv5Q//txuwLL3Qbs6vNet/vsjO/AMPQYjNM02kZVW
a0bYGWxuTC9JgU3zllpkcZLo2oxX5zJ+8k4D0d74wqJol874whuxSv5yYPjPQxode8K98e9xHNGF
sQinoI5MKoFdCgDNgo0ZOneuDGtB9GOsgnUegB5QakehrrfCVMB0LVWRiEKbSbFqV953QhtzEP3L
YASDu2ytfKJwNFOATo4cRu2w0CGX+yFvMet0oq11UerkcmrkcODlq5zQOpscmBzbs1amp0UJF7nU
9pWTpqxW0jXv29pGYJ0aUH2nb8pmjhf+PFFs1cTdyf7uXHSrEbXIE4G3ZV68UqMglR5dMNREomRy
Bjpk7Eo4+/yoyLd5rV+fcs9jrIh9c5zEL5Qe+C3zvbnajPeye5OZDDruQxO4+/mytr7XxWuE5X2f
mtboBQsWE/2oyRQyR3CVurzMj81kcxYEfQUxZ87pArNXei7I9Y/wkqMg3IMlezguKH6MLAKPxtgB
E6QbXH1yDVuVy0+V1kutPmdKizb3+LVieWLi7XHDDaq3M6zc5mEDn2rK+RVmn5Aa5iRTi4Bc3dha
0k0sEJ07RStqvtJHFFeDwSqLTb8Ea/dAPT1D1nmlftLiCK3Ey82IQxKiK8Yx3HHIIr0ryMahAU8H
/qaTATQx2nTqSne5gn5xgQvJVoszmqcAoobiLWmC5QctWBdr2ujn4A/VqXZ0WQZvyXz1Ve+8WGPt
B1UA/3isFnLW1rXHYe0fMcQwm8aKkMBRcl8GyOPL5MDWZl5fgJ7CUe6XOUXrf3RshnKY8opJ7CIi
4DtKYA/ePpndiJVPe7V+Bg6UyzPj8xQa2gKvF5BcAE/fkex8pfhZnDp2NORazOSankgSf58hxYA0
7RSfMjloh9OT6jxuH+P7JHYTMZywUHOjIDcgsCAUDCgGdjAaLG4i6TGTyZgo0ewUx0mULyQfrHki
iRuSEVV7q1Tr9BqFwU30Wnu/UzDRtlp/hFan5mSlGNeScIP7VP0Znaq9W32wRUSEwzc/W7jhIjx9
QMSoPzGxthuJHjH6xOM2QAOK6EzsiygOB18CIZ4M+78OTS/mez76q023cdxf
`protect end_protected
