��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$Rx�y�<��wA�*;�x���@�̦�W�X�fa�M-$u����n~�%���P�$��W��kYَ���P7�?UMfT��q�6�U��k�>����~�\N�(�����X�e���/6U|)�X2pF�]$h���d.���9E�	�IN�f"�\��e�z�y�b�����Oo2�?�qˁ'�͜k-�K�P|����y:����3�l�d���bl��ˢ_�d���kx�rq�mh�MذM�`aS�.�DW�mS�9���Y��+�>��!��!�T�uOB���,��\L�7m�O��W���6����'���j)n_�I����2:��$�K�2�Sʫ��l ��!���{�l����.�j4�	��很�̢=�����N��s���s5���_�R�>����ТP .W;������	�"�מԫ�����]�#7@O+?�⡾�Ԫ���e�O�\A�	�ͼ���ƹ�d�	@�nQ˰��E؁Bf���|D_�%au�-�'���w�*%��"AM$w�*4���J*!�y��	?L@7���f���ƈ�|m�`����0F�	Lĥ]3�L�QMV��j��%$!�ʢh����������ܴcZ�5��?�B�������ק@�So*�u�RN� B����;��L�1cI�`t�y�4x�%k��R�������~&�,0���f|у��������(��]�]���}�K��b \��W<!=�ͩ6Q?9�~���7<�-�t�E�g�����ˑc/��/�[u� ��ﲵYݸ_y_@����U��r~�5�X����x#)O�áb�W��ۼ���Y�Ұ��W@h�3�]�.�i��A�ְ�7�QQ��s�G�����
_��L3!7�`��\�[˵�Y9��%*�� �d�\㞮Go+�i�p�%�5��<�]�K����]��-�cn�q�����Ѱ��Vj���3N*J�<��#��~=��]�,�1�Y��g����fa'j�A�ȱd����?(Ǡ�F��k�{sb�j=���(�z$9fw
1e��[F��,�C�R�X&�����*���<�+��"I���4J�:Q�u�f�J�ì�L:#s���2��GF�%$K��_��gF��uN+3�z�:g�YLh�4�&"u��F�Ҡ,���i23Zo�����	�&@�s*��}vm��T;G�Q� {��t4k?T;9�O|�)Vq�5� �Ӎ��}-���d2PuW����+oj
��/wqLo�>58dw�B�%�qӋ�y٥d����	Ӵ�+��%X���>.��rl��[���{�0��l�H�%�Z3�JA��Ṅ�<i���h6L���˹I~ə!��;���O��ȥC�pI���~	�*�w�Ȧ��'t�_$����?��.-0�b:t��6 a��j�*89�I/�Ƶ122GF^c����#�/����NHw�k!�l�s�� ^T �ڨ�Q3� �%���Վ��v�Z�`>c�i�!������A-.wV�_Wa������]�8���(ݫ�(���o��@a�M@&49������TU���F���L��^�׊�B�I"Q��]�nݿT~ѯ#�9�d�&�tgb�^�&B'�Tj�FH��~��Ə/��1���]�f67�Q�VO3���x||�JID��u�ѵ�f�p0��/8���$�bFہwӸ���|�%u�(�4xn-��J(�����+��=�l1�tç����--�eπi[���F�{O�s�V)G�Ae�02����5!f,���8�eJ*-�ɷD���ɻ�+�X���<�7�K��wrf��"�Q-@2l��ARi���	PM�(��2�9m^_�y8�����l� �.�U�+p�T�����G$!�o��|3�w��l�W,��
�@6x�ג�b�G��bD�rVѦt%�l��g�m�KXU�%R�,�b� ��̌��P�IZ�˼�8��O";Yb[B�_�y����,}�"P�TO�LQ�de����ee'��Ӟ2am�MeJ6��_U� ��p�&�X?��s5ѭ6���؟�u�	n��·J�3��i���1�����"-��[6�/%F;{�Y)�6s.6��2�Q� ��GZ�m0��dH�M�9�ea�wsSMb��~��e���c�Ƌ2�y�5�d0(���&]N�p�hlI2o喇 z��Z�R&���ލ��g2�<3'��O�VͰ���帕J=%gy3 �nL0�A=5]]�Zb�E`BZѽ~ѩa�jC�T��M��`�s
���*��!��$���	}�2
-��Q ��-���v����X�K��t]�*�o�,�� �-���Ķ�#�H��p�mS׍j<-��	�|�7S-��n�G��_^m�3��;�3|�,����ꕡ�4P�`�^7}c"s-+M7vnD��iJEe�Q<��U�c=�-��9X�SH_��ìA��	��@�?�WI���ؔ�����	�<��Aњw�F�#ղ�`5����Ms�
��N��a%���}�-�D�I~Ճr�6E�������[�	�)�|V�r��Ƞ 9��ϙ9�� cޚ��G���6��Q<5�0L3蒗f	C���Jo�����O�*�Emh0�W;��G/'�#��Y���w��w����K=����@�������>���Y��We��h���kR��YA
�-��ݟ�;ͤ��{���`��׫�ڍ�"O]_��h��<�9ͭ՟�AܕMX��;���+��C�v�����?޾�*�t�tva�&Iҝ�'�=A��yNr�Q a�zj��\��{�2�i�
96�y��e2��_8\�`H��H�%�b��WT�:ݡ[���-����G�\�d�/�]7�!3�<�
��[%04U����.�ӟ5��X��V�O�@��x�Fҿ��2m�#���[�`Lƍ�suB��-�N���,.������������w���`1hBaU����H��z���F��g�x���������K����X���W������*Q�Oyu6)~4"(Ws�F>�6դBɰad
WΔ7pB��yt/iZi+$��?�H�������Ζ��t��CMu�^��l�2Tae-@�7{�ǳL�#�>��MF$�C�ߢ�7���Т��2zU�Ǥ����b���|�p�W'Jj��b�{���,vWx&��j����<W]�Z+ ٮ��sBX�k���VH�� �D�.u��UYL:Dk�����Ez߼��6��O��.M#:ڞ�MsBs���'�_cq����?q�U+g����$ͭy��u��Bw��P��&p��
���(���cwn(��_8����^�4��"���g�'�d)Iqp���f�Y�z= ����,~#��E�d��|��A��W�|�Ȁ��%�z��l��W�4Gu��9>S@�]���OP��
����0Ǒ���Fy�|�C�ɷ��f��0� �-=�<zrc(v�v��?tg�\c��q���w�%��� :ȇ#mU�$�M�[&�DS,H���3,���o:�΁)�u-���RUͅ����q�e���u�&"9�֏�U��Bۘp��ō%�Y���C��	]�9����H5���ɨy�C��TzFFq�z]��cD�K`����^���P�X/�������w�� Q%X5�eܔ0��n����O�t�}fP����/SK/s��&��o3X�y�1�.�=���$D�� �P�������q�Gh>���Y�"�}�9ˆ��I:S6P��mh��������s���BM�֟`�dC����3���'8,�M@��g�����(VV��yc��
}�^x��W?�G�Aiȳ�ʔ>�g ��2(�����c��� U4��(`�c�z����"��O��~(+������b=R�-�<�@�0�]<��$�V�tP��	@�!�8���܁;8�g�y��<\���32,k�����}4fb ����D��f��P�����p�21�r^d�\'�S�ü3+z٧�y��ܻ����R�9S������(�˷N��{�V��U`X?�9��rIS�o!�1Z7�q�3�V�q���Jo}���7ڀ[_^�S*Ϋ���x�#�=����&��x�ۥ�T�5H���;Dn��/����ՖjsyP����ˌ����	%Ut3Y�<Ĕ�2��{L6���>p��OdX[��n��$���ԇqM�&e���1f>3�Z�x�t$L1���l7�B�g�!�<�)NΜ��N��~^�Ͷ��HӠ�)��F�Ȥ�L����]�� Zq��	�N֜��0ڡu��h���1���/���!xvDn�)$ěG��w���1r��n��1�Q�.*	ػ!y\��́9���MvҴ��:�(��H�ɇ�J^�x��F�1���X�а�j7A�p��Mb5�ROX9k�v�)3^H��@4U��F;L	�X%�D��+��gAf%f)�r��dY��8��h��Y��n�xիë4#U�(� ��\8Ǜt�؍��Y�aP�����M��c:������qqsA* ���WB�I}��$|�S�u�1�״n}��b�Z�O����~�9��|a�_����k\��P4�H�+=l��e#X��X��)�耪>��Q��h���d�ua�=��ϫ
h��Z��~])MLhh=�8�{�,Y�3�� }�+3�#�W�-�<�w��]�ea<�[j���\
'
�Da�j��I�8��s�O�4��e� 0m֌]��oڲiŻ,�5�A~�# ��!�C3>Ϯ��Y�Qu
������]Y �ArƘ
l�H�ō[�^��N>�
-/-.�\"\����S�Є���!̂W�VG��Y�8��������GhI@8ol]�o2}3+.Uo�hN���`���KYdd�S�x��f����q	��Ip�_�F/f��O/g���)N� ]v���`p��ؐD��*9V;�|�_�m�v����GԈ�C)������$��z��<�����gP������칰�j�	�������a)x���J�-E�@�p�ST�/{�=O53?�w� wU�X�	�t��[�8��H����z[`>�ռr���8��T�#7��:��TI��nÚ�i�+N^A�#O�d2wy!�j[�\�/iЄ�yŶ��M�r�&S�y�i�'� �KNz`�Y5l5���9��*�KoQ��}��\촊n;/�+1=A�Ng&��	����o7�c��u�s�a�Q��*�$z#Ųᕺ�e��!�����o�v��M/�\�{����ռ��m��`��o�����Aa��j����vO9�Q�ւ�AT�5.��t�5���w5γ����>_hya��W�]F���K�<a(�� �l@O�-?!�||&�J��s�ED���k��6�7�9�0/(��(����R���险���0��&G�ǂ��B\i#Ħ*A�䳛�K��O���_���'���G��pmH �KH�I6z��YH"�~v��}�(<�yo7�Ť��/�QWd"��Q��KǨ}�k�u�h�y�Uv�n���8#Zu��y�(\T{j 7e�ڱ��X
��m�B�w���d�+��E�+:w��)��a���:��K�]r��,':�g�����Y����[^�G����dǙۅ�X�'�k��o��u��|B����@hpbz�����êip�B(��Ee ]����zgu੆.��~i߱%��Q_׆&���l����@&�K��}�ER�ܱ5LBN �;�X�>"{�W0i+*����x-}�8�s`�S��4���j�]�՟��?�}
c7G9�
~B~ #u��{����٩_��7�ل<� #!g�4Z�N���S�b��ǾF5���~}�	�k�[��+NV>ZjAG�#��'d�K��;}\�K��ے��*���\�]�7�%��]/�~+� y3����I���Q�쩬B5#��N!�çY��x�p�r(9u���������{q(�z�i.ږ����n�,><�~=�m��#�i��دeW2-��.���x�ob���<w�)v0:��_�lX��u5�t�4��/:�R�^�\��t�1��Q�%�\�4����&�����V*��ĐQ$c��e`vC����ؚ[#gh�㎮�+�Ӎ��wM����殅��1�I�S�5��Afg�0�a۷�ͥ�UL�Ҟݟ{9��l*(`]K�]�$=o���F��N�c�N���HV�jdSw�1�j��M�������6���T�!���gV�&E��n.e���4�q�;~CR]�{g�˫)��(a_�1?����//�|7�Fo���]?ri�#�z�r1����ȍj:��6�f�'���_	C�?|Lք^r��~�*VB읽�`�"#���Nbt����]˩�e�a�)ٶO�����w�W��� ���-��H^o�F!ø������ �(|���
.���I�����O=dM$+����_Hb�Z��kt�*�k�
�޾  ��"�ǧ)V��4�=�3����C�"�7Q���ς���F_g8���b��i��F���/&7��'�#��ae��C��z��\o�ל�"k�=�Inp�D.�'s��XE�sW	�x�Gv�f`���k"�hCm�*�a�`GeG��?p�Gj]�3��G�$�h�Q���O���e5��<o.ǾN��*hG��ϩ� қ����{��
�[Z�N�D>��JDV�S9��$����ZJ���y(�l�I�d��BG�9�f���}^mP8�	J��l
��"HW(i�teu0S�V���$��}5�TRبb����h7��C�� ����<���ZťZ�RY��f�!�k1�E�S�S�C�rD��Oci6a/@R��q&\�5"�a���tb�j��� ��Z�'z'D�����c����|9��>uN��P��gL�+��"G�w�`���*?���LB)5���0�b��D������R��=*�L���~jc�4 a!%gd���%�v�#����\�˾�����q��a,�\���ȳ��l�5o/�����20p24����}�w'�ե���P{|a"L$���~�i��� K�ы ��� �fP2�!7����R|�0�&��<���zT���>ì	͹4kՊ{N�4�j�j�Tú��k`�aD�������RS��	�C}�W*m}�7�ޕ�-c���w1�[�jF	��h�):�c2Dr��:��?FԹ� +��gׁ�o�#X1�ˈ# � ��=6��ɦ���2�� "7�me�p(��ΨIJȊU����k���9�F?d駀b�G)j�}��k����n�-�Y�������� �a0��m��-ŤaN�����b���oo=CǱ��r1�0>��S���\�O��c[�XtJ�@�VT o'�>eZ�mWl�0s�َ[�����MJ�LI>����+����� I���.ڕ(��;�,�m�5.?�[N�B��s�s��A�~N6E���W�; �� CXǁ,��kn;�ȇ�]kyn/_*\�=H���������p���H���r<��:_�<�x�y�1�����R�!�C�1��\�@��b��+a3�J�v������y{0�l�0���`�o�r�Itr$��[�N+g�z��ݼƇ�Vk�0����������B��h�&����I���H��E�S*u���3��Y_
��_<x����.�S����B�:11pu<��:/�V��uy0q�ҡ�����k���t#	O�mԅye�!���'�K&ݩrtT��&rJ�6���<ܥƽ�����B�r��"��6X �ϸLGA����Q]�|�T9�Q:���h�M
���b9`g����텊�v���B��m�̶T�r�l�SЄ A_�'D{��3���kI9� �
g��^���d��O:��a++E3uA����#������8*IW��@M�'�o���s�FQ6v�PJ)��|T^\?���[�oG�n+-:�J.��{�\a)�qPa�V��8v�O�F����{MІ���"I���������1;���Zb��V�$cUȢ����Իt7x��frE�����|ڢ� Ϫ��n�H�顧�� Y.���#�d�!��Sp7$i��ӿ�����@;;���_#e��ߤ�i+�ً��ԙ\���s1t�iY��� i���������y�F>��C�4Po�)�3a��l����i7ɑ�TT�:���ސ������NJ擭�T�c�v���Ȉ��tnǀ:�X��ux�I7./0?\Y�؂1�e-4�2��8	"�,k���̨�r�Q^����)F�c�-9��M汦�i��r�乄@:l
dd�a`�>���_��Uw�0����D�V�M�s�V<z��M�( ����Sj���YB���`�h�����O�m�u/~�@v�������0X$���p��ֽ���G'î;f��fh�Ĕ���X��sy���r�� G�_v�J�2������8�I��`K-
�h�s�$;��lCy�8k�Pd�2k�Q岦 [㉯���`��F��`��^�9"_�����G#5��07'���pg�ƙ`���*9�J�S�����TM�7���4��]���S4N�8���(��Ys
s__5�ַ)�;�~��\�,�jy�r�􉤗�0�b$�V����V��q���<��ZY���f��v/��K�=� ӭx_��=�vG�:#w���m�dX�4�<ɜ�΍2��&�w>byr���=�.�0���)6t���T�νaF	�g��0��v/�I�T[m����<gmx%��H%&@��?���8����nG�_���#F?����&7Rs�	�1{���xR��|� ���Yi�'zl�̷ ����+|�0��Y��v��j��hu}��y~ �X4��X��\M���<��������'7�!͉�Mw����u�	���!��\���욳|S��%�,ў̿�0隡R���˂���F1�7c]痙�9��1Z�Fne��Ժ���:7�W��Ȅ�]'Ф���+ު������z,ٔ8��}ӜT���{�+�'�)
����z��O%�����M@��0��fc��9c�k3Y�DUk'~iN�4��l)�v �lvH.Yax����w��y�-Ͳ�o�Nnv�O�|�^�*<ID�@|OgCU5�*���y�9�t7�:�v�#���X�V�N��Lb���ml
�d�;hI�Vo�rj���MH1����B$W����	�+io�d���AN�^YA%���.6��r�oY��/��}�%Y��A��"���y�磆i����YER���#�ځr�Y���k^�F�t����K:����|g|�$�Eʰ�`ք���`%ROp��HJ1�\8�+���+W���u:e�4*�Ӌ+H ��$�Bo[xZ��'���������
C�+/��1�HJ�q��#�B4Df�^���v��ꯍ��h�����)�fls�΍���r\�!��͎���=�1D �X��ۙ������Ҥ�U�5���z�������(�0U|�	�E�w�J;��4�����c����-@��E���9����+^h^�`u�2�@Ӂ���5��H"���O-pF�*�++a[
����k	��/��R7{N�6�H�_����:T_땞f��b*J��)Q��Q��i�R�F��<E�M	�YHm���,�۔H}��-̘�v.�1��S�+���5��Y�����GX����턼�*Ȇw"�c�͚�����#À��:51�����N:b��ȹXx�p��0װ<�!`��͍�V��U��u�b1ƒ���J�o���3rR�ͧ�	$��U�;a��k�"���d���T3q7�:�ƒ3 E`�)0壃�Y":��7 QoM��S�P}���'��~�q�����A
�d��:����+����»�h���2n�H=��;<��� =!_ar5�}s�S@P��<b�ۉl�Wipo�c����	���"��L���Qr.����ލ���e,��"  =�
k9D뿝A�}�hv���q�6��w^H�lˍ�i��,'�R܎V�����HT��&7@R��3%K�x9{�aqk',`^�!��6$&��g���F�����_iVO�_>�	G���ߌy�8����Ϻ�E��l8l��n/T�h�0��d2�i�2OT���*��X4H+'��/E��!�2�Z걊��;����ή7ݢ�P����m�����j�x��������z�*�â>c�f�Z�^�'�թ{��J}���K�l"3�e�ѿ�Iv�<��-:���&ӏ��?}M��5�f˿{��VT�&�����O%mn���
���e��Њ7�4�fJŎ�Y���]�^WU����ho���N����1o��YqC�H�/�._����Sra�֘a5��?�-�	?i��[e=B��0��I�I��egrh"�؄SC�%�}f��6Tڴ���q�@��UG��3!!�k'X��]�(��A�Q�F!�m���Ƨ�Dg�������5lll0X(8���c��ЧO�Roe7�r��,J���0�5n�xu�����u۴���$:�����ձ�Z��6!q^�+�^�����7MT�Q�ܾ~��pRhҾ�x��x�g��b��%���ğ<��x��po
�.�=#6��	�-z��;b%Hz�1~Zۦ+nMu=(�[Ag�?&M�X�npR��)���LP�'��L�]����j�V���<m��?Uq��(6uY ��H3)ٱ��WR��^z�,��hm\ez}i�n�CH>�H�.�4��?Fm��P�
�z����sJ3=�k���FL�GC�׀�.����6{sW�Re~*���A����K��o���/��$A�W)XϨJ�]��/����s�/!i�L"����i�]mr���i�~q�<�W"�}�c�xv{�~�P���d/�/ϱ�mJA�Yv��5�A��U!P�^Y4NWn E< #t.]�]���'����z������i��kU\���E�P��J�/�(��N���.F~��Ca9�\�G��HO�/�]z�W3�b�m'T�yMg
^'�_�6�@ppV��АuHN0����lh&&��E�7/��]�Gp-���x)����:2�֑��5��߫䥨v�ؖ�qq��g�Ȳn���i���;;4��r�n\z@�>V]��HX�l�7yēc���B���i�I�*����w�ۚۢ%&�C�ϨK��:��=����r��k�١�l5��`wHl���=��Oa��q�y��WS�����?45I\��#��zQ�;N���x��[��\��O�+�tύ�o;h_*����ʱ��:c�h�$�A�����n.Ɲ���⃳M��z�G'KG����ڊU�P�3J�f���v>���&�'n+Y䷼GA4�	�diY���S6�`W+��)��a���ᬱ�m����Ћ���Cs���r�o�Gz�����c!G��9�R�y���o!a�"21�r������X�c�ʧ�e3���G��2"�H�m��s�����S�r`(�bEy��Ȱ���~� ��<�z��vj��/����Ģ×K�43b���k�Nym�����=�8s��ѭ����Z��J�:�XûHwVإ%񼑠�o3�w;Z���q�<��$K���՜���/�L���3"�̖B�(͖�;�Z�7q��L��¿S�%�{��5���R/�1s@�.dY�tkYi�E�ƇG(\�]'���'�ʏ�wv@HQx�_O��O!&}v�ʭ�#�������S�G���&��L���t�c�Ü�IwOv_��
:l��f�ƌ�'��c�3���p��(�RVo*��߈;��Q�
�m��WOzlG��p��ݬ-���4
g�lenНS��>r�^J�+(��Qf4/�Z�ҒI�BkV ao1n�Y�U���myZ�_����]�P����ūi��F������ςhѸ0��,ٱ��O|zl�I�#c�6��Yt��ج���mIr�m+���ɜ�� ��X��i4��!��c:[l���P���?�Y�#��y�؏���S瀻��5rR>�ԣfX�`���/����9ݳ�6�?�p�!K� `i	L�(YN�W�-��1�O�y�9mlh-4���y�xj���>�1i{����3켆C��@�K�MY݀��F�|��f��K_U#���NP�����C\��Η��*�k��腥�H��Qձn�:^0��a�� ���oވ�j4����XmDL��pK�l�n[0���C��!̦;N���hzؽ%C�D���FlBC� �Nk�E�R����O��iO�kQ��H�����P���{a�ݟ�����V��L	0Dy�(��V.Tc�%�*C�w���Q�A���
��L�(�Ӿ���d9Uf�ؘg�.�ą�Vg�)�K�z&�j����2$f�]���_����2��z]s� b�T+��;ə4ҩ � L��B��w�3�։`�$� ��+��t��T�wq
6�R��Ń��\,���9�2�Kn)+�.ra��擦�~Q9���d� ���Iin��-91���tev �%m�A_��`�a���{O󲝌��<�3�qq(���e���|�m�{�F�_��L]>�,��w��5l�aG��)lD}��m[����7W����t�ҳf��ľ.PJ�*KX�� .�\`��y���x�8O����'z���>����@�� 2e�����0
#5!.X�FJ؉>��pt6�k-
]�j�Ft�/��r�i����
h2v�&&��x�}��-��X�G���ݬ����É��3d&7�/(�x�� ����-��dg�_�.�H(������WoQ]���w��R� ��o3���	F��Ȍנܞ Ε�� �%��X�r�	P��R��&�z��]�����p�G�̸}�j3׆c�r-MA����¥��N�g����֌v}��0��/IPp3��o��澱���&��哗;\ÏZӚ
R�cG�I���Vք��-f6k����U�Q�I2��,���l�|��SR_=:op�/Bzo��M���b�V��^�~��:�!�GҪf�N��L���2s��:H?IN�'C=ZA)*������<�d�_�5��y�gdbʵ����qK���������!'���Kj���wo_��M�Q�@�`��0�ovؼ�O��f�tf���:�<��.��̧}�x�x��C��߅?��j��_�%mq���5x��Ul��p���|NJ�j�Rز�A�Yƕ�^����7Zf�MC�<Ϩ<��c?��$�eݔB.��bV��I.|<K�S��QY�t��`Y{�埅2� ��H6�����*����lDՈ�Oݕ�BvW��J���Y="��  ��F������?���'A��	��O��z���w��F�sd�<�v�(���M��'
�'֖F!��׼<lv|.7}��%z�N�AyJ�=8VPB�%QE�3B/��m%]?)�����ӧ�>��K�."hl�D��y�ؔ�TE�ʑ�a����_���`f��7��pY���x?��t_�"�5����ک��S�Ͷ>�)0e�Q{:�Dj�D)u��"v�cwՙ/� V�.��&$�#�<-#0�A<��d�h�K��_��!��ä�����\�����n��i�霸1$6�1�ݘ&Qʸ�:��	�3?k�/��q�6��vG�Uc�
��r�+g��?�����KZ�g`�֪S�o��[�e��a��4(Y-wdX��q�-������M:p�l���_�R~�RJ �mI�S6K�׻>L^<�ӟt�����Sԙj��,N���-�U��4�m���zL0��7u��x�dsR{Z�S��	�"	�����T�1?�]4y�*7�䰆�
$ǷN2֠O6�Ղ�!���e)i���Y.A4�Q��H����D�z� !h�'2�y����Q�SMr��?�юp����JAī�%�O37Z�M#C�K6G�ŉq=[�ޜsx�LS�S�v��t�� �r�������L�4���A���9	�������*�#�1 u#�#�G�ť��Hފr�����n�Y�p�e0����FYjm��|�ƾ�[��kJ`Q��|��#��N8r�J%��\/���wv�0Y��,8��89���_�F�S�ۀ^�_��֜k|��禔��R(5Q_��������B��wx]q6�&�8��4{e�c����pYEyp�\|���
�s'�ъi�2�)L�?�����2��<ƛk/du�� ?���]�B�ϾWo���G:�x�Q�^���'ؒ
�o��.������+gޢY����^��bp�Ͳ{�AR�~���x�M�)�G�#��a��_F�bs�f���w#AӬ��ϫv�~:���Ց��u�O�Om������[���rd�H�������\VS�X��1�T���b#�#7�B���iL[����>dм c��d���l-���]~3.x�2ﶖ�ٝq��T���f����1���ӗq(S�7��|J�LKQ���+csq�s��S�4�Gcs�h�Y����_�2��/̈́��HV�,�t��e��Kg��`߯<�)�Z?�	��ϛ$���	
P<@��� �۾Ċĵ[�2e�
W��g@g�y�x�4���*|��jT%
������ :PQ��K�ZW	���k�!�_�֥�!���ַ8�r�<q�xSc��lz>[\�|��`dc�`��\ƽkO�������������9��m��4^�S�J4��e�jщ|�6�|:�vp@C�F�7r��"�N�-}��>��A��� neq�A>#�6 #�3���P�}�����T�WC��J';�5k�9|p��^1"�֢����O���(��f8�)l��l����=����ឺK��%��9=V��#� �����xar���,A�s��7R�L��?����in�h8ȗͣU�W.;I��-�/�2J��,�lY�KF�Q�zNq.��eJV؞�6�gq�+'9�U�l8�u������Y���9�W�v�U��ʰL$�����	S�G�Å���0-��Z8؜�ɞ��r�l<}��{:����w������N	7���	��M ޷�l5�1�&Ĳ�Vʛ��1fִv�X��- �z7��?{�FU���}�*���!;�;�� �{l|��N<�x�5Xܲ%�*��o[��H�^�夨�'@�M�m3��*�:��,x��$+d�fqY�Ɖ��h�C����7���B���b1 ��f6jG��2F�hR��)YدfL+0��'��!j��A�r�y%.gM4��.��2�����fa�~���
I��l<���#��։D�)�@EU�@q�ӧ'�����e��+j��)4����
��b��z ,P�"Z��;;L���~�o&�ǩC����qe��r%י�T⫸4�`ڱ��O�Z�ֳ��;"jHX���&1�[?�V=�[����`�k�
��Z
��{��]����^|�f��8�N��2��)b ɍ�<���[�������?��G�@J�-[Gպ=��j�)��! 5i�떄�㄰CBc�.ވ���~3c`S��.��D�h�>߭"H�S+V3��r$����U%ʥ�6�P���K�3�U�$8s{��;@�@��\�o�\(��q��5���f��\�H:m����*@\�~�T蜱��\?Ԯ���;
����#C��ۭ5�8@|9�N�fP>4�qtZp�8Iq��FZ�;��?��,���8�,}x��Y8��T|@�c�>�~?P֏�$69�������1_�,/���l�!x߷)�8��L�
�;������<��<Pw��Թٹ��j~��W��.-�6h�
�ʳR;G��!֋ٙ�G]Ee-�tZ�J��#̶?���� J���[զH51Q���KD��&�԰ǁ��#�p3M��>sx�i�h�3���f$Y�8�/w߹<��7��<yfI��q���Pv�!�O
3|���g�I��8I��ro�)#�� v��R�m~b��ZQ���~�B�x4*�C,ky֍��/�!�cI����Œ����AK�ZE�AB��Az>'P�+"S#/S���|�ߘ�5��������c��D�?�f��"og/4����~�h[.�q��W.��Kd�������x͊ݎB�@���,V��t���CB�f�9-���Q�P��̜G�M�ꮵ�&�N�r�@��;�G��~�3n(��&���K&%�
WXw&�4�J�:�ѷ �e�~u&��a"�L{����J�6$��U<OJH�{�`�KH�.v�m˶���M:��8��*&Fs��@3�8�dE����u�E�_4�4�<6��� ��h$���;������zx����4����)&�p%Y=�P�QL�+O���;h����N/3k���E"v^���]k���� [VU��9�׹O�zvТ��'u��:w�f_�g�=+�Y��-ʕw� Ύ�Q��g#S�6;��
��X���GOZ��B� ��N�B��h�WT��T��(��f�e��ĎJ��J��I�_�0��`��)!����;7^�Dсg]��Z�v���{R2�~�ҿ/3D���jnt���K�C�n����R�U;�1��~��\��*xRc6y�v �og=zH��P�Q��_�< gρg0���� S4����äYzO7�V[�7܁�����`7ٶm��T&�f��g���W�0��[��{[o\Lv�8���_�����\�BP�kVT{�F�'u5�����Tu�P��vr��t\'XՕ9�58��f����:��������sRW�4��{��9ZS��R��7N��	��N�t��uj��o��̈�"��c��S��v�"B2@/�gu-zbrT'{'�F=<+�Oq>PaJw*8�9:7�K_AH��<�o�_Q
r���$	���h���8���="}7����˃$8��J�_��R�)��g�E���X9~��Mu���@�n�҉7N���$�+n�d�|9S�6tq�nn�e���:����t��/%�,-�v"h���87H㋆�� ��$�tIU����
�~C	��B ��x(=� �;:V\	Pb=�K0V�_Zh6Æ���K@@���ؘ4���6r��[���V�9����M��d���o��Mnʤ�3����3\�����
�/�r5�{���{�d���+�4��L�Lձ�+~��� W���k�/�=��*OQU�P!���p��{�uެ��D�<J��56�4�c�f��2U�����sT�tS�I
�����¾z�{��W���"\|*���Pn�a�~%�Zd�����n!���$�HmS���n.��6wl�mk��	&�}�hKM7���j8w�{�xxk��E��
x4%${*$���0WLh��g�?�5z������)@�&8�n���f��C���v$��G<M�늡�����7p��Ǭ]�O���C���6�((��-���(�s,-{T����-Fh�ؾy�a��;�ӸpV��v�Zc�����q&u�%�Q�|N��1F�F${ˏH�F�3wXg r�: ��X%��-6GI�_*e�6�CHҴ�� 7�j�+�;c-�͊�3X�so������.�I�x���:Sh0E�Fl��!It�0�umJ�a�ߊVRf?|����k�j	�t�X���r���"�E�TZ���sOD�G���{ݼ�X�G�;K[�c�0�}�DH(�Hl�$׬�jt���'<g����s������A�V��ֶ�3t�> ϰ`DW�,dAb02���H��,|o�D��T([ȍ&�2��'�C�^�:��~��l�TC0a�{7�}X/����*�i8�{%V�z~'L�k��/o�_*N!q�3�>�lh(AJR��Z��˟4�#?C�%�0ǝ�7�Q�*nF�[�-b�#�HwWLH��cr�wZ�Ɂ�@������D�X��8KM"X�l��Mp�g��}&�7T��Sؤ�t�'8=N
�����Ҳgl�,s:PA_al��=tV�4��[n/�EGy�P�sUOu�0-�[rƽ���3 �H��ѷa�{�Ч�V�(��)`8�����x��%�!R�y\MT�����\ɾ,�]S7o��mO��Ӕ�|���$�
��JڐsE*�y��}ڐ�}�ϸC}��ڑ�V�_��������\?������3��>�r:$b)�~�~�u�Վ��Ug��Ho*4�
��0���w9
�Af�x&h������Ͼͱ�Ռ�J���.i֜���9)���B���,�^�����WSM��u�0�O�5V��@^��
�t�d"�& �N
3Z�N��Gh%*���$懮C}�m�~����Bc���m,�d8�ʓ��Ih��~ja�}ĲZ����9Ţh���Ț��/��E�p��@_1̌B��n�_���	P�hj��"٣���+ΩK���`��V�埐O�h�/3f�~ؒ��#����(��- �A�/� �E����=�Œ4<E��<�۲��Ie��%q���HFnzq���ܷ3U�0����g9k�l�0�NE(RI�ㄕg�z2��8�
�)g��A�g�gy��-��E`�+�KSCT!?O�*��+^��z��tn�pO�����g SXw����
�ܥ�cFz�kb���#����px��s$�l�񛍳�l�����Y�xp�D�>yQ��B�'�Ո�Ǐ��kV��W���1*f�M��Y���Zt�ݽ�"ƥx���ڰ�J,<�| X�;k�~g��N�_ٯ
�����㩴��0sU�Ԏ�E�'���H�,�jq}kF{���3������
�p�N�t9������8��� ��x�Xtd�$���1)(v�?� _}�'ጐ����ˊi�}|�w�����-~<Y��T�����Ji�.��	�W��MTc�(��~jv��]��Y��΍>C-��݉r����+�x h���`���@���ˉe'_Ç?���1z_V�/E�Sߏ>�o�_�|� �F>�COq��� ��}Ȯ*{��|�k��h�y��7.�9�^}J�Rs�C�:��iߔ�WJ8���d�����O�S�8�W�|�r~�Tv�}9�1����G�!!��.)�J�ߋe�G����>'���p�mG�}6QE�2WO�D�D��S�s�IձZ�M�p��X}��5ߤ���Z�J�v�	�s(o��&tf_ذ�-kU~hHT����UGD$��c��k�E���D" ��c9��ѽ7�;hx?���+���50a�7g*ͺix���դ�/<��݌½���k��n�RC8��'j�vT��'{N.��A�U���)���S
O��FI�.�z��(��=�v&�aN|�����h���A�tUv�w��Oq�~_����S���#I���ͷ���s���Sb�'��R�X`�Sd4�pj �����,_�!�
&Y�ӪK�bP���֌uʴ�Yh�|����=u~c��E��*詜�ĺ(0߼��e�~� ;��RmH��3[����Hr�iFOԑ�d�!&6bpY�[0�2�{�+�ަ��;	�jc�����X�/Qk��Ł�~����Cݘ9
�KC@Y��l��
|_]��B�,Н����^|teNc���/5�g�2�ҍ���F�m�����E��E��<��NvEw���9���d�'��N��<b�o�CxWP}�e�W�i����e' <oT�2I3�l��SG5O�@����$Տ��+�d�n4r���5ܩ�h�;V|3���wo��
��{d��-)����sK�pb�m�I�ìVt6x�wM[E����d<��R���zb�^���h�_�q�RԜ��+7+�N��[:r���7�_'�bp���X2��"3��bdhq&�ωUǌW�׽���s+}���|�I��l	f�c�ΗM�%�wt��b��>@����KG4��G,�*��unwh���V��%�VCA�;�j�á����]���t3Z�Ģ���#��k3gg6ʯ��Xz����ا�p��h6S����A &��{/�2hމ#.È��k��YR��I7�?�Z�w��̍ig'����� ?	EW��Tn��q�Z��~�,���� �3�?2`+�&��TK���ʁ� �	5�_5������;í�+���㠃����'	�6S���Z�|+�: �]���w����_/�f��i�%�Fvλ��E����˸��U~T3�v��pb�}���/��{�9c�B�iwS3n!��1�Q[:��,Ԩ�'�r�8>��W���&;E��6J1[l	�ͷ[(y����5�̒nl�~�`���{�P�6�X�f��8#��5:EE{��>���C�.�Qw�sCQ*�Vdl��mK�O��:cU�OG�8��z�i��a�������-6���!�"h:n�O9����x���iP�7aw�z.Vx���/s�YI���ۈ���Ĩ�����|l<�uc&c�%#�l@������|gt��'Y�[� <]��(�jW� ����oWp)ȼ>t�\ԇc'f��K�F/�[�Jg@�!%�����"�Dg����f#(��X3_�ޞgh� *�c7"Q����ҧ����8��Q+h�|�*)��$���OO���0����S�@١-onji���+{ң.{x�S����{%E����$���Eh�>4هM�]�Nu��ʀI'u6KT���is2=�����'�*�I�oS� �Pg�N�q�k��0�d@Z�~{�C��.G��> �s�#
�4Q�4d;%���"Π|7��d��x���W@Ү�W{�pr�DT[����~G�n�Αh2���Z�/�����K��-zл�	����N;%�pY�Ǳ�ۙ����,̴��`*�x�8����3+��Y�3�)�K�IK�m-{��(_��0ձ+Lr��i�3z��0��f$6��8�i�A�N"�(4bb��7 ��x�3y��/�o��D�`���h��C��6g4Qr��Pɵ��թ`�'�ٙ,ׄ�.'�����+*r]�P�p�}���U�)���0аv��v�����v]�W�n�\�t:�_�%�e)��"��3^�06P�v�<	�mC)f�\��n���-�Z���>d?�),r��y��
h��b���h~�;J퐟��/>bh�(m]����T�����A�E�� �.�#��^mORT�;�2�V;&��%��n@&L�h;mJ�V����.��9\�N ��6��լ]\�щ7N��d����U����#Иw��i^���K_�|���9&�yu��q�ߺ�d^E�K�JJ>>k\i�����q�x���49�R��񂟠٤��f�Y�Y��[�О���D?�!F����Rt�q/vGn@�K�ti3�K���h��ݶH��LM�-��g��$hp�>�9�9����`�R5�Ҟ��_�S�厮�� �"��~G��%�l ���|��a�=yF��kb��JN˧�j���ɭF�t#!Q�~����w്��87�1eG��&��[��럵���/��sN�o�fz�u�Q�$R�E�_�wx����{U@.�w���.<�6F���p�Uql9i��J�1��� p�nSc��q�d\?��07)��L�9�*�i�#��!1��00����7EF�
�gJ�{�U�h�q-�R#D�C㵭w�4���R��.O�zr̆n|5|sd�b�_���D����O y3|�-S'��qmLMLa)չ��o����3X3EV[
�>|�}(Eɖ �+���h��)�ͻ}��i��]_�F1��Z'������!�A�6�P)O��~+A�@ƟvB1P;�ܕs	������w,�I	�1�U�����.?-��=ew��STZ�.��
`��W���<�uT+�ӵ�g�=�]G+�<pƛ%=����7/ƭԻW�9�	iz4S�A���&F��w�#^�N��{>XżQ^M$g@�XD� 	*�̉xJ�0m�(=?���'�4�%�L�n����PM��V1g����Ƽ��zc�E)K��k�����`�d�Hp�+k����!���gu�'���=@���ī�$�DY@)7��^�Q���~3�,}���2��c����ؘ��w$����_�38�ΠDZ�$E�F���]��-�-����Ʊ��	m}5���/�|1Szb�M���B�~���}��(e�p��>�{T똹���?Bظ6��ryK&sS�7~�O�b#����t%���H-_�B�*T��ׇZ@��œ�a�)��.�GM_�,�K].�-������<��UC6���L��\�\�an��x��N%\�K���/dG)w=�9���)�NwBH<G�j� �q�x�/ ��Hg�0ܴX
��3CMo?��?bX[�cd��ˮ}��2�xz�"~�uIf2'�瓊0l�5Uv�O�*��"�D�6q�*���(��K/��E��>;�ZY�^B�$hŰz�a�2��V�;;>2C�E��E����[BQ��j��՘L�
���S�"}�*�	����_�~f[68_v�Pctk�0qm�."���Ǖ�TQ��X!{J����C���KV@��>	G�U!�7i&��Oʴ �)U�yN�#PG�u�΢"։;3���y�!Vb����u)�^���=�Q��H�rV�<�k1����a���.�{UC�eb� ƛ%�K���{1�@��M������Ļ-a���k�|�~����*#�ԟ��T6sP�4�}�&���%�}De	B\h�8���������6�k)� ���2���U���
<�Ω/�Xɝ6�J�>KsN�	HD���;�N=��Fi�E�sɅ�f���/��|@1�3X��ݩQ>#��j���쪅׼�x��B��zL���-��i{�v�2Co</��ex$���jF����z��&� �PD�`��y���͊�J ~�Ӿ9͠^�E`Cs���}��\&rW�J�E��H��M�����^��<�L1=�3�C�9[�];��{�!?��0�H��NɌ�=��-%�b,���!��kwM<m�%7�ym�6� �E+r�������_k�N��!�=���BuV�!W',��71����-ǁ���hm�#	�jQW�՞Z�r��v���O/dk����ƨG��kާ�����(�>�����fW��},�1�V�9ˮu�ł-�+`��,E�x:� ����|��8,Q��OTFD���j���f�S�7?ض��(s��)����I�y�4�DW.�)g_�����G)g�����9��]fƩ�.�$z�+5e֥PƆ����&���K�r���j=��s8�5��Y	A�{��B����3ty��6{�d	�d^D��~�JF��Y� ^ ('�<w�-�.�J"��l�����`o���_�,��?
慊� L�A��)����</���PY�&���Z���o4*�ܮ�q�l�/�5U�/��	�$�^���'��ooG���͊�b����/��0���m�B����`��ǅ�yVwXUvD����c�d�,\l}��#�/	�?��ɂ����1�|�\ʰ��6�5,��g���RB���y'L.g}��\<N���R�\U�Z�l�뙯�'�RB<ݰ&��Td�}���g�d7^W��kDʵzpd,�����>�N|y�D��(
�]��@V�Z.�f��Ϲ��{6��>��YM"=B��<�����p��Ce��¤�:�N�^�_S-Cp^���ӹ��^�G�s���)��'Yό�զ��J�{���s�9��3�h�#,�'`Q���u�ߋX��!��<Gb�.+�5�a�HI�N���BD��p4|[`	/�PU2Er3�W�x��Zt}쩷)eť�R&������&u�*�Ԅ�f4ھ���b�\<�1� Ղu
!�L\ځ��略��=�����5��֪}��w��Mڎ�����B]��a�!�+9�U���!��xl�NeY�`�[IeTa.2�h��$���C���q�h��#IF�G��K)@)C�u�jE	/�6Ӭ5�=�K�9�ǂ��T�d
쳗�Ay齧��2��ǲ|eK1O���!|W1�����fz�	����+�`�.e�L�X�3���>�j�M���w�9���'|`^N�8�`�Pdh���lP�>��,O��wT�M�R�F�/`5;�玚��b�n^k;l�-G1�Q�z8׆RH]_���]Tش�y�tU���-��9�z���6Ŵ���_:�`!��ߍ�S���f��Q�)���B~�. �ZH!`#�R�N��;\Y6Y�CܣAB����JV��l�ef<��"#�҇ů����u��V$�>�Ħє�P�~PT�ii��9�_��Z|���@+
0��@�Vkf��	>��b�͇�
a��Y�|�Q�=h��-
��k�kt��@��r!���H$�Z_�2h;߹F�]��������d�4By%�ϙ4�.TqK5���&[,�����-v@�C������~t��G��[@ZƋ�D����~���v�jGk%�R�MۇHn���Z�;�(ێ���YGP��h�8ͤ�m�9�s�5��Dv�ݫ2��hSJG����M�^�����o�yjn�Â�M$ݼp�t'�4o!A[Պ}��Z�jAr�=Xޚ������b�J΁v�����Z-��8�q�|�7���4�i&wg�(K���`��º�&��,M���A��V��fw��%M:��3��#��p�x�&Z>�S���%t�!胞|��r�3/oC��Q-HL���`��́-�f����}ɓ�c���l�m)yV-\0Ł1�	<�[���g���;o�9��G�Ze�{��V9�+U��w�~m��0��������>�S�V���ܪ��D��Ձ�d�u\��נ@��\ (�Qx-�h��SW���a�0�.g��'����))���}�7��h����5��C�TC/l�/���k�˷v}��ء;��s:��Xn��Yf��^Z{hIX>�s�ᖨ�UaXEL�vְY2��ir�9�
[�	�Yylaa=����-����h絵�~�Ab�KB�a-�5���1�2����$,e�ތ4������ՒX^��
=؟6D�g�w 8��t}@�U�R��#EH���.�l�5 �Z��S���R����2�ࢍ��۽��X[Df����,��7p���먝!c� |ӡ����ztqBr�+,�^��u�����A@��c�N�]�y|��/���N�ү	k����ֱh3�ܗTL�ɉM/R�mC������88���n]�.m]�݄e$N�1���S��C#Ajg=��M�S��%
���(�1݃��=�
E�A���D�p�Q�Мߋ���qTj����������X@ �w+VO	1f���L���?�4�´���r�U����4je� �>����A�m'c���o�]��o"�&�^�Y��66�I�;�O5?ز[�.� �S�Z��w���H�V��D���.����Qd������Z@�u�=5�1م���s�)t�"缸^�{ęxӏ�c�4^��6�3n0,Q�s�<{3���T9bW>�n���jJ���5�{����1L�j+V�.a,�B��ՂN~�� *���\C�m��w�a���1y����M�o2���o�+�C��P�|LME�&�MGa9šW��rj��	eX�1��8�xWyLvk[Q�	R���5��nA��ZR��7��N4>;Y���V����B�wV�����W�OK�iq��u��J� �"��5	��;�.�)Zpbڊ����U�c6A���iL0b��-���T�7ZJ���枬��WQ�(���L�ySf��J�G���[VV����~�Y�O((C��5;!w1Lu�B��623��s�iv๱����㯢@D�>z��4	�N$��+����4b]�u�w��Ҹ�BQ:p�%A��6SJr�Ș�>�"���aF�ß�ڱ�s<�NӤ�4�V��j�w�W���_�m���l���dӑ��f%�3bJ�n��ha:<S�3��C`R3��U�@Uxu�tQ/�����W�<u���S��f�M�o���c1j�貋Do真����%o��b)��m\.s�uW��.�inY,}�Y:{�n̟��r�8�[���Վ�G�GT��V�{83��KFFJx�x�9SrB\��+�9�%fL�9��|`�����<���>Xv4ůɂ�L*�2�#�P?�lH�Oi�2!�|׌^c➀�hi�C�}�;�S��A��<� �`��Q+��$_.
�
R0�JS���5�	�[��!+{��"(I[��������%�L�v�q7Y�#>���ǚ���v�N��s�!�fBE� 6��������&"yFD+ǟ���U8�l��� �>/���p0	Ea�>������4 ~�����xSy����$�="蝚�Е�OW����ู)LP���^�O�}��P�qa)�V��U��EZ��Ό�F�pn���΋����4�����KX*_C��3�-����%����pȖ�T^� ��VLw��e�Ÿ�:�{�b��0�p-����L�`�0��}�!�<��̠eIϷ���,���$
m8��C��wA�ATT��y}H"
}{���uQ�Z�Ц]���2��T��G՚>|_�2U��D�wk�P���;ؼ�[1�74Z�8��/E���OVl&|.!}ZP��;;Ջi��7'q�!ۨ(�?��Q���)��Hһ���=�hs�`��Խ����<ׁ��s�}�K�I/9R�-���f�ט=J�#��XJ�BL�99�s�P�nQ'LD��=N��W��֯�B����M�c6bxt<R� ��ӻ_ur��o���^.��9(�g�AnX:��Ρt��BR�;v�AH�$0��(��|�x)5Y����{������4\˽E��<��#�e�I������L�A65�[�8�{t�1nnO0B g�V"Q"��.> ���2B|}$��J����)XG8 ��nT��M�|�D�ڨ�;Lz'o�R��l��)3��?]�QG9ӓʪ\�(�-�=���V\#F2��7~�� �-�F3��ʍ�o��ŉ��ҥ�Z��OՁ�u҄	��hi�2R��迮m�Q�r:�W��B6�+DA�Q���EV�lh�=($��."2��Y����L|����N�n�2tC�)ٸ���	N�mP�����)C�g
5Xd�E(���Rh�ֶ���~i�xF��/8��-Sq�ˍ�6����"��J�&$����E�;����ҼV�Wi���ޅ:��D�/���;�A�p6k��zʣcw��-�BMI�4 ������gN����G���ͮ�Ҩ�ٗL �MP�ꐓ=<��c�Тl{W	������B��v[>���W?=٥��#I.p)Ej�d:��?���y@)%��Bj�ewp����ģݴ!�+t,]+헍�Kg�T�4�g	�c��d�Ђ7Q�[��N"�Z�.Y97�����y��yݭـ�6z�ju�^$��gO�O<��`q���d֧.^/0ԐXx�2O� ���v*�g�m����{����\�FN����]����Xɡ�|�Yr�褙�ar�b�� �5!4��a�l}s�i����_���|���1,`1�g�,�'A��f+�����I�(Wji�:�H;�\�:�����^�Zo�
R4.�2 �Q)'R�i��ٽU���p�y�j����J邯��kl����:,�K��V{�����DـȯQc�5�>�[R�N�QRJ<�0�̬p 0r�B�N�kuD��F��	�Lk��Ŕ�לr�Pg���!BS�m��h&=AC��Q28��q��T|L^�DU���	���O��*���Jn~~=k8���|�V�G��[���w5㋴������`gB�"S^�cؚ}GQ~c�M�����n�I�~���&8�H7�̴���f���FS��P�|�o{7��A	�x3ʛ�k����������Y
��mӻ0S�> ��t'	�]��:]�Y�pO��]0��֐C�n����RK�H7L0J"kzԪ,�g}�J_�)˳��Xp��|�5A�?
E��&|3籥�=/���w�ʳ�l�ýn���g����=�^���5X�s�$���i��Ӝ���7(�sH�)NT�����BzX�Q��8���jφ@���#li��=O�K(�Y����m��[�I	y0�^q�/�*��֦W�!� �7γ�����p4��b�_��:��i�
6~�f�d�f/x��#����X�r?p@��x�~��o�ǢH����JM���Ϥp��\drA�:� �)���4z>�-�,B���z���+o��x'ŸF�k�#�u"�[���#IY���q<OХM���+ VFq�y�����?�#��-���g(�Tq�J.�<�
G��S&���v/րi��r��~��V��.�s��Yk�I����М ��~�h<���«h�B=��� �[�-��l��m�
G@�oNҬ�Q#.�r�F���Z^lB�/��Z>uЕ0� %�mʪ"�|~�(�$?4��L����D��/k�+�nt�!��{A#���"��p��g�����x)�g�2!�Z�?�)��R��[����T�� *0^\��3�e�{&�(�����.��TBԷ��N��2��_Ms�!�z8_�荨��mX;2���Y;Q4�8)��렫'��F����=��A��E�GEH�#	B�kg[/����P�ֶ�>O{�K_,O����P�t���!�t
:��kLǰ�L�ߢ�1�'s��$���u�_��q�¹�7J��ޭ|){y�O�XbZq��wǃ��Y�G�ANeCs�p��� O�����������~gk�'Gp��.�$,v��S��5����8�d{���v�-EC���P[9|�"w�JCؕH#����6þ��lm�M��2��_%_N���s�Cl<�%r�w:5�2v���R(Y�OP�[r�ƅn��[F��)є�d�
ύ���t]M�*Vt��ȭ�ݕ�5�	D/`,�]�Y.������qL��Dʺ!�F}|/���i4�9yZ�����FQ�4���Q��j�Y�sM� ���ZΨ�Y�i�^������ar������{�N�nP
��	�/
�~]w�-�f����%4�<����bc�L�R�<� �2*�([-jj����|�Dx}E�m��x�T,��UO@�7	�R�hj��!do�j�Y�:�!D�?�r���͗�U�!�����DM?�aζ�r
���6��Jm%�F���S����:����NteQyh��Jϒe�K䐈 � @W�`���n�E^7{��KL�v#�q�#x.�e �wD�VQZ���KjS�|��6��g�`b�EO�8��+�-4�X��E!������t�N,w��R��U���	*�_;5GM�qv�j���������q��ÿ����H2��Lɳ��I���7��G5�Y�3�j՚���ҹ́)�Q����/wm�QC�6�>q�~[���o3�,��P�cM�@k,cPR�WuKS�,���O��M)O8To/~{�k��<E�+1�T�1���6��뜂/�kY-e"!��6+Oi���*��1ĵ���I�����C�c,dys6�?���N���0�A�}'Z
�{.�S8�di83��o���������	߱5�&{�;=Yu��h�u��_�~D!p�=Q��9V�F���^2p>N�gv�Kn����=��>r1���͍�T-��m��C���'� }��v.�L¦�d5\���[>t<D������S;�Y�FL}�����]t�-��*����g�*> ���9�k_�R�������'6�1���.���S9��kE��4�G��cq��0�n�Ⱖ�����ؤM��
Ѯ���=ʬ�;)��5UXg3&E�`}.xE�|<���scr�iO!V��k�Y�L�V�|'*����.���4�'�F!��	d�Eh�4�aQ� ��N����5�2a�DeQ�ߌՎkm���4�"A�?�ʿ%x��>X�ԋ+b�0io\�] B��_�f>8�]�T]4[�鏆�v�/�hZ_��v/��W���[-�\�!�|eg[_��C[(U(������t�"�i\��f	�U-�dXM��`����D� z2�G�&���3Q��}*k�&^` I��T���C4sd�+�C��J�8�3rr0��"�k5��k�ͩrg�*?zY4 ��p���FHj����F�h6-o�L��2Q�C�*���C����?��al��ݓ��_��ܕ�l6���M�+Cͩt��n<�+��)��
�\4��3���^�_�*IMH˺��ϖ�5�:q{�)���":�f�|��}di�m�ܕC�e������RA������d%YZ#�� ݅q&�&p{�/ڕԍ�u�=�S����g~�P���E��U��IG���a�e�M������d-GX=�,1�$��b���	���8�^C�|�0��,(>w�]/�[n��<�7X�:�&;��`nWz����k�/W�}�c�^�P��$ص�y����j�ފ8��y�HK��5+�C����x��R�Z4�l�C@9y������&�q�������
X梫�!��ۨ��S�����y�0�}��*g7-��t�*�J`��?%٭1���Ƕ����e���-^>�!m�]���+�����S�V|�9�F�R;(����Ԇ5��[�����qݤT�V�Tn�zϪw(P��Z�K�`������_��}Z�P�T$!��FS��7*���X��$=�����s�m`!�C�B��N�m��@:&�y��#k1�^3����.�+�ܼ�����{�P�Fڞ-j�OG����3��8��_N���A��F��z��[�]C�Z%�-�!�ġ�a��C���Ɯ�{�z� �G-������T��V[=��e��Ʊ0r�7����Q��"�r��4LC�#s�G�^6��/z�sIU����v��I�Hl�4�Y1��˯5D�v6�M���Ʉ�6����{��\�2�b��Q姺��r�ޘՓv�����Z��TڜGJ�DL�H��A��0k��F�g8��4*���I�^�P��<V2x6�1H���m���2�g�Įj��H�C�:ʿk�nG�K���-�@0h���z��2��&�#���T�]=��z��`�^��Oʵ�lC����`�`�y��̛7Ѷ�$s�Z���8�������(Q���"����ɍ�|���(�
X�����H��Ǡ��n+������7����v���vEl=�ʁ��"`��7��
o:�h엟�;{�7n�#_���X���U���
���i�=����Ä�����r���~�J���u����Խ���hOK;����qy).T4J�g�W�la�Ʊ}Br39�0��b1��0���~�w �O��=4,f�%���cY��/Bt�^�D�f�-	a�nƐ��*ћ�w����&��U��m�tb���v"��_9�c�����V��� ��;���`�-�wZ�e-�]�4=w(7�1j�R��F���x��Uk����4�2Ҭ�sP��R�q����|���2�h���	g+���3���ц�R��u3QX]`|U5� �R��|�WUY ��M��S���8 �X��n$#��pSV�72��`�]���:�j��|��bVm�ܑ֥Sh�rn�g���_�����c=��:#�6vE�SNx���7�\t�b�[���2��>WaD�"���,"	��o��!�O���>�9~�<���&����MFy�g
��_Bc�������~�0���l|�]/Y�f`n=��rL̹J��z�{X1lo�Wu*@�ԣz9D�HhL!�9�]3��_�`���x�>��[dMY�7�a ���h���dh��6WH���,�8)^�=��{T�2��1@��B�L#�A�M�����7�	m�HVJ�~@��O	���������Ey[�iM)��le��z�MLSU�A�=����y0Nվz����Ɖ�X-F����1*V�R*�G�I!_��Q�_Tĉds�w�}��Lb&�}Is0˵|%��ad�T'a��<��'��_ ��������3�62�֋>@ɩ���}������������[��]������9'�GZ@��w��rtjy��`22�<�]�Z3�z�M�'l��m�|�>	>6_U�D-ɥExm��s{w��A[>s�q�,�AVTt�;�C��y�IW	.�J�~?�h\����
�Sa)B�פ��(<���ьA$�\9Ҩ%(�9w��r��T+Ai�(d�Gdz�%~���!Z{wɁI��5B�8���tZ�>�������!�(����#ɿ©k�l��!eJ��/�� [�����L'>���i+���}�b����A�����)��"@.yД	�����f�5k�ٹX�c�<O ��Y�oߝ�a�	S���6�P�ܸgz]*���ހv|YP`Q./��'�=�'�����8�!0q����uz>2�?��ᾫ�I�c�=H�z��g�I.2�.���ll���K��V����yG�N����~��Oi'�<xr����E:������BI�����
ᮅW,x~�{W�:�/��j���#�o���y;tGm��S�k��UH�$�?�#S�\�Mf32�Y���!��g#�*^H�t`:�ѵ\��u���:�C�p�*
���w.���>e$�U������u�2F���Z�Q���Bh�Ƌ���,C�)z@��թ<��䈥��õF
��آ����q���(Kda[���؝���p��-�I�ߩO�6p��;���N�6��J�:
#ܰÅ���Ӝ?`�Yϓ�D��q�Vs0~��p����؃��� 60l���:���',[����>��l�O�2o��~d�kt�d���3$N� "�	���+@ǋ aA�b���af�p. N�ȭ3~��N�]���w�:+Ŷ�a�ݑ��ξE2^�r�~�J�-
���Sc�����Gu����T]�b9|o�t�lB���������k�<�;l�jB5UZ0�v��Vΰ������0=FST���m3�^* 5~X�)8WV��-+�X�ӛ��`\����w����5!6�&����9���\��]�.C��Ĥ�_S9�T�oqQU.�h0����.+�$g��n���E<������=�֒ra��ۜ��@�P����V�+�UΏ�"� ��t���x�`m�b�Pf�� :^��e�N�y�D�B'�k1/Z4"%Y{rg�?��O�h��ǡKyXJ��u��E�*XM��8X��?.ɺ
�RG|
X�0o��l��L���Z�a E\rqh"?�I\�r���"��O\��#��u����F��)��B3��zU
kA��2d��v�^{����>�P-����3�KB���|7�W�%���O
��S��
	��c��xd��U��GT��O�����䂦��X.	Eͯ�$��%!3���޵�<�1S�ۺ!�=�ø����Hep�4�����(�*A���i��4t���n��2�A��r����8���0.I��B�o��U��1U/�ze��q*�e� b��$�@?N�^�}�U���l�]�E~4y��g�~��:@��#1������V*�Z�d�H1k��z���4\�:z�G�h�c&%
j/"���w��A$*�'�$@�@n�%b
�&�8�ʩ�W[(�E����Δ��U�ѧߩ�%�����P�9X	�a�S�Ұ��W�ݳ�[�,g��R(-߂�+�A.�.�Z>��>��7K�㘃��7���2��wU�@#�J�T���t�Ȉ�/U�6�(��m����Ye�(����N�t�-���֧+��IO�^d
7��d9�,7�Z�����E�lv��x��={���N��6��J��n����ֱj�ZU��{�c'«o;�I�L����5`y�B	��	!hM��|�+~�
r�U�@x��j"��+�Um��6������H<D	D~��E�Fb0�A�A=��,Mk�Y<�.��>�-Q��6"/M�Ӑ�\�d�hFb�_�_/P���q�+N�s@�2�5�Z�АP>0����+ٜ�d��� ���=6�r�T�A��MR~���G����K�!ߌa��2#O�6�Q�*"�I$ӌ
�iw�%z��U��q)�w��g�E�,�.���	u��f#@��7x!L�,���Ubl�9�A��2�y�Q��TX�J�p6��.Sv1� 鸝�j��?��n�ߨ�:^�G1�ۦ~m{���L^D���IޟI��7�(]���M��ѓa$�j��/:h�m������+P���p��`�s�����
�h�勇z�|o���
)K��,J�9��A��H8�5L��d�j*�L� ���ՉEc��r�ַ��;�<������@��`h�A=2 w�Q��a�_��Q���J�J�6�e�ߌ!잾���8f��ɘ��!��>�P%qx�xYO
�鳵N���5�C�c��L�).�t���o�>i��s*)2IT�Rٗ�Ņ,�\�J{����Łp[���ٟ�7�[=��]�#���-X��(ѓ:�k��ގ� 2�)ߔrl9J�u.z#��nn�<	w@�W�@:D��CHZqmZ�f���_.l7�B��0�'S�t��]C��x;�n�����e��� ""��؛M��5�I+f��s��ZTd�)��D (�R_�)�SC�Au���Ɲhwfp�"��ӜM���E��:º9)RO#!��˞$1P^��(�j��s<��4��A/^�Vn���߆S���B�ET�#�TM��_�xxvk��r0s�5�+-L���)�(+=&	�a-��Osd��R�5�E2V/���9q���������!eϽ"+W����:^F8��;B�ꕡxu���+�9I�G<fl={�H��MZo��U�by3�6`�	R��r(��W;
�^� ���ڍ"�&q�D�S�?6���c����� v�A��tx�d����z9�KE����\n?�\6��/�_��U�#]�R�(0��qv,��piL)��X�-�pt�S��@ +�DTy\���0l+����� �f��	f��q�f��b^��l��x��腹0��� ~=vX��� � �����U�;��G#�������;=�|צ��e�
ht�1��U.lu��G@jm�ر.����'�Kk��_�D���K&��Lq�e!-Hw���Z�%`3���M����e��%��ƶJ�nb�O=��J ��>�;�A�Z���c��(�z(�OA_��TW*�&4q�Cw`��P��W������y��P`���;�F7��l����_�������^��h
b�.ϔa�C�oI3:/lC��_���#+�����#�O'��L�ؙ�$("��Ѭ���/�qdo�]��uR�X�H�űq��b��۽J� �P��l0�qM���h��[�&����@&M� {&p�~�3-���Q��JU��_|�%������q����l�Ur�܆�0i��������+b'2�ߓ?�PaȖ�n��b�é$�m
�6��oO�&�j��N�,�s��A��g�&Ƽ���ྴ\uG�CY�9ri��y������d���:ڐ�	*�1
9��gBg�fy���������R~Z@_�[\}Z"��q-A���*h�j�-k�&�i���F��F����:Y �I7�W`��Q(F���Š�,�J��"��;COpDW��ŨZr�d��z�2������hw4l�7)���}f��V7�� ��y (�ah�J�R��7ޜ���}T1|�ѭ'+O�3k�e��v���<�;���Gݭ�.g�������,��=�"0F�p��(�U����ƙ��Y�m��[y���aLp�5}�z�* �������N���)~nZ�$��/͍�8�r����\���G�nE*1���u��I�a�-�O�U9����g4����<��$����/�����Ya�Ht�#1�^*�)
EyE�6V'�e�Q�dx,�g{��߈I��A��kG`OSF�������������"��5 �1R�r}ф��	�:J���Bo�kt�t�M�ͣ��d�4���S��=F.�*Z��L���腯���RijX�C*��N�зe�6�'T:��+V%$�&}lH��d�(8�.��@��:�Ws��Ӗ[#��aك~9	�g���-6S?��X}���6���3��9�Su�����9��iOP]���o�$F>+��y�)�;��ӶNA�7�@7��2.�:,-
�ٴ��#N�x���#���P��y�n�ۦy���[�����m����Z�{����xm+b�@$��D��R�z4�
� |D��5�6���s~(W�������ǭ���P��?�]y-�M�8��[d�C�?���?g�� �U���#�̤t�2����(���b(��RUb2����� Yp/��I%qM���Iݰ�����<�ʤ���/�+�sz2E���s��p�G�I��H=��Fg��,X�����t�_CP�T�@G�݁��?�Lދ5!kCx��)��C�)R��d@�|oK�����"�����J���u�ѷz��#�2�Ja�c�Gv���e<���k��of#�b��#}7���XO�T�����W%�R�������c�+�#4�mW_OC���F��`;��<q1�XF8����8D�z+��;8������:i�_����+�?<�
{�����U�V3��O�`�tu�R���j�{a�?����4�p�װX�u�1��Z�EHH�Y�K���'�u���f�^h?`�s~��Lô� l�H�Ֆ-��6��{	����DA���P�̱J��z����G2�=�&'��+��n?Nqk�Tʢoy3�D� x��SA(����:׍�O���S��E&;�9B5k�@��^#+����UA�]Q�cw�r<85����Y��)g���S7�1���(&�UH�^������z��I>-�$F)���*Ңt^�u<DI@ �y]�	q�Q�0�;{i����*�H�R�$�6b�������rÍ+�Ug���e=��,��0N�������[�#����@�MA�0�x"�,GY6��)^9��욙�yv��zp�ÔT2�P\j���t� s6T��6T3Dy��� ����c���<�A<"Z����f�{6<��ɀ��.Q�f�q��M�k��iE�'��(�)�_� �њڃRR��f�������Э�%��@yC예�=��4�4������i�U���A���eP��� �o�榀<1X�tiSI/˔s���׳F��%ҽ���}i�K���N���3C���xm��-�X�E�7��z�N��[��t����-��;&=�� j�4�ɺ&�������s7��1=�3�H:��L1f��pİi��l�`�I:p��BT)�����[?�]��-@�� p`�~����*�끬���z��n�WjI���v� A��0	cR��V���SB�X�e|Q<N��zl����b���&'�l��Bj�|�x�� ǨHOTL{SDpX� m�|Uk�=w�6#�S�{@��>���~��na�4$�(��ֶ���d�7�d�Q}��Č���a�՗a&�]Q�z ߂cTO�{3���9��`�}):P��7���{~v����K	~�2*VB�P}4?O0��Kw��wGt��m������ʌ���r������T8�pyu��%�Y4?Or7���Zgl`�D�B��@�x��&�^�E�?)y��	���E�6�6�z$Lȧ�?'�or�����V�eX��)>-�w%�G���t�eL�M o6��=�e��t2gM�V����%��i�A����\��Kd�*d���]����z�9�������.�oCό0֤�Yn�3H����{�+^m2��������s�te��Rҭ��[�SI{7��J�x"F���9PTo��	5��m����KT9O}8��ȓ���Q���tD�W��+�t"�o-w�JM5(%;GT�X"��-<�)h����%�k�~�n�.��z*}�l�/�O�7��d������M���m��Ǿ_�C E��͎+F�=l.B�D����X��b1�����IQґ�;���Q�L��<�`�!�_�?�Z���.r:ʏ]q��T�Lpb�|�bG}�о�?TQ����J��6S�IjG|����%U��/�2%*����9�;|S�m@YG�`�7я/��O�)�gZt�����	c�9���.3[T�7(_V��
���)	:��xSS�4�*���W������kV!������]�5��-���jUn_ϭ���7>
3ȇ-Q��4]N���B`��#�ǆ���%q�6��bQt��' �˦̢A�0�pn�~�j���CF1���coT�d�X�F�	@hCU��a߃h��g{�g=
���ڏ�r�����}� %����rL�����˭�o�9)� v������OTkd�����R�>jrC�L�95FsI�_�&1�~x`d���V����o���sF�xvv���B�}`4�B�8C��j=�/��� W_��!�B�!ǧҦՏ�Ӣ�.r���\ri�DrKϺ�Ι��-��&�r5��Ag�h{A,���8^' I���L����'us4�|��hE��̄}fy� O�e��bQ��}��&�\=Nz��iC�>�R����/GVlX�(*v����:���.Ub�G��K.���73�顙,��I�LC4j۽�՜�{ڷ�b!���k�%MW��Q���$'Z[���|֦�@�r��e�U���}��V��a3VK<$��/3�ܾ���b¼��M|�j��I�2�R�s��7�$����J�!����4k�K0�VHqӭ��h;2:l4�.lF�B�jnx'K�Fъt�(Q�l�7����IW&'#I�R��s���:�bC���9�h��Ģ�g�p��@����N��E�^�Ǫ˂^�N�$�W'���@&�ʗb״�����2t܌{� Iջ�1M@~�����b��	��a�lxM���2�k=O9:�P�(����A%=g���9�6��y�N���X_a�b�����^/�$T]<x�bHT��-l��j����a��1䷀�`̡"c�}|ˆ�����t�8�q
�*]���/�B�=��ܖ��6D��h3�Q��y����9��9:��9.cq� OZ��ĩ!l#�xME
"�Dj�C�Mn�g�?�i�Yb���\K+i�r�Y��YCREJ|���B����Yx[n_�~���k�8&Z���Q�k���*ϝ���f��#,Z�t�a4\�IV:ʞa�bV�+)|1i�:x9��G�<<άv��p��G�S0�Z9i-�)4��*
����mb�͹}�'œx�}eGIy/W�t$�u����_���Ͳ�)
���+,	L��/��(��Hg�s��Lnt�/^��VCﲐD �ļ�$����A�l_�@G����ݿ�s��y��wT��AS���վ�����?�l�6��N'UV��3������u�����3L���;0���v�^H�GϽn�U��_v�	��K����.���k�}��ܵuw`ct}��=�V?��!�5M=�e��J�6� ��#��<��0T�`�j��,���d���#�C�]�w�/�n��� �yX���f�����x۩9 �T�_ޘ�����NY7;�`y���d�T�K=�C��2z�)���&���R��>����:�Z{���]��S�\����
���{�~Q�Y�6&!��}V��	�:�3�$��0�X��@������@rH5���_�oL��$�5�(ۑ�K�����KK��]� �e�]�6�e��A��M���=.{iҁЙ2*wb�v�El����z_�$�{��6kX�lC{�l��s[<�`����fQ#w�e�˺�>����*�k{�w^�1rEe�d �����6�]�tF�n-%0�iP����O�Qp�-5�QC�c�C�V��8�:�
]zAz��Ԇֻo�1�$!�k��W���,��p�4c�|G��Nt�CMj�8>	�ٌF��snY����UJ�
xe2��`�;>�$fL�{�O^suH���Ձ9b8��|T�v��Wz8�Q��D��/�I.fɴ܋? �$�%�]iR�3�f	�B�W;Ȭ� �v̬�jx
�/��d���i�}>��x+ � ���(�6�`�(�٦7{�����y�����i"�A[�X���@@���`�7�Nw)��Xx�rF��';VE�@��D�~�W�+?$Y�4Kæ��05��Y�9b`|���`�?��d��8�r�=�'5��5���;
4ڼx]ũh��g9i�()hf�4���3-\e��J�k�����D�
��)8�Čr��7�m��h�/v��hI=C�;�|�WD'����/Q~Z�{�ܯ)p���ͻ}��E.e��J�H���*�����U���`�#��܂=��cN�9��Nu��6E��v��N�� �b-���2m�/? O@@��ew�� ��d�X����g�dD��[�P�arbz� �r�%ώh�o�q�i�V���!��	i)7?����2��x��+\Z^��d��%4@@*����m�Dp�8���v���0�T`�6�%�pp���. �\�o2�l���T�.���]���W�VP.c�9�`��]
�VKj���CM5{��~��.�����|,Ĺ2$�!�m�+�El��4ee.(�:E�l�!�w�,�I����<}zT�׊���<e4�8>��P*)'����^��M੹��S�c�lo�?kO&�6����:b���'�mE�Un��u�*�dWHM�O��չ:y%W�� ��hgEyP���ߖR2f���u��Er���)�^+g̝�"����8]DA	�(�#Gf�0�����fR��[ydz�㕫��:\#�=c�,�]����㤱w�uA:���D��h��0���P�5=�bJ�VE*_m�V�\P�]a
$c�M8�hwP��.������O�.�śOӛ������g0��	J�%���d��O�~XYI!>]�A��� C����{b>~��wE����;ʃԮP�[Re�Y�U�`L��k�LU�*��G�^}�oƯ;�.��T{����xG󖃟*���w�l���B�J��/��:�����S���9QJMtn�X�>o 	w��6Z�Xf . ��w�4I���	:h�+H�c�J�>�� I�jC��]�2�������O�a1)�o�/�Ɏ��ŨD�"90��L��������F��F�Ǚc7�r�&ZўO��+e���F�6֨���x=4x����1P��i��y�eU*֌�"��>��K��l>�Hn�G��^�Bn�n(\I!z��4�/Zؾ����xj��;O��`P���=��\�������bL�$�f��앓@n�[�`I;��L�����S�dhD���j�f�Mw�e��r	�%>�g��p���=�Ƶ$=X�-l���w�P�i#ܮ⵿`_j�ݕѳ�$�E��!��4�ݒ��}p�X"��ݔ]*ͣ��@`�ç��O[W��}�s(��j�H~�}iEꂆ�4�s��$�|rv�.F��g��x��t]�x��e����ҷ�ۙ�ժ���8� ������2F�W��F��T��}���c]ߦ�Y�ƚeU�CQ�z&�f��Vm�c���?O,B��iJ��+x���2"n��]��*yv��+e�a�N��Ć�� w*x�ϦOǻVʦH���A�ev�S�4�b*ɰi˺��eQ!CجΑKÜ��}�b��$3I��R�W&��LY���`=����6���Դ=�^R7��g^�B�0�դކl� ��q��1���>�ϑ�$���+¢�jT%��V#�W~�؝������dM�y��.���॥?֡�����f��i�
y�.��J<c2u\���G��9	��<F�lu_ɫM
��SG�~��H��]md�k��&'�[��̾;]~�hO�[ɹѤ�j%Y���r��U��ۙ �E�0��~}Nz����;��$���r)=���a��r�ܚ��]zf���~��?��!�~�bF����ĵΠg:u>2��&��=-�a�5d�/�������5�H�i�!"w�T���`�Ȭ�4�a�M�l�����4S=��K�d�l�}�*�j[�D���nN������DW�!iݝ��f(�N�eI�!uA0�KY����NJ�6�?�Yy"� ��f�/9�C��3C���FVT�� z�F	��qM�]����)V��_|��#�M )8?[K�F��;�$8^	�5�*�J��"p:�vj���ն����D%�+H�l�����o AWT�9ipVǋ��a�z�| =5b��?0��]��ɶQ���/Cj�+��\�^�,�-���0,a�a�����p���<��8~DP��"]��UbX�ͻ	c�wu๷��1�L�%$ p�18P�G$� o�8������G�.�)�(��ew$B���x�J��G⭮�Oä�pM��m���Я�����ˎF�3�6��~�o�,	S7J��0T�� �Ƕ����7���XO���?E%�����G7P���_�s���� ���7�eh`��-����Zo�D�N�N�oL hɊ���W
�=�9A�C2;t@/�)���_�S��T�J�@��*Z�q��H	M_�Yζ2n�\�b=,$$����x8l����"(�P5;�����)xk��~{�ג��,�e�8^��j���TE�ƴ��g���6��o����'unY��t��s�����"�l��V��u��-M��Γ߅"�Ң�C.���i��餟/=v��oZ����a콷�VQdaSI�9~�I8JG�з���U�k^#�Oh�����E��1֟���Y�(5ZF��I�}@̭r����.eu��H	)i(J�,� ~%]�y��.@ʬ��K7 n�W�3�.�L%t[��]E~��@��pj�ޫ��B�J��ή���j�m�Pݕ`F��Lp�1%us�ۋ9�bh%pN0�Na4�,���S��gc�����6;d�'�=���8����S��1��)��\_���p��-&>��	R~Q^d�]�����%~�犔-���ɨ�e	�}=�s]��^ �@_l�C��#	'(��4G�Ϡ���r�Dk�\�F�I 8<�	�0�h���S!6�/�D:�il��j��� Kau�5�q�U4-�ʻ�)½���!�kn;���[��A�JQ0�>�5�v�ɼG�6O��qe����C��@يQ�^VV�{���܀��������e�>�+�Ҡt�J���������Bשt//�����K�(1����m�_�]���dY�`�r�$&ĥb[����|���9;��w�flŹ�K;��M����0��k)^��wJ�cb:��Rߑp�Rդ8�m�r�*��k ����8R1ο?)r�,�.�Ŝ!�k���x`j�z�K��4��]��f0aB��_������=�\:o��"ccm�ns�̞#V��,�G(��+��t����&�2kh\�'YVХ��XêVu����X�;4���n�=#0���C.�E�r�>Y����_%�m҂@�m��,��?�]ߤ[p�b���H�m�e��g��2S��hE(r,��v�;��$��`��N^��
2SH�m6'R���"�P��}^���&�`	\&��v��r��u���$!���Na���'��8�YB���#q�Ag*�������P��`�Ǟ����w���A��O���Q!�q��K�p�$lZ��E�n�n��yr#���eXͥ��(�3r�~��r��!G����r5�( ¯���G�cI8r��ZX��M1Ǯq N�T�ˉ�t�a(�����	W���Yr����H(T���Jf/S�	���W�w��V�}h`�^v.ś�*�U: �'jh���@>�����:4�b�e0`ϯ���!O���6.��rb�*�Xn���k	-d���qA�P�fS7��O5r-�ї�������.e5����x�	�\)��i�E��KB�W��#�R>��Kiⵆ����C%]�=���/	�X�lD���:[�n�4��q�%א�ۘ�{��%},��EQz,�W�w�����(�����h^�;��	p5�@f�� �vJ���ٝ�>Ygͻ6�s��KjC[r�ר�}ї�w�����$���2����H=e���D�+��i����J��Aخv�c�<������4P����;hx��dH���pP�Z���\Z~�Y��	n�.T�eM��|Nۇ�b|��wm�Ӡ%X8}0 Q	#�^�������ґɥ))3p�T��̼f�&��X�FԨDѯ��O�� �Ί�x�W=�r�����)<6y�@b��Qm�!�k�����2��i��4��`�nWw^8!��T�>�ǄO+��aHE߇0�07��r�脇t������P���<�I��Y����$TQH-j0Ih��e^]fP:8�%�ڋ�ב��nn��T`�m_Q��OB�����;�rj@C&rLVV�v�8�Y�}T�G6Qp�oV1���}�9�X^UM�rى�ek�U���B�@9/,`�e��l+�^��ݝ�>���Ƴ�i&V���ͯmg��Dd��2�86�W�Mg
+l)�R��p����	�֖�14�2���%�K_cR��ř��!cV��_��'��}B�W(��jA)slRk׋:Nz��}�ʧZ��x6���O\
[*i�Vʛ�X����.$�`5�g�r�eS�]�F$vw�/:|����$.m�>g�F��x��=lC����1��l���X�� A������%�SkJ�C\�mM��2ñZ#g��x�?��Ib��_�7�yx��|�?��+_#����Q͙�;�%��oGG�����IA~�3��'�M�ቜ&$zҔ	�j���M�̚�S6��f9�b][��w�q�Ai�����v`�	^�br�_�0U���M�e����:�x���,cO�!�6{��s� ��w��A^_� ��e� ;7@�͠��jz��8�K=Z�?r���?ޓz�o�P��[��=M�gm?�8���z9��Jr��fٛC��u�������٫ځJ5��T��5w�ԗ��,�&��3���,��_y >)���<�V�E9{,ꖒB(�jp��WӼ[e�e�ۑ�y�%�*
��4Z�/�/?��S��S�.��2�K
�<҄�
_�E�фnQ�Ge*�Q&J0��rЃ^��[�>0m^*!�>������V��u&ﻀ��A�cG0IXy�1�ֈA"Z���5�_?; �+M�&cz!�޼Ԝ؏b��^
*�7�Ukad�سʠ���11��g :y������"��U׃�}!	n�sc{p)��j�X�Bq��h"{P�/YY���x�B����
��y��=N��s`�X'&̇����y�7�����j�bz0���^0�:U&�,�-sBS��s��<N#��|���Z�@ ��#�(�±q�Wk,>?CE��f
��?b�x�rt6�_�;zpP]I��P3�|Xe%z�c}n�����/���`��Ֆ����h���z��$ʸ��7����q�j�C�L��4���$���< ]���c>Zx-��O+�q�
�/3%��A��RZf@�@�nA�U;%a���]2�!�$��u�>/#��.Qs�Px+����M���G���b���N�ݎA�h�a���P��1��Fg�X�������c��
�/�ؖ$���=i�a��� ���
}������T%�]y���(�G��1K}�<�8��klB[�>GE=i�e@�
�)$�q�53��q�Ӆ,=N��.H�Q��8�K٫bӈ�c��Y_Ͽ?t����0�����E�_?ߥ~[�����B[������Ml$�y�y�ec��61ϸ��iJ�b�$��������C�!�H�ɯ�%;:�#r�ƽ��a�<�lPW�GW���u���� �J�.*����-6hVl�O������ao��|gF{�o�Z�8*�sQ�t���D�JiʪB�5�WwF�����C�fyZ���,��d�}m����2G�p�y�V*�B��[��$H�)13��9X�ao�=�+GrfN�QjB�s�0�찕��_��̬t���m=|�x����!�nH�G~�$(�ڸ�,��;�5c'�;�_�;b�q˭o?�Ѣ?LJ('B�>�z%�If�޲�G@��}-��|A�ڋ��d���Ȣ�vbv7�Z���0�����f�5�����1��Ӛ��@C	vX�!�U�#y�]+
��*��o���"����@���M�I�vݝsy��V,� sD#e��&�@��L�Я<�UE{� �o�_N�-��+5kT`�r�3�|��B�et����d��NXp	G\@�\)��u2Q/��A��ܨ������y��&�9ۭ�>��Kq٧h���R�[Д2!�gz"���̟��]+�s��fи�ѭ���,�3�������F�Ӄ��b�>:���x�'{aP�8@t�Iʚ�e��YWT�T `�͠����������D��"�T�Kkj9�7�ss�y�(��x�[j5��E��4���q.r��V:M�$�UQm�]o�	Xvp-b��x>�ۼ�� Mj��
����aT+�����+M,pyHi�F3O�]� !����, �%%�q�!\m��11T.��K0���9;�� �[��M�ʸ`�NиMғ���5/N�Ա(]��g��m`B�hfg�cJ`D�4F��u���X����*�PN�;w��t�Pp	G��@�3c�l>���g��W}V�Nxq��r��(�-�pR���dv�5�;j�u�U�U��I��w���kpo��$M�߾�~"6��s��<ȉ�<N*_/ N@�y/�fV��>n�x��r�AU�o���n6��D/iS;UC>�)��E킒<�9a{'3���y/���z=���=��$�2�����LK%����nd+���_F�1�	3Ć�K$�!A�1<�)@KC�72/���[ߕ��m�'l��yc̝��tQd��~Y�`dp8$ߢ�jkr��}�>�#�\��4���Z���swk�d'���O���&���b�7�e#N�u`H�[Ӯ5��vjӆ ���M�+U�>�m�?����T�nT Ij3���W���T;w�w�)P���f�w���O�Cc6�6��[Mj�	�'��D�k��\�2� �)Z).V��tHHV��8��t;���7�X��T��_#�"�:��J�i�Yb��FøV���R����56�#��Xpz��^��F*,G,�;��Ўi9�����4GA7�~���oosZ �G�Z������]���� ���z��Z�K!� ���l�����6KF�ԯ�j(;"��n|�=��r�@�N�{'�C`�LP��D�ϋE��Ʋ�U���}���d:���gWI���z��W�s˕~�*"]5�?�����XAw�lK�>�`b$9�o!#�3#E`��<2eq�0F|`8�Ebb3U�������g��Ym�����|�H��鸒ڃYg@��+Bk�h�|�1;=�x��犯�J�K��$��1��U�A�^U��#S�p�Ry�1�2H��jY���/��%�h�W�r���A�t���A0�A�7�H����+eOe�{�ӈ͗�g	���@E�0�>?�����G ��Yoơ�I�]j��X�Rn�ۭ(��ar눆o@f��y�-�D%O�����!���;Q\#�r��UTG���QiJ� �N���Ca;�k巁�3k%[��T�6����tm�zmrO���fӴ}��K5�f�չWf������#�B����V��xT�7�p��ʤi-&�q���]j�����`�]	.j�;�y1��.�E�����1mOt����>�!u(�_��4`�9�Դ"��n�i+ ����{��b�Ug�efL_�4,�1�G_��u#���Jk����zI%<NN��������Lsp��(��eREۺ���u�՞;}�ȱ1����%��Å˟��'�}�K�����=~����d���zp�n6/{�Y�U�X�Vyo�T]y�Aˋ�Y��.,�}p���DrlB����|��R��@�Ņ��w��#�O}3-�@	��RRߤ���q �N�/�,v�58���b"�fS�����I1�u�YY�ȣ* 1���E�}v�8Y9��;�~Z�|`4چA����b�yB�7��@%��i�5*��	�[��|��j�x��Ǩ�$1�\�)>�( ��fr0\b�x��H�+�����^!�-"���[9����X�ۂ4�"��w
�o	�ǿB��rVW�vO�#��ݓ:S�87�E�_�icFp�_������:4���"!^m�W�$��Q��T�ܙ	�� Ǔ�T݅NpIסg��(74�M�J�(Bo9#5�Ã<�9O�g�>K��R��!�}=ۢaV���V�f�H�P�ST���j���ƕ��9�~m��?�q�t������(�;�^�,���jd��9˿�t��w�XU�,Ҿ(���P�8�X5N��^ݍ��b�����?�b��N�/��r�g�u��;_�Y(���shZL�y��_��*'�+�s�K�O�o
�B��(y�(��?�6{��3z��HU�T�� ���CI���)_�X��%�iO�8�c>�x8ї�?���Fl�<���*�m��+>��@&Bv_W�-{��Ӥ�Q�����(nu8�G��ѻ�Wa�=��kyۉW�7�5�1�0Se�	�����e�Efk��]�,�:�u˸���aZ<�U;���S��"~�U%(�b�9���
P���a�@��#M�kυ�2v�����G.����f�|��4�%d �῱��+F�ś�&ӪY$�A�L��`�(=���Q�&���'�O��6Izr��MC.�v��*ϝN@����80���A�1m4�>�?�!\���;��%ᐯ�/	�C:�x"�S*��4���jW����e�������}O���\n�l9�A.���u`r!����&��O�Õ�.�o��G��k7����u��#A�9B̠M��Q�P��a���w�H���rs�m�?
	�u{��������^%�h�-��]�,8�ЌZ��lv�����|'�N�W�@����{o?tՄ�x�o��u��������}��Ɔ���)	i��!�|���ρ���Q�;��=�;�I=L4����;W�oxʭ�lp�#A&��l��fh�W�
�f7"�]@�������U�M�f�J�e�7Ӂ�Z�O2"��*|�O��-�UpE�M�Smde�x��>ҙ�I���*�&2��)#�=2ÿ�J� i^1�H���ӕ`�p5Y�z:Bӫ�^zyE���w��/�[�[�K�|�B���_�&6�ڵ�Ak�e2�<�!�s���c�/ʊ��a��/A���
��Q�O�Q�����jn�jtNf���q'%�ʔ�9���H�cVÀL=W	��i��Wa�?�9�_�&a��?��P�W��5�{N��M�@�'�P�'��2.y''�wؤ9�k�v4�i�]VUGq����θ� �� Q��k~U���o�8`��.��J+�r�"�4~"p  ߂���x�Y�4}�H����=?�LA�_>��'砂��`}�/�1�L��ђ�5ˎ�/b��#9�F�Rd��By�Н�墡�����S�9�;eilE4��}��� |sX[|w�&��u���ƛl��rڥh�+�2~�Xɘ��Ș�iq�t�C��2X=�k�2���)�N��$Q@JxY6h������<zg~atOC���M�]K�g5 �b�Y��j�u�Z���s�2��=�{��&�2�
�.�<�w��7��^�Ԋ
��<��M�	I{"p���x����;�bj��� 	��o�0m��= 21��( ·�K�N�`��z�P��[K�}�?�E�N/�.m�lj���g���� �.�r�@�%����Z�[�̞q�u�R��9s�ܦ��=
ז��O_]�-�8��`�e�S���.`wI���Q}�����͋!v�c�16v7�NO���(�G����$�k��QP���G��w^�#�1,v�L��T���i���0-����U�Dq]c@���­=���B��x%���R'S!9��=֛Tv�g�! ܩ~ƿ�a'�����CYCw�z�ǻ���w/�����5�]�ZB �|h`���r��-lS1�L\�%���]�B��*��"��^���u����Z�z��Z,����|$!�:'C�p ���T�+��B<W[ �:C�gWGf ����g{�-]$TYZ[�G�.��2�)�@��,Tcw���)�{�w��1����(������GU� �X��r�a��R����f�KI9BJC!]c���X�.�y�d��}N�0��"s��bD]������1Cj�Z?m$}�A�"l��O"R��0c�T,�m넘���[�0��'�+{H�x���������'�NPdA���W�I�G2�8CfyK�Q?y���:e��z�N�����Q,px�S�O��b����5c1��x,�ʑ�~����6��RP��W��f��<m 2}lb+H(��f��&�>I��Ϧ�K��+�0:�d�tc�̉�U�
�Ů�Ǳ���I����a	Bgl�u�P�!5I��5�V����-���`���NˋV�?a�Dl����ܬd87�3�uo��,e�f^����8�R��v���mo���V7:��y���sF*��&W�:ફj��Ҧ��<� ak���!��N����1���q�j?��܎ S�yZo;��0���C���#5 �ĸ�1�M��23R	�r	<g~��=�B��#OG��y����Ѻ��Y�ȁ�.}m���M?i{gmR��qNf�PXtā�7$��N���C��Ĩ�z	����^ڀ�f]g�0o��h��H���2���XP�-�֨(�KH���|y��(~�v"TY�h���z�%An�N���st�rG6�| �����y���!��x�@LQ$&_��5�F���k��C�d=e���6_[�7z�/vˋ�U%.��{{��p.Ե�P}����-o#�^��ɝ�l�]��(c��Cꉍn��u7 � �Ǌl�~0�J�\�uqJ�Tb֭���Ɇ�-?:)���a(0�E��b%(	�|��c�.o�d{cj��ZO���?�υ�p*�KOrt��z<���;i�Z�`��	�JZ�V�m�ȍ�||�VnO��Ϣ՘��VA���H�؂MF�&@�RLo����O�;C��Z$>#�g��ڬ~����g��]�Jy����w�F���pm!��k��\��y|W���U�f(���#Z�*�m��^Һ��T@^�i�$��h�{��MA�'Y��*����W�n�P/�N�f���um�8��8�O������]�1�0:FpX�ue�N\	�U�z=��4������`�L�z�>?�jA���jGxG�y_��mV"CW�܋��Mߡ�ޖ�X�� YtG��4vMK�E7 VY�dʆ��1`cxC�	m���O	�ZuV{���TiL(H'�_U�0�g	;o&TgcVO�.�=�G�����1c�L�IT�I���4ހ�XB�-ҹMU��H�0"���CX2�F�4Dthf�^K�n�PO}#�7�dsv���.��^�$�	��W`r��by�P�F�UF���u�ԫ^zkf:b|�L:ҫ������f����^��T�����\\�%��"L�𱿠cW)�[ǔ��q��*:��1�{�#����:�P-!�di�wp�aa��N�p��0
q��rznw��i��wz�������1��5ϧޅ�;-����x���_m��|$�:�Bv���=F9c��^�⓬{m�/��I���g���(��� ��!_@��vaԟ&�կ"�ٺ�ro��<PE�ڸ�󜥼�UVns���W}�Q�}��%`�I$�vp�����軄���ʏ�!�F7�hi�h/�l�
bQ��±Eg�h*�U���te�X�5�)�����%U�ʘ.����5���lxbe��F���1L��j�Ў�io���$$�J�Hk^,;Zf�pEoz�fkF]B�'VfXؼ��3�Ң�G����.8����YՐ��}�Q��i�ϰںy���4����HSufs��OH�q��s;�7��A,����7up^ڱ�1O8�Ik�YOU߇��L�k)���ɤτ� �s�"L�H}Uѿ�0��Ύ��O�>y��X��09�'��j�����Z���'Fr^W
���5h��dۥ��KW�H#ƀL�yJ�2
�K� ��>'L�
�s�fw+���M� �ᝄ�=���NT����a�]O���;�����ʿI���C4��ej(Ki�k�B�Y�_pb(p	��uI�c�t{��,>�$y�y�P���q8YSB���.%e���X,��-a���Vc��(x)P6D�����p�R4>\��Σ_%�i�u?����K���E�˿�Pg5��V�M��]����b�L]!�]&Թ��i_�IF�fGPl��͂ �[�ثv�9w}�5��v�l@?�t0DT:*o���I)O��޲o���#�q�����Z����v?'.���лe�Um�����G�ȳ�)�[�C	 b-(�^�P3���7�\R=KGd�)�S�`GU�h��^i�<#Z����D1���˳�AS�c�����1,-�W�ˎ�Iެ���޳S�g�N�y�{0t]ɼ���E�t��C(V
��|�/h� T��?�ټx[B��𫂛A���4���p{�č��fe!_����ֱƖ�,��|�����ݥW##�$w���ܛ��s�G3I�
��,�>��R�S��'�s�1O`Yph�w�1?�+�3^A!����MO�D��o�;Pv��щ�`�F�B�
��S5��������I��)Z����[�g�+L����x�*Y3kM2$
��i����:s-�����Q5��|
+�;��l�s)�E�-l��.�?��^4�����3�O��>خ�<��,0
��NS~V+�<Q��?6�"���e�:$��$.L�r�JS���W{��L�k1{�p�4�����p�Σ!�*F��o#R)�o�J��뮡�%�/�Z2e~�:�au|{�����j�6]Ξ6�<�>E�~�[���ږ~�G7iY�	rCj^�㘽	9���^��[0��bC�T\"MXo�:m��9H��ͼv��u�
(�u�� 4#����HO]���V.�������^�}Np|��;�!�)H�V.E5-B�Z���Cdj#3�{'9���sy�)s]�X���LL����6���ղ�&d>冔���~��sD6C�.k������df5��k��ձ���1N��RSh5��{l"��ݺ�j�O�n�s+<\�S����3�VKZ�VEF�z��%���e����:�4�L������t��� ����g�I�G��^�PaQ���q�ȭn�IQTet�(�������C�dSf�:���j"���z*��Z�����ƺ2+N-�U���w�u�,�0��8�ӣ�
�}EqUd�E&�O?����J��.�|���9NfY��\<�y��%�)M�J�=��h� ���2�;]�,H�ظy� ór�K�^�����!g����Xl&9�@�'��\+ DLa���Ş��tu"�yB�����B'�'�6T���U�XzH�m� ��=!��+&tݻ���������g�sV�T�������Xr�M���%|��#�Y���p�l��rq��f_	��6���v���i�H)0(Ĭ����#��Kf�|gŁd�?kĴ����3�(�uFwAe6����W��cKz����NCn��߬�-��R��sH^w���J�x3�y��`��Q��(��Ke�U��e�ӷR��iC냒����_��x�P%�Y.��U��4��%�'�;��qgNE�$��P@C���MfҬA�Uk�8��c$�1$�d�S4�pa�1Yu���z�k�t��b�11т@G��Ѷ&{ǗceGOۓ�wT�3e^���h�?�j�e��I�,�5��م��;��q�/0�N^e2"�q�+E�Z6X�P�Gu�͔�����`V8��Ec%��˘���d|���gb��B��h�Kz*Pt��A�_�z1��n��?��)�����߃�2��oz��l̎DQV�]16��}��Jȴg�6n<n��|>��5H۩џ�����)I��Y��V��F
�1�Z���_��GB��&v|�U<y>�Y]K{|�
w��X�nٲ6�\yL�O��>C^9��#�ł� �}BbC�7ڔ��M��f�<�Y��wi�R�l��\�vȥ`8R������]��υ�'�c2%��wv�7GZ�L:�GM�����������X�:-�����Ж���:��I4��HB}���&s}d��^}����i;2B����ۗҒ+������N���C�0CE��� �M�bV�⥯tEZ�5$'<ȧj+WD��~��yj؈$v-*u���?�3e�X>�ė�B�R�����@�شV��2��@ V�[>��
=j���H��aR�2S�l��C|��M��%/���D��T��m=L���A#L�s�	�
a����"G~ �a��xϔ�6��n���F�;ԁT���1!P�L���7�R_,<���)�c��:��~6��4�g�y�EG�2�f��ij��C�P0�1��������B����n��F�+ͷ�X�I���)�ߐ���+g�u��a��gug��g�3F���1"��&[��8��(\�Y�\Ǖ�n��ML�ܮhS�9�ӯ�O��
>d-�-�!?0dߨ>�`w�F,#�%�==�}2�� h�&��`�P�g7��&]_r��k������}���("��&#gQ�WH��q�U���mQ�O�rvA��_Z(���}|T����-}�=r]ډ5��r���6���G��#��KHz7L^�쮳�!#I�0����K��$��7�B^�]�S����VkE�\-[��s�S8�������b���f�?�3$J"�N�x�[j����֌@�9R��`w�� PKc��[g���km}ą�;��cMۏ'�!�I���j�k&�Cf���|H�|l�Q�	-0/��iC	N� �c���̫��������4���^Y�c�ĨW+�T,h��>�Q�=���Eb���b[���X����Z���E���ݯ�J�M��I�5����,��r&�zVth	c"� {B`I��:U��x)�M���E�?^<L�~�T�r8Dp�;��xN����\�t痠��i�|l�?v���ЭA2 )�_���;�\2�!!�O8�[M����Or��W�^�����P��Tx�:n��R��x�#HO�Bk�_��M��Q@�����W�'Dy~y��d'���ONd{uk�jJ���<�rO���ļ��i�&
A�0��8����H�p8�}y��9%woq��H� ؂�+�p@��`�e"O�"Ho�B�5g��v'�����}��h�.jy}/[�v��Չ�$Is?K���Wq#7�b`qX��+r';v?V �?�D��$���u�`%��%�g��� �VA�fw�En��jF���뺋@�G�=�w^$O�4QZ�P�'7��y�8�A�5��O"N�2����������npn%�[sA5_ w7M���[�!�c�
�&�K��2���ϣ� �͎*A��0�8ZjJ(��kK#;e��)����Z�6В��r�E$��k1�7�Q!��G����3[�����7&BD?6��o��w�O�S�.�� G{n�'k]M4���83Ɩ
't���9Ds�K��DJ�A�C�~=N�d����/~"[�@dk�T���D�u G7!�Ht`��,ҫ��,�D�qY�=�r��Y/[��
C��5�T��?�;�*��GP!ԼSM�:�г���d���/�d�k��\Վ$�KN��
������;s�X��?5����{�����(��'8,9��6�@��#��d/xD��n����`i��N�YER�͓���W7��ľ��٫=$��!f򭛖��d�cF0)۩u��	T3dݳ��E�ɶΊ��^q���[lP�.!Z��5T�w��^^�ޑI�{y��0�d�hl�zJ8��i+.9�"������S[�=+O�:]&��C�&���4���Ք��L������>��hT�ؽ�˱>����ޅ�2ͧ�
��uZ'r���{-P@��3�w��=��G��cjE}*��s��[����LBb��m�^v\_3�so6_8�j$:.�rx�9G��h�c���6Ǌ²�������Ҫז�����ט��Y8K܏^�N_I�z�n6�f��b��h��^���u"�#�*�ux���n�I�!`N>�S^Q|cw������6	�!�����Gt.���%s��>O�J+���[-[#:����n�3&YY]�O�/N�=M��w[�]0�dn'���
$I+��?�/�S�/��*`��C� �/
�If�"m<"��8�/!�����J?q�+����@+�E���:de>�[�=�1��@�:Kn;νz2Y���tdb��V� �>3s��I78��P���F.yv�r�oZN�y��)���Z��q<s���h_�,���7a�+��o��~ s|�b.=Kp���L���\�s�>^m`��d�7����h��I��u�C�vS���.�L�<i�6��&�7b�t�6]e_���m�H�"R ď\�3�hMI��_������e�9,��FV��t�R�'0�ǟYx�δȯME\l�둶H�+~����έ��H���Jo����kxHNR��t��Z2��O��)k�� YP=d%�"�<C´< \wEVh͓��I�F�K�X���vz%��A�' �0T�QY��gC�l0h����&,�k��̟�:������aT��q�D�!C�<�Lu����HL���HUy��ю2���&)�]��F�M!���M���^��sK�^���*G��&�)#����B�����"<���	��w<WE�\#Bk�W3�Q����
��������鐑QG�Ea_��4�)/gU��nHu�:8�(Q��/������ �(�����h�htvC�{��ސK2G�M�и���/�S��"@Bl��1����t�n~ZJI�2}����i灕���f�S`�fU�:���\��q]0�;e���]�/�u���,�7�=$5�6��� ,D)����4��3UL�~�)�P|�|��vΨs ��ʗ������ҁ?Q��p�)v��?j*��=���H��� Z�=�!�e^`Ѡ&"i����X���0�X(�ZL)���r�&�s�A%�w�;��H��^^���ý49\/�f�xp��_Ya\Q;�*��&�m����mS�ەlL�'9��JT���#NR��̊阠�� �[4�)�td�k���T�@i�ӱ�%��#��D�����L�n����P��5��[�ݟ�Y��:�8�l�Rԝ������!�R'͡��",#b�#�f��F'�	Q�9�3������	
e�Gt��ع�	��鯀.(���X��x��ߞM�44B/	c:�S(�+����6�Á��Rt���{ȸkL��[���	�ӭ�B}IU
�F|��L�Xk�/߅ ����s�nk�	�8:�[ӧ /X��m��>À��D
C�"�h�$��.����^�Y6�v񊦀�Y���
��W���ꖏ+�M#�"[�?��W�7��ૉ���C�VJ�d%����E�G�L�8�|T��^X7��H��4��C��?w ��V�ZB��P�,��`�٤�$�:�{́
�.��橜'���|TIb�T����d�_��;	~I^c�^�B�k�5FF�~��"�d8���ݘB���� ?+ܥy�n5�z0�2{�R`႞D�?��g��_1"�xm�d���� �aj��G��� ����nA2�d�\%ŉ6�K�w�����������*���L����l̮M�6�H.c[���榶��<�p�B�k�����8:��Ig g�f��rv Ȥ����e?�ޠ��FɒT:��[���Aͽ��m�0�MrU��
�y��jdK&�c��ѳ��?TV"�ϖ^�Gg�Y�oИ�����q��`үbH�.s��7l�*Cߤ��-�(���l�=��}�*�խ�~�����.�޳B�#O/�~�� ���U-�/
���f�SK�.b��(W����7t����ʰ%�ݻW��S:X��B�����^�q^��bBz�)�n@c
�|�d!���\�d0�**t�L?0�Ә7��H�X^p��g��h8��ڈ�jp��V��;�&�#��\�_p-�Z+�MvK�V��$���N�r�^�X�³A��n����Fή,Jqv4˨D����V�{hu���16�������a� ޸�Uy}��tj����z�B\v5�ATW��I�K镌��/�5�l����r@Ue	�+m�=?/�x��֢�C-e�	g���6��$�g���3tJi�p˶�xEiLyΗ�/�v@"�{�3(AΗ俶�zy�2wƻ�.	��(:x�sȧ���쑯�i���z�����)D.n�o�c�+��3�r�@��'7eC��nZ1���j�{l-�M5�o�[f8���6��>E��"��y��r�bċ�|��^�s-H2L��S��.�XE��d�]�{���E�&Q	Y����9&T36��OFm'�1�T��d��r����[}g�ꍸ7�a�V�V_x������6� Έ�u@�D]��2q]��{ӵ�@�<�4�5n�%�����j`�Ԑ�K]+�zWŔ5�|�H3�\�^��뤤�N'�:5�u�#�	NwS��9��k��|q�c�k�	oՌb@����$h�Q ��#�9�n�w����
F��rb�v~a-[)� n�������1�œ�%��q\|k�+X�w��H���;m0�Հ��2��n/*�	���h�����4ɹ�A`[����Iߗ�J��t���-����:`r�j%4;���9��������[T�I��t���`{FO�1�%Չ����?D?l�N9E���V�
�5�4�f�;Gݮ��ֆ[�F6-�.�B�,q��������95L~y�X�I��z�_����h����G�ָJP��z~uc\���pw�C=�<� o66nĲBPg��*m�����Vs,���y7���9���u6禚*��nɧ44Jx5��B�9�ّox����'��E؅1g�f�ڸ*�Zn�V��w��z�$��ބN@L�Ɏ��*��4����3C���\�_#��k�C���|K[��������4)9�$��K��8�@�k��Aʴ�}����Ʀ8K�e����p�Ҳ��-c���r��ц1����~�|��~4��3lJy)�ciP��Ğ4]fØIL��s��)�Z����9Z8��k)Vɼg=L�H�jB+"Rt܀⵻�ID��n,�|r X|��ѠV��F�,�>�6t݁����.�s�KҠ�	�򁋆�G��NO5�k�wH�_�q��A<���0e�eH�8�&�K������I�$D0VKo
����x�Kx\���E�\���:��g��n1?�0�Д0�N��P�,76q�d�cV����A��X[�s2'��*�
R(A3�ռG�4�&L��n��L�ע�J��#�4|�HQ�o�u�y���1����O��V�{�3�Y� :Š�71�)�!�o?o�����O��C��9����{.����[��'(�#enA0zg]n~�>(-@O>�@e5y�L����?��k����{&�/�Ȓ!z� f/e��l�:�Jb�r�7b�������Mfe��}�ۧݍ&?��"mY~Dk�[���IM��ּ�� f3�U�[>��&���6����4+ŌA
��t�?N�,�f6�����Y#�M��+`G�w�6��n���z��)\
�Pb���I�;����Oa��^���vc��Yga�� F��c�eo�J��5�Ȯ@&:Cv�ݑ��2�- �Dέ뿏��~��h4�����D 7�0��B��9�m����ǭ=�f`��Dd�W��~6Pq�����g	�j�A��#k�[�je�q�"e��e��>�/;�[�U���J7��y�u�+%��o�O_W���zuٖ��1���ݩ�Ư�a&���#q������$7�mB����<�.�@����\�Cf�h]�/W>7�UΦCj�.B�ގ-*A���F5��-7�~���H���4״����ԠgqƂ*M�Џ�̜�oϋJ��U�A_��� eO�g�I���?#�;�&*���ô����R��I%>�2�s��я�� ���L���J��]���lN�M�T�X�£{��טrN�=����x�6��;ְ;�@r&
.-����J��c��?��&�h���J��$$l�(N	?E��巏\��%�7D�Kz����56_��k�:�%�Va�U�٫�m{;ڸ��@��܌r�M��}@������:׆�EqԽ��s�kd�R�����*�R�#?_�4�l��5l,D�A��8 ���5 �F>��Cw��M���A&����M���U\p�+�(���E4%>ۗР��6����E��6K���F��4��]N�k���b���/E���?�U<����K��&�0W��c�㱚�����l}c���I���z9�x�������8��oɒ_UFH�R,s���~�
H0Ֆ��6\�l꠰d���l���loDq�/I=����8lF#��d *r��� �.B��g7�g�^����we����5�b	Xy�8������4�w�I���꒽>r_F��3���d	�hCL�M�c��L�~��S��d�9��]��m���c�}F@�����Z��.��u��+�yͩ/߃�}�X�Ĳz�ǐ��Z E�iq�E�ocDPi��l��ō�!�8f�ە�V%���s� �
ޤm�0�
��ɂW�L<�� ���t+��
Zg�w�~y�қ���p	cP�ɞ�]ctx��?�y�ě�kH��=���	��YJ&Q:P��Z]Fw�/�=EG]��΄���ս;�����$��Q�O��fն{�߸��d�
���u��͵��s�q^Vv��]����~V��Sz�]��A7�Y�4nř?���	��<��"NL��
������(ӏ"d��A�Es�bT�KA���|_õ�F�v��2?�~�%�/Xl_�+�?���K\	��S��t�J�QM6�k�	2[���FW��]�����to2>��Y8è��?V�M-Řx.��{�)�h��m�o��rwFԬ�V4s_��������+���|ٳ�-��Ȉr"p�g����l�r<��3�B�����P���^���n`_DJF�C'���L��L\dy'���GY=H-e�%fA{~��$}3�= j�q��4�a�SXO���(cՏ �02��`� �����B!* �P�{�H��%V�mTzѰ�6#1�gh!B5���R�WUW��	�L���sN�
k�h=9i�6�I��]:wz�'��u�?�ں�#��K7w�˥�J��AKR��$�E�)�I�y�c`f$�gߓz�����c5߲���S`ͦ��]��⁦��¬��y�B������V�F�?q���d�w�#T��x�[G�u����g4���Z���l.N������OGU�����	��{��c���:�A%����x ��A@�<λw� ŭ1�.HC��o;��t(�$�:���-��j�wUua���*��K�ٖ��v��h��X�ڠY��D��N5G7�1���,��nc�[�9��Z����DYfKg�Mj���$����l?.�TU�r�)�}��ه89��[�H����k�3V�3ȷ.�Z�*&�/�W^�F4@Q�=�̐��+�{��D��I��]z��߯$]��qk7�����]p�S\�y��	�k�T��0)?�>��tlD|TO���љ�ŭg-�
8}��k;�,�rx��%������%�N�S��F�zX �7~��@o�Q]379��|/@'�Ik���{οY*_��|"���p�X�9���*��G��r������(��}k�n�2��y6�^{Y�K�"�X��r{4*V�T���g�r�i�z�!�,���QZk)�Z0��Q&BEa^�Y���T������v������b��'Uλ�5��oىHE���T���=�`�ue�5͚�vRL�ٺ��qz��sݽ0�&� 9�E`+����,�����;���n�g��^�t.�ئ-�D7HCV�zw>g�»����qjI��Z���i5�	��S"<��-4x�OR6}�XQC���Ώ�� S��e�F�|��,��=�2zX}�g<��	������:����6������5^Zܸ�(���a�M�:����;�HZ�W�X؈G+�a�N��S���Y�|e�ǲe:�N����X#����(�	d���w�\��:-�����1	|Ϫ��)����`���P�RC���j�cU(�_�c�T��y�����J>�O��J��1zqNՇ�?�ey�%OLB�!��TZ�ci�UV�� �o�Ou�j�7'�J�c [M��B8�`���^�rC���A�#}��#P�,����&���6;Nz%i|5���ju��}\���}+=qX[˙�\3��eX��C/�`#v������_=M�%��|ŘF�����=k����nb>����3P�E�n-�Uer���..�pS&Ѭ�[�����/�p(6A$--�#d�ĸ�N�lY��Wt����������\�ˆ>#�5����dB:*uƦ���S��5TڔF�鉵sm��?쁀S�����1�_�m¢
Mq��4���j�R%x�wŨD˶���F�I�@�^�w���XGt�&�����ӻZ"}���!e�f�(�K�����<�b�,-�x�ht�Pݹ�3��=��j;C'E�-��3 :�D���jL�J�S�h��u/sx��h��C8�][]����R�?ñՒ,>9o�{eO�P���UC�6BG�4f2�-��O��x=rs�]xc�M�V�(p!�X�;�I7�	TՅ����>:�YT���އ��y���`����>r`9��7�ClBug��m.�:�.s}�7w�����,���~z�Kt��=vg�#�#��>E�+4�,����k�\.Zb�t�Q�a)�v.w�&%>�Ɗ V�� ����(l���)�-f��uRuo�G
�V�p�>��pyפ�0�']�:��[��Lp���'��9]�8�_ �����$h�[|%J	�������\���?h�t����.(�L��^lL�b��$����T�����v_���?�h��B7 h�2�;L�����[#�މ����&�R�� b��mxX���{��TA��i�tvK2�ê�����1�PE�/4�1N���Dcښ>#�-�
�=a�d}�5�����^�;�z����C�Ō?sԗ���B[�@���/Ƞ���2���.�ڶ����I�g��Nu	�57tjr�)Ƞ���*A������]���H�T�J.�����k �-��"��[<����-H=��l�|�CI�l�q�)LθԌ{��Z��M�\�	��m��`��C�_6���[��P C��|���%;�=o7������^B�mC��=���墹����w�q�Kd�i�}��U��t����r
'NB�ІD���Ю"2[t�2�Da��yӟ�{8,m�^1j��<;�}n��$����R���*�_Z�r;˓��qNS.$|���\�ja��<RCR��_C�sl�Z�w�o��v�]���}���W�)o�m�R������{y��o�̵:Z5�	%S�0����Ǒ��DUh�Hf��9�^^.��dZga��Y�Lc���
)[��&r�-d�C����龃eS�֪[�я��1� �މ�6��<��R.�A�����kdlE�Y��/.n���!{�WI��z���]�U�������z��Q�G�*��Wc������Fl ��U2�'�9o�~��q��<�wO��r��=��4!����,��rA���,&F�"A�h����Beq�p ��N'W������f(�m�1\۫xJ;4���>Ns�fPY�*B��p�Ë����7�h��6t��&�m��%���[ᾘ� )�'�]���Y�$����N�����<��!?�/���k�Ǌ���� *��^ K�������b���&����R25�lJ���4\8a�X�exh�U����$(�����x��E�I��;S��;��#ш�p|��3��<��V�i��.�۹1U�+����jD#^>
*S&��wQi�;M����c �:�Ƙ!�ét�l�t�nC<S�Ph���?Q��D��@���=���ϒ���5�b�\M��)޴����pdρ"���Cr���n����vr���)-gw#�YY�gD�x�=��S��so�a9�Ixé�9���1�5w`��C��,:o�EY}"<�T#��M�Ȭa��
E݈��"���t�9꽒�����x�C\0���Uv�h�?��}���b�?c�'���8�6��Ǎ	��3<�I{���zL���DÎ��/B�y�A�*6�i�kY}��n۫�f�1�孹0'���`.6�� �>�҂��S��W�m� �W�./�CZ�onb�u尺8? (�V������R��yp��� �D����uc��R�yҬ	6��?8�k�ȕ�_O��,b��+Y���i�1;^�(*v0˹����� g˔��a`_��^�KHW��f8`��O_AB�u�����]����=�Qb�|�\� ��:�ɺM�a(��$��c�]{P��Qo5�OV���Ftl�O�y���*������A�6Lu��2��V;a���'��	L���%>��\m��Y	�|u���
%[�C�?��8J�T�\=����S*� ���^5����N�^�o��Vi�EG�J�ː��#2
Vu�^�]R�SA��f.�&R��
��U��v��K�e�\�fgpP� ���[0�u#ŭ�1��Gt���x�&�����93�ҭ�p���w�y�W�Ca�>e�t+l���7B���T����J�x1I'��U��憎�N}7�i-ec�j�
C&�U�� �I�v\�Դ�ӰRD2�	���yz�0�I8�?��!�`�mS�d��Y�����|,�|�%����P��Xs+�0��%�L����P�J��:Ή[
��#2�pn���uVnNza
T�#H��%SДnY�J�����8�<�b��՟u�~�3��H�i�sO6���3�t7�X?�Wq}r`0����_~2��՞?]Z6Ʋ��6le+�K�FZ0�h�#0-��1aD�Z]NV ���*Ӿ+�TgZ`�3�2AB .�D~��$uZCe�W�_�Ui�m���1�]AO�rW��EyT ����bMaitrο���0Q-\o�ig�|_�~'͹=П���X�����
����Q|��<�e��O,�� ��հ-/5ko�h�11��P:�InI�gp�:����K8�6�ͺ�ڸ����6=�NUr,f|���[�ϟp���cU�|�P�f9f��w��P,S�4��W��2��_�z>��f�f#���'��f��O/��l�}�^����&�A� 7	v����r��'|q}vw��u|Ռ�X)}������vfa����RӳE��o�ϡ6&�0���M�mQ�RXghj�L��uY�]*��nW�
]�L��u���Q�ᮖ�,8���й�q�K��� �Z_AF;�+���;�W�F}����w�VFhZ��k��6�#dd,��\�\��V/�3���c�.�C�G-HEj�AΥ�4ynF�(�Q1���������A�nX�PY�m ��J0�����E��v��C�Z�~��*`�,LPz�|r�5{c�gWu>���y���,"S�x��LZl�r���%-x�(��Q�"n�^ZmЉ���SZ���n�[�؁h���d�_R�/�C-��G�9s��/�}�W?�C����~}`��\�!��L]_k�=�[I���8�p����ψ�>\��DG�7�ox�j�U���C^gnX��-�Kp�i��/���+�Ayh9�����$hJ#T��:I?%��������u$bQ�:�����i4��aq���	k��A�����T�
= ޺avb�lA���l�=��\4���WF=u���+�oޑ�S�*\���#�#�p�v:�K뚺)d0��:囪����VռG%��`qU�?6b��*]����������Ǩ	�u!�!��F��mZ�b�&��~��{�5}�ی�i�N���7�F������ð��aLQe�!.�Va\���^�� m�K��#v�Ր!�ܭ�/���j:I���\!ُKCJ'����.c-웭��V�B�b�W�)���eM��x��LyEY(^ՙ�n.�~~}4��d�t2��i��F/�;#���O�S�e4�b�D	;O�S,����=�jV��$(�43��
�y#~&�P� ��c�e��ť�4tƠ�:p��`;J�5C�3<Nǲ�y�y�Jr����5?.�Oa��T:�� �"f|
�e#�}<��#�*e�����"-�����V�YQ_�Xڜ���x7���`Z���:伐�E���Q'��۶�F�w=:d�B��f�A�'@�Y0����Tɼ-|zO�S�酨4�xL^!���:<~<b�݁!�-���e��y��J<�B�pBVq�lCR�}ݚ��#��J;s���#�TL�mA�ѹ�8�G�/$h+l��d�ס�Œҝ�v��Gh�������/8��'E�n�0̏���a��� Ϧsej��\[9೼�c�&ˀ%����!�vŹ��i�NK?�I�%�0P���HE����7�u{��{S���3�O�@�ev�Q�A�/��Tj^Ρ��6{.k�@�e�anEg�!�f�mb��z@�<�yGMI�Ġ��H��U��-k.?���u�M�B��Y�R�me�$����a�D{ؚ��O
RMc2O9�\�����I��di��F﷥��V����&��!3��@�Ee�&`-����i"e9��	���ߛ�q|�Ng�_�Ӽ��Ֆ�h���(�s��=�!�o+�^w<#o
k}덛�DC	]ͽg�`�e�^o�äKa_�37������-mC:����id�4�?�>�u%���a�2���@Z��7&�JcȖ93R�N�m�c`��D���~����X)��#wV�h��a�w깫:+�L���"$b�ĖJޯ����^]Q���3 ��Y+֌��ª�����2K?���N���+AóW������t$���kS�<���/Z���Q-��,��u��M���.�F } �����A����K�p@��ޡ:W�Z��Z�-3�"V4J.�I��s�Ի��Z'ϵV})�M���V��R>���>�yf(�$��)�VT"
��\�虎��Ѝ&��I���զ\���DUV�Ée��S��w��/�(u~��|�xu2�}��iD����}�L�eTϮ=J6�d�ֈ�[��w-Fx��ӽ8���ƕ�4�X\�`eNV/>�����w)�z&eрVt���"����ZY�e-���cב<�4�����Խ����e��K��d���r��F�wS��ڞ�Q�V���M�6~��Z{�!��C��֩��� ;z�9w��_M��v��|��h|�m�v�xOMuɐ���wL��'�_ .���
M#Z��/�y�ej3>l��j��iS�J[���Ec���i��M�ދN8�6���m`_��,N�^�_>Dn�J��!���tK��;N�2'�۔�w>2��9� ��f��6.���N��Lpg�W�å!�ZE�H�,?V�j�l���Jؐb�+��I�O(�r&'J�c!+I��K�
��-/
�-�y�W7e"��9�l�ɍ��y@H��� ��[�&��LY>cWڭ�T�|�k���UH��YĶ*��+p>�z��Ւ*P/.X�y�j��ii��8��ТF��~k�r4ON��xZE0-M��i�ܿ�9���śD�GV~o74S�y]3;n��S�Ш��@�C �~"[lvx�~2��Lɔ(�q�NJ���SȄ��"]T���"��P�:(���^��ѢJR���{�o?��&��@h#9o�����~?D&oc������$����w�H�RP��@��-����J�ac3p2�]z�s�>��S�,Kv'ۉ�9e��E���(���)=���n1�ˁ�HQ�E"�,I
��{�=�}QMQ��1��\,�{��a%n퓯����u�l_������-c��8���$�%C�J9B��p�1� ��
����
�G �v��e�\���	��V����%9>@H���������@����)I?��8%6��9���O��-��V����P<[��R5�d��;��������Nxъ��E�!#8Vb;�� �APF��7&������!ڙ:rokK��
HEv�.����;�Q0-�6	��N�H�P�✟�^�, ,�®%�İ���w���^R��]��/�s8�p�'/��]Ԅ_������4O���Mg�j#�R���m�M�"��鏂��&�������t��]X�X��������y�����q��jڏAv.���X��	��������Q�ap�1�Ch�QŔ�3!]��">
���&����Yr�_J9F@f�LQ�FI�
�ؿ�"�{L���u�!>_�k(��F�yHd`*O�)Z���̟�QG���J�����h�7+��-j��.��#P�vs�1\��Q���'�Dn��a@�)뻩D�q�
WSTqʭ���n#�C4��qXb?����⽮�:�;���
F�`���?�SV�ǒBCɧ�*怼T{ߏ@צ8[�Q\�`����f� �t�%�����u�X�VnL}���w"����,M�n]�"綁�03C�|7�d�[2����O�{r/�ɔ���db`�xV�y�Tq��.އ�._�X�� V�h�$�T��̃
�O��s��0�&�bh$}�C(p,D���AX��N���^�)��A�na�(�B�nY	0�S�����n�H��G�drYS��(POEt��q+ds�@RtPVY|\�/�����x�(��2tS�����@X�i{�1`�j&��]�N۵��8��b�}�q+�i7?�e��fhC�v"�n�=.V���h(�OƼ�O�Uw�w=n��{5u�0��P��\w�f '� �6q+�y���=���D�I�վ��N��MI`�h���rR��HE
ʩ�R"<�P�m�y��J&&�f��L�{d�p.��)0O6����*���>|-W��}I�s�͟2x�r�O��c`F��Y��$������t��K�`	�n��o&!�j�� T�L�w2�GmY��Q��a�ߜ�<�2�`_AÓ~�q�U�]��-h�� L��&���f�{� G�JI_ ִ"�C�qëkr'� �I�p�3�@�8�~�%��i�� ��)7�S���
8�����"�Jn�^)�s:�a*h�4��ʾ_��(��j2~���5;�5��t��e'�'�I�A�6L��,�O[=1`�{*~���S�G�h�|��&C�Z6���޳(*�̮m2�i��a8��4�&��I�1K����.v�h��|�R}��s�V�e��Wf)jH�ܯDL�����/^mz�v���/�I1atb�<}4Lq��,�a���$��{�_w����SN�m.��<1������E���b��������8�^�a9�M��6��Y���y��"č��[�ݶ��$_�/f:����V� ���%������AK���_�̪�R��|@O�t�b���Gw/��XW	ԛl֙.�����/�RxN���tb���(����u6Y�پ%�PwҨz�޹�w�E�z-�'M��R�v4*�71U	i����_H�9��Wn�5�����)��<}�>����HP�P��T"����PW� V0�ݤ���6+p��ɢ{���Ȋ��o�cmFJi�v�-���4\[�@���c�m>�n�G�;;�;���MX}ۀ�<j�����Q�0^߳`cW�O���c`��"��#���n	�t��r[�'��%h�b�5�v�%��bz�O��ڏ�y�PDP�s�O%�/�Xۯ��۩&��*����?'���qY �������1���y�mF��|��~1���Պ��)�;�+�l��u燤 Q��\��*����w�J����V���3V�:R9��*�sJ@&�����u伌�.�L:�?򇡨��ݥV9$�Jb_e"�Hs:��+i�5 ��v���S�95�����I�C?��J>�3��V�yoW���jg�ڻU��T%�;���
{�Nֻe����LQ!i������λ���ԯ ����6�{�9�5Y.\P�s��1���Y��t���w\>� :�W�����l+�?#�i�����W	�7�h;��Ú�ʟ�cs߆7;Og���\�����e�ؙLqv�@�n;�#�e�$��9��8+��(���_m;���C���t�;�=#~+by��ǬR��$pN�70�n�t����� ��ڐ1}r��*��z�� ��D�\�;y[��~�zyw�ϴՍNݡˠƇ?7V���#�鶈E������=�ܥ_�9\�)CVF����f�q��l�����M]���Ѡ������xpM�'1=0���㇝��b�3�0+��zE�k�3KE�"�+OuY�I?�p�pZR���O &�������G=�����ɷ����t�	�<������ad�S��M'�A�_|5��7X43� بZ�K'$_�c���~�}��_L>���ģ�#+��uC������(K<�����b@<E#ߠ�&�s���[-+ܰ���/-����C��5`�]
�_A��474;H;�����fv��˞m��Yj��w�=���nL���qU9�Ql/O�!��a�;JV.`����o����\L2t��s�%#��o<���[	ܓ�I�h�*����{a�IN�n\S �g�Њ!o��� S�)�޷�1{>�Ђ�d�%	�DVr$D*d#G.��h	|�Ui�G �ݍ`�K�O1��b���'AUO�T�m���@��ߵ� Zi]�������m�Z4���;r�<����C��b����q�|5M7�D���/��0��o�7,��sk
/IM��RY�I[z	R>�f*B��#�IUK��z�*}R8�@K�Ft��F���3@��
q`�gw��	Ϗ���|$a�b�5.�G����Ů���ӷnD��ͭ`�ˌY8�N���$1�t�^�м�X��̑�g�m�+���u#Ʀg�n��i��Lx`X`JM#�n�����D�%�a(2���>�n0���ğ�����H�����ZwH���_|�s�V*�%�Y�k�tTB:%5���7Ij^����:}�ow�Z4�2��)v0�T��@�N{u�L�iWڋ���b�9��u��ȟ��,Ǌ�>  �o��O���n�L[�?X�@N!�x����v����!g��I�R�x�$M��^	�	0�eP�ۆ3�^���rM0��2!g�.�=�[�|���D9kS�?O�/��K�x���#
���Ο�a)0�(Q�u�g�����S�fuaEպ����H�f���R�~��y�_��E�eɠ�(����iR��.K�Ǐ�e� �Ͱ���y��"h�v���!�1�qf�w����}�X�� ��ߖy�S��s��eFNL���%u*�\}��b��M���󜵒�T�MS��4&PBj_�t�nסu�>�n$Ef��ϫ��!�W����3��'"��,)���G��	�/o�� �jV�"��a��iVS{�ײb?)�$/��u4B|��,&�B���p����O���A5�������	U��]#p&m� �d���7��O����K�-: ��9b>�o~iӑ)��XR#�/G��ؤ�S�:'JTR�g�|���o(�@���o��LV�%k@�&�@�K�0��r���:�j�f�B�u���,qBS[���#��6΄�[m�Y��dZ�;��C��fD�j~+��չ���W	�G�\w�p!��B�S�Q��mK(w�{g�'V)Oڪ�]d�o���Tv����"�|줉H�Sd�pM�#!l���C�d�_.
g'�yb������	Yo�."P����1~�Å7nb�D�ךtb���T���Tmˉ	�S��x@�\��5-Ta�ZbnmaE�a�K�cPq��ҹ ��Rh]4ny]�Ô���j��4oA��\"�s뇟���r+����n6���#��OÑ�J�x�Ph|�vQ����b_E�a/͠9,N��@��t�IL�)�Nq��{��F�a��m��c�J�D�튅3���~�q��\�-&R�K"��N�KKuZl�X�8�z���0�dT�l�����\}z��ǧz[Rq�j<�=��vƌ�:Vt7��g=1%M�]���K�~��MB�5��A���:
i@�X����n<��^0��A���l�~x���_�����U�.KeW��{���G�5��c�#R��3v�RVD���֗����k%�|R�lo�g�Z�a�����i��l�/���Zij9��F�Հ�����A�G ���MV�����3D2��Ƴu	�}'��HZ���4��.n�w�meH��S�f{|�l*Ou�k�20��@0?���B02r�nUn��yNА �G>�R��)�D��-�q�TN]^9�w\�=�y	�3��K�î2h�2w�Nk@��L����O0H�A7�Iv۔چ+O�w2<�A�J"�U�}�\w�@!��ԧ���������~�ao��?͍-:I� h�Ϣ;��sZb\T��%m�ɇ��ଚ&#�th�#��(m�[J�rYŴ��`�-o)�=:��L]��Ä1tS}���ᒐ7�fi�V�ݔ�i� ،A�<�^�e�C�&!�&��W��+=+�<��#7�X���g��s�R��KΦ8M'�8)�y���bQ2�4���O������w#�g�Զ��=��ǢD���E
cp޷2$�V�`Ue��Q�?�(�~	��A����:A(<}h3�)��[|�\���6��L�&1��.��
�t�H=ֆPCj��,��Md��͢�̭/���?St#��\�����A��(-j7�ǀ#�C�	og���f(�*�Q��gO���c�z��Pj��6�%Yh�~V��/|��П�{�D��=���{���9��7�� �N7n%gh�ז"%���o��M#?P��6�?��[��8(��PusSD�������O���n(�N5�?��o��_�7}�ģL����-TF�ty��+��!�=V<�O��u�AC�W1.)�)l���nf��Z[��o�C�X��t��K�s���"�e���t�z����IJ�sU����o\��!��U���%W\���D`�7�3��q�%��,�/��|R�^�i7~�1��M��N��#H��&�tZ�B�>uRo'y�����4���*�F��)k>H_��jX��a��5K�p+ݶ����� �l_h�������i
[�)�~ٵk��-t����b�
��>c��Y����2傟ұ�j�T
\h��y�_��� ���CO�/�������CN�o��0�	�Ɍ=�xP�~��q�z�x��_U�u�n�#*aaQIB׳'[�S��O�e�����Zxm�#���r�~�S��p�A���������pp1�p\���K��x�&��J��LT�k�ﺢ&�
�S�M�(_і�
�׼Ohe1���	m�ނ �#�3��H	�.ocl�$����~~�}�Q�3��a����hRm����ɝC�t!q������xp������=�m�Ԋ��\Q==x��g�й���ǿ ���c�9Kb�-"��S8�fS�T�Pٱc��������$�So�讐�P6��.ǌ�#R}�ˮ�֝ZsA����x��9�	Jv̴L8�p�c�����7�t%N7�l��G{����Crr���� �6ܛ]-�4�/��%d����;"(C�z$=79_���v��A�����ܷ:�3�(�i�Kl���%�E-��ry�!����t�9���GU������[�����*V~���y/�u�K�1�{fdD_?zw����\�V�{� ?!+'��<(���������I�A��Q�ioZO"Ǩb�u�%P�
[� ��q_.�ł�-ݩp�J-&��`j:�;����x�;�:���d����2Jv, ��>�ZAz�.�
��ʶ�0�@͓�s#��R�Z�*��r�C]����$8��?
�O78��?��EA���x�,E�ٺJ�
G�K-���@1���N�P�f��m���^�+Э.�xr�e>�¾_I�|J�s�Ϻ,E`Ws%��3��\���7�]6�J�[�{�f��
U��.�Z�Ԟ%(P�
hh�U|��S�g���������m@�0Yq��%-����V9�,��n���E/��+^9�����aI�����i�gn�"p	��mM�դ*��[����V d�X!�~��X��o�ϯ��ە�'n��^ot�{W9@���0dM�AGl@d|� NW�1G���O
�h;�	�[G���P�J��8�xh��9e�8��P�b����RT:xףJbSݸ���4���<�9��jTU�H��Ƕx�0�Ҍ�{���-ܟ�X��1#�'?:����:��Q� dTR�32�+Lp��U����lD8�Ii�ȓ����p������'*�0�A (�fV�������Z��E�K[r6���E�H&Y�i�.�ӏD��XNC��hN����f�Z�G�9\���g�І�|~��r~�㋦����b�(���B#:�	���I�;9�� +z��!f|�-�	BF�3NL��C��є.?e}��5p���E�i�O�	�*�b�\��y�H\(�~v��������ę���3zE4f"�'����4�Sͺ���3I�&�SX�Bc�oV��|�|U��>>M;����j���*I�w�,d����P���J;
xNf�����ҡ���+�#���݌9 �5���{�Υ�XA�m���{=�1�c��TF�7�>ӄ�� T�C��]�����@?_{d�4�Ǔ��=yۈl6e�(^H/������Tn�	u�c[�Ԏ}��,��-TO�:%�-p��sh���Q��!"���������/Bc����l�t�Yت�8�:x����DRH@䞌!dC�X~H>vw�	�$+u���-f+ ����>��ޚ`bW��k-v��,]�����Ꞃ�n�O��8�q~7�l� #�D��F$���q�p�Sr��k���Ζ J�B}l]��e�C��1�A��.����%�ɬ�8{����Fv�Q��r�<������@��xJ��󞀽D��v��-;b$��m�ҭ��m؆mA@��ܴɜٰg�,�3���~�P���K��
����N?�����r��ڍro�[z>LN���7��:�8���rVԶ����ւ�%-�Po��]l����#vY<q�Iޓj�@��HW����z��LO�~ylL�&��C���o�A��9��Mx�~b�m���"rܶk��~g�9Z���7����s݂��ml-�]���n �?h{xˌ9���^���(d/C�����?� ]s7�Z�^�K�U1P>Ŭ'�w&������	\QR�b�t����Zt�v3^�T�������f������e����:��L 	��Q��A+�s�C� ��_�l-{.��t�/D��ů�$��H�m8n�I�IO��2���v.E׳���m)X��q���EmS��7ձ��Ā�\A�ӱPt
�,l��B�{v]��g�Gk�*gv�c�t�W���ti�F�d�� ��$��	�刀�6;U�,���l!������Iv@F������z
�n+4{����Ț��^��9�����,\��P�����y&����J��5;m>5���
̶�A�C�}-K��{Ⱦ���Ξ��x���XTFQO@?=�����'˱�,e��m`��"��(��_�!��z�XO�]M���tc×g��b����g2��#ڶOD�����N��3�QSR���YV0�mz�D]�C~ߗ��@]Vx|9^~���Jׄ ӕ��n�M���J��%m])�A4<��2� ��r_���?^t��@�m3���6J�(fG+����i����g����
�s�h<�.�xb��S�\�M%��^��ݘ)����1�O�AGgx��U�KhB��Ȅ�1�U)Z�bo�%�4�)�'@��6x�i���4�
��I�xuNI���F말ڟ��<��O�-�%��Ys��zs�i0�N�Q4����B9`�j��}���OE��9�$q����[e�1�u�ar����|9ƂD�Xc�뒙}���4֏ƚ*J�W��Z<R&{�+�y\��A�*qQ��3ڬ�`Qzv WAѕǽb�iv��M���^��ҵ�C����Ե�p���i�HYu8S�@D��1M��8 h��cȰ�ȋD	MK�|"�x�^_����j�`������ A 4�P�8���E}q�r,�3礵uͪb^s��t\��w�,|7��ۥPlg7����/7�=��<~������҆�C�Rtd\���U9Qi���k|1yD�~Q+5,���ȴ�=��j�'���-b��V,Wy���"֔��﹇Y�0C�������y��KV2#�����Y��q`���͇2����	ӥ���Ϡ�p�Jy=1�5Gv�֯J��<Z�/��ѤY\t>m��0h���pj����(j�`�z9�Ҳ�:{VȤf��1Ci;�,�&Up�3�D�j�H�i�p�c>ޓ�'8�C4jOS� 
IF���⭎T��*�eo	�~(J�o�D����$��_Z6�x���J�dF��5.�I�����~��	�����Zv��V����X��pR{_�},�������Z�H� ��`a=K��y*%1)З��X���49B'����8��Q���A	�B��=paQ����4PfG����X���\|;C��<�'&�;��*h�&��ȼ�Z�vq�`/����?�w��U��p�'�A���
-Ŝ,:E����!��$u���X���.��I\x�J���h=����a�g�
B��e��kkw�th{%�d�7���a�3lL@�NŁ�H�By��O.�m7�O	��9,���.��/1��.`��6D�ۄjGh�s0N>k�l�*`|���;u��ނ���}1�a�5ӹ��y�A9����m:�-r�J�43vHK�FF���������ʫ�Lc��x �I��=��!�b��Ȑ- &����?n�*n�:͟I�5��|P�_�_�`ދ�}4m�X?��v�]�K�M�y������G(�����#�~<�pHrl��Ksb�a~�-t]��B@��0a���v�'sJL�XS�h�6�)0��k����|%�+p/�Mnt���0p���"�z��h���X�ea��^�}w�j�s�Q̓T�1�����c�J����\��U�=�~J�3��f���Z�C��-e�9��Kktrk��9�z�ɈHKn'�E�?����k�;N�Ǧ�bf�Ѷ� C�nbĮr~�O�rR�8
�O�"B{�j98$�q�����-��O F`B��1z��2�����9i�����*��vv8YJ-.��Pm�ü�� ���7�S�M/�>�x�x��j�Vls:��P��W,�����ZC���gZ���&�I��'=p�Y ���RjV���io[)*F�ߪ�4kGc �M���O�$Ϡ'93]Y�)G'��Y3�e&ZD��q���5�4ȓ:<�)Db�~<��
��9��F�9��6~;t%�

TϯjEW��f@t�/�]H~U��
Q�Ai�W��Y���ڔ�<]д��у��~d�����ԅ�ۄO0E�F���Bb�ʅq�?���rihX�|�x+����E�E��g#`��q��3�F�Lo�(U�h7t�p!͙~~&ͩ�]�R�^���ʀ]Q��?�@t�_��,����v�f8$5X�,g�U��&�XG�e�h�[�2�9YI�G�I�k�}�5MB�zU6�� ��v���Cu���N�����w*�^:�q�
���0��2�7黹���"����~����J��m��6�c�����Tu��Ҡ�9��0�r�i�"Dq����֤�v�s���a
:B<�]�!ŉrթ���ZG��M2[1{I�	��V��y�~֘�s N��,q���<Qo�N���ȁ�-��:t�ݶ���@6\mF]���'hW��?�����s��;8�����\di%�K+�����U�M�f�<�K��kEj�3<9��Źu�'[�Uu&ݾ�m��� g��0��ʷH�O�T�]�GK�\#6�C#˵�j#Q���!�
4�%�mۙ���� ����g�싫��LQUP�GM�=M߁>%)|������
�7���NK'���z��h9��F�S�a���$&\����,�i3��_4��͍4��N��Q�!T�P��6�Hl�4ͦC�К��[��� �X;�a���$�d�_j�VX��|�D9`N�$�?1�r{�_Ɛ�֛Q[������ZI@�$��*�9ᩛG/�%��������	G���)��k.EA�u�D��@"]�a3W�&i�Bg�:�4߭��������{y�]F�V�K��z�Y��E�Y�8
F���=?����%��M8�� ��hpn��$E${�z����tNնn��ïg���<Ӓ���v�T��ފ�o�\��9��}�˒�(s�4rl����Ck�4��sd�dO4���u#zn���Q��߱����uyG��n��_:ߩ+�N{�?��OJ��m�H��p�^u�m*�[V��d�b�` �:R������V!&��ӈ�08"��NZhT7�ߛ������ic���XFnj�/Zך73�x����v�۰��-f-��΁b�zK��4&�o.Nb�t�K�����^���̳��HU{
1xᖍ�ߔ�YO�r���J=j�j�����w�*_�X-:z@?�K�XZM6�~�o��hc�q�x	1T���jk�]83�F�}3Ow&����d��m����]1�u-!F2��A�R|�����8jC�������ж���%(%ʃ�[�/h�b�p��B���1 A�B��.�C�$�a�r��v+���l��������|ܪw ¬\W%+۰��k�٢J z�jA���˦�3	9�}��A�K����r�T�CZ%4���7K�N� ����$���9ҕuw��'�#'���k��]�@j?�|�	��9s�*���Kx���}�x6�b|򧒢3�'\���r�`�Ʀ�� �]���L]�q�e0_H�:��y��t����[F�N�[�hq=_:�����ܛ]:}@�i=.(�.���.�S��D7J���'����f�&�s|��O�%�˝)���s�=#��|�$7��:t����x�
(�m܌�l�#փ�='[7�s1���d=��'6��F+_�^��RtpN-s3=��Q���ila�_h������_Wr�+s�F=m�u�k\ӼAm��!��؃��-&��õֈ0������+���܍�Wꀋ���,g�,W^fO݆�I4��ԗb��!�@���2�΄��ƽ҄�>�n-e.`��������¨�����ըvAke�L�R�A�s�І�i�ȋ���R�%�Y�?�g��$�알�J�p
��[�E�43
z�!�_ϊ͌ug\�~��pZ�p4Xt)g`��P>R�`��
�t[g���|�l��-:���]~�:g���'�����.���M��6�A����G+���G����o���@�EK����c)�	��X*�Q)W]��b���&��C2�ؓ"��ӏ{JvV���%t�*��9w�1��5���/�f� ����y4y\'e��1��#o��{���5��^!�H&os�QA��s��7� f�vәTl]�gN:K<��3x��'D�4+u����Z�۬���O3V�zH�A)���>@P�|���N��s��.��>C���d�����t�G��>���q��m�s���w��W�,p�R`Do��!�J��GW&Tӥ��>��՝�)G���oA�/�ܳ
�N��0��"����sch�v$E��H���gΓG!-M��ٙi[�T��-�x	�u���_D7	7W��h_q�x�ɧ�k*��0�n 1���AU8��t�շsI�X���>M�pj0Y���c�uPz�xgz�䆈�*��z��d�f�~��~:8��ƿ�͵�����z!ʘ����*�����CW �tjU
��3�N�9`�u�W�+��Jk���ڲ�c�����Q�6�x����H�xX�P L���F����!�9^ͪ��#-�Y�z�A0E��%]�pa�}������J�)+~�J��0c�����<��c����q1�s��L�=�5r3�1V�����ꃒvR�$�A�O��~�U�/�f�'de)k�A<�B�@��B�d��!�<X�zYW�**��5�M��
���]a�'$u���p����̭�e8.�M��c��7o��c@�!@�)P�UXE�������>z�ۇ����F��0ea�p a5?��4P����^��uTx2&l���ɸ��~�ʜ��OG,�nd��9�M�����@��ю�3pK�L�dB=w�Ζ~��3Ls�|ם�n��Bd�$(A�:s���u4.`�����eeм �`~�DDX�̍͢=L�=>W�?��u��(����k�E�6kּDD�<��=�w�"(��eqψ��b;��\�4S|�7Q:�H��8*��m;�2ܛC���^�qd�)��`����D/���ú�(
�	�	��M����ĦϚ�?��ӫ��ɸ��}>�v������l:{�KaoL�4x�mB��@�T�Fbj~l�
Mi �ڇ��Ra�Ԅg���MC�����*�4�[�w�p#:q�r4�*A8H��/��{�(���S�c�r�;�s���*����pF����),�dzk��;�^qH��Z=7F0v؞O �2���w��V݄��J�S8�8u����0���d���8�@�z���,��9p��
j��gx���g��~4S�Ћp
���BU��ʬ³���_��e����N�Ø<?�СR�
L�*�ׯ@� �/M���%2����\mqbE���i�@�p9�� B9��{���/�%秅���>	�Bb'a�?S���ǭ�9]�bs��ĺ�="�|�<p��3�a[)��������{ G�e��pf�¬�u��k����=f.��ʅ��p�N�ν��aƨ�xw���v:�u��5�H�z�L�Go�H����_�_`�?��dm��W���=����9F=�L"G'�f �֖���r�\��E�Lk�{"��Iހ�VS	�Ɣ\�@DW�S��FM�D��7�ҁ[/h�u]�.���:΃�|��T�N5 4m�c/Q�:�������:R��
ukx �p%�C��{�����$��z0���?O*f�4�B��'M8>�Y��������f����=N��R+$���a
n1up�Gl�>l���D���76j���Z�����:�Q'�܄w<�@��G|p��j��f�_|rmv2��o�4,ϱ��,]2�=?�f�A@xٚ	��j	,�,�D�����(��2�e<&Yr7t۽P�wW$��1�*D|-9P�C���,j��R��!=�B�/�P�hc�kB�'���(ؤ`E��M|F�)1p��Z��f��2��rb�Go�pqJ����4��Hh��}���S���o��9�Q7R�J�J!�Z�Z���m;_��7�����~EĄ��jV�'#UgM���~,���3 ���S��Iф�D�D��F�E���I�xi��&�OL���]XăHT.�>�N&w�o^�'��T`ƭ�ؑ�������X߷	#�ab�(��[���y���37�̯��2�TJ��Ҡ��r����n�%�B�l<k]�c�T�O�e�Inw�j�����T���+����-�;!#whg�*�� ��5��*���\z�C`��MU��\3?b��E��A�ɷ�&Y�'�<tL:E��F�Ų]�7�,������@��x�^x��KÌ���z�j5Y�~�n�@C7�?z]�e�΋�ޕ�Y�đ/�N�����G�T�ǐz�	�2�NW��C!,Y���y1,�Nr�f���g�k��T��Vʒ��?(cM�p���'��x}tj�{`�mW�w�қ6�pG�;��=ܙ�i2�`;кz|\����+`me	�svVg9Á�^�TS}�e���>U�[�*�h�%I,E9�䡿�Ө�#�?��u��9y�!'&i4]�U{�O^ː�����]��GoGp��Q��՝^Ӂ�!���v����eCdP,B͊=���@������K����{�m��R����F�F�><�����_�O�|�"���(�1��
�{T)�bcz��+Q/��a��>jG�0K1�q�f�$�4D���M�a�Mmf���S�Om�qEFY�`����ž2 4���/b��\iJ�>o� �Z��N���~�ZzI��)HoF_��an�����.�to'v�{?4p6�R�2��F�ˉ���м��i���CJ/䞵�)��a�������tcL��#[_�I&���ޖ��Z��V�тcg^-��q�"]%來��6�s�Z^t�[����������3�š2�4c;4"++�*�2ި�R�v8�6jfz�A#�¼+h��	W���N�����,U�
e�R��j��&�k��N�k͍��|������L �Yr���~Ѷ�P�m�$\?��_�{�0FҔ��n��r#[�"���l��⦔~�jٯ��t�9����ԉ K�/a�A��fedT�̻��=����U�x�F��.Hx5��6�^P��۪�O��;�S���"�Y�-��4U+�ST��뇥���ҳ��Vy��4[8-ˎ��1ʉ��m���"HT�?���2�ؒNpYd��q��ά��I��A�U�S(�vF5/#I!G�������,�œ/@[�X�'}��TP��B �_�a�Ö�T7��V^#ӞE
�ܗ��C�kx���D'�;�A��Z��g�����SQ.Ex��Ѯ#��r~�8e�nU��i��w�2Q�!��u�x�ul� n��x�N�*H��IlKZ/�!��V'��	���+A�42��	�w����%7!3�u`/�j-���+C�h3�����ʡ��X_@��\ �� �0�?�AR���o{�:��C��Ĺ2��lFW��r�h�{�73ڔ�����
�5�8%Ax��`������������@5�C��OZ)�ݼ�j�3�52�Fsh���.�l?X��[�.�OU))߫��&z�[]ggCe���IǶU��cK���-"`��Ik��V���f�ʢ��Bb��ܩ��J��S��0O��N�-f�����Ǹa��!N��.�VSz��^�f2S;	�?�5x���ڍ2�e�JNI�>�N���lu�Í�-`���wA z��u��zN�ԭu�V�O�_1��=/f^��2�/�OI������
���F���id�]����-����AY�eݔݾ����cܚ+�)�����Hoɔ���UHS��Kh�d诟�=�
}xTػ���)��/����޶>c��.�Yw�����ٻ��Ծ�ج�h�ǗM��eQ��P�]y�1X�mf9`Ƚ�vD�3kс��� f�^��ZP��E�9��dc���}�Oަ&,��bL~|-%��G3�2�����C�]��W*۩׹%ס�<=��[�*Ŷ+`��o���$Wt ~ �_�=�X1q��D�7�m�t~�6�g;���,
�?��������e��6�,���d��ָOp�W7@܍�J[�y^�U{t��������i�ӣہ>̵*�߽a�}�=Q�uJ�6$�Kג�1�=�yQ��.삳���T�?��d7�?�j�6��j�>1Om#���.�p���j).P�fIRmw�k��)S�/w"�*o�E�Qe�Dfvn����4O���3nG����m���w\�h��l9��i���&y�y�G�=�&S����w�iL~"=eֿJ�B�:pȯ|��#4Ӂ�)�b�F22{7���z����}�2-}����13VJ�k/k���^���(�X#��vJ5Y�`�B��G
�ϡ᷼0�2�|khLޫo�m��@7X;n�@/�D�TaA�t�ECƏ ����ѕOy��+��@��J	+�b􎙘�L�<���;��癮�ng+�hP���I�B�����i�%<��mb֑��S�I����H>?^��5>��������ef'P�)����Qg�Pl5�N�8P@���Ҫ!s�3��\3P��;�3u��a����{�}OG��ZP-��8�՝*��q
x�����1W�8��f�zz���$n�<��\^��,��@�h��f۫h=��h,-F��A�$����]=��%o�F��(
�m��ݮ`)�ݦPd�q�?h�>��+d�Y���H(:�%�v��Y���!���M:BO�����.+�x{�Փ��U��+�OZ��sO(�z��5��A��d;�Q�wB��86���L�g �%lcЦj���!�8���3�w=�uO@�ʽ���NFA�&8$7�D:�����|L"*g�*w��F��ё��f�jP&���/R�ö+w��j�}(W� FLhҀ��,��-{\E�R�&�W��fz[���Z��k��U �N8q.�"L���c��n�����jI���_^H�]X����Ƴ Q�"�9�tܒj����}��a�9j�AF��u��%�DZ��*���]V��'tS�Yv�d ��/#	S��MH�y %�G;��Wz�mD:�g���x?g�����{�9w(��>�,ɜP�������U���k���<}�3:ET2�	����|�Z��~ݰP(}���4[��l�IV�6�x����Tu��u, �H��������3M���|j[}m��~D�E���F��E+�J\�l�5����w�o��1����l&�z��7J�bH�O����� ��]�|�V ���t8'}?�jk������)Soz;�I04R(k�/z��hP�$�ܑ�e4��:7��a��'�6�@b"m�*~�2B��
@f2,�i�U<�F��Y��[co��Dk�]���3\�\��u�>v� ڱ�E6
Ҝ��XQE#+s��?<���:��g$�Ax�PM�<�4a���N2U_D��p�_�*�=�n��N(K�s�.5g�>��7J�z7qz��2��=�%/�Y�U)J�^�hh&�)P�U,܌>���M��4�Be��?һ��4A�{��ۋX^���T}N�:�*�9���4�5A�Bu4FV�-\�5J\�Ү�on��������y�*��Xb�<7���7��b�G*�Y��pY��!�Q��灈N��t*l�6�G�?���;�M���s0&���4R�[�RZ1I)$���o��{>�H�w'����a�[q.�w4������۰���/@$u�?N0��ta�Hn�1S�
TY�Wp%8�n}[(8+��P���b?��>r=1ӣ�Ll[�,�yC���>����m{���5�H|ĉHe�%��@�R=�2��O�<]2q}"-@��7Z����ML�E�"rB2���.��?n9�?0�nԖ���
X/�nn2N��J.�{K0/X��m�wuS� <ϐ��o�gs��+���-7hR�-�H�G��b7;՚	��ނ�A������Pp��/{�6YLs'8�;���2����V�����g���}�b�Ƃ�|M�t{�|�nb���zGw��1}�4�s��x��㻯�-ϯ�� "���?�5��j>^�tRn0V�b!ʊj��~�t�GZ�#β�]��2�����)���yT����	m�
�bӚc�>'0X�h.6	ݯ5�.�y�d-��χ��##D�l�	�O��J���� gU+��I]� ��M��B�U��}(Jn'�űk�����o�= ���z�2KW�����p�w
�����D"�)^Bbѫ��hUx���������1�Lֿw	_�B���eJY}��T{����hV9`S?H�C�w�W��Y�)?���?�yd�p�eĉ�����Ep*��Ha8�pYU���������S� A%.�/����f����d4��B"�o,�w���ڹ�S�+����F�nY�0i��٨Uڬ�H�^��>PD�D	�J�(�`m�+��QL1�&��H�'Yo��D_x�joǚ�:	��'�` ��u'\)��.�uL(��h���B'��j,�0Ϩ�@)?��a6���U��k���˱]K�x �'B@����%�U�

Z�+���rn� ��+�Fy��(0�l�/)��?�q$V���F�3�!Ե��6���<�����g��	 Q���a����P`2�<9���E�����D���1�����%�_g��w�6|r�lr�*X��� .��EO���$gK{��xa�MQ2�]r.�����ǡJ�������t����^�C]�@c���y�hSk��zh��1>�M^��2ZWvc΍�Tr|��ș�-���>��˕E�'�y�"%ӾT�9#�X�(e����/��5��w�U8Ǎ��w�����U��c�Q�E���<k�$f\)��ȊH�����ZXy��@�� DC�9�MOl $�o�i��{W,����N��t�*�-�B؀'��ko�o� �h\^7n�K�w!�*�b���űM�-ɜ~$B�K�/���f����1֚)6��݆���x	��D��,]sp^3^�k]u:���=L�Gt���$!*@}�̋Xt���OqN�s��R��&�!wL��!d�{��� ��COk�n����]l�:�D������E:�3N�	��P�?ڲ�ۏ���\��,��c��{9Y��ʼbJ�?��sL6��H{2h�&5Z0���z�_��a0�(���l��}�Cz�" �wl|�8��ԙѥ>��p*�"�t�t�O�w��A� �=�����
	�F�!뱊��d�y�`�C3�����sxGi'?R���F� -��8�ƨ���(G��dgt9l��o��b_�<{��	j�t)�p���])��0�Fr9C�-Hڂ��y�e#���٧�t(<�r`M��AJ��LV8���ɫ�|��y�0!��/��4j�Xo?<n�]\4@��,v�E6�eB�ѝI� J��A�_�T�#��������>�*�M`]��Dz� �z�?J�i���¤���!�h�6�~�J嘤����}44�UW��.�%�&�_._hC�5�B�*�YY�l���}~= 5�k����msw���((��
�X���(Y^{ng�{�]�ZS࢔-�1��N~9]b6E�Y�[���N�<�x�1y���E��L��¬uu$9��!UL�U��>5Jpx��`V���}y�0QIHv������r7D{�	�LB�;r󀾽	]54�ލ��S؀L��2cq���k���Hj�"����Sx��2PW������*�� �OS_,ѷ�=��uΩ-cB���C�>�TW����Q�d�`�8�A�-x��OA��[n��{��:��9��3��Kx�x~������	�V暗���v�(����	���=�Xz�0�#����q��܇8��(7s����)-�/THl�]l�J����� �84Bow�ݯ�a-]xw;�>�u�\�-����_�����j~���7��IE��,��!Ax��^�"Ti��n&/���"~�����4��&�\M��V�cݽR��ʹk�`�������M�yXВN.z������F���R�?�|���.ǽ�V�b� V��z�g��Hb��x�X,���.�`�O�
������|H%�yjr��q��VA��G����9���~$���?����v���\�~�=�>�7 �+:�2b5MEA�:ƒ��p�TT׿Ǝ_ ��(�g��5���9�w�ϕ
|u2�GRqM�a"� �aC��q��B���J�����+���J��W�P�:�&�1岟`%o�w��\�]vL�ȷ^�m?p�h���
�&/������u��"�[�湒��K�&C�IJз�fɢZ���h�U�N 78#�bo:����� �Oٙ��.4��B�H+r�Y�J�PoD����B��D(���w�1ۮ!Տ���G@�Z���}9�DE$�=�)����w`V��D��[q`�oKԄZ���y^P-�zq��L��"yXY�}Ɣ)K̋ȝ�|���4$�x�(A���y
�z�&�&��+"�m?(�0q_q�[�+NR�c�M,��m�)���R3?*���Cl���:!h2�,�F�g�n��[yp_��>c�0<|VЃ4�)��^4�[����X���5��s�-5MԶ%�@<��TU�2�ΤR�~�|ET�>���)Ft�x '
4�	C�6HbW�������\�d�]ͫ� ���<���u��ㄞ&�^^UY�������%�XuEq�����o:�u)�&v Op��6��KA���_��Zs�Y�]7�ʕÛ��o%��j��PS�`�,:5J华ܭX��T�׭.F�.U��EE�ǚ��Lʷ؁�@<�a�/��&�~λ�Б�jR��j�,�����-u��I�"r룤��_{�֜��!�Z�?��i�D�t͙�̆�P<R��zg7��锎9�;١I����]NL�tñ��5�� �^��nHq��+]����Y�}�M�p�Y�x���h{n�Ĭ�4��ƛ���.dN��P��b����Fq�\_
~���&S2Ę���%����0����Y����|�"�c6�GM�?B�2���Q��	#Vy+�ZV�{.��k9��}J�G�B��A�@�7����Ĉ$2�q���(3yg���Ca0,^mS@�t#���B��ػ�58�r���^���sj"%8#�bb��'�æ�j�����ʙv�:�"�W�@�nvh|YQ$�7�89{0n�B�Kv����"#�e*���
b�i^��z�8i��!��,Q�M��@Ȕ��Z��f��]dBl�WO���u ��x:�
K�gY�FU�
��K�eNN��q����3�r3^����ϼ�EHYq�!.�ĺ�O��P��[
��ƀ�T%���&?��ј����s'k��~��LϚ�%O'�l��-E0�U�F�\r�A���ǔ�"��j�-�lh�:�7QU-�s��H��F�ͻ�J���?'U�'��b�M��{"�aO�~X�e`���I?go��)��1 Xl�I���4_�� ���/uP�m���g�&���+�f�q'�D�H�T�镫ut^�uo"3G� ��k��u%%/H��0B�� [�>XɆ��,��M�ϭq�R�F�\�*��1�sfq��l�\����������h�1�$R��.�&�9�6��H�o�`:~}��.3�(�*(�n�
�.�Ov%�FB'x?��R���bM�ߎ���!�t��6I�'�U�<䇝����;�-1��+�F��9�_oQ��4�m8���vO��1moc.����(����=B
c�BVI��N�ί>F�iv��<g�Cؿ���89�p<�n{��^S��� !c����9���U���\� &�Y�/R�a�*�B���3��0���ֲX5V�y7��'E�34����~j��	��i��.K]5�ý2���?�ф�p�v%�@+����w�R׮i)�JI�>�Z���F�2�nf0U����+���j��)E>�`�y>5�a.혁LA+����C��$�,:�U�A^2��~��h�pDL�}��+0�\�'<�ݎ9Vq+Z�9���*K�?v5�6��_j(s���_��tS����;f!��nW�t��G�Yb@��"T))o?9+�����i�P��gLrL��+��3��C��"X	)�� a·�J;�}�{�	��[���K�7�1��m0Vd�X��,io,稲�c�帽h.Yھ�ֳ�ƖJ���wN��� *�C����������g����r����������:�bъt��^��EB�r+�֯��[ H{������l���'��y���u� ��e�v��֐�s��܈D����FK7�=���bӳ�+2o��q�\�J������;I):��nvi��zЊ=��Nt�G��nL��2wЈW�w6�����lmu׸�+��ch+贱1�_���ϤpN�$t ��&�^�uA��L�(�AO��|�X��x�=�w& M>*`�4��)�@F��)4'0@zjjcWw�F �\
����@���$�<��W�X���������ut������،�ڢ�g�<�Fr+��;�o��i���y�Ĥ��˼h������Q�c���Ӊ�cOE��J��YQMv�c�����F�̫.���Be��S�*{���3��)
o'ɛ�F=�ֻ�!-3�[�v��q[j�ԳH,��Y"O���*ֳ(��`s҈,K��QÃ��RC^�= En��Oi��dX�u�E�:�\�� 61��Ԗ�-�1Ж]i�Z	oR����UM�-�j��`�L>����:ga* ���{�G���ߦN�N�����$x�h�U���wC�J�	x�e����.�QXݗAW�{�K�l���d�<��U���/@q�Zd(������D��3f���BD�\^%�0����̳�AW��8s���Y?�={�*�!��S0Aگ�~ъR@��_�h�T�Dm"<]OJ��t�f��33c�'��8�&$������k�.Ut������}Pȫ	V��C�]� *��߻�_1_Jl�m<��W�z��{�׌�)�g(ë��R���1��s�|b������J�#����,m��_ǸB�r�E��z�������u��s�B�!�gw� X�>�U�ϟQ��<�d���D��޽L0g1�s��S����R�u^�8�N�0Bb��cP�v|W�݉P��uR��*1�4x��x���z��ĉ�:b��B��pǓ&��#�E�]6?�/����#du)�w-��ɪ��N��_{���As�@�r��RiU��`���?�����V?�=;��tU�}P�ڷ�P3
����>͞����6�Q�m� R���5�g���mn< R7'g��ñɖ�쵃 5w�������r!0k���h�kǷ�)ޑ=d����YB�[$� MP���)�����5k
�N�~�%˛-}R�vD�Skz�*2,L��9��a���+���#��lխ�8M�����nn#Y,U�9���G�Z���i)?���L�+�=e hʮ�'�l��6Է���*��M�*x��E)j#Ҽ�Ue�V�4lkC�A��������c'w��R\v{�qP	m�U���A�͟���>�O�Ӗ��gOK�-����m�;����W�jt	qf`�ιNJ�ͭeu�]c��Z��8�Rt�gm�FORy�S�a׾���Ndߥ�J���s�}2���+\������V/+�)9��&�%��]�bh�#�WL�<�䏍�K�Aؑ��<��eJ�D+Y'h��Q���e.ͭ������?~Ē�f�R�t���~��Ԕ������'k��lx#P�Q�%�I� C=�W�7{Si�2E�3����Xl��,���$Q^�_��}����[�w�~��T���m��F�Th�f��2
�s�y�b1	�D��ߚ�G|�i��W�~���}���Հ�nA˻���o��c$�ۋ�|xo���?�?�=��?����OjgT�aנ��X:�&?�T`gh�P9Ž�$Sr��O_���u��R��~�����Ld{��qa���m�OnS��{��hy�q�gu��,���:iK�`�~�8ɸo
���lq��%LT���ϐ���k:mW�>��"j�b&��z=�-Ej��y%ݦ������3�G�=I�^$��S�_�{�����\��٤ޑ�����zQ�N�1BNf�����Z��`�b��B��0o-�9zj�W������#
3ArBD)U8yd?���u
j���YT��D��˨�\ˉD�A�#�N	����=q+4AD �:��4�1}ӈ�����>C�2�r���U8��3eǬ��tmk;KA��n�M�xZ)X�B$0V�`���j��YZd�-\��159
-�;ꑶ���fChh��i5<�6l�z�Q�? �Z4t�����/2ن��+;�<-]��VVO�{���+���G��B�#�"���.���s�E0���kI6d��IDU��2�E���䊺I��$��dS�!7K�^�1����+䅻z��gF���,|������A���<{Q	n��T:p34-�&��0^=e��AIr �m�����(�ff������]Ɏ$��#m��xo�����6���m���f�Q���W��#����/�;"-k����ݺ:�T�#Q-
E�����zZ���P�9�`����r��]�1b�z��KR�.��0���)��V.b�}�sy�ˤ).�yy~5]��%��!�;?�/)qؠ�et?4_"�H0�$�^O�91����d���8Hcl���*=���b���^v�P�I�Lo��7��_|���y�&i��Y�͔�#��u�����Հ�Wl���-$&�C�P��~�U�w>��4ZaǦ#ՙ{�*���r�����~�n�X0j01�1�Qp�����Kk����:ў�N���bUoXmԢߖ��@.��~�jʲk��,���I-��I���������Z��Ɛ@Y E�p�n�v���9/>s[�.�ς^��h��̽��Ek�Dd�D�x������B�Z_��;��^!yt��	��L@#�}JOBt���P�d��
�5~-)�(�0k�t���A;�Y:�i�r�����~&�~����A�,jFjt�x;6���5h�z���ܕȃLB��l���qW��z��w)T�/q"�����/
�~���M�*j��+�jHQ�1Vf �j`����6��Ĺ�?�7�_mM�]T�y����*~��"���G�b��T��;��~́3�]"GO�˖�;a�H{�z�op�~��m�����V؅M�lw�НX��:��&��Ie3���gg*��:z<S���f¥.��h�l~{�������f�?�C�F���vAp�]UP*s �������ZrQ�qH�6/����4ǥ_~�(�@O�?K�7j�Zlֳ1�6��Dh�*����}Ԕ���!9W����L�$x�RZ�@=���\�&�j
;�;{���*!�ѥR*�^%eX��j-],��	/'�����������cM�)iWk߈���U��p��������hݼh~ۦ��(���S�A�c��{G;{�.����̹�iA��U�`���A]Ҭ�2�.�У4R6l�jW�S6)��Bm��F�7U�&x�0+�2�ws����v� �dPU��m��?�ܽK�o��4�?2��ە��2�ɩ?&�a����'�֌}~g��z��h�ĳ�X#+TE`p�z�Np{�X��&�) �A0C��8a�4�ѶE3>��`Īl��/F�m�J��`�3M��,��
ֹ�X"1e��������v
�	�CA��V���\G�O�~��D���^�|��?G5S7�P�'��̥��(�5�Ʋӧ�j1˟�R�]�����#�;��z1*7积�F��g&pp�* �@JU��aB��&�L Mg��n"�T���#1n;������^����U3!ѵ�-C�`�~Q���]�g�2�Р'���/� |�1�Nk�Ϲۅ�ڿ�˶#�n��.L����2ӈ뉟�5'7�<{�")vV��k�:x)>��<��=�yz���Q�h�	�:�y]H��+8B6�����תo�g��DH.E�O��e"�k�aC�ͭ��RPpj>TE,�V��	�ٙ(r��A�쓜Ʋ��_Y2�W�h%�|P�hi����5��$��K�[����fF����zؑ�4��F��y�s��R���ŏ�F��R͟�s�����}��^Q��:.��у��/�&j���^��夬�~�M���_7.)��v4�
��&���!;W�#ٕ�)�fdCR� ~�̘7,x¤+a�,t�� ��5 uI�]'M��å�g`U�膘?�����rO�7�N{ �U�� �/�h��v���N�Om��BȎ�j��g�\�mq����k���q_4�r��l�Qέ� _�
�Q�r�3���y���}~�Y*D�AZv�Z�
@���Qu}hJ�	V�I�S]�����4L���}��N��"���B�"X��͙5�QQ�;�g�k�H��q>3f�F�(�K+��������(yiH�G������,6�>�8��g@��CD�?���|�\?����
kX�g�V�J������NuY�z�g��ϢS8��O���U�L�?�����Cu{����A���8�s�����3 �� D���P2gs��Y�x�QQũ[��K^a���Dr�u�A�\m�{��1�.��P֐
k�$(�B|�7��ئm/o��ߠm�����8+�R0��)�e��=�Xo�W��>Xf{��[`��3��xE5�]��fl�U���Θ��ȵ�Tڝ��K�θ��\b��śPz��nS�8=��F\� ��&���U� AX������ �EW�U���j'J�`XT�� <F}(�aU�0.���s]�����~����Q7>���5]0��`n2��զ�]�m���u�p"0���0�X� ybFّ��FY9{t���w��d_��B���c�׎�,����]#������������~\���+(Ǐ+ŷ�נB�g@�k^�9�U����}bo]��O��9fw�0��6����Ʀ���,�<=h�Z�K�(N���;�N �%�؎���6$1��F�c�zP��8��W��OPM>�8*Б���Sb����a�����{�^�v���w��+��_�W�!w{�h
}`�daO���m2;!��� ����1eh�YOOG��-.]�G� ����Μ1���G�^��zNSwi�P�Lf�#��+m��4�<y�؃ ���<f�N��x�s�Բ��o��Me-�"xyUn��+"��h�T�_
a�<�3��;����(D##Ǯ��P��_�k/6�]�??�@d�T����WɒPoǖ��)�/�9����F�ŗ��R���]�Eܬ��%<D7���ЦN���I �*^��尳,�@�ޡ�X���:!��2C2�,(a:)�����b�
�b�Q�(> +�w� ��B�¢.�@���-RX�Q�z.���u}^bt?E��G�����4QwtI 	3��}xoَ_y���``}�<Q\N��c[�@S%���bE�����I�G������j��X��O�7�Л�m�G[��j�hJ0�<���dY��X$�����=���"�q.� ��ꃗ����A�� U��b71�8(Ի�����
����b��=L&Xތ-�8�)dWȧ�&_^��7Ҏl�ZIC)���Y��NK���pƧ���6��4���F�+|8�$(���d֧�����*�W*zKK��c�bhl�2~�	����"�y�L-q8IR��u�R�e�v�k�9��v�)����2nr[��N����2|a���U�0�%[WT�_�Rղ�mջ��X&���4���i�]NN� �ѹ9����Y��V�x���K\;\8�74�b�k� X��,�?���m�9���v,O��`����\�E1+�*aZ}'�k<R��g ''���tQ<,��E#����z�*����Su�:�6��f�ˏ\瀖IxS����w{��e�� �'�Pp����F��9�V�G��?V��Z�r���H�}<����R����~T��0�o����~���kq�����sr�ݘ�;�Յ���Q55+��&���U�(��/|ϝA�+R��DO�(z�N� \X�ނ�nm��zzj�,,�M������dV��ڴ�4e(��;i ��]h�N?�����=P���yb�Z���:8I1�f�5;���oF��t�_�쏳�]��v�Dn%n<jf���r�����&x7�#P;RәtwĂc�Z/����)�ŕ&g3���P�l�{�WЀ��5/�D5��`��e�'{��|��NƳW���o<�Z�fY�s&�A��+��D��:��/�f�J6��Ғ:�a����ifL�Հ�N+I�FB�1P$/7G.��|�t���	9��!�]ͼF|��G��S�j�ko���E��FQ˚���G*;�Űٝ�?i�Br`%l�
X��K��_�c4}�� �w���+�k Q���:�?��@�A�Ϳx|������	[<�u��T^��Ape�.�=�r3+������X,�;\�lz5��TF+�0�5`D���
��t0��(��D�ut�Kٷ >�oQ� j^���}ƥ�Z"��[s��a~��䜿}{gCeT���p%��?�^��U�+k,�}�?�C��k��[(F5��&�$C���W1>���c�ۆ'��Jsir�V^:x��x)�)�B҇�$3�k�B���n̶�;�A�osq�W��z���%TE�74��
s@p�@[&�$�f%��g�]�I|���T7��H��$����߽3�P@N/SD����z*�P��j��짷`w��T�K�7�x��4�6u�`����[���ߍ�d��̱���4:��%����ݒ��@��3�hrJ�/q�5��!�A�y	���>X�l8�hو��v��������زHZ;�m&� faEDMv�vgD�� <ݗ!J؛�o!�8����R�)�&7�尫�4�U�o�-`�m��J�ISp�<Z
����V��j��_�$�1Å&���z9�JH�ڮ��PK�����Y�X'p)J�s�@��4�LO<���̖Y�=�%{m���w/��|���rU�aV�c����R�6�!�r��kc�/� �:�W-�纉�����
�g������'��Ѩ���Ȫr^�]�@[��y����F�}�ϞE��W�y_"K��!�K�Vz��LK�n3��y(���=�یQ:��D���1�q�NYN`�|,hd=�`�JPg�ֺT�_Y+�u+�v*��Cf�W�P��h�\1�^p�w#�n��� �U��V�Б����m���lxm�����ăc]���`,C�P���Iq��Կ� Q�?�)}D+�	#B^C����7��RW��a-�Q/��o�}�I0��01��4𾨞�7�[h�EeGFnc�������]��H&(7e���f02Z�Gǳ�������oǎ~��9�L&(F�� ��ro'���Rz��� Vs�c�r�C����P���.ġ�y�W3�>B��0����E}9H�����zգN�q:֒&��-�奮t�k��� ��;���1Wp}�
��B<L�q�D��ٞE�)=0��+3��������(�jX��5�=v����y�������;*ݕ'��Sr��T'WGD5=�E��������[}Ic�U��n6u�����$>S��+pQ�$��;
AB���5˵+��*'����)O����<4�ՐGYȶ+�e�t}�I���$s�H�Ni\�Q���[c$�+�ը!��s�$�Ve�ߙ'S	�������a^�'ye|�ۏ͖�)��[�ǹ����b���ݣ�Χ��^r@�q�+Ō���҇�������:g�Vz5���tJ���g�!Xr�~%ީ�ei9����#��E�gj|;�I��C�x��m�{(�k;u2�J�H��w���]�_G$z��n���T6<���g����o�Z�PH��z�\�-�<�׊�� ������FZE��~:�3��Y�{����Ի���U�F5>��a��p�4N��xQR�L`:6͎� p�y^�4�S�P�{�4��͉�gP��KOY���ɓ*Р�)V�B��+[)�&�IX̴'Sy0�hrR�?�}2\H@���Մ'݃{^���V�O!D�"�E�q0k����K0����\Å���������|����>�H����f��)��Ӧ��D��,�Ԣ�.@��<��6�����o@R:�.��S��� kJT��p&q��;��x[�ΒX��'b%kZ��v���n�%��Uإ�\lA��K��v;ŉg�_�{����8U1�TMN�(�
C{��r�>���a�{��a�l+/m�u�k ��/�.Թ��G��6@4�و%}�k��UX �k�*���η5�	�*���7ԴvXz��6I��m8j�/rBZg�O��|قPZe������~ �YV{_͛�w�v���<Jc��xprw�B����P��_Y��=����4GiC�Ѥ��\Ƨz��-!�M���=9�3��c���p�{��֣!R����d�~��������r��A+��� ��)�?�I ��]�i0�d�D�$�W.�Mk!�x�f�_]N�G5A���oe�R�����J��T�")
�)_��:Y�����8
�?`X�)\w���o��s��7X}]����	5J��d8Q!���XoNώ.��,f���N+��m�}�������}���-��a�"���П�_Z��R�%௫���ѥ��Z�����~4�:�q��@��qS�������8�Ě��c7x���/���(te��e��"����91�4�]�I����kb������Z%W����F+'K @�>UI��1�|Y0��xS�?B��sI'mZW��E�t�)�Q�n���3}-��mm^e,Gv�h�!��a��Yar��x���+�=��e�g<A>��Z"�CQ�6U���8e�-�<�����	P���T�"pI^1A��A�B��:�D"���o��I%�&=*�-��B��Cus�z�mZ���}��������ˏ!���Ԩڢ$|A�8�X��W\�����8��8�E��a�M9_�8	�P�Z����+�[hhQ�:H`h^��0̹���&����3x`í�Q[�=C�u:OF�So �I��q=�#wo�Y]��.�r�p*y�����#�yl4�������țIV�&�Hu�X+�H�z#����
>)�lx����/���nmS�j�ю��ڝ�O����ܮs��;��DEǸ�:J��K��{�D�7I94Lm�`ҭ)��0�UO1~��sx��2��|d�(�i�Џ%�{�ÚG�(�������PM����N(�
<x�m^z�$ x�Ãep��� ����o22Z(��S���tm���˳,�{,|AG�ٖm���+�B(�0�i����v�^��qQ�_+�H�m8p���Z1Q�����Q���
��,��L~8�>b��f'�	�y�^�x��	Tt��ZD��,B��/�K�@`Ym�]/,�n�A�s�y��Kva�*�EO��H^�&�(�CP�R1�I���Ǚ���*��a����BnpF|�g���<k%V�Y���;��tb�HV[Gq"�Hf��R'v�"{��NI-���#�ۭyI)rF��\�ɰ��E��%t�iLˬV"2U�
'�F\�s���8b�,��u躪�q���U�{���U���r���j���i ���:���sQ0���TI�Ug25'��b�T L4[K�?�1TS0�%��&?������x�~��,�I�言;��OB��mW����$]6�8��OMk`�cǝ?@:�ŮNk�p�O��c�}J�˚�y�C���s$�/��^-������&�]��/�z:6�ϛ(���mT��`�qoݣ?&�"���Dh�����d+��f
#L姬�e��3MB��a�}6N4�C�6P����\x��ߨ�Ҏk2�.�u�
�N�Tr%�ز�FY�7���=���E��@���BlM����EZ�ZU� ۇ�����s]��Y���0~h��{�q������^�eW;������y�`��=?�s=o&x�P�i��=��_2Fҥ����OMO~�H���i�f�]�ެ�P����֔z��T|�Z:	-]�&%��خƂ� ��d"oIz�������9��vT��$F�w�=>#��3���vwh����hW��I����í8u����:��F9����BΔ����w�H��!���f���П�)!�:���P8�w�m��2�9���^s�6}��C�>���&b<�YX&�b�G�'�n����Ifx�7��&�o5u3��TF�î@�$h�� �U(\nA;�׿�����60�1
�ֺ�>��AG�R-sk��q�D�U�/��o��Q�Ѝ>P	��FU���kgp�4=4�]�jp����r�@�/�HR���C��q+��$J�)�D�~���/��ѓb3��=;m���a����Fv�(ɠ�AL��퉼kש<r��DVؚ� ^�n�\���Aj�pY���/��W�r�������������ݖ�q�aǜ��: �=�v��e>��U~��O�nzQs���V,�D�𝿣��>;�4Nx$:���w�=�I�k�r�h�u�<c�L��I����q�[o*a=��N�0}��ÒVo���8��:0? Po`�%=�h`�,��k���N�bo�*��-�26���w��%��*�V��^x@]�XdSG��	D;��S�yWJ�n��@�.��
0��Ä�u�f��a�X�*R��q�7hpōe���1�~��L��������&}��~(0��%/$�}��׌�r��Q�Ղ��U�7�P�5��n1,)��T��w=	['���*�*��>PhD�R߫�
@��{�i@��9�Y�}M �E<3�y��=�O�B��u����~��\�N��ks��S�~$���$�����}c�!Ǩ I�쒜�RD��<T}�wBڈd�>{Κ�9�ʥ��za{'����o� z�ˎ�*(0HΤ~C���-��?n�X�b�ת.Յ�����y�7��+�\Bk�"M���I��N��i�'
�P�pf�j�>���=��yW}�x^l`P6=�
9,��xވ���EU��l�AȗOc�b:�#����4#�*�<2�ޡչ�[��Ci�G����<�f ��)N�ϯ�������P+��x�f�u}��k������3$A�1A��	�-]h��-_CI?a�Y�f�G��6´I��Pm�Z�Z��w,�x	���|k/��aN��C����6
�I'��<���b-����Xy�,oo����D�����:YN�)B���Z�+��6S9WA�r4@;I=��\���+�1a����a�2�_x����˦��2�<IyFayp�\��Ro12u�X��i&�`����حT-��x�rK\FIQ�CsEEX ;��O��"�����8�X�gl��q�Z�H���x�Y6S��9��|�$�jƗD�`�1���A~���bK�jD*��߮e"�w< �J4�a�,�s�.���8��O���|vDo�TR����m�)s���,����zC�bݕ�̉��mVg|��س;�h	��3T�"]{>�5�c��!-����!gV�}3m}У*.�'�n��:-F�YXp ���C�Ӧ>u��þ�u�H�}u,޿J!�fztN��j�(��0s<�v9�	��⧞�F��&��@Tc�Roy0�o������.�J�3�M m���+���qD6-d��i=�<��-w��C��S!r��_ΤCL�'�
�7	#��o�CT�����~p��Nh�M}d;�kJ�G�o�1V ��!��J<�̚}~��y��B]��$�zL�Υ����)�ڱ'"[BI�J]����NuM���j�첇h�U�-F�YU>�w���#B��b,Ki�	h��Z�7<C,<ŨH� ��n��RB~X��l�4*�w|LW�+
�gw�g��y���	�}��/E'L�=��%��i
��@H�#�)����x�����'�F{��|?�-炐`�*��k��/�>�t!���&���g��#FjAwngU r��.3-=��-2��v��#f���<]x�-q[��%Ka�@9\g� �Ev�kgY�Oͯ����B��LsJ*��?K�="��5^'�W�=�S�U؟���G����e����=�ӽ.Q~�y>V��!(&U����}�d),��E7�u�cU�1��� I��1/���:c��L��	ds��,yZ��hj�U]�@X'.���UP�̽d;��hS��U�B��LY(�?�[�
[ɻHL�F�����HF	e>µ��@���r�vZ���t��'%lwY+9�dr���
��0E�@U�L��_�M����n$��+�;B�!�`⌚����a~�8�D�$I����F�*�8�؆ymh�rk���iUW�o�TQ'6:��13�{zXم�b�������{f�K{��իˌ�4/�9� #�b9�wei�e�rh�fjq.�:+^�]���iQU>��ks9�y�j8w�7F�iJD|5�l��o�`����o����(}����k����D� b��No��v�,������ᯬ�\Эj3��R	xS���G��R�d���(l�����Ǎ��r�8��3%��-����ڌ��s$ɲ���2�I�OI�k�ս�E�zf� �����ǡ��$�=$*�ń�?�;�~̛�"�$9��_�T͖�r�޷}�霅�
��\��ꔤ�풧/u�u��5�=͔�R�]�$���`m��7����"��k�����F+��t� >�*�Ѱqؒ\�
��EE5��_�����?N�9h��R�S趽 �_�3E��F�*9�#(�&�yq����"��;%`�Z��R�;��0��)��jjܜ���C�I$]�E���P;�?4���Av_+	d�Ըc�Ŭ��l�C
�քn���b������<B�n�CdN�ߎ�.�:_�B8��m�?���ALI2�;20l�D�n��@1?�3�;�-����Ӌf����K�+�/��l�ϻ�_�-���EH�yxl09��i�j2��zP((,6Iܮ�xUqV�Fvؖx��X���Zh�	
H�?XW�=�tku^���:sR�9�"��:Qݡ���#�A��(��D���Ozɘ�6.���L��%�Q�#}�׆�1�"����.9�A_2�X����t�´�T%�4aeLG�+Ľ��P�	�`�$&ۜ�IR�~�&I����#+�q���gX9F���Ћ�T����:��}�e���M�:
C��D�S�~n��Iqc�� gH�B#;v9"�4	�T� $���y˩�����ޜfDEE �Ѯ���#���:��:X�㽴tC-ʧ��
�	�:dk��pV��Y}���|��is�a��^7 �_~(�fCJX�d��j�[�u���fd���LM2�A=4���c�O�t�2���Ɋ�<e�i��w���"L��e���܏-<;s� ���3ԡE��灛�p���IgL�5C�v+��⣶��? &BR�evwPL�n�G(��`�2嗎�=Ț��v�O�H��m��+�����p4 J�`�Ck4�qc��^-�5Α���pT���t-�0fGz�a����r��K�ڀ��Z(t����h,��c�$�ɿ,�$m&����:J���ْk�%m=R�*������W�h�BV�DZ	P0�8,����C���l\�E�������ܙ]S6"��m��V=e0�DQX�ȋA$�,���t:/��{��_w��;k�����%E2"��� �ϴ�Z�)����TBv�c����o��Z�?�J��^j�O����=� ���Q�z��Eto������B�o����x��WͶ)�j�TC�j;���q���[S�?Kh���xE��O�)���o5HJ�9�o˸n���*��Ӑ�;�E�rV��y9N[���βI1}�,����I�n�����&%D�&oV͚>WU:i�.�K�:Cc!K.����VT�Ѻ�W�!e,||��w�" O:n��q�����AL�!@`Q&%��X�vz9ǆ�����O���z'#m��(n6�On迹��t�nq�A����-v���	.��C��Oh�EӚt� ͝�qQL2T%�G��z3�²(��ikIMS �$ҧhk'i�DҋtDk������ �%u��v^�V�"#Z7߶�W�S������d��|��r�H�s������������m������.�6՜�1�4k��yPO�1�n�;�J]"��"ձ�`�zܧ���q:[^��z����i��L�OWR!&��3F�PT�C���9.�����Т�r5|��r,
�8I^�`��3��p*�U���ĕB^?)��{���O.��Y�`�i��o���Ҝ��{�����!�"�x/�U�c��?� ��ޕ��f��Ln����-s.C��ڞ=�=����*rڛ �3r�,�M�q��}��2v,�b�8�; ��b����A ��w^h�l�7���ҽ�r�B�%�m��'%r��T�ڣ�x��Q��e����>Ol�̬źD�
��kޯ5]�QMn:B
����Y)r�4~p��B���Zk;�PE�ع���������HT��[�mل�ec(�f���VZk���D��}��¢|F��ST��eǽi]��ʥ\k�&�����yE$ 6�!-Ǫ;�-G-vӼ��.�._�^�	"���hE|d;��D�U�k���^�8�^���#z.�O�y����]ai�� '�(�U�]!�I�V%~X�\� k���M�G7*�D��|'|��7���M��Cxm+���e���63ki��сb8�	�T%׸4� �_��.����M{��3��J?��쁣7zs/
��Q��ζXK��z��9�[�j�na`���@�����s�E�3d#�L�,��T�l\�:+�9��aR�	�Q�ƺE��D�h1y����)�e Y�����#���frM�U�+��ƾYo��V���ġ�Z�w���ڨg��M�.�{����������;~S�%3z�[���τI�7�K%�c>*��z�O:�@?-y`�bꍊ��ժ���0�X�u�?� >*d�[B��%-ңM��T�uX\�]>@`Wqc�G+�B�^����2�-�X�e���ǈބ�y������O�;�4��U]�8)C"o��\%ʿс��^�>ҝ���C��+C-���,�m�����q�����r +ͨa���7��͋`v�K8����K �x6EW��qC�֢<{�͗�&����`�MX��
��b��_�5�	�L���e�ʠQ&�{��o_X��N�o��>�0a-u&,�jF��1�"����4M2m0��k�����1'XP�EoX��Z|�z�`Y�V���p��e��@rS��ms�z��;OSt���T���d<p�����h����a���/aE�ga��jsԤD3���8���-|� ��՗ "3>4Z�'�����#p�#*v���]tB��n���3�$=/ፙN��b� `���������{kN�����JtF���B?D�5�p�K�v�{���S��~<C+{2�%AJ/��H��K�����T��]�E!�[��=�Z4��\�W�I~EN�]k^�)
`w�a+h\�:��S"�4��l��a=�?x�j�D� Ŵ�^cB��J09$k5��Y�7X���=�F���9}P`\u���Atc�dN+� [ҟK���N��� ���?ɹ�F��!f�q7��� kV��3S�$�a��d0"�J����w$^�Qip*/��� ��.qRbl-��U��ӏiOF�K��Z��kl��m.��i��Yw4*���e�[�ΰ�U�nj--إ���t������3�N1�S���l����C�����
�a&���B��k�8٤c.�L�D\4�������Y�R
�r���<r��ES�1���L,������H� �E��٨��h�b���1��傈j��j� ��:��hs�=�(�����I8��E`���D=1`�d�T4=����s�Bc�{��o�r���8-/Fd�1�ƪq~#�RR�՚����}Fc2���U`uϛ�������ڔ0���w5!�B㚬�*���!(����^�=�}xʾ�����W�W�B�2�w�u��=���P�?e��{�i��W�f�Z��JaQ��x��m�;P=�����5��g��3E���`v����J@l�xP$��[Y�s��~W(��k��~������AiٯL�â��W�L."��.7BP�e'`�4��E|��r�3���Ҿ�������+��8�F!�?�7�A�\ԛ�w��S�ު���tIĨ�G�"OY�!�#s�o�w��#'7r�$E���6eP�"�?L��M��<�.HԵ�7�m�Xj��w$��z�͋9jr`~r]�� ŋ2� ��
�L$�@V�r�5�9i�O�8v.	���օ+$������̖�A��r���"�b�Ʒ�K��7eV��74N{&=���x��� ���\j%��#�*��tҍ<�K��3�<�#��U�J�-"��hA�p��ى.F�gQ=LiN�������w :�sr����Nd��&�;�.�A�]{v4�������?�ɏx� |I��S�{��Z�#E7SM�},��XQ�R1Ѻ\�.�Ꮩ����� ��8b"�)�j.�T�{?!-4�S��͵X�?4���K����G3z��MY�tc̉��L�U�h1-m���r�+Y�gəI��&s��r�����U���љ�1��d�X�0��s�ZX9����xT+}�\^TxbB~W z��J	��=|�c��tfۭ}�B�(%��_��zܾ4��G�3Z`=���O�Z$�8V��7j��P�m5��c,���U� ��,#aR*�]�J��DV���!DQ\�^p�����9cw>���Xi���ܡq��S��|��+��xJ��~��̓�+j.$xN� ����;}�O�ߙ�Zj���uN��}h2a��	��P6IZ5)��V>Љ�\Y`4�F�%�*��!xT�7��k��y: #��1=�&��+�3Fډ�p6��J�V�/��@����x���-y柀E�}KNfֱ����*�t�XĂ�V-Ҧ:���M��\8�=OrN>�XZ{���KQ�g�!b��eZ4K��`^r����Q�!�~8e'�!��,u�!8�_t�Z(G��&���,���KT�{5�S��sn�U���α��U��X-���Y��8���QV��|���#Q�lJ�Ɉv��;t?���?���:8�s�ҁ�u�0H�k�:�eIg�W�	�H$zp.�7Gp!f����tkN�����V�á�F�4|]�C��:Ġ$�k |0/&����)l��@�.�䕲�ru���t���|R�* �Ȯ��ߌ�&o�+�R��M�w���:�5:�Y�C�uԞ��gy�����s��N��͐�ӗ�zH�I����i�5]�]���3�����sC�f�%��}�)�K> �C�1��j��mo����`���{vߢ�����c��p�Ei
�*���
ͤF��V�H���*��*�t��;�G�h��JC��c������ \h����̭�7����^�����O$R��,M�G��m�8&&�5!��W)Y��(����%s��:"~�2"��'i��_4(���M�2x3��<�wPgPg�oP\8���/0����<%eb�Kw���p��٭`�~�2߱?C�*Y��x�B��	$���8���l�}l#����<$l�E�qYc]x�4]s���5/��,3�_�IX�e)	>��c�[�0uA�d�]�@�=��[�N��'7b�V�R�$������c����t�� Ս\Ǥ��VrR��%��9�~S��{DQ�IF(��M��XEv����o�DR&G{F�f�N�Iv�W*kL�<�>�B�+C��&m?�c����/Ė������f�	h3��r��Ȝ��
P��:� >]����Q�K#��mW����/o�]�퉒��Q��!��>���tJ�.�O�����xg�,���ϫ�~��V�W�t����Y��[�@�1KG���Z��cm�h*=�T&[�����*��3f�� _�=<�p����/�-+#�P��k��e,�����BX}�x�UԼ��go!��\��1#���̟���@�U��5y�n�T�����+js*�#R�΍Èmb|������pAR��>d� ����,�fs�N��E�K\�v<N��$m��1�N� ���tȈ��&sT�L�"A��g`C��v:��Z�1���k�_�lR��7<q]�EPK`u�w� v�9�g��y$���p��DM�e�}��\9W4���`�s���%�u���$۰'���\�kh�!~�ҿ�M��)��%��n8��	y���)4%�����7YJ�{) �LT��=���c����?^4�Љ"�"V�b�gd��*sj���|f�d�L���$�%��n�_�>�S5��������Be�d22���rrփ"��[&�p��<u�3VZT��1��L��S���hQ�-�=հ�ܶ�QC^s�/,�����ID����W�C'��V����n���ͻ�]��WkSӷ�}�cm�(q�բo��KcsƔ�5��@.ZE�[�1_�]/�"�EM����,k�)Ⱥ)� ��(׆�Ʒ�g���6�N&Thp7�||<@���+�&�~�x
H7*�"Η_(V���Zh�j+F^Ӟ��»��Y��+e�;C���}3r)r�&2�{�R"�F���o��{�u���x�~��7^O��������?��10_y0(Ej����'���wP@���̛�n�F�N�
0�#��UL,�5'i�i��}&�r�U?�T9�3�ͼ���G1�fD��Z3f�<��� /��0w;v�I�5a���y\��n��@�:��*H��1�+Hv���Z�DJ4h�#g�h�,�	u%���z���5�/�v>4A��S�B<����
��j+]׀6�a�`>�[ǫ�t��E)������qM�p"G�/���8P4�L1��@nx�m�2�|���l�5�~��T;HT� ���핈�.����nl�����t=j=r������b�Tc@�"���AɅa��#�t�B;��|�2<|��2��N��J��gS?H�w2ʐ=�m��L9tP�U>v�k#b06Qya���������qQ�C����ڲ���� ��A5���{���4K��:����IJ� ��~w��p!��vF�,���* `�U��8W�(�䖧��ca����h�պ��i=��_v���7�_Է6�\�;�C��.��v�+1���L4;ƫ`��.$P�eY�6+�ڦN4n�,�8��5;xM�8�<F����'D��Dܞ�O�r�T�f��=#~�/������x9;"t\�GԴf��q�|��M�Z����+N�:���>8��;��R�Wg��*U����r�>�w�2!*|j���u�^�_L���s�y~µ:���@�ʵ�0�.�Tڤ���sF�EO1P��Y���jv��O�@b�\���=��
�g�[����p����Z�4��P�vK� y���)$���+i�PVL!8J�e&�r!?�\���3�qӨ������ُ�th칂��=-Ѓ��@Ka#O_k%Bl���\{�վgDb�f2ّ�O���Z��O����(��t��lE�Э5���J��:=�����<��\�%a�AOi��47rw���"�6��E_�I|OJ�\ԢD`I���7��qݮ�JΙ+Gݠ��|��ޥ4�NT4����3>��0�ȅ���MOw�0\�ؗv,�	'H ��"�����!]#pб!�"�_{�MX�k��,>�ׇ߄{TZ��5[ ��w��qe�^D��[�D-x�}���#jq1S�,H4X�
��l�j��s
KbGE�E���<�.djN�Z�ʎ������f8$�I� ��3N�.4�nr���
�E�x)�d<�<�S�+�]�t�>��B�ie,�V#���O��s�m�$�Mz��.t������+.��apDc[��Pp!����W8\�9��h�M���E]�.a`T��C�|�������lJ">��w�΍ �E���;�l	�a��v�=ߜ�*ѳ���C.�e�\�Nng��%��g��*Og���r��^��	t�!�I�%|:��	������u�2OK<
�\;],�"�������͇�C��dge��������t^L�4R�)��d�V�Ir{� �o:�e��au��2APS�X���
�9�nZ*l� y�<��@��.�Z�� ��9gj�x��N�jd�� 4�N4�; 4jqK�JA�4���CW���/v~�xC���dG?Kxv>M�B����=e�'V|���^tT�8��Wu��9!���r���oE��X�R����H�]����l���/\��0$�/lBa`%����)�͡�/uL��ݔ2�N�(˧�{�l�j�m3�� �H�u7��NF��;͜p��Y�?�A��f�V\�\w��g�i�wd����uT~yG`$
��N����T�����ZS$riQ�Ɯd�`ƴ|�ҡ�,ފ:��х���D&݋y���r�}+qZ���fz�'�T,�p@�֛3�"9�B�Efl&'�J�[":��������%�>�7:h�S�t�t�~��b΃��W}V����$Le�BM�ԪA��y,yt)�]�g���B����5�����F�G�f�{k�3��'�%@_�d_�͜������m<�����NK�	�s��d�m�F�_9��A&�a���6�%O٠�ȑ���|�o�t;�`#Mbt�w���͆���%���O����N�HN��o �� N���;��tg�]557Lp_�9��	�!�`M���-	�ݯ��[i�mf�����<��!c��o(���c<��̾�z�	������A������T��-T�hM�ɐ���yT���F'H�?+T0��Q��9����ӉQC1��)`�3�@�{6� ���t����RC��'�k�F1<kG�:�i���B�9�E�s %S�	�R	��fTxQ�[�{��;v��:�c\�J�Q1T �RtNE.MS�+���䣯ε�tu�H�Up	Ět�I�K#"#������ΐoDHoпGH<�˕���斁ܧ/VK�b|i��h߲4������� o�Aخ��De �n�d�S���F��Z�M�8j��lc�n[D� �(�ѵ�^���m2[��K0�A�غk��sh�
�ى �|��yK��\�I��0�W�AJV��+^G�5۷�)PEu@,�j�ӈ9�e��4�Hr8?F�C����,w ��,��M$���C meQ�ҭ��s���a�<*��V�S"�����e��Y��e*\	:2\�[�M� �$)�Uě�<��z��7���OY�~����#a� �>�\f�t6Q 1z�����	� �M���J���h����cjo|5_�*W��?�[t^�d�@�$�	@�F:r��y�h<wG��5,6�A�L���i���O�O\��$�ŭ�`�
�T����B���2M�N�5���E��>7j=�Y�B*74� ����zӽz��&�K������EHOEzY��ٙ_s��R���;瓃�D+�ͻ]~�zI!u���s%%�j�K��#�ơ�Rڙ5��Ʉ��ҐR��=E^��5.��Q�&��Zt��7��? &?`x��+/LU�VmB��2�c�7z�\�W�ؓϢ�~���H��ǿ�w�q�Kg(ϒ�7���F��y���ʇ��d���P�	��iϭ�:�`�2�c>JU�y[�2�5���K߿!��˫�q�,v�P�0���X��cqP�Ǥ0&
��L�Z$���3�M��K�s�������ɢu�Z�S4�j{	�f���CPƍ
{��#=��wݠ�ޤ��:�\Y���P��(N@�SNwN��!�L�%��V3�P�*��8����)�:�s'gx�dDf{�$���0X���gP���1h}�.Ϗ�D��E(nU�-kQ]�	e��"�]�W�@��ES�"�eQ�8Nc���\Y1�k�)��nq:Lo���>oDS����f^}�F�坂��������S��0�X�F��)\(&�۾�{��:�pJ�ř�m�Jp��	bWz�AX๊#�7��>@p��C����9��.�dڦwx5_�tv��Wr@Zq�/*���q��ڵ�q+�:}��A���Is��ӷ#yA/�WA����?���������:H-�3�[��hy��6���(�t�{Vבj�6OUY�֟�ǥ9��&
�V:z�^��@oה�Q�xT��e��}Z�z�%iO�b�H"/4���9��/ݏ[�˸�:M�������ɤ p���k����>���:�u��=�t�}�e5g�:��A�ގKKt*s!�;A�OhK#;�YDOԦ�·
D//rËK����ܗ������u,�P��a�R�H��X}\2�N��� i�c<c����"�إ['7�|��J�7О�����.i��}��5[���s�(�L *�G�k6���Ԫ�m�c��Y,ψ�k|FD�,Z�ߚE��FFR+��@�y�4�:���bN�}]��mK�vQ�����\��]K�7�_O����j�>�p�6%�����6�P��a���`�t�1��-��l^�j��?�.kO�D� �ܯEL�gA��x����*��)$JU	qЮɂ����r
~h�6�W���2-��C��=�ے��9�$	����Hjl�Jb��=�wRla�H%�}�e�֚�o�!I��|�┮��)աX�^A �CC�"��O�oͱB�"W�mL����?:Q#���F�
�@j�L�f΍c����μ+4y�y�^e�ꗞ�6ՄQ��h{�*sn<V?tM�^0 ��|�v���H G�ًg�xM�*�8[��Ή۴n��%��d����4���;��U �m&��J�|q{Qy�)R���`YT�|�9��m߭[꺢��q�%f�R�iTh�w��D~��T���TT��x�z��ٳ� ��	\�3)#�Dq&Ѧ��~�:�1A(�0�0/~'d�󣚻w����$�3�1,��K�9ݽ���#lۘ#��y�Q+b�ى����L�#����a֠*i�o~;RA�gu?R;�e<��b�Rs#c���Q���s54�-�VP��
B�P#�]K>�t����+#��S���*��`콪mT��{�fﲵj�J��ɛ%�/_�ĪF
�����_T�P�S�؉=�c�/u�DIadc-�������Y��j�Z1��_�C	��IT�1��);�M��sS'x�d�*�ƶ~�yY3]�(�+),,�x��[!�o�����Fk;��r߽L�����E���'�_����j��-4�>��@�-zm�{� ���������/��يM�	�h��e�Ǧ:O�}ߜ��6o�͐�nM+u�^:�%^�_�$��fx�	�-��M\��7Z���+��
2�ahS���Qu|p�S!�+V����{S	'I��Բ܍\��b(�\tW��H�
�Q�� �O+y�و[j�6샦�g�%)?�jANP�o!	��B��F$�N����8e�|�\܃�/�Xf0Q�$�S�PS�/��k��e��#lA�i:����N�C�S'���7DU��d��O�(/��%B*˧�~\K�Q��x5Н�J��c[���OF.�Z�@�u0`$��+΋gx���]f=Xr��[�- ������D;-�i;R;�-yNd>���s�
xx���z�w��+٘&59��E
N��F�B����1F�l�̈́Q#>�����Ԯ���KY*|���k�-�/�/W'�.���>��D������cҞ7�:1��U\_ҡ:��G8�(*uΚÎ#v��A���r�U�������t:���2Ȑ&w����#�5�4|jrz�K�'�U�qd�K���I��E��M� C]j�di����A���lM;�ZU'�Ɖ���2������r�֫�)����8xr�k�7�i�8f*���f��t�\�(��c��dԉ���+�����������m���6���X�Y�uxi���r�uvC�S�MR6'|R�B0��1�e��W��b��~��>�&6#�b�ESvG)��f/�q::O���Ŷ^,,af�;�-=џ�`�0ȫ����LAN{>�,�z-F|.�6��MG����H���:�&󺹻��jhaU����z4G�����,���>�툛�r��9��l^��'1�(*A��B�n�S��O�Y�n�cYNh�y�r�r9�|%����L.a�i��!$�?�0	ҿZK��M���+��H���0�1�����W*_�2�����Ӆ��Y�9�F�O��|�U�,���r{�k��eE�=��slo.���6�37O:R�1�����$�\�!d�PU��n��aPؒ;Py�L�֩�}�M��4�?�/>���V�Ls5��5~�x�8;��t(Q�s����^�8@�ͽT]��EEK.�O��H���	=d����9��p����|���
	�1h3�J�PY�Gt)6[���N.��;����n�,b���B���Ύ���Anz�h�+IR~��)���G@�]���:o�-��5Mw�Ƒ0�Ǚ�6>%���� t6Z��#j�B�!J��-��C�&W%H=�Dl�B(��Qt�>9k�m��3��o�z�+�#^r��-ք8�r�߽��p#���[8�oB���=Pe�3�ӕ��=fYY����RQn�8����}���t�sK�K�M���fo�&����~e6_f珙�}��(��l��f�o%`��֌���x ��d�v��)�K^_��zMt�?ڪC��s>���a�5ٮfӍx��v�
��Zv��yŃD�^�B��`�ޢ��P�k��h�s�WRixhͮ�I�-��pJ]��7PBQƕq��'��Q�����"�<%���#�1<���^����Ag˟��xJ6�����>Մ��
�o`Q���Қݾ��5_p�6�l�,����I�#��HO`ĝh�dR�3��Bc��L�n�3e�+y�R�s6�ݳ�����=�4�Sg�¶q�	9��>�[�R�N��0��=�q!�C+S����C."�A�=L��
��	�_C2.�FK�qm�L��!�WJF����7�$}�G���g.�Ċ/�$	��?���:�.�����˸�N�7�b2��a��ql��/�|qnD����ͺ�e|Uj��z���}%:�C�1
g���o��J"j_�^��tq�f`TpY���[ՌD[[i�R�g��m����������$)D������y`����q�1����������'���ϼ�	^��%J�ô��鸆 x��s��~$�j�-ևmlG���hq+�9\g�F�fi�܅7�\OY/R�O������6�*���@/��2�{)�ODV��>.�s%L��@+;��O�"��O=�Ly��~���#k@��B±烍u���ղ�O�7��0}]te�N��D>a����ځ	�����N�)��4<e0V�mJ<4b�'�M<��V�]��V�|)�黟~�nx	8���*Bl��2y�o�:����bG����r
�:�<K��YX�`���(�Q�>7��ٯ��v�7>�o�hK����FJQ��ƍ��6��MF�<.����T:��h��,���q��2�������Ǩ� '��/��1A\��K	�Ōؿ5밷�N��]�Lw���SS}��y9�[��>ǲ�"��A�Y\x�Yi�)��Ι���k��M��,�-f����!ՠ
ʾ�m���͆:	��;�ݞ�N��(�eM7 ���u��˙:]���2�EGP�G#R��X�.vj�ۘ����&���|�e�)��E]c�P�棙k�߹�8�y提�s�T?�p#�!���A��>�G1����.[�2���a6��e�GZ��"sWf���J0s�@����+��ޔ�<�'O2P��E���+C, ��W�;�𴧝<|�~����9`T�3��(g��@��g*�Ct �AmB﮳���`��J��%�;D�-;��A��+�[�I=��8���Q��ns5Y�/$j�nT�df�Ax�9(����)��
��8ol'
G�Rw�6�k�ݐ�O��γ��;9!,;u�%�����p���C�b��pC��o�h��v����L!��6S_L���/^�ح�,�zmHק��Z��x��j�ҩgg��a8�.�oST�xč+�py�|��Ӗ�*����y��6c6��CA���>̰��&3���Y���ۺ�!@��_鄅���c�'�|CU`]=�vb+���ǰ'�l��G��_���7�l���e���9�<%��[�}�=�X��x|��IcJlk,���[�1R6� K�"S���Y:����f�~�hRv��Z0ĉ�̱���|������K�T$�P�r����؟%b��4[W/@l�����������
s��\-�N!�m%���eB�{H���<��7�J��G��m^�Bӭ4������N�ΙYÆ�_�X����a=�r���d�$��'����d�*�L��4�qT��b��:�}d�ޤ���˺)}�l�[[ةt^R���O2.�ђ
f��X�4�*}}�tN���x�� ��>�-,T�y��0�_ȑ�x"k��bUc�A�z��בx��'"a#����W��׎u\}����Ĝķ�Rؾ�\6�������~�c�E�\��Έ�`Y������1M4&O��G]��]�a_%U��1
�dJ'[���	[@������n�Ҙ.�7���[僱��Y���|��k�f6��I1���F)d�OY�a��`]�F�k(w�N\��X[�o�8�3�c��B���c�#�Q�7��p�rǌ��������}$Oj�p�P�r�X�3���Vb?J���~�����2�0��o��ײu�WRq<�~nN@T��=�Q��^��õ�=������n���P?{�6�N֖5�����r�����y��3��'G�Vz��z��r�o6��?���S9�k�GC����x�T��.��F^�r���t<f�����{�b�j������jTHZhc����?#�CF{xq�"�>����z��s���s�����*������p1_����3�Ì%B~�9�T����{+��2Oc�V�~�mg���:P�2*P Ap�����L���]�7�a��hR�W�y���,
����X��?�����	����_�<��Ʒ|�wz[p�ww��zn�(w�PG��>n��( ��`�R����u����e��:��Q8��|8_��?U40�/�Cv��>�O��J��/���$ .��h��c��2 KgS9)*��#y�b�+�b������%ܮ"��%w�d�;�Kc�s�8T�6_mCđ)��L�B��为P(5WƜ��'o�����wG��)�t銈��ykM�� ݸ�-�����s��N`�j�&2�T��D1L��&o�M+�TR���?t=
ty9������<��N�x.H�)Jԍ� Ck��J�m�ô�N;��U(蛁3j�ֹ5=��6\�3|o�ͱp�h� ���*ρ^��w�����>��=�a/=��� 8�]�J���o����f��|�fQ1A��j�?�!J�����k�uU@L��G�*F`^��=�ȿ�u�'����{�T�.V��7��$��υ��/@0�lD�K�-7�ӝ�J!e�,�T$1PNJOYB�d�\��6���|�sQ�5t�__UM�x��!ef��~��E��k�߷���
�B�Ȑ�Kegŗ��_�UԒ�w�=/�\��"!��
����L�m��䬩���J۰e>��APo���T�Lm~5i�hP�~��gc�+����5P"Xi����Fk�k�r����}�h�!�^R����U���������Х3����vu���wTM�CЎ��?�ΰ"�ynGl�V%,�
�|�,*豓�k+P�F���1�8�/v�`�gO�cWe`ysY�s������.!�z�vZ��q9�������YǬ�����"���y9��t�������e�L�UO��'F�n�k�`��F�9�<.�2"=3Qkz���EBD4l�\���WO�xT_������s�U���;�"�F���y �\@�c_T[��