-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
ouoRNUlzGa3PGOXz6U0cWByh1heFvz6cGTzhSnXBb88Pw3dMgIZSZ1Ufdz9K3OVGkbFYX7lWdoFI
NwuQETp3Id3BtwPCs7k2upV1ySiott+H0z//Fxv7XgsvJKBi1Jlnmf5F9hRlDk6/UWiYx/owkAgY
F0tRArLu2wRm/saPu/tiG/Xu5mALKpyeP75x1EnDPfU8pLa6/OVEn3VVrBOBWzAh7j0rDtmfgTKw
evuWbatsFBoV9WDgilFw8wvNsxgaD9QltZ5T5yydE0y5S0mDzuQfnx+ureNBHcXfcHSl5o2xyDUc
H+LwznEhh92vADPoak6KiTWJors59qD2jICkUQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 12400)
`protect data_block
vKBrHdvxVRawq+wQMhu/qjyqNbbf8T9YyMrlD4P1IBofYypR9sJvrUgGutmfYUlquqUAo6yr8Ngk
dF/0G/SHreSjxseas7sjxww/IfAr6oymYz/NIHJ8bjclNCTf3vJuLg++mhSBsKsufl1m9/z4J5CI
9L+IspB1DICIlRW7D/OQKHdQympL0a7BaUImHZ/AGqddlXAQeecyluLnQZXKneW0PYggOiKoxfsS
IEuKGdlXGgO/g2FXq+lNYpCwyvUZ+zIbppN/5hsgh6xrKrvd2Ao58QB1WGoEzz9o4CyN5Pcb5IRb
kf8KiPSns2/2c8Bu4EfC2g+XKALiafgdhg9oxXBmRSyM91ErCpB7gvgOnJ3jRk9Hvsg8GMa+XrsS
cN+HomxFi+aZy1YuS4RQpNrB8t4Jjjxq84AmKmrrb5rKJFhXdKJAci1JVVLpDP8ujfLoF3J0n3n8
BoyCPqztHWuxnWBjd2haU5G6JMc1YU/Iyj7347+4hdVsiB95ZS0HVXT98aIMz5582kBr0thHHTKP
KRD4Jb8S3+gFSaNtq3r3DnHRk//vyNtJkyiCx9/6/g3xuD+pnG3NHmKsnCg01wxrySTLaQn+3ROs
L6g4VE30r7a7HprXcqbficirnGFueiWhKDJi4xrq6gvQ3TpZTf9XG2W64UuHquaKjxpng5k5EFwD
69/y2ka+r99M0uKSxw4ULxpTBiWOewyLmz45lr8YdmdH1/RAw+8QeKEDP4JSeV0PS0v0122LPLBA
1ey1GTPb0cAhqy8pYjDw71BvuWs9/5/HrmPOV8b+d+rXpXt0SY9c0Zs7uOKC+s6RqvNwWnO0/AHe
wD6AkiEAhCXS1aBh1jE5yF0HH8GtBSkhQd1MqYNsCPCgrV+knZpfdtgHPuwqOHQopOiiVLxTJXTW
tjWXOfkitrcDShtsGoGo3OzqGseu3CGl37hVB6OVl2LaaewmV9yXH4Jlwibo2fLDGDynWDe7wVZ5
timClBXW4vF80KPfLMz18Ugqqmw+jbC3ie7qvPBboVnDLP1jKocl8Kqk8+dzKFyPIgWHZCJRpgA9
oaUWq/LHefLLQWqXfpC2p24PPDLmzihLS9Z81Q89Bve5qTYqKEorov0h/sPBFcXRqBdy8HJblVS1
BrMLLp8xbdiMD9iFCo61C03rkxM9iwfxgObVJs4WUy5EuG8RiqnT6EYeb3hiZ7g2MjSpdAQKM4v2
a7OGqYy91ENZhdM3UikDXLU/Dwh5TOLOTCHfuDnbvrDsRatzoAAoRESjHHErhzv9TfQBYZ7bp3As
LhRopFrbijazOB+nLCBJxFBbIgMFJ+tkOlwewn+1V/L5zofsrpxtlcnvNd6AsB3cCB/RRGmXtdtd
GGyu28QZopvfCa4b4mkoTtMoQI3zUW2WEatrcT1ANoiPQXUgNhyC64XxsKioZ5vJyZDVX8A1b8Mr
TdHkFej+uY8Rv0oHSP00lULMKdSGHwLlAtAP8PobiZ2eYizt1MPkrzAT3a0w26vzzgB2BgbuYboM
lm/VyLuc1LnEqPolbN9FvxQwz2cTxucQrm//BnIGcrpxEL3cz+zlzgen2N0Wkq/Cy6xF/9ST+heB
HQwExiphA3fT7LNSlF6cyOEfqqojbY2BxYnvACJ4NlPyQyWotec7nOzf/czNhgTipYwkGtxTZHR0
NqQci/fsJ+NiacOYYiqBMrG8LdyXggUehuQQN3WTKZKf183VZEdjEn7Jy06tCmgLkdpFu8NgTJYI
1asSRhb6mELLrocCGwpZz5uma9iHs7lDPOR8mtO2n5a4uMk8uMnsxKzxzPoNfZ8LuWCEwxEq4bzR
XPv4+xkCSimDyUHLAfe5GK58Nj/CIPYIqhT7HIJ1qS7owOgA3jqq3BwWXjymbznwwm+AjI/cy83m
WQPEK5oZXVvwAYvMlm+OnGLXIOsNGQgBxFqozi8/bt0eZ518Owbov8+7YlQibRfjGMw3i4OFnZqg
zuOvhISEWOSGDXB4uPr5zMMeDU9Id9B5YYbVyn1CKKqbiiheNDaivOCUfbOyU5BqyfuXBuzZVXyB
yLvtYpKEOIEETOdJE49EB+jB4wGGUnws4heS7gPIKMaFCakuhf2+bTCwANkfxmgTfyni4BgIEts5
W9aFGkSYTU66sCC0xH3JdVz8gOmSctoggJQYqaY/XxlNO9KoVcZ+NAsExa39CgUEt5kIt29eX45+
vinqjT3P/U5jEcHpW1Mwgmga4W6VoWEGYYxy+p3YT3K3cmH4xX/ujEsgVJ/T76gOQZJ5tc6Ca/Bi
d2smBgiPvQJeumW0C+hbTOk5vIz4OnPV9VUVLuRiPce3clYg+5yFmPzBLgfYzNTftbZ5t9K9IpXw
IY9wsB/7En+bjAuvt3cHYb7ObAwQlRDGebC5He4J7dUumQAAKn2F2nGqCzTdA2BQFQ/RE3IfVYLA
b+IZgv3h1p8yjz0AwtBnWADFYmyZRp5A9kevEN2csDxJfRlqd7VNA9KRN5yW2wjS7HbWHF6xjZxI
UajAF03Jb+eA1Ap5Ju2sHgZ+6Wlblvm81aOI0ntqionRhhp2advsvtro5n664yMheFvL8Ze79v15
I/UWODt7A8AtUol0oqpTWmhVj3dNkwpphA6TO3xGPXfA6cxotTIkWLUNeyd2rdmtGRZNJiVQB3fL
JDqa+3y9rtrsq7MIH1HYpt/ak6X013OjWXRVc8MVcb7izFdww1TTKTc10DGC1Wx5AmTf5EK2KHJP
uvZ4jbHqMVEaUi0MWZHhWT5osJ6Z7xFC1BQJc4kVjHzdCr8YzqaO+WM7caLYT/NPTQ3DMznI8BVu
/DkhILD6bnIwgyn/0pQFUrQ3K+Hu62z6pjXRgiIpTw3mdsvG5fdwybfgfb6vNF318wgs29ffspQy
T2bzqCO5M47ZQw2dzUBBwBWq9ItDnHNbE2P0VQncf8HxNw96csBemXL4cNlOUx8221tp/vl6dZRW
+g5Dgidn3fIFeyYVkTt3kaZ3OVs5wUhO7V3VSeRJkZ8l31OrF9+A73YcIYyv4QkenIgmWsh6SjDY
Vt9mCtEnrBpApTlXmbakFYvqHpJUXe2G/SCF+i/91uZttezTaJ/Z4k80o51PYBniO3KzVbF+DR5I
OikWDGvxNadSjCLTjlTJFWN0nwFLDLpuA5UF4oYygmxko5dZctLjUUA1/cw+mIvHP9dXMT6G1QmV
wqR3MXmoJwnAowxLEI/wyaPHrp/wj1xN75DWHeWdRp/bjuLpGXvr2WJaH04xrgfeW2IK1bWODyj9
1xJr+XKm8FvSlYbeM30zvhsCeCShe31C6cAEoWYCmYj/n4/I3rjAgzl5BuHSC1rOClGyqyB3j4Un
YINRyRMhQYxjPlJmUI7QCMjm2sD13XvR/Fd7o4vZi6B8Ys/841JOTv1aX3Tlf5P0fJ77LbgpxsfW
nLBtQrehGEo+uUdIG7Qypw7NywxoYhwsoBmO9Y076B/3jLHDrnhMfKCsge5i5IJrrEdD6dqzhc75
BRgUyU8OYMZ3QnCJyTsJJ7q1Me0lhvh8oawss2ArfVfbPu+eDwqlLNcD2PK4buzSAg24/nHUr1kp
fUPcGNO0iOkxrHIQfdDdzi9II4sMydOwF7MoSdCRhC0TTtz1dyuAI8c44xt1hSXv9NygMpFZiteu
tpz3X5M3Ovte/QbqszWFPJ9x02IcH8iLDe4W1rBfnifrKHXHfdgDz8MEo+O5tTvSmJYGuQj7O4z2
f8PUKplVECy4iCuRnePXrrNNgsMnxPOGBahIkFUY9epwPi/rkzThwQxsqOJPiyuI6RMQunOY4iHo
dH/GRFQHLAaPT3J059r3oEnhsg5DyxoLTx0ngcE0pVQnL8EXMNEvOC0yMkiDeppevyFGmBV9hNOW
Q3QTGdHCnIsLmxpT51twnWg4bdMrt35LPUorXwNkaByCkBuJMJBedgVp8h49o6EA3hyKnZmnzlMN
SeUiLRlpio9DJ2d9ESaY1pTjbgvdOQXdCQnUqdSODXlvsqREeDjayLnjrqKnHV+Q1euZ9R2PFSnV
tZtBzheGdKBMxDqqG2fYHeuDGAjqXT3H5x3OIcafphu9qWhod9VQTiz0BjiZF+TJoYsizT43osJw
ij7SWEZ0AEam8Nnlu6sorefZs3mDGLuBedH3FvN/WsgEgFb52bbuKYnlFM6qQ6cB01QbTP+tjESW
RuDmFT/uh9l0eZ3fpNA9GvILfiUlyGaKND5NPmtIUSyTwGNhRka36HiojcOq3ck5Pi5tt/6ITmCM
jsUiSMF3AL8SI2QpEnanDD8hnsZB/+PQtZmObPnIb2EGauuNeu61GB0+PQtuArecxB8MbHT8C8RS
newEzFaVyvRl5AbT9iu3RbQRJeYIwbaArBcwql8L4fMaEIDTERYGB0XAOTf/h2E0crxO0dF/9ARX
m4HMEQGBbazl1VDNBZh8z5ns5BgnB2ek8SbrQUhzG+nQW7aKkqQnVBJ2m6fRLeNXOJK4+r1vqg4V
HQ/+sXVK7jjxYPROdq9Aala5J0RS+thykynti7da/MzfcLXcqbDQDZOzkIxEgyznSF8uRH61oT1j
oM/wx2Px+kfrtnPBn7Crw6LK1v5kmX2voLEJcK11cOK2FIa4/8yKF+rf1+EGaFEh2RtHEycfcWVB
NrmjTuX3Zyz6lRYM0F8HuK3egpEZwTX+z+XeFuH+2XWHBfeEC/tsVVtVQJ7df8bPdqFhnBEebLrz
e8zob2zbzsWyr7KbSf83QWKaueaqkCjTOGsI2yhghFNiFMqo8F3uhhwbEN7AdXD1haZqj/m6gC2B
jJNUU7OdYy2KKAwMpIJFa1RSvhUrqIdGv+/7QwUS+HW8rQFqIkIH7u9fWj6BzkLoPH/2YvmbjQy+
iKE4mM1mYLl7L4+muvcJ5gMSF9tAbWQjIYhDEThJ7WhhyM97p8+exWIOa9a/FlQJTrmUZNPV7lzb
tYNTfYoBuoEtljMZmLEUlPRhTYDxOry0qbC+zYD3TMmUBfT1U2WCe4rq9F54y7ibFY2000BIEqCt
7yjIjOMV+Km3yVVeTH2p2yViyng6KoCZ2UkrrKTu1jlBSW09nP3X2ScNJ1/q1phm3hwupwnliBLt
Z2ENzjO0mGzShxEBMJ1i7nH8zBOadl2elt5ee36WuE6boqJJTAjAs5zXFtVB6mDaJU86q+v1hyLZ
1ThFSaBrwzacucSVxE6j9Po9Iytt4MP+ai7cm1vl4an+T/2uTBx7J+cXpe+AMzZMkyoecqus8C5s
uUc+YXm3Hlpgewl1qeaqRCfXAUOxmvCAyGWghLTAWwK1A5W2D3bBYDaF+99SFRoLtTIJ+a7fafba
/2mkc3P9T6gf4s6Yn/rKVkkv2segqS7E/EH4GBlUaLUOYs32J2XPv2D/U8TdPpzb/VWQ9xUb3uX7
4aiTLXt1zt2EQ0k5y02fYht83TqBNf5OT6bpfsAyRscnH2qyJZrbdCpM1iAB+EDfZp+OiOkb7N7Y
tcuKdlVC/w1ID/15dnpmchz7vl6noibIxHFBVVTx0yYTpsCYVjOzzbtTZadjSa56Vnkaf6bzAdSs
BXiDcz3UjcPST/ivoq/Jep/JyVsxQE4FPDITGNt+xstdfDWAqjC+M3m5ZJZzfEE/5UIBGRYOg07A
77bhIanV2FJPjvWgNhZPpB9tRG52W2FEqke6ly9A/ixTzRETTqdf7yey8DvmWIfbcz+Iyd7dGqeg
rwDE1SGJVXSdseQVZLdBfWmuo7EUALA1oOsgf8fZTAw/YeM831HoR+u1RBs2WgyuDk+wUOuLVNzc
4/ie/bWxu/b45F1giCXnS/js0ekWEg5XVBJkpuZ2OMwIoVxc3L2MxtpFMb7pl4ie3ydA1uxIv+AJ
8XesvKp8MSX+WHFOpN005+Zia4nORcYTBHpFhX7iHgBzaXCZsD3QBuEfnu8NdF1HEyl0X1OSc8/o
2u/A0Oxq0S44W8BmCQaRuSO59iW5RFjrebAzICNaZIki7klGZXoFHenNvaGDYPF2rmNAS9ke0zLM
UsaTEqVStVuoLjoqSShTAQT2boOBY8W/jKJzcnmzDm9hTbHe0rH5QvPmTvuy4cAYml66+Y2mNqFs
bPT2nQFssWjox0H9NP0TodbqSh3DbgZr1lI9t1X61FjMBmlZW0UfrcMlfhQHtlpQC8iwuYBCKTg0
Ysw2aZ3kRllbGYshyRxHozi0lj1ZMCOH1FvijLh7hssgfSRHDRtnhnD8V0Ds4WWhMzWk8RXkjRHX
rmf8x96TZBBRFSV0k9ageivFupOiFcbiVp8cn0GKY3HfzjwZtqnOQmh1GCZgvEgfPWGt+hhdcdzB
N80HfOkYAR04qhIc+nsBwQKkB0pcw5jZNwnFlvdl/wrKCZsDSN3QGj/9G7+IE3UtUTsF28IAqUrQ
Nz4CW9xYbH0zCMNhiLka6jjSh4DK/LJltzpunLu5NdMfpyVKP3IEgko0ivQUtEwME8rtM128ylNf
2BsPZ2GskCF5Sz8Q+bSrUNdifMBZ0jAS7WIp/k6xfa/TeqY1VOaHrNl+VkjVEezTKJeNbQjnyOhu
ZyAriY31I7WD97G2MzfNQF3z1cPJBhyrpuV+GdXTXg5Re5jAFw5ixaqY4/PqQMat9gFF5G5YuKon
qzFmanSlPuwe+XPm7xP7Ul+S9rA5vmzwtqWwue0r4gZGuUaf4x11USI9CR7Qq8KIUYVjOC9wI0zB
wt28IpjV50kZYNRqiUq9tK6OMjTYOT5/1Bh9pBRI+qVADsdT0eRUDW9bI0WnCtjdZbEgB1vaZUFp
QntzL5Uacsst8m55p+IdpNsm6ptRRfgYEIzVdtfYrk56Ry7fQ5L7sMs0L+JobLPWNHCt5w2+h6Ff
ABGE/NhLiG/fwmFbD98gainGNT3k2u8Vv+CBm/2vVttLZQJvnMq49n3zsQJ3YGAviv607fZsZyFO
EvdNYdlMG5SNr14Yuv5OXY1utG8goYaTw/q/DecWgUAOUn6bdNtGDvo6UJur0hjMrRYHns3PElMk
C4jE728C8xdPPfkBo5LJYI72EsQbmhEHwjzMkoHMqJWx01X0EcHYhArmMw8KZXpFlVb+Ql1UuBdF
ayRyXjWrMjO+PG1cJXXPcTsayn5o5Z481oZLJHfl2ikws4KZvDz+OoPgXiVEy+K/oeFuWDmWNyyL
hQHWBNfgYYkWrIFuIM5Vkplj8O/MIeeBLBMO5TGK2g5i9JHYefKQdymcjfH2oJ58PTUlWaqu27kF
XV6bCAG4C3Ajc9kf5C41R4ti019MQxeXXWPf9T7SDSXotDWjDJ1H2VTQBSK1m9UrOjbIMfKrMzZP
2PplhcFp8L8e9tOHR+jeUwP5328gpkKb4f1xZ5ltGLL6hizBwBq9wLFa0H5+CS1b+6wWMwCIKws4
s7rDUpvvFukQ3aJ/X/J6ZqER7/RpbzVi5v77tgOJ1SZNXW8zpyxCNobs9Vl+BhH9OepoS/1mkIY2
qpu5AWVEBumkyUcT1CIlcf5DnJkVXhJy0pqNSPyPST+IzFZLNGNAos9XMttkkYBUXjReA34wBXn7
/jI6nCq6vYZGzJL5PlcRI/qijFr02zfxN2QgBdRHbbnn7FxuwXmmAuUE37EMW9MnL0/fNquA/8Sb
0r1SZ6U9wuH7dGWhYF9xl2vf1jUM8gedDuZ1vCSUaDvIJvXxehMdJQPHGMDMTa3ymkv9WC7Dt8ka
npCdiJ5RBz0DOyRhk9fIK63Kw+99ScorfAtuOSGlSMZxUnGJIHMM4Jl/rIC48HO3ClcNtqym0vWo
a+3gjmRYae2zsjQezV6I8ry+KNVp9tqX39cBPEI8+OUpeVZ5iP96v1pYNlLHo8dhrBb9S8odro6A
Q1LIggNW6YJE8EFwtbNLJRMihWagjtbBZ6DLooGFtp9mI1FNqzapIzcIv6mVtxlP1SNofPEfPwRE
Q88dHCYcJrtizDvI1pLfNH0DLtpTFn8mr7WeGCbJjxs9r8E6Tp66wuVXA1JjAJS2dJeRPH5I5oaE
n7wRY9/n0WK4ePPcWkOQaYp4nZF7o/P3+WcX8RiUFBv4go7RvHGJGJk3+j3rm58EAEqsQgjEsSPq
cQZd699lfFash5TGbR6RhrvTVYXZ0t3J5vCYjsfAHZW2vJzesR2h46x2LZMgotdIw/LuVYfZW+X5
zwGkeymstm+VTfhJmZK00nbY9FJW806tsz2GFpL3X8/iPupgwr3BJ6CCmTUbTTV7C5vVq4/Yid61
DYa9jZyhaomCzYCB3FmB5Ok1Mh9YivObJzHce4wnOEiXJdRfGQ9pvvF6EyIRkDGygDzO6osjb4fF
A2zdhYb37KbSXp17VNjQ2N4wmd7m2XZANv/Zr9legvSqZ+c2ud5VyhY8wqpfYsn8E4PhEIlpy+ZQ
HdnHqxIFzZBw6PexJhBcO53Gx2eJxoFhwviUnRrdhoZYp+yEhXA8FBCxGVvzbawIHx1uBgtnIP6j
h7bep1HvMUBCobEMLYVDcoUAUmJR4Qe62b2/PuR+KoGrrMcW/ouCXmv7sSeBfwaAcw23KGKsHKxV
PWlBoW+f9xbhtELRDNMS/0boUsOEoU2dkdF1i+iTN9e/TOkcd0dr3ADGn6se5ojXWNYFCzHODq1w
WdESx0BbhX7xXc7mScDfUVR6cAAjJcmbjUkU38183ZqQ9xEsoeqAWj1w8a50mxpPvQheb8v2g4dm
mKV0WEbN9S7l7YS+Cym/+8YPMW4Sm3sCxesSy7iVkcQGhu/vI8vPsrhIiqQO803DrB4XR1HjMle2
Bi2OmDTXyAYVK/R/MtXvFY5bUQYXet9hmy98mW5VgusLqy+Q0x9G172G05qFl0ZQm5ucW9GvCDJ8
deRfUocwKy/Bo0uwUwbTrhFle49PLKOleKYbsi8Py3imahslP9q3huh2wBDmJSSIq6BR7gvIm4A0
aRZnVYH3pTQi0w2WtCQh4uS33FH3dgcXxK0njadp2OTZvvP+RBtNhMiLIn4+NoFlp7s/JgHHTfSA
OViXZiTxfXuym8h327sg0+QWQbAhQetEKmMBK5e0BM0lkMEFt/n89EvsqQusLxR8mKn8uZmzBmwc
CdJPvD9ppuPVmjhElNuxo5cphQCIImxnhksNFrDCE2OUImOGsgtNrlbBUIdhMp9Y6iOylm6HKD6T
x3uMkznc48x47v3pVG8O1VKB2xMCaxC1R4Ik6dc8X8EKTvljK7stIf7W6QzHOEMX2ikWQ1IHsN+j
5K/wYACNiVDOrUdUgqOhsLuhclXY33wnY7K/UAPXbWKLAZjhneRZWrC9F1JFOvisS7s2EiYJTHhC
RZE0egos/A7Rh92sZMJgM7aMHzv+Dbom2cJ6DPrJHL020YdSddJdm/0wtBTT8k57kc2VoXbpwN2b
RARcJqb7+k1KLdCj5Aa5wM86LgKBTUEm2QK2lEXozIppPlk/qTbGcEQJmHRudwpJ3ujgV/+N2gqt
a3agA/mCrMm/WkLOydXKLko52Tejy+hYYlnNOhEdxQNA2WGddo6Zcn/wSnApYTZFmoEVlbmYJ154
4TFa9JUYX8pSWW98sizu7oNQqQF1gAUSLSxaQQ4V3yvpu0cRztw0DazQGc4HMw7gWnEVSaf/MOxR
Y2M9FkuzixyRwOKSpGbTP4T2pXsiXmLWH2flKYjnSsFIbIh4CSxPA/Qdd9geQgylftbm5u4pELqM
GySzuafu1ajtgWQHq0/IR9GsMT6dRSSCTBSGuxsPkGOJPqHvNoOepcBng2magYtmH0Pwu/xvtIRJ
1RNlGXaWEr0M4gYJcTYSMRCSt0Fn0cBLy5JRHadH8gBp5/Vb61nJvywS9LbpVS6Gk+vQXtTqCrAz
tMkI4uTg917oz+kx57htuUTyjijTVKoULLBVtlN1hE9JntDO6e96oVoF/QuMwVRumxmkzRLlHxvu
VCiF87g8EDzBZcICFTl92FvnF7u3olnBBpcMCKFUknR2/3Uc23A0FfJmAF5UunqDqVii36cp9zJx
hMA6YeH96rtDX1mIeXty53qQxaXBbpcGXtSNYo6jxy44KxCOiG1dNKGU3alOnGWGKY+ERKzCgpBx
eefmVrNGanoTml2mkhk+gANCQ606eqvW8rjAex0H+rRJolg5JwtKKTFn17RMdEm/9GN1IAGFyO3P
NDOsDFFMTO8t+TI+WJ2I5vsQZ47/qmfGzsUxPisik2J5vQFJfho2jKFtLQ4v5KI4ZqiaduGKCAnm
8yTovdQ9qU8JgPJtuzgoZ53J5zRhWfxRURVnjpu2Z9WqjB2xXv30oWxuBu6G/bkRnd7c7Muk4sVs
/sQMyOkgku5ksWBPXFgmxyFZOYQxdSGMUJyORFngV4TwMyfRnRw1vvqxtgjoNrN+25kLl7otpq9t
Zf2qpYN8sPO27Il03EclVQjeWuLhALi63vKLsLu4yrU8cHRpMkCIrD2rzavkRO+oTqR6Ur3rzBer
qQvsq/E6NLfFmHRg7B/omHRuJnHJK95wUFkTY63vAea4Cm1rOGgGTyhGkCrKsYNsNiW75AINFx1m
agAnX6hZ5ucVUHck6T94CbBMomEjgTS+HsWYyG1lycE81hiEVVtKfAy8e4ooMyhSfPN/oqnwxn0m
kgxV4aKhq2lo3/BcY+Rx5iCSzoFbCwxUuW/7FLdft9IvE7Z8eVK5laS6tyJN2Mt4Bn8EJSWnBbDf
oT/aid5TxU8HIdC+ptAF69CbrcbgWm4LMqAM427m/VPj54Hw1txH4F7sxrNUkyAcUf99BAG49fkD
hyCqKgWHGgi/Pey5rKsI2zsBIWvFfUDYThjjN5m4phChNxvddyeaITyAnRv/2DtfYJRsN0P5dQBD
T8nubwxn/ocYzbALJEdcAe1/qofZA8bnLeLtyj2CBbWHfNMJtuvNwCqtlV6U4AaiJ0SOlYh2I9OE
YtN1JnIxJKzgwkN1suiCprljvzUWG404nNjZn3L3QvjNicOB6x0XqzSGmxlxsHLH90D0dXZeL9R/
6BZwAvcT9q82Of5+q8FkRdMxCCqu/9JJhVgZ7UzZUjwHKDtrvir9NiDNmUMUAhf8jJ5LnuscKeF/
NWY9pqU55GWMYISMxrFTDL/sYZlyV3ApInVLhD7chuIpBa5mhBQjA+B4N9wOD8uLRA+jeUwSVQd1
xL4jaqjA3Af0/55+sLbnSkl7sr8mEyqgjScJLc1+F7CwOAjLiw6Ws7mIXIHg2lMiIC4lpX2YbSNh
yVpVPqWov3j/FfR4pxMuJQG3XtJy+0UpVxnkgY0A6Sl3oc+Pi152ER6ChYbFLncykMXIUhWQaFJf
PzqGY5iPpVKv3/0bixHjF5qunsTkgdQKJa3nHbp5Ec952RlAnqFlqnKOElQOlqM5/2JGEyC1uoT0
b+VlTwYRcirhCr8KD4tPZ9q1JQCdV14izUetfwXcjjkdLqMz4Vuam5OxMogvmdYQw+NINacxCBMc
eLX7/orU0HBrB0TEUEVkKiTlniPh0yeP36+dxLtk4pZyfWZy5pAUDj/2Fc9T9kLO8Gg6qaFIIQOo
MGxh4dtcQJ4Ic4Q5c/73CfbHLGdn96/j7K01FVBKCiaANsra9gHrxo3ndmScp4i6BS50t15GXZ1H
fOn4mtCnTU2SWGEtomGjUUzHv2wtNbTZpbcxlUCCaRmNuE/iH5rCWyjBfwymGyl0PHarZEHrM3Pl
7jkIy2uyohD4utiFK3mFm8tQlKx3ipUgZjWTH8Xs9nRmdl1znjER4gNDjz+cUvAk+T5EqYL5uWgW
3Ocnn3YNwUryAQqN9Q5qFR9fKjr4l4AYVk60YSkX4QENcNItgsTxxapSzVujYeZiy8dEtXhvXdJH
zM4XLmvQPIFndz9mTLY6CkHU12uTa1uTBXyi6xbB9VciRk9gmWmQuoRrxLF6kQF2uCjYACzkR4Gu
pUGzvQ/GZBwDdK+nJnUojasuemtBb74KNpCMjNJIgqlqKlOie0VCe99qxKSlZOHKp+ZUQ/4j+X8N
baDprSdKKRZ5kUQPLfB0NXDQg9o5QbNTIdtkZMxMSeyJAGV4ePrqSKPv0VgqTLIazyPmmbGUq9co
xRD+R7QVn39CwPzFwF9UVtdaRZL1ffb/rGfAC0qwch1eWis8P+ciGMaboarbFd5OXxTokDufqPlV
tzfFUPwZXbNVMMRxT5ykV2kttHigW/L3QBKJS1tKXvatmMnW7mTIJp3bNLWYPxeFfuwocyLid4nI
dWqydMHz8OhRPcImmNpBOHha1z+9s0bc1P8/EAqjLYj4jaNnahGt3qU4EXXzu6jm7vhkzcJIeFYJ
O0J8jByQIZk3G84I+v4pWNwx5BWXewviyMkoxNIRJy+8HbTTfsUUigFGkAl39GU4h+qo97p+7emb
ULHRSkJXrywb9mD5tuY/Um40ohUXnjQPGfnovd49LPMyKaoBUdmvZncTy4WyIn9N+jHwyZm2DSSd
N8F2vKmSutbbfgDPCKFd2SVXNaEJ11bQaogYs6dZt5U75WUk+1dDdatCqm7LQetZSuwSlPxYx0Xp
s+WkeuTZ2BjQ81zg8g+Le+SCwlae3bKFBLXsnIYjqRcj/Cy2+COFktAUGXI/5iRaE5jkXxrnA1AK
COx8YizP1Z94/2r9N7MtH43qWls04B2pBrf0n2t1B5HT2/+x0ZtAwnEOysRuT5eMZyQcxINJnCva
SHFCAfasbBxR/rAJufUpjwm7APWkAlXJ2J/2O+s5FTY8h+WeMa/IH2j8FThirNWc1lxFxysWQBMO
36bqfGBF6JJfSFzCJZ1NHwQ33uHIb5xQFMWwwC5jsTpb+bMWh/Lhqx5C92jtUDEd6YqmSwpvdcQn
hmvtw6Gfnx6TbL6pvYUSvEvjadQyMTwfBHq/alis8V/2Xfp+yqdX95JcHP+CXCrFpfz+8ULJrhCJ
vGLO+Uj59Iy1E7MLF5exIRqTrhzMuocvLODJVYHPKDNcXLLc4PO3n97qs/CZf9UzDUMZCIwEl+dm
Vz5Q+kw+YeAvXvBb1JicSXLjLNrkWvv3uJ8cKnZv7tNr12MtIW731m+9EZYhCcgOF7I1TNyiYY9r
TzgAxZVu4nmX+5cCV0JrhLPNbcej/MkuS0+qk2oC7Flne6qrkS5BgXhQES83TkeCXW+8ZdXkkmhq
b38W8IpW6rm1Z0tjXLNl46XyzB+4q70AuGA/ElKcbbMJ6Wk3YUip+xfRMHZCZOEI1O1ZpYUVtqBQ
HT6k9XfuBhI6SAQHvmY2jxWrkg+3gCH83h0+mz5dAaa5mj6Puk/3AcvRoOYKZNl2N1tKmeIEGhWq
vTGHKNJ2to5/GKRzhYhkEBi+CjRXosLVejCkxzKgU25ahgePtezDhl/SBi8saWBTf6WjNfT5NJuA
dfDErN51hAJ8BE9l/K9k86TG+mS2aEsN+BwUT79Fvd7fJ63xzkKY41XTL6aiqeKtZLN7vHrWi+wP
B+NUXwDYMjTBW9dEm4Fl723TZoEY+jfqg05Es4MXmXX0ht9uExjQ8xv39EI5Qlc3nAmjKYpnfuSI
VaWLGE3F6ZJp58P1jkV9BKdUgGSd1AxWImEhaSWJNj9QECVZvXmYQvp0FS5joNSNMdjLhCVllhrS
0tgjmXBCzsu7ATVwgdA5j/wQSrCD8SrMB2ii0CglZaRjbjFxWbso847v5UD5UonwZwQr39IDTTTc
OocaQ0Y1C0aVCVIN2uyd+UCd63k/FoPmOcd64lmu1SSyNnmp8lk1IpCXubiKrkEN3TR70s+O4GCz
gE1nT8YDwl9yAgaFOx/gbOucOUaq+FhUPQfMcCPx2RXb0YftwhapmTLAkf8/8bIMByiKwx+f83Yu
kUYMqhubdmXbfK4BK6B5vvU4Q7Bqr7GBE9E5SIF5dFk36Kox2KiSqcuoimj8totYJjiCOdBiuqPl
9UiLtQcduPnG+82m0wlXen8dTcxAG1I69OwvvjQdF6ad9/4p0h1Xq4wuDC7g3bhGWb0E6BYedCog
mJ4kqH912vaFyE7pKqZPqXOekCB06nqcKFIgsfiGQ5d8VqVPGc/kABCwbknrTjBpgYboAzHmqEpy
sF4AbctCvOLxNmKdgscRbVNWR4+x0d3rzwmFHAOOpwbM0VA23ogVjIuqZjJuy5kLXJtMGGOvfMHY
mbg+fNraYd8zc9N3jHHAB4Lrf9HcU+WtaZRc1MBgw0a86gqn1uJm1F2jateyYTjLgr77n6E4hv1l
qg8LCowkzmTrqe3ldeHF1x9ycFLivWzC1KAzmdAcJlItE2dtd9Bngr+4SCVITlPLG6pH0bE14HnN
b9aYu6rkYz6NX/bR8FD3+ySB2nIf+OOsMXhztWaqOgDMQAPVq6CkoP8/sSILzA0OPzERPbOThdWR
TMcS9Z7Sx4RWDgk1/efUh/vu8PpqQ9kdGZD6BlPM3jaiJ1Veefg2Gs2m8nhwzEsjEKpllvn1c4qp
Q87OnCS7EMrb7W8Vd6z+zfqMR04fgFZ6kB4Q7Y/ndurvgsSQzfd0uXnmxIVXvWQTuc97FHS6HsX2
ErDRKE04BtOABzPKIa29Wr9tvM27E/k5GEcCAXAC1h/jCdszSxHGCfNeHRvl14hums5zwkkCqWlN
JtH8l3PviMrnysC9eO+H3YMQjIKhPlGViBpR5yV7bQ9uxO0gvlAybJ6xanlTmd7LjoN7L3xAeIoY
howu5M1MuXAJ0qpi4Oi5MdH3jloXsulkpjwjbEcg4YSQdTVXdTn2LA5VJFu40IqsQenFmOtXcrmQ
sNZXz5h5xCdC8yT+WVYTGoUI9Vs1eJ955/DdCD1HI2erTkmf/c5AtaKhbxSCw6a0lty/VdieqkVb
qGIxQhurf4l1CnZXKL1xLaQxo2h8SgULxsA7rvA1HvJd425VVxlzzwbkUPvBDXp5zrM10Vduh84P
HwrD42PQU6ajyucDZT/6vtOOcHrXXI9DlQPbr4R3z5Qzt99hfGTljwXdrPeY8LrBYLxz6/fWS5lc
AtTl5d/s5YNeaFMQwhunylRugWaUuNH02xLRgIRfe7QDmiYPdZJl7tO42mMDpjDCHz0jZqLxKAoi
jIURyFgtxzo9qwXJrWfwSxU4T9gf7R4KLcwUAg6GQOn3XoRkoX8JJ4xrA/dAze5G0URkqJV9tS48
/WEqvGTlTLK603FKvo82OgRWVRoEvXfVqX28XyXj2rLdrCTq3yQ/9yQLxYdg6E0LlI7od5lW8uJy
jG5wvKkrpuAP/+688v3E4PU5udl7PTo9mWKVIA/M9CZ1UyiRP57H4anAmzHNksAgG8oBNpd+1aRW
Hyd86mht2pX3+8Um5ssl/bts6UOncaBktEx60ndC+Iz2tyLtjRra1ju95ByIu0LpZgybGIKiUY90
NdIS++AwhFMGFeIo3u3MbI/r8ZU9vceolTRPI2N/h+dJdfbHByI13zIy3I/ToQR7liebBD7nMrx5
CfCQ2Gbp9lb7PPc3XwAx2EMlxh5xd3B8/Hd34+gfA8Bnlp4u2OCkasFQdiMS/kNtfeQqgyJXQKXP
f4nmVXP2mWheBEp7Cg157ACH0zpQ0lUYz2FLsRHj792KpezJ7ep3kLpss+SLLmj7OW+eUf0Rli87
D2SXmvClZPEIYm5VgGV0WFPKTrYJ9kMqrsgC22KxpZduVGVYdvCEVvIT+zmcGOycseuXtnIlSv6h
N0b5cP/PTbN6IhbUKaZzOfHcLO1qrlJNPV8cvFk/d+m762XLEhzngcKkBKSfcbXVrHV6r63QLfR2
xDTj6OzuO15dW6Shnv5v2kbJSbs06g4Ae+cXZPsoNyVBkwDE9WI4bBbIF9lIRRnnvndp7y6HYnS1
1Fs6xrNzmaEa7AGw408rLocnENwR0P1OdqC5HMf2PHGshXodBrEGKp/VzqaNFvzjJqVUnetKRqHH
XfHisxJtWgySHV37+TARKORFzqLBYE08yEJfqQVu5FSyWGG00D7CXJaU9ugm5BBkIrO2uEEZhCPg
y77qOJq8iCmII3Zk160U5ITYe4rT8RXLXdZ5C2ogbf/GbfOt74XL5Pp7JnhZ4Rxw9clNbZnnFDdJ
4TrZgrbgF6WQjdPFJyVPj18ZyXtnLwG0A8U6D1J2+9xgM+BDNmxJClrwov2kW9WL/10H3X4NkDFs
4xHoz58uSu1t+xZUXx7orEH81KO2McVxmDvc7oIQ1SIPxTe8VF07e3XDQloe/uMbV+W2f041t7Pt
LW+oAecpd5LBBltxm4Qo0SmbH6rNs/RN7XXzTrAAy6m4WO/nC/dJsF6QZF9wO0RcTTqrOiUk91yR
3K2YndD66EecnahR+IHZD6V20MYYjcN+71GAjQJ8+bd4opFfWofeiB9dcfvt+RMB9CL7mRMEx7yV
g8q0r4LuFrHDSZ4p98tWH0xIYmoa5tCPCvUawdfxU885gf/IErS0uO1DJCBSFec8NO+PpjUNo+5A
p/53h9etNUSlPXgUkfBlSORtvf3WGfpYqtNpC7ahvYgOQVc9S80p6Dml9Q5W7RdCSOvT5bUacCu+
VE6wO56GYdHR0p90/YjH9992Y1GYee0F+A/lpuGkKgYInLjYEKYq8BECm1VKQdUfh4lbHRqCXw/u
TuGm/FDpqbjdao8AemcfiKR9F/aQx07rEP2BJFFchQ==
`protect end_protected
