��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$Rx�y�<��wA�*;�x���@�̦�W�X�fa�M-$u����n~�%���P�$��W��kYَ���P7�?UMfT��q�6�U��k�>����~�\N�(�����X�e���/6U|)�X2pF�]$h���d.���9E��WG��L�X"]�Ad����ľS���8od����e�GT?y	7�������ݵ�^��R�q^]�鍦�����s�ae���h��L��P_���ާ��YЭF���'\��68�b�[����w8�[X��V�F�0͘3����q諵�uW� �h�u\V�?@��_6G�_�*�G���B�絉�f������[�G��U&�����~�F��AׯK1�`c��[<��FY���4I� �#�G��x[X�=�Q1��`��R>(�w����R�O�?����7�,(�H\�#h(W�EH=�������yq��Ѿ��aF����:�U~m<|��.��0=�P/���4ǆ���T(���0f 6�����!��ݱђe~�xѸ����v��YrGʹ 7c_DP��6��~�m6��;�Mc�b�pZ�p��<iz�c �8��y�s&�9�]�'@3*z�;N��{�B?�|AW/�`��iY���ʟ�OTܢ����
�[7]&Y&�Ş�ŭ��q��r8��[W���s�/fc �@��ʙk^h�G������Ld	���A�ы� �o	b�T
&�з�G*�&V*����_��xv!4�����p_���Tr�QT<G
��WR��
�rH�EX�� �f�����!| ��n�L|}5�Ŝ%���u��Z�d�1̣]�^���I�O�l���E�jI&E6�ŕ_:�W_��ǳ>��Q^��>A��lUX��28��Xd�>h�@�;�� ��1��(�����/�&([��}i�t�\���Nq9.;��.T���'��(�dI���>{�z���#Y�5k�� V��]����Z����x���-V7����~��D
{Y]>���k�k!��	֤��`H�JC��$�nK���NDi�
���Fs Gm3{9a�v�] ��BŦ&XT��&@)VQ��T�!�ݝ�f��+�j����>wM�x.����2� ���l(pE��:���%��6c���Y�s��#d0ϣ�/-?�D�Z����ۘ����q��O�W�L��J1-��Mބ
^�FA��tX�:�b����0ek��E�����_ٺo�����:��W4����hV�Z�D>��.�5A4��u��/�V����������Si�R[C�b.{rfY�\��'5� ��i���-낡' ;�I=]����,~6�
>�U�]EňIOP��z*�f+�qe����/��K��9�w���י��Ԑ�$�N��◄��Me@Z�=N��\��f���ĥ+8ܱ�(�d��J��ćZ2��Q������7^D�9�fwt+e�zW9�Id9���������۸��SQ@��>D��Z�"�@i}�X��3"�)�xt���Q�z1���r����_��ZS�[/���O0o�c�.&�&����E�Xԟm��$���=A�ޢ�#_I7��
�m���Y	�MV�hOj�$�3�L����y��yhNP�i��O8�l�	�L�n�'�Uo���3}�Ӕ1bh�a,FzNgy��:���\[2�?R�H��+��.��FC��Τ���Cӟf���B	zkP����Y��ј�3QM�=]	k��ޭXjqoq߇=�9��o�1Mq�]��"�V!�]!F�2��a�Ř���85�y`n?��Q�{���s˺fF�^P�q�I�i%��U�Yl���,��P"X~rL�v��K����'QIs��G������7�]�����E�f�C�$��()D�_r>���	�ܻ�ߦ��k�(��1 s��~��:N����-B$�M3�h�_�S�EoLm����miΉ����8��cFSad�k�ǃG	�F>:�K��˰�1��c�������+ٴ�w���g��y`�	Z�y:�B5���D�_*mH�_��p>hb�B.���y>�s ��F����q{�{��1�By-��;��rQ�D��������M<Gh�R�;WDԱtL��v��)�L���o��ʴ�ʼuRFg*�u�T�ψ�%�yG�aa�5涟Ul}����Xk�weǪ�4�b����q������m�K�yE2�B�)�"�AF�*�H�m3D9����X���%��=�%�{F����0YȬ� ��|Y7Z|���M$���H�t:#^��P.��y����J|DG�_,�O��_� �K'�|�kY�Z�}�paN=���~3�*g���~ir��y0�Ͷ�x�t����|By�.�0��?]���줐��_P	�(�KQ!���s���n�k�*�'�����D�{v���Y9E'rۣEeR6.�%/��HX��*�m�$�X���q��b�8bhc�MSO[���͓q/�\ɘ�G��ۄ{D��������� �I�t��$���/��i)G���ȓ�{�R�W�9�z��A�!ϻbEz�QJ='5TA�G81 ^���&w7j��CM�00�F8����O*��|E�iR�]�VxT�K��7�4�j��g�r�µ/�e��oT*��
�j2�����o��O�ms"V�.2�}+�m�G�l��VH皷�$Ho�B�����,,�������u�gF�J�ͦ�P0�LwO���1�ſ�;c� ,� c:����`Y��]��oYo��M�@��@�lWX��r�K	l[��I����q���F!��^�\2/�w�ю�n*�3��Ê@1�Md�
��P�L��U�I�}C�{��~���]L:� ��j7^L���ϳݚ�� ��@o����풛Y�Q��몭ѽ�F�a��A��B*1�<3�]���Ҫ�]��`a���J��}Q��ni6Z�������3ȋ~�i�f���E;(C����@�
��� ���a'���6н�۳1��Fr����{%�5bti��U��~0@c��㧧��)K��XO�e�m������vyO��0�s!�=� �����_��I�'̷��,P��T��",7>Y� ����C�/���^�_�S�D%�y�V����gYny.�!�\�K��Ɨ�����H�\�~�R�Z%h�;֥�il�D#Ӌi	��l2�B�|�H��~�K�.(�:k���b�tW���*a��>>�v�&㞏E�c�$f�3���:z�7�۩[=�i��ZH@{�Mڌ��-I#DV+{A0&$��eyx	TRi� �ݎ^�����HD�ƃ�j��W_�Q9�S���c �>B�Ɩf/�U��+(B�kc���g������N8�t����#X'����c2JI}_7�5(�q�X7�{T����t�|�zN4����J" H0�ЅP�dp�4媃/���,�M=T���V�ԅF������Xwm���Ȯ$n����;n
L~K�T��~��|�����)R.{��g��%���
����$i�7^|�.��1��=���R"�ʤ��''���D��з���w�
�UC�G���$��s2!�UC�B�?1@HE�G�K�Z�@ў`��&�r�>�_������c��^�S/�T�"���B����*A~�^��rH<��P�-�w୍2r� ��uf��l3����J�W��Xq���.��	�M�[ܮ�&�Þ�P���c����IFhe�%���U]Q��:L/��w݋��N�N���[�r��w�5_9����;NP�����+烺H,k{٠�xz1�L����IɿP�%��c3��R���E@}/L�;�d8�-��H*��x�]gO+�"&e���R�i��� #>)^i" \cS�+M�.�x:i@ҿ牌l׬�ͷ)�%b���։��+�ڃv޼�5d��d�邺��=���E�#�U:'�]�����q3�K���ݝRl��CJ��=���@��S��u�/��T���ԡ5!c��ċW� �e� ���7�U�r0���J]����%��mJ�2��"���B�.~3�O��c�Z�����]��L�V��+��=O+��y�O��D�"v��:���t1gj�A�'��r��㒌��/�C��Ϋ*�D��ȩ�K��2T���t����_R�'٢�"��2��
��'-tlNGyɍX|��=��)L�	�U�}�НA]_�)����^�kL��6�M����GqRt���|�z��!*抍�2W���M����%������@[�	�@����
:{���~�- [c����&p�O�	}M!y3Y���ŰW�\hh�0h��ژo��6�0xLE�w�43�Q+&��P�k�BR�bc(s�﹟y�O�s_m&wV�>�\U��{��Wz�F~��p�6�<��Fj���G�^��"i��_������Ws���.�;��H(Rf6_�kR=��l���qs�� �#��5�jP;(���V�Wp���
�ى��G�ُ�#���N{�*7K�j>I�i�|i7�#��V�߻��vr̪��y�m�_�'W��}8q��e)�`R����З�������	J�M�כ����)�E3j����<5Ӥ��"�w��� Lt�D��ةڭ��k�<]!���.p5�>[�w��dj�x��z~
���+S^aR�,-��A����2�'y�o��8�tFKq�w����,£��Rdd/�P��l���Q���)jê��bk�P���R��x]���l^�&H�a�@d^%��V���xI�Bm��g��n�4F|��s�5�+Ad�.,�K��'M.{>��ZlxXU	FWg$��%"�וP��W�D�cO
�����^󾑆�5�Y㶢M�<�w>
dF��%2XZ16����kNu�h�}�V�w��3ds���������q^��J�SKm�j�)�I�|��rK��+��4�X�	���(����y��S.�!l\����~����q̪�AU��%�8��%�C���+w���J���8���AN�ϛ�E�uUD�3���[]Yh��_��/���H+���]�7�z��ꈁf��$:�Z�M$��z�V{v����a����w ��d:�v����� ��ܑi2�j�=�`e��#Z:e����� ?�y�\����(Jc��E#��ѥ��"M��R�o����D-��y�����)TLu�f��L�,S�N��G�bfă�^�*
9��ܾĚ}�u�W��F��o��n[[1δ��C��.�W�)ŝ�t��5A�
gWk�����1�8`�� {�|��L �
�P��ٻ�����f�P2d�T͂?ꉡ\���>=�)'GI�^���-�C�%�q�Nc��, lcc�5����iz7�^ �8F��]���^E����
�E�~�wܟՏت.����y�|  �{�4���N��C#�ȥ�q�ޠ'��	��Ԧ�Ա�Vį*׈y�˞��E��i��v�9�=-|Km/���|�X��X�VuS��O%g wv^��^�]ۂ�Ж��KL�Z�[���jH���a-AX�5��P�<&y�+"y�N,�ۏ ܑ�B�ލh趵>S^#���mo��|TeQq�~KbJ��2C?��w؎'�=~������[Pr.(�xe �v�m�f�V��=t�����#*�%�6׽�)�r<F0
�׮;��¨yy�W�1�׫Ȧ����kn������ɑ���ƞz�11��5��M��^��6ߧ �V��ڈn�#-����y&HE0��D�N�?���Y#��V�Haz��k��Z�]G�b'z���r`��_t�\&6���/q��Í��Rx[�F�f3W`f�D:ͧ��B\�bg�_��'|��;�A��y�c�w����v�#��Mih��gOW�̍
�U��w�m|B3�+U_�ĴduG�b�1:	ޛ��8�_��f�S����Bj���I>�V���Y}��;���;�Q�������6�������<��iq�Ƥw�9p��}������٥� *��1�H�c�)>j�%{;�+`z@@�Oϯl�+t�z�/�`;���E@	<���;�ASJ�*� �@1�g��8�]2�Q�^��rQc�c��ܤ"Q�h,I�-�<�H3?�7d��*C�G�wP|�t0���ڏ�Bu {���~IU�2�AO�ݶ�A�7G��fG�q�t���_W4=��+���9D�,�L�	�ՓeIR���/�T�;��I��06�k(�$jRhTA� �O����(�n�y��QV@f��@v?�gB�+C<J�;�d �߰&��)$�~\��	H������^�+�U�9�ꚨ�p?�4��?*��˥��|K�H��{��q�j�n	ĭ�-'_Vo�{I�$J����8��&�/�?��m����-<�.�Ǫ�t��+5���]��+�U}��E�$Sk����=���?B{t=^�O�b*�B��	�SL��H�z-8�e����l���+�݀�#l������w"�I��G�����I�u�\]z0��4F?���ItO�],�#}睕�6[����,�y��o��uX��VdQ ��4����{���1��.gȐ=&� ���m��~�w��eEސ����B%���@�"���`��K��[p`Y�&z��6�x�u�1y��\A����c7�+���1^���z��B���?K����Ӣ�Y�҃7��0���k�w��*A�N�-���xf_���ҫ;E�-]�b�{�h~��=��D¾�y����aZ��g�H���1/��9e(�&�^�Fb��x���<$lT�3��t���e�7��g�,�|w�{�@}	��'����\崧6�'r0����q���:��~��R�s�¿2��ԛ�P{�q�iԱ/(�v�qb|d�������ȫ�5���<o.�_����N<\�4"��
���K�]���p�?5w�����dI�>e�shE��@�r��~>T��LLl��qd���bђf�wsN��a�)���Ô��4�i/4�cT�����UV�T{���[m��n�CT�sRV���������{���[����M@&��5���8�@�<y� S�:<��$�aӢ�%���R�.����_䬟�R����d�>�m��
��ٳ߀p��3!j�9vp?�o��~F�W�e��OB�,��W����ZOE.��m�W�uҫ�oB!�:��u�a��2��bq	��sI�A����;l,���e�1�?�@�0$�N�X�j��E�RǨd<d��-��/~���/۫''�i�&��D�����l�W?�e&1�q�.]ʴ�c�pߣ[}	1��|���D�ɦ����#��,tb��1�!�`՟�Ȗ�$��K�i��Ҋ

�i@6x�h�fM���4���ǭ����t t�XG�kg��<�Xu�2D	Tw'��ڠ�S��vO��]��?Z��my� �C2�M?X�̃@7Δ��,�������@I� H@�l- ��E�F,�?�)���ߓΣ�'�����Y����6I8׊�i�S�-XP�]��e�_I������4�PGn���2F.�U����W{5qn�PdV��e�qQdEQ�i��X�dML:\u��;Ԥ((%_�π����� ��Ҡ��ÉKck�(�W>'��o�ϛ,P�Am\�*r��Bf'�-�×yGGm�c�n3�v���mJG�i�B�V�,��gG�v�[e����C������%?~-}Vw�op=��X����/�Rd���z0�3ǋjOQg/�c�90��"���G>Ϩ��>埫o��5 �m(�F(�0?gos�@��&$b6�����d�v���ᝃڡ>*X	��Wx_�ѤD�[�ye5��or^n�`(퇒�L�j��[��q�#W��[�V���o\F��c��S��W������2��(�_��T�P�`�,�vOe����a��Ĕdf��r��o*�,8G��|5}�0(R38�3�/�	���oV��"/ ���T���u�X���'!��<"�8U��̒���eД1	�<�@�G���ߵ�ԻB������Ղe%�W> 4����^��T�c�ܲ�J���x�7B�њ�� �5�4�\�_9�/��[��H�������5���97�8e@�� �)O�v��%����8�K���1�[1]��ng�����[p�	�Cg���(%�8a�h+ӅzbwY��-w��C��C�t��&g�ϓW��2��X-@�_{ߣ��x��,�3ϭ+w�ѫ�Fe*�?JOp���%.X��G*�r��Ҡ�=�%|X�#=�yȅ�jO�F��{f��#���YU�RXy��	x�D��LY|>>���w::"z�(5%�N����k`U1���4��|����	�.�+�t;�	c����f�����^��3.�/�.1D��{r6�5	�Z����k\O�ct025Ja��B9e9��M�3V�ݫ\_'��_e��VSP�!U���M�"�f�|g&J�:P틳e������Ǹ�G'0��<�G?z�M-%��dF~(%��a��FL?˺����c0����������#μ�Eq�D����=z��zK��֞���@'Su�u���.D3��1��e�%���}��&Y��C���[}�"5�O+�����g��&��]BmA���c!�-i�Q�O�����^�Y1�*z(��+"a-���U����	�t���SK5��7C��?�� ܁�͗ذ�O�g��� �K�S�_���E�B� �I���7o�u�M.�7,�2�P\�A���Bo���DMnR��u�?i�;�HK-xΙ���=(�F��@4�٩*Ӡ#r�QK�-M'�O�tcת�)��kH��sR `��Tb`��ݻ(X�H]���������pqʚ�q
���؆�2Gȃ^����d��M��E[��������>��?S�1%�:@?y�U��T�ĝ+��*�����P,�'�"����%��r�0�p�TXg���>S3<t9z�~����zv�Ip_�Ce���Tdچ�j`��p֫;a�SUO;���=ިs���`}N.��%�G�be��.i!�ޫ`~�=� 4��tK2o\;�.F�T���(hG�ˊS!Rv�&���+�
��6���m���˰1��:�JY�mH��7���f6;�7U2�T����h�e��|5�s cTQS5�J��8�����{�"��'�w��2(�8g=��MGW�m�0�.��E��Z���%f(ٔ���x/�E��4��'N+8��W��.wUDg&W/�Lv �Y�u� i�?-
v����Y�v\f�^�ٽ�t3�ڂ��+�5ݣe�>��i�u�B�$Y=�����V�:�J$<��F�v�P�|J�X�S��Oɯ�@�玺��/l|ZJ_ ��P Sw�,a��-�4�`�M
-7�� G�I���`۸���R��9����m�42�O���@ތS�rCC�����4���@ԀE��v�j�R������?ٟ��g��
�u�e�e������K5�6�M<v4����%	�+�2����C��x��":���/;�|º�Q`�\��9��g+��=Zn����۲�Ud�I�d�1��$����W3E�*U3E��s@ca��wݱt�a�	��+�^B�p���)��bb��5Qfh��}uk"���OdB�׊� �m���ۘ�D7���w|ޗw��6����3����!��η*>6�`֕�"���3<M���C �nr�&.v��3��\ͣ]�ܼ�}��^Y�?}v9�M��/:g�����*HG�L�{�pZ��t#��~j�ٌ�ՙ�ˠeY�LAu��yf༱�V��d[6�x�~��&��٨����$͈iN���U���R�1(>���?��&���7��e���:�ڜ��^��Aw6�j��8&/��'-�}Q����������R3�i�xv ���}۳��.w1_��Q��$�*F�����>���Z	���U%S��HA���Rj-�+Η����4�c�Q}����~�Q7�O�:���.����C������7CB��)Y�=k� "����.%�T=��\e����c���p(����{��^�HP�މ�,��X � ���X����m��D�����+���(W��P#'��1�E0W�Ĉ����t�]�Y�hC��Ⱥ��Lt�V_�盆Z�d�N�b����z8����%�����:�a;����K;�'N�9���܍+K���H+���� D(Y1�� Q�����������#�!�LIwdGe��V�	�Q)�y4�I*$�ݡ+��Ƀ+ȏ[X��D��W�����8�w'�w/HQ7:x�f��Q�CA=�B�B�q�IF���d���D`w�B�*ǥ�72����?K�"�����"�e�"'gP��* ��)�� P�P!ZA��i�wEU���W��-��Z)%�;=�:J�"����l����a*�>��������v����#���l��*ۨ������Ws����$�&��)�{'@xj��m49AR�D�%�xI�\���g��j�q0"t����'ǹE�%�Yy�`��_�2��@�S��k`Q>+�Z)x�T�ou�b�`&�`V����F�3�粚a�4<�߬���ך��iɃ���U@�!_9�	E�Op����=�*e:��l��c�.+��<l��*LG��C�9�G�������K�P�ؠ��0h�e�[���=^I���Ru͞莉s�V�-�kM�}�`	�,��e}9jR���7��b�7�q�i-��F�lJ���)���*`>�2R� �6�r�b���&�np����`���P{�ߔC��w�v3�� �83̇��הc�.Z���mhz�ty���ѥ/�l��)�ډ_��4�^Ru�7
o����J����	��O��}�\��P�o���������}{�cwp�Di9��8��f���㧇��S��(~w:�����޺�m��~FiL��m�%�K��L�]����!‍gotoj�ݞ<Zu�Ê&m�̋-��d�G2��0Vk����u}�U�J���A3	�M ��s�j� �{��!�jE쥫4Y�^Y��9P �"� *eb���U
ݓ
�6�m}�q"�W4-Nr!G�!�Ē
NGA���#{�~QX1���U<G�F���6(�@-���d����$,q;4	a��QI�d:�s<�M#SI4�6�㚰H����^��X��)�Mh�)\��+U�1���7Z��$���}�y�5���F����]N�.9���~,��(^&���dwi���?��	�hG*���+¤�?޴�{������oZ�Iw��31)�}Xu@w�@)偕��y*�K��ȉ�p��u;�0w�����UM0��W�W*a�+����H���e�).M�A&n���j�(�,QZ�Nm{���W+���}�������}hq��c/�],Fը�l3dLl'�n�x�9��,������v�y3��Oũ�oeBALL��.�Qu�>�ɲi��h�� ��o�.w5S�^�Az8��Ir�;Ĳqv����瞥4���e����b�fd2~{U�2O�I;�A�P /�gp�����;��R?�	E:�ŏ*��y(�eAQG&p^�ml^���!�o�Z^�.���B8g�,5k�]zޞ��=�����uA�^�C������|�@q��?�T��
�ԟ�@gZ�6;�΃}�;Q��U�֗�mV����c�W���KP���^� �]U��"n�0�a�	�+����v�&�!���^���&5�J;�\�.*�Uq܄�.�V�NB�ָ<u��(L˛���/��z��?Į��+%���ژN�5	����G 4.Y�\�l��yz�!pg�=��e4�2�;h�N��q:P���r���<n5I��_v,>��4l�^R���k��xm��q���y?-�Q�q�q�$́���&����-�&�U��\�v+ߴ������C������=��
ɝw�â����vo��O9QC����cWEQe9�r�6��OX8E�3��Å���q؝�c�5��6;�d?{�]���.���4��%��Һ�/����'TE3~t��5��~Y���2���$�?�X���R��w�����ǐ����=>�<�U�yu;���?��A��p��#�Dٽ,Mk��41L��^@������3�\�z�9���l�&�Bc> Hb�]��B: �jZ��_#<]�0�g��ҧ¥�%�a�bח�V���֚2rfӢ���Wl؀.J	LWVߕW���Vp[�A�&;0�#��8L�"���6�XnX�2�5-(�������5V|�4��������D���l~/�a�(DbZ��X&a�Y��l��e�h���ٯ��p��9avAiM�`�֍��~�$P�ܕ�sE�%y%������\?rn�ھ��n�ڜ�Mg�N-C#��;�����g��}�q$��Pn7�$��A$��);wУKKú���E�$�5P:|/��c:�x���e��nUT��>I�b�*�=��i�,�`2�h+����őZ��o�Z|enU������GbB�������͉��i�Fg�f�o�!VF�nxT���V�p)�Qo�An@�l���,�ų�1s���M�;))���i�*hv�t�U�����'����g=�K��m�t>lg/�
�1��>�B�
O�q*�0�4������P�!�T�X����T�ɀ��)P�`{h�-"�_-�IZ�i!�8�q#�K��������pƲV����PT�|kxFJ��`�0�X֧zԁ�=�N[�kq����ҳ~���J���v2��Aj*$�	i�oO�d�sg��_0%qo�V�����fJG�c�=�X��@B���u�S����iu��k��L�f�;>����<D��8��)G`(��o��U��G�/oWUگ��c��H��K�Z�9�[-H8�/�OsE���HTh|�������cc*�s����g��7�u�&1 u�^Ə[J6�-��%���x�˿N-�nO�49�vl�>�O�<�b�u�?T�M��i�Z��7ӹ#�������)���ԂA� �����1�?�u�8��O5d��tLJME��U�j%`@du�-ҋ���Q�o\P��.�%A5-�c� ��ye[�����/�� �_����0G����(�1��Q���i	��D�xfklȧ��)��lq
���ܨD�`���&����#-`6mJ�� 7v��BwW�k1��������O�f���Ng#�d!Ԟ�lJz�W%$1h\]��I�lQ :��Jt�pw+�8pK�7֛'�bڽ6���YO�*�|��ɐ,�pn�j���جj��*��VC8������G��O�MR�nW��
��i�B)�*�v,Hf, EJ!_�����Md� �Ne�R�nk魵>��a��y�I(��[��b� �7�G#'��w����FQ��;�1����$�sv��L�3�/�i�h�:I�okxe�K��5�y��$�@5ddnl�����'�+�X�����ٛ��?I���Կ���xŕꃎ%��H� �� ��ֵ������y��Ǜ���o����~��p}�ep�i��։�[+̃�1��:��6Ds*� >�o��1�ٷ3����ڈ���Uʟ0��k��Z�Y�F{���+�p\pR�]G QM3@��{�
!�B��N��1�+���+ᐁ �u�z��-�!�GY�%�G>d�$�F��M��Ҳ�,�Ӻ��(�G�6	�:!����Hͫ�<����9���=��ɐ�S�o�ҿ��7���!��� �x'v�m�`��C��%��`��1��� a %��R}����'�B���c��xH�n&��_P�`���!c��>�-W�~�vȦ��6�Y�4�r[�k®`13���[��@�t�7��'!b�2$,� �mO��1�:�qp>��|����1O���jI����4��s$�D�ll��L$�}[�c�4601]iUʘqQ��������٠!���m5� `N>�k+*�{XW"�m�k3V���A���p$���2
�	���y3!�㇅ ���*�ݲ@���4N#����wp�65�"TIg#��C����|�^�Ǎ�\A�"��Ɩe	�P���7��ĵ��p�5&�G�jY�͞@�<��XzVy`������r�L��c,�2u��o� ~,~�~��'�;�=:���o�� �ӯ�0��K����,�fb:��g���6c�"I�n4\�_�F�hx�]ye�t�P��+���FYk��s��#1�tQ`���C��&��c�@���@�Z��k)��<^��4�-��N�?X�	#���/��/e�75�${mH������t^F���0�iMi���+2�S��JІ!ZMt5��<��3��f��%T*V������^�__�����3���-�Q��\�oB:�:52�C����M;2MF?���C0,T�~�)I"�g���4�H%�JySu���o�2�q���b�ANz;�*1D<���XR~朦?�Tr!n����B�dT
�}uP�H�4��0�t!w�Z���C���v��X�My�C���Չ��#mǌR� ��Ef��V0�O�T�R���n,�iA��G�\�͛��+�L# ��)>+���,��hX�7lrN4���Bk����|g�}-Á�3�]��/�2�ʘ��wh���G�-f���*y5&���F��݀$gh���t'-`���CՋ���h$�Q��i`Yw��Tx��q���U]|��-ռ�塱��P@�)�7s}��@�\�L[ɧ1�jt�J7,}J	m5���W�`OI�ן0`����M�k���lɵV)�/J�TM+����d�c '�^g�oCh��hix��jXAtn�����,
�W�ٞ��G3�}A�Z�s�\��%smvW/j��o������P��EE75����BE�.VsG�~���!0l�ן&�G�
�*��������dC�Z�$�ǰ*(��7$� ����v^~���^�8G�mo�Ӫ�j�OK�~1e���a��ݖ�o�Ϥ�'\p����j8_�������j下#��,��1�zO}�t��'w�'t�����Y��v��ΰPL��#�x!��r���\���h"'����o�A���2a�+.�i�-P�ݵxǉ��vv��40�'����;���ҽU�gK�ur�^�3����
��!(�Xa��V�"���� �׌{}�?�c�ulI��T��hN�'����,a��l����� L%rj�����hΠ����h�e9�|��_c!r/C8~%{L���:V�4���qJ�����P|Ij,���z�@&2���T�a��g}M�S+��P�����%Q�H��g�*q�r�g �3��U�Ytk��q��o*1ff=��Ŗ��Gv@B@�A[��,�5-%�s-�J������l��	A 8"�ZO���W~Z�h��z
���Ӷ*�2��?����}���Q�z]�)F�ǆ����Gc���Lj@巻.�r5�y�������e�~,��e0%a+�U�!n!dC�kh���,_�UY'�a�8�����@�q�^��,>��ǳ�׹�������c6.<������B�jX��tj{u�3?m`5��$�w�JU���"���to�u�䍪Z|ՌaD��>wUF�R���������ɜv�5�M���q�U��.;p�!�H&ޟѡ������$]i���c�嘍�@cfP1ވ]��"5&�L�K9}l���7�):�pOC�I>�BK`�q݅EQ��I�-��d�����z%�.0�p_�'�ᣚ��6�!������.Y<ڲ��fޑ|y�:ms�*72�WJ�:�x�6�9����Ah���S�({�"�2�(a��W��Z����d1�/�թ�O����+Jぬ��=cץ�����'`�:���������i��D��X��ghn����4n�TK*�G� ǯA+�6d�J���N�d���{�w�a�`��q��5=�)�$����4 f/�@O�&�:{�+�����*�d���ҭ�?�@_~�Lo�Q��� ��@-ztF�H`��rY
��d	İ��)=���⚀����$E��a
\��*](��'�t�4DL�Yogߔ���&C�����s��J��_	�z|`��	p�P<��]2Z���`e�/� �Q�n��4>;�b��a?�O��L��@��[�xG� �R�=Q�I%�j�,qˠ��#��_i���>ex�{��X��
�{r�lS�I����1��k��P�蒊^/�whL���:� �����4�X����dm���n��z�`���� �ҍ�D��;��82��%�AI�tYGk6xh�={�n���[�K�m��dn��j{�}�W6���<N�I^e���98������;D��u��I{���U�&�ƨA|"D�:�P}ݛ��B�~,�]Ă�w�u���)U���M��b�b3�Z���o�篂���X���_w�MT%]C�e���fd�1���o�1�_
D�.�a����f��j��k���)f��!�U�[X>�_B�̨�M�w@~���[���\�ZEm�Ez�+o�0@D6�)}׹�oTR�6�M�d45��VI����]�do���w��&�],�`�P8K����n���|�W�R�v��M��x��4�9o��z�+�~�3���avn�N�6d��9g��� sK��N��&>:/e�P�\y�LrP4տ��o��W��m�O����zQ)��e�P����\]�ϳ�Y��W�j�HKi�����E�%�a,?����s{��ma�GOױ,��z3����P��-��{e�3(�L��,>��J�m���4����:�� 5�P�C�n��_b�m����YE)��]��I��� X+���>��G����D9���$���o:����6�3��i�K� ^3�����"͔��d�E2qLF�C���oL_	�����~��Q,se�h�s�m;���ʛF�w[���2�o�k�ZI#��w����z��^���y�8�}��oQ㨺��l���8z>~,�m�+��w��>p����l.�>HY���B��To�/�/ig��a�̧�Kg>:eEU�֪�@'}vD馚H�*m����yE섏Ӥ܋]����+R;&�?����A��?�p��$|��xbL�;5u�"x�HU/�²��c��7K�G������E���$��-�m�V�m�y>*f�\}�^V� ��ʸ	�Z� g�C�9��y1�F֒�R��H�P�ڽ�C�*87i׷�P(�ǚC�t��O����i.t�����r�i�䔂/�TwU��G���"9��r�y��>-T"������v��v(���,����Lf���)i�/�z%"KL�u'����Wi :!��qCA���ϵ�y0̛���t���C��JEα"	d��w��=]��H���4 �8�P�o�&���� t� h��9�ʜ��,`�*Kr&AT�$�1��)�:5#{ip*2���������Da3���s����@��Q���1S���-+��E�_�����j*8����ݽ�Ƕ��Dy�w̶ӯ�sL�k0Տ�&-�R�$A$��e�ʓ��j�MQZ�a�f�+����3O<�U�_�H�
Au���Cx@�� ��<�FӜ*! ��gI��nW���Rl��	�w���{�"�L���ݭaW�u�]D���jdT�s��u�*l��{u�[$4P;/.�(4��	�1xׁGX\����<-�:(��8`{T�f&�K;A*%T����b�ދ��N�>�	�Ud6"O�NO�#LX�<�Z��:hlZ���#+��|�&��$?��z��:�5���U0t%~)t��*S_k����ꯒ�{���z��@� Rt ��<栙�+LNJ�`r�>�Sh�rQ�y�!U��jG�ow`V���f���� ;�+��)��4N��F�~t������ xMF�F��&�-�5HB���v��w4#��c�-+����OL�nt��	a�� <����e<тf�r�tH����jW��8��Q q��Z;��x�u�i����8����=n�O�&��'/b�o5.ړ�z&U:$_I���`x��<�j����W�n��,S}�W�����k���9�Y@<�ׂ������Z����d�O�]��t_��e���zP"�k6%1�� 	9'�2d�;���A9����VC��K�T��J����d�?㲗ӷ����N��Lٽv�!}kZ�I�[�;����	������c�������J��m`AV7����t�#�Ǩ�$�����xM�>�%򷎁�=-�㤁�Ԗ�PS�tːF,��x֤�Uzx�Ͼ���<:s�.uĝ��(���'�m�氋۲bt�w�8���tv=y�0�7��m)w�v��D�@0�r��
D���w�8�^�o��vm���!V�.|��)������JcM@���r�Od��^z_��J�tY�{���H�a`��'/y:N�[�U$t#���°W�5���3aX��k��ϡ�r�"T@�9�M�_��la�T~ ˣ��~�7R�rTh�詪�ga�f_P�L�2,�X�<FB�µ�{�%ڢ�9�]��mTB�ױ�FP����u?�x?6C"A��0����A	V1S�z���}�`��à����?@�x�Y��2LP����0aw���*�y�:����Ax�Gj�B�&V�,r"6i�f�j��@�1 1�z�� �E�UpݵT�i�A��H�g�a妑�\yc9JSQ����U�c��Jg����*n;����`9�!�s����������)��2'1ա��<tS�g ~��?2W�,�~VFKl$��6�P�tq@�P҄+#v�Ҵ��f���J�kY�ᖨفDl��ܼI���J{�k���P����3��A��SS����F[�$9vFu^Mh�������[�Ӛ��#Ie���w��c9]W��vP�g��`}�%֗u�&���8pդLFUݚ(&���V]O��&��j�ll�HfSA��ce���tO����� 7���[��������գ�ܱ'áG�$ݗ ���^����?��ql�F�
*�����YT��C�d7|�g�n���O��aϞ�a	�# �ۓ�OSr��&�̑@�\D�8��q#Gt���#b���12J��\�q�-w
�8�w�7�##+���t~��q�A^𑋋nT�ϊ�х), v�E.aV�H�M�΃Pf�]��7{_t��8U</7x��Aâuvq�O�w���k4Lґ&7��	/<���C6Jb�5\֊2d%8�)\w��
��޾8T��:+Hʝ���af���SuF�����U<qO��؊��wPM"w��+4jT���0D��l)����!1	����B�B�y��#jp���7C�Hf��4�����$I}La��	D$�gx}/Ӱ��g�"��$gb�D�O"�U�M��/Ǚ�Q�p�\�:+�^{�g�d�/��(4�tY���gL�q�n=�c3i)�n���{`��޴2�$��0�6����߮?P���A��<7�A~�&:%��[{אzi��`x.�ʡ;֓�T�̩����{&\IOM��twz �7���5���f���n�_<1���KQ��[cD�Ъ�JSs��I�1�ܲ5������_�	��:�O�ߤ'��]�Cg0�=��R�Xh^�;Y�fL1� ���=�]�/�&�%����0���i7�ho�q�Y����������.�ޑ��$�B`��.<ūG`^X������8_1'D��L�������Qۅ�B���4��h�͋�@S|S��𙉃:,}�.�)��\zz�֢Z�jMW�P3����O2��-D��i�8xf�GW��h{I�XT&7��9���������MV	�.m��Y-���w�d�[��(ߏ$�D�Iڈ��M�T`eZ{��@#rߥ������_�өoyu|���Z8��躕�Lj�	W-D�G���{����35>�˧�_ �8E�j��-t��O�Er�!ק�¿��3"@c];V�B�>�Y��&�p�'�69�b	_b�0s�3c���t�����A�56m�a��/����x���C��tӥ?t����V��F����g�,Oٹ裓�Z�`_V�~oQ���Y|-��D��
^�B���H�B�Y�}R=,So�6J�7��KM���,���ݕ[��"J��&d� v�$9$����	�C�]MwÕLnZr�R��Ҽ�hVC�*���
.�u���0��H�k�j�M�Ҝ�=
z����<�p�ّ�
�e��R�t�ne�HA�������6G+P,4�-c'�Mr�"��ya�6-���Խ���	�-��N��\��9o�Gcp�������l)	ۆk8w���Sl-��0ExJn�dKp���d��򿳣����ʺ�	���<��(�
��ixeѾ�f7aon���Xj�	J�#�Go��Ƥ�$�5_(�>+J�^l�^��G=��r��@�`�G�(�<d����X�]�1��0P�}���N�bHA�mI�ށ�/YlN�I�>�#���2jUM�&�Jtl�����NH�B�3`��ᶌ�m)�����m,,	 ���C�q����"����<-Z�yDT����^ɽ\�lǢ"3����M^�Qu�l!�,���< �
G�@��i��O;�N��"��g��w<��8i3��mP��^�B���n١�y�ϻ�&�e�ǲ��4[~����ѽ��"W��Z?k��T�^�1@5���kߒP�+W����vB�ހԩ��{��a49oդ�,q��� C�1��$l�%K���=`�"lX��DpN�R7ɭ��][Jqow-��JK�/T/����xl�	L�D��ݛ�K
\ָZ����&�BI����,���A�7��S}^�U�T8�g����D9�w=�
�F���6�u���F��^�Z�=���F�5)=��
k����_俔߀b,��:�(Hb��h�+��aY�O}A�t���J�.�d��>g��srΆ���v��91���n��{г�,
�����Ad�j�YՃ#d��:���`��O�`),2��M1�J�5��  �@0�����*��ƿh���_dK�V�4�[PF���y؀`�������"�}FS��&�q��Xd�!���Է�QG�EZ�<Ch~p��GMρ��5�)�����ƀZ?|���pvUQ�a�oGw]�@G>j�+����G�zYfa]�5��5~�[*X-h�f¤����_AD<Du��ݪ���c:
�!���"��ʷ<f@Y��|xz&��Ks���y��O�B��pu���@ci�O�Y�+��ü�Bk�D��A��s�%���x:
�����ic���P��!_�Y��D��~QC��Y@�,�n.;�;�S�]��h&B�,�1����4�gL�G�tRǋx|��wzݢn><�f%�~�{�9�������d�+�<j�l�I�6�?~���~(���5��UK?��ʮ�\���6��I=��jsIpPtj�R�����"��*�g3{���EK?��	���;�,��h~tD���g�� ���N��+���&��Qc�� l5�|�y�3�w9f��g��sn�l5YK��|���F����'���0�y�%�	U]��X��7�3�R�����+-�-��˥�-�M��bߞ�'?�f��[`ٱu�z23�(=,�e�`�)���p5�Y�b��-���o-Ø����~���n���㽕�ZF�Z	��N0�ɢ��q��Nȧ�DB[=,�ѐvγ� �̽lc|nC��>hH�Rz��)�e���l�ƴv��_�ځ�m~�t���rt7�E?]�y�9�z{H��<��X�`&]2�ׄ$:�J��.{���6t�1�C=	\zJڻ�pBd�w(����I�[�k��������+|ST`����]�p�Z�@��ƙXP~seh�����F�Oz�N%���4�a��bo]��S�r⚜}�E�[�G��6>���2�3����a3�
8�Q������:���Hn-VR0h�T��1�ت@~�D���1��Ἀ�`��h��ͣ�Gt�a�ZL�p���5�^3XBAl�TlTO��~=�N�vc��Рߓk�����S~8�?;%d����������Ӹ�!�[ZM$t�b�K��q��1}��d�O�9����}��d�0{v�ϣKz����0.��g���X	ĭ�Q�[������#,�ܒ�`���>%���?D�cZ����[�� p(/\�L����{傎]���ټ�,�һ���E�JE$3#='-n(�K租;D�$j��̈�/�y'6��5��/�K}5�P@H@+9#��O��A��u�h�mL~�UڃϦ��y� �/��H�f��r��aÝ��6fh��VK�&���3I�O��e�$c�"j���Xn��L]��D�JE	h�3Бo?1��-���f���8mV�Om���d+pu��(�|b9�c�]�?��\Z'C�M�����G);���8[�p�b�/�Iw��O�PO}jq8c-iq��4(���f^�D9m�Ԕm#�t�VZ�yQ'��h�g3U@��
���8���8%4.qT��՟�.�M��h�v�=�B�����I��^X��I�$����F�_Y ��%$}^��h:y_�F�SM=��8�t!�0|�-�q�e�����{�K��b~���s���k����R}"b���	Px�����џ�(�CsC�����%J�������ωܶ�S��P���l{��lQ�@'=�i��'�`r ⤁�:�ؽ޴���o��������l(�B7�	c��t)0-��D5���:@����c;��¥�<�¬p	 @u�gr_�|�m�O`{b���j��!�Ū]h�
�������s������'�؊j��t���g��^v��V�`�d�<�n�ч��c��[D���:)��]��c�?� ��ц��"
U�T��0�׹�v!_%@��̏j���x���9�Z?�ᵃ'������^�>b?Ð�Pl]( m{wb�E�̡C��ֆ�aZM�L��S�,)r����K癨S�\�`l��l! ����d:6?�)��R�(�Z+%��:/&��<a���1�a#3w{@?����d4U@5�~0���1��%�/G�;��1o���2��N�u!5��vo��[�zHiu.Y�}YN@��BY���6P�i�*�6�9�Y_�[�KUUl�c���|?���8���k���#V]��	���&�[٘����vvn��v��N:�K�F���lF;<��ohX���4�;�#~�2���5R|c��(l��P����C�Ņ���iN�s��B�eI;��.!9|
̯�o^��.���vO^t���ք=������6]`	��dP�9gY�F��xkt��g�H�Wx���e��)2S��k݋��Ўc�ӈ(5e�ḡ��:0���a� ��B v��B ��`�u��O���}�(te�(���^D��kZB a͢HB���Y:����P൮U�wAZR�:/2�3�����Y�'a	>M�C�/����S�Z1n�B�u�'��%�+���D����ɶ��t�޼��5L]q�qM~���T�	"��w�����9|��bPJ(��w���2��QG����R.-b�#Fp�q,Y���]r
��_1�GJ� 0��%�g�Q]s�\��#Ak��l�W��Y����㯯��?Z���Y�d�����n��6�_m���G.��?]\�w�>8��cC���J��`~��Ļ�BOe!�Q~���/Zp(�?o��\����TZi���T��QE�������mtyx=������GIc�_�l�6,� t�T���7LFR�{�J��W8��΁��O�ܱǵ����ډ��Kq���>4�_W>�ſ�����8o��$x)���u9��J�5����<��+��>��.���`d��d�=K�n� �	��lXybo��~8J�=�w��"��'��+"��@��	.l�&l�5<p{����~G����Y�nE'��+9��.�A�3�����@�qb�5��R�$.�ʈ��R{ܴ����D�����^�XMǣ����>$�J�ű�B�H��3�.����Q��ޥR��;i��gB넞��䶶���֊7$�)V��ȩ�D4e:��|� ��M;� ��%wc6kzlx�?~�2��Bk�{8m��6��`�\��Ӂ,�(3�f�����5�����n��,=�<W�zb�#t-�4({�G�I�rR�F���Ƚ3�
ߏki��C��yԹ��9�ۭs�l0t�z�*�*s�ۨ����?n�r}O�#PZ��~�������P�zٶ��%�
��e�wv��w� ���`x:��$���W�\N<#�O�1��0N�ʓ��iuۊ�cB�{>Ϻ�����"���P��&>�+��rHon�o�7~�- ���τ����hc�QP�J	B��_�k��)(>��tYJ�bn$'�2�����+�����2�h�����Es�?ñ7A�� �m%V!������ݍ��սE:?��I1#���!4���EkoK�m���CZx.%���R�H��(��S�O_��L<��lp3��5A��XJ�a��,bf��yb�S����,�/7˴����n�ݛB�;uΆ��KY1�RS��
���ih�
UC����?�n�R��Nn��|F͹��4���/*}x���6>��-�'{h?N2��τ���7�����f�0�.���n���n��H�|�֭�9)!:��r_w�������$m,��z�Y57�������ly�q��b�}�����VC����`��?��O�݄�#�Z�x}�}����aoi�L���������i�?8�б�{}:�y�_Ó�9j�j�Ez/t���U���j������+������$5z���o"����.����_~,�S[��k�:D��V8ƶ��LD�O`��
w��U�<�T��J��>t��(`&�ث�emWpH���'�6k#���^��/��UO/dM�w3��5�:,q=�׎fR�����X0��"#4�2ݞ@����+���o<���J?+٦�AC#��d�jN!���GNrdҼ���n�Ҷ��(��7?����
���c0����#ﮩ-�<�4��3�0�t/�f �{<�La��B��T2���Hԉ�/�YT݈oܔ���zU4�yj�_������������g���	Nv���W$c��n����7�7�܄�2�*�Z��a�0��;��/f������;����6�p��<� �D�^Y������_��3���D�
�E|ѐ�xg%��۫��u���/��\����u�E�r�1"�[��љ�wE��A���x8i#9:w��l_Еw��:?;7V���ѡ*��	@���^f氖Bx��]���~H���r�	\N�{��|Ќ�d�^6
Z�%��Y��!s�n\�|MF�Q}p7�6Z^��ɣ�g�3!Cyw"w�)�`�#gAjd�X��j�g��L׷��>:�S��J��.+ݚ�r��ъ���Q��9�p�l��?Sj:�7�Ȭ`U�n7g�B�s�����VN�J�a�+;[L��ȧ����Kg�1�i=
ˤ!��++��E�{�F����~)�[uo�r�HG%�17���4�b�񏫖�^��_�t�G���G�KLv�D�kS,���:I��>�M	8>EJ���2��?q�q6T-���I��IB&�lO��@�"�Nih����+�x�UMXa�W�p���_w͖X��U���5-=�#�1�j�m��Zߘj1<���������(���	�����������=�����un���jU7��[d��8���n����'[tg���ubۼ7���i=V|���G��a���������(oO��Bܐ���I�Q{"Y�]T^��3~(����Hi��n�$K@ ;?��J��~��/�8�Q���|1�a�^~ʯĄ #���0�|�j�L������������*,yk脿�e�el�H���C ��!~9 zgQИlJ�iW�<���"�˥W����A�ׯN��7г�� ���D�]V�{r��48�U],��l��[�D)��TO�3�c�Lfq[A���8�z��U�&�? 5��<ڬ��6!WBU}>�e>M���N.p*b��#^ʛ}v�-�1Miʵ���a8��B�RA�h�5t���V�<��`ؠ��3��'�;��ȃA���.Dꮐ;T�r�M����`GX��pQ9�lZuP#�G�̩�,��{���6�w$�RG��Ѧ��z�\L�Y�������p(���̬.�a_Nj0ٱq�IQ��Pq�&�KU7f��Ӱ���y+d�Z��9uw��j��f�{�P�eډf�Ni����DB
�]j��b;{d����:Z7J~�#�	������)�o�zq�����(����L�������y�c=>d>� �p��y��������mƄз]�� M��g��d0t7������N��	!R�������D�ҹ:��'n������B��`��1�k�Bw>�X�cg,dp)R{�OU%0{{���Y�ȣ��i����]Ð�dc��a��I�����ѥB�ŀv1y�:au���3-8z�Ig��1��cX���O��:c6:xOT��N:�裴j��U��r�w��D�C)��?мsN˧i/.�S �/&�ay'��_A�a<�$j"�{��嗑�3����2H*�݊]�c��w�CD/m�So1���g��2څ��u�>�w�ו����'�RW��A��zd�߯���`�pn�v#�4���|���ׄ��b�iq�����JY�:h�W�����J-_Qѧ)Hz[O���wѼ��݃�B�+U�R�z�;t(g�6+Ð��UOb��=�����#A��e��ɬ�����T����$�Z����m$/���2���Q&E�f��:�>���-��L���8���`;�����f{�U>���@�@:�/a�|�y�4*[�|ŀ�j�l��&&��''ʛ�X��*�޶:7����g�GW�?�v��)����5��:˞F�T6���a@l�����C�	������PJ�ɡ���;4V�4� `�=M�!�?R�e�E��X�c�t{U��e��C�)U/w
?lLd$є�}��f�1���^��S���5��`-������Z��6H���/m�#L䣜����B u���	}(~��<>��8*X�;��j��7Z������ /s����z���h-7���d�`��n�c� G�Ȏ�e���b,��'�`�Hh��? g���ƀ+��vz;��f�GL�E�nM������̯�a7)`#�9��>MY��=7?F���~2�44r�VLv9G��m�ݵ��}�?�N�����KPT{"��T�o@.�*ks	i��8�3fX����뾣���@c���dsf���Ј�l>*�.A��Z�����@�q{ړ0�DG�z�~�ԭ5�$Z${����\r�9��$��q��2�s<x���R-n����Aus��g�;��o�,jg��.G�*e��pNڥ�Ǿ6��j�4xnjw��I�c��
(1��9�{�O-���+�ƝZG��Y7�E�kM^=���L�������@�d����B�Bya �<���cG�F��!���]"� ���Tmw)��<��FG�:@�Z$½����uj|��ڼAU�R�ӕ����8?fYY#������/ ���ϴ�?�OB�+�VZ3�?�+���~e��HG��!��\Ms��f�ʅ�EMI��K�݈�p2��_��Kg�oVQ�[�la��x}�[���H�̘�B�&�I���%"�v�x�$�WHn�]���	Ö(���G����rY,�߯ʎ~� _Cb^#l�q�t��
?�BP���~�lžݙ�����q�75h�1�>���R��3!��W�/�yqՒoYv��A����<F�ƥ=�Q���晊G����EJ����,y�,m���iF'��@q[���@��g��%P��׃���ڿ�0\�|�N�	T��7�8}@��:,QRtƃ�{��G���R��K��Թ�7Rk�6�R�7�Ct�&�s۱H����t�4$�8��z���1+��s���^9ܳ`$j�T����M���]̠�.EN-�����C@��v�H�e�2DŅ�ј�h���
�����"MY,�Y�v��g�+ve�p��q���T �����py��0|�L�2=���|�Ul���X�����>"=HN��}���������b�����r����r����m�䨭.�����j�ǄvM�����ꮄw7��@� ��aq��ŏ-��T��zuX�;��3]��&?�m������v�P۱�Y^�h�B(���Q
��}/�7�+UX/�(o&(�K\�22�/b.�Bc�I{!˺��S����	�Z���m�����+PM�=���F5�:: 
�0�7�]�vĲ^�m0D��(Y*���r�[	v��E��4��0���E_�(�;ݓ�S^���uF��r�n��q�A�Fw`ą���m4n�ߍN�=��ml"�,�U�4V��I�9�����J6z�
��(�'#��H��'Ɔ���`f��SCǯ��Q�J*2\��Y-!P�>Đi�߻C@�	�{�Ŕ��>�0pz�|�����Y��#�a��j":���
}�je/��[��@CwQ@q�"jM p�K���h�$��Y�i��5����b����R#W�(穎� �Kl�ybb�f���K��:��}�f�z�X��}��i��R��o�Ɗ��DhWoz��I��D����K	�0"P������>��'����s"u���2��{_]z�h���
^ ��ė\�A)n�����R@�p����RL�l�%����X�tҚ[P���� f�J0>{3z��N�'�:b��27�>Yë��R�*�FS�$��aO�18�0�\�9L�%Y�j��nHYN]8�]+��of�!��H��;J ���J�Zǹ���tꈖK`����'���!B7s�W�>爇�f/l��7�|��97��xg��,.H
ji�>K �ӜWO�3"���p@ҥ��k�t���g�"�ͺ�Őg��Q�W�1P�]�hlACR(�͢��m�1��sy�Xj/�=?<���\�Џ�G�@8��t~��1����9 xi��BL-v
�o�^��.���G��l��	��x9ٍ1�PL�G���s��F�ӴE��ě�� s����T8�wz�����kQ�o|�s��#f�5�%��F�!GG�x��2�,���E�e�'�6���9�iW��p�`:F[����/����X����y-ǽG�:� }XXk�@�<R�~Y��������c�3a!��:�q̜x8�"�}�:�:�h�@��w�g�9/v1�"T�H�h��CZCIG��d�aG|���k��>���?���{�#؄	Q/5���z�>��m�kw�D��5AJ�g$���j~K~�j��љ��'�7L5���#�۝�*�Hl	�����h��<C���m�&v����V���VX����uG��z��ϒ�����X�,�.�w�����۳��z"�D��^\N�(i� ���ũtdQGP��Z3�����_����כ)�v�#~��)��_����u���-(N�k�Q�����%��r��*�(r�CH�z�5���2ۀ9��#�i}0K����ֆ䔕G�}l
�:��On 
k���Xh�[���`�~�ѩ��&�#��&>��+L���lZ4�f�:ζ��u:����|9���F����A��1��cV����M�����_��(U靫t��q}�9��
����j���3�����$x��n�-��
�g��	~,&)��J���""U���s����5��y��Q|S���ɖ�!Vq��M0`a"���V�ZS:/��!�ƭ�Lbk#�1�XE7Nj��ktbc�dl����,��m�	<��h`5^���Gq!v�!�i��\3������w=� ����/���m(+���-����`�0�Jk��h^�OB�U�V�����04�[����ƼIV�H�x��Ѕ&��{�Jz�D;��u��������۟M�����<��6�@����"��nmin,�>r�W�ެ����]���@��\�%"炽'��A�5��0�5{8�=H%$���	av%��Q.ھ�̒��y�+ꉃ�0���֫���Q3#�>e���;s^��&�&�D��(�V�p�v(�頻F�Ӭ�|�>���?��b��~ZP����_[دg����XC'�JJ� T�|��A��]��rA����愔��s�<{:²!�n#�r�Ս�!�AѾ%���c�͛�LC\����E��k0��x'�����u�2𢭋�d���������O�q�<R�y��.���xaYӃ���C�up�nZ�r��}�6��j�M���}�>A�//�F�Q1ֽD����4+�b��HW��=�?n��o�Ք<#��a�����6�	dFos���5�M
�m �6��A6��X'��t��R&��,�(�@�^Cj�:��Q�Fޗ� G��G$!�je�߽6$�q�)M�
o�WP����Q'��yNX�6$�<gf��W��4��)������o���k�tŬ�\R_$\�f}��p
(�)c�l�AS"Q7����@��v��ߤB���l+��Hx�1�]0%)<��l,X\�U4��y؛Bhc@��'LN.��,�+����C���D�&*��M�}��ވ��BϢM��^��67�5�~'D��W��[A�B�g�=J�L��i�L�'B�^������D��t�$:�l͡��怽`����>&����(4h�;s��ǨҲ���a1ʮ��t�i�u����!D��E�
�<^	�m���CF��<�N*� �ظ`!Y����Z\��=�ي����ي�~.+�,��( 9�=���H
�#�kɈ�g�b@��d��k��6N�1��ʈ���G�G��78F�?Չ¤ˍ�w��~��wY5���[��2�1��Z�(N(�(=����l�'��ױ���"�T%�9�����U=*�'CY��F��g>z[���Y��b��,U��\Dʽ8q0U�,fB��GE�����1���*�+X�����ܗ�̙aN�h����`��Gv�x�
��>�rP>*a�&���Y� ���Rh={ڲ@�\bȲ*Q�o%0A�ۄ{,��o�VX���H�_�R}��&�s6"�q��o����n���* ��T�,"�g/��U2�xL�p@���Z�|���Y��/C���7s�9�L��-��w7p@��Q�ap���G!���3V�ڜKRN�Z|���2�����]�H6w٬4���G~�(�@��J'��s��"g`K�ڣ�PU#���%�I�}"�i�w�[��	 �AD���M���?a��/��J�g�Hz
��ƃ�l�4����g�U�w���g����8a��4 �W�	f�h���I��������`,��ڕ��veo�՘N��Tq�,bKI^P��đ6rJ��-����I�s�������4�li�w��������c�D�Q��K!1L��\w�n8&ѿ�;m#
e�D��{�1ޘ��'C�� /�*m�*�vd��l�~��#1|M<y'}��ܼ$4��:u��,��݀�J�d��RVN��x>1퓡PYl�:&���,&�|��hz/� ��tPp���XqM�����p�K�A�b=��M;�����u�o�~��&�f��o4M	:�q�ͦ)K���9�Κ&�r4d�,�,
b�yE�K6 �ȷT�(Ы�<�x��55,��U�[��ó4y�����܋1�"��Cـ�Y�T80�����;���3������e?�����d�cĀs�"�u0FH�Hk�皨leNzzm[�U>�|��oN[F^��d�����,�ҥ,���"�B�7�y��#��i�[��@�d�4�'�5HBk�I�zp�ͺ_�T����m��#>L5f��ϓj?Ij0���Rn"�	�u�<���lPK�b�%�2Ԧ��i�'5�X,���M��56�"I�SG�_�Y��z���ξ3-�Rn�U�A�]�J@�}-xv��-,��	׊5&��-��'$�~�ʿ������h�8��������jsn5+Wf���
�H��]zP:�K��黇pM��,n�ܔ��_�lH�3lNAxO
���I�k�-ݨ�t��D*�C6�Qm4�c�a��j�A�Uxr�ʒ�����5��]-i��o}W@����u�z��;85�����gV�
��\$��We{G[���6�A��k^M}`S�:�#ϻ���\N������F~�u1@,e�	I��K�A1���6�dࣤВ5�[���i�W�&���J�ZݮGҝ�S�A@�
H�}V�eRǶҿ 	��6J�����ryZ.�j�v�A2�%0�@Ġ�47y�ƮY�B���d#C�8E�#l�>�!�`�A��:^mwKg)xT��S��A�0�|�JS��#���V�) ��@y_Pk����Z�(fZfi����v�4uNĥ��ݲޘ��/7,��P�]�������޻3ub�)�2��Q���l��Ӯ���~����$J��,��h� �q�j΅�>�r�����d�W��t��<�r�f,�˘v��u�=&��u+�9C׊��]���.m����U��<\D���56�k[_bIŽ!���!sa653�\zb����AAx��찔2`��i�̷J��N��C̭İ��YɏߺG�]�H	�.�@��������mCp�@�47e&���29CS!u�+m��s����:CM���[c�s4Y07��'���̬Q�(Q�hy���U	�f���@�q��q����j�z��.�{ҕ�-s�ծt� ����E��]E�%�R�k^���60�V�D,+�M�<��)廣�-��$(o��A�6��yc]�-C^Y�8Xzf
M�g�F���r�+`Cap����*�s�wxsz�W�_Y��fl�r��oM=�����xs���Əg�ƑWZ��!���*����⫏M%ΘNde�޼ �gI@���u��I�Fq"�$�)�Iq��*�6\����Zu�wl� ��y3�ahk�>c��NU���y�DS`��%!Y�uꢫJ��?���@6������h��猡�K�%�����)�g��D�����8F@������Uん�����oOSM�ǔyqN.j��0t|����;u���h�Z@���Y���_������S��YE����$ĺEG�06�N��!_�e�$ھRi�A�փF[��79/E��͠fEN`Y4�&mH���jn����zV%݁M��tQ�HuqnA4^�Ur9���V�S�{o��o���1�>B
���K�	�=u��N�km�N����C�1�뼨��y��ROd��?�2�p��1�R�.�$�U��9�����\3�%��B��ڃ}X�+���sm`4��M��>����|,�k����1��=���'��l�,��c�0L�Vh1�0H/�y���{�)�-I�ȰsYS,�A<i�1��#&����<D����MnX)r��$�aKܧ���į�G���|�c՛�/�pCh~��k��M�7���l��W�SV�(���;�{��?���C�·��]�fK�iؼM�K-����HԸ&>J��\�,��c��O!��j�*�����������y�r����h?�b�	.\kU-��S'l�����HBI&��Ƒ���(�j��1T���v�ߗ�76#�]�2�f
[�}=Bf��p��KB��[$�゚݂�r	d�;���!�^9}�>���������V!w�>SjȤ'�����(�SI�z Nۖ^.�4Ko�'�O�g�
?�z���"�V3|dv����Ȍ��8���f� ���\�$�-�~S�������>$�����u�����X��*�����̚-Yl�:N'�J(v�;)������ʛ��E=_��l���K���FL��yv
E#�q.Xp� �m��E3E���| C<c�l��{b����<J�����90��u{�aXB�����ڕ�嵝|�qUb�	�$#�5Ƒ��c�Z�xg�q�@萌@�EZ��4��ρF�Ƣ���'r�id��Ip�[o����Y]-φ#8��A�؀{�:�"d��Kd����r��.��6����"�)
Ś�or[(�����BD����Fn�C?U8g{H�&��{4�[��]�$�t�9T���I��f��)�L'�]�gh[X�������/�qo���+�\ �wF������z��Ʌ���=��-U�}�j>��$��h���Ĕ�*��n�VI`�>�#�����W̅�!�m쩎!����3c�����&=��9ҟ5�Y|�"H:�7T�Xre�/�8}u�7��(}<�g"���+e����Q�(��G����]$�`ħ��{>�@2�ߢ=h�L��Y;�.�
P����8�Z#��׮�|�i;�r@?��Y@uR�s�+���'6N�u�57��Di��q^|�W]z��-��{o�R:�[�Z���])�hxڷ��͓��(��t<#�E����*��8�.�{�S��0�c�:@ �C�P�5 �au%1 �����"���r����c4/6�筶�x���Cw�b�ן�x����A���z�}�ˮuF>�,N�mw2�orIm��l�o��8�a���d�hM���������+̩�҇Q�n�{�y���Q^&G��Α�1:����r݄*� ��=�+%a�.d����X��u�������]�3zQ�mn^���+��+t����\ꊳ��_��f%|��JB�r��W�l�{5ttT0��- s���2���m�3�4Y����Q�w�|@��aN8*I�}^���H0T��!\,F:/��vi�>D��(�N-��3�
��<��D-h�=�{�U���|�r6VL�.��ԩ��sѨ;�|�E��V_�X����<X������k�1�NB�r���
�"�R�ջ)��T�EX����wFq������1�a�z�ú�?��hfZS��RsT�_����	_	4d������vΠ� �#�<X�$������ꔷ�F��#ڕ&�6�p�?��~�1�;�T���d,jK��.��7jZ�I��/��-K�O��R��WK�hx;	˘�f���������bg�&֩�쯥O��U��ڤ����خ��/��<���Xl<�銹��[�Z�)Z�29tL��\���X���Da�e���A�������/5��j�����;��z]4�b]�+5�^�@z�r��Pt+�g�M����W�r�����6����}��+����e�!P��2z
�&�w�$��fhV��"�¾-�5VN���,�Xcq'�e�����g�4e�*��^.� n,��7F+zH�~)y���\�U�*�9@�S@��.	Ŵ�
۪��w�Kn�*�8")bA�G'�D�b{�p����;1]��_Tl����3�4�uc��c(z	w�W�O�>�(��.�_i@̔C���ů[�O�n�Ԧ�2���a�p~6�:|�|7j��&i�~m%�Lo��:�h�E/�r���#n&���cy-	�����k!��&�˵�y��7���EWa	��뿓5�%�k�3ȕ�|���rH_;��'��.5m���d`J(ة���oo����h����]�ɯM���"��������n���)�#���+-�ENS��6w�5کZ�n�;���Y��u� z^"�yd�z�c���a2[��n�S���ռ�zX7�{
	ڶ��z<��`�J��΋t���Ut!ľβ��W]K�g
�K�S�b���&���Ч #	OԩU���c���2�/��aѼt����ഘ�:���o�5k����f�˫�o��gd�Ю-�:��%m�3ɰJ/HD���R� %y�md��>.��_�/3�U������]1�Ìg����u�	V�諩�?c8W�叚K��؝j}ĺ�8v������N�ۜW#-��:�?��U!��ԑ�Z�$�<ELS�d7 2�Ɣ>-6avS�BE��m�i��
EU'u�`u�y���ȴ�˼\��\*H�݉F���Sܿ8�)�*��-����P��
+P��/�\�ԏ1����K���&�Vc���l�y`=���T��k�!�*ݥ��{XB`xq�o��������l[���3$�k�_�� �/z�a�feXl)�<���&��ʬ����� ����+��M�������i�!��ٲ��  5��$Z��8z,PL�
ޘ5��#4\f	O��wΎ7R�DPxD�߾OD�ģ�	� �"��{���8ǿ��}�
j�ݢ�Ryq���Ҁl��CM����!��V��UXva�H��Tc�W��!c�ѡ���vH���iU��x96�Q�j^a�	���H��B�Dk�Q�L,��}��aV�zN�qݏ�x>�"�p�S(�:����!�Q�;/S��
GO:!,���is+�o<��q�Z�%� ���"V�P6�c1u/�R��v9�W�����J]��vJ(�yC�D^�m�R"���a��0yĠ��EUGl;�!�%���|��[��ݧ_�>��:��,_[�A�>쭔4�臭G��O��m��"r\ej��z!�a�ཞF�(�o1س�v=���-	R��'zW�j&�6�Hە���`��䇎z�"�P-�JΕWX ��qL��A�����,5���"�ݩy�8����@�Xh����ζQ����6�ӳ��k�5o\l/4�C%B�cͩ�L�!W�#w�%`����Y�1mj��+K��\�k|���"�hL� �����O��%�����+)��m�`u����n+��o*�,"%�~*�T�K3qp
���w���O˳�7Ш�.�K��T>Gls�Y�6k��kF���1�}���{NSQ��&��T��Q�������欦��L칲���O&�ƒ��?��I��]�`�!�O6�)�F_b�UpP��t���6�Of��Z�j-B>�;�%4���,�8�������N�.�; ���'�m��$�.�ή��u��O�����U�U�D�i�!.��	x�6�޷X�G�]Noi}r�L����j��U�:��؀i.w������C�aKc'�5Bv�1���@e�w�V������V�C�q����	�~\�1l�s�۩idc��=�q%>M%Ț�pJ z3��'��ӽ�֍d #8_���1�����·��¦Ё
���H_��$k�����KdD���u���HU�ey*�FT�y�UC�r�9�ŷ{�]�,I�j�n�*Y�OϢR�8zlvq��7x�&B�����D���8���P�6Y#�>��A�V�Uz�sUD�����bi�J��i��q��m��E#�[a��	�V��E����gI�:I�8��>#�B���]+6��1�l�|�.���D�++\��_?v��mټ���S��U��i�*:��`�p��^�.��p <\*�)�!kf,���Nd\��W��Đ�1�8�k���1��z��˻�&��ʽ��a,�#���D�};^Y��5�� �&x�Uˮ{��P��s�{˚����{QXY\���EJO��Sn��i�.��cN�� p�t{@��� Z
L"��%1�bP\WHEU]%̆�� ��-Tq��o̯o�{>[C̩!Ƈ6~I�×`�_j}xW��f� #�癖ݸO�1B�䙗�z�U��
�ɜ�3$��G�W)�Â77�x��Z�L57h�9�a�JNW�!����1�@M�y�T#��������Y���&fM�`��m%I�jPs��U �~,�XBF:!ȴ�| �r뎋�I(�@Ptt�R�GB�\�L�+����2o�ȝ��W���?�:��J�=���d5*����p��`ۗ����{,�8c{�bK�����`\|Riw��k�r��aX��}�tw�
F��ÀaO'�����O~�ߣjHδ��bF���d�iq4an�W�`�*�v�!�5�a��S��*DnB�dn���"���i�����(��_G���z����9���`��N$�2̭���)�����V�3��˘�������/�2*��^��_�J{�U��|�Z]�J�_� j�Ll@�QY!�ͽr&����oxr;O�TrQS��vV��5��
���D���wC�r�k	�Bި��A��m:������%�ZZ������K�Cd,s�hk����� ���S�k�z݇��Krm�?|ȶ�1��P��2�^����<����ϩO�6E?�j$e�������޴�s�>S6&[-=@oi�YN)��i�:�u,VNĤ�$J���9�z%#�G�jlQHY��dD�s�!�m�z�l�a3W�;�C>�����vIQyG��g��T\��=�z<U�)��-H�g�]�Ml��OE����� ��"I�7���&�I�|Y/bXį��6�
���6js�#��]���%�6��`��=1,A,<�Ng��.8�q��%p�
��3�n�;�!�@�����'�;��~�Z�wwJ̉nq��Qf3̵�$���ͮ�̸�����#/�����M��N
�2ؒ}q�W������3�?��F�\�Օ��+��X��O��Z>�_�
kaq�&J�΋�\d<*P��Z*�?Q�Tt_�?��G�y08x�]�uŔ#���X{�)��3��F#�i���L��M����0����`��e�S9��8��Y[{�N��&,ϵ�&�A(o��"̻pva|����0��rq�#*pn<����ҮU?gC�A��@O��|�b�Ji����Dp�����m�>>�-����5��h�2��Q/�F�b�{<�a#>�:��<������Ay�� mA'����WLN����ao�!�u�'�����+RG~�M;��)��l+�1ͫ|_��Ϯyo�0'�JQZ���?Ο�x����"�٥�|���L��!���s=;DK��/�$��C�Jȁ�_T����/ ��\�ڶ9)��gt
��m�ٶ�F䣎c!����1s�M�ç$�z�pK�t�'��N#s9޾��iQ�f�.�GJ�eRd�X��X �FN���ΐ����E������'Uc'�R*�FC��,��W�P����;�Z���`�<{��\Η�!;��+�G�Ax	c@�,�.�(�S�$u����#�����60V"�w���0�za��=���!�s���M!$�<�a�rG����<�n�}Y������j��Oow#P�^��to�"��aq���+��g�y�9�iV�"��%�.<��5�YB��� �b�u3,��Z��s��	��0��kؚ��c��œ��<LE�jV�);/�Z@_\9�m{;|I���HoG
gx����1�+��^6i
6�vfz���	H�p�7��X��6�z�$��:z��%J�R\0Ǽ-�� Uy6?m��C|�#.6	�T�*l�í��WA�Sr��.�~��$�&��,�u���D��uy�|�Ԟ��@�X� R��V��[�	��<aj_�eh�b=]{=Ա��BW����P�r`K�j���1YUzu��� ����~?cFϡ5��
���BFۡ[,��xӐCT�q�?o�R�8�S�T�G�����7�(�a�/���Ȅ��Ӎ	�0�Dt�d��W�	&PYVT���L��n��_�h�lb�.w�mb>�_�ֺ��b�F��w��,�&�����G`2�����'�� r/z��ٌO��]�a5�mvD$���G#U��g��]ѩ�j��@(>T����/��h�$����w ����D��7]U5Ke����.�Z�c-<���Nu���ޝ�H�5|�0T�U.3q��rڷH� �ج?��MHJ� ��(Ġ�b�l�5�gDڢ�6*���,K�9�S��dx34�QUcz�R�k�eIWs���'���&�T|�0/�D��iv�A�XШ�|)���>�Ӑ��cDUiq���,�g�k�E
|\��K���v-3��׉4^���Ee��;l|�5JM}֫Md�����Ĥ1��2��~��	��Jq��v�z��Q`r�����-,R*u�����V�NGLt�G9��2�T�Ոs�}����]��LN�Q�+�$z��_�yC��>��axf��r�������>F�=�?�wu�$�	--rb�,jw�p��1N��ڽv�ה]TP?R��[G�0(r;�9X��Fᐼ��BV��z����F��q����`���GC[+�}v[�#�9�}0�pa���4�J³���[6'���u	�	��A�Q�g�`��z+��v�l�*TEP�t�s�[�e�V�]%�
�O՗���*;�1���X�n�7�%TKa�\���G�����?O8y��E�z4���4�I����l�n��JC{R����f��IF%�Jz�ߌV�����h����U�� ��A����ki�tnܑ'+�N�8�\#9���ˀՍ�O �OS.��+/�&�!�V0RTۦ�䷆��R(\!�9�����R�cs��J)���,�54��i�Ē1�M q�Dɀ�16��G!�y�|������oy޽��.�&�jGg� � ߛ+��H����ш��/��M����]sR~����U�C� �+</��\�r�e�]a�A�<������^H)��6Է��Ş<�<��0��@oY<��N#տ��9I^L�L��Y�=�9�C��.���_0�Q��$z(�'8d(������N����b� \:!����VN��F�!�.)AQf_K.f���-��/�F��d���Z�4�Й.n�����J����o	�P��^`M��6:l��)�y-�`�5�b����GU�1)+�L�b��V+��n�B����[E�-��X>��K�W/�l����KsA��z�8�H1�!Ei�,�W���5���>j�6����I��_�����(Ь������e
&1pƻ�el��e��ޭ`>�cqV-�9���Q�ݨ�S�E+* ��Z((6���W����D���z�Y[I�_-��ͽ�D8Z�d�|C�wPO���q��l�f}��ϕxw0�s8� 3>2�y�9�m���M�����[H`�<)J�Ŝ_��R�~�&�f/θ�`�}�by@ܐ�ٿ����
�}ۘF#�e�pN��a��$�7��a=ѻ�^�e!xHa�q<{�`x��N��<�����0��,�b��S6FZQz�zh����o���H��+����4�@�����,��o����}�s�%��g��:p��֗W�r��G	εΗ�}�;��*��K;��qk����[U���r�珐(���7@Ζ��+(�~6c��&���W0���@3i���F ��3��$��	��@m�4�a�0��f��m���֍8'6w`�W�L����:��'<��i8�M_�qe�F�n��>h��$��km�����/7�SY����)}�̙kK�?!�g�"���]��5l��q�g1���[��H�� �w��n���Uѳd籲��Wi�6&Kr�lͯ�4��z_��{���Տ?�Ψ"1R�����v�g�0�g�8�Y���;Mĳ��鷽1�/��K��7�z���C�A����_�4�W�S����|V2������9
?+��������i��!���MzU�����+���9�@�L)j|���r�S��Ty�g~��'�]�����B�$˙S^�7I�aD�
+���<��D��@��`=gJ��[��>�
�7��~���>�k��@Ĩ8憆��"��%u,\;J��c�(�0�Vb$���.dڿ��nQt�Qy�G`�VS�nuR N��@��F/g��n�qpM.j����R�0?�����f�:=XJ����$-���s/���W3&V{���h1#S�'�`��0R�.�V:�~�Y���c~B�����څXIx��a�ÓW*B�3�S)��3�3�kF_��|')���ka�����m� �v����3�t>y��N�y�I�J��Ӫ�!F�v3A�ʊ5���X����1N�n��j�Y�ޫ#�/,`�0�}*#neO����K|$��~�j�����ӿ��N����TA-���S۲���������O�G >�7��@�P�0r���b"��?��?�����z, �PA��X�ǝ���P�,ѳ twUޣ��۱�T
�X:��<58��%Q�	^kY�c+;W9\�u/�S�ا( U�S8+�s[��D�[�{��|��|"`_���/ei�J�����Q5��eUY�_y���IZ��ܠ4�񢞩�T	��M�����_$��_�V�(�� �g� ܿ(�â*p��i��r��q�$K��?�����D����DՖ�3�r�V�љRb������4��ۣ��3�	����<jo m�X@:.�P���gy�ޕ%�-m ��\&��5t�<u2>���4�F�[�q�7���$���.V _��]����Z8@[�0�=4Q
�@��׹pɴ����*gl��L*�.���?�D(��Zϔx���R������L��)��U_�G�)� �kώp��	0}��s.�u"�z�8}��Q�x� �Yt�t]�$'��9+�R�i�<dX-�!otw�oI���7��mt�E&�����Ύ�)��]m��%�*�K���c�ʒz~� 6��Y�>]�n�fx�pH,�#Ai۠����w>� ��F�H=	rz�"B蜴J;���@ڹ���l��*V��F$"�J5����QyZ|���`��]�&���Ku��Iun;z%{��#4�E�C0��$;��G`f�S�C佞Sf�xk:$�%f���m<d"�G��gG���kyS0>��b��� g��X"^��T�i�bT[F*��h5C���W���mO�>q�fE�h��8t�u�]��O
�	Z�>��p�6��aSza�%T��-�}���b<!��!S�OP��0;�7��s"�5�r��}WV�e��p�w���x ��`LLRxH���З��K
����``�TRn�*Q�6��9��0k�ʗA�%|�e��anԶ����8mth��a����x� $P��V�	!��HlX��#Zs��u�)	/JA��m�b��D=���h� A�My�w�L�uS�$҂�Ɉ(�%J�v)(|g0��{�f�V�nz�+��?N���ƀ�,>RY_���Nv��tͱE�yˡ��Zj��Ɵ����g]~Y����|���@�x[�LWT��{��9/ɐK���� ���[X�A=��v��ԑڡ�M��P�� (<?��A�_|x����?w��`d����b���1M�f�
Yk���?,q�{��p����
ٵ�Ӣ|��l�X/���A�d�A�){/B)D"���Vbp���Wٞu�����eH��Y���YU�G�f����� �7�gY�s]
�o���Py�@�{�a=䕶���[@M�g,�$
Gx[�)<����y��쑈��x
[���\k]T��Э�]��)n@�W��E+b�U�o���\��SZs�9�֐yA�y>�6�_>rpԱ0v5�@W���+���U��W�0}�2��"� �_P��~��?/K���E���_�'~B'���|� ��5�gD�e�:���sty^t0�>�\�`)]d]������1��W��R[o�؍����Ti�V����d�_ b��K�j]�F!��'��UJ6	Wd�m���3��(!Ʀ��S��'��M�#1�53\ɞW��o�������Po��u�YH�ͪ���/S��'�7W_Q9&��E#߱렘�Y����JVJ���nS�`j�.���\.xz�Q�2_bQ;�Ʉ�x�[�AO��I	��0L�����b�����۱�H1[L`*B�L��8~I�a�mnN�ዢ|�����u8�m�w��]����aT`�yktv�f����D�e�4R� ��^Q]�v����Re�a9�x����>�jaq�p�ꑭCZ5��$�� |��PVO��[S�#m�����h��ߠ$�_�1�?�����@��WQ'N;�K���mbY�@ u��w�Bs?�j�k�����*�k)�a|��.v���J;N�8֏������û��H8��q�X&�о%����w�x�&b]��Z�Y�k��&�����L��;1�^|��M�y�Aa2�s�a0m�
f�ڡn���衃��>L�k�\0'��X����D2�p�y��K4zu��#�Ef���b��FV/0�1��d��	_X��A��y��đ���?��Id��b�D�sw��.���|[��i�|͌�����!������y�TI��Ԗ5��𪇕(A�'��Ri?Lp���4�ĢA����Q�%�kra"�I��?ma>��Mc�<>i�1gX|]	9���М�b\r���R�Yw�Ӈ��0S��]&�����1�X��vS�ƊϏ=M��jG�ѝ�t��fj�Ҩ�_��_^E�[�~��B:;6I�m��r�����I�KwE�xԑR#)�B�Xa5)�����-c�f�Z��D�#-�+-�n���Ez�0��0�7��\(ae�������Fr�-��[v:��9�f5@�@S{ �`�j�*��H�(�6E;�uAR����Q�y��`�:�� /�d�~���H{�%���jGv4����Eѕ!f*����3���V�g��G�ݣ���2�����9'�O�ת)0_V6I��'&���v��\�q��r@J�ZQu�T�>س4�l3��N����/r��T�"��\�P����1���F��� ���g)���hkRd�I�.+H��J��#y�k�
�{�b0��^	��9>U��Z+싯�R�"���ʧ_��[��ٯ!I*�g�ig�-326�X��ҧV�����n�oLg6	��˼�{�2�v�'�5/��.��ٵw�EE�m�_�h��f\V�M�Lo�FjO���`k���_��q ��f�Cl����m�C��>�9	)Yn�eLzKY�
t���If�����
+/���� �����czS����	�߹�t6�t>N�t��h�@��"[�5��JFby��{o�����Q��
E�i��j�[��яS��d��Q��� ?����+�z�~T��ɣ��jdn��9~�n"��m-�ŕӻ���S��;R�n���8��uyצ��D�*��7����$�o��]��/��b��~gD�'��*Wt֊�0�d�B"���g�7g�HQ�����ʗ��Y�,%E�V3i>̖���}� |%�� �!\��lNht�Q��Я+�p�n�_o'�U���dV��@���=*v�<d+���x~(�P��.O�{�q��(=~v���S�d�;L:�7}���q��[[D��25�F��|��7+���P5{��TY�q����t����WvೖG�.���+~5�1�-_��^�̤�F�µ\O�a�3��v����p�`��т���V>�����(��rߞ�PD�p��[�-���ۂm�@���0u�;ɩ��
�M�d�8ݙ
-\J^�}�\Ȩ��5��(��RCv~���M�8X�����z��W��)��(�VQ�p�:h-J�"U�y�.��.b�u�P�)�ӱKqH�H���ɱ4�����T��n��k>��%�2Uk_��~��9���JrK�8�0���9UQ�#-ԋ�R,�)c��um0�9<��s�v�.��R��
�o�Z�w�k�0��f�gr���A�,����Z�_7a�Q�*ՠ��(��lh��i��@.���#O����D5�0�c �wf ����o�Wζ��"�Z.hR��6�T�}�PO�|-��y'Tx�H�1>�X���[�ƨ����r�>���3b���DQO�$[ ~]]�����B�b����
�ʋ�� V��Rm��j!B�!�\Ξ&����[�=2`�R�#/��Bk��R�&pb�+}�������a>�� X��K�@v76d�Z.��	T�ɣ���o�~���s(�B�0������-Xt�e5�E�Z��`�}I��7.�'�c�&Jy�b��zX�X�����^6�z�a$1^��^RL�z MKL���"=��`����8��Qvy��u�YT���2Z�ɂU��l��p+iZ>�����
�뼿�+c��FA���z��$= gUp�HN�C�efO�~�\��e��7���
��� z[m��Z앚yZҴ�Jƅ��"[�`�@�7�P����G�(my�Bo�
�3:��O��č/bk%�ř4-�X�b��,�8^���;\U>���'��x�bM*�2�� )��쉎 �}�a�//��N
W��d��_�t8�s���}@3��V�����~��ڿ�~MC�5vI$�W�t�RDg�`y1�T���!��fa 'Q���T)��/7�O�.|;Ԝ��4�LU!�:�ਧZt���KL@KЛM�L`mҌ_[1�`�8�^��Q�i��ᓕ���0�v��^*�L�a,Ce&�����آ!ɼ�����;	���f�鵃D���p�XuN�py'�M(���:�lx%\4ɐX��[P@��y[?�1;6\U4�(Qq�Ŕ|�"��O��g$;��Uq���/U���nfQ�o3�={�ڼ�i��*[�v�ñ�pNL~�����0��R�m,��U*�YfGs���j���>�eY�
]DHO�7�]��Vi�k�e���Vd0S�P����衡�Pg�p��D�^��6�P�T���W��6���e�lBA��{Y���y���?f��
��Q�Eo����.p�����#�I�㪐��ǵGO=Y}%�����~1a	������6Ƒ����W�/��9e4I��NӮ��v|�:^�E�׫�r�n��X���GU�S��v%�qVw
����N%�݅�����5��$�gTma��L㮷�y-i�c���1&F[/K9�asu��q%'��"�"	�z���E��F�\Q�tJc��;�x:[ ����k���@q�.!yg�)�s�b/�������T2���$�ޘ�#�����q
%ܮj���`z|2l�P����+���(2RG�[�����tx�B)�|����b�N����ƎKܩ��V|=27�M�/B��`l�>JF_�,��X_�����o�J���l�������4����p�S8I�gP`*ōǶ�D�y�
�cd��|u1n�i�3Sǌh�:T����r��\)�j�<�K)u�o�����'����OO�J�l[����˽6Jo���Z�n�A\U�]�G�9�vIv�|��P^��)\FWt0|6ڬ�K� �pw�2���U��=�臆_���F��Æ��S>r!Stxc�f2�^ "��2���U���5��BU6q�kn�M5i��ƌr9�<��$1�F��+U��Q�#��ŭ��7j��nz�Nu���TTC��5莯�m`Ew�!��l!��~̀�hM��_��H��k�'O�Y߆4=>��<�Qm2��}�B�wލ2��"�F�D�ڞ���sQ?���_��>H�+'q������!�.M��w�S�Y��MN9z+��yfl�{s[��m��Z�&١�S��� ��uU�OՒ�[xl�n<����[|6C��fdO���M����U���g��x�eZf|����S����b�4Rs���
'L�"���b��%���M�=\���K�kz�;�-#�9'�w�D��fŀ���\���/Hs�Z� �
�����d�EyL�uXL[���H��Se�}�������ѻ��Ӯ z9#eosϺ�Dsg��Z�e�+nN�� �n��:Y���DJg�O�X����������A�ƥ¥�gW��r�5�u�[x�����g�Ｊ_'Y.�8E�=���+�vy@�[L��t�7vn��\�~��*j��1H��Oz}�ӫ
�s��[��vV	ԥ)E��3�%�ڷM_�t���
Ɓ�<�Tԛ갽��:9V�y7UJI\��LO$�����.���ǜ]��eW�M�XiX�������PG���TܦH/���5��KH���ֵ��b�vb�bZ>��2+vf�BQ�!�A݁u�c+km��Ȧ��6Jfm�`��QXG�5�x�:�~��5�˖HH�JF����5AF<#I�E<���0
m��@���~V��>e���ٕ��t煹���֦+/��Y�ˇ��CS����gVa5#-:ۋ���4���L�+�N��x��	��+��¤����"B�nx�F���E��8�Ji�쨗|��qX'� |w�^!����>'��N�P��i��cز׍�k�Q�#��H[qާ��Qf���W��/]߉щ+�=�3!�Z/��X����چ3�ɖ%�"G<���r������v�u:�f˙'G4�J�3xC3�n�h{��ǥ�.�Fu6E�hj��3��qP�6SW��L�XS}�'&����l?�r��t?m�3���9�./s��ȶ���Ә��siuOج��gs�a+'� 3��&��׈������mc����E�6� (TKϏds�}��<���<�'9�B] C�E�&�7�q�^6��tg���R
��o�H�_��8<���n~$]����`hu��qW���Sr����d3��WB�F��
vL,x��4�p�h��Op
���"���t�F�R��$pIJ,�)!���{�A�����5�x,�ڒQ�K2�2G����9��١;��^H������o�����Z��T�d]O����8j������^	'��7~$��XN���1�����AA��р��3�=r�Q����hdZRf�Z�P/�VMC9����z��e����ڔɊ�B=��*N�R��>PҌ�����c��$��Q�wx��s#V���[-ږ{T
��f	̻b"����8�V��C�)(}F���&�|���l�E�����f"d���3�+$��#�j�tS�� ��rTC��1
֯$�Nˮ�ߎ(���r�����I�0�֍??��K��V��l����8d�,Ј+Y!F"������!�+�ʩќ r8Y#��*&�{7>�n���R�uI�ͭM��3p�An%#A
Fv=�g]��X��e�;��bU��`w]\7���p	s����s]\W�t�zn�B�G�n���ӏ�X���@����Q��"�Vul;�g�O� ��'���Ii�]O>'1@R�[K:4~u�p\@�9�!�LaaS|8�Mޡ#��I�2�:J��?��d>���e�D�+�����!��Fn���5����wѲ�ao�aA�%�@�:^�L:�\�7���n����<&����=r���0x���Ə���� p�J�{
&��fQ��I�0o��/=�"u���:\DXV�[�'V���lh���r���2��w$i�����1X+��~�?�Ғe��P@ND$��y���ǲԕ�(=���X�P�&�7�x.%���IA���ք���q���PD%�nD.�D(��N�9���6�\i��x$dCzT���[Ⱥ��I8~6�#L$&⨵AY($��f��{8t��]���'�7y膼��2��1��Р�6�NJ�(w�����ށw\	�d�����E�����G���U��FP�����G�-��f�b���f���p�������>-\���3k$o:i&[��u��dL�(Cpd
Oqu2,[4���Z)q��Y	�u[�}���	����/s�*��G�Hpe������$``"e�:U�y��܆b��-tvn��Z�&����z�0L[�-ox�,�ZK7������K�ys����v- ���[K�j�;m���t_q�~��/�Ju�.�)4a�e��:�37	�@�yN�A˛��!?ܖ]����4��ܢ��j{������Wi�$��,%���\E�X���SZ��ʂ�e��y���U�攨(���6�w�9t!���~ݡ�Yq��z���H�sT{m3����P0�,��x���眻����N�<>n�o��WD�v� ���!$#�b�H���	�'���U��z�� ����a�߯�O�h��'�K�����ۄ24+EW��ۻChC�ei,I��$0�r�+	��׀��uS7�!R��77A�
�������\;j�܋�ʋ�u-��^�7��>�B o){������1؈��_n�eHGw՝��6x��GD��P��fX`yꠦ]w�_������^�1�f�a�t��jiN}%U���<f�P���2��~@}����I}� �gI��׹Ci���1������v�P�:�\�*o�ǻ	ǌ�V`C�S���<�~s��ˑ��j�I�����yS4��Hv����R3!(a��T�ڐ�n�ˌ���81�� JG�=Ts��̵���ϓ\�v�'���-c�=cS>�Y�t�?����<x�Ќ�ޒυfo ��ջ<�v����3�k3��L �Lj��8aY.�}~�=��(�a���Rh�rk��)O���*V�~�Щ�5�L.L�U1u�D2����0�9��ptr��+@��Wg�VJ��b�.X�e�VL�S�\���=Ը�BW�A����lF4sg� T$���X?	�����^��&��UC%>Y�PT9R1��vJ��&{!�����-�����9�(2��C�����bs�E^��_W�~���$~��.���M�UXWvK �j4NѸ^ ��;g"`�֐cɹ��y{���r10��[������{W��|⬳��u ��xk�{�R5��M�Qu/��bb��i<.z`@s[g��!&(h�Q:�L9��~�@���=Ev�b�j��>�\�ӵT�-��̻ �?qF��s�P`��%�����|�D��W���ז��ap��QT(�[�+-��Z.�&�5�,R)�'��#=���2�2&/��k0�=�����0^����;�{��nҌ��@Y1'���6��.���-f!��#͝c~a������%d�T>�(i���9��R2�*ʪ'�nYn�c<-�T�uX(�|�'_�s뷙����3DX���lΆǛd�`!�Ԓfc�����1��g�j'����c�QJ&��5�����@?�4��<�AX�4.!��z�wdbOA�`�1/ɧ5�L�Ttu�V�h/L�(��-e@�v���S5���҄n����׈s��6�!����*��%�a!�wT�a3b-M;��,��Eyf��2˷�x�Uw�<��GRˠ�W��l�HYEn��S��&/��nC�4��9�����9b\6Wʲ�=�Q�`���kI�AHJ&<�X��Y:�½�'
�Äv�-mC5Q۔�%	�g����`��Qd ���C�����.Ͷ���`�<,墙�้V��9M@X��f�hDJ� 3�8����0���-i#�U��@=]���]���)����lA	3{;HJuC�;ċh���C�&���6����?���k���2�+��+�6(����X���*~����	�K���Ӎ47��aR.k���O�4�TS~���F� n��trd����h@��==�|.`E�K]#�z���4�n2���**U���@�P�9"#���S̫J0a*����T�A�k�����WSc,��#���9}ĸ��@���_��!mL���K�N�.\�Oj���;H�}��G�������(�� �'MJ�o�{�6$C�a��f��uJ��݈�Ҡ$�w-� �+�� �.nM2"�Nu�o
3Ǽ����g<U=��'�s�Q�Ɍеą�,����G�ky[�y3�Q�}��%��2��G���m*v��YXy��_~S�#�RL2�v����������*TL�
Cu��`��'�Dg�RV!�^���?7
"x�/�qh_�E��f�~��g3��x�SBL)=B�Q��b蘆�0���Q"	�W��J�b�"���'��%׊@��_X�:/P� � ~(���m��E�fh2@PT�����g".8�UF����~(.)4wv���[I��J@�f����qC˶{)��{�%���-#�Ϻ�@���%ɝ=�Fp�88Y�ٙo���`=<뒐���U�=6X�:>��؞x'xPZ��JW�.h�G�<�0w�������>��
&�{2�}��r�*��7�G��!�4���zEz�"M>e�� �ʓ��3�s[R2-,�6dQ�/h�5�Z��X�Vp�1��#����\բ~y$u�f�뽚[U��1)���,����Q`������u��f��o..	��L!�$ͲmVy&l�mΟr�c��0�魫~�\�RS_��@�#�e#^�t÷1��8���jk9�װ�Ǔe���[��И�n�Jc��m-9P��^`�(KWF7g�\��r�L;�Gf� &Q����Lw�|¥H���3����hu9`I�yE�4�>ik؛yL2h����RNԲ�u����Px��bU�0��H?? ~� ���C�Xsf�Hq%��_+�!(����7�ӻ���O����U4tx�*I�_�Ϧ���T[=^\Ң�/Ի9u���הE��a�ii+���Lm��Rẁ����f�LADǿMJ�����"��]���1G��ɳ��Ʒ��'�����oQ�]d.����(������V��jS�T�&¡���h�����߆�<ܾyB�� #V���[�	������s�\��F�BB|z����o�Y{���\�+A��ş)c�xF1z���T<p&.�kH>���ɛF�8m�Hx��$��1q��2t1Y0���p�C�Gy�̕�t�QAPn ד ��� ��x莝�N�&� �Դ砌�O�����̽O�a���[M$2��t�/�zΰ|񈳾�U6��y�Om��7�2t�C��zE�^�n������)}��Ŷ�#���ϱ{/��qU���B�h��R<�dq�!p�:�"���W��YKK�r��f�o�ؘ\��eu[����f�Ð�{6j])_Fʣ��e,���U�ܴ`���a5.�������fU���/�~�H��	b����G�5�����#C�K�˨�ŗ�M�/�V�����j�`��;�\Z!ۋ�և`�A�-*}�������T�?�1R�b�� ���ֱVp�Ym�P����fB��{���q��
�ȯMU�����Z!}�U���+���u29q���-�:�Z�E_�E\�=g���]A���g$oiy�ɏ�[M?&~�ZnG�_�E��@ÊA|��iݯR�)�����na����IP&�)���g�y�a�y����G���4���8��+7�I�v u[�՚��K �ײB�E��[߰�P�0�a�*���#�>�}�|O�Ka!{�̩�സ��EP��?9���%��l+�����;�p��X$ 16W�. u�����Ɩ��(B��4R��,�V����gY�_��7�F��$�A����t��j=m�L��[��*�Wf<�SL�W��!�]`kT+%$<�5�]K�ꪷ>?M��_���|����8|�V�i�����F�k>��n�/���'U�'/�(/u�|J�#XN%5�q�<���v51�%|#���Q� ��o�d3�|��p}�GD5V���Q �'D��*׺X{�T>N���k?�䪝 �-%��~�J�AMN9���sS .h75{�Z�$��騧B]Xhx�o����a�H�y��O�%�뭍Ǣ�4��F��9i6�nG!hL���ᗴg�!S{
xg�uPh|s��K�7�|�fm�"gMPi]�RR�vB7����8,���L>ʵc�Ud�R
�c�	U�*�^�>��%�  s�0<KC��X��9w�T�Jq�����_�`�Ϝ#�4�����B�����Z'��+�uP22S�����u���B�=|�O� ���K��oٝj��s�ʮ��̓�}p��G<,$	P-*���%%~�r;�ؗM�`NG����+���#����0ei��6[� ЋoNQ��a}��*�g)��w�(64�j�����һ1����	e��G�r� ������7Hpe}�����O��G�|p9���9�l� �V��"^B�y�r��sbH2�"%�D���u�;(z{���=�GIeh�����.6I�Ò���[(��ɸ]���*������㞢�dq�$!�{`��XS�A%�����=*��_5F��U�K��SQ���r	趡`�����m]օ�Î�$.:���i7�yE8�
���@,,Y*?��ɴ�Dp������G�]Fr�=��wt�	���);V�Q�8��q���f���! dr#��@�4ά]�0�i��#��.X�V��2�E�V������M���b}�O�M+X��`Q����x4�<l��q%Їyy��eiM�4��ֳ�9��Ԅ-�o9=�h�_��A�U&��b_�&h�?�V��m���P��p q�Jnd?�\�0�/�cì��w�~�������Z1�c�V�VB����T����sֆ�<K���)��S�jj4'���mEŬ!�7@�n����P��,6��8�㒱A=��!-���j���܍:9�AZ��rҶ	���*G&������N� 8��Nk�ͧ+>�wb��j��ݓ~E��6�S�QĹ�h+(�I��a��w]�l��g�]&��>W����Y/=�
��0�{:
�h�҅�Qכ�&�/A��{*ю��	�]G��s%ë�]W�s���}�EJt�2U�7]���kX��h�J^%�����?�wm��ry[¤�^�^`ntq�iUw��ǂ�1i��ݶih3d5@��5R��7�y�..Q�2t9)Z�	�{/s&o5+qB�ۥ�7��i{��-|��ps�,˶9��y����r���!�0�@�6��>=��Wr�!�H�WԺ��\&ɳ�.�-���o���W��[���0S�JTVB�V�i`_�;�Q�a���j�ߊ[ꖊ���K-��a�������d��*�/�&8n�o$e塠�S����^G(��9�|:*V�s����"f'�Y̗3��G�9Q#O�������ە
%��_�Gl(¢k�u8v8B?�����=Ү�6�w�CcT9o������P�\q����lB���[;!�W�lE6[�~����q@���[9�84z�^�g��K�1��bfP��&���]����Î�Kzj�m�iY���U�FY;6�J�5�/�����{�i������~7"
���� �\M��c2�����n������M�S��p/C�T>2�1xh�wl��\��q��w:��ޅ��0������:�Zs��O ��_$oRg�/���F���ʐ�6T��!��lr�U��/fhl���Uw]�q<��%p5�@'��0u�G�ti����q����O�W�ԃC;�{F�}�I���FF�!V��#U7�m��n�n�T5�_m����4��q&�@>��cF�0�)���@>0���/��<a�Bcs�+(�P��5����@D�
�3���Z�K��:9q;ԙXL&�`��,F�=�
Z.~�]x�c�<�q������+<(h��D7��柌c��9��~W9�E�����u��ҦO��ʇkd���:C؈�fsΝ�|�F���̘��,/����خ�e#5?�q�K��?"bZ)g�x���_��sU�����J���	$��FĲ+i�C�oH�|��E<4�J��T��_x���zvL�Ց�M�����Aњ�t:���ʟ�T��H�(�}qc�7�5���ٍa��X����D��ʘnx�&S�Fo)K ɾl wD����x�,A��o�ftA��Rх��m�����E�z�L<����wa?`I��Y�X���ҙn�;:���z��}l�,��L�|}[pT���Ҭ�Q_U׎5:���GSQyW�c�q�Ih�� ��^BK�8l_�f3�q����U��[��귍�T����ɘq��Z���2�y���a-���dU][)U���Q�ʖ{�����x1��ϯ�1K������aN%m%�s�o��y4{hr�C*^�r���+�YN���8��p���h���a����#�]�aneyʗf��=w�x��"�n����)����Pp�D�l	j�	j�!39|؞G2����ɩ�i'�32���$���M�RB�mI)����D�z�2Ѷ#���Xk����9�+��&��W�<�F���>���U��s��߭8�FĮ�u+~LiG�?�fGV@���1��S^���~�N{�������
J����n2�	�+�H"_�H<�A{v9�*�i�Z9�̱��|�3��@��ݩlIA�I��l�����[��PN�aQO�f,m�}5�.�o�7JF��;G�yp��	 !���A5JO����(����(JS��W��S(��V�S	���]��wZZZxl�V�!F�E��c�ˠ��/"�t४T��O��pS��\l��	ї��!�_��n�G��%��?P KΖ��G��laڈ�#կQ�Z����-���L�g7ъ�������uwʈ�V��~�ʛ�aRt���P�ڞ���/̐��+�H�Z���j��z���m۠.k���ob�v�:��X��/Ig��5���|i�����J�5㪷�c���m������3~��!�ޙu�|pƥ�yɧ�PY���{�˱|�΃=�o1�$ܽ�R���	K�F��k�Ѷ�&����v�ވ� ��X��)���C��4����8�RT(��V2���C����}�)��i��'fB6���$u��WԵ��B�X��)���Jl�;:󑺯����+Ç���*�i�������J�jVo�d��$�c���.��O�D6��.$�)jƣ�2\**�_
��]	Kh��J��Yk2(�:&�ĕ��Dnz>�5�y����&6��:��Bz%Ğ��(m�+!�fA������z���Jo�f}���DM՘g]?ut�\�J��	O�Èq��x�H-��t����9Aޞ��zo����I��ޜO��M����@�v���@�����q��ڡì
���4y��v�V]�s�ː�D6����~D眿���W�sQ��.-��(�%l���]�Ŕ�yO�>���5�m֧n��.=V�v@���C�W�e���A�ظ�L���J���R���P�Ő�Z^�]�3�4w�i�{-G�R��\b�=����\k��/g�!E�r!�� in�@,�8��.����8�rTy��sH=|��z�Fi����J�1���p��Q��|��m�	�� dء�I����1��v�$Bu -�G�d�2z���ȕ2�x�un�]9nx�������!L�ix"SX_X0����s3�� }�Zk<ߠI_F���r�	c
H��h�kz΄h�ز���L�C@`N��0@"B<�w�#�b����yY6���6D��X;�
 h	��h�����udy�]&m9��)�I�D��c��:�T�>�l&,��YO��'��ӣ���(�KJAg�i8�6����rŵ� 1Iӭ�|���Hr2,�})��^�@3�j;H]qEO�u <�9�+��~�n�.OԶG��=b��-�ǝ��ſ��DZ@�rg��S�M�4�������~�_l�uƏ��&�U���W=�+�紙��X0�5�1�O ��_I��d��{�o�tOAIq]��Z��gs�l���F��gNM]NF'�tc�yZn-їt����ø4�#x9.�T�چ�v�O�D7+�}7��p8�ǟr3��8Y�@�WA�)M	B���\���\u�G���B�X�؂lO�qc��9�}}<���]^d��==\9�`��̫/%}Ɉ���}?e�1���w 4e\*�+��6�N��P�����:pg��w�q��m���Wl�õ:���Z��Ն��U��j�3|�j0�(6v�jU�:�6�|���'��W]���}Fc���ɺ}��Z���ܶ�Q�ˊ�鏂��r��~WW^�:���:�s�U�E��
���H��CSc�}��d	�1�ː��s.)[�dmd.�r6�Z�2�+�҉ �E~��d�toһ�w����B�±z��b�ʠ��F���]$=V�P <�uG�Ӵɭ������X��:7�ǆ���>�MdZ���j�'�1��ϫθ�l`����g��K%�Fļ򮿰�">Tm|XHͅQ�L���Ōrͨ�B�=LD��n;��t��w��A
�o���H�_��s�*��v2%�p��O�Ļ�����AI���ٗ�1k��E~(.�����2s��2L�\|0RP���p��RNx�<G��'��K耙��;ϳ�FBy����k..nh�o�Q)�j�X��6�Ǳm�&� ����D3��Hk_�Y��W�����t�v��2ݺ*��XI�kB��$L�l�D�1�o�`��i�����»±��z4�
���?�d;B%�P� R(�5m�������r�H�_j<��V��+j<^�ls���$��z���(1�K���(���wh�`����i�}���cZ^jHZ�ҖHF�mj!��K��L���	j�g.��g:��Ó2��,� �	&E�l�c��A�ja����/��1jo���ra����է�$]���ᡷEd3�Ea��V��+�ЈKM*i�h��7Q��az&�q�w�XWa�W����a�텦���E��%L���

���_z)�NC�7�X�K��  1�#8��L�ǖl�������ž�H�o������)�0a�y�T��`��]ۘ*��
�#����}Y��[�Q=��w�Q6�f��>I)C�1�nFA�o�޼���ׂ/��q	�Xo.�'�vx),-e x�S��X�t���d&&���j�|w!jIn�mq�ߍ�#Em��~:�0 *�s����Bo*n�?��:=����Ә�:c�X���-�)?9��#�U/���?�ܳ�@�H>E�5��R+�����rਥ�n ����cU{v�� }\��%��C@�GV3���'�7%w�.M�{~�\5I
08�V�L�Q.�Hm����">�_)��y����� �+�������9��R�R��y��k�7�iO��)�����V��`Iu�8�1k
��n��3�5Z����%3U5 ��"Ns1z�t�N�ƶ[�D�ds�}�tJgpf�o��ĺ�/2a"�6�~.�����?>n��f�O�y�E�4~��R*u2���sy�3��m�����j�ΆP(r�x884G�!hHC@,�Cs��3q.���_��C�R���(�?8��ݛ3�Y��
�fـ���kb&
��l�b��Ydb�O�=��>[��Y���L�k6��uZ�X������'pqQc�6�plS��Υ��wGЇ��9v�}�������j܁U�;�����d$���a�����uZ�,�Qc ���g���vbQ���S֑��KL��l��A&u"��շD����)B�ΰU�j���&� ��]���K�iְ�l�U����<���lr�[#�	Bz�%^��?-���q	3?��ZB5Z~p��S�g��e�gS�#��?ۨ,q��X�4��(o�%��K�t�j5�&b�\��W��S����¬ZZ�P�U��<[���Rh��f��P}���<��0��ޢ�� �� ���TFCf�i� �:��+���H��)4YI��W^{��q5�j�Z7�?��D��qmXr� [#%�	Z��N����@@/̳�oG̥C��gR���p*֙��F�8p=n,金
�\�����j��z�[����:総o���iu��j}U���~�J��}��������7�K*12�vkRw����]+�9��?=y�^��A ��R�{R��6r	����{�J���~���ؚ�ѿ�ؠfm��T�5m�1�3+���A�%x�>�s�(�J�F�Qp~T|UgD� #aa��S�I�HQv5Ǖ ��y'��J쩗a�m
����/q�\�Xk1��@[�H�-�#�4@�$[����ݤ��5V�{��RWG��M3�c�H�����ת� Zs��<�7I!q]��a�qc�� � ��v���F�~����T�} �ۖ�dpj�ޡ�בe��@߷%A{�]�-v��L�X�nvF5'�~�}����p�9�ş�(%r��c�;�����l}ӱ���|���G�7��A;�:�EJq�q�S�2�e$i�f�'O�o��M�=}}Bm�����0A��bsa��%�j�,������Y���bЄ'�����X�ح�VD{7s�gRG��,���a
��_~o ud_��.����-8����A�l0i�"�{t*���������*�ᐇ�L�V�c��|Ml��JGU�.���hF��Jǐ��uc�9�p����0ȹ�>o�
��^���-�����
%\,�V�43#�W���Q��!Ck��Hi��)RH
��
MpH,�~1���U4|��?	�^��?�\2aMlH�������T(�(�c>��p�Μr�r�YE���\����+L����Yj)3���\���������;;��%��J���8�&�@+��*�k�c-|���g�|}"cff��
�~��Kz;�W�>��@�@�%6u3�|�I�'	v0�S�i0��k��c�lߊt@Y>�~����1��Ǣ�bgF��;�j�� 
�&�-��p2�3f��i�A� 	�D�c�o�:p#�b��[x(������S �1=p��1'6��0U3��`R�7|�\._�O �cȁ`��Q���5|�\�WJ�h�l("��Poqu.X�s�����',Va�ɁI�<g_SyF�r��7��4�q����3���;!�f����'8L��T�į���(�cȄ�m�J�(����;�9�=2�a���c�kp#UjkY^R͇�����*���l5�x_���=�K�v̜�I�6s��)Ka-�qg`�3�5���Ff���O�[�-�Ds�Eه�:��q`~�e�����pYd��'�4vf���!Wx$UL�u�S&������D�#R"�ڲ����;��>+�Zn˛�Γ
�F��FW뮨�V��b�Bk�^��19w���)�0�]��1�7�u��N��VA�kw���M1�>N���ʓ��Ǹ����}�8��?$FJ.4YM`Q!ա�_E�����s=ٯoZ�b}� ��h	�N�%0�$�|��P_��y��V4�����S���e�
2`J�Ҷ�K�������'[=�8~�_";�����Z]ޔ����d��Je$�}�7��q�pTQ�(�|�bBoL�0b��qv?(��@Z �y�բ���$D��%z�؋�����R�x�Ԝog�u����,ǔ,�e{t5�>�B�لJ�V�B�NM���83��V��#��p	������(���&�rT��F��h�ٛڙ��q�_����8X{)��b���k��(�LF�����S5���kٗLs�t�&D�҅�Qz�`�b�pj���IFS
=m���Ov� ��H�tC��`'���k~��o��?e*�Ԏ��8�A������zԂ�ҳ�_�Ɋ��"�};7�@;��� ��0����=���{��+(��O.�X����W3��Q^W��t�`K#18M/þq�S�� )�
i�.�<G+�����ӝXnA��xAj$���و2b�	��gP�Y���t����~p??n�"�vn]P.Wp��,9��T�;[Sگ{~�f��<҈��A>=ֱR�4q��zz`��CAQ�@��;�K��晶U?�<�����Zþ��>��i����(���GA�	/�΢!1DI�Ƣ�%V�8�윕C:�6�r�e����k+�*\ʹ�d�Gh{}\0҃�x���H����0�sj��$�y}�������I�O//������\(٫������D�i�ZȐw��:j�����e�f��Y~ү
�Lj���Ԟs�x�u�� ]`�7Mq�3aΫN��O�ui�bC�.��}�n�@0ps=l����*6+�:NUp�/��~�{�o4�����0жlW�2
ͩe%4�T���F��_"��Y��I�ȣc�
�F��
!��[
"LA��ti��KQ"ua��?m����bf(��Q�/,��X��A�L��"ƺ0Z�,+��h�0C�z�dY�XR�c��~>��q	�;F�gfL�6��5�����}�_��ׂZ�HSs#����ށk�E�������p�O�S�*͝?[~����8)���Ŕ��Sy��wsْ������,jG�cMs+��x���me=�9����{�B"�VN�D���P���Pֹ��u����z�j�YXc_��oi>�L��a�]���_�:���؈��˦�?���SC�T��J��RQP�|
YK�@͕r�<�3
��>���7rx�ܮ��u C�0��P@��I���#��iV%�a-��@�`�,b�wkrR��j&ƫ��e(ȋ��܌��B��{:�gԫ�4�I���D��ݎU��Z��\YeH�Ȩd43�O*�t�atÕ�a{�/�@aR��Q���AQ�5��1�Jt�5BƨQ��_o>��u>�]Ԁ�@��$E6
��->�y�ݝ:�܏֔��7����.�]�_R���m����dO�����',Ε~���a����d����Хtpw,��}���>���)�2qɊ�][/�����ﱩ�]�7������F]��arri��]_�w�����f(a�kM:���b�Wʽ���J����xor�A'HB���P�|5)�]lyX�(ݨ�?.T�e?6��|�uEF!	8���2�OSiZ�������^�Y��	v���!����|���Ț���f���W�6�YM���\X���I>}L>���2y�|.{�����S�Z�&/���;m21��B��zi.=��r��	h�����f�KC�����zf`�M�/E��1��ǀ� 
*��>@͏�j&qu����S���(�t����Ȇ�m'p����4d:v%T;wc$�,HU���Р�	���~��ɣ9�+K�'`�&��M�l�]�x|�Wz��'��>���)�����3l�k��b�j��@�Gx>I����#Y�+@����"�>D��cOj=ns����l�6`���ISU�<����϶�MkPi|������  �!V����$fF�r�0v����(hbvoa��i�tg&C���������4���i���p��;,�.ff~���ܠ����-�ن�,��[����Wen���}f�[ro�md1�IT*
+�b���Hn��(�:2u�N$�Μ���L��x�Fln�np<)�	�	�6柠�Н�}*fRŵ]:�M���4�&A��
ω	��A�zt�=?f�����g�In��;�	�}@��~������!�]T�kP�+������8[�P��
���+�.^Mp"�A��\<+r�<��]�.�u�pH �_�a���.<�E~9����[]&�J'=@׋߼��f�ĥ�r��鿕�,��E�A�_��׎��>7��s�ަ_�$LO�e�B��vA�Џ�� �qٔ+N�͉C�	'�+VYX�W�~�ٹ#�'S� k��p���r���cY�F�]Rr��a3n´q=�ΒM�o�>,��L��k�*��e������xx6�z8�k'��n�3���)�9�!���1��4!b���$/�fj��+�U��t!�O@$/����	���ׇj�D�@�n%B0o�Io|�Bz��d����WF���S�_�p����I9r⭤�*PKA�\DR��#�/�1�w��7OgtÒ�f��}6'Q���D���b�+e��Pv_e�T��G��Q6m��v%����8�喼~�l\�T��kX��#����~�����n>$ y���������-����G�������j��X��9�V�H|�4�w/T�p��9�cS%(�|D�����t1�co������1|³�CS�1(���ۯI���sf�5��v,G�M������9unQ[�[���HF�·��c}o�"�F�%]Nh^�#�d��)����٢>
�R����0���hM2�ٞ�����B�����4{Gـ����x���֥��?i"|X}�d��B C��m��h��j@�CC�ˤ«�Ek�z�������2�h�%�E�_F�5Z�u�˔ZFn8�=�9������	��zv�aE��������t��9�xռ�`U}�sN:B6,�mӈ�ݠ�3߳��.��Y1n�
��~��5� t+9jI�VC�W;]әSv1����e)Mgg�5c�i�E&�BB������QE���FwGg#gV?p@�^��2]�L R��l�<�u�!���ԨA@���y3�/ղ��Z�7�>:wO�olm�����a������Q�:z�o�4U;��?�����dp��M4�;YZ�)���|ȯ�/�g�ۆ��2�xT�gL���p���$\K��Ӷ쇠`;M7w1$=��/W�S�tw��lI�!Y�Ok��_*E]k���B}a-ȅ����`�2���IA�.^(˹�|���H4�YېL���EF�J�nG�H���Ȩ	_��¢q��@"�=8�}���e�Y��~v�7�[�7��O `�:���g6  y�h;<�dv���f�z!"��������k����aU����iiLJ��)�A��ǈ1���І6�P{Ǡx�ux�5�'n���=�1s�l��z�i@*��r^���7���/��lΝ�Gb%-��`�'ȿsG�M�e*�Ok�l����=����c�`��vK�yhj:��uo�����U��<%륗m~�O���R;�4�Ǭ���$�L���{ra�5�*w��f��Bٶ�U�+�q�\MH9���8����y`�KЩ���!��dច:+CNO̪R����"���dJC�8ٱ�H|z��_X ��;��}�yPπkV���F��@� o�ɯ཈���F~;8�
�w�=�)	�|�V��t.%��qY�Zm�`1����|���Վ2q!I)��0<6{^��Qh�L��Q�Iʼe��f`ٝ����;t9-��2�	��Ҁ��?K^�fɵG����6x]X���=r��	h�ZM�Q^�9^N��0q�A�E�ǰ�V�1Uo㉀/�f|�RG9��}�#j��
���y��h�*#g�sm��E�&�{�F����ʿl����J���"�>�ȧ̶zC�I
q�@/!��[u�K��%�L�?R�����u)�����ՉƿVInJ����
�&f!,Y.��`�BB����.��!8D���"<ia�xʀ�>w5���ٜ��ѓ!��'[�@��|�X�����`t���@���rc��O��0�DWݣ?܋��U��h��Ĺy&�
{�M��Gz��h����}���Q��%��	"��S=<��� ��֪��w�u���V�RRhN�+3�[iQ��xD�`D�#�;�Ժx,.U7�a|�T��V̤�O2Ʉ��i�)o[_�];�3 ��$�j���mT�6��4��p�7pX��(Ѩ=�@D#(� ��P���є,��e\�jB��C;f�CK�5����6����� #�����9�"\m�,����r,��ro{z�+P�sC����5Y�ϱ����Z�Q�1(g>��5긦>&v�<Ŧ@��:��~��ߣH���F�����r��r7�E���v¬�E)+!���h�"5���Oa)MJ�˧�x���2���I�ZL6x\G���9*0�%�æ��D�-ק���4A�}Q�;���ed"<��z!�A?��.0�fA6�\���j�:c���ݫ��"�ɏ�uK���'���| RM�1��hg�M�a���{į5�b��B�m��#� �p����2y��|�D��'n��R�d����ɤ�x��#�	��K�{o�!E��6�1�Qe	��bP��K(L����@.��l	�E�SC��(״�|f�>��pM��V�KXD�靊����#�7�̘̫������N�/�s�(�FU��F�)��D��P]����� m��r�G�1��cc�����䦂,�-���K�����EyFU��V�c�MQL��I�T�b0�}z5��-���,B*FAs�	����f$3���<���.#�zH�D:M(Z���e�<�̕�E3c�h�O�����R��,4��8����3w�xY��G�u���o�
��c�[fy�Z���q�>�"����W#�o|Gs��M�" wh@
Ha<*@���WG�E�z�ͮi�z�$�mV�|Y)5�l(-�(���\�yYdf�yk^�ܽ�W��m�\H�_��߀I�O2�s��~Xg�|�Hh���r����	><K��K7�<������q/z��C��m`@	�H�^+�Y��O�,"�i�k�ë�9��&	΁��rl|'/�E���c���=���,������c�L
�c��CQ&��3���*��G���ߑ�t���\G`׉2�t�fKдo���$���?�H�#��(vU?-���}���f���t�)
�	R���֚)�H�Л��u�0�0NH��}�̑���~�&�(�cXEJ�u��
�͖�eϣ����J�Y��l��2���LK��9�\�c�E���+!6 L��%�t�lXku�;�+Eq�,��ǼWPz�8慠ˉ>��)lg����O��Y�����Λ3��WRìh��TƮ�i%��2����iX*�WKi�0ˁ�5�>ɉ��}�(bi�ɢ��5�gUkdL5�������Fܯ���ϕ����Җ�Ƭ�{�Ź' ��L��@ݴ^��.���ҭ>�T(�Y#����=��sw*a�/R�`���g�.�*�~�[r��n4a[��\$LW�_��LP���TqD�����k�x�$���`��?�������yA�\�Y;��*�s�Ǿ��g<n��4ظ4�˭�KzA�;�kR#%�/�-�0ɓ��TF���"��т�����7"Ѭ���lUk����ʄmSǉ+J���[�з�~k��+͏}>�ע;K*~����ߐO�L6Fm/z��=�+���~�X�-^~��Iȋ���?y����ކ�Ô�0+,�wߏ�y��xg;C��H�k�B���m컐]�*v�'��d�#�Ν��{_z�W'��Z,������l����ɬq�g�P�Q��u0G,o�z�u���{�O`A�1"�C�n�W[Xi/;���#j�.��K�>~ά��u�q�2���h=�e��Ȍ��U�ڐ�ΥX�DH�8���m@6[�1���姽��<��Y-�Th�<�R��uZM%)*]�K��C����ND�8<�#m�pr��ފ�d@�C:Y��݈tj��f�\�tb�=ϟ��)���E^�(cQϜ��}X�j������L������7������{�2sk��ˇCΚ[����~.��T��2�'0t�`�%[�u�a�=����Ė���p ����ch�E����Ϻcfq�� ��ʰ�yfҊ�\��8��V[4.祶���+�U򿌰%��+��@)U�7P��/`	�t-��װ��0c`�u6a{��C���L�v����S��]5��61�{�~c��.fِ�`����-9G'����{��ڊ!����ļg�Cn@M��`�H�q����/��ӓjl�<��>����#h���J�Y*��~J��;(�uh^vK�&�|ar���3+u �'ߨB�����f��w��l�}�V7��.P�Yh�/#��?�u�Ɛ }���IyKY���/Fsֈst��ݷ��'M0�+�ѓ� C-�#�͹�p6����h�t�&����\b�Z�K�28y	�Y�I�c{�q�Vmw�!R��|�R��2->��w;�Z�R�'��>	���KWDA���%�o��:^lM�_CNml3���­��X�� ���f��o4�9�ZC����K�Zk��^;��ֿ硒�O�W��5}�ܗS��}�ᣊWi�P+� /����|�%���iZ�Za2%a`d�pUg5�������ci��[bʠ��Z�u���c"��W�
H�*#lj���Mg��y0�!Շ�j�8Ҟ�^�a���[`t-�U�9������3{���Z8�9l��+k��߯���]q�3ԍ�ޱ�)�z�c���\�ʠ��_z����rad%R��ݢ�j>5�6���[���A�)���gB��Yp��� ʋ�ΡPi���Jœ��dv��TN,�����7�ô��f���n�=Zx.u��ǒ�Ni��rN)`,�-ZĒ�0sLc�it�I_����5�sDD�?�5����̾U�H.G l���@,|�y��)V=�)�p����s����("U�����J���6�&Zk�̺��\yP����^ȸ�����媣�x����[�<ԍ]����yj�����Z6�u�\��jf�[��ӑ9�Y�KQ�`p�T{�'11{/�F�\PX
��'�J�����@rݻ�.]G~��	O���p�H�JrSh�+	I��W��-*� ��K !;�w�M���1F
	:�R{z�C�Z�;a(:j�D�d�9�����ol�D�Z�����4����x�A�����^�ۥ���\�B�p�4	���n'S�a��:�ނ�œ�����]���������ҸsQ5`V3p�#