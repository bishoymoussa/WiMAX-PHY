-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
ksPrHsBmy2T4jpSLdIY09EGqmhv0luMVREQ66jhN8elLesq7VSxZzbFiur3e81KA9dslPSfk2BfF
UaSw0fZpBjBfuWPZDPbf/hBv7yv26Ui0pbOExEf6kzTEWpVd4LsRHZWmVVzkd5lbBY8VfKZopPFQ
DU/ejJdYrqZ+Bp4IWiTIhJvo0PnS6D8OpqWDEmEXc8/y72agHJb7n7qJBLF0IMACjxigFnC9kEfl
5ItmrC5W2aCN4qtWqO2mDsRJbmP/r3p974yLeOEtuUAPU3LxsCk9P8N/AsWhhj/luq9FPDh2BP63
l5oLLzF3Fj7xtdn4+ST9REd/mLlZYlFg2LczUw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 40224)
`protect data_block
enncrfKFTg58zj3nhNNnprmubdbv8YHLb1ADNplo3ZrRDBGZ9H8cw+QEFXpP9f0GxuqbhEIWLuL6
XTd0eA5RDocAzC0JumDkl71wYaulRHMt0141seRsmnIT1WFomzKsAWxgI/GczUin7ajcHPpL5ouQ
H3hRn94Y6VW0uNhb8RlZVQmyDVoDozeRKDpBmRfIMe1/+/hAzGKYmNZ8u7wCqSUxeTRUJQ9oEmY7
iNpDsbxetcpMqG9g77fzTLPzyvAEG/BeAWUUoVPovMZ1JaL3kRDTbg+7zNsHLDVchQC7uui0BcUg
zp/ONG4bVggWliq91fEYfVmi3/+mvyBifVBzz4qFOQsQOFC08PPnRasisDd2crOoEe0Lr7Qfd2Ug
ssFuGbsDkx4K7bo6ZKaW7S8kvrb1jgOeqgOE2xu/YhXk9Uivv0Oci7IbusI0p1SHRABHgO/Mljvc
QcSrcjdGMXOpxtTTISrFRD1Q8oeqfMIbwtRXjHgtMoKXuLqzywqTIvlhD2cmkuy1crX75fJEFNFu
RT3DrOLohjn5u1sZ8aE/ScB1dQ20gcnSQEttjwzh7FSsNb4pFkmSv/1EJE4qOFtPzND5AkFsDumQ
vkNicae4Sl99ggJStSY8icg73da9J4OqsUknFGzo1uw35JmYO8NCajbNNIAZlRBvKQOF3sfP4OI9
qWWwdaBrGauw1RCVoU/DcfiXjbwWMYEi3M8TsF80cAZh4IwVEjJKcvltULEz5F7j2mf5YtW7QjdS
3T7hfS+7ZdZeFO391nn0ws6gEKyw80z0jkIDID/Bj+j5Q3xj8FYLA2lOmFkrTGMPQrvXZHQ+3QtJ
I3lQaG8T+EgjjH/9ouf/wyzZjAEHmfEc/28/pqV5wS98193e6Kx2/svwkCxVcCQVaVqGubBtIbQ5
YmXkLQhB0QRXiclpGC49tdcaUP8xJfUScfzvyO6pyP2qIG2hhdCKgaNmxpiAfZqJtrJR0j7+VQV3
MhHd5i9iMkdTsNCdD9NbsJ9rF4QTT8dS3DxODKL4WntGDQAhVEz4dDAK/dPhqOLruCQjLUAh0311
n1rM4UVsH+3ZMygTa5V7LkjVQvL9zZuOM5A93TXIWGr5ZqcnlROvs2+MF1ze7TQXYtgb0741GEwR
p8sUfumlkIl7ma+FRn9+ZP0oXdaD8YcxZ/oOQbPsVVVgfTMtW1Ory2egZkAv2g2hI2je7YbBEBZH
saEDG9lqeifGTedodO71ARBp7HByvr8EzOsdicX+EkcEj3oFh4pdEu641LdHyZwqRvcuyz7zduOl
DkZlRVtpTZhBrvfb773SiuRVNCahNUCXOxefpgT+O+r4Ae81LjqkN97pVmC8SR1At9d9e0LJvC9w
CyBIc0/CREbf2+8cOaXBTStHnE6VAfR4MPeQqOz1wqydKFzBO0guCNufFHGTh4TuYpJ8w6KkwjTz
NMPxnIhSirrSUNpcmVeAdde37O03QnPaSZWXmmAcjmwFGUgckK4QKzlPc9kyd2gDvfP6NNRmA/rI
opJGV9R2B1MLZd5N2D2qKNty0PmmEjnGQt4tXB8bHA2eP63pQhY+HI/vbJGX8aqxW/PscA5I+pRJ
PwTTSoKGsqg7cz8WiYhu1sbCyAYO0eIvwsdp0Piat7mWI/kyjmT3CVXMsOxMJxk1CYeABoLpqWSl
77bipLG2rl2o+qxZwbjBD6arPgm+jCdmxRoU+Yxw3eWJiaedySUBkndUCADTalAi5vHYjYEbfWdH
dpK4fa3t0GSQDaYGu/Q9H26rn2S+UbNXYmHqV9Mv7gL/U+TjFrBXCnVvEmxcSgyWL5RraYFB0jwN
P3E0rZo0iM+9E9K96h5IAzX3rc36FlDd2rZRktm4aozSCx8DISeHkU6xweTBYzjqN8763FVbu69j
zYK6sl/LTL2Q2wYUkFLmmWZPdn8ZsNYYYAstQ5ufQok1yEzCOWVztjLNh7s1E2jXNzv+IGCrpbAr
D/GQmP3I6wVxYujBq499i+5EHuPDBNQ5p2cRNiyt5VZEWjTMq9Rle7vda7WPaw5s49QLr48NaH4n
XY/+FcnD4qd1ZBBdc8P2hBVxCg9wz03PjZ3hUpH5wYG9MYbZO3BcBWBzY7TAXjWD7kUqRO043FxD
3gfdyNEZUNAUF81l/3mBLe4W2vuotEDgXwXskWj4qnuW3XCufhT21EVDbNcHccauSmiNwYWXCG/c
Nv5zUV8QX45BWAvAzujT+yj/z03DfbxdODnk4YZclKulJMttxlh9YANYx7L9awEuRETyEplFqAW8
tgp0vpzoAvmDU9XzwfvBmSp7bagGWPmuXCCS8Om27iY6U8J48uBOGee/InazTAV6pRakk42wkC9C
mGWcHawljj37260Y+m4Ls4uh54fen7ZfannGJOQrmit6ZxuUphty9ltK8b2YBA37Na3bO6WYiSxw
WUEK7vZmAmYs5pnHW4y/C5Img37SCHDxPVtAq9tBYd5CGTIBwaZERwmWycBv/5g7UhhGhLcCcx31
WMoVg8eZVjtU+zjwMiNQ92NG74WOT9PqpWvoC7iV0Y9ipvHBMAmNXmKy6ES8DQkEif3AggQqfdja
JHHykEZLRLP6qr5GOzKPcNaPNvz/qYnm1c77UxHLLXE/J0SnbbWxBCR0P/BFzs8jMAt5cwTN5rpL
E3s3p+soRqIapKx/0Bv9KWZXK8HQQhzlQtI1dlB7g8JAOFbg5O0wr4+8QxmuXXIIkWgxXXvJvatb
0bot0D0I0vaMuTAM6c7XugtYE/f4xZaWKiUlbFJpe3A3fnFPiWVBKoIaVazneMi71pDUXf5QMkRo
2Gd9ZepOiOAgpr8pWfKVFOoDYbgBdpMbNUZuFl/JNd49/E9kvUxaQ9ixQr/TFTE17evRbTN+Jnk9
GXBSMiu08IqOOCD9vruuvyicp5Q5VF+scaloffnzA4YsBnEZaQTADQ4+u7oAxgQEmZ/xugoEYsvN
r+Y93/gRx3Xdea75PMlhY88+BrIf7/u3vRys7VnPasxrakyJaRVX4PnpstvB3zcZCuoIDnvhitos
dbiWtblOS2oLXEPma+vJIk0BqiWFeEYflTG2eVMW3adMg9COusP3b3kOs4rE1rZPPn1vS6XOPfaq
jRMh9w3JqxdDceFFiELXdi1BVCYBEamkE6N4qDN0nqB79xcdtWumQ2faXYaonKp7NKyEUvzAXOnw
T9dc+pYQsfha+VoEmRa46UdoGTC6x99Tlh1y96aA9EJyzgGCOOZyPC/yjqdOmiW68DBMHJHof6B1
CJucw+JWB6z2lVEtiIuiTXHfT8d2GLfqWzNJCh8CNNQOUcFhnRbB6pN70LAkjlQCpqBx8T7znP1R
RZbjfMC5tOeOg+k4uWvOUTlgNg/HxW5OFuQ0/L6W9Q11xcJK98iCZsDDmO5Au9eOryf3Kiec2bsD
5x1To4vZ8T/49mNEJ/Mxa6U+48TYc4a+I01fu9w1yVYhi2q+IIIv4I7ZQU3z+BGqCQWA0nwADdPt
hJ5M5ZG0oGQEmCte7AQ3TSIMohMtFkZ5MkPVw79unEv6ZwfjKs+pIM1o6NPfXqKWelF7EoORjx0q
G+5PJDaFiHEDxnYy6ZYuRw9FxAZpqtp7qeJrJCsTOl9ZO+J0vKGLZ8hSlRECG7J63TWuDn6dIjzu
PX4hE8/SaTdcGLr7TL74AANYr4bjVyeOj+W9ZFwXLW/BRPwBMypMXajqdE4yTeBRbH57SOaDQTA1
mu/lIOBkX4RTmw+4qhLSG0WhZpo9uxzfm0sIOS9gRmMF0biW4CjM3Xwzm+gwBzZqW8Iobx6njdWv
fzdUh8NcgeRKz1hDBWg/6qSD4v/vjoZjGFeowYtnEjAm+jcxr5qDze1cSlr63VsPSkeJtI/id9u+
+3c4vnkypAG+jHEORpErUndzy521LWTdbXUHtfpENbK1664EP0AdDwKrcUvQksRqS6Dw/1QX6/fD
VPVhnwGetRg0CeAmzmXTFEhio5OecYIa7oiebH7uPHXLyku7zUIhtq5X0+pL7Ob5RXtoe0uD+sHI
NwJsPwITIm5rMn1kR56wqspJSu8WhtsZo+vTnvbx4tuXbnu0SjB09UfrvSh8ZASroWYWRMk6GWIS
u9ZUxjI3UfX9YM4Dr6+ruO2mLeFhsxuEW3OFYW6Ev5aoVcT64Qty3T4O0Ep+jQITQqqAa8/lofmw
ST2LxCdcWtXMr+QyaU/MtY3qL+Lw3IPcGI9jvSJ38l42lL7gBHG9tXjJ4AwFhjXM/cYmuPv3Zo9X
tR50f3D3FYQOfFwzZPA6jx0H8sNfz+MYlT1f/pndjZB2AB4CZ3JoCScyTc+00tM6vqNlTgCh6Yo2
A+SyzQcJfkG1XQx90/Mf6s7uxhqH9I9LlQMZBpLLsGP89lzJZaGSgFAMPV+yrMWK2kpYoqukIfe3
QkI4gZLq2hrEJrkAzf4jtUjR9ca0QnYPIfOLRaX5KsP9sQF6+aLaciE2z+jjmdxVHsz9OMr8QhvK
jUQuoi8lmVG1h0A+ZJ0Vl1ZryDIBSlUSdpgKMgB99coiPhXS2/PeLcxmWHvhsKNLXmzImjHmjV/g
Y9byuSxfIOF9J6HN+PQp/5eFSxUncILtvUxitCU9FAbYaQT7s3uJk43cYZrDB1TqhBUzwUZIivwD
ALSLKE//vSie11UHEjr4bBIxEija0CHx9csNwvgRQygEwof4iqFWlH3yZwpkzkLxdIfHW1AJDQd9
HP+pP46As372KOWWbPHg9GCZPbBJqm0iYwFjY5tiE1IjbPl7IPClzPiM2leXp/STRIte13jL27ql
A7s0fvIpoONEuY8gTlxiildR+CbnfYAVXosSO26Mpvh5pkzEg4AyJmKBBgzPZ9cAVxYXMesjW36Q
vsCgdGlvWaI3epYeq62fq00m2qUj6TA6WvgZDnXav8622mlsNMxIEN7o6crPJQ9bwhzvuucE5coz
sHwJ/BpjVVP5AKUQeOdfbqIjsDftB1jvHfB34oh2saHqXeUc+EewumxtsFNh1GyUrMakdyjZkBJp
wgvreYkuTvzYGdBok/4EN6dbhCieC8wbxDgWthHWn4Qmf3xSLUJLKXi+H5GbinKOM/GyIUr0u8cX
jj04ilX/nmjv9K5rjCDGCYs2v/a5uKmmoqbXMvSO0Obq0cuuPPJGSF7T43P2PArYXtXQOudGzqt/
DcFgd+KCJq9+qbsIpWoZaCO3YNbrQRf/riqWtyHdMG7VQku2cCn6gy4MT548awxi3S/6NE3a1aol
9hO09PhW+XUd5WoVzb1lXXn+Gf62BS/BNht2yED7TlydYz2//Ux48AR9BFDWIDrHeA/oVA+Rp91d
NmkyzhJql/aEDufMznyMQDWB/WWGQj/pF2TtLmjefd7Xj8TDPO+lWGhht4jcW5fr4rlUxPlApxAw
pvS81ujAH38ppX6amBcDapALBU0wVyDd/9gStdQ87SkrPXL2SZs4v0Msq2EfBe4luQWCQFKHiC/u
g81RnudpSfG245LbJnV/htInKe9Gsjkc1tsSu3p7teYs0ukefobEtGdixe97o8yLEy3H/UEtv8dI
5K4RTOhZzs/2BwXmF99zQ5snIU3PydOb4Xp7yAMbg29yPJT38Ig4qs1NJ7Vu5k6b/UGntTl/jm/T
6XCHPUGoB47BFiHdjeEP4VqSQVRBnE3ZgTEoECdQrgw/xiZ0R/PDktiXkPFmRrD259h/nBmew2SL
IYF14UlqEj47ORyuUw47hMr2UTew9n53iqG3IREvgPQ2sg+JwcLbzz8COZnJyzd6kyTtIM4HE2Oy
W33h6y8+bGXR4ANF8GzXL1DQTbXdni3efWIqPSk+aV8ONR/IvRMAlIDDiUu9nD7xPKuswz0slZP2
4Hkoq0HCrBKLSRPp1TKZFjrOCEKKdS1ikB4/zq57PFFaBQN6G6eWQYSCgQDbFGFPLMBE3UPclqUM
27p+96q3fvJ7lNMlZQZQ65J+owJfpn4D/nijKWUrrweR6kMvVJBkLPhmoAGaS7tmcTbS4/VNd9p8
+4WP6/DbPti6tZvul3NYa9v2MgJ9QSMMXrX0gVp3NQC4lmfZVL6q1BC8JAg16LpcVLB1X4a0CHrx
0UVbxtJSWw3qRheJBeXgiJPpLlo+KuBXmnZODhsPlSy0K3jXj1tQB83WGS6BAUVBcNh6Nf3okRYE
QZUhpiNITL/KhMLdtJvKI6C2+xBes/HtVgnF1i+lX+75ohBEuYE95VvhyMX8fsBttfrdCw99Zosc
umJBT3MTZ/7mwfeX6n28Dcnd3oonOjW/Rf+5aamVKx83Xja/mMcZgcpr1CuTj9DMEbr3MPEMtcgt
QqDQnel0vs5/Y11tWr8uesC2M/ZZubyVFiuJaXvVihEXvls9Sq7/lw9K8MAJ18/Os8k0Ior8jdTN
8C63j5k0bekKs5kIpgF1/Kmvt46I1gPAT9WogYebYqYFVc88rF4HFLna0lBL3qEi07sizFaC570k
9iy41vG/yor1Pnm7r0GUj0jjsP73mrW2cqXR70RglX+1/CDsIoSxUkkjf6cNoha13xIvOxhqRwQw
fZ+oF6nhxgxDHMuMWCHwb/oPPizVVvOKk638/oGH5efYS4VvMY89pZV1EYVUi6YdAn9+NU22ZQh2
puyHfEcI74/ysNVX+whW40xVqmdZh/FO6oHtx85uCvGvuNex4JWKqywKeeI904s165/vKNX/wdDZ
njTnHkLiECiuDozDgD0m1rKQA3+jR/JzroFFRujWzH9xpQOJBJD732ltgCDinjzNRhcFQzJRJvqY
57cZjlrhChCVTv5wvIK1Ambzp8hbVPvYHZ6jFMkOHErM+SCmlz/GdBeYO0rfiYOqI9wx1EB4joUX
6fmFz/EdLixRi8BSDlsJMHkOOsNlKFw/VaPMlLdkhfIiOnprndoCDsUlOF8yOp1EQSDdXKATqLI8
5bRO6kbTukczPayyXWwnfjLrQBQ70s018mXrQ7i9tC0pPCcuv210/9Qrrdn0Pdz0OxlvsW6D2pJS
O/nQH86UdEQt2+7NBJR0jO4dsgRrFjHAchKifWja1zKmAGtbyRYHW04c+mQmmtBfYP0EIawLi2qs
imLCkM7LIENgu/stavoKxVikPI2q/iKOGg5j7wC1yWB4wPFG+jpF63UrbEf90Q/O1d0waky3bEll
IhOoHWbUioRmaIsoUfscxuAYonQg9+o1aR5xaWZq0D5jJWTs1gTNrZDq7qeb8AYVOV6neZE2noZf
94Rrzj5Aq5MPdrLCdDmClr0HUptw8LQaRVvBefgBv2sU5LOBrul3z+0oX0SrX9qPgReBXa0mlwU8
3qJhJxp76xMnTqcvMD1PSUAOUzx3jsJxb9dVxhi1frY4ZHIBb1IJ5DCW3F0aMZiUZq8Xj/01i3X+
VJw3v0g082qmDpx3Y8+gd0RQC15R0jHUkK9jwlkRTaxN+ou1pFjHL9BHK8roFRKe02xGLueWgIA2
JTg1bjzt89Mxz/5vYvRUJzw+UpdmVEplN/Vpa9Ahmi3KN60nzWe4HWSnh9BA+Ae8ESLU9caZOQaQ
0tKnRaiTRaV8T4Lh8tN5OtJOSRSFVF5yN31TsVughQ/wpAVL3vxGmg7nXJsbn2aHevZhtK9JnNc3
KDq42aMRI8e6WUo9w78FHHhctYsSnAsRoWb5ADKL5PxdAOv57osUUmX49XnqYb7/4bXvXyk84+2q
6LHF21v9b2kqoNbUG8Pp18Fu3rwjyKSnCpkb6AeI0mq67WZdA5cy9lu9sAeOF3o6xXL1ZkPvjUd2
Ktw1eYJkfnXEOoLjakniRLtCkICBm7INtSooM0B9lhoIrcAHBXjbHX09vYynZN5SV2cwx4ba1vKh
z65Y0CmvvnyETbnhh0gGbGfJnzJEH4iPg5zsBnoIEVChz/9vUzuMgHy6yWkrODOkwcoQdw+n6iBr
Uco4wVtpjmjv7NGZeJvCgKzzIgloxRTPeNVIcckA7XNfqJdhhYJOy+Fh2yLuITkKqp9rJFwX4hAZ
995e86T7jETUfRQ2Y6oPJaCg2az31y0Eh3OLCcYfhiJ56njPsmiELK48hT/EwXIh4B8R/T9AQtYN
H5lL4nFQBZZFzZHcrUoSioPMwkplSM4wGJ+Q9LLpn9atGTYLQkyQrIKSWCk1UEFU2uIAOtslr2sG
cgNDmHOjgV67ab7vdI+dDT+khsE0+0pPFn2IPNa+qqj5QaV0osqqd7pcWFb13spd4v3zqy5osK9x
ZD7KElEBdO7GWvlTjTvuvGmI5m/pKW2E9wnOQPaqY2KwWeLdqPUwoQnZwF8RSeM1sVasmUbEJInf
Z41+hnWPFNuni3kvffkWKDNFJmHUuCpjCOJaQgdDIprBj2gTcfPtMUiwjXijUq/vR1heWGPvwklX
XjCboHzH06u+TZhe1SubM8i/N9re2DeF4INQ22Rp8wcK2XQljUrvOr0/tGndODeiO6MR/GO1ZY1s
Mwz3k1lRFVITqVY68YbTbqBXkocfUoUiQK2didVF95AMZh3aH+EtvSj/DzaMx1fXJxM3i5dJ6XJ9
+Ktuiho6+I/zjfs+E1tK2h1KwhOBL9vClC6cp5kjL6v0vlaHY+f6BgmLH5LYAGqZi1+8e+KiSevV
64xgKsExId68jsHSCjpllHO+VV8ggC26Z66pJUJArZIsmUI5wnwp/Vn9k/Nlp0NlrpWLHPza+T28
2Ze7zpk7i4+dBFJgvjgKQmmptPKOFylzNyN0E1Q9YC3PBi3FlGc1+B26H4zrpRJI2CSmwzSgSE0K
+/kdIaWJWfy2YbqEC74vtBK0PPr5849ivgWxsf6pVbEZeRhAW9v8Aj4ZHPP+f2h6WYKIOSGFJu+G
Gyc4ku4UrlpQfKpT8NrAtr/xcbSNMCIkm167vBG/04UE9l2AZqIP6X41eZOQY/YwnBUrXePS5nII
7HMxAd10ZIuNU6Sfg7iJQp2524WHPhLBx6YXjqHmQUKdmVMyA804wUD2Oly3h/z2t4BGdtJrf5f/
dtUhAlziNA4fS5TS5JD5kvEExxbVWwIDt44xxpdWed3BBqu6H8GSmE5pJxOO2Hs0FgK5sMfeEirI
kPyd+jV5NLn/tf6Ha9wTqmsCyfhHRdzGLAIr0DNZx5Xbpx80K0VSH59ibCz+Q3OkREYv8CI5bNaL
CBDp00s9EeKUy1NK3j4UpFQ8FS2+YEomKdwBbdJXdqc19lk6uBNe6mmIA6FOJViNU9uof0bmWi21
HY0T6rUfoFFFcWzys/s+iT3fdNT2XC94xubttFEnPLsD8GkL45ONIbO56S0JBycpRznevYNTmF0A
70ej+xo9GI0uKupNAubzel44B/S1Ht3tEYavrhNeFLzMv4hfTWUI3mXbwRVGwQLEu76JhCHof96F
U2mUOXdzrZ7vSrW3zF5+CNQfjYw21qrgrFVtNm8hdwfey0PgYRGYqFQTwaPWBoz5r//xIMCIJwQa
muYYIO9zNJmrnYOEhJmitybFxHkWhbRPlv+HIe6C55UUDxTiKZ9mfMVmHYwpYH2rculcL2bMQwiQ
uZ48cR67qzVRMEwDZkjlrlUm8CS3mrWRSkHjnf6qH2oc+tE972w3sq8/Y4hMDLUKuKGP6OIKUEs5
ZiKywBB/geAlPAHDeVs9PnytbxtkBRSUOf0ho846dmz+I0mQr/5AZeFW5zXcC+eoWYtrASvn9jDz
flAa82VJQAUv2Z5eFGp8/gM6l0bSZTbxU6WZyliPdAqZlKo82L637ruSMbAbxnCEfMnla/4imRdv
ms3O12u8OPMINgy4Xb9pdqZqKKapRrjhobjmI5w2w9Y6GrFiU6Zw2ZO9mbWKWGN9A/hwBHAvNLUu
LJdoBtnodlrTuy4E2ZeoJ+nBBOPVXqb4lC3hXyIBpZzzG/WHalRp0t7kKqAkejXg3ntjL/U3Fw3J
BrHshIgt1dHYQC1WD0Ao3GtlhzBIbVsxb/q8b0e0RIc0n7hBts+RmTw5Bl4crWwr0sF39Lh8QPgX
LOM6JKRDASgkpDLcQcDsCt3oWdZ09tsD1Q0vp7IWIR22JMvujjT5UMK0VAr9zC4vz8IKpgG7WdeX
LUp7KbNryqhTN7e9ThKq9JWCrmuf6bodLv6VBnmdq9xnBsCf9IQbbdU4Ra+JdHV8BvrXp+1pkofP
Wk8uPKL8a4w8ReiE5dRjwnRuRthnCAfmOm2x7OqYLKPtwIIV1rczdJgXu5wIT1h9u/WZhaAM3vmM
1Z+qvKGFCbZUxaAFkJMbOeXP/ostVUht/My/u7Mon3+NSfb4XM4g1AlgVXHsje4LVTb+X+7kBa5O
ADPNlrMSVMo6lt8kYHPP40OUflq/cY8qpk9kfmwdv6vfSfb7XIBNhITX3K++bguLEHXe3klSeXFY
O+/rv/0wq9hnPgBu8h1HZl8Z4ct0xck2wYozKURxpHoc+3bVb2qR/t0gy/NTOtxi4frVt5Oe9ObH
m0vxXvqewq7CrUmXPHCSoK/6C+77NWVkZMGFJH8jgzrcwE+mHmN3eOi1nX3LcOyQ64LskAy1J94w
3qzT6te8kYhUwVWD7cLhLgzU7jgc0ZfD1gZ5OsKihoTd7nx1wIymaErxcOpYp0E1ZXL3mvJKRpgI
d/KIHsBodP0jHe1fd44i5YR79J6rXd76ItLtZCAyhuO9vb2Kjbg7onZ4apwXVu1t2mzVu8Z1mAg2
WRUnMFuwSjJTrSVstbVfjAAaN4YKkOJO2D74RRMAe2OY8cUg9dh5W75PQ7j00Xa5Grddqihh33kc
uG/VcRjWQipjue27YiRJqVhuF1S5UYL6E4aSbUN8iFIub9qgevIla0FpRDDgKF2pHn6TC+QrwUd3
FftCRO7bDC2Brm6DU4lyon7/H2LL47+CS1E5Xpi3aRokzWe615ZRGvSx7BpHrxSNCrDoLeWKE/tB
1F+n7Irz76KsNmeiGcsz0qGVzGn+zokLSP0Ca/xTj3kae7FGtKKbpzr0mdYFzfazUw5W8fQckKUn
Ms0HfYewAKDYKlDLLoxgGV5pb0jwY4qfhwj/f9w6UwRcKVOo1zGT++UO01aDfcg/iT0xTKAdkTSx
RWk+Zes/w87BTrSsq5VhD5eSMQ09QdbeGydrJaXcb8MfYkQOrQqGM9UPgwRDl9RHE7tOjzH+Z87K
OSyAMXH2uQ1WrHXXk4j2r/NprHtsiAfA3ERVgV+nX+eKZ8Fu3AGpEaU9HNIGL2349GDgn85vRxth
AA+qG7kT4fJ/cpX2d1Rh5lbMht1llvgfmPKKueUYC07jVEcFENswl14Pj3/YtnPGNCIAazuaE8nN
9+GL+4sXoFll+lYnzt5Y9WxiC4fEeSnneG+IGGSZkrmFhN6QoXrS8Ewwaq0wLLDDMmo2JcUd1Wj+
/xvH9JQrwEy/8JsWks+fsb7xJVUjF86yo2vRtF5eGrdPoJJy/K1xCDzX+nd9Wil1iAOzFGPUzVc+
dMU8Pw/sappfPKq+jcZraDnGmc0u7Acip9TUBRyIchrE5thFI8FcVhpX5MAJPffL6ucmvEfOm0bl
z4deLZxlAMMfO5tO+iLs4TvyOjs4vBPc4BwZ6WNv2eaesQwf4r6rkTMojY6HzPq5Haze8isgesvm
prZQj0vpsNnVGUG5Mo4e0OjkCmAYtg5WQBp4kpkRS57wmZf78/mQdh3V6MSDE/2nF3G+X5j8E3Rv
/aMKWbPcZcpTLGmmfFFYY4wbGncO5ckWFhsLD8kkfcMPtTgSwy9uCK3FxXqAOyXRycQKXN0c+xXv
PyjjbpPhsxT4U3v51bwV2pTB+QShnftw18GbZj8RnL2JZ38nDKRA887/0JjhMv6ocOwe+1jI0nNf
Pv8o5HQ2h/FMuz89iRjSKGbgeAF5B/PrrjGk3+WzlSxtxDD1H/AYpV2A39EO6Zok1SNGqcRiTJl3
k09opPW0DevE1cUUtc0A3/hXjM40DKLzoEwDhrO+6HfGPstOyuHGqH6osUETrHcwEEY+AhFqAv6T
9pVGWzx5udBDuVEAVKqoawVA0SVrLOdqg2SXDs5AK0gbvdfxzLSC1NSBW1+epTdpgIj+y6TDnqdt
ze1Tto01h1aA5h1MZmw+PxOFKL8Fqpwhr5TBuDN6bcWICmvfDrK7k/m+tCdVPTnwqyKo84IufjN2
a73Kbnb1gbXovI+YI7cVf1wgimB0OU90ryl1BP3BDSDT8rcdOjG1u81gReFoRqkK54rYk9eyTMDc
vTGJaoyEsKxS+bJeSroJRzCfVN6XhqyAx9qcIB/BwIh8EB05GiGWLLsiieP6hZVR4cn7O8NAzC6e
Vccq3xshMe+lXMneNUsVBi7b7GYNMyyuD9hRGk+rBYntj+5OfmvEZXWvo3v6Ycc1udotKZxCv9fh
gqbZ0EXiatMFyR5C5d7ohBvLxRtmGKxnThbpip83jyuK0PxElbh6PAAsNM/atAsoddvHzZ6kb2e/
U/spzA73nItK04CSL4JHflhpK/Nlik0yEyhnKSosDDRixL7thjmtPek5RY5fnHWT18wLzOkBKcVs
s64yBykkeTumnd0FqK3Arur5b7SafiVZ95wXRjrHrlix03/plOuqZdkaRlJvISjZ6be1sKFvQm3V
G0QIO9s+MiLxDJIRBC4DQ0Wykc/9GIroo3aLU353B0cqWxvkhDL64CDp3mLEjiz8SWTcLod+ODX5
0jq4dWcVFkLlRS1Wmt35RFjCWfOMAt69bmn8DCcteqtofKk35y+yP8aHJee8an92dkZsA3pOFIsd
0qRqo7ZQc+9rD7C3DU7OCG9jwC+0XAnEUPJrHZKgWDPLRzcQGA0QMFtqhWcrIYk9aeHCEIgNsoMT
YreAgk4LM1YtSlrNbVYupi/efd0O/caV5rF4FYIzxgT0d2szVYl+YfXLzu8u6CEp4TRU6e0Bn2yK
ZwF06R+0K7qwVTUwLh8ICVE1BpWCWY6W5YajvjSKP3zmyDT7I79DznsbCLOdBZ1aJMOw2mYyijoK
b2V7LcWH8E6lciugmixhANtRvKMc8weBXtKZuSLFYZ4a7oVgxn1YO0Yx+OQqJakxwN4yI+WlnoyE
9xPnKKwngzrMcf50pD74zAanJrbE+eviPufc41ILx7lvSfJQOv65iv36+7TaasiT494BzYsvKDX/
d3BKCYdBGD//O410xpzh9ZUARcsJfbPSQk6CBMK13uaTnjzs+7iv8v+9RndGSc+FVYVJ6QOhFXkP
WFsyyxQiTVAPY6TPFoMuIiG3ZpKpasZdHz7v6BxljNaYF5+ALraqzll8ugrV9G4CzQNWidhWQzkA
SD3oWpwfpxFals/3EU+1D6zTypbOu1cgD8umk35jIvq25gZSRteGsgjVyifmB76t6Nk6Wjf94aC0
LBS4MlLCgV8yZW46fK21JgKEmlK8S6NwATE1mwagZ4r640HwhkW6eLXP/t10sOVQotpY85anUwwI
D5lvyzcSQtCfDq2in3fTwpl1LGuAhPWDV7DwaRjqehvwO+I4dij3HcChomQ9URfbQmxPyz7eVNnC
0CUshMj3pcQPJbCpxqZ03SKuZuiGDK60Me0suTvo/OPEnK0eri3tswFmdtPjtfHXEer64/siXcXJ
kMqH0giaZH2MYMhFp3i/r16LI0jE8c+JIXUCYWdx9reWek4KgwchKf5lY6Adzd98DikqkU+0SJJM
VOBIx0KpRojHFpOnlIhtX8csp8uBzaP+gt6gWLQnEi2LuSjBEhIZw9kqlvA1vfUB8qDV2HhbjTur
YrRRY5PL0Soqds9QDM6afWUgV3VkJJkkTGyteyd//i16om90BxSpqLEfhnvnLwv0K2vTuCpHwU+0
wk8fs7ka2Ol0BTxlj4ZQ7ZPWY4UKi56lfHordWrXmflR/dMNrtX1QzkEI5iFWmjo2wya3C2hjt8Q
+7/CKTfYAlMTWPhx378l3g1Wseqbtl2PEwfaeXb5vY94cduzWo7i+0q3V2OaPmINZAlVQeWTGcVG
DWSAknxmgdbz6WU7ZZqcbLNaJrQGGFGVaUGhluoDaF0dozLRrzxzxRs0wVb4PB/p8yFdz/6nQeIO
AJgvwK1UMm6aGwytS5NEYQDal+Etgu7AffHrU6UmXFRxs6iIhvJEnUwJ+zV7fZvhBMpqrKDJhXZk
MMdUppemSqI6a0b5Sa14eDlpJMfNrcXpiyRoFJYUenY5iexcmMTgyfTc5GBHJzQzvjoqRTyFdl/P
k4WT4u0pudTDwCeGpNI5B6ZFgjavp23oQ8qT/zS1u914QJ/K84dh+AwZGZI6NkDbHpseMa+JxPjZ
/CGv+SD4kkPC/nFUaaYT26+kc50UCYHQL/0novkaMcYdNRGKdL+ddq2AtDISoBc4rlFEEdOp4adr
VzVqpON7DqP/hNe3rub1EPPiKPjlgRzukQCnAx5ZOu9bxn8d1UtWMn6SS5j45ZkxbasuyWaxI/kx
FeSbTd/zkxpIJnmnNfFyLBHJPeLF2d2Mx6nIVsW+zUh4LH7Y3qGG09UBg8SA/jlfR0sOQIqJXTz9
9tNzQq3B51Py3s0reOTYivW/3cFPgbeLiWek70ITlInrDY8Q0Z1ZG93dZqgz3TNHZ+bj3v+bpAi6
DsDXRQjwmWOexlx7yQUoSH38MgZvmIoWF8eo5cUmFXhGVf9MRDEvs/pJb3oCLSCefQhxSYIyezBL
3uEaY4AIyInLtr3X+qtakjmvwDYra+2zdPoISPikFpkm5JlvEKTZvpQbngkS2jPH0Yl1Bx4iDCPC
dRpweKsuEAXk5yZ7ho0Br10cTym+WcKvBeMMqX5kHdtjWNeVrGP8Dsgo5BJlavBn8Yne3PQK6POF
jEz19hKC0bOoxEEqEJcz/4ZX+FVRDtLU3MTwhEmPQXBCswhUKlA2ubkMtDMgAfnee1LCg3VokeSz
ESIMZWulBWeC5p+DG7a4GKp9OWIes2HyTF4NZhfYPzSR5Hi5+MuRIqm9D6Sw00axzlZBtsCZ+vuK
eExj1ccdKHaigMs3izd8OLThXq8yA9aRF8uaDQa/WNCGJZjGsfzGLKWQ7eNw9X4Xbn4FJZbxu3Ig
8GiqkHRC2BlEKJ01ExUM29jMR8j4GGxPUO+9ROBixqFARYiUdCgw9IHAlXW5oAHyBrn7rENI8phc
VCuap8um/BOqSFwiDZXDTsQkkUxdlI20fBiGpqNl3KqBmGM9rTxcNQphs4HHY8HVaNyKJx1b7BHt
lDkWmTCujFtL0CFgOc/a0fBPpMxRy2t2D2cbiBa4A7XBl3I1KzzIiRzBKIi9U4vcbn4cuxJ7QftI
katFFo5fPDtDHacew1dpyS2bIrAyPPLs9Q1Ejod4TF7xvnzFEMQrmdk4Ue/6CqXsrFbkvSASVA01
oYO2nIpadgPyruOP9sdz+izPgWpQ/V1hfg9PTzBZPQHE+tPYLRyFzxFJjUjRYHtOHmwtnTTdV7gf
2NvuNzK9nsRbA1tOU7245EmBMvPsFHvucQe+oX+8GOwHw3tANS3APK9x2N28Vvp9nfbgnwoUBoS6
2OmygDLheGmupMOjhdsEnkc7jtKowUIoSv/0KKXz3ihZmTC0NN+1UbHLYgX7f+rwGOn/kHCz9ENr
lPV9GJ3PU6KE/bkvGzOuAA4iMG9J9VrbbOSksllS5ZrwqCLnN4GztUwQJaDomXCuMvv/trtD2atj
hdnvcRnioEHkHvxffQQAuugNkTkD4+2CD1iI66Q5RrJOJ8VJSEKuW/2CTM6DBuRFrURV0SYOB+Da
dijL9ae/AnB9dND7tKKgifJB0t08C29aadKW1kibXSeCdYONMBorlocc67N+XpL8J196dQFUjm6X
x3QGGbtlbk2A8iJMi7/mzfP99IIWEWZraVjciXX4AdSOlQlwe2vgVlGw8FfHB2EayC0tIbAEqqRY
ZnJ7cpyPK3PIdX7jZ1QzN4BrLfmdeUBHOgIvuG3ZkSAA+3r6WzMTeA/IOJOMAYstSRuXsm/JF1aD
KBEBWxmZfM/JuAEFpwx16UUitv95zkxhLe3cAEXEIWlezpGiBjdbVe5rk5lFntWTHd/cY0MW6udT
Di83TxKoVMrDUfCtYyxzU2CFgRlWu9DBeu8IRq55ER2q/a/AThDokxQ1I5w8mkkcSg2Q6LlPP/+m
Gr/bQswHgsurTEoowNp8G95o2Kitj4VuINSAbVCkkpUnsP74F9zZDfXqaSeao/7XR+WqavgCiTtH
8q7o4P3AUfey2CdMjIoj2I5FQ1UMFoJhLdobG3POCUWs4/vh2vwD1BkGAHPa/t5LbnCMgvTvNslt
nx89REyl3nyMG576oNiMXXmgLAy3uNywO1K2goEkZOA1o6rLe1JsTG45QOvx9vAMVpAqAc7Ok8gf
AqwpC8M+o2FWHf4hqkc9e6rIutkpRTHWRleOe/Ew+x2kauC5/qObDjwZTjk8aIVNCtvGyOug3fh1
NkleOW70vTwbAW6NJPHWEk86wBV+0Gg9IMuhd23KWJ0UYEHyYATyIt+8M23Ez8Wwdb3ucBYP5chX
j/8pfJZoCuiaSyV2gdwqWg3UsbNT2raa8R38V1FIQrVA0982LWQxF0yjw1RPkUY8oXGztEW4XNeJ
EAnMhNGzTLf5oo9oGdKIE2imLdO0b3egaelRnfuyN4BgzAIvFyWNTzbzqBuySE1Wg/wLxEkicMvg
kbnpW/lZ6LL2Su2oxDzrn/Phbq5WpvLNpWQGG9vQ2LSpbSxroq5At4SNaIRcyh8oTYpWNFyMjgpA
KxtnN0HuxHK0WBXD5+hoJFJvDsOkjdg5mpOdqVD9mfP3x3BsV1ojMwBZMDPQgRgIiEhoSce0sM2l
MOmjfIkhFPY1R9JiSJ7sgsTFViab67hQ8Cn0FaExa0V2bCw4KqlsQU2vOoD/SBmftRK5qPZbRtkI
hOX920zMEDinx877omi7w/qumDjCZXsP+1CsyjIg9La8mPBN48sk7H9H8fHtXvhKjrIe8Z8zTfvE
wGQztZkd4fjMxJ1cB3JgKIYpHSFStYfF3MXRM3M0KPFJW1Ai/SHZiB3wyUuOpn5RF23hVEW3xCK0
TYcxPx0krCTQS+1LS23BELBGZCSW6LYxoZt8Iswdi8PciM/EcUKqjR+iElfiZdN92n+yIKbuJUG/
u0rtbhocIoZWMoMMrPkY/feNMK/7JJP/HU7XGD2k2maOqaQ6JzLexkN8qy8+ydRI9ufdb3mRMLZe
h7VKOrqKB8kZxylLgn8J13qqJjZaNEOeWuAXVndcMkAWOd90H6bsMqSPKL2nh5pBz9hAbXOtxGiq
idphZkJbx3e+ZmFJ5eMMLM+symLgOmG5eZyYfQfguH561jcp25fd5QeaKYaaH1ErlI0ao+57+31W
rMUlh/oRwoPiF64eBMlkrAPDAnL2Ue6NV+wDVq3nl3LAicP4+G1Ke9UQngfEsckoKrryxELikM2g
WZCRj1YNzuEibLFFE6VZmL5P1Iy0phb2YNPFXkhcXt6ClJaVqDZshMfiVfvuAyy2mxAo0/zNWqE1
hlCaHK4j1prjKCZbV9GUmRk3y7BJNhQY84Kjr75njcT33GiJmIo+YulTxFpL3tx9UaUuzfo6kaK7
xNeasXS9xs5mjLtFiXN0TqQjuoKVWgt8l0UkzjBDCcroQbs43TUK2F0vYXV25Q3q4oeabOj8zLTw
rhx+Xhu0BqXorPynpBTSXXdVVR6ZIPsyQRJ8BbuLDLl2YteS5HqVq5PHVy82mu70vmDm22LDlgtC
8QWmt893S7AnJD2rD0YIR/RyvL3elCGjdvShKQxEcz4Gb6FTwUsF7UPDvfw5LQRZUmKlq63Bz83U
WZwvF5a+w7AUtU554rBo84aDGNAomk2jbWoTk2ee4J6UKEcDov1rWVaPcMxX5L9p/aVkUKorts55
vCR//yKD8wQczgYmjThM8t20rYbi/PITx+s4/0NGG9GIuLxKWPyOB6UNxVfTJzk8UO+BGGTPiTAO
0uTe6MhbsYJcl1KeiL4WG3h7qCaXtsyYjRahsHzFKGj2LM0Pjtve/bSt5LkEVg5PwHtHWQsZpzpr
l1jCO7XRf7P1u1im11eVTIMY1BqWJXRzQ4b3LG5R94vnSi+ntVZZCoEAARCTXyK4ciwVcDmSwvrk
xMbC/MYz05u/+yvMJSwgbrasYkrK1/Xk6xN/u6NZNQcIQ4haMf04Y8xX40XATVziiA3aBrScyTos
DJ8XcaaiNLn+ppTH7Npp//J3lK01rBzb5Vc2wtsT1azOWytqAdix3Vo3BhMXsXUNsMZMKQYxuwYw
IvH8mQaEfeenFIIi6tkE5VyL0TxKE/ktoJQa68h2n+PBb4mk2PaR7MVPCUdWpucIfAQyOmrauayE
ptPY16vqy3Vt03MlDh+zsU2eXUBDokksvH4YeGj5bGMYVP64KpwSxoNWLoSKjG8XmU0E4OX5J9Sn
ySvlNOSZGA6ndh9Uv5fpBLm8shAXnWxA//kKUIfnX8kk8ZCxlQlSlV7UxihhwdJ6wW48OZbPI1uj
XVMMVQPdgOedtbnbLpfEOqNEoPnhgEWen2ugFSHyKRKLfEsdbmTlkz3MX5AnwvpS4XayWyF5E98m
sGat64+Daq5+D3X/JzI6W20pJGs/+NEkFJMfVzJWkbYDCWdEFpp6ODQ1Nvj1nVp6jiUTUAwReQ43
gFzpc4IcjuSXA+832iS0Wp1gbC2H8tMaNNdrfrBpawiIPNHc93Faxi3f1Ng5w9L2xG3ysHVQp/mX
tt+vw9AvW+81M4e7b47LYwOS38eGJTdjo72G4wnyuxnaRI154GFz//k1E2R4PgNQWtJ1Dcsjh576
85nWQhzDomqHkB6yP/iMcT1lY8qCQ6kPip1849y/8Sty7AYdTHJbJOJSozVK5g9axnL1soEFppJU
uOcqtWn0myl/TXP6HYXlisSmJklNaPMK7APd413YC/l8WEEdLB3u9d0TxZc2+mtaR28qiy+oQ1pp
q+gV03XYQ9+1/7zDNF1PPuU978NmiUsrRg7JYiRw1CQt9xj2KsdeBIts3wao6iqkwaac1Has4ZWe
sgY6p1dckXDIbF7EPRL6ZzJsL3xQtr0dkmvGexlZ9sf1Bu2uwm0W1H7EeSBTSwy5+KC4elc2G5Xn
9BuFiXPAK8VhhsyWBQOxeb8D8DBs3hV/q3+wd4YcEgx5Hj96Bkrdy889utWYcT57oqgMCB4KxK9S
58qh1RXD+KNCTuKpnozk5UCfD9cBWEyNOvStpLdCFlOO4Hvf9QFvB9GXK1KitmV5yEyNIwu83OhN
JoM9U7pFn/A/k6kcPhMO8RRHUEKgdQ3VLmNPdZB7zpf4Gy7UxKf7JgIUeUyS9KyzVCJaFV4F/Z7e
ZBUfEqIZolPzsUVrQe5R05bDApbKEMmQ5Pq2Lf3kQZoH5O/ZyQYjjiBZGCkUPnxuRUKSh3yDk7o5
p21dhEKd4KlDHCRwpwgdT57uI2Z2h28xQ+5XiE5cjwUKXwsLl9BKQs4P+fqLKAdJI//RenRoRUoD
ccSb6e1nsiovCaAK2RBGObPkpxAzdWQOwneJh9+DIAXUXGlRoS/5ukrpATLBPNptAEAh0q7T/Szl
666ueRlYWwAdKYDiwed+ELc8ETQL6266S5jeTV73CZQ1ZGkTBX/ioW7laHgU3U9bwRe4+VQz/WS0
dXC1MKu87iQFSFkdYDG1wg4R3NnvVrKTuhQyMDnHjkNtnEh5TmhWmNTDfWdS/JHIt3PkIK+ve0/J
EyMN3w8jDcmlJ5VSzUY+RZ7vKJWweu7Oi4saqQ1h5ohTyjVhhP+Pwf3Orpizf/KjkRHgM26F4xOx
Gn0FDRYIXPC+6XyO5wTbl0yKrqQV2h+KDJP4uvpjUPkfgdZCK1dy9pPM6xnimKvFxiSW4hl9Th2R
Nb31/ZjIiG1gH0PhC/sbq5R3ypkp6fLxDZuzTxFc7EHTpQlrz8V6s7YdTOvofYPKYwALw4RN34Dj
SCoey+DnzbJIQ0H+e24Ou37eyAzN1C1ENlhaWDjVxjU+exWYXdr6IrLY3smoWJ3weTGd0AZrL2sf
F5zJE4cmWsgKacsR6RYYTmbJLzgFTNZER6QV4ggS2wVw8cQVmvH4g0rSnkNt09MJSiSIAONyaZVt
KiP7PKEg+YgNYTzfg90rbpln8yik6P05A4BBGUdUEW7hUveIoQIp2t4Y4fJIEOTW8P4hOzXqyTSB
vleLAEjIiPrfmpywxeb67q/SXual9i3FqQ1/eRBQ4UjiU8JRxaVTebOArqtSdnQpjEBfrj6RdJF7
9E7cSMUxipozyiorOkilYZQ7I+TBj/Btz968wvnYvscfSQTZ0AwIPCMMXoB3nXaVHWX8DAZYEPNQ
c5+BPYlfOcnen17vKS52ezKo/BhlsfeMcWI0gtmXpRJZYx3Wo7P+G+ikc07ZdmW624Yxe+5sNfqU
113puiS+QfGKiQ6w1MYHa8iXkwiH0YNJ/lFPIqJ5aYXTewYDlh8ArXfpJRVixIdjYEjrvAVb/7iF
4PKy+55CFJcYV1SaA6eWGe/7kZvzLzrJDQfZOKaWetIHzP8zo47A9Lk4XCnvhaEg5vZYnOHfyOff
O86HnsRqtM6nx6OjaJN/O0k4bf/TqxHZm50B2mC1Kcym5zq5tQhNn99jr3Ed0Ld5GmJuRG0Ka4k1
v1mFuYDnwtzXMekgR2o8oF5+Q7PS4tSf5pjTrN7tv2auOAuBRquOite2k1YuJaOHZae8YEhiJ0Qp
ehFEkKk9phBO25KmuyDy3CapwNqpmPAQNtoRdOlXeOvlYHTwkcGvM5rTHN15GFkT/GJYWXzJC3BV
VJXeTKmhZgBz1fXzwBX0Oo0LTFjXenxx8QTVl6PsYOyBh9D/PJGA/EikSfYapuDe26HZQprkrCtx
kjIV0PToi9wgmP1kGJxK/G1eVsQ0/oNYSona2hJ/pFc86IWt1pczC2jEdGQT5zkoi/friiYSWr3A
SmyF0SnjR6H9eMHQ4AtJDNiwvKFdfiLOhChU6IL+cOl7EM2vfTVpAwXTulE6asJ/yhkZUF+1s/OJ
VZOg4nytHrXd2vmLb5JixMYBLQhmlupYuSzEDpj1S8AfUnMQUA63uI4VC+EjQeN1++3cjlX4H4+u
McGSNzrs8fYetXPcEqyvLoHM1zf+PMnevCAtZ+yOCPh8Csqz+FQZc2tRw7CIZv0X/e7HCopvV/FS
no9atUO/xwvXgzkIkHlnwKZrt7EaABYkRp9a0jZO55KI66BOQOOk37g7IJ3/HoQ6AMXD8ZXMVW1a
FxkAABsmSp6FEk9EJd08MdUftg8lc9yqwT35NO8AE6cvawar7WSR6Iornck9kN4KC2P/G1IB2nNP
bnZEBYLcJSdSGwCJERBYXhCB915F3k1b7aUI0Kk4IcN9Cu42u9OFDHBToXmmMLXDHBKWlisns53W
Xl3n0plJ46Yt6OxTT69/Q6cxPUNR5auhWDtsKn6G/gJ+6GHkVNIYOim2m0a0io1qq7PpbY+dA4QN
9nw1TG+zmH6vuoypEJBAxF/JXGXJY3U8x+S03JTbfl9S+9IT3V8lCC4u72vKOgBvn1LYq7gpvaMz
npQ5zhqSTLPjY1s08gdKcHrCgCN0e3OKLcg8yy/T/ivrEXaS/sLIQxYjdMStrFSrJXLHwWZ/Dgzk
jqCncWJMd/2gtagZZvSbqPPV8IRk/nwt9r0PXf+vDmDus2c1dHB97Bz/xds65jjreWt+LBW3eLfA
FMx1UFr9fNjxlWEuaJVkrYfB48mjvFxANSDuNcD/CsWtljsdUo9ThjMvepzsjRh4LnDUZrBeDWH1
jq287wQiTD6jAvPOGHqnFMYb72m6YFz1ZAA9A6lzeW47SQ2S6EySnp48uHjyraXm2v2Xzp3AToiT
H7z6ZScaP4npB4Z8aXEfvZqM6Skh4DbArBsKYqxUboPsDBhEQD4BD1B3zHEExYQSUOUrEVykDL/a
cNDf0tOPmx61tqHvejzwl7TVXD2n0OtHs1xg6JPo8r8/18pFUmSMTD1lRtknYI6AwNcfEKaHUKe+
UluFiCjTaYZyoE7SevdtybdHNnbzVNpz3dsFONlYKAc6Jqdk+AgLwp29RmkYgTobSAmnKaABGCeY
mZ6HlS4ZhgAwOWuAY++b4LAEwviL5a101Z1GftYE0kJpuTOOLevY8mHydLEFi0VfXIK/09tRfp1u
V/S5JDxCUiyx8RzaN+AyivFY18p3nfsWK7ate21fMeX4P1Z8WJ5RJveNMDe4BlAgnLXTEk9bWt+c
ovR+gb6G/UPyqiT0zDIroQt3Vlg0aLNuzUhCFk+ESlYM9VyU4J6AuUneUsiKbW5gxHILg+x0SJSC
pNZd6RuVME7GYS/7LqWHR/XpmsXWs3lBogZFDJP4YyQDHOAXLda7OpXLcbJ3iTe6MisIGbXv+G7O
Ve3jY1IuDhLbxqZDp5lSJChdJREvKH/HUTu0yRIlmj1qbr9dufsJu9qQ5nnImDi4Ozi1878lYsIB
8qjOSLLobjtb4cHLa/gU7zxYHNrYWLOjqFkCRkDSq9Fk61NzVGcfsjDg23bei7fR0ateBj7hr2cw
lwzNKZ9u8JjDVgJe+QcGNPdi+2dnLBtS7zYGDvWehGTRAcERQDMggBBf2Gaj7owypOuDcGt/2NKn
C/NPy/Q/W6hyCqAIa0fe0W7FEvsVmSDperofkp7UNJg77QCOp0RNi7cgGlLJ8F9YHYEwVv59yEGt
WkDyGF84MybcyYrEpnuVOlHpRrbSL9xrX79J20JdkCHmaD4HCQXPn9lC1iPyOBub6BQ5iHJWDnrm
BOgs5U7ejb3ElXHu894k97BoeA1sS45m4Y2/TfErhES94+6wtBlD045v9ex23iWB61va0ejfIMB2
ToJCnsvKwzeUlN4NIuVBh9FHVYkAeGWUO3HzJsKCmN4G4IADAnTbuuOZt37vNT7soobhZxfRDaLw
j4kKbdxNftdGfxXJBxQluwY7eP/kHgrbJx1h5gEnPLGKYNM/viBlTv/tgzRuxQNwo6H3jh3lzv7C
gvOxF+1cp8V46LCPeoWAt28u5Om3gHvWxMeDUa0rwo3VV0AG2fRO3DuWzVrq+ZHk/me3Sk5E+lcJ
AWJOwp3HSgYn3QRwk7TNkN9Rb8ot/CwVeegX9IJaCWf/ChvZijw2R3P7sEUc8lPqUsfVc1hxh7Nx
sSAYkMBlPsbqs/8/SP2M3iRtDGD6RCZ0CRfL6IjJSCtrv5f5957oCdeA8R9zOHrreWSo8IX0lgtz
+p05iR/R4pdwN8Yk9u5MjDHqO94BRlqH1zkue59MWaTTHVGa1ggSMX+Ua0RdX6T8NvY0ZT6sZfJG
lp230YpuCeSRGkTc0vcTMv+FkjTTjrvBvQp+oCH6CM6YxdCILUpr+b8+ireErKyySSsAM+x2vm9X
aqXYv1MHEYTheo4S2o3KA/umjiUjP010R/MxiYh3cjfmENgiHjS5RuG58wZeDEMJ8K+U6E5vpQqy
lnw+TK7CgyDsgmWmpbLhz9fCjCul5olB25fvPi4+KPXByStzh7c81dlti5nwaZQl8i16jYfcmFqF
0j8Y7aZDAQN33msvK6iOPy3nZg0qzR+JtsHPf8kwFSKRPxBPRHbRn/+1UyvrfcMyN9QKg1eXHkLs
wWVgzkHJyu6QJdS4Co3npb7zSOOfo56P7/ZOrv8SB2lqNgEVbbZ3lo4/kcty+dbTtsmEIgsDfJ67
Oh3/99SjIgSitVAV0Ozx7EifDZLUkkOXT/TXgueiHIhPfc0LSO1kmKWshktd0UMbUN2PZkVCLzXQ
E7AWSpwBiyhF3xA+fFDaDTIHVG6t5pq15JRWcn3Rb3j54wXxwpPcvH3xW7LEkjvoX6gAKOELI6Bk
lgKNfEvevAz5yVBqpHt4G+nWVRzowjUBvRjVhWTtKL0sgaFuK7RW5xhsk/e4S8nuugBioXrkC+nT
knbdoVw2hIfUAytTb4VdzoGf2hhHit4GC41agJYlEZyLf9Y+rzfxDIEf6+Q/75P0qjz0tiM1BIjT
hskmhCoZfJr6OVJ/+jMGiXXhHMtN2XSDePGjXCe1HoErcWXnzAJ+RquGVZ43cYA2IZygOXRENA9D
u4NQVdmWXAcdgMPGdn6aXtvdW9xy818VcHMOz8i2UkhEEsIJPqeVhJbo1C6DE4j4Vq9RUNV2avb2
JL9zroa9YWwoXvAP4QJHCQn8zNjxNg1PJZbIrgU2DcxqPRRMDImjhjJTK2hj7y4THtxCamhswaGV
2gkrjW0bzZtQv17dSMuMVHKN6BTLoCfGZb/Y5/X6X0D+HCczhXFEnBtk3TXS+MyuNKercBixoFVi
TqRQ+9whOTHSg1VhGmX7JaTKZa2z+szV9me9DkfNFmJL2BACP/DkU9pHRUFaV00vZeXYXVnJWKI7
F2imu6rXFx0wOEgyfuuHqvuP3EFhIMp7H7p6ZLWr8LzlaNdQzEZEET99vLt6otWZaHQWcc1gjMSf
UpbkCueP/GZ1SMEldSRj7bBWhWgKQK2ZWHz/DhA7fCe6EIGdzlTpFBdl8X3s9t1LW1/DpgVb1IEl
VpcwubZODVC3zNZYkI/IZQzy1f3NAiUOaF1z68qDqwpYW+HqoHqqmGr5VqTSJcstE+OoPWUBVIrc
3PWZZalbjbhKXSGyX7LD5Sx5eXSXvrXs/jpf9AeCdMDEbXdf4m08U60oREBFZX1wAc2TjQTmDpRM
C4R9jqDOxgYmSJBzZ8D5H5J64NqBhUmXXQrcRDtWfJsPYhj5Qzjjd9dXJWaLjmW/KqXPKHa/mAA2
TZtT7nTVRTyxqTwqf8P+OGrS7YTYybVOXIRGiiKzIPlIEXtcZywRTQOVRM7sQC9k0odVy2sa70Ga
vIoqDmVFT/Kxykp/EXdu0mARmAuk7rRF15slXUG1+2Y1JiBiOARhmCPz++1iwUz6UaQfVoImtfW6
BPsYF3EmH7Q6rzAXsLz8fBPURKN7B7WKG7wyXoCU5iriG6/pn/I9kxmR9zMjA1djOsFvL/CFbLcp
H/tP7mdaQWtaaMcSE28wvuY7ujyE9DRHvguDHjZQ//MEGyOQRFTvnEnxSVNcAo+TSmVzgmxVMNL5
UuedXg7ttBOkRzL3jUQmEQd/3CVGWGtmgBjB2tCoQKQejaWSNLD+SSRLXatXYuN6O7DFZdPNRyU2
ysAtCPhY4T7AXPezLXsX8pcnRZK/BaxN4EW77ZmtMRPH0zCWKCBj9SHHiA4OmQnJ5fK/qiYHtU5N
WDYX9ZKhJJN+PSaJwDWXfGaFlCNIB+XmoLZy0QQi1sZDOD6g+iH2Ozi2qfPkc4nJYcicWJskyTua
180nfVyyoNBxoMm+r+E+LykXx12yP/14DXxJh6m3It7Nv3m+vHJhjBa6SE/be6E3SWIvax24lJvG
zy2KpLWVkS4QZAPzWpD6xLqOHDOWSPG4n3BErhhNK0nS+rVhl6wcMO0ZEILg8UAYjVtRtVj8OnE4
94njvRe5SYhcb346PuDX3E+05ohj2nrjy79MzxDj0664wKaJYhsYNFpVKAysJVRcj2cWGbTrQrKG
Z58+Hc7LEjIvCdp+vP2YU9oG7ppdOYno1q8HDP6kmVlGyowRayLfx7NiYEfR6TuSQXb6ftcOrthG
UAm1HxDo437VuL7PFsQcNxoIHzasnf1sIMGwMu+UpHaFFapE9K71XaqH/kimAtfSqqXE8LHektrF
12V1Yrr/i4FxrkcnO5YZK2JGhURvdwwJFEoCwSxfZ5deVRTtpE/bfgHJJwYEZNkBaKFhTFQ1d/+3
7jf7hfOfAf25zaN5OLplTENcBYUprNkAyjdhTPS2ChvMwmsBVYWxMkpTRqrEny8DY+LKzBBkLZka
GoWxi4WZV5cq5SIRzWMd538iqShJa7cpcfY63F0G1DQrrpKykscADX2QC6kNqpK968wMsdv96//g
ac588NQEdssrj5Vr2J8cnkGwQvJhIvqZsqojNgAYGSsEMhyE80bObyw1RrdX/ktYUxrD+poNxpI3
eEegJ4DlvzL8w8bpUXu7ek5tLje35T7aGIQFPgNuH9CZ2eAiP/rCaMw9SygmV6I3AL7CqTmiVujC
WV4dK4qoy+ehhO5DxnFtChBDNMQkMG3EMw7uSdp+OkhFFdRLHPN6sUyi8YLECOUAxbXak/Na6QTM
ai6PMHocP51u1QBS3TAJNqvO7QVCK0PL8GlArZghxjLLUo2sXiBIFVwdVfxxTY5k7Q+dr8hGMx1j
phzbTejagS+a2qqLtlD5FHr7lIEX4NOaWYckdIsziM0bNZo/+TVreclmNTIEGK4wQ4tyErfW1yir
MYFyaUPvlRnlT1M1Fykmu5Sen47Lbi8n+WEX2DtkddmuJm42d1hNsUrXw1wYcg9lKgoRiKgYfm3C
+5c11L8k93Q+MfHPvjTccHk9Oatau7pvxjw2kIghKl5xG9fvJ6ag/J4OHmG6gvTcDBZXLCYpEASa
B/esESjauqK/rq9PaZLGJc61e22EhJyoVr4czPy5ocvo8Z5TNIdOrge5qQSV4/tZRwpBzczxnkKb
1zCbSMF1AGsLJprtYv5LmfTCHfOkHPzYpAYS9Uj2k+ntKdcNSAFOI/7xUBGnKVDGzVWG6sXe02Ue
U6ukEWvWuol/X6LcV3f2pbaYxmeP5Vh8OKzYbLGo2iGbKPrsMnsNLmdeiZy3O6nsU+qHsUs9MEUF
2NRtw4eLeu7KtsKtj+qXFPP/Ho0XDzqG8b0FBCcs/LrGYJ97xgi/Vgnqy4Saq3Xdx3mAlKzWKoMm
8wY+S4GjBYWCDH9CiZ4fmEj8YBU1BqVY+ewIbtb+AKE0FtysJv1Xb7JyTBz/Z/e+KKnk69yGbN8f
+ZrdSZJuaYg63VDrSgjx2/aO2xYU83bwa1ob/qBAJGXhJP0J9ogk6ZXTB5W9Au/ZXX6qwKhFtMHH
ix8H6CwDM94YuizrnL89EYQzz4IeJXA4UWC930SL4RJIjc8yGcGemgIgDsoBHVlK9/O6KZTWCk8J
aTi4mM9LIDOBINiTRSjT9PMEGAWrM5vK4R5TLPetAFKs6PJ415xGjIBEYtiyO3kS3Cjjvf6WsdXt
9PnhDI5WRKM6GLjnNCpdW0FdPd+MTwm+Kbv8OaHQQka3N1STbsoN4QJAAP2M47tDmjOm7j5rFjuc
rukOugyZ/0fh1DiBpj/f9rJE8Rcfui3rXKwRxraKFjnoI5vWasD0TxnUBdFKdHIetc1YJJqkvJ7n
idgwI0DeZAYmxliw0s6Ryqtn7l9LvHTtzrctIktlIYUxUzYHF2XHDO0AYd94dekWoc7m8t6Fr7k6
VK21a9+kiDGI0HTwNiWvQgVLO/7NFAovB2LXj+zoM1184ubrBwaZD+xmuoIJBzmd23bP71vKOPvp
xyz1hl+ZsX4HseMtlnS0Mew1W6U3tkG8YFlt2ty7t0yoMShYJ8yNogdCbxYe8cA74HuLtY+cmcQP
51ExUvf7ifnMGKpZ/5CX6mCNNlegyoldUFl2d71auZd674vFrvFvi0T3mTpHFq4vLhNT9Gcw1Wyl
4lTDXimTb9Tmjxmu5qx/udXlmj3HGvAjwY6oasaH3i2N+Q5iIbc2MKaJ23MRrPUWR3E0V+TmnoVI
iP75DOe5Kv+aUXOqk0bve4aV4l9RszNv+olPH5dNRYUlMzGWaBfCEoniqPr+AgGc0GE2SRlndaNm
Djv1L14QM/sbrNRi9BT3GoHnvL728FkCNvulSWAAEtrRw3HPniT3DXLljP0r3wFHnMS0cKrqTVs4
llK9Kg+hBvcOsVc+PsiEdGy8Ik07nMgD+ZNXu5V4veQHjbbmy4MgsdrI9R9N/v6tAprNxHXdk4s2
sLInzB8KSO7Ra7s0BnEkZBUTQtRoFEJgIqvlyLa3qgRIC8Eo85zFMibOnT5tMS9x7RVfYb4YTmmk
LWiFQ+zKRqblRut3PVmRU4PgT8t2n8rjg5zTC+YZWgVPJ3X2Qt5qsu1jYvVgArbm3S12gzaozBm0
iOk62d5lLrScu2KUxXYvNyE64zpdjUa3P0mmW8fAmkX0wzFUSIjyJmDzOEeLMX7uPsr4ZtB1rcwZ
3ryW6CQCu/QuyJ9D68cDph2jYVUDNHyJ1m12TN3zqJN5JDXyn0qVq96xHH826IkRic0o1QajbruK
Z3M1rFBBDvQqQMYQ0bIW4VHN7onc0AFFYvT4O72ivU13tSF3RFzVK5q+LxbG/id/cSonF+pQUN2S
G6JI5XkGyaoc3vaGhR6f6uDe73XNSMajCV4Z0BYu9w5Xzl7rNix9X4dYuZXYGd4p4icOoLT8tuM8
rzypABvig0ccixckRqoRPWYpXTaVMwD6C3oCZwiz71HovxQwTSXDW8lqdzP8dQJ3Fno0kAceSidu
PFfXY0WS3O+zTDYoup1y2Uyk/1HipvOp/n1sfTFnB65UUliqTew/8QW4JKECv/i/B4gBHzVmF8Oz
EEYWxnSgwyn7OlbTw63CiDI7U1N5GRsTkva57/c5ihKNYauRQMI8OiSK4NUkYuRwtZl+iRXFK7Q3
674ChCab/YGGLMzizLRXjbZNXglwE9hRxMQI67yDe1f3MEiZnEY7CR/lv3KNnTiI1XAIcDDCBrTm
U17/ALFje/vOD0kiobTUUo5iu3ASgvKps/J69VlfSixqC9x8YQA45GI715IPa0kA7YTkzcbeGjW0
SmIs1R898o8Oy75Kxf++HVpB34QXQhURiDTi67JUdUNiph2zLRJ6LBOqcGnaSufoPMV1OO341AjA
YWY6Hm3mXpVtFnMfDcFbynNWNXLfkcECJ6KmP6XFgiyfHfJf6HZiZkhFy6oFNzl33CrF/83L/Ai6
ycTWVeqwePs3tMgGUXc7ftwiV6QK7PGzxOubuAG0/FUW0n3QzLJQRpwJKvNZkDv5vRVzl1jmZCtA
/9X+2sP8hfuuQDuvF2XHO/yKzGSvn0X8Rovk/ec6AG1/JsALz8Bw0QcTRMF8/YtPF/Z1WZv76Jx+
g53Vk+9yAxpDu1sqn935lkSulzMD0UmdKd1wfyMXvI1q50quZ17yV7mIxHgyJzvbGr97rLTx2H6G
z4clvA8YtMNiwEyuGj0BtUO0b1rHDbUrlJds7/EMTxCbiUN8Dvxx2MggxtPIITv2elWKeCf3Ki5v
OXz2dKgyPh98FkFDiYIrxdeieb3B379xBxJq1DYA+4V0BcxQYRnce7b8XuBzNsIETIGtQlUTPjB6
6PvoSVzTK8T9EOb8O/chm2EQ71frESvyz+BtR3jC9ftzIxZkdQmQkd9RMxIi7ZUQxtrs1Br+MoZC
kjagM28zJL4+SH/GZ38wW9H1viB5y2hAF6rlZWdUXc/Rwex4NYILqy7e5qpQueTKmHudvKPVGJVw
va3Av9tqvD08Oe4vpN0ocL0Vj3ddBhkTwbnJCY77Vpssk18VeOd9plj99a5ey9HiR9Az1VgGZgUi
leaRK3I8W1ALuGL2p1laC50RcRddjeYhzFYxD1HLqireTsRTUkLCpVMsPBR75S6rixXjZwDbST6a
AvHDscQdn3umylb1F3DGbw2qms5vN2ZYUjr98wpE8XRdP2Ej2TxWNzBTIjMX8dUbt1o48Qln+G/T
pepAgtHbvEKUgVnkiIFDrwSgfACHhb0NYhR9quWQKKNHGKzLDg8m7Uz38RBcrfTjUtdiMv+aRX02
QRXZ6k+PhOmFV59s7VLXiBSc59LzftRR8FlheAFZmzel4lnukhnG2FCCqCS0/qP8uk5jdNwLBL9P
58nqplYAETOinAW2r4VlppIx0NThOrUYqUvvZrqNWDE/s9WE030QSFvLt2WaTjttJ9aAcvWj8YqP
Cl2RmcHUpU3glO57EJ/iUbwtZZDa7XkSoI9JBFTB4Njiqi+BCvXdfQUXONoz3y9mjC9biN0XdGXr
SN2Bm4Sk90R7ggNO6rbi6+MCU5WFSEd+iDdRG/mrdjeIVBjIEQcyp2FEdXWY9hYiyzPsZzOR0wLZ
VlV8KUfVZLSSwqj5VYL/3EcDGET/ByBqkZrAtwtbtngB0nb3pKU3P6pmse0kK3IdPcJPT3CEbuDO
dJKJ2kYNuyYhUn0qCGfDVm0Vvt1u5Xj0UW+iQ+D7fgfL7FEKcQIflVXb0iXVnoPYemMg5d0HDPwQ
Uw9S1gQM7B3bhI21/QZs+AnH7zhN0rZCMTSlS0RUJSM8wWWNfOdHJTuHGKYCEizeDwVkrjdJ5Q+p
TIRy/mSn3i7l7bsnCIlrleCp4NbnVMBAwByovxQUdPWehfLFrKeeYmQeih5vmYy2D91knQsSMRv7
JoQddza5XkMiQMi1poJs7oQjZzdsPvj1pUwqIXHcUcsz9Jm0ZOpHUJzB+Jd/aFaGNm5FZyWSlO6z
IRj6A6aXjaPsxNefAXXDB5tc2RixrfUIJECEvTnOkd/8UNxUAY8Lj4xIN5iETZT4xBZLt0PAARuy
uLkAuYZcgaqtKxbmeTj3Hw3t0lbHUHtcwM8O6VD6qZuBoE0og1f6VHeoylj4/N75qahuTDS6FHdf
kx83rnXvybR/ECyFwA7FNW3YOxXhUvi7WR+hXviFYXTWlnHbZ3UvIdv1uWIIU+8HCIN5zuELeaSx
UFZI1DuLKygaCbZNYDK6HUpp+ClskEDlEvSpvKLBK6uDJlZneHcbjLkNtxscdSdRno/7UB2EJ/Ks
OClbxZwyTC5usi2OatfkxSLZvKc0HsJaoieATOpt4TJV4F1YrNKie1hhKbq25ILfCb7cSqMH2Oxe
t1jNxJYYTcL3JS8t+TBCM9qQZkET+s8733keYWCqVKmfqLQEH+vgdEY7Le6c+Eh6HWCeWXYUAM85
mlV8eBftj89nD7wX5wjeC/35QpD5cQi34buG70IqSH6PltKPve2S72VmW/6dVnfCBRs/dCY5idfi
dY9P8KXwew6oq5NiJwU04QrZ3W+sntyReAuiA89GtPukOaNs9Q7fI4SeUA7VQdoI5LO8BGc2sHaI
gd7TVoA8vL1coW0ATwItGHqkxT7zI0hJeonHg37MVWNPKAGbb7KNgQ69M4LWZrwXud0qzmPKen6/
jLNnUxdiqGuD9uItNH1kS1iL6UMzXwP9E4wh68mzOTSb66nJVWWcKsGgQbJEcPyTSnRZUjT4x3ay
f+1YQincgtviXPbWOqBhH4+XOqoMx+6AEmQ4p2NbPH7yfsvOfvDahwkRAhOeb9Coih9KNsDTUFZv
E4SRUhLiGhi4uM7faPQRF5yY/LY7AdyQp7PhhBpVE8HBhuKEcsptZl3tNtQVIkAKbUJHxeWHOphg
vZaInS7WWAwPtrzPlH/uLL8hOXOoeGOtOzdM1xFgTXh+pQnWxr192xgzsz5zWGEi1yBGb/IxfJal
q69ahchB+K9LM+ciAg2CMfHdTX/lEC9z+rC/K3zMhqVSUsdcxDl1tVYp0AaxiVFswkzXK0rI7WVk
3kM4l8qDh9J20CVEudlJ3mlvgTTXWdcQeELH4gqC36wrNvHk+Pj/PJ8XNXbIFywVFJo07KHQiUoK
AimCiheFihBuwKcExDq980F7rQt7HFChgK+G4bpskKgCUHQB8Ds5e2EuX/Cx0kXinM2mN7GBGZAz
YCQdBXFedpzKqsQ/GawOJM9/ky25UxlXPREAgS2WDRDKqTnKr5Hb/d9+flA/uScX/WnS7m+Ljihs
cf74c9xDNzKWMAfLDTLU+2kK4H7akYLcIc2CIFVYvXP0GjDvLIv9t8m+CAv1h1nn1Suuk48VV+ct
WfqISnsmt2IerLPzbUXc3nPzggFRsSXZQiVKMl08BKEdWTcsCgs4v9eZbdm5wDpni5PpeFjinH04
vE0r4mZoTycoTtijxNq3wbugTcPXQiorw5X5Ot0AON4maaaUUFXOSxIgWQ+R9nGSheQif21epzBi
L/jRywVz0Ack6EFZhbUklWVEL0JkzAn7cfFUPkA3s4BYk6VQwP6UJCieeslxrk3zgueYQjeTT3nZ
qwiRsqkRKVJ1UDRyzU9VVeylY1HUeD1dTd12Dll9AcL2XgckwvvnzdJjz2nx7i9gUDSHawefJDSq
MMi7o5P4qgKdFsVdwT+O/QMFFtFlmvNZ5w/6LzQwbFBJMIVhHrHsYl2xAhS5eFWTQPdQ79hf6/q9
AUlgugq6jG+0C0EOAAd7UbnhtlwaiSm3ZXnPimwC9TnAtIjfJxn8oCM13nReFjuIczeliuE8soCk
In5czp5YBGYmO73dGumAhxdFcVpsuTbKYQH864XQSvPGSnFfasxsWP0zrrO0qFxEqrJgat8c9wV/
2T61X15TfO8rIFjyl/He8UIbKMojPsY+q/tS4OtQ0h9gL7v2sXpPtuRRwmH4BiydHG8Ci2lDar1X
un3AkUNxL5s3TI8J7KmT3WymBNn54WviVa2okDyPfbATWbfQlR7oYAgIIZBxcUwtQZy1WxmgdUyD
xN0XOy7QJoTFxH/La0IGSY7kcyvJNb0kuAvlc3TkV0RE5JUao5cN7eXz2ObzvV9OAbFFckVJ4w8D
6HDmbr58vwvK9Ga8aIptOUSP9GR6u/6bTRG9Ob11Qu5/q4rQG4khnpmVRPrBzLt2a1+aLL36Np+5
wNzQ6EMQQPRgvDmQLwk52mMwZU2PU2YKg7w3ivtFWVjqGalsK8fcvF2vFwv/CtBSDIbtBi5S5QmE
8nVdummRZIYrV1L+pQRAmx4W92lM6o3XHQG6v7Xm0FVjmW+XaeS0wexL+W3VfawOR1E1fLdoJ0t6
7XueBoACw8UTv/sae2JH09y8ogaNZPG5rJuXeriAuq0yvo1E4g02t+oF4XkjuRgLIyhNounsbac6
nQstyPHK/S1xjv1iCjTpfbaaHAEJX9A+sDWwDLR5aziQn/k3PgxrK0vdtPe8bVvhIggJXvHdV8l4
w72qtoYJyX5yJavzoVuXq8IZQzBi4B5Lbl2X5uef6hznt4TKxp3rEuZqu8rY/9pXuY8q7k4SUGbB
5O6uLYLtglIOoBocd7A12oCQYjbRvZiexTVJpAB04QoSBb5PbD9tLnpRe5+UOcaElszGCqcp9X8N
UDIIxLLiFGTn/yM8S+BnxDuYpeJ4slaHMkOB2MT1n5c2bgMRvQKu6Nf+f/Y2szzt7/Hn3Lqp5toM
5MBtl/I+O072JoyxJhRbSJ9ks2ZW5xa+9RdMgveDx+j2i03rb1OWRH+SUB50n0vYRid3x523ii+D
IedSFU4rlKYC+03fx78q9cA651WVupUVGM5KmLFqaI7NBI8WqjrafAW/6rJStcO6kC2w23MqMz4+
7uc5ATF534ziGdbHVmTAFpNm0PP0DDBVQHM3llEeVvBRKRxzf1GMbNI8bcd1Qor9n36IKzPx16id
bFk6KJlv4IRfjINmVaT8JQDIXwyjtVfQilptRLt3aIjF9bRstidh9x5fjvT6bJ1Rp4GImb5zG0Is
1aEyO8hU9GbEFfqhVrjhWHsmR8RK21WKz58O78xFDRS+GhxbAXNRvHbX5TL7PassG0qxL/fUwT8H
vnyM/g86KrKUc8XHbdKSEg4Y7Tnd6nnihZaK1zb6eAUY/O+bM6eQ0WrrW3gxyxIE4lp5y5ib9Zu4
57rkaZ5fB1lVwkEO0jSXs1gNgU7dgtQybGRpbLN4TPKV6vZxpajKB1VXp1riMWJghSgfiMOEERTK
IRGQXpZ1Ooe44nIxk1e8RIWwkWocBefTg3fBsqbGfnKhhMS9oNlgIcnDmyEwniyS+m9jBRCWrdwL
Y6jVuUMfHTttet6Ys6ItV6cvI20gDZ7Hr7upHmVGqMRwXMZjmAt+RXHto+qcDV7FrC4XoDxFcXDd
+LCfvRArbP26QHF2ts5WZT9WlR9I6X021xqsK2ek9MDXd73ooWSyXPIKC2b7Y7+poMxYo3CzGpPO
HpSFOygyk3U91hpOmT4STQBkPF5MCbp/MiWyTPGHodVPs7yIiWFOyk+qzqzw+mLzN2LtkcKRhzYN
ViPPBLpiNCJGlqe2LJZXuUBdbyjgGN1bHud6zv0sYNfqbbCNaBxtNvKYZGyQp9PBemsph9OC7uW2
Dso69xVwaqry9x0fNzgKUUC1tllokbbjUtAC0ssT2GRHhoT8sNe4ojPF1Itqp+O8LyI7iRe1A9nB
MFTuMYl7506cwt6OTKGQowESEhXeJdZThmj128+ReVrVM3ZBkR9raUrmRIYOda2H8A085RdfRIhk
EmDRPLmCkLwnifVpe4evzhTk+SlKQKK0+pD9Kd4Cg4DjwRkrEc+5XY+D/DkMo0d6pyEGVFneVFkv
Jfq020T1i/5d1ogKsEoDYtaizfhXo2A+Nc3+VG8BNbsfVKFT5QcHazwzGr4tb6a5Dx8YnVJSZCfM
1p3li71UOq9G6f7w2a3Jz8LYsegpz2V7+aM33mWaV1rkQ9QE5aT/nesdkRnbu3qvOT5xqLduPhv2
lnbv1EIXPWVPBYUm0gT9RWUVg76lQnDPLviq5v7hBP2l7ZRdw6ubM6gemsZ8C290ql13vCgt4DHP
Dxd+6GzlglKLoCOj3pus5C2GlgAmpHlTSOTfbQIbBT7tItCbhAt3oYmkargKhgAxpb6s8HMcbhO6
4TZ18CQ4Szi4uPFE2eeZam2dHXVvNTe/hzTNiP5htFmeHNZ1tOKLZEAPyTTbmEs/mSMV29k7Z8HI
+tBlEGXP99QuebGv5VG1yAg8EOL4HpLp6Re9JQ8vpkfZkyg5MF2m5wBkz+RwI/e7EUyY0b/7aW5K
itZDeWvMBrfrjoDCaow74Db7BiCwo3mJgxp9Samvf5CmdtznkJt5DFEUm69sZPQOf88olRHyE7bt
H8xalkrsNdoRBQIlpiMnm2PFUigLtkJEYhta2T41jXFWK/1oPerYOz1f7hTdB3Wi3k7CbK0/kxxP
vLtxX836aQ7wltfIx4VZEg2OATJcIBHYo+9a+fjtm/U7va5oIe4wRBtU5CJk3/yVPfhi/6MqWkMQ
sOi3khbRweBH73F0ymwnHV9rNTcb5utHNlzIyooG5XXfOI57F3svUxIg4H7u/TtV/tGkPJtZ1/AF
Awdue3tvC+sltZFuzLimKYp+GgqvgY5gRCsAdkPpTeLcxEoirExmfpCbRJn4z9do99V++SCygTjb
8cu+KAYvXOKSQVP0cGwzyC/vAA91OIMfT2Avuac8e1Vyj+84/ODT1fQ32yyNM7w9TAAKbhf/r58/
XmGUV5BUhNvzJ4hwnm36bJsCeADGwxSeXGGP7xfQ1mREZxXp7PNFpnYgEJXX6o0VAMjdkjf05R92
YErfYMhHEMniyYts1JycKD9QorgMw8AaN243ljHlaAvY1CVJAbYNzlD8q1EzPBr9HVG/su7m2iNu
oYHzZ3ZdQDyXEe+DWf8pEDyng5aZPm08jupD+cg2HbjFvH/ZGyl7KEydR5RNT++LJWyhEF6YTKGk
UhliHbYTigUDhUoUuQdDmF0m+1lyp6db/3+TuVBQxdaio7SxV9sbGx+llWbhSbsJFE+HlewG2WmP
VD+H82FmQksbyAmIvulJLGdTywNxmU3IxV7DCTgO8huCDKRUZFH5j4g7cvxB1MQYbhETBp4L/p8E
isXheFt5cCbSTQP8BcNi9SuLQF9uHCNL7qBlMBKH/7GeArtDfM/rJ6+4sFXpCtMcHUohdo00n7Pq
PFvMNbMPtX/13bxTsVdEbIw8LfR3GlGRjCao4eRlLbZnU4Z3pJulG1gYBQ7e99YsMApI4HNfbqRs
MUkwhL4/wJ/IEsXcN2mCgEmE01obmCSwGdqbjCGPakvHP0Mw8yI53PAn2sS7+Xz42iMfwAVm5LYh
D2+/2qDOUUKVGiJMRzzzlTwVedDqvw7ub8Tc8/c9VOJ1ObKyJPS47HGmKe3J4T59U/VezBK3Y5Cj
6LIuXzgVCBIBWm2gQUK/7/gr7SNuSWWIodkb57pJ4cK9G+qmC8n3hd9RT0g2sCjW3cTXW0cCWMpJ
RVZSg5QFNeETZXGg6zGw4iuEnSwFfo+iZadoTn5SCec4AYuf83AttTwvWhD+kE5QTD1RjYGsUgcS
9NvJfiKaaQ3fZ7v5r+20BqekzAxdn0YUeSjwnv36BDRn4Evp6HlI+r2LTh4MMXf/pNteNC4aKDGq
0RslpPPtKtdGp2P5lWihcyLXRinbfz79j08R8qt9AWMQk4WeQFmK9p70EUtVty0OUrsE8sFahVth
5FBzz0J0P7HopF+HkxPBZIBON2NiHzLz5wWg6DvEtdVhLBGYNxk6ABq2WbMb4BYXBnTnQ6a3oqE0
Dafwk67ff+c1h16YtdtjJO1m3TG7Zn/JoNGaZJJk0trBYOhba/C/9aNnmcv3Nvk8/LMmSrDYGrM+
Ek9fCQp/WyC7TgEvO0krt44wmDfmbdT2hpmQftuszUqGLW9ANsfUjFrIgCtUg1GiZZubtpa02CAp
zokDJNV+iy5TTfvf4DdbgNI/DvmyOZzcckP6HdMLwqWP6nulJq2K3b/gpgann912JykRMkPLFzdx
xxP7DpdeD+iY6kYOhAODDT5J6rlCFSb4BmMlzN16lCIxvrX6gFifR9sIZCe6ND2OSHyT55js3HPC
f2mOnkXDhYqMnp/VburUiuYloou4bCa38YCujSao0ZTShyDYiJtBIDifUgFO9b1JjbwXr0WSJ+E0
7ZUx77FaLqT9y7wF1VucG9ZGGsWoZN4s93TSbZOrunZV0X9Gdb9EKtHJq3adfblqXbUWTSYFfsVj
5MHmJL8ZwF2tXwF7VcH61e3kMCiOyCgW8a8usucmpXAVE14XPZtdEh5pWrXgkwidMYWcGhhW8Ucp
f0wSk01yu4vTAPYE/HNyPXgZ0XRN+b7GGjG0ktO4EaK6W0PxSTVAoXD0WVANq7vVjr1Y8mJ5FBJ3
nMMTJfDFwUgYip0MRfVM++vZWoZT5tMzoHZZlW/bm+dqbD84fo2HtihtGHl9u9DJ5Gz4Lh4LhNGD
jPyMNbCABhwatqRyiWxB8DTMm7+BiJ/UbNj3Rk7r4HZbVrhlNUApdMkR5ujNXYV3M95qMOjJ95fH
Yds+om7v+yZ3h1OCZIMtS20p7/Hn6Gv8HBsJ9wZKNQb1leDh9HJL4s80wW2POYjPoQt+0JXsYx7B
RiitTO91Wqw0NR38o4p3rz79DlugdH2a5J7CcaOSuHNntFhuZ2/bWpfLzAcWJZeoLVul15RONas/
ONO9u+A8/uwy3QxnJ+/gMasxNjoOuMd8jiA6K6hm2ZXPTjNPO1ypfjr1tjj/KVw4Vm2TTULQpuqt
7eQRO6gBB0cGIg7iDJ3y5DFgU69/dx9X9UFO5L0RrfJ2i0sHoGlnrMEhmU4Y9Pe6ysoH3HKjLcr9
brefmG9RTKJ64BnXd1XB4menRmHzSpXy9c/zM+Ba7TVvKHrbZVV1QIzM8pnjDpw/mYtlrSdbDlVh
VQDVoxspkI5Hn2GSZIlQNuY7YlveU6lu/HOX9Z0bReqNSrXCqceCXbD4DZRgdOfC0hj4bRyaO/U9
BvTvpplZng1vDO21c8nkW261YmIy3jn9lbvVBN7dEyI7jUPtcsEZU3Tff/2sYflOEsE+8VsCE8ua
1As7+2rnu1Qx29ozWf8qCHQ0R0S5pmU8OdAhZ0NnMnkTcJrragbovDKV3k97aKH3McVG5+kVv57T
kGQ+8jRfFVMYWYrlmbiA7ttdiB6Yh5D0lmpYom6/UmUx31v9saIObMGRKT/PTwzzGPqUrn3gv3Bn
p4XR+/H6zFtvkw/SJSTpz+QIHj1dN4ErCBUhKk5LBlHjD5PUicFEmCjQSGJtJ+rVPUXTnwhuRy2K
iC4Q2R0vDqymmkN9rxN9lLLt9tjjWAi+cG5JiAZ6mjAsai3oTSu/TfuVPE5D/31lPcCOv65SnWVN
ivkoshLX3UrLCvaS+Ybbhmd8bpJ6rqC2s1Lv5wtvocw8ibn5n59rVwC/qgWidE7ysfzqk2+EHUuW
SHByHat/yaVTp47rN2E5sBB6fLd+hWXG0WAF+Dvbw9XPoCzgA8y3rFYuIQoGgATpLDYzGHcBjvvG
edjbv9qDR/UVw8DxhkN2RFvS2Nymr3xka8m2d26puWKAHcp5b8mbMeGnkKwIlEeHIOM2iMncWvjn
8Yqp42rVqlAon5akNhwf6aol1RNipPsUenyNNIHJ1H14+sh/P1A6XuqQ/2aLnuCyHP2p5pRSnL8d
jqRU4YOGgdWpfXQEh0JRqim7ZD1VshhueVZzwD9h8QNNXa3G4R5GbEs2cv4R9MOCvWtGoqaKRuUO
5X2OeDWYgBKGdYlndQ2luassJHt/v6VD7M5fBA2piwt6ODVGwcwvJpeOYqpBvnYh19jPxPLb5a5R
KLCrsitwIPoL3YkTk00BoUavjD5nNNTFhr+nnyUPbyFvkmUro8BvN5/LZHejwp8RS/gWxj11x06T
m67kZ8Edq7mGie+OAdn8gl8Mxqy9pIku4w8N3iTUjP0hQZ7oKEt2OEufqJKfmnNWSD7PTjZDK4ZU
EKpT0BRyA8Jn1IkRoa0NDpFiAlYz2C9nuCGmipZnXatX7UJ+Sw8FnioT3lq2iXqVOsL2+OjSjJRe
xI0+Ym2YPj43WeCHPXK9HzCnXvvE+X3TzylGAArTTj+pBkzCp+iw7y8NtgfvkN4UN67TNJVf82HS
YPNCwEwifMhPUHaXFXxghHmATCLda9ojq5Pf7repa7+UFicboiaPXeqpzJXnItIRqm4zDtivp1t4
xjjs0FDpXBq7L6S8cmzUoxtib7DknSeYgahgcivT5DEptJB+xkJK+YIbM3mx1AJQYkaLAwLPxo5X
kQ9SBZlb0aiNVzOcaspTCAp5JlYdDxXjrbXP54mM3TR0kxibWYWwHcGy8Z1wIHraXmzsCg8zoP4i
3d4xJ3N3bXsHdeTvx0KCMDWZT++mJqkFjv/nDVPUySsjY+WjGBkCu5+nW5eg8ciIpd9np1RRaMm8
uw1sNjdNL6+apnWTgqZIp7TysU8LU4nQDURsTBIywZhs6zwL9GdGv7XdY2ToKT/g2IF9JUuHJpkj
3v1rDboFsw73Hw4dt4LMOX16gMhMs6W91+fb+hudok8sUK1Dutdj6OX1b3CcKh7sHL2hxA5L9Fvm
QzrXGCzdZ5wwZpSrJCcFIy+eiTFDsOsZu8d888NA1tBSryIzbNcfj2qsu3q0BbHcgJ0RjDMUIErJ
bXgPeh0JIYIMxcf+SwFjxnq4EBuj6V0C0mXAyri4jV+CxrtckvMUPCC62lHu6SwvW6jFa1xfZdne
eTC+YIxJqd02lfJ/ocG5EwBOUrRa+iJ6vz/C9cCXtuPqH0gM4I2XJ7EUaM7nY6kuSOerfjBEpn1g
4jr+JRM4xLvOtkH8CFjEJTN5kKqmMIxtVZKWYGkPrHVNZLOMxjMtIgVt236tI0KOnCydRSEbHHj9
uoWWUpqNsa50voWNvyj1sZjPYBfN11kijXUmRbDLtO00KpNPCz79SF+4FDFIUdMisYt0ycKfcTPL
JlRgHJ6C/ZRTW6UrLQuFwOdt1x5a+GcMVT6M6VDmKD0pAOVDSanq26ksql0d20Gsp1uzkHKLJGwU
BdKeMSURlC1g0IRJ2ekQ/6R8O9UJieHq2gODwXOQu5qeW9tRiJecqJtkMD3DfxNkz+6I3K5TIj3q
MnzJ3+g0s0cgXP8JGXVVtHBOfFazkUagGg0Y80RY6SKsHQdGVAEmdKngPbYhUCYS4F9Qp0opftvK
LhXdpl1edKyOFih7Xq87jqWDdjbEd9HcE2J7ZN0JsJ4GXSxwpcTRyl+Be8JnHweEPOsC+LnpEw5l
zkZVWPdt5v7Q8Z4FDELfdUxNlxlCYzYGab6jGtmrPgatCctYKbM+2e1xxt02f5BJVWn9P6slzOEo
ftTqH08JfLtGxeBnsHfgZHOOfHHdwYDgkOSGdXrKDrLH4RX6tW3WlVOoFK6PV3qHZl1Qn39bYb8C
OJPVBY/rNlK2BK/RtjuJ14WuQyXS+H+yp2Q9IZTf0dUjkQD7VbpsjfKmJtu94Q9/NOUFHhPkc/41
VN+2OzPA51kDhqcJcgLPlyS6lWfIopq7wqJBBzuO8plH5tuhQdFtbgtwl00apwXM9berRU8uTjs2
hF5yPS9wjINtI4zok7p596FoYDKUpSjaw/cn0TVhW6paApVlSHg3k4oY0legHPmr+I03PjFA8DyC
DjfTkWbmI99BTzeYfn8dJsRMWMvlgeAoqBFiMrHcXuobjZU90gW7SJ8maH6MtXa6WwjhvxHSnQ3i
zCTh2bT5JY/VYrD2xQFi9nUDTvrGfjWOm5uo/M5YE9EHPrJ8wyOvAjMNxbijiF87jzkcvHM0fbn1
Cmc6Ceg2CMGprvO+oCGQXrq4hqyjL5sTKfVAXxCv8BPSSVOJHqt7zXZGkFmOvwCN9zxdxx+3HbVC
tPfCttIK7a0Bq9gHMryVA5dYSiQ55Xtq+ldQQqg9G42lAoh6R0rZyiSnJBQzd21lDh55uWqqTV+3
WFDyX2uLQdjEp2+UYuQhVr49+rk8npmxm6H+K4BjEmT89PHF/bjrnb8BvQjI9ge+6jS8lkk5kiqR
cTlwbu2tRApiv0RBjx3VebbNeBJpcFKzmL5r29IxUv9GB/bezQl2sNcVBFMbQVeHDzKueDahR2hc
keDOcwNfO4S35Rfe4VVOhCS4O7HyP/Kijaj09zjTj2wMYv8IOW9W71HB+jtsP5WsMJoG9wT14G3H
XmgXou+cy0Y18zf218L+oeiD2d85ruepzOlUwWeGit4BQQDXSVEhpZNzF5/k2b3MBkqar9tn/nCy
B8MdvKdx99VH5wO9YtgNmzdZmdF0OpSstx7/DjbwtAXknJ0q1qTpYKnRX7q928QXRu3rQYF0a9YD
lkkcybca1L/yx4Y3rsDtyuKuwYLVgI0Wij0Pu0hrkgJlqBAROXaO21rbuFTlkoMEx15yANZcAY89
pX3F+50VZj+54qJyjAr2Ew8VaAz9Qkfxr/K+hh0tue8CZjycmCoN5IM21WuaprvpW7FHM+gmWX2G
kv+R89eI00uUKTuioW/tcOyZhXYGXSLskDKqb/yD7gX0Zm7jKDkvUcAYIjukwLzCyaHUceYEvfrh
j23lUsJeM16/gEsZtWx6b07QBsGY9+n+pyiGEA0HKtdJaDWGI1e+a/0C+wjGZNyQKgNRKe7K4Zlc
PRoLmT0dCxWYj6SmQ/op4eQtHmdWPjnItJ2b53W6WAQSj1LQ76H1o92jwejsOfCQ2riJJu7wCkAr
gER6jam/0HvEOhhmxU/vGLY+R+YWIURh/qSiRtlqEUA0OkGDZA9vSAB0K8hHHur57JZQX5RjBoSJ
dyoUqucEGyjWIdqnTfCms2dPZTZ613gN6WFN8DYEnTMU040tcJSfXhxsnl/LSdHZabJEPAzBhzV9
VvzNTe8yj8+eO2VGK52WJKnDIrSyrl527tS/nzVfUE7GV6Vk2WTfaRKi6ZzgOuMebPRGWmir3igU
tkDA1AjZQaB2LPQyQGSyOKUBDGqNAsZJd0JPNWxNxs7gqncCY4FV9sfV2NNmXpD/JX4vUP2Q2UEj
moB+pBmPxzpVXxwb2OAI7VvzH5YWWUpavAXGS6Uo57qLBa+USanInm6bFt/CgUmzF8ZqwtKSMVcg
IPk4PBgnAxOoGSpWARJOc/0ZGCQsZgzbWVjsMIta6yo5ydNbnL7dkF87UkhPa26wTxl9JwuFK5Mg
fuEkWKmM+KZDw1l0sg3J1srUlMKsz/Sz5PYmy6dJOF650F3oxUiKntH6baDpzbgxFwukrq/kPFiv
X2O13i0EYmvFN8YpXTkhEbt1XX2gObSwZSDX1roxKuAtXY01W/bPq74oNydklSGkizsiQwd0KY9F
wt7kWKAFSdmUKaf5P60PyACIAZRb/E7tiRL3chAgsIqTD/KQPcWhtf/PxBf782dVChBEu+EkD0zX
vPXBuraKbCFLMp3K6ElpSIEvivLPC+zuAPJ3wckfqss/hnoDTamyFvHL1u0B8fh0A1+SSSpaOP81
gZRQ8bAYD40hHWqsQU7nl0ClJvgxgUPoHR5TkgvY/Sx8MeprSegoxiG4+11AUJlzzq0Bh4BBL1l6
sWkZeqADkj//hby2aU9n1ayud4UXSf/smhYsQ9eBRz4xIm3VkbXIvwAQC2iXF54NblJQ7sq7XPXP
6YauhILq6qgjYMrX7U9yokjcAzUmCMv1Eo0ormE3YnNWWPgYgGig9OxgMCFGJkQY3GodCJfGcUeK
Zx7QRkbyarYJmP7EP/V7LBhRydALfMQdXphbLXgmkAO5MF6X6LAptxe7mtkbj+0sGmaMpi1I4odL
09nk3cBVy/Svhs0j6RuHyf0zBTMYEwH9vUB1Pz6hipRb54gRrfqk4bonm3EQPLQxro/AFNu10HQI
DVvIBXyg+/WT+GgSS9AMqrDjgV5w0LziGu/HP2M4Uy4o4b3pyz+u/MfNAuBbjgJWRwwIs8j59ch6
H50lvw1IbJ3mVQqfjz+Wq1SSGZT9+cu/OZxIaLuhJuHItQl5BxMgTPIVDUPOEyZkmavammfZDO6Y
H5mURrGdOp5zloXdxa82b1VSECvejZS6+z81mxPEdTDTghofzc8i69Mcw+15AFDC1o0m9GVPdqy3
yfRnKjDU3lCpmA/sSDhkYMiKpqGClOxApxluutpIxUptlLWdJzpa6MvCeXSosVJ6FG2lf4hKSIsM
Jhf3h96uTHpPoQHbCipnHeZP4bzaTZTKwAaDqjisSxoX9jdO4HUeJliAeTga8BS0eSBdJKd09Voj
nL5gPU0LfaUI8wwKLFacswWG/uGSfwGZC5fmHhr2AL8UJ0klKlHVdJPfBsV4pQzFBNxyTZBBDh8D
DnYk7vHPGM++8Jn676kKmJegVnZqUfMGjrGTwZyfJ7VvnSZLjNaImM2qMvsnx0d4iiQegc3aVyol
ApWqJ5p3hN6a20HJ4h9OPmFNOhY/m04EgiyR3nbp5Nwi8W0xLujBLfGltajPT0SWcCyy77uDknKX
Q9c0kdM4YQ3g2OAOKw0s0ue66zS+n4csON+mD+23ZbrfrhYH4ZsYLkqVkLOZBvZ3QA7hutZfMvFb
usiRvV0NRFskuRNJBz6GwzmAwUsiSTzRmlKUXzKdd4QrNw2D5map172+DV5CtAc1c8Cjb73DglWv
co3ZBddIByfQywnYYxDB9LrBptW2wBfr4E1eF96ehNMeYtgRQTi5AGbs11new+14lXG8LhcDqIpw
jzQW06EWb2VdoOpIOw/UJ228c1oqq4lCcsQRRwafWEWARA8LIJKt4PrxcwoV+k4NzOZ3+njpkwy6
6gwTbH8R4w7WAP6felnanzta0/zNoHqS2YXlioiUq+TkPTVx9HhYt95XcqU3/MKJduJ5YYd6M89x
omZH9XmdW5VF3lv668co/PlokRuGLSrsTr3MY+y53FARrPg6tBY3EfzeQ+fHJszBselgaYBVSEH0
gMsX/LAN47coU15/EeBQ2xgkohC9zubHiHbRRx6UBA+2sRbT1UuDuAdszqv1OGBFQZqRN0Wqv+71
G0SiKTVQ8h7UppGR0elP+MrU9fyKsnAC7rQnwg7zkVUk3mhlIEgBbWjBw51/J63YODPaC+sLG0qg
QV/fhhenkGqYXVKI0yUorrNjXznkC0kU6OIwq68ZewvLtXElsS2+zCo24SM2J/wZvnTwSN39vQjL
SxFPFSoDk9BRbFntsekpXyPjtz0C40GZT+uR/68t7HuK+vn2cNmlMUfBcETrjp9R3RHpNEr35A0s
zVqBBUK+YAX5jEhIzpFMDtVopcWK5rPyqTMDtH/1GJlfselO0sYnUM4ZqbNNPWyKMKZOB0yPLMaq
FwutNVP7HXqc07B8hQyOGSnf7b5oRGjasy7wQd8aRi1nU+DY5dZmKP5qEGfNFZ2HIALmHGfkznhn
6em7e7m6I7w+a4m0ZQ8KtoacXszbgE6QBHaa4jVmOsnGVL/maABgdSWjTHelR4Fxvu3xLrL1+3Hh
CO5WQGqaziYF51TnvdlGSwWoqQQa6+4+POcfubqhRHjtardxNJnz3JHzzqvAUZTedt0hakAoLNoH
s6FD7kZwj95VNWIU/wmYhj+pqt9r4vPsRLICYcebp0NjVVxHIuhWNvwy03lFDspSz+JypYfYRaIM
fJX00DzO6FIPafoFCLkY14Ion0XsBGLZuMUfWJiLCkzYoN52lHIwtJklH+5FvkULVpAeMzzLBLVp
E2wOr/ivs3Y6Wn85aPGC4HcoAWbaADYu2LwNFjTkIrsaBE+8p7g6Mow9slrncTZVkSUGMaxTkm2a
E5gKrXzzWOMPpymJChlxo2/Jrha+lrnZ8Ahow5GxhRQHsEEqVpO0BNjkIbAHQ7N4oEf5EpJBAAA5
h12MOVhVCNWqXJkigGdTs94hcYvflx8OWFJHmtm+VUIXTvbQknFBHu66fn+nyPi04eOR1Au3LgTj
540g6mB/q6kZCwHbDKEoEejTCNr6kqwROBAwJw1QC34CUTLtSdolVdf5Mu34U7EX3D+x0Le8YVML
zCcGcHNGon3AmvE4eE6nWetwA/RzmUpKNxDJ0nDFDo1QJlyomwclbs/aIOBtDzdBuMbjAJnSyigZ
YDE24t2uL4M9W2Gvf3HbH1Vcbp4u3n/HvNYz0V2IuUV9K/BjrfNlyvR4rgiDOjmH6mqyCWnLm+dw
XwXqaAVeq36LpzQwbvN6rnfUzl6TenFq1SJId5TP/BwEASnuYceLYgpfgHpuDCLGUTIY29n6zph3
q+6Xp8kyKWZdcaWh6xxi1SoHJAgKDUngh/AVYcfaYTv9UHC7Vm+Ubovb2fTA5XZKKSS5xKMHpA4K
3X7xhox+JLr/mzd6UA0lmJQLWio//dG9WRY1LlMB6E68cSsD9xIACKH2XRgeRc96eQIdA1nNlBjY
r6YeQF/LFZVyklRGYSYqgCQXXiaHnOw/nxNpZl/f2pMr9hERV9I0/MeEB75VKmjUud6cX2GSKhV0
1gQ2O9vq1ODbMXrdnikjEqI8sddQQoGNvrPUaXUGwN5QbA5XIBZ3Y/f2NxIlOaAUy0VXPV8wqz8c
LvgiuYsCL+6awbZLqJf1kwEW/z0qdSxmRXueRn29Abd2ZrmGpz5JIyopHD9U2BwA9oOGNoMvniDN
KzuEOgm1xUVkiXfm+dEZdZslslqqDX+GuJ1JOSf0Fl1ImINhJxpHjmvQExUGW2F/ZcGfAtl0/dmD
cFDVYBICv5q4clQ90uNndvBCp47tl+eGYPprQ7v6fp+qGDBbujIbnCBend/ywGsO7fby1VjIja5o
Dk8/XYWk92QekZr9EQ0vokymsEagGpizZAIkB4cEeFqKBeiF0WsDiCPXmVXDktRzQ6wnLFMg5oRJ
Q0/lkuyQcsQMsZPcOhMyr41+OtOWOK2KN/JyJMfpmRDRVES91c4mftmL7nWckp7a+WfBUvT6fM+/
/X380qAEw/doO7dyXuDbxxNMt/fUgLgR0SHNN/u6gIvHMg6GWdpbTxAJB7xJF3J9shAtyofwaYcF
j/haRN0GGKt4diNdSCotLYmWDnmLcqN5HDdiAMX/4QUifX4sYZHztSJA5V6uZcX3VBjOTDyowaSf
680Fx01HVpAvOLmnyyjwW3zE5w0NIsVB1kvpMLcLa10dFOeSzr/QYSsZKuvt4znMFZ1YqZhem9vz
ZVoRZz3AEadLJzFvCM83OOFxFwc2Kh7FG3OFF4gcoWNPzXhXSboysDL1A8F4fLxN7wBwjqd55xIp
90PZ2o/w6of94AIKCfvMIxqhxQHT0AieUPCnCm88K+LRLcak11C/eOlL7rzpauDbyyq+Sk8WIeD6
ZfwylyiUrm97n8Aiovgn708Inv8mZy3SkRgNADsfT4GXM8DBgpMKXESaOvoi8tSYyhvQ1AM6aD24
8zOa+aGluC5XcKKqA0edcsO22l96+EIWMRU3R7RG+9CZraH7St70w6H0USyMAd6DYkcbVBM2FapI
8R19GfPtwvcJvycSskw5nQ72uQIPkP/Jf6tCrAMmEHndAbxLjxZQeD73KpopqXrHAizBw3rIkuh7
wjYu066NsRtq5BnFo1k7EkWHtEGiQK67uGtcxK1vj2nCCMP8TOaj/t0tNzvhXKN5O2/zGN5GqGgN
ImXMU00ARaOdcJyF4LNyO/xAwEKr2kZ/wz9k1DHZHF9FPfYp43mpzjFbk+oXRelDeABdSK3cAixO
uVOrzd4ipp1HikNw4rCajK+zvvRy3Qtx37UvdjgPs4gRdo9zlRwB/2xUKiWMJ6t3nMP3+vPiCVL5
v67000AStL1BTOxGzpqODXCX3JyCMgLjkHLJ8Xm1GGsKqYMZgPBhUGtoWzQR0dg5jPgsqXRTejc6
+UQS2f4HaBMDfiufyOBHVH70ZsRDqj2Uc3lWt1256FpUgoNq+oB7PPdeZvqxkUMgtb8VYYLcCg+f
OZ797Q8F3OxX7SHjmYq5w9743y29V+/wVY5TxUS4/MT1Loq1JZInaFYpB3xoJuBVSy10Mc+D/Znj
PhY+N5nsXpyOWT47CTlMlvtL0AjF0e3+26wsIUnXtK1+7y2nXtVWhTULWz8eH1JEytTKdZsgrbbb
yAIvm6izy1sMl0nkuHxD350EKsmk9OoYsJ/lpcP3W6tbsis34FHxoeN/MwA7SQilsW2hxd/8Wgzv
tjtbuotBhbYAQMYj0lMKRcL06Xnly+lSOvfjxkc9EoWbeIyqcOYqgDBVX+8LtUue/Xgh+vkkLa7u
S/3jzj4dlY1+SiO/9pFhZg15MUXX7YfBFZC0DxL+hSFRaFT0gys+AZdROqwnOixTavuvKY4NzrLz
lxsHxDEw3ITNG4hK7PfXUib213MwpjrKdPfOqv9v247gW8i8e230HDpyU+HDHd9qs8H2MXqB74bj
Js2jvWG08SmHksN5UR5qLotckxVAuuPlMCphFqaixEzFuqedb3ECxZkFrp/0JcmA5ReRM1H3l8Q6
soaB2R1V8askAZukqLdWQgkKyhdW9NuQyPEKHEHMpjt+fsPMpVL5CSd05GJhIUJ4ZiH7ra9EjasN
PxG8oUaV/yKEy5+TTY0lUuO6tLG83WRmNdcQz+p4vXya6udLvjzOCXfAkqB9rDidHxpvZvbPykK6
jLqDrnvSvpPf831BaQAQxoZW0N04VWYalpgUxoKLwYXqWoxS0KBy0hqmgqfaf08y/lOIX+U6Bcn3
NGLlzpmeWQX3JqMGNRIhJVWpPpxkFGy2bIcAlTMoYM+0f+jqrAQqGEN/uu7D02tFBYDjW/77zaTU
J2KaPKCksOMCwFyguMhVwYCj+/FBnYxqbCOEH6ueMEt7dZHa9J2UtVkhytYFndHiA6dItlm2xdNJ
jeX8v45WsbHW8RIatoAvvrDySiWFg1UwEiIUL0T9Vc+gwJnutGWCbwyODop47Zd+lVRJG0xqMxKr
PfJtd4HkhOL9VY8XAYM/Nwi9zJ8S+MJhX83Jv/6jUC/5DwTCUxix1z++VWOVanL1Gkgpa6cCUBfL
I2GDDrYJa/iadAJ6gNzOiMhN7GsRYswX5wq7FpHQ8iq0truUYPFoyoGMW1FhSIVBZQkOGlpt1Opi
kHv/AOD/dWpd+iBgT12/Z4BMUTRh6fd38TR7+lZrQp3+VJreWEVJ3wLoWBAcfzI86YLa0JlCmj4d
WtAn95DTMguli7cFzDvIsHO3moRO2oAAVFiV3O4hA9qccAezOrsPMY4gORanbPu6CshwIGfhA5Rc
GvXB5gY4VusI3o0UAda1DS3QFUtkgEuk5jQ6ddM1PSDbqrdUTg7tBrecrhQ/5ze2wsj0FLnDdyUj
oo7UpNEvvwJ/2N2TidweiRPQ79uK3dCTGncUuTK4MMSiVq+NxWhROXzZOn48YnDe7Ww5T/UOImAL
d6r8M8V1VRlaHTlxk7WjA+orUi8dQqVpNEJVKT6B+9xSiGHYXv4NjsAYxRtPoEoSpKcoIXy324Ig
KW8CTaN89bWLNanypqUK7++hMPVZgN6jysZN3uBRODZRCdhtRytSXUMYVKNfjZ4Enik+X6BkPZIj
k2jd53FMCLFV9Mcat3xqpRaok2HbW4YBs3/k/3LnnOub62MuvwLRtSDX2ILqaQ9iLCkB0TW+u4ca
J2uha0yxBft7AASjNYuHzjZc4EtlopjwqFcQo4a2qJ9qm0sa2a+1x7+f+4Zd3RYEmBr9qvCeStaN
XlBHDIUgnmWwLQUWZXPHcMnd68DzFgdLYhw999AYgbsEseZxKZiNLYHl6jvZZwRnEeZyNiawLPAl
4T2y59Ebmr5gtUdTWlsDt60x+G3wxmBFFVGq9K3Y75yEl+OntpR3ucX+8sr277WJlNBSVECcbKev
ghx1kQaRvoMXZ6e8AIgcLzGLE4CTO2x6DVvABRPeT/WWMja5XIcDdhQovAwwVkBnEx5RPoILbzIy
yJM5HLM7NR7Pk27pSH5hODjuNFuOb/JzKWOK+ni76avzoaO0Auw6Y2ONhv3eyKFUrAKSBCcqAtqY
zEINpx6LbvAv/XMmYqFWBgyHXNo2Sd14EMy33SLsQ22tMWxDfdk3D2VeryVGrQe7tO0+/KOhJWam
B+vaU8xKZHoUn6OHBaG6b3LR3fIbnMk99FgIrQp5dosR6YfGub/wnzKhMGqkuJmmmcFUEq9PgLkg
rBt5sIB+y4eBWsrP2EYNzuOHLGoSVXkGnXpflW1tCOk7BtcZZ+tautkYYn6SBidY6FQcdh/rRIri
ssviLG99CbgKCyQStOrxGtLU4vyiXQqzHoxJQlh1HF40qNmzAdfVB+dMcVJy/sw8HaBdqP5Cnmy8
+8U/DDBVtdzRfsYX4wAycgV6Pz93ytQqXCI2VdrMXHkPVH2xJEEOptpYG1LTYucx6+/yOHetslvD
B9C906prUVaO3zqHMRrTNuV2Bnw26EqPrkOOMz8mbTdQVshK9HZGOpT8F8al6IQonZxSgknKyIbu
FaPyPs8aDVairrWaUOyjRyTFUlvBEWqS6JGs2UmaQPJrItbcJXYn2mv2xZL51qQPkXrWZgwb5ujO
NToYG3NZK+p90HxSe+GdrDcQwhH87flm726LA8UY7G/LAo7eq3ZvbuXuAQ+8OBRjcakojX/ic8mp
eAw7R/WIA9DKVRl7iWIPhiUd0MUX3ij/E27FYzk2uYSDRoesNuACv4b8WXtGnSB4Os8X6x7Sic9+
lagDKuEDP9geWob8hr05SPcTpACWY7fEZ8Csp46ZHhQ/lurKOrfc4JZo2QANJxAsKA5vbKv9NqYh
7rUjujCyh3E2QgPNffUaQ5uIHJfgR7/5yYxLM6T91WFxsoaXKZ4DkWBS0jgp0iMaVspz0C/EyXLc
MyoPWtgAN+UqPpOguuwYiIuOB1iSmelrtNL5Js6KG1p6QMyyJLpGD5ZNeqVvci+q1XloFRSR2qGE
WjhEawIKXbg/9tDR2CDupYRUrOlAaaSg9WrO5PopmEVqPDm5At0hgcsljE+n3oATdDllRJwiLDh/
8KyVPnSykguPwZRnYjY3TPSd/0yy0KnRm7ya/m1aXjW4F1xJSFHNbivXXtrTUO5rvtrag+xE8dcc
/ZDqsql/CY8UjQLOsiCP3wRAfPSvAFuVBmu0VyRG9xtxfJLNBhBJWSjPbO7DY+SGsdttnTeytvdM
Z+o/Yyq5oBoHChWIU5xIg9PVq5v/RB6gB6VOEpQyZ+vEx83UNhdt1Sb4wea80Ygfs+l2moaqAbGe
MjQDwggcJwZdT9TmHmntcWl0NH13ULBG2oCV/06NwY3VqFzt8ITEOorz5oka7OivkY1rsIAt9Yih
EYUmdXmYMTU3fIumc8WSmIz8acQh/2Apfz3+Nws0Dmd5gnWdDTAcGdWgP0Dt7A2nJCY4LJ8iqSpN
THb44lSuSh+QDje1kXGEPpTqpskfM8cHG1J0dUa1EBcJvL907H9luVO1Lz58kZ1MWR3NL1eLaasy
K4qHVZ45rkkzGAqG1yuSavl9BxRZWkz5Y19PY9btWRRZBUzRskmJPXl2wPK4mssyGNnkXlW7f+VA
W+ku7ZqPkQ0Uf6BTEjDqImE+XhwZ/ZSSNBToURoarInaAgFmTFVA5B2KYfVGd2Sod7qNYIxVYsCJ
qLL9TWiaWn8cscrivOFbZ4sfPeqHgDR/ptNRmH+eqHg1PGBtO1PyiMU16TTX968BOe+iAHtILSz+
mJEjh5XdxRheDLKrJ9GmSmVOls9IgHnXKUZFE/hA0odFw4E8IyPA0h39HNzJnqRQoTmuJyUjYz/7
+VnC+6L4I7tez4YNcENsn8aABz5YPdr05H3FrCAPcZt+Ug4knoTcu42KOaVECK7ieBvPqUDZxSQ/
Kdpl7yFBwc/ZVRaltrPP5sdr6ExulwbFHS3GGocrQdYbZoQxE8tJC1bB7aYCp5LwPR8EMIhzmn+N
ulDfrHTRBcDgLgv2zMUuzlxvTPViU3wXITQj9q6BSJk88FvM+sSlhRhZxgM140j1ZPqdgENwdQ0O
vSYiU9bFoTacT424WUu3AGGDekFK0vg3IIIGoLh6b4SRI10Zx1pjlwZk0Wroq9S8caQqvxyLWfj4
VcQVrcNIdgivGlSlW/o471Dt0T7M2kGMRVoce3t8o+FYcw03YlZI6/u1bslpbzxFvHPG2nX5ftMU
SgujRiRfSfGFzycLjeKrRmINr5gBqMGgO31o3gQMKX6iSD+B7Xlo6yZmf6MOU2mLc1646amWEEC8
paTwBlQ+l1R66VcnRKBmRJZjW+sogzr1Nz5eNJf5Mdpk0RBfhsor5BP1h1sOcM6uS1qPyzFUSAlD
WPCVPMDVT1OwqkdUImpvkni7fpXd8TbTEy3TyzejylEDW9Eoo2sJjRkBR+jug8RnJdYuG34Gc2N0
lKgErcQMxPanvgAVfHENfxVO9WEFoPZUxH/ETeA+0yy6ANzVCmKHbyrlvEnsMkjM86KA9AhM6I5c
lel+gCuxOvetFZVOsSlDAgxk+cI2lXq9eH80rEe+PJKdDg6ku5dI1PmlDoLfqNkmmjJQ06zfAtu2
0hdF8uN7GInoGbEzWop7lauMSBE2qwdp+u6Lgal/h3dIdPiSNgHGoXHK0u5DDn29+Bwjpj6ap5/v
w+uZelJUVWXnoXBnr3ZQFJFkkP3z57Rv7XWuqubaNoSPX+BAhCsFp+Zc1B5m9a3+LtM6l8PT4ugg
6P24yrGEOqOWn9vm0IeZoBE5y/xSN1wSRICyNL7uXiZr+fOahhC1LIPCeEr+JYPTlQy4xuj7dQHd
RZm9W+U5q63+yu0k7ukH/i8BLYMEbVnmS0lUgyyF3duxFFp6SZbr6Ymu65bS2hdhdPneNNlVN6rM
DFShL67IJ3YrAbRrzSvmeGsG43eLMI1iwituEYWr+RWKAD9gRjqlE7/m116JuRGqPt/5AWd/VqkO
5sejE2HXZCCMcQSk03uHMJOLzhmDpmgOPY8qWB5iP1e3ccEnO2yn5MrutoGMvd3ur0CgCPEcjcqM
jzSww0jFQbbmJOAGMc3jKjNCcP4hak8HOeFjOtdqAE/Hy7uy2THBOoxzHL6PX1Fh04IDRrNKV8m8
DEgplej8W0diX+jwmm2HrZVD8ldl0kzrIsBHMgOHK5NFKuiXDJl48OFfOEv37FDmOtKwc+EN0P+U
SKyMXv3U43yU1XEgnM/h8bNYFzEcxuLPd8WkcOqQnbVNCsRtiTTH8bEvdkCGVGkpa2kmF+PuFgHN
to3Xw8z6IrzEQfAY3Fha1pS6kHoKAeeeB8h/HT6yg6f2lyMHzY6Jbbj2og4VJV6nJ9qKmS0yJnBK
R14ncum2dcGkV15IfmejnLIBZzdcbLyt2Hq0yCwmuMM/r5b7h360Y0H49FfiNY+gZEBKy0j4rC/I
/FAhe+7TlvuNe84PXfXp3qyMYSzWREvCBsjk+gfczmIi7hmT6U4/wdCW2sL1lDTFtpnm6xYyAsa3
PIa4RK1IH5G4oN0YrC7pa5NJyBKzA4lcgoBsYHh3jJyn7xmxcGQeDQODej3qC6SC6Ga+6M/Kfrpb
ckEHX36EEWyNS61ArZOhjhpNiQRRniAgteV+eXxRglr3YZxyOjLXu8P253Mc6Y5Bzw1WDWReGBzZ
MzwOvhKBX+BJEvnWccvoQq9DJBgA3mWoNDNx75/H3mwH2Pf4Ltl1b10lmrUY88bpT9Ahk9evWfmS
5C/2Z/7x6GImgCszAn3ZEMqLYLd7Vr8Hc8yw2inpGu7DXKbsB0S8IzN8f1ahfNpdqAufkLrLkeJh
zG9bFSVcoJKlZD7uJj+2HUs9YSdfGxp7TuEI8BSBtqHEMgPDAQ7raOGEabHqQBMwdWI+RoEwtWcs
/BMCeXfE+gJ07PvJFPmiOm9emE43Cv3ZXX8nwSHobD4Od29uce3q1dc41WDE/B0s4r48ObvLZjVg
h4YdXwMzBXAbVziCbkOtpmkvV2PSmw85LE1ntUUrtLxOT23TCQV3GVU/vOHB1DpqX33bznV4I/28
FISZHvXXA4VQCbG8BjYNDpxmsmjH12eVh+5Yvi9lxKvkOT+RbdXJimH+3F7VYr6PKU/7Wvu++9LI
ZLUBFK5blKJ6vm/6btkujXpTPUI+Qc/o6wrmtN2waPTR9ioeKijSlTBo+Pc4Qxi78YMML7UmX76p
j1Os0ewwnvgpEQaZLH8SbnXdBMtePLrUQDYPhVVFjsgvxRgg4OXImWI5MTap8MDqf3U3Ta+pC2Xq
bmJ7GU72jfS67nZVW2GJG77euXyrQstkrnD+vA3PWRnRZYafqsQNiy8lxyaKQXTtPGVWOr0zDj6g
iiGCO5fiQCpuFhp6kB/0oYaY4ffbAVE4JAvcqWm6FO32MYD+EieW/VRsYEs5QFDS2EbOJZBKrtH2
k2JzOpMZt6GcuYpr+UphDHiC4ZaOIurQp1v/qNLxRVVz/O+IULo4eDDnmrPlBJCN4U2+GT7ceg+G
ceNJ/cFKsDjBrlV9LNOdepDoP9GWlVJ+66jjLSxue5j54lPSs6qfDYCgyfe7snCP7L23d2lMj5E1
IesKnUtR0RaLZNx9iKNcNzewTfvbVguErnF+RMHvPRy6Zy4SyUihmUQdIjWO9+oOGtAu/ALCvpSi
1wdbxHamLRY+kkjxAQ2STALaniMKHxaFA/vPL9vlw/jHPJl37IRjQayDIEGZrDqraez/PkmGydVf
AvBIcZergKVegz1kfjSvaZMclwbBnykRrjZCC3Plngbv453rO9ihJ5oBE7DQZDtSSQ5Vtwk2OBoY
/C+ugdqdy4Zc5snC5q90BJngypFjknwL8+Y/GEhC2Zsr7h5ipGX9IXZcCejMG+z4MuKRdRaQ3ZdX
sJ5DDKG7nQE9IALi4y2fGyctrwfhcCxVLzlAGlfXxCZjpYban8qEeH+JFmtmr8MUFu4Wos5AJ5AV
PcXbmmkjGv6cG8N3hdnLWlGLWmHRtVVa8PJDqkvgnRnBZgNBU6YiByKX2MepZWZNCwmU6ieFuopv
sqNTq/VIO10CnWtnCjbI8U/2Kh67QzKG/96PQogDxsjgomrAyqDu49IFbrD03zGxMO1/F+scrvFO
UhhV9nuqN7p/B3skTq40edFoKx2hbo8POhlPf5g2ctm1J6mZNHffUUfTUR/e8nvNWyrENtycjEf+
XLDeTWxVlV4TzedTztenLwe4a4p1OfAdv6RQh5SaXfv+SNw4wzGYyXV64cPfA+9dDDp5iMQ1BDJT
BZtuwAle26003xCHjhrJZxflqgltQACY6O0s8Ldwhq6uiJ3yaUEG+XiOkeqPkgylmpA08cxh9iQW
BnT3+kK3t9EDOlZopB6KXstWOMz7y/nuzwEmejLmi2nRlTVItuaGRqQwla3fpAlCh1cFJsPrVDjh
3/rXlyDSppEdybhijgytgx2q1+BG7dUqwnacUpNmHMwyahx4udz9O6XeolLKsjJFx3qlYBY6Mq8V
YMn1ka2JrZfPOwQwC+CE9B24tr/5Ryx4hCfyoCatcmyfW6ViyIWk
`protect end_protected
