��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$Rx�y�<��wA�*;�x���@�̦�W�X�fa�M-$u����n~�%���P�$��W��kYَ���P7�?UMfT��q�6�U��k�>����~�\N�(�����X�e���/6U|)�X2pF�]$h���d.���9E�	�IN�f"�\��e�z�y�b�����Oo2�?�qˁ'�͜k-�K�P|����y:����3�l�d���bl��ˢ_�d���kx�rq�mh�MذM�`aS�.�DW�mS�9���Y��+�>��!��!�T�uOB���,��\L�7m�O��W���6����'���j)n_�I����2:��$�K�2�Sʫ��l ��!���{�l����.�j4�	��很�̢=�����N��s���s5���_�R�>����ТP .W;������	�"�מԫ�����]�#7@O+?�⡾�Ԫ���e�O�\A�	�ͼ���ƹ�d�	@�nQ˰��E؁Bf���|D_�%au�-�'���w�*%��"AM$w�*Vy���-?aU�׊�4��L4 K�W�jNd�P�D>��R�қ�r�a�����K�,9�ZCa��MG��~��¾f+'�(��R�Q�IYm�A��������>!2m�B�נZ��&a��V��e�u��T�ǶM�*���J\��m�\��D���-y�R#�}KJ��2��եb��X����
��G�|cd�q��B��#��sj�cj->�����B�}_бz�C���t��161�Yf�i������������l
L��������Le��3�;d��*��M����ZKH]�xV�[�R:����C�?�'�G���@=I �=��goY�0w������5�Y��3���Z"��3�,���ßhFtZ��e��>)@�Nc��w��bK��--
���ͥ�R�y89�V^���!MNHH����"�y�� p�$k��|�	�iV�@� ���چ��I�~��u�
�e;��(��K�F�}�b���x�����a�@� �.0ͩ e���{>�҅�|��ʘ4�[t�]��&��m9}���-"�5x���Bp�(�\h�s�87tN���(�e�4�(@W~����אo .W]5�:+P)�0ʠ�9]r
?�VX����fdr�@���8��VwM�mK뼠>w����R%��W�Xy�>z{'iP�*�YlN�˛���b􆹈y������B�mޖR�8�\�+8����e�`�����D=�'���-'��u |������d���a�Dg�FiN6ƈ#���k��KQ�ζ�m��ph�����1���2���w��� .��x��\�l֘����G���P�H-c��G*Io��f���/|+�4��(��_�u�7��$�scW٣!ʵ��p�AL"�����.�S|b�z���I�3G}�\�QA�6�cl���Q���DfV�T��(,фM�Ƣv}wmmR��Y.-�_��"e�����~�a���l�z��x�jGb�B�up��U���A���Q��Ծ���0P�46��S ;�Ƃ����]�!�H�D7����ɕ�Δ��fFP%�2΢��)娚� e1�o�E�vAʍMl+��3�h�;�w}��6��_��څ�lg�P���w|VQRI�C�/��};��s)1��m|̓ )G�b�ƲB�>�}�AQ�V՝񈙙��|ldQ'E/���%M�����P�>:mS�$�ޛ7��Jy�B�, ��ކ2�/JUщ�>�n���@�騊8Z�DŴH�Չ���]�Ͳ��3'������s�`yL)*���祤�{�~��B�97��셪�O��X���*��0ښ���Yl'm��i�g�nP�]F��?L��*H��򰥁阀�ٓ�{��9����l������+�E{��(��|d@��|���4�R��w���I��k9�j?��O�l���k�XYS)��V|ԏ1ȣy̓�ri�m�~r�C���aV2�{l� L}b�](��q���O�ڇ�Ԣ��KBʺ��0�7g�M�cͻۍۥFBHp+��s�.��C�����:�sZ�k��%�_�*�$�K$��&0mUJx��7A�}78hq��w�Gq�����W],��Ą�z��<N��
��y�0k�z"�r��R�%D�|?$(�Q����ܱ&s�6�[�A�u�ڞ(���@oW��<Е�еˢB+M�ʿ[�|d%���7V%����m<��y��CN�4����6o^u�F� Tp �XJ�A�y��GW��<��5����	ǹ!�e�?3Q�0�/�b�Zʗ���[��ݳ5��KY,���k�⒎Կσ���Vm�1p��dȕ��MQA��UL�|�V�J>����[�zD��YF���,���&J���	����O�Y�־��_���U�8��������
������)��k�����$�a���B�
G��j��XD��&7#ݡ��!o{4X���M�i��6$f�[ 3��F$�N���`0 �������B'��L�}�Gs�ga{%�����q�'�d��oK�a$8�ox�A���	ׯz!�p���:՟��j>X{&�Ո���ū���·�_�Cc��.��M���lL��䋖K��Pyw���X�P�a��,̉U��(�ft�ك�i��8bE�� O-LW�P��+2Q�?Mv�{�H�a"�\��>me�OL����"ݲ�t�ېn�����L]R�k����A�`0�I'��¼R�1O?L��z���<t&r���Jٍ��ZX>�����g��������$�[����{<�{�ΜS���뮟��3IAs�q��|����U>O��N�sr�2���q7j+�1;.�v<�T2��'��b��� Y<��=aS�a���H!�&oR~����sT%>e�?,Ų�J�nO�U���B�Y|���3������,�;WA����VKB��F��y��ך���&��o6�Rƥn?|u�<�=�b��TOr�4�����(�J���{���o�[Qv�&>3��򛽽&rY��8��1D}x�ft\Kx&�@�1QD �����Mp5|����Oen����?����A%����mo��؈��X�)�k�	���qfT�w6�����1G���zRs�]�d\���㏿�flt��\P��e����#����;Cgm�cL�n��Ҥ��?w�D��"������3mp~+)ٚr�����Ya9������[�@Sl� � {%�c���rC�Q+����y���*J�M8�B	4�vʶS65���C���"9�8[I ����:j�K���l���./��)!��~�g��W:��T�ٟ�}#Ⴙ���ȉ-9F���t����m/}��=pA�����C��*� [P٭)~)f���/y?L��mq) 	j��Fd��ԅ�ZX�������kø�C���^�Wu�y<�/�ҶS;R��:�Jso�mQ�D�.|7ez����N�� $�=g+	��I޸�%���QU�zzf~�z~hL�����2f(y�װ�����u�D��Guk}�_z�����s��ݜ��2<1�P����	75�ѧh��*�k���Œ�f��L�iL����H��H!��.�	� ���HDI�e�R�8�H��\�����c܋d�t�=l��4�qƖ�w��P�p��S�h�����A��; #�ku����O��|��V�B������ˢ�tjA����F���'�וT��C#���(�gGѧyXX����B_��_ę_�m��}��J#J�!���#��X��z<�.xc�_$�a{�U�I�D�5��"��[>�����@PIl7Y���_̳�M�m3�w�w�7�З�s�ޒ�d0(n*	����hz�	S�#�ǿ�D� ��п��U>٣O(ύ�ր�����}��Al!�Q�?���0�}��_�z���Up��4�x:���.��*{��c��ܫ���s����X��g��\Q 4�],ʼĬ�~��c���^�/A���6�^��4<[|��/��6UG��I����K��L�V+2�02*�J�4pl��[��v�5��� �^n?�F&����� /�U�4�j����:�����6Q%{?p�75ε�����Y�9����3�'�S&�����xO9���/�N��e4�0���ND��"A�4d ���;%��
�p��$5�R��b�wq�:��+�~���#!e�h�i�vz�7&��<��S7���;��P�-2w�$PX�T��ƓrSW��&,C��@9�n=Y}�&�^�%�X���Ԅ0�$���mE�߮���[�c+����ң�
��4��0��?B�@4�YtZDk�yd蓼g�Z�Q�^�z��MV� �^\O$U���债�`J���_{�S�nA�T�G*;Iz�vCͽ`�S�o���\�X9�J��Й:�;i��R!o>�˽mt9 ���J*�f��%�t���k@�֯;z��w$���fz���4l�d8�M��[��>���DtR@}[>
gd#�{EL��Ң�O q��g�a���ܒEP.hq��V���UKL��X�~��Q�v���4���;v�}�+��%�#D6)nX�}�&R��(��1]�H7.�օ3��Ul?�e�A����Ŕ0���_0�5�#
��ï�Ĭ��,D�?�$�zVu�=�`j:.h��� 0�SKmJ �	%ϫ�Ͳ�!�(���ZhYw�,Fe�x6%f4b,�RÑҧ�l~�F�2v3�L�ES�ka��<k���p��-6� �.
&��"ѓ�R��EV���F(�)sq�]�.sI�r@~��V5���W?��C���Ƿ]�D���6G�_M�����j.yM��84Љ�%�Ou�C����fc�ײ�:_��<�)����h"y�����YT�a�Ȳ��a�&a8�S�pNX)Ug$�ž��O�As��31}4�X �J��"������g�k?`��=Љy��G��I�ȸa�Aa1j3k���q_���ǖ��DFo�c�����>d���R��e�q�-$��r�T𻀊�)B`�G�q0Ue09�<`�{�6i�ޘfL�QP@m61 m{�x��,{yqQ��zdjV>eQw��m����n�)IZ��
y��'�>� ��q�wѺ�I�b��%�{3�'�vx�xB� j0Dr��>�^��d)�����_ٲ��`eM=�L�̧7����u~m�;����z�[�V]`q%�Ha3�d�T�N�3�^d�k���J8��'@��K���!Sy���K$Vq���	z�<{7N����>���&�:���O��ָ�J�P�nx��=p6N���L��$�tn����4�Y�]�˻<Bن�bq�,��Qr��3=ҎKj.�em]Ry|]A��=�g�0H����y�m� �v7�|�M#81��7Ʈu�nH:�A=w��7:M6&����>��x�n7��S�J��4�8�%��~n����Wu�6n���/�MEDX��ӿ��~�L��-p�"������0�f�o9��pM"��vǀ)En��V�+�̙\�2����A��+�E6�*nE����!��L���
=Lt`|7����oI࢛J�bM�Z%���Ě����E�IP��K���ds� �ݹ!�j��s��\�;-ѵ�즦��+q��cf�`e�ĉ���T㥦�мg�^��0c����c�p��*e�p�0aK��6&Ӓ&�L1ow���]��NE
��4#�1��ZMY!@NZk��0(L�dJO�0f��8g��3�IoC�7�_����c�Z�P�@_�ޘ%kp�(gw�����]�?~�l�[��{a���3N��u@�F��8lN�V� �r[˂89�D�4����~�jx!�NƛbA����	iS�7*g���W4�
3C����|�Zŀ=- �y�C�PJ��ؖNr��PI�w\=*i���.˄7OQF	� �}I��u'�`yC�G�>�:�+& =�����ٝdI����s;;M's@�[J�<����|ao�Q5�� \ �Ű��+�)Քa2^4��^Y�?�.l��@��w���-��QC�y��]̦Q�l��REÏ��=�-oT�wn����� �!�X�<�N@AY��_ }Ρѓd�$���(	}M��M	��c�}�{I_c��8x����x�\P�[�E����P���������n�G*`;1]/"�J	O#�Mm@ g�=�Ӷ�YRyx�-�rh�
O6Ʊ�I,�C�XXD��qd%K��޺���6
��]�Q��ήdQ��?\3)��4����R��R��h(~��OR���0>��ޓ���'�|�˔yr�{�P����?�ub�8�0'.m��s?k ��ǔ-6.���s���}��HM�G��z�,C�I���%w,�M�jy�����l�w���1�c�rݬל�.���Ǡ�?#�M�'��,�G�	Ĺ�k������L%e�!��?�*��`���@��$Nn����{�,��{��敿�Q�jK�G�K������`޹b�2�2�O��J��Eh�~e�AX[{�'�	�K��+��(�2~4օ�����h�7h�e��$�A}L�+�7���6�5�{�	��ԧ��	i�࿍D&/gS�#?@VF�Mh�;O��l[�I��R3\ؼ�P�k�fS�D�gZi�)�D�4��A�ٺ�' /%��$?��u�>����@�5�e�M�+� ���E����[V"�6�4��FEA�8�1�;��_2�L�X���]���[}�h�|V�o�q_���\g7�b0RA��́������$/J�1ߨ�1ɏ���if*Yiʮ�O_�w5��z�l�Ͼ���*_�^ �Tqd�Ǯ#���>�=�em�����$�7��/����WHn-�F�uR8��t}�k������%�뙤��C%O~�����H��Z��ALN��s�GEn�/"&Zf��t�)HaS3,���u[.�g�������G�#��3��;�+)���Z{��%Hl�R4��1&t7�WP7F�.�wx�9?���h��y9D1�z!��^�����=�ڶ_a���*��(*�?��d$<���Qa�y��&�{PH. ��6��"w]lK�WLS/�~�ҟg�D֠��N�g٥�22��h�����u�%"˰��R�0V�o9>C�2��^{<CkȬ���ߠ`[�7��CYT�h�u��T���8f���	�-��b*?&[R�����4�;��x_/�����x�l�劶������W��m�Qs�ɐ��`�eT"V�"!�i�ࣾ����BoX�N�Y+�u�:�M�,\(��\F)������9�ʿ��.�Q"�);� WF*�.��n�ũ����4\��ğ;����[zl�Ġ��/�Ѱj���(�8[�jr�m�	)$�5��0�٬lE����T��\|"fzQL�|�8�IW�:Bę��jb��5���Wq`��
�+��O��៚z2��;k�|��>�~��<a�\K����p������-��0ܐ�'��҅ړ1��=AA�9�
R��j��)bd���yh�G!���dL�\�Ӫ3�`湀���'���#�vq�jO�`����|T�6al:#?#��j:��.�	����CR(x��eRMߞ0�0�����(N���9�]B|uC}���EhChm���I�OSޣl�T9�5H�]+i��`1�����
ba�}���(��&���?9��gP�
��v�D)�wj�@?Z�7?��#3r�G}eL�����6����%4��1�)�,�yG�=�'����'�[�����_hw�Z���m�:V莍fc���1�4�5�j��������P$}�^��$-3iܓ�k>X"�a/���*9�7N^��'�ԏL����L}�r�n�8I9��&���9�3�z%��3�!��Nz0A<,��+k�t��-�(��M��n,DH�8��j�>�*;�@�밓cg����}<I���� ��X�$z�G�#����ݺ��&U��k_t+�1Π����SF��J�>�@j7��'ԗHV��k0P$b��M5�ng���PG�V*��p�x�����9�1�NNmַ�4�`���-�`� TU�K0��ϻ��-޾�Dcp��/��� ={Z*���z���4ܔ��\#��š����h���3ߕ=�~c���>qsBw��J�����^m7Y91�Z�jz���� |����,�NCi�_I����twĩ�G���W�T��){��`�Ȣr�BO����V �<�	��o�D
k�>2m�{�l�W�a��޾��`�C��������t?A�fTb}M�κ���T�_�zޔ?1��x��M����N"�AE��g8�� )�8!oy �476�2:�&��;������d!CJ����i�,��]�3 Kn�c	����؏mYx��3�"�-sƮ�$����P�p��HF�p2g��8�.R
���l���V2�/�T�z]�:F��2�O�Y�F����aES֖l�C�v�����E����*{`B�/�����@ǈug����96��'3'6���?�ot�:m�8�z�g|:?m��������	Ot�:4�Σ�DȤ���b0j�B\���BDy���(L��b��-��c�`�#pǩ,8��Bht�]Q�C�+�x�w���N,�����Y(�=5�e��XVZ��(_Y>�cK�J�39vy2���}���W!SW$h-墅M¼��x$|N�t�&���n�Nj�-�b��^��~�rm�	�8��N�hR׾��Ô�
���̏��"�?���0A18��Ơ���\�Ot!��D�R�c>�3�Ϻn��_��� ;�	]F��8*.y��������<yi���5��������@gѱ����W[�8�iB�/\�Ì���s�nԋ�}��l�����i�N�EH&,>6���HOg��SsC��N���V�Rh�N=��}�O�I�ǚ廿~å>-\Ne	'��Ūq�W��|��"<�&�ۑ '$�����x
�'/qsTZ��r3�
� �+�L�W^��-�vRы�[]P	�[�9;0Z��r<į�pԚ��B��s]�/v�\��ک�ex\���$���ǭy��z/gO��a�KJ�8Y�����4����ǦCq�z�$j��6	h�ֲ�kj|�w��y�ĸ�l����=3��N��h9ƣ��*��ot�f�t{��o�	���Q�Eq�o�$Ӧ#��i��G�V_���m�>��LC�����ثV����~��Z��k�Ԉ_.��}9���>�o���
G!���%ucX��č-�!�Tl��.~(�_�$��Pi�ǯӯt�7� z7C[��Oѻm�~;f��5���XyE*�]Dt��o��AG��)0���UN�r�݇_�d��M\��YH���ؚ�Dm�R.�b�$)o	 �	��s�ʅ�g/�µ���~��ݗd%D.��^��l��gE�
�1��F��q�N�U��Q�&�G8>���J�y�c�8d��?��3�+[w �@H�Ti�B�f��xP�5�N ���aBk��i��� ���������B�l�����0��N�#�ƂJ��gr0���j�t5@!��\��T��h�x���M��l^6���~�Jv���C�:�~�8I&�J�8x$��f�JɚU�=dV�CQO]潥�U�M�q��0�/��t0���O;V�����7w���e�����A.09�G�>.
T�X��M<hĻ�����D�S&<gT����3����Y7q�x.�0��{3ߍ��S��>���>� �iN�&n�~+��+��Ay־y3 ��s�{�K���O_�3UM�� 7�H��<��ʮ�t��lG*�A�ʼ�[AQ_��;9�ʡ��[%��ٴ�aҏۆr�&k��ƻ��&��27+H�%�l�d�����@p }��C��bg�i�{9��^�WA��BOt$L�#(�nml�t�^�Ȫ�gT�U���zR����QM�#�H�ƺ�mz��Ҡ�*2��L�1��^�a>�l�L˳�W�"���<��r�*/خ�A�c�N�M/?�&��,�жg�}�	�)��|E����
���UQ�&��J���ޝ	ywQ�T����8�w`��.��:�us���7�_�_�=������\xEi�*�ҥ7�*n�w���gC�\���Ph�����s����5�K�� ѕ!r�9�E�
��y]�!F����`����cl�ܶ�M����f�Iwzh+�e\��ݏ7���c`�4ژ[Nۀ}��0��J�n���@�v0�I�c��>���~�gFm�1,������>Tڅ��#�� ��Qu2X;�uYIr|�p��bi�z��/��_���oA���&�?}���(k���6V�-2���≚�[�oV1�ѩpf�mí$m�X��ePE~ .+�a]���$�}˃�-#M��Bι����E,��6�mH�$ci甽��ϵg�I�ސ�Fa��)��3�Z��x�����ǡ+S2k��(K#�Ҍ�3��fTک:�>�K�{9�wAvt�0��Sh�Av�+��<��O
�	�ë�bD r>T�3{�@ `Zxt�	��1@��_P?���qȹ�D%j{�癞�u<�#�S�����w��8�9.ľ>h�ށ����d��Fz���q=������0X�?���DA�,���U��Ƽ�i���y8��]r�7�J�1XT�<ly���J����W5�3�rP΋��#Ϩ���� K%r�=+���5�u�|P �E��Bv�
;*�T�\%�����I���"s�-�|�/5,@!����܌�� ��ޝ���&��� 4�˝�X�~�ϓ�� ��v���l�$:���N�J
f��s�li�6��2���E�Ւ,��~��c��1�xk������,оVi�����~��p�2F�8�S������-���[w82����Q~キK�r�����Kaڷ���Az)����������D��!E��؏D���@ 6}�@��B��p��_5e6�t ͠I����[�}��Y�(���OOӰ�Ǜ�C.m�uIk��,gM���P���J"r!"J#�wq#X���oy~i��V�;�1W'��Չhۦl�x���m#�F��z��VL����\wɂ�A���*7���@Uf^u0�i5o4q��M��a><�^��׶5nT��Dn�l0�����w��`��~i2u�P0���4�"�GG��f�ڦ:A�l�]�y7	�A���ѓA��5��l�u�h���@K����Ep�� �UldR��=��M+8s�b�dx%"�q�죖�ċ1�Q�����R���tX'L���lL���t��`��#��� ?h:u�<��r���%r���aON�>"*��#����nٚ� �����gE-љ�8ePFQˁ�?�Nj���F����$^<g��Ŵ����l�:�8�T2,��M'@��'|?a�3]��������JP/#E��A������D}�52���P9	�&R��:���$�Gwꢮ�#����wR���A�^/L��/���ʂG�_%E�:�` [���~n��I�c�����3�1�a8j4��W�V;j���d�[�&(GM��y�W�� {��ك�2�Si�������z��_�O=��s�qO������i}��T�klC�9��I('��4�U�ts�D����^���8��)7�
���z�S7�#@F�,����;r�i�GV�����$�g9#ߨ�g+Z�`c9E����T�#�D^&�<�d��".u���
����vUȟ��a��sp�f8��B)���Kz��4�>?�@��Հ�S�G<\�d9)��Jc}��EDRd��2j�S����>PEa�h#��0������7P�}���k����j�I�g���ӌ}��1&���XB�;ca�{id�wPxR�3�ޟ�-{={� [ӈ�˄(�b�T�2a<�������>m|i�mQ�B���gw�Ԣ6G�=*�5�]�JSrg$�#�����4�C�@
��>��ڌt��ȹ������G��T�X�I�3+��A�����|Aƒ�~Mn��Z<~��� z��XƝ_��Y���y���!��ԟ�Ev�&�A�X� �n���NM����0}'Thڀd�F�SP��Ӈ:�4V��-/�S�;ۆ!H�`�o��-�l��ұY�I�u�xU	0�r��C4uh��$��mt׏M c(�A@=ӃS�l�O� �i'G˟�L7ΣC��6��S��Hϯ�C�*ZB�lk?�t�=v�MLy��Q�Ju@nN�����jù[��#�������@��Kl;�d�&�p�,��l�f�"<�6|���4�P��8��!܊�.���oe轓IXa ����)5�_cX۟G^{���86��CZW>#��N[6m�N��5L�*�3�!k:��|��VMق#>��<�r�i�;x����,	2��Y��߷5�Y�i�_���}�BFy���6�/-�҉����M��㉒�&�a���¾�!.I�6�*)H΋T��>j�Ȓ4�J��r�}�w��q������p䗮�x6�_������3�l}Ө��![K��+�k�=����A�_L,�M�ь݌����L�*;���[�����Ƴm�L�2!�9>(�U����E��`�t�۱6(��E��OGQ�6Ԡ���}������f�c��,�h�Gei�J^�w/t�A����5�������:��;D<N�|<&�'����YC�6.�{��ř�(�A�޴�(<�tM.g57�
�D-LqX���>�`�p0�����C��O_��|�4i
#�la���$�����)X;�K����a�_������l\��%�`�8l|E6y��;M�B�<K�TP�K�/�:0�bߒ�&�H�5H�8z�M���3l>�W��I�Y��6���x�
�~�8#J���H��H��Qɘ! +�(�{��B��	,I����D(�){
lӹ�(Ű�DH�A�=̪~H�����#JE��z`�=s�!_oL���m��\CA�I�%�T���*��ӗ����?�L���A����-5g1��/r��*F���	B��dN�)C�
�0_������:��k�h� Ѻ�K�&�G?=1��������*gރFXK��
����<X��9ڿ����^�6����hM@4�}�?�Y2�n�3h��wؔ����i��L�V�5�h���_s��c��[�K