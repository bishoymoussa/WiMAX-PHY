��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$Rx�y�<��wA�*;�x���@�̦�W�X�fa�M-$u����n~�%���P�$��W��kYَ���P7�?UMfT��q�6�U��k�>����~�\N�(�����X�e���/6U|)�X2pF�]$h���d.���9E��WG��L�X"]�Ad����ľS���8od����e�GT?y	7�������ݵ�^��R�q^]�鍦�����s�ae���h��L��P_���ާ��YЭF���'\��68�b�[����w8�[X��V�F�0͘3����q諵�uW� �h�u\V�?@��_6G�_�*�G���B�絉�f������[�G��U&�����~�F��AׯK1�`c��[<��FY���4I� �#�G��x[X�=�Q1��`��R>(�w����R�O�?����7�,(�H\�#h(W�EH=�������yq��Ѿ��aF����:�U~m<|��.��0=�P/���4ǆ���T(���bۧg*@������yE����)�Ց�cQ`uy`�8�ce���ib\d�TMc+%���3���5��u���r��m��^�v�h�n�@4g�����Ks��9ޜ�f��:b��nE_�
<R,4�~�h>����-̽��h��ˀ��RQA"Nb�U�{���w]����O�Q����ߎ��*���θ�/"|�C�����f�`����1�2�㾫��Ԉ��x�dMb��4W���J_�'�K$��&���·�<2��6�M�[>t�s��։;̛�	���h4C��ٲ���y��dW�l*����w~��a�?���Q�Z"���@,F�){� �Z?�Ơ��ݸ,=TE=�F����q�6q|�d�lKa�i2�"�ô?�=|���P��S
Zi����Enb��i�U�W�׾�Lh�[�#�k�ځ+�`�݄��"�D�{Ѓ�|MEY�ܿ�h2�E�gJ��;M���ҷH�����}����� D�
��+!�m��mL�0��۝-��z
�� �W^�թR�0�e�߯K�]�ǟ���2G�6�;t��v��pI�J��eށ���-�}œ�Q���_2�vѐ]��\�~�i��d�Q�������}v�J���R�m��E���fӛ �RL�x���=�-�}v��3s�^��~���Z�Rb[�A�6[�^d�ew��	77��i�� �/^�����s�}�!��!cH����9�՟�&TL��rv8�ˊW��T�D�:�URP��&��Iay��a$�� �-Oo�r�]�D}��9�:p~�a��g�0�~���������ڇ`I�Z[�"�����j��7{8����&��y<���F0V$hS��_F�ڞVХ���]�9�P��C��0�s�H�70����7���~�5��,A�i.y���UTQ?(g������5mD���4�:�	2z��!����dI=q1z� ��B�2��j$��1ߦ�b22�Qn
Y�b�W&�Ʊ� L<Ok�1!��=3I����c���$����3�ݖ[W��>?���hJ���@y�k���N	4�P�z�D�1M�$Pr�W������G�T�''$�Jh	���t��)��.(���L[8�H2�T���DyMXL+���*C%���-�k��C�:�\�������1	�î��@��*�0;U�"�d�����*�����_G�ɦ�sg>u�/�I�=�@�N�ư�g��p����#MѸu�X�HP�ġq�����K���q2@��(�A{��SY���	&v��+��B#���M�&K�!�,�4������M�Ǌ_b?^wVm�{��ټ�������Ap)8g�'�o*Gz���.��[TdD���n��;�pu[D���6<���Y������p|ʫ���'�rjq�#��#`���<�q��pL�sh[��/�f���a�Hc�����Y^ŋ�_��XU(�j8-�H���k]&������:�$� R�2���o�������CC�$��O�C�F�����%@u��AfZ����W÷s��ӿ��%��j̕%���<M=�5�"����d��AXY��X, -��|�O���}���*_C�����5�S���k*��=�vV���q!��0׋�5���@ ��J�G���_���>���Y�����W&����˩�e��s_�Z,Ӌ����̀��̸S��x�&�������1�q%>�o��V�I�����HH�7@ͦ5�;���L����hA���97�Z�y����3�H$�nEc_�b�2ބ!�i�ɂ��5���ˮ?te��YJ]��)����\�- �X�Φ���������%?��d��%~�����Nv���.�\2�@ρW��b�V=BP�"3�=6�¹5H�l�$8�4Nyj,z)`l�6E���\��\����\.��/��ik{=��ݾ`�I�1<Z ��~�2j�'���H����7	�%�;��#7�O��"gOH��G`��{���cL�M�ɍ�h����g�9������Q��_��{�?�1����>p�(W�$� -8J�b�T���ޔPJP.m�Á���wM׺5-)E��8�Rǋ��3u�',���v�����g�=�{D�R�B�����O�E���VR3k�NY1�ü{'z��O=����Ә�n�]�DCmaS�&��7����a���$4�����sK�0c���C�O�m�x7�{�����׎���Xvx�m"�'�@B�Ʃ1��
|�\�����"���	c����x�A|�L�ѧ�<p��K�H/l_Rn��-\3�*�Z��b�D���w�[=�ۏ4A�e����P���$@�$�g��6#��2{����i��֠f���"��.��#�>2& h�m�
����T*t���U/9e3߽fn�q����Q��7<[��^���?�8�������hRWF,޼=�����f�1�
y}�����uQ�'`��(��-��DV��$�̰��)�����(mc0��t�#=�`��*�aٍ���?.�@�q�E�B�Z��.n�t�Xm��kH}o���(�J�6%��;)�?�(P�cD�Qq7�>�Vq�H��Y�"��隙�*BcӨ�v$�ːI���i��eߥ�	��BN���q0Q���-���n���R�+_O5� �֔W�ۆn�@VK��n��B4�'�~��<̈́��L�v�Z�_�_��.I�|�>�o\��<k�>o�sz~��7À��5O:�I �ĉn϶����W�jd\Y�@tO$�9B[w֡���گ���F�V�Zw�5[)_�����/��t�U�,08�Pɫ���7�X$�V�����ј����p���A�/�(�|�ư;љ���������Y.�i��M��в,�EKg��;V`$q��8�!fw.
r�{U{�^�Ay�~�cA4�R�\��M�*�<`5����"�mIHd@�e۩�-�.�pM�,���~a؆�K��Kj�<E% ��'�(? �19͎)骢y��Ձ�V Ǒ&P����,�e���3���x<Wb⩱?��}�Qy�;������E�|y<"���8�M@_E������`mth�'#�$�^I�V�Lq7����(yX��$�LR�G����n���Z�fB_��|S�%�D˦6	�s
�;op�F��F�=	L
[z��+9H��Ga�b�<�X��ڍ�]!����a,V�n���a�KR�{�>�y�,F�1�!/��JC{���[A�2N�0.��9�
��g�R���M����Pv]h�^<_��{5�퀵��=�D�S��������%�$���=w�A	���讈��4����UC�"hnԾ|�f�d�̧Pߤ*ޮ�@��Z'�pꁔu��CA��g8�;�d�m��6#�.vg����Sjhc���������9ɍS%��J����g;�z�w��S��a�� 4^���^x�Ɛ�T���Sl��z���䣂%��a���?Hn�C�"�E9y�4�6��K�kR�L)�wo�L_��f��:RK�d��Њ��~������j�5��pr=�� H�̈&c�ct/O���Պ�p+X����_#���.%��Ud�}P��3��	�'ٞЈ��pS��6���6�^`(D��}q�����cMH!�V��5�	�>gA�����������w=cH��߿����z��_��	TQO�#�N�_q�`� �s�m7��W3�@X�D���<6��S}(��ce\�H! o�� �ad�e!����9�QLy2�E�6F6_���Q1�x������U	��@c��j=�����VNER�@������A�j�=���1H�I6ا!�fn�F*}7�� T?W_^�d=�h�̭p��;{6��9��_tJ�>���m��̠���E��O�h�Q[��'�9
�.>���RX��`��*��b+A��X�>S�+�	C�ͱ�a�����򾒣�Vժzʤ���]�3���0%Ő��ږj����1^�P�_��Ë����	����A��m�.u_��jh���Dh_��S�݅I|��$v��cɟe'3[� 3M|��dc8�߾�C麯���J؅�n�Bm�� C~�f,�����cpM%�2S��0�H�@�J���7eٯ�PZ>Cp��B�e0�)����Mm��j)��.��%٧�=W����e��H�F�Ń!)�K�T�W�s��8�Ix9D�;�F�t�-��چL|�+mΑ�,�C?��?�t�Hy!"���p��M~3*�{��,��3��`�EHT��߳����k#أ�4����ȓ,P>G�cx>j� e��$A���ufԣ��+T۝��1o�?z�7h�z?�
��ghHB��7�D��v��c���Ɔ|/b��<ަ҄����ڀ`��v�؃A��F�����Ny���]�j#c���E��&H�O�fE`�Ή��^�ƙ�`ۡ�q f@����p���Jc}OlV�hBUHvt��{w���O.�G�qWlɩg��>)����"�#��!G�:����{�v@���4��irwX��(�B�eH�!�ՙ.������T�����Dp��G��t����}������%b&\0��҅�FC+���7]��q؇:|o��d���-�i��b��CU'��w�Y���.�я���^[�,�0W��v�$�AN��l�Sw|��`k��ڦܮ6�����z�[�7��]4;��[]�!�|��f{�ZDO�4vO_�ȿGu�U�	�g,<6 �~�k]s�)���#�[��s��s��STCh�J�g�B{��h3�9�����ȴrqi���`�8�A`��r�_E|��g�>��q��T!��E���~%� �;n��%���:%C���E���y��7����p�[մ��lX�ۑn�,u��M��ZB��RfN���de���P[�^�0�X�Vh̟A�Y(���;��$����	����8�X��<ؒ>��%�j�*����&��#����������u�Ԯ�N7�����V�,��λyY�3~&ch�0:i�8����w�%��0�/�w���ܖ�:&Y�5��ϐ�iN��b�ɪ`�j�"��oy9z��OЊ$fp��:+�F����6"�=b���0n���>_���O9#G���C��hzۘ���ד�ql���=�&x���Pr�N`��a�ɔ8�����,zލ�3�9|�v�1�9�h�J��	�5ZӸ:�Na��v5�S�PF�o����w5��1��������Qz�������J`����3{�`��S�٠��~S0�p�}�@�A� jʹ��qP�'�O$�#�jH	M���z�������S{
Y�����݀�x,Y�rn��,f�3{�&��Yf�bl��� f���e�=�� A����8I�\�Z�)�����W����ma����nC����/`�"��w�+t���p>���.;���
���� nT� $����L���e�2���D����x��/����ėF"�it�[|���b�n蹊	�Z���vUmI�ɷv�p,)v1Uv�C�{�:�#�O�ܶ�I!_stMD6�p܍ڮ��_P�z��'��Psb�=�ed�!�� ��{}t�kxYQ+�A A5B��8:�2����o*1�j�� I�
���f��Q.&���=z�ͼ��B�v����h4r��*��*�ٟ��am���N�JBs;i(^�H�mib�Jw�x���A\j4�7�ZR6yS�ծ��x[�r�z��EMu~��
�&�]���K����L�=���&f�|�^8m֖��׊�9�S��9m���lM�<Db�3%^�un��`����)D_x��\��0H��ɦe�n��=x;�*h8kh*7?HV.���
�A9�X�����<V�j��W�l�3�QgC#�.� ��<���W)���Yx>��hU�
]�1�#�2G�ߍ�Nk394U'���3LS.8�FY4��!x���C{#��rM����ؙ�<���,pj;E4����AW�sʘi����v��$���fS�3_�[�L���bRV�#�0�\;���3b�U	�EP�t{2	�3�pkٷ����\;�^��9�n�J������H$�^~C���'?.~b�0D���w�/"q��T=���`�gxM��d����2�O]!�n�-~�\f^?C�twh�<��_�,��އ��}�.��u�80=�^�Q���8�:�E裷�����,5ctG�l�S?N	�6�5<u_��>�[�Xk���/X&�+�Y`�I3��V.�����9��t!�ñ� ��nғ����r�x	$�Hq��|�g��Z\G8�N��(cE]k��?jH����j�q�l�ߍN9��D���!L}�q��C����\��Z�Q"��,�\�7��C@ˏ�"Ai��"XʨGZ�X�����ʌ��M8,h��DB	�?PpC�.�l������I%�I{��t_�W�D<��e��S-q����L=4J��3Xuƥ��lGZ,;'�VDH�VW��j�*6R���x�3� �T��(F���EY
������c�l#�8��c��{�ne�� ��72!x5���ol�����|��-�/(s��-<]�r��;St5���V 9�M"���6�%h�����&14���iXn��h]���V��*��*���m���;����-a� �nV��d2_�GXw/;`�IZ���F1��8����,�o66N�gЕe�G���T܉N,��,�C����#�*�6k�$aCcQ.���S�v%W�t:+TU�_wP�e���|��F21�Ʋ���Gp�fFc���BPٯ�AVUM��)ؾ��M�9NS< �_��mnjHk|�i�6۶�GH������y�+'@�.!B]���Wؚ3ǽ)�7�g^�d��_'�7|�Ԙ���.����2E^�B�W)\tx�.�W�����s�M�g�JLo&�N�~�*�"�9}��k6����Y:��`���~&0zZ��)Z 0炻�̭|�R��I��dy�Q�l����D�;�9��>!ڍ?o6"d���)�_=s���ԏ1B�MD��nlB$�s���(�gVj��q��>���!��8,��/O��g�1O��ѝUi�ƚ�(e���77vJ�[���D���_(�6: $6��y�Q� ��������.1@�?V~7.{��]�r�u����LW(��*�jd���C3R��+;P$�Al~j�/�;���~�0�r,Qg�yp���Kp���2��9URL���b�����p��ߟ6����'�OQ����Vb�
��H��1�k��`����a{g#��Ãg��J:�$^���R�]mG��-$�Y��X�E���/E�_Z��>#���དྷ��4��F(!�}����A�}Osn��/�b��Mv���4�Cg8�
 �F17��N(X�JV]��9��N��d)��<O[�A��냳���J�1�=:>r�<�fW�]�ȸ��*�-��mH�-��%7gN���i�E��	�͕���P0T������U6�P������~*Y"8(">�N-�8��ȋ�;����J_���h���8�}�p��]�1�����Z;�����ɟ�AQ^iر@1�7��ëᘌ�UJ=���+�̣�m����E����q֊v����<�u?���s^gM7�)'2p�~���Ifק�_�e*��5;HQ|Sߵ��E�9R�\
��J� wDU��.(������[Q����QR�4���g}C�g�֏�Q?9}���x�zt�P~�H�1�Oq��Mt�`3B0N�c�!�|�h�h�)s�Еr>.��|�q���v�cʛ�օ��
��F�3߄i2��>gx���t�9���$<h1��͍�����"�/�V���{CC/J5�TV�{�񂚡�?�J�&1ϝ�����nP�w&];����E�*��'C�������c���u�!��)��m���{nAq�ִ�nC�s	ں�[^�W��(�i%G����78�)��)|��_�O���Q�c���6�d�U
t0��}���OQ��ц�V�s�L[�f��1�P�KOc^#q ��1�N^��.նy�V�/�-z�(	�MU,g��0а���/����5��q�.����+���P�7��GE��%i�|���M֊N�M�,m��:S*40����-DEjXN$7��&��J�,����Z���Ae����P�n���R'RI_��2����7"��m�[^[\ h�Z����^�����Uu�;��#Yg�l}����1����`�^Cw���h�xd�*b�_r�ʱSq�&�����
tv5��mM>+��F�r9n9C���ǉo�mMV��$xO"��>|�(����@ν����,#�4�s��O)/wI�lm�J�Ǖ����Dc�:�F+A|� �v�=�3�pVq��d��̹{�W	��/ ���O�_
8M�#+u[���j���c8�Ok�Q�񚶑�d��6�+֣�]2'����~"�q� 3���7��呮j(G�\r��/8q����['Bfgt�C�*�n�\���I�O���g��(���pay�9�q;sc����
����$�nF�_�������x��Xw�J�u���̤�J���"�8�t�蝨��>�A�ɝd\P=���C�>&�y|����<���a�/���sbEBkn�$��~��D�������ml�(
�b<���U�􆢓�nפ�D3�od6Y����!w 	�U��E˳��h�����������q�|��}�ծFXA�x�;ׅ�] �r5�%!�{ǆ&�������rV��E��|���V~(\O,��<�h�%�1 ���3�gN/s��^ƒ��
n.����f��Ǻ��1��.;� un���ni�.�2�p��=[�J[�m�3Ɲx�΁�-$@�O時��P߆9=��]R8!{Y���Q��4���6Ij�
�j�n�5�PX�9d��,�AH�S�$==Z�%r̨��-��\�<[y�
�c�v���@`��s�W� ��<�<9��Km�D� ĵ/�d��[�Dbu�cBL���h�|a�2�J׫&P����D�Q���^8�I��_u��<K��X��O4rHU���Fi��6yg+ �;�A��M���N�dQ -$u�uHC����97V�ju�8�}NH�4���I��|�Om$I�B� ٔ���O��~X��,f��C�*qcI�M��^F�?�Mt���Tɘ�9b�6M+KC@�Ja)$�bnv��СQ�_�f��͛ީ��4:����r]�am�3��	f�X\`��ѡQL���R��I�|(�4��d�1��}�YT�@�	j
�������E�b��^�'�[p)�hu����I^md��0<���<ȠNt��Z:�=N�/���������,�Fk�0B��6r��X5[W�pn�?�~��5պᯓ ~���������W��+��DSw*���-�ў�	��tb1�V����)X��k V7�"4�(~n}�]P�a��������m�"g�?V�=��׼���#d|^�X������o.��^��;{?TZeáڽG�܊�U�Hn�5�kV���r^�|�Ԝ�ϐ/l��e���a�e@��M�p��n�N�偽Hi^>�Ӥ���z�~vC�1�YF�ć"�"4�g�إ����cB8[<����kxMN�A��݄-q�Bb��V�����d�w�"�@�.㳌�����}ͳ�[�]���#�{�v:�g_?w)��F�Y6�}ئ�f	��B��ı}n��mm��3�W"k��t�_'�'oQ7���+[�m~�S4��7J�Z�3��������_#n���>�S��wR潌s���Ԏ&�*�h�T���u��KKçr��`Ȕ�N'rh�:�O�=x(� ���#�mzO��N�s�~�1o��\���� �_����ſ�?b~���nS��A�߄x�D���%�D U2�9�H�Z���Ni�Efȷ[Rwp�(�f�|'bܒ���Ʉ^�S.{̽-b��Ӫb�x���G�����/�h�X�ɳ����=~�'$q#��LM�{�rx(�Tb��|�Ti!@(Pj?��8~ף�:	��,7��7��)4\Qv��X ɷB�d�F	�a�[r���eV��]�A��N!�T�e.�����q
�C���:A����?C�U��Ոy���b��v�D�x�v�E	w�����UK�w���/U�g"�c�Rj�˛�1��@���Y��4H:�nZ������_oZ��5g�r ��x9�iN_m��i�bdO������3�`������I��,%d��:�C��gdQhi�6�@���S�#|xY����`c`