-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
wBA85q4+qB3b5Js9cW1qISpIhLkNeke+jHPX0vVMKF5Hllru1siFoTjhKZiBedfd+ODhN/Y66vp5
Ang0NHlR0cKN2P2keRlIwmhGut741O70Rqkko5caJ6NnKH7WNBcW+/dvgFS8Jg4CI1HJgGixB4Nk
2GXnmJLArdk82Stx8ld9GbqCen4FclKx7yABI+UY2+oltnd6NIroiJ9UoDMC2vR+EgEFbybsiRsl
POcv0t8lqJzOYUfODthpSB9xPFSZ/JTLy1MSxezV2vPSRweezTOE9AVmn1p6seYDjKfNoeoskgw9
DSdpTt3N4Jd+NdxwhWgveqUpQRJMsZY1sdq6RQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 8352)
`protect data_block
8c3Og8m2wYTBz2L3IotO37guXjFHWFnv9ABxxlbuU1GlNL0FhebItwKAQplnDqrDax3WlmLvwpLw
jWY5wGkzyuuqitLgNOv4aOz3TFt0nIIDUa6CRhfBrJ7y3tHpUt1aUJJ+fKjTsTCVRTa7dFmTEKEF
+7IXzObGzdOyWRK0sJRt4CClNGMC16nQu4ORL33NS4qdAEvZFSJrTBiGZLCz0nsklpxdaIQmS4bN
0NOKodn8Qtrq0ACf+VLr8Pq77YnnLh1t8nDkBHFNvzEosZtS2tgzooOCI2Cackuk+Wq3XcDxPrhB
9JMMw4s8bT0iekq9vQfDvCOsT6FFMvsVZEqsCu4uwofEONZ432HUdFpNVhARTm60xbn24lboXGhW
5v8tyITIjEaNL1mOCDheyYFYagGLy+27gHAjD499dhmffP7VcmLnFBO4QJJAvBU4xNyl/WB+UZxJ
DckZWlXIq6FtMUowHjVd4dWHn/IPEUftIi9NBD693UPSah0qvIUMbJtvgcgZb0osqTXVc41D9eVP
67Ut4/aOtA7nI9gcR4vo2QumOxLseYcsr6YlWr0uRhgk6heGWIiNWFlZJwTIqsGSnlpeMQ5RZxZS
8yZh99WwUlNiomGPouokKQN9IpKX4AF4FrYjVyeeD0by4CYxXwS0yrK0goqaAFgMcGF/P95QnrR5
EwwFLA7QmpEuIXo5Xx1PlvU4Q0gT7G54gJ+IX5t7a6AocRxXEERNdNAUakBQ7HrKdPvYyZsxXKkT
HQ08JedrksAiEHKijhyWTVbntyjNtApYAIXve39xsdWgePebviz1r6xUXe6RbAbXv+/hWxhBMwCt
g9fxre4XpHbW2XAzKZoMMggJLiUM1DOx1p+lBlSa47u3SZjuu25tYwmRwiggImqHWzjmBbmKZaBs
R4PcE90ocFo4yBUSHTLjxpLwcw1z4H9RC2v08DGah4DMzK/NilwGPcwXV7He41l8mZpqPITQSB3I
Cbf41xlBICyBge94fU+yZf4yNQtMljrahjph8tcaWF2ypaJBoqm80uweM0RI0NGfTvSn6guZA5Lq
8HyvQj3i1fBwfHcDEIm8J76qWWjUUW7MfvhIdIBerIZxbcQ0QXlxdAnPsCDG5EoM8nMJfY+sLoTF
lvwBY4DqmEnx9RJUjyZtH0zjAh2m75H/xaSF8IaotlSDKVjej3CTedOuJahRZZpacDuE7+dcku2I
0SCTr5QIlgGLDCSzLWHMFxKxdcWGLElSBTCdGFtCZXTaa0yHdAoj97ajabH4cWXHYpd2TmuEJuLu
zjpyxtj9vosvqMQ00/Vh8YkuJv6B0Ue6evI0ICnZpqr/Fq21cpBQCyYWHVVE6bhsvj5pH00pEdZS
NN8hTNOqY1xXWa1brD1HxTalk5gdZlxQ4ldkPTai6BhVwN0Qk/GXBb6EKjj/XECnbVFPXkSMMxPO
15Q3J9IPgPkQ/gIbXJzuapt3EstKP9fngmF9HUkSsSfPy8AMmAcaJX7Fn+HXt/+KnsIFFq42UjNg
cPatRBRk7RWCBI6rxAjUP6v7UqQyOU7F1iiFw3J4+KyDzetER9UFTO4gjQ+U1mQoMIvd46KfVor6
z7nOzSMBBKRcPbf2/kcP4XdX8wxQv7e/KofvG4192RK5YIUZMqWJEviSpNJwo0w+Qr2hMGYGcfHo
Ov+/cqjhjwSitsIN8ixMRmh1MxA4LnHxQFvKKQVc4S4xe7Qac9FnUJEuzBZ26Oy66XbkU/4uHIep
y/ACihYOp+huQHg3gdgP27ph8XqdcW+cRDOATwKjgsdOp1LHSyJYmh5ht4Xfrz+fS0bjiBf2hB8v
xvudKpf2OfnKa9eNhEBrFkzgXMRMQn1oEDRRosx33aqNYiqmMt/O1xZALEyEFCfEVv0NXsqVJj8u
vuNWW8vAYzrpJC8LQfCYTC4HYc5c+1gcsEbTu2u2roGJXqSPmdeZNfYJzRVthyF/oqe3hNpDRpl/
xr4dGLyzf3UaiEn5BFaYONlJ6UzwYAGOAHxwEnYW6IQDQlq1Dkq44x6Tp/odf+uyV6mInhVRub/y
4bva1DSgRnXAj9U4+lVGVLNWxFCc5c95yzdnAwJKDPstjct8p1U/RJPTjp29+UcjB1qkPcvUsQwl
A/coJWaxAAFBIaYL4Adv6sQQK9oANw5AVf9yjipDbLYxvff/E0qmrqj1bbmH9fGr+4uPSxfVb+w+
mUEKOHlw2Nf0ItQztN+7eY+9NptbDYsbHf+0fC5SH5SKHghC44XInScakcGZqrVArRALi+0qAUpF
NHlCAjb2UuaCHPrjHbMMURZHFBYX3/lpPGW51ucQ0gpy/8oYGBYC3wpt3DNt0zV0v1Z2G66NCQ5k
hkoyBgQdUgdq57LSwZ6LJ/89wEZwWtBwbr7l9kldSxGIKJy5Ovm2SJ1xEJtcmXaUw0ucY/gGJvSu
MLke1VMGxpIpgj+IYGpnbdiTh2xxZi53L/9Ovd/Wlg0HgVHRyQLsVPwzDBgR4dzflM32CLQwPUmQ
HEWWP/uenZ28JCesg/Q56aYbKFxsplnaq7NVwLCDiW1aE0tHWvKkXG9zoflc4sHwMI04WChkrmJn
KQ8efE33wcoX2U6sgwerTUp/LI5TCN322qnJqzBsr+aUOO1sgGsvo6KFgVX0c1fE9RlsSUmVySI0
rTBivNAThp0DwQOqbI/yyY0Yl7DMFYOMnn2SzD59yvQHgJf1wzGbVRxIm+Ca3/Fby9OpvIwk4ZEM
0fQpPTxynEokZnO7HSrrbfeHJCA9d1MGYn/c/ZolCz6ys1Vgp9f/yuH6+lJOLEW7ew1mDJbJQMTe
9SZUD4zt5kzLq77HmWwJ3xiPaL7iPfnOfxloS31saIzzHqExjICZHaS5uvQWwXwdV7GxdvvtveFU
Kx0/nlmtt+62TwZqWe4uRWGWx5kWTFU6bGtR8yLVV5e/oY9x/aRdl7RuwhNSFUUwquNbopFV70Zm
86FDktLZYj5Jx8seM/FZ/5VTjjxodV69lm6S8acZb+kI+jHT7163qLM9v1g+2mJPVmp2/I0kl638
EJ94OBD2qFUFTzZquj1PnDLIJfDyb44hKkdIuWyBdZi7fE8xAM1qmnpCVmrNYFdIdk5Yip4VjzCN
8Z3KN1Fmj84xnGuAo96tKsCV3wFaceqsjnYvIYnPNIXN0ZQ7gaic0D/8ZmtLvDJW7leykrL9z3s2
WW3oB/ZFIBbfRa9VtAwtwy6KYnJw/0bcIcDvyAI9xEjm3kVmXuUVdV1aaNRLeD9I9hyeqpsxFAn7
gYbQy//4V/f6FLQMM+DGVYJ8LsydOuuM+OB6nLTHNaIgNd6QtM154r7qx7Gg9QomYr+DzyySwGqq
Xbse+TjGqJWCmi+H2PprM1Ub2TZmU5AkhnXYItCUnH5Ybz5n+JWI0CISqecCHLSrVx/wyYGISfZi
6dRs5WGAkin5NBz7PtnTTEceiEYhScjAKBAaNjfDD590JlXN1J00VfjeP4XXqxLvUMmLx/uyOO3j
S2IZkr+oaXBhHq/7xZueiqCzaLADD4FcunULf4wJA/9m35uJeCiCXIg4NZGfyT2wz/8wQsHC/Otr
XF9jy6K7hQRfzWUVrdpKQZwqhSSa4/tjqPVaijowOo1cDmB8nEjF1voyAXrMluOKxQCsRHMF0KJi
aKEijUZOV4I43kEeeP7Uen3eq5uD730+TDWGS3MqbBQBzk3pLTqygKz4XHuNb9PHyEjZraUoaONG
OmMKcfJQ6i8NxyfPgvnQ04Cp0JlF9Lj79topsbONf/4n0538W5oeu+TQuGoafwqeAtiRS0eiQ0nu
+iDLZy+6L2gWZ3PRLbrtavobKiMbr6Mt8MGzQmALqtzHvZVm/B9mF904wbp/QoLyF4H6fdYtxyzd
/OfuNMM6fhQk1iNLCxJd8D+eIGLY4OTDknm5JmE2CsYfdF+2Gx/mNzQddOwJnoR/Ej/LiWffqLVq
nmy/4y1PRwH8YRMhUH1rm/9Skpy3HJe/YWkXToIDhNmBiGJDY/r9EVViAFAPWMk1CvyYsw2USXQm
6JOvIzKn7hyWMl97VkR/Lj3+/qS17jI9wXYkaYhmD201MJtV5/IGwG+LYsAByBFuL6NupFWmVFl1
qOmq+q00+FFVQKrhJNHsP1TWf0dEc/xVx+KtpXI1gMhn2Npkq+lhSllneuQQcU+5rrdSudj68k9c
SGqm/mbv1YyXNx5npTU2pFxafM4zJXItreOuQgpRwe17JYubQhTDwlmOgsP3aIUApMksZ90Er71P
iKXBOssWio1mEg4p8l7QGoiZYVQFOi7+nmr92suAAVroIFwIdZ4yBHN48Iqa01TCO0Hbgm9gHa7U
gCiGtV7/D7DpSEdabGs99OTnI/89yYoa2YLf8S4Pv5GrEzA8WyIur2Vo/B1356T7qV6ycd6pZ5V/
0HCjX1WGlWL08BsAnhUJrz31Q/bEk6g1IYZK5v7TxOb23a6W7F1xwI4l677ZKHG02z/bl5NxGn84
W/n2IbkfcEBEN9Jw5zYKqM2bR5aigJVR8p+weZwldkne85mizPObG1GF5palGFrpz2aAZe0GIV0M
SvrJXbjU9ommanDdLNevxw8Ehx46Agxl2ddLYZxopocwf2RpfUtKkMUi1MPC9piFmdyGMVdlBowe
B/VmaumBU2K+Sj62x2PDR1Ij9gj2CS+vi26ir8rP/ofly5HNGuUzfHV/dD1kcNjupDuusZ2dl5xu
gqAAy4HSiw3iOgouXO/z1FEzN0RUH5+I0AGlq34fflLyIRNkgh8ilsH0MmDA5Y+U+ik6pMsW65FM
hZcP7McB0KZqYYE995wISCzGvjR8w8f+6tFi9yUF3fLSG5fGjq1dBcAoN76rLqp3xswdj7TbusCs
hzxSD3FjSl6UB0nlgBcFUQp1TAutt3AUlgUCJZU2018ip4yBPs4nNHnvNRw8pTeDKsGJsfJgUhYh
RBUMXmD4xAnshA/Z3IlakzTpJlTlxO/XtCIcOok/FUnImcbXX3z4YcKUyumNDAehtxnlc/c1A56W
GbFArraVtgVUYoz+TuEtM8FcYu8kcXDcogLLXGbXmOXP3HCl292BUUWOsS1cAS5GBqTWvy/qgr3U
qstrdT44XxXIQrUTOSMgZ1SIIpFvi3jb3wmO0xPINIuuwIP05xmBmYiiTGUzuGgHjuI8PtMAtHT3
jg8DQKqt3XVHq9G89BQu0cHdJ6Bahja5aog6H5PVngET7Ru3FlSId+glnxHUOtHtOgAft1hXNC8d
h3lPHqi+BZWS2yqo2UkdOvp7wtntJh0F6Pbc8T9w/VVDatz06dBXk2JLADsqm1kwECFe4Dwvciqt
0Tkgg9+BATXDeTF1fNCd1SaI8zX1vnYjS1qdJVkzYhJSy8kik0o9wavwNFBL0tH3AygJ+J2wuYLU
yh0616Je56z5B51l18YZgsAUV4OvGMMAJQpKNW9ThYHYNHt+OmIc05tY4T5Y2C/dXNIzxfjhTOeH
Sq8rBkOOObxYuV9Rk1QpbGO33O2ppXGNF352LD8Xn2YQzqoS1yuRNmvcIB+ue5793X8VdE757PzY
bx+3g8wOKJDxnCbz0zOHY/oDYnCu16uN5+3x6/fpyA0NUDkPnXTiN+QpW+3s1mwZl9unDpNIWjAo
7mmD16PC+wdQcUBC2xM/66l46fUKZoSVkzLoHgNoBz1/YhytbkzZ1XHwjbko7BLi7SOvzF703G5H
Q70Fx3Fns3GupglbyesDtg9aWmbbka+Frj+vwoE5oDdeBo2iuTXkgBGjB3DqatjzW/ovuHwwTrFU
JtDzfiGrSlPBTTy8vWvIiNqGly2OpYRaUx0EBhuFtApwNmuoBlssFvwSaTYab/3RpX1XJb56ZVt2
Z2E4wmGDioZMLZ5n/NZ1TkmWFC3lwiCfR3QYePTY05XYTAsJCJoDD6WKvNQdEv/CVCAhbrNB2BJJ
f9qSKZLYTGh64y4Grk+HEQKvWMAZTrjqKcMbv8B/+X8pEIUUj3YEKYMlLIrvcFrBC+FtN1/NKVxp
lmq+z6D4dM9IqS9ujf0lvoiVf/hZ8LB/R7tQeWYPUqJfkgjc4uxpFqausEOpW4BW3fmdOsZtcWln
0Uyyyubt9Gxm8ihsxoiRcVM3DTVkrLTrjeom9wM24GXVi1qlb285MboK4qxRB8XUBLlQF7PLblRs
kHHgFQjE2rBZmyjdTh7pBK9EwHsckW7HCI+oDn7lIIpDSWU+wlUogt8PcLridy+QhH+mtrZviOjD
pdK10SKyA2PrQ5fk7qveA3GAJGEEqNZKSt804gxQ03lVmyrQBSNJq9oRgnGB+ngGBXHfl0iWzxSE
FMqbwNrN9xRxFjmFkS8VdciIjP63ToaSp70U/xI8tpFnI/VoM6l8/SX1UDTJw0FdNh/4Y48oYR64
7/6FdzsazuweSt23+p/rVre8BveCjmQxNkiDwSZRzDKa/SFefpZtIluzUNjO6oWYW3zbIjdH4bxO
Pm8XM3Or4k+ttFQfAChio+MXqargc8UojIbthcUwqKt332La6zmeRL0WXWe+iFQQOz5ZSDX7Sobx
/AygujOmELFucKsfftQuU/msQZhjsa059Zmty/Nyc0ASMkgoeb0NJY7ywkB3wgqKJj96n0DX+Row
XPk8QUBN0dG6iZTKUOa8Rmc0Rxz4CfwQV/ulPnKtHIcGqGEcNI359vYlEuAbZs/QCUEEA+oImuby
M/EcE3zbeKPTZeb/cABl+bywedK1zx5UkNnJIkBiF9nXWb5+WvTVyofiJLTMkVkx2/Ro5X23zq2Y
VRiwJlAJ9FkUKakZYI00wJVfJ+mi6/BGEFIGopBdYqCfRpccWsUSihtRCzXdh7k94Sws/5JXtubG
BZtXFpu1Yp/jPGzWujwNI70LIzkQ2nnZNxDt80/ZqIPj0EJwEBpHrgS39Nvc2rMU1T5TnepNYq4y
01SPsnt+GQq1laKlee2AZORFBvom/6p5nE4yBKTpxflnNiY8x+qOznlXBMy6dtjIag07boF7VSb5
+AEX/nCw14RXozYdgIIKgaSS1uYEnIC0H+PoB4S5e/QhxY1WOPdyFW1G0oqTEVgTU6QONfj+WszW
aCiGW/zLxnWMaeJb9ng1R0Jo7wx86gnTwXqBikXFV2QFOL+d6kViWWwsGb/VmQ+OqOFON/b2V5Mc
E0bS0F9nc1F+nRgG2qNnCH6RruVdo3FXOYhrpa/cCGKK6/7KJr6TEUe7PLMd9YSalO/vzAsi8N80
cqWyUF5iUjyf+QVIW5IHZLj462NBcRyMz1TzlFKVOT513PB/3kXdIgnZvIviAWsL+xKTNOLsok+B
1ZV6EOuFCzuBdXc5BgcKPI972pxiEaynZ53VjbmQCC8svKQSiIOIjBLqrc/tuY0wo2mU9aXlZKxu
SQxCjoQM+ols1pja+T+/bv/NFRxiV5JKQHcSA+7GR7dDbUzyRb85tBnoB3c5hGyIAk9cfx8pY/ZQ
muUHBcjV29rvpD0aY4LC/MsS+kHjcU0CbZr8EupJHaStIBolC5EbYXg7xHI0rJtNB0kurRTRHLMA
86t6iUFQqFyndQcwQAFJdW+1dQXRxmk2shm7YV/yW56zxbbLTH1eKOWf7GGB/kf0N4R9RymVvzlY
STnKkiuofXOT0C0fN9dCYmvqi+UEUezuX5Yvqx95tYkKnOfWv9GVdioNtJofEC/HsVTUM7+hC2Py
ki06rtjPPSDn9Zc8eGyxKbaDkctzIJ88q6aj/2NMytnoG+8Dy0ju6fcY1hXr/DsVAbvhUU58q6Mv
xgul7O+lEeEDTkdCp/VqWg9FLJHBScu+hl/pXGC+xAZEy5JbA7gtKtvEZ/t7y+sX/4vca+AKswgK
MQCBfgcAGGiJE3dp/O5fcGGi9BlwobXD5QWnaWRDrbRp8acomy0jgf0jZTjlVunT1RVmphmVQ+q2
h6Vzlj/4Lp9152IXFPWaAJX0YjcyORqKCTd1jYgqvaOcb4mcY6ZluuQCHL9xh4SGRKcHJGPHHpsR
sb033tvB9snb5Z2i4tTEzjStB9usFc74FmEKkHQLtIvOf9cLICKR5Av4E2JO60kkpn4ECNoKxVwx
7N+wKYPQSKOj2FMzA5VFZbUt/tfbzA253HqZfDNDF10BjmHfjHRm6EX2BYYLMPYxSyvJvRmSpvsS
3esJA6pgIaO8APHG4V+skVx2rdsayfxlcH3e5Ev8mrlZbr5jsCshZb7T9pcMrTc8gHg7UYe/Kjpd
GD/UeXcJJ1vj0orsn05c2fQOl62IkMe3pws9GB0eVe59BXg0yLYo1f1Mx0nGhbBvfYRjGER89TPk
3c69f4pFmtnZGHVRu5zj60gjKxfPDmUUvkJpiYvx+SdPinehqkC+Yy+Rp8rLL1gZb/FcZayFcdEa
WhpQdLfJZw20451W8xmOBf3byY4rJ9Japm0ei51v39KYOufjBdlou9YQ8t3ZGUqKmR/XxLNa+Ym/
3SGGNAkZnTr4DB2bealCYMuuzDFSlUP+DIa4qpa0+GzNuuTTQOAB4GxXypAU3/D0fQKBOyWDyDxy
oLgX2j3Raf7tMSWX58/RucHS46BVHnWB6ZdrfINk/VugC/13p7UjZX3kxdFiryAUaqhJu8X0SeIi
4QaQIKqXPHpZoNzjJBtFsE06dxjZM/fz0AoqoHCQhNFCyMuIY6IDpGwDdtRIAx/Z4h/HuneEcAnF
DnvSL5t0E63rEHRySsKIxje3HTXlle7Hfj1siEoWhdlDSrBlsm/fb+cuUwrfOZNsg40kRq3EE9D1
VZqyT8k0RQVZkD239vWpX+QpaQRBQDlHCqUkJ8gayKBVTlwYCxjuAWtI9PwT58xE8iaUViYE+Ret
3hRzC1mczusLVWbYNEQQcRBO/cyheNi3Hpd87ow+EEVD4EYAAQlHO6IGeLjXD9kG0xoXkYnAz8iR
dB+7TYLZU0qtoIz1y2g6Q0NG6KPZ3az2gEiqFynTvefnqAj7ykLuIXbCF3qOOu0bndc1qor5TpqU
O+bW9JTmgjogEa31S3SV+xh3M6VYKWD8cuUFjbvviMNAoLI2z9oYZJqTKdsvxtFPeFF8Ea76/pg8
Xu6THpgTn1NJEMtEdY67AuiofEBPYrgqoKhzmiaS8TVh1s5Nz2CFcTEyIxRisCqtsWmJbfziAHZK
2P58KqJYZT+khQPeVKwflHUxvOFiUdtN0A82S2mXJLQZCICkDQe/1a4s/DWyy5zAyLHoMTirK9ew
UD/rcxnwFplcriwkprzbnU6SUB0cY1Gl/nGhjb8EjZIcWYqxwun8yxTo3o1sFnEx3scScU1zCl2d
fgIZ6QHdq4A3PPehma+2g3sMfxxZOs5n5+zhFZggM0Hnx5Sb1jBo6mj8NCNyyDnlDG9AgMu5Sd39
yZur1zWVSSdAzqFRz1c5qnd4mX2ITHTHSIH2WLsGv+Z2lfFOnOK6iYTUlwTK84wz1vtrW7Y0KLdN
U0aME0jy99N2kwcOeKIEPWR6qbeeOlvt9tdKset1PsCVMUutd3dimcBNGHP8NPR5k5YakXkKgXlY
hZmlC0TO1iKt/CdN5sG9pFWDbf2eGv15DrciSrGzzZS6yML5yn9siPO9tCSUdaRdTKtvfHRuSSn4
zAVSJ2KYGTEhU84JnxfeUcwf6U3ZoHSLMR8yqe2fZvpvsBjF2WWAbqy3o6K0y1S0SV6bJypViOzr
Fs7W8FG7jpVt8mI9Ra18P8DeTbue4pSraecFbWanENS7lFo2X38sNwErtQ9eeoaCxl1CrOLLrB5e
Y85yVY1O0SjlP0HxbUW4JetXxa2+/vXj+Y5tgWpi0LVY6z0asNYWq7lPy/EkIY2oi8bF1CCy4Gs8
GqtJ3spoOUMd8ps4Lb3YqhIUkFbROV6Gm/k+fOUC/dDK5gb8WQ2mzd6c3IPsU91WcK7uHKFxLQBB
c1kpoccyAtEEKX1qME9+EdAOpMdiGKMc8fWgCG/dvTw4gihtVE7TL7AVTRM6gqdMHcN1V3gMv0tx
UkWtu89/omApz1kAF17W01Sy4VLjp8hMXtQ/Q/qlT2a8A4kRFZWj+57Xy+6gK1UV1GVpl98ck+1+
xPIBwiGzj3PCw5Khls38rsf3StrLudwnNiKUbQbttpz2W4OUIzzTh5nxEFetCriiKBEHidsapnP9
WSURjfugBIymq58wFRJeyXkyi2XTZtH75Rl4wI7947XAgrsIoBmIfm0e08OtWoung6iU+CqjqM7e
f4rlFJc/OEH7DIyf0g7Q2JpxzHN3EGT+J+7SHbPaneSxzgd0q6IwMIDwyuEDYS/4HF8VOa8c5D4/
9thB38jIdjsTlk8s3issqdYDDGo7OW/VYENVNHWKo6vWSdSkTT4SJwrg9MjyCRIHyHWtipUqfBsm
AarWdAnh831lZddQ5B2mN74rrJz+btPtIk1sG1vU/rpJT8zKLc0FVaTnsKr1z8WsGI92xhHqfx5Y
ajAZafveUiy+hWFcRy0HAF2gBX6iYY2eF+suGMw5rewKmopwFIz6ukKJKLFphe1c9+HmPjyvYjkd
lQv2BQ9ceGAKHcmisjfvLEo1EEgKUY7wFRZcvGUfKNltlAJ0b1QRnT8uHZjrn1jXth2Z0+nFvk6F
dPkrgANAQYzzJJx2KtM7r/aI3NLheuTeZvlLjUkCLpnyT1dS8w+kNgCQcz9XINmM5mRez1IB9Cc9
KMCIrJ8DPhFO+cIisArHF18zIdEFkcb2qMsw5YdV8VWvonokwleHXM1hYcqmUVGRdLg5YOrms0eE
DjphjeSEI3rzodhFO/S21n1ntKWGSKweKHum/1D7hjwAX1TK12mO595tj22+ZnCNnEAg6mgDb+W4
Q0VTZ1KHx0GyvcNDM/qwe/J4VQYkFEbOA5q8Pw12sc9xTTiMg28EznwjW62CQ0rOGAuey/4w1/Ht
2EuJn7bkBPiajQbHwTZwV7TS9sHccx3r0yBi2tkvAVlicOOLpkcsoYmzYjOrgZbdwAvhgsmSkUen
XpN19U1PHvwrAGQKo8pCX00HPxVnPenAHzc9kujs/ai6P+GX1697ABq03bgFVQfC0A1TS3txnFmd
IAo4u00YvkjcLFpoR+N5BkvePUSOfwSyDohUb5lQ58TxStn62z7LPqf+q2Ebh9IEWQlIUsH3BSZ6
5P5PaeYV7T456E3cS20QC6LZIGjGaj5lAi33yt98
`protect end_protected
