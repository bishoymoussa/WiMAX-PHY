��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$Rx�y�<��wA�*;�x���@�̦�W�X�fa�M-$u����n~�%���P�$��W��kYَ���P7�?UMfT��q�6�U��k�>����~�\N�(�����X�e���/6U|)�X2pF�]$h���d.���9E��WG��L�X"]�Ad����ľS���8od����e�GT?y	7�������ݵ�^��R�q^]�鍦�����s�ae���h��L��P_���ާ��YЭF���'\��68�b�[����w8�[X��V�F�0͘3����q諵�uW� �h�u\V�?@��_6G�_�*�G���B�絉�f������[�G��U&�����~�F��AׯK1�`c��[<��FY���4I� �#�G��x[X�=�Q1��`��R>(�w����R�O�?����7�,(�H\�#h(W�EH=�������yq��Ѿ��aF����:�U~m<|��.��0=�P/���4ǆ���T(����ɷ\�.~Z���a�L�)&i��S��tߣ�V���7����Zؽ��l��?��;A�&�9�(F��V��]\�渫�s,eJ�x�A OMh��˧��KZ󋼀�v�mi(\����t�Z����H�C�H�������`��L��6��Ł����2V?Y�+��6�_:�Ĳ�бr�� k`h���9G��Z��lU;�N���5����a|_�ɍ�%�H��B�+y�%ţmf�t�Y�"f�b�2�yZ��Π�k�6g����>���x�$��!�S���n)��#G�T������9��dl&;K��?|��������&9�{���BXT�ۻ�{��	����<x�g��� �����ߦ��,:6��HQH9f$��~��k<4U�Q�a2e��	0�s���ZF-lq7���[HYMx-,q;uct���t�ʒ �;v�:��Ĺ}HƘ7~hI_++>���!C�e�(�SK�{�QR�y���"�0U�8S�[ȉ�T�|��62V��3�84�D��E-X׉��p���Th�b.�==)��m"%�	��.K��J�$n��<�~���{������^��j�kkrV8�V���n�M����t:`�'�肻� �c���h%B��V�ޯ��8䰈�e����k`�'o~k��Z��'�G������D�����]]���6�ƩWc�Y�ǫ�����L�X��H9�_���'��@��_m)��	tG�ܓ�;��
���ӻ$��)�l8\yz��<�<~�Q�*/��5ku�b���5㛢%X����[��u��(��X&"�����Ѻ<E|�wS��6�U3��7Uv�*�s9虖/�[g�SL~^R%c����V ��V�\���^%3����r &�y@5]\R�9�����>W��p���c��8�1��$mPT�u��o�_�A�6�r�^x[�ld�Z}jXn;c��.�:��?��E֏���ؙ�,� �x�d����l|�\ND�Ija��@�xE���_�w�w���p��pE�Nއ���UpU��B[��	<�ˎ;�*���(Q�̻+%�U��9����?V�W-��Q�"c�fD��.[����,|�=�4�u>]^g����TXhn�	��Zpa�� P��ڒ�'��G��ѝ�hK���=}BV��%�y�^���t�ڹ��݆9��6ձ���[f��Y#����A���ڙ
�R+�+d�ExzL�B|��P/����E��84�xY�F������X9� ��6V�"������g�y��|��^z���)�*�,���&Qot(�u`��FT���E>���n���b�	��U���G]j�#��I�v;&h�R��Eڣ�Ͷ#��A�G�x	5��}��f.~ 7�I��-P�E"b�q��yV6�i�w��Α[?j���M���jY���5V�i�kG�v2��#B|'(i�&��D�ڣ����1�-�ۧk��)01��L��=oh��%�3`�I�|��� R��3�S�gف|T~���d�S�f����ȑB���ߋ��ʱs��9�ҫӋ@P:A��[c��8���q�1��@}c�m�K��.�:X��Zv"��uU������5����\H�թR]�f]���r� ۤ�5$xQ�z�>�~�藲��u"y�R0��{�i��B��N{��`�Lhu�� ��
�m���D�H�Q���u;ɢfB��$C�4�V�h������Eۤ����gP;����(&n�v���ZC�J9�vd��+jZ����q+���KQ����tj�nW��ӧVly"Uc��Hne'��<�A8:�:@�{�亣��j�j7Y�4�E���߻�sL��h���}؈����i-D��hŃ���T��#��K(���Ņ��yG�|Mˎv��1_Y�7�,��'�G`�F�t���!��;7���9OR��|l�>�Bw��E���z�u�6Q?���'g���eb852�Ż���ѻ/#~A�Raa1s{$�K�����jM��J6|fB�鿵�Jm�u�c�K���r�gJ%o�8[zz����v!�ѓ���qi׍V�Q�89��g��$2�i��i܋�o)?���O�%G3oA���V��f=4�����$��?��}��=F�Y�Fqf�����e�(P,�E�[L�rv�-���ֹ�Z�=�6OU��dܪ-(5}}��!�_�$�.�l�X40L����:qINq�A����)�;�J��n�4 O���G�e��UD��x'u�̱B���V�aL5T����G���r�Bc�/�2��HW~��^&�Eʡ7o��G��y��������!bN����;h�� F������聘�;��1C�8�dT�$J�ye�䢚u�H�FYd��� ʿm�^���K��Z���A\S"�6海^�a� �����|.�g4*D�]@�������:��%� n3#^�`P�8	FT X˅��|@&��i�ݘw��'YZK�Z�ͤ�a����ي��gA�Ŋ�oV{Y4�Ku����u�T�H������W<���1fp�\�~�x/��^��`.l�������f�)Gt�՜��h@��9��E������X�Z,�l�J�t�ci�w��6�)�rdx����y�? e����XIH�h7�	�ʦ/K��eq�|DWg.-Ĝ��a��Dh �� 	W�4 �ፍ8a��h�Nq�4�k����"�2��,��Ϝpmk�i�5���w�q�ZT;ҟ�2qug��Ιh[�>-�!�� ��a7��t]ܿy��]�s������}&����E4!?���0C��+���+�������7z�l��;��4��������T�O��[S���ǟO&�Qn^S�+���N�2�鿈U#�*��h�N6�"R�àw�Qȿ���&�͐��6�~����E��fcb#0��woQ)��S�Kg���r�#	~e��"sV�.��@�ke62dP�%'����[�D�[sb� �1��iJ5��tl���o	�����KZzMid0��nvl�����>%��UX����^�����Tl�<N�2�l��n��F>�1��ȿ��;�q�]���aR�c�"�1)xjS���1oi���]Z��|7�2��O2L04}����N�3�#x,��2>����8���)��|�Sq���{��=��C�
6������o<r�B��4��\S6�I�Ԯ��
�����x�=�#y	�wr�vhs���CTxBү�	L��*r���p*�lt�B{#q1�Ŕy�6�~(�bfqK���[ �{��}nB���($�VɊ"��[�?GS��>l�K��r��Ud�<Ǥ$�!$���eB�kmE{����^������&<�qC���#�[�_T9��V|v�Y���v�׆��c"0���MzJ9*t0 -��OD�p�a��=e�ں��E��}#��rU�ߣU{}%�Dбe�r5��f�x�,��@>D8��|�����Z:f#����^ner���ew9�}�Z6	�O�N�4陨6�@iP�럖#��'�{�$^᷵MxJ����6�ݛ��Q�_�t��r/1�~���@X��s��Y����犖o�OgN��gI�L��������`>��"�bhj�w+�K����Q��K�d�H�t�!�%N��ޔ���#lpW�%;�����:�ddÜ�A ��A��$N7P�O7�M�����qaj�[󸜔y�n�O�U=��,��|�>b
�YŐ����C����^��x�0Cϒ��dJm`*��"$S�(�ү6V9ĀPio���M�A�oHb�M��W�q�d�p�����^1j}ѧ�;0Q�QiCW��%�a���ӌ��(��U�XlT�g�ۈ����I/���Ba�M�ڽj6��b�lԑߊ���J �׫��U@M��_1xp�ߣ���,`v�Bbe Ɛ2_�y����|�)V�`����[�r��h��h��B�V�p��G��0�[V(E�v�*���+�v�0�כ���)���v�T��Sy�c�hmUe]�R���)y���H�te�P�m�_�y�����%`�8�N�ӕO"�s��\��KԲ/�il~�_s��݁���y���|��� (X�J��ˋ&��*�Ķ[�v���<��h�D�鰗�W�>�.#!���yDQ/r�z6P%���l����%]$�LK<MN�\&�Ce�D�L6yH=1E���Cf&;>-p��ۧy9j�O��:T騨Mݢk�1T&p!Qɀ� �utNS�6��\���2ҁ\��?�i��k�ӣ�4(�p��25�yZ��YOB�`k���kQ狛sz<xB�U�p}�����M]@���u.�s�Ej/�?`_A�i�%6S�0 ��p%Y�'ol�.���X(Ȋ,t�~�@��=;KH;�g��^����s��$�����L���8��V<�M�#@�5z8MS�9�z,F0U���c6�{��:8�w�����w�I���ml�Mi��n`�
ZŤ"�(�A�A�m��R��9dli[�7�*�\c�]�p�Nv�&u��=�%��d�M{_1��<�>nO@F�%�'k��ڞ�y��F��9�Z��������ǁ�'ss��;�.�=�EX��ݠk�B��Jk����v�� ��YZ�`%���-ngTvA�
q�E�ߍ$�͌�����6�,K��7����X�O���x,M�P�GF��)��n�aX���\����R�>G9hl`�4�|k��$xe{���;w�I����x:�j���lm��+����'���� &�F�F��C��yۦ]�_��@z,��*��Dq+��L-o��BxL� ,�l����s�<�99{�93�᫒�EN�{���uP$�<*ilP��Pc��W���T��m��i�5F����A
l�W�j~1�,�2�L�=�Հ��{~%z��T��r�Iq��"[6��=B �?}w���󆄪E����4��m��g-Q:���y���
�%a�KŞ(�	�H�;�l��,����қG@��p'|�Gs� zv*������`e�#)�3J_U���q�������!վ��&HBM���8��&�9q�����V[ɜ��|��8�o��1�L
�n:�+	#q.�_Su������X����Xg=Bud\Q[w��`����Ҷ]��!�7!LXq����7~x�i�T:IE���ea&,.�4`���4b��4U�B�9@��A�ӳ�h��t��l���&n>�� ��o��1%�?�p��j-��z{1�s���w��~�㳟j�_d�L�R������Ur�y-5_��N�����3��43���l��l(eȭ��ﴐ�\���ܲ��lv���l���l);�U?FG4�G���h.>ZPaY$T�|ܐ_�:Y��<b]���o�,	w�4/�gX�F��$E�-7�k���Ǳ3�~���5�߾���@��@պ�r�P\����(MJ�*0���Uo"�0L+�ܡ��7�e Eׂ��\�C޹	]X��JA��BIU)y�-#䢙'�I^�_�]l�T�Y������O�������m���sH��ZpK�G��6�ᎩzD%{yD�� ���g_Ь^n���o����N;j�?+������"��)��,x���j�F��G�P��_;��v�M���r>��M��ښ��p�v�3��%����_�3D0�m�ZOfp�9������F�|��r�	�$�w����n���X�% {�j��~�8�[��k��SPM8����r�^Uoj���b��y�BL+t2�wҮ����U����n*�>v��d �5U��R��f�R?v���"�<���m�<�͠u���5">��x4�bbO!EJ��p���j#g" h�4E}�b!�UU�a�~��H����`����8�a�@;T��[DPı6���"껀U��2C����ȹP�j��#�/�i�0l��o�ќ'�{� ȗl��ȕ�O	�)�QE�6B� �d �^�w-?������G��hZ�����aP;��ם����t���#�Z�s���c���Wf�P/{��7l;�i)B�D֛�úr���}�m'��w�#�ʒU�%ϞI"�n(8�[t̙}C�����ș.0a�t��*�������W+��i�d� )aH��T`A�#���F��� �=o����כ� �@� �,�~��,��(�fvH/��!��e��$�E��]ǳ	�p����o~��'��¡��'V����os�1L��d3���"�lC����B��b>B 44{��v[�+��2V�kQp8O����l���ڌ�˺�V:���!�L/�:6i$���!��KO�T��s=�r|#����mo��ܘy� ��#ŵ�$N�(uk"+=|+���F�ԦA^�l�yif2-�>�� /p����,{�EF���P0����g�b�������z��¹�VB� ���M�1<���eT�%��vh����N��Z�݇J?�:��)�N{M�����(��|��w�pj�&⭨����.��?2�=�pAHa��K��2í� L4�'�~�G�S�>��
DOf}��\�0����}�W7�d��3}�d�+�`XZ@���*��r������,�x��uz�Ʊaٯx���	(z\�,�3%e#z����׿������y�y�j����P�۹H/*J�֖�SS��̮%o�����>}�IP�a�vYu7�� ��b�Q�wR�NR�F� t�$�$S� ztw~+���o�r!�L�1Z亲U]se�bH�����4d�k˘��A�z,� �3�F�5�V���d��e޳�;�G.���i�Y�t�G�	�Jx6�D]3�"NL��o�MR�J<��XP�?� ��ܬ�t�?'&�ݴ�>[�/6@JL��z�ѓ $:��)j�u�!�ֳ@	�F>�Q\���.�f���J�M���,��*�0>߈L��Ec�oϘ#^�v�[/���s>J�}�����rs�[�n�p��%o�w�k����ਾ�W'&|%L0F�����b���y�	~�g�l�N����<�$[F:�DVpG�V%��K�ɓ��[?U��R��M����}���;����[hzH�a]��]��ޱ@�#�4�@����٭�5�g��2:G���5����X��A� �a���Z�L�7)�`u��yF��X9��r;	�.v�-,��_]��qf����KcB�*3��aԻ��C��9�8��WU��0P�<}��\=��)�K*�m%��V��o!sÁ��R�&"ez�*)�Y'l���yw����5�Y�6�A"]�-�1(׾��{N��`ю��O��q��ON��+?ϟ��\���=+��Քƹ r�R�eũ���JN�|k������#"�A��x�2+��������t7��hj[O�zDÆG��<��w>�|�I�CR����_�	��T�9˶�s���?K�� �K%V϶�aـ��S���>�(�H�lO���s����RC:�����D��J����$�@��T�P����?K����n���y�^M;9�ȟ��?���j���E�)?L����eڙJx%i��dl�z������Z��� 3��Cs1}*~�r1���{��4K���]���uÿ�RB���52��R���C[.��m:��pl�?�U�#����&��:��W��M�VgO�;e��\�M��Ll�n�X��	�ő��؍'���UlfV!���nο�3�W�J��n����tԠj],6N��t�p��-��ʋ�4|�+p�����m�Bޡ˛��8�=G\l��C�(�+wl���C������P����P~'�ҜKƊ��XP���4�.Of,9����0�矞�JpeBh\��ݝ{��L���b�����2�n�[��ƴTf�$4κ�O�9D��Z��S_/�Y�k/�9���F�Fl���_XN�����Y��ظ頻&F���/��t�Os��m����o�;tͬ���W���)��/6]�s��]�)ٰiU��SL}4���}3t-ܥ�<&ҼKThhi�(�\��_ū���L�@�=ĄÍ��TJ8��������!Sg�Y�L-��%�.�iv<�rb�����i�
Y�d��Z��dA~�&�@�kmQ@ ��}����b{¹�v#t�q?Td��B��OHQ��25��<�t�t�F��w��jZ{��FE+4�7�X�Q�d�2�0�`J����� ��ҩ�V4�z�c�AIjk�7
�W"�4�ߺ� �F��%�֚HbAԠpH�G�uA+�F�_�YN⇦$<j�Q�	h�_�-l���*F�쯛�ж��P�f�[��c>UW����a�T��س30�aƦ	ʝɽ�*+,�'��veh��"���� ��J���}���ܕ*C瘻�їI� >%|'��������KZ^���Wk�[��;=K���_�f��w���z��?u/:�,pK:���Y�+����;�8Ϩ�S�":�2W�q�Q�JT~:JN�o@�[��Rk���K���ÿ4r�t�qP��">�/i��2Į�$}���H+C1I,�S7�f8�������c�`.�O�)dG9�:o���p�#y)Ԁ�;�~,Vzxz���(܁�<�q��I���
Ұ�Tg�M2�3~�ߖ�m������ڦ\b!�jt�?b��|��	��wҾ���'�z�B�j��i�*'���$=�����0�~M	�0����H��0�ד�\�'��}��9v4��G�"5�{I��.��h#$g���+!}�_�d;DA�m��Re=!4z@�#:p�;*��~���������dbS��:��T�
<��>1KdXH�%�ХJ���J�i�QY\��pZ��}y�1��������%��O�ӎ`��:���K�C~�Y��~�W��4��)�08�g=�P.ԇJ���ܼ4�g3���!�-�_X!�w@OH�����5�u�n��~"�ץ� �\�(�x\q��;@@�Ř�4 �'���W�]7�gJ�η�g�/���;�3V�l�����t[��"qm�qk�����u�\b�0j�]g#(�<�* eO'U��,�y�XA*�J�PZ�F�����4kW�b��Z�'�\�D��hƓ�+��*��s��P��J[uŮ�}�c��:��	}xF�v���ڢ�a��ز��1�7��ij�b�����G|�� � �6ۤ6��9�۪ ��jǗ�!��`|Jm!��h��r�I嬏a	�0�>+�3)8�4[�A����4��'�Q���b%�C�Q�[ ����K�SD*�V8�1�W��m7��)o�@�:S��������~����*yҁ�t>�({ ���&�{^��2٢�:���+��_��(,��a��Z�������5+J��Z畽r�o��l�S�䕿�BiU�9�6lԫ�?��x'���͕�5�����x��M�<E3#�O��`59�O#�����ۻ���3V���1x�������ҚC�c�➑�n��/�����OP��&��� ��D��"0�_��(�;���	tE?�^���1.g G����^�F�y����.=/m����|�2�:/��v��D��o�L&!K��A���;��Nں�ab��&{/_�/zW��!�?O��7=���-U��P>U�u$���h�\����{7N�vN�[e1��*�X���ZO/%*�&m@X�����Z}�� nf��q����Gv�yW\#S�iE=N��?鮲6�`{3Ɔ�(����jGc�U��P��v�heW�H�'@)`���f1�9[s���ި;�=�@���lA�ɚL���%$���[�KQ�)�}���b:����nc`"wn�rs�`:�Wm�'s���ҹj�	�|�A,o�=��#�t~=myn�w�(����-G��f£s1�#m�~�:�;,�r�"	�[��*�M߳E����~KNI¡5�u��{b���v��
3	���j���8#�"���TG�Hb,�Xjmib{e �=�
�S0Ensf�$9�>�if򏜋	֞�;@BHÆs1'c$��&�$��������ѩǈ�+����<!&Ɂ[xǭc|䪎����b׭F����&̓|3� T��%r�φ靉�EHT�c~�Y%:M��G:[���Y~#'�6L��`K,adD[��� 3��A��������(ِ�n��Y��od�w;�[Z��:��FZ/+��������*
�֐�l�-�?��3���Igj����o�^Q��fR����m���m[��4#@�ZIb�Ƭ�ۦ�٫q��y�k����-�B�1m���L�����h�c��^4� ֌W�o2�?SJ�2%�i�|&�ИT�:޳<,� V�;>6�T�?v5y����J�����m�y�'�0���Q�D=N{������F�I�A��떜�[T���0�
� V܀7��ҐY�*�毘dsҋ�=�.���`i�Cr��`�TM�	;��k�����]�	!;�������$}9Y���V�*��q0U�7����m�7NE���-�Q�ͯ/X�A�_j�\r��{��Q����D0\�9�U5�A�ڛ11\�ҥy1Wm�X�B���D���[���+i]2Q�'�81~K^�:�d�׋#b?ѝ���)��zFd��73�i��2Tl��J��R3��x���|�Mٿ?B�u[C�E��R�*H�6L%����&��]�ꞆQ�`����8�!Au��Zn~n�z�����X�� H��S�庖 D���B�P���%9�b���47$オj�h�u�N��;�����������������." �Jr�]xk�>�eI�o�5g^�S�#�Nw �l n�-��*]]}t7�F..���>�<P���-bD����H����O{@��\�@�O+��Hk�I]|�]�o�8-� =�gV-��C����q½��M�:
���o><�=<�"�/����c����D��Ҽ�o���<W�pz�(�Pt��E̞��zk�r�(u�k�ȧ�m�����/^L~��`��*���#)=ˆ�qt��Q��%����
�ؖ�,�`��iU�+|\ <�vH4�4�`b�����#�F`&r
4��<��S՚/ƭN�g�+	dǉV��Nx��&�t�Qv��)p�,��}>����ig"�?�D?�`�~�C�2i�rxQw�������5��B��\�S_���$&� Q/����MU��_��� �Q׵a�K��^D! t5�
��q��'��S�H���b9���0*�������~5br>�ậ��y^�I�v�Nh`v�w�ˈ����@;
{�Zk6	�"�xR��x�(��񵤨_�<g?+-���H�PU���|mZS�{��$�C�eMݹ�[@�ȯ�OCx"�
�fW� �b0��J��d���✺�1XTat�ϮY�&B�'����$ڷx.V3�E�����E�6�!�"��*�*�(�j�(f�TW�߫���@R��P6��+�cIc	M��Wq%�R� (l��ݒ��[��Dc��܍S�L/<�\g;�W0W_`,����.g# \��6��Jn���c}�	H`d�fm�,ڡ2(�o�I_`,q�]�H�M Qu ��q��#������h��2�Vl�������o��ߖ�7A�_x�~���;������l���qY���}�����t|��h�� 9���ϸ��3��vc��oQ�]������uw�F�ωR�M��ˏ&�An�̏�sA�J�q�<u}q�Z�|mݪ��rk��T����3<��qJ��d�ĩ�n�$U����h��N6��0ws2����(�� {r��ATNy�D��&��L�LA�+8��T@j;-_wD�>2!��4�Ϋ��XZD7�+ω��&.3o�-_:4L0e�����J�/潋7�����"��<�Y�4 c='��,U[lh��޴�#�@V������t�Z��
�7@�a�C����_{�LJ�c����T}V�7?J�kh����� �5�ȼAVc���ґs��I%�t�B�|'�8�&�b���Ϩ��E/��>	��bqM �����Ws]v�,�Ī���8�I��3�v����>�1n�)Ni	d��y��k32�d��=B��xo�;�/N�؟��pn���_��%�+Tĳ(�I{0c�!�5���j�P%�7F,	�	0�3Gy(��g��X���|��t�]¸�M���P�wfAu[�����G���JÑ�%g���	�JWEǩ8�!ܶ��tA��ۍd�r�&�2��m����ʩ�B��,"Uّe���c�fl*��р��[�������`'�+�r"p�s�>��I�^k�X�( A�3�{��?γ80��G#��t%vM�JR�|e?4�RQ��K�oYm)�U[V"���u������ꛭC�g���NmC���"��Ʊ.N�WP��T0vص@	�ʈ�6"W�"�h�t�џ���u��~�^m��xɐ�̍���K�3��֓�=�]}�����1,�&���V[^;����� ��y���	��`p		�j�N�2���CR�e��ޤ]�z=�e:��^U�vg9�s;�e6*�jk'e���Ѕ�����G����r�-n�7L��@��T|�Hd
�A��j7\����HH��gÓ���+����{fŁ�EW��)���Ig�~���K���P:��w�G�,zK����Yt7aH�����B�-�C���p���t�,J��L�i;UE6`��xj�)�-�[c�s�	���E��G��}{�_��ŝ ��:�����j�(��϶�h�?���lei��'B�hXqp"���
��W���S�1��c4_!�@*�F��wk� ��"U��-�.m��w�X��ܼJ���`ñ*�C9,�P\t�0?���I���;��������������������L%�^��a���7���X��|5+;o8��ܞ�j���7��p�aR |��>�3���t[]���4�>�(��󽌙cp��`4��K�p�b|��m6�|K:j�31���T���gpu��6�^I���ec�#�'�v��H�^��g�2I18�n�����Lzo��e����G]��ό�~|��כ2��Xv��>��
���M�
֡���\H��_\��HFrƴ�?��f6�\.�E~Q߷>!$�[��3(M�Aӫ5\:Hg��8x��0�_�9�u� ׍Nm�?I�<݁���L��Y	d9��	ϏG{��6ɰzb�$J"���f
��{%ǫ����"�j�o�{�Ds�mx
�a� :=ˏ���d�jj�ו�g�M~��C0k03�S�˓�e����m���ѡ��2m<�����6���!S�w���%���.kת `ײH9Ps��y�k~/�:@p8[��6	@_�k< AI&��B�mp?��}��Pr/v5�.�.��A;o%�v/[�2IV�fI��5p��}�4f&��KȌOHj��>�`?`����\O����0���2��(�y)e�Sqɏ�Iq$�p6�f\dz���&�_���я�)Z�x@Os@ùz£Z����P��|B�)^�S��<"Rs���E����&��6��Ht<�+��Pe�|��z��Q�c�����X�����^k�C�6[O;�o< c\
�� �!�G�}�6ů��.^hIVOK�*�U�S��h�j��u�.��;ܯ�^~��T�ia�F���;�����t��D5q�Kp�p �_�B�Z��&Q����J������x�n[�?ya'xZ�y��|9��6�JŹik�kJܵ�!�/�S@>X�TrX�W������`ӻ�[q(?"��f�1[���F9��������@6�s0J&h(הxBk��dg<z�=C� |��6&̟�2/7>�p�h$��[G7P+�J�6Tؾ�g'�n7W����8x���?�Vx��p�7�ﯪ=Y�eAJ�;����t(��9��^a�"�ɞSbO��U���y�M٨�Ywg6�K��H���0�PI;���o�od��Y�0�K��G����T׾9�#l�%��d\\��rͿ�?�P�sTV��f���3;>K�]-����R��K
`��0v��j���.ò�a�i4�-
��U:�F�m�Fs�z>~�gV5Ms:SZ1XqY�ed�c�{�r��D��rDF"ų�V~x!~Ώ���6)2{�gw��u	�ev�]g��:�R�H�yØf�~�8��(��T�!1��X��![	��X;퓪Y�����JQj�p-�-<���8�/��Z_�W����铑KЕCv��-�1X���po�M���?���E�Z��r?�Q��a~Rl�ڪ���L�kfsw
:}[���NO�?��~���ptC!��wE2�'�>�&�3�N�����H���\�����y�W}�l�n�Xr;��"�ۣr���v���Z���,mN��6���%u�&�L�3���9�pڂ�p�`'�(���@&��㟦�-%��uȾ�OAS������J���S�#�Ɯ�rԓ�eF��n� sU*f���a�����/y����ۧ�Q'��NԈ��"��I�*����������������u%8>Td�o/z
\1�d��q��)}�4��9%�v�o���ȣ	�A9�����B�i�5����'#p�n�Q���ٛj\�h�T7��P!sGN��I쩩k�	l#����5R�q�$�����8�W�����0jm9)��[@2�}������͑L�.ֵ��Z���<GvEn�i�L:_Y��^����E9���Ԧ�~�hz�z#53��P0��-&q_p=NHK��I�i$�R�l��;@� )�)�&3��g�c
썅uU�7��܉���j�"�*�����u�-�;��t��p�B�hb�ٱ����qxJ9��)�e�b�����$��0�l�ZX�蓶-0sRa�Z�|jJ��mHڼ�e�e�N��պ��68-�+�C �_�
D<����Cp@J�ժ�l3����w>��������aX�/�Ub*`O����&�Q����Vc.�˼-|��e�����'�5�u/�c�����M!?����Eɀ>�����,΃�n^�^����B�����ve0��ɖ%��`��������=z\O�b��-�ݰh�ب�+A�ĝԍ�d`Ă���>aj�Bx�[Ƅ���6�MY&�^����&�ٳ�\Zk��O��!�oZ��3��Y��u�8��*������О,9�����n��&���*�얦^Z�n$״ƞ!�F)Vߠn�r�^�>\>���v�b)�Ԋ�����I� 9t3s�A$���'jm2g삾�dr�6<��77Wo�ʒp'�l�j��u�Ub6��ֿ�X�I�\����gi?�I#�Q�J��իK�F�rc��gλ���H���u�V�� ���`�"���o����Pe�2������#��K�֘t�a�:j�#�V�l��x\ϝbl)I�u���o*Aab���cs��U��2�0ѯ��$�����J5X@;C�Ŏww�R��XщҡOF��cu-n<���E6tS�W2:nh>/��LEE�O�� +�.��SlO_cc	��������ǑlT�(y4՜�^�x�ׄ�����>�s���xe���6�Ϙ�E ��d��.ѓ��F~�vB�*iἼN3�zؚ	lT���d���sێ~�%�	�DEu�O��+�4�,q|/�}�f�!����œ;̻�[btI(b��ɨ�5\�w��!^v@7-��>�:��GV<e��kr�$��Y��|�d�"'j�y��Ag��!,Nוʍ�� �g*�x��7|I֯"ہ����ϭM!A%�M��Xa�:��w���P���qg~���&¼�$5���:�o'�E��o_t)B��g`jĆ{~�O %TO&%�l�oŢր(��e���+����e�q�uT�Z;���?n|苴A{���9��$��3��e�(��pd>|�[׊�z�x�k��ij�-��6N�U%��v2�Iu- <4'�]�k��a7��|�|�9,LAJ���R\1�tH��ml�ӄ���>ta�������I�#��{�os3��f%s.	e^bm��ZW�Hl.��L&M�o=d5�wk��`!I�u�j�̅�W*_�ɋ�p�\�g��	Jc"���g`���ΧK��e�yq����V��z�FG����f��������Y�"�:�X��L�\�
�8xoҙr���q����	KW`Gzy�M���>�FY*��E?���|S�}_ڕpD�:�.�_kH���w�K�ʃ�F����D>B�ވ#u{��9
y��<��@<����vԆ��#���ʉ7�)z�[���D�U������Θ:P��?	ѴN���g,����n2o價�w���k��
�VB���r�=�z�ʽ`��Uy8�z�v�d�b1��)7EC�M=��^� �g�Kh>�{���Q+
&a��/���ӫJ��Fu%Jo1o,��y�ӽ$o�5Fq�Y��нi��j����G���y	��#��ui��������A�K
��%{��Ȃ�V��E5x3��\��#�n��c?�G=Rc�6�Z�B� �te�t[���>(S����WW�Q����[OB�:ؚa��B
�x�9<N�8�'��Ɣ�N̍^��Þա�>LcZ��C �!2 Yo�#Л^?��r��;��wJ� �d��g����M��*��J�5�|}-b�hk���E|��� �r��l��s�Jb̢�wo��{pw�O�<2/�Z�����ە��g��%ў�nR$kB���z[]��r�>>���q�����mY�{�:����]�p�L�#��j�!q�c]ڴa�����Dy���Ps.r��T��}�:5�:V�������ct��
��ꍦc���%."�r`"�����T�Գ�m�Fl,�]�$. "��O-~�>�LJ���"�g�u����%��������`X��-f�E�ef�a lR0jӂ�O�t����r
oI���W��.y4ǳݢ�K��n�HMzY�81���s��g�Cye(|9���Y���.��� ��`����㱜�����,[����~-nn��7O�n�m\�=j�z�c����^�{����S�վ��J�ڋf/݀\̬n�q<�w��b `Ъـ|}r�G	`^��u�.���[b,��'P�$kF*���g�'���Jt)mi>���r���oi2����s��>4�=D^�� ы6'.E5�K��^��`��;�u\�n���A�V�T�8����u�~��ק���K<\�뿏��_�*��tQ������Ӎ)�r���{�� 78TƬAU�_�Dc�8��v���q���D�c{k|�]˄�� Au��2џ5D���	j�y��Q��1��ֹgE	bD��\3�#�/2Ϊ�K��~�egx01P�qD\ɢ��=�B�ނ�S�1c�1�V5�tY��H�Y��z��[�l^���S-��=�'�C�����T��z�UH�`zSYU9lw��fE���Qg+�ORY�qpDx�Pk��8����'k�ghh�cs2ƪJ��%�4���;( �e��D��c�'{�2	���5F\	j�<ad�2qpI��%J�wKc+��d�*�3(�r�8W��^�tq��{�9�N[����>�DM�IB����G�U��|�V�����Xl�>D���_����g�)q�uS)~���g������C���������%�OJ���a�0@��yo�<��b=�>��>E<��=���v�N}凉.YD�����u��3k�1 �|i3R��Ͼ�eέ��%���V<��s�N�*��c�����������JQ��乂h�k�NK�P��GY��n{�&��-�I}a�e��..��^�������P�2#�?θ/��K��v�����Cz�k�
Xݓ{$f<�*��&�Y�3T������e��
Xe�'���n1)*ɡ_-�/,�T���K��/� �須�-?��!E3�\��vǇ9K�k�>���� �L(�!�:)�;�!���q�5Y�,����
��(J����Xs8�R?��NT�u�Gǳ"=8W�L��֠��i*��Oy��7����Ui��^j���~�LɊg��fk��w$F��G��~��	̘�jǫL��N��vJz��/�_�mJ�Z/�Ra�a�h7H�b���L�I��s.Z���.��D�u��!Bv$1�Y4N;R�6O��{
���S���~D-�E��4 �uG�}�].��\u/��ES2٠�Si�Lkя.,{Q��P���:��.G�:��������%�@��&i
��g�e�<���6y�n�"�R>�(Z"��Z��[YW$�5~YC�˚|��\�$�Q���s�=����l��r0�v�&���b&����K'�SR���4[���N������Y��}���!�Ո/�+��O,��j��c*ⷺ�lP���:���'t������D.
�o<%.y�7���i (-]���H��+<?3�
��9�=�<ʏ(��]0�1���Ⱥ^!��r�J�B$�$ͅ�n<@@[�$�FxT;��P���>�H(�������}R�`t��=�I����=15���������	i ����|���㑊$,A�2!a"���G��U���r:ż�э���2-cD�P�O�Oڝ)�f'�K~Z��R5L`�yU������x\� ��<
������̐��/@�r�踉�m��˱Q�����w� O^蛭��h�E��Lt���e�)�ݷ�������·�2.�����6_Z�ƄDb���Y�nLC�Ɔt_���y�������aPJ���N`�M������O�=��2�.hcU�L���Z�����C`�r\D�9)����p�p�bZR��B��v7���������x�鄍[fv��JMf�(瀙j\^Ŭ�\��dk����="��Xe,b����uj��].}bb�l�9��'�M��Т/o �}�H1�^����� �x�ob,j�1���<Rb� �����AC�w�^˿0!�q�ڋ&�&[�UcG��-T��q?�xS2�1Q���E"��k,��.ф�oS0Y�\u������Yo����ُ��ϛ�r�n���=3�v=�w�i?j��A���Y4�_hweCI���^��ĩ����c ��=���7O���.[�G{�u��.�F�G�M��2���Y�G/ H�rg�|�T-���J� _�K%���j��9;�N�Q�F ���%6�^�.d<�����B�щXw�1=��2u�����뉄R��/'%�y?ݘ��|]ܜ ��m� &(�'\Ӻ{W���r,�P��'�5�~���q!�����ߢ&,k��B)�=j>���
)�no�!��)M������̨x2�;��'�"�%���&|�x���⑛8ŪZt]�E�u.������Ŀ�V�8�
Br@9H��W��ܞ�ip�L4n�&���C䡂aV{��՜ݷ"�v_#!�j&F�M�K5uĨ~i$g��0:nY��FC��f��\7ͨ˻jcW��Q���\�����e��6@V�mj�+Yy��l�IH���}-@.Ca[�l�gp� XhC��4�|JNr=x���;��L&O �H���`3N�`)�#��hEN�1��Lzv]�;���G�V�U�$9И��^�k|���Öt�u�=�p��N-v�	�r��.R��П7�Mx로n�
������Q	PH���-#7�����Y$r^3Gb�-���.T`�畩ӷ|mFUI���S}w^К�l��'�!-����"�y��H=��\�gu+��Wq�
?խw�&�#��R�jk���K��x��0c�{F�0K@i��gT����u���<��	bo�Wѐa��[�Y�R����m�,N%Sb;��'rO����l�.�|��Fu�uy��E���<���+��A>ƈ�e�Y���'4���
ȻMn���uo�� _	�*�ȷjl
������=��x����:������	ɑ����w�:m45<��������(���KV( ��S�	Ս�o�ѷ�GMxq�\�h/�L��8�M.9	[��B ��0�"�f`�������u5t;�+��/i�9��Y}�/���xM�k�ARS'��W=`�n�d������$�޹+TцQ�9��Xw�2��	fA��:���d��Lj&��&A��-����v#�B/��$��g`�{����/�U�0cM�"_�͓�)K�Q�F�c�а%u��n����~�$Ď��U5�(�]�Y�|��
��>�~pZx��2>��/��%��EM	����i*ay�������!Y��_����1���u��q�Xpu�Ow�O�z�I�E�xe�6D����=dxhپGж��Z�\L��f��_�8�k~��C����(!�.�u�QM�H���{� �C����i�"k�R�X]��aA�5��Ki4���>�Ɖ:D��-��8��DM��Hw%�J�F{>�v�*g}6n���ɀQU�[5qxIԇ%q���2�Y���v����c��=��ƛ��7�B�[դ䱣�H�����
��T_��A���'�%�=s�7uZBp�v�	w� �%҄�J�{�M���h����3�5>w���N�k8RNUjHٳ=��A�]A��ᯫ�?�I7�K�$�`���v�=Z�3}x�d�.|�I���#�@��l8$�y(�f�9g�Ґh��A(�ڬ�e�����@x�b��J�y���в��(4CY�	s-�X�Vv	A�����\��=#�Eޒ���]�о3�=f�Y����އ�	�Oit�m�b9>=@`Häңyؑ3\��.��i�!��l���K���xծ�#�p1�yM	��$*aC� � u'��	ɑ���$��恓N|g[##Bڀ-�h0�ն7h��=��j��j�6o��4D�]������;��4r	��\w]�����U~f��,]\a�@B��E l�r���@lQ�S�e�V�Q1@��/�H���G�/�I~q�T;'*aV�T��w��9Xp�c��+� ����v W���R����=0�F�b�G �D�e�.+F����@$=�fS��Z?�t�͍�E������Tt�O\�
����p�Vk���&���� �U�
c���6@h�f�>�,��	��u~���L­-kE�oy��u0f�ۙa�:t�p��@H������H�&�~b�4J��4p� ����͈x�0�.��K��h�>��l0	�s��W^��m��yA�8'�"%��n5e�m�E{����W����5���ڬ�W+�~�\�B¤�a�$�ME���a�/)>ė3|�Vj�G��������R<#|��9�ոn��j�[2*��;�uY�jnv	^��[�6��{X���2y��s[��~������2����7+���+��R:I���z*?U�,�p=Z�|1_�&V1���[չEX�x�P"�6�^�G]�p0����Z�1@`�\��[
cpEt
�ϭ'�h�%]g�Tߐ���e��G�p���[����	�����:K-1��T�nB%7�{M��"��x񱮽ٙRaz
�8�����y��� #<��Я3R~kq��̿M8.F�rF���r�\���}��3~�-��u�#r
'�?ݦ&@Wv����h1����`�j*�4Ub"�$8*�?=�� ���M�'�c)ް�-�@�i-$�U(t�e2�\f�����VJK���R�1�NoN�ޫ��H˒��t`�� ����R�v��L��r,�
�������<���^�K�$�4�>Z�7��$ �fI|^Y�k0u"����s���g^k��~�?���ފ�̤G}�r �;r�;�g��MN�@�򴴺����M��=�nW�cMR�H-��!S3��5�����̾V(>���
l;\ڦ���/��5������������ad�6XI�Lpi��l��i�^�m�h`g�<X��jDr�U`$O��$m��܎�qP��e,���LY�M�R�E�js4�[c� vخ����P���l`�h`�ȪI*4���,SHJ�V�	��1mCǝ�adEOb� e�����!�w�ŭ�~� ]W�/B���c���%�cc�ܯ���̷�X��P��\'|2����B7hn�ƹ6-�� ��W���=p��w��p�:g�����?�d_���<%qz⤞A�IY����'�����o��8�Ǖ/o��G��?�!��j�wD�շ6�^�qʷA��3b�����O
H�>	3�/�.���x��C�s�f���<g���a��NCbzˣ����k�bm�J�N�����?X�(>��jr)�MwSo̤nbf�6��ȇ3�w���S�C���?�1)�vk�j�t�:�%偙�&Ǒv�qG�'h��ݣss^%U��!VY޳D%Ϲ�o"�/pXD4�ܺ��B�9�)x�]~
�����N
#��-��M��Ǵ���t2"�����<��`�t���bnaq�w���׫Q�=��o7���q���D;�:> r���p�0UcG�[��u�-�5��?�m�5{2�F�|u��|��4y��J�2���-���q� P.żC)�D� $�O+��4�jR�)����Qs�������`by���ɚ	��ʀpav�X ��S�>�6H��NJ�zߣ�ưV^D�)�� ����,���\�FÙIE�=��CR6��6>dl���;��(�|YtB�u
7�Iu�ܮ�|I]���L&q��M���j*	[�)]��6.��������o�뷐[��Z⹊ց$:�!�v���I!v�\D�13�Ў���B�
�6�p�G��x������Sm�����q�b���]ȼ`�`U(��c�7�;��OPr�;5q�>�Oe�n��+٧i%��ڣ|\���Q��gJ�T]��oɨ�A�Z����n��ᯛ�d,��������\I���P3�mg����G�}��/"<#J��COm�R�j���H}&��=���z���~{���Z�9X��O��xR�M�����/�B�>r��<yr��Ñi�P���!'Rt��~<�E�s�Զ���L�r�x^d�<��������G��2OE#[%�6���E&o�N�'6�0��;\����ug�W7ٸ�Ў��I����tK�qF�Q>W����?�:8���,C���P=��IZ��L"�}����s@D��cAb���ȜTC�*--�h-e�ɋ����%�*ʹ�:="���';��
�p��|��A''�
�����"PH� FV�~'!�)�|e����HP���F�"9���?����7��`��qN��'��[	Q����K��%q��o(j�O��v�[&igR����N�U3R��ߙ0�'4K����o����2Y_M�պ��0��x>�<7��	��Y�=���o���{wh����<[���c��]�������
�r�����:e�~���К�9��	�}U�	 ������)�9	Q�=�j��~j&��9�[bH�!X�{؂��7�n����\��YE�^f[AzX�Tzć�-�轳��n:��ˤ�&H��5~ہ#���2��b�U�]z?^���<ALG��;��Q����=��*���o޸C��/0c���v����<���(3:�q4�!�l~��u�Nw�U�$&�);0q(�H������؈��g��8���<�)����Z*�(�-b�F|C��L�m�}`�̲��E`�O��z9
����c�� !��Dr���yip9�`�t��-�Tx��T����R�g��UV[��K$��&�1�M!.Nc��虡���T�E�>�=a��-6w�U�
<�V:�/��B��Z��J� "\8o-�`�:^f��=>K,Bݿ��f2�	��������|=9G�'��6^��U��X�T��?<�߰s{���Fo�m{*��`u1�oR�z_�������&g�'u��]<yzM�3�;2�n� =ZV8�Tr���k��\���7��b	��SZy�Z��eq��"��b��df^5fx���/8��SQ�:>QTGۤ;�}X�l�4�][�J]�z_���L=yz "3�N�k-e.U��OZ�p��@n�#�,��+?��eI������d�Y�34��(2�ViX��H���?J�6bK�\6�]�`�hF[�4���O ,1R�ǶY����C1p��օ�,飞�+�aW���͠%�F<�=/ϙّ��w}\G�2ˉ�<$�=��M�`�J�+�e�>��A"H1Ѐ#�h5�m2��y_'�H���ꑤ�|�z�~v�9W��k���)��Cyބ��cF�����Fr�-���9�]���[�`�H9WîI�d�~��cT��Q�2��bd$�C�`�r��"������Aifݨ�ȌG�`�=�gQmjޙG=!��6s��o`�?�w.��h���1�nFFN*|�Z���Z�7E��=���k�6[���_�KWY7Ou��F������ ��.��֟�θl��*��G��gQ��Л��n��C'���G�g]�>�Y����>H9�2f`�-�u"G��ܳ�����d���"�����rJ��q+�?�)��N@K���K���c�L�S8�e�)L��& ^�y��k�{�,����7T���ѳrKd���Gm������M��@��c
HО�!r;m�*o���d�<e=�YC_4n7��$>��mu�K�~o	�y���*58�3���&���Z�(�&�2�g[������.�.�$e}����/�iq|A:���^�Ӛ0?Mj)�k�5e�
׷�R�t*}�/�æ�0L0$��Rt�&KXy!x���R��J�����]Õ��� �'K�f���W�W�3��� �#a�+՞ïN�j���_�j�
�n�s�R��l0 �g_5�Yː�6B$�a8� d��a)�>e���9<tԏ>�y����p[�tm��b�7h�� P2-I�nW�rm���L�C����м�޶�~�B����B��T��������b�4Y\�l�����&�<�k�/
S��+s9��e�S���ӣ&�9�@'�۔�"��<iw#���������>�oF�goᩗe(@���/���2-��|^gj]d^r/}��}��|+z�l�I���0M����s݃�/a�s��"��m}7%����t"ښ"U�>_��e"�����[w8�.�����1~�"b?���>�Ҏ�zN�c(O���%[�u@R��&���4��3�o�,IAMn�z?��n����	�Tv��Q�J��w�E��Ť�˯M�Ѳ�t��A���ڸ��� ��Xm÷�����+�T`��H�qN_SF�˥&��5�1��5�^7��}lV��-��g���xqrX27���vn%A�T�qz���ș��@0&�'���!���|�/��bB!�o�Au�K�u�Mf7K�cH+cdL }�s_w��E;-O�J^��ُt��_��!!�<�T,�Ԟ�<��W 0L�
a�Y��1�W��1|G;S��L���3���m+��{�n?�b��w̚�2����Qq�u�,�?YX�Iá��n��K�_��R�D�)=vy��<�x��;���Z�A�vt�"�E#翼��u3v�m]_�ܕ{{���D��'˟��r��@�-:�"�m4��<�lE����e��Ȓ�q?|�M��))�4��ݏ�Wg
pR�~(����H���"�t$���g�����Ȅ��A���,�A��*)^l/��us-,5怓h}��V\ʡ��j<an1�R�=�A�9�(1[�{h�U���������츚�u�c���O_�޲4%���*���P���+�@hÁZVX��͓w��aр6��`؂�V-[o��������@u&>������m�٬���Ou��k?�	��!�����`�Q�@h}�u5p�	�#)N ���k�6��6�ª� ��v��l^ǭ8W�\Yޢ��.0����`�dО9��C�Oo�qn��A�m��W)i�i@���6R��ϔ��0h��~��o�F���R��K�O�S� �H!���V{L+�.�����"~� �nnT	L�!���H�jU����id3w�l����"Y���;kh0�b�(�.�R\�?8�'�6��byx�n�� $UՎ�Q¼�\rz�]�A��`qG�TG�p�Ȑ��T���W����{`����?Z���Ksy3D�]J����6��S�J��������)�{��'��MUZw;��o��F`�� ₽6)'}���O�0�s�6o�����l�@�U/?zU�v���Y�}%��,���tY�4�>T����'!�|�e��(ya�h����%�	���Oh��x����$�0\��	Ypާ�a���R���%X�ny�����J�b�5<S~/u�?g�$�03uޛ�j������Vm ��,��K�����L�# H�� ��}�e����jn;�B��h�1<һ��W,A>D/���D,rP�\X
�	I��Z��L�9�ӡi0A��4C~q%�))B��X(�DΉ
y6�4���=1���i ����z ���E�#Kx�c������I��F�Kا� `g�i�x �����WM�n$��I��� #�%6/��0���BÂע�5���.��1����˺Q�d�y���APm�"�o��������k�����KL��u���PD�P"��+��8�p{V�a���xn+���Ʈ@���'��\O��ݿ �����,=���E�U	Gaem��%�DY��Fkm�âv�o߅�����kM��ݓ��`[͎�qn~wJ~0��5X5����%Ĳ(�J��:Qi�F-��w��m��$����˿�����Q�?��	w�V}?&k��s�>��x�K�ſ�V%u�ζg��`���n��`�����#�X}��G�_Ǣ��Ě&��άJ >��m��M�C����Ħ
���' TyK��ٖm�0�{%�]^ :P�[2�bx&��0�:�)iS$ml�:�����Gw�w7E�Q�����{Q^]$������p����u֊�������-�M��⛍<�+M\/�;h�1s��Zɫo p7��݃�)�1�Np���Έ'�{��׵7ح0Q�23�� �K݌�W�XK�rƃ	>$¬����ٲ9�Z?߮nQ���M�Ӌ
`�|�>xrp�}E�2p#|��І�%dވ���k�j�v@����C�a�%n����5)�����29��D�[}wu�^�{�~g��M[���I��V=�w��;�@ߟ;�7l��,�egA$w�/E��dBM9P� ȹ��Y>�drN�qܟj\��6��������њK����u����P�d%U���E�CX$���> 
vd��c��NKY@w���HT��ѕ�Y?gV[���kfd�1mv�fP�����7�e0��خ�?�����ZN�#��׫��P�E�g6�54���vi#���4���g��W�6u�O�aU������������*�!>ʋ����]<���
tu���TT!>e�T:ǼT��F���/Z`�b���c�S��Y�ڰ=�~J��2����Z\+sĖ��Tp�^�c;iGh�~��>�w��a烇z撥��y�B��nU{LŚ���DOT`4;kC�ާ��/���M����=;*,�ʊM BǓP��9mn�̃N�Uֻk�o��־M���NG�1����u�ΖkzT���b�u�xy����v��>hIYT4yR���{�~����B�N�5vo>�����&�8���x�)냪��#�=��TAY��z/�ܑќ�PX	�*FZ���A[�-��)�>R����o���*���N�܆�f�AQ�	W#���2�<��-�㿷�����8rMCn����F�pEk�5���:�G�t��W�/Y KP\b�p]ޒ�x+p�8�"K�C:��
݇�l�VQ�>�$*'}�)5�	�U���c��G�sh�Q���P��b< �����6����,z�	Bȣ���ר�sC/Փ�彬���-�i���(/���*%]�ր��im1���Vz�Q��,R��B���4��q̌ʮ��-C��~貸fssҡ�$H�����7'谴�x���~����~_Gd�o�b:��+���XH�m+�4���^�E�����V]i�����,l��JQ���*�����U[���J�y��Ru�@�152}hz��XO%���Fl�<&��R�� �<��{�{_�_��\���%4�{K�@�qv�jLF���t2��O_�k������SZ��IdzY��\��	��|�$��S��c,Ӊn��-6��ڔ��q�>�~ɗ�E�|�F}
RAiFg�9ay�J �Q�S%,V<���x��Z5
Ҧ_B�c�M��� ;��6��;��=�&7�h�DgZ|lΎ0:4��011�
9�;��,�b����CI>�S0�ǵ�=a�au"m�$�=�B�#�]Yb,�6�S��N�Rmi4ď�
_��\�@tU5�Q�]\����x	��0U�Ҙ���X��@'�Kf�&��i?dl¢��8�:��v�w@��|��,�o�*\�CL�u�mv\�z�l�(#�fѥU�,�|�<���a��X���I1�Y���ԃ蒶}����[�^D�9�?�X	��e�<u'@t@�}d�E�����TbX:	��g��H�v��[�$l��Vw!�|�u��ۼ���BwA�����b�=s�U̏�e�v�1��f�R�%����J��}��L�D+�r�*l�G\�����ǿRLJ�My�1��խ�e��)@����T���B[b�i�җ6��
��i	����_�;G&D&J�z�w�t[�!c��7;L�T�s�`�p�?\�&���i��2q�����RWOd�l���Oc�8XT�>(0�����:PR��`�gmd��A�k�[����3��P�����(�p����i�S܎-�F�"�-�,v��7Fz��Fܱ̰�Rn8S8����.j��O�;9 i����{�+���bk�do��W㌃yƸ��R6�k��ޫ_i���jP�a��+�(��zǗt��o��U���I'U���I����S���h�tLK�-�ݛX�p�³l�K���C�M*Z�1���n����,�].O��������*U��r!#j
t��aa�1�Quu�|� �9%lP���tQ&�d^�.*�%dM���Ü/�n=9N8�Rn�΂����t�j������Zr����D�:(0�̮v��j��ſ*d�I�&����3��Z�{6|��ἁ�^x�_/<�)���=²�l�)��#A0K_/O���.�ČB<Q��ޢR-r%�/w�A�o7�N#��ê@�">���fA� Y|��z�5�-��ò�@�������K:
B̠�^�"Sd$~빆��)o^ 0�-)m�#�i����H����i<����JĘF�ـp�ⰻF�!�I�]S���\o�5����=�i=q���HL�=��H�@���E�a�ǧ��d>U�<q+�G�u�A
L���2�+�����be���QŘ~$��������v
�6�������j{�b����Za��O��D(bG`Sk}$��Q�>�bSb�y�\��7;�Lf��>� �N���6��i�:{�hR�M����Y��n��0�+Bs"'x��g��+*�,Y5FA�m�<�BX��ϵ
q��d/n���w٬���`8F<M��]]E�[��㰙�j2�����y�-x$�!s��^�%�SQ��}D��M���o>Ƿ�6X���)F�2��K��T���z��;�"��]��0{��b�R}+�s>2�5�qg׵A�K6��V�ȯp/�ύ����#8��8��!53�-����FܨXʶ����)�����D��ŋ���2Iٴ5ղ`(y`��@�����'�e��]:�[�YhDU�{���f�L�l��#je��c�Ps1L�}�~n�ß}�����*��>�Ł�䏏��lCkg3���.v���
�yv�ʽ�f��ګ^��'�u�����2������s.��Q^�,ez<�C#.������:��Cj�Q�SQ��
9���/��r����t��J���	���<�+�ى|r��n��{.��#�aޙ�~�?_�`�8��ͥ͟��=�U��͟$|i9*��v9�7�mEl>��a-�]Bs��~��Ϻc�-��=�	΢i�K��G)ؿ@b��$��B��G�\M�
)}�SN�)�
WQ�kq�-���/G˒�s\H_x��Aj�b>��-h-��g�
��&�Mj7{K����'�HAC�����%�w����w�<�ꪨ8���bc��w^	w%ev�5B�H2���[�g��mS�Z6�D��'�����:n٢'�+�����5S~
j4W��WyI���?vC�v��|�n�9F.�B����7 ����14~��{C�Yij^qr��:+����R����y���#��A���wܺ'ŨS!�	��1*vUЮk!�v�gX\���ٗ�Q��+,�>F撧P25��E��ւ���@(�k.�F��W�*�֑�ܺ���b'�"�S�x^��;��~h�n���;�g���p��T�Ƕ��E�8��z�(5\����٨�gJ��
Q\��$g�sO!��$4z�n��]�R���)^�����*���h���V�=��P>�P�$��g�V{��d�#J�1�|����G�H��|�Hv[I��c��[��alq�:^ E1@{}x����������ЂZ���]N;��)�J��ғ��+�& ���y}��J����)�K0q��T���f5�,�6.�
�^F��Z�����] ��]�s�l�h���/�MK�N^V�����M����15����X��ێ���3�+�k�z:�(�$N��k��>4��E^��j���
֋#Q+`�>b3�����v\�v���S�%�Dt7dG�i�@��_lm/�����A�����=4U6 ��^��:>_�މ��_M�
����o�Nm����p+Es��T;n��J���Qd��ê�e��j΢��նl�;�qϋ���FРY���K��QSSa���j��������8/5	�~fi�;a�J������O[>ܿ��D���J����ȶ����w�㉔	��B�Ɔ널E�
��,�҄NB��Fߕ�$:~./צ���]�����.�M6��5��6%t0���c�R��f>�PÃ��!2�L�o��#7ƵL��j]F�������5�dc�d��V|�4�yc!1�:��3O�EjN��h�x��I��^�ȿQ��V���{mO~�J��\�Z��B�vm`���Q�g�4qS�jj� ��S��s�]�51%L�TE���^�&[��r��i׈�RzR�T:��T^�|.��e�y�v�^G��˃YkI�N�Dr:�+�����@/Bj*>,�7�dFS&fx�$eON�w"�T�A#.��F�G.���+��P$%��w}�������Gu����ӈ%�"���� �k�D�ߠ��ü����1��39T4��\I�P墶x[����O�� Ha8�6-����y��笠s�(#�u����~��>.�f@'#��F*�G2�\jC� ��텛���u����Uݮ ���0�rhA7ѳ}�Յ@�s��J���'���ꡙ��^�83:{N�ɽ�����,tW�|���NV7���޲�;ο:��Uμ���g��^V�\D>)k�cپo^0l�fQ��ὣă��/�@�opPR���c��f��wJ.UX��0�� ��Y��U!���7R���_l�e�x9�,���i��f���yl{d�-8����F����y��!v�%������y�Z�e�h�~�zZ�c��ZM����Q�����˻w#>�]}Wy�N�b�6V�)�o��,t3l���myA�Bȿ=w=BǾ����ݔh��}8S�i���D�:2n���ő�,G��D��k���q݅�!_WsYc`���@2���隔����C��L����A�lԴ��[�p����\�Wj oΈ�%�!tp��C�Xp��2"��<"$����l͈�Z���qsf&�P�zCL���J���{|it�I�K�л���!<#4��5'���L��4S\�C����&{�l�p�����]kw3
4{���=��L��Z
N������1�����
n`�3�[��hVPa�K)�AT6���������g��` +|&���z��xY�ތ��;���4���"9�K��_�c�o�
��c�
{n{�v�����R*�@e��N���;R5 �{�MsG��ċ5J���=��#?��,W}-�e����Ȩ?�)w8����̧I���W���y�h��z�Ů��e���$Jp$���\Kܸ��Z�ꉭ�2X���$��7�G��%y����TB˟_��w���TS��M^/�������j�Q�f�ըm�Q9�J�%,�"��ݝsg�+��;Kd�!�yg����mW&�e���X���=, N�f��~i���8����p;�;71�ę�;�H��#qY���Y�"sN�����h���c���\@�T�K�%uo<`RG����f7؛^8/���!�Wȝ�v����'ޥN��?��Zk�t��09�VF� �z�MZ�Հ���<Z�D����)�) ]k�iذ����D�*u��0Jn�z)����n��Y��I���8g[{�kf�F��"�@���I����(�Y���i��+�(/õ�K� '3:�?~Xҫ���4.<0�c��S��O%��Z��C�C��H-8�q�7g2�@��vG"Ky�F86�ݯG�(U.�׮�u*>��[%gE"
bo��Щ��M��D��|����#���6�����1.�8�~I����}�eOV������X�x�t�.m�����|�~��eV��RL��h��L�w� ��8$��Y�O0�6�"��]95L�ͥƋ��m�+D�!�I�mb����A�C�%�!�>@��'ή��&\w\G�&C��uT>D?KO�c����r)�hQ����#�@�����[�6�-yI�b�zt�l�����Ub���d^1v,3���&�a��&�?Y
���\x|-a'�[-~T{�O?�+�a���|����!+oK�m�N��ًvl�SC6��u�|#Ȇ)��j���g�^����'�L L���o70�'`��f�㧄�!'RJ2g=����)_����|�����QLx`w� p�@To�I��}l�0�ò��]��i?��IK�.�D����"���ud�Gа��>b�B�1��or��QH4�śMi�$ƚ�2�Pq�]�y|�����%�rh���M6";�+��TO��t.00F�OTM��|��ekt��HJ:
a5����`/#�~2F�|x_Z{��3�B�=��|@7��a3 `F�վ�x.��'��Y�ZCȹ�-�*i�[��������i�OJ�Lc����w
��?o��������!�]@����hV�G�Co�?`�P�U�p�k��7i�-����'�j��hlPr�o\��]�
���k�?c>`���Pi�{�&��/B=��u3�<b98��1M����O��@(�H�H�b�
��h�$O����5�-ig��E�8��Y^ cԑ3ƈ�{~l����.>I��+_[��#	�eF�YG���D�p[�Y�Qn��0Ct�yF�FjCf\y�Y�p��V�(U2Ky%~�3R�:!���K�[بͮ�?���A�_�I�W�g�]#�ĉi�!]��y�EJp�y�9.�� ��[BKςf�~]sP(�!�{��}T��{|bR|�>���y�2��퐭��lO�nV���#�-z��`D��>��2`��[�G��0Ŋ��H��׳H�@wK.R�*2�<
��7�ݦc8�� ��|!s.H�s5-�<�(ᄕm�=(<�I�U�Tzp�
h2t�y3H�%C;�U?�̊v�gT���w�S�����"��Ė�ɖ|ɵ���`;���<4b�iao6F�� �o(դE�p"@��}�-J��Ŗ|�2Hj��6�\:�m^�\����/�+�Ÿ�9��z����~$��?�+�j�������Q���j�x�l��e�c����0��5��r@V�r�[�ㅐ�~��R��A������3��K�.�?�:�t�Y3������"�w�r���_HqӐ��-����\��)a!O�E�!%oMa�</D�L���v���j�­[����찖�c.U˹A���ȑhms�iṱ��u��h�ZJ!DPT�ף�Д�@�P�}ƃ#T ��h��P���!��2j�_2��2bA�?C2��.�����I|;��˪��F=�xft㽛��#,�<����a)i�b�s&Yy��
�i���&)��~�a§�5{��|���=U|�܍�}|�2ن3�~/�̝���	d!\m���%8f6,�?:����:{�ws��}u����M�դ����g��ig�����#08�mJ!^�Tn�\�S�3D�+j{�������M1���<x�s��'g	 ~�i���[jb�t���;c`���}���πHw^[+�A'�voVqh"�P�������o4�v�����{��n(jy��ko=����jڜ}�;?U~N�w<|\�ٌ�$��3���P��+�;>!̃�r�,ح�V) bA�~��Va!>�[ ���)�dY��v�F��|.�E�%�9�P�p�a��k�I.罛["sS�T�����*����a��gw���w�G�O�g�b�4&�o����xyl��bԃw �|X���j��,��W�XoSͫju��$�	l�4�.��,k����A���+�G|��8�X�"H��1��z^-��lN�&}�Ru�C��L��ɚ���1�r{�ZO���/���(�TK��4��Y�M��k̿߷e�WY՟zDh1+k:�wK� =�a�0��� Z�aJ	C��fs��H��8���x�8�N�{��kq�ēʦ�o���M�d�g���c��@��-�޴Sc�)��/��^�"J| �7���c���s|�\e�Ԥ�m��������8v�ʯ����S� ��W&�l 5i"���89lrߑ���4D��b�=������Ƥ�S�n��0})��rO����XU+Ϯ���� �-�{��v�c�l�C�6MX�,�}�S��4f�|�I�cAf��:���%��R	�"�����zD}�|�U�7n�E���6�b`y�jKKoU�gp�iZy3�Ńg����I��aɺ�:[�	���f��k�� �e�E#��ա+��`�����v�b�۾%6�Jx���/{�B�(��C\`x�Qj���]e��X-fv�}��/���UǥH_a�vBF?�D Mg�����Zp�}A+d�� w�,"�4L����x����'8o����+p5Nl����Y�e���Ғ�+nA4�r����=� �

�ʹ�'Y+���%�����Ί;�k�{53���8�\<���&/���� ]zI�>�=I�/�90eH��ƅ/��KM�c���5��i�{̉sGa��!�a�˧Q�[�j���v��͕t�L飓�x��#e��*���9[;`�����{�g��;fvfyW�~m�"F�)��%�IGS���!p���	}��d]��>�7��?(�r��{�@k�Zco�������6�I]�ΰfŇz��mH���_����"�-�yT7�B�k��^P��_�o�"00Ko��G�'0�������rN�<
J��o=�o���;�u�Z��ݡ���V��J�d����C.�"�Y�@�����@�y`wE�ty���#��\/�F��^g�6�����ݧ�\��PfV���r�8�Cp/:���,;$D��6I+ڊ`�^����A��2�<���3Zٓi�"K�C
��s�&�~�kܚeFb���+Y,�j���d�c��)��l���8b�zQL�D7'Y6k)�2��B�K�A9��"�PJ��a��� ��He]P�\^��o�d.���G ]�����J�3%���rV9'�wu8R�Bà�Q��ғ��4����a_��/@�%&��ޙn_�6-�w��Wm ?�؂��I\��R)z����H�����*�1���u�NZF�Jmia~��	x�,k��OV�e�W��������r�1N�������.��ji��<���ˁ��>�݉�T�3��yC~1�yS��Oj�l��a�R�_dT��F>ޚ��
���N��19�g�IJ�@"�1d(Ю�g.�¢��� ��*JǢt�!��NX<����������?��+ =��������W{}�?����MV|�/v�p���ިh���k��A��ch���Z:�9����Ts2�Ac՘�.B42�(��o>�h/a���˘�s��=�v��F�}�B>�E�^�9k�G�`Py8��B��P���ޅ߇�eY��Jf:�7.<#���D��0제F���HweQ2��?�iﺯ+��Y	?&���%�U��T{��B�PY�ҁ�\>鶃����щ�;6��F�Ʌ��e�7Z�S�C:�nop�B��otc�m����ga�A5�k;���3����614��^�|���;^�!��F�e6��S#ojO���R�<b�:���8]yp0;�����pX˝̓l��P���y���V��]�M04?���1�Z���hJv�g�H�1��;M�>KZn�� ��%P�R�l���:�M1fF[n�����q�+v�L�6"X��x����~�`*�&2Y	. ��4��Q��%�ޞ�E�(�F�:%O9��!.B�n�wM�b��4.z�O~����n�*�]3p��4�ů�:v��>�q���� ���`��c ܰ���^��]�$�g��;��&l��y�dZD)�2�R�U�&<��9��W]o#�UW�Xy� ��clKk�w!��n� ��lB��֚L�9ZQVro�(�k	^XY?�|s�*�`�C� �,c��E�(\L�~����ie�5m���&�݄�úd#<��2�̂�(k�C�F~GuM��e'}�1���&��#�	��)�Ը��b�Q?�{��G|�}ո4x�ؾt�AEX��Y��\A�k�Dې���x]�'�7��`o���S^�j��T��x=6�@%:�5x�䧲��n�v:=՝)�yO�	���P!�5u��\i��j�t�R��z�]3�}6f��H|e��,/��2{�CV�s�y�=&�����
klvSw�+ ����b�%J���f�e/ĉ���;-|s�3
nq��A�z���0�g�0�n��A��p��39<��$�r��hc:���i�D
(~s�������#Hw
K=����8��k,�{O<k}��P[6&'���`RO@{Q���/U�ׯ=��Uz���~�%�+h"_#��0Qψ�z��:ӐN���ü��I��N-�����ܔ��w G̥N~�=@��=����8b������"Ϥ5�59�-��,�\��
�`�7bb��g���MЇ���{��̔,B�r��:���6J���@�Nv�)hw.2#ޅ*܊R��ʌN�J7U\�Kfي��i��{�&E�-4�,�v����k۽Sn�mG���!!�_��<�`z�j�׾�rN�!���XL���U)��Z��j6!]�,��;&xb#��[��%�?�dN�tv�Q8hr4dQl�y��h�X��y�̢����w����%������Q�x\��YA]o��Ӟyy	�z>�(��2�����܇�Ms\�������ڥ_+��M~/���SBk!X��36G���Y��#�߽�U��(%t�"Q�S��0E��Y����悧���N��϶�>�9f	���c���o��NW���#?/v�߿����%������=9�V����Ϲ��w�#�&��.h1漵R�����u��C�D���ȅ��9��R�PG��E���dcL�D��ke%�������@��/G��p���ԋ\�	�2�r7�����2�9�
��\��x,1l7�qJ�gD������'�S)��`-�x��}`uq+!�6��?$Fz�1���R�L�;5�H�-JPw�5��On�)�.���s��T�&�Q�<��8ޏb��GԐ�hԿ"�'���E�e�J�Ꮆ�U����	's/W�֥9��	}�������Ј�K��8(�Ր<�a����,�����sU=�1'�"���I;��c�C��"ġ[*9�[B���"�V#�~Nw��_�X�"´f�$�\]��(C���vt0�yH�6�Jg<� z��
U#��V��Q�h�[�E�����(�l��.g�uVV߽S��'�}.XT��kd(��|L����
#^+�׃�}Z%[W[�+��u�?J��->T�6�R�1��8���FE2%�u�
X���V��x1SXAr^�8���N5�����)9c��jY��l�	&�� ғ&_zO��~!V �Ica��^����Y^,�&�s��þa2I���� 6��)g��owy��o��'��?Qu��V�,XP3%n,EQ=z�����9/rb�#�U���\�$G��o
��N��T
Z-H�k.��`�p�>:����y��IQ�nO}b_N���Chʤ.eV��I2{�f�� ~��N���|a��;�
�d~���v�	I��+�˩��#͜-E����:�����y�== #��m��੯U�h����2���.�"�����Q��u���3���P8u���jٸ^�k� �o#'`ހc]�d6��9&Z�D�:���1Y��J���M�I	ޚ��|2����LȲ���Z�y&nvG]Ժڞ�Bu��.�����[��lT7;�c�vA��Y"� D=FŢ\v�HT׍���R�D�"(�(�{���*z;y����LH���u-�:���m73N�9���'�u��A�-��Q�M�}�xE\ј_ZR%d�+�3�[�90�2�vzr�6���v���B���/Ot��1���K9�ˡeTM�H8@���H���'>�S��u�w����Ͱ��	���Nyb�	(H�>R �1m3��v�ͣ}X-'������v��'E��9��/�1����x��:O��b���.�FJr7h�2Z�h�ҵ����|"�Z���#�Ꞥ碅>�?5����Q��!D;`��/m~#����w�N����B�1�@�m��*Г�A�t�ʷ1�+yCDs��!ҍ�O����
�|�XQ�Bu@R-E:�o��j�U{ a��G��>�,fv��� ���1�����D�$�i
ӇbOp�����:I�Q2�Ņ��3�� ��J�F�"���I4����K{ �[���ˠ-�W�055jUvJ㐊�~G+�pi��]#�SȞE�	K|���#7o4�C����|�GG:F��R?��x1�Wo�_|ք����R5L_^"��`�Ck�a�"�7�}~?������_� N�Z���E��#v=��'<4�JZ\.F��K��:g'Y�����p��x|����d��H���\W�� �h���x)����W����]r�ǎ:\B���9n$�Q!S��J�������������|J� L��b�/O�16�^g�A�y���o��$�������TL	�?[�E�ל򗆄Rn2��)d�.���)���Rޕ�1S�WRH��[?�e H�0S�&�3���,����k�Q��Cހ�"E�& �E3~�Э�N��mR��'��+I���!7����}Z�DfZ��[G]����E;��զ�����Lz�sJ8z������KM��N�Vt�Z��K�W�2���}My���;ȣ���V������{���Z?�D(v�.#�9�9G��Lx�a|`�cخ�G�0B��[AdU��:�qT?o#�b��^\�Mx�='W]�����w+�S���P)5��*��eV$�s��)b-U�������k��s�g�?��V_�y�/4�W���KM��
���Ԭ��zي��=lW����xG��ȱҝ��H��b���)��!las���Åit\d�+'Kp�*d�B�ӠO��䢏'i�%��6[&���:�)�j/Bԝ��`��mi�P]��#2M�O�]��=?����# ��&���]*�u�+�
2se.��?�1h�/#�������k~�b�Ò
�['�:x\-���XJ�#C�`x�r������a{F#��Z$rw���T�����fAY/��ǣd��V�v�:69E#��s����6g���u�Y�7�S�3Jw�q�&$�,�z��7�"I������*�sx���$�Қ@�D,����}�YK��noaC�x���@�u�,��7��ɽ�<��?B�~ɍ�C_�4
7o9B�@{���;�ݕ��1/��,U�J��3�7X��}z��3!��'�,��2��eɣ~7��<l�5�
�]1|c��(�I=�Yu� mNi��j��?_���"���3u�Õ��C�W��4����]���߬�K��u���_�Z�`���o�rxҨ�UF���л׊��q�߲*��%��oHɇ��<���c��X�4��P�A�8nD s4XJ݄���Q�/�F��M��gX��ƕ�ژג��w�sGD���"�@� �Ysߥ|U]�'�o&-&c���3oe"�M	�^�@Qh5����)�2v�/�������B��2�:S���|���K���Խ4�i���JaDo���xp���CC�W�@��2�ىě(�_�����>e��B������#�,��=��W��z���T����N`/�:��(W�*���k_G�!r�4�lq�]������K�(��\c`:2V���3(P�ӷݬb?�*H`��/(���Y����3����ܟ9p.� �+-�KE5�~-�Y������n��6������`y�\r��%vA}�*��_)̩���k�9��T}r�Í�Ҿ��W�ײ�CvH���TOC��"ѣVOt��>��������X��I�69?3���|"l����Zh}�ݷ��I��y�Y�"�8�H�.V��]Z��~��в��#quT�#�
�˸1�������-�g�X�2܃�x�p'1���j��nC�,�m-"�{N�{)L���5��9���.'i��-C������N�D�N��1�R ЏG�U��k\	cP,_��a��Ϧ���_!Q��F�
�%�?��g��ַ�M� �Dx��:����LE�6pE4�TB�SÜ��uO�0�TA�r'�3�`K_�5S��)�M<��N�R�So���gfcF��y�l1��2P��4�nc�|j���]��Cb����'5�y���I���1Kt%�3hP�v�.(Mī�����2�Yt�}Q \_^>��y	�,=�FYa�M)7���zS�q��UH�#��iv������Bo>�ƹ��/^��O�6�.�=2C��7lO�C��a�#gF�`膆�h7j�=ҘY�Jl.�خ��:��<��,�����?(;M?˚/�hQ�xܘ|�}��)/�d5�[�h���+���q�/Q���;񲪇���Lſ�i�1|t)u`
r��D�ѩ��>��f�d��}n��>_��__�(�C��apg����>�ךW�⮼�@>˃��W~'%�^s90��U���<JI���@��q�����Z3��lp�a[�^6���eS�9y�����#Y���-���(?�ڧ�[��Xc��a�C���l�w#�R���ۚ>�P���X]�|����H�J)M$���%�5u\�-5B�]��޺��}�n����kV�Υ���7��%�M!��5LӃ�g�,Ԅ�6> ]�oe2@�-4�bPysu)URޢ.k�Y�I����h��,�^�/���'T['��z�V�S�2����t\��Mz�	A���w��.�/Ec�	�dXM[�][�3��|�5���D	�N����)�'��?�,�J��!���$Vg���[�Ȋ�>�婰����'K�qS��Wʿ�wz{*�9M� �򔺜)	,�w��w��CW�r�xDB�����r�b�vLJ�R���e|K��.����;�D�M��g?�GV����*���j迦nV�9SdTu��Y�w0���[���A�to�:��W�KLXn�w���"�4��W�?�%����𠿖�����k���.�k�A�m<g���! ~��C�V�~}nm���s����O*]#=��Q���>;YY�l�W�@�ܫ}S(�<��l�+��O���-$k� 39xǊ��`.Oc%�1#e�R�-�휀�|c�K�!I�i�L������r���`�Ѫ��������	JNC���	U���;�	:��1iʐ5��.���[sɗ��gi�M�1���	Le;�������H"=ެ��~i��|�T˰N�¹��ϟ�PJ8X� �G=��_x�}*{wz�Ƙ�k&��v��~2�8ؚ��,e7�,y��Y�`��Y;Z�{oӵ�j�[a��jJ�Ch�l������r!}-���X9���������2Ð*zS�¯��)�Cm�#��r׎A:$/�?f(��x��z�Q_���.8�{y��c��2@��9�BiWƿ��]��X�xFA'01b����&�>��%X�y��j�ϯ����k��F[�?z��时4g�$6vNWK8�/dX7^�I�7�5���'�5�����}�q�l�]���C	����n�J�aE
����ܪ�Uֹ]�$���2���/��2V�õ;���/�M�w
"o�D�9�(�'�+��Xuͯ�k�<�" ;<�z�{��K;nқ��ʀ��q�A0{SM�N^�4�b1ov����� 51�G�'��*��Oڕˏ�g�E�o��C����w�q�a�\��/�M�_���4�ic�#��hs�����v��b�r\��-ru���'+_,��>�H��n;J���)����5�8ۥ�D��>AD��^�3q�����튱B�$������LI�Z�h���K�T�q��t�6i3A/��s��g�t�����
�W8K�1c�I�1jӌI*2��P�ً�������1�K|'��4D���� *v�Q�X��hr�N��=5���6�2�E�+M�~�X&���iI>C��Z ����TQ\R�/�JY��}�u����9,@W�I���+Ʉ�!D,Z\y��[(]͂Vt�����Q5�w8��\�U>}�Ʉ�V��SuJ�M��#h���T�3e�aU����g����7<����a��3���K*�e�j�ّq��d��_I���;��/'��m��c�>������N�HPg���Th�As;��PII��~o�x�61�8e[�� �wRǛ��}�����c�ڙB�[��(�P]�1p�~��F�p�q8L��i�p~}�gҎ���O�|��PL�����Z����k�P�I;�f�;�<4���GC�bf[���B�Jz.>�3���۰](���Q���ns�]ޛ�~&�s�#��"�˒��s�ZZZ.��ӈW��6'	b���Ԗ��������}0��Ph��u���&��f�a�|ɖ%GV=�H^�6Fy��`S�	��awU|�w��WD1����r����C��Z���=�h�TQG�!2`�|l:^^��<w�� ����m�<G��/f��m���#��hޏKÎQ(���d/�"h~1�>��l��qىY�l\\_#��HI5~R=[���k�^t*��>���UƲoMP�3��@��h�gg�U��\(�}-]K�b��弃a>B�� ���J�dX%����KHŔF'�Uu�>\��9��7͈��N��r�b��ʑm[�J��)���js��̚�֏�CI�Vm������a��=Zb�'u�`n5:IB	�*C<W�+`����yw3�Z�q�F��J������Oʞ4�5��¿�N�?��i��;F/��÷v�Y>���c$wT�����*M�F d�������=e��sBHƝ��r����:�<�$x~��?��؀�iJ`*�����{�<o��a�@Q��our��&j��t��*�{DY��K���V o��NL��9Iq�D�t�b7:4��iݟ�kr ��㯋H�ufx�4'�&`��YN(��Y�� *��v"���\�<4 ���e���n2��QjBX�u� !Fa�/F(�!ͷ����!���"�67!��|�k�1cy����}i����O�P�l���z��v�� ��C^�]�q� �,$�8y��7B�Zi5 �r�Pf0W�&^���A��ZZ}��h�]XNݍ�eN5��
����ȉ(�z���gx��-�翁�ߪ@Q)O��3i3���9�ڶ�vİ��	�s�=���p��_���W�U���Bln�����`e��E���ҙI4
}�4c���3 M�YT�./�(A�ݚB+`u����rRnd�H���қf2y�_r�-}�W������r	.�I���;l�!�]͈�:�J���sT�G�?ej!�Ի��y��M�"H���Y�>ɻ��ژ�c�k;8<��ؙ-��q��}���ɒ6��4p�h���}�/d���e?V҂U9�bOYc��A}�k;��&s�^>����v��#㳶�����H|I�gK�y2=C>1�Z�16��M͵�c����vF�y�E����{lə���fz���f�vΚP�~�e�*��VL!+H6 K�Bu��#���r��N/Wp����L}�V�	K�"g�-�R�t�?��1#*�����rFXv���R�?��Ă{��m�kgՒ�%v)O`�<��t�D�Z��͈jTkr"��Ѳ:�}�-U�#LW�b?D}��I��F���C�t�Ҟ�yV�bK�,\iĸEQ2��槸�z�����C��F���J�	XG�]��򏕊Z#Y�OS���ڑ��F��=���'啞 )�p#�rH5�ջ&zRV*���s���z��q���t9cۄ��Z0b���Q�Չr���_�A�s�g�갉��|�(a����]u�/D8�j�K7��bP��_B뗉W"ϳ���L�>f����8��ާ��yCղnL�h�B|��Ka���KJ(��W�2��*��1�X5^��H���%�(j#�j�2�C��\�	�6t[�9�S�F��b���2�L�qI�6�Z��7'k�(�/�fܣou\�n~G��rN�%�awɀ�`�����h{�U-���-��d�����
��Ki��mu�����;�?�D�I��r[�^����Ӑ��X�ӓpk'3)	�j�-rv��w�Q�S��C6+��$��%�8D��i+(u�&m&u�,U����u�p�	zz��[n���C���iX�{c6�l$�%W�"��ť�`>Qv:PIF�����K~C۵�e��ta��9ޮ���T�V Qd�l,�\*��ķ�U��ʲ�"d-�#��v��.N@�h����Јn)��c��$��op�j���#��K9��m+�#�OX��p~q�V]� -���wAi}6f�<�:�]�D��4�L#�η*� ��Ӗ���0 .�Òǿ'�\�߈"���]��n�B� mA*��CT�3��{�.d�������7j���+뫓�\��j��31ZrOG� l6
mj�5	���zx�r��P]�@��|R�Y�V7?��RG}��#���b��W���rT�nlf�G'4c'P�h���4\�'o"��>�l+����q	D|��2p��%w$�+��<��r�4��yl=5ߡ6?�r��3��; �5���
`@tnGם;,���#��w����r��TE/z���ܟ�8l)a*��ϣ5�#~F,�l&¯nW�����:׎�ؼfX5f
��Ӌ#:��7=_���l�w���[��?���
һ k�H���|�l����?)��UF^�1e��K�;E*��~��5��ȁ~�;�f�BW�&�z���;!d���M�)]�%��Z�]��,�����-#�� ��V����7[�w��Z��{`�ã���;����z᫇Ӝt���=��s����F�����R;䫓�M��n����~Gʥ��mne�1a|�}�����?��~A0�2ĻU�+�#R-�uqV��@�nQ_���6|�2M(M���5*�K���&�)t����s��%����E|�k�Ж��������fO���2��4o~3oȁ�}6@f�|j~��a1w4���\c�~Qaz��i|�;�&�d���k�[H�M|Ƌ�7���$y+�k���c����tV,G��gq03u6F��(��	BU�N�*QɈ!�#U�_��f�ޘл�6�ՙw��%p�(�5�z����"�$p]i�::���.�y*����ﳡ�w�Vr)�N?_Ԭ��&��*K�U��e[�x>xH��B�"��w�ݎ���e���7tN|�|���M���*A]���u���Nߧ߇D�+��������'=jb���4�,6�������>P�6�w��践�^�
]�_˿d�'�eg{��T�4�/��|�0��A�����z��?�2_KitD&��I�m���Kk<Zu���ﹲ���&N���y����f�I���Ts�S��WU~���M>���ba�zXcKve��$����R��H��}�3�S��ǤbZV[P�����v�$B����EҀ��)�~IXYv���C��ܬ�T�
�!�/�zB���{��v/��J`/$5P��_���8il;�pH��=�X��]l��Ts�"zkp;��vy�K���("7ݰ�"�G}���gB~���'���f����tw	�-���a���ʹ/]0Gh H�ǮbjY�%�)��"�G9�-prCZY��g��`:�*�@	2�C8=�_��2�kAɋ�r�VLW��(�:��<��T[:㾈�
�~�à�8����eI��O���L�� H��y�x�l�{v#�t���#2`��(N״S�>��+b���!���6����Y�a���6�v^�����#�.�H�ۺ�fjN$���!�����'����aZRo)�F%z�/�\yĄ�n%�y6��?@�\�:Y�u|�K|Js�Y) B�AU3H>J�c	��f��s�#l�̸'&���g��:隳���+�􀼬���]Auә�lߤZSw@�/~I����b�'��6[��?�7��0�d����u����<���ۊS�L���a���ԖTkQ�n�1�d��.�4��s�<ֱv5��K�4P���H<�����U7B&�#��$8-��S�-#|��������d.�>RF�<�EwS�0���$���ڦ�����ᰜ���Q�f����R���bO�����r�Yޞ�2��| ���^�vR���B�D �uV��06���.�(-��m7��(�󛖊���V��(�19n�%g�����7�������ElR��Wf�t�\�|@< ߌ.k`09��KZ����Pvm��e�?m�~D�o������IA����xz+��-�V^��v�V���c�hJ���uNV���9\�w���i�t��ij�=���^I�s���-�W�$��Yb�P$��r#!,W���ȿ5�$D�a��HJ�(-_�OQ��3wJ"�,@��ٔ���sId0M;u��"hCx��2N�{��O90G�����xs����@	"s��$�5n��r���_B�e>�He����K�]K���?�,��+�xJx��_ �9Xvԉt����\c��wr^���W2'���+d���.J�{�����O�f�!a�c�*��ciߍ�;˨���JL�o�qw�)ﺣ�%D�&��K��xQ�T*�1�����5"��G���O�xAPN���Ec˪D��?��KS&����V޴��Ѳ���,U�A9�{3����e��D@h0���SJc
ւ�D�P��%ha'+�@!�W������d���c{���9h�Ӝ��Cg���OwF ��!Mb���ە9�))\�W�S㥐�d�&)h���[����ra�'2U�͞I�!�\��"ݗ!U)gۏ���2�K��f�ww�?�-C'I��G�&r�`h�,	�T��-U����} C����\r4MK[sڿm�c�j��kM�)���?䔽�
����D�Գ�/y�.,m�G#���!g��f%��U�TD�x�W�:�{��ު�c௜	<�%���e���#Yઃ��uM@Y��#����w���$��'�EE�~�-�,�,��K�C��<�t��4ĚH�H�<���
2��7�H��vE_�,ш3WoB��K�YZ�M�Qz���L���)A���y�� �j�x�8���y�����49��Ot`rRཁ�r6D��� �>�������y�tZ�qm$�u��~�=\�q���@V"U� �^G��į{v�-�uuX��J�¼�����{�|˥o�n��r_˭X F]+��z@�s�ȑ	�#l�C3鹡k��������.R�"�@/���
;��򌣢���#��\��{�5�s�YC���*C�QL��	����P>�xI��s"6a=8`(.�X�;yI��.��T����{_�.�b|������Z�iWB��9�/����5�i���}Xn�sD�Pޕ���	�+@���Ff�6�X�Ӥ;�T�M��"���|�a6lo�0A��W�}�ǀ��~R`z"�ޠ�#��xyVZ/�a`	d`����%�։U?�k<1���e@\N�	���5�Z���!�ۘ����p�����j���g�a�1�:H0�Ov�MdE�ߠ3�lg�faff��)N��[C��H���*!�E|�:����s��0DB�γW���1E\X��+G_��'ѫ�v��{p��P���פۣxH6��D���X�n���`�˙�����w�k1Fą��S���[�cpH��b��hP<*n%�w8 =���o�I�g�!\m��>�Hz�o�1�����h&�U�����P��E�=K�����k�D�:PkE��V���&�z�טk;)@'��ꀾp�]txU�s��ZhA�/�#�����~,ԯޮr�U�Rt��_�H��G��p�n��zQ�!�F6&J����]�	$[͸��kj�a��j�I,syٚ����Go�+� ���".\'�t:Ū���� U�B
�R{�l��"����L˶��3t����:Ƴ�&+�]��XѦk��!ø�,�h��L��5�P6h�(O�W��~*�97d�8���N�on���a,�~뻥T[�湷
\��+���;h�od�*�2g@ȦW	0�ڝ�B�@�6/���e#�DUz�_��,�*,�ggo��>�h�}Eȡ�OF��ʢ��6z�.[��Ƶ�ۢ4�lǴ�@-fl,�Şcϝ�t���u��t�b�$'�(��Vt�A���`$�
L{�Sb��l#�ة����1����旵����������6�/~=[(�Ն�O�ٖ��!����RƯyu6�w��+��-��ui�V��P��4[[X<�m.y��L�f���3��ֆGik����n� ϡo�ضQV�)܃�mS~>��q{6���nSj�{���؜-��x���W����4��Ma�lF�OE��S���{ƍ�U�i�4��ސ���b&ߦ,ӗ"LŘu�[�A<rV�������d���	�gъ)�L�>�q��x�U��N'Op��\��3�-1���?���EKLÔ���u`�Z��$�Bxw�"%��nxΕ'%Cg-(آ��G�! >��o�B%����`ܯ��w�?qW���/���R�]�{�Ig�z	z.�&p�#S2���n��/yZt��y|�B&��#���,�n�a��+uO��d��l���8�V�V���04<
H��҇nU����fҫ,�U�t��T���*�E@m����+��5��Vr��Ĥ݁��AXJ���z���j�!IM��MA��ɆO��8,w_��1Y~�_Z�w�R(f�ӱ�o��s���mp�!��#��%�-.,QfM!�:�d��_ҡ�+���<T4���6v�ږ�c�~JD^���[��pz�$���u�L��t������Wth*]*��[OJo��S5�sJb\�>ιy���=�_��% ��f�V��Dḩ�i�ހ[YF��O@�7�"�j����:�AX�=�x<�vVK���fE�#��\�/��ÎT��42Uw�ac�'9L�(�d �_B����a<�^�J$H�6�m(Uuz�g:h�G�v�C���%,Ӑ�tn/�E�$�� ����p9ji�rZtV�����n�y�8=���	bd�>��p�C7�� �E��8<p ��ߧ`�AA�2b��9���R
V|�C�]fM�|L;������K�GGp> �������c�ֹ���%�:�*��1;*��jٕR�ι���5|=@�R�3��Ap�L1@D��;0�_��	�5��1&�Y<��}J��a��{7,�cr�	L�7K.ް����2_�	�@����F���ݢ�/�kj�$L��X��?b�?�^A
su�A$��	���h�u���V	J��|S�.Z{H��$G�5`�@����V��|?�����{��TD�s-,�N�aΟ?hY�m�F�L��g�;�{}[@��xLx���@�����?��ٲ'�ĽH�����=+J�o�9�w���W�o+� m�`(�|	O��h_��8��-2P��'���ۥrw2�ު�7j������=w��Z~���"�+����ck����o���I��mY�;&�W���ۗ�4+��� }�F���\Q*u��RF5{�t?M@�[�8ԱR&'�~��qt�!9��嗮CO(
�#��a��Y��-[X���E6���{O�bi[7"��D<+Cd���_��g�cd�{�9���P�bٸV��%i����k�n(�n�����ڈ*�笎�4C���z
dJ�O��ۜ%�n]|&as8Z��b:�*��.��ɩ��"��i�K�
Zl�-�Cv#�g���Tc!?�"�?�n�&L�6'�����!z�=���[X�r�Y5�m�tZ�ш��w%�A�9.�u�B�A�,�J�	M �Û�`'=�VB��Nh��#핊����
��]�=;B���~�YV��,��s$���Η�|ǁ7K3=�%bC�1�b�~׊R�Pq�h�$��2���<���C�Z���Y��G���$�s���G�|o/2_Y�����{9}��r{Ί�bSC�1ȝ�v��\Sϵ�V��{���3ˠ�Ȯ��	D�}�B��|�����e���2/�o;%�tw��Qw�Xm6=��¼T�S#W����x��s��~v/\��Q�r���ɵ��Q!��^.~�m,�S�����w)6��&pD�@�a�4d�?��s嶋��^9_p<@�;�<c�C(�e�K�1�	,����#���O��k�{l�Q���"S�ڒKA��©B�#�~�5Z<��_��x�9�t�9S��e8y[e���"_W��6�$V�9
����es�{��4^�3n�s��4q��L=}�'��Te\���`����Kz^Ir8��t4�ҕ�9:��bCN���%Z��n}�j�s~�7�������g�[�ĳD��#���ֆ���a�ۦV�jf�7cov	�C�A(e�Ԑs��O
S��F���X��dH>UdTEu�_��;�x�kK�0:])w��8����nZl� �ti��Pr槽H#��i��C
b�4��p�~��n��;-^J%
T�9п�,FV8�"�D#|b�Q�B��
���Ђ�~e��
e��wA���n�@*UN���߳g�S/���m/��� � �q���6�j��ƒ�̘3��x��5��`�ƈ��!�l���p��$>��u5�$;�� kÑ
yF��䧡�v�s�Gw:y��UEMl�y?5y��3B�I/Ш0���H��_b�,��	�q�$�����CZ)�U�M.6��SG�0O4���y�hC �jA�ʹ�4C�/�5���~#Ö7��]�Pp�9k}K3r��i�0ҥ����!!{����b��;L\�Wm����W�hDUT����F�2(�z����d ���h��qx7;K�����������A�