-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
1gsg6A+lOIbjhd8utkL7g436QzUwZcknCgV0nBmVstL3mBj4kLgh72ACrbVbIjHCxQj94lF3WSTd
whdPcmaVNV2Sg5iejkYubVUrOphTYfBB6g/epljrYPfBTsTAGd8EgOpVwrf0phv/1XYMI1yHNOWE
HdasqO167DEgW8MCvR2jay8qiJNtlevX7FhJ/fMLvzTlDnUXSOgCCAS9yQfwywPCl0IBDc/6havg
rGmuNKfTWrVWac8R4R+0TMhk5ki1UzVE+B/zNhZCDe7TcUouQ0YyCchUImtswxK+0GMqYeYl/7QM
GXPs+idNcWAzDhOgqdIXwpyllhDbJQdwKweBqg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 13456)
`protect data_block
osnnTntMtVhsq9J4tw5eLoGkQM4LiSDOR4C/p3iTmZ5DdXMUhu3obGdfNOkropdQPosiHMD0M+xi
J5gzTjfhl0CB5Zt7pPMg9pfpbsZWPA9dIMzzUZASl9Zmbh/GrOhNNl06gHHVsvJpI4RFSelAjLt8
MaBFbtkL6zK8v9qg+bzUwAsEsVvXTkcqaPKVa7zoyFo1NiDYrW1uJ+MlLJa8lRXfq1/zn7TcBllz
ug5mL04Rt/xiPjlvL5prrysQyIn7TDiEVwxFuZoCLEytQyjRxzZ4lScfyJjfctU8QLyDYCeIRtz2
KFI0+r4wNj65Y61QS6uJDi/paNl4lQ+fN6XeCWnHfCnYER1ocFVFjwFLCChrfVB4AXK8324gAzXn
JH1BMDlNA5qTf1ECwETQCFdkovOY8GhZObu/zIUtYSEcMwnAxHZ7tTBQ6eEIpd83eDQKbTnOpxH5
Qvt/3GaQg+YYtkG8hfAHcvt0ISDBIisA9ROJIlAzEzvW+ZJD6aJCMWUGjHlp2nyT2nmJB3QzimA9
eQG2LLl49ZNAqAGPTjmaEL5vYtlxnncXqwzx3wfJBD1c+2DxlTckGDXhUREi394C/4r56EG/iVB7
LhEQMbbb+vD59o3y8BBCj5lvS8jF41XaPQPZfJVl3iatxFwi3d9kqAGf8xL+9IJwzmieYgUmF8Yb
E09yY2DSfsD++R5rOxrmf2IFW4jPboeIetDYke6T+t0bxtR9uPk9ZULF5c51HN00xEbiGAuk3JMj
Ru9ulbXAdX6gse2wiYsEfuMAGSMvLBLunDSjpouZHTS1FPsrXBRQIYsMTaIDmkZCPslQtuotFz5X
IO7AJ+Iv1wV7ftmDf8odAM3Hgd/HncWvE6oRI6Vk7jZB4/0+wR5DLVTDcUtotGjmtWeSISf1TUnU
jEtQE2p3loPmcrAzL7x4AZcIaBsB9nOBP5nycjzMQjIOP5zSAuJuCxitu5KboxTzkD02sPvGlzvX
taDHF2KMIXzFseVujTolA3YcBeJo9ejwor5Vr7/fCAqVO87w4KVlqX4AuKL3SvORsyBJxE/+IpiN
baJQjoTydi16919jMNMT3i0Uc/OEyHbaB9XO7dOcKovZzPiMW2DIs7lVEyINSV0rrsJf4xDqNU8m
Ccg7/UkwV4p/4EKSETptxI+Ztfd9zniXC1dLzh52dx41M4FMcoJkq8z7dE4+ej4B38HEuALUNUUt
r1qh1+k/ALCqk0B9DGez8hncG/F/A5Zc0OZ/HgudOm5fxjTcYYz3B2Q6lrVwZVxiw/XFHKxbXG7m
W1pYv/luMGZ74Wq1fJHBUVZSXAXkDNHcRHiQlHi44BYH7x8z+K4DxLvzCqQlwYxeFe0BsIG2Cnfu
32cBy4NDGUtP5eFGV1K2/LpKK59792SbN0o4GGkl8fXPbZbhm+XdohHNXk0iTWo6XOYgKPiLXPf0
lihSwnyXfYBs0SEkkMZugb39IJnQrRwZ9TkTiZO+APfCOUV9ESE23f/loQub2vFBx8z1YeEltv4Q
itMWBcZJnKjS+WwpOfYwW33lAdX0Cgj8TyMpywIEUy+RM9OKLf9LQ9i5QDJ/XklSxAT6LBSvFzE4
EpcdTK0OKlAkWvNJiWcxAiLuLygo0bD65reC80fAoAWwgC9O1WX8M/Bv6WQYvnm1bn5YYeukN6zz
EPaGr073q/cdc7EEEE4aFVupLXUgFdaxHo0pkhxkJB/b3lz4H/3Ld09KP6JBvJynJQEP4DLh06Y5
Pq32KfTMiYCKZT34YEUSkQ1vXRQcPnEh7xwTCspp8baPbbGFY0KQ2V6ddhILKPUlmpqWZvy5s7be
j+j/AtkYFQVNfQ+9wBgU0XEd2Aia2cfbeRKBayJzWGPCFAGhxdYhpxt25dPRN0AA/zQ/0AgVgEp/
0DiVwLNoLp8nNbFSHn9obZ8ydAl4x7bEFcB+jpZV9vrcq6fA12IDSkEzbnn+n0Jb4FILjuNjMFj5
+cFOXyLSF1F0bONqZyMfkbByU3bqxyMH5jZFpFS6feUV9A0BTqWLV/j8E9khuq7ke8UcsoVMMPYQ
upfYR1SL9VtGQrVohvKPWfI5Z0s9gUrO3ao8IyeAWQftnkiXyuUNAdcXv5aHKzBlcWrdYLT8mT2y
FkU6RvJdC9BYJWCsjiHZIs4vm2jFajpFLNjwA/kGLmIdLqtvH1TR5NS3rny5C5lmYGM9cKYGW+v6
isW7T6drZz/1w/o2QiAt57hTHcf/mFPPN5heDQ6wdIKaFHlIgf/tsC3/oJNCXBzD9ci/ntpB1hCJ
s/RsrZIfomv6xpx4ebfbLceuOXUWgnLpmi9dLvvWFJt5a42x4PX/HdOxvCSTR9M4CDD9ez87QfIk
5lHyDrVdcbqnq1RfcV6gN66o1HR3wSa7zk92ykZG2CsArr/TAc147RhNPKyKcDNbemp+BUdgLZM+
bhFhNyXmfsP9TPfX8YAYpYZrTuMpvnVOWOiX8fi+4ABMM+SSsry/UFL9OdkJTwvySfKmI7ydbeNM
YBWtfS4coUJRVdC6yJO0s72B7Io+WMvY4BDh9kK98Jmo/3p6Lt5ZqrLvTof9HICfZpEK4ufPWkTj
20/JcvcXOMiDij/zzYpr7WCv6cFLUsvTJBidkbVEu8DJ+7MinUnImnV4LpdE4/5x68rY3pefk9YC
oWcur+OJsUnkMf9Zps6LHelMp8wb0/YtqDvJ1Jf+M/PcwuLt2RAC3uo4A8iVqV6gmt2ejVRRvyZn
32H8Ox0Zs70xi3zVcULDgumHEB5DiPFHUi4vjGa0E++YoZv+wpLh+t+yvS1/1o9r9lxHWEcxejTu
baXSomg9CtjOcHDmfdWTmtqMuAn7hzKzyftZzL/fMo292tWppMXUUZgnZit/etQnG8ihxXZQ0m6u
D935Nya6n43lFjX7QEXxRHwdMqvwRPL1YpQIWPZIt8iCv0vV1CnDYRRFo/SRwZhh2iNYk0uBap+b
gKspsmrj6PLCZ0nciK1FJHY6e/AjyThi/nOFRwNOAyTorqw2g2RpfymC7DkrwpOhEA/NqUjWrU5l
/FbzSdgk1O+e6Jbg/YHdGC8nyILxveo6bwp3zd/RDhfF9Jzui7Ye/qpua32HjJpXMJqG07uK+o0A
j13ndHKD2SLuvdw3rRjc9rpnEnLu6IuMZ69SxGVEV++TaCVCL6xVGqXt95AJu5uVa2g/ZJzUUTEt
pDeeIPTUHDqJW6xnEhjm+84n8QAH+4CqVh5cnqIvcvd65WsoCgOegPQF6a5KWpzi/Q6KKm3FslLY
HIK0EBn6X8eNAvOlMJWxZy5G76qkqcgZ7QsQ613hQMZp0UB+clNce2JPaKCevzxqnbmv3kF25N4w
CqJDK8aSS/sWpDyyhhOM0pGJk2MwIyBtlxaNxxLMpNVmSt6vD95+6nopwadSdUYGNchiG4fNjiYr
GtEz4s+imlKeQJfeYGRfqlA7ti/1YqHO60+AQbr7U7FcworJ00xi2jAzx73GMtKebnZ57+NSY4h5
gWpn+rPVVAuDWCDYsERSqXgNd2pBxmRwhEGxkJmo/cwZfztfOjADQa7q4G+tz06JEcpfGddrA0yq
0G5OVpD21C+K5syWUZgjOTsFo+cAAw2x89z82DvBObhdx0gx0tyozRlhFCVosTH/ZObCcwD52cQQ
gTSj6CYvYpbwTzOqF88M5VpmCBwpqpYxLPLoSfLw8qFhqOVLOwIcuFnJ/lY+5yPrO9zCdscY+3vW
CF0AI+4+UPEkzs6GwSBM9BCfiGH4EpS5tpU1wUh5koNg9bnvjxAAbl8yQArT/AKWsgA1Lt68/9AZ
0EJ1elgrJZGKQ/PXPp5XPGJPQzl2pHqMZDFbew1QCIBl/tzYKmK485LtQvwFdW+sJ8I71U6YCyG5
I3La9yIIb5kHQWxBkf30LUFahDa2fBymhncECqroGw0Bg2DVbbjTLYMqgIwz+17FnaPtcFYKNVHV
0S7pLKn4PYi9qF809RegGfl+bUl9mm5EfM5pM0FIpfJ6HH5ytJilq+3X+ZIq30eMql7wH2bmG1JZ
ZE97/KKJJhnxZACsCyioZH2798M6ksNzH8/Z8kQ9Eg/Hr9GgYTTDDp+K7des6pQviYKDpNDySUHo
RqS9xOn11XnLF6iX2CsAbuy0xlrWVkq4CI3H2yaWQR3CnG8PO2zusIB6gzPTh6B4AHdIKgL0lzOB
01STn5IF3bikEhlMlROpJfe07YDp6fcG26swGbbBvLoeu1Jk0s2UkiQHVv1TGgKx51+gwwxKe0Ef
mDKVhkTpG7yznAkIAd0tdX7I2jVFFlkBB6nhBef+6HlTiCmDZy+vCGJNYoSUtlunZrFjfRR9z25q
mNJsG2Z4mupd1gcjF2WkTDNsBT7QJNDCtDWNA+Jm7PS231fbQisjT/7ivxyMbGt0ZSZX8ZYVgoQ0
puNxnGByf6gt+fjoH1UyxDut6jXcPL3H5Zesrg87ql4rdph1R9xhXksRvx0FxLJF/5A49B24SLRl
aaN81/Fshm3qWkpNDlFVDA0mzayxFH/Fb7xFvfj8YEFPfkcq0vfL//XpCkVFtU7FLVE3W+GZbfPP
GlwgqQywHODTBQ3cvL4cFy4YYr4N/QZjqKLRUQsb0QdCX6RNVhOYDyW7EQ70V43Q59QBqzeT3zoM
4aWscSTLO2fv93harHlqdCRHq507i4pgBwqO7h3C6YMNWv2t8hiKRq6lYr0dTm2YBEZz9UoomM3n
KxJ4q48KdU5vi/Lz+ndPOngyPfsKuUoUHDUJhC7+voxReuxS/lxubIT+UuozLzJIgf+yD32icb2M
IHQFZ5pyiURyrE+E++O0tU4BMcoZZ36DmAOWgCC0cV8iiHCkNBqSz8nyf3hJCf9K73urQ02xxumj
1vaxYuSLO6d1njW/tqrSbzOcC5le3nyQ5JE1z9XHgDlZ/xWqE/GRENV/jf3fDuDafL+ltsfRVvX+
8LSp5VHI9iG4fXC4SA/OqfrOjLrN6LY4Y4hiJrdgNJkyq5hwcAGeWzwHRHJAsu9BJaISPHOxhte4
YE23EZuPu4xhpTx+igw8TmxvrmAPdsX9UJ23o8AB6rPbQAhjbnOaQqLOlMe90JTZ3wf6zN25d+Zl
JQLWOOfXDemtoXxv4AW089E5hRFuozsgQMXv8fNaLUVbu73X+bYCRPPtVNPQ0RqWcETcZqOvKU5q
HwNJJBxnLRRXUqy7+o4nF66wG5CJz10PF8XrzMBlpxkcf9eUYQwk8q8CV6xoYDLc6XxNRPB7B017
wM8VYr/GMjl1TClXBoO+4z+JLt5BVVkjkz2frdX6nlq6yJC8lizj1aa6fYlllWbe0cY5JUcK4atH
Wrat+tgITd+Ui1WS8aqUUqRzNZEiMKmn6aabVx2V9Bh4dyYKrRoWZvVbUiU5OJkQVWldhYj9eQ0n
qi5AazYSUgNbgc3woZnQNJ1OT8+PqvU2NrI8AqQO3j3wHur0SNB/xhDiAjP+vTf+0Trq3hX3oUF/
h413/Ma0+dfWAPaxhUa/3uTmLTerX0TMPDuLEoQ58Xklu2OMrsraPybk6EbKbwsZIeqF/nz4PBGY
5vAkQa97ndP34uSnVrtzOK36qeOcTaiEXucHO0EsJWVjZvU2T9VHM1JH/qdUDVZqybGqqwaE/OW1
lehA8Bn3akfhWpSGrcZL+DPNRwe0POexTZOJJY2UftkXRyBHWqnmMiJOJJAMOIhNskzuc5Jk4dcm
qOKtZ1BoyGJ3F7qA/9LsK6wsFjS9QktGpXiyDBAyKklFXqgp3vaQ1uTVjL1g4km7yUMSZzZCDH/6
8QPTGw6UkfIe3855QZFXeoq0fKtc6BTXKiZCtiuRzkgePMjJI6r4ZcFbUFGy9YoxBLURqkaIu+Vy
RqJWjXWyoUxELfeeQFhsV10FAlcHpErNXHENCLt8+qlAs6IVrrIv8nmEwTgZ1oPYk7e+JnWQ7cUz
xZcFzRT9MOaxO1ZsKnwBjrzUXHAUv4moGORsYcukHMkrRwWaIcMfehjJUbGahpSE+NET0zam9/0J
SNGqmKLrAQiKcqTmzX7kFVDTOcfuLrfVpy/iVHMbvePEQOfHlvAvTLVP1+bdijREXG3P3mO7Bl5V
PRKlXZo1t2kT93AY7eveHuMvTQjdsLLCegvryNiLP2csqVaYxU+g7zOpsrk843yIm3G+dSdqaneX
80DlRnpuu1D529DVY2PeEMTCSXP/qW/zDjcn8rxTG1knoRJNYLI3giTUUNSmFNS5pGO3TfrluVy8
TRbcWr1jpb/iAoCsX9kY0jvsLZROO8nZsloYCqs4ERdTrJ35YMt3tVt0yYYtZyF/qqLFfjmkfMjg
vSR4qpFh1S0wOJuyDNT6SnT90HeR6Lazr2nUZU9at0Dm0cuyJhAXr6/r7UJL+nHxvrfUsVLYJTq8
k34vdX45YIg11axkPgvb1sqsRYWnVhrmRYQI0fJZjSzPOjKecwCieBbMrJw9s1Bgie/Cb4oN/mwQ
xr3QgMTcuTMTHrvETinmTuN9xdJ7zei8Lrgumy1Kqm993Jf53WdMNpACok+zynl9eWVODgzjfYNH
dC5y6UvSbQwe9GiKjrpTe431U+uvOKRXoz0zq38L3v3o6EvxkJYVcvZ+zlm9ZCxCIotZyrm/W8MZ
z3CD+fnbcLyAkj2Sri5u5xhdfk2tNgF5I6pVB5wZGp+GYx+JiVsc09f0cv4cF5cf+sjlaqedrdJF
CoYyRFi86ArOTsQPcLWQWnv1kTshQpIktrbnD4cNKQE4DCQ7F6lGM/JgJZaRocxwQhV/PcJGOOZs
vx5kYM41elYkjXoChsrqkNUy7Dx2pU4kDe/WdhFz01dCILkE2L/KpkDEA/2fXrdFV+cX+8Po9f9S
s+LxZZvBLOrRRaCRBdZJ1ZpQqIiQTYaOp4VBavjyFum2tejiFLwVjjqIfjFdARCt4a0V8keKTj8A
bB8CKn1v1H7k7vbubIpj/PkUB6/PNNFXfcsSe5OxlL4uPzBRRrAUZpy4wx9oMiZIbQi2i9280BKU
Iw8i358wnZ55fmIZSpSFnso5GyDLqKh18fN5eRXKKaernJ+YymkMAYL00NhrlOi0XBvPTxFLZxzH
ocL+d1gjJrGiPG1myiFIeFu5GaNq6yhulz9xmngjCoOfU4K+2MsFAQQ0DtcgootG7dt9z4m7sZ1s
mCQeGSR3svyjzY7DmOAbOTRWEfOKhpgitW08DWpfl0xCiNEepO41SO4s5+rtV7kirpu8fx9r8Sz6
Ndrg9s91AjpLK3djqgLCNiPT01L1PrAXiPfWe1595jlgV33FsHPGbhHg/R4oamW0oHqLPxTGvyQk
VWHO8xJcsuLwA0e2yok3LJVhAcFPaEmoIArX2xuGqsEw9lArBLkPnmAkJSQ6EFraJs71E62VwBXU
OPvPViUTl+7iSOCo+U1Ud1pg+340Xr1f1uxmoZKxEdWl/FO5SUegGpsp5lLFvWt7epcPjwO5wctg
b5wZEJeLE0ytKKHaHY9wZkaHTEOjUgoOr25sAbFCMMNtZNnda8Yr8JWpCsFKVyWaax2SZ9FQJ0n2
hgo74nDf+rjTH2O7hNeMZvrpD6BkqCe0Y+GEkOgfxroY3RAcQtS7BNTq/4gm/lzl77sIi8c2jO+t
AWJ2fHJ9I0KdZtK1waa9T3cVkfx9iUts7WXpkOxVfCz8V5zrTJdAHv5i1mVGzNqNFL2M2F0+vWOD
QCmKKONeVWgWSusdefvoh5wQRsE2IrrdgUv/xvDVG893cEROlK7uAN3HjLoBWCAJxhrqiSYNfAE8
6vxsfE3xSrxFMHlSNSr6hpx/DwZ7ZesQKY54I6M5MpgmWBJUnK/y0KGrcvyKNWF+MwpSduTINZTl
APuGiKO24vmZ4OgoI4i5cOFS6AumMi+/xMq9UGb/no/yDH7oh/e0MhZCQrbpFVLLBzj0WLI12Jcb
tRFywGlFbzcoeFogMlHzy8DKuWbcm4D1dF1OsJ3yqhfAWxJ97p24GusXNvJXfdgIfp/IZc1yB8rD
TSKT3DKewb0rHbLXMwwxz2KBIQeWT8qv4FsBQqasrPEmIxD3JywaEil7jH6e6mmOSiLRWP8IuR6G
GxMs6e5UZzk8UHeJ3GIDsYeq4gWeD5aOwXTJIZwhJ4U+BlUop9FeOeMTKZG1kr+vU0uFS6Cyh3Rd
/UxYGJbs+/jsiUD9wF20fw2z+m1EDOurVXBZoRDFrwf8wOwAMlEKHw/WHVCcTDeSWA79J/KBym2V
FnGgQx/JnxovgmO+urV3Psq0oe6kfFp/ahmkSGfotMBRvhe3ZsvAAaX2Ifz1q/qzNjAOUrlWuyup
1pIWUZHTpYHV6DG30nKOwELgo46BZRWFyxJ8o9V1Vlb3Pm9gIIC4EwhD2I24rdbFMH1aeXO9sKgO
fJdVyIzM0HTfJh/dqSoi+nVheEwiFqMFhr29z6KTfH8hKZo5l9nrzFMiiiQ0TRX7Si6MgiUpGqZi
xIEidjydDXkNTAhsAFW+CZH0qTL8uLaMzx1FV2B9v1HeX6przMB0htOqps1BzzqEb2lhAh1rsNHT
SQiJso1K3i3K9V5RuYSLdGlBPhvSNihmvfUYjhxL0yBMq90tLkh3TmfNixVua/pFlrftBJupZEK4
w6RW7Tjc5La1x2tsp6RNUgmrwg+4oMhJuir8i641JwVercPKSqpCVI1pr5XX1lnGmkusFAKkNoXv
QxxOIPH59YiOb7louAOB54cC1Lwc2tBBTPxUaC4mOdApq5HLipe0l6pnMydipvQgE0+k2XYLHbj9
CeSM1YVLVsjhYmwS/pQ6f1BaMLgxIB6GF5EP1NJGZrQLDWzfGd010iDJC61u9A+0PETfPzF/vqzx
r6IrTMWQFWrsOXbbtEu+YIBjAY4PfRTZPRSu1SLT0RrQ+umxQStr+zwIPAeyk+n5KGp/xNtYXItu
80W5u5oPUiOR9Th3cF/s+zPrM6FlI8s0Gb+Y2zImvKvjH6jTkj1ub9Cc+ExCRBN4NgpVr+zCmz5o
boYp9XnerswRoUi4cf+M/KuOqBev08fPpDOuUGqnXoWCdCYlKMPbPt+YePTQCQaMrI9RsOGvu3pG
dom42FPH/CAp6xo6zPoA/zejS9yK6S+EHiJBij/hlpxXDvbPxCDUNWS0PL5dYkBlDQpOSemc1YP8
IQy6jtqE0tLMpA+rG0zSZhuHLo8+wNhehY+K79p/3RfGX4EEFZPW8kfgxannWNpEX2vjMcDicJ+z
bKLa6/uX+15otN3f6AZTXELQ/lEhrhp68Zr0bdC/aOGxuYjmrO/yfO2vUVIq1NJ5Bl94/R6rM92H
4SHiPG1yL9SgB9YSeEnAi1dCZ2ZoWkctrhM3apu0uUVXhkEFGeg98NW9GV+bW1Hko/0JaHmyaVeh
sPmykWQ9iNGL+qg7J/Fa5dLBCsYOveuJVi3mrtbt2twDu2m+p+jD/MAUyw4QwYoWAONBzYcoXnJP
HTktYQDw5R5BLBawyrcyUZ3EZv06NUYXCsBhYnj581qj7yoBkrMcaI05C0aYruSu6VrL+JFJT30e
axAD+6tYzpnGVyLCNlDA+47HRkth9+L6RHGnuR/VfjrrdoWtkpwKYexV75msu2y9/NFxcX0ez/FP
ImmF37xRGPKj30MI6WpccApHjja0B1rgl05OzozUWcO5L48zf2muy8a+jNEoXLY0w/cpBWYePryS
Wwoq72ewTKzqP/U8qlZjzzGlxA+ECN9DTf+JssGM0RHvCQZOx5uTfA9qXK8uH/dthrGq+41kZTWS
w217tWL/Sd9vFq6Iz2dx8tntIQoF5GxbW54Bw1qg/W1QrzP7fgYmnx/9AYw1+nUGEHiSxE8lH3Pk
A+O0Uthpd8I742V/mgFeRles+D4VChxcDPoeG4TyXeVfiMQp01AxKND78klMHi2j9o4vax7T06i7
noT4Virir7pL7qQUmC/ZMNIdaFFNr5FfaN/iuBzvGTzAxD0yelFj5j/dxvPvMtd8FB4NPEI7658G
K8PCm9b8QWL9cAszs014iQ8Ec8Lh5HjyASglQG4vmWidldtEaKIudxCFcD9ZpIfSAE1vs5SJraf+
GVC9EXe4rdNLIhZAWgP8S3sjjBqZ5e1zlRUJl+JJFRNLsnHxO21Q5cdB+cume5slh1vugf5jeQAF
L23fZOS2rkQtCmJcYFkEehBX9K7uEFeUVa6VxmdOSvKarp8c9kNntGGwtuIoI5YlB0/+Bv+uKI7C
1EpqauRs1AweP70rykICXATittJ3SF4iXfDzX/YoYsQ2HyCQIXkllL1i8PMlAvQMrewGMyySxUuK
4ZyDfbCi8OBpavz6rhQN2b78lJBPZiPeOl1MWyyUBY5dRZwqZlzo96W8SGkXOBIXWlaI9Eg/ogm8
75g5b9B2IB/An15VAiHHVp8Zc+p0twIvOsoK9cLDjxP2LIImraPIlR4cGCj5t+d93YXNFnFFbGYr
eNgTV4tUxGwkhMEw+WuzUcVR90bxxCOLwYGd+CVK+wEY/SK5P3lYUnIu2wGzPISSx82Wuls7s73i
HHg2Uv3lP7HpHzH/L0ooQLPO5VfB/bVUcB2Rl546sUpcxUHPzk2q+btOR3ZrafCHTSFNqjT4ETFp
pOT2s5JxE+s4NSNhb4k/qaRU2MqIidDbjWWE6OeVDZRH/NA6go0ySPqVjvBwIPDuz1w1nSoER1Yz
3w47th54DYaxfSoARz7ZohDJciMGNaWNC8GzVLR8nfPCC4PvORFqGS4wscImEUo8yoD9pdw5dx1+
YMGcgMGB54IhR/+51Yvh641k0Ew71RkujIpILsFxnxSRNmON2yVXeITrvbW7ge36ngD3dtAbbpYc
rL89qZNsN9JGAyBJCq4EKIBvKSKRbXk3Hud2nkfs9OwVntBZrbvyyZAv6qju4cObcTWetSyiYPlL
lLOMLpi/Me1uBbj5zoJ5Q5R/MJbsa7O4TYNLBXsX5hHQEbRQZNmSnQ5Y7IM8+9EyQyT0TyKGfWzj
+j6Ry6s75ILiaZrd2w25MaoMcDD6LXblSwkPU4o6hU0PJ+/oW8buUBeh/BK79UtDTc7MlY8wrPcH
2A3qcMLKTXfVAaltKRCRlhCtzNQNRi7HkBGBmHk3N4SjJ1ogzKBafPDWbk+7ATu0gT2uExwg1o+y
Kfa/87mhomjDXe4gXhwgN+l5nfa5u0KqEegUGHatS4RuTozOE2O+q1fxZjZZin0IELdHxQI8T9g4
y+1yV90t8aovoDTz0UWZqF5pVYpArDOKSrAIVqcLRdeO5I8WWtPCuT9Fkt7P7V+ADoctFhZZAGom
65RZYjG8cwQr06t8PWoyARbhHgLB31pTuAlt7BMJJckcZZZEfzEIK5gQRZy8JgzvEs8NOp1uMc45
xGBG7lDVQNzhxMVrDJtHxbN8L7IL+MVc4ea62fXy18aEF/wdLalzXqZ/WsQWqeFiyu+31fxc9fMV
ezjJBShV8TIm5VPZbrmL9k2fpjLZ/Gyda9UeXkaelNtVtVfBb1FenFv+PsIfZgM/mbmnusUozFIF
1jIsdm1BMI9YewxS3p0ryXB9wJJx3yzjkLELDn9foalEoymkGBRnpFBvm0dCds8rUsmJgYVZGBuv
bft/HiXBcqzpp9N6ocLc/nuTNQ7lSD6CZoefqp4vizNT7HsyfMcmsZrMK0ecLOc7gP4dj6rVuU9e
HSd5AJ11b9yFJiNgVrgLWN3UzUsgOK8th00yyoOY/+NFK69YJceU5cHclwuIqDH6UYTHZHFOXkMN
ppyyvBXbdqc1wJWVXSXR/kKoRInhkCDIstIhN3kzI+C81qI/h0RwQOwVG5Qn9IyhtS8WHf51DO3l
Jrd+t0/GAbfWS5GovkSYSG0btxcUD2PeE7xQHKY679gyblgDLLVjfNh/8mw6Umg4lQ3bt/ubLMN9
kY3HXPVqR6F16fsyeTb7ay0vDHxRasSfZIiOYvZDUz2uk1mNRELZJpdnwIOe5VF36Y6N4oaiDeR/
hs+nNHMnbt3GRs67j3gXT43bUeTo1uBsCAzW+jlv2z8iW68I6RPDdNKXONeCS+4HeAlaw8fevTKU
PX/uLKzC379AjHKfpT68GoPOdo4Ao4CvlW3aPp0Y1khAquX1MDVJoeCkZt2eW0ZymVCBUlvqOvah
hGH9EPlYlspETyg+QNulGJ1cAAqL7Fjqq3LXbPnCdyFko3Gk0x/Tcaym/RZM/uwuw+5Dg4KzAAS0
aJiJxD8RjRHT8P/2XFQZyTY3013SnKsO+BF2CU2ldYLrH3T8GCvsKD/vMxbjEA8wdSN4cv8g4rah
BakDDQYvZMwf1LPQhABL/l1aZbOQ9wx0di1NEpdwlEPme0UhBeeZ7kp8ocUECDvqg1rtvTKAmP0+
4QD8/xSu33wJfLh8imzjS9qxrMzaxq2TYtYjaOvY0qMM/iIHJNEmW0GYa+KZV0kHmbPchgH5/OSu
AczYiWQDzJpllEAkl+UIc5RR1wR6fxz+p4NOTbLappCd0SP6tot68ZB8aJce/wGvICyKdoDTesXo
N9G0GnXm7iuovH90EPqmqrCDt942gItkLx8+m9ZjkuFc7kjF+tJzYCLrS/NmRZaq4gMZEyS3UgZd
rfTkBM5WjsVWxYtERT43C15T4/EPUXleRGFAu5bhPJiSWusAXzcBbfZxCElOlodQ232hs6e7V1CB
CpoShpYBZTc6jzPq5hS2/xj4+eCNB2u7tlWgyErYXr/BnEuHwd0EtLx2YF5WNxtLQ7RuYGMBhGRP
5I7b7P/06ReMDtNBJOMxMSYv0fk6LIXuzx5GhPBjGouT9hVJZeaybtlziZ4cW6F9FlTbwgVgdh/v
uCOGcEt8sQsLu6UJ7C60Rzp7W82K8vUtKEI7XFAVu5M9K6Niov73TafVdo1I8CZ8sQqrPB8By/3K
pg7t0Qunlayu9a8yPJ5N0PCvZjsS06HWToTt0r7bbnVVNaK+CJWLrHgz0gejQEYZyf4CmQ4ZD1Ag
lTX7elSL3XnFMKXzwDQ1pT3q6t7SUCIj0oglLrWOKuTdyJI6deJrZFRLHcq5fzLIgsSYWVVV5y8M
F8iK5KjJlLcabbqnq0jKv15OxSfKxrRm3uTf5ltBCuF1Cw/FRXdtthFZVeWYKVdfW1n0e8Fk5wFl
tcpBOWsdeJrvnAZYBiLAbpL7mAeHK4aA3ZAJCewzqU2Lze9HZeXaULjtXxB5gFOz4l/G/CgbFuRg
WRdTkGMmQoCrWXSYAbO9pIBFTPVB747h+IrQlt97JPqlrvMwPFis5vGF43jVOW0We1gKfA5xX4zL
4zkUBMjCcd10C3EoCqFnjXpdve2SEvS1U6TLW69j8SdKSEKnTgam3nXnDMz8HZwdEVrDQikteyjh
7KX8VfgujLFprPECECO29sJ0bnwBup7MDi1ojGWr9s41IpToIJwMFLv3aOVn40gEbtXfy15INHDm
HcOgT8qdUQ1S/XGSMhPkAx3gg5Vkwt8Ie9biYHzYpEY1TyUITAgvb5vNtfsVUaR3M8FWNDy4EAep
CV3aYTF/tIdCebnLZwtINPqJ+RcnK5IgAeafSxwttmO1IWc3bFsBFrjPd2bb4U1OZplzDE0ikJa9
aO29Gj6/v/nmR0869oag/RCi2/QU3B+Yvu8aI1bG5UD4l8MpoB/kcBd/itLsRA3wfkGkNcsjJ5aw
dQVr1ciX+sPdYq6n1VEBpeNiweaaHCKTt88Pu+a3p1p2zrOA7w9Rq/kqzucf4B6MdKO/E9z3m453
ppv2LPOXtmqsyRTrHsx5beABbOIvW8qUEgsbceanPcpxJSgIU22UtfjhWvt59iHEy4S0RTGG7icT
MkKbrmRosuLIvRm5ITeBuju03zppC3kzYNaobubPL9xU6hdzISnBhhLaKFsCBGtzp0oSXW+T5vq9
t3fdsoY3UqVFfZ7HEMrtC7/7F1nVlodiIjcueIyWCUPsP3+swM0Tdukzi0EjH5HGfxapmCOHck/q
hTaXF/VFvfm691jHB7P41o5kqYN+/pHioM8eOlooRlHSQtDbP1r1AS/3wdqL0y2YILAeEpudf7uk
ladDflvk5elIQ70R539qgmRYTj3Hp2vir8cdt6e1vciLtndEUzTgNereJJ3PRiWk829htItsny1Y
VmXPGEBQCmEsY1iI0B92XUj4ookTf+16/djA/POyPGErB9g4SWARa1YE28uBGRLZbvseLXi9pW5G
K/51oxAkOwu2oT3108J6MIsjnD0JfB9266gWgmEL0vP2TrWY7VG0VCKpOXC83lCtOfa07Rc7IS65
rYrWqbX59jpQDADqtZJYFtUpUN15MX7Gji9ldMSMXMCuV6RFG6NYF13F8zaVItzg8wq70hIXL7Gj
6riSHFLrAk/scYvUCtMqk/kvomhPU7NsEbg9m4aLL+dOOr0E9kfRR52OtwwZDrQwWOzsrp+R2oAk
g/6lg5alhfN63Ut/iPH2yyiud4gQAT+9x74m/W8HfW1MeT1mkhvFClt+UQGRXPVDppVni5dt6ekK
RO4I82JdnK0BMKk7gUAV0MluxNJ4NG2KN4t7fIsm/k4R1G5uWGBHeydcw+SB7hksG1BD2W79Nt//
gD+Pn86oqBPjbkBZWaGYFCWdGLC8r7rwaAyT8Z1ktSs6SeEoeEID2GgmBj6zGruBxcl/qSXOV+0Q
n8nTp7lJTLqjsj5kz/z2Ql/28Q8EEjt5QeZHCyazWuoVlyvev7tjW81yMGzQiaPonqYavL0ZFLtK
XtBY2M+1ajDEESqUwNPHKXsd6Fa/IV8eCVoA0uJk0gwYjAjmSHYELA1jAYNLd3Z3PofwLErwoyB6
DJkCtTPzfma7SNurqmPu2DN9+zM7y6UjkCKgZ4NTAehsRRRJN/bsJI2TCJe/P+q2ErmtJwCNADa/
7XeJWLOLjR8Kkk4gcHgmCTB/DdBD7lY6zgzFqjC25TJAsO66PM0N6MnLTWoW0vpipGmY8i9gC0pP
Vmde6TX/LLovrVKCFL425LZDo/moYf3GCcxzlPA5lA7/joFYoVF8iqVOjwXoA6Ck0FTqibLCMQTx
D/FdhGBxtKY+vH7Zx/d8RHehH2K0/zhX9HMCOmbQRf343rKuyb+kT6ZnbGXJrg8R0Dt1ZgQaTv00
ZduuQz9hAhNN8VIRvEgDs7ZWgxNi4peXp+BC4UrGmKDjbES6ZMx+MIGDVwVin6qW1C0q6G1JzbQZ
k+eYdoK45mQAovj7JIApHsFpa1PB73esm3iwD1+qKoGU60u6rgijJQMFXYGx7qmdHAArtaEm5rS0
Z3r8Zbhm+IQsJVuXdlz95ARNTq7uj2nEpTSgGOuU4DzWuBiBMkW4BB6QMF+kVPyuv6fEoGOwA8SL
jMUf1ACd9aN21JmnZt6UJ3s8A+bYJiVzUPNybpg28ufCLDhzxcT4Au7CCQx6Nl+mWZHMMcgId8wQ
Ar/Jocn8KOEl3cN4GPGyMNEtKBaG7Bbg3sh6ueEkBFKGLZx3KPIGTXZFa5fmszl/CYkO1A4njAzc
zGgCx0qDQJVN5QQ/1RyD9FlhBv5DIfkQLuAksRG7CoDNK40DTU5qti7k0itNNy7+REW1F6K2tM97
i54sjBQRJnLirrJ34zidH4e012MVtYvOvdomfsR8PH/gKYzarSy5sSdqL9x1EqRSSo9fneidM9Ta
RVi/Cmumqhcfk2H2ItuY/Aw9kCiszLe3v3A3g6a4WOs68baq1nglRO6XPRH17LfEVzkNkEQcVqQN
eU4COYeEIU+/kCewQXBxEd0IPXZUHea05md4zsgJFAzyTO1OPX8H8xs5Jl+QMjJoUjlA9MXiNgW0
ER2ByxOjZi582eKWBDdvoDDxFyGb7wLw8+QzILXMd0NVQujJqd0tZnSpafS4g8m0FFpp19fdCwW4
cS58fw8+hCTtyFfbfIkhBNupeFCkZTATfzRSJ/9QgaoyxoSWI6hxGLKjCKsotVmsRiX1bsisq25C
H0HJYIDKz97vE86WuW2pluj3oGcgmjqOhrdkI6VMY/Am4Ow1dRJdZr+NY6mjTiLgqRpZkZLd7UtL
a/AMHVo4OkC5WNHnj7pbdDAimaHk4KXqU1Hdl+0prn+iw5Il53LFINWq+BM35dqPFBbrbJ1kzoXt
XMuDPPsedf2ux4ehyWACc50S3yEzxmDVenLaV0NODG95HTDaF6tUgsW+k+h8IlHU0p8H4U/oP2Fa
ox9DU4OCzUG3vrMgDsg7fAMdxNrrqmyBKTZx2UUVeGM0UYKZPfGrpyqZ8i+7H9J/xGHdfBz8GDhX
d2Go8izduhv+gsVLwuz72JPXbYXmlrCb2RUwJe3grOwFSPdhBwbLLSqzFJBFfMU05I5G/cCC3p09
t3Gbjoikh5fLaQNfNkG7o5O7pmKwiuKtCayMj/trmQzFrkRQEYZId9QO3tgNTd/Dx8zEYM+pjAFn
vV7SWIH3M5HzfUZOHmWI9zwNYTehHw/BBrX7MNjf+1TT5ukubum4kodu15uqiBGP/Q+BIr69g/cJ
RxQpntlAZLCEfpew2hSF/H99kWGS3Y9kAyClfh21Bq+kciOAgnAdnNFMZZF7ACPZkZnyDigKdxKv
wjoJU8D7slgnUAJbiNpR09PGaEYmGjsC/TYRehe5B2VQ/5bbd1TFF34yuArKMtIaGhANnfd6zQN/
5dwBiYFRGPjkchaMrJTShLfl8J9xDCsuiBRkh/M7u02Yq6uTv/zVIntytvpzgJ7WMQx0gSMgNoAc
Li/aEfjnR98w5TF7CRrUgJCNhOGbgGQx+qDcCCQXTBSB+ywbAucY1Uh2oy3gyuoDOiorNNbz9f2M
WzKs4oDSBeWGTEZcUcLjN2a9KafXbRWMU9vY2Iu/PFcZhClSbENqmPAM1AgzICrVAuNMLgkiqrO9
I3QTupANePPIJ+LK6Laorbzlt/pdk8b4EowbY3TsvVhXDscwXW82HTzA/cJeFAxAHq1Ne96usHSV
yc+ZI+nFEGiKMcyrxIRSxdMICpX2eetA8w1XJtOOTQKGAuhLA4pmwi9y5cnPfIG8IrmEAXYI+K6n
qYaPBh3fiQrM5OCm+ofmcpvC35q/VdCedFsczpsru4eJUEW0Fpq33daHN2+IyyVcnNqiZPbfAt4f
Gd4j3I2HkIoeuGEYnuq+yyb8od3aiUcz+RLZ8eMSN4zjdGkLBMC575P/m0K4C8+8oC+gzuqGbxAu
a6dl4qpGFoC0jEyd3CW07fPu6W3ivpDtLq6v1OxEbx3E8XujrYnt6QWMYCVkGvibZPWA3Dxf5DFe
eMCl9mGFpR8BeZJlk9j2hSaiyizoiIJRha8r8ZljPhwtkjECqu65jkZfr8yUz7EWaq5zKRDSioNy
mnP0a7Q30hiqZYSP2AE7r9b9CNzajyag723r5skf0y6lz35LozJaon4+ljnoEDNw835E5+waoQnd
XUmYB7akygtNpVh7hKQXvCploF1oEMDqVnZvN8Dy2yoBAx4rPCScVpAqgJ940jK7hoqeoCSrfhJJ
aCoiN/sMhhHbB6+QoHDGRu3D6HGjxOmO7yxdRpSVLxgUrXnmIyEmXAR9sgh3jlF4gTMhVP1yaTer
clZf9E1JPPb13l3S5uvUJxPY8N8Iykh5xpDFU+BlsvhXvBZqgn4cbQ3s939Cr2qLx1C6xhm5kRE4
hMemJSein18CywRMfm8+k6su/zxmB58HwnscLdVDTHpxu4DEoqDmJCOIyyRTvahsTE2CrSxTxr+I
2kdNpPE7seO8mGW9TPbaS+nGcFA10mFnErhmqeA29PqCD7cS0SXqfc5jdCz8dlGP0R59I0EEk/Y0
zL185pHMr5ArGi2jqIy+WkSIGtqe65iUG8YxlZNf4HyA4apWxmEwMmIXE/TEqvb9q1JmbjSrQg6Q
9RcCQe7Obwk95LXUAU6VVpOhkIeFRmuSv9Ulc3dOmQgkgbxVoY8r5lxmJFq6egN7mGndChuXKO1z
BV6zwc9oMVVYKRUu2JPSeXgA/MTMHcgh19lgTDnRKENU5e2Kj1XhlsxbcO9EAcOz+DwBfWRgriqU
FC6T/Q==
`protect end_protected
