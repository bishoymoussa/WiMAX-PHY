-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Wdgu3t0otr+lgWZh4JKiMitD4FPzlUzJVxpFdALUn5b0EpcV488mHzT/qY+F8FtxamQS79CYTuUr
ASEKQyrBAE0sKZcqnPAKod02h0/wZobZWpskCmhqgGyHCAvjNE4fJozUQiTUiVXdhEyKy65IkUe/
L3TovF/CM0tWeal1rR+q1FQI/sbJg1XM8rHP3l9W3eG5mS4EWVnoIq2ybDSH/6M26yvMRGk8K1AL
KniUkHt3UGd/IOdmA5MXU24dNznQbUVQnmfOOHyiM7vDcVEiqc0hoZTaQ8onGO1r6DOp9g8xgL9K
VpSqPDHvfjws0E8HXJi/tGPrKMjM9DfRefFOFw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 11952)
`protect data_block
9FJTyMR9KmU8DXEabVzj6YJWWca6G/Ff8aKQJjInJ6FBgMKRr8z1K+rEC9ElPGW4ushab+62EdJH
dObXll4HiRl6zEDJYgSDAqxBaMYqLmlp5+mtbZe4E/jkNhmOicyuulaB2IYV95mGQY/GRchbOAYR
k+GUOv664go6F/RTE51f6TgNMPi9OdZt7QOj3Jf2nIMFF0aU9F6TZtLYUkIoPUoKhQqimSvbN4Wq
7RZkmqs0eOOJ/OIvOBJzhBAFFe66Rt/+q2/gpOBRucFtt3fHMDkLXptFQ+6v5ifwODFslI9mNrIf
8H/Ni3Ev2pjEX3HNtfRrcZdfn0VdyeextkD8kK3b+ymgsgG6XMv0PeZ+pz2lTeg73OR9C4nzQDey
f+v0XUNMhdp/BIttJlphPBSzJEEZMZXBxFceXdgdWJ5jKUE9pbyuA/icTFWFN+6HCXxZpuKOkdBy
CSfgo/cEHxaIvHN4TV+bac4x8fzuB1uSJtROC5m2Pc7Xp661QytMLy+JJIXvuTm1/utafyXZry56
2SSmCVhindxMu5GGthJNp8tXJptD9gYZhbzxY5Nbaj/MI7aR95mOSy/4dy0nVsLXkZUzjN/6PJSQ
kL995y9YqlOQOcN+5c8dJOV5TIyRAIcQU/nLSJJda6xtjLZrEoMId/p8l3EOIyrC5VKvxf0MUQbz
Au2y6sfSs9b96LPK1CmolS9iUZjGTjiEsOx5PvMQ2X+vfyIwowjcF8Ab7JLZQezWzVD/eExqyywe
8KdhIrqPo1qmQ4l5vsZtR7ksYkJqP4yyrZCrwhQhdfwB5RizlsKf54R0dulflbQiyhWlhMAGGG1p
kSi3TUQ5bCAPUy5n7ZT+kn6uMnhNE3GdKoM9jbUSFAVCyruiNYStBGZQdJ5EWswp6qrpo7jdal3u
xMEIjeTjIbaN/IbIkjCZGrHeAClPESUeQlULxM8KRtUvAqu1q+Ox4fo+ssreo3pKTFmmkWYffXUP
yiP3p6dF/yX/PqLSpPF3fwTB2+lkRCMYQpmwDNs+ZGWYRtbieubjiSwiJbBB44fwBRQBWoSfK62S
fi+W1/KH5Snv6Th+HQo3489zzOFSBXjdr4QGrproGE+yisDeuLVmB9sWtZjyDolYZaA5kaK1qi8w
QfrPEPX0Wo4NEt/XrB3/Bn2IHZdq+D0BqTFsRuIWt34eNZkIpIUz8fOg6uedTtVK4WgYcZdgdwkS
CHjG0GuDoUuNg0IQP31XkpLvrfVTZVmzkeObEjRwdXhDxZFSrXS8nyPHCPdwPzmANHDeK/qke14t
p2ZplwxaaeJVIQDik1ozLQifcGQKgNvPjTPegEZLZu5COK5s7AzsCOxa+yl/Yhr5U5QxKVyzavKd
2QoMou7FmYDu8U3rswIH13fxy1bGdTVhJ0H0MQ+YFlwCKFQUoKXm+2wRT1fhnLy/yZRmMU0JAcDV
Wy+LiXLhF1f46d378vCf8PhxmJcskPldiaFQFBWGsBC1uDQilRSQBCuRJS3IKtP6wBf52mHChjA5
0UcHQOBnjR49U6XhAz+49VtpkwFAijAj7D6dYQ1nAKgadAvn40shqntiaS3uL176YJiaanGiKdgX
G1yb6KUrcpaQy4mw4rhQLXN7IM6YwEpSDq1ibn07ZX3pF/Y+bc3ujAwZ+eMtbMGWRj5WB0iAf33N
E0iI1UMhZWZytCXl24kobvTexbp76kgUljJrqkEoce9KXnlQG0bnDyZtW431zY0i6VOkB2nmHdS5
Pc58qJ4q5p2xDTJsWZaBrHFlnX5SNdtAApgpriGrB71pf+7TZkWl5wtRUAI7pnMA0cjwg33HRbYl
GlXx+uq/32dA044b5vDsOyMCd2CegG7t0eJr2uPyNL+ypDspoqhF1EE3pSZwUSnmfiTRgAL0AFxP
lQ2YTWK2w0NRpApTFh7LR8Sp/jmOXgxiNFS+XoPga6gzUho8I/HbXOiakcO1jVynBdlhrtQzfu2v
CGRPm80bPbYKfA/Bh3TgFjyfMgmxNm3IZT3l7u58dd53f3O9hLblWibDUDuVtyDobgdPlPHsj8O3
2STTx3wqBgW/EKokUsnMyHzMBOxoKkGknF7UiEZvgL6+XVolCZkcb3/osetnZX/cLsSsNEBcl2TV
gDXex31UhDaPDIJN/deqlp3AtSV5v76zECyZ2qJrFBurJzqgMRyFp3C6ApkqGcIsFabZBd/T+scF
8/H7nRLoCuHZJYVrS4emZmlBDEtNZHjC9LG6yavX1Iw+sZsFUjNn2ntaC9XLSrwAIAJJp29nmKah
VGRwl+Cb6fb+qlggD2mhJf4jg6B3EkW71on68yVnVIajRd1cwgqM4ZawpvlE32YrfLddnyppd5Ut
ROXxkApKCxEB4sc+rvPPCJRkU28/3Y4VJTO67s8n1JUhOj0FK1ae+IjT4g2dKYik/fYsihp9ilez
gfmIAYcfEw7I9rv0Z3EFR7IuexJJMgM52Bw62CymTYbPwvppBVBZXZ5gpzqkVjgRsgPqsrfSm5+Q
AX4DqPNu2XLTILRzIQ/kHUsBBNJm3V7RPcICc9oPC9tGwyEoFDS6xmSUosk6fv/SHmuEgiDJJEe4
W6aDbZ3mbjsKnDieDPrjpM9hS9k6deXHiTQiyd5xrceLBge3VgYLUPwDiWYeFO6AiOBy6dc9Lzb7
EpgRQ/hxKS1D4Ij4GMVg9hofZWRqnk4qQYw4Gybdn8bYLE4xQeL7lpM83n5Tf5xzExNYkijvvY3m
exkZEVDcgamZgE7WnXdQMU7ULfdI2jvxmGvpsddM7w9yGaRhWum74jxjFu4n0E1xMfjU04kO5Ssr
JQgbDHPPtTMQ6UuqkecVHkXPHEaDXEmNNdoX+6ZAxK2VqLE1UwrPvgK5ygQpyIQ2gddVNcCZmP90
g8m5MfumJpcaz7tkmwMg+k47SsFMT/kOeJawRgGSh+8pRrkfnib5uUA7Ue0QfiY1Rhl1w82n6la9
iHsqe893wUs8NmXJiizB3UVanUYGF1OlXr5wHZEtl+gbf64hSX710484kFIdDQtpxGNK7bPlfcc5
gkNinRih+VQHuSihn1AOPxYanj9xN3IlobNJeJwCD+ZXeerrTL2s8GWZ2r7Z/h3HPg4XQIvYTGW/
QW2R4kPR9iHAaYqFwsIPtLuBb3RJw63E5LWe3YGl9TOiyWbCATmSoY5OY212sff155G8+abU318I
uWi0M1zYATHP/h+sU3dB3kqQijuNI1Qu1yrW9NH7lz8jGWdBVn+tThdCzBQRYtM6MyMbr+AvRi6p
7H1OVBfXgGw9UCSZVerMbDo12NCWbAU892Q8NPLLQwpsjFqrkrNNC0/wwkZxbS3zJZBcJvq75Jxp
h51gHMU7a0DQnCsyEajeNc9wr+cK3mBY1J9lxJf2l6vXZM+mrdzSiHe62jAkufkW7bJoEuMQf/pY
mRuo4KNBOqzP7BVQhX8oEN3h6ccyIxNQ7dLYskqjIM4DoPmUZV2/wORKATFUH0fhtO2GdDnjn2vr
7hOFgveuP6VLbO1YbRJ8NXA/+QXfoj8ADiaDa568Qi0fpoQErq2BWw1ZHN7/21flhEH967pry0HF
p+bbutt4LiyGaiFWSxrmw9u4WXXNNbpT0S6HTWnKzgFrkIjTR4ebgn4oP9nWd4XBU6oqHfDV/r02
l5cPQ5KsOGM4oVWYNhknw3MS28RLli9KsKzbwqV/+g5F7jHZx0sz3TZ7aEaAu8n8MgcckGHYX4Fs
Dr/bOiVZ3/4vpcSUfQ2LJCefZf8czeJfINH8q/E5cTw9jvsveJjw0p4CT96XRnEBaiVdDIE5lFDP
Td4r/haGRclFEb7zxXOhfQ2Ndl5vziC7twihae5CS5aASKAmljMSjLiJmwSrk1ePyCSavkbKuer7
BWZBTmkmKMsPGHLlOVlxY7iuflJpJ4Cy6zUcKCGgTpXAVLxQ4AiV3P4OtzL0IPmElgSlS7DX6OEk
hHV13Q64ZshUu2sBqg84xHCG4D61Hd31IAP4MyQ3lEdzo8oa7c7+pFWa/azYa+EPAR85rbXuf5f/
5qFUP5EecCKhtfCfV1kORrq+7pTMJwUtzJRc/pgB4yHxe14DCkJDYwCWuY60xyncL4T8SgDRxxVu
nE2tGe7TQ50fVPuszwTZKhDW4PDdXQiX9kvC60AI2HoKgSbRgxR7iqoCWM9FU6NRba/jVc4QvWc7
EEI0BZgQ4A43wmgN2UFcUHl92lf7MuiD49pnoWINueb9gw82XXnxkfAYqvAfQMm/289kDripFxXu
PR5nwOXpG39ZxjdAemXWaJLh7noX1tzaO7DPFOhpVJfKBn8S5uvim3zJlUjrWAYVGmzdGAi/apDA
W54sH3NjGtxyjTSziUDJd0g9WCu2p1OiRRUfxz+Kaolr2a5prWvYCzzDj3W0Win/nHWI6UEnxXGA
j0COm+mwzsE24B1/wPU4j4mFTtmp5+oxLUT4s1ncHwtd/ZKsKGWMD5Q5HZxdPwuSwX7KfC3K8U0h
qPmNFhtpTEVC5qM7HaagJzwVTCLuCqL4a1q/XpFZ6H2tEgDxDUxksKEjAaKDaLDsGniKkdWsjdnj
arW9IXBkSboFcUvZy1H/JVuKlrm3CKWcuTj/sDfytx2zji4c2ZNbyT6Km/pajdkeGMopbBLIinma
yrhLh+aA9ZXN+fqEx9IvxHam1yqJn+qPLWyQ3wr2LAx6Dv20MWwx7n4QFpI0j1R+Qy7Q9O/6L/jj
M0PAOZ5oug33mgVIJWtPy9Asd20E2s1/JE7MU+bGE42IHLBKtkYFRLK99KtaRNGak7PGX8F4hukF
gryxmMjV2TIrAoY+lP/vXAh9odMDsyHg73YbgyHwOxXGpReZUzyGVEHjpNB9vvBSKpAfQasKO3TW
ls4ViDJjasakX9rXD0UGLwLpIW5WqG8114BZn2ePp7dw7whkj/tt/X1Mbn8LxLyyBiK1QHql7HBt
l/LXdAQX96gerefA0OYS2258gC/ijThj6FLolrdHhDEB7xOMgcOriUS9y06Cku/lZLboTMjSgu0F
mDm7kbNskweIg0DFgG1+FWJlcqW33W8y0eHGAZTUgcheNc4RvEKy/7/w+EUD04UFRPjci7exK4kV
Lzr0MPf12CQizjl9z/d2m0dx6p2NceRui3E7VCYfi4v9sglm/HHVI2JWUD9cX5NIGly8ZCo9A9jF
1Vq0KGsJkuhxyJwPA8ywf/ZUqWQAk6RrItZhslcMx0Zm0jLC4dLZt/TcPeaEA3JbE1crGfi3xsUe
LwVc2E1iaG+qcG+cs8eWd4PmSUvhu5DbW7559z+jVnMn/BwCEX+oeGIYAWiGK6fOiaFXJboNgXpL
rSl9YMeaWmhk4BBITeF9Tt+oh3yZVSUY4par2jj1ZiFjQx3z7vh5YZzLd70p7MfnAR9n80t94K4g
NRUtTPmINIh7QVI7xlF2fQ6x/ODmXSTQaCpujWG6YS/psSdKQi07BKomViSCGJ/hMtq6i+Dc/eIO
0xsd0R+OSinggZxvKh58Mq7u1Jk03NjN9S6Mn37rd931XUCdvM3lw/ubCBLm2FpcmO1vhBGLiZXq
w8YHNbATROvgCkJbVHqm1QtA5EVB/t4F6EZzCRzkTIg6UarjhStoAxmzsYza6RHOFiukEissMkOV
jBMnNwiopfRSoMEkHS/tl8jEeBoFuZUwC8Rr0Rdi8nyalo7jeDUWr30+lMpjleu9mydfwt2qJj0p
SSbdSlip7nvPtWc4srmeEhkSAUXe9FEQOYaeWKXmC2+a0jXOj8u1UUCBFnrHJCl3id29gxKj9E/a
g/KUJi1J/F0TRAt9hADLQGe9ozIW5KswHRFRqxvCP0RHTU24ciRUsjuC9FRc+tsPQzj78sR2lcuX
LO8YPvwu3wMtj5Br3gz/tYQkaGTG3G/4uWadWK5EcAxRIUnQn1AQHc9hWPlgSmMrRMqMSII/HSme
jg+EweKMjZOw9n/xxajS4IE9qQu7E0mHbxXg+GrGpsZovom17BvrfQS3mO3wkbJrpH8lpFwHKh63
X7/lUAIXerR0WxM1wFVTpsqPBjEVO9EZ5n3agSBWIBroae0lwi12Xg4xmINdK8c8MttL9hBRCTxL
oorOZ1s4uHkeKZI+c1L9VlgLW/r/H+CU0VGcvZtyqvI8lhkZ9/AtpQY3YUHvAc7ZHFoHWFQlew9y
dxC4lhXJJFRZB6KlWS2UJ9OsxMuQZqCX9D0wXFjukbEP4+AktHK2qpe6r6KMOC9Bu6Rhcy1R5bez
wXBEmYky6A/NTmrYNyRk0Zwcw7RHISJcxPQQmSHS1fPvHtPadQyZgeMKtNDY4jAVjmUKy3R/rWT4
nc8wgYdGp00WzxRTrs4sFk4cCh06zOumTIb1W0sYuzVQMrE+uFHxl9v0PEbkrRMewjPnc/g6JvOu
QLqGpQNErsO3I3kSIthCYpVMYASKAMb8wN11HSS8au3wRTTDzsmQfPLrINaIAVWxLVCW/8NWtOsg
DHSUZ9C9bWkVNhVLXQND5T8zj6r5VrnADj/ZerHhfoYc1aFS2a2uA9JsC0LtYecTO+MmfKfuPBcP
XQTqP24SP5smv1FpKAsPva/6mkVnpU3Vkd1kuGVhDNNWxau78g2HhgYErcOvSCWliyEvZp0mckwS
HDETCOuAc9GF3JHyt6mB7/+Vq+LzDzKoq8VU1Ioa46BqnZ3X69mLgsjDtJXbAuM5Cc3F2bzCHz57
Pnk4F8WCyiD5e9ffwxyLirmuS2tlb8Cwdjul5J3uNFgFQedN2vO/SvM/kDtHtmRytDn9BIOERy98
GUCe7Wn6TbP6rSXnSABrqxNeHDls5uemrXIVg/I42d3o8FQkVcYf4pujEaxLkaHeGTaT4nzltCt4
kizAllTIxhzPZANZrLp36sU5n5I7VPd5Ctw8rTuowE3k8Uc1sEvamGrU/CVDu7fUK8lb5V7Cm5UZ
YaaSVSZt+se0t5X+p0ZZPWXKkzO5623a7pdyTMCmzhaezf3wmBPW37PAVJJKCMlux53MtrqlDVHr
WlrmHaw81Kept/4p5cBZ3d/i+0/LXbmN5gJcKubi4/fWriATelI5atF64PzD+pOXvRKL2E4hIeDv
ZlvXB8XUNUCh0ueVaUiA+ub2PrN4iGaNOjxHtpG+ek1LwNYG3gl4I6kmYjijUy+nYJhhycJeKk3g
5RuJx+FhijGWefaXPF9Tfys3mRzRi2RsxxVzXKockqX7mEjiJIPX7665mtuxRfejLPA/rD52xXuS
wIrs82ROAuN5RKl0bK3G8E1MLAGJ5ErWkvpMzMvPDd0XhaUMO4uERYm/iEnBAKcPUVNjmlROrVLG
BwzFHGUHkRmKd62k53J9uP6/3OCWFhV1OBZDsHbjaZQ4WfDzDykTUUMT+pca1bf0Nf8XZ8NmBRvN
ksEiCuUdN5y3SNNSTig/WKJO7PaMRqJiAkxJMw2e6tRK2+8ilTZNfjQ0i2ntANwzrIzGX4juYeko
FdzSCv2LjYIPmv/VpxyYqDr7QPcwVTlnVvPT1tsXgR7cNqm6nK6nqugP3E2xbR3VDq9JA7IRqN75
EztsinFirrAuknwlR6rsYN/K49qHXhI6QwMkMPzLpWOgcpCmqabiQs24GXJJqafHjwle3HYtNsi4
pPC7S5Z2Rx4QXbGS331RKtv/EfcFx95KE6/qfrJj45UwwN8N5xulB2I2MH6TEAOZAcuBKgO5QpK6
xpJ/ykVS1blrpuhurVpmW0Gg48vw/7IO8N2onU6Lz3KP0gZk8bNN/wYo24lHXcDU9oGiYaDxDRoc
5ihy5v78BK/apdPKZJPZO69c1n5CT5hkTKhqXfeSsae7gWYWzmkV0OVaAYFVGB5kV740SRFnYa2I
zhFuWDJZht+8ze1Nm99joCSvXJ6I9WhUD9rNgBx7LTeQZnZYoevRhkjyFVcmXcp7NTadIsocPC4I
V/EikzpxjeAoA3u+4iHpzCKZPR64/7EIW/4azhNGivfRBZkUk6vnkehN0Rmn6V3EAiCsMUsS1noP
4BHeufnuqrdmLpktyZy671b5aazRhxm16qOHM+VCqR/PR+odTW5tYXSKC7WPM/Eg8FlonbQZrLhy
cwkG5zm+NuteLRaSlssb7+1amYuobg+uHfhjLfLsJU8B3SfGs5mrEfncCsvi+tDZmyKKLcJaCXWf
JY9xfHhnk4DIWa3rek/UilSg+32UguMIIFCfYuwpwkCUEsuIF3YVlJIqSA9Hji/Tm0cShzwZ8KT6
SLdXYTZFi6T1c+WxSj9vIGtMyVbrtuNALnOM4zj+4TV9DrU3wlg4CcfiLKk3dPGvDkYYHAZYN0Fu
Dk2t238soIqg+Dzb1xatpdivvmqPMQmutNxOfgEseeZk410i95Ub50OfKKb7svfuqlGX8AlK19cm
C6Nm3ymBWvNohOtNhT64xBSxVfKNTXsHx1oDFfr2KxZ+fMJscJNHNcs3dY9JwjhnpgS0K++QUBsY
GYZngkf4MyHKVf50pFqqifjRFA3vn0qzcG4DHetX24N2JG0BTsXzmL1hqDbPhmLoKT7UG9fJMrKd
fmhzRmyoS/to75bgRamh9msZQVA29RjotO9PkN0eb/GBSqINKurVwXJuojRvfS9boSphrf8oVO4k
GHW7LbkKCg2i4+nMqDUw8v9eIHi0iXgwxS4BjqD6zFvj3Dd4sA4KTbDYger3UriNvYj2EC8qWstf
V69FCYRNJyg33DXS0mLV8H74iG7by9jz5vMV0Yw4rgp/3Sqfl2Exg+xoF7j6M2CTIBC5WfM3BVbU
y4kZP+e4cTEk3y0OErBnvCCqZ/hufJKeoopTXAFsEH3fAKLRe64owH6kRFHQBjrunqTxv2nUyS74
6OJ3Q//qbVzjjnscwxjqhnRgT19Rbp+l/TNo6kXbmDmTnx/LnXMmBjP2kso67s+VndejCysFNhXb
VrB2s6jWw9SnRVaP9/HZrZngezKsqGYyV/hBEuxaw8MVMMHHM4P/SkQAUR4jJVPXjMspb06UyxfF
gLZfOGvXkgCeYMHN1Httb54Vw3A6N1BI4JLdY9r/IjRqZQDOBxjBTqHZdtpzSMkOw6RFY7FMPnmP
3+iuq4RLJHIoL0WmdKUUl38bEDblzwE/0GMqkE+vEG49TtKpE3gERUb8/ngVxFGG0LlPrN0lVllG
olaI2QrxkZacfBod4NX494GGnG3WoBY/9vCJyCIFCYduNUn0CNfhkhqQd98SSGor01rFyJzHzc/L
eWp2ZMpG+B+u3lORdG033V7yG4S4pOUwcTypGJxh+uOg1OTwQakjSOfG72OX/3fXYQZTM0MIL0nz
Rfhw9O3GcX+xQI/1a8h38GVnXPk/SiDPHwAPqCoGTPwUBd7PVQLAjjZLogKLPotuPw8XCtUTLWHu
sqreBzIaVxqrXW8F00fyAat+LJNsH1XZmQCFu8vnC5dAmcWLYpTmKHQ1uJT3iY+qmvWQRJ46Lhr+
llyS+VGRM6Kez9Ej35f0IrXofB05R0or0++j/54veYpOqCvnX6f6qaeHWCfY+yX0+KWFRZEU3uk2
FjN3Z3x8iR8GzCIV4RdS8zAXUKdKDM45Zor98Y32K8qOqbxgxffJC3m870aU7KoH6QJYHPMGZaHp
QAHYGBbRE2vJd3K8YFa0T8ATD//DRsIQpLSXCjODqzobekQuSeLGCSP6XGbuWYDEuCaRXxiBxzfb
tSGIY9WYih0JjX/jTcYP//Th6Pb5ZWX5ikwkbKKgqdgHfBjmS7qAaWHql504FtCQ9Nr7bl0IM7OF
Pe8v3PJzU8eyvEhg3b/g6++EhQ7sW7fbJiHAkDjE8wnjPl2ikrEdragZcdwK1mDwZ1XIrVOoFqL+
LnIRvok9+IQpBvDkIc9G84WDkH5EizQF2ol9dO9GnRZVMy17mnjVgrjncHP3t54HqAB0iuBMaH1S
pD8HVcOMEb8nXVmEOu11iNZrdxOztoihm833ZClasf8YGPJLx2T0W/u2bWbeSs34PoL3D+Gl3AzX
XT2rspD8+z5pbxNCTP2kI4ialBpSz8SmbNQDDGel3npOaBivE0mHe3qBlEWSbKovo6AUqM43nDjv
bsvAt2qjKlYKln6F8/usg3APQYkEz/32RUApoQclaTP2G2UtSHNgWqwxCr1gFhpgEMy1VIl2Ed79
UFDOWKyYqQpLcy41ml/DX1k2i4ibbeFrtknOkNyLH+ptO5F9/duypw2B77DDkQrEMzhlGESgu3IT
HDsKPJkpqGrdf2DJ8x5ZUsSE8pl/I5lqK0Vj5NybdS9gG4OYwZXjL4ZZseH8nyM9B3JPCV2u01h+
Pt5SgxtuCx9k+KH2rwT+lW0d/jQf0ae8O5gVdbJeqZUZNz/z+Qp9OddHR6LYBXi4LNxk7Uqws2G+
0YhNnykptyANJEP+qX2FxkXRKIu5J6DdX9tSWRArSQ/EjIqq91cg9YoTibvkM4zKxB34OR+1lwpk
GYmfl0r8TkgsdWtMWlUuMlCu2R0r8Tcv2vRw+7cJA7v9Ui0WfL83fipadAd0j8tWfbTVXoLaVGtK
pWiWTxnlR16zY74Po3XLt6uZ/X9EHzoedkwn1hhWSsz4Pd1mTrpLAoS52oum4vVzuIt3yyMCrRva
YzpexC9sjvHQNSiTFdTbpI1RXdEcftkODyag9I5luFG04XLV8E1xfRCYxjM5hEqRImNtNwn/e/7r
V/hyjggeHlo5FOn9J7g+M9prgwkAwUPIXesTU36A6LYnCtC7KEFgNQF4yPmM2NNY6kOqJ+yDwxXx
TZOmMamKkUd59lxV05cA6110oz+Wsdy5SaA2kCaKBXxEy9BMPB3rlbMEA4e8VfubrYlHKhpcwWnu
4YM5WHaEPzWR+K6i5OzOSk5VGb8/Mkvdsz3EQTvDSNJ+6LDwKuSnI1qD+qsE8q2JaTHZQ5+13l+F
J3Mp+e1N31VB8OvhW+c+k+pj9eq9jZybOBxuA3ZXrAtH2ClPfFEMjXffdVV0zYZ27tE1N5C6+xvf
L20JtRNJckzkLpAwAYs0GJfThkyBeNslNEy2KLGlIYeVWN5mZjNKca0RUwfFnw8aPXRf0dBwMrnu
o3OefKedzlix6bNrVXW/WWEQngXCDtVISBOE+5RifVgyqDRavZoEGKZEY6n3U9HetpH1iui3IuSx
PUcvTUCBhmFeNNbb5H9DOmKUpD7BCs0oULswCQQVvJlZpDCT+fx/KJhdG10iMU9Oraj307rDXnTf
z3NNef722MA7jwFf0L4mqF539nDRez5l1eRraEmJUzfxF9GQpNScP3xOK+rIVliA2BI1Uv44+PnB
QYutkaXgPqLTzORHkhB2kqQDr34Hr1lzJp63JLOJU231kSd6GDIC0VcZNH0neuMvW6v3FrVyDsLW
haJneU2MpwBGC4qU6r75Wd5BkWZFHR/AdwrW5zRAQps3enWzC66y/4gURqD3RegxfvMOzcp8JgrZ
JEJ3+Jacua4Vf6Q9D5RyVVhiTQkHYPS5+qgiBLtlGyH1DO/XE5hEW9X8lEj5HlgzDsXK1aI9SaI1
YNdF0dbSWYfTTO7Xx0JfyHMaNdEnkuovUGmvQCwuK4TycGZYOcyuGSxpLuQdFlLzC3/XoQo66/9d
gb5JkG3B/PgpEOGAJOO/eiRU13l93TScbN4RF6IjG9ZDcmNHU1tSQSzYFRQflyalzq60pLF3uc1m
TYB2PQAq51tnh2gjMtCT4M/If9hnMtC2yKW00kHAH+itl60XW1/XkTFO4lma0z8GF0A0cAA92DfP
tHuiyeJmG7Gh/A16uOaCNWAs3dByrRgvZVXvoECaQx31gyMWk9oYnfx6KztVYYO+Ogg4uVpfeaMw
6n3kkm7TpkcYitF1h91OyUoalpT82TWdzaypvAYA63AKVBpUypYllNWlb/iA/o6iN/OfrcckUe59
ItfuD5VaUGrecaArFuMIMgsa5dt0vwcZ9Z0wwAb/Ylo1brNiYblhHqIN0ydpF3pLUYhb0O0tcU+j
Wwr8kZDvWsTrNcKL1oQVP1ZKIzZ1auoUH2gOMDI5XbNUTC/lFqkyRxlFP0VAWDyzCUF2WmH6YZLv
vZlv8P4SoY8weznTtKqNCzRIzp+u8Q38oS2j58o4HAZ/Hcz+EA4AXlWiselZ3Dirt7nWsZCdE3E+
t3s0IFohYDlNoIocJtEMTyArp2pcND/Dl2fQ8NSUDRAX2QzydL/dY8bod5Tm4uYYx+X7Lf9W+Mup
1+lm/PseLtxmTOdp3S1dyh9jm9F2liW742h7SEfR/RbyLvylj38Vuxg0lS25Mpyr6A5Rivw+y0Vm
FvDyG62JWOF3k2KMZdhCd3RgpnMPSurIS6bkFvrSWhQIiAa0vlrIqEMMzGExxIsYqGqvkscYDgUc
Xe4/8cIVHN4uXeUSrBsNalzLIZ+au/CCCYdwHtaHeR3+HSBldwxvQl1SxGeLqKbATh6H0OSEEjG0
lJLyNS4v7/BiNIviUnEOvcsYh1WGV1UuCoJ8SoOO+J2+ntCHG5bhOfxzzK1Z8bk2y7IFjmcmDH5Q
gZq+q1vZ/1Kvk7gOD5FT3Sf8Cz6QmCy8q9RPucu4bx/TzF0OlqOL4r2OpeN/Z9PkSGwyFs2VJfbo
tMYIP/nJC0czZ35bL2e0STex8biAql+FtSAB5NaOse63unwGqLEyczI+xVIqQadZmTGf9VBm4+n7
VbJWiHeLxdJ6+UqnB3KQi0Y+6KsKEl/Su/A5AXxT09PF6jQbbc4k4o3p9fsiK/5lBgdmtYFQTxTc
xEk9w4PQ2nXiTie22XEKtjQSLiHE0acqrFGYLNcOjL6jSsPvq4BSjsJ5han0OLGHscLGAS3bg3mz
V7IzIrFd2TeWJlyzFWf2VwYQo72zndD7Jq4qOZTvXMq2A9dnCPYYynHH6UnvTwH+onB8k7+ivNzY
cuN85VT5EAYnycJU3ZvXwUm8bqf6OYIkI2s06Cp1sj+m9yeh0/MZhH1Nsp3O90zyfad3eAx0qFYu
ItTXqjgrcvCMTuXj3SafdBIuniBJ42UUZ77a+Ln36jAm0FAjeYmghzblG6HN9ZlOJnBcBhoIKI+8
otVt/8bCTC0cOZvXax+oW2C7yUdeI468l3TwN3Wc+mx+9UB0OXwn/G7Eix3rx25+b9DM3vEYxtQp
ZjnIV3mHfIReQZrbZyZG8lm0Nd7HY8xhgeCqxahj3qFiLFmxCc9GCH0SZGqtvW6CQS9mhZ5FWPJC
Nt+GYJW384SMkx3xDki8lUZmEo7jTjh9lhr11tZ8aHjN3LAOAblLtA0dum/wOM/h19w4/St+l4a9
uIGkgIJ2VEMTzh6hGML05VVDjYSkpTk44ahIQDrKGewYUYqH3YMeCws6DePqz/veBYmISHYEW759
yokJQ/pDA08gcFff/JRAi04uZux8qb3WVz0bXD4T8A6I84ZFYjqyPqLAW7c+GMBHfCaAi9EquF80
CRBIYGRgzgdtQkSaI/c04zn8TQfb1sVgLd29IIhDXyFvF+H5Rsqk+14c+t7A5eMRClcPoGzQ9wKH
TlN44t6g1aNlFnHBGaKd1ko1asB16b/pD76Y3OMJsDsyLrYQANik/mChftzoKtOc0Ks+BsnWKmkP
6CQB8d4m1sB8gIf2G6EXX0a7ABqGrV04Jl7y5HGgsPEBC0S1O0+JEmSsGLpZxO8NTULQyjYD+CR5
7Vmt7bwGxh1Z74CSGlN+k0x00jJMN7oyp2nBu/cALhLJ30F+dHBYiBUBw8Ou2DMkkiXkrEQHJxyQ
yue/pW7tPiUqNrWHopVQ+7yePAnIHPzlrFT5iahiSB5Qoq5U++xA6l+lIRLjQAG9OxfO+UpRwnFo
dIhmPZuODHUomrI0eTeC6pmiWIouw0YPXz+Td2+dwmBRJJK7WFZeiURCuLHtmSDHih6Vrgr9Daon
uIvxBckI7/KeQOd0Ut5LJDfyx7oCytjQTxrBJ6AhyOiTg3uNTM6j113QWss/qZTKPLs7Woh7JJGp
KWD2S4bXZz7LpqFkISrceD4Ddxbafu5M5dQaYpxvfvjwm8xcu4cHCy3cNnUXPBPOeitEj5Y29wkO
FI+zOnT9D4i00wnvmqj2XyvB2ZWfEug/lJI1l8movpg/Q9eykCPQ8TkxVaJEjwwGjANXgZ69CwOf
9N0/dLoSNHW6VvXUpdwiH0BA/KkFUqrxO6s8xGQcneW3G7gXQREHj43cH/LHmhkJDgJJGClm99Nx
kbBHs5vlWdWlmsxgBd8ao5TIO1h8N5lRRszGtkELEt9CK2IyokcxQ3hKzP/Tsovz3d4bCo3sNa9h
ChJOo17bETRbpLcKiQvLISywXmi/83lg7m9W1udXUXLR+TQCQ15bCwdNdTOi/OeCEf0UAa0p7jeW
hBYpE56lmNrBFKUYLwrAxcFmx98yPbgpKz/HCjQkCEudBVZZEHX6/JLeCxLtRBEEKLicrd8Qyikb
9unoe3FGpDBLMGsd7xlSdDGxh+U9xyAy0Ok7B9QA2eQNwHShw8OoMjk5VmHY0OLGgCUioqkn2pZJ
xswfH/S5h3qvo9OnCY3xt58wgKS18kJz/9vR2brWNpP/Y3VQCr8zXzd3KOgCtfEEb9dsOmr1K3I8
hN7QXm0aBtp/AfOMquIT6Gkfrp/Yrg3VqQYPkb5bPxIuBEbMWt9owZfY3FhyOqJtK0k6ViYDrycp
bj1KE+P2ouWW1uegB8rBoQgB16tn5v+caJS5NM71cwoBPVpyeCBFJB4x59zK1pJKtz8KTEYPbBdh
HMPXd2/oz/G9rvsbkVmO09whmOXapFwF4plrWj67jLILY830ntkfwAGeBlHt2oj4k4+tmAqt4kHs
XjUl0gPS/KrXzx3LHibtPo2rW38Khqe53KCnyl/bJx4jCBuwXHoWwsNoPgiVneyrDDes6KI+1sxD
YmDoi6RqFyQ/WbrvRWfpcmQ8rUj3Uv11CWOiyJ/U9al6E5dBIYjuFVK4cf/wzkljxEsfISs9huV6
V7Qk3hcE0xwRJNa3gKYYSakdAGUhlf9i3Z5Z+9W7QoOO8/cAsBZMGmLhlG+8CieepvqyqODFJrdJ
1jM0/EEvLmzfNZHSbbpx/I/gEMUA6dQRHW+Da6PD20cuW7JolmKeXyjGYnOHbT0JmjCJvZMnaUN2
Km2bEnpAEWrnvD+N2Rmgkm6cXpAzGB7diXA/6f6TOymfL2tiAidG3saQk4KN5ltaC9qpt98EdiT+
l1l437eN5vBQoR5vh7PpISV9Po9U8jutRM+xk6aRQAkheEGAG7tukeOZLdl/Uw0BR8O88Zo8Oebm
h9EgB8+jZejSbyxU6aUoh8qEyBljtX1clN/B2Gz83dLTdjpEAfSZczV5zCA2/00OkqIv65Dn1xJm
3dtXI6AZEQB/LMsEddxQF48u+JHFfbT4yGsaKZzjvubQfR7Q4JgRmNMTwZFKx/tn9Ppqot56r0ms
Iq4tMUO2k9PpUaoLXhI08al86WSPoRU/9+Wdsl95CzL9XAj4mMkZSvHuMCxgTsXFLzzE/Nbbcdqn
fA7HfkjFV2f/VyHRq2kHweDF0H6vBiSF39XskthdyfKbxcejSyconCiOJ/5Iyp6bGe+D7t0qgUwU
b+07VfNOt6SBI8ild0vqD3CyIQ214lnKzuNtl406sW3JL/AGtUvU/PYOFV7zGzViti6QKNT5zGHW
fFcVAroA0Ew3LQNyYoUUPhYToYnSAjy3ZoIXQpj/oVEoYaju6TDQKXt6uHRhyW0D+tMJp1X93LJI
VPGTG4FvMKwgkwcq68CiJS26mr0Qd0oPiY5rfd8AAEV0fcrGdfD+RTzQQ3sNFXZTc9FFyGCeoqtw
OkbyjJjgfR0S/qbaSWeTgFjRcCgl9RTR/j5/BzOX5QqrLtizaxZ9LVTz/PrmPigN2a6hCOVURk5x
gBi9owBOD/wXtS16dnq/E5ELFCSO8SVLTMmUqpVrXiplyDyljNQAbvRPIzmfyU40MuEES/d5+i1M
9nFKCLCt0XVIzjK23wqSvJ/3KrHEOCKjSZlCnKoJKD3nWpJwFNUi
`protect end_protected
