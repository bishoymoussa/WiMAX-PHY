-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
n4Swb6q8JQ9KVRJEEH3/djgkAq5usTfBFKRwA820uQbwpW4Tby5GWzbLaHrbq+wQM5vFAJvocQO7
+FCTjRIP9t6v4X++bwibXyKJ8vZxoM75ksVzisUEqI3JDncTYoXGa7q3/39eldKwfAaFW7fvYD34
MKV3fhBAHX9smDtVCBEs5qR9rbW09v62XKail8ynaVcXppsnUJFDPxQEmrJl8TDRAaAZskbIGHAa
FVS9z92T3Q/eu8JaP2f90TZros51XYUxdrKNpMeBsjCbvVU+s34ycUb4HZHPgdergJIbDUrr/Hng
ehzg4Y9dKLcegkiid1gBbyWzFSYBASFJAJmSTA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 114656)
`protect data_block
jIjImvpJvani5IKK/3liiJtyPQ7HhscMXSfpp7x0yfHd3FD/rIVw3+/RQmTRYi7wTruXGie7lxoI
xfztlj4C3wUrUrul9OykrO5DjyfOUitkyBCu0khrKUzCG24IygOWt/HT1RA6Y7VqyNbyFYwgVZLM
Ask+21xFnG7G9E5dB4SElYwhw4Y2Stv4EoXeK/Pu62QB4rEKBUcl7Yt4V/U9ljFVLq630pdC8Z7T
vYq4FyOS1ao3qA1FVw2Igez3bixmwAWp+lPafowXYuG5qU48BNpZBZeWoPPjFivJjOKmerIDsykr
mj/QZggf9Po0y72n3mE31tgQMnJw57o+LcN9qlOCNsbeKbgNTt9WnQAvVqJjsJdS603WP481uwYD
SOSFNvoU3kyeceSwIWCg11O3R7l35q9/S73b/RTHvFOJGaKa2CYeRVgA5r1VPxbRt9EfJx1e8AuK
mgDyWJ/Sk88yR77sJy2uvdxLZLI7/tAzdmj8lvT9DxT/bDbn1sgjJg88/BGmCVHHEt+cBsCvA3vJ
TadKa5F6vEjD1tiS8uKw52fyrEzePjhMMIlSDkCjwex1VpbBEYC+enhqmqbvYfF1Tz3PtxZ3LYe3
fidzktB6nA1g2nFcANd864pTVlQfaK3QWUyxExlhvcd+7/ykKILIMCYFFdJW/OFD49cB4GbTO4a0
LuOVp5P8otOPBDi5XZgWKWBSYqqffODw9Sye4WCEUeD71dLYPB55OllTLde6VBfRinVHWfJswnqp
GLfSHEjCzl1m3NzmfbyPo4AObw02JVVgoW8E2lN4GuxpfgdozBOTYKgnZK8Nd9Eo5N7jNISiDOQ+
2+OH5Wv9b5C9448g8KNigIk8p6POSQLa3AfHWT3b4Y08+TCpTBRTaW/c1Gl9Dl1Q1dnwq68lwdHo
jPzBDCl9qA6jFm7a/SLJwR+fs4gdjjfd0IyLPZYWuojvdYuiX784GmYV1FMZSQUeEqjQOLFt5Nol
OHINcPcrR7vdjo4Ohs6luuPrN6JYLZy1nMSdTOub+WhDjEfMR+lCpbTDikOMMbXkOsnBASpKQ/AM
L2f1EQ3IZAdpOM2gyPCeqXTsSLRFtzmBdenW+7zfzbVJ1mQVVASzpgtFNb5JJ1pITrvpa5fNqSqH
ICQTWa2lwSdBY1aKc59R1EeuATgmSMZk8WlSF8bPebLdbR0Y3QBGajGO22RTkDsFRyX7gYYa+ktw
yILEjyo6WM5Hkzc0NH5vHZc0F82tXL6PD0NXpcuUmTX+qxaEZs0+VTg5Ev4gq6adCgEwqWe1E1fv
TU816SA4LUgx90bpcx/Q5WR4Ri6mcoo+Y7/wWJSO8JOhlJ5ayly612t0vov3kxbSkIBsEJtRWxt/
a4DbtvsLnuysZARp7Xy4/8PIqiEGLfBH2fbh1niyCADNnkKRVg4qGhNuSrx+yhaLCSvtUYiwyRaP
N8iYZvQM5OcQXSzIluYmAXooLCIHqGmV4E4TLz5qkDCmrbuBacl7nI1SMS+oiGnZ9mRAB3R4MfSS
fGI1nRyal4RKJimvY1jqK+2F81W9hFTYpuwZxBFKXWQAjjFTpZ2UpgtGHxoLlnypxEXpqAScMkdB
FD+p2CShiHxBE1nZAIDuEAINbJFqB6qSE7Zw3PQIAuN3UIw89WlpkWePoKK0a6AHmlP3XOek+WKW
sP3W9thgdL9VetuxI3pziSnz8SaiNX3j11G2DtHTyHmxvqfUH2kZIpeh4D884woU57poANww2SK/
SeYiXhgpGS2CqinxbS41GTj+ySAU4WiA9fbBmBPJdVOlFpXB7wC/XfTEL7BLgd25xdcdVDBRx0aS
7KOLJpkAjKh8UGrjP7Ca+fZaw+Tch0clZR37EiGCx4fg03g9wrcg6ndLQM6u5H8NwjAeBaJfGUNI
TzGpaMdEXWxerHkljAdha5bQEr3ypTViiJYRcL52zb1cbR6i5ryPJ4vn8b0D6lzSRtXw4WuGIxhs
5+0wcgY8JHrFbvWeFWI3rH4y+aELAfxbyX0/38e7bL9bUa4T83A2ZCiyy+Hu2SQcXbywX0u+Bf7o
T5juY+baZrhJsPyOf3ghAPgbYt5U+fUIbqlmqiSA0PGE/o20JmF9fK9BOHjAU0uWraT8HsmLzoyw
gbK57zBX1+M1eMvN0Fb2X4+6B1M8Dx/h0W7fpxKaCJzQ+KJI80QZL735fpaOK2jPXvOOmpdMO+YQ
/F4nOCj8fe5awdU++vI9+hfxaH0XHcb+32qSOIB8C51Ddqv7AybqRsP/lzDudIV7cwks90rKCO9G
2Td6Cz43Avd3c1UKV+DpPankp/EbeX3WLl7yA6b45jCpopmNO7ppZtTjEk9XAWr4ZtvexzRaNHmn
b3c/Qnk+WSeqmQvOCkTiXUyXicT0x/aiRm0L72dkdWQN4TMjBrsEaIOPShJKxWjh7/36K9ObebAK
HGzcuRbq6ghdLIgeCOx8npsPMq0YZl+RyYFIhsQFokP5WYASwmRNG6sltexF/8vJ101AAOQwcNSf
x+ogxRiYmY/squu5hrqyAzI4d++jhmsLz+N4DP3l6bqauSvlxNItASbPr96s9nNV6zQijH7PMGFU
+RdsNeSvw9KzaqrcbGI0/ltO1KDkS5oBa4cj+DRoZ2/f04Im4wDlrupRYyPl/N6dQmdgK+ErP+p1
hCNt7ts0Xnkk5AbeTuUhytyWsLjLVqjFwNnmk59xgbn/c1Ykp8lZKV/bCnea5d4epwtWpuz74rnj
FqvHn8sVkOqE9++YXeARl26c11hXWjuJkXor1szK0W/yRAFeI0aiX1P2giBwirOuNGnmhfeCzPN1
91PAwSEK8tStnyVTy/ELakcLaNHfjGlp+nL6xOBt6YgPcHKAaDwVuH1wvUT68EmmNTq1fWZGJPk9
s+5ldgzbXeDbm6KGHl4Pwp4KBDnj6wcScoJGbqMZzVRDvyQ0C5lIsI5jck2ezQoZetawVOGpq0bZ
LfDoYOmtqZo6SDJrWEy3NGCitgiKK7lMpsV23XUIjcqPJ37NeF79d6rQ2+JHwMApNG8E5lrMG52T
5CeaRLEKvQvroyK21Ab+haQb2U7uF05z03KYG2clU34DkGOrVgjzkG7p0C+dwhSF71D9/PjkrMkG
49hP8Kd53+5LkcGk3Nh+aGvkdS1Dnv0m4ffDuZF/JM3JtOgsTXUhEFs9asyeHLVivM0P9RO9U3M+
VbeY4ffRb+YYPMwVwl9IiRoMY0GkNyvyiIhcz5O8s7ep7oZcnDvz8B3xVsdqRqWKq/47r8vukOrN
W5dIVJP7OAhV3P226N7FxZYuDb7p587sz3Xd5EIqJbhb7ssOYyRhPgRJE7xRS5ToyKaOYRhKfryY
q0NP0G4NSLa2m0VhE7u8Yy+8RS2k24BNxrc4gXaiyHHMVXIuV7eXFcc18mE2r5VXyg0eA4JBwqen
SUmwriTVtwQ1h7Yl5bJPHuEEdgZJPDRuZMYkTlz5DlRSFk70MogqXlaE0w46wAfs2/GXP40TQDLh
v21Hq8xgC4Qe4kOAIcidAXXZNsaBZiLH0El5tnVtjTuSZo1P9WJyBNtUHkj/fdHQbd7pB9QAtS34
OWFksaT7tr3XyXaSWp57dn95Ct3K4v9rCrurgyTwAhRqvR3gXVv5hYhN6Rtl2JbTAXzEEaxzH11W
XIP1fC7Lunm7UR/j4TYjlAD8ykU6OdEfYAmVXW5CtwY1z18f0y+YhqCdj1r73iyGLfyM+otPGybR
N5hmIk0W6BXLe4YjeP8o2LgWOpgMnfx0BFyhrVLiL1Rq0y9n5v+qtLxwh3OZfknazxxaNqFVw7Sr
VDiLbnZHENIR1RtZSaYHXieNbwbUvRj/NuVy4uzXA6EpFCPYJ3xpWMf2PkxJpZWTEMhzAPnUNYln
n6PeP5K1EuBLVKad46k4ndGUfVy5b3PNxcl2ZdJJGl82Y0rqBDuM7e/R2NpEM1FheZfZCgmW7Uw1
Mk6VXI4wC/xTGDZg6J0tOaHbD7/40qf4glUVHN8j3JS4Ejl5W+sZr8wt5urzuFuv/kNgUCeo1yqY
ioGwLBqyib6O79meQpUeR7Ys5B9khxrxfCNvbfm0i4Q5T6wWCWOZtrva5+p2ckUoklWqd6k1MP4c
AvrDu4rLTbxEdHOEURkFCH2U8yrnzPmr1dWqHg8OypBhfFH8+Gh9cGzzPGCX3iweuV6h2YC4OBIX
JRtoSU8F6ybavwl6nQNq/EQcvnjl2dEFMraN4pqBGc0Th3tAk5ZhLAPkPIv+t2oi6EjVe+Vn3fDQ
Qj3hB4wcITeA2MXywTDtHbq6zC3iWTPUeKpUvte8XH4WS7bdEf7Hbj7kyvUYfUCkHcC4tZqUOkSv
SH/P0zlxImKadqez3nr3ouHFU312+wCYEn3sfY0lhvEank0Zo6JSfC8+IWGryI7T1f9KkexinJE0
WSwfozxJZJs5MBqMLfO8ctvJ6pPbGAhXqczPkNV6hX5WayjcNA1/LEBsbD8Gtafhc+dHJLgiscV/
4b3Egk2n8m/BF1eicOOkyj3i7ylGk1oIwlT9KkPRObetbsWJOA1eqLQ9mCOwRTE2+oABRJoclXaM
cpTdrb0ha301vZKqmbWxin7/2hv5h17GiCdPQsuYkZa2qx/PeRgL8wCsrRj8o4xo+5b1tbeJrXUs
848ydYTG+9N2Z6FgQIFJtd9npMJQ3YQh2rixPZeZaV9gW0bPZsjEgdfXNH8rN89K7mq5PLZ3Oa5H
a8G6DlhembJt6ScB6QL2pOvdln8Ck2UtY/aTEoLM3LdV7W6gqZDF5hp7vuHYRZ0tsg/nCwGQZeUA
yMwb8yc+K6eqlxI7CIdbsP1CLyM1k193PmgaPlgvMcfkR6RaGVgufJtrxpMDSqdgsAc9k0uABywV
zl6FT6FhxUiTFZDU6iZNaPlS4s9y8YZh5So6zWnAMRq22k2OEPjXbGG9EOIiztGIp90nZT5FomjY
zNz+BiJOheAxvvnnB9ukR79WAOmgzGxRf8QDerpIBSSLdeOLC3nqqiY1coVLMhis5W1+HIuyTTTN
GiIOiTOIg3Zv/mji15mB2dHqp6i3Pjt0mSVpgAaBlBf2h9SWks2QihxHWY8isYKZzLyY85tyTVL4
FB3Eo+g9+canTn3sFga+iTYn28Nf03WqQal6dWpDlR1XEtyvD/G6lJa2XZbrS4SThyMTvSDMpyFq
HJNY27txu7h+PtZ7a+/TucpuzDt9AJdh+EwSpsL+fDGoFBtl6N2gbTzeMb4mt6FCmWJA2l5DAXBV
kHfOF/on1Mr4h0Ls6f6PBH9sGMilHGW3QCIwTWTxTcs1tdnjtJhwiF7pyxLLIiXncaTHtP7VIheH
ZpI659b1FFQVaT5+IlgKovG661Crj/BhCuuS+X5SopBHhWDG6/s+dZUEjypBjWx95SVj2cHzfp7q
89nTZFmkCZ+dw2nTujMJ40ZKFzjKRpreppQZ9sppKz3o94lmsw5IdN+/EIAMKXrrRAfX/znqXb/S
vilExXGi1TR1SxBZmRsF8unOPFHP86nJGQCw+/GvXZxRpoObeE4W+SCmI8SAjLgso0L6FCMiMDpN
dnlf3Fyb37VrUPq1z69bjCCmVJBwUe0hcFFKbcImXAMEroJYN7NzhdXVpTVNDCfMY2KyewQfcrC4
hI/1BMPZooDEZbATtZUJW8wxl96+WIbeKI1gjpSIGLp6bRKJEdXQM5Br0Mg5q6di4qJLTHHN99AG
xawIt1eO7e2kgMFbH5k+6L+RrjFRj5vVqdybr1hhWSAUW2hwh6kFT7npOgwVT+8YDyhGUtitf0kL
Jd/hJUtR9QHAuWykBFrZL62NF1xUgLJ4M2pWlnrTiB/Wu/+ebqglySYtPqB7hXVTUYwjlOK0iwNr
J1dd/LWWe+kG1Acb9nbiEHsquz5CIk7MQObOPlz27jP1Q+qi5m7pGgnzIRdiQxGFDIxRgmJDoLQH
rkgWey1XBh8niJumHpj2hgPRcCCD5UXRHZFDUlF6pK2Zqfpla3drMVDOfERMtuSNJWyAAbt7Y4+R
qYNc6pykyhXkAtmZIPQNaCP04E0i9BbiTThT+VcsGLHZe8JbFGLbkLC0Wk3gZ3ZtBSC5eZ3y1Isp
MR84jyy0ED7hHNl/Q7u8EXpv2CPajUkcIvaUfQd1Qrf90k/Yx9x2q2LfItcAtFOOXI02m5Ki0Lah
hjdpjcMDlao62XlVzIhrm/rJAEZhx+3MRwRflw+7B8sbPw57abKDekr25ZotXUwWzcS4XEhNOGWM
c6MVcvWqU12Xajdvq2f5RFmF/Qp2We0z2Pv3U6guoSUyDO3W554OPP0VQfpQE06hke4zSBS2WaZz
uMM2t4X6DCkjYshaJF+6onmjGM8cqaB9K7Gt7yeWQr9G+a4jbLtIjZ63LbwrO3eIwCeX115l3+aP
iYGHIdcNRjaJ6DrvY8T0Mj9/sbl1PfmzKBL3wliE8zTLXfoGVQJFNQrg2uLB+qPfzO/5UqqvqEpd
3ZiETCTcUMWtu7dXb9JRxEFTZm8o6K5XiCwZp6mkTUJmLDYkSOhts6tZXA+qpY1/q3HhTb8m6N/Z
fjqU4K5m6r4cltLlJXp6/3au5KpKozshJdYxkVuR716GvI0pz3GtWU3bIhj6EERtuIvHLGaufyum
aPgbxOIbZ3O9EYqLCBpSh35Uwy8sWvge7nqLhh07VrihZoaALqDJysrDcVF1BkcE3cKnT4z+RT2u
XnwhpoSckysqsjd1I1P0h1tcjwiHKdMN7kBw4L2pm+5nbyml4SFrs9LBVJTr7Lw55sBjqjFV/zOG
PM8NtN6ENh17mRqZYsJEtLvqfixNDjmjewDcdIYUtaf7HQx2B3G/nmQ95v0qAUwRufPGuRef0tF8
FpyhM0Zsg8IN/B1bljU04ENudFWTXBvNth0SocwBpUQTcCvLH1GO/j0tDrPMaBmlQDyrp4PkF16U
OiDlFL5FDRvCQTy2MzksbeD1/GbSQeFcL3Co7qz9dS6BB4sqvRwbLd5iFpk+L/HltGXLvj93WwUt
1CMWtuH/v1aZYxvcx/SM8V3dydT/Hr8I8XFB0HiAu2lBxd/BqLGcxwar0tEwMxZrnCDovcTqEnY8
NS9HJi7UB6mAVRh+Q+MGOEVsteLgJx6iI6+DOFO0jQydg2nsXgnD267OQAaYIsusAmJtSXl4sOpP
++il5cets9zKDmS2iGk3CihXNR8jBtp8hyrkp0krVUyoAcR9rrdr0jGHLCA/gUUSz2PM/eeS8BTV
AEtGjZ75uxg47og3gBzYw7yIBmKX5Jz5Xa5hTtPstapH3tlthqY436g58ymO1S9jeIagpPULrbyK
BtYKzCn3srIxlbBx4CWaAfYECBJ9QXZw+f80A3DHwMgVMwhapsfB0hdsMEd1c1Fj8WIeKN0eQ9NX
vgj79OiU+A3oRorD9XuXmPx3UBuIxaaotke3h2+uoyIG7eiX4gvQl6pOcCmb9sSisvMGFq3eOpzb
UW8UgjiDA3EBLsk9PWqx4zyxupgkAdI3y7lkgzLIXy3fFzI4Gk9rU2i5FgVYX3wseAY6AsDkcpv2
nwxl3kHuDspathIL+J35pVdTKTkCfwKYSVGoprPOXp/rn3cB2p/frKqrOX+/MePahpXUcVVjhcP6
E8GQo+LBtBjkcSBtvkoGdB4fowN3aKxQit8lNOZgB7+cA7NmM/VnOIV6ajTtqBsMRQDJVoxxijkB
gpqqwmteL/6DvN2VsZVzNHI8kJY0IywKNnn07mWYf8rBHqJ0hmesSeQzbTcDW9PtNS3tpLH5LUhs
o6n5FEKRDqJzgNsaqZZlOv5tdrbvbVfUllqPLdAoc0axXZUiiAgXd3Bvov0b+qafvgUUkhLkwfFg
6PXqpI3okm8zmkAEuYs3itaZzaXyX4FmNxGT3BCUzUAV41nShHFYWHFFn4DhJmm08Tmp0YQtUACd
/JOR9BHHHHV1HrcDmb7EwpKfBLA3o1PZB849L6pHVhm3Zgm+x+s3nL/V0tRS1IxrHJQrLVIPKLON
wt+5TN88fMDDDJscjzfPoRx1XN17ELYx1v2n3f6+leFkUkay81qwwJvCgxS2psHc5cujFJMqmFSj
rCHezmJ8qfEV3mHk1rUhcqf9QGljtCtTU6utphogglx0fMRYEqW9l4sqqbow/Z2eTF6pYLrk8IEM
d8x/dOGnl9syLkvtsOl8aq/LBqm6c6xXFPjtEuEa1RtlOKhTlQoZ37OKs0/E3XI/523c+naLQN6G
vhopKEDAgK75qQiNGdcoBwOwrqnWC3PnPztRKs3bqxlmHRtg5chLt/ZAx4aid75tAgUj5PQC+H71
xliVH3H9bARirV5DoMKx0ZrTwa7gQM7RhKkT03ukNBsiPCoLB8YFv3GWFkP9rcmyfqx8fW3vEsl7
o8FZtIOfE8KD0Xp+w0woKVa7PyM7Z4ggIdw7IUwhNtqJ6U4bkd5gE23cDH7agwDxXR7sruL9dIdB
qozkb2MWnLAFbGgZxAReqLAcjIdtWo3qhsu7X4YPYu4h+zs5I4ANGqgcj6JdkZiVVAb5TWxgp6nt
J9k8x7xEJSm3z21bXz0oTeAE4KmwulsvRH31ZMqJ92BJJFBRQXB2R5Dk7scd/9/GuP7hqU93dDoh
YwIWF2p/QEgPSW2QAOg6CE58NVNJIzzLCzRP8E4j9wn4AdE6E6TrdR+2JIchhSU8M/dMb4u9gg2F
jSPpoii0mtdTgDLqUA0sYeg4dhPPJl5Lsz+cWsMfHxIQ/YCbU7hosnotQ4xcay2WHM9jJWK68VjL
u8FZVKywzOSdTikSxwwlrhq/lOf/IvzeFgRa+monFtGkkd0jsX07TzwqNdMsWif8EK8iMDxmFX23
yIyhfTJDigo4s6nEanaKCVuTumgx+nv558SzcGPdFHW8I7DG7JPQmid+Mq0CfWcP3IWa0z45xLQq
972uwCcVDSAvJqZFewlj7c7wT61CLIZWCdJ1htjkWRY/j+d8+YSXhXVyVjS/Rw2RbIfTLvFX5GdH
yj4vafWGG30SWDmyp0o5Zi5zKcYDWG0WQ0IkhyJrpe9IoLGc40W9tibQtN0UwhliicyojiqcZkVH
+djdZ0ZqA8cpE+PHqSoiFESFDeWSvyYpDUH7/eNTO0OX/dO78ibmpC0m/7WjTuogPMAjgVznt3Eu
lq7It2Jer5m6Odtli9Tvi6uBAOc1IxLZ814Wycdc5vaDZjIiadLrN0Wv8U0xhsdpAd9CR8U8PyOb
G4jnn57Llj1oD2eZV+cz46BbzSMWxCev22i9Rf9XTIpKlhcyGHT+Nfes3+EL1L0NAlFgKBmvGvlV
7mBg5oGAfVmISmSd692CVayt0c7EITIgab9IwlpRZW3kHIU4GvRT/s+bpZiNDtXgEtQFpjfrFP9w
wmHRrfD4S5zwQ3c9M94FXK7plzppAVth23DG/0I6Dp4Gkei9du24NhIXNQTKQU49MW6Q4m54e+v1
NBdW3RZyhgO8W3/C4Pqeh4iWF4Xyt7ScPiJFTafupBXeS+O9aOb2TG8WW2RFE/iSu5cdg80Z8VEy
T4nhccWlDtwehBj8lmAT7qmM26pFGNzJaq+0llwQrcIXfOPGpW8iZdMB/PA2ETMydugg41sDqo2I
wzx7r20hafEIPi81ysocmYqlwfiHi/y0ijIbfkGWjxFC64d8+szKDBssSkYMgcIDjYEXB6cKivJl
+iV96m0OZWsvi/p/q7JJuiy0jsj8EKgufkK5U5BkXnlZ2e2dgWYuxv9oWAbiwXLnkome2RzxPvz1
Pw1IVXomgZnSc7qMpBXPb6YiWm9UzicvhNVb6+zCmE24LBWTONHZkYETCjQ9NT+QebLaqm24bsqK
g6zlEqvWwgnJtqEuD6iqhzQ7XE9Z/C3W8iOOfzrfvaFeAwVFLslAogKRQpw51lqgdEBxnRZ19oXR
aQGWAxpQ4Fnd93Hmv7rLOjgGWjjASxgbpCj7SIMVv0fjsDzq/N8LRTyu2/VRELlc+MpFJHB34YVg
n8N/lUGrDmnQbeHeKexq5Fo0dRLl1hGEgL/VlGT/L2KSvLSz+PE0a02f9RflmOOOcYw35z/1wGYd
jochBSL3XyC62bIowPF0zFhFO5gZe3s3hSEDOa79Odnqna13HJjm5zmpIenodOOdYB3j1TZty639
+sA3+zru9+V0TocDsQqPlPswEUjKoi3Ld1T25bYMvBdDnXVtWSoj79IhArK0pxJEvTLeKmgdaWRA
jC5EZXitzYopZBQjo8zcHiePEbDLQJDNd7I32NCrej/5AK9H0lTOd1eaNOrO2s0z85oe77S4h+RZ
KWsir4ZxW/FZ2GkCfGWl1ux1PU9MuuwFwyDowMS3OyvN0tnOJuTS55nTICDMGVqkCjJqyiSIe7hT
KwVu0eStmfpT1V7aXCkSbZnnSB8Ozok41XAHjnZQSBcRQiVW6cS8MnTFtYz3iiFUkZEFwG9Bh1Rj
8SyiLkOQ/N0Cn6hjEJLp63wI7Q3SoUfdGK2YPQp+kwnnf/OVyLVEOQv3WbyUZUuepcpsXMaSX2ze
3tkKgv63hTOsKOK2fhIGb4uxYPoEhyAHEFPbKnssQetbg+T+B1LnGiEH4OZQx5ZDZ9dPkyFu6qJP
jKkkUKLvnYL8+P5yCr+Kbp74HqNCbO6w5S8LaeL92Bts7ke1cWPSwWix/pPfwZCYjw/POInDJykk
KteOuieXfC21tK93l73Y/ssdEkONsAgLb9fGCI4oDhjmXr/hFRZoxg5aOtZPq5Nb4eg2xbunZEuP
b11J8lR30dzlyxD9aUtm5ptXMeQqHWrMtQEeeQZi9Xwdy94sDJ9rJeEbIgcgEHbDY4ta1Gt0n+Wf
LOpfRcDfsBE5mhBRCKNzzz/DenlV53FB5VUNgUSad8P6RKYZ9Dt+wqGqZHqZZyfND2fuCiyqdTeF
57ZrNcKszRhxMP/xxPJVBMSblQcNv8OblWnuCrYuvx60hYHTbHFyo0gbq9BF3k/oOaaoF/j2naAz
+SIMzVcHIpyoSLHcKP9X+iLeXLjxsiJCYMQd/zs11D7uO8Z0z7DCu/YHoA9eO9vOzYI3o49SLTIs
9oRcrApr7FP+DSoAq5Hl8QPM3X7PcV1KbIGRU0Q+CXJopMfpGlrwipYVCiKZY4qfpSM7PtY3m2FR
PTLZEz8NfW8pLxmhqvyX00w6iUCvFqxyDdxAcQwgZ1Cd79hnI2Js4OFo0NoniQy5YgGPUH/IC0pk
0s22NhwCuBCv15dbL92+gXsQGLJYCB0LaFPHgWWBHkcxe3WhvGHeAJ3RavCEGn6Ue9OjU2jtmDSU
EAqUGeVAg2AY3twW3H7F4YaZw+D3N2gu5Duo7cOkyYnhY130W3+kJ2Lf7Nal247CI9lK4wp/iVim
jVCiq8NFiP59VkQ4+XHMRfFfJ/MBi4RXmX3C/8kfeTcLJjddbFH537/TEch0OD51eKoc0dlC9/9D
7KCO99QkaA2bDLicJyVrS7ueAUxJwU1x7fwSP6E6oDbdL3WwUbaO5cACPr74eWAIWyS2id4YTToy
r+slXyPiewW3ihEmMMtO2vkttl9GiQW5wBaswVOlZRgqAcuF+Er9YdZGzTS2KMCJprP0kqeNLMvj
1IwkjDoVnhpLjg+sswHcGY9dP6BiO98A5KJVXt+k1TZXYNaeQJ1otDqeYcZJC2lEeV5bZRW55fw7
aqRFR4gsqnQgq3qoQGkO4NBkdtH6fMjglKyfkmj8HptuYyyfnE07Q3DswjDk0zPuycnVxNfQQQNP
Zz+3TuFVbDiHF1bpywWuzdMQDUzxglFMjukila0fyQS5axh2Se0y+ur292UyyQT5xKKYbNNdK+tS
v3ILXTk3XDq6efrQDqdGLUwns7txb+fRHU+WiCqhKjk4cUjvItvOaeODrmGOu/HeutRKeGvzxd/Q
R+1im1Zwa1P12FqtawmVCwNPJDT64L2bpBRjZ+tZC+8OhqbD5TPPVsfdiryT1Izv00BT8/0e4s9S
RAbr0klJjHXFtP/DTx442A5Z4G5kPlmf4/LiJbVbZ2oAe1BBoX5t9LU8prS+c1D7JnFxhG8TKaTw
d797vI+cxFPPinHSxaG/AhcnqSVte22/9LkMXQnaYXC4L/REHMI1f8QdgcQbZJBfy3/QeRnKeUUg
HLZeVOIqdw3j3jlWTxW4w6SV1if01MK1r/grow9gfeKGuPH7LLrOxnFFVaOeYcLI29GuiZYtz3PW
DqQSpYQFBYSNIzuRlPXIQJeHoDgHAPt1Jx4l930rQ0/mD8sOICvqfF0IEhoY578EaxmAfxL3y/Qo
0CuPGbx9I2Yo7Iun6uhxDRAjm5to1dFdwMWnMaRrYhiKuHHECI9qzeCCmMY01f++RfrYXFA03ZRw
1WsZNCfftFHcJzcsSbTEKIinx9mz2JrDh+eU7lYcaJz2mauQXYDEfN1gdO6ZUmWiHIz/3mHuuJtB
eDYdWLUFXc/eJ/zbMybCsPOBZHaL1j7GdmLkY/bdQWjZeXsEaisl0eX/bXTQbsf65eKfHXkRzP3K
WDeuSnfUSZOVc//UB1N2TY+4sFRLh60FY42e4uukhnI58n/+CU9TEduHHqz0w/uLDJdUPXhozLv6
klmFFuJOiZJn1H73/Jnyc5yghlJuG8MQQv/pLIPIwBCTvDR9aXmXpLCGw1dwTfEUJwpCBd/b0O88
4lpi6CXtg8dRl6i6q5kVsXK4b3VDiKopLhd4IJIPvdOqj0bYN6ZiAgsFC0Dj9BzAPem2SqW8Y08I
rExI31rVJy5XemneXHelbUS0fRi7Ut2OVOKpBE3Vda8bIpclyHT2eLkSAg3MEv6eBmtzr+ZMX5MY
KEhFfbR2mb0dmCzjXvLpDrpZeUSc7gplEurLozEPXeLpOFJb3mZ1JrD60Wdz/Su/yI4/ACU7V9v4
uzD1VdwsiRuKy3c0z0iWSdZT2EaQp8sE+HibqB2epO7dA1cVnDAupn6fbwlz8OhRiGkN7mBFpAET
ZAQaEFIhIFRtvlHzXYhlq4pQag8dJE5lZLtY2CUBK9W26AvCFtPpQe/jSGtyJ+8Jokh6gGFglxxG
hWreX5JFQTTpPqOcqEH+Ths7FjSWgVvZzQSR1iaZGCuD3P3x5jYZtjgWNM+tMudwH0IRsGXT9qe4
9UW2P14AwCexSY86h/4oNg5OA/NNQu0a0vdiOwOs2JyYqj80hhvoS4FpNXHZgxvSI6hp6FpUqICL
KbbloeHdHYB4fkRNmqCIyS50mAFMAAfdITaVGLChxlzJPMddq2BW6YgXmB4DHohTRrJYMa0wDSLO
ob7dZF2MWaAh2DwRfEnkuw5VatWWPYvhBDRkBlAvxe8yVk31f9gWnLEKgcjYkgKHg+Ph6fYTnSCW
T+zLR81Yxpk1kKnwpsKGkTY+FP4yAHtGqHxOM8VKh6IJJnTIGWn1Sp649p3ZzLMhKs/aSuxnnB6+
3BEYFVxsMYFondNw/LIY8tnnmysVrPl8jktWfPiqNHqgYlmjTqpa7kYty1PWI8g+ydAJ5I5Moctm
PuEuN3D4++L73z/Y1XvEJhe529DvIujMxvwhGokXfV7oGxH2KdgQ8/9IsalCnh4f4WvG7z63DYbs
dKKy5mX8fpdQpOj1W+ARATo7xEFtlZn6E36STBYXGqtXnWTJnXV3T/r7VdkAsEweUm138gEpgSbj
axMw0+bMbo/es3wVa2VV8ioLm/AMkrMH7hVE7zUn66fbgCme4axITVXn7emPRcBC7LBsPLW6ps7Y
zF3kQFoYefCjOCL0OC24iq7R3kZ4RXzEnJ3PpFX5dcPqUc5z4kjbTq7FuLg79quNHYLtFUtHkWGH
O62kZCH0H2JmdO2XVHdQB7nHeO1pb+KI2dTaqPIV1U7tn12OoDR2iPfvt/XCDDa9dhTKg10l2Z5g
cKOqtu+Xv/dr+eqFr1Q2uqVig1vIM3iChclcGmg0KXJzdrk5XO4bDVBTGNs5o8g2sWoUQsEaSkSv
ldTyDc16lbBb0AVmwTHXwoE5XK5YVvQpmYNdCH12/lwEgXcxWmgL/9rq4cExG5W0rfpzD86/Bkeq
vy0ewmCqAHVlIK0dBrDEelfKr1Y8JFTTW5zcziCHC1Drs4Gr4rO3Kz6yhxOOEbIW9Um5yt3ci7I2
xpDb8TNJeGvIHbdaWX7Mxr8ezZ2H+f0FXkwStB9IQ1RTSdB7RBXc25dix5lvPFVFOYR1hRv/1Uq9
C+etLWdm6gcssy0yKHP+nNpG8k6iQAJSRCgu+0N+DGQlxW+Bgi9UCv7ePXIaJ6Y+YomsdvkNZ9x4
RHAFfjgKuqaFFdXpWdhbGuJ7DJK1cHFCsK2AIBTKU/YlTjyNp79vSYnPhojH8LfPgOg1tOvkFlON
pyFeeAaEyWE6WRER5t2RHx7GzU+SOwEVHPj5Xtd5W0SWZ82iALeIztZapIQcBQS4x8lPYcn9e2xC
JOOj0jO6zEx/hTha5T30O1LX60RygLgLFFI3GknGhRtDzkbJS7eedjzytTCnse304B1Js8+Hy9DG
sxgzAd5Al3ONWyyDcXh8qeBoVYjIjGUAPhS2tllRNCk8y0tHO4/xP9HsLDnF1PqJWGny+o5l5+Qt
JTFQy5mnzwsdNY7S52Wt9m5jCfOEPa2+HPo8BFsQHGFUctU38NMv9EFW82UdnsF22yqr+CTVSk49
afqvg85Slz/MFbzqdHLU/pMujd1qr4LbXTbw3OXD2b9k7ZtU7yaiuGyvbF3pH/WJr5v5bniSTz2Y
I9IHK8lgzbHlmHkpqHRSGXKKaMmmHrpy4FQmwhx2XJMyl0KO1xL/Ryu3huszpqf+p0KTqPyyq8AX
QCuI2f57jiJufnzYRGaPj2vqxljKMf+H76S528ns5gRwS2fqj1uT/lZ6nWtksbnrC/t8SfH8U/wJ
Am30iTWp62Gu4aTdAYegkoKFMxAikdrFg4GsFQHHblnOfizu4YOHY6+aI4WUWnsIDS3wZjY+BO4p
OF6/5QvrR33RPF1lHgQ8jMvLpgyAzJxtToAo0Hd4favO6moX78Nyz787tl2YT8oOO1DKj22Ym6tQ
K8TqcgHbevP5CA0hpuwN9f8O4ArAb18ElhKbtSs3Je2SwnsTiUdz91TdEKQ6xR6n3R8PLOL2cqjO
fClSCM1sOabSfhxTfxl8b3Wx4zHfnbNq08W4/kAEjCRrUqlfSa2pkvhkdFfM6PRAO6fzHU+edMDD
aLL4StPGDJsbJ/72Zq2z9wMYQv2y1i6XzK1S0cipNEK70mBbvzrjKqYqjn4QXhlkLhv/BKY99L5M
Tx4AxRXP60VoKlv5ErFnJLdQsumxH1kU1/Tb/vXZz6D4P5bpOBQqFnV3stgNfVwRRztP6nZh29y9
7QVAkcwgzgNxYuwJLtlGaXny5oIII7EzpbockuJNhIubtWOfYyWYeFWMAoVhMhdoQsWOnHkn13kA
ELklq6OfAOQKO6UaSGAW3eiFScVZzlsqPtBDQ+p8GCAstZ1LtqN0JVsDfgkff7xbK31mHxg/C8Yx
LKikfJcfZWZjJvQ9EfebvLUQfkmxMMKrCIAR/z4owmasa2MS5PLtrzORkJCrfX4yHuN+oPI8Aof+
NI/mk1i2Zok79jWK2Fuqbk94+YFA6EckK+rtOI1lmSgpOzXZMKqZhw0zKP0WAM3pWEqT+4A/+afc
Pp9REdpxxYfckTr3P1QlP62UNSRrkRvMlOzjUK4yOU3Jd+4f1naugi9gNEo6H77JjxPL6OKonp3k
+cEzZbEWqqlK8e5V67fNQFpvM9zplW6Uw7suSG0C10hAQ/Yq7xAb41yGDy/Vf1MNgXCJpcQabNcK
6KKr4UpUjpzFoIY2BSUwarqg8cYdkdfLYOyEuhm7q2j6bBssAnSOLUKOJW9hWpL8xLQDlh7f1LMI
ZtFlupBDgwOCraQrSnT5gzjihyTPjsEgHkZA2JgjrxJkdUgmPkjwwXa3cIht3W48xvEeFuVOR0MJ
nITupXPv9N09M49XT8Ztl7PLUlRpK7gjv1HS5kKRvNGPvjp/QW/QAFeceubqrur9BVX98mbMJp7w
VlKGq8ClPMw3yasbzSMMo9SErxxS1Uggq+Fl1yeWKCPLKl56QlDftUO79nEsKSP3EsY2nQE9qx/h
FdNMofT+0pOz1LU/fKpIoDckXAwg9IDvgRCBMJawue3bupnjfVkJKdUjEr+pQ19O82g57px16O2R
ewLsorVWedz6W+9g/5mlTw66mDjqMdn+RYcpQiPWtiluWLmcSwngeMT0jSXqyrZKQ+JIAUPDABjb
po80wo9U+7fNOhliDksBMxiKIaMpDsYwtiG61rFmeWsyzsdgh50ChzS+RnVk/IuuTwLV1gDCeR50
3PIHcPkM6RpXf1pQRZ07mi80CkCOMPg47CWGaAEsf3FZLWyi7g7GYQmz8Fsy8hxi86pYbiBOJWPr
jnySNidJ97Isghb9d0kOt0Ea6fZN+t97xs9+VQk3sXW768SuEu/jY8DqoTCQJnBXgkeq7Kz45fvc
LJqE5xzpHFow4Swr3bn7cH5ft2efn+0bhhaKPa0ltCygt9I/oM9lkdr29Y+LHWTLiNYpREOxnW9C
1WHZcbVBIo9AO+Ed/iLUY7kqxON+u/r+1ryhW4SR9EmBOcd9tJS67d+8ja/GUvkdjh2HF5ZEpdOA
WOUJqtjmiHgpq0QscdLoem1cZn0mnZOQudeVFM2ud9RGyVnmCsLWvyTcFYZBtrWzH94ybH3z0sNf
NILlTw9UFWxdGcvLNcMz+QgUjCCkX7ZKpFoS3zvs1XISKo8l0sHg7pH2f/Y35He2RnQ2R87nqjJu
wbx7pTX4+G0BcT1tNCZfGKh4xaGuJFNhMzHbd6VGNxHNiceUFEYLc1cU9tje2fazgbwgo6p+svEE
bN1KTK+/G2LOg/8goxjmoPdjX4Xpd8Tr6W/z0tcDF9zhCJ4Y5wv+/NTN4CXIhf6ds7FH5YoPc93K
B8BxpvTBdTo5c2NqSg/VGsrlyUOwCjZlqnhIArYgMYb+tatenHaxw2KbX5Z4luby0vesk7xEuiNb
4/jfkTAfjv484PTjlGVO5xvK7+7XRa1wCo/3VzQNGPFHFOYgH1rUQUW40lZAJVJal1gp4lLnbh8h
b8Tt3vEaxYkbGhBD5xejwLTBJnZIPSbnKV9V4bVieih/g2bIbWdjg9NJ/L2T/B+KqOPi0e7Zt2Ev
UQInZxHGLBrPlteqONNBGJqgd4JGYKFqJZfzJZKJ08yUbEdWB1af4g6MjYZFypImi2YmS6bjbAtv
yFcJKA+VJIL59kP6CsJEdndL3IEhueofMTElGMdO0r+Nv3P0a2fFsAoWJiL8agCFlymK4NHC/9GY
/RGIdw7R0S8nFkvQ60yYYqtIPX/PwcMxy1cISSgEdsRkUXL7xtLehca8x6V1gUUurwn2tt7x67Mg
qignxuVUk6rjAh5G3d1tNLwJJdR2aVFgwNfigbq6+lZI6Re7P9zJRXX06Qj63IdKad10AngO9Z/f
XalcnA+wM1ZQ54HB7DQ+8p6Ki2St4e8devhNlzRSXo2SjTazPozsykfmHIKJ0WTeRlcEhV/Jlenr
ZtM+3LF4icZPP5drhlK8mMURbcKTibV6ipXL35Wlq0sY2MXxBO5zM4YAs/oO+2HtsPwCrNHO3TEb
W+jVhD//NWOLot0O3WGFx/wyRM65207NMuzV475sJDxfIRdu7/eSwOhOi/XRZBx41q1VesgbBGce
pK1uht4UBAXu69JqBLWbcTb9+b7r/poUL172DSL33AXNSPEKHBWEGGbpEma9XZgBUWsVOE3B5zZA
ZNyHUSKtUWhlEKo/60zR43XGv9vcEorxJVtH6vSRoG5wU4IR9mG5wjE0b9T4hQIT8M/66vfoZdQk
QYwmEPk3qae3WVhg0HnmIxfcLwXzEC0VIYGtZZ5xCYXDXn0Lk9KdTaa8l73rDe9PIvixC6ZuLW3z
DxfMYhKWvTnVEzZWx2UfZbPFSxdIDmQsfmGkSXkWa6gKwBJcxvWLpF5XH4sskECtbnHBFYU1syKv
UCL8U0/ixVRqfdYQ3DbHwMkOgBld21powPsGge+u5lMKYJ7knmCk0uEOsnSFLzLlMoqOs4wbg00Q
YTsBEVFDwGe6O8d30KFJ/N/JfGxoI9r0JLoLDLj0/CxCcvkSOI1DCvU5B1a7HQYE/jhag7jcoH8Z
xkz5Mhh76n4wpbt+ZdMHqEoYK82VW0cJTtNRZcaYp9Uk6KGaXaarZ05neNhUqvMLXfQsei9EFBuL
kqJjpE3j0fE7VEePWTVg+R/vZ2cKC6vk1NxwSLn53EoZu7aGvCPZKqFvqEnsJY26VoympqYii9tr
Kn5E7ryZWuFyrHVTSOgkAORnaXfs4vEvJCMdTIWdsCxbSbxNngQYOm+J1TY3lvTNmjV8DvIcryqZ
nxJG0wqSu8s3HvwQjxCJa17QObNaUb9W/zWSoGAGx9SxDEqzyk6P+yWchoZ9gRMiit/B4yD9EjXn
fdeX19r5AnGxmHlg7HD40Dw0vdf5NwKlZD97un8myK/+IBMvUpzwK4zFOcwlFBsmn6QLJAx+fWH8
Uw5PVYu/FbudFz7BoCHz214Rf7dqUw2IzpwLW//wS5471Yfx8da5yMUrRTgAFW4fMnrPryico85N
rkDUuqVodLfGI+L886WeElNz1J1lEab6Vr7oaorD2Fj+/KNINq/qG6kqfDKQKPWnAzT/cR2zMXCt
MaqVFTdwAsExnCEA0gPTrmUtlynLAAvzHazbq6Qla7vz2Wb52I3I3F1Ojn39NVHpJXlxuCLslUSc
nvmyzFiM5oD7jC/YJRZaDjFmCyDR5zCLpOy4qpsA4xVLF4rhcxplazEc4TQdbKgOr9SegOp5FoJV
UhhHjxsiiwBYfWj7rVz0ajWuax7awpNCNK2g1+9IraXoPBHdcTbytiekywHpxTefCY97jGg/mQek
RRkTnloLDuU3Oi8opXho7BSnPXqU6X4HDXIeTQ8D/c3B2cTewuRZfIPy3EOvLum1TpaBeuRRtFsY
6PN/jd89eueQ7n6q4w8o+W+jJdc2GLVCYmdWKw9sF5bkjJ2GtL2wtfvIU+IoPlD1OBvwhmlScseP
gkqPBrFBH6ymyiMDzHkXie7bFzApgs0CKX5tOt9Ce6Ez/l1bA135W6lEwsv4EUKQZMFX62G2ZOY0
0tJUzSh/gcuIUv/VTO6nwe+TzGSfa2M8m6CECjr6s6qJgWwClW9YChUlHTg1aOt5CoV7+GEzE3MX
Jr/GOeP3CRQKzGFOqS+VtkRPTbxHP/yVF4eHs/p6TmXyVaxyz80cl8XeARXOcBj6z/hvA/Wkw1qT
hw8kx9Nh5bw8DYtgiouYTbvDzL2Dne1NTs7ViQtLYDiFXgHm6d57bvtNhlV+IzqUaObADXkY+5X6
kL/F8iFnSQuJkTUnGDllWGnN7L6Uq/0e2/tsxRm1LBvyO4a32onBNPVAKqRRzG9Gwgv/bgyjI9gF
Pfc6T4o7H+HzkSg8xi+iFHpkKcTjCRrBQCZr2UMk13we5IPG/Ig8pqntnOgza7TLKqqvRKRhx0E+
SW0x/aaElQnniVEuY7TYLffceUCekyEUMMQ7dZlXTIcS+OR/KwNe0yflI5/64Yxcr2NEGpvPJhjY
ERygVgENb0OQqLs5XEFgvggGI/m2TulLrIKVZ6xlJOVc0cyX9LIxgHiiDZ0KGuGOvgjvfxtiNUC9
HsZj5yWejCAJljtNaY2zuVJ/fPQ2FGsSgS9aaY2aN47laTKZ3Jra5tHI9Bxueg5hHt6P4FtkYizj
sQTE7I9Sa2AX/weCF8queoVN1ViVBJl6sHFppd3dhRMF1/1W2YsSWcRGPaYxuefzXJVLPRbkugVw
BtFqqFJqt1hX7gQKOCS+xmBb1BMFTN+gbal7FwBKumNqyZB3zppvUSuu5WWwiLnX38dxU1yqemBS
bLD3e0x8hW2OxzS8PGSl4qLajj5uCtU4xuer1ohNQjCawzel2eoADVimvWQ93Z8+RAlojp9B/oLP
lb3YoS4DVI0Tq7r+K40V386R6yomM3Zpkz9496pYrKol/xToAuclv0nEcagJ1HZtIQIKoRN86mZq
+HVr8xuoDycIlxJVZFUkTFXwObPgA0zJdj2/EvqSMkHUZp6UzXMxD6tODsV2q1jxjleOL6+byf8b
mu/h/2RZlil5gXsvBP7JSzQC78yHkdvwGtLrzmgywcC8VvFpZKWAQeOHXgbAGErBn5zfL7JpkCVZ
CF2AvocHs6jz8q1qKgGkDiLvj11av9pprFyg83UHC2ojK7EwI8LN0BxkV8cYXQJT6uRAEoK01mMd
NyNI4aDD5kx/whPc66e1nGI0DihgDwpUiS3gn5oSlYouQyYgEezsK4oxG62IBdAu/BT0J45SRBGa
QAu5G9fdts0m31ZrPP+ZLxabSFrUeMRdtPCGRxarQHoAUjwExyFTZT0ked/BiuHx9E/7Gt+5FfLU
5kFHPzJte3+Cvif4v6XTg+IS81GxnT9cduHQ5eRy6qapXFFB8KHq1lmUyUjCJU/VXIO+VpPJuFly
D8Cr+VCICdW19JM3Cx6+FCM/dvFJ2eBnvWFN5EuyOuDhUdxI44qrxqE8yY19TwIPLdn6h3YZRQtr
Tl+h1XdloCvIqhvUPIQgEuefG38do5QxLDFASYIFt2fGW7IcyXIi51Uf0aP+NdF99VHh1zaWP5We
THiwGYih0KKxMdoXBS8olwNvneRL+MFGDXHlY/OYnH/O72u10frzgJINTrEe8Pb5KR40Jh3Z734P
bu4y8reTZjeXwdWTrh/wntBPVdGX8f4wDr3w4x10nKQwyUTPDEkUGKZlc414YOVGskEskXwOBzA/
tF6jmGAs/vaetyYnM63FCPMbR/fA2vB11idPH7V2jMwnxRfPKrnNVpZMbpf/Z+u2j2RhN4WeJcPb
dwQOhRzdjQP2dgMiIQbBQi+XYdoV8tK2EGc6w8kQ4RfIsdJ2WZ3owiL4cvHGKO8/tVj0Pf+yxZV0
vr5MWF2DC0WSjx7xbukkhCTUyNvqyoH505Mnq1icnf99I4J9n+q1GFaqRTQ/+sKohmrbhGb+sDHP
Tc6z8w26WfHt0aOjbPNW1qDH0LDmZ88qoTjYQBFKogJ4HfwmsgNStAKbERHoz0bQswkC7tx7tBHq
8kilmh+ZKuIaRhUDcMEphfJUN+S+o3xuYWTMBnWZ5Dfxx1K5DSQ8ovLcCuzfPqEYfP76MQFNglgS
QeRaKKb/SnXHL6/wpdetSwacxwTSZ+ggTqKGUR97eGY2BzLiggfNdGj5rxARD3KOOdJ3NlryOQ7P
SZu4gYSYZGEzIefVwSqM/oqilbyWlQhbi+RuHomZwjqBCDb2OJgiLH6xBn8StfasybJRJI5NKTMm
VpMsy+9XKg1/2+osstMACUToo+x/zR+legmdahBRcNc9qfcdT62iuwfAeJw/tT0VMx5SyOwEo/U6
uSPrMDsTEARQ6M6KwHeWqnqNAgM86v9vorSltoLGvsY6GBPY+EFfMKJDm6vmx/6t2yn4beRWhxoQ
6BYacIqDYj7/ORRFZdH5GZgN69wZ1iHsHNTe9AfsfUU6NnN8rtcPEORibAa8nurLeFQc0K/BENv3
dbvwYDQFkoijC29Zf8Mgu//TPGlYiCqjeK8mZK/pU+zNjy+ydkiIpn2iKNVkrWY0aabO6t4FZQlW
STbqy0bRCTpLZwklGoncFgBufjV26HpBdqnGG54t487WhjwjlD0ceSh3N/oyp0fqhD692+ZvSZzm
Hww+qzYMwxrlbnIbdnvvL2ykzp+Cc76HrzOhHymO8+a5P0dFc0z6TSik9GfAHsTASADlyrjh8JAm
Q2E3QprihIr70I2YKFtOUszvDDz/WjJGnpHfSWq0NQ5JUtbw7z370wcB+PlPm9z8uB13XhB+hNxX
fryHYm/DzJ/JEcGQ575p7j52trgHq9sgm9WmNoWa2PLy+F/WrM0/E0JeCCkb03owtbJXveUwFmWy
BnBRzCA+HEPNNEefg9JAJaHnvnrq9dbK38MZD5t9HDwg6c2mILJrrDyafavNRm1gKBrhvxWKQIZd
TsD0IxGyTEbFD8IRNh5s6Mi8YCNEuaVmMh7i7RuWEwxOr95MGffesI95uGNQnbstcEEhPLdOlG0z
EJ14/2pM/P7xYC6oFdZMKzgIasm6ap00rR/7gvH9T9twD3fpZebi0C6Kzv/gthXUM4XoGxGGgIBY
pos9dbZOKibfdPot7aaxsLATKl23peUXF2Y5Oin0sHG9jOJM0gNYw7faDMe4wK+Ogpo/KCqrj01A
CngoUMtCSC2cModjNzT/q9tXJk8jubSNaAPCvKvkPP1O4MPI9lRS/1zotJEWH2N6/oKOaHDEOeFN
vkhMyK/yRGTi2tDQq3CGE3yRsgjOaPcGxy/XD3IkAt1RMY2j/cXn8AHM60vQ/o2+pJxh2Tvk+pB5
yoNU69xOdDLxNM6Bgm2EjlcRe1HE/malg6XSBX7XdNkjH7dP3GMmYMzJwojQZHnKJZPyiURR+v+3
6BecILGqWgLpcWIVZjIRDXoAw4GMLNqeRIwSSmvH5yQ+KW5UZ0Phe39sn+nZt6qUwJ96R3CIjLCe
yab2wxztPji7vSfIXwgjRuD3cZQDDbxDdS1VnHZ9RoeMA/hK0VLYK/a9uE0xHiSLyLmOwuAcNBoh
AIBJrLErqZsiOq4oh9ZTFe7IFqb94Nu21b5cQUPeCralkdrzPj77iGnwMPlW8Hi+LiaoG7BQVF5R
98e8vqu2xiMwCqMkymx2d6I3mzMq1hqdx4K0T0RCKgD0YncbcrqjvtP5q8xJn6dly1+hFM9OryJA
UO4R34QY5NWM6XsaO7Pd56lMS4XRDiytZqoB+1g+TjM366VTMOn7DEdS+VltD8xqdqjLN1fSAue6
cv27dzLfUXq69iaOfM3e02VCjjNMyz37hWxIz7YAOfobW34uTJ5qEa78k4/mcsaIiyTT7ZpzXxqX
Lj0ArySYAeAVF+xCNQIi/baKOjX1dX5eC3B7hx/ykflLSC6bJoKsENDE2yRRJjFiwDxGZ1OYaOBP
8Vj11LaeikiUQcsO+r6LEQI1jDsdzybrv8Tqkw/iyc3MaWOz47tMqC2LJyTCOG/lfCIy+gWsWfzu
UgpjaUtnSu+gUD6YtnH8wnpgsy1R34ebCPoIxeHGwtnOwF1qfmBE1/1+MM4Hypz0Y2uXmlZANe2O
WsorMugpv/pF0VFYsHpg8guDaT0XCYf4euYQunzzTvtlXvyBshGk47eGTUk9c3ux5eyG7HPQp//O
uIGGPIa/TDr9UI2g7gYmsZJAfWu3in7rQXLqXs6MoWw24vDP7amjzXzIxewghoBgkDyiWQLwiWb1
wYxNxB8/Tho+PXc4puvDvWocTfcxPH8DxutO/lAsPfzdX6fE02GTD/3GEqOP67rT8cn0GW9RCNM2
0DocOMdRykfcPJyQuN8lLLh1eOXdVLgKbGWuJTYmj5k/vKd88lRu867nmDnZaWhy8EVUfQTQakx6
ZAdP1fQaSF7WfTk5o4mskDH0bio1uT0ccIRS/YXtA/b+twFIPU3L8Wg/XaDzn7Ne4gdq+f9GhWQ9
O813/eWHsq8X99cgvyVVPJoaiRBCU7IJyH5hjegble60tTbI2iNBtqlAUsLOsTYi1D9xiJBM0eJ9
zpnqYLaiSYFVre44BNJvoz+G+6rLebJvh6FSLrhii6QqOJDZkp+QWGtnJ9vVRMRk6OYhpDd54QMH
TY9zs39cpv8BH95n1OD3/ZZaN+8mgbb91KIBXhKYI1GJFQNG9NrNLT8tBXcLxM3di3dKbbuECuIx
KEgLJZh8ZRL92DXsLchsUTcGPi4357LsO3+qNDBNSW41x5v/5N397/Ek2VOB+VK9fDANECBWXOxt
9vYLskDnLUeN84vnXtCiHVK6WLuEKZl9z53fJc/vdTUn6Do06VkfixB49iHLhyyQO4lSsjbn0kkl
9HVmDbzDKxQPZuSJlNqsPAp5SLttBc909NnXOolGMJ6tmfi1UR+f4PIpDSk6kPdL83+U0mTDfNgl
NVZibLM8FY8fqVaaRGdjsicYAALlPV4Y1gpRWqeSN87uoUQbKjiO2xwJJ3LPaRL0GMHjZ2LG7cfK
kE0AtoTi+8cdd4uyja3Hv/eAoBGVScpCeuD/gli1rP+bKKmUd/hCVldVGU38w97BMFQCPfhTG69c
aHiw3zAQcoSJBprbubz/zm+rjChb/k7ME9RoVut3/SgakZT97f9GMtnbIYo0WcimX/2VwyDUexJI
tO6qrmbtRZqq0CWZHFYBlLNBCI5zS3rBl/gmYxH4V6D+o940+TVp7tmWfYDe/NUNzcUpDokzahAF
KRecL32el5hYhtj4TKW6iIydHRqPqPPdce3BDfoYOwS5afm3jWHxOrgs2aRlKdvbGMBsXOck0k6l
3AAcvfkCieDXLG9Gz0WGBgh2XQANNB/nf7Nmmo5jf7UEfMqnAVW5JslGPBBIrbydFMI8RKAI76/l
qasGU0dN2stKYkH3CJv/c/FwX7yCgRajVnGF3ggieaupr5oYr2iKoylBKMpE5Fv5L5zZuZMw4Q7l
QdUdTH/KHKarzHM5zBjifF84F7KnBBLVPRf82b3Vvv6IIwVZCdotI7FpbzANxzIaKuw1WyOoon/o
TPkbEN/5haVOlSb4KxjphZcVV3nJ0GUL+LMki2vFKLVKTX9sSrNYvdz89ryMVsMCZ9Yy9kVh81O8
ySd02TIyZkTlpSkkVoCdtdmJ7l7LXma0maDYnMv5ncL3EHBZZYc6jBIY0jQQKJXfRAIHv/MKAKqN
8XFNQ9SPOvGDoc40cVDn8ZckycyJ9q8EAt9noUUtt1q7Lgk/AjTnZFNePThAVfvh13l3t0ftIxmd
GDA5GWfiiHGVdo4SsSSMbFjVAij1++IW/nU7el2thwrWNoQpPOPB/voHm5C5TO2YykCic8Uo0bLb
AH1G41RjSBKsHyU/Y6aRt3B8AHgwygNNre3KNCc1IBi/9cUFp+yy2WhCMAr5CffdPQTBhURsUJMz
cX5gu8ApkLqRFcjM5lEx2+2V+WSDhMNfzkQ3b73N0BusetAC2JmJldc1JCNIOFU9k+SUkT7i1aII
xAZutqjSMIOirQA5wMCYbyNmAi1e83Xk9kHkkR9SXympDsYPcrbjqdB3k61ybpG0vhXE/0IjlPdb
zjP/JxwPBVqSuCM2I6/AQqs6XLvQ7+DbT9kFSZYiH2GpRGmMoCCvq10gAXW3T8zo2vEzK+q7gz78
38zU51DB6kuR8hEm+igvcnMQ+MwRClfSqOzVwpCLbihRWBWFgA2lORrXIHAopUgbrUibywyejUK+
mVV3P1vPJa+XQPuP1vPpIHh0kc3FVFFdl1/F8pP+fsO51R0Kdqthw8uP7ylMAWV7u2U4oxX+Svbj
lTLTUAWCJ1RSDSgnKJ8By6Mzqv+JJAnb8tXWPEB7gBWNhaKsbB9zxaTdnlbs9l6bR1o6U1kBEGm3
G3MxWAFqQpNdBYXNJDM2RIwkeDuKJsKXqmT0REWwKw0MFXXztTs+7nnpAklTSlYz3LMaNiLMuZsZ
C5t8gn4JOOJw+CnqVh1Lv+/d/j2oxc8QeFjl86+A5XhaDY04ymJo/ViQpQ11/3uXzvLLlp6srb7h
SLqc1bD45PhHSFqeKhpEVZzuxO32aOkGarIQQEox1ErhTYMHDbBGidpQSaflz34rs5A9LTHjzRC/
FFlCkFly3j5DstnkPOjcayoh5sveei8AYPr/csJxhMYQunmF3WlyNrMxwwh50+SeFb/cQqrvH+DK
LLaX3NykJiZ6UmuNdB97WFDauHRnZslA9smsPz8uaUjaOD+NlisNaub4z3V+fp54MWrcVjvRYrGD
yVALil2d9/79wJVoR3sV3UVCcPh6PDJY3VGKwrL3LOdrIeRffI13QrXSHcslL/Y3s9t44bJBAt0s
UV3Y0RF17xIrhgCKCc8xsFQxdekPMgI414wJdWSbysqkfqCRK7vGoWcPQbigLmPn9LcxACRFRNKC
4AEB7opc6vtL8PVzjuGd7mZshky+ICoyo8Y0wZ5Nhq07uRVqkQjRQy6HKxYsS9u/pBa+AQxkDhC0
a8urU6Q+6UAsCerv/RnJXtJmQZ5IQZEfYrydxIYp+kO2W9R/idFqwyyzH06vMQ5BGy2lrjEVeRUK
RtmrbUHH8mrbB43UPy3EQIJ01uecIbO2Mgs/F3g1raBP+LAgbG8Pj9lcCWKrASKt5KFDkeX/xu+4
T9UbufxRmEYjOTXMfqBZK5DPIxyKDGr/8uw8/iMlJEgBa+ONDF3ZEybJCCgV/dte0YNFuhnjSQAO
dlAk1eb4YK9diuy6V65k8hXlKCnfOQ2zeUbt+EoHWDj8N1e2LVMRdSlokmI1vJxoIdWzya1kRpfy
PXkehliGua6ECRqtwAcAydcxTrGuGsBzRtmkux8tCqQdAdsVEvhCLagdSWNGbVPOXvFkvX7XEQCr
sKq68TdOac2RuqHOSRW1dej4+FKMX/1Rx9GItAbD9WDRPAS08ndYFpP/DPgQtnMDnmJYRPy1Esl7
mtjgngs1kW0KeSD8M8W9/OU5yX7voVIQIQHW0tYG29B0hZ5wrcoanflmX9nqy+CvQuFzVug3qOgz
kZ2MtxEmugeavGJvzGyYcaq+MP1LpY80M/pobsPtFK/thziUInr3B47hBw2SOyt3zetWyYaCqkzM
0acxTlCFapBQGpdGL0pYlFPKFRhyTi/JPVBBHpzpyNj7Cpoevtycv3CPpLcW44C1F5PPxKqhAB9n
fAX0hBkM/yOL/BNrif+/54pmMcHFotdEFrB0KdmsAiA3mQZAj+/oIuZ3wDv8iUMmpBdP7KLcGp39
K9r1exzJWG4qSpmr/Vt9sabdZF8pgbcHWNMT/quBRcYuNPv+wnKnPMRTc2vElESPQAhNBUox84Os
9rQRI7M2aTeKT+0n+MVj+Pg5n9V6G5wYdZDkRnhG4Fa/XRSTC58In5ZQujKuufPA5CxiGA0HH47a
ZbsMHYp5N0d6gtpAcbGPz/kDQr1TEgJMETetqzpC1JiiV5Mc7xM7OKmOc0FeuKL4utSiClRd45kj
JYm+g644ygXN9r/SPbXw1FT3IybxTheAuSaER4TfV63XWtYu8VOGJ16YwPtY4xAel4sFgdEr0yok
YIiY7nlkQoSdr6oH/Sw7vsM8IesFRQ+BzIeFF9O0E1YkuSOkZaENBzDQtrkpwEpvlzxDQbJ5P8NA
8UiUeBk5eltuzGpiWWtCr4mUm97qsFx3PbiB9kgLyrchKqNvVCZfAJTnQZhynCEl4pwqzFdB02G1
X7ZEyxI9oVd0iTYWWoG8AJjUeO/gbAX/OqnlLMpi2y4JPFQrkTMFakxlMi2nVyGqSE3AS1oyBAQR
LM5PJ0wt2AD5XvdLuw3WkzGUVZh4UzfSCGRuAd1M4udq442h8hyDPg9f9s/T4ikazjD6KOHmbBTX
WrcoqpSjfgbY0VBEw7Hi8AR+17Lnk/4t4QWHgBBboYxqFWc0snkL6CAvh3bFESg2fBB5ZExYZIWb
Vgl+tsJfuEXpMnt0lWCw/r5cCgMvPtlTh9ueGJWohUMweU77RUsGTbeyT5cIuSRYiq5GBTSAOooq
Xepjnw6RZjgryFR335pmSpXev+XpOgRteu57v1XtsXQ+0K+P+pGFkooaBneuXuFZbj8Dy40lDhnS
MdjtO4kpsJUz6X1CMtuClolPWa/oarkaZYy34X2i8U6Ylk02BAa5J7wbt8Rqka8cgg4B4Xuj7bwg
SzEkZokfqPb82m7Zp0Gy44pKFkqYf9xmtteFS7KciYeMouBrnehFhcVhR9MHllKL5ZU3+APEJokp
lH6odbrsVqijbIQVKUZ4cNbOhE39aCWDiQnIVH9dfKjUdnR1eg+edstBneDKFvQ8+LYo4MfAiVcO
3ziDV/nhBLu9amfZSAAN13P2AYVlcdgPVaEUW4j+6Ui6nVfQ7qK+ZNdnLGBvEFeriFkDFEXBKTlx
9mzNSiNwtT2VS3mCjBSXDybJD+5r3hIbkbHvWZF2eUgusyOnKSn+5GrE2CmAZXxQw6lBhjJL/Jy/
rA2VSUtjwjTvqqsW0deR2yfmqXh/JWxW8tFOjetXnu9EZqL43izkwfMv8zOWxfXuQ/PRWW43dheh
XRNs35RcwqW66GAK4L67CeOXphWw9fkbGTNKQLhVNHPSe/OCJSP0H9Ju12k8ykVblSC62i4+PicA
8hKARnZmZ5Fihs4jgyElUME2C6TUeHNdKWhayloDV1TxaPZW2LDuH4VkcTsmxmNCUP5CHX6Hqb2z
HOMuV6u56nvOxmXWKLMzLW3xLi4l55QekbADOE8LeRYDG961ZXmSF1NcdAzkw+ioLUqt/1svYKEq
zTHF6peOL2NmijFyY2Skq743RM9lmKBJgrgX1/ww60XZe1dgUupDinAzeIOgUA2PzGXMB5IqffQq
cg+LoiGo77g+zrTA3thF4niKfbFOLnQewTY9c8eLdfpLVb1Wn+qDdLQK6bugVg9lOA3nqUV1fLTK
kClRKCb+gzVKThE9ZD684YDBkDcIBz8SxGFJwTIXUg81MCYBrbQUOSBCkNGeKrwo4sGjdM13Rw/w
XjcQXosbPxBDPVzu+i19onQNCvMXrAPLqVYhChAPlt3pZmJclLGx4Gd4oC9fLYJcE2KxTXa2yzUC
eQJBxOjikA+uOdnD1XVSysilB/ud0K31JYxXcIK1oh++YkfQCjr5BIWnX0YRBC0YTezHxfKPjx/I
Iv272vbdSxJINrDQ7o7snyTGBdRx9yK73hqFW33/JVy2k8f1Uq8yBRhFRxw28avXfkpLfnKJxjqY
Zfypk4RnJaYyK74begQznNheCqAW4AbNFfPc+74B7hOENbmnyC7jFyNkAdFh1OcvzmREQ5uH2NhW
TLlSRRsOIsmuRaS8M8OuaOR70k7KA9lWCC6jziTaYwOws50zRz/G7EEltjfp9qDU6KhdVHfLwBgW
JjzPt0OCtkK+NIDxArjlwln3aeqyJpj7g50+/MZreTcS/ZNS/DpK9c9jdCY8KwPQCWW57YjNfzTW
MLSL5GDnoWauqVfpoFhdQJcXcvFgOdUAK6AGzm8aXEs6D1PM9S3gC+oVQVjXozHoXflalbILL2gu
/juIRZ7wvPAqLhFLjxJJ7aOeWzWM8XfEnsP8NyNxHFU25GhqXYsVp2Rz3HaubgE+eJAJmNJKUJ1S
DMuofDqfteJ1xfaj59oDrOFav6TQoBy/1tUpGFkLewc6AC+1ky0dfmBXkgGoWuW5xmgORgFvsWky
mmAQjkpgOnW9nwv5mmAtt+TaE1UtqY/nh55Qrtz7/TuN/+P4aY56F3mQEsbT1OM21tMEfMoRQ2Sn
yfbWIFHGVP+9dwPdKY+PdAJJSGCWpa0d+tF5toFfjpZwh1K+QKp5/icmqlQz6NZNFp7uj3/93RfC
47TP7DGlLb0jCYv+hw/H2tsFyFH3zW2J1iNIaHHDcLFO0o8Ycu/PZTWwyM54i+tN8L8Vtmyti7Fg
vqkcMxx+ViccPeIKxXZzaDmqM6NF/XwmDKBv5sxCeI8OiNaytMtZMu61sPi3bvsNoypzJfYi7Pqk
XXnWmZcQFxskpnDWg0DlpfpcZ8Wdln6V6ZdGcu0Ft+Czr0LelAJ6FTFofZ+1Z6YH/tgryOWIR7fZ
dAlugO8ZBvJvssa/+m3yJetsxLDLrr92adbD/l5smgKl3Vy6mn5EKANX7y3ragLnZqB11n8StnwI
GeEmf9Xw7Xuj23pBQMPeEcfvqk6JaEmrfFcOc0wEbp3VJ9c8vjI0Jol+dT4zXRtophT9fo1GIgYj
xo9mvHfIRWlAQAstFRBsb7xSWQdI43BuRtCajPfxS19+AQGv7kKd/hk1MuMSU9GDLSblt55Ku6VF
ojoKeuDcm0bjWMhx0AiIIy1TBc6IyeG2h8VaLzCFIsMK7uA5Oqp+pXaB4WwCbdrxG4Ni7e3e2tV4
+DcOtbbYhOViYctGOPJB+m3GHPkRHWeVooB+nKxqceYgOmShgu0m/DzPvw8sbiAf+wZDYURSNMoq
NN6duhb1pkdye3zWGf+GASFryPpTk63q93QMTMDEm6m8Ou3A2quxSCo5EDsblW/yXuf4GJIE+r4O
+/5SZO5rt3Ax7DewP+1CiX45WPkCEt+lwRJMC7H1HXUbg5s0Hg3HZEywkOhT5k5nKvJxWIthnp3n
mv3Vinm+MzTmcyPS0KbifTPY9AHJmYC3kSjopAiS5GQKvE4jw6EUC+Ulc2pXcqx+5rQeDhdpcmAV
+BIeEuxAZsxzvTbNo5HPqRmEvaWl/U9l9RTMJ6qRpVJi/ZLv++gyeyjv6/Q26i7TyKhnoLdyiqOQ
a9iJ8csTCipWdkBGokcRZjHEUvwqmi7CxqQZGNNVz6Z8PpXIYOrEU0Z166yAWOo7gydgPCCKSsRd
/Ua6gshqXRQkaEoHNksu2YWyhwyXruAdHMUqjgbJgJXuxUu3mkXbY8TU8r6smCx/W5qrIvdpSXfj
2py4EvbsRaWxbVjYD/SyKqqs7ERz2tUKCpchS/v1g4Txgv/ABzhnzBS1zdUyaM9HvGL4G/FKSfp2
b7OcxopZPkNP4n7Je0j3iK35mXOXO+L+OmPxn2MrkCtRD0GG3dsuL5XRXm91vDjoCi0B/Dsf9y0U
Qf701m+MN35Kx25f+UYNmlEv5+RQIcRjefzNT+LCg1WBQVb7io7i6EEk4fDjcujUO2tzg6xCR8Eb
+f56K71kg1igW9cIeqKdBBz2qd2XSWsko6XWpMaCnmW05sYhq5Dhx48bI1OqmSsipVVFiA3Yj5zt
YPPYafXCqHA5En+QNwI7OpQnkE2Ont9C5GXhSd4ulsOfaLadiKYPtQu5othrA1ub/QTgYDCy5/Bz
ss3g6AVzOOsK/MlnGCD0b46ice2wHZ48nVyUkQuM2/dW5ClbthhU/AuDItUC5GqQCvUpeTK6bNk+
XcS8oYBDVQWV9rToB0ve8ORqbBkMvpCKEIbKNmYXykO+WGRJxYEj/rkyLgHXZLu7tD4H20CwfmAG
qEDndMTs+RI0t+Lj3H0eMVFpuKr76HtWv7s7BhYyPkgSbBavqrvza8E/X9L5jio0vQ4AuhaISZ8n
acclVN0rnJGFni7lLP5HapuIbxzZsVQAZ0OyolHvMQHfJQ7pfZCyn6/OXBkoDHtsZCiMhmFPycRQ
M2cqbHARiaK2qnKsyhvjobIdQffUnHLSzeJOzqTZtnWnyjm6FXlVdstlcIHvFhICllLCjy8e3b+F
6UDHIcNPa3xEiFwfRWZW0szMN0VQowAmf2jM1pCH4VlV9gX3t8PXW6DbAoz/xhx1vXdtBCm9R6hE
xcSxI9XmcJ/6YmmCLW3f089rbUpRsKaQnVE45608CntJsBFQakMOVgphiMLSU3V4wn68XpTbGTmE
TH7UeiMZF1gd0YUUrGgFqfN1n1PhcTdPheFTF8+6fBG46Zu/NccoWbCcp/UBJ/Gm/aXxpNExnZ3F
WJOFvSOmqRi66W3HOvO7JKkX2oCV3pOLGhGn0FCWZ0uYC7oc9CdsxkZ3w1qkj0izzmKjGigwtEuw
ZwSxrQYuZkItZgG+esZV/r2RYDMzZ3d17dAnKafzH39KLZmuve76E3bbEpad0Qbyg7TGj1JEDXFA
y8v2PixAcxY5iKBWufISddB/Umv8jb7QEuh3kAEYeXUkAfgs40PDwms3QlTaypnCAHEdxFljBfIz
1V7A5tTp/04RUdjlbxsEG3L23SgfYrXXFu+vrN2VKzHZqbICOmC+1Jv1xsYlrKUsePTTJ72FE3oK
nkLI2XCWAvTZvYrCoaaqzAcW12VtVofCL2LKcCT94+KkPDpgyqOxe6MPAZis6Kx7/+oKB4h1MI81
e/CO0B7Rw6W37ZaDcH2rzyJmWqMSPdxtQ1IuLlvqFDdAucKrw7CemUZQb6FvqqJV164/E1wypjau
qX3dZzji+Z3doHIbicZK6hAM1TGDEf6TGzVwWQ48/d61Us7APrK2uEKiU0oKToC+uzwJpubKa7Do
MJZdqByzvJ+D74vXWSu5PdNEx8ehe5IyjmxpoJ5JmK0s6AOylnt3Zw82cJTsYrwOXcKLz3Vdi4lF
+joH2I8oylc754KCB45sPxpoSvxYwkB6MokiliUzcwK+U4IZGzzw2nu+Uyui+AHLHbyooVwej5PS
4pP4nU9h1wB9HZlLIw3/9Xz9l53cHpK4bdvWVc9MP80S0PjvwyzAlxKOPAfOubZp+th5q9ryVBD8
rWYRPyBPjHQXU5K8Gyz0RPh/Tf0lAsKb5DGfgf96+izKtDUGNarKkbqzWxLuYu5Ud6tjPx6PyKg3
75vGYmyy26tkDQh+grqrLYN26MRDODIxJmZ5e56WUk4aYCVxSYvmt81k8PXyL5J6p8T+AT870qQ/
oJPkjA+8nX2JxvXGBsMAskoL15+XNBkAylvy+Dgl+P/wPEXsoOAkJEJA1McgWnf6UHtMQFcAG0s6
V+wIJ+zegGh297lINssEWQw4kcSkOdHOB44K2gJT6G6Z+4hp+3pDuOxGPjG0lG3QguEp2liZgJj7
ou5lpPTxlljIt0yhNC9lSCT3p+SyPb6t3Y2q392KvfJGdME695igDEebwE/FP1DIo7xEonxDEFWz
HYiEashsnj4llexSWxdiL8V3APlQ407eDm3Bxn7hLWLxgAMMf8rccej/gnpmemOZNpJXIeUeQysN
TMnBEV2yDMMQuNMtBN1W09ExS02kuKjoLfXsXxv7zNQyoN1bJmiclhSNkMap1Ru09IseHpmbsY8S
zX7k/DbqgbcgjUiIu9owpJZBnoau+UVUV78+HANJd2DvXCgVAO/sYl3DoS4NpVEPf5MeXRtJPdu4
5ZT6+pgxOFslaAe47Uciex2C9HS/GSQIeRt585xJ17unYu660lEh9DNpJ6k7LbzPMJ2W0o2dMhEU
gP3m3yMQwmPpCASconCx5PmXl67ZSnvbt+YyOoKdfDD0zTV871IsGUhHBeHvLISXFOzCsMtBR53l
KWB6hbRztmdkTJeDqD5FiefUKDvNir0ixpJdVGTBVGxp0Nt5UfVBV+dJQTVlVmsk/hqw1ffpjFvk
jdpAuySgamKfrcDP5vPrnV3Ya7L31O03OjcGMKpnWIBai51Rw19Qt9wNEUP2t9bIIhIXB9yyxwH7
ux8JsSUCMTBg8B+XaYL/Xk9zxAO7esi8quzZMMYag1Ih+HAN34SQt8Unko1iQbZP5iNQE5YxnmLo
fqZGMUa4PfLUzSxH9cPuWUaPAF1TFKddBk8EBRuRTExs7dgYwSqsV7f3olH0+L92FqH+ArZC0g+V
dZSvCM/FoOf81VMVNcW6qR5g48Ap8ZmM5pkKOKIXU2itI5hHXQMPCX/wfsQiGx0hMfMd7J6+iN3m
Et1D7Vm0/nrrz+PfqQ1CvVk0ipyiz752WK2gGv53bW+Sit8Wfqx/btLpgUR35VK1e4qAr1I0f3Ff
PWMNi8juViV00l55hA8SlsRbiFsy/z9FBzN6mQeo351S5qc3M0pJvVS1GZx9Hom/6MHP/yTSUQJa
1X2M0lwahpIeN6zicK3E7m1CDYLBDWM9t5UVe9AIjAC/OpT5/MVwpuUOnQFT2wo/N9xihEV7EePz
yBS3nXs/gbFQBBl+VSbxIt7E/N0dqlZbLaeXmyFSxMuPk3vufHHl3I0f1zCQe1wosDCxe+DXuJce
5jO2yEGi3xQXrnkD8eDewtJkUsELnPoDXoctW/HoONEnUWfpzg20DMISXjjDzNX970X9eEQvscdX
KMVY/p3a6NgataNyAzzbaOSoZm7htTrEahni4vK6PktKQWmNkhdybUbBiceSOvjKfBYPj3SxxIAJ
z42aWzLZFBx2viNYB4d9FaHo0vvGguEGTQY5K55JySRR123ZmVeXORgIYQu9plIYCqTXniMuQNJA
hUMmS1I36+CbWN1N5onAgzGB8FJIO90xKqvbhyy8llJzSRiv5WmFJb4vRMbMOHFLxm1xnnYUwbNr
Va1ofkCXNJ/407cglqIk65VvBW4a6Qqmt71hPVgdshapTRu51AziiY/u8UvawctVBKGeXNxeRnV+
+ZcamI8b0JzJp1ow0tpBMxGWk/F/rXR4TyIsF39xNJAqbx61SSkdX5Uy3yUGQ4gHQK6VBppnOQvb
j9fqWKtW0iqmny3I/OUSG5g5h7rD/wcPjnbW2fhw+ZyVhjnnhaBXXvkGkFeLq3qQ/RfSuiufTK04
metZvG0h82D2eKSCSOXfoxWbnp8vnpA1nhcI84aaQlkPn0oJFBTGvIf0HeBgJd9g+VPgzOi3AOIf
ZwnfXbArnqGQGOjBzQ18244jgpFbDeSkaEIKY+mg3rGDIfktT53nOOVDAds2BsQpDDVqFYbWVKeS
moiMz1Y2uHY+zcFEpZyxjmEDvmOgtTqBNPEcE1xS/E0TnQCctMQltQ6NQstUDkVze0A6pPh9ZqiW
uTkZUKuortCOI1cDNiPn3XEEGKB8TNAxTCtQIoBwydwOdjaNr8eYdf5seBpgkyL+zdPrr8RelNE6
YFnOxM6mKPgEYq0xsjF6q82dsDeHSLr+rw3pBojvJgEZz3k0lqDTY5FazI5wNelhH1yJiWFnpKYY
DMir2LMaykJbbHIgnZliVt0ANd6MwbJ4a40FkAljUekbcN7vCtMaDDhCJ4JxSoXk0A/AgoGjTRiN
nLcDBSpSuhU+Uj5uZXlkpN6A+FeTOuVNGP0wXGRVO40mhu5+z16rJZ0BljEWZaKj3iI/PnOtg6O1
ijN/u3Vsn6gBmruk8j6HaZ0MJa9p+moIIDgGLbF1yscMO7DmucykQtyPR9H/A/Ab2z5XiCWiaiB6
KElRinVAQKLqARoL8iPNo8ZPEHhl1AwWRH9CoizdZMaL7AgXUZ81juJAJGYPlbFnHcTUQdNn94j3
gOtLfzgxaKwgNkUYuQBrcIRKByI6aj/m6nM3m5inO0aRqZmMw94QsOP0SM1um77SXgywMXu5MJxd
7xq3TWCGZ8/qIZywPSvJpdzyxd5EDdCXFye8gI6oA3wfGyNzePA0TjQdV0MJq3GTLgGQBa2kVllj
ASyhz2AfE2G96bJCf6fs2Chzg0lfgryUBRH8ktqVzhAoBHASIEJm3ThuNI8UBScF04se31xXSf0O
g+BhF1QQU0ohbvjR4aqeAMnKJ8N5AFZv9/F6kSxnLofbcwhosWgIcZvCjEnUnagtSUCMqakksJQL
vy1SYf/5FMXe7ztVJWtqHQqizRRVIh931ac1LE0Bkokl3uaSNTWlwu9GE5/idih26EThtOmuic8c
f2uHp99LtymEOp0ShLrUKgKRxQd4sAshJtlNNZnuDBfzqtftu42j96rtksopY84p2Cn1jBnDVhvO
ytfpw4lzMva/gUWNKDnDUupoPY9NZ7HRHsNfkpyCgOWto0nJJZG88lU/kJd0PXv1j6ohLqkloApL
oTi2UWIsrjNzj/41v2+AEIFEsEgF9I1oE2J3T4SVRk2ICaVFH5kmV2nVGWIfXpxrZ9KFRDz9DEKE
F773DeCVNadAtcwFe919+7bBhSWTIWq4tm1Pfdjz1J+Zp3GHPGeihOdRUIcB/KOVfHS7Fd/peSsR
wSSQY3D288hk1UqJ8B/3a+mphsahMeRXdk9JMQYHOwlBpaMJ2EwhFrzTv4t5f/OfDcfKmK2IwR0o
XwkPXZObvuOcRDNoh3FaqvEpNqjJMJO0yUNjCUWVagOdpUPInSn2G63GGsuND/1YDhyBS9ziqIF4
G0RXs6dO3bKFz1ovT9wtMvpgwuFVqZ9vV7wS3lxyY5IzpcBjEyjoxo5D+Az9XVWz4Nxmr+ztDzQN
mRd3mh6FjMyKRIGZg4GELBnDrodGhjRlMh7QPZknyotoQ0022//J+szTWGI/7FwZSSTbmjIfMqdo
mvwOTfRdsbi++EsMpbjB6rhIlDJQcLbLcWCo/KyQ9DhGIcQ7BNrBFdKqVUBHh/wMxbwal7ZUhsVM
y9AeW3H8erCvQfc8p7gqNqdcD5m+KEwtNhfCjhhvkZcdArKGkuo5A84TrA+u9LcRF66OQhSKggm4
0nuwGHS9ubAAsC3gLJfp+yCNoLgsewyssS+/yNlMqbcKkiIjKaC27vKbWhBLR5fgLlcwFuX/7yub
9PAJRBCo34pReMC2Z82eaIMrScYMpUHPH9xzNueoXZMxJmtaZEPcjNs/9xNEHphwHiivb/UrrqeD
wJ8DhrBkaIWS/43o9xsb127yApcSERp31o4TDARvnW1rlavSWCOdCZYOhcO62XnLZCZKIkqSt7S9
vRuhnNkcGg9x0J6gJHliE/oCsY/Xx8gHdfkDE/4tB7vW7qU9QwF6nvVpLmNcpugEvp46n3YQ7fY2
iN6kMCGwVWuLbi3rnODNeZ+rrH7oqldfbRE5nWLmvDWHCIQpdqDwQCgSqXIcQHJ/fAJdlyZsyj2+
esTyVPYMTwjEK4c+JbK6PxCrlSkBVXaYN5ghGhExGk3go4jPXDM9U8uUB8P8mja9s8MVII0eIDC6
Xk+plXkqFT+jnZZizOpz4EASiTM7jA8RCUNXrPVuzLQyoEvre+vksoXTnG9NHUEz9Jx8My1eyKah
jEgQPJoswAYJvGJHeHKlxU0qaMl7CGZBvgTyjMUafDYxL/g3KrDGuCEj6bOiN5mTT6uOwm2gsNC4
CKxiNotIizn8RbvmohHTMyAfi/5MDZYqQyw74FKVdoVPMbjL22y/ghwgRm067AuUlC8X4ifmzrik
fC+y03ULOno0J3LKYrgMEXdRPCRx0na7DrAdAWvLq4Y36j2e0oGeU0sBG/QLBoPPxZ6BdLtAI7N1
7k0wLCUeCOky5VUrNlcVQ1y3rRJsbvRYnESsGro5PtJpfVZMlx+phJqkVrppnmMbDc/IKB/t1nAU
8Lc6gajqku9G7VOiapdlULy7YruqnTL+kqwlDforgvcxHK7pePlpdaK5dLqeEnU5Gv7Uld3hrNmT
sDwzrgAuEgYVTaX+zQx6X56j1edaOXcjW9RcjCB6g05Y0M0WVbZLjglqqSLjeyaTLMdJbOB20cdh
shkaurdHxZ5kJL/VG4tfuafC+ORCm+gLAOZT+meplOEAC9IekLRKalB3/7lUpnfnLz4uJnBl1IoZ
Y6TWV/ObW48sc2oB5gkKkZWAMnBfjwtPQHIO4VGOezIXrLkdFGGoP0HARDGDDHtJixy6yW6r/c1P
wyC3F3UhOCmHQjmM0+RAKD3a7cFYsFD0rj4DYiwVO0JgLvIENDcRrW60tBDCPEejXtw/+w5LaD5L
wtISHomH0CN4+mxOYsLgKd8JMlWi+3MKF3iH8L8DitauM6TeqHaBWApCajLQ6VVOP6hSYkg1gVQT
zISYm/IRLkX4qSr3HrxOiVqONQnYMvnzkAN4+IzcqTF6PCT2MuCjLvempawFG1NmF7Sn9tGE3Git
3E6unueRAZDT3lHKza0fRCm0ZZ8BKanp7vk4Xa4t0lN9S4q03UMWjdmigd7ohE6ZKVOYli+qOQ8m
Bkhox8d9EsfLyj0Ez7jsrGsGzQ7UtDiXwSlKsNJWZBECNrHEFFTcn/yIgGf6IMEySJXMb3MFtxP+
Wp9hRx0C7C9Q9PKs/+HGxlGk9u2wFW0d7b1Z4dqhPCFhihbKJv/4+9imonP2OMwkUVCDOUkJlHM9
HfAam3J/17RH9rPZPEpv19owydgbNSemz3Km0C20AipDWWwTr3XZGudCImUUo07xYHVJgfTsf70k
gJg5NIK5S/R9V6l4L+6IE9q2FXgrwAdIj6r7ldJ/FNilCX4ddnMXt7JG8PtwjRdoo6nGAi5E4TNa
LrDuCrhjZxsMd0NqRDVZT14WqDgFTjNPhSVSB0k0DXI1qn/LDM3HlI6JmiQOgSpwStBmOjDAYng+
5YXI6SUdXDaN43nL02TAzjn6SXJ+bjDMm2IaFbOrxrcAf6kY19/vPPRhssNLPZTIP+8dgvFjBx9u
oYKJnMiHpdmGjvF4rgwH8xeglDY+wo2q3rXxwanrO7iNgFQZb+JnqBhImXMPmasvd2n5nxOmAvI0
RAIK47YlXOLCEtI4jPY32gFTJ2UoOHmuKwJlxKl1IH6IDJEIzsXa41EyNv9GuHvu9AvAY/fvqJ+l
pJKT3a5KnLu+ajfARetiUiQ/gbq1pVpQ6Pw0cV7MvL2IHk798w6DUgbYMwdj38uvmU6j7EK1DSAH
m7oFavUJjtKwVV6qYl+1B25EdXyJlYA4otSSAnZKeqWZ/urlcKS170TLGF71eqW5A6HLsj7hcUGB
BJK0WJFXWHcOAEw+p2MRYlW9ETQosshvdQmzZh+fWUS4bfJYetG5Ylan5oSpb3oqxYqjlFalqyLF
lkoQ5ZDrDuMJ62ozJu40e963SgMW7F5LSrcRkE5TAhwnriwMeY2Uu8WQ+NvjgOENKvgebjlJRQy1
TQyVTvvp9j6Tz5Bs+aLQbMtVA5XsS/uCX8oUdklRoVUI716jhQdKkOdO7oFoNbYnsurR0sf5YGEL
6k60BYL8lqimXUIHTzJhqnPsKqbVBJNumDZzWvjMQWEx6MOUT1nQTNSLGGXhGP612gUG82y2i+vy
gQf3pY1vBvvEMN0iAJUgLRG7f0igGJx4SE/rC3TdgZtq3OIk8QG0FgpdINSZ8EhfbrSZmaglxUUo
jyUqrkOrcAR56eNOBg1TWCZJevk6f/qlgbmjKMQAinp62V3YHnKanSVAh888BVbyJooPfFYDbOr8
tkmA5BWM8YXCodN/Hf9GOg7v6HOCbtUyfGkMUsQ7Sn/v/gllb5Vjdn07JJmBP943nJUpbt89HsSc
fXNDAEAijG3e8CCAxixaitpg4+FtYEx7LdC8kzpyMiLUqbZVGXgwJ6TB3eXEFpz5rSBjG91+VUJv
EjAGBFhjbUDOY+O4MQ85giRnI56DPmzQzj0US8O+No31LnoUsiBcI/xcQUm1/onSUXwLgx3jM5+P
shdsgy4jgymynS/zeLB2mc14TIDpZ13bnEy/+WDEe7XLVsmrZFFknx2ehjDNXytx5v6/SKcf9Ian
T8jg0Vt7DkArVyeFOCEOM/7x7Svlw4A7nHxOAMUbYC4fpclIRPEX57HaDNYnl2ivVsFGSmuEkjEM
+9Z5ciiVqU9F2jKOXFMqZU2d2SWMHbrkHqDw8ne8aWhQILsoWu5rJIbO3Yz9ITfTAY3lPq3bDldk
IUCKO8xKgestOPHMBXLlnmHyBRHCvlCsuWXxzDjnYP/DFGJ2BYanDG1su00hwWfTKwJvNA+RKP9b
sa4fyRwwwtdU+fDPICxvOng3shaOv0OpNWRTO2nBeYnRPoVV/5AtjzFQ7Ydyvky8rqyWFvgCGpsu
vRl65jnW0w2Wx30gfMOX2F3UDdVtIaLA/0Z+7nqotmXhVW2+GH/pF3y3e8obu+izTXV2/KkRW/yo
Y2KDaJST+u782p68+pef+X8Gwdbp3bRspTwTBXlbU5uu9XT3OD8RsuZ0sSCzxdLKl9b2b7Om6up/
ytPwgpoX8fPPzbeZm+D4ptoxU6LzpnNKehl4QVqrhgDAy+feqpd5Yh3rqPeaNDh1pAIcI0jIiPej
WLmNiNJpDyN8n1cWWuqwV6sK9t5QxztRqXmTd5a3zNbrd73YoZ5ChWiuZtKKt9jNxlE7TNyH3E/O
J8ic0BckT+FPc6QW3lPtDNJpScyA/PgLpZv2BEVHdALePsxCqxQXLPbxKR0IlfI+kRIcncznF/ue
H1CMAAGet4ldVDfSLc0OvjietX6uoMkVTnNwkpB5Ohn5tTSL294n8UAsmN+Qc/E9/3G7ODcRU2Xn
vj5qjDQfzZXNEEVHAXfV080rlS/ysjn/lpfI7a6/QMnz2cFXMKbxeKO1XuSKwON2TXPwD3uriT/w
55bG9bmaHCcpWAcq9lds1aBhV+p60b9Z6Wyt1M+RuE3xVOdW4J8yoPxtXyUEyE834vqb8bhdrPI0
YdWn4gRYpTVl4QeWGH9Jtj+G9UJFEzXdt067QhyzRTH4PysH4BwiuP4SmZgXgVr0LmG3VqPs1Sux
b+XC/aiIG5OIwlFoHGfg70E1veXaEFCr/8n4W3DjSOsvukAytIfXEBgQGMkxWaZTdcZwzNA5NEf/
LGz1I0Y0GPiIWXYktmD9X4QZxAkl0bjEiF5mjqL/CeFUVZR0LLlnef/M1pm+SJ7IHzDvCRRzeDdA
BoBezWypOjuBQEGjELWt+o1mp/cHs7MLqAeoA+ofrheB5VaQKxkzu4pLxTUVZsFoEZMeOtx539ye
cb1cnQFYUEMQLhYF59dOzZLGCh2pP7CBgVhP4ohBUUzRySee81WesR/lePOZjc2DvB72/Zj97lF5
4oSVJB8lIX7dPJqf92edmWKv+xMwMxcL9bQ5YAAzV6Y+X4bTyAuMugi+Hj1g4e5rASn7p1cpS/5P
bAnc6mtmOxqjkg5i9LfbqNe28loGZ8xHyU6ujPhkyD3/qni879MrOdZrH8GGMaEsjr7+UrHA6gqJ
1OuWvEULVxy3VUntwcqkNKr7MoQx9dt782cpoang5ZZQn+50z/I/LuvQ2iumybk7t/VwXTMJH/FN
/7IVU8y/yv/+6Xx8vAZTnnefkGwKn5AZFqbCB3TV6F5zosVcLCSAw88+OjDb9R9KX6t6assj9axB
KhdfwjY82ayDdKa0aFOCgDU0Ls6kP9C7O32W3L6XIRiiFaZr1OrZMVioEopdcfgI/oAWlKEYRbOG
I2bBoyWlD3wnm3m5Jt1TUzXQ40hqTqY2xcibg5lRn66kFQc9AAhOAcma0d+F9E/Rqb9+ltmk2UH6
1R/K+7RZZFx1fjBSNjZbXzeosG3qa8P9A1s7G0abpflBhZ53vXgYN3eu9Bt1sSRV6dBrTCPxTV7F
6co592bBMk3GN2xzpoL5soYHyivkb65xGLV+ohEbOixtp1j+rTcL6eS3orO5TIZy0mPG4ajDOhkG
aWZAbBJUHiDwJ4ZB4HxQHTzyNH/KQUum9+mlpLMoYYsv562TxuC7j2dplj+cQi2prBiHbxi9GwrD
4L9FJiyFw+f/9ov794rs/kmTNptg102/j0vdW6WMBgmXkDK3Wf5/NGgRduHgQxkMUl4ifOnM6i2o
2bGkGBzEtUr1zJFw0Ao/0O8aOpOjGWC0IQrpuTk/OCfw3vkkwhNkFW5OlgiKvDjj6uV0I2qY0grz
pPOFI1ETay6ZjsHsPsZh2zbIA8tnfg6JevDXZASLGyLKqViku/K2cwfuTBk5ALAYb2Y60tT1WDCT
0XSKeMR0XjnMGvbxfywoaWIackjdVMexDB4SXdWQHvmw2Ry0L03c8hT7QdMYZXX2Tm0WkaIrn1cU
0cdo/zY2EELY1GS1/NkO0KL9HNGIx1kDQjMisKOEjAFGx1hFX09ErwFOtIegKFM1+0N81AbmoLMC
pa38MYc3m0L191anD7C7bRkjpNLiTgXnMR3opGX+AeMvc4ksVFsU1DqN2bOurkZhLZ609pzSHf9c
9F+o1xB4jK19UgXWaXx9K8mGuFHxpV+bklsEOSZEaF3fnCPUL4npqxk4AUq3U0pQBJtj6npyee2C
/cQdERHjDdDWoSAHz2D33JtJxoeZaehcxdy3AXD1nkI+2JagruWr7Bpkguf6t7EjWxGmmKbTm1cK
ZNqS01NZH2zeuM3PF/3z37rZwJzm++5t7l9uL62ZCabrb/8TLeblZt8AgNqO58qBawLOp6mijI+S
32152nSDkWBg+yughIKZNIDoolLmD6YlFmdnUaCcfiktmKsXY6vws6ORTyPwCyeO6m5+vHdZA0yK
dGPDF+Rbf4bBKoHCs1c0pavC6PotTulE5e6tmaYnde21m0NGezIiJ7yfzTMgqntsuAlcQwAzOs3Q
jGfk8o4kkH3aDZFBL8UsQKeppCCn+H9Mp++ew7+HZ4lBSsS12mjsWPW+zqazOODOgZ7BFr+pXvEX
jy0fcMZQhfTyyqp5+WC+df4IrUKanOtS1qAbpiNLPjlvzbgoWj3JXo/nT+1jk/+zhVfUY7xVDqND
ftP08G6qq/kyWAoRdkH3rxAhm/1PDyyr+V6WiEYhmOChXmx026bNZjz0UagVMr2tQ7aLGHp5fSXy
iQmoOs6/70OABJNCLv0iNhZjhhjE2GxmQFPlKFOsQSknARze6+OUYpX1pmTI8jDl2/TaYvwtcWSa
N9vcEGZ3wFqXYDtqt1Q6+kQcIm9arlWGBZLVmjdVaOkhnFfXL2jeOomfRlSknBUtnbMrESPI98eo
ttj2yZs2Q3Pls+jdGAOfWRIKbBQqaMR8KFkFgJCQyztnvLUs5C3DsE180IszrBD2P+FQXPqtNZZp
cdc9jC6g6i0oWBvKh4dQYEwDe509ulPRuL+chsrld1CvM9nt8Op6leQ93nS8zozkppEqCnjL+t/r
aF0MTvwuoWe59KbIwCxz9OOfI4lmR4azWnjFyXQpxfiIQ1uOTqqNaDA4GmSIml/LO8Z4z4su1rmm
Vk7LtV+/GOmlDlEYULaPZPiVJUQqG8EPlXcS5cFoeB6SCWmriZXf8qvj86Ulsw9HrgrcOMgYiqm0
rqdYkRAlrVC8eEgFwhcQWQeQKaH2r3Pe9E4/Jo7e+jFKbioFhZF34Jh2zl8PDQIpvdCG4fTQsO4C
Bw+lkpjksz8XyIwy3kaFn1KvFJQLNH7pAxZU445RjcimeV85NADnVIbKXjRXrxSwQWtTYrwd0hGP
r/BJW5ng72ajovaLQwwgNufEQndPaJhO5XQRFbVIwyWTRCK2jc32npn1GCHODYhfGqDgWIPnj2VR
ijn+Oqe9dpUXVG8N5dMmPzc0NFq7ipWMTRLvl60dhDQH3/Tmd0oTpsqZvj8ua7orfSk8XuUQ2IrZ
PuJiQfbJIv0Tv/hCwshdK6DrKtL/704+miQ6YhBFE/HW10bYRNwJJuCkax4OPZhZy9xI1A17rdfo
5FJtG6vJL3A6J63bCxPjrBctqc6k97jp/iI8+U4z5cvwsaCdJ9Nk2bHwm4qdQKGI46P37/tYS26Z
BHz3a9qXwFUOR4uUrrb9Y66bVwYsDJYtD9HGCOmvehD0N6Iz3IP23Z9a2uAmLH5jr+zGBPiA0tnR
KkPMmXfuNMtOVMkG8nTdDmPIJGDZZxNnapm1PYTFTVSipJshMT2sX6kRgJWPuYu6kFdIgPiRllJ/
w4VLMiBFTUp84PB1RPH19OUmIAIivO5btLmrnNHoQU4JrjUAIO8XXF7d6zkwBmgQUph65hJ9OXnv
76YpsbN3xUzc9ml+4nTfc1lqH+InVKrZPUmyYy2vxPZsFWRLpUXbavkichVU8SQ78gXOTai7A3cl
A6D+ACckTk+hO/lYGaQDkkSUSvvcD2qGjHnQHTYhY2h6OEAEJIvYCFYkpTJVJVY9DOWJV64TuVJT
i3YDes32xPww2DJeoXy4iedysKHaNaPPIULtIBTKtsLF6sbAewxEODvZLmDLH6FMUbhJuYaPBi5M
acj1x3l1oEeC/3r6GF3HxvtQBJYjNJBkAnodElYQCOhielGCrXUA40zsYOzV509EN+5KZypigBYj
21YbKynOelhf2zetpm2QE3TMnvzqkj8N1Tc2Gc95B7BPvCv/tgxDcLKUotJv6kvopzRZqfONUm87
lhB09dSvtVAsigfWQWGnPqM7SxKNQtE3n0cVJt2F4IgkH/tcuJrJIBlgflqa4AgvV51O7chKoaua
WwLVeLGuRXqShfjPB4dMGdylQh8G2DFSvjj7JfWH+0FwzikNR8YvftRBJ3jhMLltha0aL2cMARQj
OLoFIrcoNlWrkCE+hqyNrXcIqKbv469s6HGrEJAZsiYZOEvv5cgV9RWlgghP8Ds02ZsvkjJYJ8NH
k/uIfMgRH5rVbXn3BCUk7ytcNeExfsh2Fx6+6yIpiTpTQ39QfeKIKvIjqzxSGLZ8HtQJB0ZjvIZ8
29KD9jGFjKxXGVhNSekrj9vLc0SV+9t6j5h7h5xWm8aUblQyvecePNQbTUPvrOUtR2jrZKcuha/0
aUNMOeLvuZRw9wa156C6QpnfTQqabQXWqQKUQJc7zDT77Ka/6fIdu3iY9/XiyD3sW48zmf2zwlpI
MrFxbNGMbH01l4fg2GSN/a4/jEb40tlflQdKkkow7bLDO/tll5Uk3FBORW4HMdUERG3g0Y23NYYM
Dnd0N9N4Na6CN+W3r3oWtUmSxMjkWhe+6lhIw1MYzPWNzfl8xOUwpySgNwEgBd9rF+q889IqmYvx
k0yvv7asheCejpCt/C7Wh2QNN0OoIYFbRYmZTozLI3O1MiyzTT2KWgjoTIt5Fk1ebnmGKrIoPcAO
o94ZS2MeFmbjMy7xBbbRXN3VC1Vm1dL7NMJ7lL4y0DF5orDRRzh7nXQekBVABi1hld57Rj6zTYJj
cMXNUWNW19fREn06UwwFT7s1jj6cZhBTj1diINZfHAWk9AamKtbPlr4ZscqEKmbZ5MZwW3Ep9Jkf
4Y/PABXqXzsaVIghuu22wNmhNmfrdv2AOCA7GVoxn+NLtXjs25fX+OCiNJhfh2JDtN3d4Ijm9Wtd
hzA2sX0FiVfITUY4rlpl1fr4e+QEzEUQPjC5Dd0V+JLi/d5IwnoLKgdwlmNT+lczcQ5GcJC59o6g
MQ5ykpvCEQ3r64thmRX38JMxmtb+d7WyxaejZAnsT6UxaD6+8uu5C+nOPFPyoHSJi2Uw1Xdg4f8D
yFm162nlV9yTf0hssK9aEMPCDeO1+0t+SnGVUi6TraaT5nW7MFakAtyqsJvtEyWbSHu9VWQImrWw
FSoAHtFExPSZ8bhN7LugTmGHt8EVXA00qK4E3dM8FuXwPPkSjBz+FZGQ2cWsqRlH6Wdm6g5LeHxz
HnpI2tsfHs7uViIOWxRXIuZoa5xwt9Z1KgNdSizEcBC5O1vhjYHWsKmCvsF6aYD68ngClA90RCXU
3JGbBphFUJawbyjaOhTNH9+5M+jDrhI/disBr1x6beNrFnESdaUBUf6QH0N5UJhTrEtea7t7N58O
/NMHgwG5qoxG3uWXBM56LuP31gBbAB+cz+F1p2HWku9pluQaTrwPKmKExjIHpcswVpabYq2WHo8Q
0qbfOtof84L7GrI9msfVmryBUCMakkNpeez0CSkcazJMQ+fXB3Y0OeTWH1DO0XAKY2IFHHIIRvbs
zj2LxnPLB6plJFIzcMJmmBc9nvJ4CoTO6xUQ3LZyJsDHQDaB7hPb9RDIWnQtvD4dGiEnSf1d6vwc
dxkIOCHrrVcHBZAx3BUlM4a0fipttEcqJxYfqji2LDPMzDoa5/iztiUv9Xin+g3Je45g3ecThVBh
EDVAa7skc6YtvPkr1nVtMuKlLQZ4IHXB2PVJ+hD93E+gIDMaLrIW1ccRCzj6bCAMlm0m4/fBB4/d
IzlT7We52lYHGzdaAQg6q7AcdOqCYEOUsTTEXBNpZBtDlqMo5wqu0griNS+SxZyDNCjeUs8OFTSQ
L82v7pyu51QSYQr4jwyxhiQYRj1Ypn/3uhLYAZOtEAQ5leJJDHj7VgenTf7KfNp9/8zZ1EyVfR4Y
tAWaj76Gv1YZc8DZwxauUWYsEdIBN4wtu3iZ1AofoOUQgQQ1tsBI2e+77ozs36Pw+AbJ3Wsgv17J
mihLAXSoZDWgSxVVQCWB7uMLlxasJnFQTJC0SvLlsd0CNL1vFqK6UzjuxDvi1UBRDxH1isugcG5n
0BeXlJQlKDcCz/LiTEsybj1qRssS/ecTWOMYvE802mkqDyI/9MhLxvZfUn+Qk9C/Njm3fn/SUyuf
kyLqh3ja4PTTilfmsasZBTSayr14zzPR4clxocMG6c7tjsrCCUp2FOvzeMH40mjrpENWsx/bShoz
F6P4NQ7lHOJBEk501cyZk6W9ibOR5cyv+eCe9ohhqsqZe1YE9Qf2eP3PDZmPL3hld1JPifYLJHQf
TMhL/F7tault7q5JVjXmv+EXXSyfZ4VPbxqwqXWXb1kT5eEsoza95YavwotH6xp5YZhzfUrBqXcq
pYbftPkw7L7jMWQ4neNMTCgM1XClKrLVHi9zaHwpGU935uqoLMNxXZXPYcmFCFN5srjc9gq+IlVC
wTKoTFBnLr3kk1dFDhZfc3PL+Q7n5HQlEjsT4DUBdy8O/hJhvZsMb16TzCDgtD/0WkQVnNGjx4Ea
yU56QhQI3M5hbhtDAO4w20tgQnHeVDJVTOIZX0bnlFOwKJ0q7sgXNm8peNzs2BHyBEvrbOEJGxrF
/AVJ8SVyYcAKYvHuKU5/TLXmMIw52SCuQFpAe5Ze0wnf2plY4yGtoxz9KxT8eaJUauu5N6NbcouU
YyeWEHT9eHyfoxbatqOeRNfSQT9Uq+5srHSHLdnc4hBWiMNdjS6eUi+GuWuqwxrQKjrZmXCD8dGa
toGkySwynU4sQKPMNPauXpSaB6qFjHt7D1OkaeLBa/3K2gfTaEiIqHHtRmWMrFOsNGI4XbmM1ODn
wL+GIyfeYRDS/Kpy5TwSlz2PjwIQuk8awyXklU45ZREL1Kqmz9lF6jg8Lgu5rpedSUVIfqsSd637
pkXiivs+E1UYc064pVnc1IOV3KtiyoKPbZTU+m/gCldj4hDXXgLCA9Td+a1hDxSccLp5hjFtPzOr
1xm2G/ATYio4ypWGgejcAm7dokI7Q+fBd5Am0vcV6yYML7rsb0TsPFpjt1ypLM+i950VPTUl3o+h
5gOUPmg41AMDCXdErhA4d1tDvDs4yjJjoQHtwWpS0lRv8OaLEJq8noXStPAYexhSBU/jNC1uz8B8
mg3p9DZfuKEFQ+sSX10WsyyyYhGCzEfN1pUQv5irnU9KLNFMU2tPO6hCSOTiVJjNnFygwOp6Vl2l
tJNoxqgTgjyn4rnDq7bJu0YC4kmUdGboppAs+RZ8FvndmMX8D0ZpKldx4orWDw6zAAPKXOEYOXOY
ZdwXtu25TPcEJDWP4MuTMXXOEd19uw7+7fQogJp2QSaauoJQYfEC3ibirW8aeGBTip/53QfiV8Z4
8WJs6o2Z+MEUb1VvUn5CCPIlzRYwhcVx54m0H9045sUQA9d/+svD4lmoNpE0ot2IGoLkhM2eGPLy
Jk3W+mit5bXSDQp8Sb9FXws+avudiucpckfvhmAQGGQ90Qd7pIJPFEuZhVP7GHZD3kcEyekn8sV7
T696GQ5KY0oXbYo4lRpCjV+GoDowSqxAq5qz8sH/PE9YqtDsaPX19wP/leTlwQ/OGy/W1YWNl8fl
b2zbPIm/Ydjf5o82mtCVthKg36AcV8f6VgXr8PIvzPZ01+1DFeQSDI5ZwnkfXM0iWudS2UvPkw/r
1NtGxjgwgmklvqHZotrtj4XhJtqE1U07EpcPq/vIrEOc8Ewr1LCUUvJTsEO7n0mHi98VH7lsZc40
L/MBk46TPb1hpZf/0ZKr1zASWM3ledbqYDWT7Vr4mJGi0zlbZiQyaMswaivooM7o76JRX8fXeYZJ
6QI4GiQsblkiC17gZ2NBmaFQkvzgismRwdME4mjphkqWrLp/91rB74g+gHZZCGOvSclQQpAImwlr
N/m0xFxVipKbMfSr7/QQuoN2tCAKLqy2JoBAqACZrAdpfy/4G7wfuEeTSQbUM2UaTcczF0SA6Q/j
EXd2Jg8k0ZisbwOJgNW+p5QwrewmfuD8CwzJqE71adxgIG07NtBuS2ALPO+CG6qGZpLmwUnAr/Ql
+xzIdn15sojAD8LuMdJAVa0MXOWxhNwSTMzz0MlDGpXnPUh5WErfuoprEs8y5feSXFdBYY2v9Tcn
WCqsatxFI99wiXY3v7f/9bdCmvrQe1kDSBVF7y5+4CB+eyOI2F38c1DGz6lKS8wyOsM4o6YT/zp9
TEraxBwE0U99o/rr5CqO/1/GBsVwSw32409n1L74TlfJ5Fs1HFN9q1kL+brUfqsPllWZ1sdNkp4n
cSUqrKUo05kC7KVT5p3jKHMDkQNUMpimJljEgE8C468z1j32oGVlE1hzWCq1MCOJu09X1DD5IgHe
fhwRMNnXRx/mMbxltelV8U2lFq76rQauMV8UGpHLzBGDEDXATByE4eeat89yGlCmh/ciLA6qOXnA
ZZLneYvYwhel3Zc/Jn8wiB30YPwpOBfSHfTKtAbNIKlgG/fyoJlmo0XHefCPDLc5wUiMr+a9mHQh
1XVHXLLsZGRIz9lH9qxagNqfuXky1EcC2utwaxqPSyn75gdiSUtqQLv5tENShQ2UrVlVcXKAumRO
PPkHWGQl4QNOymJveJpQ8sZlTMAcuilpsvDU1q+/D/bOZoPjdziqKUSIcsYkNFEozF92aUG3yFWe
f5YdKMPkMas4iRbM+5ZyT4Vh0lLZ80y0TQ8q17ErcXjICyakRmVY2Vy8MtQi3ZGjlrXPev54BS5M
k7eyyuNPPUiy2zO1Qs40+TLcvyWdEUga1YfdfCKPzGHXZWRvIvIDhHsX8nUuJvvxvldqHDRtebmC
NX3sr+3K/uwZCiGKPWgytk4iy7LgY4hXGGCAkL5mXJNTVbkYfVm7ChoLMP9vEgex/kiSHsCDLNco
9RAxbQzcirs6t1AMWjCt5rOZLo9L9MoowIrzAjBOBK/MSWbksj5gJAfZtKWZlkslecdm7iY6u8td
rFHxSEsHfISTi1e5QnOYcvSTLXh1Z9xL65qE1MPmfA1/Ej7dCb8ntpLctBkvZy4HtrDhmEwe2k0c
ahImp6j5u35FJ1bWHliwN/glbxjL+mIkafN9DX6U0ayHqISUxMmP6yshexFS0G149mO15zTFpW8k
YeVj1wm2hBopI3qVnQO2ZBN27XH4bcu1IDH7cAMrGRBmNblU7xp+E0nCbDSANOaF1+d53zObwN/8
AJC/BXj5fo5tzrUbGzTmHylNWb4RYE6YJ9UTwqAdlfUygEtiy4BJg/5p8BpLenEVnJzZ6opoPCwY
HvaCYIrDF3f0SDq03k1s2bshB0vAxbbrwgMNRWKFCGdg4InGM3HePZ4glbtVtvWtMOI1dLhUV2CL
0skq60iOwKxQA226mjmCv5w9KVEYyqdtFj5i5Rbr34n1ULCoMJTpINTET+HIPE3iRIyiioeU7hsJ
R2OzOp5IrV0mXMAvJ5iAXuy+K4t7FzGmQgYC13V+tFDsTIJZPHYt56+IscJ+eTvDt1ALjcLpdQ8l
2x7BQNZ9H3yNcBIs5Y6QPBnXRO127kvW++2ivnjCBt1lWxVTqsuiLgxHFhHvRIlPuBw6Rq8mg7vq
Cz9C7RIpRS7KxnxzGnjncWpTtcFjAwUn9/NQZFdCaND8faOPZAC5bVfLJgfUusREWCTQAVlDy4H1
ir5cvVcpW/VIeorxWrIQl758kFkyapgHiRqc/hmuMXq8RhkDx1b7M2ih/5qcK/ZUy3imqG5zc9Dh
bSSfYJQk6G8goeMCeBiihDFWSa3qe/RGseakc3Ev9t1eDsMO9mTOPo4YdRjHMDdfhKaQU3cUFhAb
3TiAP/jz0JPzcmxkYCdvcbOVcKB+PXhEVk7DcoI+z745Zl2yiMN1Zpkuj+xlLFrFMhdqlPEWHzgs
fZTyoPQ2D0qdVyuclxoVTmHqZfLJCl2eIXCcl1oe9unWffoUBC03P2YKfIRxKWa0EXEpzuWKlWSe
EvlNlZpn8UunXFKWD+OhI26B2x/3Tpa+4dUwIGzEatNFxVst9rI3OZUK5VDyfu3iIt2SHSneLMBv
VU0AcMVrFDBJMRVbFkqfzxYnv5gJuNXX0s9FCechJGCSq1fa1sHkSyGUbSl+IVKob4wQsexicx5a
OxhLIehLRtbnOVtI0FyS7JHS7rNjSDMDxvZOpCWHjq/wpsNXpCZIDkgvJ2AsKRbUqlQDyQEm8aBz
TGm/GY/MKCp+jbIa2Px8/DLAM5oZag1B/yBc2mMvZzbaZzBo2j29JAasxE4r0mZhDA/qGiaZudSw
MwtA1h/qo7wqGLUQM1Xm7hLsXtfTgnFwISZEMos9t+aAm8qEfFm7Tjqn3fo65iGHzYsD85f3My/V
5QgPZsVawz4K4nanWiWOdM391Vzy09vsIfQmmf34p0eSkuet6rJy5f8otFqYEfzqoSkmVDmsReCV
bnYYjXqZbqrV1w4AdSYFMFI9RlbCon9B6k2HCwCjOKi2pMBqroGHCfv1RsOGbxHp23Fjzd+yf4ga
S7SGWoAjd08ziF/K92W12lUZGIwO3K+cBTJ9U9O82pBN1MVBYaN549vcJzsrgqwOoiczibUrPEdj
LXie1MdIU/WSKaAEapcWF72sggo4cnbGiuA0f8tKj+wMcAYRTOAyh4VRO7K1+aUOx+nid/t3cZBq
ppfzYtcYHRF/6bbcmj9r2mkA3/GujrZMsgWh01cglGcFE24M3ZQOrlEQgexrh3akYOtZZ+2ArJ6y
u7jtDEjRovC2qfYIBjfCyxAQx9kGVSQOapUrGjpIkf+1mcLsIVi7fjWF/6R9zpR23O6RM1WP2x7W
4j+OG2tVFuJngiTW6twpqa6IRZeWrDWFv+mMHs1n6Ww+ywcgSQObnsHvfUeuaujj8F2GwkEVTDtv
9Nx2z7eGKeXMKvP6qQjJU47XapiGmD9N17AVDb21gUNunbUGbtvQVZ2kqhzlM/UVHDU7Er1lM9n1
hYSJVNbIwvlJfmuz4PXtX7/pnCOKho7hV1ZG8I/d3gQsLyqW4v7eiC/hhBCHdY73iNm5sWk5NBfs
II89seqQZfqLpsGwacWch6xI4lcJgcVh+QQM5p/a4NmtB2Mm3RIhAZg0HX153q9HWk8Xc0Y82wB7
DNm9OSfYYSxoGQmthj4pSe0nr2hzf5QtRVXWY+ybs1CPyXoljxFQ14JCe2c0kowglu/dfgcH0bNH
4ZhOgBlrN59w5osPUo3gYG9Ex7zxGfYZIuSUH057cKqtJ+cO5Ajz9oSqaNpfeno/0qAcVfDFQALb
ophms5WoYtLvgKgq3ejO7v4F240nhOZtirT2wpf3C6eo2Er25XRmMfKcs/XEe5zSKOPctZqnkqdO
4zmH7n9BCsUAmpdUR/5ctBaPEe40YIlT1YUj7Hq+i+03pd5ta8gclZyW5pdWEuT8fMRpvwFxSnek
drmhnFF1Cv5OT7XvNolHiZJ23YEvqZJV+eFSYlljZd2uX5+5pILv/zOCAtssJ8bV3ApGos9pwaG0
T8sA+q5XIIPxcydnN07L8LIivnwKY3kGPGwaBbYR2C9jpBro55apha8C8XBmewDfydWq8oz8Y2EW
uC4u+kWaicJ9KUmRZ8mG1Zll+zWiXc7VHCndSkRYIdZgmLOpor0BAH2czyhRphxy07+33sdc4n+M
o29YLHjg9poFJURWOdKGIlnMTOBBl+vh+Oc/yJAqmn833xWinxf69NbdZwA4BU4BX9fED/ZJsley
OLUk9cO5DjE20QnaDg7CVrhD+k2pwU/H/BOU1Q8hFBMw3PRoCRJ5iT05NiwjfTDOJ2XNgRv+YEeN
rL3F7dhdN2Iv6Z2hVpbNPfLZDajQMb7noGrCL2rWwZc0xniOuIHAgQztNlw9MFcSh0pxYsZooH6t
UvXD03hjdsi4JhPEXWlqX8KPgnD/ElxwOjEs7rGm0Y0vw1X9jABy+/5pBf8lF1cq4jlRRTPcS6wA
6pHdkUnHqNhLcKwBnjxe7zSi99uqF4Pt1mG9gDSu76fJFKyd5yzk9vHSjKT0IcND7gdxRg+BcVTI
qJYRcvYr6Ya7o0ia3Y5jGJxpY6ICHM9VFPdV2U5nfUg5C8a53rrdYiZzI7E/dRKf7oIUhVdTk59j
NF7BM6yKpaQPWUyuG4L/rakNOfp6t1/mGEC4O0x/phM9K4DWf3kYxxP06cCAUDeAur5TVAGBGEOY
siTxgo7Z6BuGnfVZNiJcNOuJUhZbF9cQTnc0iL3D2jhxUBFeupO+qmrikjGSyTcwGcV0PcFR9tIg
pxAQhJzTV1cuAaEHg+YULZ0EfhLrPEIcI3XRlzINksf/TQ3oWImqnTvmkBHFtri7RXz3cnf6gH0/
NNbUBP/wL7sY/crSEnw/q52i+35moUbyD6I2cTyYJHkQxhbJXO3BE9xiF4WyYynHwBIUe0/TWBxf
UybMCMe7Rw3Y/82xw73b2etmp4v8xyzY5bgjFnAmzGQTCZ9WMTQzvl8vcyWfzRbO03U2OqkILYW3
3m1OpFTOsXSq+jF2TlwT1XQe/cnzA04+nS/e+GLRQm/wlQILcLZawoa2wsAOajwQd3gj7OfEhN7O
HHuyMV1AhV0y+Y3gKM4XfxNE36K8kT7eUrD9jc1dbX2lNsVh4sXneDXRjp9HES2VHy7BWdYNun1b
tQpRETXN92tV+EsLLvcpZahd2tdkI6BI+5H9849GAhIwCYrEKaKfpiRqNZgsYljEIwsB3KAyb81C
e2/T6mB12e8l2k/bOhJ2zm+fzi8Y5H+7GEYsp4mOj1asv/7sb0qc58ZSiQtjky5RsXkB+T2Wkuj2
910ZzuQq2Hz68qkH1Z6BhUdvDlfsdd6TDT2stpiYeBpNXPRAwJ8DLDrOeeb1wxH/bZbovRu5HvQW
CdivVAU9UnkedJ/hb2C8oe+tslrp1kGvq8HVTwnkN7Rn/uO9y29ihj5Ew4oHBrZaOrdyi/Wj2DRu
QNc7BBOaVez30m9Mchg9OIOGts6cVs6AnF7iiyUiQB6t0W9p1nLTDAMazgCeYNzcfhyg5KWAtkxA
i5b5zvkatI7R3Xp1sVGWpFq1zqrSyTPxLXYRlLe+5HMOe67fyxBv25bmkC7laAQSuGnnhj5MuSC5
TeWekkOHMWc+JygZaBjqhFk4/UrudHXjxIDGJYGuKVIJSRB3Zxmk9Eu/JXhYsSCPZnCUm0EJ9TXt
iPUE71xZq++b+qadx23lDljOwRO7q6LMqSaKIBxcqmoXbz6l7kczWu80pHCVar+tFhBzSf+Ty1vV
6osXc/ZjmstlCTwocDlTd5yXEnde/SPoWqoXNKt2GlrxC8P0mjPmyhlLB7tpT5MYzlLBI0WOvkuH
HTC4AceT3h0ePV+k90h7m8sJTe10oRgSPvwq9GEQtroPnXbg8bJQgH1xb5QpaxpaUzzESQxzWRkX
8ZnlSdwhcRnVfus8Dc6P0fq7AxqglgCAhKer9HQY4We0oU7p+e/wT2W7tRjseUmnuSg5BT7dltVW
/HKgfUYMmS/B9mu56O88BWqLPkJG/+V6xRr+whQK+2mczuzeQjlIIiqYUJApBH+OQPnnNBbmOB5Z
NhgkcKpN5MwpWIKLhIiGMLzkj13Y3Qf5ovRw0Rpyzc4BuW2jwp5/hq9YraIvt2xguYCVcVPVkw++
yGbzmHG3DzejH0Hm945z1Taxy3zUGI0UmST+ai/phlWVR4zX/fzgk0nO6tZOgTOHw+YhLqeFAik5
0xwoXr9ukq4BooudtoLob8oO8UJeyS6rxvXrttcdG3A7zw+x4HYhcG4qC9sOoEWKUyj7GJMORKxB
aoI1WsimejQHaO/C+wRG1X5TG0X29/Euo1yv3BKWEqqAEq2VTlQBaant3+GOoPLZg5IZpgme8e75
VXhAS+kL2bwqB8mIQQHmJMF6eEek37NiELo4I5/s/BQIG2WVFz/XvL92PV607+bFpWi2lNIxEqBm
EkmWEOA8jcmVeGao9AoRJ90NFwzPgWBbj41hEdgA0sMsqJWs6s+aHyAMkQE89MAqdkMtqMUBPP8A
iu11wPQQXFq6/ma2vclfJai75pBlXb1QgUfiwbR67EV8IvPx9iBH8fV0b/Fv9mAeT5wHiHIeXb99
FlCrqyfinqTXO2EaWwlsSdEf0NtfCLTXu6fFhJzi3Np1yGBappLjeWwCb0mkoEspA6uR6qe23uTi
Sk6UJOeejJTd46433rblwj0lswwRMkOVQHxEW3c7rCIIKfG2DVz79pWLApHNOjA/Fxn29ji1YwhR
I1lPODfF2hlyuozP8a+yrvwOzO2OKcj7M+OZuOnJxVFaenvdp30/HlSkYTOEhaXS8ftXUs1PV1W3
IATCp8q86jCHi8PqVRV4NW12JNIvGAFZUh08Yr06zkeTBoNoFbGbDlgNCIM5maFF9yWi6sgqVhnj
9peM4I0i2gn2ZKTdP9JEZwlDi205R+woFtxlqU05ALrSmWXEf8ysGDfx+7XLuVbM6fidoJfVvqjd
7Jt6jMoOxjwpAuR8fvsL8R6xIM3128tZJt4QuiZxEVUEv3oxH0WHm+T5mgywHk2syXlABsg0UiMP
ujU1JRkxA7BNjZD3wZ6R01uNeVE1tXn/GjLNzcmRvJ9yZCrfJqzzBTsYJdhS7Cwympugm0t4W7Cf
dTHUA4Oc3WzztemaE1NofcSUxFNH0Mc3mwFMBf7rYW6hWRbgBwSrIx+0qoJ+TyoeAycNyG15O+8d
uqeXoI6Eukd6pitJ4tIKsUKHOVtZWSCscr0Udh/20oO2U/HwTVVMPuX6mw2P2LJ4FcuZp/BYJA3N
JYKbDBTR/KLPoa7ecymZS9eZEYRzpAo4JSDmEQWGn8efYfeVyvvqWDWp9CL/kLg1MgHG4mSVXCiA
RrEobqpLjsY0Cnm93UaoHeMq4+z6D2qVbF8xidKtfnASyDUG97hVs+lQXLClFfqPjoc04NqDMNZD
xVQFSvO6PNLqCC7Ci5vp1Cdj/tZJ+lrz1mPz2SRKgyJO8W/8peTP0CqBBJWTlLGDvb3N58SpZznK
y1f3s4kav0ZzzI8QdB7Bp5GIxkGz+NrWAl6EgPqkT66lHKN7HYGk8qRe0pR+5XTtm33XHnNxQN5v
HcaSDkD3bO/modf52aZ5tLGb6M5yOeDd7bozq4RnEFIKC/uXGqkW6gT0sfrHJ0qOqB2LBEF7tkLu
zGeyQMmatsUoZNdUaOWx9NW5HxhcWft1zbJs/b0dApouoMT8PQop8QRGHZ6WcSvLpvAFfvaysDr1
oW8mbz5jFx1vkUklOlcXM1KO6WTUiJsD4v4WkQAr8rn7Q4gKPtk/TAHDijuVoMbSKw61km13wNLe
t67XJglwbWd9k6lltWsJoXPiivpb3qRTeLhBheYMkRH6jiVp02hPaid2uIoDn9lRdaSAeimCqoF9
Nv/Mf8j8NeJwu0CNIO3uohcDbnILdUDuW9C39KIhWbNOfs+Slp8TdrkCH5kTW3i5sKa3ZnedRBqo
dhpzz0QXA5t4mtm3SJDXq3i3e8pMIRZe9RB8fUkflV1c/amnX3UyRh4iSUeNwFFP4GEbjF5FkyWe
+AT/sugAItttnr1svcMAdjO4LOgxIDwgPad9zLHiLtmOtq+YVWfsQTi3iHbUR3gSzpMv+94b0g1j
FmkoeYIV983nksWtr1z7vTgBjljG5W5rILLah0jEIRgPLmLjlA2cO4QPwbMsH6PawVHDuOpPICc+
t8akpP12SveUjMsI9um/hGyD6aDeyVtsqsYRMyfZDrEaggxWTP4cXNCtdlN3RXC3pDcvKw8GrtK5
oaT8gNxHcXcPkdsjB/0+iVbmT22lbTt+kf+7ESoqtm3HlJ9jWzzwjly1w2+uLD4g889otskldi9g
QT7AKkockAU6ltpLFVhOUfPHd+exUy2V7cUE28AICrg08woarUyXE087YqKPxAoeJcxCqTK9yfHj
ZkMsFXxh05pi0InFe/rp55eb+dpb8bt31H2FjPJhcb+T+Sx+l4PST3hfCGJHXOqNlOV50fa7lJSB
9IMf4RHl4ZX0NJ5JnGAMPzdKXOX2sFqvtwj/cxSP2LfHXqYfzQdxUunG68V0/z/czYzNV1gpUWb7
bRCK0mDsMva8+ocAtmPM7ectsldR/WBXtVAlnDQ4K7hsZ1gtPG58/qUr44W2ggIXryhEXS7LfCsi
sB26YbtoXuiGIpd6eMfbMOfKjkWmKRVstfk4G56WduN8P7IxDkIZCdt8LHMD9012OYGbSyOwbluf
BPyn0aL04ViaklN3pC+QpQ/M/5q4kDiZxLXnCTl/Dvd+TLJG7WChAYd4xAy6BM8hEFlOIqUgwzdT
HxQz/KOI6lx+Sen/+nO0IWLzSbYAUXzEgqp1viQPpiquc7dsUL3GHlasTAUC7lI7uHS3TJ6by1OC
KE5F99u/MJjUHAdLh8lq5wqPLXlPXGG51qh2/rl43nb99GuEn2z0yyuTxGwLK6wdiuPo6xyklqpu
voe5hmuflugL09SxewjjNWP3Nd4jD99zbLlAbcL84Iu+zU3bubUNcP2kKf4X48rN7iSFl5rQB5ld
Fv1DtHsw6TVKOfS2i94UP/XpEKAxr//V77/8AOv/GUhUWGQG7iq7cKagYyZLEXMy7L2cLZQto2vf
qPFYM78LAPp1YsKqJFFbhNvIKNBocokkmif2O8V6H2raLTIZKYmXzr3lfQB4WQdgDuJMahI2o04f
tErTtt7LEbHmrV19Y0ZD4InmAKz5PTcFOptEOxnGYAOxArMwGmE4g41H5XAJHOkWop8krroNTofl
i2gajdxmdRUHtmJ3GydO5j94DBjtqUOaqETvt1dJHxe/fMlM7Cf5QtHAlCXQroMt2DQBgZjcNfVX
sltYTKKLmXEur2vDslToYoTSDJjVRMo+lemU0JZPErYmeBBYAfT3ozjMKAb8R6j26VjtqLfXnL0w
EU6HY4D33FvjB4cJFHdxI7dTEDNJZagMzdaes5cW8475EX7l4fN7mf5NnNHyy9P+xaJRMtsDksj0
zSWlKxxu4VNQfIoOPPr3LHpQAafWQXPyRjvfQWZcBE1AO1eAHApMjMjDA4yCGN4tvj2S4b70Hncd
WxnHEWGb2KTMcFpJFc15J+00YCWxL95Y8b6fWyjNFa6U68flPZcWp+U+hcn6MbS+/y3OJ/xB9IP4
+yyvf54kmipi0c6DoTZ97ZRkeOIyrtvaX2l9HL8d3Ozc84K18HBNXbDe9fIjF4vlA0hO3ivH8hbd
dvtG2BUiqnuJuqtfu3Y/2okh1mIc2jo9EFFyCj2GhvXIvQIOq1Qs+2u+kvQgTQGp1K6VvGhhxRz4
kg1jo5nsjPnbCGApOieszs0geIPsmugH8t8Kg6+mXrcmfOZvh6d0SOn7MeiXq9piTbtd+1AGro68
0X+TqxYw7osmXUII1yUCz8tmY3FERvYMxtfVrYewwwgnt33GvVwAPnjD5GycL8qx1rTkiR+OA2PA
sxfXeZCKfEtWZEajHwTLNYkD/se/NcOixX0KXA0YgEY+JlS+00MgGDKqgy/ZFnXOwifdtE548kSD
Kr2xRh2Tzhtu2Vr5yGzBAMtN5deUSb735Q/HL36J4GMZ6Xs+r1QGfFeMMKJO8mMsVhM1IBqyvQy/
JObCO0Q0MGZFthufftHmSp4uSClTzIlDgDHE/NCXVYV0BSng5PaJFWHvtwldOYtLtNbn4/thqSbU
blD4j2Ub7YASBZYnlBvjYYyrEKgLyWJZyGYdux0eHSlOmrdZoIe283LNfJIHc88XmA7rxMkZkXch
YnHXf6uvfbL4MDqQgPK5Nsek7cJeHJhvdzVakgRBPcvfCV/cfJRxXYpCL7MX+H4pDfF4Y8+BJsm6
XeSYbKHLtz0G/dxPCboJJ6IrM2MFZuIbFAInFu3p6//qsIFVQNOzEhKxKZ/Y8Swwm/DSRixYkBgY
vNYj6eqLPPC75r494iDQkN8uqz/iUuhHFglIJj9svpA6pV4sRhNr/Lylek5trJk7T8F6sq02/krq
MTF+4c+Jw6bJBbjJmJC/sgITreiGp4Qqc7QwGm0GxABummnk/a7CY2aaSz5tuz/B1oqzrWSNYGTu
5F77fs+zh31YR9YT6BA08vJ4OsiFFFQInICLlL6cPMoa498zOk2TBwuwNKxDTbgsKtI8WTMuFjXz
DXcf1YPrVad9iolVI9Fkrfu1ILR6+raEcLmfWfcLCqK9mS6/L/FKTudviQn07R+gm7rrSrye4H2Q
KduIopqcBfWuSguvVFP2xwz/rBbx29jm9P9EhtiLlYCHrqM6s49rJ/ExLOMSYTOXruoh6ozODLdf
+6u5OsmvE38oVRH8hWKFJ3OHN3euaMs08XSKtVcX54edecr2XYyCig1jg2vnbQl/V1sET0Z9hwu9
Jd5PGEp2gaB0w5Yc7xgPpuJXrD1G+Q/oIIHJVIYwcFmFGQtxzzLCRtF5q7YFJAyWnniB5W0XdDM2
RzMxE5G2KbieuKLw+1BA0vF+1TrGX0RXQlPxKz2+5rlsrOTvE0/JKhTNs7jhgX0iD6+I8NLasDWV
5GzmN6O+HOQVUTy5GtIqoutaB+si2x3MG+tj0bats0ZYLu7dmij07LOzmLgatrjZYEQ1IGMaLnCn
7q+VeYiP5y33UXdMXK5y7nR8B2zbsNZHjZFaBezUL+VIsmU6khcTh+a3W0+ZZ+91oiLXc01MzId0
YgVZGMuv08OhWR9sBb0faAUBTXAw5n2BWFEPofIcQ41Fpg7U3zDgMUnz2oRsQmIvPs9K2r2shL8J
dUH3mxhxIj+R3FRAl1aS6twbHz8vNQpRG+zdc67Hx5vFyLJCTZIaHmSb7P/5OWTPOYn/+A1W7w58
uVW/ja4hW1I2S4zaqexHa3bc9zbD8nO0I7AwYy1D2boRqyJkdJ2iAXFLX/ypGuAFKf84Wfzv65wh
4LvGIOplPWuaFv6R9hAnkvTQcjQ4/Cge8HV7ww5CEwM7XENhxUZEgkBgGyJ1DHfcvXUYTfIbKsSd
SJcgtAEjVIOOcCzPtmlhTLEeikEs6zbT/1CGFqq1lTtYBWbm2MqYXo0E3DEVg3ozAU9itlv+o2aC
ETEilhRqOmMSyOCJAwMgD9tAxoKJzHVAxIdJhtNJzfywAG8Mld/CZOntD+a2VBWn3Q3RTeKUiPn/
s9SF24i8DihuHiJ3JIaAEAb2X8r4HCx2X7VznUuT0zGQqpHZBBm6QlvDM4V+QhH+wqWu7jH5KjGK
bGVm9890VHSF4xtSOUOssDy8rOlgmtx3gIDNtxDuHf7vOZb39ywSL+56ZHMuti1GwMpfoWRxz968
XzTWi7n7sCCsi4CHXFoAD/5u5yYtr41EcvzNR65t0q+Xi1q1I6xqUs0y7155Ep8YcRxdZidst1yN
FihZPonp3iIYaE8MbaoCPsKWdyB3oQbUF4SZbLmx7G0S/tXyoTlPmLoX8Pm1gI1X4dtqoHaoIIOq
ZTjUvJu0DGJximwyVSRg5Sficy/vsdAvTHGVbadBX0Eujk/AHCyr6k84YFWdYbSzae3X0Kmd9hHi
fw8rQOeUXKW3vHTpXTZooZgfTYEt90N0F0Ud8wz8Kg5c+yVFgar9bpEHmf919+PnBOzX4fhwUT1S
UVXjIPKykqcS4LQmH+kcuO9ujLFRn/Sp9NBnFeCJ/7gH4Z/uOlZMUpf7P9/elWZ2Uq4pGppxPAhm
1fO+OZkdW+7agKnFkTTCII0AjzIuXeKNi4ws1tEUID36Vx956KgVeddx6CY8XLfiRqpNrgdTqt2v
gbzBr51Bd28l3QsbICrNobcFhkI6C28/VpmIvoYS3PVeQnbVrgBQrO6+envsj4yhoi6cwMgIq0dM
gPD7EeZV2ad8t3J9nLbP3Mblg3V4e5Ts9VhfE6SZjV93thwvi5ON7vTDhFO10aKd8xVnh2qRAHqv
dR8QEkUQKfClAXniiz6D4ctb/2U/byquuD2Wo9VkxB3UzFzaPKKr6fhSLzkOlqK9D0N4wRnxz7BS
kZMJhnqNSgwPc8dhtqnHVos7iR36ZXrinJ9KpqNONY0Ndm3MzJB57aTTUFnKoQoHF+n1mqDO2zjs
hxkKx80U323EY0mE04jphtRvER1OfAw8AqGPol1UYdoKL8Q+MzAkLSaUdZYYSWUhl42MndwdCUob
+AHy8VbT/fsB68NytC0y0yH+2x29LDp3zn26GAIa87x/lbku7Jkss8LaZuYpSX/xHzFaDbIBBUdu
yLIayk3WJSj29ZiXv1l9+k8ZwcmZoLq32ZHA9d5rEKt9TOgoiqdYQSjLKCrzNOuOi7dtPWtwDIpm
5lHmtfHAWE96enOcm1BBGQ6k3bwE8GZkr9y9rAdHCRXogwIuuRPm30Gdf3ksUlZBjr09ReZ+1N2Z
3gUaEgs4UA9lOz2gsbqsSLDrUzEapN5Xc9CQTo8IE2ByTj3HucAylk4cnHuqlK43xfYK7pstR1Qz
VHcJX9A7x+bYPUWHUL8fkpD2Cn35SRlErDvua0I772iJajXWX+m3gpXE78LR0RNxcMRTtTl7Qlnx
kAeD12JrDn98XWUumcSxYSFFOmKpeFimmklv24HHRcqXyxzEzjHDHDlC4JaXtC/zFIWi16CN0xIS
F90SccpYwmrxO7bkUJgBraMIBJDJihwKy1t+oKcACLTeeEfP1ZlvHCEjP8t0SPOUeQ7S7FXTI3K0
A7/LUQOQaTtVlJM2sGpbXfNUL59DeXjqfNVa2+zA+VJJJF6Iy9xS420QNc9+5lmFZFdMSB+/yruf
t36H43XzEczI1lGcBggc/cz1sS6fzn+IFT4xEcKK/9i3w8X6RC0BrQR3U+7+1RU0Bjuo7FqiIkqw
ok4Nv+3PxQfZdfdoUK/jpll9r8ioAxsMrtKRKhlkzeXzRLfo4y3K2n29n0404aoiPqjJbrG3AWtR
ufMHXv7Vyel4TfF3ZA9C+RggmdV88eZdgyXv+cTBwNQB2d1AIay0C0NQ9n2UO9CsBz4azxB4LMqt
S95sa77QLQ3AdH8J6fpurvhFLzrk2yJqdeNYCkOowXbjUPpyVGvZUkEYVFuxnEIzDz+w7ybgjje+
r7SXXNUmemMW8ko/lNfN/JbQd874vqVAbuoqCzhAdxr9xyzbW1uP7A6biyHf3Q0F5ZgAt78Pok2z
BEYeAQpl3IMy9Jt2EReww6gY2mZ9U+C03HBwrr6msKhdPLVd1vnzxjZnAJ1Wtg6mFLNtzKz3bj0j
V0FDdEYI7CDAiElIBdX2FxlL8vZmQt0ivg7g3K81/iPt64OJdxgkZSJlj+SY8rR+J6ETer09Mzci
M6fiOCDbuRZqX3bZt3NXXfLDWSlaUFCXEfnqYxikPA/ECCD/jgj0h+Y04+WBvfuseD/MELZO148R
TA/UzUSsJujKNXxrUROLJwtN0zE5UV3gGzwag1iOzYYoAH9AvchrXOTZ8eHm7hEt8PYiHKajFGMe
S6RLU5nsDf3yo/XgLq9yy9TjIpcWnLwTqkwY8rzssqYIi4dvY1nZMyqM94a9wZkB0hw/WG6rscAV
N18df4BOuVqG20cHsNQHoamuvUnETVzqu8pmmJAPzeAxlp7K67FHRu0u+Fe2ZkJqTZcHTVDsVrER
TL+SHj0P63fH0a3Lin0zhXlqyDIZA9TpIECK9Vk/xL7SuiI3U5Mb7cmKS1t2hN8Cb8t8PNw0dBNb
HY80g1eqgBpqQOJUufVbS5H2g9UUa6uFQ4PN7X9lzsMlaEOitP29SU/5WIEl1xD3ZySTCxlAl/E3
+GZsCLOvXDBj5QXiGT5Zy5y+EnYtF0JH7pcvU6fur9ZmiBOCYD+/zZRSmQyweUvdt2n3BWgcgpol
AhwgHY1ERVtUMJiUTEFXz9QCgtIbf9FL3KsMKSKNGJufWChnelDZ2T+YiLUr1YP0wz7Q2QO6b4zD
ak2MQnRDwwqS+SmskbyJWyU/Xxs48YWlz3AzCEZdoc6z4+ZWRi50DGkOJnNf4pobUmvDM/21zuHQ
4Nq9RqHMBoXVQ2+I0CWSiF0YANs5jOFLYZVjh6xKgE6ITjxq6a9fkFO/FcfSNhV5Dxx89+/geljm
6zNUNOtZoQs5IbKGciy/wwZNb8lngN1tR/xZNDmgKa0P1I9C6SWTLM8t5l4OHI6FeXYY5eG0IJVS
EbYRVu8IhgRJXWm9qWlWgkTvXkoBy6FA3vADtM3ztWZVw/OsFb4ODWR8nIS2FuzyaucgJHH/bYD2
ZWzbMli+YXX7mcYQBu5bVz1lb0axoNkRGJDwIuXWaKGa9+5qgnnoHC/60bQ0HnSwqV7MgfcbisWL
YEome6LkhNXc9K1WuIp0ktj6xDA9CQJadJiRbLXanX3CkFgHXI9Sc/9G6jIWxaER12AbkhNigYeH
i9uOcU9/qvUhsKhl8fK8dBhGcStnw8M/8lBlMbdH4Bp5Lv+WXkrSaGWf/FdcJNpi2g2I64r16Mxd
patUT3OJfYlRdJZF7tWz+FJPhdgUwn6mfv+TKZDwK7fx+QSV3r7Zpggd9VW06EEP6491UuJcoA+F
2uVbtz+OZ8LEqJJ9LmkHITjux9BoN2iLqbjvVoM+9vaRkpbDXz6hltdgNXI6Hk42YmGkgkw6/aLW
yDOO6Jm4mNnAMDa8Kmsz2+rGyPer7VXY+tHo6t1hRzxxqbO14yX+ZMfuXXWvQyvwdsnbbO3hMiC2
Y8jlsMRhHtxf9c4FFc/833kuTJJJPzwSCGKEgzsjEjgkf5VtjCMMRMk9Bc/BsadCeI5h3Tw2mUL7
02REZZ5P/701TFbo3Q2VZ8F6ZBn4k1fTKIYKQBDn0YyIGeMXy7sa4TIRw8WIinwr6JFzp+TGug03
CvQvTkZI36Gl/DCTp9D1xCBgt4SP09X+H25Il0rNVA9JmpFopZpwraxI2N61cgHmhKOEvzBl93FF
4VCZE1EPEWhHaQbR/q6UytW/T7dpWzLMYnc7az0jE3Kgm+nU1cidEStc3+JBJwgx+5ODQZ0COqDd
iabbDxhbNP+OiZT+4GyWFbUAahRkV58laYPw95VuvVWcwmZ1oZjN5CH850GUPMqP+9q3l4r9KXZO
qQAC44ud/hJ0UKhMOd2iHKUt33l7/0aIRn9J21FoeGGCsh9K7jqY4xm2enstnIompg5ZU6FoRo3g
9J7DLrO71hCwfgb+ikd8IqTMHxBdKPfmolI+Nq2UFAazKCRVIt8yrVwwGNHzEWeKLuVLp5ZuD+Qh
XDuwVxbrbNUIO0mRIKcq68ki/Cg7vqijCq+ZfNQIOncb4d8G+LFniAmt2SfaLXyM1Ww9fL4ae8yM
TPGmLCzuwKnw3/ZlbgSU+LHpCwgplUEGM6dM8tMfBQTjdPTRoed992YxYRtgI/QOsMZ9CbNGjUEf
qzxGvJO16iy3QjtCZNw4FfuR0P8XZKRTVHWOEy04lZfew+OReI+hFtM4Nr/MOSfl28IunkFmswXu
0zhNKQBfHrf4E6qHyK2BIROCtq72hR5GwmT1sy0dm309oiIitUY95NOKijx3XLfjUpRgTKWTvmvv
mbgX/DFnmm0N+iqCe/l/gXe6FOSdfm7VVnjYVytex4CjS8Vh+OSSUSuhBZ/R1fgXQgyY0vc1lquf
uREjE3Qyuavbe4rrFb3StLg/Q5SU/MFj8s5E/vcDDrleSDSOHnhq2/qPIY8Jywa80NKrLPan3pcy
06F8QHKzPpTRGP9+6BdWvFxSrIfvCu8vrRvAdHLlz0GPLSk28G3e/c1R62EiptSMyJIMXW6Vol/z
9LdIsJHjYr0RQ4NKampRQvTkomcYk8vYmhiqaYeaWsEdlOoES40GvTDQR2Bzff6OF/dMAkgqaVNv
RT8FzcZiporrO1WBAiglH5mWqhgnI1qPHYj9PskUAGTpdKpOxl+SgFJjwiTy34VNsNd1g3OXaK8Z
dL61GTnvejbd7vy7aqnrTg9e3eMJXGpjQ8aA8RVFqnVjrce3KFiwC5L8HprEG/+Tnv+4+4pNlAQf
RT+xi+UHVhVrhMYuXt0otOB8hcgLx7shILXOhsQhGwJjRGsZXvg3HYx57hS0PYoRqhiAk00emm4W
Y3dUoCpfM06OX+sq6x6RSsG8fE6BCW4DHL+g0EF/u3KIUjVCnxVWMzdVj28XvyYOxLs6OWtuvfe/
jY55cUFXxFxmqQCoWYxQ96h5LILcgFct47V5le1XIGfvF6YtlfEngYZmq04a/2G9e8HSEfh6jLhy
OQcev0klBnxn2xL4Y6BRYiyMgxtMXcYO3vuvsq/ntRIrJQdvZrQahcnYDyVHT33hIIxZ3WvJaKoV
fYmvLVlTyK0g2pqF50Gz64nHwkSwQlaGqQE9GCLPRhevLZ5HT8j4lc229qlJOw+udl8i+T5B4dci
eXpPvfPLfddegg68EZYgNB7vC/36pArn+rgPipYaDoAE5mAdMOE8SBdmVVeOtLlxiw2b7tanuUin
D504mdENFbM2gWSYJw69KwBuulDXYAy8Tm77rytVBratALvX1D8BVMAZc00vynZY68FJic3ZI+OD
7erMhH6TSc4OWCKTnhc5n7NSanXv5Uop9CUTUFF2tgLuzQmz86KiyBOKaRRpoA+4OmQNcG1z4tWc
CgUI63FfCNBSsBM2p+QTdrAJONtjNLfwQj8WGo7u/LzQCKhLcr4+gM21D+NbkNQdTda3IYCOM8Xi
PTO96euX56GSYmeh1qjuLqQSOV8jcXmzYCMk+riQ2+HVZbLBXJngbk39sGALfZw/FIa5z5rMgUcN
EWXC0L3V+vQPOkr7I/7gNwFUrEZuu2fezkcBkpfb9Gda3o7H9aQLmM7+T2Z5lEveJKUmM5QJnJRi
2vDcyVEtTP3KD+UPMsUnhA+VVwq9yC0UcgRvv10GVdB46IYjOa5OJZOVmOL/zyuyNN/M24KN2ae9
ivdaqloaNFvwj2ekNXQ8hQRUigxAIaS+oCdH4nHcx2F02L5DfVyOx/QF+m/7QnFU6Ti4ZUySSy7D
+W5YEiaBeGOfExmLV88xLEk5R5O0sLK2OuOrQwdUOER9I8qwbaT9q+xjql5Deph4lmgMmvapVF0U
G95pk1ls/l9Tt7WrHTc4kYUYAThkgrmXE8pFASTsHPhOPA4PVabKprImiQ4rLSJPxQDoWRZF6d7c
z4pu9ekPX2yfELV1eP1GLqj9AIOCujGOiP2AsYp2nvR9hXq+GJGFyLzvivQOkX3EHKuk/rHJZ0pa
ITKB07K9xK0ydiAnTn7dTt9ycu4vwhjSoYYIJc24uqY1rOs3SlOG/YRBbF1C4g4YQuMZpb1p+Zvc
NuCVBqajn8cPrwiyjkqiHZ6gN42GRLRixhp09FVVL0q4Uh6SSjXZYFKbtsShlsLHJsM2H3t4lSR0
EjcHDOfCVCEW1U9AJJML+NJIqGjcJ/onCWQowpM59BCJfu3+BEABx0ukB/eZvgNAEJnOH4ga+1F5
c/tgj6lKAVTLiH0f/1YnDoE2mntqVmtgCGmv0WIFyj1ky0jycM5iHpJUC6qdn1qWM8ceMfN85Yfq
T/f8dVqglZReQC1JppeGILUL2u0qj17xh6xxCW1dJOGKwcw0TKFkHg0q9TNBpVzDyWOFCrjc/QqT
MR3G0Ep2csCcQED0/9u6Lls0Xv932e3kWwkYnoiiEEUpFf5S9H6lfm48Xmwny5HxvEcs4y4pY598
oAmvrvJ5XaiW1S02g+iE5eG3F4y+e5D11bTaO3tRFk621Ok8uthbWR/C6ju1rrgV+mwhWT9n0x7Q
FXcEmKlGABot+oip4TExQpT/SOzWbEkjX8PUVK0V9/NsKskVA82x4wPYKFnEjk5Sq6i5Yezjijo5
4UA846tVZzeZFvnT2HbXp9CRbAA1q9k0WTlhZANvErwTMzAeNpWwAJxDSlTVjLFBxk+8/dC9hjId
yNFGgtHMcOnEDNSW6d6TUgqR01QAcIsVDr9awcPwEuSTtqrUqO63+nx1X/3JyKJIqaISDNc/Zwqx
Y6rhlEVQpmpwy7rUjLMs9OEzNhkAgxGV3xt/wp7sILPBfV9VwtXFe7skts6fH/uHYRzWQziQxNv1
XkNM32FN5ULdjm5WcfS8OadaMyR61uDdqA5kYOWFNiYa+kooyCcFTrWhoS0Remc3Hhl0hxJRkOgh
E3fTT9TEQoxyMYe21gXOWsnMYxunQcagloEES+6h4MrLWNFJVRnbOcSyya8bNM87FwRQkUPWAT86
6h3yKgyn7CHBoI7gy0KGQM2qW96kA967mFSXgWtmM5MVfvun9RMoi0Io0w/AKnEibb1aenPq4L1K
vleLjYP85l3X0VnG0xsGO4OOt4ajMp1hVwRT/MojJwIyCiwAo4fmEj5LLxjFyzOVkh+hzTXiUCkj
KFYnZOYuDEAMvqEzBWrzf5Ofmpbcxr+v+mAHvdZ6O0ojAqWQwEXWEH/3KMHyA9QS84ATzPHoOVXf
qbbWUbgwPUXUBBP6inFdMZF4r1FaqUuyIXv3pK51icmcEPKL+jHRaEXiCtZmbqo/LHhCMqTvLYCh
EyzGIw+Tgq5mO2KAdAyIGUSvfUtsqHYcjJ4yn+LptxoQDv9hHhhIUq8Z6osOkSqD5DvvMNprXSRI
baGrsmE+7Vb2qrXVP9JPaLcFghs+lWShi0kuGipm4JBOndIv1+zHp3lj5Eh/LS2PBUAPTeX4mISx
yn7CTPGvhOIm/WFWbWhb2HAu38u4WhujEhegMIBhN5JwGQ+yx94l8wsxBrPmYf2NFm8E0Deif7EL
EqVbANtuEM1ol4hKpRxIPXd2AmOCFhUClaiGrlDk2Rt9nShBwP9tNBYOsaDtnNovl0KnHApSWrsi
4jYZxA+xJxnLNXgsLknaDqFb5FlsxMSx9y65GauoyVk/ohtTkRMFDHBYtSiWnJgo0eya+hEFFCqT
hK0d4oUn7MErBqfAiElKTvGaPXyxxZbDljGIifQEkGOwCYdMGaS6EnIMQnbqy1yhEVOVUmkPBttM
XqJZR4uno0O+TLPI+yOUC6uOHrTiIkAp6ZdS6YV0EyQrK3AmFom+9qV7L6kF8sjCpx7fPHFhagYR
R6o2taieYBybKFKbTo6NVtIwhMIOjpy/zoP7uCmvrVtG0bJEf9NIELJ+eIOkWJdzYn8X4ZU3hb+d
iD49CfP2HAUc2+LThQOOFJFhX22ff+DB69vycEa/zG6ZiiV95AjqFLK5WEehPmyxRKFFYFOEIswf
Cdq9kkNjKPfqsl0olXvUtmmGhL9lMW2s/1ayax1acYBTlyhHecof2QtztYwq7cI3qtPKWi6aLf68
JWbbA0NBkyogCPO0rqwD7u4tzDtsVyYz+N7s/8OTTFrX+BsNlDwCYO6OxVqPrsKm7XZUcBMUJHHm
QPveHR3M8y7eIL5rmFvlsqPwre+c9LYoO+m9aHy1aeDsRIqlfzNxUF4GVudkmx/SXcZQJ1ol1NZU
Q08imgYJl+YpaMEEZQe7PWtsc2HNwa+HowgOF/ovBT8XKQ5M0uvKABIxLym1XvK2d4IYf+GJAd4L
l+V84W9d+6gwZeIaEUPIgVpXO43RRYvYKMYeBvKLo9nW4VZsi1Lk0g9OXPC68Xb1EqIwpld+oiYX
4klgBk0Qq2sEgofhyNFkNWcq8uoheqJC5LwrLEnLHrnePZIUw9HTHOXd3qQcMDyNXoHk3EBA9dFA
kvjyowJcrtfTX4hHqBj8CnVLj02iDkPprRNnWv4074BKoTXPVGVZ5xnMw4kES+nK/7GiN9UY47Oz
Vo3JuevN67Y+gVISVRwbfWUMnw4fSakKRxySE6UqP4+BQT8WDs2NBFOLcUbdFxzNCNYELYN+CPNM
2GG2j8+65pP+1NXlgjMFb/HzjyYqNUI/IM0rygS8wKDjiK/+ZjYIIYPhRkXuhkFScQeYJm/esSSW
N2ukoXMf2jGL+b3acFPA58WyW7RMOL7n/YpV1DXW+kjxGl1uMqJjlGJ/TpOH1fy3tWelnpav6PZL
ONO74fCDzWBbqxKxzeVrcN3swJ38Vuh4FEeXPqkr8k7ixaNNfmBpQD1B8xaHFwRfWXhnCM3gwOby
WoBO1iS1pqk1zyqQpAQSSGgoF2+lsQflD8ufdMEumY53sRsUgedO0bBdCgNvR2hDs+jBWy5ihkng
mMRVENPxzRdFT5zCNlh5eapPRoXTyyxIDin2p5PyqEHZAzPAFr0ysNzaZz001Dd0fJcuPbL6r9mb
4zfqdI/NcdqhNMEtF1pbcPXTvce8NClahR775pGAtI4/CCyG4KrxBx4PGM9vujc3vSCtB3Cnky0F
PkDAlwZN3jNsHM3byteOscgYW4JXQsYcV998daOzkAvZRNhfjBn8D83UzwC2c1cNS2l4K8qNwx8u
JpV4H4vjZ4mLB1KV2xlXz/oYao3sX4vurygy3hb5bR1xeIZKKK6ZFrnYg/ErzUC0ezhbcuA1lYF6
bll2eYhZqGJgcuGLQszYQQ0P9TLyZOItVsHINEioDYuwp2NwaQhoVfwoF5VUya/kikn76AqRUjRj
SDN9q+KxsuMtRDI1wHZt4rqFBTpXkZv2pQYWukLy/1hfh1sEKzvPYFbAihWOTibM1Pzq2mnrlX4l
ZaN2crBt5G/CF6zdYIRCgQHZxh5WBIJFsL0WKJ/jsaOklj9r+sTSFHXAs2a1BfxQvKmgmU5dF5cH
X5576gnSX7a+P+MXLOn/OvQcVZ5r36QaveWXGwv8C/Id+Nj/mvssJWp6+fvRUm5hLR17eqB0K9jT
Ww802QruKKrdfPyoOFCs/Z+Wj69pAD4tY4skt0KIhv8sdFVPgRWCXy3Z4cO4TWvPz6jgG79NUJJa
K7teBcpFHhs1a7wo0dVAjrdzD8FwU5e+ewnkXMaQDQHPVjcSu7GThDLJqxHAsNILFWZx7MOR8YP/
shdMV5kltDJo6OeMgHVYa59whsjoNJ/K9X7dyR2JcgHK01lkgYKpOLCs4RGWIs1ysaUdvx19Z9W2
BSmz1BFoXy/ifZUSojK7dcrdm2qms0tEQr/3eXEpAWdzKL+jy4wMJGJpjojZF5gUmUEqI8/eIdBj
J5O2PtNbrEZU6Rbs3hnIzCTp4v+sozpWXqbULcM0drmRoLKYRr5px5eb7l8n2mjdfo2PzHU9uIWp
eF6fIl7TgGmSV9/CjiCWl25F3Yw+SpzhOWRPLX8AqWVh/oRNDnm72w8S1Wj2ixdoPwQUgh8v//ls
PqMxB0G+GexigQ2KSBvmyLd4SMfTQlhbZZdtXEgJTfQBGCZpiXNFDUskJd+N3qSkcI6K2kCGSW3D
DCZ7m2TIzIWTtMjNLlfyvFiHfUwYYPshv6S9ZGUTKd3QNuHr/J/EupQSInbCQB21M51BOlyf1ZBm
eu/hRndmlyALCpNUFne+N82+9DDxzETwB3L42o6xuAj7AtgEkiNKeodp2iC3zhyrNWveA7guiLjJ
dXw1avFRpc/K8O31fDaZjQN4ofmkUaWEd2tLuC5LHCSMkaGdjohvHF5OjXKuHZ/fEvTGX5bVDM3h
cXIknSyY/skCOQfyEJ0I17n3qGYHCpIL81YaEdWA9LinS2YvGo1fbFwWeRIa3DBCKk6I5sPp/oEX
RVC2dBNDlrlQ78q+xDWc64v1F+k17LKTy+8NFOaGWUBbe6yAY1BvO2PYlA7c6WdqklIYi3nyfL9d
Gj9XKuN53E2eRZM8TLM8sqMOi3sXgEcCKX8U3Yr+SoDh0O73znEjR82uTQwTiJtjoc1y5dQXAudX
YeAQgmOuRBd6wqJih/2PJJ8A7Ou/6JDWglVSmbKfw/dkUyRs32EPrhdWfQTGi4Blt+aoNKc1EdrU
Ci8s866hFnW6D2cJ69peCz3lO5OAP1B8cusuS4AwJPb+o1Rj4Vm+Zka7O37rJ5YrguA63j1W7YHE
pLPPVoizp2U1MSowp/zNhBDbzlZ7wgngNFrK1uhIGTdEz7oXfKywipbPcvqC2aP3/QVYaKPnjJrR
9ktjsM0TR62yjVrj1KMpjRyzIgLO7OhX9f+933eP/pGDhPRlbvmjFPhLiQ379e9/azMb92mhJtZ6
ivzzmKvbaCOgJFcsNOA/E9dlUooWxz7BiKGItrLj5g2ssLt11jEHAdfnOGGVTT5nWcivwitqJ+DL
jfN3EuRCkWilmrbmWdCYaqKlZttk2j13Y9mR2saveHpJMqtSwjkHIoNNW+z7ZJB3B7McqoOeSFng
HN+1s/fBkgjB41FYcCRWhbGd21UIClpRTbpFsyt2ynMPS3+IbzSlVC4uwuGX02sOZAC4T2y+Td7f
I7THXUh61S/cQx+khR8CXV6UFtQ4t4paagLd/MpxKPyqkplh7Ekz+HVF9jZZHSinQxf/FG/4OcI2
iBWFQ1WIurGKjXG0as97i8GUmY3Z72Q9owWLLXVZ6pu8AoyVWgUXJ9+UAZC7fCLuxN4dterojwlr
l9WTGm6enHb/k0EglF9UAGu1wb6g+X9qsvXva+InhbAHzemFQTokaK4IKoMYBKDr80K9LCH34hoq
QpPPk6kW154h6phIguId/NRxiPPjEFAvA6f+gbJeBLEgDlldH0iUPwYbjSvy4OuCwTCcH7ugH6T/
QM+nJURQ5eSr97f0+uNXWwvAE+EcAv1PmD2DYj3GH5QKI/piqJ0sQ+bsRksMssjBzAnv54VR5ini
SMCqqBkJm6jFbl0znzEPB6hpqhJQKLN84Vq0PmfcwoF9OnUH8/mgGpX2IWWAYXDO0cjmmaqcMfFK
2KVeRc6O1BgKsC0XdaLu+CZadpTrbHY9WWZWa5EfwEdQeLGsq92wWNR9aiojhFsjvWbgOke3skN7
FR0dFcHkqrpFUGVGA7QyvTKW6vXcDoKlEeuixhsq/EHB+CFhvHBvL5vvTsZTfdxS0M/nUvB9n9XT
59RKsn2Rrf2AQ7aXS2kFZjltwqunDjVLD67K6Z58A3uH8BHl8dIkMTyWUYAxjKavC6XgwcR7FOoe
K0tVF6zBgmvWr5E5hxbKhAr5K5fvjTzL8D8AEQgB+vLCdUbxGNVBI5FqiISiVq9gP8FGhl7sQh22
ZfpxUKaG0Ce4KzDJDDLVQ8vHF8cpxsSJoRL1Xmd6GxRQeyiNhyurdqVD6nMrDE56Wp42MlmpSEgI
3BGGt0h3lOz7YBEfIJcabkJ8aW9KHB9sQRFpD5Ift8WBnzZkvNM0b5FFCCsOQKxBz5UQs6lgasNQ
Z7CI1LuIWJY0gRspF3Q2Mm3crBeRxBWebgts6V8+y1dtAFyfedIcKkuVwoWuze8zFX1n5/oVPQku
ba0dl5FxNMgX2KspouUaXXgXkOUhwPkCdVBi5RwXsOuEYyLZ0r9qrRwH5gPEashgES7C0NEo/MP/
6VCHGgNmhKtJQQ+Bcevpuyidf2K/f8/ZAX5y57EGIJV/gIqoI0A9YrHaT47P2ePsKUn2Hq25BGqV
4uVllYUAVU92MUpb19d7sNpsuRdySyVcpVvy2/G6rmJ1ElPh5mdyruWdYPn4OVwoPMFBlZduGBzp
C5uIBRS373P68EMfW8z72izUH2k1vVvJb4o2ZwusLqp6FO33ugHhGYzmQnF21JoBvm3/IxGc23r4
k1Td/p5ng8D/jcW5Z0xCj0oP8ti+A+Nirl/Wr0XOmmY6EejmwyGnCqfVMKUm3K0C1bcV61uQmVuS
GPdelbGLqc5VB5L/GTPcKg1LheAdazgU8Kkb88AcZ0hXoS9JKKv3a7y8Rtlt2mjrC5x5+5NwwDoP
yW0z/ofMiSLKHDtq5PiDWetJLCQDcpZmuQcDdfbOG6qN36gfitsa4SaAHa2mv+Nj79sKW1aajk4T
X0nPklz/wqdhEcXGotpQO7fAvktuHNfkx8IgXTyCmiPixHh5V4c2VS+IhbG0fwtdNfhTVAfSR1qq
PYIHa2LsrxdP5e13hqNVxdvDH8lr3UJiiqC1i1oiLghua44FakJWKfP+fnHiX220IPDjF3XxE8nv
0HhzbFFgxhwkhIEgsJCfbky+XbP18WNKAl27Vx2dDMvhGyBzD7YYeSPIyTRjYGt82cIW6h7oq7tE
d9MqpLdov7zKBPUmKyB7pxIhP1TtyorEy7umczpxoloUA2lzR5pXTxijZIEvd34Kj/dVjdJqNT6t
NdfwJy8xpAwyO+/jMwmvHNNTgyUe3JfnYcaGQ+gdk9Y67UuPiKuyjZoNa5opPS4nOlW+0T0ZRLNB
7kvOpOLKyJ89u0ozKffOzz7xLVH7SK6xRZeCCUEl2AQfnzThqW9RpFcrAFyH/Gc5GmZ76cG2MFd0
Ca74mvudMxlIN4OFVnF+OIsEFIBuFKe4XHtljKyp/tSaZ5jWyAnnozu7ntPNJIYUnEwrjbWwWRt8
aOquCnZ9vTx2dhcBJSA58jkwz9Yzyw1U+9VvJSAxidn+ltNDSq+5npEZqzdp6pIrksABXquSbFUL
7mI2mHr4uoWLs6N7a2YKQEMpqf53OdbmfRXO7Fmoh8HNsOzgcr4AlR61tkw1DTnsnuimSmMbNxrV
/1VQP2i8qUd+L+CMiUIch8H6fa7AoSRjHsNBvbbNx9UwDy7TTe2N0JPK2p7RLqvlq2BNq1zBsqbA
20NyF2MzFUdRdZSBZWi2GJABMD19JbJ66Pgsrim78U38AFMTumHxCAEWHM5g6H/Xr/wuxjemmuFJ
yuCSatkquRGHpwyCJa1mvAwQ7VJsjY0/VTHJ+GRbU3k6L6L8tsXe2J/T44Sr6rMvAebiJp5vqf/8
gQcmwVZ9QI4RsmnnBel47RGRBcauDBYxcneSbsaoLOvHJzePQmbAmA6uTMzPvXoM7s8pwcQ7wlNP
BXU3eYda9iaqbUDfuKwgKKR+CDMxcm7m4ej1C31YYuWuJu0Bq3THeDRWc/uITkQORlxV9TxdYQtG
z3fA5ifUFptYQWgMjKRqmCwlNOHLJAF+LZvKiRrFoF4HdXdBFo6k8pRMQ71RBCDz9IijW83JT74G
I6u1lYZBWxmxfIPXsuYNMfDveuHxcOaCVwdycjY/SQrJSgyjen6gFLns02g+TuucQaL7Ocsj6TFZ
YVu65krw1tPX9/R4CfrpFhPPhmEruAgw7Vw49Ah0I4XGiIPfOpfqBtc0y9YWYBpop3urAWjM2Otb
X7Vo/K5/WguhTSsCMHKALHSOQtXpodKwcE21fdwEfharUDZV3nMypxP4LSlxJeV4PhHMKxQNT8UL
LBJGJMGb6VeCKsEEyj5Gpl0ksaiwHJ62hmg25NYs0QRZBbALkSHBS4IJIEpiXgaxxPEg+BYae4xX
RDDTc9s+R++tikvziEcriu+yL8gGsa75iC5NVF/0uasQduVU9RAm7XmdzBWMqt58T3onsAgNTJb1
j1iDZKYcgasbTFR0qqjtyMHbqhIz5snU2h/RXxhlTJEVRf/2W6CAPKUduRucogxFTb6yYqfZwGTJ
rkrZ5ybNcG7h93mC3rl5puIoHKC+4+u3cdEtw6SMaIjm3YKyTaRVBtFStoU+VHUcTvvQq2307ayv
CwxvOCURX5rlQdkmCPdmya64oHEHZxhnfxs2odGfCwrSPKCrReTyRJINOUAmb2ZyEnbZLHP6BAS4
Z5vi0h1k6egdx1oqHPs7cPEEw7VlOUmwEMfa3EPryu4mZR20EIPx5gth9k/V0PaW6kYfBjuZcMt8
DNoJxOha4PVF6YaSOYgui0wGlcXkQlhbjwAvOd2l/pz8xS3ebzVjbQ3HjdLITPRWifn6YP8vVq/A
RXRlTPzK6nT0yCeqwe4zathlGKjBhKNuRrmWHHUOzG9MW/ypQ9plspGVsa9gGW5EoyhzWUSAagGM
69TZkvVmptt9o/O4glGtJ8mgwzcu4jr15w1epAwtoyurxP7EsMx3NFd6Ap6TXejpNNEEbZ7bDTwI
wqO42aQ8Be2gy4GdAGQbnh6uVO6Pdj79zNHqneO9qwWBsFGmPmrWX66ziN1CdyoQ9+8h4zcEyge2
hTXkXDKw2YwHHhsmfsMprA6OO4qgV3zLQJfBPjSLahQqawuob4jzsl1E4jQjWlVSHzTy/bx3OCVi
2Tv2ECSgcfQD4sggQ91l3+uQOoOUvMOiMr5AkXeaBUAoxWtatDWCc+0CC9D7ybF6V86eaZCdcGe8
eSAZr+7ljusR+5EvKAgv5wTeL4I5XNCuFbdQ+c1FtRmx87vmirnnGwSaWVsavLGKXczEQ6glZwh+
Nrb7v56p9lE8Qeq5HWMMds4SRc4ZE/mDn80URrPJ3t/37MqqBKavDmMhzzZZ74ng9TuERM6d6Ipw
h5DXfGPLEpyxgpYSG6w2gmZEUJP/A2uGb80mYrMwIkPFy+Xrz7Kk+sGdN39Pgep+bjrC7JhEhcm/
qvENPkgZ8UsFN58iX5rGn3u7MAJN9YLP4C6YAip+/w9E+/SFtHRfQlk6c/Ng9gZlvM1mVei5d5sG
u6ft0QHHb5bz5PhBzTzHLnjPYt9TarALDImZmRn8B+V7lJ5dc4yU0gvXqik0ET+YIPgDbr9yXf0W
sekGyO+ZU1M5qsG586VRbmYHOBuUwkvZPrkTh1IErWMiXJH2Q2/aJPcH+/Lx+xFoKY/4OhDbb7Gx
n4OV2Wotrgd6Z/v4r6YcjYYKkIwCgtFUkikScX6DIS/MucBooIlNzIs6BtvLP3H2KBy9VNQWWqtB
jLItquPRRWH+IwQIAgBFRlZ8rJW4FWOIEL6pWqnA4VFsrpzupsvEmi0zn4AyTp4YiyJFpQauCwGt
fyvwV55B46vJkcvSvmiFG9t85/opDuFQfA8UmdImcRpjUWBStnWDOnr6qX7pRmxqw2fz9VszOTdL
RatO82GzIEQfxoGYNHJ1063LSZUasEbmXvsfNhzQdaGukzvXYUIn93/7vRcyrOcyKVHMRHLm336w
eSkNVbmni0DWz4HqxaUwNd6sIdh2BAqCOTHTOEiLLHyxvQxjrt+5S4MADOBaXTZ3ccUeIZb4ikB7
B8i2ifmPSKTNyAVyJlV+hRrnZMe73SoE2YO4Nfb9FSL5F5Ksu1u4FAF3K8gBT7d1kOgNBQLB9PkF
jsxcgcHPWaU3UCTohqRlGokIFpGs3iVEAg3M/TwWoRkPINg6NdPNp1LWPzTklnp0z2Q6u4Iu7fdS
y9kwiq2uIB+Xlz8JOQLZh68gb+5CjPQG9TJTXpnfW2U1carI9EId1kD1CdhyHpJjrgxrBeF+AzMj
j/EvObz37HLYU3zdNhsJ3dPpnqs5EkFiKm+Rhl7koO4fEQcWENBCVlTFmSmiqSyZLvEY0CiddaLT
GbPE3qzeCyCuoh9AHz/CeJXnjJ/Wm9AiM0oKRJ3aDg437msVvkq2wcJpxk+0gV4Yv+UPkywvW6OP
WZNGedc8yICuuptUKWFsb8ToOToiK9apVxgaDHdTahdD30zDLPnnrWPuhCm68lT1w9r1cx+bKI7S
Sj1A5LCV+O3A/Rl8SdWThZn1SMnXDsDybjcyhI89YNqr7NxGkSucxxyiFeO5pEnHRe5+1bn0NDGU
7NmHoJ1j9xjWIwTwiD2nuArROrrGXnToPvaCYblKC125uGjxcMVjVe4sExLw0O9KchHAkdCk6p8O
I5dc9ewuQ/4JL83IFHwSTcHRHZ8PTUQFldqS93NUS7VjkUWb49jUGxVn1PD6hJLkBDz9pCC2Ekqh
/dMdi7wlkAO+hiWZXwm2ulXB9zorOONWW/I+CxprWtZTpCYYbzEVYkqqXnfjaWdBExfEFUGd2JQY
/mXduODvCtcWJG+czKvlfZBUwNE3N4g/u+aCkgeDgvv2oLdPnQ/GdDQWjo2MO0o7onPFTyL0j285
gw7TPe/CRt6qFadJ2dkAnhweIAYcBCUXKnpTFiLPwSyaPgjan7JC8w+MqLPAXCMB/nHS7SPwsK3S
xU78+lcaci9/xxUC1cZt3jyUH0TiSWibhcgxi2MQYaVOS8ngovmWuIMpFO9orvFK+uSnEV8krVz5
loBcqKUHxKsGuiXo9SYn4uCCxEEn7j1YQ7Fqzi4deMFHkDq1d1xgsNEjEobz09iBVTR3OjX10PR4
mayIpRFjSVkt/DlHeIw2a2CW5gom0+2X6ZLRX1Sx6BscbJ9RWxfHhfeRjKXYMlnT6rUdR1buagkP
YL158ZXcxx7RPyKtTIYyZxHEsL5ZYM8d/hGQgd1GsyNo0jUrNSjJO5P4U/5idxMsg4gMzJpmXKeo
EE9zJ5znMIYgulc1r0tC+570ngwJcc5xVizxQDR91GaBOGJwcOzG+d1FK1Yh5FQn5PaO+Y4mrq9A
OvZk8dKgDddPQO7hZ0j99C3Xvs5jFVjVzHEzxnPoUBTcxlBfqmkB/3++U1G1ehds94UbwtDHtM9x
u++8uoI4dv3kPmhV18jVkdVGrysVGMAKYLgaA4td/aq3ar34fQm6LKluZbE7LD7SkQMtZsmZHviz
Z/KxoJXjmf3EV291H1QndbS2p2ny4j7UzosVRijp9QYRVopVxv0Xmw3qjp1lPGtSMm0i8K/g72Iv
WX0imeO/Yc0HUw8XMtSRzzTxTPAWhDN0DBf3xMSoJVU3ihu/SVZzSWo9Yor9wyIyLuq88xUC/0vC
0jEUBfcnq3LclmCExTBr2lkkCuMR3eDiz4zXBAk1i+W37DXf2Ci+I2xiv3KC+e6thvnwwRPqx1T3
fjCN39RwZCf2Sa+rcFfn+KIlq0o9fw0+X7zilUOH6oi3NmUMcFXqx+8Ea6PMdVMfSnNOGoENfzMr
5BSOHaZibwJsUpUNNae+DtSqrgfm1EtX8JDgbtivEp4BAOR3d0CFyKAljhVQy2K1zeB9lMKAJtrr
DXmwd4ONnvQJiqR5Skr7Suod82fy3wFkW8szKdITNniPEtTbRh7cWP7CRlmZwtgzCX3gKSAABSHw
t0D8ftTHvARWekvawb6q+pBXW8eKXW1iYCggeuEeTNL9i5boZ3n/uv/dml9ofLDJK4dEnrF9uH8f
/K+N9eyPn9DQ3fBAZxmaxBnokGdmyXlHfvB65oDBPZRPu73+3xmZ42RgeC6ix5nwFMaFpOTa7vBo
xo5Ycl852v3Xjdi3nzPtI0rtS8I4E9ERAEGkHd0O/AkJXLhRCNpaIeWnXBlRKoLSU3tkKqA1P+eN
AikjhXz/FIfAHKs8g8ufVy8a5lYuzLSSCYe+Ln++Rpz+ib55RiVmBD39VLyosUo7YG0UCBiWkpxU
CaR10CrhsyaPqSX5tae53bGuIi4SAvlWF887EF8CmGLNuBt+liM5q4Z0wyk/2FDFtWQwjV5MxlAl
Wr5INtoFeB7gIvLbXFybAVNCETuTz6xE2VBsTTnPW0hhqMzU90I4oNNbbnrLrG+lFzMrlXLRLESM
4jlMKXzeBFMELrKgLXQngv/RVPqHI5DnJz5whJyQBq1UzydnMizLAvWmOUVIX/4H7RRXyOLLOCfX
bYnH7ouFTpArxQiBT8aQ+ui0y+QT2cfjmrGChcIsko8TwuHs/ZLNT3ehIB9Wxmh2WRZjEloxHQPL
ZKljhR495abpwfARXYEN1GRFwLLepFyMe75uqkqJeRJODV2qp0rBuzbTsOztnfZvfQmK+O1vEAP/
jPdHRhJ7gQxsNijg9SESZZRFNU5JH/GOdTwLLfT3IG/Fbod0rtoDVU5avvKiRY0XK8Bchii/rB/9
ozSwg3Zkgy4oLs0h9FEyzi5vuDf/y/sDhcsmINzrVTET/u8dBamMO/mD0pVqvKzQ0SxiIjJbmZOL
qNj84fAMBAKf8UoI7evOQBmATZ0oNDF+3NhgVH2pyevfGYwhqKU44WDZS7iKDij5yEgc5SbvLYz7
7m0ZP4CiuwoQKct5mIHsFhGluydC/WuAE1nquZDt6WASFi7a7Z2MMN70vPhRoBVJ2G7H3uhx3/sF
D8WHcmkfm12bKYc5pgmHYODC7Xl+nY7qkKGmsFhnWKzPuhRKoI9919ybhrjnb76DKeLbYSO0jdg/
R6qOQ78o/xlY9hPd/leNUkgUbx/gESRI1nLZVFY8w1nYRDa4jCgrO3LtRbli/wpI5YDuhEyVJOqC
ZQqAFRGQtGCRF1VcyR0XICATxC7h3/0sMtAhF8SalnSZvUn+Rb/jotBAoNaA7zjWDaJEguK/2ih6
YJOfZplkIrMUlCZ4/D6G52RfZ5WBF+47JUerpnTZiNbsbkVZDBPufiwcXV2AVZc9a42T8228+1EY
tbVs8PfEx8fa/gs3yYBJFA8I3S17r4Ea4xH6bXl2qF8FtJd0/gKqrhGi40reFkmMoOXlKLuHpMax
htVcnuGhPl7wRVvdjjYwzUTi+UlnXfRlWtxEC9O0lhea/sZPb2IU3hTiY0UFP37NznPrxtk7UNn8
tgwH7R3fzlqnwzTNrdrDmq3KeunK0YxZmQemQYvMoI+72hulUPkUjqB1eUtusZZ4ezfJ1MUgGU2S
VJYehtVkM28i2OF8U9VySjq8EOoyJGmM+0Mg4vHTKJxyKzk6hrmftNXiKFYo3mig7299S7XlI+Pc
wkN9rVJRuW6HOyvWhEUcJeHmeSaVOewHa+4ID1dfIsf2tu1WzhXWX3hiAzPWa9yBp1Dnj3ZUOUGd
ILMgOUxp5UoTMftTMc95ppdZNv4oY5N8Hogk9S1yfwTepdp0Za8cQMWGZgNFnRvTlGWlcgRP87zL
gmPbm0bkFnIja5DIKES1k08B1KZC1qHnteIrvjinfk3vASUkfG6yq0VtC9r7MFq2808uz5jv3Wzg
qeGnz+1a2CAWfspB/dOz2fVAqlu7mLpLTAChAghgDDPlU8bIy0Y8Xnpb8+IQyVFNuOS1tOjBJ1HZ
X3UEm59Gy82+F/7a6pJDG0YYWM2cS3mQaHT+5+m9nPJkfMYlmuSMOqwOMl32o1GwWQzXfa/TLWEz
TrDuOYdO5UtyHHOEgX4un9FbztxR+3y3LCxrSElU9jdp6JxU2O4tuIJlrr1DV6bDrt39VfkSosiI
eHlxDorVSz31/cZfVui/iwja72DpklHNC4z8KgzYVcbc58k55QXaxR4h15Qk3bWBYdeBhkzlP8j8
LevKldyzTiVaWeyDx3nz8VMu9MdlYeE/0fbYeaf5p1ReeHI2ksVQsRgI0R688kkLEjgUGIITpL3l
qQW4FJG4OLuwNINc6uwUaZ6Z/snigvicind0cynAUruqbDul2Fe4INJ6gu8cIqZjhVdK+QKbh+dZ
mAC5f1kzA1gBzkzk4jtm1ZEZtQc/PoCDsEyKGOSwSqRH5NCal9vJhxYjFb1iI9sOq+bFg43A2CMV
YpRV+plzqiuI7v9OI20rXtBbBk4KmRR4bBfcpxSiQcKV/ffnZJRpBjFL2Qj2AeyqepEEY52TG/qP
sL/+300AZwiqURVh7TCVf1Z7H7VfFEdcjGPL+HG2PBVYwkZYFnnsFMQ4n8xHnRGTeOi907fgCgWw
tZOpL5ygnamdAHmx8iCMuXFIVdS+rjDx+7tZ6gEmTTJ1lxRCECkKV2lJ0OG7FeGwA5iE5efoKJbi
TKpciBy/z0O09V488hxZ+8yxzZrUyxLKFGPTsRCdYrrsYLMfqm9YA9vHGq7HORPyh1p/y89oxT1+
G5Vs1UhpFPhLdkEMd9mj7onqsafNctlwCqHJJEOerrPWuzW2PLxcWNx/Ef2NCKfeBLyY/RdYSNYw
vTEZTzDSYO/6Q0vvwKG16LKF1nn9r3ZhRyyJKJDvkQAJY/G5gs4b/bDu7SmruRT5srlpOnbMX/Ks
HMPSa4ZX4g6hT6MIfrzOrlKgR2/jOfseGA6fqWFB+HtQ9+XkfSXC6f0mMsrEDCqD9j5hrf29dHLr
QialVtjhJd4G0RtLDr9LNO32EOJ57HYTzOkmfpO5CD1qZ+0blCGxoeFrw7AXNRo7DrZvy8cGqRqu
guV9P8kh9zRLm0AotEgupBmzuzKeiG0ifPKRcTm/iUMGNEnh9orZQycRHDAVqTmYeoO4+z+RoHPy
5+uJX+VhK6iy8crn/MNkn1Z2uRlu8pmGpTFQOd1wMGiYM3dhbTzCfj8oEgm3gbLgZ66UyODv8Iqd
dA74UW/EoPAs5YSxVr0gUQdzd6QTEvh6pE0eUBiOeZRQAGyIKv4ngIobMGQRybK/M5reG6QlY6H0
OLxc/Mux0v1IVzuDApbsqf3+6aqTm5CgQhbj7DNTQu3tq7XgG9n15XLNDSNODPOQ8GbNbqd7XcGt
pWPs1oxb8ZdPgrXzyLRlb2u0J3AueCk+/VH2+s4BQnQNzqFQj2ZbkAndnkCuWnWzW08QnHG5AMei
48J1lymhrm+mwHSXVVPlVGD5DixOc0pH6R17t43T0mM5vWvZE5M3YtkR7ifxlQbBkdgsC7oVU7TD
5pVvBjswxVOBKnQrD+Aw7eDcfQit/4yVuj4aPOsFnqYvjeTNwvFLv/3ts9kVqz823lXNJRkGg06A
dG+/StjewP65UZ7vLjdll4LT0hC3yvpmYk83G7ygMDa/QCaYnTgFtVR/7Xz2MEKLAsK8cpE7IpjN
PqmPI8HwsvBv5oVjAqVQTQTRsdbTCYlNPCF/oQGYmTvbsm7metPlenkpIZLRkPhqnHlLZIQYPHbQ
evWtst1ubomWFn4vs5C4lck0PAXuBR8neFJMvVT9RdKzhT5kXmSt9iJZhC+qfnIOZ5iRqUmmYpf0
zphcDWqL7+U31w8chk/6Kk/R+8ah7gwDlQHGuTp/VVos0alVpBqC3KIs9EXf1zS+4ZWFOUIfHh0t
l2FDXwKRX+DOWm3TYenNKbH4g6mIryZAuV14oefVXyCCn3Y8fB4GW1nvaT0QMCPhaY/NlgZWWq1n
4Tsv2Yfbrr0biE9KpoXAuu8fQFuYNL72sCsMpOrzQBp+aUouTkgPSFEyYKX9xiSNs9Nc7KPPfJE2
tXTTRh3vY4gEzP7jiL2m+JyvnyDLOYXLauVAzWIOFEIty4kU0pkYkV25DnYBzdFVpURDtIs2M1/A
ZJDITXlmyuEUYbZtDO48S0Rq9GFduGJrLJBM4aP/MW4sFrucrIQYD1QdBFWHBbnQY6pFAqVFBb+z
d4iu5ze4o9kTT65oloyF2bitfaOcuUPenvN9gIbYtnDazRXfFErqptBXQ3VocWJ6NkfY8jA8W2Sq
S3zbP8NiaOWfa080JHwMwM2rQS7BYX/CXivabQDHghY16dTYW5mlheoL5KnFRd5T8PphF32s1JWZ
5AEB5AynE/2j3U9C2b9KjDhqj6Z7I5aY2hj1fUk/3Ug3vq2FjphjiEl+lZowIuHzpO6Y5jOUnHiZ
dcpvsAYO2NHpZGzR6TNxihEwsK7Em5PqgWGZjtkNa22t6WCiV77nULT5S7Uym7Yks8SRNtYz2LuW
7LIr6QRurWxgzphxyxObYse8PDwsMiAMkR/uiFZlj2Ryc4mNb5ez/1Cagq4BKKXa5eWWyT0Wwwm3
77I/Yv2sFxY1KX7bVe/NMxZa35LjVIbdq8mFZSlckBFJOMsszAOICMrwEGyeHwW1EJJqH5uqJal1
MKofFF7nebDhlbSY4QHxfoane8hF/GZy8yNKM6P6Bj+LBU0lx+XFLf5bCapv2MZylKh3TzPvSOc5
9t715eSCPsAV9QR3f6ivLhrefmKTSHZDHa+3ZnFPKj/n1wOR4ZNSL1rLQrccb7aKGT1MF2Srwt1s
64ElDSfY43YKR8i7G5tOvjZbPuD7XgX5nziMGtGS8Pi1Bg5bJYy4sH1fhDiHMiYyk9w6ezkedjCd
vIGCOUDipHMYc+qdlDaf5rFuYEeYRlhDQAEUkeWvpQ26UKAgdGtPKClqL7g/cy2b6lT6zaV7XB00
tVJCjYVtUXTnSCkpzOwhCgyhIxcqZzA/fjacj43V6ozwPig7qgjlmKdC+gajZav2XfChk7TC2eQK
9UF+lLljL+ZwR+zdceDjKLb8U+JIciEXdmN57zWp0FM3FTS/p78CDPV7GPmDZNeCE+pv/dKxKNIY
zAH6xCOPiA9k1lYnCGkTJFAPYckEh0cjxyg2V3G3eH8tJD8TmLGD77EBvNSNG6D9NcA6DyOIFw06
5ypcMaF07LCVa65iLAKzfpHfdO+Dt5/bLH103QcHi0LPIccUgA1IeR/z88t2+UWOphQAXqHnET1s
kknEq5HT/Hn9uzRKxehkeAPRtotyqyejZUIyzMo8JSml+8ys1dFZUSmLcywYwIUCxZFKrce7adyL
9pKMC2H8ggmLeKqJBS/H1dLxXagqanrkOnnIsl6DzdOuGkzsjKeJvB1zjVONqBlDDDJwYRLAC651
iUMyQOtBhnrv7cAbIsAfigYvYqVFUV2lv5sjGakkGgKWU+fgEdKrFKc0kaYabAqrFEsiAiXFqyMU
ziC3e5s8MDP5xguSujN7WQlgdvwZriHpJuSLAG2YG/Obc0fHSkTFasCZvdVRKP6NeuYSzpEJkDRw
5CyBnj6gakPmYKfu4uofMLZE6e156VUotPXcN+CL7yyGJ+gOHUlunACgYzMKVn6qWVLtuyShpTA+
q7rnW+TQQpugPds7S6RM3iZ0yAEi7tDBXatXTZkztVgBZf/djntaHLQs3KFcWZHnq6a/MJeNGtdq
gzFmh6gc5NlhUPyU+BWdmLDok22ZA7WR10o1aEM4z1Ejg8btBAwmHhWlhqxTvMuCsnQDeqCJ/ZHb
4kjnfN7MXlvOkmiaHWrA29gtK2u7J9iudZRGBWgi+3Rn+ToI+SLi5ev6dYsQerYvGCDGD/lsGC3j
yD9n4xPQS/uSPJOxR29sYj6euxmI4jD/hjoE+K24Rbr3whhBCQ316+UdhMeyznO1IANrP7YYFdhS
zWtbsLHjhytaVQdWtVrGf7csPDS5x2avoHcPHNMX452n6AaqtvCwvX95Q+G/p5xZh2bFb+T32Mbw
ApDLk6Hhyp95uSJx5qmnY3uPipqJ7SJM/Q3anjGs5EVSIpuOEkYU6LdPaJAxzoWRszjhloeujW03
JgGNt0VmYpPJySjTNVk/7T1eL/QIe8sCuohOTKfvX3fkesZ3lHFMsJA3cDBY5Tomyw0f3dyShDv3
xbNi60OBZYxAJRxuRCfT5V6gIJKM+STHwnAzFULPx3R7VX7EVmoQy/O0qU3rr99TLVe7qah3MsMB
Qc4dAAyLSybwL8/sagT3xm8lhGVz+2n4roCV+O3xbDaLi+fHOdLugGH0vB3XMoFifB0HwI7aO9L0
RX4DAWyvNmMSCLU2JW5sH96XexsVWHPcldO32TEBiDsIRmPZ85CkNQTITIzAhHmI6ieITFdK+sbI
r17+Ws0yBppXdyAtpODGLkpL6TkfxAdP881Sg/OmlXq0YpDYwJxGWY4Xto+W6baVWI6AxGJ9o0Ke
7C/Q5cl/2Rns7nLdNdAbpUCoFRbJ/UbE0I/C0MZUQHEYMj4l4800KiR4cg7m5C+U2ZsHJbDrZNWr
0w5ag03YALL7J525KniH9bpjPsatqoZZKVJ0bfAfTAVSiGUGlNM3/xreO3DnGe8fqaMMXtJX4G1h
WVzCv46eGZoWE5yW/E2V0dwiqdKwSgs6y3WlyVNm8FTkTREN2yhLpmPzt6Zugyu7B83xX4fJRfRK
kvhxtC11JLS72gWJmOWzrvSVpRfOHWncnB8o6RFyc5uOZkHSjHXMFCelgYh4r9EYjzTO4j5O58ER
Jp+UZP5dQ92FGPUrisBNIR2K713r7+UP65gsNn+yUA1Jvchl0ksDkb53tpj7kVKvUWzi4DVwyZHj
AqZscJrhk5ZHpiEpjV/9BPTeG3u3J1jWj1s6MTC2oECBXF4qfU31j98XTlAjBMFN0W3y/rJeiZtQ
7dg+yWNo43cmtNVvNqlUGE1yEICoi5uX4PCb7YPtXdD4bmtzl/9Wa1wthwl8WEgeLtx8ntKXrB34
uB7HjPkriVMLqSWqa+gzop2HsIkuQ13TOl6XuqdJJ54x76Wly5LwyZ1fEirQRrt1WnqwC3Lq7WNc
l9qOYrLiTubYCUWfuoMXUiNISBP2uAvf6GnqQin2TQRR3Hci7gJyENZFblbXbvgQi108EvhZivD+
kp1lURm5HY2pQzi9RPBBl9WKCqGTeK1DW4rVJtgPCKC4X9h7C3dIcmu/UYoTrT0u5A8cxZcNdIHi
c6Q4/QatxB9zAe2frlZlN02YrhuufZbsVHpRMxm9gV2BTLSwlMZpgHMpyUWmjx3GDm7R0Mwaji83
Jv6K2qvlCuK4h2FrlpEJpWCr7+oQ+E2o/qHIPadG02hk41mmbTF+ivrz9eua3unHwFllR385FMlF
PJMhmQjL4GOhvgrp6yRubieUEAv5uWLddj9n7UvUaBrd2uvVQe8T32T4WgqElJoIsHWot9tbAxGF
56T4+76gSVJL+A4E7FnPZxuWIe6CMrPcCAFC0VcTB1xPNGm3M3PdgoXrzNxgAZAXfu9z2Detfdx4
54sRcQgdIy33VWpOAU+mfOxB7Bed3mEASgZc7K3vzOAiPnQg9C2nLLY62xXV9/KzyfpD9A/3Pz/f
9V98gfaQi+KRE75ZyBcwzYXIUJyuERdh59E3zQb7M6OSTMrVuV+G2LKvVebydyD6pyR4jQcseqrq
oZ11EobiNKj/09y7lDH/Mvy6an10xLWUaf67RPMc5DqUmSCMR0ss2oFJe7ubVKe5AjbDP2XDuX9L
eCBjEASyR2wV+VhyWK2GoQ8O7naBQPtVaPt8w9B1DZgXO+uUqmQBRkiTkfeNprtgUCGIY7u5MNJa
GqAOStxu2e52fwyfbWnLcZu3icWng+WKdwrY3gzicN+JCJQHc5OTCgIRcWYWjIyvSwm6ph6x3t41
Yu+6A7hw1JM4uHe1HftUz9SJLZ/CvS0HyYn0VaEfolNrnQct7ZVqD9IuZmNg+qSppwst0XhnRfxZ
CrYYsBteHTXDTzSF1sEoEi9Ii0q3HZAC/8LOnxwtoELPwPM5R4TsvjJMBliU6ezO0583xSZuxjkc
M0INqhQ8QBJ6rs+X9/tSjcnTZFZjsEY4gzR0rhQW6umLf9D6SYENQTmsaJbOuQi44WG9O1HQgqXy
RaJo7jjEt9IMXhzc0ymqgff19u3st357yqjk3zVuqn//tpvrmPIC+0MXx2k3i5JU0FvWYsdryD+U
UstwxOJZmdEp+L46Pg3WmR49ON4/mJ9SjSCQXka+/CSUT1B/CGRHWm+UlK8m/viHEuIHHRFJnDKm
tLvu5d+eQLlYzDjr7ts/25oqzt3Eh5Fk4wQ7OcQEGQRI1tyDaG+m8Y2Y672kAMLPcRiCtv6nC+xo
AkWZv2/RdBbZp7ZvYuR5Ti23QdeRKFvHnVsb0U/vQDXV5rwbJ2WuuIwq0u7z+LbkVyGTZfdTd6kw
JskjgaQ/3ouXq7k3u7o4minHw2ILxNMSNm+k6ykRe4NlN4e5mzNM23xp/ow75Jj2MhczlTOrzkQt
uVsdVREJ2U+ZEaW+Hh5j4lMTtMalfhI2qKRkOtCK/+opYp/7IL9Yo+ClSVjDqfb0URx1bNlQVIib
BWqwdBWH2V64ufgGofGEEYCoLkT8jQ48J4rOiqefMrkFCJfZEHMSoQd1BfZVnHNGCz142wY0Mteg
1HASu62oMuv+eW65jyuxybxZcZnrDmP2QDdJrDkxC3/n8lzcsrwFOfJ3YKJ4anM7fZpxhhwjLxH0
MHyVyhLHViotonvHiMM1ahceu56cfpXmqwCZwppdCdDOfU47dZF7V+D4EeW9Ek4WLpf3S/BK3IMQ
kWFyy5T2BhKs/M/fudnqlIl3j5+Py/HU/YS0r5ec91QJHIZRbd3VcysgseD9s1vkQsUfutcoUYFd
0yWiNU5v2oq9VjUpnENFP/v4AkTFD2NBAOTg3r06rwFV1Ml1ckR1IbVP0ybPCoFuqm8JlwnHtZnl
RkckpxDtMlsFQU6xkKMtMmsmTCcgO01m+WNAobVAT3FQ2wA7nTQ9XzEjzlDv8z//UkqOP6PAziAe
OwrL7w5KS6fSNGXTU0WaHgfTPSNWykF8VKt9RGFDd2l9NK9WkW9xN7XF+778N4WyyS2nFvxzuKZs
MGkUasPnzdIFqncvE8C3BeN9GefhM89QwwR+wFEHexExDObWD3sTovXBbVdpnTUIgR5DH92ilcBF
mKv5uO1hUuvJCFSFyxvSLA1k5N+i4IBPPxd9MzoppErfMCW713Ez3+9yUhDyscvEum+88Qha9IoH
uQoGrCPRDRny4rChCnpb+SnIdWU1cmTqKTNaUuKSnx4T8nD7f+R36iGaz4pkg7O5nUura7RgCSoM
vDdapY8r6TYvJOpqS0iE9oLEpYSlwX4N1S/8UPCY3N9izU7KVCJ9hWD+PYwY07N1w9oW2xRyy1+S
pzOBY0vusk3cLNM6xjGC7wghR7yzwNHeU3m2P4b0Q6RP531sJbFsBhXxkLL5I8/DamymlL79lRLL
6TW1m0lHP/6gDlYxQ75DbFeozbom3cMEs2qIPbSVhcMPp1WdpEVFtwZV6qXorM+BnYil5t11lh3Q
qtAmG5+k/J8zNJ2NWn3yTbsAuEvPvL/vw5LQYbbd0IFiUfjtLv44C94Zdwy9Ex3d/hAubQtvUcS7
6yZQHOTMF9X162XEcRPXetpVdqNP9Sw89gWbgZ9/tMWNgOz+LEFcbVnYRauC291Ueqhh+Cc7gNLC
Omomoqmr0fc97tu2fvcmG3Nady2nB0GhIhsdg5OYQD6l4cfIMaN9UVS2w9dUdukvoir9LmY66VLm
Hhv3jNCM7c22/uucJiBoHsz82axHDhkz87VfdE7TtfNkuBl4/6TyxULnTpjBlcF7cNFuBN7PuLJk
ZgUjgjWfd6TE5NYpIqD9/f8NzY6rsHh8vbZVJPV/XBsH4QUEyUQj0JGA589/nu9xPuS5LglssNQm
47c12b8BGDhEpjhRo5MLddHdA/th0/C8JHrz0TtOk5nt2e09Jc0/SOtGlj4z5KgUR+l6EQEj8F+O
XJfOR5f5KqkCcntrNyx3WDP2+4dXjZ3gzRdZTYvC09Z3rZu5myiFxjbLmp5eDO5GImVepH4UCJ2j
/5ES3IVvO0Dq3Ear8bGnQE36RGkG8ygNyU3Sm5b3iSmDYm0QNEQjd0WLnWC2iJPtp+zb0J2ureer
K79q52NJpg6w9ZSd2E/jBCIFB1bA+vUDM+tTwoipaBWqLF6tX5KOWQ3YDSgiTcRoCm+X85yHVcWd
I8hjAbrGvU39cZ6+b675KL2FYuXTr0FK9hFI3dn+cexT9KqzAdo8iD/cQR6DlC5dhvMcr7FeVpmb
4VkgbRCH5DPWanvkgAVGLH8qpRHtmlIAouvgwL1nXyIjgHceJedyQ+LSZkb1yaFCbR5MAxIMibYq
ejBfIPaqfVJaVcAU5WhELR3Zwb0ZIAEu5eynHzZYb2ZJLMD4hIy/cmvoV2QL7EIQ9JNDtgvPYBsK
PO6/9iIpyjhU7n7Jmdpt+YP0LOwxsALOmB/0dbjFkZv3jknryiB8uDX2c4NNFv4hdbMK02MfVTaI
UA5tQqOUIITTDxvWpe6Y0JuxUioY7LXgoiinW+zMn3V+XwoFfrHi1I70ELvZFXbMxQM+zRcA72++
Bw7Jjlrv9aOgPvyyhiXnOtVN42zp2U6TItyMTp7djGJDY5DnNTx0R8c/ACCKTlNXhrbTfARGv7BI
vxtnaQEDmUYnRAA7GyZUavONrHYSvqmGAjzW/XUjfkreFOV0fgDVIzsCzKHQgSTUTGfsWFNRdfEc
XjGC55IioV7WKgXux15xBgqhGImxijUJ7793Yv6uCmU1G6b1OkI3Pju94XKQEzITDLip/A8rEo0F
IsVWH7m30P06uJWxCX7UPgmxh4DQTNuOsbPQabOQ1kz6p2L94zNKHexBoON+ig1XdXkffqGA8W/z
98kn4Vgve2durkPkaLyosykNbBZnV+V1Eet3MXR538p4bUNSzWInegCLyPMHFRNZBfOVKzAzOJqC
nAydFk25xn+fXnsc5BUyMdIwFZw+20AvmUcAdVlu0WNuqNZb1AXNFtQDf6sU8DK3rBVSrGSAw22m
RWLzLkIWSxydRKvCOzDvzP7UBdLWq5huqvKt5tHvtHS/R2Nik7IgdoNx/ORTX44sGLSCrnvhgXI7
sBbbUPJaz6UQVPPx2SiBZSCW88Gk+B9OOrGpwavFpa6gyHEYXIh0Phv3Sgq2rYIY5davSopld7Z1
lhQsYK97JKCABUjifaWfjtnAA9RNEo4FIYxXFa53kSvzNVR16ILdFD5NLyJ+ExE4aPhioRNIhG2B
wVFO4R+8fmWG+0XTUVjaTl0Beb13b3F7LV+hcwSmC9mvuKF0zOMfdwix58+QOdhj9WsInpuli3DM
ExVBlJuo4LkmYEOjMokoWq2XJYEh+eCONnfuGJU2divttvVQSA4KsFfC2Mfw7Cxnupf1iyDbTAqY
Z5zD0B+BvBWrVpFGs3c837UtU7Y2j3DhH9YD5MDepQKzIZREYBB9XtzqI83T80+otossNxhri52G
Np0azUUHJyfz6XPTMntkLvXYsfZYm2SXoKigZXqFrUTR5Ij9JoFiExBtRCQGblL+hqH6D9OfaAml
B65GObRO9TDz/P+E1bsEHz1ENlPLro3FI33zxolL/LEvCxZlTbNPFQ+IQGcY2WX6P5GL1k9rhdA1
Mbg2paTCDyz2WgLDI4GWm9BI2aWdXCjHHE01YZNsvMb0cr/I6fgnS3XuGzEbrT12MaQdkofBJSTM
KNuPX1OCfJMh/Pnj3t+yTctrjRv+IxhtlDRAd+YQCA/+G3v70YnyIZyNW+SJFf/O0R5qC+Rjg1Z3
bqJHnAB5nEvEo7xsWl1v6D0C1/cHbEToqYMul51pAn7lSf/EyNGIJbZxtOy+Y1mV8cOe4MJ5sFqi
9QMeuy+kmMl+GBhqeKUK5FxgB89M20GHazkF5wkpU02Gt08KkF58r/mOqosj4LdakbRvLUnGUdBp
qsBkzmRwr3wR6TZiACHsQicFkQ39cx35dGHNtK+N6733Kgf1y4UB3brP55FdUGYcYgm76b8NqjYB
MNU3gvPHmkqaZuFzErtfm1QSiGFSBXK9UxRuVzdWYdUwHxmtn0b9fK/LQXdCcDbUm6GcfpFiAIRw
f2e/g7Ek50L+TjBCD/o8hy4/l93A5VVl5uLpjJP/rjQNYUSC+IL/42xFaILn7qnPQFOiaqkFK0pI
mXrqSViPjwmx5geR1+5Yv0aT/CViSUn1KvD2G5geZghmDwDz7YDWxeEnGhSkiDg+c8KOGb//UIwf
Xg0xDXNelx+qjrQ9KHN8J7oubzMtnGIRNyOhiPiAs9PLH5Xz3LVsZkAfEL05UOvggmXlInt2fYVh
UcLFE6khaZ0Abd8xJbGg7k/LYnSNMst5YPjMta1Uo4y6LrYRLP1Pv2OF9CEFz7thoG10yBFDlxtD
s3NB0+FLY67xsHj64chjNQsfktG9406LQRS8ai6/3XMlkn2zdHzd7e1Abnre3nFi+nzWCmCKlw3U
kej3fAnBbs1BcHY3e6qa6QIM4IRdFkiTm19T28rJK6ZzCemzPyAZds2KzNUhdhFqigXuyCpECdnv
puQPGvRNj3UpZrqK4JzrRNXDbHkH6lgGFkEMDWGhWG11rEfY/NLFOYO9GcDcNwXQl378VuSgTQ+3
7ts85KqjaFR52OnSg+q6DNxUT1Z+JZVit7I0pdXGfQX28MiptlabDPHOauNP8NGYOqzVuGnRYn+D
nQ74oYD2PXYusfj9CDBpVMbpU9zVvBtMAq4QMB5Ie2CTFmGPQqdzGM368pLyHfoqykJn1uMO3Mf5
fa0J3xgVTa8DT13bDghQnfGD2ipJF8hMtAoWiVnN1iQwPTjoIE0gszBk1/ao4HDHuKy/m5LYjeQz
g89qxM/QMhBmhamnzETBm6Mre2bJAnYsum4l4mHyZTe+CnepQhO900jyZlNerH+Ut+3h0a46atK2
CkqUu0UtIHEWC4Ciba/SVLAp9laauQHU17jQpOrjQKuEqQgcJk9EYbcj3z4/sG91Os8843i2rPsk
zA3dB4laOGV2Rl6IevQAT1S7P0dXqPLcXBbQVkrIHWYTlwvNFj7iN+7pFdDNfeiNQAA5HzJfF7n3
3lYrf/wQIf8PdrC2NcLVzpCGxSfpTZe7uQfWMueBQuFw61RI02hpxwSE5TqzflqnIfnurz9lOIDz
iCk28UaVZXyXM1ENWol2SDwMXrQ9uuLPAe5BjxrPKNjz7HejKlzTkrcWoAR1MY57jfbDFJTbxey6
dTFYxtPxiOTGXh7dwTtxFH76b92LrLpIxZPwQi1O+n1nHTcGFV87fPkxVv76dOSKN1LoPlRkYvZs
uSFLOoZTI0+yI0ti83iFQ2sv0ijRut3MKfcvkrv14K53il7Kiuqevkpdi8p8xYI6qFqvJcMr3Idb
bGgIFTxl7dk0BDssumWsiPM+U5POHpkzHwdYMv2pCpDFOJK6J9H2Q6HXVwNm7JvXmizeDcnUKr7Y
JKHx5nkeE+bRftQ3xJe6sVNtB7WEJ4zmZWel+5HkwZjF2nq6jFDG0bDz3FCBuw8g+HVjdGuAGndC
7w3nWKhrg+F3WDovsywS9h5heIrVAEjO3tu4dGIL+kRxbJhfFvmHo2W7+i20iPdAKNFqfW46GmQF
2Ym17upz8as71Vq9k2oGq1PdycCNDhHxAbK9Vo50ukhrNrxJovnnuwVazJIB/cdfeBg1aCzFw5gX
8Hc8HUaEJLd5bxv7cB2grVXsuI22jNiSpofJ0geOUHLnHwgtMU7NbDtA9eQ2zgC7fcouYuEym8Nh
IAyYcFCF5H8URcnRA6Tr/OqecixenCLWXGpGfbZHjP2oaKrSeo71QRaJpDa1IOa1GmGd3o72pR7k
46h2/23uSXTOGvU0ZWRs8/KnT82A6Bn54x0q6NGHvYcWY9aVL4JLGyg2WQH73uwvjA5xDd74siNS
42Kj27pRl2tUxmoEIO3lF4PN9ANTZdo0SEKyUx7Eg+uycS8AedB5p0fUJDQaZljPwAaaN+3BtkJG
yw0N6S8+HZ1vgNLqOssnK9ig6rJZw+zt+SwZeSZbh68DzQ3eVlHkWkYtwOpBDriHVdwLiKsQia7x
gyaWvGLg+Eu+3lpXrlolBI+zojeAG5Gl1whGjjV7RABsCwWBAkSJTEOpMtSLzY+2vqaM0FGGE1HQ
52PYgI7VapRSCgoN3OmjVgBe4SKlDTzD+ts5knpRiltk1p128pHIeT3MFbsoyuCyYhck3o/Prh7B
8lk1Xh6EI9SUHyS/ZUnS6DFxfzw2RNDSpu2N+NzCU9THn8l1o/DDzQlaMezhifnqFilLDcvMp4LA
0SG+0Tw5EvW7TH/PzjH73HGYdi4ze4yM28LQER+4ztEzFxUbDoGKwd4KKbOShhPd+lJq+XPTzHxF
zUf2WbToLhm7PPQYFVR6A3p+cjX7DO7wOHkJ94NxXAWm2atciUddgPWCTTASJZcIkdzZni1coyRJ
MnCBu8Gy3CIWbyi1kA+m20howrTlDv04mV2uE3KbUdV8WLimc3Ctwt9qszwdZzdMRSSm5qOMFN5s
5JQLYo8foCXCV+i9uZ1gqHDDfUbfyIjVEB9BURjPjLRyeKx65gU9s4XlEssrhdRiOTg6jts9BIza
W48hxRgONIOLzPtgTCsfokUForee59gwfKagXXBOM9pHjXo+4fUUTeC/KGW+g+huQNGCtvjhO9Ph
0KCao4F8Pl3AJyRzrvXwQdRjyrmzrduQ91XxRBnZc2lp6AjxmzHIFGI0fuCYQXjsmZeVXSgWW3Hq
F+O5EkW4ZsfSUZ1YBOnonyXvs7U3TTRniYHJStLvBFf5s3Wj8u0zyx6KN/tjF6AZ/nFtA3y7inm/
yAT3KUULa0+/ptiWf4aokef06E2rLB5NZs4mB0SEHP0aU5Xf6ZtpVjBfk+apQfG5OxbefB0W5rbx
lI/dIQxVEXY69Jci0RVRRUTkZn9K0HwCbFHYDYezFrZp5bKecCc+wMV+609zALKU0i+YzXnVHGOm
S6T8z7xMHmnHKUNRbqhtpZ+K4t4FN7qsIa/51crpRI7+mPIsT0g/MTvEbEo4oGZ7tJApRBMrplDS
4d5dCoI0aNS++Y5c5B9uxEiYsmp7+NJ3GBDtVutQdbnB1fdSitBBxk1OxaiXOkt9clTePxAOTpO8
DkrUF2xZh9zrZtFlTIsltaL5aUntLDj5ymqtiZI834crS9cV8WCfqdK1y6ba4S9NKrDV/qVWfmYr
/E0cg7yTILtPmZabQIMndLtyhKfa9ua4HDX+sli+oStIxMlrT8D2iKOhlh8OTfpEpWDtMw5z7DPN
Qymdv5ePigkbrJVfsEm8R5paI1jNJy7vBxYkqAc4ZCogk/mCKiTFg6rRYY/BZfQHr5oX86Q9hIh9
wjZJGq5SGtojoycqT+SpZuBefpPiKnEZG8gLstWwekU7QdUaK0Cy5GEBhtawXMKHnEcdByWwlDRF
xaImZSHvE1/LEeeZQJhh5hyjSChygCYBZjjWyDZ4ez3YNQ4hmhKw4do23oHFcQTKDTzc7taSdDmt
Ob7VLJI/mt2kOhp7MHKoac3Mudd2YrpKgsTYjRrrXCFejPfuFs3xqItwE5bGF8yvptRcXAGYYo62
Pl01SLdynPaQuhHB8JU8m908I7kYzokam+edTmPh8mSp+wyhCNuGaqxtTKDK1MWJc7iZqP4IiAEm
ggkFjEnzOR/LbVjZNyyGOVZTbeiaw/y5zo0szAzX9WGUsrjyiLSMQShqQ1eM6RMFRnZB3dbuy+V8
HY2zEmIa0mI//3w/7y/+P2jyfYL68DnDfCFgsevfknD+BjRGhcmQcAzkOo95nU4AVzAD6NCkg5HW
h2m5/VycLf2m0+/W3f869HZj5PkYpKfEe9vIShZOm29W1w13vbCR29TmFZ0k4uqR9WmGXpNT061i
x/m2yg/gQW6Aj1qOXjpsU/+bKGMPVf6XiMkpRN3chu3rtnT0c2T5gY4M2PcmmmTzIjcdYTkfbM6y
cdLklBxSP7eflcZyjM4g+2u6PL1a089xr44/9XeOQtidwbkZqh7B2Umg2pva6KReOTe9+vx7iDp3
Oa1UJL9w3jmd3nSruzkFclTxRexOoPMfIK8TVJc6BxrTgyYAsG+5ktNa1+xfExwowdHZ1G/j8ljS
+/K/nrjmYXNNqdxivGS0fAxrYlxwHbd86rYYA306X5hf1v+C7rlzKRKAUHSvKIUylH+StXbO7Lwx
AHfRYsgx3va+AhY5AWFqZZta/2/E2f8FWkWemeHiFrTOH8gempaGtFb0GTZgTsFIlJnpWhqBQIC0
m/xr1mWDiD1KNepa8mL5hJxqxB96h/gEmXh07iqbcVq2MDw2FWolfTcIY6yLH4IKQ7B6HZPXofXL
SIy/ecZbtMbNzW240uGnPKeFikFRb0kx5fZCf5xweiV0WvrTXu4RapwwmSkVJ2GGgAUoqzcmProF
N0nQK8Z0cdIWqxzP24SSrCtAIJE+TScTcbI4agehg0GM3fi8iSXcPnayiEEVrDMnNxBrzmKyfKAW
ExGgRozQdKO0YslqXcRg2nr7PHraAeh2iPry19x6KOg2gE/X115RzCgau90OMGjDR15LpKWx7unl
p83FdMvUrOgahWHjLAHkApfAZP0aaBybQzuoFCwjJD9erOtDweuBTqNyDYSTI4buXs4lWdjvIk+6
y0ZLCQQiodyf0+O5l5YWMQ4ancIL56tPxAXhow1TK41LSzzs3BBXE6OKzGbl6vUC0B10wDDEHcI9
qtim2MvIz2wSE0nfYY1jpTfV8WxwgBNOq4+cn2rwF5mm9+pBm2V+eAv01pWgn0ZTqhgwV9COcC2E
wEuIvpQGUxMGzdloKkcFuI2VF83/3XV/Q+oEp/0epLnR04BX+6uC5AZRtATXiKIdf1f8IUpF4lMa
HIhH0kZQmCHzP+EzPIjDYt1MLM6gEwDu2WQRUyn9xzRWoEP0wFxQHbBk2YkrrzB6Ry6EOpc/9u2Z
FV6mbaJNpP66bafCzCZcMzvU6YhdOjH0bIPL4APsTEUrQ4BdpuOMFmujWCjc1sOc1Woav61GH8Y8
kh1eKA3PilSIV9cWV6T6PFBtz1/RGd5u0shYZA1z8IBowtNCCnpXSznmnP9TvTr1Fx2oqQHNEc1u
V15EZyYgZvSFgI9/5xj5+3vJIMlA/WhjYD6qA8BARHydHs7q7l+4g/mFTdXMrJi8DyuAmfvj5Hzr
ThRfKJt9pv7eqZhiDh4xsRGAm0sHRFkAuhH4vZ5yHG4SXAcdsRUecXveDGx2ukf4o9j0Eg5yQ0Ky
OrQsbIEnyvxz2zQOiN6XzBSQNSnU8EepM8jf9Y3F7/VGXByOEaBwL7e3+83bpqoPbHlleYBAYv9N
mC7DMq8CZar36QJ2PZyyskyZUUBrQMSft3lNC7/YebM7JiN+DtbUQSPUgvXdrs2s5S2mT64w0CY3
XhPz/bwE7+TWByiwhv3tuGEjVq6sPl1sGWMXbC2/Ygl9CGkmrevuFjjiKchh9sYmjbq9n1KTAh4M
5KN3RInuWjDpRoRRVoGrd8STvsB+zHwEQhj2bVTkrKx9uayUEe6g2n63tFeJGVt1nhRrmdKg3iM1
xL3/j3ODdzKloL1tJucx018XQqsZhpTtwYvkWp+TdamxDbX347wnvWnX8427Q2DoItdM2vREmqDM
V9nv4kEXQ+TzlvyXGc4HHJBQOBwnf+nRbejYiDGp7JHPDmLE85riuIKWhmnZ0/l32OfyTsige8S2
y3gf11gbNm5V+0cr0+ZhOqkUzHVFm+D9IJp5DScxOk9ZKyEpiCzMqY+pulK3RHTwPDlhZC6ofWhS
z3di0baRDGiEXQQDRLipDALwEcOkq09KJ+O0qPAcUvWB5KNWcRHqkzqmzG2zrDOPj6wU5De8MlCT
iJBERv1YFMoN7Nbqh+jbWcHeHi0bMYkdmB1oQsUoB8wbpxf8+GzVF1fdC8zgUlmBJPoIcbxnjsEN
o6hlkpHzdlIBtf5FfvSqbcTqazLW2T9aXhvy++8xWoLHLVZFCnQcrPkW4OQEh2GREYFPl4cBQIYH
KJbgbn6bNBZgm71PhvaFkML5WjYrNjmPMUeOZcHPbYaL0NSH6T244XlRwRUMRGOKqM2HHYvxuzAb
MVzIoPo7pxe/pd1/BEI9wDOVDlOQOtvjK4K5y59BrSVu9PxLK+zhHcJcwnZwYYpcNP8HVtlAt/9Y
1uro45LcvtwbkHx9G+UmXWZRK8lFoiAzfS4YIY0hpAdpLhyUk69HHqCsxG3hDfRYeWJrTcMciUZT
ku7UVG9GCIYpmnkjW9YlAO3QVnlZVLdLbTjN2Lmorz49o1dIWKynwucVzZ1IK+4N0hKJ+rHA5CJ3
NH81pFaGrAgy1pn3AVz4rVDEX/aHluJI2zwCIhEMoxX6+/QYU3ESSt6yqLPEiVtNaaBX5IimrJqE
EWxjd0x+Q4u+7hjLpE6YHqKKrdjv8Lp+g53irFtRblENOKttZ+xYDvchxv9w+KS+yz3qOc8ANqgb
CYaqI21xn5CwdZDvzpuL1GU29eWwpzlMs6cs1KblO3ifqaS7iVEF0teXKrGsCHOm78L9abGXc4tG
lmvaAczfnRlIKjkGHklfwzeeJRpzfUHI8fIZFaFDJ3h2FP5MjT2Mbo8AhVhhYznItfXL8YxcV5SB
0Hn8SmYDgPcL17hu6x7C1Ru3pYOaQisHd8H4TCYchcWMyzoDHViKkQ6zfuCO1IhdLKnatAxpaZWe
K5c/6CQgHak9woV+1EW7L0OOAXmGdKbvbzwl5utF+HVHef4YJlRY2SBLfZ5Jpu8MJue4cE77gn1R
AhZQq6p44iP5ld5IiMWKgQjo8Y3LAZ4DM8u8fbahzij1fvlVWMsYGADRDLPC3Bw3CWu7ZvIKnkgf
gQOeMJl7/JZYRPgdOY0iTNVvsjZGQkMKT0XwwDIgHtRJAc4A0fIuu3gzlX6v3JUHqI36JvLKMkrG
V0zVQO1plGIDr/iYwWJwAfei04xcomdkaxbVWXJrK9yXIBS2k91KQu7jLNoHBoGYzZielgBj2l1v
nlWyasWGas/kW2WH0mCRnDYTDA2omALmXIirQZMMk3NI8p3Jy36572WQdMaY1reqjI6bIyX5npq3
OyDd/dM1OabCL7ML078CkvQu+m4MGnxVB5x9YNgQbkatS50GYK8xj9aJhz1Fu1ksoBhr/LYFysyA
7AAqXh/UMyNVYhEuiQUCpooVSMOhuR+q0RWKeG4gKC1IUdx1Lv7JS1q4Mpdvr75qQul2UTThPCO3
0ZLQx4qb3SE+4jZbgZQ1472JM4/rLOVSaQ17J0jTOFujTYXDAPPg1awyjQOVTaANZCBA/z6Uhb0Z
D2nYwPKB+iRj+XjbfI7EiZgyy9ygK8ocm1d9e8sJwmf4qoIiZsxsIBq0r/caT+PuZNZmyM4JW7DR
Or6OI9dBjzDFQmi+9SNc68vmXK5IXxFrBL/Fn+pc2QNqDrkKOAo5zN3jx3mSfePZvpmyNQRG2sKT
X6nl27iUJyc71MYcHqSSVWpwEqi49PtlIDcU+kBpwXlEw68zY88wOR3ZJN5HHo6R0TmagjUd7RdC
v8GNQVvMdoAv3c8Viu0V4xvswptINEmqOeP2l4IO60qoAqC+VKtB2lwh8/WqW/TEMJc054R3BItC
6Nraniv87sf2fvR5Eqb4bX6PsKairQnje0QLTUyePco8v7T13XMKKN62KBPeZd/S+z3FypASqQvE
LxUho5PuEb0luZDGhM+LLrFAEcjUaCFHESFb/zG2lqg9+rijvCzsjratYzcoZ4tIcfGi6TRTHnA8
3cUQoqU4Jt9h066tZxxulq6+Fpma94GafWPAKkzKhBZZLujNAlVs4maBfrbsmEpcqwwcz2XuvS+i
o0yBMMnGIUCwVcl9721DLzz3JNKwr9YWONPZUhyAZdY6+B3JCY/ZS5ZVFYSI7jU9eHvvX7Nv4JnD
FtOgSWbozCNppkopaji5uyCZynwQx8eyt7hI3GUnN6H7QJDTgSuVfGOeb+78CbH1a1pHT+0KY0Ua
0MX3xUE9loPb5c3Y8R9EUWksnnKLjNcqh8hgVmil+NcykZ/kUb2S+w+eTDlfkwJzzfIahdQ+ce4j
IdxfP/NJvH+iFq/OB0eNRAEAbLIkMQxF/0SXO5CxqS7kR79BcVxKzT3EqM289PqFTyKHAv+OoZet
OrKhvF9TWCdMS6eW3gSu8xvy5d19E+zImDkCbqRjhdLX9TduIRyC0AHH0WBXhPeOTNaJMXlTNtO1
45e/5Io7mHKcltfHvLcOnB8hCapI50COM8NWjTtTp1z425SmVcvhcKzsnf3yP993Ermk8wI3NeeC
jO5cNhzqNuVv4S6mXIJ49InLpBOaf2dd69LhBaXUnBKDZMSB4ZZXvkx9rZQhtuLpG1W6vZhWl3Fn
kbI8SrCEm/UBYy7fC/7bF4D6eo5mCzO7jVO4ecMeQpfUEYbIvaorrIeTQ29UVpDmerqg2sZL8pI1
wLfO6zIEwpupGz9uhxGIS1a+ISX8gxTf1udMKs2kJvvEx/RektUAGJyRenCYyOUelF2S/SnN2soc
kBU6sdnaIRCoeL6ds0Kxu1RC0sQLLPUZHkSGcGimhduGZuoIAK8Q6H8LHnywRHuakSBvRfF7qjrf
2pbCRdKcbwbYESGj0O89pOUZdti3e1jOaNItLMgx6W4sWGcDQ2EsTf+eFs4GslcEekZym3eUmtK9
V+9PgVr5eH4sBMH4wzIu0qrEocE7XR42CW2o/QdAs0f4w5YqDwuDGQuavCalmyubNtBS0fvO1HW5
2bAeHRHoN2A9PNIkpptjUGXRoihzKJStMsPpVgq93Qu+LVKju9guXgNLs9IgDAvW6Vaxt2I7brMm
78k2SXhhNspRXfAWFgBIxxxv3Wki9zDVs5ALcHgXIIb1HXfjnhlKmHcKlKCjvx7PFzZsJg+bEnu0
mXpan32SCkBU0smQQb5A5nPRC2Q6ltGEZa375fPB4q0z1+J99OCbSq+qITG8JB2lP134b0Pt9ScW
DEENitW6EZkhymgNMHqmTBTAzl0ExSNPlZ6ECRybNK4y06ZG11XH3Ec6O7iOHKCsujvjWRxvtTCr
EM+rv401fd2VBhrPP+ZGweY6HNu5bW196LUuHDA7zv5tZTjyWe3CqSLqDg4K+LDe6w+pUVeN6R/c
9OFbYYHIS6VrjAISV5dJv0K5o7+PFHur1E9r1wYOlKg4w/uhrag7/UkTvZCYzvUK3yo1HY6UCM/R
lumWNabXVOZnimCU0KSN04x2udn4I6tY5VNULdSRC61ANdWx0ovVEqcBSC78kgelDi5lVKWT6Wf/
Gm9bh/CUwaj1OrrYJBJQBQ6Xi1Zfw5RoAZTz1fINFsgVNrdHO4CHdqc0egOv9FhR/gMQ1FY0WzVn
wO03GeMiSEmskmc4eHwB1Qzqx7ln72UC/5ZU2DBDVLr8opq1yJiyG3aQSKPo1E41CaTVMseOEski
YX7m35Hq1249Tg8IEDEXS+2F4u+vUIOoY9oehfAqp5Lk9XdrMsSK9mHD+jCdpbMDVJJCQDJQM86i
rrsul9/VJ43GkPn1KJtZDF7KRamIAM4AV2Hjf6dPJvRSjYCYeSqgovu2S+2qqmMObkxQvH0Ur6j3
b+3gZplu91hZ3owROQpg2gsF7nWdhBfA+C/RVm0bJTjK5GRWFuAx0WICY4f7wUJXlHapCIltGJhR
+1mT/3L3OZC2mqUUwAU1Q/3dsMRS1aMiqxwG+LTvTelRhsHjsYsUWyRv9dfcvTl07yBaYtOTy8fm
UhqveqyOoNyuvYpNqGRUUD04CZO8J9tVHII+buA+tIOpr+CRlxlEhaFxW5/RgoTb8LXqNx72uzDS
duueEgdF/ND68yInS3TexTYy67mlNRWQfoSFusr4oX6lwRYYU6InC1UnThFGUmmU36jHJmzWWE1z
VpxNkSAJRCpdbLpNaatFrqXY+3kdUnytkmh8TcDHhS/HUmnwirM+skJcRWQyGKNn9LuvOsD3bS7C
x1P1Zuc2k528mb1wzxlLMIiXbvM/7sEWZNasSkE/QuhXHsPgXaxQfo8pV7Mwe27vjZN9t4fhDHZf
6UN4KQN5GC7JrTggRR0dvGdWjaZanktcOAWWpyw3wD9pEqEfybZNSnfnn8A7wjF/OcXkXGD5wT23
qsHSiYMXMjHT0dx9Z53qOdl2wkdTseZ4AC01k3v9A0VFx4CCbanxWf+vFSkvQqITl/AqNOQhYzEB
gjQQwr45m3X5q2nim/id8SCD7MlsqYQ05MzdtcgT67ogwq6ZUHb9UGuqaAO75zst1+UB2sa09p3f
lxpKgOeFf91ayZdv4tf7DxMvoyxDW/k686W+acgEB8kLZh1auEXEtJXtRqyoS+UgzShinF5oiHY4
M1XuJYQg0p34wBxfXEe1iIuZ4UZ7pMfVRqbRjnlTJHVhcbtwSPHneU31IOPT+NOPE2SGgd/zfsVX
wwYM5oy5UrWZCEeMNXEJp0Nm7JY0ck1qJJbHxWUZOEcyl+X/eqqcaxA4sHlD6YwMAfaHN8K3PrDX
3cdUtMg0zF3tQpgG62yZdhhCXvE8e8uwmohy8LcQgdZ/KsZqKJVbFhQz82V76souzw93loaPRA4k
EyOVOZdJG54mDRGesvn1XJddP4rL+LwG7AUe8bBCanaFxNEYBOW9mEhUarnIS+k1x9epQEr6V2Fe
y/o1QtQIELLRP67fZU3aFbGCrWH1k/vCDRjbSEEfJMrdvzEqtmkPtSx3TrRMywaUvpzJBHgTNTnt
73OVMBNByKlMrX3ijfmFrING/wUtD3eOJqEu6AcFQUjOqLj7oIaEAQzw5C88ntKNdnk8UGbSrhvH
QH6RHouKoS8CaDZkcS3I+sIHpyHFwQvFb4NMRtniCAYh066GUZtt1R0G0vow+aL1L0tqDvmQ5DHW
3ojNuAWJPUduMlEmPY3eyik3Cy5gp1Rix4P/vE2EuE/Qqu7pZCJJs8niLmVEd4GDvIgA2SAkt06P
eDgBcMnVKD62SChdbdzbM1fmqiPo9Rdb8VshYlRiiE57IYY2lSjDjDFQd0fVko7kApDIUpuRs9AU
5GgteDFu0DeCpxHHttD8V0pWiHg0sQ/hTfgBbRETSBg7FCy3ksnqAH8dx3J/18HvVKkYd5NjWdSB
wa5z3UfGnG8nhduiYa7nzj66VecAwY+d1ByeTTcd6apb5wm1XuS9aZy3Pqop+ZJ0Ko07QeZ1f31H
Qr5MJWj+GA7WwoTIKWCeBsW4DMz3hSNB0vuH+hUkbDGCNnsHpYGN5tpC5yz9tPw1oxw/m/h/4ijI
Xkkpo8DGZA2J/GBMfB+gjpzLo2ZJyJNL6UrZZcP4aDuFMNJzpb3keVWyyWTnLVbd4TacS+FxPMCh
oL2bZVEaBq0t99dKpmQC7D/DMsJhOusq/RnCnin6pXWNBJRFZR7bNxbak6PTTyrvBR1zfXlWnfgR
luQkDNuAPoes1XzvXivDt+fTSos9BNmeXCcgaUqLwtK5XeuYxh6wzGJ+i1AVVCtVNy/cfJwIezj2
KP0jp+i/oURoVl4waoTn7eWhNQDtYydSAem7pHgrUmqfXhruq91SmF6kvD50iHsU1XDi/wwdHx/C
gcj6TvH0zT0tRZqiJ0+9RdCYUux1Y/8bnSQUv+nPe0Ewcr+Z8rioauqg2as0PpFX007sZRuklNX4
PNAwHjz9M26Wj2VNVD777ZMzCpnw4rzXLDNOzbrPueJEYNDR3c44wl8RVocxhwo41Sp04UPj3m5n
1p3Gdx2XTXtcZPUQskBzkMwDzV6pSltkMkjzEpOXNl2ReqC2x6HAMDGxETsXoGCvOYoWKUS/4H2r
/sBRdxcWfqzyZ476dDhJoxNuPaX4l/snTagNqYkOetIHUd/DVoys72WQQZFH87PsmHXGtA2qlXVX
QCnNQz4BcwvW3Sw/3bfh80Mlb2yTzi9uUoWkdCsgtIDEFQ4JjYeBJE3TQXWtmyNq/xusdU5HfOXK
vt7euIke5aiLbS7a1nqTVFhCkroj2xw8R/M7HExdEag90tJOqE4ibHqit3Q2q75N7AGr1zjHMR+G
0b6f+NVHaRQEQfVyJQT6WPWGLIFZeI1b3e/korECBbjBzo3J4/c5gkOFoQoTX7ZKxH9yrHprZezI
2x+EDEIPH7WSSVwcB95y8ZhNm1CUgsE48ZGx50C1KGlgF5I7awxabX99poZLlkbEsQu+h1xhgYfp
5Q2Ylw3ckCo3yC3skCZqZuEKTmvDn0vPzC3hdfAGNhUpaHxinjEdhCmdsflR4J3LGGI4W3EyD3Ps
we5fW+32SUs0xI6KM4bTjJfPvr/4A+rLxCEkUavc515sAwW5MK33YjPjrivictX8rFi6suEZBU7m
g0Gwd+c4nPzVYZeMF8VJkiAeaxp1BwqJYekmVW8sJ3QD2m7naLS07hGprx5k9m8bsPlFZchfOHPC
B9rEK8k0rAgg8LyFhPr3OuNLPxYZLlujXkmayTKDIj2IgI9jgGKi/O+nz81raRkf4N1INhGyTywf
6r8z1S2HGofIwGGdVdG8uve3qElkSbtlAiVLeVcIkYggC3QoLrgYYAlAjKoT3eAZwRk4W9Fx72iW
/C+NVd479+uXQq2oFhfnmEh2oRymOzgm58pdwLxi2FnD3pWvoorFTX6abDV/z5mtWdo7d6avP96Z
EbohQHmiuFU2pUcxWK9ZRo23R8hQA/6ZNPQ6xzLUBnswa3HDVqkGnWZF29bl+dHkHcEnC7HgGl5Q
UvIruB+vMKgOCA2Fgc3MsgsmhfI2QTVf4S7Y7lBeahRl3vDF52mDHo6006sAHxp5Z4fz7N8pfFFj
4HKuK18cABnJVK6AymXp/X5AfLenBqs1nGQ1OuHJIpBXp7vhnJXOxNUHKTmb+8IO2GyCirNxnpAY
+yRd3uA48jcd7PUhml7hp4hJ0pPu2Hp0TxzIeX3+axozPkr5Tlkl2LUWIFSWgagKB7ItKzFoSS2X
k8C8D7x7023ipF1ZGytnaDznzPYTiMtp+ycUTj+dwTR2gpVH6juvTOg+xQvU/NHyrB2JtaCJtUxx
ekr1htoGplAmuRACVNwjhBevdJaRsdhPjvGxXL9WTmQXJ8hCqw0VzTDXRXAKDp63K8a3GY94kABf
UeIAdEwAi5cq6wBqKi0zIP15T2p7sZN/Su5wbVVUkW+XsYMNbuEaVOvxXD5eyzBe3JJ+biGxdyGm
6SZpO3ME06nelwAf2Ii6jRpMfEImnappa4SjKC6vDMKvDwfRGk7bvnmyTBvD0TlO/gA6r0vWoWls
ICp1VL2nD4YiBSwMgteSpAPHp+eqkcBzCoxH2kZXJryD9nqO/7qmVP5YAh7XEtYLNNqA99FJPbnH
yDHG5ecen3cumsiEjDWktF0m+itjCKNqXNy1NRzMveUXZtIDk0iOESmdK3ZRAqkvqKrGVXuQgJBO
vVkB02MKe43xXpHZKnCeexSM1+ql+gouFf+P+H7Y7J9kd433gk2OR/9JB1SuFpmAEzvYH5H8Du45
0NHEvQrXsMr6gQDxDs84KE5XY1+YfER3rIsI5mB0W/Rvbfk+gS7S4AkeZLbOuHcRZxEQZ7v//kH0
xURmHWfj6vH0HoKWh5e+7Jd1qq0Fia1y4ibOm/+9feh9vin6ajb2TuKRdFpMTD7VAosR8kB6o25i
7hUX2l5iHNcIhfofpKjqqm3mWMakubAQHMj9B5kdRpDx4WYlJ2ZvfY8CvJerdWUbC6sO5QFCvGp5
tpCjUd1EwVzhIudldEAcORqHkaGTP3Dq8c2PhxKHwuVw55k/GHujLW/8cBY5Lmy1ZYH6JB1fIFvW
rsYY78jkaItzbdnlc86gFV2trMEcIoI6ouh+vuzjyBE+mn6TdOUHWMw9ZAK86tqZw9RUCuiAuvXt
R99yT4tkbZUqLXMafC/+tnbOwoBx9yrovUYbtfkzC/1G7uxWXXkBEfrgLwXcXJkt38SrA1/DYM62
5lGdLdSmb4zBbv2KYckr/x2VVsM9rdUDqlkErnHrGIgB64gNzls588Af8HjP5uiRQ5Ut7oACLbtn
BoGUunm4g5io0IcGdyrAhAIKwShq8zXzNdzSQjNKr8c1o45FKioNBKa0EK3duGXQ+zWPTVuvhY6p
2C+KYQIeRwAUAR+ARTY+hvKCiy+FCfoA/Vbp/WR39tblgg/b1vjZdUHE7J4pkoT1jOrHAQPb7Pnl
z5oOr4QQ2996vxEQY53viyGCA7YNM/YO1xxPup57mNqDuTLKYL49ksenSnQFwWtxVGYUwDeZ2+UB
koOBT95nYUiNhNt9EZtnfBYfDdZIUQEaOVZw+m8Uab7m9CZJC1Efmf+P5jMOULwyxQjbLjGNUEAw
lyjotukQodzmnK1tyK/xVmc7m5Hq776mWIM5tmWTzQSItL468SsxN43SouVkvO7ul1fCLlKexFCi
KYHWF2zCV4OJBeuqYNbDYEJi2JL/4nF78WZYVR3KoNvOg3poPYxQc5mNv0SEgaQe6H5FI118Fzfb
2MYmsuKy8bMqGp6XS2fLFpmVS3sOhWFBcfKfCM/Yg4+hntFKQNjKLbG73tZx1Veb1sHfg23sIBQM
jmp3XIcjz0erSZc69MSYMvDzHd99zSPuZI+EQP3Ii7bf6EPMzYCzNiNV9Lwh1/ZDNjMy2zSC7h1y
h/iLnJrn/NpftoztdoW9i31qxnrU7GsvVWkofAOqxFokx+6ufcTKftODscRahTBNtl6IWv+xN1PC
oBxIwQREVjZOsuP6yLWpLIocSgsDOII51ZZbvxsuIcu3d4RWAtOsmK+KDk5sv2CN4aSOCd1w2R/a
QuHY3NcInDvqZkabOST6nyGqrdBZxQuvfYCmU0AnJBpSkJibAgwJt/ebkKpEuoCa/NEeD5bw1CG7
EQhqO/GvgZK2ULOwo2VbxvDB5y4xWlr8HtM7VS+/HcFITBbcalmvFnADsDlThaexJTQnLdEyXOnr
/RjgzdD6cJ0pug02UVdy8I5gthEZoPDZbYAE0Jfgp8u5pfFetS7H9G7hudgrBTapva06rSQMBBwH
ZYORIovji23lo/BGGzi/xB92hwAVe3b5gt6JWOrtCKQbqrCg1RXz3snghKm1e39a4trvUROK3VUE
Bzi9FiInxDl/sazRKl9m/wJ4OSF1glysRP7WQg+S4a4aucCYCyZV1PNuGFkJOXGkFtYXhJDxnVwe
di7lF1f+KDDqZC6pdUAH6RnutjBZ0q09DtCLuiQrviHTtF7qmAZ5nujGawxk7uuMxrW6jpBshNTF
3jD+0hYaubFk8YEYAU8ZKxcabj+AEX3gOKBMbzCFTiSZ8WSjcG4MrbEt+N8mjftHE455CJH/w5rk
LHtIPy+T9gaorldnRAXPzptKeEv61DAumOcPyuz2AESiCUEW6kXvVHCongJ0CojhEK5AgUF2Nusv
fc36SCgYhaYeIwN8tIzdAt/5p+cKFJZxc41P1YMB+Q4N5HapuLjbnDWYH7dcEsVYKS8aFDN3gosF
gulsQv12MyOgDEiFIuWK9sWt7MxL07wAfXMKjxtj2Oun5j34vYnlxQCq4GpsnGultaLa+ldZc+8X
x6reQC8zMvMZQ37QKdNE4GaqJFn9NPyvoKd+Se0QQ38NLgYOcBqkas1BcWp3I9Qx1pg2r8zRfdec
n1Y3YdWNRVcrCaIeYxSfULXkorqiJwropScPKugvpRBOLuIypGfMO9svLfcOGRGxHIo3l72A7r0I
7xjiBwzWF4KzjMFuobNB7aRNd9pw2J7Ec9X7V20yV3ji3515yUGJ66T0hJj/9EgPMiJjubwbxnZB
IYoElGvmu9oN2jlohTx0hhXBseAlggUMOFSCvwzqAI+0ky4z/XeVOGubacAYfsHbSKpX4n/h/JY7
vsrCZx0OrTAylEHz8Q6fJqwwl6OsTmOkXQ1/QkbvwP7ueqdfpIbr0U39rba+H81mSGW5c1Q0UJD4
jWt0QxjtgE8elo/iuUeaUk7fPWT0dc6Uenk05dsDIAMC0Cc66kJvuNs59jszih30Yh2lWfpG7c6Z
nDb6APFoOSR45GYBtapeSE0vWxLNIUsV5UnB2phuYcJqPpJ/RpcuzCUxbqkKalkAaHaz+hffhOtK
DaQ86kgcZjt0l4UibY3xawztq0jdLgrNA/acfBZ2dH4qUA43Xwz74w71JFIpAvRzSL36+yT9rXfk
60kI4eoieYgohug9iC/c2FxC1f/728fYuiDbgdS0adJIdJrWZru9gjvsHlcQiyNQXSjUY1kHpNN7
j5dv50v2OqxMFT/FqynH2ag4mEhVaghTMr4PJ5Geyok0eZ9jBGKzIXjW3z+KTuKCiOvG/wUdztVU
IgXkCSbVWfNCrsaixasK0PpPdkkfp/5BBe6zd6vj3qx/LxGJGh1BOEh6nuFaOdwZzZUlLVCLqk98
QXkxeEx4u2yDuEj1KjIo+GwTCUdjRfhUxEJIU/zuhx73Nc2ZNKxJ12szOmsKhDLS0C3fgL3aZ7jA
vxSaNvzoUzJjMW70wrUKtI9QbEb/CsqKU7V3OH72tXRuBxSt4EGnMqRogkaRarWCp0Pe4BNZmSvQ
tjfUgAUWYF98nBSi9KRAUOB/iayR9/oE3vNE4VDsCU/ICWpmZeIatlixCfReAQsc0oTDKFkMw7+k
j6v5QGwP+s2NXb1Kqdrrv9q+PTrmNKTWfP819ftR6MIdHVAgUMyFjW2PRtswpkC4/qiTATi4qsUO
XjHCcEOeGFO8qIbrYvqD/xgigiJ2R69rEe9lSyQfcXP4H6z9zLhcctWLUH6xGFgPz33Qg1dPJekv
8i8QmwX937Wpt/XADJDNvFUB68gT8c1A2ENnEseebKkvlsbHUP3qjok2AdHu6E5qYsz2G2MVG5ow
805JCBIiphmS/PAtAN9HAvdhaZjcRL3yOvA8djNrE+kR0sz30BYjzYf8IsIhpWd4g/+wOvVGzkFf
IlDPC9pDRJALdLFX1jaAq6VAFPQXGzGCG9KZJDEx6CALF+76mAl6A00VAo8O6rksgfDaaHTqUKwM
ySL1yMVN8RXRgjh3WW2AoolLX5vvGT7FvXoilITY2n1HPon60kTcy3BbCAoshFtXKn9a9c+gVyMx
8tLOT1xoEUNz2+wTdXDOjTbP1AfpeogM5BMa5xTTJdk4lvNmthYOt7KjZpQNfLl+CQ24L7o5e+Fs
zQl97rvpnbX9aBuEVUhUuI0gM/yWYqp2RaEE+lrXzH7omkNxi80tDcImB3Z7Tg3poO/mq4UC4MOL
eeRkxcnPmiowC2Jd+ENfBsuhcU7xSn7QdnpFGI4vhBhF3R8edOXHt84Ubh1BlhjrzhLSK5p7TLF3
lTugiqlg8KIJQJAmzTqcdzX0K6UIuzHm2CmsTvoaJL0nGc/QmlklePKHNnbuL0r8wq8D+Gn7J3It
eX5FvCTMQPQzLSkATdBJYUw6h0Ryj7/stXqq+Sg7RY1n6rSGi3XIHi0RBoPPW0ql+AO5Ye4sMiwV
UHHcCzlNzNH4oh6KtZQhhv5B7KLkd6vnr1MVjHgOSy5wZSUB4HrchbOS/ykJXOrza7Eqypflb3PU
/QFVEoaiX+hLEf+Fr6esl6OENihHdsIxJIa4IH5R3JYErAO7VXk/vjIr/hi61j+D35gl8vF//iqB
yANeiVtBf/Cu+5TOOlNMX0ve7V70j5ltG9QkrlOmp5eDH7h1tJDg4sbpoLkFXtF2QRg5FPzM/3um
MyWzur9YQpAy7yHS4kxsvTh18Vwvh/57zk23wkv1fiIftlOeNfP1WBeiFesDU2W2P6oVFoic/zGz
SFMwhb8VCpQZg1RFVDHinE148hheiq4Gr6CV/8cR+d11fVl1MSGuX5Vpk728+h/AnFgA5RyIk5Lg
3IBkl7IMlKARUjxGGrFuzmhzWP16Oo35LF5RIRIWMlM/iFWViFwaUktokCHKc9uey4jX6MQCb/7L
tG85CKDXaEKByd8C/UzdGRIX7xcYEipT4LK+TccmUYqgTw0mY9Xrhl5WdQVtcn/wJKvpPlIK/azB
Ug4ovsw66cVUT7riPlpyd1mb+J/dwXJ+NY1FKRarXJ/aahCb4ioxpXpsJOxqjxX04JPfa9f/GEkh
UB58uU0FAK6s48ljFg1psc9DlhNlYXdbqgHNNeTZoVh2zAH94IW58bWHdX9ymAhVsshLS/zTmPEt
qsnhr2b0k+1L+GHhOvSNLH9ajIkjp+CV8nei7AONfdj4xETGk9B1fD9FA0wRmNXFhSZ5BdkNVxg/
OfV4fqx4xg0+kFz2cj/ve0Kt0r0JHgiDEPSp1uUfTEyjKO10Z8a6PUfxj1j+ENhYrdiQtM+52FOo
5nATFqdjgiLaREuokHHljhj5z95iUiE1JApEjXaO71eINMT87/2J82r85+ZiCYjstybGCZPjluTq
m8xn/+J4bn/rRhwLHZDAZ4MAY9JrwIeabvLdUk+Z8xqjbkqhviCPWm4yBj+QvzY3JLLpVVY7aNAR
fTTZRT/jqehzD771QyKBySjOc/MP9A1uA4/+p21xvq7w1kuGo9sQqj7vmf+6BqxiAo68YZMlXwX5
YMVxjoaT0qyldSObGCd8D2VW7RobQw9VDPZrF5wMHHYD+r6I6wPuatcB0ZcTLtGVsHG2VrPOL6Uz
zDdVVusZ16qJDIg5cEnQA8TKCY++78XUoFvp3vOG8elR3Adx11YXvD9U5pNEoBIpSPSxXd19+GS2
IKlnzTBITLhvK9k47B4SK38NpZz3ZURF6PeDBLZZHbz944gLR1zO63T3EHxdC2efrSyUZaDNEU8S
cWRvlvqSa49j5XbmC3DG6a1/foUFDv1S4hFYkuIGTuSAurjcyVg5aPnOAXnmtSgVtuDe2P3rjrZB
UnhJLin7sW8rWFQ+fseG2o7+u2u53kiC/2KHgJmxKOS4Iw+WNrJYXvUM5m0oN7HEAiJjFWleu6um
GDPL9I6PwUZQNE0KrHC7X1o9U3Yhdo2HrNJrK+Q0qaH9opCzqiEFpbCDu8OvprGSKDGjN+7eYkgI
Y4FOAw164CHYqjZF3UNvs8Qab8h46H+o3XlqITUVDbv64EiZXM69aKh+Q1OuoDQp+mp4hsc56QmS
9/FYgHUlmHu4QZuj6BsG7UmuigcmhaOFbF8s0T3fb2UbjcBohwiJ6Xvqyx+u6plCkUwxytKHI+p7
4EDeM37ujhM4l9PRFqrjGsCQoYsoDxW7vltvYqpkqI7cJLtKvvnYLo46Pv5gy2JEpByZc+bIAVkW
4aOOQ3wlmIVlnBuRv0Z0ov7fpTyS44XtaKj8QzPz0ZuEggmSx7i5FgqjFN9S+uIZIgRBve9gFOeB
qRPXlwKA3JGCOYLlZsIAi/fwzLcjREp39ETHvraXLyBaSJVNuLB12/sPtK9iy0c1iJqkYuZtvioM
/Gih0SXNzcGj5Z3vWqU6SfYbDTN5MkLmrOluNamVi2/u+rgBb7V4Ghv+QwD51/PWvnsTedQYS+v1
xNl5eOBcRkHMygGboj6F7XPeBoy77RbJpau8gTdK1y2lcS9jf+o0oj+Tzt0+rju2W3F7JlllBaUO
o1OHhgAY/1KZ0Werl5aSyPdnjS6qQceIDdb12BX6dHetsv6wnEeoglhIlYtr5QFFO/+mCQo5PN8R
pkQDFHGbxLjlLVkTm+VXi1gMZdNFV/ySwLxER0BW5xAEXs6QK/U6fTRNl7riW0i/jtU/wLAnho68
ojPnwvVtKPq8JhEEyw+kVeoRTnkGNdFKIyL3sLOpOxnZWMhNFkN9F4EKUSG/8NuPSuAKJwk1Hyfi
/HzA0IpKoqFfpbBgIAs6+QrYIFBoguTmhb730QSNGjcZnSzv9P2YFJ8iW+W5+s6iljUZG28ZZ7Pt
amATekvD30b2QQwZsXzfeh2uUlFcqGPMinfWexf85SLkPXnHgJa/zqApLjI+co/Ed4L3yUnT/oBQ
F0JjhlMLrVmxeHgkcHnklK4jC3kJYNdKFrlSZLdIR+0xy09dqZFT/T+ju2ASidLSC+XJLpsjorey
2pwh3ROyOktx3NuDq6ioTucWQwHHAL9aEV30GCHWJj2CgHBVxStBiO02+SgReFJw0lb57gqPN8r+
TBxowgR93M0AKoWVu05q3/M/WkoND3ns2sGA27QrXHgEjIjbveftS6igkSov1dHwVszZ+i1rfM4C
W+ZnCXn5dpZwvDx3YdT1mNYFs2uBo7+0N0fLNyAxVljPdGDx+Yoqn/oaXXdiktwzsZme8vFt+8QQ
/bJr6U6B8MWtruWTOAuswhcQT8P+ztxSwRD7dDqB5zuJZKosijhHDXBJ8aFrzoONVd/n34Usvp2T
XOmL3stTSiRecfo39C5INAHmzQfMavo3swPXw+67Xzc3kqBFyTxBJ0AoIaZO/PQHIJNIOENne2IK
zJRyEkCVjcbGTmgxjkoTtMwdimVW1LEPvTgog4kq7UGLOyaz31YGyCxnrUxlqoKgoWySirY65sdP
jS0EFNO5yAEL1nkgKc4ZP1NPhjvuLcPBT5U8C4p3QA66RrCFc1MCjhU3wYt7Qe+ZsMAFayr9TiZc
ux/EtEUaojwuHci+0Eo7druRD1vlyjwbX+/FIakweLSlZSmgp7izz301SeZhVRL2VLdIgyi/q7sy
M6ePsRVcvkRsKzgcArg/2KNT4dNTZFwk1wsHuYqychd8uWgh2OwWQXxR96kNeaW2Q+aSGbK4ks1p
Cdjxkrn9mi5ZPxQ/WIf5Fo+6CjDF2uf0Lp96IbRqLLxLZKL1uwuNAm9/r0Jg+9vvUpaRkqCuPdNh
DKx0lf9+5/dyq7GntDo+2XASpAn2UYu1ppRTO+fyl2hIhHFpJrpy5d4A6p/afHojruL3AbpR3HP6
4qsesigd5CGQEMqjYLdsdWF0cqegKAM14bowfCzJfZj0aukU6XeBJs6Z9Jt/U1/qrSDKubSnvXL+
eUBRwDzYM0avC6/UE+wApcH5mtsOhyJqRz+wFG2J74g5SiSTjG8HQLTWjUlaxwrkfaVr0qsvrEZV
kiLOaOjZsM1zOXaPD5dm9CBRTQpvOlIS8u0+bk2dLMQAwU7vFE76JpEfnxFDvlwg/xfuyEIPIImF
1tR7GHO3PVl3NrCSZcU6HafjycltYh0tx9GiQzuFzX+51lbq9bgU6l7zfaacNKi2YAbBlgPpMDdu
WqTYyvRNvni6j70UZLjgw+Dl0ctZg1rtSUvI1K4u7liJrt5Jb0PaoBw2D9cHZ1d1zgoBHgpcA/PA
m6AI8nu2n4T+s7PuY6j6z9LeP9iv7Ic4B8j2W4RaasWcTrgqxh83fek+LCN7D61wbm0nyyew81hX
mfaOk1xBZ41CGkvP5MXNB0/GVzbSaoVZDtOBV6MvzegBJUyXWtI2oJ2c1UZSiRE7xQNXEa5iNrpJ
rPrUu+RNRwj4bJxZURKVz7CBZF6dySNMH3/S8yAmggagmByUd++VX7CDLgjWJho6nK1pbMLvWfiu
sdS1CthSCv5X5BFa0DZnkiu4RMM2tTdZGFGF7tiQg0gfagYJS+VlaIybFBvZzK7xZiKHNhUPgCmi
9lmakSdEImmtjQwnsWYHEW6xelk/eZF/KLkQzSOnbhOigWtyJze9Ja08BKihy32IgFhQ1e5AUaF9
XXWAI/+NkD4FoAQbTn0orGQXMvJwzqKZ4YDpLw3dqBg2IpBTv4f9wDcISAmF9FNZzkmQ70vfE38a
jQ6j1EtQCLVMQ4bEOLq4pPEehM4NUBkNbwuzhMVby9QYXYDuhOe7jnA90jZCLK2JrFFeNUNqQxMN
hxB4FfgyRrN74yF2k9ZSqyjrr/K0+axKz65piQ5MgT0CZuoLMdPZPZg7m7HMy9rYsA7+5/X7GjYm
6g8k9EvREl6F0Bqb23hXb56lhX2fydBgW+qvNlsvskYZM4dQAD2Dm1TAc3IdJe1WzffzkRmQFm7b
BCi0jv7aH6zjO/z+smwiMI5650PsiARy4l84Wt2E8BdLeMTbltF085FOLW1woOZsJW+PGq4p/SPK
4zClvuDH8kGITcebH6hXh3v+wbxN2PupVjFQY/OilMT+0kvKpJjOIBIiSStGqTG5gJCWsNcyn4qU
DxBLu2RFc7wcK5cUZzE7E/NmlMsMjfXiv9iLnT3uObVQOgAlAP4cmsjKCKWCUtUvy7pN9JjNO0yq
+3QHV+1wIQH72X6Fqhb3jCzLFRaLox0Jj1jr4CVjjy5jPmqFKOMbQEhWSlFpeddtogdW1LmFjXPL
/5AcX3+hMtQK+OKHJC9ylyT+jntp1h+4wmkn5QDFaagDGAXhgThSWZmA+IfiQWebYErHN8VlZDqe
iLUpb30pBHiMSwqeVDvyFbRxfN3JreZr+LYKBrCCUxi4lVcLpVQf0DXFMTEoVPb71V/9P5YV0Yas
CrUHRKUjdjX3atLHlZPDz/xuO2w/hrhiDhpkU/h1zy3Rr9UytFU/8YAHEMmsa+08IMZ/ItQwNyBV
9bUsA0pcQK6i2ezvPYq6J5G5hjNpTcZGvEH5XbMepfLjD7tFfrkFNBq2mrRrdDYw+TxVQCDaJ6eq
D0dPytvSEsuynOaAxx6JIytbajCVAGI1+k62vpFJvZ7jYmUNqQioB1cQI2XAh4mofaQpj8iQBL3b
voSr4GlqV9kFBdndu9zc6sNCCB1F9hcHMfMpH17jc1ZD4WKcHRvAxsQlmftEnWQbQCV4m+xdbQys
qqk4rAMvt9kmhwHMs6iPqMxgO5uSlE3IvzJSY4sNbyV54STvXZKPhNlwy0gS0cmK0dsLaFmijzch
r0TkGhRzHe9XP/+OwkK+Ujei8yz9PGIcURJEMRKW4Y14vRoIJ9lQKRekdJAld3WuUFyHCgHQdPNX
s2sjOVva4rSw1LJagUuDgIuiRVlikJSL1wUb3jvA+gG8aWdC3LZA0KJ9RHvcez0gZtpdV7uqZ343
zQBAtiaqiZ4gcFXu4o/QPcl3Rfvwct/XjmwssJCL0gDjnSFwj3SjgBKGoxSUzs7zHtlYIhSpnoZK
q24qPuqj3mueKgcslDmljifYovxz0DvtBtKhEeawUfUIKtODIRo3vibexv93CKpgN1akew4aJPLw
LV6fjcdM4UwUXirqHJCEj0py1+JzKFXaMm4/hs2NMQ2jEjJDy8Lbk4I8gwJ1LkwsGIhlWPltXbjm
Ux611dnUyAR7qwvgC7gzN06gXXGOsHjreTJEYba01J1hZqsnMygwQDeDfZh9KGIYAVg2dUhSATBu
9gOuw8qTofWkIgPytbdbISSHcJUQ52iKFc5AtOIB8D/KGq1Xraa8C+CbjiyvdqF4iTXqvFoEuaoL
EWDY8BKE5lCyphy6iQoORnEBH7XniJjFzpsSTnrj/uxZjs8cWNBIHE8CBNm5k1Po7WVvBnZNi10T
E7LFKrb3+xiSLqjD7O0OMzHbzzY7/GziwXaNvvZZoMP3drjCo1QgTIU2N0yhemBq+sVeSa9lPYoZ
wu29rfLf0gJd3bwAoWq5IMO0I/tdl78/BzIhAuJGvQZwoqRAju/FXVEUppJkUa3+2DBPEVjYAHT7
JGcT+tn4kPR89OQMIIvWdmiKgrLecRkPIwIrZgFQgDSfngOTU/DRDmqKAgldlbJ9+mVS4BFuEDWI
QxSTNK0UvdqKepi69lpMxiJnibKiwmvwW7+AwijJHEaN9bITghgMkqabJ0QQ+sZYtYh8FiuypaNw
vkE3CzU8Jy+y+icd6fU3u2Co7YJZEoC/VHCYBDlb0YO/DWAg4zWhGtC3LHxNPTD2eBWnFEcFbyS3
C8tFo+Qi/+VbArkLp1j9UrtRTnd5JZyvIM2JunoGXujHZopUyrFCeJExHBlNRMAZKAS6kLHAtb1Q
KCkqQg7tsW9KLHlwZOAdxkopXRuyMGVKAeHvEPW1HqWKqVKup2d3get0brqMMOhI8mEkcdCVjtxR
HUxpsZd230liK1r52h9HV86StOudZA4RudjqvjEYxe50kbkStnngAsTMykXTHl16VImEyr1w/CU+
/wvzOofsEyfYH9a621ZyGvlmcoCG5xMsBeE4s2ON+8P3wEzDKWFxqvInRZHBa3gl5iZ4D3XGgYS/
/kEET6a3tfDs8+N+EtqvhhnIBbjzZ7q1+2h1YI18cJw3m2MyPQtOZZPAymLs/8L/d+Sxz0Zvrmip
Y7ha/jGrYkHWz/djlbDI4nqX0I0+r3238vbuzAPknSWMKskGtGsJnMHv10GvEyZ/uXF8VrVNSUWs
2e7yH8vMpMV4jcpIwd67uYGpl+5sdRFCTy0irLk244kBxce5hgtoUsXh/kk1Iy8wdpkSrOkfsDCM
BseS/NYz1mx6lhOMkbavjzEOdbO4yciwwZTd3hp+QLcXlsPXryP61EkPo6ZA98dG6L6z46fFvuuW
FcWJ6WoYs7vKV9dQLKPznoLzQyZwSYv/N0Kn4W1xxqdpEl8sirFYFv+jDbZN2C6m7mDYT62D2YmX
xDBx0Q77aXVHsYdO76AQNx5dpYwFO+DOoLTtQjp9qa8Uv3AYFoQiGw16Jc5vs1RtVOzVnSuXVN5d
98BmVrt28c5weGV/9R/IftibGXT35tAnL/H2xhUD5+Yr1rv+myVdj204sbn60fxPQUktZE21YzLE
vydF4cyEVJEuZ2RE2F9VCV7zRcybM6EH4lczfH2scRj85mn3RItp4CouQG7SsLytVOOKkemy7iHb
ZtKTJ8qkUNZioPhHwyi+utdQzDmS+wwOvhfMQtIoYBcemD02PYhLkDDCplXpwjTVo4BuRGt5u0kV
Nwo7v2P6v/O4lHrUg7yBao2G4vTA0rDtfJ/Kp3OFGbJA+r5NXCf1cv3V8V/SSS04xqhS0iiG9xVm
ZuUTv7eM5H/phhXgdwqZ4tEde4R20P8leC+RwHPYu8Pe5lkudZsaorIB1lYwFzQIxNSiwiKIkIY0
AH4WNv2JpKUQOOC6U5sxaoI7h1m7zdoSGx5MOe5CKtsJ/43seW2uZ6mxll/TPJzsHapjwNwpBZsX
18JOPGcZqeEIFKrGGyy8lRldxu5Hbqv32APxh/qqcaRp0aFxgVncw5VR4tWslFwHPp9jY2IB8vmt
0m8rSZQV3/YLg9O6C4e3o2JneaZYSXeKqPfx68SNP5ZGTEuh/G3UBq7P34DU/0HWSYveiXB5AVat
9hApXrKOXjaqvrORALTW8p+gobPwCA9MS/1YY3RNhlEO/TRPPywjoNwDMe0wwPOS0CFB2s+SQJLJ
s0ncO3LNssSN8t3b8jYf3LVUqXokGVdEJcYJUNtZk74Cdh+FK5HG8qPNNxBdoRPYClpAV2GU7tcV
EHeyu2g/2DVBmUNb91ouF1rWLGuJFLB/+dXELzliw3JDSJsaKU0Sx1fQkr7JhO0PgPSscfT0yWmo
Ebs/X0H0+2quqFMRbVnyjYAqbKFCYvv5Gz0GA+dreTOnaCUwOfTly9WUL2Ealnp8Q54GpoyfbGK6
SMMJd6KF9LcWUBOvq4GkkuWouRqcXUCg4Zgcdk4uo8OvrpN0cn50OYK9DTU7T5jKS9bNlVHyvJJR
/gzmUvspIfGzA5Afizdp5gQJuy6bhvp2EPugLaKBVHhJ0+QX7VxbzcF5XZUUtMTYzECCrBPLr0wi
FpxUFt9lsWMFOYRM69I+pL5LE/oUUyT3dBeYvQRBPNCC4O4I1D0b64wSlQkesSTAeC4BZqJd3M5o
rbUTAVnrs2zbTBO2FWT7gXUq+xsWDb+hq83A1RSQ0nhbGSbDtSawlTV0aMl6nrs+0/fqlAVBHV6J
G3RjfVXGnr/QRZb2tMPrwiJk5u3wP2Gr76gLebUEqelu+4e/YN6jiOVurnVDk1Ul3maPn2r82e6Q
IURFSA614TDDtOiz5a2evxp+QYvR0ARcEWTx3BCfGrnk/SV/es+bVpfMvae5yK/poOJTnWUBHYd8
N5mrBJsULWEVqqbpjdkAbDNSY4/Rx/q/IW9gdiXf5SaOWKOtZPZtO7Cgh/8uYMe7AOtVXAcki4DO
IrMjUZgEeBmooLZtllYavBAJ9cFLDRg6Pa3cGJ+pfpgVD1pxsQiJFbXsekpDnKin1jtPjWqVo7/l
hRTl1zrTjmj1RtKLajTjmCAbb4vyIlcX76IGR/z0z4g4/nmR4RyiDPyu/01NfLX1SsQz8qmLxZUj
+Eb5o+ljHsQpo+UeioT6BqMBWknA61FvukCQa8LburDSE57F3g9g0M5NkGFejuk/2cOpyGoBvVTm
hHaeLyB86VGSLyAkosV+hKqgXIqRzWTde2mv2/LiQ5sqtBbQvrjP3tv2xvrAG/naTjJ5GMdu9+Nh
8NED1yE+EJsMcje7Xcicl4Ai3z8o4AUObdJ8FPfjUikqmNtmK0Z3R+vGqbGNy43xJ04PvoHstjC2
3sFVB9A1EeZoZa/Rr2sbDt2t1qtVQN5w+R1Ha2JLbFlEZiapbmv01Y5hmGHAR7fCX13yAVrA2auK
22IuPuCDh7qLJT0vdqKiceD44Dnzh1+C0X/lkaKTjCvltlahAAAdI1Fkgv1vPoMVs1d5cEluTvkn
BFi/bwA+2zKbC368kHwKpg5WjP1nq84tsILbrnlAEqbfgM8scDiDD1kYZijReKw3nRt07xzbrPBt
/5aeBFrvaillK+O9coZVJ/hdPSzoNlh5KH/g6X5Ienmx43i2b1PavdUxEhYfIiyfoLkRBlRG5x1l
cZ5bI/qfPUTMyK3RMnrLOf4mgMU09XoR4zhVe49CUH/N9iofpauUSO+iycNArhbjwFG5Yu3vlrbW
IK6PKtqTMPLJdvVbwd5kBamNrFUwuxEXX/iuJ3e85RImeLLjSLNUS6zIx08eaOHoYM/uUnbw6JvE
B4EI3WAf+x/ZXc5ac8wIThYS8GOIj/hzR7SF7UURs7on9uiR8z4PCgoeI/srxj2xvRE84l1ctyS2
HZ2YfrTDgZE5/aB/yF5lz8E6zpcHwBcDT7ScoHl5jXvOzULO2oQM5rLv8ymB65fa39SoPhEEkuvs
Id2NqJucTdm9jrh6q0rX3CLyGGi5cHAEis3rjA9wvV8yb7ShoGULj8OeFhHXY7LNdYfsseqK9eMp
LUGnnAXRUdT85bwH8IByz4xFHpfZWZMPxs5lJwmcUs9BHBJD9OUd5bSsEV3HayBc75F995IaBYWv
o/6zF5+1pCZLi54wKjV4+NIR+UDkxtmxTNc3Cz5QLM7tlWKVYpGd8L5ZM5EroGdPhsBJBTQxlfXE
oLNknInJgZxEI/+URQkZ7nCQzBVr9J/nG7NvQKIQRHeLqjCZyHZUSx3QuSDUrqycee7ZCbXUrheX
45TEZ8l2DQT6i78jJvM0EYz7jFCQDKEIoZh6dr+xn5knpEZs2kyITI5fyGGTXbITEeoxk+VGDV3v
XYLHbyd7J4h6rk5MFdX/wPrfmEPORhvi525eqJeUcqbHqI+yVwXVNB2tfOipxs8NqRP5xdTq+zzQ
Z+Qzd5RR4HZT6QXL4/7nyQZYneTE0QwtEqx20lvzVBYZqRkuBKr7TWT5Yrh5lb688tyF9akA/IMl
/A8PjyG1/bHgDy4nVr7tdmpE+YEbXFZXL+mxBdqvm1Ta4tyrHHdswB5hFsNnKeWol6dniKYBGe8x
IcF6bQTOJuAeJISB/sgzwUy9dtM7mbN2yT+48rA2Diurc6mxmoAb+l2p+VQk9/s66VEPqWo7yYEQ
LY2keMoLTN3ACLKPzNfCtF6901DA3v2QL16tIayO+lGZYSfU/od+HPTAfoi+SbOvqKLpHUgEf4Xd
xUVXSZy3+uCsuI6uUhbZIBWqp9/DARVH/tw5IVUbeX3vjhATSw7wNUy7nG7GIn2aVjlx+kvdSt5y
00kXJ8Li8M5ssu0BtJa6UEsBQQoKlnGJDHJ8xM1HK9tjtxkf/4A2/kQ96Lw6E/gq4ef9p82iaEWZ
l7nsKZZcjsowioPzv4+vQn32Ng4KjV0GT32yeJw5r3c3m0+wAyFGd93ZbqeZIQ3KdLoEvcQXF1kP
oNfY9LgZv11+/Z6oopGTHgKQxaCxZz4KfxBnFOtIeajqIsy2M1qkspsbx7XfPer882uNPAVt9ehU
GRfZqvsEVPSCkJgOJuS0C6fE3m4V8bG3C8xkiPajBAek4QcgqGW+CpMLo6vo3sw7jtaJr2+hdqyn
u2esQwqIqV2jImbg0DGejlF9BTlQ7EqcpttfGT5RKmUwRA28ZmijL+0mFZAEhicX8r7Ri1SIcz8J
HeaTnlhRPN0FHySl9CWCXt4zHs2Cf07oTh6vgcHGkg8FA9hj4cLjYJE67kWE1/KTULabgXGS6hmT
LRdf37YlDd0cMITsmXF8wfsaJilBr0ClFHx+xpFl8Yihh8fP3m2pV4o5KEEp9ujYhRcAQL9Y55oS
raWt37gOKG5UZTA8YFoqdL08Jfngo98SJTL29hRgJ9+EUOYITEgAxiie7dahIrg0nPuNSp25ipnv
TyAoaG7VOYD0veRliNI1W9F8qOol53CIlhq+qwG+m2pmv51cXs4mpYy3bpZ9VrcD0qZbDat+wua8
oebxTYzrldQGjmiyLWQtN4wTzmRxV5dQK2ql9UUFzJuhZElDM1vwzvWp48TeEjA/ms1ALTohRZ8g
mQ/v5MmFKqfUYsAwQnKn5JL95ySfAXXlrZLpUkTcNk9Skw7y2yy9UsvT2+sgjUrbKTHhvNYEzPI4
z42g0lsToYPyDMmXWo8xnMrCreeGI2R3oyK68/AASGp3RQP9czEdaj7HYXXPhxoreIr1n0llv405
zaVe8MZ59cql4bZO6I2b9RDPiTIofb/AOD5VYKp3Y2RRg/6gUntOECR5J6bxjMLXmAKItbK7tiMg
5cIPUVSUH5vjqk/BuArR3EB0HUUv5eR9kHKczAMPqIslyWEf9y8ti2T7aObcX4wKKQyXZZBjPpic
eKHIH46F7fWthfaFuWnm6+hs96yJidQo6tPnSmHtyas0WvSiOORhEQ/Ic6Suj+fL6cYQ6PbWJ2YJ
zVAl6/a5IhMh8zccyHi6PNW+BGb59EmDP55r3wS9W9O9ksYnqBeG8wRL7eq5fz6ce1hx1Z7A/YM0
rVVWOp6pddcSZk3+/MbGV21+7BNXLSF7wbHVUwe6EEC3Weko0litgTc2FsXFuj9W67Q17CUoquKu
UwQL5nCQtXk+SzkloFmrnqoyrFpeBDhCBSxNaERt4ofHqfBIiV2tROSh5UJTcJV6XJdSa/P/V2d1
mCU6jLr5lxXl1vEkjqt64c2bRTYNxnjNzvU9VBhhJoC0+y433VBtg6L7l4QU1tWWe6GR6r+TSmZY
OcXd5Ar/nCh69Q5DJPuaws0ESCKEiVvhPsIujt9dqkzlnWPv+ggU0sULGbfG3+OACwVkw7KK90Sn
BGSkeBLjj27U+jMrGnu/3eoseybWQmc0P1U42lJi0QDf1I0TTlxjiQcv80KM2+g7Uhz4TFL6q0YY
Cjnq3kqz+ptiay9pPnkiJCKcn98DyisgfawpBhWbOwGgd/cb+V3soccY4l9QQX3Qsi1eSxwhq2e+
aXXqlj3PjhSFMx+dyzm5/uBgcp0x0YdkyvRUuq8nlbAE8oIXzm0LXcfG+a+gHzui9Wn1JDGE/YeD
Oj52a0T6wlouOBrI/Mq2ryM/+dnHaZB9/f9PGc41e+//JgEOo3Ka/WcyK7Scldm2L8fNYucGsVh8
V3n3LttnhnzQMsXjeMjZe7zzXNZiHiqn7ngPwndrEfJbWlFZMLXUj/CxH0kjM927ZkO9PK9MpD7r
Ky/ZQ/Ria/iZtPzH3/+EGSXClT2If06ZsjfzyO50oqJ6jsvOOLLubi3DHq+a7aEQy0y39c0lFdCk
rRHDCM0uWjlIJze3DNloZDFQJnBhVZlXXX+qhx+sldRTeFY3mkWWsTP5wSblcQxZKkdbgcIbRyiX
BNpvLn9O+HRsx1iYHDHsptYLKDny+Sl5Op6vuMg25TdnBOE1dry7ByuElwNcu+K3A/dM67/WySLq
gDvT0NhxENRsmS0mcUxGAHlEZ0vWxBpZDA8zuU3prqsL4mgWdKKO9s6KNjnL6Vu9hx+SGwefjT7K
cq9pyJLsFmquFmXhUBSm4afD+oxyjOvCz7sk32LqQJfB9NkQM5wYLRhLdCCIYHjNpCMC2RaIM+08
NZ4PTtwYSxZi2LcAIuBa7TM2HecN83ZC9XwNVPnQsEiO19dzWD0q+jmzQ5qzzMhQZiEHa1qOX1fu
LF++ixZ90dIYdvm8Xvhrui94Q7MlBLZ+ZOMDl/5pe3b3B0w+Rt/9ZotHbm+WYedOEp6ZBwRhx1ou
xyGQrjEW5vM8aaKlwdl2rlCpF8nM0JOP0o0XtIT6cGYkphfL0GXP6SQzBfL5kUGmvqsAi6Leb8aO
8nLIsrnN+nGYMtRHvXQjz2PSII6wpYRkRJZDGTVDeslAZJkXRe/+mBABRHp9+v2USwgrJMrTcrGr
Vri67n6D35EsIfjO2zl5ajdsJ/5TEKR9yED/A9yOsBRSEg9tJyfCKQpkvGvx+iw6ouV4AwAExTfr
D+6VwwKjBhVKp6Qo24kWZUXvpd7Zeuv6vPEoIIgyn8CFewn885DAUhBMM1llS8cwzaaLJhbR9/T4
aDMCotSX92i8An/GcTkLhZum0XmsieBVQOYkQ94GsDWkHHjImC3jAdZJqS0zbnuWGSftQtJHvLk1
AAKz725cXMTO1j5ilqJ54t14TFNkXgK4hfDBwHzYumGzHcee9c0twRyPSNXkugeIsE5k3yIyqhgy
nw+1ie2tGsYGm91e2NX05Hr9qnhw9omFaC/TkaBD6hqI1i2F41hBJCQ2LW1BxwLGtY2v0mrlSfVD
0Y+Dm5oJlIuGcpvGHo1PRxRRGBkdnZaYna+ooEmP7evIpFdfNvcbae7YU7UxO8NOAJXY15S32Lvu
g7Qtsce3jRDLB2lfkQeYE1D9SXHX6f/qEqXPhBI0jgH8bPMz3rcVxHFXVCoGrJgKqB+KOtKY96aL
ah67THRkIh2xcv/I420Q5u2TPpBreHjFccLEgark5jyV8QwS0FsG2Z0I6zERPyVWpdWZ3Md6w+3W
0I4Ke8EYadfu11aYs2Lr+nKfl6WCRS4ikhlqNMnwZK4SJXBxDP9aQv2ZDPmBJjrC4chG6EsDN5bS
B8kj6ka3HKx+6R21mL4GgUG7XT/ssdbWPelWS8fO2J7nbK0is+CiZZMwHE9rDpIjMPZf+2hgY8ga
OIET9wFB7m70kk/XjJSKqvasamBR/OG0UGyZ99YxcmlTp8tp4jiXwo3OEqkwgg0WjLzlZ18NV4+P
nSRceu9RA61rPQ0iyTpSEWpaLuCVV5XU5A17IlDAI2EMQFLNI/1WvtUs3G7EL96VvSTkPBUJ8YnM
bxjj68dNxEVip7erY/A8Kh/7sA9yyd2zyR/wluwPyfT05WpdAP73rrrrvnjjFXbmKmHxhdESIo1h
XJ2oONHkutYlLyF/jncI3ER0RRpHctRmHLPbB1Y00RJ8Otw0r+MgyVmQvzQDsEzrEQrm7NXth25H
JJKW9YZWvb6teOPGhvX0/xYR9G9hc7uFrcXfLe+26Yure4iZsgnS/stVxsNK4pqbSQXOkXywXUU8
sdfGuKx6Lid1Zs4oHAO/pgF7A2/znup4ixD04+rI3cvXrxmie3nrAdZBI9iSkQDOx6mQtsUbEE+r
4OAGLftZtS6wObX9S1NNQxvIA5fl8PxpDJvYHQFQ3OgUrX2eB+GFcO2d/X4/AXfddYEMcpBz7Je6
yRNs/aB6If5oG6xTB8z0kaEej/mhKCteebwU8RFm9CfeMFOGJ32NeF33H/Wfxm0HHBJqSJaxV1jV
gYwaThK5aW3hJoN7jpSObpmcI0vRiLGxSewJyE/0Op4Frj2oEKRssY7SAnYCamF52AClswbkka6h
gotw4oT/4c4qgj4Tc2FB8HwO2rJDIK+570sSSHu3+EfXdWCLY6A0wNG+33xbn2/g2g9qrP4CML2p
Y+SEHRoPLGrKseSj+224KNn/0Yiu9MgTTXLAW6ox75lqiE+PxCGOrkL/ntsqst+PqsJPaV33SRKe
97vVD4ngwHFJBLwm2fIoanFFp5NFB6AnGXWr7TfR3pcL/BQ9ky5dT56bE0CerD9io9sqwLNuo0c7
o+uG9vsSAVN5UAoXDu15YKSRrUKy8TRQmyMvJGvnYmFaHRKT1igqQZAoUfDoduiFZU1hqsR8sZ81
/v8V3By/bpSj0IoWjPs/pOfwAq/49Cv/x6S8B3FaJhMjPK62cXgx8VpQys6umffArrP6xFnJheYA
BD7UVUyiw5oLiaYcLJhvDIG6r68QZJd92pXvSSZwtOrvslOkGwWOa7FuB01vieiwYC0yuNkJhHtA
mkQnlYUFfopBgG1OQFzpU3zn8hxkOFC0Gm87lL7V09iqD1qRgbl4Jn545u3g6KCS6WtVQgLlhbRA
BaX+ZzagShpP4mE05Ntg1vjpOCcPbkS1dgNrwtWwbbv4Kjj7c9A5VXCBMgEgVQ6FRFUAi5+NnrdL
CROLBmz6nherFalKKez0z6DQgmeknb/wcyp/qRdJzS7TC1TODedtpNv232sH1JTJ7n1IXZkC+A+i
/BrWKdmtagDLqr2t87uezzJljo0K8uzXj8J+huNPKQjke8yzWavgkTp8uyuJZHn/FDgSq9Mc9XfG
1rtS2sCVcv9hMPDaTkN6XCH99hQI7rdTT0qzxxu9xrzGB3jCcEvWuq8c3RJM13SKXRdVVXEK8HJ5
ebTwEFYkt88I6hAEtYyhmkJDaBMU6CbJdQrtbnlxP5in8XUOt+CO4uV43c5LaUeKdWY1hYGaQlEh
cgHz3NNgtiNpGR/CIWClXpcqVknp/+SFubVSrhpKxGRwLiLug9QRl29/JXSXedHrplL6HnC1Jsu/
kGJfue4giVkLIZJdjaUrLkkExW6ALTgsJJU4022QH3bvUrtuT4wWp7oCb6/9K4iAH7zjOCDaqvMs
PifaArbGWusbzGZ3Gi7y9V/6UYrBu7y7D2xtZ5nBCeVBpflNoXM0wXKHkPHr++OOfGbkFmGuihs7
GqYADI0RdMOyx7jS7KJ1PzNExNDA5tcAc+w0eYH76icShjXje0K1i5AF0oCmlNiaITusmWz3z1kO
76SH7EN093MXGyV9DqFFJkjLUfHhwWNdvVO9sKfxEtQ0VKc87ENCr/Mfmx1wBNYgco+4opaYvEb7
V8xB3gFCEm5/GsWMjF415oxWM9ng1S1dfqpNHPx8+i/XyqH6lKdl8Phbd929eVqwL8eZshrB2SO9
t+p0Ej+v3N1Xuc8nWo2Q3yv0vs2PWTKrjM8Isu7osHABxLSpt37iYiKCYhDJnArx4uEJqUvqdGXI
DdoYUULfCNRnT2ziC7Y+PzhWpZ5TLjaNHO0ByzeTL78iKARKgqwEU1hug+oMovMJ4lTmRWxyCQAf
gkxwD00o/DoRoTIp/GZfK2AfvwmpDr8VFcuiz9YVESzMSwGzS/5YxmjPRZs9Jhm2LPVCLDzbCLqV
NUOztKSNdVITHueSYh63N1zbgyHEaG10vO++7zTXQSfqaIzgrXsQspZkekTizzD061tPLS7m+rQt
IDuiVppp2D1Heq0NoRQIYBcnPmeBpv5YR1S4z8CrYWVznF5IxuMRIU+uv6Nr9KSvM8mqvDzKBOJr
jSEDghc8luo0dMg4Fvs4CObxJcP9Na+vjOvS5e2SCFVmW/YVbR7ZCzRY01ZyTOfPvHpnjv5+y0kJ
afydszQocjA+7mKJUgXOYS1gp7+Cn/ZJDPDLZ6055xxFuxsnSaKH5JhUNkfrumBpeYH7k77iFRCn
Rz5Ab+IwsiSAp0KJY0mzEnkuEI0C1LfYcnfatrFPyNCbp/FdUdWw8TFP69CrXLjylDKAY8noai7Z
aSpoXZ0FnfdnnQS5HeegVnPCe++2eOrHigsPTMOjUOJ97wp9AgaqiiC7Md7ahHQnAOq05ud/BGGk
lTMoHvwq/sHqDiLovTP4YMCV+dK5Y0rPzJOcDiDuoFb5OrZew6UZHJf3PqQuzBgWy4pqFokaLzQz
VC2ClI78Y3u+dJ6/x+5Y0XamwHyDQJwjesRmuYsZ/SF8PqfxhzZHt3zGU3BZ6+y4SneslkGG3gcr
1+91MyE9bbFjZkJfOM4Cj2UDRXbLOopOcIy0gU7SA+7+lSiI+PD3qy+Qgnrjp+0f4+oDY/gNjcT0
pIVCSY0LJR+/cCqWcCY2saudiCT8WEyYBkXm3CimWG/E3vUKmZr+o/brZ5z59ADdxqVHnREVXIFB
AEu7E4+iwZ07w6hbPiGFhYqrUsr4iwW9ipklxUV4WvEbyXWeFqcVfYEZmdMQxRDx1kOQ5NabQj51
z1WK1OGQIna5+XbQsKRVvg0naBusA/2gQi/kp7BRe7PPxdx4t26LLGktinVNHAxVm796kfg4xGA5
t0c2StyRxI+QiDsFY7JwsbyeBIPhpK/oLPyxu8qvRaJGz7T6eUdnAQph3NqoH8KFgjrY0IqQjw8q
PKGRcX8H5TVGlD4/nb/9lwGcDM7pJh9L7XFmkrn2QwxZLT2WTudRyA5clbqAen2+U69XAcvZ/lgz
wjFUqQ4mYH8ruAChGLA46EeSzYedGK/cDuR+zEj5eCqzMPsBVC+nUJUDR7T/6INXrkMpOcI2Zaxt
MW3282tdbrWj2ONV4mtzN16b4icv45id0AkpcPv9YhgNDrv3QAZ+LLrMf3Ykxo1VYsGaWbOPzZWm
yVeT135tE0QqhpElQ5KI54OK44Y5ryI3TlAA64Z++YauOhlDx0Cl3u5X9D1KWJ9NYG0+QyusN9XU
SmpxwBkIGTNzUatBe79Lf9iDwIxEr91Gcx22fB8ozRhDMa0ChCjIxjOsoHPnnBG7bFoa9DdjEGfn
JhYdx/zCJ2wbv1JbZ4O5Skb29gYnmZOqUt5eox+t4V2bL+ioJml9Yoxwk4MGaM3IOKQX1OSYBrwJ
/oAiqLcWdWvieFMxx42CUI8oiuMOrSg9p1ZPsGrjdGL6lzAYS7NC+r3x/r3nWuE75cud/xBy+BZC
qIL1/eBMq3XxL1hOnS68EnPrWF9Mrv4TOEpSeK4P9CoQ5mtUnvt8Sg5lvspSaoTiZxvtqXLz4kk/
/ryWVsn3UgYa5KEdGeEothmRz/q3RPhnn2Mw9pk09ivlZAVX/qHlHbgX4cOdV/a7fyr5lMQJK/H7
ROxwGomdU6rICjx84kzK6vr5O/YXROs1CHI/ShVKqUSOCxyZyalJa6SsOJThJln3lK1vsw4xI3mQ
9jyxjMj08e+6lKyK8Mb+5J4pEEGFde/jU/xdS31+mHkKlAIaC3OUfuK0NyyFv8i1PdkWKCCRyhUD
X426KoV0udbPdB1U3i2csg/zpSZAjIT+Bac8s5cO4fnDHCeNXrEUP5Vvc3nlaRFAzd/huOIvxYt6
yPJwICAimLBPQTSXHEg4u/Ew4EfPGAkwr/IITOLIZAhaszfWiT1bdHHJ5Im+UGSxaN2IAGI55Gv1
XYF/0osQmRs93GF3P5uauK2J9PqlHIGyyoFAL75TiZeACPIIsKTQr9nfGr3/wyThFv5ne/677O9Y
FQIzgqOlnO9lMB6JJWXALrfNYwiXuY/EaqARHxnCYhURP8RpTTi4x4pEiClO9b5rC7rMTEbK1/zC
x7zIjCMWYA6gRALQIAurBNylOAZ/3bo21u07qce1xHO7ATwTVgsQYPX7OsYkN+TY+Pw+XeD4uUXl
5SbKYZFkSoscms94QLoSseS4zuElnh+kyuX9TJ0jdtowLiAJO2zAGAwZ+MtY/4ebbabtq0v4//ge
NjtlbV4BsGGj/Hwxjust+Lj3gbZd4ifiTrHRpZwFFF241HXgJciuACCrn7Bi2vkgYLmA8etIyQg/
xOXMtblYpRt8T4JIPAYMD1sqzNACzf6gsVmo65ARyn3Z7BO6T/PNYJJt/BDd/SWV+ccRtnzeBufa
EaGQNWQg2Laii/xAhpX67/+JFF260jalaXNZ5rRuavj7HNBRKiTw6utj5h0D3Ns1s2PvWo7uYLvj
D9mBbcp6z8brVDV8CdGMZXBC8u6BdA98Z7c6pu0oNXcskLNxR3H8XOhWVLYASMG8FVdx8PKsbZwp
ueGAtitQ5ZBBsaxeCxg1/4cES06kCis7hRLEXp/TjiL6g33eUJ/UFdlYBqojhQyaqs6/EWRvWq7e
jW8ri66mOX94Xg7kV64H0aZxOhy8AxHiJXbdxP1UVGX4BrCqzPIf7iIk0gg/R5bnlcXXjcDXX4oP
m61jaEJGf/Hm3XQ54bnMM7ya5pfJSL6c/2CWv7+dHVb2NMeJpP3E3Q76d4taf4FOyPgKxUnx+5x4
3LHkpeKhnwPXxczYiJ5NkyFgPlX7R2pMqtRgy/CSgp/oCZ0n8vZgbYjGIOl5FyCmUEZJi3pwfZ7v
cjxAYNC2+p5/9x26XCAJd3cuYw74XOFOs8CGidZUxsEQ54t0sSS2YzRt8x7lwIYwUhEOxNafO6za
fBPZLTRo7rAJi00pUVYVI+VkDrybvjITYULWVsllGcVKkn20yjijl5zDcczKyIDFTDcLmFvDmb5r
szzGcE10l34EwUbxlLBKlKVs6Rt8ByDqkoLvHXGET9/UW+bwJisVp/jYVepavk315/i0UFAWvW6l
Z4OH4tuFac0XI5eXLQo0tiqNQDO66jWmmuOJ48ZYPmojKPfib9Xu7odCpO0/Ubi262X316fDhHh5
G0NVkyPO/65XOOdefnFiaMfnB21Uqvxsiwdm/PtULmobeshLp3Aknoa22v1PMJFtZWFrbCP2bW6/
ob6BDVaD9hs1y4xl2mO2fKcbKK1XfanRRjrFdJvJyBw1K5jVJKc06GWXRbnA/ElHLeSlGKAJ2yC/
w0DWLATBGVqGX1inkr9GUOL9eR1uw5lPn6B/n1ZYowPrjKYjg9ln1gKCmXzJuWmTXn5seQDSDIDJ
XAkcrnAcv4jTH+64N0QMwcztDxo6koWBbLeypbyDxXrMi9ylVYvF2UbCmXK5UmtLyJTm9Sl44TTG
80I3pnBmbpppy/aKF807CqJbcsowHHXvnnfYym+hDW8yHS6crIDo0+pQDuzz25s5R+Q4L+nMPKOe
UA6HCYzuc9yATZKt8XyVYmXvKIpAGedKyb9hdtIQjeKspYHh7jZ2+BQnywTmeHnuvmoNzsFfy6/M
FN22n6MvANJxRQXrG3v9MdOvyuo2UahDaV1q9vSHQdz8AgSXPOljeE3EFT31z8KxCl+5UeQR0FzP
gyHspoALHINUVzi1wDJYH8USKV70FFskN8NghjsF7OpgC+Jc9GVBiv/tf1KrOeY5tj8J8HFhbCqS
wk04elVamAqgO1bsF0isEaS1zkmZ1TEYqQAvmPQDwoakOarv6H9Ci7OuJY1R5LHMslQd7TaxkU56
NQ/67/i4KKo/ur4gU1RynSsR8xNsTYHacIasK1vmUpJ7S8QAWeFFDHl6X4zJCCAHaiGA2C+aVRg3
3d8m0M6Ag0/08C/ODGmhxRqJXnJb5wBJbvliTLBD4gJB/fgenAHaz83m7iq4kL7hOsXPMP5jnNc4
HGEWfgri/DaJWoBWWvrRRVNR5PneXyjPYGC8M+6KtArhd3DV5BcWMPWrX+lM3I+oeo6KiWboEGPP
niLnLNxldDqI5GDkwoDS2o0eC4d+/e6lEaeOyWC7gW0uqTGJqjPgRQYI64Zd8LPUvVGYd/zRZFc0
JuCOllFy93aqdH5z0LurpqKvan3U6IOhG+IxGVV+HDbRawcE4nddcNAyhsLbn4+rjZVBsBl8pzyJ
q/WDY3dMtf7K0kDL3YUwZpTKTjpPwDarftplJanPbea3bEZfV45L4cLzG6rb9IPx4UJOYzIyutTH
oCkqj5YF70eAxPkkKfIUr1v7JMB+RPYe8rnfGzUG6ymoQQ9PLoaheUDMa4q4iIFipdVxeHb0a9bq
DtI91cLvo/cTt9a+H7GLhNfMZSwaL/0XDwaiW4Yd2OhAcmeWP+l0SbnWhF07yeCl/AFOM15ksgof
j4HgYAUE8RPC9B9BmfZrAHZldodgtMS0BRmguBUl2Ap+Vf4fu308qlW7Ov4WhuQ3mNaNp+t3benT
abixjYuBVEwikgIFxhyHDbg7SdPkoi1iBIeJib8A1kcGr5lRjer40eUXBH4iA8l+/Kz2V+iQSSnk
XNu8C5HTq9HPSc/FLRusbeg3XXD/08GC2Z0GRJwHLghfyK4U+sIimHTjtr1o6J66tlsdBFykY1nv
vV4j6pOXC2BYfYgV/bZ3LvhEC584Ma74KQ5xFxE/aF8YDyGY1zWPW33/v2e2WB+CBpI8GHemLVJy
OagcC1sX7/WZZP3z/dZGkLcjZyMBlJ0tb5iCM6eWY1H17YotILzfpfbMLW5vLyJ2O9OvMHsgJrH/
jCXWRZkj52DVG3g0kCxmJJmcOMhCKeKLOxVM0wRw7t3v0+sadqZrT5aVx6+Kr8R8MMVP3lkIRmwu
cltKSqNHqw1LEfLQx3CateI6ndF3C0IcTBm1x1fyzB/DvCOsq52lPC/fUlUqkKKJVy8F98TFR/XN
dJGbY6F1/ggf5PN3H4wiZ3FAAGfcf5yoYjlhTEd8XQKA+WBWLrQNodjWVJe6wnWhs79Lj9bX91eV
vPLdvocimkbINc+DN3IikZExjAgjvGqudVxmlc2TZCxYCsKgRtoUOsnHzOAOwZBkTI/J9MruicdV
uzYkTSYoEegwraQazKgVp6zbZtgsYuRguTp5wcXRZ52z2Vm7HkagdnhMr+TGI7upx72/wt2WUJ8e
E2gIN4BWwArL5aCGpL4F+DFDinyTRpZ/jKPxrIecGmVMha4FBHRdvc0NYkLkr23wuZhZBW3qKSrB
bljlL57uIgdCe3t2LJu2n0w/cv8UePttxQnBBEjOc98k5cR61UUW2tVPbJsMehGUDpNt2FJ1Jna3
umObc4yagPUhl/iuhFPIWmLqX03SZhAmSi5nLremMq92XX0YW2LeRjHB4jL0VVIDT4cZJ0EHRrvM
3NtDkusS0RDYl4eDbw2cvzlPwYkLRr3eAlbgeC4CHn83w1dIWX7waXt+T8usLyIBFoYkRYvwNOxB
jFwBp9IZ22itqg8biDfoqvGWEjDVj1JWJmjw0CoX+gU9wnF2aJFChB5yJDMxUK7sts9cpzcmtafM
VB6fN9VcPrd5KDpXRDWTFcDqv6aRSreLKwUfCGtb3fj8T/qinIv+pfab0cLs0FNnwPaodgi4Jc2u
0JRx4fgXSxggHJnofWLM0yqoovsivjg4XSFIwhZoUGIbMDha0/3M4K3a/cSfhctotUChZSRk6ltK
KjOry0ZybkXWfrp7eQiR1WJId2ZcXBs2eVZx0lgCiR38XNrh+Xs7xXW4bsLb++6t+8dSnvQ3Uprc
tTQMcsPNJBmitsoZvfyC/BkxJfxXDFcaR/N8zwKsyCOB8O3ZO7b5XpaUrXMA6zo1sOW5DxXfocRH
Fe4fT/jlqqZaNVlRjD4TqGOBrATI4Z4Tz4QHnY3fKl+RTt9KtMO+V18yp7WLtDYK14hb7oR/NkW7
RhvQwiwQPGXBadKvIl1x4ylHgritXR28lehozZ7YOVdvdSBl8xpqKjZ+qWsfxUfw4YYyV4N8r084
WMEMNuLzep4LAtGDg9jYMZFNFKvjRlN2de/saBKLcBJAXsUfumxa2mke9Otg3z4gInoM1Vxc2Drh
47yl5tFyhCqS3fH5dmS3CcOETaH80HaqffB2NaoK7s3Pe/u5tAB4hN+n1TQf6DlVr0nS5Y10I0aH
rjSLYXkgI1dSGdph1UaOG4hPEvu2GHKXkiVj5sJrq16XiVh2qZUCdxnBggxnqCT+3Kngb8elCyKZ
1JtEK3k4heJ8MtIfcXBZDu3Pw2LYXI4Bfp6JavzfAFEa4LmIv5r6+bK24azczl5wZ+na0cC4D1e/
wKcYK5jkoSvaqW3/Ehu2rC1RhDhb2rbIQvfuf0++ohDZcFRBZ+eauUtA6/2YkJ7NxEFKlcw3QM6w
dCA0IUXjXJlNCMQx4JDjCwd3u4kjKEUeYO/eK5qEZDPSIAmHq6kO6l5f9uGPWjxgTuU/NllytbPO
kfO9m0o8CjZbH7qLdlcUtslEhUu7nC8+FdcwLHDkWe1Ss0f5wIkijoOU28a9hx0EDMo6d1rjueN1
rdXWvvu6WTFDOXxZKYdSeAJOdwSS3p+75rfJLquerhzBU3KmMVW5MCJWoDh70aWHoHhOQyiN0DOM
qTrn7sbGDGp3ztLKD6ip6/wiUISdmI1bZWijTPErr5whFhjYoBj/bQNaOSGoOm92x6ZUpuBW+gce
pXhAxwj3e0SQSZJsK5ZNvLudYtWlBbBfPXC9GDzuWwtPthDAzm8nNTNW9LC/H+wdqqDLrT7yhLFA
+KSY7A2gonJQCBDek6PIVn66A92IrYXUL3J2ckrPoyrMuq55zyjQGtmVP6B8ndZiDMU6EPAWwvNq
TVhqjVWIPqDE7wKbBQCdg6rSwBTokh/cvgPH32h37lMevSmlR1EXEnF9Zv2uekqwiPd9r4+iPf6V
RBlbHs/6vLtP/+7CCMahTfYpnAD4jMkSxese4BhNP66SQaoqEnhC4PE1lrqeTYEL/IFpz4J6lH9W
rhCYU5NNmIT3xUbtX91zDIuta6+lkVs8rCwbHdxqOHuQDdnF7N19DnEOylQT2NGMjBMctW8Xl8Jg
XZezwfQImWLBc1/1hNnHgi/IQMItMDfxSUOUu+hIkKeoYpSUYgvl0PJ80W7NJm0R/L7qLSg7vCgb
INHBtL2eIPoHekNU7Rc1WQc/1lEnVcRogU4RKpYytKxKC9Kezk3zTu/JbBaWv2E3JvdZFulOSyDZ
N6XVZmRvQxy2jAn1y8h4AGpifLqlkYOmcAWzSkMM53CU5O2snscIuAMMZb0pq5yMga/QBlX/7uiw
fuoBiY16iL+4a+2d0loqxZQGl+pswDIdf/21+6OltHn2OU1P7mSt53qdBmz59ILSjIFcXdJtt9w1
Zl6T0XkTHe8A6gMxcNmctNh1jwq8cFUjeTYT5fl3L29M95lC1cMkaLnPaZ4m0Fp2uo5D3nMgpb5B
qPa3sbqd6YF1YQQ0z0fYqqslQyBjVBi2YZnCyqczVe/vCXtDdvTH+bkRBXwv7HjxTynMz+5mBalF
IZfiEV8YomDHuPj3MFqyli4bQ4OFhzaJzAhZmDhFQBhm8OEMDYwS8TrNPuk8Qb44Eq0N1/vBpByJ
Ps/DDGyx4e5BjrwRZN9JrKnbf6DAr9GAlzarqHQ9nmFUmUmjMxoaS5+ExImIiziDOHe6YkXH7lm7
JdNqCKvTKo7rlLdmSZhcfXisUeBQEpPLnMnqEwqcp71QapqjDfK8bAcPsktuSIM4CW1ytDwwZ4xV
BwgxqcCSrpJ6nBLwazNXcsjZkFgaJOyykDqnt6TMe2QnafeyxLVIk7s+PSoUxxR57BXLgkusIYfK
AtPHzotX7pv6f2smL7budvVjBGPuyuHMt9SkbW9+hbq6hS9GMN4jfXWNznJc6dzXW/XdJK7pLmWU
CzAYJMAcdOjRpambuI1SVAOsLKakVXQlxmXdeX40TV4Fot20BYJSphilA1gRtAQVak5kRXfy4t2F
J6tRlX6lmETugzFW9y/aAZKVOPUXtPS1ODGPzvx+DAMHiFlTZwxbAiDUI9ZkJt+zvTUP1xBxeEh5
Bcgw5Cv4gffkkE1DnWBxEcmtqSWXoSQX1bzXDtIHKXMHZ9TZJyTGQNZaCr8d/cKFNLFEKeHvlVmo
D0tiUa/NLaoDqraBm0ENA/tVnnwpvvN0fEbdL+qAbinzirHKVaQvZaMiknh0iG9VuHoCuvnJywHK
cDHqV1pd/9BkXZ5dUdvdmsxkuvLvAI9GYIg/Ldrz59BEaVdwIoMJmbIWGrG6CAqVpLxjOB/zisbc
if0XWbu1xg7nNwxKxvT2AHlJ7+5BesURNKjmsNQZn7tVVetC55bMEDakbINwWb1s8stmVGdpuoZZ
FZceDRj4d0CIR0RYcI6fkil5NfFCCsnKLQXTMha3ya39310yLM/nTD4AY70RrEphilwlUrPXvBA5
SeKVEiP5MYGqroqFejiT7HDnsGfE6zg/3j94U8uqx6ec5bbEGQFiqzMANG6X/WK7lsBr7doJ4utL
NjJCeXfMe0BVfkxWkyAcT+sEIHM20tMtoFrtAlTcrUnIESWcFHyoew9NNtqbrOtHulsDlnxJl29R
SX9bhQngoXqxnRpZRUR7ZYpXYNkBSB/A1CzBhQKC0+hfIpX7SLXb1+Zm2hH9RpbsblTsIdYBoA4F
vOUIjJWOQLqoU+JvREGA6Ewmg7pQUhRahakFPepKDc4OD0VEusKGdNgyl+VyDq7FhzXE6PSJvy2K
JdFEwwFifro3ilbIN0aPu2hzyc2duhuAst708RnEGNUUjt/7IhAfbBhatA/A4q6qSu0sOQa9qTbo
rRt6Mz06nOqUPJ30TfRWkkqCWu1OFkHmwUGWjW2c6XEG4SaLvU09+ZD6S8tutakIe9922EsyMn/w
GVEH/bBSr75Qp6WNlHW8/d8UzdfGJ+DIytWyFm8ny1P43LUgPDsEQ3F8/ql5vnlPKEwbQhdUNnYP
r6Ew9wNe4/jTGtvEQHiPNa2pkpJvpVvwAeKloLOLwPMbwyixgjUGSSO6DNIdeyrPFcKLD9e++RZn
dhZiQAxXitYPxEftkFwai+vlPRkxRvykFCmd82Dj4NcphGqpPizCo71rT13ZYS0+2j45XtWsCMIL
vQTASUUo+w9ElBMxywYZn7Y5OSplVFvdSUUUHa3aBp8PSXxHrqzGvuUEsac4vsMdoR3AcDDwv1Qo
NStDKGpk6zasNyzJ2nv1CIL+PNydHanveHy+NgEjqIbgqOzu1GVCvskkga9j+b1zdukPChI8CI9f
dmHZwegJrZKmgBNNG1KIod1RvqZSnwpysw6mg7z5sSMLF/wVnTYtqT7zsDznlMSaotFpOcbreBeX
NQtBu4teDQ8lFjSm6Qlhbn02eGiFLyKAQpjKWVMhQQfcUsuzolAOD5Aq2kGkvWrovQhQ3JhWbQtQ
AgvK4itSj0u+cz3XK+8hPQSFS8yroY9QIeBY7E68TcLy3N9ZGHxYn+c9QgufYvOziUG0kO2qJJqE
xtu0gEnqZSO9880hCnWe6LNDMLGyGRgDaqvjXqQp+wRTG9/U1i2JOHoW4DepwdDFHgWBOokPqBcW
Ju7Eb6XqdQv1cpScLVkh02M90klqGpkrmSyMDliFSVm3OCOjJIRT6SHw1F148UJUKvIGKaWSnnWx
k9xszCftYFIS/GfEl3T+gUgt/lKKiSI7oEHQc1q2hv3AOl3DUedsEFsIt5NT+p1jlxCOWsw/nN5e
d0KGLHGe/UA3QODiCT/WA/UabmSokmvLQqyCWJvRp9bpD5lMqcJDiBvv9HyibN2obEKeF1RHk3dx
jOCttZpNiQZW762iOy0lAePV6HvIhL1IuTd8L3AoiE+isGAL/cRBOzu9pkgm0/7ysxH8bFWXYuPF
9sBRdb/8zMTWxoh7UQXa1/x5A8jMjGZh8Ym1f5M9KZzsfB+hdb1ezE6Nb4QNVDf3YjewvElMHCBj
nocIRZNaglhjyYsp8/TYG5x+6iu5DqAzWNAqeZ9eUB5nvlhNYl6qWmxST7saqf1K7W1yd1ks1TYF
g4VrserQqwFbtQ1LOFhV4reW3STVuat9MRm2R93X/35AZ1vmw04BIeqE0vyxhCYRbJvcY2L04/Qe
ivwXEnhD2Vq8MSZYHqS/8hsjlrfjYQrTGFasr/2hN0Zyhb18z8xZPoVO75P3muUDVXQppMNEyBuK
dLxzwcc6SmTJW6qiYCaTvsyItpuAa0u4ThM2mPJ9hmuaT5aFaegc1MlhgkfOW6wBOLJMmiFXMln3
N+GSQ05sNA9BupQCz4HCcdk3d1LByT/ciGHI7NhEXakRFoaqzku5nxmcOCvnbqGW0NFLRDdBX1Ah
xiiCZYktE+PCkj5tvnyzTFfPwwHpWrI/gXQavXr57mmJNpDd38j9D2MCn8bferLxDrWAkEXkxVgk
+AHzeKzOvL6M+q8/5oNvUcljgWurFo+ceTW+hHvQTPjgDFbA2ubxk2m+Sizbb95slnL+R770xPt4
YeGBJil39D9W5+cqQZ6We1My9ioDU3aKMW8Si4Re/AxQ5rdGwIGInezw4HLfxvolwRKoLJErGmgk
zRYA8kpOy4M3CWp90NN4FPHmAvcVsqzMlrG8eyDPrK3KlJ/HeYqWUxC8JZNTWwqCtuYShShec3hU
JkiOPRolnKKqkobTzhFn4BH1/M7FJV3jSWXQ8dFm69ggV9bLW+Btkji0Rtva2DJ61wEcB9a4Cntm
QP/Ty6hEkL5XOuNq1H5zEn+r/63/6e3Y8Pxh2YtcU1bNYT4/tIVi7687HlNuTkN8iWBx5vIL3oL2
9EkNi1gahI/JXJMHd9RbNxBNJfQykcGxEvWK57rPzyVUcNZuAAGvYLAfH/ae54TQl/BZ/4khikOL
l4CvaHpenodnyLsJN7a0uKg12C8psQqTs8LmyY5WEeGQVMtGoeBXuOvAptf9R7ruTuOMD5Qto8a7
w/7sQZjCz0mjqUTJaWLOaJJdc1LPJ7N0lmk3w+hQ6jvcb/Qmu1cHIUF4ejdYdDZrudN3Zcio3BHb
3Ffhgkd1GTQmbVti9vE0qEGLDM/nG/ugdzNyf5SPLeu9ZYK3E+tBK1AkK1fNJLwOjfJc1uAzHDAq
4uIMgXtd8ZjUSk36jpARM0N+MdaiQwSm+CNqmqawzjZKsH4s748eVW56IgVKXjOKedoDAg6/tPUi
likEeBoPkRNfzmPtUV6xpEGGUbFiVZj1SIp05E6TGqUbuWvSz01GvGHA6mneCDPe0pCncQHzTDpP
x/2cr+ksEt2J0S77HYZrjwaKan+vSrU874Hph2bqtQ2/4igwlOTdhfKqQ9hesA9nrHT3DWiOezlk
ys5J/fZf3/XylGjryYLHMEl+o1psdLg1tOKy6nMGKDpKbMZil7JsTMCiEmlhSbimYMiQLs2ZgXhv
TCeQCwyyC2U3UDKecy54HUQRU3qkhDVRS2+3xCQx313tcsRFduJ5gE/UJGt8B9arvukGDxrH6qCp
bEZU5VH4HQWGVA5ejy84w0heE6uGxgFghpYCD7MPIO6S2mHp3thxkRbv01nksA1Yr3vjy0GhNJTw
6RI1tWeV/D9TEHsdZt/zrzJWRkoRkFFNEvhaXuVu7TrB6wYttb7jSalIK1ed8lVlDAJON1JPNIRz
r3CE1WhqXFf1rAhfEi7s9KgaoY4fWvQKiv4bfnE3ReavSgtDR4yBjBB/T3eXdi1WMCTyThU60KVm
+uWkARDkkQXdoX/syZmgujobTufmCSDG1ODxiYqvK+3eI0WT08MEhVQxUUizrve6ISegesBfkNFI
ptEHt6P0GHUqSpgziAp539Hh2PUnZI3+PPMFMiNlyTskV+10ZVuUorCq+VAbiAB9ZuttIjuEyLmA
NpklYONu0FJRh7wlfMEUxbKbFE7ui1kvzflEqEHGdbSCah2RI8bxmzdoR0hVKojzPVmTLL6I1TV5
yKjf+D83+ag7zbfKpZjm38jXpu0vmtydhO9nC68indASu9jQ32mZLLOUWosHYCBYDkOLCTODBv1V
hxC9EV1gV9bmeRaRvtZaZ3jZfoqmA7x6mAbMLwVEVEPqN2nxvoqFUYFoQOo57yu7an+HuHAVYenT
oPWLaT+cUUaZxeWWlSvMX8qJtEUhu9FMAnndI1HKHeQ5JQ1YelfPOQ1L5jKCCktnOswXPMwQbNhs
W1zpLDytJPYh/uVoQGWJeR6ykeH7bk/w/9xmdah/fD8LnCdYoWXxYOh03IVXWzkJnvfpmgcNVW4R
ozbIjKAES3rybp5iy5NPEwoOGIIjAlcEGwvqp3nMoA/bLQ/IfUrxMhCtOPPK5rx2Kz4GQci9zncE
LAD0I/wAF6MrwJziutvAnG33Lh8+lZdNTvH0uhVuqK00S4qiUsLODRlzmXyEbxUzzMFB1wrnekkm
PRy9b3fjN2bT+o1OF9pMbbb4o8oGjIfvbZb0COJQk/aBBGfq/Am09gD8wQdJZLEScnvFzEQGferi
GYYF9M6irq4yu+Q2xtVZoyaoe5pe6mu6hoPUrwl7UDaFqLdgypH3SjGZgiUrKcdSH3iNkAL+sp+p
+pMyE6/pGxeBdxgW+/2oiP1oeZ39VDGIeM5mdqMlEw1FnqF5KoJGrVCJ7x7fk4dyZtiw/rKtHJAF
F1rfq0qa++g5+/Bfi/8mTQ+WIBGakL6nmVV8FRg9DS5TjjOsP9lrq0IPfsJY/uYgS09QgqxmZbqm
X2UZMlzucKhMz71luGyF/XB7kTJWafGvM6AiaSYVdlIfFS/eDuTX1PbJomu5h24qfXu/KxGJWYXT
RE4Ka5OPF1IR23p5X+j+PeI033mSYpkVLGJ3ugBVvL9/Q1FFew5cFJHOQIcdNM8eIrGDSYW9RiSS
YEWhNW9e0xgmJMfkHH31tXBC1YHEFOxJYE65q26SncrFvfmfTAqxkx+dG+rrkiPmH9SVXl0jGlf7
i/BKf5oQKJxFAOZTiv7ZuxEVnweOzuijztK+7NSH/EKtfjHsEDTGbjv7HkzQLmhW4LyGAYsQ9xJw
h6nkI0hdrtMKOtijZ4i7FhyUh1EzZ/rUoeUOp2nMB/XxW+nJ7i8P5MFSL8gYkNhMyfv7NZSnjLa1
OkwAks7FOorFAdf/NV3DWEvinka+d6MId6HGGcZ6MkL+wyGJJdsTJfpMqV3JmiA7DUi57Gl8rmxm
OgU72eB7Szbq0rid/QKAgZcXwWWI4vwbnlBOhEqJC+ZXQOyRXc/YLwwzWD0QhjpYRAF/6w+ymkm9
eV9VX13MGf9RCgruy7xECw7lPpldBcyRPS++lIPNvGUKXwfi0H2fVu+mIJgkvEAVq811LQFuJiOD
nF420JSkxUIsI9q3ImL1ka0NaISzsG7GvP+5DIDuqOtBP89aOV9fjWqaXP3TS939oJoISYtPr/fL
hHIQCa1acfoYkcGgSh8M/fBeej4yILeWmcwzTRWRJqd4/1RqytNHUaghlAg1UJ23qfWAokTLB1k9
BcrfsYggv36VhCUNx8+DUx+XQS3PDsaTiur6/qnnITjd2V366mwNtLgEddMmVvnVky0SOJdFiftC
Ch+njFZ3CvAKyrRopGxy4VyFQellXZLTAnXWKLnqNLnJOIIM6/3gmO2QY6DoDBrNsaAfypzYHUfs
cB8XwK1fXGuJKcZ2jAWUIcjmjEnBjx7+6K7B4kD0w3cr60ZlArBQ70EP3OsTuwtDDjEQZOfM1Asi
d34sBndPFUHOn4lk8ozxK88hPx6+JIMCeAA48V29v1Ht5Fd+Fa0/qOEb9tBewkDLVBv3Gt+wESFb
aqAV6ZM4I6AUYWfBqaRWB+usbaMKo97KGApjUzuxZ8+C6I+TxAF1RHtp3j1faOJc17SxgYPPjf7K
BlV4ygf3mw7dfUmPgRJbDAq0npzd+Zleme+2aVaJhnf3ncqGi+XOsWzRKVGzpwryccVETqo0rKQV
5tqt2POY+7wpMH4KtfvsNJ0zoZushR0UDQEdp6zYlJMZGHAEQ+VSD3V9JzkeoE4Ce4ZnGqKwytyp
R7GvsDj0pZlp/2dhuoTgXAHfHB23CxgCw0eu0C/1pbZsVMarU24gINQ+BnbdvN/u7UiVklfwlFrD
/tQTjV5Dsyfyfy4YzDEC8zHioKPr4D+toOf9Qm83LVgyEhQ3nhdPrkYFAxWotjQ4c2atnI9CafbX
a3zJMuJwaD7XSKoexia2iPft3xNpe2dO3X7d93G8YPbpYB116ZKpTe3xu9amyd+uj5qkdfUWXjTt
ZOebheR/0dkURZLzojqd8EK651huMcvJsf5sMsNp1C5BWukWM7v308EM5GlkRdCNHCG/1Akv/iW7
HeAMylyRLxoJsOv0s82i791tZUA7r9/fFZZaw+yA81HiRdZtkYocopaDiKmHgrlSq6S2Nv0YbcSM
/trJeKhaUKxv206mfTzzDTvdRxjxjfc1+2jb1OEf3M7+TB2JX/WNo2+EP2urJV1KHcCbOPxYm0o0
gWKTfoV1ksOIcVcsGLkBgZ2SbyOtNBznLlykwdajp3RwtKzpLFIbgUimwQkCKhcftE6wNnsn/mYy
W7mgmxDC+3Klo/wehzIhB1atb37k8pCkGGn6sllijREUsuS4Zs92em0Bk9u/hKs7y64lydaDfWTF
d8GMdbkH4dj37gzsS7gjJQNS9f5gXpGfWAjMZQFIbNcNQj8xNiP0liNTQa6y6vINw15Mo7yej2Am
KxPtQ0XCVVolegCu/hnDRaVF7w11qI0abQj/uzwO3tlH8wzPiRED422lPNmtYWbp/gkJuAr46JLZ
aizckPN1e7tcC5NK7VwyDfdJViTVTXyQfDikhAHfCKnhaNV0PgPFYJLiQF3XL878dVqeAoOIhDzb
6ClzpG6pDA7wbPbdOh96Q0aEcyk/W6FJXg5cpLFRYttRVvTraDutPBzv+1cDjxzk8kxFNLeT63H4
2j5z9pFxojP1LpdLHxPTrgm4aLhkYGABC23zbrLx5hE0sEC0uZUap3dJ3tGAVxHypNcSGo9aceWe
d+tNVEehY5/DtVMiqzHzTnLny14JSrtSCKGtWYTuC9WdH4WbWY7eqljX8/jOMiz9VlS3FQcci3E6
Vd66mvs7MVwXIIHoatofeB4r+41C3zn+thIB8mVi3RBivtn9MkuTrEcBwHSE/kLDN+3xHaHeL+1P
/hm9sbnm0hFVWXWFlcMC1RAXt/fH5Yr35bP5o7xxAw2HS+CuWhZVNaCCB08As5mZr9hO1DtGHAkg
dLCsN01zICK7yqhmRibgz6AdrEN9zpNSar+Ucek8K6Q3OG6l0xZF+DBGkdQK/Fr4Z/aNqToCtCkJ
b71DTslWQxklaPU/6x7f2oHTVIm3gzwIFvgUYhs66TX3X0us+AoXtkINjXvrLRDDZTZAvgYemfMj
c9YIuGlFKmkxwWI9BhysgO31MwFqxzntb2fznc8lBbxaNHY7ClJ3zGgMH1i64BhqIlExFl7M1nLp
x7hoSWxPi1JOfRqAnKIrYtdlfhmIZQNl8zCGkzyHZ3zg9txzXN2mjm8b6xvFSW7DW74sLkXfYJJX
/RUyPr5fDYLB2jjuEVKOQtJwB7S168vqDE9oRP0wLKEQx/y3iIDypPeAsqRn3FbIgPmT1xWQMvIh
qFVy4E3QTbE/Qk8MgnP+/iKOz2FVx7FhyqWtnYV1X5+082zGyZtkCTZ+rWwULPHJO6gpcD6S0i0L
x+LWbyuuwc6gmUhe+ng3EwZTQzPu43+0mUxLwWTK41BFEPT0prgO3zPQYrcTPvWr4maLAMRnmEDb
9vqyK0idOc/5D0yAYYIYuER8IbGc0FUPbnp7fE5rmESvreVOVaCQB98JmTcIBlwWjLe7Aq5kIyFQ
CMB8uiB9fOIQdCAOfYFQCfivgmIFKZrXs9O7DBucRj/TGbSI4qC5sBZGhyNz0/ltB6CZdPb1yKe9
TpjC2VqQ5vbOinUQ8krt48KU/wJ528LQLdx7KENVZUMbngk9adjzAfzq3T/3qW8SFdjY9zGyHksv
4hO5CQ4Zj+mk+1Aqxygl0A9sKS2EZG5aybxy/BHno1sZWBB5FozFGxK9cn1a1hTQF+y4njG/IFcB
Gzh9UAx+d+urazGp6nXQyRNtob+5qqFn5kcXYx+WhUea9eGVBm2GxUU014hgeQx28akTwsAAhji5
1gc1X6zsjsxPIEhjoDETSSdLqILjG2clBLGHN4VgFJXhH7eUsdGc+0pzR9Avs2rbZlYBlZkfzfU+
QyKlj5vOFyN0bFjMfjK9SYZnuZ42EbrHZ1jETx1UZwPKY5KKF2cfm3i8fTs+JAF0EWt8A8mHLcX8
yWKYrDZ8z3HX+NPzUqMnZLpBzNeHx9V+3T7zkbQ9dgBpI7Bq6vs01k0xXOd2Utz9xg/ZcVPqzLLZ
jNL6XRK/ACkH7g/zthAQGu27PzAg2mDswYGhDX5LKNEVa0A5KET5+a4GUlEErZcTnXQxftxdqNac
VpErtbTfqJdMlSMcyEevj+DD0e63wZC1bkCR/ujVJgKhmz76R/bS/bwRUYGt/fQA/hlsEGesiUpn
KNLLRVo8ttakpY0DwDbhfdP4zL+8FnG5PXyNndjK4ovCuyL8fR8Im5ma1SDxpEv8R11rgL2rGgKy
ZWYMhj0YiJDDwczlkI4BUhI0g/U2o45yuYYQtbGeZJjz4eWebWW9vjJZWvr3cdqo5BCkiq+VUAS1
Q+df7YqbieoLSWn5/Tkotyj3GcTKmvy0pGvhuZHx8/uf6UuKpu+THPuTFvOyYeaTDSVBZpgkogS8
RaEiFQ1yP6quxlvFFL64tqOSXPv1gcRuYbLcK8hNuOj+zBiojbqTgP88jiHBmouLm5V3bP+BlV6l
aerdJ/LTYUZ1vy5W3EvHqfod9bQSqTsCycBvLl+Q1SPGoMt4mFbyZO5fJx2zdfLHH+2KKmAev0ut
jjx5UEjFm6jfSEQTP0AgnMZtl3+hO2sM/ERADyIWrBKiwe2PXJS3qpFSHSgaNuAwabQCZAjL7CYB
eQJ087Pdvo7x+cMrXvqOfTySVvvEaoT327cMgoqavSfVGSVfYqMWdDkkvLrwc7w9K9/z9A6AaXDd
Ra+uzia2204JL2D4SkscYI/EttpTVklumWJ+PWxr44UPBEHm61aT84BkIawOApAobIXTDXzFTcdS
xEbRPvJYTFLZ0WZmNJSzsdVOIYDc1O0SAx8n/y1ej+ujYpLeDCziIW/Zl1FBFg8COgsgPOl0zT0/
USCCTCzkiYq5stmLtsXfgvT0fZJ6dt4VZ0Ed1MLeRLA7Z9CulGFew3KZ5HiIeUZeW6LD8Dvzyoyf
TnyHFrGJdXzK2qn2OCrh+X9pFzYV9oBcWctHlOhpY07csbIjK4zpXfd7B5ustZk+U+neNAVNp4Vp
UyljI/9rlmoKWRuSWFOWoDJVgE00Wd7hH7FIm7/V3utlewVQg1J+snPAVRusK71XxoWTHIKBKGRw
lE7/0275WLfL+TJiOHPveqlKfp7/GQDYJSqpcRveF965WCQl3nbsffv3oF+fSp0qbto91TV+VY/W
1JF5EGJ5yze3kvqTMab8vm760K+AzXkP4NTxrLmBeemvOUSHvLPf40nC9t5/oetHw8OznMrGG8uw
804WngsOcQrfCBCY+geaVglDeYoRPCAN1cRXLHyEjq2RuOOrTyIiCHSA3DT6ox2vC5uJFztQrIzu
Nvi2ODU9XH9YY5PqsAHoyZNFv2fog1Ex40hDspOd2flpYxQ2ABjnSyiAlV0+yqWH0OsSByD6ZB2j
wf5mBgqmCbyv/aywCmJS2PkzaAmnjCxwxKixF1Wp83jw5HeDq+xvHdBCDloJt2h9yEmLd+rfVe1Z
8u/djIWQ4mFJFMVlC+YafHdpK2c2gBE7sKKCKS2lMtSbfdErl3u0PI/O3/4uM5YuTS7I6aAQBiOO
LI+2tmIbt/s5ncP1gYUEpOPKzEY+iSX3Ne9JMePu5nUBk4NlBLEBS/KGIL6zr8N51qZwFzqVr96D
df6dqMIYBD+jhAu5wdqwADaE1XIrJUEBFbz4IR5ds753n7F8ffmZlYx+kW586iT16yce4eJE124F
MNgYOHAMgGY4lBI/KlWN9kMFvVhWJMnFO+WB8VKCrH9Rgz6Md8kh8CR4wSzqB0xhuS1ID4adu6FU
PocbIKtinFHHv8ot6u/UsFbPzkUFOoNRJ0TeZVFCkNgwXrbzXTdtNs6eUanNTevmtpSINKOqYHYf
1othpGwIOdVacjcK2miAp3EuD+3aG9MQ+X7LPtiI1hdnJb30oAypwMlgHinnViFLIHngah6T7yEm
pU+UbQefXaqq+V+Gt3DWh0cq4FZkdy+WTf/KeJuKuAulcSa66u6XXObnmGMryvuLaSv8/kBOU0gr
J5YMISpWs2ZqGqFvpAsqvKP32T3LsfGO1mNy4Kdf0RquoUFk3pflNa3yP8It2NRhKgKsCMVdpJpA
PwQeoNE1ojhQQ74XntGdwBcgWXga5bJcNjp08Qw1NoURu9xUU6i+CXuIOs0wAaJoqTk66W3uXKwL
rm9G+KpxDso5/ffkhGH2V10RbbQ2rrk7g1zg04zlxyd/wbgPvLJThCykVO4mjxlC9uPsWJM5nlAy
AEaAzN7y5hWzwmFJ0APprrRu31w2arI6JL/X81c+zTDiqeLUyZyPr4HlmCz/95u360AwBNuDpn8Q
mCW7e7Fe4mMV6Ox/bYtVI54w/0YjxQPTBaeL6oG9bJANPVCH9W5ZCTwfNSGTPOYBwJBAeFJJ947R
KXgyYSh5DvM9it8R1uByGFx5pOVMO9r24AGxJEbT3Hpoe/HZ+8+IiYONXFqFH5NtyiHwU/eJO8Xi
UWyBTHfYjBjXsL70fhwstWC4slXqiY+ysEjl8iGtryv+7GAMKiJO4dxsi7kfEudMD0bpAmgw0DJE
sz2ascVppZ5dLY2ckDKbpoeYphNdP0LMzxgL2oq23SFSTg1YMWiUtga9nDOJAqdNbKNJo4mH6kwU
LtGDIDaED3/qvZo58zQrLn+Ku4CubcWDCuDfdVOA4uMvpgIMNOa/ZFqE1RzO9pMJg9hudP3ZfHMI
KIQ/DNlmEeRO2C9alXbSFY4NO/ETLWMG82m88jD4B/g04XNPsC8/LZwv8eAxEcTBy9Izyur4hYaj
J5xBmJOqLQU89IP34EnZWRzA90s/kBFkKm0OwF7G39lWLl+LojDXSrj70OYl/IRFAlrJOWJ5G4M8
ET6a9/a5gscDDY3Ywgyf0YiRMdQXA20aNv2gmu2pg6QDxoXSWeH1jRzaud3fu/9jD4auEdejh2Pn
6fKKX4DwXrJZ4lyizNSpOaFq/VjPgHj5AQRMRJ5cQzIHMsNdddDQ2fABUrF+DppVxDEhNo96M+Mf
BOxgYt/02aym20Yh4/naCRwwAEti5jLZttPmyVHtlU6yMuyzVKorJL+LhOj7Vp/QGlihUjCapAR5
gfbnA3QTbSCPjAM+z3WJsuuLQ6dy8oMK2iklXvl3VtG/RvJYWXQiV7NFgd/29GFnOByUm3lp7T1T
T5NQjmdHDlRo5tV+8TpPmp5g+UXc/lQ/CbWsWsBWNFZ3MAzPKwrQfc4rh057W4KnT5bWIqVjsQax
yeXNiJWFHAhj3MT3szg+BVyWfF+dlV0PKGyLGJAiuSwVmwNJQ/BrmBKmxyqT9tW5/uyDaAqTxVoG
swLpxTC6XrDNjxF2t1BQqK3LQf0jNBWVzldVXhrZZhWmifcDt2EB8UjfXw2fqFzjPGg2hoKcjHUC
gbRwVK4djfEPT+1AFBEK074tYynQKH14U+9Gfxx37KbXHHprexFL5gtuE4MQavwkD5fuLql8Jn6b
cyLs7st2UN12tjxihc8BfrE2F3LkYPR8BTjGNZt+0LDV3/rkUofWS8CWitaWuExQYMEJeUcKQm5L
zjdvLPVQWMK2my9tFZ5HPlodC8Hyt42sodSlLUFamem9irDyccrw3GpXR1V6xBzBZqNVQ7lB9sXY
SKCEtyqIiwXZu9QnpD2wQaWgX/LHo7VCyqwINBSDAcSiuxrG5wBy2KGDX/l5MUjMXHNghkMRPzbl
F6SCVwgiQTkntIhqtm+LWvoAhGXq+Z5vgCVWgc0W+ZtJ3Iht5W6NLdPZ562WPDYi2SMmlr2DHxts
UzXMCbPTeR2rzkaRf8MAsvtqmGqh7/o4ZPT8YR2bMKRNWdISb/0L3uWVzfL2Ru3BygQK9kgCNT60
3IwRVzTWzpu9jmbPLUpgu1gEl4mjpp/pQ0LOLf4tAkWSELoevBiK5hZXW/RQ8kTtr/p09Xvwlxw8
0Jg21R4rKGQxv7qeu6jDmqDeQPOd3710tQ5kjbbf5VG8+nUpEbRtKC9rIEgXdAofTyjLDADPokJh
I0K00TVe1ads9Vg4jMY7H76JzaXuaJ4w4vdGSGUWaUYPnibGpc0FP4s3oik62n6GddL8Vi3Sf6zU
4k/1DGKRtUsGCQPzoCs9oPGN3YqdRQJtjiD+o+WKfIp+iS6xlibtPzGCQFwUJNT2ynn7Xm19QAcA
Fad+xqpOICz7QOmCuS/N+LAOQOfdpl8JP+LtL05fDqgtRE4eD5qu4tQydlfvVFmSoEe7YEBdJQXA
wDyUG4ZusfnLsAoXNHr851lEdwJ9dfoOUizu8PTatUaDeFFk2YIM2OoniQvzJ9cvVXpJjHIUxsFp
5L6gK+yPKIWzoCTpUXf+qg/LAGOiJtdPJPRMMRAMFGKCyxpWFYDjmsbWHErHeYG6HaujETklFFyJ
6CV5aI7r2pWmInuRIjUFmY0JRTn/DlFCER2ToLDvp5U/DdtfNnv6CahUuFoTStgSqUrNbY+fglPz
0G9Bo6eTqD3YQ4bB76JJBPNWh0OR7kJO/n7BsWcKfLZDmDXDTifNZvai049uYOjn4XVJo00+XAmO
15bSQnbxHGZHV8t/1tjzub3aYfr+/0jsHWNiD9GgqAqhxFmzWMmt7Qq+XcI0SyJNuA2FVv2aL1S2
1qiJ51H7u1xNgOthuhNOtRGOGg2sHaZjrHRjfA6BboiAJ1i/ED+9uV9qvcfh+T54TeRx4SXTyaTv
70oiljD1b6kcAqqtdmvduzMsm6ZbeHKjtdd/0VuhTOKfUM+DDVa2H0CG2asGx2mTpHGaurTol++a
A+3NajAzpY577NtpRQ9XETv4x5+g3uNzO2l/JekDpkG37ShChnlK6OKpAuos0qZp5Ds2iNswQ4Ns
UN06mKmo5FDEDj8ngIpvxF89d38SxMXM/NzVJO1UMz2UuZrYYtr7UsgV5enMPUxd9iVGxLOZ5RVW
UGWCPlpEQjsL4BYWml3s/Q7g/UFpkidyj4xGys6kE4yCr+FMBhezNvldAp1Fm4+nf/XOIaIy+LeM
4fwjy0zlkF0uWgRsDGheRpupKJCgLrjjVl8UwS7FgJLstL1t8npbwAAGF81t4/eWb7dBs5xmCnOg
3cxv/9aEiqdgmWdInhjy33GlfkH63hoqeFDLD+E4l19yuBAa/rPDKtKg/DZALrI8b8pPttS8SS8B
refMSUgYnujJ/9nWooMZY8rI8aoGikPrVErcNhtUkviNBdowKoRKjoEH40lHAIPlM4L8qxWU4FMP
JwpkUTKybsQct7etH+/YLJuMEU1AS1c2hGDCE4xrnBvb9FcjOPOT2pH/gYQOrLFBOx0G43S1y1+w
9JJ2W0/IOYibgqqe5cGl4Qjwq06vaLK4yK4kaEVpZD12bksqXePhuvIOBRq5TwVm2EXC1RoGppVs
zHa/yO7iJVRMeyTFTSYScuiyC+MRj/9Oj7wYrYM5KdVNaI/JDcnQ/7NoiTLmDfjtikd1BPx5WXeX
Cr4CHHX1tnbbnPcQdRy12t6p1T2zWTx/oTpUC3kOb93ZuoXmf4sbw2GTS5MYN+bUi9CyUAMIP1jN
PPXK1/IfeAkVGEqme5FQa5k3zi0Ib6LmtmUUPbRvRVG+XvmfR7o/CMcInxg0uVFnTLYHFYFxnrPn
V0e+x3FusW87o2v61GgPLDNtK99n5YaTdXVDjBzqPyt2GwlshpWbTcRBMzhwAcBnB7f7xUfxgH1c
7PVWrKpJ/qv7G5eCLnxZR0AJ4iEPYJBnQ7g+XzK6pSOhz4V3RI3r2+rVqoIhL/ihOdbAzJcBo9Mh
cbuYd1R99eLssavvEzwALg7SKtBTAjYCGcLjLUCN0raR8ndXqpXR6iWIC+RCONrNJwliCCdE5uSD
Qg8rqLF30ZIPqRVMGfTiqHucPtExBC5IFlsaAdDhONkkOHw1PABpRZC+I0D4IoGTca6dDVF6z82O
OSeqw451CthIY/3NF6e7IUZ7CB2k6BOqC8eaiFt07YX/W0b+8OAcF4r2nU3uRDJWTSo6J/DtgmYz
f3ZuivR3qD9Wh/0ySBa5ncbiTrDNEuBFifLetVhu5lNpvEVxuccLeYZdGKPG7CfDXZZeFjGLBiCA
RvgK5nXIs1wedj4nHl/YfRXEzoHe8cGlJbtOI/IUy2rKkrCj7+00c26Gz04JWVstC73RbPypEgqB
LZgTQBmVYQskaxzDs4X1xW+XJO5BbxsYqQbGbnD+Xyh12Pa/BLJkHhgLjWqABzNRmq2/SCfYrMGH
ptKCa/sY117GbaW/vCUxVzHnAAetgi3bzyCPvsT1lZ29X/iFemVDVPR5PnU0Y19pkGTgO+o9waLX
dCqs56gNAPSjsPqat368gwWmuH7c9YgmtdlBQD+DIIlz9tW6yLaH76jE3uZAt1dNDRT7NhKnUKFT
q+dzUaysNcgj8EHW7ONjT475kcPmbzA/g6YQhzYyXQRT4PjseG+T18wFHo8+FWXmMTljYdReXIRU
Ts/CJUdIFEKi7qnYKH4dP9RxTdbac/xVzah9A7iRx9/jgI3dY/PH9xPBWYh4kHr08HvLjbt5O5tu
LGRHOa9D1aumeomhYa2MXorhnWAz2WOWBblUNOgctynOVZEGjSLaX3QpPiAmsiFk5xKS0dXZK0HY
7ZWx0Wdk22xtqYkux/iOFjvRtrIdF53h2lPCwoJB98s+DJkBIAmm5gYDOEK+Tbk9skWi4z94Q51F
Os46fSiAIIZ7RC3ug/awhm9ffF6zQe5TPrJcQFygZLunnUyNaddxq+kkdhqOkMqGgN+kZB+cxa7l
4/JJzOGiDi1YpNfvnoTy4Zy93S65PaI0mD2WMTjeZFKuZLKdBTWZCYHtvuCmV+SiJ4oo3hFq9HUy
tHrwNX1BuUyhkGXKTW7TA81dJPwkkbbBzpLREEZtPY3Wn/sbesbjVQMsMfXlsVehgfhXhFXABkV1
s601Q7EBQsuvgB/3sEnN8yEkX6zZ6kJCDQyKUDUxa7jzlKYODH8UvYKCna+JaBV7tmMuVFLwixQM
qMlUMCb8DCK2L6HGY3eB1anhKSwXBcpsXLbBH8p257OC8y/3dcyr4ZuG7A1rnZuNUThP33r2as45
13FIOpGc4E7G1wde1atNnlRpjTwhStfXhKLkRzrgg/QSUJgG1PgkEc7ye/2pfAyNYAPcfUa/QTrC
pSMd/qOJgIqS4gIgNONWhRQVidR6ECZ6mTYcR3kTz/5K0gRl9RPBazwMQDnf7P1yW4WT3tdBeqbV
+bcXPiFOsP9KYovZtinEVuWA8VXcK4gLhL8zZiZwDKVxYZQvoYUTOLfDRFqshP/8uJiYByZ0w2rk
+JFHMQfeHmteomgFhd1DDy4ronUPz/oFkIZStVVPGfAgCgmKZDNNUFR78GF8vqOHdXwAp7xYuE0t
3rKJTPd2hwsa34vGfWfWmSOxaA70yPHjycWRfs1ZnF3rrlsoz5srM2TsqrQwFzS6kvloYUAPF7ay
/W+5uJfxWeX7QQvNUPcLWDaH/yd5pCvICIuPl0BQq389EoBSKaNzk3tVO8+67bjgDYvwK4R1Dbrl
zvN3p73coe1ZruBJHCZTuEPjLkfuMbf67nOv1lTlVxkl7wzzzLE3T00dsUrxeECymeyrXDB666UL
qhNKrWuv/kTsP6RPrdR7q1Gzvfh7zLjTAbYNCu3BdQI84seA5vsgpC7d1mrJjPWZqi8NAufQWBUr
aT0Dt+OF8rufEp9TqyuHJ374H7YcId4MMHK+NDnHHj15lw250l73lLJJfH+GC4qy1coDawGe00kc
1fybZHXpTm0s6m2Uu755D5ZRMl35zNWlPsUZFven5fBSIeO2TLw0ZQkBPbZ4NAJexurpf6TRyY71
E1FLNlzkI62bIAnv44pvI7c765vU3Pg4+vHe6vxfedGDpoF4EDicyp/dOa42xT9afBeg3vX6tia0
ARkZxgxgb905nMe1IVl+crO42C1So7t93EmyZKtXZshzUyuUd7Nsg71Ka5veSX5sKJi+ixoj6SHH
5IqnHvpzIwbfllGXU+e8vKDK8sy3Xb6yK+PXT5vur9Kq2SsRx4OupsMM20Vh1aIgJqPaeuA5SVxR
DMnz7tfNKG8vCGbwA+pRPgsT8Hx46wU85i4uuQlcHXsVgyinxgltPuItNhOlJ+1PVBplfpf2+YEe
bw/IHoN4IRQ5On3MCUuGp2UuYKWC9zQIKj91RbWJBaYZ/mGaOs7NCiQi8AJR9cWT9oRuC3/pd2KF
Xl8RgsfOF5jj1XU/wHr4yqGGB4/PHBCZDCPJemRFFJMwQOw9GS9C+oLQMf4yth+ugBr4Z9ie5vP6
5yE6IM3OvoDMio88OlIHiyBouPElfROwZpYzzFwgbNjPn+Mw59ptVdMxkOfq9M4QvM+SdJ37QLyi
6IsE3OF/awHMubB76EqUkGeQtS9OTgXgSjHEiS04EsV1gVyS+Kq3QBv9xfT7Eap3ispStim4cJIJ
RjYt/p3LbZaV/DduKYxvV0PL/9qzurSNvP+ttl0eNYgcpNlkb0DkkKRVOzD0Z1gutdzecGVZ35qv
bsEqD+yM4qkoMvxz/a5ic4SxPwyRNtJF4VbhJHgNKbNAJP6WnpcDLJmvdfow4PspodMh2imISQ9z
ONa9COgGwqahj/t5edvR+ZQTu2/Sdm0UNobiwyIapo18wx7bGvnoPLidG+FY6RwEOsfQQjQd6FJt
NEmbI3rf0dboB9cZOE33ugm4zpRhxxRBYAT5BkLVynxC6RxjY0qvJbNyYXblcQSaoP4o0nKzX24o
0X4a2EwboVLDAc3/HG4dJAHFNe/Sv40X6QGX3Zphk43FtwvzOokAwJx/6/JU9FMJ4JOJggtKRnC7
ycg8gA08Qnw7HyYikEDoQkLUv8p4YY7zmNAm7xfOvvgzMrNCPY4Vc8R2NYwXmngYiaEtuWqtUAXF
MqNKifxZigADAc+eDzCiu1oz1gNAQ58dsS78qeQRFqJ0FNdQuWJdCQ6JrAVtGv73uIAR0O50DJjQ
L1Q25ZClI7lJfcuWuHnJ16RW77r+dQV9UA1QgycJwfgNzxYRjLuXkyx5mijQ62d2vUMnFe7O0NL3
NfSWhqWgGZGQmADocKYpJAqwON6VwuDSYhz/X+bSZiqffAhGLafajA17MnHL+ft9VadSH6BFcvVE
vYliibvQqQBpKwX2FCg1NyqYGgtxNt87nr6OvQOSFmlNJX0SdwoRu3VfaDtQdksy0VrijC9Z+NTz
lvL+NlIfU7cZRtFTk2+7KdMqnHEZ3DN0uCz20gONZ5VcK2dp9U+sJNIENYJMqmAWDEFC3JUl4ZRj
gW/yiOJSTbJUPE+dzpkc0i2O19XySEn7g2pb/047x4zqmOqweRhr4Br5JDkkXzZH2U+08l7u1bgN
Fn/XY/MKvymdW+sq61zlpu+DqmmiODcbI0s57EILcEXOCfLMpKQ8IHYgcS6pxwyD/5QwjIIOdLpt
qXVQ5b6sqU7HZ6gZvNC/zTBobjK1IdzRdOWJvL1ENeHJMcScDW8sPA/IP5twzO9HgQL/pU2uzEw/
NcimxUMa4rGBKgVyCFjBKiwQ7avOj4PhlRbFJ4V/52uxwbR60d2WLwAON/hroO8bxzF27mhrMXH0
wZMs6dJXdHnpeCQPWaDmM5K84rAJhlfhcuwfWm4jSte8NMyqjzDN3giH2T7NPz2ENnpZlPW/Q/Hh
j4mc/wMDrSwXXB4SPDBxgZV3Sd382HYrKh+jBVrf5d0U3ApB8EglZzfKx979g93U2TmFtPccaKko
Jgv6sX6K5bgdKpqE/brLgCjDiZo/9h7MA679tMY1F1gYZU6hWfzpqs80TTnWt31xVQdsAADOcCsy
t9l4vH/1dU6xe18Js3MoX7ucNHthqNPMphBktvNoC0jEvRlDHBs4UTf5kyHeiHoDJdzLT9LbFygg
05/uO+FOUrLDLZDOOV5eJZYtGXqFr+HWvUoYsrHAYxV3w+YVPkK5mny0TqpnQU6RoXPX82PUdoBQ
6bcUcu7VafKjil56qqhvuBf+yoMfI6Vz0H7nb6lCR8gd/k4Ivko6cGcDygQKlW9es1xNS1tEGVEE
BPGQAfn62V4+Q6V16gaPd1AUZjrbiXuqXcrG3QB+zqcmGSUpc/FfQUU2CHaaKWAT9fh8GQrPpRgE
O3YVXEt9pwnQBIsvYICRmY3vpPG6YVckSKjmBvd1A5solEWM0Mtw56TKcWf0HxUwEPhOx+cVkra+
vEx157jz1SLCWCGSBZy0H0vvW0sToofmZe8Anva+F9i/QlAWFHbuI3e5fwY7ubShgSdQpMJtI2Io
ZJDgNmX1jMtAtq/LTEHK0w5PerE58CBAFzFVCli3aMNASOozELccxmNEyIaqZZvp7LivvSdUCJ4q
rDgL9PWPc00Tkcrj36ocFf4esE7EVGs9FbgawR10zLjBQdwOG9QQY6JfDsvNAiEILX7uCtq27RrV
StiLINBaLe566IE1I6Ii7Ypx8+1mFGKnzzusdfohJ8wHA0YiFdFxBed5bgzVq6IsA8g+lyswnZy4
013LGFOvexCqHqNofel3DJ/9LzksJ27PiyVnUGdzfYWeQVnq2Rps3raTOmM8ovC30vXM/ulmH6Lv
+twj6qzhCsMwuhDJPOxuFX+u0zEewJqcIZFQVccIP1POzIiUmR0cW3Yn2Mg9ytPjydXUye9rbwcU
PbhPFOXwo2nfaPhz55q4WpgkEFGO4caWBSl2Vebt2Ms0QIm5MzoTya1zsepf1F1neIc0CD1MrxCF
Y93rMtiJPlvMeDjWYooLThmrz9ZBiB9ijxuz5jMIgl+7xYVkYxxbsaz8/XHmYtFn4eWVOSGPgb/G
p8yPN+T1GtYHLn1o7qaFbZn5vWYLKK+GunM65eDFd+NhDC68toYQKRZCjheOc2HDC8uqrQUN+2Oy
xmHzxuLq3EkFcTKe4I5ecru0zu91OOc9opEXBPyrr8urUK4AUNB566la9afVVg8Im6BDPi11vXEG
rZyLEe9wqJOMYtBFGcyBVnGequKjAoccbS7zVSbcj66n2c9NQCg6hvuzEmu6a1i2I84kzBRooYlK
jlWF/DE4ag1tq6gZt+e58qQ3OfIukFsibzmLltxmwSZIW2uMZtKiwtUTNqKTUJKKjef8+aRpVGOT
mFlo2ZCwxaaiZBQhT62VQzq+Q6WFOkEhXCM27f8zz5Fpz2AtfqcGFVsKMwqzxSbV6z0d3qX/E0r/
l+nsnA1/ceLmxpGBeXIqOXyo09zvvrM+SQevtdi6B6rYtiFfPCweaLA618gAZagBBYp6YQIUNr4n
6X2D4g4pOeE/e0CPXm6q4kMXgVQ8iZniqS3VvGuwbBh6lLKRdIjYzs3gJME0bfuH2MdrN5vB7NIh
NvmUgkVt0vU6TmEB9hDVBjpEM6cuA/pj9WEzZQURQYQxguT04m9mhTFRC1uVpvAItF791E8l0BwM
Z+phYLt1litjDe9v9XexRCVyfbE44/O2Z0ornYZ/iO+dscRo+vaMDH72/QrmRLusMA7QKkWjNn/C
Zl1d6/8E7FRisSYaS125EEhBQwlv7V8QI50e04Js4jJ4ATVsyja4ESUShTBYm9QtcecAdW4JVuVb
XlTbT3lVaIi3886hnrsrvlcQ1Ul5ArrNt27u+kZC8Y5XHlBOWYVT8PA4/t4AsR7P9/mOB5ZZquIi
Cl65GwxO3JUj0DlzavQx0qZqAl/3P1hJIEytO7K4thptsJ2iOzPfgeor9KXxuzX63VkuMa0pW9XP
6r7BYvvhMtlvZHK+mRxYuzrg+iDGqUxbpVCxHAaXw2jTwz7MwBiH+5/NnIFPnNBahsi0uuyXFHuz
IhudCe3+GXbHDMuqZl/g+K+21lCqekneqt0z5KLIGVtydE5RO5qkQHqLe4OrH37taMhOnqtJJlL3
+tm+RzKfvW3PEr4Gi04MdAlhFCDnBYBYN6iCDlc51F6LPfCpkgH3FySy1PnG1SxxElLJkzvtb7UJ
AzfE7O3QMbC6fprBvnkMHDlRNn8Ujhyjlmpz0DhFFmmKJ0RxCaHxSSstBJoXfvPimEk0s1WoBCUz
DKTpjRo/RwxSwMTUYgk6fCEX//FVCkEq/+csZzPqXEe93IFFAG5YIvkKgI5u8h2GDqX/8pNAFJGT
HViAcIS9oyCKCdstAlFV1uh6cldWoFifY/vohEINg6ti0EAVrv4T2/rYEob/CImxD5UkQl5blXcG
RLqX3mKEo+bQ7lbYUkblZB72YIX7n2mNz2llfpL4ZXwOWxZL3vFAANtE0LSeITMDWeU0PVKp6gcK
nDPvhbQhdCvVaQMhfPqiqG2u6L0HGOpcrhrQpB8UzC870hNEu44oZ0oIA0L1cGCS2c9mzRAVErq6
/suBPOpX0oZLHrPGHx3zaDFB6An3kQGLfKUCr4kpGQHEel94un8pObmQR0TgoUHMO85ng+Z35XnC
su+tFvRSXLAYCDo+qHODCBD1Z920y9xIwY210X8yzAotAwOiY2Lm5f4H1+wDiXHaNtknf7Xlqnm2
pBnkq2LGL+rgsxxAH7SLTFYpVhTzCes/5EFk6wrJGn9YEXtBQfBlJg9kIjsvfHWcdLkEW9chkRxE
RNSDt1W6EP0L9hzR1uApyLDx78PSELX0TX5Fp0eee+EXDvrGnVFL5PJ23q2Uped6n2NqWF9+dilQ
u0BlwS/LhuJIVGiIXMSyv8csUaXW6A78jznaQIZGaV8JYchI9xEyxaA7E71aa6Wj7OwEq2srZ6Z3
1eYvjzxoAYtpYv6Qizhl/IKKN9VgcfkZ5rZAOExVWzEF/fsciG/ziFai/989+LuG1J+VAc1pI90r
yzrVQdhoGuyfukEtIqffQWRf1crpuLORK5RR30DDaBNn6kc+uHz9fa+g/f46HFGZwP5SuD360iRP
QoCBznxYakG+ywcdpHPIdsBkKyqpkrJbnuXY8mBMPuxwJE1MtOfgs9WDGEWDW8WpvjYp0f2HtySj
fa/PWzJR4w1ap8neVcRMAQtnre6r0r7w30S7lEKWYXQ/a6ia1lLDIYm8KhEKkS6OjtYx+LrX0eB7
Y5uA/KSIfsv1mMR8qXHFTfXggdEYV/qJnSJeS6ZOKuso0KZiSVfMLKGH8tHWUCdpWYHycaGfZvcy
7L+UkxmpBH7Ol77jqDyiTAs+Sv+YRk0gBI+DMEvtbcbr2Os8WTNWsyqqjoh0OZCSV4O07zQjfE5h
To56AA5cPnh6o26CmJsv5iW2rQdka6hbx7pO06V+3PbpzZZYb2+4goVooyCGbgtdPD80hzRM4jv2
dHHbcJP+sAKbutI/s7zAMIuRK7ghMiPr5zRDaei3fAukxiQchz/ehbVcjzWoHBhkSsfkedoEFz5H
Apus0TIiBLsvK5RAfZf9PX9CNcHs4mOltS9Qa47AJzNAfeVF07vP1sNbJaSRk61dcrZJVQZ0mVrI
VgtBIkWMlmw/hQ5BQfjSoyfQtOr7Kzho8A1l56eiFZR4f6XOBgxPGqNM/5DPP+xfs2BvKt/LQYKu
4pixQHO37SDYteQsHqxrkc2FsPVBYAWjxZcoDl5cOa87hqKUjTpZy9CiLGccuOfRPpxlvLnzdGO8
dt2S4GhXcjXzmT5aGPjgcDwXJG31wHKmi7xRFSNcgk9wvYt4UnOqeNRQvUnSbFGiYnRpsAGwTHqG
K/WYBUpL+pptRHgNBriNkZdge6wEWNcaOyHyGnRnZ4+9TubKIMwElCLSGmBX77Gsr6OI106nXZR7
8JjZjbgsS3EQPfnkwDM5YX+rOF67KB1dRBW5otL9htmYlVB/6jDoy+k/Sav/+a63DHmgn4N6FeOO
860jv8URIUoDRL6zFRQzujhd6iYj4HyGSMTPfDlLjcF3xBurspnMg9Hiai4/J6BbVTfFOPoMmdHO
T5MDTr/8x8+VoGe24UBGuGixPhhd9vVvGEEVc+IDlFj66aPqWkQtmolwYfb6cpae8Vql1PJrWVQw
8i/T7upWuql16AdO6lGvpQq3OPTyn/spTud4OxkanBj4yiQSWZ1GSFqC0DGOXk89fZTw0Yo8cIO5
m+IksdKnxTffg4gi10tNU+o9/IjnNeFuwo59AVRpSaEeHq7ppu5tbGOBomyimxVO39u0Soe3L8bG
dzTxBEMBLU8LwIRmKCT/M0VlayVeUcJxzrk23nQ1ZzSMMfk5e7ZPnaeW0mx4loJxzNJbvNJFVF+F
eI61OFambW1Hntp6wqQ0dqijINDEs2H6QO8AYtIsIn30anXIycNuDekSYvwLh3ywaP701Z0ych1U
NMDxQAL9nc9PvYpv3FX+T82F9zNtQUEhXo0yhMrSPz4nc2gqq9PLJn4UhAyB0pWCBTk0SMmjjTkB
oHPuMXAjB/igAxf++k7f94Rxr7QVkyOL/VB4TQat0pexdxk/6fYK7OrThYk8whTCpn7L4ha/u3/j
Wec4NMNescS3SWZrx52IHugmOIkeDTk/XoyOHckvBpVsG4O1OcxaMGyhO5mZFU2WZP4z/xvjd+pN
du/4kNECmzwjVJaXqngEfOFaomY2ooomZStlacYVphiOlja/p/xAtuy6nEWkoR3WLBqIMWuEbTh8
/fgoqJKxMywg6ptk8MJ+pTfEyJFK57iLes0PBHd6wFZOT8aXODtNoWqh1NirCQufbtvTPe2ynvM1
1UbvzvAX3Q/5KMw+OnzjQVaSIHxrsUl3Wu5Qw/1XiQlZZQJVp1XfpKzaw14EwFlc0OK/OnSjm75D
fgJJMzZZnMFujH4kk+tiMwuResCCoJvvEVd6kHr0E6Q30ZSKEfOkate+XD0ckw47U1yQ2KjZY9AG
kA5rrhPoV6DEpeoPCUpP9PcyfuqQ2oZ7AaHcBa7TPz0/dmb/E7+doiKWQZhrTGNSNOKLf51cqXfi
BEMUK+/0O9f+sWBi89gyz7jejm4kBxDbYeTbpiE4+CP77SRTvGHjNN2o0CgZK9CKKo/plfkdXbZD
3r0QflZUnXRQFDKYRgUFfKwbxy3QodXoFjWs/FGxSYwZiGmEzBFGv3KOKSg1UuMAHQp9w9vADrwC
Us3YOfmS/TRokTyKGqKPjDnlwIsy4p9mK68G0J10zItavjzF09wW1Dkq2Z6PoIvh81N+d0NLwqR1
gek+q8HxWlHNbkribRB/XDB6A4wOH/SPjJ6f2OmE95+Il0ND5QmCWjFK/YC1zp7nQKO8H30iPN6U
0na7QQTeHwJjlD3vCnjD8juEWCuJwffHjJiY42U=
`protect end_protected
