-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
SLRINccuQXkXAciRd47IO6v7iltIlg7Zp5uk3ssMRZ/S1dZ/G0hyzDC8gJzL+miSkuykpWZnANFw
UnnAiNstZqI0gtBtkxSE4Y/cV3gqpa3CrwzT96Uy7eVy09gll97llj7j6DeEsQymwKf+E6CmpWqE
fmAEsDokGIDcdlknheVFlJ5eXIJsssD3PFjYWy6wUuoIQHTkmvX3v2MZM9wNYr/wWZ/APUcXyIsP
ojFnl5NfVZOF+hlyJo4FO2d4kho1fD9ADZv/iLSdybAosb2KPquKc1H9tTuouY6dnuHBsdAIeUjD
rAGH0GGjG7hNtYdqkxRVoEp3nSNbaw6na2zf0w==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 56272)
`protect data_block
zabfonKO/QLvM849Q5shIeUZ2Or0YyPQ41w5+Rirc8bMEGOgJKIvDxs6iKvaoViY7HKmykuoCZWZ
CKu8S5vRLoSV2ZOACRvfTceP/ZOF0fhykxgSe+uu6y8l+C7l9A1qnxDsJgw5CAFKWCfvLWVn8Hm/
n0qO7GHCWA5C8J4+LapSq8pljNRkpZo3iVGefd8VvrICtc7a45hhcnE9R/DcwQm/YR23z2YlNFKn
/jUi+FZsvTfUOYxuUjJfuu/5YAmLc6TJhzZKKPp0ES36nP9PwIiacSoSP1SrURLnnbUs5omIHyg4
ICmvVTYouMfDaHCpgz7OydmTer7xSC+7cJCXWcD9m7h914TMvJOR5JW90ppZYLG37vJ1Nl3Vr1Lh
0pX49vRTy1+z3KOx+6WjvXX8vYr5TQKS9EAUdUcngEPzEHHGXcLQbR3ZPcguGYWRncVSktOyRVRZ
D0EbXiVR+zxC7fMXedFbzgzL5Yv9S0iOnm0fDJcjso3tV4UkfmPR1KcVIuU+/vsqISl8fWOf++j+
q6LTvQ2BPEKJRC9PhQxMKWuPmgEGE1HXAeojQZHa0sZ9GW/C0nkR3aB9PputJ1UkeKRIwN0p59Tr
gEDHnqKnZWvmEfEX/Q+kaJQiBT2Bti3j2L2cporByhWGQ1SejHyTJaivm8HZA0gw4JBhcTKAR+Zp
vV4Zk3WShZchUMu8sWidTVxakdHNjsjwHGPL0Y5sSpDhWWRnGyZ02PMTVcJz2GKz2QFPHVFc9pdF
zPRbQ+BZaf/7kc1+ja8rTFZn20cwNkRi4IWudCqjBT+OZiUDbcwZRoXj3QK2yRYDjt94GlMYoK5k
2tSeL8Ayj9tlfTKe9CRdqr787R+BA8yjkV9cFRGnCBRYv5a6Nl32Jyc8Zn4y70Fjj20fg903NhHY
X/LoMIdF7cv+I/S940y66SbBGGOit0E7cVV0irWPGzRwu9ro+2JaGmU+5JS3zhxlCbACn1K/3ZBK
5ehqupD3Szxcyd/H9MJMqYDGbMqhRhuZQD7ndAsEb+vp0JC2NrI9UmQkr/iCusbaB//NYbxOl9fd
ThXFO/h2cqNvUSi/QnEslzx7doDGD7BAJaEdJUr7CJWdgyEpz+6e5y069cyM7uRPmKHWIFIIeQSH
rwn2DoLxLl/djNO5WZTVJShR9SdDM+TK0MX//+MpEkHQr5oxcTMaLDz6zEwNyyhimIYBZjH/kLWm
k9W7TGo+Yyl19e46g8vaUN47HpqGG6dj+7OkoCclDh03sWq4XC2cQfsmafUgs1MvHPpclwbeyApl
ntWuIXUTuLXzUT3z2tUK3pqln5kysYiWl3PE1k/bvWOGrE/jiimGFj6gYWZYUdZ8hIuyiXRpoij5
j08SdqQ+wpUFszh0neDmYN0eyovQGH8kbNzVIIw8MiDoZNmpo+txjcX4h54LMBbY4VCoNjCaZuKi
k00u65OXpv6UHYptf3wDAmUCjOXYTxFJbXREJOGbj/6Dkiac7Zmbr+I+mRb/DHQRVhuHf3bJ1vp+
1fltp7dn/aYIk4SLA13AdSFwNV45wfAvF+mN6X1tKBqAXKNwS7JoSidYyIgDD5KMMpcaeXob2xp2
nzOTnBHhBGwKN5sS0FQW1fCtg6FThecg3bW2/ldyYKACPYQ763AAnLMtHVSEu+yl7vWcNrJPyv5H
Q6hEwp3tfqJHNSocxXGoSx87x1dmlLAAUmFiQ+Ip+GVt6CAQaDccytNdiP2R6skHTYNPHeyGKE/W
LxcSwZUD51P7BYeob3iyrDO6LrJro6HQ9+PljfU69/vqh28/e6g7wWO2t1zitZXbxSNW0BrIiX77
hFvZSe0FJ2ppdByGTNr1tJ/hB5yEedfs05LigXYqfwml/N6ZaLiSN7J+bdar+RJJev1KEdlrU5BU
pQYyDtS6FO3Gmxv8JnTWeqvQ+77ZVKUU8kTSDcceRpqPUmuSaYL2U7GhMROelb9TYir4w4Lz1xCo
UC7dd1AXSxqHoXmEsy7Zhc5Yh+sX8mO5fVpceuOIKUEX6lJ3pJlykAS6QFiQRSKCJKAZ1I1agHnX
HtQwq+dlShFjbbtjBKkO0Au0umFid7ZbUgOJ6Y+f364eKoatn6adnsI0399r4SU7RDhG9oM517++
h/U1/QDZqou6/iU5ktB5qnnW/MBz0WeeZ2o2bv9yi1jlzI0hgU9WMi0HPdUydExWwW6uEojJPXV/
rNqjDHMFODIHmxyIP49SWIHIzyzO6iQb0NJpG9ik9+B6rSFztn/bj0kK0P7S/OBxZzjW2JBr8urV
EwOhUgXE6rGdIT9IXqRmh9Cq3wJxLU8dj60K7FLmc8mV6D2DjFWCwaTQfrGasuojD+u9T8NIe9Mg
fsbIHApltkIhVvRe8nyd17wa7/wrYAYKlHUrOHRbrHHLoEsIHDx+fijCpJwa+t4omwKzdZKSSUN+
c82VX7Iu3Q/5RUeK10Arz0O+P4qAo7ZnvAnqIn8i6VuiBuROfLwT31fK1smW/22EYYHAkhsKphXz
+RnYsPpFU9gfpwmIZQwx68y5qPKsIdc7LXyIZrHMc/IirpfOkjkzjfuKjRKsFnXWZFqYe/P1Y33B
VCOtGcvXZhZO1jPkLPT+NUKiDBJGyRt3A7HuHwFVDDcJlp9KCFM4ENT/fM2utn2AfWb18dV9GYHZ
8C45d8De1WqRvgwafu8lWLa/Yv28AIHzC8EbBS7rThZ1IXxg08Muz7CgRr1oc/2SWR50GoPncqW2
/fC4/FmNQGYMEJLa/vxdXS8ehSEiZi0ge3Jlx98gGYImmnDlyoYEGaXwfEUddMgAnMM1t7Xugff3
NgiPbLHstmbL4vdU4fcPd5hM9jU4MYCavspTZqLDaIaRV7/pN9v3qVwQAv8jem+MjZrO7PD0GOlT
RzE1RD+asjTdDO8agqGBEwRlqtwY2e2MO1aAuwq22T9T4vN4eWrts3LkYmvTg9epxtOjZCOi/hja
X+isMNSXCqhq/rAkgwTCpiJLedQO3P0fW9CK8PvGAgwM2JGH9h1NZghw7ojmCosOCjc0Osaty3oL
ss4O/E6G5c5eHE9Ne3xMaLmU7S1X9OJz/k345vLzf35msgRnXsWitjKOWEQ0RDBNaqFuFg3gsWQN
PpbKz1u6VBoMxz6ucDpWjP95caw/6k1Izqxz3uknkcqQTAcgLtX5F0nJtjwHGiWmKRbktemq/tMe
i03y3mVd8crZr3MVCEJAlbRgH/5zoB9oNfzOBvThmkUuF2MjiNqFUiGdkhrrlBzfuhtPTJVCdj2C
oDtMoglYENlwV1y2LZmtne8VEMq/s1C9uJIddlQ37LcG2X4/o7AacFIG2+JI6fjBr5cYI0NdeC4x
NIxRmSy1j3BKZRTUnnkIExyPeNph8hzvxWOU8vHweVPyaHmG7HjCgpqwQJY+SHP6m3PXhlnQm0fO
rY0/vjHDQf0zFbws/M7oWmt34QF1SZU1RaCddCevjT3WTTPx6fxyHBmX0kNPbS3FH8NnxIEuKqyQ
0ypFXEKUNmzmS9udCICec13wJc3lJNrtlfKdki+/H8WFrXXBSXoyhjhH0cYfdDwJZMfWaIaf4QsX
fT3ECvxbevN/FguHEvn+3dj69aFMuF7gRloIveqs9dYWm9WbTo6ACIwnssxoHA0Jp6IYwdvHVmz/
eYZt9Gc7k8wxKLv283xXPouC57dhmqs3MKVaAs1RL7JScgA5VMU1l4vXkQIxTQAIfjSdG3T81b8e
WoLCGC6xmrog0PeEl4eLQl5+ltmwMTluUICCpC6VRbrkFioeIO7ahbY5Ve2Ic2gZc1Mm440RBqeq
PVOFbbav95091aSfCLR/VbeRilfFVjBGjPomum6s2Zj43QyH8YpeyqvsQ6Oa7q8cgtzjiOxObTh9
H6JLTNDaqhPRsB4MdWYJh4RGZdhxXYGTOTUxlGOsx3M3e+MqWdBq2ZkCye9zNPr9g6n0Uh1x6se1
Q2JTLGDnLpL+nejoebnXiBtCSeHxBnBDSs2xgdO1hOlOtcnlhlPi6sIidNbKUnghmAoWZD/XKAA1
U6JuBM0DDGdqP6uCFJ0ZS63ZGRzYGRvR1yHG7qarzAgp94Y1sWzeywqDEPZk5dXXDSlsT2lC4RPA
1hFpDON3EKF0gUM5rjuWoknNX3l7Z+RscCWMxeV8bN5aSYhWr44P0yR9RTrUehB0BBUrgo0N+1xo
B+Es9HK74UwW6Dx1WjccAzPh8rkhJTq85DwlWrcf06XvphOvzhN4tcLnO/4/CG1aR3TtzspDfUlz
BW87XiqcZtAFVpyOMjOrRzzaS4DbWokkxTcveyjmgeZ8jM2jZ62s0Mqkd6MfXv7gsc0+Nn1nk/Nb
5PDOXN7dIsMwnMhGe0YSc30MTDTb/kZ6bxPnDxaE3LjHQqcdMtNHmBkhhhCCrn45zPpsXAAtEcA9
m176FNu94BdqFDXQ8dKqOzbDJgi72e5gGioNFqdWud6PrI2b5Q2ggUJ0qtxJ3ZZbgQKrHIPmhOxv
0JUszrLhJn1C+RIB2gfHCGwP0jzSGuHDTqfDrDE6KPTZ3okdbGgnoh+vxb8BOK1nNOAVPJ2sdsVT
zU9md4SnIoHrH1Jqs+absEsV77Tc6qAVRui4rofvc7LlMiFrPTMOX8h9jX2u42HtoTQcDh9oUDj7
LQi0mCO3mh7vhtYJO8Yrm6VSobDdfjIYqFFLTK9Gb65vo5iC5FYX72P5RF3BGW/wvV7TItutHGlc
taAtmBfsmSvPwwptjP+9myHuvspfQ3+T/k9NcL+kCwW0pG3MsSLUNzG8Pc6jmWtERM4CGzKWU3jX
y+m3Uj9i5+qzWNpHvKNkNfkNddmud/xe0MNPMT521zJZHTDswoKrxSBdYuekRSvlsNR+dYovEXxN
cd3kO/v+prG6mftfOR+8+X7HJb4whJJQ0JYdqkUnIhgWpi2vcR+/3jvMBMwUKCxmqaFFvhUnpcze
tT5d5P7adosofzXuB6iuD5vO/UGzxHIIRb1hxeAAfZ+3Ra/XI5HY0+5ae40wUxQocR4l4xRRDeM/
3Q55PZZtkYrq1TIj78MEYf/I/c88BPmU9aRgUmepDEu4NyZWkENXaLidTVK9eVGCKbb3KAFsrQSs
Tq03kvMWk+JXMZY73C/Nl05HYrkmhZ30/AA7bVt5zewVLZIGBBXvX2+bBgPg+J/CCA985gADxIwM
WPFG6ElC6nJxB8X6ARni4zvE6I9L2I/nEx1EgYMtVRTx1wZB63MFPHOw7YTM5SW6zUMF5pWw11gN
Nz4WanT16V3lsRk/f+REn0mJ50us8TsokajtFTnYWGFxg24i3PVGQDaLm0c7Hk1FEH8nUgTBwe8V
+oBOHwuAscTwcZ3WXFB21Z/Sg90WXZBUntCNPk9FAwYIIVCQffUiZh+o93EobZQOpgmunfKsSd5Y
BLfbysPTSaJ1gnYRxfCkv0/OiYnwo98L+/agrn50/R7l072J4a/jMCgIlpEokaYxR96UXwFbWHlA
kN6mXgdqPAPE3VVDnyz6dhq/vhhJqSX3gfhZwQy8MGVdQWHVWfDfAiLPDbsMO3+vQs9bK2YH/1N1
JxZqk8ZFwkF4l3LfnIZP/X/GFp480ygCwpkr0Gj10sBEZrwHQltNYJhBYtcdmiUxzO/C74tbgd4U
TPAsnGl90W7CUsTQAx/4NxgMkFqC92bUNXMOrasxl1CFLC1PIy4yD76yhNJXNp5Ang2tijjv0xot
Cn01WBSUUQGfPGuVpfx4FcMxG/bBhqElLEINvq4kn/cHzoJdaN1iiNkUj+wdPZxbc6SmioDfJTWa
0qv5+eP3VX+FnDO6bOmx/9az1nbpj24xoGaMW4IJGxnfCROCQkdgLgyk1DhqazVwtYiJPY0s7+Q9
S+lCtHjMvjJ5BLVTHcRDhapzwjgTvZQCl0h0Bq9eeZ01510wpNYEbCYh5Avg/7hvvIFDUXAIQHTQ
r64dnWcYEkUmk/R3VqgM+LteVBStvC02MQOxHpwaV9h0o16lnlyrB7zQG/2jaZC+CG4hDxj//ikP
ThZqFF23llf9n19wmvC2J4Iq+wSujd5Ftj3S3ER0VuRkWJxV9ZpgvCH4w2b609dWcYQ/4C+4879T
Cm+r5Gi/xTT/+zIGG7Kl8IiKQoZFBlwmuWqxzCCH3gtDaOreTVq9jh29FJHCH0oa7bF/psG2cVJL
Nw5tOgcaWyUsdDnDa6UW2OdeaQ4ud9ePPSrIN3gkyEhK41awOLs7QZ+NCgwXS96lQUv37uGaoRxm
23sndhjtrJ88bsOzXH6qlPtci1KQFYaQPTjWdg80d67HOKufFecmxz0y6XGTwVbLaBMYMc2tF7ny
1qLazZM+Eo3jFVaMfBq6sqZM3lucyUzYNV2J5X+sLDSPUmmEQEfT+VrrNTajb1I6A66e7bBrK5sT
Ri8jMKpWcvxj4ex6rrDgfoCeC2qhZmz8Yiwra3xf82VmlD9S4oxj2mkfH7937eWHh1iAkvhKOAo9
nc/GmBYij/yyM2U6vzSLFXDYL5evhTShj96BoKKpOkuTV41fDvbilIoGAVZd/lRK4dnI2u7yzqfU
7sDL90EDWu8qzjJ1ND36Fw2Xf2yBAGskhnmYv51dBwevqWGMbAbexh7RX66dVw8NVJymFVwhHnJp
r8iMwpyZhPZ1ZPvIpV0SP0taCW2L+9KEyM1Pv4vZD2CEmm+pH1WNr3zwhhBCk5mZHASAw6cVDTbb
QKNOryS2dlarbSA3WgtUd/lC1YUO/e5Ey4DZC+HTlzJn9MF5yo3Y17sAc609rDyaSfxkak4UnvEC
hwsroWHNVYu5a6HsdjtB1Bavb1OrkKVXFGXbyOAELVwOuru8ixdXCmkKpDJZ53aAW985jNSAnVRv
ZAj++W6+eFJNCc2xHqO6moEPqiE0idIxeWabPHI96C0VwL4iK3OTIrlgsXllbXtT+rQdSFfAlbQP
c0ZoyPCJLpHmyrq8emQKqtdQKRfiDePgGtSs23hHTDhSGlxW6dvtCTMy1o60GLxXWC5yyFOCU9in
bl9oZiuid+HLPnPoKA8zVzey5CxjMaMp+o09umzhSx9Dir4iqcha1SYVNi+FD/FrGEQOjaHyPNrA
zCcO4unQKJUORMRoFoNvc49hUHt6zHulrEMU/NH63UWGpPkQDxUiM8TsnfKCX8y8C2DysMn1rESR
EbgLWB+fP6K6UBJZp74xfZ0hi9JQTt5lWnk2eWQK77LtirLcrCchAQyZfaqNLGbIpSzmq9AzvV4K
51chYapJgpwW+7ewTfrodFRSzSRL/35y1LIn8oR5hhb/DWockWESjUzpdNmZBQk/ruG5t0K4FXMt
yu3CFobL3gMUCf9SEg5TCmfGw/A0kRAH84MiNMyXQDDzk7BLQ5rNxSNtIq7MgZ6pM6ZQGT5cBMa1
r9P5/E0Ordo7u8PokVlWkUnC1uHz4tr7uW6OXaoSZAGoCZPxUj61DVWbsUEYVdRpOXrGVdMi2a2a
pEvebR05s8Yjd9QPEgbe3vGGB5wZ2GaNLbCzbrtLSHVkhJhIaC7dJoNiBzAAeO7dB2yePCUrAqey
hfjMbkDAURB0fgrwuW226EtBeF1LV6Uc8Xj3Ml63oNBTM7sZn7KuZi6jxrazCMu+nxS3nLi470hw
Onq3yx8jgZFrjkzZUapXnqTVpE8e32ci94vFmCicvwrpEeOug5CcM+mfSbQRNHOQ+oOcWdIDxSDy
9/BJSdbwK9E8NwTHM2leH9k8cVlIPMvp+XWdG+4LrE3mkfYaft2kq698QqVMZ+2E0S23d2n/UCEk
84NsnKVkOShTnibnWMix9Z8ICzoAZKn7rBKH+VqGzFwnbOJkAyBb92F2aPWE8bmyp+xPzYxaeYun
MnSSKXp/1Vb20FQvc0MjXAc9OgZqeD/Zb+JXe+HFOmcqZu/xN0uniwz+OeOa3eL+fmsJquiCKXcg
4REBBZa5CTaVB6OKWb15WMU6O1vuwBmkgFUb7jmv6+dLfs0oCfkHHb3C+79HF99YvbRtsj/3DzEI
wRbffVNp4PC6KoGUwkFCNe6mEpSKZN+5tDHTzBN+L5fSdsiaoFtfBj2j6nGC+P77eS+HNVHoqHFq
VbBAmUPoFD9JQvthFnhch66gHeMn6qwbuHtviPeXN1NxIvcf8KbBcGDWCBqs84t5L7ySzl2mjgzj
VHnN2Wsr1NlYmVXPWQ7jAcl6FydHrsd8Pq1D3tHqvPOG2gSRQU9hHqLhFQvYFbHYRd7ILL7Vg8GZ
nm8II/fzX2DeYubmbJn2/4V0HbwqiN+EV6TWhriYYGzNlMsjCp1K/zSRio5CWcpCRigMcaiMyONJ
sOPi/heZTVoFeJrVeSCt5QChhKvvZKGJyogw8WJaWKHWFukdhBLE49Zloy0Yu0fKy1bx6nLeL/YA
71luhfEiC2yi6L70D9rg7GxaribYsiYQKBFSF0r8dYMnwrjHVM/oY+Amm0T00SAUyMJx0f6AhPha
+9V7EYVQpxyVUucZVsOv9PselVL4q0PcgbdJaXD1/vrT6WjpisxXAGIBnNjoDhfTTYy+X586iNTZ
FjiV2K6UBc2c0HvNq8NSLSZBnc345EJ5aM2nkKtKH2jvVl9ERb6ZASDWOuL9ri19RKqJKV9SB385
k/HJxA68TTHaZ8Y2BS0Wp8fAzpP/DjvLnzd27hKxsXo4lHzSZbUlMbQ5G9bYOz2dZtu6V0sycnLa
05fe49idD3e3CYA7NprxzjbQngJqFAvTXpKP8Y2B6drMtVYuhId67kMdZxU8wBEwiTMqRZu+BCoM
ci40b15Ul3rPynSQ4rsvDfYOeqFCLlb2O406r4y9fXJe2gyNt4de6opz6IFy7oZ/o7NjF6ORmUSA
xJWao7RNyoHA4sSf8BvW/Rd+C/SsFz2Q3dx0L3kDWswWAJgUu7SCw9G9NSgSuf5M64DVnnXMou3M
CBRelCiEeNEeofynJLEiRvbYL0MKEKpACgWiKFTljqgTgvmD1OGkeng5SvZiJr7FBsm8SRpuhkEe
ot2oO0RHdSCvM0TsocsJbhDCQdcJrUO9f6w1xzy2Nnw6o6gSvKgt9Pn4cajo50WPQSTRp1wcXieT
GpL7yFaPCHcgWOFJAhEEjlpT6b2a6uYORUYpFpAnRDaye04SX8vMl/x+wBHDsUTXHmSTGWRAZcPf
Vp9uwPtQKMna9dLLs6A4ePqvCQHN4HUfdLRCfa2yDh0laihXAYC1wbs5CNgF1k1J/ThJhiG/gMqF
XbvbKBMvxe9H8i/6p/ww8gd6piyyMAN0m/fgqvcNiM2w1FW3W3o6GlWMbHT27sRFryZ3iuuSzHhe
ab62psjJ1g68+CXm0EOJQiNqsV9KO5dczzVWULWAK2dgwvu1EMqfPIMRzaafSb+A9QcBE76V5iyQ
deEHTxt5EPhnhSakb4s1lp8iCmvELTCsGtkflq3NYIvBeolMNp3AZ9iNOcumuDDLpmxx7N7jYiLh
aLO5i+jQgtAPje5cxnmd6FTZLpzZUxW6isNnEBJPeuwa7HlmdsezduLnrBf1Hx/bqTPKg3coSuwi
wiYlqKktUhlJ5tZny9J1RL8/v05Iw7rpo5GQiSj/ebNz+Tn33xfnXvitGNbphb3FgLPHdIHKIO+P
+sr673ZKJxJyhOijBdfp4SYv+tnICu9945Sa4BcXlQlVq2Nz5rbpRJg9uWuvdJKY3sIjnBeHvK4d
lGZXZNiFZRPDKaiRusgeVYPvag/QVMotfBCVZf+LKnHJx2nQ1XSun3WEoJhPxFwDkuBLVbYD76tJ
XgnLfAzGUskmS02cEmgL12AMClDc8KDSz1XzCK2Uf5GA2RiKnVPMiN2t8lilUOVlfPYo7jzdxTzt
08g/ItXcmBd4KyrZOqrrC44QzUWUUd/WdxxWN6Jb/udOGLmH0QH6RqhaAk4JqlMdzvueYWEssgSI
E8tYKISO0OAWIjOkExas2mYAugGX4Geq9L5dBdNMXNHWA+ol7hATo6yt34Yf1Arsykb4QgtOPo33
3TsAFaAngRI5AirYrSI4uQvLyc8MEz4VydB6dU6lzUJ54ZaxW2pSng65VdZ2ZO6bzwdEcFLzrNX0
qMcg/APU64Sgt31fJ18ybsiLhnCs6FApv17+C1kllOqNUQRqD7oKp/hTcv8t7ZEAR6Q5GWrXU0kH
tXwYh2h2BhMmte5cY8e7kQLTGi9Y590n67vYfKKvORygy988Xj5NrbOCnrxU2XNkXCir9+MCeP7N
rV7n/v3xQ1MFg9iHvzhdEaavwBU9fCG/Sx26EcU/CFfR2AGYpJkhlsGjkIdbtPJyWDL1bOyWqTnr
W0HM8XKM3mov+903QXaOIcgyLcNt4J3IBTDPK8QgJGXvdmiVOsoMy72kbDcGoV+Zagl9cnNmtZMb
1cpaNoMSzGlWqdzdmkRJktyfmyv7jt08qSuvx/lv9tTPX9DDmnyclISMH+JWnMUqGFvBXN9o0utx
Nij9RME8UiwSvPqP55DP/KjLrdw5YXXZeMx4Wf4ZwWU7fYe7KLldx2LF6Ila1i5qNECQnQwK/QtY
AcVCaPPw6i+c6nreNmkZEcTFaLZBDynmh1YtH2E4O5ZtFbTa/gUpmsZGV1SrLYNEjK6YKVO25Pa8
sMwqVQVY/Nuz/KxpjOwjEA1pEB+DzkVO56bydBbQtSy9ZYBRhxD3izO+iJv4b1s6NlxheQZ75C5L
VQogyLEJJxIf3kfDi/YaxIqFpifKYMcv5tWKc+kvvFFL4ata2h23AuRl5MEP84n8IrJKt3AnC0Kq
WAHchW5yQ8ctDGqLQmSLq2HroIg/z8sYQL2q4sS4YOfj6MxhKOfx0rvOUActBG1Rfv/8FN9gf6yf
VI2GTCuWqlk6Bz5v3Wt2YF3lsYy0eOHNIcf/jb4UdXOB5LbVBHVW6tqKoP02RjKkZQ0qcNxhj5sz
YjeS0FpiUI8phoClMb/3oociywCVU2l/s1tOhbjNRQUqqZbZ3uNpa6p1D2hCbYL/J9g7S9zZCKrf
hhIm5ROUJvmOLSazdZVlefuIsftcAXHOMn4Rv5PVuVGh4AlaPIltlpkfLP6Ps11VZErdnoZDCBC5
As0cbSTORCC5sGe/gcBOI3D5UT1AEpZFqwK0W1poTZH843kotmcsC+YcgA7aXngPMfx3iwY66NTF
P5rUFgoUYYn9u06+N+1h/hhbtqtGaDq9aABhXCPjGf61SYhsNns81RwIeuyogKUjdQ4u5N3JZ8MH
PY/Y80TXAx+2jWDv2InTT5tSKoAUwHnpdORn6N8Jv40pQoZdpHjgjgYAe8udKNlMsKEWJPClQ5//
ybJ3KhooXyE55la9LL+H3I8ZPlkUSEYuPVVl13VeHwYpw2BY8My8EWwfrlkQbgKWFO8+T+dP5rrs
Tee5/jZu12ReOzuuzdBbTRCTOkkNi6J4GoOkvLQzVeVHbuXRu0q8tAzjL9+JwYWxp/ooYZGrt//2
BNcdf8np3w8b1diUGzApB7+/LME5wlWaG+RP2q2W3iWyMkZmnz8Je4nsiy2oWFupJLwl7IzlDz3d
tq3tFJUwDFbChjTl433C3/+EDxQ4vfAK/pdBdrmg4/dQ5LxKnxqe0lWrEDV+OByXbVZLxIVsgKGg
4E2X3dKYoE49SDRCD48jNlbKN7BoBQZ+c5qe4GvGUHUKfFInTQ7DHhdRKnWv9zWgYYNH2Rr3ebmB
nG29+3YJIiO+N1YW4t6bgI7QD90vlFbaK5Qyt64qzApXUHtzQvm6EOYx2YNZ2p4wh5XS9Vs3PtJ4
K1AQoPFyDlJjOBbtcBCc6m0f9wIAHxKfn0Y+YN0mW4zNk7xa4aE27Hz8bB1SsV5qhO1UREFTNaDj
oqenjDebovuHg1kLAVWrIi++LtNjReE8lf0uLFwHgMTYbeKFB0+bjKdgyjBRT/M0xBVSYqd3Ut0r
+f3ZTt1cVqFg+Sq7FLuyii4vZocu/1Pr3vwNdd3mZ9++29s6LAP9QnYbG3dSmsvyRtPIr6hKwQDx
FhLioriNNvsrwAFYL5t8Kn+WzpArMS1lxQja5L/KB70w8Fx5+WTybCnw2GhRyjPMFs0rlaY9vacL
cowHiBA5/2zRnseUS6oQaGqq3h2xr+cG/mVVJtZXV8j+hnR3OVcICpRSRKhWzCwNwSru2lxhFwLx
u2120HOByQCYv2AuUHrZxX/xQmuDuT1fpiclxbnmkCl0vzsqamSCjoJxcgkK5NyuGUYktunjeDlj
cTkYDbWqFYubS4yW9UPOEfRF1HMsRqXN5bL0DwGlLCVePD/pgTGeut4OMILZsStezb+/INh8YN3h
/i+09UVRPrYDwjICVi2RwxaH7BnDebtyOUWzjlNrgf8lcXAmPtIOpK6g5IaDf6EJ3YQuVS2j7IG1
hu7gvXfE/O5MkGAb6K3odMwqQQa5RVcykFzb1gWNr/JH8tu6Cff+UhFdtanc6oCDaNOwjwM4jpCU
Im/6RVkrziMY9aJsL0ALbm0+wEEGxfO0RPxofLgCk5/5JRLMpZIDF5Emsj1Svid5IvpbU7Uk1vG0
fN6wawmacEmzX3xW8Dw0EL+PtQSdiFD9Gm86zHJlotk6hFzI3TMussXGW4A+OrsJrESQfZcp/cFd
behB04M0bIwYakHo0qL02w6DalClmEoClueAI3R8OAoj21JFBgRawtXruWhAbbU89rvqcJO060lU
PccRTDI0ARjbvEWPqzxC5VZ73Mx7ETUTWJxqMs//M7QYBiUFNEW8vRlo2JaferQ9qpxbx1yn8GR5
ruO5FMPUOJrzmF+/hlWN+9y8qyVcPh0lCkkMPCXEwlWFPkAeTdcSgHvgjskA7YK6zqgp0VV1i+I2
j1NlUQj7lVFONScul205q3k0XeEASE7druAPFXoFca6182e3CdnvRiyaTS3su1Cc/tUUVGGHWeWC
kROZaJqze3dWrDrwDP2EsgepP91UMchCqe/UuHn3PxFbE60TO9E3CK2xNen2crYdu3e/yFi6VC0a
Dgr3JodOcE/C4IbPsmwOv/BDi2MzXxk7e7LNgGjjaJ3LzhKFbm3Pa9NS/SESaHeRxaGw5gPWCRCA
CBNsoJcgP5n9cXYtCnC+EYj7HjvmWObeRx3YXBYHKnUaQ/p7eyTK5p1F/J4aOY5R7OxEA7foCyGh
Nm1oBv1ZETJZ5KiUBGbMkMXCSU5uU2LL/iy+gqX+6J6kToZWGczKMjbl5IJX5bBumeOdu3NoFYeX
/jKs2rbT4Uw546Ry6aoNTJx9UQq40NchUmzkG0v/l3dwrVgqMub5VPHiVwI7nMJ2v4+6RinmYEap
bDOCWVzaBV/PnnGXVBngr1FfVN0x7WQHEPGU9WFBl8mSiSUMUi9kKOBrxwC4kn56EXXWf2mVDYoo
x7/EcFkJBsNEihJ4nbAvwMNwJ9Xa7rgTbCwdlK8Lk6MUhgeadRtxmNbUHSlr2RQo0F5R2bzkIN/q
WOnJ3U4oJF0cxNf3iSNOi0xPF3PDCxKJe6cziE7ui9oEELZfr0Uc9ortIeGadw3pQSO0yqvvbXW/
GlB6eitSvIsnZ2RlFs3FXiVeO+CPm9dUbWiWzrHYiPPTl5BTfM8LUPEvc9cNLcoYxoqz/Kr0fCdL
lB4o1rztbqRadXzEaISu37E9NKghGXdckpbDvW0LBxskzhnDhL1DdDJf/PCoSVcdIvDqeRKhj7mV
526xaUCpOP9jRsca9nhViFdKL+GdNV0y/yMI13PPPdm9D2IN41AnRrz3d89yNKhEWJTNnqEXSj/M
8eZtd9ioi4faOCSZpydJnXdw3uHuP9NrsNfVw29wPdg3jQPvD+QIgZsUFgA8XY/qF0niLoWYlIL4
AUyzKS/rwOO/y6SUD94MiKRyTTjRIHt7Eh/Id9MrcfI9G1GBvdU62xI/gM1UukYX7KtM6aGLUrk4
7enQIpfCNwinDhJTRyiZbMhfUiWf3Q5WdKh0NN/uuezRiMTIuffuREMxzU6llZgJWvDEg2VC9RlJ
6DWVXs0V+u1PywZYQWc/9j3QCKMAJaQ2WSGlYCM88WKbwZqyRIueKf26U46OMK3YdwfoczudhtDY
7GB2viPg4MErtc2iO7e68SzjWqqSj9P9GGPUxmxRk9dONbfVbeuENWACLDmABSx6+Tm77wZHvywk
8whKfNeYsx5myrpajRxs+fXK7fIDZ3+rW5eMF78x9OFUbANnZydiNZB/hW64igPaRProExVgckbr
7wwyjuyyMk/hPchhHnpwOUCoeNztAbWsFT55fBYSw1QvON7MCJ4s0TaQBokvo9k3eq8ck/spZJ4O
NiQjJAg/Fu/++rTADJs5pxp4aHub0ig7+vrPAPEBfZ55jXdsZDY8peFjCSsj0yJuW88zzD+uVpvJ
EBbx+pwwLb0Kw0DvLOIE4dssCk2xCnJfUV5fcvg5CCzZzR7qODomM0QtOGJzUOoF89/PLE1pZuNp
jxhP3MSm024tcv/oYOZyEXomJUCs467eLg6pFa1ZS3P/grsZ8zR/uR7T3gGbDuBXpIKC2N/q/byt
s10E6cQGamQ6WM+DBPZkiU76jz61Mws1nhs1/En5J0AA55PWcq0jl8X8kYmYMZexKYIrizX58Dyj
aNr1hIfXD9Afy8B+aWX45PlBQ0NtON50rJqxWtCfEbuqQlBCv6Ieybl4zYlHK9Ol3KpynL+t+TW6
LPeC4eU/sMstLMI/sIFzrGumd/WkYcuScBTR8FbHyFeD4gug7j/8V1Pe7BRZh3Xdcx3RKqlTPi0L
w3hn5vYSRAMPJ0oN6/VhKD74nYQU67EeosbhsFi3/hrnxE+TQ2DruuF6zSJvWbWyabpDbPMRQULd
2TFdRV8Qd4QCX29jDLQjKB9pCNvideryYc/1v6uclA6wIahMwkuSLMWkiaw1c7EI6HPUIZzvRZWs
6Gco05ESNbSdcjKIFoxHrzNUPAcGrSnkmiuVVisPStheU/LFGb1SvxFMSyRHJ3iKwWcx1Y1qcH9O
RQF4Uv1oMaKS5MfNtTYrhLOVhJpeSAU52lmjB3gFVQK2KUAFBEQwBl0xlxfT491mSlrSVtcFv2bs
4bdsuCF0I42j73boawMH9hMk/l/BOyQ7uqxpM7cTJQGpPvq2mR8k0bHfloaa13msCoL2fdAWhz9J
zdsnYNST4NR/QpM4t7t0X2IQ2tiojfPA9sGiPIoVdCyT0124+xOlk5iWqcvMiNvNi+sRowh9w6o8
LOnzlULDKYE/dy/g3SxDnFsfLQ3x/3XaMRAMrdqrTM3hdnQwqCv6ebaIWdFsucy0vnSANZOHcdee
5NVC6vgUKT0/Wh8YR0E67SPnVsZiB0NXQwlxeoRUMs5qYJd88Sue06PK9vVeDnLl3kFW756vR5fs
WC9ugkYOtEePAU51uqpysswZg+OQ8SeRbRdDbzCfIHI8SzKa29A/gpVvfeSkFc5qfk1gktLcAV87
fw3VTuYyNvGkIUlvBurQodgqUreC06TfCLasP0r8Y0Y3o4uZohgRMntzyFs76aOR9WNvSmEtwUHJ
7oEYiuuqP56SetpTlIfycbF0qGXBZp/yyN63mJKEhsqs1+gwyXhzmXSZjyq9sEwJk7JCTM43ON13
HyjoDEB4Fru5LY8hYrKEffH3Nr5NYLE9NGi8VTWyA6joZDV0iTTX1G5W25xxmKp6o5iKpkqxBZe7
ZHUey5H4DuEBG2jKGUQOizr0tqycNU3rMGI4zT0plwfPvvIJbddiRPPXWLdXZ/sc0dk/6ycxgcE8
UrFv4REU5ENds282kLaM0L/DY32zRrLepxCnE9x4h/YCDeTzk4V4Z65mzO2G4nPetlL5VuQjIoXL
6YvC67KLDSAud/lR1L3ZXHzc86DSqlSyVQNx6AWUL7gNYF71SH2CL6smApU7fisvf7OOlW54wEMZ
mfLO4ZSD3heAc8+VJLnFunb1yHRm0AQ2O/26gELYYysz+udxSl7aAn5GisTVJUKw7kLEchT5TzGi
a1msajPya10E4CNtx7h5Nuxbg40oFIaiacCS4AG9RT4fB8xF12HUWbS9aMFsP+0BaQju2FM6ICS6
JU+CWIoqeMy3ncY9zIuVruLisSKxiYocAEGxRZ7BZ8rMK+pjVpi7pAwoKN6zlWCjEpV/eguPkfjI
qyURGMMR3JAmskSaXjX8x8eSn3Unxxd+JEC/IA1KUvJDzZKWSBL1OoYRvsAY37GbxaWQEycI5NzM
l9OIFf86Mj++NeKmHZjhvp2er71gUyCIpdrE127g05kyYz8/mxTEgARVpNrUDFImGkynUBx00A1b
IrNdejxV+Xx5Dvk6uhzMdX8i0pTo3k4Fh3GfW1V5UD+eb1jf2NBNRloP+9gA1iZZk/Wb1V8MO9vZ
af1IjOtqWFMYV0Q9t2aKNNfx/0HHm2zjqPqkeUKNib+BuKik2iVdwsLUavvSZ4Ow2c08HblE1Xtq
UJvfVgsHpJLMor89mZqlfF1rl+Ot9CKeXK12CIe7u9PTldmZF2sihtXrYN+tMH/STpuIYWMc1vbB
ROnjfFMrRIWVSvXMNHDXjJRAiOtj6pHRTK0XzbRr8Oi8yaQq+MTHbBcPTmn0ywoua30OSVPz/9i8
g5LbgjE+wCKwoTySTmPtOCmKXZp85bRQzN6Scf1r8gv9LweI3w6i74ewhs9dxU30d4Bv/4kmAtYq
Css5HZI3K8tf553L5o5XznG6nQOJvNvKcBZdcdaguEy3sp+iWQlKHOU9KtIOkhWNHLn+LAqWr2RS
2iX9yP/uJT1h8EL0BCTETcMIPl9aNlCtlM6hxw96mJc5bOIyxK+NbjHCQOM0/u5TLSpi9lft2oiz
crl+ghPwbB4q9G16894VYJvGorhHNCn/XqUsw56wfnNjETcp7oztSBFlbAX+lGbNmR2JQgoCwDeA
y1zCKfeH+JGheVMPRdLW35LM5R1bRS4LZETZZHHF2r0xKwdZxrbBc0lTULL2kHpjS478MdqQJdtU
eqIKC0+aEMGYNpRg+ERY88nzGHVDLz/G/+Jv3v8Da4rmipRJdjfD9k2yGjOuh59HNrUoLe/9T9JM
8WVJaX05BUH5Q46FKkgMYSDTKi2mac7BVADR1yG/RoCszMarSwFRhM8Q7i/BOOTtEpboYQvDKRqm
q8BGyO+K+VeLOEsWGeBsfjQOJTRRpj0v/L1hnDgZ8itrggwVyoOGF329kA9ys6+P6K3BbhqJ9ip8
Jgt74rFx9mIsX0qVs7BW45k8PAjhbqDsL8gqXRK/X7GjhH7eWvS8GjqcelEZcOQ/RzEtKLiAoLYd
Hn/dEQ+Jqle5tqofFZ0PP8CBOOPFEZqhrAYTOwzRTQbJSWCe+cfFJsetKU5yvTziGZ6R8FN7VYZD
vXoRpuOoBQJjP0g8uVNYaMBs8IaDTgUpsiOaWwQTloWjFFG1M2hFCArUHko9cAh6uvko7hcUP0TY
00UiHA11gdedEJk76bdEyXuB8JZGQ76RtfMnee8Sz2q/WdPFNnrp1foiwO7WMHAVb/RlsaCZHZEs
4FeI2aPRi+Dmijq2A9O8kclWdf321mjq/G8Q+YoWRI0cNhKbhnj4+DIcuJ0nc2FqPNuMmQE0maMR
CprJSGvwLC9aimNszWnjQRYNEuOoJ/fV2k1m2dQK1DSrsElkNaUYXAiUSDWFZKjR9V64Gevd/wXr
PIILffEYmIVOBNreb8ASzLUTiP18q1KWwE5NnLCBvu8JpKHWb15vYljJSM7iWQAgQzsI9K3yFSxF
UVKT9gr3H1/EZie1wij2LmxWHOgBEi5Rlb9uy4DLODQeCmp+Ioha9hHxKP9cPRKwHC/450dMveZX
boTyAmB5icKzvBtZYqYuiwJkM+2XMNWxZlrB5FfLm7NOA3BDv3JhoAvcF9bpWxhayzYUm7VHfmnN
iUIgtqBWFBe6FxROXxOGc4PVLO0wENnRAkgk5T3ln3LhkhWmpFkscgOZbmdT2kQva3GvrvPVJScF
jCMSIVLuQ2o1JXo89tQodkLj5/+r1YYErCoMvkBwaXldH5OqEoAVm688hEGo80LHVaV5G3gb2saW
oZzdJMg747JEBncfogrCmy+BUWQG4SxQ9FI81kjzw5z6dQhWZdrb4009VZ1Kqpbwf4E7/3cXkP9E
Yvt73y0wlRBcAMkooVh4UdGD1K4+Wn9IR7Jdugorm8xqseS1JoPAXSwRdMy8f4lrx1FL0Ut5f5W/
4XmX/HFyFioRXpvcFgvJEFf8z69j+yRkEKLQzdW71fw3WktzgVQvTjBM1bgprclwQyohEKlgfhvh
cMBIOFtTDtk37+PB+c8NmQ1ZttKL7T40CBYAU7MlPRmP8ROZkta+BQxqRYJDLBhR7FCp1tJBWxKV
ieKfINkFfkR2EKc1N6Gn/GlBa6P96/HRB8URMNWOhaSfpk8GE58xRmy/bQgAVFxEeBrJ+19BzCxu
lgZ3KBFVv/1pBk4J8K9MCQ2oG0XLBTPUxRGxd7R3A3+50aGTQ7lmVCtXYyer4I+usB6yaA2Yny/3
piqGd9Je0YAbkTVo5hLV8QMB77jZNdie2mrumFljU6YePtfj1rcS++vOLnFL3iC1k0D0fePe+mv7
kClAQiBJvcspzAguf62HpGnOLlh51oz6k9lobWK8kuo2+CiyvgO5ji4DUr28L1N3+zUIcNctLjLW
ethWn1vrF3/5/ILG+uslzBlv3ssNS/Rby1IS4Areb7yDAA2pznrcbR71TBBDBHdIQHLA7RJxmthM
9ZoQHpnW+TOfmuSnnpEx9whLI9PNIOzV0V/dqujE/1qgHhDzDmGp22fEVpDXLq7uLDk9sN8LmLJ0
6zmWXALy0ijPKTa4jySwtBbzKfRQUEjeWOWKivZlZXngAbpoVFoT8QtlJNbCUoKFY++r1xf0dJOT
ucpfH87RbWxutBx1q5ftF04u+VxMLHkvS44YgBVGAfYHGk89jRjxbtzhpvJJxiWSslMNpSB16FyO
zfbFHF9sz41lc8jMZ4PoKnbWlJtjjruy0tYE22N+WDu9wC6svtWTgbg6JIky630YHJqxzwvx2iDd
Qt5iUXryQU4Lr1fFRdJf/zz01+CVIdAN46nxai/eciRXiFUaPk8vASgUmCN4o63KB6i3FbgCC9vX
0F0jYhAb/dJqVybsLlfvOdnKtaSo50sxpvfq0KPtAk7zUeTSG5/sZuUjTXypK3FsMCkTvyjJeUxC
Y28FkovXbZ40z8vSt8GyXPzo12pfOMkg5po3PnxnlN+lvaCMcEjR0Sx+6mzYnGlEXbY4iJQygLkE
8d7BS3SotzekVf6pzSF68pS18369CA6/gA3zSWLm5BuATFflWlJFGY1kbiCElXvh/NfHwCRN+TQE
6vU/bz79QoVON9Uixnq7Uz3Dk5O5pYtlfWS4INf7eFSMKgusjPYzEtpYa7mKCGYyyFh9wfyeNiKD
C6tGtDy+duiGnay1Az7KGouxBrr5NMZwd0Cl8QkOKNST8iwWH+v3c3FWFjxj/0Q3g4XgIYD8xhOe
/M9ccrRbGINGsb4bow/E8e+PHRJdxT7du/1FPqAyqGrdHmSe+k8AJrAtQPgefPbZBVRZJdFIngi5
OhbLJLHZL2pAOr3r6HeQJRzsf3gcbL+FOyzJMDhZQfQ7VTk5Hq8F/rhyq+UGoJGpNLiRMDbv+Ywm
pU6j5csciwHIicsYnY5XxVmaCout2uzu281vNjVXQX8P0Iu/4rPcmc3IMAETOJ6VMb0aUcZoNXPf
8tnUN/Ow6UJSzI5/7GR97OzoU5gWvhbYcP47cTIC+/0UZHF+EdruhvjbM4F8bgArC9Ql11kkbjCy
45DRK0DpSAFz8PLizKutO11G7PXERSxLVwm1rtz7Ge/RzFxPCd6TwodeRgo2OiHD+5257V6Hxrop
5shmsKNc34SZI0m3n+V3TVgf9OgIttMnDzMdvmM9RizvGECjxIGBpYRz+hahMz1JmN3cTMe5lz6o
e0ArSgKpvKDhwye9LGkM3URqE0JVzY/hf5wP2PMAAYcemnZNGkOspMi/umo2MZajQbaaQsQryQLZ
sjmrCiBT2NY4HMHlenCSchN+qcQudfNHcEos69YV5TFKvAZjYk18Vpjpcy/WR3nRg1AD5qpAWPPF
A+dHGmRMbME2zT2YRCqOLjX3ILZ121fd06thZB0oQNPw+bVURsvzBZVXAS4MrGXbv2/VUXz/yvA+
8iIDXaR3AZ3VjuxStSKPOQl/Iv90W6lBeJldrBH4UOFvH5vnJnWb0bDDcrQfpICo275fnzbffIcn
TV7cryRYShVg/oFVFSlEYKbxI1NxtVuy5QdhqG2/VuS6eaD87/k4dcOuYzS6hYxAY/okQQWFkMqj
hF0z7jE/DzzSRW8nFawTLIBK2QJZYLuYJ+H70vs2HmNbjbWVdM8U3Fs8boExve5kq9WlCSYc1k7N
2gfL1pUL3aoIt+hzXxX/oXZWDF2XELIhjXPAvrUbHqOKf8YKs9i+7bDKpAfO/0pJxwVEZRumHmSe
D4tUl7fpf3dTjUefsiArAGOaGytzLMCvMaHMnzT5PJiuysRJm3wANYqMcSb54nqZzZhWLWdY+L5j
XxBvfIm6DhiGORMAad1yc7TWWVdpefyqpMfi3r9ySxjgsrSykGu8YXnIhbsfA7t+71H04QFobpep
pewqO2mil7GapKLGw26Wcf9v/KDfj9k1nbcXZT47qhjQW4WKyHxindScXwwawhQpoZNwwh4oj377
IsBq0qnNfPUfLbxF/otGkuelyyuEN/SQ7NLSsYl+Vb2PwY2ALEI51m96AYJxR0V5d/R9iAXPwCU/
W8HScul3sKDoYmIHSPrDAgNC2q3nSJfLugMEZeS5UVCMlhrp66ThgjNRZeUNAG0YePowLwLW/SdV
lDdUVyeJ7LomnzTXgDbPBCyfxO3CWUsEgWER4hBeMJs8T3qo6UelHOr39fMQQVP6HFC9ShC0UJBL
rbDVcPs4p9mO5PZhtiptd0kEJYL+0OapBgeYi81Aszqu+xgcVUQHC3xPrMDS0lFeUZ8FM6N0RMQo
gKI5IKWo98AwOGBP+9ESX8G5fOKxc+TVBdzg8oPqOs2xLwB295HeZ4C3Hu4kgZh+NrdXZ4zqT9qY
5/H+DijztYDhE1oNYnvR6Ne9vA+6mj+z2G6gfpczXLAtotdjmsRcflp68xDmfG3pP2MNKL0xVUKG
/kuX9EgPvc449KSH3DPyDMEiMO9u+FqIyiNO4fnMBv1oTd9YznJPDTBVS0k/fDJFe6R098bZGu6I
E9PflmEAwAnm+Md+jUf62ui5Tl/K04wRVheK1gvQbXogkycgLgNV115u52nmUHuS2q7IGCsW7Tw0
ce8JGR3Yc/4IJdzV+3URsbKl61lgxsHBEfgQ5NGAfAPzA3a3Lhfz0acQkpqTWG5+se5llsN2E2yt
EUU93i+keOeiKOusFADB+3LJTbAbOmX8kjgYqzkNHtj9m13HOS0wNla0k/5rRVbRIG2KHav/cbn9
UEuV4WKCVz2RNorYInQUpVZg2HosMZzo4OQn8HU7qjWFIaA96vxfFjzZnjEaAhan1Dbl0szYPT3G
GXDvOlp1dPxWCCvFvYuKI5Dv+H0Flelvijlr5F3ZQLf2rArrBqHJ7KMyx5lqcDwApAvTBJ6KzIrp
FJ5F9FKxAOv29MAI+02sqaTua/7OrMstuRUVVMVHFXtj14ayha2kmQJeIKqIzOXuYJtifnVCHMD7
38IYvqj1Kbakxc8QYAqnvdXz+vssB5pZKWDtLERmFJLhBPVaadLnJG9UYaXjUZf8CGlyMTP9s2OT
+IqAb/dAfGBRsL4uBMprFOsl8vrbzJfuC4RhEV+dYzsZHhi3QaUQ/qHOL++B+zNWUIoOdW345QKo
cpfwaITZXondxjaXvRCrymJD6FdtUueHFlx8mJAW6lMTG4EIMWqutUPPivfWVMdzeIl8P6C+ycrY
Q/foTQ96pQrOSsrbBXXXnEW+IDPvg7AO8CCSMZcV1ktrCLSRtT47jMCdpBT+NbmXbtYKNjZJqskA
a79KxW3Xl9+TWwKu5mh060dQItfRzvlGz2foNG+cGrCIlhzvfE6/buouGzcCBTnGaG4eyBMjjvGe
Nv6WXite8pZm6y7eAcKF3ieTsAnsPeLKRhXMZ5ohkh/HsBgkrO4WGkt6rAbdr2X6lVyWm/INLwkR
TvRbpqOKth+klZMnjqatBAcR5nhAXIcvOK/dPCghnndMRNyeEBe+FuOyII7u6m72IQw7t6eNEGeq
rUr9n7HvNrc6qnqRv4QyrGLHbbvvoN56vqx309jSroeqN/v8dFjF4by+B0vi9hkGOYE7PZNX0nrU
snmAb4yJfYGRDLCEuO5Fhfav7mVFy7PSAKXVzclhIz9UTLdRRhfEoRfywcvelPJk7K30PIikCyEK
veHdfEpO3MtOtYLZRNndjbunmbzdLsPb/DfGnT0/thC7rqCzwjwgSZm+PDK6GQqzlxVJBB6nJcPj
XdN/iR/tl5Z+HfWgmbqwSKYBupbSbjl5+Syu4CIGr3VOitHAy6mdHblNxn3WjVCYvf+98WZrz4U5
iYWEkpqhhhhkMrjb8ibIXY5VAfOM6qZ6lm+0cURvry9HNVONBy4CdGiwve32dTPBsryto/mEFayP
yDi+bLK/7awQC+Mfhoy+onINOpPWm03LSuatx2oTEOTUfJqUc6p5GVFmA6ydvKLNnfBo4OSOqWDb
2bh1/t0NK8Mde14YIsaeV+hjDFrlO1BrSdPsWXN8xR9rz24jNfvoMjigugivZDZV4z/dOjcQqL4c
0oBkZnBFsYRz3ZeJy5wL5FxUhhs09rDM8y84PRvB/NB9LuMgUcPXSkzjN8KLyByAsRDv+UdIVo2X
SRnLflcDz5t+DV1cKnwqX/ikaMri/Lx3wcrwaZD4eNEuy0SjpJL+1GzuIooU7RDwInVcYf5EWqLR
DPqSCujs8io9r4EE62SLBTxOuFBpWQ4EHh6JSrxQY9G74VxuXDBF5gyWVaDUTkSU/m1BnhzikixL
HKWFCKv/p9cX4wPE8+HwtT/DLHS10DXRUSGAdrZNi2GeTOHG/uSC90o8seHVyB2ubWQ+IHBBwGke
2+69ymxjdUeKQTXHH5K00seTTlU1veIhaogv9GaKv6okyBPEMHw5pN+EPSyKnEgJqs73Uji49LPC
wsl/liryKUCsZ3A1LwDYPSNvjeWr8/S42hoJWiFQrru5ywBIDjJpPeSWfsoNZBK6qgNVVSw3UoIh
zxRkGIO2Nu46CaTWP6UQMXtedhzyy4tHDIZPQQbSnPetUi/nea1XIkygzbzUXNaTuN/f7whyGGPO
UhXoitkCThkvQZEp7Y3bFJetAatTUIMRk/mI2wUwvF+9sOWxMgkrxPG2RTBh0yowhyDce+zBmJu4
SfP99zpxRBBmJ1iXAoELnC/GyqUitR3CJ2/W8D7XSuTpnQuPUKVMDuY+qEqz03h9BJE5Qoko2NtY
Q610+4roUgfutPP63MdpeGtcOst3J9VFr6Bxvk2Kq/WlBogylrKiys6a7IlqW2rYN15Qeyokgh15
VYM7o6khOnn09QrB5BlNRys101+3bs00/Gt4N7cDustu2l6/bWaMAr9aatFazWSJPb4tdGztkDFR
W4MHv5ECr7k2I/QiYy/kl+XZBnRQtrrYVcQrMO74J+r/05q+MG6OAPBqoP6g057xVV3U3mRH7OBt
33/KLPz1KNKSwfaRrMXeaK2s4ZBQEEBdwC1cCR2zpZLbBDLXSFDixTX/uGWvwD2qN7XHCwSzkJRg
4tTy2SjpnO3SOOdA8yP3tV8N3Z1hG71XpQ/XD6CJEU5XWScGgv5/GzRA4oiUQEowV4doV39m/4BW
WlKUExqvTqHrIriEruZLmZYYX2Yx63R7stKk0ttDoWipGgXf8P/zK0L+1UBOVUHciKa/eNdd9o/H
3pTNW0lGfiLoujaVsnfu/31hDBecGULj7vhOeV7OchjsHYIlikq6oc43JDNblzGFn/RHp5+UMsXW
6sOXAukM2nLcAp2Q0MtDu6u6ZnZNpYdGTEsAqawMKupsmsojz9ruUakqGWO5+gnIeDO+Rrkclllb
5opp3oBUDBUzebyQf4bBxgpKLt2Ac3ttFqMfBkvPu8WnCS/vgQXdq0B6EDOoW+7tIF+DtgcJXFux
B8S4w88zWSixDz7/tB/bwqWTRLBcYE04GmkdfoQonEshhDkAqnYGezkpkluPkNeBXNaw3w09UaPt
Sw641Hzjibdu2RRBaxvDIlVulCw5KnPC73JToJO6O8E771BtAvcSGx5ABpkRi0yn6eXscfY+OP85
QK+GOaRFzgcDKghdasH7F113UqZ2I1FpGwhPpjIWJ13xXbNHXto5N9Ki4lEpXY6ChnB2Ng1zCxIF
JfHwgfg81fzPON9UxRIhhtVZZ9LadsIsvNF1fuC9dzXERWnHA6Yj1SHsRBCHNT0pj9pUnD4jHurP
F0DdU3Nw5/GjOCLNj8yG7eyTbqfohWv/srzdj4K7FN4wtVRLuHCLhE7OJggcpN5QJeRkjv849e81
Gr7LIPufsgN813n58w2cV6prSc/vKFPpiQ8n6J3SqqIs4t7YpBnuHHC7JsI6qX9utKO+YVnujquO
jSmoHOl2rgVIZYr+vTxtKCQG0wD5ge99DoEAuX5dYGQ4bTF0KHffUZir9Q5iqWk7mt2lXKzTS7Jl
XoD10Jg/i8dkfTh8h+jmx97afpEgDkbBgxN5YCZM/e4xzbIIEBLzeNCh1tSoqVCrCNV4tjROLTGS
cViZQEHgtl0SeuvnT0NhFhftnNjEwIfYXFN97BreqiToXwVgaA2U4Eyhe70KfhqxycZZv4rp0Tdl
wyKJlMjSbYnlHcYuG2FQT39m1tNQBpH0ieKRPwVFTf1C4Z5XY5jUaakBE0Vtt+KG9BJ9Gy0C7WA/
Y9KW04oIWFFTMrT1YR15HNVfAmTRFztdZghnjurAC0HTB91B7JEpUDxif+/iaOxYbIY4KWm/Kksa
TpfFTPh3NVrAf4PNLLDf/Xmh35yODclqnTGAuoF+UQKwNclx5JGUgKU7Gbn7o0Fz7veu3G8jAtwy
06dZCSNyU4ZlvKZPuPGTH+Z9Drh9NJh9DoinaoZLxIagR7p5FP0ttVfEXtr8ZLnbt9jMSevE/Nly
cob0eDavhG58DBq1czJw+pu0Vb0tdRiE1eM574Y/OB+HuJm4GNvnDgJe3np7yUMFuMWlM3B9MQFt
GVh2ZhMLA7p+wvcoIH63Z0Sf7dTGYsbcLryCdu7vpPCClqJXq+zeoep/TqhYw6d3czOnLn9JahHg
PzEo2sRbKUF3DUGhA6ULWcslY+74bLDmfAFpzQy9Kqox3uN3cj65+uXTBQf6GUkl1zcQ8VBK3m2H
s4GHsYj3AqF+UJqjnF9SN7P9D09k9+reV+Y/oa0Z2q5VpSC/eSw76zq8W9ozY9+TLrGH3Eb0vwor
keUr/OKXM+7WCZUSdNYCmf6YkFWKLRAUFF2z4BxbL4XeFguEP8PQ+EhfuUaCyiEglTNXWbM5XCIJ
RnmAVm9h/Pch6joUA4gsd6KEgfsjrnMfib5LFUUDuTuUnSsgr8MFHe5dknFf8Ga9jx1OaTivAGEj
2KkhNtuznHCQN3cVAxoe38w6OTuXpRSxQfp67HEUQeC7Kik6xPDYZof6FSwHm4FThzCPYnEm7Gfh
1DHJL3GM1gOo+tgJLII9xNZZqy+0LxpFFYN5MsYbsc4LwuPbp1X++D7xC3PlVz2XZi8yNC3l/pqa
jfpYEGFdn/AwVTKahVrQmi9/EpySOD8htmz7pR0ApqitwmCI7/zrd5Ma5ivzGSuQZwX0Hk22JVRY
yU3Seswibo23flyYSg9B4gsfJr2Z7n/foUJ/ShfuaQcqnMU/3tgpir72JVc93XTVQCtdZ2hKnLmz
r0kzkAvyoaxXvk6TCn51X6nz/t0l5xbagSfynizlSKXlTAwSKeUZmll0bKCgRACsALq0MfxMeg2V
hGA5X1CLf6c4yCJqDEIKs4U3GnC45sybcftXGOYzC5X//kQhGP3jPkPdAdDJVy7O1kqt4F2LZl7B
XrckZBVnGcXftt3BSBN2HN6UjTMWUbzmSKCxSzTbkiECt4zIhnXoSpEHuKImCArLrSVk7ZaJY0eN
KkxgG4Baalx8bVQ8PdJ+cgs21qCz/gVq2qfR8H17GyVOTSGFMjywmuWC/61I8p0FNLMjN//qJ88f
ybj/PoAQBBXDJQazBEgoLC3/BsE0RT26+YmVqq8dFAYdM+i/DYE8DCAOEKsvRE83vJw9Jb6zfaDQ
trpKHfSrAxrIDfWFSJl4Nlx9Riw9dIX1p/pWTNs5rkua4cilO8DYsk4Wt7DyHkX5PrPVgsn38u7R
JCI//YI1LXwbs/o4BGeweTLGnvVwV9hwSyhXZtFcD3+KgmHjvLs4K71+jdy89vyNczVbyN6P37G0
/3jmxvEI1QCwZ2+HqS4BBn8j3Vyj+S89lpEb+f6k5RDj/3jHa8xjc/FR8qj+Zi5ws8MjKtcQ5T4C
u4KSNqxfhb1drSWbuSp5PPSKNlgBUKf2e2zNJjG2zTVlJ3/5SjEo4jqDu6BXvEGPPq/EAlofOCcU
dqCJusbMQNlMsCnvrijXBBz1EzK5bGYlpKP8+Ti08jRdoRCNs+DuSb3vmY0K8ptVXST7uLyPVjGG
Ta20YM0XA8cUKis7atCGAhq6stbFA6YkmbQzgGj2F6v4xPBo6dfZu/iACk8SKk/A8S3uRFjFUHkB
Ve9YlOlVY4sEn+zColx1QmD9xwGiDKgt1E/vRSMXgKiXAxvdEdN45cbyxMXrPehY0n71tJJvUS0V
4R4FWLmlutXObFGMUuMDmkQL7WZa9D5bLthkbWZgPgrt6KQdp3ziRATfwzzdNy620P18HEDxf/cw
/cPa9djMMAISB6mn0ppM86o63oJCdGcmP3wSADkHzB3AppPbPmk4zqvJLk2ZZl4+mvfET9dwwxye
ad/s9DuSvdyxp74Nuk4BKUy5JMgCC4hqmXgfStOdSo0QimXic/mGUqdaZUcj3O36S55NXwjXyjBP
d7TVbRnoXjw5LGoYGRx6HyO8UDkInpvAgdd6cClXUktPrXWNd6gAQHk2oTeH6oxb/9F4Spb8fIYf
HSWsrvDeM1fVFnKYYns4vig0u5XV7pBoq4iY160QJZPV7FbdkiDDCjbc3Bj4Yljsks/wtqOZx3m8
lXwv0w/e0aMzt1paQtRbwcSTpgk54ymxmhtDkGy5xmM+bo4CINoaQZBePdPpJVUbCADBGzDAMC2S
dBPd6ZNecxFQEugsB31LDAwnKQrnaTELMT6sJneCTbcrejR4IzeE4vxLx7IFVt+9GgVZC9pm6fbZ
F9rSYu6WfMIfeKJHq9mJsp2nfka7PVDPs4U85MB28VpPDkZQds3KlEi7qDYQg/EVlL5IW7tPl8vA
ieW8e4mzKuOLu7nvI3QOdJy9+PtoZ5ymgPg0EeyHYh0pluSpkNk+Jvagx+O+PndWvA9Z662HBNLw
+IE9/qnPvZRpC747jiH7x1uZDP/A2/nq3UlRrxqpbIZ7f46OaQMbYq3mUo4CmgNxi3teG4nSjvS8
iLe7vdG2w8MFBgMp9aRz/lZY2XJ9FsbXthibcjMKlPatwQzNdxLXV957TWM70TiFn1dpCTGOXzjy
noUnO+aZWZPrUnj+mLADFxk2/kpqSTpI8hhnjQFzAo3B6fopG4ZvVkvjFnK7OU4G51frcACysfH8
hJrjqC23yHnBo+V6LRVJzGVl/iq09C/jSgvGx1YyHAW8h7xVin4EcPx+s3ETTmm6upY5zomteHY2
GZhS+vzqugDS8YSTy10ktF6DiBYG5+y6FXL1wi9lKkza0IZgpexKFGbYVX3Fl9BsMY2bANDRWSyq
FPZ5CbKW4QlVrdDUUpShzm6KHc+7TIabFHNH8dy0FYLm837W8ngSVZWFaoIjR//HJdLrhGCv8znN
5EYLHhZuXmTmP6u0lSdUA5X9bLX6P7g51vzJ3kfBJypA9myz4vEK6crw+bwdfDPkqv7Sw1C5Ifyf
+S2ULfq3OFXYzcSzA2NEH86k3pMK5Zhwx/fr2TmJxoopfGfP0rhDHAXewFa38yqNn/wl1DPaNYlu
QRLw6U6zm95ehaTFP60uQ5BPpVYDB5di9Xz2Uz43MA0uIHcfFB2a4qMse8pytndBnwLy4OvLp9dd
eIOp1HG8aoQWugL5dfXQic7FJd1lk8xzcAulY9GMvgyx6IYXZTq5c5jxsEdYgtFBRcYbx2ilkfpg
qaKOl/CXH4KnHVzzLRSTO6TZnzjnoQzFB88FEtf8kpSGQ5GPKdB0JiJqjQvcwXo9ZqMTBGxiM3aW
9upjN22ZKnswrMAuRihF8dCg75B6uZP87lEUJ7hogPPO8e8BHttIp7WRX+s3J9sC1xJ0phpEDYFT
fPx+nunSxOEFxNcxxBO6OmcyI+IwWNYgXxv1Xv7MsMRA1oGfb2VC0TQwylP4kpm+bsoxR6kYN26f
nGppu0cY5UjiK/iJUBsbbWKnCSgQQW5P8D1piS8d05l5vPYPRQHtpAcOoN0Ql1PsKfctwWUcF3ww
pVsy3+nwGv1uQfh0++WpQ7uJsNQk5z1TZBqbMp1uDAKR4fUSTMEr6Vlch/dPZULKSKjXCWv1IeKW
38MfiLOJ/IL+ZrQvS4y49spAL+RFHnjHU9DxJlXgAbPHfYzs0sE92VzikM9s3L1qde1eCBZ7L95B
alSQ6R5T66unvKmXhX+VnRD3nk2xZyLxoh7n7t0b0VsVTGv1bIaqCdf+VwI3aHq2FYLn+H1DbsjV
SRKKWk9U2TiLVmlUrfeYYpMLvz5+eh+t3EsWtz3UiD9TOvbyDD17ij6S778pmBsRWXgnklq9iSLF
6LlhFJnVE/2NOMXAX3bQldnNV5Lij0RxVKIZgfJzaBcAbEADnn28YVFiRQyJM7s7t20NLdeWZfH9
JAmzvrkxXLtQ/WznnpjB/8ODl4GVaELw00FiM2mtj++pLeBPd/d4YHJKNzps1+ZkeBeexo+xW1mR
AagY95HWIHrr+Zr56gYU/4Flnkn9swLvg65DlySS5aAAskziVyz+2Hf63FRowpC52KqF+U6o9yLn
ZjMtG5GpRxgjnHVd+53/vXjrDGnD/p3apRkkrvCMT9AM66dUPzrg/eVSpHiOF8SJ4Ol3j5f7Po9n
f3JTPV8IevAqmEdIkXC2h6LsXahQK/4Xct/piZBh+Tci4tLgePWzApNjyFhdA+WmpRKbTqwJ6MuK
62FyTeRwOnVMd1Ljs7AL1jRSoEdrJIQUqTy7EQT7C0gsF4MzbiZ/K0XrEAQ57h3hkiEyIdDpbWzF
qXB0ut/zFM04fQEbUcPRiKDvd+fXErb78WoyNt1/xnbjfECOa+iptGpMXMo/B42+uzWgcegc90a/
423R4hReD3HjCjmKluHF2OX8kLxVpNIwSYp8FdujZJEiIzAAf9VHlHIOQIqzSX2IRcQEA6y64G/9
1nEx8ApRzqKmXrU/sjfbTRAiFyJUqR8g11FzkKRcZGHWWV/XIELUqqTk/QvcPCMFGoS/b3D55IAz
v/Uh05oY2KEHXPxhu8b4aPNnIVrQ6pjDJ+IqluwIRrxQbpChXUda7YHbnD6Hw1PSOsTT6W4qa7oZ
gbSHqbpqECwQWEKPDZIHtXL4pPxoSrV454ySNmLJ1QFlAMc280FKwNpbrwqa8ebXcWlsuSQ0hPjG
oXW8sP7mxoBjPWhvy8pPPPT33W8Cirrio9nXV40ddEO0EaRKhcLPr9MEVUXc4p13q2Rc//UjTlv3
+RLApD04fWHDwZ58HhjwhtpH0cwI6dS5to53vubd2DqPonB+4urD39mC+oJFD+H626VsCiVdEkZO
Qxy/puTqJDTRTRnclMTKJSC/4vQ1nZeSYUfu5j6Trb3OImXTZZkBApVnEqDxikmCOb5VTQJpjOCg
KQDE6Rp7u692DxUC+2fMTTF/F95wqk4AVo8Ea2FjnFGpoL80zS73Pgd1w3aCuvRVv9XR9lVzplqa
Kz+AFGf2rHSkkaQODifreiwoMybm1zKqVm/1J0XLgGBYDo4I9/tcF5Pmo3veMGbxNM5IF2Mnjk+4
1nhOVN6JQeuqowIs0fLt/hpGs9C/+1GWDiULOZGuxp+b23T3igHJhhwOW9eQNcRCZgbYWQxrxjcn
pssVj+ACxWdT9em+eCpx0uc/aefWJPQYACmabiHnYWdPvpNxWvvd30duEPBjyE95xr6CLjpehjhm
JAJXvMTcGPzPObCEn1MoHDYPquWcFkW30LMMJXpl+sl+hfoVzT5uOUBg4QLNcAdgOgOFhMUaW56g
pl544ZGE18o3AMCKDS7I4Di8aDhpwtnOEplFcsqgsW+4UIDQR2xSSodcTIuUvDB7dC1VYkCq+Qi4
0MPJGF3+BWAt6X6KCV5EwLQ6x6+6LX+IPRxi0gp23cU16+T92cbhBGkzPasCVCrKrsifSxvO03NP
7KKMa+vV37Ka38yRl1E4tlmMQUgxEa7FBROqFpFknhGOx9kZyMlIjfW32cEX44AzWt3m1H7lcxyN
on9CezASuxHt0VVPhsdL2BYimOR5yVqfZ2EuT7p3XkiM4NRrWKHYLfvKyRlj78x3OhSvRxqSp2tE
iF2UCNWnDuWt5aN9kxU8VE6bIXVL0VnuEcli63J7lJxlKQEmqgXhOx5A8fkw6aAwUYRuXOGdmBd2
nzb1W/7dWkt+3ruDHwem3reV+VvaE6uUBqIK2Yagj9LnNivUe1YiEgvIhixGFRi2oTugprZeBhUb
CUutn7rDt4xGb6XmvrnR/7kKbBG26iTgRpRa6EiPOMtCtVog/bEdK8EjGZSz/FrRw6uRejC2lKzt
W2FalLEINtDDrBuqL37rFtI+E3wBYXzL2tA3K8xgPN5EVHKWuIvv5VoX18YV3PhNO1qFOMG5UIpp
pWpykp0a3hp+CRxxAfuWwADbi3Y5LnVAjuhRdJ0NVOzwF0aCmGDDANrZYrJWoN/tJt3citUT6D9w
qYca0LyVNpyb3XAIMVG0p1FjdoEiarc90OmLKqQVqiOt1YFk64/Ks5qD5y6vzpKv8JxcdiY9YPPW
ff3YDEhgck6JrNrKeySwAfZDJkvibDdnDnT5RkwqhjdFRt9ydboxrcG0WdWc8Pg11XvErqc7avBN
e8sWnf3cj5lwRxWSm7bvW5llrEngiXZl/IB7ARei1eIbxN0yT7b33epMgKE1o7i4Nc8dpCbgc/12
QeQUyQ6ejxicsXExd9DBYOr6YwAy262BNIP/du3ByammDxCnvOQUON8GT16Bc1wq6jntRNNjabDh
thBISyv5pv7oeeIuS+lrHsykzplNr80S8L30/yv+bj3tb19sCLaN9O6PulTM8zdFKfq5XrLIs5Ja
rcMBu0XtaGldz07X9Qv/ZDg2z6EUH5XILjmKweZVqgZS8k48uZ28BdGm/r+strvX6TQXnX9oBAYG
Aq2ZqLmmU498WP29nYEjn4IzSIUFILvzuTMx7d54/A1A/paWMfabr82Uu5ZF4HwCloXHvFosYeL3
hMtKpsIQQV8RlhO+jLYAbxuIUVwnaYKhlKOGoHeWA5+0UVlIyLxyMT1cfOgf+aywKBdDo4ADMeh5
FArMmaYqec+KEl61jto39Wuqq/bSBYGD6FE+eSBEXMmYiLbI3xnaZ8vQ9oiXCT/7Z9AdtNW5uVeS
rVso+rqS8ftT/4gsAXSjtdXCycre3DcBa1vMc/Y4YtX61PYaAhh4JysadZqYoNZlBu+9GOVE5EPp
vhszpG+TtDHHpr8XSoMKfN4tJjqi9ekqmAhgnBBzQQsitIIYgbwGqli1njCEy978t8d23BurFahD
O0nBfQ7sMlU431xhawVlrBH8KsVHrF1VHT5aYaPRG+wEIvgN10LxgYtiqqTu58bpUyN7Nw1tkfsJ
a5MBGfLd8qcg1H1LXsO5fQzElgf38f7Ya4OaGQlEURrCNC74RzuidjyMKyveZDB2SGrjeerwBIWK
N0pdNRYYAGQsUXNQG+mYu4k4HHEyusnViQiuDJ4RLv9rvB1/10Xg0e2gZ08n5n5GhqhQjpwTnl69
dLXBb61lOFfVxJz+dS4j/jZhaaIEwecXO/AQcXbj9pQ9WkkF0ElPAe/1XRaSr4Pm0LSn59kZM9Al
rZAw6gwoF8Y+52mbP+gpKy6OVaT1XLE39BMjdal4T0bNY2JJ5+pzZFbMP/JEZBUWdqxiWHA+VKat
b2aivd8aGC2hh0iu4X1pTJYsYYbnu4kjvr4JQiyxbflJJcHD5psSqaQT0XCaTLXauqQzs7aHEWQI
Ta2M2oXohdn8tJF6rUrmRvv7YjHP/bH/y21p+zDmCS2Qx6KKjK2q96dUIMtF3jNpAJYXvdSc2ggc
ULM+9JNpPMJTp1s3RksT+vFucY5r36AVDIOYvTDXpO7R5vZlGTrV8WQoHh4OjQKtXbWDvLg2eyLX
xBejlP8GmDHGiBG46QEr6FzK1NQx81n8fyQ81w5IOFAhV41bUCT+sMa4XM5fsQepH84n9aKhowLP
OYfmuZKKn3jNCJpRCZHL0FEMHCYT4v110UPDbc0+A+h/6BlC/cmXwc6vFLOlypLBJUuJngARqvJm
OYvKsPpuZ6wauBfnE/rKwbo12PA+mW01mu6I9DNKjXaEnmfJ4mIQ9HNOdAIv1D6Pd1/qcRXEvpFt
hHrIYbQa5r+ub7lRp0InRr71qlWisLPHiEHhNoPEPjKHPBZb7GQOpXpTu8C2JB+/FkVXnj1CuK61
6z8px3JXblh8t7D+VPbIj4A1+MslHlw3jmcx8mVN5hmhYC1WFPwLmDLCeKCuweOKfRCIWBoEcD8a
/F7lNWF9C5SopYn7VbSP4h4V5SBk8T4AFhcA+vuqN7cvcSL7H50bvccmoh9xF77x+A3zeuWkzbNd
AjOrxuCosGsiUCoWxKTl2eU+ONauDHZpautxecxcArgkBbQEjtUcCfyJKo4cARqznBmv2Kcpm/cn
RYkF0to+RF8k2+YawsCVYaiNvAI8qJVUU6Nec3XbdH7Off0F66jAEAKf+qDWN4SBHU/m9F50/36K
Vb/GqlrKHFhgDmuRmn8SxxtawUU04VNMi2VpUq5WKWmmp730q40HBjQ6Pk3ob0GAiK0wotlNg318
O5Psioqqwfd3lI+P5Pql0+DbY+u1WUcVCcx9eqh+27sERaJy4q9hQ2Ff3yXfMMg5rhai4bhWBSGo
2uGZFg/IiOA0rZXvIgzgC2szcuKvw4TIIznk5Ald3NtZ2iALD6jOz73Q5wyM4EujOexqtfIZ1K68
V80Lfx6B2BVnFEID/J8ls1+oRpIkP0d6e1IZngYM4YzL21imBKFLsJ8eY+5FwEja0L/awAVOnYLK
lhYmOL0vcjjH/W9qClLtDBw33KH+8b0/lsajeFOxRR2ub0S1D+WxRJkpC8iHmSeEyfPmySsTxLNr
Mswoovv44qf+eA7Fl5O+NEuznApubUuCZVBLWH1Taf/66gQXMV592ndCaXN4TA+RauGsM0NRf3xt
8ml7CXzRh2mLZMvDbd2EPOmaMNQVTmUCH83OiVgjVbioceoWhJEK6VsWpMEpok8gAcmsiA1CZuMj
ujw6POptZvpt0QXCzZWFhhU6t9K4XRjogI4cIs+EwdmBVjl/YV+oAAf/YHNKLls9tkhChR3MiqVh
ou3mHq5WHnErUhq9vYhNK7dUig0IPqJQ7upepcIK8Mpi03XsWeTIo2Hfau6YXWlDeZYxHE8x6ijz
qaXBjZqBqRlg9nlIKi0uCoGOccDrV/U/iUsQcdN4UrREUiAK7MsHuh8dwNBzt5VzsuiKmH+6st1q
ZqNExtqPL+DYEAdV77yzAi8oXn6PO4xbW+SFTeCB6VMdVKcuhFZ4MUBVPyJMmAILEqcrdeYSbkmt
1SfXDEhytKYiIMNQ80P4cwp20twgd+hurhNxKiy9Bio39Eo6VB6VwAgHOMB7f8yzNkvjjlnT3Ry8
zTpJ1NlLL4wL8H00OYzIVUhaR7WZZLpPMwWasGGTuSyvVv3lg2QssI9L76Cz79P3cW1HWBlvQrAH
FEaasvHEHp7PXRIrogcIZsKJB6BUBmUSPShlHGB9kp6SOBC3LUqFHzqAuBENkAm1LFQwB2VuvA95
/IX8V8tl9TDssXEL35db2QmiPobed/o2cF4ipJl1pb1ML8dqmbFSG2BXb0NudZW264RgEn87bNCn
gGFJB5ahOZXF++bMpirZeYJpZHCT39ZC1LU1Arr8Z57BazHrPtCq2srKJJSwzJ+FeYCw0T8NVq2u
e5y5I0c0H1fHyMvn4MbXSZJt2FmNUW27k8+vzPXB3DY1KQm2v9/CTBHelaZgIWHWra5ZQ3SLqmGO
9gMSnHnx7iiDP/BtXvfIGzSzwgcdTJDZsoPIibrOP68gGWcZpyH52WvRFRyvoWCvt8NLyj0Um2d5
0233qi2S87zZT3H27ySt0dD6j28tV3YjoutlGPxHph619+7zls/ykcR+RdvcHCvSz0JYmM3wJHLC
Vt6gp07kvywq4mpTEUXjytpCH5MTRgsRtzER3b0Sh/4K+EWyj+n/PTC/K3rIbE5uouv/GqIS1wuc
cv5/3WZpinGm9oHEDDFYVpbJ8px6EG6FhMTru+xl3d/6567ijSwX+BUeFpJBdJAqwe5SBGytwPRf
/Hk9WynhmzUV34HTyZnfwLOxT+VyDyUecghASScQv2GrvcsXGqWdjvS6z0ef93VL+AFLwiubn31I
T3qe//v7Wxt1YiMBvHLzLsaWpEDf7bRyhQf5IarBu03u4wQ4PLo0R/0C7jQ90Fpq7YWKQbSEDecn
vANyu3oBIoGqLB2W/QNsknEBusHxpJ/ozMJ6xbmCRWp1lxulRR9fRIEFSn9PlNAHNE/enMoaezqo
u5G8qczRiFDP0t9VkLV3Y1nizIoZbnQ7Z2DppxFzYd5uhukxU8ChEmqLgfRF8t9kOoCbc1GU5dCf
t4t+6uOHxrxxciqCRU5sjslfPria+7SldH9rJ5Cf57vDFGIeWw7Tw1lHmhxnPKR7TcnkdxSiSuvM
pQorr0DJ527BFpVOn5PSEsExS7tAI0STle23/Jj5xIu/P89/n6ZWMDVBjFY1GklUjA2LCIDXskKA
nCNGpTf/cvfxeUv7v/Vi5TRbl+8t5fhwulo+ChKiykNr4p9aXhThcbOKYoWA60V7o7dmn2uGRANa
8OrtdtVrxGm3Re+Tbymv9w883A7Qrubqoei/ALXfDICaoHBWMdm21QTD0Rh8EOCUIkZGhzR8uvdE
NNWfnlLkUoLHGCnhrCDUKY6nn4r2hJHJjjK7Yf9EnxrsoLuoWP7BSDHGqeB6N05wenot2D3G/7aN
DpPy7jkcIuf5gldzDRUcBNH0wJG9dn4w5x5s9x9NiSO8SyDI5PW8HJLe7SuztVB04JIaT0WSL/BT
Pt3o6j5h+o9yTsArm0Xj6UrtlIPVFPQrU743Stw7Mz8VjwFIk1+m9+pkj9k7nFbsS1RqD0MEpehk
Nty9S+ck6GqBEk/CQKRWoaGVMa2j49EyUMWd/VNN1bffZvsMY6mFXCHnPQaKa9OILdVWjOpQ6Xgv
9tn+O0Qg7yQxtVeGruH55Ul15a59GbstrBMUX/ET7qxSZa8sz2iumaJZDLR9VAZNJAJFbx2vHu2l
XCCFgeCq6SOUUIIs8qiWAwNEAi/EK5HDzt9sQ6T9cME5dD4Q50b8YFTwPomgCwaNr92DpcJ0zX1b
fZ25WaCW7Tyu18j7vYT+u8GRem9Y+SSzZ7bqH+pwDpIuAOV3j76v4icAwLF1whGEcEJx6j98lMTm
f+mOhyJoVw+2hOFAy2m3Sca3ygnobIYLUqExyj2jB/LYTKHTTGJNFxWl6yeBHLhgKIpF4kmE6LAZ
PlQ2m4MXE9VbtfpQAkkEFpR5rJVZ0wqMkcgLkacXL/eTmE04TEpLMzqcRLEwSB3Tb2VF3yqOmdVi
JeXUDgndhcmdzgrsoBWo6u6dsyYBM2j7T1VW4x2pcHtP6DC9jnvhokdiH+BEM0xufy05rt8T7WNV
tkPWo0QBg+DktYOb9jYUiKgIAo3SaPz2hYw7Knp9896hqL8bFliJKmranjF7isGCadujhPL3pr9C
VpBhPUQtJKxjf6PKaw0y7ckL2PLMSmrga9gamqB96cy9Si4E39o9dMkxLU4163AabstSt1JdWOdQ
IX/cNGxaMIHU5bEVuOk1+E4Wc2AG4uYug865t1BheDHs3LLWOo1040aaaT7uCAS7fglT+616qAjB
pWU9Qd3Qy2vrS8ZWePx58tEj1VFhzd9HR27NEY7SDWyItCh//5seiwb6MC9nu6KLy52wkz1RBL82
WVmR4jP7eoKlzyqtNYPxURZ2zDbbpV4ycsiU44bnMqwtkJrlFFllZ5T6jhvgtyZntn/1bjQZIBYn
rW+NWwkKDFLhUdukIOX8O8W5pGhP1SuWidROhTz2OzF/PFWS+IgFQSe9zgkkHEgDeSxHVfCbDJGI
yGUJyiwz+61zmPQojoTsY++4/t97HkxbygLEvdPpAwJJZDrzLpxpPXIats+7E4BIOPphxR84Sg7R
9LMrQoo6TE10IyP+Uv93sH6WvnMN7weZWzXjWX2EbKF+HusVw6CrXC9jmII6zSOSq0skD5yVm1Lg
RyNj2ebGXfa0Li0F5IZcUiGUKtstH2aXiP0SgxRcLjmxtzU7vk/+wfcd1nacYOEsyaJCP8DnonLk
m6vdqzg9CWQdJqHSHK5N1Zke3KkNOGLPMlK8y2MnY9dqYc5oR0oO3ScOAkggdDP0wi4ivWNuoBYe
ceRYNstZ9TgVxBQ9uY6v0QXT8gHdbztxtqNMTDVY1FQRNpIdMiICaMctHrK09oXwJ5/VkfAujhWn
eVXPqjZ1HG9K5Vwewk+yqApwRO7INF2oRpibIHm/fuJ3phQ7a/OKKLCzrayWHOYKUsnyEP5fLwr7
7a24EB0JDqjHvuZ9GVCc4Zsd/BiNvT1/yKiszOhMsQQdB0OfmaODQWPsdzPRj5mJWFzCZQrR2e3U
RrQRvIWBr4VKSLT+jDi4ocZVivwAx/r9pFSVldJhGs7taZBuTIRbPZIMWmfu/s2deswL98JqGBWC
tOwp9N2YVrjzH2eqxJ+92z3+3YgBchkewmpRO+K0axjNHboHO/bjOjgEq7mu3Trp01ITjaKjjNZS
hAOxL/hPLmyPbHVoUOpBZ2DZ973YnTHKYA4dWgVwt9TdSBU7/HGyaPKQYCgiZc6T0zvd9WBZMfWT
eG5MhtqTORWlwjCfnPZwP7IrhHYZMR8OF3F05Zk8oYBjTbDZViwcFUgifFnMb+fI+ZM95WlRyrXg
KDiBFUPVeawjKQ1GLsKR2byzm0cqVl1fyVdKe1qnJTvrh0Orc2W63Q90Vfw7P5A6vtVRQOUE1ywM
nDma0WBjOHdCPfRu0OErfloWNUd95iUEfElMRZvR8k1W7Tbo38cyJMMIEtxcfDD/lY5E/1Uld/PV
cUMNENt/iwJ3UQhKVaUtvmQCiMJy5bIJoKhB7rwO6qYKTPixt+Pxoy/iF+2TLYp36ik9zTQmsskj
qvAUO+FLG1NsdusXSrqUDzT8RCgpwnP035MAkrQYp3W5EZLFV3T4fv3VAnY3KUgSsM8+ahaMXiB5
FM844DqsDR1TwCwkcJPbf4JWR5ewM1fDNZRdD01n/DQ77w3SlRdarglUV3ublJAhGRmKj5fEP43k
4zVdsx1bhWrKavXNSRaPD0XONc9Yqq6saBh5nyOssh0e0BDCCK3/Eba+qLEt+Nh2vlZ116ltmVWf
Nx1hEZkM7GeowRrcpc5b18svobocpI4uGwMPF1ehKmF/sJxqZfLaZPT45kfA+2rJjIuq9Ye6do61
YXGtMsYC+w5u3wh/BWLrdcCG7auWR/GEGVhfGF4Wx1eszsu6DqcjdyJYHyeqOYrZ7gJ1sx4kvQVq
LjMn0SFF/VvNilHvYjzetk3fGV9isYOsdaBb1Gnn6qkYFFQarNjp/ycVYZTRre8o5Z9LqPuf4mQF
aYp3kccFpAG0iIaGF/+5MRBsZATGLk8yR+US1ORcR+AQV64CO39qwMAgswr9cspzu/OntbNqlLtI
UwZGulnu9QtHPGJKnJcNdzFVcD2m1dOBzjx6JCp7YOe/00ruPYr6fgdklfBAnegsAyWvy5a9Ewk+
A1H26LorZ+IwDmGkh83h6dbJPYQh2t/upk+GOrXo0LeLiB/DooINLQ9XiOq+DWFqT8pGbpelCDoh
s6x6oq/hhnGdGf1whGrdbUHpHAHJ7WJCLCNKc2NlzqrX7uXOgMpKT87Klf+ZkZ+Hu4FVPTSbb4rw
wnPy9YhpH+C/Mjy7AabwXVxd7cdO1X8iA1k2AqdUH+9+tkG4VDwMaaETE/wsWVK/BLvQxIyC5qVi
BQoYdzUPVAqzbYl6AJGXjRTh9uYmaYIwVgHewIq90FnoKqJ8LbO4bybbyIeAzNLzNj42x7jZbcmA
2TcrgQMMwd+eXFzw11QBrEsRCu4KRu/aM3UIGbjfitaWqSX1vPGrIbsY66yE3iKusJqUEN/vGnRV
Xy9VQlYAXiDCZOlxF7kFT1wx8VNXr+3yhoypAsYDOQC8A865+EIt/IX6p0RI91nwp/GLS4+mBCBO
HNd1eeIFvwtGqu95RK10mJF8Mz55IRMsbKgMZYQOlvwABaRcje1EXyydAPEKQh3BmAj5/UNOKFjx
kvWyetiQU/A7WIWxQQSgZG/XQQ2cfdmHzqqBcEUqC58oNEqCMVX1pzJoUJkN6posYQWrOOBL1Au3
sol1OggFmkQj9ucQ3yVrbJifkC6FfWluxQhII5mmUReLoswVhkVKDxMt/j57XBXC1+HmbHmBQ6yQ
vU7Cwuvli1qUYO/TYLm4CPMtsynHI0LAqwEJ7SLxlAo6+Jla56Ki9IvmRWoN11gJAx3gHaxGLu2U
DCcyQ6in128kg3uLv60ucXqDzs224z/rTSxBAVwv5X3YXWEK2qZzGS2FRT2SLMLY0/8SJJMx9BlT
RSeenDV1GsqBH5Da2mM9VLyiu/svnTncOnzet420bMYX7+fzwtxNdnHqfB/3Pg6GbrdIBm5RvxvM
W140CuzpFWvow8DWVHOEAnTXoob7+ZPujnojOdpJJf1ZuxR9j8M01i43TrOZ+LJWKWwDi396jwhP
n4wIfbcJuv95oMlcC6XLOEuYOQ61lDtk+Wy9a4oMDxE52j0csgyUJ0qjuxPdyy8FDUlMzYZCZ3Pb
jdUC9z2FtH9sRVTMm6AfX/CAK3NZzaHyJE8Y3v1+DrGV1kNFQasXoQOlhxi3BpfVWqZIhyFpjzTV
TrSDa07IwHDtFHa0m1vl9Y2auLAD+788dS7pZbQsc63UY1FLIpN5H86ZeM4i7t+N4P4gDXd0UURa
Ud2OrmrGfJBg0k4H+xisXqzRmD+arQUCl52X8oQlB/+izVhFhgqkxpKpJVH5cKb2Uq/wMWgcuMqi
Vfyhhz3y/Rtribx3w0/Nc3effZ89HRqTEu9WgFAkonl6DZexZiR8r8i3uX3OLj2t1GqV9XcUZO1j
0Utb0VH9u+SvMk4BdU9cM8NL/S2lshCp3b+Y1xLWF2xC5DttYwtBtcEnbt88YahQD4u9xTTCC5iN
/b/ELM7DFLBbC16wnjZEoPKhPhQKsFwuHM3ZBQ6/1E9MYaKfbTolzgq8tsdPc6LX+he9qh5thJ74
cC7JUblSZIZ4ICu68OxqAhlXLU6OhHDnQX4sk0610q2rmfoB3NzXhMDSteKj7LiSWkPAQpcPssmk
G9NNaLFzp9M3aw2MLxV/8xQw4LSd+tvYd5IDqNt1sKxTJNqtQejxAt9aaMqMFAwJT0YVQYLOu1sD
qmQglXYhyAyK7marcz3RRi38iV2BO7ANZ0dcZlZ0XbhQKMj1spH4HRzVbVwDMx1tPVIn805mLaJd
ij41XJDipZFLqTao/DI/xU3FZrbF+Uxb99Bkkca5ToioNT506B5VFPVoUTdu03b9BM8yhYDeX51h
2T+/gg2z5ATppbbM4nDAnPejZ24o2ReehLh2JMYxAgqNxJuCD1Aq/6Y7M4NgXvG8TGpvXdv/hD5L
74mgulBCkxh+8gJlG4L9aXzeVpwr0RxAyCv4qv8jTW6bq90ZrTYxy+WmlP3cVLRnKcMbWh+lyIMe
DBfyyUP/RbbT6XmXX0V+LSBhkPf7AX+D7cMwO54fybl8QYBvyHSn+ZPnKN2Oyfz/+sVniCVLqUx2
CJI91Ye81uGl0pflqlJ2iR1ssTyR1pGE8RtHIP0jYvAqYuCd6avKhgof2FVHg3ba/DfyAM+nMQVs
qLAV7Hcg9lPVE4mCMLVAjTNH6vUX7AmMsUtqeTz0dx3xW2NKS3vVVuJOR9fewZPwrP6yWBtUJS24
Fnfe7Ey3uLae9sdHW7mMLx8+wNNzxolLTBKth2+B+FlsaVReQIfynlnhlKet6hFcP64c7DdWzMdG
l+tN7zpw4B+Ot8tjyM1CKDbwp4j+TU2sV146xjQgY8RoU8+2vBayso30K5Kc0Y+zd6GvEfgIM+mR
WzlmvkYy0RlckV7xJmztUA5QcHHLrK+X0xPgHnU27pEyF6jaEP57RarnB/CZaMgYWE9Z/Rv8pA+U
lcBUUl106gP1OJ5Gb7MDA1QLuLsz6ke4JeWI8oJVepwkqq4XGuC01W53cI/6LVn+MEqxIMYVFArs
FvyVgtvLA9DjapfnfJloj7vXhX+muXF2MJ0amvQVI4nQfZTgmSaiZVs3xqN/fctb2jHcs5ZY91p5
tUUE7zsyoksOimu8a/gzVzY/DD78zYOXh24ZNQTKVfai0NMJuiwa74LvogtiBfUYeS3+BtFTiN+e
SjtyHcoC27CDR5Q1trXi1Nga5nZoE0I7RpkHUqiYuD/6Z0RinM7avsOENs7RPa5YLqZYntTQk3X5
xAR8aPU4lRQaII4OSX3d+tllzOPUGzc0BRZaZBZAViAD2kZQB0cUTj7sfpHBD3fDlMezkGzX8YqE
HQBKPMWUDUnMQwdz9tau3L7cwGV39XVVFeDad3DsI1d+01l2b5GCXaJDQ2jXiT1f5QKzSNpmnZOC
LFvcGRve4uPGrtSzrQfktMw+/8bJfVAkoeHRt+X5vwrNMc2Dy2K35LAfiYtpxSdJuwr5dGFBUmR4
cpZkwoKPxFSdBYl4MOfGLjrDFvFnUPhosXNULe3PfhwhK7H9bymx39Zz3PTbM6jD03WzZ4idW1uU
XlXNXTyw8lTsiy3Nj2fWLTO07zMNxfJgRb+cl7zHyKGYrHlhy+JCd3YqIb24McTi/GIl0VwWr3qf
U3KjKg43xjJJsruIGnLwG8yz740Cxrt8PbC4YrQ+jRv4+Gu1eDsQoRNgTq91lW5ZUHNVLQ0nf7JQ
6HMOkMt5HmOwxM28e+Y+5BacEv3+GoGpcRnxw2BjFr7evKmMC4+gADp5s0h1JjvrywTNCk3pHE53
gnw0opSmpr3I+mpDejw/CisWgwW1GbAHCyxHNE/Nq/YMWwGN6gLWqzwOmRxbyZNWoXQkHWrkXwc5
EvFXwZtggxfiMj5kUD/vTbhUSuWQRMe7+6aMs+E0QrrYXMnJ7ZvcfdN0BnFVezjpDjNlLPT6vckC
FRbUmpo17BilvWoGudLcUTVzcMuvnzmbpBK+CDCl9LOXMWmL9vIAXh/weBr1Pxrvwv6GgUpQkdv3
zdQ6LtG9ploEU7kem7fOzJbDt2vBcGIQfdgE74QusVp39eukf5fV+qiDy8TiOald5iepzVwqOs7+
fi+CUzyTx+bFTpv9qNYL/TtjPpsQLdYW4iGOD0IBPi7c9iRZUjbJ4EW5FTVuhBGkqo7kcXUDuJks
tIZZJ54uVb33XL34cdr8r7Nkt6bINtq8PXNxOoTKxtLUlGDIXURsHCjoDxHRBClH85I0ktHxNReO
k8v1YcZ2Q85GEePjp2dkvzCnsP4+ZOM5MfqY6m9+1ohrQsy4vGyXBGjzzXEWMi+ErVPWONsQlBvK
LOh7mh3GrglB1hcukDgWmqG897FVAELc08mNuiopN1hCyd/YHcN1vk133wAfUl6F1DkLbYb2T+tQ
brUzcbja2SWyJt1q9QyI+XkXs1LE4LbcZS8Q9JuKDKwe47zwRK0NGf2Qp/tTtSBYGf/0/+NDCgIM
Rpsy8za7bUPjaSwyLtwhHKH+KLEvrQDWuCZYmhXy6s/TQkrW0aagI2o+PFfUTrgh9kmT7YbJ3LuD
E28bSP7C4HNtJ+6mOWuzfa67j4xf3kYiZuWELAFZUGF0bDCSOZJrssFEN2OM0HeN7e/lcozpw1l0
14lKIycB1haR04/Abhx2LLWYLJNWQKoOfhtQxI1vyBHxRLX/J728Zo/rv7WEp4wNzRGCMV6Qh5K4
g97AAvp3ZqJZOSdzXc+lscJ0/zYphDrBKz8HAyTINUJljOom+Fj/gimlT+MtvFp+8sscpa9mE4NL
8g6JCaOAKecIARTgwy1A5qmQYOvK9Z3gMh9ckE7PlzTyPeGXZIU5XftHeVBM3azvOTNTj/uBMyOE
ZiUUvhYuuzBdC6gMajNxrcE2kmfFefjN3vawdEQ4D8B/Jl7tvLkooV7YYhRo4r0rWkef8mPifMvk
pwaWkAStGS4VeBeGUeMMcSXXQ/tNAf4YVkbX58cyXALfWPGZtAtW3APyqMLc7xMAy2QTcMYBv3+m
bykPS+jQJWbVDZiL3UDqOOYFUmigqFgWF5fNU13VTgaJMGFSAtAJTPEVhhZEhqgTph1iiIAlIe94
VPcJfP2sb4Rh6auyuEiYQpcEQ0aKT323c+wtm/MtGRfaSrsv0l0pQqr0R1qM2pz35naJ4sdiIzkH
mmi9Jtr57NJzJCcKYM3Fm0R8X4YZH+kaPbOdRo1VRsl69Tavmvj7RlAGed5hajzm029wPJeVYe78
IvxdWdmlgHRcFS46dLxnWhh0b6ak3kmDVKC0YXTNMq699wNiPRdBoQf5IIHc4rCF6aKpvWlDsSEE
NbksO+OdTu53hT/kVV99hqXkM6eQhJ4bJMuYC3LCXaVHKnzqVA59UKhnjJql3yfZYDGztfzCxF7S
b85BTIPt59gGO+lxgXJsUBNWWO/6uLtgfSD3Q/mJRvVA9s2MqOyatxeJbKTTAl8Nc43rWixU+4lN
5GjZ6KZlmXoPdxRfCWL9d5/s8eFjHDoRT0W8O7yJLlvqNoqNPa9eB4ePHp3CzD99XqkZ8ilDbAqc
O7NTcttnmwNAD4JLP4st9nf7ohV5AGetRG/bcK4/yl45TZQYdru7NGrqj/YRds0JsXdfmPXVnwjO
H0RmxoN5uVFj1+uiTsZRDzuX2YY/T0YE6fn8Kz+WF75B4C6qzbyz1y8qdF6i+c3OTgDKsY9lznzg
hmj4QrMWQWdyV2iVEyv7+83lrxZGATlqFkUMyVJqOcnW2W2qvPpEsxwPFxmGy0pC1z+pOcLid/YD
7mkocwItG0mc0xFjpQN30vJP7+WNB/Y7EsiSwAdhsLYFRzehHBlCWvHt1TCMmU/QDSq/Efxny4Pg
2wDLYe17dUstwuquujTGOrrunGHJA53gcUnl1Xp0jN1T56XysVzJSHJ0kfo5j6NCda3WSrujFQvD
RAqfXsVebFLun1XilqTt+GOoTVjUBqvhXK1vFm8LjZuiImp8avfdh+7QtTASovgc3U2TFLoNoKfj
ci8NN3JgQluchrwK7TlGP1h3JCrugCUqIjtBDd0yu22H+GUsmGddn2zBKUNh/VLk2sO2Q+uMWQd2
LZAIW9Ah8NcE0fVVQJycPdPkFSXxcmksmKiMv6/w50hTJ7TPzAS7x3w3M6PNzy0PYds3tUOY+bZn
HV+W/Twa1KvLpleBb4yq3qBNLN3mmr+E46AdhPDXVFRlVVqz2uhA7NbcPd1uRDmcc1EbX38jWOs/
iOvyI+0zVxtBpjNrDSFCc6YtsE2jXec1FQOtO+rybioCxyYxCMKqVLwZIRxKcXsG83dqnxhOUthM
bYlhpIWKZJFhoemxIu5EW06XJyX2d1dwnZy6f7DX9Dlv6pIpmB8TGlAZXwUkjIlSo6+kufA2RoeF
EEh9Cu207DY5rDQ8an0DWNOeslI5Xlx9tbE69m0uWgBCMca5oQ7YTQRjbeB4JLa1397n3X4WFXny
sWEvuIszRArVHlJcgE/c0ub3pD4js07idUAs4uVQoWbLC/xXrAKFDCtln3T0kXUlG9JIZ/a1sbk0
bLXIxhF1pP2pOhjihYB1YLqs4pdCbu+D97KAqe6tRFc7X/+ZzpWg4zaIp0fhVFyvJF/F+u3jtXl5
pDQ+YeRTag3gKkG0SyYubnbQ40bRjI0Nx/L+fh6+SoO30FHXSnmj1ChurcFfyxH7g+PEO6vsgoV5
LuZQFuJRMpmEw+UZWnlaYBbNPRXYngk1ocbDY9G4yx3kRp8lNTF6kDScs7YpBuciXAKBehVjJjzv
W+QxSltPJKGsi1Y7uscippWmsEryWIiorZsXkgeJLab0EgVxDYWgsl2MFvbQzGAJUIip6RS2vSCc
0+ANk1SIwhLOQ3Zy/d8ubBdFXbqNsB16PxtHcIwA+rQQXrMzZ9OZXnG0JtwSD5xeQuXHblPA+2v2
2XDC2iK0kkXIa9gGgJnae3wW6vYi+ki5uFCursYOc4X4iHoghdB0syDDuFMZ1uoiRKmofeRiHy74
PhSR6UBp8Uoa1FM1bU0B4SfV+9GDq0unPRp2aTk6i3dcT6tsfEDjq13M3RiU2JQH81zzU09uhJ+C
W0ujHKu4N72MRY+6AJ2Ah4CO4IxX2pxu/CE+MR4+6ko18LaSB4LIZ30DTLW8jS5hY4R78HzsBu/T
uF51OgZDHHYq2QPjkcb5wD3DUDnjbK1kmhCUX+09JJRqyDPtnCleeaeadzZA83EP68RcnrUZ6XHS
gIV9W0hOSXjc5WINSFHF8GODEOolSAXRhnMpi2/mpjO9N46lZtQuTSEbvidYflmgWc0qi23AvXF5
zZZaU0Gh1XNuwSgLBroXD6Jp7yNpg7bvfc1wNbIP9+5/ULxMoEBAfl8SPd6Jzw0/kAhtSHeOBysO
pisiyL0UAHm9ndki7/yT+MNzbG6kSHmz95fH1vR6M9D0gi/AxXDJOvh7zL+04fveO/5h8iShaU0v
JiqkImgjFDcz1hccRSD7le2GnaOx1t2KeBFVBOpzFEzbKixvuMPzfd/LFWfjqkO50wgVWJE9N5qt
HpOVFA6NK0zWaYSnfRqRUQmcPW5+Jw2iWHXkrPFdz/PJ0r8JDZF3ueKCfuXG4iV5Eg4RttQALyfH
JzVF4JJpxJWiGYGAFcyV8tgIR9HWMs5MaW1JW8oDulBzYay5mkTl+Q27iE/sQxyFj9aBUfTfIEI7
M/ZboOsNI1fXizmgnvjfojhcDL0hAK+icnF4fMYuEYfz02ERYBdCyPV2Afs+ZF3GGAX59bWUkYi4
SGvfcmUQdcDNTrIJKjAIaZ+N2tmECNf5faxI2nhqjPuxPNbser9Co7GuMVcW0rWEjVnz9wQCb1Zp
N3kUHKvEaTnJk119idT5R855Zi5T2cCf3zi1+iNSlA8oIoWcdUzG38Lx62UqLhPDuzc4KqWv1dw3
xJ737r2eUXmrQzKYRPNNdwK1wp5zCBBNnnCD3/n9PePqrzyy7Vp/3UrQYwYZnPp82Lx41nxiAjsl
lyE6a/olR0qyJbnKjYBShU+hTfmkaz3FxxLgwd6rNNKc49Vnu1NX4WZAhcfoL6UIu9Yyl/EtMAzf
4XE2hdEW9CB3LKSqDGCEdu2c7eKIjPDMI74VaDEE2SmdTRcnLYYD/hqADorOf7QLL0y/PNH8sKLP
gumj/Yoms2B0liWypMCyMMptlj7KsSNtwmHXgVTrFBH3/T4fNe1yYC2HwjL8mvM3VS7I45sCCo6a
U+S20Hk0lGu5cc/2OjpxGPAbMwgRDIdG9i/Vu3zLDZj2Yc6+RaQ8EZeToh7xVJFKYXolZfaU/uBC
JxcPL7TvuXfi8kfXF/h3ky71G2iIXobGTAP3pC8TyrnCxFpSfTEBrD8CmsUVkV6S1l3RnldEiZ5i
hHWrj7r9JI0lD93E+t7L/WjSQsjwuE9K/TMxMJdx2ftlHQbzSRDye3eoHlJuddepWexKb1YX7GCY
uX2LV1AGBUuU0ymFdg+26iJ8tqzcSbQQYj9siXxKElX2X4/ck0PGbg7zh0zPyEjW0FZ2aLoR9OjQ
IjPcxKUFolhN4jKSVAf8YJ1W7kVOiSjgmpHw8lEEcztrsxk4vVwafp5gqG20nvFwZTaiRNlD9/Qq
EWZeiP0a28RP8pfPCoMltIOUQwvO+jc0VZ/oRwmgBkzZBUW1Gi4wFWOlfpgHUboTiW31jxVCTEHQ
92lb/EivABDH3iB5xZX3bFIWWykYKaF9mgb7gEYajivnDxPENxMvoOtc/NkbZYXhwbzoWyadLNdf
YlnyGOzpZJTZeOm4gobM5YzD7sbUzYFBWuC5WZCIi0vNur9rNhjk87CKo1gafvMqRTVQEttFFP03
risa4JNkVeV6hSNixgJzXsuj8UVoyDaXk6IYzWLQKrCdvs8P7tZCEStuo9rqhdTRpgTGEKoTcMrE
fwr3JAZ5JSPjeyFkcyEMMcEVkj6iAXAofYFvWjvmQHbeGeJipM5qHGKiqh3gGYf+Uk95uCPsPIKw
R1Vh1MZkbmlNvJxte/YDqbtze6381FVajIkwlcdD3M0E39jib6koRoMPZpDaGLiFslPiKfb83YIO
qBAYN7P5oYwurx3Zc4+5F6pjZxI1+i2QWztlEF2680thTBgBHw2cnP5Z4dIQq6b4OkoeD8cWdjd/
YMctxke6fj3rgIM9P6dBdoDg+ygEETxZ/35o+e9OHK9oOThyvl0dpIbfTigcrY45CHLPs/aVG74C
cpkyiX55lIktojcPgOUhJDoAdQND82+0WEUpo9587VjYkIjWriYtY/JpPy1leB0icLW4EadpxswY
OmGacbpU+dgH3Y5mSTMbSCEH0mDQGQAa9rHAqlRcR2EXAvvstNbhLq6BhtLKRBWSB+zShYvpAXwR
hqdu+HFsz9qrlB4GsJUT94BLv92bd2GDFJd/oT+fc+d5qaoUwQnYycI6gMICkzvrVv70J/vta+va
mMntnAM3VRLk+v4jO+UO+0ZFY9vB8BSmBjKxa3nVFwkTmuiGX595ubaEX3nwfR6xMh/d2isCPNil
olj8JTOR5ECJ7eS7Q5ia3lXMAkfDRct7ylcm6pDCxwwUrzcj0VgSmDGBAsaqmz5bkIDSE32UYFgF
gRx8HyEC6BNTv3+LlIhNXThMaYGFv5WX7ZVM0KwLiqDr9byD+g56vO8ex/ImA9r7lyKDv72RNdBc
II3UXFNglINqlYAveffV6iGTii2sWptkJzzQbA+QE45i7OO1E6LX/cJcKajZsRLxCmG6V/1cs6AR
9hmsV+DhwFRNYn61nQVonKMY9NTrp31KFIsHpwudqaBtjcdmxyNXdGZYASRklr4WXXLaMW+IE144
5f+5leuvkNAwmj9+HXDklEUgsHfM1UHTIWlWXLWiRw95ngABQh8xEO5+p5vEHGdjbwxeWp/tGLz1
rhMZYH2qjdR4MlV1CRS7CEWX3pEEOfltqTvd9nC4cJaov0Nf6efehloOi4AvdTHx9y/d6+l9dcrI
7VTGxPzPAVtJ+To24cznRbhRUhWTyOizT+sBKs+3ydyaPEpvHldUMas5YKTAUK5uUfICosTKyzwf
wn4LYTn3M0InqLJC/hARTsQQWDt3WA1RUhMG+NoCTAA7NdLReEGb0nSGJqcx7e1j56SuimmyZdsb
N7mjhzU6faX8+NobJyIyMDTlaux+qNGJveI65PGgsDjJuX8wFOU7zOV2keJjnBlNY39Do+TlJ0Ev
isMALdqnjXEsQDVsW9wTFnPOpf8z0DPLiQKmAw4xeTc1r2+QNLUkZuRBJKPFNKBPxQctwge/C0iU
Bijhqzjyppm2Vff3xqSDScTc/2N6YRiA/ezLa5oNzB5WDy08DWCgpmHQCROwdqYciG6SWFm7MmIq
rb7gYZGPC4NvD9aud23WCOBNJtPBrd+icbnQFUbwIEbp6A6Gphi3SKhCjYy/JVeAu1OZ0tI0Vhe7
9MkoGoOwNIBmIQ2gNrVlj+nDlGgwAJUxtda/WyS3oc1svv4gCxIEMw/OWFiE1qEPR/UFdyFt5qGO
klz+6SBZJ0YVWhabbmh66xV/6Xq0FSDuiiNMCoBByFlqFte/lpUNsPZBW//mc2wcd9PyMLKQ3CU1
/Iwup49cQ5+AU9mr47elE8RC91n9c7HIoqauPw8LwblWsQHC5xC47AsG3rziRSEIQNtS2F2Ga87O
zUacK2iA7VN6CErOweF/GvZR+M+XEvfR00MKJk6ZRebgkYF8/7xfVTaBpoVXqopkfJDj4r6pKQRE
nuhjCaHi4nrdWpBNaIV+F/wvcqOOecG009YAksTZD0t/awMzyvRPZsTzDbK01URo/gjjnlPhDsYC
DimdJ1gOBmhwwtdPbzJL4SBC0NIvMwtMjHBSrvMIoJyZDSZDbOT/MGtr7vhBDhyrz8woM28lHWf3
OzGZXW+FmT4HJNkeotvfFse81ma50+8WacQUUMjab8Djj+6BgJmPvFukPWPSM7C7BNBc9Bks9uJw
OtmyF2CoHSYDG6D0BPUDj1tDtIYk5n5jmGKV6iP0LwEG3IClhT3EBDptGvGIpb4RcsSIYJ+NgDbX
Wr5CRlcIpDhUJBuc2UjkjwjD7UIuNrb+/K5W2RNCxb0TX3B07N0y7Lc1glOBcY5ViMXcdrlIf/Lf
tZO1P/imtgpuFBiNfp1BCSyhWcV+Q/ZX2b71qDSEElJpuz0dqRlmDQbjPZFyD4Xm5aCMiWyPqyjs
5az65BgkC01jj0Z7YMyX5EBauzCfFkaQIPGfhjhQQO7cWMBdiucITGQY5XR3TZ9w05Xd2J2ATXwB
qf+yg/MmaPtWFux9kRiqYCWgdI0Sp8/zCtnp1O2PdqaVUe95m0cqpf/OWwZZNx66YQCm+7j49Ld9
4G7/GlyE5tRf8B889+uRRD+1R7Li9ymZuN2agoFqmLFKrTWNam6sRHYfTYmraGSJJAy4YqGYHVc5
K0Lv0NTWK1Iob866O1ePv0bgWQtQsEXbWNHQYajkVOd0MXQYidjh/HjeSD13bqkPpnHtGvcCgDVa
9Uukqm/LL4tZr1qYu0VtRwwtH90lyQa5C4Z1+LJlRuZzuuZAiBuBWt+hQUE4dXwBbgS7wSvkt8n4
bt8FyasXExtNFWYE4KIYUFUlq6VjKfxersLpGf9DVLPFPrtnPALvQwRXI20ecftCjV+/6gW0+vx9
zZsXVUiB31GB7t07aDph7EDlMQIIl1BsI90GBUJuE43AN8p/FR4J2/lIXLYkf4v8Tn0i7YrhvK7g
0tjfnXXOo7zFOKXLvbCRP3ijxIEJYn3hGueXbFcy0kkrwcgkO+1NU9GMPjSD0NJdkQx8qSXaKnem
43BVCmJk37sg23wiQWvELwMBKBwJS6n/SlcTw+NZOqZDc3oTDA/enDM3Huc+3hS9L4S85XFZw+Oi
LucH7pvTJP7ipBYorIrD/iM6F9M/aw0+SwvW8duIKJefdbSAI2+B1jPVb31rJtzC/QT8obQ7wME2
ZmhJZ8xOKAPhTpNHFV6Df/E37T8VDpP7ikyYg4GO+6EbL6r6iyCYgphgJKKk4OqxxLYwh2ad+8lT
ytP2NMpn1QXEcEQmY4uzMIm88FcgUHGmXbxyQO1uenDzvD8DF0P35fD1xm6bIrdtqQ9J+s5KEWDy
zFMIohzNZ9c7+KMDE72ldIJoODUdvO+cQ4Wnwsjl+klmjcuT+orxbrGq0L9qdUTwyLmdnHqTnzoA
mWnrdSpTtZ65nMLQiJP2s75QFTm/mdxbyjIYypZJQnHVErJ4JZ2yFUkDR64Fb5XUlaXd8yRX6Mya
Y9Y9JMclxzMraxOGtbvq1O/y0IwkMW0JSCKgfODwD9b0ARSRFmsY/l73NpfY8Nr9pzes4TwodIFy
6qJQUUqGcvBUQ/eXivJ2lmCHnjUihgNrub+sJ3YI2YK0KtgiSHW/7YLMeaXK3SytnXTbd2qZzdfv
ipLv2dQzqx/5h+qF1x4QOHqtqqv5F4gfxR+uY3RkRLJga25WaKGEhx0Tw/qkGFzM5peTL7NI4Idl
f0Dv4o1vj5jNAZGS4W/4YnabsgCGVublekGKlx09U18M0Z7fYOuHwXb3HtTd814zLt7ydO8MNgJd
EJcTiHCKi2nIGpQztJb/D0cWT0kvelzA+vsjs8oAHBdUHVWG3GcPzn+MZNWraXm5/DntiCKDxUTB
UhMjJ13VTo1Mr2uYNwjDPPqILqbHMW+4ZlWNFWaCaRhSjD1iSB5bJOPh7IZI3jv5AF6eDiSoNTLI
V3yeZOj7/j2WzcBE13rZdPsFwBDHpzRx3YQoLxTOd7fWvOR5AWCcc2hTL2k165oquk5F+8zGaGE5
Z9npX1wXfIpDPICdmDn6CWLeVrxPGF/YmpAS1jD9q3KNPAqj0spZULUV0dH7xispFvkvpQtgxnCL
MKceGo7y60QhZn77i2hjTCPYdsBPwuFbXYMdfuRAWbZKGiLItzI3X9tJ0VTd/dXxrB5/07dO8Qs8
ajIMJxfMK11Nb5jfZfz5XTkkpNC+tLoJ+WzFOrsUu8VTljPp8bkD4WRqR0nV0/o3OFQ/TMVmXU9w
Iq+oJEm1J6h1DOcw+4VndpbLqAy3OuE8MWCeDu4Imjrw1LJLu9mxJs2FgZc2Jn1587x/rAdqD4wb
MJDGmCTh/x+0i3Fm8ENt+Fa8lat30gFmM9PdjvSxwRFDn4ZNR81Vq1WwUu2IE0LZxh74R1T8cY9o
GsvH7OmcjiHob/l95PWvrIZ3QlsxFkRQ1NqKDwCVprMoYjPifGaHwCmH0F9FDMteX4HqDCbj3VBm
QCCs72kSLX9EjuGhrUY6SQI9veAadmUXeYW0ZXObnFYFf0dDBnspWC9qm2jwKxlTUYxdgVrm8jpT
gharZVhOr6C7yqMgFaFiUfbSjpvF0ZKvnRX94xip8AnhoXp5qgEEBcZ/wEATloqXTFfF0HjkeluP
/aLEQg087wGTaqsynr0rdjEaG7chw35J1/eg32gNV0seWOsrtBGnjkE3AvFdnOI95xLoJQX90aaM
SU+RKwK4r9K3NEc3FHh/YBrtXVeEECfwFkqrTQXZcjJ/KfDEdc2M9KcgZctmPX4pn2SN45xSOARA
VaWHuC0m8KQODhFsz80whvbP4uTTREDNHVxCFuVkbj2mRp/kePLjkdw4tvSuEbGB2eFUrxKQsDAP
ZqUaHlNbdffqXdGzWLf42YI5MdOfuNy5wm+IhgSTX+zSSHQ5lkUWfnq3UjLsKoQWIKC3hbod3kQy
MFbx6586lFMHI2k/8a8XneYcVm18557JaMq8LoDQR3R4TQjHDh48AYdHwVBOitd8VYyvENIF7EpW
FVYzfYb/r+HJMAkx4KcVrystMzsetWbUBJ3W/F18pna42DJgZCwEfy+xvPPdx1K9Ulg/KhDI5uVU
A1BQlPAMbxjn8bPZysOp5wzyii7kXOjtkjLGoDYrdJAAXTDy2g+4OXkejTOxwsbpK0Q67wc0V2sp
8gEU4LRfUr01kyEVTveVypzAcskCBmAeDQsud+/Ov/A9Z2IlapFb5FbYRJcNLCv8sz/ASxwBvRIk
9DQDJkci/1uXB7YDf2I85WoJYEOeAIlP3xZIKA2vsq6qPaHtHuyYqFQnZoUQdrJmK1cFV6E8cb24
zQmepuzr8afNxL6LuvAKq+SpftovzV3DzM8lO4Dd+FKGOOReqZWTi1wV2uuu6w9c0MkHl8JfeZRS
njPPc/CE04TQ6ez8VILtcdSOXrShNfJRRBsyZK9Yj9QHBG0erVwVSosdTbMHQBkkel9R4Mt84oJg
GpwnpGKKbL1jmLlbvQiOl0wFJeRS9PLVSgTOpT2+sbl9Fpo7VT51SHmQjKy9i5iIaq9NaOCGp/QE
v6p5iPCBTp7xBmRraovzH/Wue/e6jCGr4dnVkbzuVeHNRMI0MmflcYA8ZUinXMJm2JhtzqwmrvKY
gD961LldjTs5vOyGThxJihMBQjM1YEh1KmWEC0BtpGGk9hybZ4WjucJRgX+ghLl137jeac5yjaXZ
GWE+cqLEC1PpzA9d82rLefCxHvq4G2ZkErGT6jN4ZErtqLDbh6f9MlVDgHdwwRA43uR6kh/qWT40
j3ny9+NFSNH3mV7IY1hGFzirM/VVetvY1bvZVM1RadxX0wkG+ZUHpHyWoejN6JXaXF8LdVSgUz8a
ZVsERUUCJQQ6nOgzdJwJ7AG5r/ReeKyo4VPfKuINUrB28Ug4pbxKYYq5dLM2hvP57Fss96eBxmi9
aszjp0n3KwWWr86pz7Fbv2ov6BawCvbLPSv/sExmXQwvHUZvzzw7lAIJHyFuBDkXtM+E3rcT7tao
ktR4H2tETvA3SV1GifzPyUONawhi6+flqUHUlTvh/1Rw8cgPQTQu/Ko7UVexYGgnEubIgH6U5VIS
HhdBLstbr2Pe4iYN/xpPxL+Q5Jz8z8yeWlzoX9vr6AVjfLWwT23C8Lo0JuSmPzxz2XTLnip4pVKl
VCcczxUEjwIhwgD0iD5UCxB2KTeS1fVMH2GfQ4S3iCdNky7sAHBKZB9TgFcF3+1gRQo+ukP5Rqz6
+aV8AYGiT6scPcdedm6CYbjobATsatCVfyQ2Th8FLB0tjSR+w7zLd3xVsS4OwnNY6LC7IudT5hv5
sqb7NWRNQ7fncfI8SJGUppuLuYjD1cuPifyJCl3QXBertSNt1nAND9ZbTD1BQCCvbPlusFX2WMn8
rk2MKVcySeZxrdrSpyL92vG1P5Ht/AF2OEIR7nNRTwVjLvxXsYJ6PGXd9aUJqloCSPI5moUbL6cT
OytE0vbffSr8Pysn/YSdDcAHEKna/hzqCezEwULWsUjr+roZJr6PAY3tHMGvUzH4W5lhsAO7LgKh
n4CM4zFXimdZUpwxFF4def+GtWd094Yqk3YM0nDoLQcBPbtBBp1ruN7H5+YTLdHbnWK5Fy86ychX
X8sUsO8uBUdHAWeREO1UpbATMRClW8Y4ONemPOhWSouBVvCnL8cBuAHY/zJv8EUMzmJiIIaCRMyq
BP6GKjSmHuqUv08DAJTE3S2WcrBsgoPBIE6zAKWwiSfKBc00Ki5JA9AD3Vs8hwZmjLi/oSpuc2UC
sz7QJXm20Dx0X/IcEBL/wH2OhI7+Ac5bOEK0N6u0G+7vfuv7CMdpaXGMkbaltueLPEM2DX9hh5pn
gxJXx9gWAJUV913KkxRobvtr84Y0ymAyq4IG9DyjkSETevfbBzp3VLJRTiaR92ac7jkiopmnCLBw
8Yu8YUiqK7rHNYY7jt2FqkY2HZj0WpBaFA3Ouv5Jt5a4N5Fq49/w+i7GsOEMmju+8LqBpMt5rlwV
PdKlWSy66jlGF0xSzgHCRlVebP9JdakJRJfxQ8Rm8oKbvqniTGrhTmfcU5OoGY5AC05KCsV2jD9q
a4FbwQluIE8z98bV3uPY9MSFD1eD4UOBKePOQCvchJX4HJQX/S5r/X7giRhT2/12l3EBL6HA7xzF
iX+BvNMOV3AQQ8lwoJPyOT3mi6E6Lh80dIAvLzDutnHApboE1qZkVbQcoHlM4spqn4f64IFLYx+W
l1x4Bhs98J8Co6WCcM6MoJJJK+9O+acBHibZM29iXDO1yM+TFiSyGMC9BgexBQtI+3HoHqFLHE2C
lx57CSW4npmtB9sXSKf63z+n16Bey5kEO8foTSQr7qh+2oxtTavOko2lB6xykzp1pSsgFJUPCrQB
BFkBYi+fgt1wpo/HlpXUtTT+0LwIM3zf1Cp5TzMMbOHJDym3vg0Gz1xa+Gm33aQ31c9k7OfJ322O
ej/dYsdpy8zOQ68YjVuGvEa+bpDovkfmICBTtN2VcxvAQQslFPHFrJcY8YSiH9AysgFcz396+6qv
U0/4/qaso65O0uzOnRrR8w1B7MXaQYeFlj0McTJD1Ii7xJI/y9s/zGcaHdxHseZqsLC19tbB3S1m
u9NqOHdlV8K18m3dKu1m1w1oip5il2wxDZVBA9H8Nprm9m4YyAde6zyRy5s/CKS52dF3AjHo/r9z
oTJGI7cfnm45PPDAgqXK6cPXpumo1+J2DeQeD2jK/Ht88Tu7YuWxmpppjQTIV1sf+c+KHmdqXBaF
aUREOy0tkSwHHvWY6BO4HqkOQMLYcHxY8JMolW/xZ/wd0d/3f6aYOP9NiR4NSNTPSwNy4pwe3rRk
deRO8kEV6Mo0NLULhtD1HL2XFPvjoPNg6acS+cCVFRPVVSen0A+A5vJHJ5R9BCkNBktmECMbDrOJ
G7SnHeMzesKSN2Kub6FuIdU+2lQhrCfK76z8zqjg5TgOJur3MtSddQzrdVrrGLIZnnAEv1m7aksS
XK+xRibq6CvBmgECuJLtLrfp1gAiSeMlJxBZhmT1wd7+g40F4I7BZVUPiJmf2oZfodmGayzmzSEO
iHxdQJiERkOsnbnz2y3qprIJT15r4u0CKD9pxuf3V8C99Iek/dCLOnenI8iC4Xu1hzGYxPFeDX+P
kaWwUozOVd4/9kiCr7T+Wn/LPoHP2C1/fd6CchvxHfj2ARFTfOF71PKANfBT/9YyIvpSIYIpZu0m
Mcep6ydsymfv4t5BvSDVbd/32IA5LGWnNqZFjVXXMU2sexHy2LJcpTQToVCkRVxg0RpFyQNsI9VD
YfrRBrQL4AmqPq2ERHpS8YZ5/3cEUWertZuM6OnA5xEb8hd5oZHgajE7YujEr3m16HusQseJI6tU
Kngxm9bgnbUcZ29I4icaL+HkMaAW/tzU4INThoPjq7vhNXzmjw0BnHDpHUXEftP7aB2Msav4QNpi
KTyD3rxhYIJa4K+Hl0w1qwprjS+32rdi2TO9hmXQAbvUX+HvAdpYsUhWhvixgydpf034iK+EGau1
A/F9nRZQ0RE2evB1chGHe0A6FLcB8mIWiYE5UZAY9reN2pJ1cVcUQrd0NQ4AKPXBcB3gRhGqvV53
OBbkhth3OX/Nx1ynmRllSr/iiviZTiSyIUZWfIGHDN+tZMk7TQ5KrO7S9H4L8rWUGcMw+4WYFH2V
mGriLO2VGsbNGOiiLnN53MlntV+s38NV0xnw59dxRRsoERB2E/z23Las5igHn8afKrR3KaGcpCvA
U3mOITS4aF3L0Fo4g0BaLnniGQmsHmLXCvk0jvz1Ny/6ttQQZSunxyWnnxKZhtGoA3MthYzQ1gOZ
5tMzna6SpSUQZaClfSi4rDdqhi2yNsbXm6fPC2oDB2PjbYZD2VyYML/GZA1FEwssiQsSiNX7A3aG
NvirHeesdhgvWBwvNmbhqRTwD4uOOmzuRCbhhXVPAI85FSfegM0gz/IGzEcCRM1LK8G1ehJT+WEu
iuVzXnmddbo0hgfIKKSy9ScGYfLg4x+nP4Lbdgpac0AhU5u1J1qgrVHPxjVEqVzeT7MXIAhoHrKI
9gSxWli/4bBoHglC8ANvkzhgsrnoN9W/FHhJDyyKqWqbiae1CxS0Dm4wKschAdJQzf/MfUjS+zWm
FzH80/p+PSeUBAnxBKEcM4TEocsT/nV7GgXAzXKGNmtcdClTKGAzLzF2hNfALmBSyBpM+qEzVB9P
Gpcmg+JYnPWSsYxesua8WxtksxUg08K7Y7Z+r7voTYSbqV2deX9vMvysyKIMf99/Lw3jKNDgaElE
v9X7NmVwN6kX+rdKXa3QnECC9he5zgjxKk0Tcbu3CH7mfMAT0eNViX6/+Uj1zfMpVb6dR621SIQw
WLalngsQ/aqM9IxfRG7WCX+uIir3k42x6rguvqQ9bNXtbrKqpXd9H3NYWihqE6mkVgUs7IQ0XMwR
J7BEkGP4yW8aMlxats+gr8crbCu13GIgZFrIb3Yy/zljPOI6Z4+y6L582ffISEravYo0904R9CIR
zfaq93E8TPGVbp3EjaoTR9qX3fmfN6LMjfPNyfrMzrVw197J5qK2tZTn/FmBxf3B9dN64lVTurV1
Y+65l5i11LA718yFdvE6neulG/pAWgP/8IPl8WBGk1SQd240dEXweOyHmAfFPJfsZ+LRk9y735Na
jjEh+eTUcD3Gyaw3y5PTjFnGwyIsGfMm+/avg+pQOxV6dy8QIdV1H0NU8fEYcwTqIc2xyUjhWHoY
uvHef1qjqx2mWLS/nVE77VS1diHaHy6pPWOz+vHdAeX1H3E3Cr1c6a1pxjVFocG4OuGa62jqjJWP
qxzP4qQi1lGh/A0O9QfQXkjpUlhYjag8QTgJAXeFYRAyVKF9k0k7weXpAZ61ZjTvcPGc1MYntLVw
P2W2bEbNFVJJyykh3Pw/4SZ1tSCoEg85JJ4Kn0+NHjO29xvfkjy2TnJ+YNPtWHLDT7sDUUuANTOs
lwL2jK4890M8Ck5l2rseP6gCd31c/qN0CNpwQ+fzh8pd1KXkj2mapon5YOTmQ4YZHbvDM4RT06ND
jLqf0Qaw1wgCyGOeJRcANghl6iXKbDYRlCIqWCxwxpWVjiIDjDMp22/pITrHwnlwHqKUPMf+o7dI
ZTX+VueCVN8qnJ3LP2ZLYZx+N1s0ADFOd0hZQ0/5DWXMeYr32VpspjXbqhRJn8FpMeQ9HMIo8IEl
6YNWngb8ojvo4U2D626bA5zkO75pjsvgZRdpgWgBcCeiBws9wwYneSteB+ZYR29gg21rm/CGwi/+
wETvqXgEajLX1wpmN7dD+DmoBjc9fhNZoFJiLTgIP/3K2/zBSVEWbffspiwqavgIY/Y0r7a31exh
oRLX4C8ALa4nkwNBGD+9k8mXL29Xm7hSvfCkibyaakcZqUiW30ziKPpsOiDA7R+M+IvGB/iM8vuz
W91Zi/M+dQJDUmrsvD+eojH7id6u0I6D/hwf1gifrjFs/Qd40l0NOHgeGN6W1TOVcqVSwhpppOU2
YIueKUhN5dLcPL5onrZTcwWven41epBqPDL8C/HN+LfGIu+sfKeKQ4qvePbT+uzz9R0gQtqpV+WU
WzrZ/yUS4NHQQ3mplbkvH+P6P2JGaM5bKiZA7Nf+OL7Rsf3NR+IQ8bFtAkJ9psRwvKkiAmC6qY2p
cVIElYEbXKqjT1UBRdDU/1RPMK8eqTZ9cAucNiBaLCQBp/G3Zjp6RD0gNFSmK9wUYgmYg3hlteDI
Hhxz60/CXSmb51fbbfy5S0W6zi+AShZtMZp5FqeBW91Pq8wnGzfP77ZH1cPkn+7Um3TYa8s+MPaH
4OJ1C8WYs8GyTxH86wh4FwZXRI76Uapjiy4YScYqSUrOeMDc3Jo4RnkFZ1BegRVbfcmgfJLpJZmY
ymgtYCSIhVH81f2u0PhH86Y+JoWCoTIWZNmETacbXk7bNocGLjunb9b6r5hNEeMguGZAm4VnNBVt
TbZyB9JZGWsth+Nem4ZSuUhE+eIljFlMD/W5vh5QsgSYCs7EabG2vkzyYf3Fx9DHYh8OXrNOe7Kj
gJuHney+78cONRoN4w2hWESjKIv1ARmCOcFxrL0I6M9WLQSeUM8UCeNOV9h6hxnq99hkYHyeo+Mb
tvdrYDOvgSZauzoAhuPEhW4fW567nSkTKmcHaz1oxB/59le+v5qefXchx1cWIYRlFAYlp2INVjyW
kW49lLkbWrdfFDcdBAUYqwIgsDDwabBSCYNgsFjFq0KRRx8Hm2D97meKjzoVyudQfqu05jmxwmx4
dDSymnnhyfKId1HESQnXXk4XZ/skxEovbo0JBOVTk+KtZS1Mmb3ZBo5fjxx2lqRKN8drck6e2LmU
fYWKOGy5xpA6i32oGpsBltRtOQsVuoA7/mEz/LIrm1ByojqELDGy5dPnBnv6AIzDTpFvPcEpjDDk
kndvp2cndCo43QmZnp9n60Av8KbrCiXbGH25Jhwj1VXFJCqJLEmW+C9nHfeNrJSAbW4RirsHVkh8
LhrzOGDZyRbvlJxnvGkFezRDE4g98E0+3bdaElFT1ZsvGGsvTb5bN9hfLnDvrWXB1U6b3Teo0sGo
qyAUFtS4AcWITF90crxp2zlJCVjQc6prQw8NRUE1V2vitDfx4lcD+1SuIqMBCuXFeeLtJ6D13Pqw
1OL2S69wouPLciMjOcDK+PMCSg3f8SuNYzEq45g0g6CcuP5ewTzC6EHhnpiSkZtLtJ55LP5YqdNr
OgrrbQtIYorC96kuvCzc3uugXtgVIMk2dXi3rrojC2WmZYHpDpNuRAp5+KL9R7PyMW9axSQ304xe
pk2J2TqDrrSPN1q+/eQ2LoJBQ929V/Z+j6HA8neg8nrdHE63D1J92cVEohND0ADv/qXEqfIvw6iF
UAr/QJE9qXh/2kx1vC78zCijFut04i745BDE+K9JpiP9fCDM5uo2QS35hrtkPTsMQY/4ZyxmcVJf
6CEcg26wHPCP2SVV2C13ejtNuvF+oiNXAJiHZXL7Cpd6XK/6fAAuy6QwEpRoMkTKBRGWVdauQoYR
jyTe9Xnb4xQKxeYQHsy6YTdkIV2d9h3EuSWg13mihTRHMba+v4dffW1Cu+Ce0fIUHLbrIPS5WYwf
5x5O1NXS+RIxx6fxzOMEFDf4a/+tf/6tEMQw/OoWbO2SI45KAnp36ualnMX4ZVYvyJ8O7411DVgC
huzBMVztjtXWgXLeMmF4MbiMGg9b9FiyVUjmiUO29m+YELd5WVN6o5/VCdGKtanQwlwZYsoWbyTe
PPoa1CXqUJDUWincyzKJo4OZXFfaq3jW+uQNv8w3sx3xCIX+WqokCC7dGcW0F8yLWQLaMjKeEM2y
rI5cqTK+HF4fyTJgREAM1A5wMdaVD2Hdk+CiAp9rhf7EpVdYrf8ut5GZKpFP/d7wZQiRQxBCVIeA
E8bYVFb1GCGQ/aBr+BHeydOewdp69vjghVc1Llutp4999mAlsYdvZHzmTMXbLRR6rexywYFlD+5k
5WGwdHXlhZNMUOp0FaSucXf53qBaxbDDS/B61cNwzEZaJA4FVo7RtAZpbalCyIy659OT4U5sJRln
LsgAdeR3IkpO/urbkWQgo42jFZvac7xcOgCpXVrc+KC5R3sHN/iYsL/ZQVcG0mFKU+3oKcDvFaSJ
qSgB0iIpQU9r1gglYBEfzy+3H34Snk/SXrkbcZCIqYUS38QOf+ulxh1m/12XlfKDBfl9aSwWHOzN
Acjn3AWS3ZiYaQMb/a2SVcZFbXaEo5o7WGE9dr5PHvY8WizfbX5x3pXP7hXqBUIYhJG/heqoH3GU
22t6UNvvdKj9YTnLPoAMJC1U+ai1k0Sc0y9HU4wPbyCjFTWhy65tjrxUo1eVpUp1Y9mEjj1jH/ok
gJHDVpn8je72wpC01g7FQdj4UqQHkAhzgGxDHiNRykRUzJnJHactByBtbhnIDiaZcB0HGNPONhSW
hzzOxdAFhLEKzZG73UW8tbVvrWdYj32joq9VuyIFeKI51u7EJ/Ag32esYGgDoBGDVSl5EJmCKJJU
vxfdnDK3fwdCv6moy5xvdnVnDrrZ81qakqz9+Twlm71DV12L++n8d3p0OKz+5ZO5Vy+KHqwEW3Ws
QBqVuvZSj88ysepDKHD8LE11v5Ibh4w+GhQkO9pwHiFwW2/Zkr/v9HIngdCi6x3nEuOrWs6Idl9m
R56vQ40SKOLJMbZ7kNGtGhT5VMv0Opr2vhePpp2/4yK32T2+JXB9xgAQE1AcJRhRmr0xzEgLyJW+
e5YK7TIW5EigjOZnFMvTR60lm4+228EqiP/2R6vZ4wKHHBRId/xEyrq2nJ/f6Qv/Cyy6JofXrdcl
gbL8P6SpxO0qsdkWfDAYEXspQA6i6ChUvFxAoRKrvb00AfXob1H6UsD2iOAc2dE1lgd1C+OnuIvo
LOgsYIKtQlfWQGjSQQyF9095JsY/v+2sI87U4IyyXKmcZH7OiH2mwlHx9Z9DB43fqAqfF8mD3mrD
mTI2GKj6vzhHsn4rQbPq5XdYJCK8thIOzLwj3ObqaCichjhYzp1W53zCRRVQ87YVXnCgoLUOkgtJ
TJ9Q7rY97nSsSnNS2UtbVRQN94EVn0XILAJRRUmRYX8gi3s69oByrfFUsYyPu3pSJiJX8Dtpl/iN
nq49onNSK3eEUJBPUGD7uePbw7bRzUiS5PA0RiP02wAF/A3HkAtUEtvtZ3pykS9PO1AVaavMtzqO
X5l0K+ocs/ROohUteDYdEARinIOlumaOrQmpEBLz8P1F0msRnZGTLiDe8/aDeuNGubr160NpCjo0
cYOsJ02PNDfSf3KEGKEEU76Qanr/cEfEo+uu6jBWEnh964tHJYNRdR8DtMGanGQwWKV8bLlrRpeB
Fkz85rT661OpfMtWRFz3khfDvs7L725P+ENkPEI7ca9fbJpGTDlz4fzyKkvBZlLo4HO6ld1wb9ak
aQBQbaQC70LfS4f0CSwm3V8Gm/dyvlP7jlkuE5D6rKZkB0momj7h9G8r/rHeCZkUjj9bK7aGzEyS
h55jwiNQ9olsI//Pp/m6PwPkQYWtmRwvuqIc0Zep1o2a1G5rVmJtuWDuEpzx/vQ16R/Tjcs8FIHk
AYVIX7Z9n7lCVE3443kUwtUJ2Gd33tCRgcP4PZMm4sQfAnOHuwOwmVVwVwoboW+HnFuQOPTzvIKL
VS3rzl7k+PzWf6bKBz4iK4Ri1zVKJ0dUuOjTn6neS6PEcKRIQnBZvQkI3+8aTUeI6aVM6dGz1UFt
zwyVAkB4gJBBvRPyJMnIVmG/3DWdZ5x39YnhlWjiKUkd9apxHEvfa0o+T015+7V6wvSN6b7Am6y0
XVgplo4KjBxMrh2JUySE79JuP3t+irWXvtMIrIMJDFnC46hoUkWdrBmbbXKryaJzg3e6mpFL7PsV
rt26G0yqLfiH20yHei8545Mk8gmjAC43nByDilh7kiFQlwAMkFVAoey5qn9KpvG8cKGXqbkHscr2
xQDCtDOyfJ9eAhmQlWh3PtxENd4+aEw9g7j3sexfmUtWt7vF6H07zBGJqtakSIsyECi+WJr0zum0
sg/5SSaCNuFjtfxngoM8b53TOcf1yxPDVl26sXXAIaoyZnoltPYvSDsKI+czasehnSa8cfzzqeVs
c3gEx5e9AhtEj/nar2YLcF6fX4cpWSCo8qfEFEHxtL/MzTqRHuYCoG/leglOv7L1fhmI7cBHuPlu
in8YSxCwtI3Xj352C9nC6bnxDSStukYjJTh4JLyIe7CKdsKFOHzRTjw8rDxAhz5e254B1BXIDbeX
Svz9bRFILGqw6OlqjoGNxcVUX75vkdJvy9gOn1CHOjF1sxtkCuVkequhWuEVVHjcqX6I4X+fiqo/
GLpKOE8ipQaBx0vRC5Kgz8a5hjlkM/pGjIT1LEmZqXj/OJ/zJXkihZhebAVDqOn6YdAwig9T71M3
JCpigFQG4d7XSehoMlosTkDBV5WBQmcaMoIuj+J5ewIpFRVYPWwxzh1gs1L4YoeoJP/ycrVp3Tfc
0jO/pKWQUs8WU1wKWiijWIr0dE51FqQuJTlqrDwybyNIHpzEUPGyhBnjO+79QxKmJMlkQ8BjdXFn
CO5MpbReXY9Y6wzRE64TcI5wW7rOCqkOkKeuUjQxgSCqfrYKk2EsMHhNg+iz7+oYJ+KnUk3KXQjq
Fb6GPAfNRFkCYyX8wgGxfWosDglUtV4JjvExCbyfNUZiQ2PqQ9MsctSbGHXu7uXAgwsX3jw+p8iX
h8C/2iyZzqFqmycFEdbicqUl/P5PikfmmRYov5UnMr5E3pWVufeAh1K/jZjCtviLTvmx9p4lhQk2
FpjIVuJ2TNhiRy7g4IBb1yDoeX3Kc6+XppkSpjPnW2gbssE+ye6xeUYc3bcyu3eZO4VtB6IUT7RK
VKY+bM07Ll0vsC34ea9W5pqab8Sl+d/5rPuRtmCS4NhtWEQlCbb4WnUi4gEFeUEyc43K3E770NJa
6mRjj6vf5MrZ3AegI9P502oCOg0jtg37RWeyV6IrhqcCXsHGIyffpnZDoS+CUTz6MAqAuk3drv92
xNOTtcjeN7sG48FkhlDbUTpvyU7fKI2Gk8r7UH4LwV5aVmCjenfynnjEX1BGzBkR2pataf+hyFrN
bcZcixk/bB8DjXWkkXeVZTfsrN86aY7GtmWUwuRrrXXXsGqiPVjyAodnbeqlj9/nUVcx6hF7j7uq
g7YrCTu8IztL7hplAQAsdPW7CWIqL7Xk//5l0zkygfVSrOcZ0NuA2MUGov2JD9MGAthvzzb+fMRk
tMEzAFWw8+8t1xBKwEFLkTVxH7PExNTxFVBPXAuJ5dSeu+D9VySFTpXL/hc6wwyDSxqVXB6U1W0Z
XVtSq5XN+ud4+wgSdbiymgA6QbRmuIgKAU/KH9klSYppXe8oYV8fPIEyWSnfNy+RHQWLshuoqZip
73KPM8rE1vxnM1O7dOkaAn88QN5frCjsguR8J6gWTQfuv0KGIeG32eW0lra8TEquHgTfEwcPcuI5
LCRPHQs5PtI7uqigAVjXcg0rLQjAg5WBC9sHwf0VTO/I5RlTOa7Ytf3/PvQHh345BdDjmL9j9fQt
DNaj5TVyy0iUo5Haz9Qev5cEKzLA+i8N9EAPEn4M9wnZVEc0RsGjPEERCEXaUT19YfhMjUpP4+rr
MSYGPX70KzAwzcXlaSn/LAtWglt+kDsPQVPe+CWDcgehv1FANZvbiRn6wtDQU1vmXCnIFO4zD/i/
zmgNveXAUlluDpitSeMwsda4G7oj3pIAApQtHmNtf/PyZ+3fQ7gVoqcmGMUA/GWby7vSh76O2Ejj
NiN8cMw1nCKAWMBeBiHvJwGRyWD4iQ3JIAZGkRaVcd84GBWvXLWknwKnjroV8Tbxrgt0OEUs/eha
lRTX80U4/8eWj45mrEjWDrBkXDKMqPCK4QiPtoyvbTTKKBzUzF8ZQhDX1mvQ6PcIGO4L94XzSOQA
/GXRiBxCjdWZZaqAHCHL4ApsD+9XnBm3xl9keBn43Nrir96zTPGMq7UYSlheHUa5Z0RNKrMrjWq9
TA/vT3vPqYuiyvyaHEaMF29i1jDhzfsw65GL0v0I6EklRZEZLE4rDEfxtF0EEQ40DuJ6S0L1MKxG
acqhgTgdElzQGGX+8KJ7qpra+bpWfo4RlTv6RZwv6jwsyfE7ojGFkAJW2c90uTM7/IsxW8YMwpJi
Y5YUmK4WWTrk+V1jWc+kswnLfsnM/bJrj6lnMbbdoi6Vb5VGByUCs+EXWpUDQgXniHVtl2vIJOtk
duOO3gF3ZKHE6kmYHvpszrWaKHEwxnmgbftQcb4nVpC+lQb34O1N/Fy/K5zNH0ROIP9iN1xfQuXR
ezyfAD+kfoJ1Hs6vyg9znMpgB285UghYO6rRhCixznPyX/XLaqLlf0Dj1liUYOqVxkzOsLz6gfEs
NLWrf0ay50AHimTyPf99n5DIy1F9MI9ccGMW66RQaNJJzKOa666EMMp9QM+TKReFuOgy61CBQNS3
+MvQnpD/7QvRHpE9lFJlEsLRFV34aRwAYxIA5E2IvFBajAZU0XS2O3j80wVAJjofHpETQuCZFOjo
r7mq4n5XvYthcG2W26HR+G3QlKTtxBEtoxnBi673fj/ZFhRlx8mkAmqUuG418id6Qk16jsmW3G/J
iFHBpBvzBOrNPt0WnHJQUO/riSxELd/6pr1HMNKcVs09Wl7G19HjGJil3SVlAb0jsDQ6u/xvQ/XB
k5I9Esk6m5iR7doehSIyFhHQehqmUWAUW6P1pTeUwsUf3u8qU37nES9JKGQa3xjGfXZjN/DnGa+K
ksPPLmQ2ZE00wRfM5iqn4UWSYUlnZmXuCVTKvDODWzDqk3zNPIzM3ZlalR2cM5ajsOTR8xEGXIQ/
GnPWT+81QskKCn5f0NPG/s5CzgptpuVJfqqGKXk2O3HrQA+tttuoHEir+GGcA7xAdPrSmWr1kolZ
lZAUAbukJ/zaFeqR5q25q96pHfNBXahMTN+gGE0TKvD2nQ9jRcFy1CUFXagf86VQWj4QTmN0OT8B
D9MZ5AvYreSX42rM6ypTZRQKtrgoxjFoFNxsxXL6lbpnUs9LFSc/Rt8lPaKpir0ptBubDJD0kcRz
kKJd1crrmTdgTCTcRs/gkYYiBUHUfvc6T5q4nsLjAye3o4kmwFTzo6ZNQ63coYBl5EGd+THAirPm
EXKMMdjv6rts+vBpbaTpZSvNLRMqJW0t4GfdoJF1e8OduYdDVurZ5zeGv7ka7WsOpZsjg7uMWUMW
jbWqUxZt5sMeMl0pOs3Pk6OqYRTOuI+ZsjjdHl0u7ZaPS4DEHjKvPMznMfw3u2381ByPocM6eYFS
napuwVbqLRTLNnKPLEIhwb9Z0Z60pqWPfOLRrGHtXjvIQC+i3ISpdp2WYnsE0N4vEb6d1RTD/Wgr
WMRMvZuHgINytPOyZpzPuw0GhCAecvSmrpNyKSVAJdbqlje276ZbBDzblsRswVWVqmYcfdSsdlfs
zcmTMzzYPKZhZRhe5YyauWJMQtgtchNKBSkUEE55zixd6Nzsg1sQgBI/B7osPgZSs54dezMsT2sA
K6HvmzIIqYAjuD0GFL6nXmc+7yFCzW+AVcBoijZs52mkWRZsz9tR9BUj5OZ0owRimFFI1z8QNl6X
klBWJt7kG25pkN35treOF5JQXERWaqyELrYobNI9YWIdNa+dUftvP6TKY17bEr4NcieUErz1LmqY
mAC9UileHYhIFM1IaK0JM9zsA5l7tyMDsQKzmn4u/M8rAEU3QI9zwVjKAxFZV8GMZqz1k4VMgoQi
Qvsv+Rt5n0JbK2xbjJRfgy1QlPAmuRQf1Rw+T6DMSF5K8j5ZEs+dO3SjXZJJECnNiv8WDkM4r22z
YFjxNvSyZiT+Xyb+Z8j90rNTmIYFqZPtMXxo7SEK+YhGCG6YAm7EwD6+1nnF2G55vsuSOlrNQDpT
MTd+/YqyifS6i9NUjWpIZIKylqdW7FLSEnrfq5fIpqgJLBLzAUkMTRttCEAWmObsL/dX9B/h2wX7
vwwwdRkxxR4Z2nBcQ1yT2nj4xgR2tJt8aayLkFZLHzi2dvDifBfFesDRBQQqF817iAvGHTuHoVwv
xINg0O1nWsSsOcIVti6DCIXYOjoBbz44oApxm1Z2KZSyKYX8nIG+0h19g8ZnDwv4oAUvpS9IokRU
Bsli5E04OPAzEmUBnheHDThT9pDgnvYZxOZcN5RfuGqrOVdGU7QmlCseshPT0ogwRI+GRkKfeBAy
NF5hrMNZQQFSKQ3hNxh+96Vtj5/IWRRbgxRvfxS82fz1ssrHXVnBMIgMqyCvDoch9pXyny/9hcgZ
utz11yDRZoNHYG9k0labWToQ4LoezqlvNg/ePzmbiwP/82yK1dyFiZ9APFP46X7DHsLq8QZCgBN5
Bx11jcGoMLxXFBIBFZ2Qvru3de/wP5/4H6+o2//9BIJubx558xiNDjjmKNb3rbqnlX3PHWiBeGQ1
TevnO4bjL0OW/GZsv0SjyKin9HQE312ADycsQZT5W43xeSDEjWcTfCPCM+yKsHxRfxtcKymQsPzO
XRrOq7WPwLSjraaNWUpeHaJ77HpQD1Kb9cV/1whBASCi7ftPfx3kedu2oEFij6AKDccdYVdUNTXz
BUk8z+0YMZL0YIkRZDwrcz/BcvBiURBeMX1kBvDLbwQkxlrOUPfo6kAvAbqGo/E3qWCY6hl9gKSE
FxM88cXim5qG/oeoATjLO8X84bC3DNzb1GsSEZvWu1Fok1zcSQc8Wx3U5BE1mCuOxHIAybqhYoE0
vqd7eapYPn3lW33RDsiJ+ysJVHQXCP39mSuOiV2DYiTavqQkrIxRf5CHsNYtirYD0yaEFYrrb+3I
cgKBrcBphCX3tshMoRDJRJ27Ejlew0hDqIP7gH5Eu0pfs/oP+7P+aLQKJPn/DU4bK5jOA1il6DI7
NzgvWbC2KVDOJHlr12QNchOXL1YW1e69Us+dqLPRB0EBVA6aKzBiqSYwm0Wz//Q7gAgCQ/nHcn/k
ha5p4VGHvTc3SmYrR6Zti1T0tOjtjp5Cs98/D071CIaHCy0/49xK7fRCgqaxgvyfuS0Jw6q4QgsQ
7bjfJa8/2k147vk3trgMtjLHLV90X6E+noy0Gl2hnPNqBoX9Jk/Femj0LaIjeJu53hRE/ewc6lC3
oNPXKxgHRa+yjSVX+wiIhoOjADS/qFqJ8N5QYZ9X70dN/QsAqeR9OCZImqJWXDTILz+FYVVahJ8k
eh6wCxJXs/hT992BiBUtoDH+BmBpDE6VGPR7Oj6NpABkSQbZl/l12HlX6Qdsp11NshJYV8GwMGj1
DQKCgdV78mY8lVvK1CIPD274OyGj/qThSzF5K1Qd5IYxEM+Beh1BsGEJTAGaWMgm1HtAp0xg2EGD
0Aut+kM1uTlAY1jUmSSmWWN5Yn9LSgDB0M592FtGjW6e+oR+VTuZ3KXJlGOATA44K6mnjXXNXyrL
tS1B/nZJbfRjhvJG/NDtUFrJ79Q1FnTT7p5mdx34Ccozx74KBczlsDkjSrUcN8UkQCPUArzHMJ0O
YLYfozaWcHC/h2DIPul7H1FehiEvZo0ZqfoMes4DBvTIFAymgn4B0kk5bSek7Grwb7YlTS1jHWDS
MskhjBSSgKUxwOw46ji7yzXP+7Krj76jPGKevX+LDFp+bBgqkyAf0Fqo46yrgFNI58wyfxN8eFje
uohgydJsR+TEI0YAhFVBx6TAZUm61hoYs+Vdj1nlUGKNc1nHOJCG0N4Rhp24Vruw96AaFX9MOwZK
4szc9Kclo4nANWifeStdnMM6j3RsmoOlPIZgFBBCVq/1pYTW0IoMgWOpdCKkuHLgWGRqSkpsJHrs
VZZsG/R4Xy27Ro9B9mUvMYHk1vvve/i/QUAa6nUsESY+uezTICVSnqL8EhengzuTcq3RvEuwwbrJ
9+B+KXajehjfz3b8Wr8i2kElAc43CSkPsYqY0nCrp3NvybZwZ5HdmXGxcvYujyBZ7Jy/lcWhPDv/
pBeKnb9QnJUNOOydCrT9UQz5dodcrkG7+vnb5aGlEUn+MonklQSa7ltsX1+dZJ5DJ5mDgErJqIhV
ZIzN3RtvZ6ZJrnmFcJoH2nJZoNs+Zb0RlFJkW9zaVrlUcarNL6Sqz2ciXZ4wmwPN0xwYMPA4fRoW
e8CWWeifKw9jN1G6CVdHkNgAYLyFJJqe2Jv2PLG8pWCb+N2n2lsD99/JWSLVz0fJZUoU9kERCLyi
pY4NqXcaiJLrGnBfs9l0lP3pRQ5S+TbqD54ecZ3RV2auwM+uh9ni6eCzE3AupHdLsMKYW72m+K+E
RDOnKZaBT+4FZbd0rFr/2T9PFQFXP/ciq1SyWCFVpf0tFHeZ8P8AW8B29sQ0JblebSLBIVIRviYb
YPTMP83i/gKizb98UHP7aboR9E6BYBs17+6fuzeaW0aj+q1D7vNzSK40wPlbILKIMSrWFQsLbZQ9
XZfM+721GlLiZ/32QMUl5tJzUuE7oUV42fs0GCSNyD8X0180qwxtG1RFtoXh/7vXrwIeksQPxl2x
hjWIwJ0+T158BNmpCozajhxQGcaK8GmHaFaMaOejRik3/osZuY3YG9nzUF0/XPMeQDoJYazGf5Lf
cKqQpRcQdNen3ssKObgBs+T0Vr24+zvWqhlsi0y3iQ2psRTEbvIqA7newRQ1PzGbZJi+HUVZJsSt
ycft7SHRKtwWA+ca01IssizCPeF7w4jJeAwtGhR7WWKlALMgZMXp9W/ca8rOYMupyAy1z4v0c7Ld
DzeVa6LDpsp43OvdP9Nr7/uR9r8E+0oI/3W7NmupZeqPL98RmfNhQJK+IB28EOMvFQUFYGByuHOL
DU8K4DEySRAxz1YtgsegdR6N/8IiqxineGWQ8teQuONI+N8yGyyLcXtUjVYjr+NnAHOzWByb+Qpi
hp+PjyAeHB8IPtmKbjtwvX9JY3thY0BVAH7YO3inocVD5Lle9YpCinT6cp8QOj9AHezUZtRdpWFZ
mqIa20HpabXUCabqVUUXFLZGu8ctVnC29oox+bUN8I+jcnUJfbgpG1XfbY/tmjSri/Xuhim0nNKt
zHocd48nELWa+OuVxWkhhvpjElw7X6qLxh8GQsalZ46guFxth78kXZq8QpYzc8qGvuaEXpegZbb2
l6nQTBa3ecmW6EYVFWhh3F2REaBG6sDPv7wWqrK2csJp8Vxa+vGrVmNXHS64Tg4swTaN+cj+Y2fe
FcfDESv9XcB3c2KDwKHC1SmpjvolRyvhJieFwEgMifWyPjtm8sV3vdZJv5Ao+ZL5VtoVujgtRnQg
D0taKORyvDblpnRqc+0VntrIRXTMUSFlJ2WHRaJP/7C2J71drpdMkSdsplJmkIWanCMYhIklPVcf
v3f8vaxl+Wvf0AkQ4W47NU5qkmR2EH2txpb386/Oqz8Rbk/d/3+ryhPc6SHbD8cH8Fnr0dh1fqwn
dnoegJE3jxvmbbrkOT2HZzpAevMxFFn4rmDByYzEo5W1cu2m6cODxuhNEvLedX+5/XAnRlMrfVsv
nr2IRt0Q8nyKYmrBj/LyAwkVZNzgygHVPzXhM2W5cl7eDm/3ctlkeCJipJaBRMdSDmfi6xnNov6a
a/+QCj4V4stIuOT0hp1PwxleymYu+ChPkQkFDGokhWvOc0p0tfqnjET0Ly5rnkrun52cIhaCJ6if
sDUbbs4GawpJ6PBaKqDlTI/nIFehxTcBic4R6t68XUtOSqMdBPcxPzyH63mwmO3RKaq4+Al28E2J
l0O1Pe5GKfeZvhBIpXsz8xk8+yKb0/LHmv8GTQniYEFmgkfn6CcGP/GBZnN+xYCw603h+MOCCwWA
Ae3d/C0l5eHA0uAgrSapo6tRWHPcAEDhU+P7WoaM5BdE7AgMj3Ypcv/fbqK1rFhMmQ8qNfF3vHe0
yMhhn6Pku+quo7QQTveg3KRuEQr509CzjGzKCIO4yX4OXkWMvW+vojvotk//LLU5yMZ80orD2vMH
hKfUK8SvU3pSQDLv59K/GI33TM/cjoSnpDen8T71omL+xrrGAIqh5uUzXjwAMg2sruHpxwZCgpfc
3dDeRljgewj2135meCFmm4n4OKea1B9FoL6o4ZqDoZ+w9ffkZhc4s44tZsDJ8a6y4GDocYkP6SDj
iIITYX2eq1gpj2Gf5YVn7lK+tS8B10O9mjKcJsoYKtMWyQWAC7oM9OLkueCZ6V6YJzQudmV5H8sQ
nMwQFl4jWjEp/iZItZ2P6pTke2GbRv6cXA6YDQ+ABGgC2fqf7cCP1lLxQQO6LA/DgIFY784wXeo9
1CY0TxuW+r7TOZiIZsuLcdXV5aMDhM/ovqIEnc2ydZnoPhL16/DYbTUCVmtqR6gtdWH1g/JE5Nyb
gzRoYyztfseA6hyzK6Zcb1XMdGyLrtblisUnOcW6pCFT7MntHHirQEdHJUTuF4AoTcEHX+/htbqx
r9W7GNEuHkQBk2FH/uOEwCagK6qj1LNNjAe3XfrEDOZ9ASEKL87XJNDf6EIuhhcYs+6juDKJ4ART
S5j8lf1Hw1tjEDC0aZb0A0jyvc4nYM8o4k0GMmyYib4dyCsWfJPRCcYXumdaTA+bbTShsNkOMKdW
tEubQOX6/aWXkYkCi3UZwpdpVLw65D/yDCnMN8WHQ+LJNclV9fC9/qT1TjLJ1MXztLTi/trqsKv6
W3xI0nKVqMgH3uXc99tGCAJZK4vfOHyQ599QqqD2GWIrp4rKawsaP7+G4QDiauRlaFAbVKuYLP/E
SDlyKowmR/Xam91NE5utblDeTyvjBntMzPV6JviBsL0ErhuMJoeDrgBI7Z/02ff/C224HKacvLBE
UeHgzR4v6qeWfHuAkY0d8XVsEJvep5XK2Ysu82+32/Dy54OhdIN3lanyQvYTh2WfFMQEAXV9CinD
Y7hKPgIIdQgaXQOqqHjRFhqo9+SFsBWl1mjzED7nc5JuUtOYYy7oXn4Enhw7KvBvrmuRNP3627F9
zROHmeLkSwB+a0Ns9eVs6c7h80wFwLA76hb4HVx1s5OM7osS8gzGOlwp45ftueQFgU+DZfAif0o8
BPSG8fjyf/PFEIZwsmVqUE0eh0ka3vOYUETorvy3SS4I0NCccfbTOr8urjK3zoQXoMBrojoGy0gi
Qc2ZHgIbZ+fp0JoXr9RnVpN3WqdzRU+kKkDwDtjvSjiLjULovL/68ESyYD3ENO9q+Fp4bXyShWF8
t/ugPc4sC6Kbnwnq57LNKEzGgqK5FrXjiLZJIEmYMGCaxghznnr99LJN3p1mqPX9KHifJ/dw2pqm
end+hJf8bKufGE3yIm0y1cet1Q6Y+cRWzfuAO2J21YgQQk2cidTnxdJYKFoy4IUuWflnWofggQiv
7UQaxJSzyTPkRj4j5GHC4qFVXLFaydrv4pkXWEEe3HAC/8BPR4QJFUqPn90qHD05w9L3Jsj70kkz
9I0+faFY8D1K/m+LckBaGRL1yCFv22ChyM/BDCjeN2xtus9n1gcdhRKdzt3wy12FfN1kqi641wSS
d+/rfBeTfnSX5AnZAFV6sPJkLAhe8arQV2jDeOOX9I9HWmJW+nP9dj57wtsxpv3dQzQPCHrNkjEJ
c1ThETYnbtjpxyahOumFGQo4uw4syaEvqEL34y73a7A8C+Axi4Eu3oi4I+MI6MGrqYcFOtor7Asq
hdrVPukg2WKezEyEiQP03RWZ7FVUYd/FOGSmagt7dRLnJ5pmcN3t1EWP5Oc/PrVddOYodlRfR7Zy
WHAIeEtUwWAMmf+zQEqcd0oPFBrgwm5MmO/zR7HLObtx1rQFk4js6PVT9btYQ9qB8v/v90T7sPPh
OVxux8G82HfzUczfPypgetxbhE4M6M3abSJogapy60zRH+WTJiDsyMrUxV20otUzF6py/vEPOoG2
ibqrhj0CbPbdNQ+jTlTEJ2zpVgQFL6NgwaZQ2dXvyVZyEwFQbKEu8/XXxh10vXT3o+Z7/ip4odUJ
tTJrROqI7oMVL8Xjz2EoljiyP//lKDv3KyWkv3WwesMhX8qZVgx5CCPs/xLy7H0VIjE2wJd6BM/i
FNI8loZaX89IbXCqJlFg0BeIUz/YXNCyviiw5bHRjcSAoFyCRhWUOZ6RlW1S70T+yd/r6MUKgjpo
MNkuSfjrvdahDUJGUKvrxQO5qGRblim/FT6qA+2+mN1ihH591hfLVe+GGvxGm9L6ykV3PymOR6h1
B/dxgUDjwdPNqKDXHkqOVNVnam/1c1GmK+BAXAg/2yMPjnW9BBATnzoR1rwpMjXbt/jyuPccfJkK
sM2xeB0mNoDOX4i6vwPFB+lHlMDps1GVhMrE9FcnOgR9PwwWjAxz6ui6GE8ooi6ktPxKm9XCCdr0
31Z9f/7nO7RMXPxVmZdQJ54e/2T6TLNEAtjo+Y9xh3whuOprzb7vgPYgmKLihKdnwBrGVUtGFdIp
2K17Y260H9aNVkOwZVsGF3VSwGuDtC7wxq4VyHFjy7BJmeNsW0Td3T86VZg0ucQfN/IwcAXCVKAS
m+S53D1gA5uJTzEk/Qyw9mDCUWfqiksgVRVC0xOIUr6vICOjpHnnN0r9snX69pPn1h+rAjBPaK+b
1mkbHrhLvjBLRr4DspwTc9Bjja7CUgzhA2TDA7mJJgeILVAHp7ufIkF7CsCL9v/p/pepJVud0ceP
6xGlaBNmRCsFE5QiBjcpbu8/9jTInS40tPnrpZ/ngqxV5jscLifXQUd7In+PeAUIgKna73b9gzrE
H5IndPfbDOV8aaEpA/WeaqQg0vMvDuvaAIa39CKQ3vCIBclHcUZV1+ti41ttAYtOHhpWlArg6pSR
H6gusYOIdoLV9eMRE2t+pCtdg//vE1Y3SnN9ujvkAOripp7WKeKk+jbsT2ERJrs6XIBionu6feEe
IfOF2p7pczkBnhed0soZgI6ehPmOhSvtZe6M0GNtC3BVmUIK7Du5Q4jL3FwE9BvPbP5NT8eLjGFW
YAcNTevN7VrEny4c1j2uMC+4z5eqshPqAm1CTokyrbHZKeub62SNZqcTORt91ll6D6MpKYKm7GZm
n04WeECUdZDuU0KELYH9gVhIIX7RNepTgGLgAbdD7dlcaZof58bxUncedHzgLc6mQ/jI7/8t/oY1
4H6Nb8uMli6EGVUGaL03aSju5P/qj4CmZFvoxCaPOelFqZTkHDPWS9IqotVGFH1dZic+YbiFUo2t
3POYe+V+BKtO/4GM0YJfbyZqREAWu+KE1mIq3jIbGxw04LRAXMVqfPP4qtEr6HrI/3S4algWWDCO
NyCiu1n5HnXWSc2240rTmrMLKteRHZnlndanqne8WJJFBwHz83f7tPrByLWPnVOXgWiXYMZNWQly
HcTG7JbjeMU5rUX+DzahPn1QIYsO8hQuXHGcbqmR1Ag6urgGJpsSxiZh3g0hngQwX2rrlnMEV7Iz
qtdpOh1q5vODXLncAIbnBuft/4jrSNge0oYmFWI5N5h3S9ex+coAjNMfuPdw1+Zpgnd+xOyhc5Q0
FSDwxAW70tjzDzf2mMss+/grEPiaq7BzoKGac/2UwOKIflrxIhsYXDIGUpputKb1cjcEfcrrNsWf
7t2bTzg2DCm3yRCsQcgI34wbS52Tl3ORtXuwwM/tA4dQ3aYQXwgKumJ0tEjLKhmQOI6WefQnr7nM
/DzO+U6PSSlMx/YfTAMNuv0Y5FcGE4OiCP+g0XS3gdOMsZSR/KjQ4neYIHqMcLLijcU5JOZcPxa5
VnH0neUqhd7VTnG0BQCXXsNOMHw3bAWpdMawzd1Kfpf8WBWTTAVlff7DCyk7MX7sBrpz42Z1vJdg
gk8VMCtL+S9C21CCulN8PaB2jEnDO0DKtQxPawaiEccndDFiDskJqGuFE5rTuv+ckzB1qMY5U87r
XAks4CuhHelvLN82s3XJxjtk+lhYx2OoJFZn9vQTmjEQ2YSLys5GpWv+XhCYyLZhT0foq1UcloQi
ITTnZUDu5KkCZhpatkzjaVY/FOXLLPupPYSe5pIqpmUDTilcHFnmC//K7qzfMComntRY5fEOKIkG
2JYTfrjayzQypKnRQe0LcwsBkHhFrmxr6CEb1/drEtluSBVE0ryBL0Dvsx/rN/fhzHUtU90Tk6vD
1rN8m8geuxEXHDAJHqAjMwhye6ADUB8jKQgZ7o5b5iwVMIJlOPY7bwUrqLI1bhmc8rapef8vIZDe
9Zu0FoXtcTD9oSBCUXj394KXNxKZErBtyUxVCMwiwD4pJwNYZl/B6JjcQOThL5Y0wLAASQY8ne7O
jSAnlyuEtey2NBxns9sHq5d6TE+2p/KoJ5QZ3/k+18uYQJJ+kydvDON3K1hUglAnk4aNpaoEb1ID
bAHLO3wbeSIlWEGKjGHGoLBKhi9Kui8jVzSrpkE12MTE/NTjYXNQMg5zHQqTAAUxh8wREPXkTrFC
tl2f5WKlhoBr9w/LPhyHY3gqoWHmUfKv9Ojr8vLwBIhc342nKNEierWTwyH9x1Ckm/wujfj/g1As
Iyb5PlZI2y31ex6PTAu6csHSj6fSYLRAsn7sdU28aSfVgv5wVm1XamsrB8Dw9lhM54yUWIO53tLP
nrhCbul1pNH58dsOdFLd3i2denlO+0FjxE8QSAkpZxJaJ4sYaFp3rUnFg2VJ65JXc52PgSkU+MIs
e8k1Rm4ALObKwt6IZurF4kc2RmrqGHAJ2mSbVtnyQKlPe8pSjnQ+Ml3a2b+ruwB6CQh3HArpCxvB
KW7tA5n+l2ND3fhNIUpxWvc6AeGSxk7EfSEW4JLDNunXqcJdKV4LypwQ76CpWI4zEjPcTC7qbKXx
/f2qNMUUbfsDHGrVFP9PMyb7CRcrRh69ghOxaXyTcNVDbJ8PJ2xJsCnVwITpbUSxKYTYiXZlcX+e
P56ggw3+DdTJ4gtfHwh2WIbAGpN31kT0Wwnpy/PWGT4+YZD5QX03kgkDDLnpLfFREKO8/HjCLQ6O
51eFXAsyuPaeswOFP8zgyVB6Q2R4hBaX41Sae2xM1ceEB5WDD/+W/rXHTOTU7PJKnyGNrXBtp25N
GWaf3ywjZ2slFd1t/c8Zj5GMbsWgh3Z1q96vwnX2rMx6F6T5bFk5odur95d9JEOKkJ18amLjUZUV
pPCZvp/S1D0+Br/j/FVNOdSdZFDqx17JwbFDhWr0UdDQ56LcXdsNalskAFco57rzY7YD5e1oLAL3
c2ac9pgmzj42Ip+aV3BPjk4eocmSCFu3oDKmN30fiheZ/Yghmkv8uIBRIo6mX15j+3qEnS/yK94+
ey8aN2NZHKQgY0+pF802oLIpH+vh1dzhbLqfXkJkUb2NsDeJ8OO0uiy6juDZ8RfZRY4jwEk9LRs+
+aQuZqZT0a9XbMYUr8xuGIYrGgnecKIh5Nz5kBjGvUJaTvJgUU5GcVpMA9A09geRSv0VVKzXi5qT
V7AbmQvcpfck0HDYv2qLWK9bb2P9bXgqjxMTti0uKVz2Twv4+1bxvD+NTIQLL9Rx82GzHihjU9wu
cTAKdW9z4LgTuMrIjYSxAHdQvwr3ltJ+EkqtcoDMT0mWlgOxDf0Jjk6aiZdMMqmaBU1sC8BgmijW
1JTbCyei+/D08AktTC7bXcOtwCSQWHosdsNSvIvc3PZYLZyoxpGe/+aRp8dObagUuv6I55KLF36n
5JZiI2pducY1LaHCE7kEvQC+701WNYs2nrEzIY2E54OUGnCFSjZboQQFy5beAle2RupMSfMdAy+D
OvMd24e2D64RVtfPxUVniRM+KrrfaewsQT2BxqDPjnUTlPjh3u/kpjC28kqAP1IJCVM/twGR7Gw/
DMFoGRmxog0QjQDGfa8td8bh5rockjfDmcJ/p264+pcJC44gSxB+Ognm3WD50mahdaJnnSZGiSXU
YHhN/eP6irzwynL/nagznvBZB6Kjuz9F8xDi9XqV6kCvZeJREtBJXMpUyi5d9DfNppOtDvTQZgpW
vtjH8PH5J2n/DzwRiVXOCoTzZDIkkkt2L1evdMi7dcMqw3nTWtb64hnxg6fJ7CLgHPYFd1RlE5dF
RaFfmUJ83qFWXHIrS5t0QrAYwh4t6pVaNUGbCj/4wtE9o/F+8CwdpxmgxSvBOVCD9dUSX7pTFq91
XthOaV5qCW5ApYx6y/Teto35rHCgNy5KT3gKM97NixpPSKHzr8aJ0jmo6wY0RNMCFrpjWKZrSvSH
8Y8uypLwys81GeMGVHhnW3YtQpWglBzLmubvIGHBecih/3SFIJiUeWfNLL6SMKBkpH5cEsPr0QVN
j982r6pB8PVCjdxG81kTsQq15LCKIrsxmRu07DFMdHSmnZEc5fAXS4wIcf4IJbygLyIH5Kt3m6J4
SMIFKOjkUih7Ig2S0iDKRdZiTDl08BUnOVOyDEhWGfy6QDQZLZNUlvXfIEY8OpKHWWSLAL8hT31R
u2TOLwSSsIfnNNSJqA==
`protect end_protected
