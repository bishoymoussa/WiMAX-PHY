��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$Rx�y�<��wA�*;�x���@�̦�W�X�fa�M-$u����n~�%���P�$��W��kYَ���P7�?UMfT��q�6�U��k�>����~�\N�(�����X�e���/6U|)�X2pF�]$h���d.���9E��WG��L�X"]�Ad����ľS���8od����e�GT?y	7�������ݵ�^��R�q^]�鍦�����s�ae���h��L��P_���ާ��YЭF���'\��68�b�[����w8�[X��V�F�0͘3����q諵�uW� �h�u\V�?@��_6G�_�*�G���B�絉�f������[�G��U&�����~�F��AׯK1�`c��[<��FY���4I� �#�G��x[X�=�Q1��`��R>(�w����R�O�?����7�,(�H\�#h(W�EH=�������yq��Ѿ��aF����:�U~m<|��.��0=�P/���4ǆ���T(������v��!��Ϫ��71n��������.���Z�x<0�G
_���`��?^j)���gZ���	#����!�bJpq"�j��T�҅&�t�,�W&ѷFץ_\��@�~���j[	#�i�Q�t���,��i�m��D��]�_��i�9ިh"�5��v�%g�:�6���"(�lȎ�A��!�De�!z���K�n��1K��T�R�غ���*���C�T�BO��$��6���UA�+¬D��*�?�Tny'L�j�:�i����s6���o:�(�[���X� ��%g�ڢR�ỵv�i�^���B�B����u,��>t/��
�lO�g֥�=-Kw�-���T�F<�s!WO�E=�X��Q�`px����o���%�4O��>H��!�3)�JZr�;�)hyn��DM�.k����o.Զ��vJd����
���xɹ;�*vX���ʯٕh]���t��#����P,'4U,��A�[�3��J/���̂�$���o�A4;f���ʹ�l����1C��N�/�� T��tX�g3_5��(i±�J����\	Ug��e�+7��^4!�1�bG%����
�������S�Ng���6���'׬���g'2V,'���J�l֗s)�5�Ȑ��}!��{�'\����Uw|��|�
lF1��VaX����9�H�(A�����m��=���t�$�7�Ĕ�W��%�z�I��N�Z�z��YQ:��t7�����^�ծͧ�ژ�aN{�zR�4.ڇ�6\���뷂��`������6�@��?T�I�6������A
7V솥y8�����Ǚ?w5�Ӡ�۽ޞY1�TjM����RT�®}+�ɼ*�5qE�w��C�62؊kKx���rS2�Zn�|�)�F�o�5LMd*9���eR��*~۴��>;���l��"��2���⮠��%'�;�-�[3�`�'�X�v���Q��lGQ�ȃ� k����~�	 #D5�Ǧ�/�֜GD	�_o�ii�K�3�k��J����A�O��$�嘇 *��NS�W�	�ϵ��*����u�&xL�,���D��w�7���~VTe��� ��ie��l7�G0ړAW{��Q8
���a6����zl�IX��I
�����0p	꾢��I���ߚ��.6d��!���X�@�hҗ��x.,��W�@?����*8&f�o�O�7i�Jp��c6�+��%�������eS��[�~�I���MZ\l�%��py�C�<�|;Ѱ�)	� <��(��d�M�8�c�L5�j�����[M�2��p��n�� ��[S ":ΟZ߇��ٺ��i���HOa>@��=���3�+ od¸c���B!�&B9�H� �H,��w�z��5Ay��C��F�&/�&���䤬	tw�t����@�T5��g�����YҴa��j q���g~^��,�ݼ��9��P�99XѰ�j�ԣy0*��,�����IXq�z�uf1�x�F�y,���i+3Q�l��01�0I�".eZ��8�,�N���Tʵ��R@0\����|ߜ�z�Qu\��%v��������O}�K�)X}���u|ƶ߲FńI��������/���A��~Ug�.I3��UT�ᬺޫ-ǳ5F�x["�x؝���/̜�L9d�8>0��4|:��F�B:_�j)\C�ǈsLk�S���2��}4�^wD�ڸ��:�:�9"��q6��n9jؿKl((b�x	�"���C�˩������ [�3�,|s%�a��g�e&�o�/K%���lHR�6eT[kI);�')J�Sf���ڲP8�9���`Nr3nDD!`Ѕw��a�Ϛ��k"	i�h�rJdh�Ly���BI�]$���Rm�X��e&1	k��טQK��cw8�Z�Y����L�=����pz��J�jW�������mk��.;����0q\a��*����F�4���S̽�,�d�D��l���v��K�؀�i�^9�Q*����.�
�o��VB.LX�\�	V7X�|��ú����ur6)���x�)\��%�Qu� ���s��<u��%��2�f�M0r���0M���b���ih�T�M��7�ܨ�3�ǘI�aO��*��Q�E���j�|�9B�?m��A�`ׅ�R1���1톢�1*V�����x3��5���s��Q��v�>C��`�9���2�p<�l����cee�ȸ��)	
�j�~MA�
9U۵�8���f�t��U# �'J?i����/3o�v��b# dI>p� �m]~��h�tU~ֽɚާ(�sg�_<xZ�r���q��A�o��g&�џ��������5."�񷪀Z�Ny�-�7)���6��,'���<�H��ƗԚҼ�)�WZ��󣇙
��Q�d,���P���`�[��A{�=;J��zmdն[pea��Q:| ��t�uŀfb�C�*��z�;�	@��ۅ �����MsY���Usfg��-�'����m�� �^ ���#� p��"�c�}d
��{�K������V}�?k�#b�̶G<�u��}A8q�DAԶ� �[�¯�a�T��,[����B|�1U�q����Ty�#V��h|�1;�~�ak��r9$e��Ɉ_���_���Ǎ�ʎ]n7�����%j�'-3��``�����	~�٭�R���G��@O_q�TV�ST�B%Ղ���B����S�;�uE�����R�}��	J�S8���Y��v@<N$���w~�?�?xYg��Ag�a���ʣ�����W���64ck���'�>⡤T9�S�+~"����X{݊Gĵ"foMGFv,�!�A1�³������e��X�[��T~�ƈ��>ì:�`��&�A�"щa{�J��w5鷖��]М�Z�h�*g�r��)��8T�DCmg](��)^luT�CO�M���"+ʿ?�
w�4M	S�Z����4��ur>ku,-B���H�u{���E��&L��7qkD��}#^�!�� ��j���
2ȯ�9��<.��6v�x-S�i5;Ӝ���!?�Y7�f��dsKm�V��(3�g��
ϕU����,	����X�Y��0����K�/��j�z�4����+r���)�w'���h��oG<�~��k�B������������|���ě��ux;K��([{o�j�3���,�B��Dq���_v˂�P��/~Y�7����B�dE2��t�4g(z�T槻�Vm�Cc�l�4K�d�9��cwi�&�O`�a)��.����оC�hB?&�%�_Fq����;�'64B��U"t�.��/��R�!�W�|~iBo��9�gbGi�ޢ�@<��Ϫ	c�1a�%x�Ax�����?�.:���J�(�W"{�­�qE�hD�X@g2Y�N%Ɲ��s��;��zC$=2k@팥r�W�:IO��]�zw[�%��uԳ=tgY�oMj�Xt��w�p�}�n���M��M�ċ`�2w�Z5��d�X����*:�4��⛛�ٕ�`�ĭ!�*�58�b,�5��u_�6De���y�
0��0�Yz���{B�*!Q�wG�§zC}�56�
[�*�g�!�0����{e⯞�Z&�x[�5�qR_�"5(R���Vy;�>Ո��1Pڿ�}����bڎ(	��ބ��}�|�e�ӹ"��y�GPz$���P�G�^J�YS5��;�C��x����F��{��x�׵���Q�K�ܞ�;Ju�~���7��qc�Qb0<&s�;S��'���@}k�_n����C6��&]���e^�t��$��{z-���ߴ��sF>Yy��}0��4��,tx�X7D�/�x��^����終!l�����0U�FU%-�ѝoэ��{:��3yŔH|��2&�m�Y�Y>��� ���mt�����8�T�'+��H�x�R��BЭ�;��/F
��b�'��,oS󼢘�a�R���e"��Q�Z�G�=��V��u,����(ӻk�6�.~!۬?���c��l��E�-��.-��&$^�C��=� _-9�ֹ$9WZ����-����$��R�e�v;a5��r��>_�#��ߩ�?!C��ȣ6�0z�_�MP�+��ka����_ߋ�W3��{z��?���`�E���}̩b��1���{�5�(����B��;Bhs^c���C/>2�ZB�ҷb�)Ҽ�٠�6G��@[�@����.�1��LQ�4�9'���D2� ��w�)�� $�X�r�+�:H`X<W��c o;)7H{ތ���Þi(�z��x���W��@�PF�O̝�/�3]��L�'�i�`�\��F;N���-���2�yz5� oҘwk�(-�����~�ua��v{v#���$�{ #o:[l>3����y)h_��ŀH����2�s��S#�h�&hW��>f�8�T�-�=�@ϻ�w�@b���~\Q�������Z��R�ב���9p~`H��8��5���~7��*��e���e�f����t�l#��Rٷ��/G��|��v�<�h
�)F�����9̛><��M�	���u:���`�V"L�	�˾�,�ʹ���"�56�c'tc��\VV�[��+z`2/{�����݀w��{��ф�ۇ�