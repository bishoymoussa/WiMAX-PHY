��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$Rx�y�<�f��p��}Ԇ��c�Ͷ�Vϛ�6L��q��9fNDjG��E���L���5�\Kk����(7�������y����f7E�Z9^LZ�'��X�E�h���mD�Jر�7'J� �u��u��B��A�^�Ԙ��V1V�-�G��Ɲ�z�������<���Q���/ ����������,�������'��H��ޱ��vՐ
����[�Xs�O�.ݬ�%\�AVf|s:l������e|E���	 ��#�o�a�
I�0�i?w� %��F��������+$OC������&�f�I;���"'�,b��H吖����F�M�籠��`#D�@7Su�Z���S1��kb#tD�쪔ᅠV��� mʧc�+ء�h�]"N����͉���^h��>�%H�9�b�!ӻ/|���3V�F���k�-e��m�>�вڼ�Y� �䖞��f�&21��TS)�ǜ�X�!~�l����ypWiz/�(%'0N�Q%�!+v���B�ج�Q K���qg-;�I��>xA	��Z^�승6��@#�%�x�l���F�W�&���1i&1r�	�t<������[f�\��t����M��tC)|R��E���6c����A�D�J&⿚��Fs��=��L�9;��A���nfR�d=��R��';���Rs+i�k�e\U����XW嘑�'r����y+c�ݗ��"��`�����{i��6t7VEO���v��%tQ���w�3j�Bh�}�q���^z�ţ��|�e�V8���(?�^�Z��:Fv�C;Vr��r��Y�
��c�����(�зdh5 J��2T�bˇN��W�	��ɥ�wj��l�g�Le�a�^(O�\��R6���b�p(�l��M�.�A��;C�:��y�E�
��[�9���^��h�fr RhB�����#YYN�a:���Հ.�
��s,�\�@�?bT���R;��XAkk�V�M����=�0�)>ʐ�S��6A��F1k��uz��{���8"�e��~�����x��#��l�$�)���l�j�Z����\.&Pl~k���ғ���5�T��Z��f Zݔa�1t�>�q��GR���+;s��� �<���0hl��J�h7W 4�:��<5��$�����{[Ւ�;^�j�\�s�\b�~A��GY��a�]�f���ܙ��ZH�m��5����f�Z!�&R�eg)tn�K�h�=�d��*�9����d�1�j��q��V�S��d0���C
\�������M������%2���3��:�N"�%ӔX�׀���)�"1�}�E:N��S���c�xF��.]�!�/�d�J@=nz�.|��uA�%8E�)㈎jY|}Xc���w�0�������W��\�t}�o�қJy�ߟa<m/�*1�?��M=q*)��(
U���u������q�'4���j�Q(�����#�����P��J��B'y1/���]��o��H��d[��\����-gz�\�[|�G���
M��o��@�&у�K��Kڅ�����n� ׮ƨQo�I�(��r���Ɣo��yh���h5��^�[�ϖ�c�Y���r}ը��rd�"�!W���iݝ��S���Y��Zɯ՝Ƶ�ʆ0�ٴM
p%��Dp��e֤�YV��U��kTK�D��[�tkh/j]2<[��1�A�����9�xsqB���_�y�N�^j��`/����/�.Wy	GX�jvFt�6Z����p��ډf�W:[\G���c/}�}�۸��Q]�$s��1-�1���� �ǖz�sEJtO)!��G�e�R� �.��5�*B�0 �U�4��*�|�(8,I�2Ͻ��.���V_��ÅQ�1eR����9����]�]x�o)�ݿ��wwu ӷHt����Z��\*��Ds/��!�j�� ��S�S���g��z����N�H��"ܟs��`���vI��r��=�Rf��a�6G��/r&kJ.OG�D��/;�f�aӟ���Q7�1&["�pA��|-�h�K.+�Bs�!k�ǅ�����լ�Zà+&`zI��b��&����9o9����DmP��㕶[(#_@:���S�k/O�����Pe0���$%��#�NU�	Y,�U���C�����k�{hs՞pI���h�Ć~�8/�WG�y@$�zǳ˒g"70|��.���\B6)���²R�ը���{�e@f�����9�׬�H|��v����g���3!0H��6�#�I�0���]�
m�U�57޾ �A�@ 0|V	~c�B��[��h��6��Łf$QJ��B����c���8��U"�{�f��.�^�n��T+W[�k߾����Y/i�徐�����db���X+�I��g ��L�g�ѭJc��ρ?��1J����՛C���N1��n�$�r����6,?��ж�C��&bq/���%�O-��u�٤z* �
AE!E���7��^����gv/Taވ�B�Q��f.[���Ef����z�����.�Z��~��U���m���վy�iݷ���s�=���j��I*m������B���J�|4�M���RJ�:�<�����{�c�����nAnw�ܨm�W�{�G��Y�	c�G'����F�X�.��N�sVI>�� �)��p�7�!��0���k�aT˭���3VC�5�2��K�#�=	��Z�Ɇ�8�Q�L	zs������{m�Zj�E��i���3I ���c����b�B�υq�ҷ����h��6����G�x8y(m��C�*�)�4��2�Egٟ�C�u����'=x���R�snB� ���
̧I��}=�3�{Y��W(�Q_���O�׼�g�.�hBBɵ('tޝ�i&�����G��̵�t�v�������C-	���V-1��XGtU�"�O�w�٩��F�^	8�7Ȗ�������4�K��|WH2磉�<wN����fJO=>��\U��Q�*�\/�:z��,���4S8�V�Bb�@�}�l��{<��Dn��t\_�C V
�2�Т0]�K�a�ƭB�)�H��P6_AF�#iz]ٽl��奲�Y��f}�InQs����x��Ź��ѻ?���
-e"�'9��_�0�.�Y�x�g�p�wC�8%dH��Q?��昢.�^�$�C�|Q�[���.K� �e��\8Fe��&:�+��Ɓ<;����S��/�!�\ r;�螤dm��3�t�٥��ofM�y�_Ò&ݟ	}$"�Z
˿�e��ڐ��Y�{��ܘ.-��mQ�zr@�����±}�)̓��?u�5j�>Q�7@�܉��%�������*+�=��By|
���2��vK�{��^��P���k�v4��9�;����+٘q�M��������7Y�����Yi��3H<W��+�4{`(@ٗ}_�����Wp����W�'�q6������6p����$u�3<f�*�<ʙ�E��?����� ���~3��(���^rTy�`p���d���6��NcF�9�륟n�Ä]mD��w}����ē��T*���k�_]���حTo��Π��VI��:Đ0�k0��-sxKG.�yͳȳ�D���Ei)���Nv2]}U������i�{|��4�x�Ө��C��k�C	�V���[3&�;� �{�K◨�=����2�-%�?�%�}c)V����i����,���}(�GPjFQ�Q=s�mCN~^���iC���P�i�gBMt�	`Z�XB4�At�3m�����V���Ug��	S�_CwH�W��=���&,̤�D��@��*X�-���ް���y�<�eɄԛ��v�S��'�F�-��C��-��ʮ��O  ��5Z�%29{Z����]I���؉�q�G�XN��!п7fG�-��r��ą0��jG[a�BS����l�]r�~_'>��8� =�_;� =�I8�_�Q�JQP�I�k�Gd8_�T+�Xg�����ο#�����`�Ֆ����#I�6����|̑c��Ƿ%q��	+�2�2�5Z0�V���iQ� �����-�����T���ьy�b)�M4��v�o���k�o�e5{4��+ֶd�ʰJ�e�L��s|�d����j��v