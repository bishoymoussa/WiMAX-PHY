��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$Rx�y�<��wA�*;�x���@�̦�W�X�fa�M-$u����n~�%���P�$��W��kYَ���P7�?UMfT��q�6�U��k�>����~�\N�(�����X�e���/6U|)�X2pF�]$h���d.���9E��WG��L�X"]�Ad����ľS���8od����e�GT?y	7�������ݵ�^��R�q^]�鍦�����s�ae���h��L��P_���ާ��YЭF���'\��68�b�[����w8�[X��V�F�0͘3����q諵�uW� �h�u\V�?@��_6G�_�*�G���B�絉�f������[�G��U&�����~�F��AׯK1�`c��[<��FY���4I� �#�G��x[X�=�Q1��`��R>(�w����R�O�?����7�,(�H\�#h(W�EH=�������yq��Ѿ��aF����:�U~m<|��.��0=�P/���4ǆ���T(������v��t}*���I�6���|sL��� o����jP�Xfۚ��u��5 ��<sKa%Mx������_�z�Ì{V�P�����@$W)�}>�^�1�7��-k��[�����p/�z�R9x��|+% ����b�.p�X	E!Wo�|rF����7f�$���[��2��L�U���U"ճ�����w��:[��Ӈ��H��Az,O��"Jbqkn!1J� ]�?ѓ1�"��}��qP5BD\g��6��#a�b�x�������x�K�{.�OF��a���s_���^�8�㲓�⍣:�k���y��Loy�w��-d���:���������(e�[�C�$c��h��G΂zȡLD	���lV��mrbp]|�t\�y���+��9�ݜ~ �JՈA��&������>�
m��~�Oo�r5��j'5�rY�\�������������~̠��ƪ��������6DI����p�V�+	��`}~��9���R�������}Qw$=���e��ok}�xћPzǤ��Z���7C�m����-"���,G5���*9,�?U���]���Ck}]�b�$�F6���h���0m�Agx�}�FG=と�����?m������`/�B�ƃf4љ���}u�^W��{�]T�$}�'��V�ӽJv���Q�'!I/�0��~�`�`+DlD4]�� �c���.q���b��ǧ0�޵H�,g*��Ͽ��y�Q�_,d��i��Z�2��3�+��Xa
������
rOX�[/����Z�G ٻ �K�g�f����]g8���d>|߹!,~b\iۡ�l)�}�+P��	.�A� ��?��e��X�K~�ug����1ʃ�I�����<KT��E��0j�1�f�������I��'�K�(g��2��!ǜ��j�u��V[B�k¢?q���4��? �k��l���S�K���p0P@J�@�	JF�c��ߙf���1�Hvl��J�s�eM4��w\�/�����R8��s ��7� *G��$n�ʊ��~�����H�5��d��[v��v"���;Roܿ�̼,��9�4JD=ib�`'8�6������y/z̖���/�����gP#:A،ki���|�A�ɻ�A,�ó>�Ѷ�v�5pF�؋[DV�� {���lF�E�����v�ҳ�z5a��`�!��s+:����5���;u�Շ�`��T�ЀF4�;!=�m?�IuV�`B�;"�!���W(.r�����d��ݕ�2��"�2qϻ����3�ʗ�rruJ.Шx�̜��������~��	�LM{���:Zl��0�����J��twO� ��fa��2oύ��}�$�S��|X��`{p4gt�+���r�8�̆�>�s���'R��ɬ%۪y���*؊8:tuo���.PH����RGUh��y� 94@oc����:5��e'�*2^{�"�8R���������7�NxM���Gt5�l$FA�=^ ,X���]�Q�n�{�yt�$�_��yU�d& �JW���4U� |�E����d7��$��Ż�R'�Ī�_�� �&5Rm�������<��B��l��Y>~dƉ����p����mH�U�&B+���k�-�Zd�����*����������#�k�|�� @(9���F�/��x�G`+�f2�7ђ��4�8�) M�/@t��E$�Xd��A	��&��=Cç��_��� F��ADFTE� Բ����Hc������ ��'�g�V�	����c�h�:��.0��D��*j'�t��<�Z�>K__�^�-�o��k���&&�:ר�{$��Q(���x��P��﯎��8�>�����2��������*��l��qp`oN&;��~:t���ı!���d6�DT�>�Cʄ�C���^�#T�5�ʘb\��n����t5�Q�2�5���w/Ʊ]Sߵ�i��LbXp/F�5�����Qx]&��*"t�C�4�U~�I�y�qT ӿB���zn
�f"x�@\%L��'���͠w���a.__ƴ��E-�7�*8rr^�\H��]���Ȯ�`�j��H��{=@k��f���ѦL�=�������PO�� _^�	LD]�/q��$���UI[w�!�qU�m���~�U?����g�����9?'�\��-�-����Фa^�7e�gK�-P�$��3Y�٬܆5ȉO����Sκw@���uG�����,*���������t]���hP���A�|l�+�j=����	�+2��7�o���h�Z�ppſԡ��fl�Ә������T=C���d���@s(o����3��dx��TT��� �i�jĨ�t���B<����=��щ1U`l�1����r(�T�Ϳ Zކ&���!�Brs�|�x��E<z^�l۰r����i�7Ct�;B0��q��O%�:J�V�o���X�[�,�4h§�v�馛Ąe/�D�(�7^���)��.���g�M��B���[6�b�g�N�,��9D���:�eD̳oy���mY�lI8�k	W���bv�ኤ>�<����N��3'Ehg�^�,kى%{r����[��9�,�N�Pq-��"��璬u��`�u���y�5�ߚ�] !�s�:�mE`�����~ugY �Db�����S�Ƒ3,��=���sG��:�+�r�H}sg$����Ņ�a�v��Hp�X�%�R+s��^V@�ko4k��#'�&���{d��ҹ� ��0ZK�(`eiU��8���A�	~�����~(����XHu>Z�����$��雩�������R�?d-�B�&���n}m�����A�� �~��EκK8����ul�cH���<x��ǃ���M�?	wF�齃J^K�~8��gU�hyiz,�)�L�Q@%��Si�<�ȴ�b�h���k�'T�����	J���������R�ECv
��qf ��Lv�D�o�<Ƒc!h<o��G?�����}"�'qt�N|t�&�m����fiG���5� �>m�E?��&m���6	���m���i��Z*`�+��{~�)�ѭ�'T9�����S3=bd�۵c5N�N8������-�p�i�k�
��7�[^���>}u0�vz�{1G`�OX�25����p��o�"C�����Z���
|�'�֑�;��+�3Dp�?%UZ[
=j
�X�zI?��0ܵ�j]�,�l�SJ��O��}SN�ی�b�O�4#�5C���̷՞ߐb&�c/��da/��ת��,��gm!�":��>��'���i#��.2%J�s�wK�sה��{�jׂ-h+����L�Җ���fi����dN��q.�����S:oo�m�>A����Q^!�A����jC��D[D�F��܅����Y:'[ÁA�;� �@�݇�����P%ŗ�����=߼��r�����.�*��v\�j:g�3ylm���3�����xZ-LA�h��aߩBM��օ�2��/z������8�g,�n<lHҜ}8��#�h�YA0��I�Ű�c�"u]�C$�M��~�^|x0�{r'�u�`���vB�br�;$�͏��k�b�nU,;4$u��w��S5�r���������+pϭHq����q�71��$ΫӸ+!� �7'~J����BJ%���C�Ά����IS�ȷЙv	�5�L�vN�w^B-˔Tc�]�^��"tF�$!�t$��AU���k� ��W3��̏[Ә.�߳:�1a�SD7b�qGo����5s�cU��͋E6�k�x�����&�6��7i@5���o��j`/����"��T߼"�Q4wj�"G0m� �>°�@�-؏��.�E޼�_��Q�n�=7ނ�gs��G�����t:�f�HGx�3b�G��:am%g55��,�}I��Vù��^!*���҅�gR��<�>��o��t��рk6S[n�_����[�^�����v��-X6 �2ƕ55`ۆ��AJ��F����U�*z���!�>��C���3Sul�~���AY#9P�@_0��c�̧.����ٞ]��R�s�E������i1'����������>�I�)�3���c�M�*�@��_6�����\��'�Ĥ��^�����e+��#~�sh��-�
Z:�ۗq�?[��/�J�JhJ4��1J�׿:oi0���巴�&7o�)՛��y!�����C��liLX'dL����7
F�9��?��NKr�}�̿��������A\J^U������L�8�|+H%=����;�֌�k<������I�W�*��d�&)��S�$��4,�=����;�j��%��R/ov�l��5 ���bX�����W��e����Y2un}�	t".�_w߿��,+b��T�Õf<�籼Hb4��?HLvk�B;/��m{���x�����{��q4�M@!��$��N������Ing̘�%���-|_*�fp����	3ӏ��( �&t3���bdȥPQg$e�sX�3>�a�5vh-�]���T,��ϊ�-�Tޏr�՗�z^����l�_ԇ4��z1e���]	Qh�ۓ:`[m֟BY:��Č������͒fc�-�
��P�*��!x��n��E��vs�t#���Bn�|��q�C��8��g2s�q����woo�w%CX�(C�zo����M4fLI��<ۅ��b��I'�ŵ ��^J�����W<U�B�z0��K�|��	�ĕ�٥cߚ�}��Y��A} S�\��+���I%1)����e�L�Xt�� Wڼ���8;�5�:����uS��q��;/�yh)�^��@>��R:��w0�J&�}�Rk���Yiy�\��-�U��[dN��-�2�>����oxSi�?�6-��Bl$�V^�T�B�qOA�tM��y^2�]������U���5��#�Q<d?�x�˼�5<ҽp"/�W+��^�>�z����v�����N����O�D�A����a�Y�<Vi�=�]^@������ojo^�Lg<r�ƃ�:�x�.�;b�"9w^�/�ҧl��>��B*�dt��	LƷG-x�xp[��+��};��J������8��T�v]���s�.���8�s�_���X�e�f��^�Wк&��=��j:H&�Jݭ]�~��Ȓ��'�����J�LK��\���
�U��zJ�a �9�]\`�c:e�\)��L=2:�oc/��)�Go�I? ������Ї����vS?�(�ه���z����ר"E���4]�D�k�Fc�=��.GW�BJ��a���`�͹�T�&�vIWT��w��G�G���oNg$*�9?(�y@0�^�-����х8�vS8C0��U����T*~(��貵��TD�[������\�z�Yr��h�Ą��x�hd).w��k)!j��[��W�F�ө�ވ2Qic�F���K��H�w`���eOO�k^�^�O\��*~��;��l�+؎�ױ'�������q����@�Ю2���1���lۨOP#/�`�C"\X��ߔ1�jS����+��MV�~�7E�-���� �9����L,�x�U�$�A+}D.(t�r�����	��u>������w�5Gn�����
(o���4����m�*�0�`E�O��_7��EN\̛�8;��#:zZa�s��i��!�c]Jό��eh�F�<�A��k��D��2T��P� �vwf�T�`�r�d7�?�����7���]��[��� 2H���%A�fl�*�^;>� m�:C�o��R��k�^/~5޹�+���1�W���s��V)�l�˒�}�G�X�o���Z�y�V�2@�#�"���B,���C��,�����Q��̛)���w��Qs��r�>��1R���R����X���[����B*4Ř~�����A7�"$��'�|�{���K���^Mc�lɆ^G�(q���2��ޫ�v@�D]b�qq���}D�CU�z�\̶�?S?��j΂kx�|�;.w'B$�qB���'��PN��<i_7��/��Fz�ܬ�W�����@��s�lLp��<�&��;����a���������(k�B.KU+c}O����bQ�31B7Ǽ)2~2�������ܢ�
���[�Z�A���g�H�4�
��ڇ=��I��a�Aa�tƕ�!$��[��6ޢ27��2�.}۹c�c�X�\S��ҍ�;]'���UMpi�C��ڴ�X��3[#�� �lA����e�M��B��%�����fͨ�&�F9u��3u�� ��\ᳫ��� �@y}dj+�a㣎'q�i�ʛ����	�&N+b���,�RD�"^u.�$�i�n
U�����I J��L��z-��l�@9dw%�xb�,
.�q��� c�}ug����z��ߒ*Y��p��� ~� ��eZ�&y�F����{�z����r�^t�N�9���蛸��ԻJ�p�X^����]�n5P\���AN����$5ʵ�[z��F6E)�0�vC#���R��*M�Z;,�g6Ԍ����+3T����mj_���yuz+We���γ��<���~L'�g��S���