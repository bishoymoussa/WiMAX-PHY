��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$Rx�y�<��wA�*;�x���@�̦�W�X�fa�M-$u����n~�%���P�$��W��kYَ���P7�?UMfT��q�6�U��k�>����~�\N�(�����X�e���/6U|)�X2pF�]$h���d.���9E��WG��L�X"]�Ad����ľS���8od����e�GT?y	7�������ݵ�^��R�q^]�鍦�����s�ae���h��L��P_���ާ��YЭF���'\��68�b�[����w8�[X��V�F�0͘3����q諵�uW� �h�u\V�?@��_6G�_�*�G���B�絉�f������[�G��U&�����~�F��AׯK1�`c��[<��FY���4I� �#�G��x[X�=�Q1��`��R>(�w����R�O�?����7�,(�H\�#h(W�EH=�������yq��Ѿ��aF����:�U~m<|��.��0=�P/���4ǆ���T(���=?�D��D��Z�W]K�[�+ӊ�W�9w�S۩�[�nf�"%���7RV�e���q�gd"'�B��Qң����z����q'��(a��Q���MZ���R����s�)�>�c��*hE�3t��j�(�홻�W�t�����V��- ���;S;#/�o��8���L/�;xX� �g�Ro���T3���e�i�Nq����I���?��o<��K��o �1��yd��/�� �&YV��kJ�2%�{�|��+��}[���D�>�S�ŭ�<¼M��슭��O���W�3EchV������yh&�_����ӥ��~>�<_�����+�C,TA���	��1T�+y��~~��k u�E,�+����qro��NW;R^2���a(�8�줔@�������2����y*�c�0���j�{�)P�g9un.7�D?�.5��!��^�Jne���_��n=�5�`��i_�"�8icf�@uv*�ܟ�B@�7�S�*����L5��ϐm[�pp?|�b��3@=��9�n����-Q����r�Y��3w��R�`6:���.h����{"F���{�(_v��Ϸ�C�D�e�!D{�ш��/��a�w)�ɏ�s=�XyWC �ȩ�����El����ӐR$�J��k�x.3���~f��bc����h�گ�Fm^9��k���_7Q�Dͯ""WU�h�Ĭc��d���W���j\�Kڣ2�aN	 G���̴A?���+X��o���|�_�(!�}�?o����ypR�M�_�?	#}�����]}˩�5� ��]�����Z����YY�Z��ó7��N�O@i�Xݨ�&hE7 ů4�Փ��6�|}�i��u)��HU,*�98!�kǒ�!�
�^�6bs�Kd��F�'F\�ͬ�=��=9S%��r�i�Kp(AF�lH�o�.�'w��P,*/4��Ķ�#��`<��/@��g����� 2��g1n�8��w*�~��6��N�S[}�xd6�:���<��A/>7s�ti���Jo�
�����ݿ(�3��#�O0����F=(���w@̺�����64��Iu%��[�R�dpGA�a�!�
kk���c:��`�����}���P�Ha��� Md���/T��������Q��Ln~1����#yz��X�?���5���R;��1��Ӥ_��ڎ�2��ˬ��ye|�O��⦙2*4Ԩm����(�