��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$Rx�y�<��wA�*;�x���@�̦�W�X�fa�M-$u����n~�%���P�$��W��kYَ���P7�?UMfT��q�6�U��k�>����~�\N�(�����X�e���/6U|)�X2pF�]$h���d.���9E��WG��L�X"]�Ad����ľS���8od����e�GT?y	7�������ݵ�^��R�q^]�鍦�����s�ae���h��L��P_���ާ��YЭF���'\��68�b�[����w8�[X��V�F�0͘3����q諵�uW� �h�u\V�?@��_6G�_�*�G���B�絉�f������[�G��U&�����~�F��AׯK1�`c��[<��FY���4I� �#�G��x[X�=�Q1��`��R>(�w����R�O�?����7�,(�H\�#h(W�EH=�������yq��Ѿ��aF����:�U~m<|��.��0=�P/���4ǆ���T(���TK�@����3L�m��a@e�Q ��1��~�7z�����_$T��6�E����c�^�^Y��Ր\ߋD��KG�����,��wm-`g~�0����z�k��8�-����S�\��6�0A1GL����Y�޵�mA�qg�i����r%M>�sx%���l�.鼪k��/r+y��Y$��U���Ƹ�WW�л��_P��g�$3�W��vW��'��յS�R�)����:!��70�p�31��g-3���x+5ܧ~�&)j֘�S��f#_U���]�V�s��|��o��[�E)��Oc2i�'
�u���Q)�rIFʓu�o�,��s�!N]c����|�jLJ�A$�r~��#�V�%~�����H��Y.����bg�B� Yz�� �F��sG(a�O������xqr0�����wQ�}t��M������;��߉�p���!��rn�hz����i�����~e��v� �jhk��������CI��j��]F{=y�8��M�ufz����k���0{��2Z�"�r9VU��/!؛��r%P_������rH�sƿ�ByJ�m U��/0Ճ/��N���������x�.�}�8r������-��Z��q�:_�;#Qa�>'L�9_,f��8�Ԗ�q�Fbe�$~������-��iH��h��3�*��U�r��K
��XΧQ�]�|�)��i(mH���F�x^��ə�D
sؕEa���8'�/w�,��FOt��t��VJe*wgg"P%�wՇ�Āaf� ��D���:���DY5P�)�8;1��+�z��;}y1P���9�#Z���u�*��ֺ�� Q��Cls��4�jx��/0'����x�<1ͦ������SS��������B��D�1��I_��8eZ�J�����̦�\&�E��q�G~�v1��,�w�uFd�p�ҝy���-�*jZ?V��蛩f6ߪP�ͮ'Iq�6a3RxI���� ��?�4�f�%��Y4N����晻�6��t����K�/t�]��!�'�N�:��D�9�����{6��]al=α��kc; O8��.��E��K2����`US S��A|������#�]e*��{���]K����p����G<�)�.ӟ1"�M�e�@��j���^:�&M- 
-l0�dwn#�T�� �4c�=���p@3��lr���6�WǊ�w��7q��S��0j�`�>��s�!8�|�婨���Lⲯ����>Ǧ1p$����Nrb�������H��\���ӟ���t�(�'/Ρ��?������<�q�����⺡O&|�듲��Mcd9�[޵���@�n���s�a/�!��\(S�}�$�QXҝ�%y�8�F����v�u��uz?�q��8��&�x2K02oD�P�R���)HS�1tDK@+�4��&�Fegl>K��7�/�T�}:� �I����R�bpsk��i�R�[�Б�xUj%��\`r�����d�����]��tJn`KkO��J[VW�g�ѩm~�������6�~�n�4�md��w���i�6>1�`�^_�O�{���!�j��P�#�Th��;7�(O�8��t�͵����C޷uG꙾~�����Q��u�r�mФx��PwE)�M���5��X�ze�t�r�e����C�d�gYwib����e�2�<Zq���+YIp��~w�gs���p<����\��7�V�νA|�X��x6{�ܾ�z�\鉒�7�EU���?4�/�QM)�#�zW)D�6���O/���!T/iU�,�b��N9���N.n�e�fo�P��0%�݌�}6�Ƣ�9�S1����M���9	�<�~	���4u
Ja\����ǡo��z��8�R�G�{���n4�˄�]e�-���o�� ����d��Y2�yf]����.u�w�QCWE�-�p�&C��} �\_}?�����u���Й0?Ɂ`2�I��Q°�V�"�'6 �l墿�"���VdN�u[:(~�ڏ5�&(��z��ke�6n���y��"Ia�ܒxby�'j�A�A�t���z�RC����v ����0q:?N��<0�Z�룚�"cZȮ�8k�J���h�ct�,���gdGH��$,Q�4I5��a�����{���C���a�@[̪�W� 4e,]���������VP�0k�����i ~�3�bL����l��!��Q`g}��8p����ϯ�.N�ї��~A�_�89�/��!
�9�+%�5C�=�]̀!5�è�D�:�k����ںW����յ���������)�E�oq���4m˧�X`����c���3��W7�X��[�&y����o��3F�6����~s��ૐjis�V��|ZAY�m|�5���d��mO)������[�:�7f�h��% �1��9ۛ��O҅���3Tf�.Q�����aAV�4��}Ì��|e�~�;t_Әy���dZ�����[͞�Ր����E���x�J���aR�l�,��dFt���Y��<[��(�ZL�\b� Vl�ip��& b�f����j�3�t�sg������z ���:oF�7 φ&�l�c�Vv!�l��^eٮ����s�bZǀ��S.�C�|����4A6�C���q��}����D5���L��ѷ!`�h;/�EG�"�`��5勒�ԡ�OK�ߧ��L�[�pk_0�y�8�ra��`���~Un����#Y��U\JGtT̽�J�P�`���i�E4@&��e'jm�t��]�-�4;䢄9S���ٖS+�/El%��餉�w  !�l<0(���"�p�\�\��!��e�i�ΗH�]��|]��c�bzح�9�
�;�F�M�`1X�Z4zR}�-�E�~~St��iY����᚝�PX�2�~�;EJj������[Ea�C�(VD��a�`̂���\��2�p�8t��FU�V�Ss�:^�[ܑp��A��$�{5r��d�l�2v���Aş�w�̖�Y�$���ѣw6����M��|�:�0�	w���^{��`���U���D׃6�`N����r`Rj�W�y�j���AG��K��C�q��o�O�g�;�$�F�Ծ�Z���0T�G�S��As]��`�q�2�&���ښ�Ӕ��I
�����d�:�Q$���z�T��nB�" |��3�.�d�sdGJ^r�ix^`]�'L���4u��yĹ�1��ݐJ��DY��8�V�KJ����E(lh����D7fU��D�T�;���'�K42c.�Zΰo��h
�d���T���&��i���>�2p,�c׶��[��ۧ}�՛]�r��Ή	#ƈZ��j�۩����-�#tμ-'S�b8F���p���ݓ4X�~��Xg�ofH�K�����^���4��群o��v�e!��Z��L C0�쁞 �>a*l��g�m�T�&N�xG�M.���ChlL�Xc~@�B�*�G�d����.�0�wj!�����:�;7Ќ( �����c[A�?a�m�ZP?c���3�.������ja�4Ĝ���O6�3�(x�Ь�d:E�m�Y�d
w%f	I�l��=Z��W}}�M(�KJԼz��n/��C�"����pb��:T���c�֕F#��u����0-�����*v;ap5&�A/xu�A�<�8����G�'N�݊�u,�[�Y��d�(2�)e�xvwQ�=�u�]L�����y��%d?v�s�ꠎiӜ(8� �׺��$����W�U2j�[�#`4���Կ6J2�/��s�i�P�{�0 M���&�p���ǧ�,�L���r�FGv���djd��IwI"�D~�2U�N�Ļ���8��}���:��]߱������7=u�佯�@�s����0��W��5 4\C���VQ[�냴6f����W���ǿQbit([��_ce�h�J�$�Rp���8��Sه,����q7}x�s��š�n<I%�i�l�[VE�K���J5U쾮 @���5��(�ls�ы~��$�e�%���@�qݜ.#i�*�+ժ����b"��_�;$�%&X@Bm�}��]U�E� �,���l����
�)�Pg1�IwrA�)2�}���r�����H~�BC��N�1{7�-Q�V@\LN�cN���j��On���|�=��[4��������QR��}pX;Y϶l>A
�t������5��Z2�O��� A�P�$\\c��ю�1:xWqwCw8;L6D��o�]T���4aw=eKOoe*2xiB$~��FI���p�����?s�k<��J�������R�3�=��A'e��S�'!W��f&?�L�A
- Ғ|��hY�
w��]Yp�Q������������)0�D����L쮎�xq7@┦�QΥ��/���H�Ϝ��m�Ecn$ 1�#M���2~�/��V����0.�$�	c(�B���$P��C�������PG�U����s8s#�T��S�%�_�hS|)���C_���ν�/���K��!	�Q�qO��|O=�����1�^�uf���0&��ī[cw��zbD�!T�L��nE�Q	*Z��^�߱��%'�ߋ�{,�Њ��0�DJ�Рa��Ǯ ��ÿ�����c����"y�*�m�� �l'g� �J���Z/0#��?|���>$� ������nK�M��΍�1C��7|!I՗LBjh��٭+��/�!KK��q�s��3)�=>@
�������Ia���1��D��LQ�w�og׊������V�N�p~iD5�\[7c	�y)/���Bj�+ją�<3A#S�n�Z�Mk��6��6VJ��?����H�#`�~I:ѯ��������G_Zc
�Q6i���	�e
�pLc��l(�mJ�tD��5}�� �o�An���d
��?Az�d�,l�.ˤ��������2'�� �p8�/?j�q�D���b��_���������K07�1Ňd�.����\'��B���.��,Q]�k�g�w�����o�*{�����str��VØ�s���xg���2Lm$ ��(���� ����߅����(�?g���%��Ր��%���ש\tY��;���=�
�u�u)3�L4�W�����m�u�s�V�B�8ND'�3�	�R�j@��/@9�j�]ꀗ�5}uCj��������>��T+ �G���u+����T"��\���Aw����7NQp��z�7���Vr�]�|/��b��38��Ȧ��{�AyTe�j�/���C��d�S�	�CPj�4������0�hn�+��9;t�/��F��u�@�a\@�w�"�`r�|�1+�}�c�QOb��Д���: ���R<�|h�$r`6����u$,�ߏ~@.z>��s���%�RB�M�P'�#�As�||:��������AT���� ��O�n�8��'Ӥ���>t��o"L�6+�B��?~��A�(��b�`�1��B�.��30���H���J���Êv�!�^z�֧�]�u��fy:���������|�ye�v��1)E�S��(�Pn{;���{,�� �s�A�(��	��bt��F^�
7��L4d5(`&12�5:[]���o)$��_�n��3tT� ��[��$�yIB�L���">�W����1�8�уtå:�G���Wlړ�z�$�!�2��H���hC%��v׵hM�tu�E�"F�Xk+��aDUʦ��EY4 �����#���m�w�'i1�t5�%��@�ޏ�|����U�����e���?��:�f8�FD�j$?;��UB��8�ʕ���	��l�)<�T{l��sSSX@	ۣ%v��0�v��V��e��p��8 >���E=�}����v~ ��D�EM���� P�2]����1�ց��P�&$��P��"��d8��-�M`1B�R׽m0�:JJ�����3i�@���d�;m;-�:�-o^��hV�߾�� 	�ut�ș�z��Ei�_ߖX�-W0�O�]:^�fK�Q}3���b�@h�>ொN�6��՟�S��D�*`j۬��h��ә�
�'|?�kZ�"ZM�8x�nj�Y�M�~��P�ᄅ9�Z����)'�����ĥ� DzP�>+&�P&����x�ϨJ�J�?�:�r7�8J~��W��N��#�'����Ht���/{��p�4#��u#w��CNС�\���Gdg�4%QB��K>�5d��%�2Sw�����s��^`b7����Wp���+�=���O���z��a��^"^ppzp*�"�Is�9$}�ca]�=Zg$�p��9 ���w�zEu�H�խ�OП���z�D}8��`��x��<��y#��E�*j!��I[~[� ��Q�?ez�SQԵ�׏���w��$��w���q�T^ �4�̧�3"8��^�|�9[x�r��
�kR���n^6t{fWƯ-�c�A����s�1ay#��͢��zPrT��V�K�7G����(�;�j���e뭯��+}����3N����6�����w�1(dF��÷>@�F!;�amg�{�Z�U�Q��
qǛ��J�io.������	�XG��0��VB�v���ʋ�����6�;]��GO���XS�>��!�R��U�,)!�}�&~`�U��J�*����:���,vC�\u�3�Y&�,��1��K�#����0g�KD�����3����=�N�O�WJZ�n��x�C���c���p�M��"�Q�Tً3�/�s��% ��^�R�H�xa,���m�	�I�\q��f�x���9�<��+
JZ`#	���ӥo;��� }+��0i�$!�d�1v+����XL�ϦH\>�z��(62�F@�(Z�@q�\�~�[��F�|�4�;;Z�V��}
A��v	���%ရ�b�,��M*^�ђ��A��M�% �\�M������o%�?U�Z|��(��P�G|%�vE�w��#R���`h����ħ>��CJQ���!@/Hey[���� ���`0�oq�$�r�5v��f��~�fS�%�ݕ�,���Ƞ�J�TgX�>w�	ד�5�zf{�$~�-16�,I����!���C-��gM{t��R�R���o��=�Q+4��U]�x��oV)��'�,��+�;�/!���,.�,�j��	�N�v.�I�ctP��a� �F:����� )AĴ��~Ĳ���B��gׅ��׎B6���¯7"��V�搆�����axK[�Xo�s��1%���96"u��/R���'�ag��kt�Mӛ�_���I�_�CjS!�8��K���YvН�7�ati��b�|��>>�5U@2�3p�;$�]�V#���?'kJ<�zARA=h��NV�s�p������\���^'�z4�$����0��9�M�E���5�+���G�C��s�zfG��s�?I�l�x.tĤ�i�T*,P���S�wS�!����l�b��F�n�l���vov%(�A��dP��x��47��A�L�P��6�.�>�7�vq�L���a��2MO��B�bcb�y;u�} �A 5#��𲅒Q��`5�1E�s.�� �p���5� �n��>�f}v�)�:��T�N��e����m�5Tz:��D!f+�N_���
%Id"��������7�l�AO�S}K����w�ؙޥ�d�zO�^���Q���Bz{�t2�	U�4�G
���ݫ4Xh����ђoL�D�vgFN�ZM�w��<�MjJ���!0��nx,z�U�GƘ����XFO�B@�AV1V�o]s���eD���	�9@q�(�Ĩ� ��z7�(��K�j%$WKR�sb���ΔG�#>�W���Q[��-=�c�Y$�r:����h��q�Ͻ����%�����u#.)�7�Ԉ��;e�	q^�7����E�lr�n%�ƾ�[�fb,�3C�Y�Z�uE����'��ʧI��x���'�� �>�����;j���awAc�8P�eK/@�Q�[N�FaA-���#T�D+AdK]��́K�t'k	,]�7VV�/	�V�cL^hᨓc�.2h��� "�<�I�e[�%��1�\�_����ڸ����S|�{օ��&� !%�?�e��d,3��}�i��Ϫ��vZ^�ੴ�8�v��|��R#]�2�{��0Ǝ��%2 ��4�DC��D�r���zA;�UU����Ww檝�A���.�i�;$}cʤ��_��О	9���N���l�+;`hkB����^�A'����-�&ٗM½X~�352������3LD�$6�}�W��P(�d�k�.������B}�̍D`�6p��-��0��mB����ʌ[��IPfZ���z��I�:��=�ָ-�ܿ�����Rۀ�h ~��p0T����*t�o��V���D��9I�B�� 44�׳"(����+�2�~�ݥ؏w�xb^�Q��o���R�>vw���S�0�ҁ/ⱍ�;��kU�r֬iIs���ܺ�q�i�0��H�#�C���A*��R ���e�.��`x�;lVSp�4E*�a>�2�Kc%��y���E`־��������Wk�����\4���fR��<�Wn? zh��ș�AQ��h�� �E`�M54>P�W�h��&�4j)A ?�u���oF��i��/�r\�/��ӭcº� ���9A�i{t�>d+����!T(��Ț|V8,7����vu�5���3��j4� 0�4�f��?�YO��e�x��cP~�i0`-��ӿr�#�U�DQ��3^�qFfľ?�؄�燐�E�����$Z�4��%���t#��
t�鑃��HL��1�co��eݬ!ER�S���sQY,�vPޔ���Cm��:�H���f�P$���] iF��֢�(.�67�p鲞m�3����V�6'r?0,��/�C���:ciE_:� Ypd�5K@��n�`KD&4ܐ����*���eݦr�����s�,)Q7X��<�
�;�� �k�E�u�p��^"G��\�RS ���2P��TQ�g3c��P<�}�3�T�X	� ���.j�2^��=����	�\������x.���8��i'�nX����Jh�(�{�ٖU�f��!$1ʀ�PC}ޮC]ű8��*���E*����"MR�8��y�E̩������܏,Y��;�3�y�"-Ϋ��A3Ip���a%����|[��"3c��a�4�oj۬@:�����]Jx�kW�AՀ�������'4�_f5�h���K���h��#���M	�'X1�~�$���-�y�1|�)|�=2�J6��q�PޤJx�(�	f�ݽ|*����I)�U�ܵ4��HD�~9��0i���v�!2!z`��wSw�&����`u�_;GA���X�@�F��S�͹��$���i�+�w���?���mb/ĕifU8�� $ng��,8A.���4Q��;s�ݬ�a�@0^�n$�>Q%���.�b	�R���<�V���3�Xd����֯)9?�H����w6����Y�y٣/ ���B)��4�jy`�3����f��v%:����GyGP�*V�V7kEw���ŷ\������ t��ע�����z�q������Y-\�L���`��"�-�p�����m�e`_`;VP���-��S}tWฐ�M�K�T\U`�w�[K	�c-eR�d�<Q�c|1��cM1Ii����Ю�W��BC{?��Ɓ�bD�E+��������q���2ε8)�rc�1Ւ���x�R�,݊�YR
��(n#��_�q��Y��ˈgτ
���?v T5�ɧs������$�Mڴ���#�GK�Z(�(:�R�Y�Sk�۱v���;l"��l8QL᪃)+��(�x�&�V��Y�y�M�q��/܊X�}�h�����Q���7�U�\z4����gd��K�� ��:�}���_PH�#�;/��W���-�op|�G؇��2��y1�>H,��`��L����>���R?p��B�j�r�\f	]:{Ro(��Z=c@���K7>t�?�$�2e��lkM�ihD�xx��7�-��jc�$!xD{���m�#���e9;�����#e�xC$�Ld��[ٲ����-��gw=��7t�d�@A��f�$�#�N	���.�;��xf��70�l��^]7�g�В9��vN��p���
"���:���0q��|��#�«��,�tǬ]��D�}�����JO���j|��VM,L�:!����wn�n�͋���P�z��p�o�-[y��e(�ҙ:�c6ɓ�_�%<k|��#e��(�4�H��2v��am�v�U�M[�o�P��:k�Մ}KwK���q��J���a-'�;*h�_Է��}{+�7E�9E���"��cޥ*��[s�+;ϨӨ0�!��\�[�,�%�@4W�C��B����%�w�9�����R���ͳ2��&J�e�ރKu����t֚M9oEEd����������M/P\�y��ܼ���}��Z�����:g&ˌ�P��Jli�ж�C������P=��&��EJU��):��v��7c���e�c@��4M ��+y'�pr�Pz� fMU�t6���Bx�$�����a�C�I��eh\A>L�_�Ι�;��5H�S�����5�b�&���� �"{���ZѠP-�����ᴸZ>Oc݀J�^ 2R�0I�5���4ZO�k��'Ab��8l�W�����b��H������QD>x�l��2�`\ev��
������,G��G����<��:D�j���w��lW��O@�z�����*�
Q�MU�d��$e%�<����=�����Q�:����O�$n��k}r�+(!bdeel�ud��� �A�<���K�߂-~��b:}w���y�,�.�zdd��Pt`moWL�#��^E�E�#Y^�7�%�OM����q���o+ �K\cw�:5"���4(żt�/�j�1ݑ�a��Cc�z9ּl��J�>U�4����g�4��~��.�AY�ۧ=�H��1�
�� �����B�D�Oaݒ��x\��XT]9
�H�a�*|t�9����7aɷsw��,3[�w��Xi��T�,@Ո��UlD`�0[������	0�p�rL�f��؃�6�hm�����l&w��A_{vY�-���Iے��U�_����O'!H�B$�
�okq�u߈Z[W�ÖJ�6?������A��5��J�	sy��!��^��u��

	HL `[Ⱥ@�������%&�T1�j�#JWՌQc-.A;�E:]6�|Q����b��)�\,j�)�(YI�����n���y�"����)W��dGP���
:0�M�������\����������og3(�b�/�dk������1�s�1M/�\�X��A�ϛ0����녲��.��${{J�J�3�SjIq(�_g�0�B �`�j�M�aamW��R�iIH ��z�-�k�� 9M��L�6�"���<��/�q Dע�� �f�Dۨ��}
(5l�����h������ꈻ7�%��K�.q?���^̩r���k`��t����r��6�zy�9t�4O�%ѻ0'�	Rl���V�*��JC=�:J�b
n+��+�b!��j�5r3}��D���L��Y��C�L�^$���X���9��lE��Y5;2����4
W3`K����E��^��u�Ё��ɚ�r(D��Ou͸����؅��֊��j���|��{b��M;^7NrG�1������2>N�"S>$0/����erW6� i�-bU/�3$�AP�W�=2�~ea�g�Ǥ8U�Ž?�\7��DF�xUj1�O�H����kj| ��6��-Jd��������
��|��D[����g/�nLw۴xK0�	��N�"�6n�$C�W�1P���d֜�r�aZaK����9��L��1̙��o7c�op+�^rVha��Ӛ�s7`�<Kp���M���V���,3G9P:%se��Ε��3]���Օ�7��"��x��!��qS t�3;���:;�QҒ�[�6as� ���xl^6.q*��a
�)��^����r����K�y���n�E��\\�bx�lGM�픹9��!�����x��Ҍ������d���e:C���,)��� 6�hqTa����+� ���G���5���UK
�
���Rh��;��\�6MV�5�[%[��)HB^ᠡؐj7��t��	d$Nn�m�adqn[|B�)�*v}M�p~[�o����(h;��oU�w:����/
�6�*��恽`PX%�͊���z�E��C�ο���t�,sW/
��k�����SrR5M'��ZИ������a����Y��؋~vU�����v�0)p;��p"4T��'J[�� �ڱqO�uTD�U��i����"P���.����=`o�9*�{ԱR�&�T�R��q���2����03��vȏxw����	m��ב-�[�<}�Kŀ�4&���t���@h 6����e��l�м-�/�̵�C/�=����*��X=3��:HBQ@.ot[tl
`Կ��s��/��Z�M���tU���4��U,���M�%W��B~�����|�P�R��O;�)��A�O9{�?!�_r-'b��&��Q|�0�]F��MC���6��&ɘ��
�DGg��bHg�/?F�H�D��O߻��E;��$M&k[>�/Kϴ���N����X�U>M\H�P;'�'�CFޜ�M5[�3Ԛ @�
��b���$�V��
��C���:[h�&gM	��;��"�KCRܕ��Mu-�Ś1��#��,��<�K`%��MQ��1]<X{�E{/�ᨑP[{F혾��9�86�z�7�&�nmrYx�ik"w,�FY�`��L���S�ƈn�vk���i_��*ފ=����k{����WW2�[����%/�n�u%G�A�iZGu����o�]�o�E̥@'�"�?��� ��$�'��K�K�UoWB�%����؉���>7ZMdb��C���kA�.��~`�X�tt?�i���h�Vۋ/���Γ�(���{��!A��s��Mp���=<�pY���"�����c�3��p�&d��:�K{A��ӈx�g7K�6hĞ	�<��c��*ĳ�dDm$DLr	E6>br �{���"�d��:ǟ��"~�z�������O��iG�����l�9&���O
�/��-��-�E�ZUG� ۑ�û��O7���%��%�'2z���\y�|��R�uTp�a;��׽�����`��{�������9MT6���5]�ˋ9�Z���،6�tNv�ZK��o���Á��9x)M�Z$�p̋�,h��G�`6^b��t���A��'��h=R݊5�A�Be���I��HW)U)�e�}=5ah�JMꑟ��m_� 1���*Y���PM��i����G8�^����z���$%��w�gZ`1XE+��$��ocB��Z�#��]b'�p���1B" �8@��%��K!�4LKӇ�β\T���W�>!ؕ�s��]�����Ց������R�K�[�M7"��r6��E��k����һ[T@�3&�wdu�$Z���=<�š\`�i͎v��OE�o]��M���P��S��ŉ���SQY,Uk���_c���8m�k]��s�Q�|�/)K�@��Y�-��l�9��{qUm�!�_7�E��#�SV Н0�v�{m���� ��
.b��i�~�P�˒��W-?�.�����ӕvVj	�i���A0����"���UI.h8�\��0�&kTX�
�<�g��v������w̥j ����e՗��+�n�Ǻ�un�v_㯤�)i��	W~�M0|G�2Tj�9k�W��R�
�r���Ork����%DZҺD�ZW"�u��vL�����3Obv:����[0Ǟ���W�!Pp��X, 㙮�EM,!�_?��U������e���@nC�NEpu���rU|&���6e��Ƴ����2�Go�����C�s���醨%���,�L�ZӃr�������?�D}ٷ�#D<1�d�%��nߪ�����A�9���'�q�5����g����==�P��Ȝ��l�J3�ܒ�ef?9���m�g�/~)՗S�-E��p1=��<���y��ԩM���Mb��y̻��f��0�$�ͧBW���NٸL;��&���lz���D���W�~�y��vb��*5K��~"��g/6̂� ��Ƭ�J�bU�<B��ag�n�1���®4By �1F�ZrV�~|^y&cM��!P#��g�͉9���\�QZwV�o�8b8ohM�����􄇬 &�p���c\�(�}@]�T> T��ԛG�_�/T�%� ןg���Yqf�=�S�(QNFZ��x8ߛӃ#�B��ӨP��v�#�t��E[�c�mf����j,�X@�"��B����^�<rx)�T��x&�K7x�&@�EGz�8�&XK����b���`���i2�L�����J�U�`|��"tc5�z�SD��Cx�y:Ŏ���EC�F���}�CT�	����<-�3�Q$�x4�k�����ys�1�p6Z�Hp�C���i�5��|ه����7�T{nG�L�=MK�ʢ6r
T�������6�>z��h�����,F����t}cU�n���� �ˬv�wzsZU�*C�l�٣�#^�-N��ʍK�k�"�i��t�&wq��[._�(�$̞M�ڊ��y��s�)�=��N���������'H`����g��KSz�yr?QT���&���Pޘ������Jc��D>���;�M:y����LcR��l�2���X�Cq��2�/dYa�n kǌ��]:K�+�Mt.�e�M� ��uz���������o4$��恡��5&��H5�2/ �b��>ղ�W8�wc��v�[4�|+L��#�D�������� ��ƛ������f1`ձ�O�j,0����냌H*���y����倀�O}�K5n��A��iz���,A�8˖�C���Ŝv j�>p#�ǎB)_��;�c=�1TK�˔��r󕱘b�@����ȴQ��@U^���<]�9�?���cl�UBU8lj��7Qr�<ٍ.�#�Cf��i��D��k����7��M�Ö	��Y�t��ۥ�����fs���͒��y$՚�+�n�QO�F*��.	�;�||��Q"�N�+�=���|�<��T��-:����Lw4�������)b�?w����r	��ܯ�z6��\$ �W-F]��E��@�UO-�
�q��D��a�cid�M��q{�M��͏`@��E�� t�^���r�!���Yӎy�]c�0 ����	�����nBߍV��'�����|�34����Mѓd����@㈧H�8���SLɻ�Sr�3�G����ǁ�g�C�i�|>���lK����V��y�� t�Z��`qۊ���mPK����g0���O�l��w�N��\+Y��M�cv�6�(�_U����yJ{ѕ�����G��V��@ۓ�r	t�`0�$�Ü�d���Yٖ��T�g�v�,���I�'��1B'��@��Ѥ:�B��%���e����b�<kF�&��Qf������P�H��ȭJ�����RQ��,��Q2^�����1�Wx�Sľ�,�,̘B�����Q�|����W���M�S�!�J�]��Yr�~�E�Ft뿙�0n
�p�j�������٬�XE�)8��#�Кqp(_�Ff��ی��