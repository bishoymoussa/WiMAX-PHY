-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
WB5Z8juNRd9AQVUHFFURtTIS0ElJ7fVbpS59tRhgypbZwq+oTAR4Gs/haJ526/LD5AtlxM/AtZrB
jaN0u58UbnyRbNDH+E94egmiW+qJzYhG6gA12+q01tQYC/YoGnJ3PM/wfV49RdblA2I+hFBvmOw7
MLiyqMR7z4IreuSFQQcn7rahGJBoei/+5aWNi69f+graaJT+mXnjALPCm92D+eDtrUt0jKnChsHS
UwyyieeG1U7sy4I6rt40f7AXXxBVU1R61kPuGjcFqDNIgbhgZxgRDmifzcYGXSTV33HbGeHmwGDI
/92lHFh4v65loOKuRwCg1bq/n2SppgMnWVRcYQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 10752)
`protect data_block
xDxa3EnuGvS0b8ABhrkZx+Wy6xYk+lFCfagpQmZqNo56AUs1JRTi4zEX6OunRvfJSB8nndVAw45k
1yZq8QP5YwiBroDhKeTYFHnJq8W8DjEa+UJI9sxrhFMOBX9KjLVgdYqMntBrqg2A0IitxucvEieb
j+28Uzfov7tPOT7kKRpqfb6lVOizWlxhkwbdigD9uEI9QLXTpwN7k1RPZ/tJAzTvxiFfZBE0lSH4
PGcpGxj9YY5CR9r/batkvytRQSEnhpq8I07wTQdvabDGfvpjbLV+ULFc5iff/Y1wPn6Nz00VJq2p
5JtNJPg3Bq9pIrBZZifieONkVxqjrc/MajuEQT7YDnDjHHRVWuG1MpSdUv/jMIXhtYpNAZprkw7y
fJA5oDxOwjbAak/AZPySDn+wahlfJW/tfrEzVJLO8vF97/S6quKrBBLiaTuwyrbCtHh673AEGKTW
Dzy6Zi2no4C2BIlQYzm7yiT73Fx6IaUAIcoJQaLSxpIhhkagcUeFFvWa7QN8UcO2eAqvUE6EyAUg
2brZrqfelECSILYagbhLSgkcGw0YBsWBW75+ys4KQqx5BjgGhCEjYf358wpmglUBhsXQxP5PqZFz
hWAiPG/PYcmjmxSCsaZRlUe4DGbtmkSCv/RjUHcEeuKaBtmpiRU+AYFHnJk1A3c8+8UctjM77SqO
+12g0BohLhTVaUahCP5oRNLu5kBAF/1FmofU5rBh5HRHEpAI13Du8xOvBLzkxGJWLukFTQmTmRrZ
Q+R8tC4kEQAlgq1xDt4FSxdjozDQJAQrFLI7yytbUNYzJc8EwP4uOOL0Cr5spx/cxkJfLlaFPFbf
jgbqqOH1YE3OS8Q79/oRg5N3FSmJGmMh0Pvpw0z23sNUaNorrHqkU2+TKCOSR7D3GYa4+uT10ga9
DdsCCW7AGq1BRCi3aay3bDxkV1cYb1oz2V/eIE0AkpsdLHCHNgrWmWwRfz1pVftztU5vK+lriOKo
iF3K4LWkOAwu1jMhs8cESb5F2sCoIb48fgDPqmGqyR4MhIlHVA2uS0i2UnRR5fsB3vd9RUhV6M2f
UN8UIs0HnKIQzwLk+dyYTk77kntyzruLtCZnXvMPbHi7XYQksOg54PSpCeigzmXJ4ZsdUZ8cByi7
Eoyj6zmrmwYbvRVx3NpDVjxIlEYWjohzpTcOChZ+VpDQFchDGM3ilksB5MQzM2AVKcq9/Ls230Fv
mn01zpQ3WEiS6DLTht1y0lO/rWuvsqLZCskowtS9SodYhMstu/lyqX9/WE96YxpiXsniKU+6I47T
cw3rYstvE5Ty3wKOdENShsOG4GpsYK4st0UADBbQumnauANkX8VyxR4zpa6m2UC7SAPVmz+DHLh0
s9mLJ4cALybWFX4YO35zXK8GU2c2czgz0/4gp9CLKPxS7guUvDTN8o4/5qULvxWCnjnTB3lcpADd
OOUbnPiOQcZTImhlvxlV+fLwzp0gGNMOixWB3+jNbxaC41dBgf25H/XUeAc8bLZGOJfBWds+5Q/1
+IOs8bZQfXV+hjzokukM5xDi51WKB5KHfGOhQ68n9UKYzmm541OyuJG8g2ePO0Mza+LgMgckVIFS
UKevpXjMCDqtqSVKQSVtuTTHe/U7CUlv5TE1O+yGpBWe9lQYhhQZi68J8PxvzRMnNijeXqDBDxHJ
wj4pdP6e8dEpG7FDCF/Gt2lzBgHod8AJfIo3ScP4e/syYqSkHitzHKEVFSSYr45VzEcC43j7aLum
3IiwumBjRVmVl7lfkaVWmDcBeyO2mC6QLw3XzpSrIxIdUoxKLrXRW0BoEnCu7W36I2bHYr8NeSL2
+IMkxh0z3EHl3aMsDWwK3aiKCHonlJhhvsJEQbJFMMx3oCi+GlGVnVyh/ObI/vQnItFWScyKoYZg
1BQjST30ImcutfjUT1qAdEC8wG5zFGNXZIDsq6SYYuatNC9THB6lQUUJTGJg7IcYFrqATxfKT7hM
3Np3JudXpZw/1n0JBHCm300ua51EpUUnhDFctiQxTtXrxF3rpolIRoZ8e3jUd4mQUPFFWTWcNxyC
zXeCQvMp8IXwUX5885RU4bDTcM2iWrcbU0Kc4yUb+EVgecNqyYkPxeEw9Hygp6Z02P4KkVfSPIP9
D3Pz71vHu8VI9StzDfiz3t1DCx/ffSj8z7jYHVYcmyhcprVi2itNSzdFun0YyO1UrHSnHw16e3+j
4zkxNwzPotH34bmRsEcEoUdUeSvLS22QjVNGrdc/tA8r8z2AwdWTSDDn51HN5SkgJcHTvs7EMb+W
CxHaMA7sNpJiWQkGZMpNkKkZK5A6wL31J6jZz6NzfgcB/KMJ5bz2nHIxSx9+6l+2Jp9xQNncL/+P
aoBG/CEbcYJOC0RsMUq02nPrtoG1na0ZaVrv6gUlWDfVqJ2YD6Cl/t1HZ0tGhCgr5GLYziMpCrq4
NHHqDlp5+vAKOf54w9Qc93qZREapftTDY9eF4kza02IL14qwZ0dS0WWRUfL+hrpO05gBaztKis0T
Bc8RKsRpiCYYeqGuW1Rl4Ooz6kjMV5sE1BQifGTJuKPPI6zkUOszivvZb02vvwkEBtRPAGtgGkId
ag33VNIvHX0ZitisA814Q803FU5mefk+tzRLEkMYlsFpnQ2b6wNYVuKw9CeLgxej0wA6U7vjig5L
mHuBHnD3+Y+XcoN6Z8Bb0L8aQkszG8rZwc4Er4zcSA5HRQJ3CnpWtzjphDYHpjj8MqlryTov6qDf
36q2kGMB6wHggboTGVi5jF8RA6AkNXQvMVZsOMcICTgyBmxgkWwYRVmAEZutynDX43LLB9bol7vG
msVHw542yDdA3pvkDbcH1OG0w6lxGFhyirUd17zDq3/7Jlmbihe5FB0CjgDtqXTQAXkNNt/sfFFY
krJiKFCx802TeeO9O2lf4UeBAwswGOGWNe7Fyugk0LvX8ftPBamzWTjugpU7gb+dC0oIY3b7O5uM
65e6i/jpPBSKQ7LibUJ9kTgHMb/MRCpK//1IX5fb9PvDKOOQb2BHcdvwWEHtJOT8UJJSl39xpBEb
TNpMqD1cbEWcZ6uQF/mVloH7b/lpdxxLFGUmEebx+B4Q/ICcTeSXOaUsQEC5L8xdQ5v5JsZW19gB
GwCGgplycP4ttfxF3j8jjqCI9X373d+qUDkfrZLwqf51Pl5TsxKmq71Ve1Qd1Xwum2STzGQC/g8P
Ff9+AUBxRwP4ysJY3IJtBuCNdVCTIh9/yCBThKv5KcWIBeUEFL4UttAsjElJQC+jq0iYQEK5RfUl
DHsXGHndLA7B9iLy6u+5CSAFJqXmeEdAfkkUkql4o5MNuuSRUoPBw3QDqONphBWhsZKdMeiNvles
G24Ke7RgwtLj/yfFPEO5UPXGIQvYVmwFsgAoa2Oh6cQKAYOO2l7Py18Gqxr6UWzyOl/1+rpfrNFT
TyGTi+IPRVMESz8U6uXKOQSFofKBatq2KrEYFRBoLDiCjqWxhKsUDRVozI8/rzxBS1E5wcNZS1VS
Je7knbrzIOER4zRoEWXrhb+c+Rl4/y49BZrIXT46r7vh/Og/Lr2lj0fq7WoTCoW/ifzz3U7gQd/F
POYPUXeAwVNPe+SbXea+kc0lk5toq8YOeSAcvd2DczLlSgK880mDgAT2mWzSbq4LP6/ivu6D8slR
DkbgDGyq9UtPpMX3yjBvb/1b6M2sSmYkIcFsbZYnG08wwX1203Qt25JQzwRON8XhuRHNbOj5ctCR
ilLeJ5nBKMYZoW1q8/gI/jodK/qcCRzSax7eP9YZe571HmlSbggzIit7pTNYTBbhcaZqkkOdZ6S2
x2qkuXJTOvvfG1jULhYi4Y0/JrfXK7hp47O7yoW0PUTC8VrbdnXbYm43HFv1ZxWXkmPYUxHorGBP
gHy8v7/MJDRjsIL8UF+5QGOPrW+MJlEOZdm8Wv6EPmd5o2KEyP6Vjh1ZNvgvfzPzPa6CWdijk3tS
KUbqemPLLf/mFU1YJbYft7qA8YHRSuskAozoZWWWz95c0FTCTa/9rPot4GWCv7BUxSNZT/+/TnWO
V798ILkt6nGocwr6U8T4FgF8t/5NF6N/uGUY87zWPS9eFds2pHenncq1D05iiNuof07UaEjToJNF
lLHXcBbr8xG/f/9UBYGd57z5X0uoTgXSniw0pMbVUjG2HaLWnVx8HDcams9x3uTapNG1aXUL8k6n
Lvs21ka7fXQ5OmIFzLH+GP9XezS4Jg9YzH5tO7CxKuATXtlnqqE7rR8tXepMko4LdHdJUYG+LcMf
WHif7OwpDbgpHN3SFXtAYBi5H0UNA/ptYyK/xEIvW2DbIfcYsiJwCpcvM08GKmmJe3JBxNBZxTai
HpJL1LBeU/9AemlYXRiUxwpxFos0kJn4PYnJ2BsZIYDXCn+zK4FSOTM7himvVMp7VclNYUSDcXmY
FDH65t73ko5mElgn4VG2NAuVKXSfEYHNHqQecy+jiMyDZYL7TaT66USXBwS9QU8/eo9XcxKdenR0
R8SgDXX1ZkFLperb16lt0i3YV9ukHpi2B4wNwor5Yb89J9pifYebC37cPFk3H9VBU3AWnG4INlEG
LADCtHo4E+H8DunaLr2KMwsEGNxWODuu3BEBqCx4gU+wwerMwfXm0dFfSlwohR7YN2If2IoNZudo
y08X+g8tbGwFZJovOO6gjWAXJ4+IkoinwfMXa2gyYCznXhUGASYm99Rd8Ti78CWzkssXaZSg8pxG
pfJRsYUAKwELITFRQ5b7kvkYlXh57skpCfnXmyZYBGpny/kGXcdzyiRshz+CcUSIVXeUXsO6+kp3
+0YyEOUt4QDZ+Z/ato3+rnz6APiqwM4p1pKKAy6pNN1VIJmygKIQDfyAAHuPLdribMX4W7Rlqb2n
8nN8m65WTqtgVVxaNzR3UCpzfGSLOKLCrl78ROOXYOsNcE8WC9d3hWApJ826EV8Rs2S7VjhN930c
H7VdElH6hu73yJG2Od+lxIeiHbejI4S/7En97UiKJQwVDisE5tQgD7ykEZ50/P2Yd8XwmsDIwaFM
c1AYfj1sX1T+ldU+AZwl2Vv0tHs+4MVttXH1vOb3YFXj9ax12bW+BO7Njh5Bnm2ZwfoMubxdC5gJ
ZohxpdUbybKWSiHqbiI7X/s8P0nX4/kz//1iUH9R1sKrVUJBFS9iHxcH8ALxELaOZYHXBJUat//P
ag1rFWPjcisIFAZQvW6jv9AlQvMEeMVZjlevVN0U5GdDwqOfleTXwisPia1wzQ40CC2K6drnNfaq
N5grOEHkTxSQx8RD/G3MfOKAi/0YB0yBWBxd3jI9hlpXWu093tNic8iezQLwT97i7Dq+DPNMklZv
DAsgSkgRNfX5EVyJ/w/YkvY7CuFEq79FSZZgnCXQD8FSAFIVMAE8Ga76vxT6wSPgPAYqnBRH10wg
4P2pKqu3s17/5rkof+0NhpUzu5L46oJuHSAvb3+tFLRyO4kSRRvsscKpKIh9QFz4JN8YsnwO03Dc
g8XsI3HJY4I+y3ALTuje4vbQUgQNyBOmOuBqkg9ZKZqeWGWaLiAXCRWFeukm7Sx45vl/iv6NDKmc
wcnggDY0W629dC/m2p/O7WKcroxmRLRKiThZjTLRkGVEz1EoC32SrWO74n/7Dp/z8oScpgsKHArj
w+LSZ/lHYrzwaJ2nBpmab0kmt2Sq7Yu+NCgPqYoVGqEHkBjw81lMPNs5sOdVjpZAEL621ThmmIDY
BhBSxa8FrbCqx4/Jb79GIJi0yvZj4UqBYMWLJSCA59Z8ujooI0xTjHsN2AeEVTlvxFCO8QNeVwp5
zME/6kQiD9br1+riKHpsObbMY7tHY8l6VbJdQD2/QbTWIhy9ms5bBU7+N8sUkhUyH5VdmOSU8ZGx
mEL9+/HagMBBNjUkij7DB/9zPj1vMjQhkFz60R0EPKsW0Tzm7lVup7bAQxZKUj+jYaXc66jXx0MT
IE+3aNcBUKXbEqOmJrVWiXEOJZINAfMhSqWsuFIrZ8+xQ2sAlimkqxdjg1YFQwNCejVOsSzZcfkQ
Zmc+l4xeTHs8wC0wR2aW+OEIMBfzpMImxueXptKPyrnqvLwn8cMuhgTJZCiQfeJKChhEGtnmtx4m
DzQ6H9dzl7g74xEFU8novpzT7BUgpEkk706DVAFhyNmE/AJEblglOiZydie8IVJTBxB3VXuFxsmQ
6n6wAIOsJVm+Mru4sCCD0H0r0+bpDhkM23bhwmhLmt1jHAkr+4LA454ulRZi/suWtbCxnBtekOIS
YnZT8jJ9QBzzt5RvuwK6LT9PLYah+kJpz0gRGdRkfhQJYKAcI8WQSFeI3o7MedTGadCW6vDxVL6t
l3NzyYqoLi6oLUG1bLyeT5JIhFpBte3dTd+usWOXmGB4jnxK9+AyRoFI/zowmP9325tpD68zYZIY
u2JMwJlbtTtVrRaIYXfJrcDc5nYns+PRVGVyWZj+2+cgcJbZ/Zh9n94A2seZymgWuIktgc8ay5CE
bkGyGewf4GHpboKQ6G/I9fSoaxgzcUfLv1JR1iR7nr5NQBZk92ulbwnMuuKnupcjehU4WXj/6+t3
EsKWo1soWReauTe6d8WW+POXb43eL+UnuZl7LspGzItqQIFxhiMf2B9C555QG71im+7ERTAOl1S0
e/Y82LXSPHSxgeEDMUokxdjucZn83BincX/OUjXbzodcMmpcbxW8aGSQfaoxS79/fZdiLUemxwzK
rZe02rrwEw1z2yE11QaxHnU5CXvN3zws7yYyciDItmpggcuk6UY7G1AOJ9HPIp/pIoLgvDiBRSbG
KASj+RwJB+Z4tlAghNVziGCcZW2JKqPBGXdtNZ6gogF/ewEBqrkhRbGiaKA4B0Nz0YpB7hFGpHNU
w5shg97mLiYPTJQOZMQ5aN7gz1nzZCo9X2orHpGeeb4+KDuiN/vqUyT2kr4feHgrkP/rPryhU6LV
iOGg31wKmH7ACTgeBRmvJnQqC1++lWxZFVQ7YBof+RLubzsBxVL7WgIS5OYt6agd7ItGJaICuuQ0
X7vE8E0gdMqrgaT0ye+rTWh7WbFfUlkN1lakFEqSRS5KtTfGpIwm/RVgtMbLGtQQvDryNqGCg4AC
iUXqcT2guynXF554NHwvHC2EYhunmWFnieAD1HZbglmjjgQ5dDNrfR8qzNQAOC4z0NFj0ncjUjWM
/V1pfgCVFA6+mIpcp752qOvEtppM7FixFTrLtWoB44sl5OjWrP+nam8ZAg22PJ6wv2oA0vsfTgVn
B/36jBq4o08hmFTl/nnLT7uFsb+YOcNsSq0iuCfhxzDuLoB38Cs1+aQPuVNFucDqdOru96IczH3e
x4CeAthMz1nJK5yodtPkocueTjvoZz851fxO3NFd+Vn5LMHhbH7cgRGgtiEsuB2XKpdlkHjXbPN7
60eenaKskc0XggUafU94PWklyXxsfKYPAQwCw/PrNgQCSvizK0a4TnCgNTtFZgK07vHrqSlfOqpH
HAhgcMrlW0PAuoWFTIoWHAJXi5VlbucwxMA97bYW4M1AfmBHsVId2hmu/Xk/sSgpooW6TgmHQRB0
W1nBbz/yNGsNXNJrSljTG1Fr1vLmM6z/zeKv0ohHEGmk5M7e2kG/5anGltllVTCbYUNABdGnB3ww
ag76SJJbx85R53agscEmZKZ7SgQeBwUsjuqtfmLVOpN7dKAjD0zlKbfq1PcgonKLCS6HI3+QbrVu
jWyWCEQ0EOwzfVD1ru5eSinkGP6XKxZ8TIU2AEuPFS47WewrhEO1lO8LutGVeVPfWnpzAqa5/pfh
ZUjEpinPn5ge9mTK33LXWT5MA4inUfTy1Fi7y64pODPBJxAJNEzsbphYjg6QAa7hEb6Cz9mmj3cS
JjI6Iw36p7Ch4Q2IumMsXkhZ120mQAF4tRkLwWBUB99RBDLJqWhpgO1s6JhmZNU2DbUc/bD+ugQQ
G0k95ArmbObWpdgP2ttgCIfwZ/IGYhHtWiEiGnuV3zu/3orNDbcE+InP0rYG5lA9SOZYSXCScZR1
2nReV9HNIqheQbq6SLehCG0bcXeQVlhGUIzcfyxN7AWDLlWw8Iy3tc3ZXi6Fncm9dEkOlG24DvVd
IAvKRtYqSja+Q/YE1G+bDei6o8h5Uc4j3sSjO76XJKw/UjLfrfPzv5PvdS6VCf9+GmgCqzquVvlP
zFZ00hbX/IItSCPbtYsKOBwoeR2bnl3Q/jjbf+ef9mQaXAFmld0h/tbo6/Ub+VmnWKnkkVBphv+M
YQJ4pHKwssVfY/161EPrrQltRzfqXUZi0LOHbP6ZZuWF1H4TBE6M/0Sd/Q0lJJsda2VAfJRhyu+f
pYRiORzMM313T26dYpmUcKq7ICVaibGAblr7aelqmWC1sGngtSyE7qVHlOhufQmk55SeUD8LVr7P
gWqNuXtBppOuh8IX+9yIM3SFAqy+UYMr06r0wY46Hirx7TVblvOekreULLacH7tUp9wSAgdNLUY/
xI0MX/1o4phnU6yYC9KRD/d/e75J7NXnTO2Ejh9Spfp1fff9jicqPKb3Ws4lTMlW2LkrMVoJ6XzJ
t3mU88a/N9SutOBkGum/GBeLGjb6JuI/GKiRLkyUsfMz7ucj5pygTiT3Fm0IagGyk1cfec56svPk
s4bXuMop8vbBJsSQUwCE9j07IyNpT48yRJIwluDXrzX2q2wdsZcJZsfln/n2AmX/okkOew4lORGZ
qYo0Fu+Mup6i1YFKQDeDdrmHRACU/DJ9G1JNbDv4tsZStbRU2D5HRk0QP9ueWtgFuSqRg49J5ZNr
LOhEpQolkaisirpYShCi1klhdowoGoL56H9ocgOuv4yp2JVKJ3Ngsog+Ely+94p6h/ZSJdNCgZ+f
bfln6zS78IphE/3ULBF6n70wlLNqg3xzhKMb5foUr5gYlwuAv3MOris64QxYGZ24GJI0Wxz33WXl
JEpUzJkvBExw5QVPqp2N7EvAd1ZbolyURpmuZapWfILV6VPrksPdwdAz2KOCk5oClIBdiuHkrTBO
qO31cBHVKup+0O6vuv/XQ43ET2uN0/apnxTt/Jf1dhDJVpg80OREWTIHh9ksXvbUy3BQbHAGrzWc
OfWyfjJ+aEoGTvOKRjA8h1F3XQwbzGZw6UZpCz63p9r463jPVSQpNWP30EpVjqJBukULOmsBirNy
lHTMBTHeUib8O3n6fVX3LmUPc11bZZp8YLSPAhkM6sWLAPrO3+K+qQB62i9tHWW1k7yliXluYa3n
sh0zm5gjkfYoFTJukJH2I2MysfULD6aykbl1BddyqN7u8vYdQdWpU2jMo9bV64tuhfZzI9CSaDyc
Hx+AxEvv2zLCBFv7ZIvXtlq3q6usBIJtL1M3gtnU63GZ1iDm3ebm6d+6dOcmzba/pYQUjKQpSr0O
tRU0BKbSP+FY3BYqf9x5Lu74B8AkMHMfnrmnaI8AJui9eBZr+n7CQ4IS1+fle3A62GQY7vCJ42CP
j08pc8Pz0fHPRHbvZTB9uRS6ST+F+mR8A0R2GtTisKPe1wbwRD+Oo3OQjc7GuEzz5UnqKlpCnfku
q4ZYbqNwx7YKCC1QmCPJIdhxsXdJFGpIZ8k2n5f3eG1/FP0sriMx7XSfzkoZlx2G2WSfswjFtWbj
iX2RAGAnnEz6G6Xt6YzyK5OBz8Ec/FuPykM06g5Za8LX4Qc+zyl3livm8wB7fowW0ve4+InI5C4m
KJKJHGuZ6RuptDOLDYHr/V4ZGi1Sxuv29TD3IuWzT2ju8bLdmyvq0pI9FL30wwxg9GQ6P8fi1pB9
vxWtNvyagq8V2wN5cpHXPfUESVhIy9qUu+2AIl76BoeWwuEbe2sLknh2ADVZ4UMfrX6q0718oFpR
ku2Dd0imy7aV2F+24IacEk1cZJ5T1NsPjxDFzMVDptZ37XCDpwrom5w1qCP89LCZlIAo3tq5Jigt
68ZojG1NwUItVYb+w5RXWeW4RgRvZv422RxTFRIwYEeFYQERr9OjTULlOUPWOs6vv78YQ82pT0h6
R4JWAHPHyfKDeC02Wn4uuo93tedUT9isc+cZEkT7F6seNV4VxqDtWbcDC4t+h+4XqExP3/y5Px/P
Gva98ONETa/pb2z+kAbHysYvPJfiGgdgxW9JFySxxi6q1YE//8/VYowEqDQAfei9J45CeMTdma00
raXzm7HXaoaz78wHVS87Z84FhjMLmKuCtCGCavyj8QZ+mmsgUnxD2nyEyGql+v8urLgn6VPz60Sa
P0jJH625onGyJdB37typLrUHrTp5xiZd2tSS4vW8GqyQpsVfBLrHRP0EIZvzwaxFtsUGQ0vvDNrQ
pdB+jcRBZodnTjStGsaezfW4VftG3CnLdSEEPw9xXkw81m/pJWQKvqkTlmwQ+DkJSu1KFwkjYuSD
/wjV/S4J3YIGRNjXn84RBVYPlzu3g/k4RwOz+PiDgy892MT4H7/XkIvbbl80DWjeRlSX6LhUibtA
xeA5+Hcbv62rjW4GV8eZBibC7oCovbQWj/wqbhXzRQHoWP8uwCowr9lwyrgb4S1ps2qB9uCWQ3uP
MLFKLyyh8QU9sl+/hPy2/sACJth4ZVWd0Vqrj6WhETRkzX2hcIOdy7sXqim7EfMKBCsq295D5jVS
0YA7CU0NBSYvxaFWfRS3Tnzih4OWfyW9jm+G0DorrwwKWhRw7ALOh5QDEdB3aFw5av1sFVTmKb4u
O/Bl7QKm/SGw8y2wkYvEEPc9NtCSVayCab8CYLAC/CSk1OUkalRmtqLJXfMwjKJf7hA1GR+vmk/o
ZQR6uE794W3EL2o1DEzUNX/drMf5R94+KC4b7DylELlUy9WsZ6bFWSOWRsf99Rr2OuDSjZHLK/vU
8TL2nJXPHgG6oHQSMPCcoTFbBsnQoHyO6Pmu7Fubrq1YerCpuOrDymQlRfNs61wN1kwanx9B2E4L
IA0rP8l0/lMmGCYBNyolHVz6BbcGVahtlt7hxD9QwzeEKVqrwBix1zOnklVPAy5z+y5RKdbdHJZ3
FMF7J4yCYlPraJvXNHKqLCEf8nbaVSqGbU2hECgwTqqLNNoCXBxuaG0A2SmdcTZD92gRIrvNl0Wu
7ra9OhO9782FMl9fjnUOcxFupDE36Sl5GLek+xVBRZ2fsVwupPXgQEskAlAzpDn8tLLH+IvXuAGq
SA0BpI/cuMP9fguj2IUC4e3xoaILT/QUfBLYz7igVf8LBjKeahDoiqH83aDkv50EtFunNSBQfuGa
zx3axqXZGXVo2HoSYodqtyJl2ngGHsR489emQyY05UIgto+vgM8FDu+QU97z2fv7AWagg8AqHnMN
Id0J5ww2rF0I6xIo8+foi6LM9wD7RhRujpC3O5QNkcfaN5NJGmtDDOQJgK0VfyYZ8iykceqfhgRj
vjLbTyhnG1q6h2WDzH24zC9DKH2R7f/VglOYRU0uAcp9SYQfVPpJA7l68D+wWeLgR9+UDTVJT+qX
ltHpqcNptrwrL3Uh+glMuc6dgnCp5qNhtsY2IzR++gJPD6Zb1nLsLe7fNd+fk2HSfb6vrfBMwi9+
8Ja+YwfBSXqJ4K4baWeWweWFHsz9zpWtmcmFJji9YKypuNC1kYH+YhrTi/9CNf5OKMyMEemWP2K/
NNiuoN3geROmse86Cw3wEJXhylfJoQ5qLAcvOoPDWK1xkrSUHDzpTiyDUP7rc3/f2jsAHbOVicuo
8Mxcgcqcb9Mesd6UZmQnxOBsjZVyT/shRhosAvTCY6Mjyx60opU/z9bLViUc2J1BJh3ip3pbUcQ/
t5QOu+an6+Fi7Zpj1uUhSy/KeALonK5WmQEHjlBlyC3HJUqyrc2jgapzROtGykXcYYBxTL28/Ybn
3qVSvhpUNoqwuhD75lNguuJjpI4gPWqOlDOMJEfcEeeOHvd3ABdZ10/FWpdovayKbTlua+sgCEzW
v5pIPOuj//ZZotjdWTTCZOEgPlwPWyN0risrty5phHomJFQaVKRlJLZnATXSlDcV1wIy1Qv6+awn
yEUHnMVqhEmmNCsDvAT9hSSTNe30BgquUM4m3awQRT9CsyuIyEWsa8eH5czvGwVdV6FJSmiELG2a
JCeTeYzhJ+vk1iSqihjdDO8h6J1aeWwwvGoL/0NFurL295ERMcb7Qd3lVc6uTO4TI1kmHjmBXIL6
3OvkTq0cK3sMKrJuSfvcXbw7Hz0QRa+QHBQtFPVfcB90LpkPcs2bSQd/pieqFlLyvn9pXd7slZHI
sFF6OrryRzTiSGVflamazdiCqiIFUdSaD8Nh0B3VRdURaCWJfvUJohxrkRdXH3hruBA4FKbg6fP3
pZ0gaDqhHmB6cXFeG5vSJYixIyq1d5XWEk212QE7aSP1M8hjyjIEqPPjd9c+F4sBgVgHJaP+9JmK
Gm/YxbDVf+b7kjITJSQk0iQ2q56L5Qei2M7YvkLvwR4MMqSdrhIPS+VZHHDYA2UV9qYhY0EOHxDa
+b95afI+rNmX3m1aycn8nYFdw8uDLbJQyxoZwxQM5iuKtKuIaqzPL+YUXkPe4ju0vETVS28MIpXS
NxBG15a0zN1KIeUUgj9ivJhRzx4ULwBOxsYUHanAk4WnsdEwQtJaho4oI96lYgqqS1GwWQxXopWa
qlpnEZohxS7NgASHx8cMufkm/zcx0hTp1w+6RNRZv9rqFX1wOFQ0IOcIsJp3LbfL4XXbzmGpRfdE
BN9eNwBr7UaGU8eOipKlwJKK8dbbbXL5uS0TsdvxAeNaDIvwqK8jjFqKQKoz1oTGJa1n+Zafiwx2
UZZ84QLomx0/fl28qZQWfoLYFeMAXdcPuein3yecA08ZszqnnpYZS2PQijxF1+RDyg7Gmm7puxbt
PtkFJGq7HFGkH2w/qJvGoHrV28TjBhxYXNuyU2QUKlSVfxR9VIRtAvw4OmGQAoc7yaa+GLcEaHDh
kSxsObp8GPoSuGakozESoFZzv1FZyv9xQiSW6U5tkXgs8+id87QHxwQjp+QYXxSEWvAkAJXj7gJd
/VnhACvClbKRNc5soDBU9pdQXNR1SL1mr4GuyxjQED57D7+RxbAhwlZkXJ11G33m9uXJSmMLa0DJ
v/Dx2ZXw/0Dik+TwVf6aAe4KIvrt0ZTk2rfH8ob4w6doR4ES6Gf3Ig3kZnUKi8dlRJ+j0eLkL1vI
8bKZZ04if4h7J9uIycSvVYpddhDSLZzRqc1MGVmbDrqYqCT9acr+nKK0wtgLo32MNjUVVqgXohjN
jInlFYv6+lrb903DBijfwlOnuvFR9L6nbGwkPTt4SPLXlXrezhhuoytj35OgZ156/7ubX6m3Y8r0
RATL9z4Muq7q34c3o9wBBsal/mhIflV5cE49lrIRBoOf8hBZnGK40o4xbv25sGSTEIS6pT5paJPl
b23nh83XD1ckqzcMNm1rGMkiMmPJvvWchzQkwHv56JxCVIU545+HiGNzaeAMDUUhoZMsN/7rncAL
JnU0kIcdyLrlRB3UYFbmsVF9NAarZv1A5wVImsQw8i6151XJMGVehGjwxGPzLgnBsvmMn8iK0/4V
0x4aEtqVYJxp5wi391CS7oR8THxUipKr4Xnm5/ReSFSR2L1N/UDDn31WqmksC+5/nkQF2DIMtowk
7znEOXSVCsHUBAx0Q5egVnGCV37t1IoeQbGb61yJ+peO2or8W86G0xS+N46M0yoCynlbmwgkhebe
v7gWmwoKGU8NfH+AHzSTEKljyG2oUdbpZUUTsiUbNwyC4jIM10brU1fiM6rT+kXtwJXNAXTxcfS/
zBpbPMgaI8YcBGiOL3mRhaQ8AM47IA9C2AJnxSQJIMK8hmobklQdKNA+YEi8sHczF+Vl5Ein4BQ9
z3scKLBZf0/IkN5+mmK6WsN0CQNHYQVjf4jaGblKZaL5Gdn4ohGQ7wBePOfgxeWzB+LdBDRJCWdn
2s50wP0wmEcS0ydiMccaWP4lQJOVZxOT7a8D+s5CuBPDbUHyuSx4S38mKjA7ExJMy5eZo/IBeM8i
7X5UgifrxeoLFG/Gnse4ECg+DK37iqv/mFn/7WRm40wS8h66Zp2qOcGCYEplyM7JDaKkjH0TTXxz
LhoILVWBoYwjaIk9/As1j6nWwWbBOT5Vq2auilu6vUDxjU1GY+RABZPsctaBr5+W1pGlaCrlPViJ
jUQW0I9vDxFQhxx5zu4oGwOnTG0HSI9Ql+gbA24xP6v9knllN6yLt11esujVcIsGfL09u0VkYGG8
XwEprkrwsTpBdmxC0XA3heK/d2EF8E/4NFwNMpYhDZ7YyFaQv9cJQko7580sy/H2+GaAHiPtvJN/
0E3d7g7OcqN6PjeTu9JMo6UQA3ysMz3yxKDBcMTEGLSTo3jHr3wKSbPWbcLcdfB9bweJg5l0I6Kc
IxsDWJ5p/HRRQGmsT7rzsRcpR4bxEB16kcninujDperMXrnV
`protect end_protected
