��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$Rx�y�<��wA�*;�x���@�̦�W�X�fa�M-$u����n~�%���P�$��W��kYَ���P7�?UMfT��q�6�U��k�>����~�\N�(�����X�e���/6U|)�X2pF�]$h���d.���9E��WG��L�X"]�Ad����ľS���8od����e�GT?y	7�������ݵ�^��R�q^]�鍦�����s�ae���h��L��P_���ާ��YЭF���'\��68�b�[����w8�[X��V�F�0͘3����q諵�uW� �h�u\V�?@��_6G�_�*�G���B�絉�f������[�G��U&�����~�F��AׯK1�`c��[<��FY���4I� �#�G��x[X�=�Q1��`��R>(�w����R�O�?����7�,(�H\�#h(W�EH=�������yq��Ѿ��aF����:�U~m<|��.��0=�P/���4ǆ���T(���6̧�w\�D�4���)�����iW���o���j;��䪹�Z'W7mK4L��b)�W�N��!YDH���j��XH�a��:K�	� ����g���KO-�GLH
���9���i��(�
*�T啪�j��*l�S��gf��1��ky.�&]��#xD��~�
�'��������f#W�n�?CO��@$�v��K�I�e�d�^H��lp,���@��l�ϵӯD�rd �S�FC���NWF7���6cRB	G�[�&�0�O�ȖPgj�
�MS0ﲧv��� 1I�)��SU�����fXg.�/(��\s�#M�4���k�;�@��_�a)c���7,4��Q�H�Cr����Ȓ��S�0�8'$�t��*�0��+�>ʕ�y�g*�,.�w@	Nȳ[+}��.ݩ�����.` �_L.��g�'>Ƅ�^�/.k�*� ��qsN����#*�>�(A��E�8��ǫ�2~j���@��	14{������%kA�"���Xq��G��xwA��#�Z㲊�\,���	�PQ-C\|���٢|`Rd�L?���v-Ʒ^��N��Ռ"¸`��k��Py���$@�~�ҳ7
J!!4����bL�
,g��S�X���fܢY�8��<�W�;�kB��^Ł��q�����782,�*oAj�zU3Z�l�Z��U���'NI�ꤳK����٪��
������piNw��P�oEcb�����p�~�1��fp�uU�!"���^zA���S�h��>T�ػ�Q����,�������}6�{w
�r�e��{p��<\�Ɍ��,ɖѱ���k�j�lK�OѪ��B�:��+�)����X�c�P�S��������@<F�UjT>F	�Y��,RAf���-r��l�a���Hb{�צ	�nǻ�P3�e�3@}�h��������<޵�/�(ا���iɉ�ks���1r�>@��"��c��J��/Z�؉��NB�i��\��qX�	��7k�<�5$����d���]��M�>C^r�d�}���M�������0�o��HK��*]���c�!�=o�E\"t�H��4'�*R�?l飨bQ�5�z��!Z���	�Pfv���� ��D��Zh�����\�ڵ����"PX�|�����ae���;=���N�䙗�1�Q;�Ӊ]Y�L-��L�)�dC۫�c���[��ާ��(xb�3'cD�6^�F�Z&�]�����j\Ý�ܸ�@�OZ��Nc�r���%aĊ#�k�^H�%:����ew*z[��\�4ÐC^ZraYk�a��"��t���W������a����2/��k��0��sz������@�L�ˏ|�H�}�twjk�)�W���^���`ճLW5�u4`%X�^��������0б��=Mñ� �}*Pպzt
Q�T�5��7x���p%����j	:ӛ�"������vSp�Hr����삞t��,`TB�5���iR}��t^�1��z�DX*�Z��%7��F�n6{����|L34�ۊ��� U�} l��6���^��"����@q�2$���T=�!�3G����� �"v��p��k�����ɫ��F���_���hc�]�K�W�+�� �z'���H/����`�{��Ri0�}w�#_�
�ZL����E ׺z��I'wN۬���
�$p[��V ����1੖6����k�%���sc-�йV��MH�������Y��s�=�`��T������	�L���5�^VۚH]"'Bw!�1ڕ�p,�ᕔϟOj�ŷ@�t(ԅ������~ZM��Dj�F".�}�x7�Ĥ;+�&MwĖX���4�8=B4� �̘��\�-�����ٔd��q�=��o<�f.�[W=ʵ;o��dO�fV���L9��ZmH4�����B$/�&�����*&�ȕ*wb�Z��22CAU��E�A�Z�?�i����W'���1�pY��*��
kJr��པkl% �ůF{s����(_0-m�rUŕi�^�[�P)
MB�gB�1u��'�x:�?�c�������x��&���7?��rLA71Pf�}
����J�v������5�Pvs/G*0��A�EvS{N�!�/c���!���r��Z���3x�Ä1�u|�P!�J5l�C�W���������c{vЂ�rS{�m��=����=���*�$�el�+�DR��2E��hZ�M=�k��=e�&5%�0h� t����ޗ��ruZ� ��&qA�ׯ��q�oi�qxfk����#9�i��4X�4��$�0�ZD���(�9��je�E)�j�0A�����[ɥ�1�S���%��C]�rGn�'lc;)\\�"��(ɚ���(?-�J�K�TB���0��:2��ʢI�ൣw#'��"��DaK�n��#�;�I�"��JU;$/94�u[$xAxA��`pը߱m�:�.��r`���qٲ��n��U����0�*�΀�R�Ě�����+��}B��P������Bu꺱~1�Iۿ�w)25�̩[���������������u�F4�x����Ʌ��a��P%��E�2�u�%d�p���䁚OnJ}�NapC�b��
y��co��=��9�I�z<�D Ô��>�s�Q"'t��Ừȅ�RBǵi8D��d��Ƀ�];����2��i�R����� Y$��rux�@<�V����Z�k�Q����q��#:����{��y�Q���.��81Q�x��j.���O�]�^Ly���xx��k�Ƭb�6�M�;��_`R �T'��=<�;TB;��&���Z�\��Y����� YN�?Y�7!ڥa0y�ܓ8�	��� ړ�����d�	J����.�DHi�-XG8X{`B����[�D����!���ǀ�����2�F���c�[���u����y%aͱW~�ܲ �ts��`�n������S~]��K�S�ǜy�M��Mw����%�a�έ�Le7��;�0��,XVg�$��}`�h�����*�il�R�Y�N�����v���_k����Y��%��aZ6b��rHT�a$&�/8�������յGm���9%̇ඃ���i��J��!��M�6y[߬��j�QW��#��y	7u��
�F䩻q]���oi���y2Ô^hb0~Q�΀�|Vz�V�C2�� b���rV��d{��:IIp/cH�5��F쭆E$ )_x�ecF:�5%a�0�j����D�
���F֥?In���5�w��}U9��jf$�I�P�IAG��G�(T�B�eyd��xG;�Ԓw9�d���T1�[��o{I�.I����=���9|�jq���_'�n�D[Dݷ@"��(���p���]�����>!�;B��W�ު5�݃ާ���[v"�a���F�!�e�Su��Z�!C`�`�f�f<��.�:Z���P�>��x����rW�����+���XਟՁ��,��0
c��ȭ{�%]��F��)[�r	&�J���)$�YC�S����l0_���e.T�wY�C��5i7�h��!Z�{��M��Is��{�OI�	e��e��d#!��>{�2n]���!N$��B���Q*@��b����CR��x�]p\4MS�l��4�T�.�~a�
A�d��k��ZsG���cEtݠ�h��PFt6�g�è����:6=�٠���7�E
���1�%i��s�5�m���di���;����%�����{R���v/�&���[R�^�T��B�63���h��ׁ�u5��6ᨾ(0��K@p����f�����[�*)�?��
ݺуsD&W�]�4�Z>M�C%��l�.�z-�����I�;�H���ӈMRp�[��&Ua!Ȭ.OGK��p�1�SH��+�NE��}��pD�:,�Iax퍲#���/=c�߱.�H���1��/��o�ާ,v��ɝwp6���Yd��#GmQ'|"A�<RR�Ma}�6"���C)��0nz5��f��r��������1����X�ڱ���تťu��|��a\zi�,;��ې�1,4�k����RNo`A����+��$`B���\Yh��GE-�U>RD%M�V� ʔD����Wj�h)2�l���hb�-�T��ũ�1W���}��*(]ι�2�rs��J�����WO�%9�j&�m�*�
{��6^�!�#�x�����\[Mb��HU��e�a܃�@w���7cV�n��ا�ס��Ӧ�ʏ��S��I�f& �#-bK�i��c��s��ڒ{��\_#�F8A!�6'eJo����tR��O��3X�6��G��~g�H ��ދd�)����	�B����U�Ȑ:Nˌ_��&y��z�*�q�U���J��� ��#�:��WS�̠&��Q�/�'(Y�ru��$C�mb�{��V�����G!:��{����4%�	Zd��[A;t�,L����L~_��L��`S3'�Ȩ�c��&����ly�J����F0U)�tp|��4yL�w�ՐQ;���B��^·&��i���o5��b��h��T>q��Bk��
�~�2#	{W�k��i�Y9d-G܅MS��ND7��<X�,�È)���>�_݆ćq��(��S �&�fd�3{k�D.w�F$0F���+��yks!���l�/�W�iʊ��$�fcP@�t��;N0J^�^HLzo�����N�y�/�bN�nJ"d�3��,O�n� �H]����+�(+6aJ�5�*���
o�2B�	��Z�U"~���`;���MP\�괺�R�� q�έ̎����<f�c*������Bs]��t��{q�#f�#��1nXEe��3�Q�_�2F�|beǏ����(��Vޚ��P��c��C�ގ�����CP����tH�0u���h�Y�QKPT�gQ) E��z�!!�>�6�����E�� G�`c����~���^�|R���Y,H?Fz#&����DW�u8]�����8��/ۦ	~���d�rE�Q	z�_��GJġ*Y�=f���FZ �k���(�T�j9����\4�V��qF5�0�*�8�DW�G��;�E�ֶ��'��GU�NQ��_�\_+��G�R�(�8:Ƒd��ݥS,����~��5��=��f��`�IT�eB�t�Z涛~��.$}��A���\鵙���l:���>��	�`o1��������1��<�y�����.I3�H5`@�-Tl�h�2T���>CU]:�Ò���k&���AS�d��(����Z��e詒(2�.~�M�2 0�����F��@�d
2�:Sk>�=G7B���S%�����^����.mg��??`eh��5�R B=8��9Av�����C�nD
���硕rߙ�a��
�;Gi�&ZPu���ル
6�������R`�M"'�[�?�cB���'x�<��@$gU���|Q|55��-e��᪀�W��[�E�{�̊��#y�i�ā�p����hͤ@-5'��5$�f2����������g"ΔL�BB)i�PMe��O�#�i��i-W��3HG�d��"�� �hS��?skߓA8��HJ��#�K�t�h��������-\^t!��`7Uvr�\�{�8]_�du�IU
�G�4� ��v����l��w:e����nx{C&�����0�XZ�'v�4�`�,��7�$��t���p�Ӣ�I���ѿ��r������cϸ�4j�Y��&w���I	���H�I>�����a�- ʍ-ɽ�2���?�y(�{T����"*˔����5t�1�cͩ��.y���#�P�ݻ��1z�!k]������V��V3����Q�Fz�y�A�N	��^e���T�
U}v������u]����,4�~q� �VtXN�����7x�xn�@L�9�'ms���~�����3�Z�䲜�ba�n���	��ҝ� Ƞ崛�c:���-fM�*�x��V����~���w�����#I���~��Nc�Ol/��122J�R�Ȗs�W�l�%rq�����^MlvSl�;
1�8i^��W���6.�JԬ6uydK2R���C���8ܓ��[��3�!M�H��?آ	^$�Pz�ԇ��)�@�/�;I���Y�����ɞw��.��9�ęN
�4�n:$���l�*�1�!8���Zй�`��g��M+��߻��pLۇ�QM�&IB���9����㊹�&��T&�`Ӈ�A�3WO��k��f!rz�eyuK�ݳ4D����������J]S�KSBP�3��8�̠���F�hA��h9�ׂ�Ŷ�j�˾��?O+��vؘ�Xؔ߇:5dF����ߍt�Rׯ�G9́�Jp>yf	 �����C9�����^y�=f�$��~�܏�Q�x�#�=Ĵ�m!]��W\>Wl�H-Ys;�j��y�]U���h���0vq�X0"��[D��e�pAa+n�4�/��򈯘���)X'���m�$g��E������}C�.�424@�9L����?h.+���N�ڔ�#����_I㦕�E�E1�|)����]�KĠY%��L����;Jg�:�
7X�i�S����)TF����1�W}���e�7���#ҚD��4� �
Fl
��IAP*q�A�	bT�6�*-Q�˸��QA��ѵ�Y�(->���ڶS 9wM�*'���#�c<�T�%�8B��{��!w���i3�"�℉u^4(��%`F��ұw8��R�(�4�cEJq�����_�����k%���U��%��E#u�g����d[Z	�����3]�f��z��Ũ�c1
A�k��]mR�&��#����G��q��f�V�Z�O�f�ck&�hriL�l`���@ ��!R����+���nl�]��\y���e�����(p�]"f��e����������J	��=����j���~g#��7�"�sJB�{>ʪ+���)��qLu4[�HB��@��w`8x����1�A�9Xc툉4�͌�qBF�������T��Y��O��*�۱�Tr�r 㩥���dr<";����b�~]���p�8�1�e��D�![,�X��Ҁ�Q0�<��s\��ط�����<�ݹ�d�u��Tέ�~�ƫ�l��=�`� �6 ��cZv>h΅_��'��A�Pk�.�=`.��K��R����QFAAf��T/H�N��o%�g̲
'7 �+/ߠ5�7��x���oi���f�2� +W@�^q+}�ؤol�_iۃ��������a\��0H�E�X7��Ol]��o\���`+u�8�-�2� ��w���7���?$�ɀ�A��9�U����ޱ 8�E<�����c�aL9-�>ZŤ��"~���0l��@��ʗ�Mè����b�Au�y�u��4��q�h2�XX�X�
Y�j����l�������,6�60��V����o�g��|���)Aq��s�R�OF���7����N�6�Ta#�K��-�j辕]ҊׯC��O'��p�>�L�	�����v1�?�S5ȚJ�c��;�*m�\Zu5�������k{p���� 2�펤�>pr�t�P�CC�p��$��V~g,ô!j���@��.�O²�������0J����l�0% 5�SB��{W�J���<���Z�4�u����v~>F���5�t��$U#�)��F�p/;�D�ʨ�ĤMU�|"WHz�Y $�un�}ad8��5�m&�U������������oһ�� ^��N ��ՠf�r��QĄ8!����� КR��#]m�H�4��}䗇pE�_�O�� E@� F�6P���E�L�ln��b_0/Q�8���♶c܃�1�Eq��c5]�	�_"���G���{�q��3�A��H�z�P�`��.���{�� :+yB�Xa�u� ʬ�I������t�jB2�Va�x5���Q	�"��ІM��Ѭz�ʔJ!]J�n�iۃh�4��F��l�'�)��<�C�v����k�-�?Q+<6\�.p9��
A~J���g
���[��	ۚ^-�Q0���>�b����<��`I\�r�-K���)7�0��lrI6�(�Z�;��e�X�=%���E�Ԍt��u�b���P	Ӄ
C�?��.�Ֆ�<�d"UMs	o��/����n���f!�����-�ڀ�'�LB�Ʈ���"�2��Cէ�E�N;�z�vX�|j/��O5A�tܯ��MKa٪��i��`��1Eª6���"�����g��+���A�TUv,�]!�gGYv��]+��E�&��������g~$�ϵ��4p�h�3j[���a�[d�q��\;�)�_F�?��3���l�;��Y�2Pu'�Pg��օ�
-�.�1����⿝�<�0�*�n��x�-��������BlPp���Di�\���Q\䈚�������	�.���mO"+ڟ������.N�����>uM��$ާ�Y&�ΞH
ÚJW�U�����6�#����w$_�쎶�JeK큫M�-J甤|�l��,�(=��_��� ���9I_�+�W=�,��B=�^������!w����r�ܯGo��G�Ȩ
5�|	��>��>���>ĵ����]��9��Hl���d�-���ph�w��,3~� :쌩Ϥ�,2��Db��y~\@�^��e��$��E������7�g�a�R5��C��fh@u���!Vj#�
8f���U�2�1�҂gL���z`��4(s�!ï�&��~~��0��T���>����Tx�
t鰼�$��d��E
��7`^����	u�Wiнi���VM�Z�{h�\']������ր��,%���Jb������;�#���
%���Ca�e1��Ҽ����r�{f^:X:� �N��]ڄ��ͼ�`疻�KWfvL�P����%g�.7o��6��%%�}�*k`���5�u�J�)@Xׇ\`_��?�x�͵$�yP���TJ�<�;��M5HcK�r��{�ս�6�7!�>�c֩CJ����wi{-�\�}�6L������k��0���ե�#r���6��QD����L�����_p�&�7�v�>N-�t]�,��N���y�v�P0r���M�[C$�<�+�D�L�3����#,v(엩憮�C{Y�m���qjdl���C����T���Ǿ��8�	k݈$�8���n�H�'�9h������5!E;��1���ڨI�R�ٗUE�Gc��N$SۆH��x9��fu"~T���$H���v�et�#b���Bе����r�]IW��$`�����y3��%�����c���FG����Xc��]�a� c�HQ���v�_�i�{�$��<x����ʈ"Q��x�*Jy	���G$��3��8�<�ן5�,��!q2��a���&g������ю*K�� +� e h���Щ/B3C����L�E���050��b �z/�<~��ѯ��,g�S�o ļ�`R�./��TP<�Fy�+�2�$�}*A�.��*��>��1����iX5V�ܚ;������+t?$D��S��.��΂+�(I(���L�_!
.�Z7z��ď����Rn����Iĩ(bw�L�!:�W�����xZb^��=-�N�&f"�ʥme�P趟���]����^�"��?�d�*E;�8����0����<��`e��{���e�3���2X���Ɏ�ߙR%�P9x+��z�+e�#Ϣ��0�Y��Ξ��
��t���u���f�~8�A�VaA���p��N���<(�3�3�Y��ƤW�-%�L����vl�HV4�ѭ�[n�.���h_�EK���Y�v&y�9@`|�u��"E��`�ƭ�~+4�f��]��?��TBD;?���V7Ӓ[��꒼� #���H�kUY���د�+�(p����,��*ũ*��0��ގ�W;%�n0�	�7>�����!t�b18lF��>�`v��w�DS�P!�L����jw9{)�`��0�#�Y�$�"q)؂�c��2��������:�ڝ��G/��5&tQ`Jy��E-�&��-oͥ�ԧ:�����p.##T��'��h�T5$޳R��=���R���*lΡ��5$@��,�>�8�7�X�m����W�{$��l7 �x�_{�j�O];1��w�ɻ݋x)�:��l}�<2��Qj�t�X���N���t�lE��&��%�~�@[��"�s'��(V��!!#�̸K)�=^�	p���m^�ޝ���)�������*�pI�3�7��
�r�B�,R�V��
��XCU��ޘjw򊋃&�e|:/Td�/��L��M4�K�s�];����{�����"��!�%��@3s��NO�|�R"��-ǝڽ�E�q���tSԐ��5��:c!�vָs���sD���/r|���m�bJW.k�e�\�|���Q&��˲e��6�����s�R^Wָ�#�EX�X�Y�kL,�:Ѹa��~��a�!�?NͲ��
�����J	:)ֶ�R�%�G�����$͌p^�o�:��u���ѹ:z=�!���|�c	�b�!b$@o�70e�� AȁF���<�r8���3l��aya�%&�
Bl�������2y��m?���&4�����d����	grm+�:	�-��i�ve^��C�9�`6�3�=��Aw�B@J@w�P7A�`#�ʊ���-e����S��ޥ�&D��yo��\�m��"�W� �2cVH�RI�f�:U:��JJ���>TF
W��{�뀶3_1�����¼���Q�rw�?"Z.�a�/@	>6�.,]�h3��r�o��O����������W�Jcu4���K�ΝLڿ�P�7�x�,���9��՗�:�XL��[�+�2E��35V*�-��z�d{�!������ h�yYbp3@�a��LV���S��e%ׂ\������[��Յa��<�Y���3U�D��~��*N&9ja�����]�G\��{��w���E_ı��/�9dZCq�/w���ӓ��g\g�bC�Y���������x���_�H4�Qf�!����*\.]��5c�0�b�"��Fի�mǤ
���I�>��>Z��y"��������O��m��&~m����C��M��U��}R�����@[���,��r[ �+�`J|� ���ޗ��WJ�,]z��@V�Qo���^n��Xz)e��2T�$������ �_]�����Ԯ1ee��_vɓR�b�oCx�|3�D@(#�5�����;*'���q��#�Z�9U *�]�E���"yeu��k/O;�P��;4{n�����몡l���g�y^J�5#�smǵ�a;�u����j��s���;�fLSm�+V�!�^���ɓ�ǟ���}��최O������z��Wa�cToQ�����pr�0�Q�Ϡ��:���}�
�1�a,���<�Nip̖��՘�Z�B�Y��e�,J�X'���x��K��e�=�zd�<�VUL��<4��w��={%V���ퟆ�'�v�tEI\�(Z�A랇�{C�.\�5t�ó����f��
2�@V4�cZw����� ����2�$��(����Y`�hRƴ�(Ch
�H+��3��X�+���,�/����BE�"�eix,&� ���d7�{-i���e��q���ZX)eu#Z����$�R�=�sFMm̦늟 f��8n@ޛ$<��ω9��n뫾����j���/���b�|$�Rn��5 �õ�������s�)F�["�BbIt�g�8ܑ8��ͬ��ﻄ�y�ǽ��I�z^��F0.CT�	�	���d8��z�M�;8�ݮ�E�_LF{I]b�eb+8$w\�L�/ / �V�ԧQ�bg��	�ÿ�\0�����Q���]�V�<�s{�a�Lf�!��h]�N����b��Ei�
|#�"d�;h����@>� 	�~�!"�:�(��߉���Uʗ��Q�PF�(a�Ʈ�����|'�H��/|�aX�h�~�ʤS�,�`~	��F�B��#C`��J�r�d��ں�����3j�����~��e�k+ۻ�N��C�MS�f\v�2t�y�3���`}�VwH��:5���o2c�8�+��c�J������-b�+D�6��|l��wd!}Z��塉SbSjB�����.R����5��W�	I�r1����-�r[�XT�`��}ou���l5������Q� �3�îX�8Ϯ���K�,k��7"�%n'�rM�)�مa&Q��uCE�H�5;of���<�Z�9z�i�G�`�����n��%Ļ0�q_�<O�:o��S9�!������J�@��ҳ�c��+�oӱjMكI�H��߮D���.]�����kGj�d.6����t��Y��e���"��F�(���崆�aRY��c�9�އ��mԵ��z3`��0�J���1W��#6"�a�w�!�%��yUU�s���O�-z�R}�����2
�}|�;�ʯ�5�v��V"��FB,Y6^� RTh$�,�+��S�s��ΑÜ:�޳�5l�� b���=�5!�����
�q��:���ⲇ2�x��1t;(��Ѡ�{�}�R�|�*�}��U���~n�h�߆	P-'���O��n������$�^S~κ_Vq�}�sa�>L��u�̿�EG��F���{�Jٙ��67C��a�t>슅�N5�	���!���3�՝�]L�w�$c!����?>;rD)x����yǸ����G�4��r�x�a�̞e$&�f�T���KB��59C��M�R]չ֯�j$u~�q4�.��Om�_a�R⬖ _C}��	h��X��4<<����}����x�`��;��|�։�@-�1�[���q�߉W���4D��1�"����@�o��k����v1���RVv[�t�!H�Ad�6R�"����Ў�dj_�l�=�߰W��c��+E!��0����1c�`�V@�[�\�<"�`�!�Ot���6���d�d\\9�)����ؔc����ޝ����t�C��B�-���5}� f������\�;*���A�W�q����}u@���Y��,M!�r&Z�J4��!y��F��zt}%_��Kg���[�z`����;߫����;�b �Q#�B�����eSj�Q�E�WX�������^p騢d�v�3nW��6y���H�v��@����c�ۋ�'�c�f����)�r�C���B|q���㮂O�%3�4�33�Pyv���ŭYR8���&sM�ҩ^r��-�ޓ���	�D�%�Wٙ��N,�l�JWL�n	H�m��(�~�n�q:G�򨛬���z�ϓS���7Y��A|K�Χ�ܨ����1�En-WT8�0q��3���L��QxX�|�W@#��.�=��4eJ�w^�)����a
���@+�"�O��cOA�(v��J�óM��](yIr�5g B����`����L�$o9�8M��5gj��3�����r��tq�8M��Q�yV��h~��Q�q>av�R����\ǜ�,V���g�zV�'�!`p�nC$��$K$��FB�hR��ٍ�A�˴Y����Y
��x)�r�x.�E�.gR�G�kH��ܾaj\q]�l	�)2��7?�}m��ƼE�f��$�����7{LV9���7٘ݴ�@�M�����1���5���F>UD���&��D�u�ɖ����<f�Ďb:`��͖"���ĔQ��Zڸܭ�wLI=[�r�F�������Z���Z����xw��J��
TA�U�}���ѴA�D�gN��ۥ�|�-���1�5e�vz��b��A믐���ͣ9��c�5�� �a&�#UwoZ�)�dQh�Ώ��s��p�D�
@~������jۂ!�D����N�c�v����M~���7�X쉼4$lF�5�2���f� �OQ���G�$�O�[)8�3�dA���n&x���8��Y������.�7��D��B���.�W�j�~ݚ� %w�
[8���)��qA����o���^�w�a4M��"��6փ|��I�K�b�X��~O���������-��t#��#�>���A�'h4�Χ��������G�n���S�aF���.�p�yk���dF 0eQ�����G�N:;�lO�S��2 �/��;Pi��kM�����R���B���PEº�W�5b�P~�!ɼj��(�M�,�.���廲Ҽ�F�s�����+�Q&X3��%D���T�Z��J�������2Y��a�X�uF�f���rbi��~���=��J��en�
?o˹�+�Cu�y�����lj�n�~@�̀��5'�����볙H����h��oy�Wy���LND;�e��$��D�[6YԸ�A,�PP1o��Q���tV(��=����C���5��h�o��Wڸ܊�Se!��?�����/uk�t�O��Ĩ�8w9��u/Ai���жWl��*��!�&d�˓�n�T�^��87��`�*Q�0��љy��L��E�YL�h��XS9�S#�^T����ǩ�$��0�Ȕr`�c�B4��o��=�'��υ����9��ZM��!���'�t�4gړ�ٱ�;?�T@q2�3����4dؤ��7�bE*�Vu�Ko3�4�ay4%W�����T2��R�ªV�L�qN���+������u/������J�k!w� �N����e[`	��c�[�S�#�59'�0j)�j�T�<���s��M;
����{?:��i��E+����76)�B0_�%X�Qz����9���=����w�b�ǒI�IFT����%�J�0��f�a�V-�hB���Q�tk�*����k���-�XUss� ڧ� XuzK�K39��;N[_�f���]B�5�R(@O�IU��	W_��_ô��+yVf�T�hU�u`��o�S�������i��Yr&���q-GHf��3$�h��	M��[3�#��)��q�gi!%7,Px��٬Is/��uD�ǿ�:2��f�������,ǀ���i tß��-rE��O�F�N�*߅�6 �}4!PDf�����Ѣ����Q�c_��w���Z��*wWI�8���G�w?�Ε�=���N3�HX�����'�X���Y��Ry> p�Q ����'踑L����׽�����,��w��`�D�H[a�Wuz�x�	�A��#(�T�[S�˧��YtF�$w����{m?���u�'��;'S+B�62�=��M�&�-ک�ֈ4m��V����+��SN���7��G�FkR�l��`���������O�,�у�1�;=i�7r�*���ެ:H�@��D��0��Dt��İ�:gq��h������%�l�A�̨$�!X1�+$�I�h��ɜA�9�⟓����&�G�[��>��ZB�D�v��)­f�T���U��B�w0cb;��t�H�� ���#x0�3>[�ҷ���۸;5��T�,xA.���KzΩ���]�d5� S]�zD�!µ&:��4/���3$�Ԧ����p���@TX�ao64�)SjCek�I�����?���r�W���*$�u�(��+�cx[��sgF |#)���N���ޡ�3�S �2�H������I����[���#���g�uIzOg�#�wrC��~�@.i��=��oU0�f��#�<:' d��o������Qc�r��$"i&�h򍙈Z��р`7=�����#�Cޣ󄓹�r0��bj�I4A��ҖB�]c�\}qV�(�`ɫ�"�C�rt�ޯQ(o�S���^0=A��R_����	`
��
�����.��d;'����V���u�=L�J��t�L�OXȄb;�^ �Hd	�D$�t�[����hsxH-;Q�A���\�դi���hٻK�0Ʈ���aO��g���K:�瞽�D%t��iU�Β�&6��c(\GiG���#:}���G����c�WWW%�����މ	aA\��n�Ԭ4 �	-;�)��
��ۮ/D8T ��J�-���Ix�e��3q��o�m
g�ʍ�5��Z0Jh��i���UشQp���^1nc�j<�cw&�i$	c�1XD�d��L�;�P�w�@Jp�]p!t��FCt%�j���ߔ�����׋���!k�ά6������
L�R����)��E���C����Jq��/h&�5Z0x5S,���3ۣ��{~H�� w�|�b�-��g�N�I܃e��E�/�#Jg�9WI|��1[2��n��2�O��� 
ߎQW��m�/�q0�|m��Τ@�P���-U-Į��6�`�煓R	�z1�Z�rǍ��3%��.�.���О ���G�`�a���-�6W���+����!���
�]�Æ��{�B���VEiEpcpI��c�I��]�z3�����Ҷj��q�5��l>"�~<ik�2Hh~���J�k�ŦGa�*�Me�#R�K�/�->����A�2�b-��h�y��'<#���/'��:A�ԑ��Vߵ���2��P�>i�%x���kO�-�с�URt�1�By������/��Db��@�*����)��Ě̖9h#�.8�-���X��yu�?�:U!�X�[{�|����E�3ى�Ls�P���{�JD����C�f%���j��SnqfP���$&	�_]�d��|��xƟ��E}��s�ˢbA�n\0�o�rb����XR�Za���J$�f�OV�7@��Q���ƴ?o����L**\u�>7]��ݍg�Bj7W4�d����h�[�`�ⓜ�9�iI���9�8A�;��������:�](�1{�q������E����X�uu):�[�z��K�/��c �ᑭm�W����@��(�
aT6��n�;{̢���CpF�s���%0]��c��{$;�mI
��HD�g����(��1�P�C�V/�^�6M��@�;�_c7�F��iLH�F�"�� �����������������6nHa@������y�I I�n���Q��tM�+�rK��&�;/�]懡�+���������֖�`·��I��9��P�ݪ��$��ݫ`oS�騛�n#�	M�]R�s���1����#�me��UQ�.K�~1�3ا�:�|�	��A�
_:�R��ࢽ	��aK�L�o������~sx]8R�S�
H(��;�j�Y�J�Q.�nEs�u�iz�y�W|׽��Y�=2B/V#k��p�˶�,�����2z֧��s�N[׫�7J�{r{��#� �p�,��"4�tn`(��n�}?2'p��O�������O���PN��9[N% C�_�x�T:�t����`ei��T=\�q�^� �{~����m�/����f����ۨ�ߏ�:S,��&i�*p �8j�ʉJ��e��UӨ����ݧN��?�'afr`�7<ν��E�������cy��
Z�E%%0�_o�b���Y�"���ah.���؎џ3$��澱o"���}#�c���a��{�@������[9���-L4l�]c@�i�P����<�I~t�2�E%��9��B;�O@loR���n
�9g屷:h$��[��!qYf7��-X#�����$r"<��\7�i�Ck�Td���ղ�,��Ora:Iw@�m��Y7.I7�2�P@���'	HV8+-¢��Z[��t�f�6�#���k��w�$/"�t���ÿs���W�\z<>L�e%��r�U8N��n-��{�	�+9�|��m����yK�3��E>�sr���I��:3�82�&� K�6��-8P�b���v[@
��������5wIB��$�p�A��]F��Gw���� �}�L�H���N������-�䯽xu�n�j/p���`�!�*�14�� ����.z�N�Tڋ�^EN?��G�����rK<��F(;奋w��ƈi���(�֡���c:����Q��`;��I�o<Rb):{�8�ݽ׊��w%lWl��mW�	?�U;������G�^�� ����v��e#V�a'�hV&2#�`���s��>�u�c�;+����8�p��Q��=��}]�c��Q�꜍UotT�����S��ߠcf�z|j]sr^be=>k9=���>����	8��y	������+@]	�sqQk���W8�t�[��8gz�a�����Rp�\d�S��������1��˅�m}��ߟ.D5E;0�sύ��Epdj�V�¹�lB�6���s_����%P��4*�+���#p2��ڪ���	I�$)N�#}f5�D�z$p_�����="�,[2�ثY��>���u�˧ۯ�5�d��-���#A��$(��
�T.ƫ��j�{�5�_�e���n�AOi�8��GP �"]�Hͯ���ٮ�%�7LT4d��SX6N漛��yR����<����|6���P��$�ZsB�lr�_�����$/�m���	���0�7e��W��y�Z�dQ�f�YǍ����Hm�A#?_��iS��5�:U��x�.be~q�wI�=�_nQ$r��-B��H2��D�\�w�@7�Q�J�Ӷ�qnl�z�f�
s�k����rM�D��]�6^��
�<�3�D���it)�3�h��G��ꑺ>~�g�^�&�b�~
Ҽ�4 �wtg��!,q��o�b�ٻFR�	0����+O�,�C���a7�6}y��k��u�ђ�kI�B�^2@8���f�Y�EE��xS��l	8xU
��٠��_}a�u�JӪ	m+����f��.Q>2qfna+D��欪������Pj���8��w2yP<K}ȁ���Ez��{�$��������w}omI�v�A�f�t-�x(�l\j*��P'�)f`��ls���Pp�}����`�b����ɍ]h>ǩ�+j%�A��-��4��#�����p��R�~h�ٸ��D*]���}�z���
Y�ٲ�{�a ��v��ݻ������P����Y�͊18!����I�FR��� �DN���`2�m�I��1�^#�Cʣ;��
lUG��r]��+��yx�hw�>������ۊI��=�wI�{?��$�Z��t|wU�?P�h��f� ���c�R��=��H`$c�������,bvT���OC6ԩ|d�ϰ�#Q�*�ȿR��u�B�����mY?n���äj[�UՑW��#ģ�6ju'I��\g�Fo�4"��zA.��m��8빅�|��{�6FhHޟ�f1���W�v������4g� ���w�����?.R���K���=Bţo(ڏ����PO�P3'釆�6e��)�W�9Zwh�����f����0�S�X�|�IZ�z�v~e!B�[�b�O�� �r���WY�&,����	ll_�����m�;Lۂ/��i�ʜ��r�9��*@3���)���@��R��)܊7���A�A��å(^S��\6�f��2^L_e�LQ��F_bT-{Erf��2�����0��q��Ɓ����-���_�q��ꎿ83�ImT�q���`���-j~�|�eVV�3p���L��7�w!<�c_����;t1�+���h3CD^�ǩ�ؒ���SEb�f߃.-[Ӊ������@�Q����7�pԾZ�mqI�t�|�Y��)^@u�6P�;WN^�v�`��k��Y�ZF.���f?��BPg�ު�8�_<2�Y�ZC��γ�33[�,$�Y4���oJ�(��)��ͮȸf��?S��N�Κ�"�.q�c�E/F�����֡&Ԋ1���,�V�M(߻�~�΄��������X�A�~�ƕٸ��U1��ͥ��t�S�9�'�X�++�*"��P����;�T��X:��N���4��������{�+�9'o�!�k!�,E��0�:���य़A-KV:?��r�z����r�Pw@@���a������}����y�;�X��޽iɓwC3�)-_|�O�*����.��$d�-4�ԣ��~M��giگ�%�R����Y�i��iЃ�'סC�<���&�nfJ���V��} ����	y�E�Iϋ~���B����Ȃ�
U�v�;��&u��F���F�4��GT��Ɣ���L���@����J{�[p�҄�ʲJ�۷G��UC �������8i\�r-��.&8��%�N���gN����w�ǂ�.Y��2U9��@��.�E�>�!�0�=���l���Z�ނ����T��G׮��sf��7E�Y��i�)�]����2Rs�7a��%��1&�Q\�0ȕ{®��"3�;v����[��䀹윍�ˏơ&�Rvd�xt�cL��W�iA������&��X g�7��IoW�B���lH6S	�0�����t��C��n��CoWOn���r�H˶, )��D�v�Ɣ�)�yE��G��$
S�P��#:<��ʌ��-�¤��yJ���|ɲ���~�Y�;0^L]�R�A��������z6gú�I�Vq�����UWr�J��d㎑��Yl@����]�]��xm�]�w$;f�C�D�N���;�^�lB>�z�}�;�f	�8bP�!x}�a���{�B���~'�/�w׿�O�z��8Pk\�&.�$��WN8���	��!H8�N����'N��պ���~2p��!-[dCZ�!�B���Jn�,ީ��g��q�U�ï�@��&�m���`|�J�O�l�Y�r�q��;��,}|��πXb�����$�g��{�����f�x�wCo�&P�A�:Fě�PL?{��ڹ|eԕ�G�^����^��ZN�����x5��r�< .��`^��m@غ��MZ�-�;��2�����)�c�e`q���J���Iu�S��.cU�=����F��_r�u��>�����Ĥ6������9��|�N|t%n���(k�G��,�hv��@S�~��T)2�!`ɫMYshY#I�wRWOY�
��m.����R�R,ɹ1W�!�d��^J���Ė)�쩈��ns�"0�fQ� �E�Ԝ�ys?��yD~=D��b��4,�o����h�Uh�pU;֭���ȫv,�ƠY��:�Ej�P<���s��13q�1�ǹ�RyUy 5�TÖ���W5�Aq
a�7�;r�mq�������7��
�Sλ0p�zZ!�]H���bHl����Wnx�Y�����9�/v�"v�F�@v՘���+	��D�:��J=q��~I5�g`(�Wwt���O8��:�a�z�y��J���ԡ�� ���kן,+�_Y�vPT $?�LS����b�e2=�T��Ѻ������K�cu�"f����E�W����2�&�Ȋ��Һ�5 |��,��Gg�'�]"�X�6�n�K(s�CU��l���S|R�[�ɬo�)ԓ{,x� ��%6X��eN�/)�E+s�����1Jt?A]P*l��/�mj�� f�	��	��J�G�g�P���������V��Zd��=��0�l^�ϖbG���B��£��F�ϼ�f4$w�+�>�$�����Cx^�bT��މ^s%"����-�b�����y��Ij�I�������'��?C��`"D�QKf"j��Pսzf��1�[N�?fB��e��⎙��elQ��"��O��}QKg�jw3������^۲̷�!6K���	"V�6�W��1�7��wk�z�n��=i�000 �gT�sR�j��;�_��J�*`�6�zR�I��
X,3�M�6���%v?����
8*�6��0�nAB����_�$�6�w���e������s�h��Q9��E�#��#�`���x�8`hJ⦸JY/�J�΍A�P�kf-�W�2�r]EI��F�WH~�E��t�dڡ�-�U1Ԍ|�� �p�%Y�ٗb�ϩN�H%tɣ�����:g|�q7��70�Ulg�ʹS
��x�w��,�9���Юs���"^{�&�Z[���l ��j�@#F��f�$Z�\N����(��#!�V��%8�^(|# �7k�15��*���͹K� H~��uE���]W����G?�)kn"aG�o�쮩dz�m^���WP���u�l�� �&$��y�G����j_��H����'��׻�u�)�-w��u���p�Qv�aG�%iWM�LMF�n�?Kiͤ>�z,J�E��ظ�(��:�����Ϻ�y������l�ah�'�������վG�;�Ii
�<��v_�b;��[t� K�����\�/�6�<��_��q��jI�P�&��kj'�5��Q�N�A��_�$� zIN L�^9
�K��qr�?啝揦C���
	p�=񯼷L�uJC��}�E������1K��;
Z�߅���c�*�^s�2�P~�%^گ�J`I9]TF֒aKl]0c����͙@�E�Co�BY�,]��lG�V'��Xj�ڂ�6��Ifv�*�r���~��5Wу�)��"��-�XZ�������(
�������M��g��R�ւ�����y^`5l�>�\�Q��1�V�PM�E.^��)D��������;�4}�1���nH��mf�|�2�5���I`m:��)�֙}�ާ�B�pxK*�ƪ6jG'�P�k.;�iɭ�f�p���Z�A �������ռ�f������뗩[�����V�=�9˂�y���d9�i�y��h��v�-v���Оuv�Ϸ[������A$
t	��|�_�P�⪒�~��1 =��0kZ�JGF��\(_ttΒ>X�=$�b��Q�B�;f?-��A|F!ڹ��Ё?x���um�b#���F����n���6s����o�4�梛�w�}�M�
��/b����V�������an|".�1��;0�#�~p�4�p��Y϶D]+��_����I�KQ�#� ���"΀4� ��k X���o%��i���f�l�X礽�;7ü�5Mޢ���}�4C$|����k`C���O�w��g ���F �$V�
�ќ�Ų��Ka?��{(�t!Qz,��AhܦEԦ�$�ѳd��4��kl��L|<(�Ly����VQTΤx���ߔ���+��<E�>w�:R�<��y�6��N"X��iߴ��[�L� z�2�jɽ+^}�i����]+�~�b�T�8��d���n�N�Uo���ǚ�d�)h+.�2`��������R�nxMY���5�Z�U�6Q Rȳj�"B��+���U_��K>C��`������i�:��Y3�},$�9*|tL��]7���_�{(�w�f}�~@����u����#l������Q�Ͽ��-=9�.]�����\��]��G����@[#���M�[~s��W�|�����\�`���DF�pBTILϒ̶~�Y[�ΔU���2��7�l� V�l&���96A��Eԡ���lV���,�vf�!�FL:�;�a���3S.�r�{�?~}��?������BS?KV�z���w�ӭb��L���UZ~��Sba#}��o�{P��#��ξrm۰0�r�e�Yt�
w��ّΑD�u1�̋��`��H�n�{�?�@����ԓX;�HX�Km.`�R�YbGo�r�Az�{��_U��nHt�F���9�9;��e�{��0ˌ!��������'maCR�[�-��_�!#A̘[2GXk}17�VaqQ�N�����\	�v/G�@ŸL�î�2�Tg�ɘע��O�n�w�..��?@@'h�6a���|��p>�Oǣ�ɕq��c�,%8�bm���D�J¢�Ie��-=s�~vy.5L&�J��j�K< ���г��ց/��N��f=z�Y�����0~������g8�DJb����CE�|�Ƽ��ǵ=ެ��]w-\��ç��;ȹ����b-n���zH�H�kǽ���!x��*́Ec,�x�$��sW���t���GY`�̀�I��8���%���"�/,���:)?���]�k����6�n��.t�$t~]�0Ӣ�~�"�4�	a��9Tr��=My���X#z��N��W�{�5/��x�k����ɖ�Rv��H��m�?�!)<xS��Mq�`I��?�1O"*wF͔'zh�l��v8.՚��h()3��+��!#M_H̿���/b�L���@��]��i��B^<j	I��j!�.PF& +���|<.,�H#�wq�%��&�A�����8�&K(1y~��57`�O�0TNt��)�|�yB�/�J��_�'�����=�g�ؾ��M�X!�:�QJ�?[���-���Y���
��j8;v��g�v����>�x�`?��[Zo�s=SȔ(P���g$Ԍ3˲
Y6�R�g�d�9�Q>W������9��(j�y���[�:�im:����P�{P��ڇJ	�n�xu�c��'��6]�5����R��#-A;iu��7M&}�Y5؆kT�d��0��?3�G�v��W�&Ee��@���`�A���>�� �Ձ��(�T�Ғܩ\|�_�%3b��T-ɦ'��H�X�I�<�6��e�ɢ5sv^�E�_M�MQ��"���	;C�N$E �����p���F��|�i,!+�2�� ����\�
9Y��.V	H\L�	hcp/�\���9(N۪*���~�)�
֢q��|\�P��3�|����������g�9	jOo�����~;�`�tNQ+
E��A�?Y��P������p'-��z\��1djQ�fv�@�D�z,fj0�@J?h��b��L�T�Ű�3k����uc
4�a���q�a�s��v���@�aH��i.�h(Wu���/�#чa����O���P���Πk�߸$���cԮ3D�l�#\u���g(NQj���{�C��n����yͲ�`2oIS`�Rs�HW���V����٭w+B�o�����I��xh���pn����iUh�)q>��l��{D�x=�/�T��?�o�y���>/���_�o��	��za�B�����>#����0)w��Q���^��v�=d�����q��g�i��Q��z$��&���*�79);��bu[�μ�!��ƍLʭ�&�dð�K�����~@�,ix �Fc-�9GS�, ]m�f�e;��4j��9�p��H��ic߼�UE���蚸���L5��~=�y�O����ہP�����o\�Cz������H�%��"kux�/G�xBdv%2��
���
���$y|�J��|Py�TK��{�·��"L��购���wW����,�`a���`=���'ʮ`�H !���xR���� #��j4㝇�0����L<o��',�י��uo�B�l�h$r�<RL2)��_��N�/�DHڋи@tB��}�4Aj# �EY
�VwIY�!�Κ~1���a}[Q���u��3W����Ӝ�4���y��é��MݤQ�\��C�Afd���A�y��<�66���}-�m>�C�ܶ�PIs��&n:�8/��,�0/�k
��=�?���sAO�>�"l~;��Ҕ25���憗�8m|��"�Y	�>}����j+�v�@�?����i��>z�B�w�o$ʌۙ呬�r?(,�����O4������]��[�&��|T�4m�gt1\�b�3��<�́S4d�%�Ԛ�W�M'����Z%/'�#����9��?�h���^����\D�������c�0y����~��ױ���똶Z2�����}�c,�\m9��@���N���
#}����р�w�6~>(d�6$C�|T���P�x�p�ֈ��V�RZ]����B�|��AXf�<3e�������1��N�\ӭ<�����mjp���Nu�s��-�Q��=�is,LH��V"�*�(���_�
̢�/��I[K�b�B����/C8.}rT_&��}����6*�e�&�\۔�uP5����
��u@�u�}w��ܶ�;q�g��v2%A}�A4�a���h��0����t$�����	(���3��� �����3?v� ��Ev�|�7 )� �<�L��w�.���lq	T�-����k5YN=��6�Il[��U¯��e���	m�	�J�r��Q��Ό����bg�y��h@�0~��D��(�
4h�B�n�Vؖ�Z�b8>����Nh.��M�H#S����v#�5��ø�G3)h�ί�M��$� b��?j��[CXn4j.�R����.7fVď�
ҡ�Y�|�Jil�i��<:�����E����%��$	��,)*ް��\С�äǐ��Ҧa`��7��Nx $��wJ>�mKh��n�oz������6r�F�Y{?��@��(�r���꿈MP;(]�ڔ��Bl-��س��q
-�ix��A|�˽|16,������_"��F�l����5 �&�d=#��o�ц7[��
���K-��`�͢4-����]6Oz/��8#@.�@_�zW�P�j'�&48A@e �=���ɊBĊ���f2c�S���1���I߷k&���=���7I�i�!9�֛��cT�s�z�+�x׌�M9
/(�@�K���z�Ϸ�j�QsU��M�Y�0��7\�Ќb$����i����9�j��/����A�|���"���LpG0H*�s�Bd'�3b�t��h�|y�.��'�>t#ҷO�g퉡H~��9I��"��#�UhC��u����m����.��Y?�=�6\{j�C��%'�O�H�c��=��B��z�KJ
>���M\t�@�$p?��	m1UYc��e�V�L��ɺ�y7�~^�����I��Ts��wIy��r�Xw��%��j��}	4V`���SsA��p627삆�8���F��Ia'L6~N����
�-��#��~�&=zVb�Sԉ�� X���°>MPs?����\B����h��T.�����
P����$z��";A����9�uv}���?�e�.C��������碛B9�ak���Vѿh	���;��ʇ�ݗ&�'L��19�b��J�Y�=�ᄽU�Fgb�fL*�٘6˛�6W�@�7c+��݉f]d��&�m{�.4���[��꼛�U��A��'�������Y�l��m��{��E���\~�8�|������1_�K|�/�FX�'�����#/p;�/[��1'@�#b�t(Qc�Iu�|(�4�2��_ZM�Z6�\�%L����R�����9X�[�����;�r���j>��������Tp�����A��ۄ�0,&!:������b�� ������T#i�%�h��M���R9�F ���}�1Zӫ��o����"��XC�ko� �lW`X��Pv�J.�hA�R�}L���Y�j�P�;:nXFT�Y����c;�Y���7,z� �Vz;(����Ȭ1zjт��9���0�	�-�)׹���Z��/�E�����~دR-'�A߂����
Ɲ{�z"�w��x2��y����iի-�	;������'Ս&o �hm���������q������~�H�7{VH<->CЦ/��S�^�di��y����{%H����`=SH tDhwYDQ:m��{�Ӎ��H=����FX!��#��Ww�;���Q�q�;aCz��3��4Oh�}bN���F��l���ۂz���rZ��"V�s #�@,Hj
�J�-�̪���-]���%g�4�E�:5���<SN��{�c���aLz-�;���#��� L��|��X��u����gk��3}�
a��5M����nv�_�o�T���B3k�3��ķ���/ST�])�(�t]s�u]�z�s٠�W�+ʲQY�
�4��GU�����I�ţr��������K�0�7�h��ք�F\=k޵�I9�wzA* �����({��e�����jTZTA�hz�=�K�s�@l������\�C�ۆ[a�n:�Je�t8R��wW�W,�up�a}\}�P�v�ro�У�Ƀ��NV�;��9M�U�� ����45��Yb�����w����[��B�ʴ^˨ȅTX�Mx���+_�=e&̗!��q:���ਝ{����=��IFyp�f�Q��N�_���V�f�E�6�*0ұ�g3Ѩ�$	������k+�1�×6�p�+����C'5N���&���.fA��gIB<k���-`}�t^2 ���Z�,
}M����}Gsԯ�s��㐅��ٓR�g֥�Κ{��z(=���&|/�����X�pS�@q��_���$���n�E�ҧ�|t	��.䵮\H��EU���ԁN�9�ff/�?���>I�>��@!��
����T�C�ψ��ї|�ɴ�!E�X�
|���ե~��(��
�Ŝ�zv${�������
ykk�H��
���jP����S�"�H�zR�w���Ǩ֨�)�����l���E�gnϪ<���s	,���lO#��(���;��{{��-I
�� {g��'W���l��f����bN̅-�X��j�-L�0���%\���$�S�	�Zb�/q���+�/����n��ϵQn/���uٸ�|)U�
�&fP�S�>��T:Ȳ4���4;[�xL�����/V˔�� ���V�A���<Z{�̨�	�έ1�᩾N*���U��j+������k�So8�BV��	$��������6�d��U�ǉ�B����߯��?i�7�k������0!�{j����iT��сh�!H�#g��uܩU�>ϩ�L���p����>&kʹ=1�zm�)Ifw���J]���x����<t3�c$��X�9�Q��x�G����Z�6	��W�������V������ؚU����p�g=0!ԅeR�K�Hxgg�f��	��C~�w��LRV�H���z�:A2�
�Le�;͓x�\ˏ�Ib�/�ح}I�iu���mI-�8,�R(�}q-d�G��n�1�P�]��z�߮U���컷8�B0�6�x2�?�[F'=pC��t�#^�G_��a�]=�S�|������yV7�op���M\�ɶ�8Æe�I�홄�e{	;���-���n	aS,���w�yIG�7�͋��H&i�n�i�{o#j���-��k�n���fx�A5of�K"0�:�ȅA��	v�d��N��Y&=Ј�M����!_u��/vV��4�d� |�k2���]�����C!��W�9QQ��Ƿ�P���Sz��Ƞ����l"�H���lN8�n�m�s�	p�Lsx�O龌G���U5)z�#��(����ݙ�b@�9�����01:�J!���a� �Vu��M���0O�1����z��$�-(�k�Q��;Qj�Y��ITt��iX�NP!j5�&77E]g��3��|�#�.ɗ���v�; �����',X�5�wG�k�fg�U�`8�JK��эmA~��	S�.k�06���{}��S��h�=�!�y�ۜ�Vצ�.5�Z*�cup�qq�m��2)�t�_7�S������K��t\�=��5���E����o�e_��tp�79����Z���$T))�n�����RᱳX(��ee(#!4�G 3W@�'�Y�}��Z$l�!���at��͟"p�l٪��5G�iD���!�ۿ�c؎l� r�"\K�)7#E��F;��m�q
�,Ai���Zz��VFp'��\֨�Ks<mW�΍���1��0GpV���'�yI����)������D�D��P��b�SKk�mT�O�� ��\�,��й,B���Zc�'�U�QL���׫�i�HxY�!̦�:p�@Q��A�B�3ۓ����`��V�Wǃ��K�-Y��M�� ��/�������{��#��|�������X�Ws�M���Ym�wj�G*nLr��0+����CrJuRs�h^�u3�Km�}���#N��`��g�X>ˈ�A�
�E�4��	�86�Í6gp�����HJW��M��}�ܨ2���Ҥk��T7�3S�z6� R.;���o̖s�,��{�$ BJ�c-�B�t�Y�7��$.�� �Z�fD������,Ț�����L׫��GS2u3��O0�7�#p\�K��;��]��eh��p��&�)͒�P fYu�+*6���5w��${�Q�#�͜w��;�JC�R#��t�8�����`��b���3�jw�t�0D Yɱw���R�"�m�J8{_0��6��l�ΙWqS�B�㙎nF���2k���D�.oP@U�J��k�*�{��z,9��t:�u�^Էb����GI�k�2��+���!��? �1�̛\l&:�uP�9����H�م.Q)�Xs��4��'F����UAK�H1!X ���aϻ0��|b�·���x�]�Y����Ԁ|�-�Ź*ҝ�p]�d�H����mL*@��m$���.1r 5���0h��C2�z1�-6�z�8�)xpI����R5A�%y��ĦoH���)�C0x�2CO�N���<t��K%�K}�&�7����ѮI���5��|z��&�{��ޑ����`v�`��R�4���&�%vⳏ;x
s�9Uc3���@���ۉ��{y��S�4����m#�+�~�U�����gz���+��]����E���2\���ʆ� ��e�r����o�:�֘/)y�A/�ˠ�gD��p�M^S&�Nв��ЂP�i��|T��������JR�[߼�p|=�z.e���T���Æ��LVS,��K4���	Qj~W�@a�Pv��������k�[q�:ۜ�5{���ɪ�� "�3�
��)����V �V�'kJ�=���u� 0�[���������s���ys�CQ.��?���9�C �P`uZ1��/��-��e��T��!ZH�w�lY�bZL��>�e�u��Ϲ�.z{�
G�饮qi��0�m�l�M���w)��k��a�}C;�UV~�� �pZ�P��9}�M���:�U�i��En	�'��q�� A���g1�U�Z�`Fb$T�Â��(B�8�C^7��<�_6�Q����Ɗg\o�S�3�(��$�<ԏ�}�H�<����u�NLT�d�(��]K�45�#���
��$S'����|�T�Eԋ9�e��c��}���+l^n�L�6�YRp;Vǒ��{�J1��'Bl�E$@��l"ܿ9V��F֟P����Dk������`��ُ�סk�ӻ����&E�K��gz8эp��>No����/��֓s���*2(�Vo�,�OȽ_%���eZ�
��󔠪���X���iB�5�<��KÚi
�����	� )���0���@�pD�dS��O�"{�2{�3߭���Ds��{_���ڽ�&?�_G!7�ޣ-�{Cвy��BhJy�$�j����v�+֣B���D_�E�~�j�q���GL˭du;?�I��g\h�@����%�����i11����]8(4���M�&��-q΍��bo����0 	Q,\��c�d�fZ�*�_�ݐV�&�]��f�(X~]��-�W�wͲ��d�x�r��v��Ԋ������)$B�Ç �i8��Q������{h����
Q�� BM<쐻�'��(��c�]>s�0��+Gw���=��P�}��+�O�K�cn�c����n7%n�Ő7�7L˿p#l"%�z��x��PR��F@�	Y�O�Ql{I���- C������k��5V3
�;e_� ؊$��q�2	��D���04�ȷ�>�3p���f���t�����(&��@��
K��_��E���V����Q���x��޳��%�h��a�B!o�����h@勪ncq��Aa�;������=L�B[�"Y����|1�(������fH���~~��:���;-
�={<���#�m�u����L#9�>?Şr������$��
�+ "�ľ���J�i����P�ś4jP�L�g8_W?�wpS������B��Yx�j��W:^�Xж�y�(�����`�5{�3����J�D�*{��#u�ln��N?��?�1��"�E����tF�]fל��NLx�0e�K�����J�[��T��\Ԃ�H�F���/w��)#�_3�l�v�%��xN ic�OM?��T�t�
	J]L��V�+A�H����k��;�oy��SC�i��S����$L��<{z`�=nB�:��z�'�۱�����	c`I�������e*v��R��E�T�[-�]�#����#��qJZ|d�.Ӕ�Tgj=oK�V�Cc�\],Q��Ug�]Y�ۘ��7#���$$���*�0��e��@Y|.�R�w�����k{�������U1��V]V7z L�	Y����={KMZ-��f�����ϵv������ծ8e�����_�Y�3^���k�:��H�%Yc:@�W~�ͅ)b�t�M�+%>��Ƽ�7,���塝y�Z��=a��v���1ϛ[8?�A����n��*���*G5eH{�p�}�q�Z�����a����1�-���ϳ <;[,��z�á���)�{1h��c��li��]J�����`��<�=�[p��Jƛ�!���ͳ@�ؕ�v.����Z�?��X�n�t�����vy!�t �QQ���gj�ˠ}�w@_�?c����3���ݧD�x`�U4�|���6����G��{�nNt!a�8�u!�K?�R�c�F�&��Y\��,�k� KM�}1,'OUR�ư�ې�����5!�"Ɯ;���Ti	;)�3�G�#<��"ش@\ږV�ޥ���׍%8ػ�ڜ:K,OFq���5��3O7��7�� rY��4D
4f�tN��{��Up1Zڼ�oe�}v����-�n��K�hE|#������Qq�*Y�g.�I�Z���`t�W@������c9�gt�8Y/yj�b#W�Íde����cǷ1i�k�6�I�����یC�?�+R8��%���׃�W�{F����UO��GG�+p��w���/�o^V������!Ml�:���z�ݼ���m<}wH�|� ����U�q�j�-�X�Ԇkq�c߉�[�	��%�?�?)ϻ��%%#U�eOzI�Z��oT�W�Wx��oS����6̻�k��O�چ�&����\v��0��־�vV�1��8�CԌ�ӎi6��3��r�\�l��4���>�[��	:��j*�N��p\��2�]�M�l�L�����8�e��0Mj�c <�uE�Q�bZu�p��U8b�-�滘|[^C���j���\���ӣdQ�4���N�ld���v��a��:�.`��$CK�`7��ِ�1_�ǒ�k�.��C̑�j6I����Ϙ�c�R�߯ݵc�/���#����Jtx8M��a*r�x����GhU)j6l��'���i�P�
�8<��y�x_:whH����pIN�Q��S�U�	GĵO��՝G2���`j���/k��)�{�B����	b�BƜ4��-�ZU�����;lf�S4�c� *N�y�w�?�i�Ztť���B���<0�5a�qL��3��)/���JQ/O�[�< &�y�HР��hȣe;� m*8��>fo��ƴ:y�+$�,����P�ن]4s(_;�
�雥V\�nݾ(84��`m�N���\�AK�OC%5a�����.���q���9��d�~Ii��	�@'��[o)|Oճ�!-w�]'��;��?!+*Z�-d=�VT�|��#��x���,ډ8�Q��dK�eVK��Yʖ�+%�f_����$��}�wD(�@I�L�n3֑�X|Z��%�p���e�ĉ���/�����i�Y8��6P���0���8ٔJ�F��m��/��8rP�7~��DEtIg�f�{���7�-Q��X�.�}8&hϪ�v���@�˷j}vQZS%rRpdsʒ�k����i����.+�ng3X�
��9���+cԳ��6#.)1�B`�麻��(յ���[҃�)�e�b�xu� l#O�d��Q�ۼփ0�v��B5�,Y �C�fV,Ŋ��гi3q6l,E�&<�ܐ⳸�Q<��!�	s�ډv��4�&�!	��	��km�\�hh�To��*�x���k��≷��yo6Y�83�� hY*��z���@s�nਵ�I>�2,}���n����_쏻���Y�t��uF� �߱�&��D�R!��8G~�uw�Pû�<�(w�k��t,&�CR'�	Z�j�����mY����2L���Ml6���V?�� FhJ%*k��BKG�����K�"�=�ų��!�G֐b7�jf% �sQo&���w���:��~[X��-8�n3R���w�T���P��8���K��q��f�����S�����À�`O䑤,� �ϣ�M��rW$�}(В�p�C�O�;�+�b���<�,X����{e��
�PT�_�^�D��7F��/�����S@� Z'>���P;�B��L������PG��ٮ|$�\X5ə��Q�FXv�ׂӴ�ٮI�ѡ��N�,�d|Ae��/s�Y��*HL$�I]���[�Z�م�����r����_�.m���#�Ag㮴}���S�����n��t����
c9C���,��1>�:O���N��W������B ����f{ 3	�����D+�3뀟�X݉R/����Ч�� h�����a��O����&]Bt��VC�X�	tp1����6�	�{�ݗ��("�7����� <(�j�"��J�>߶/��[_S�L�:3g�%󧨲�yWo�&6:t�Б�0�9΢VM����m�p�ʅ{xz[��F�8Ά��&�=��HN�����/���fI@���<~Z��͍'��^��Q��"��;���ҕ`�"%��!�A�i4��o?0	<L̩�삙��7��$J���o]��B�������{x�4G]�C�N6��?VbY��BvNp'V�aE���Hj���~�q8�x��f�ؠ�9't��<��3Ƈd���Y�9$㱐=;�������ɔ�E�����@��Kx��_���h�3�6տ$�|Wk�H/[���Pxc���=tk��G���QIuQ���C�nr�Z��6�wT��SV��G��1mĩ#�_f'���c�%g�p4�&{`&�w@ �Z�y3^���K�^�̧�/�tS��K���|��rU�G(_ i�Y`�;@q(j�ga�o����t-���˫�|L\��б��׺�.oWT�L�R"�m���s�Z�M��?�e:lb�*.{���b��G�4݅�2��^�#���	��N�Xe�q�[5Pg�.�؍wI�ۙy��x�n'�|]�x�[���XH]�L�s=�+ P�]����D�&��K�hw5�-n� .�
�j>oQ��-E�����F�Í��u��[k�g-���-M#]Q/�	����QTH$�2J�o.��bm\U�QL����+��gw�����@���ä�p���[�Nq�T�	D�(׫mٸM Q��tZ��A,?�+|��q����Kۘ<n2/렪ʜƀ���ӡ 
�*�0�S��؟2��_	HT��	���"�Q@D�;�zs8`4�����.�m��6]��(S:� �8ɮ���& ��ڣ�P�Aù�"iY�T$��ghɢ�Շ�K)�t��@�	����q��-���κ�*�?�@c�9���w�Xv�a$�3�O#����|nɝ�����d�ۦAZ���jP
���Ύ�T��1T�L2�x+���\~^6&�m���-G�����e~�5��qh�� b�C8`A&�SE�������ٿj	�����Ō��������^�)%B;[C��F�uP�
�������~�+��=fT:y���x 'c���� B�	%|+	h%�����j̢]��n�5\�3��8�K��r�զPv�c��O��k�C���pd�b֧!���4X�<�nÔO�p�.vY����0Z��b^A'z��U|Z���*$O��J���v��a�k�S���/�V�t��qnX����Z��/ӄ��l�gp�D���@{��V'.Gh�|Ģ��EMv��Ftx��7#F�:_)躩q�Y�R�Ӡ�.q!l��;n^�Θ/���8�Ԉ�1P	�ü��0�<��vM�b��=�4<�݌'m[�^[�����W��p�Z\M�� ��^�,0�TWk��I�缉��!i6��Ɉ��͉�+���<��6��ƩZ=7��	��k�-��D��~8I�1*m�����
��TMb������9�nz��2��y�n UɁ��I_�8�$`r^e⫅����0Fʧ��Vp؞�?N��e{@��z�ZJ�
J��[2O�:=�9[��,ab�}D���|)�k�\�`�wi�#�[p{o<Qd��C0��]�B�+�3��~�BR�晕��c��>��3[S|G�V@'�[�]��=���,�bd�uM�S�ZF�� ƴ8�!�ƈ����X��Y�1p�k����KR#䤵���z$���-p�P��W�Kj�J���0����,Y]Q�Xݨ�Ώ��L��I��]����ٙd'�?��z�eUƙCг�iɊ�X�ka��4t�wL�4?)�{b4x<"!dVo�yo��o/���J0���`v�~��ȍ�E:�9�*OZ�� ��q<�i	�]���G/�CJ���IM���29�3�)F-@A�w�>�(�@�D�m���|5�3�,/[ԗ[oN����~��[#��v����2�G�/�J��џm�V�/����J+�����i�)�m��Vpq�LQ, �����qK�A��
v�e/�g�8	��<�
��7�6�@��&o���K�zg]��mch45NSa��R!�v�l��P���c���m��*	2��ǋ�Н<�q̈́�r�9���u0x���XCco6�����C�6�H��X"���K/�5��}u��Y�|r�F����:FX!NUȆ�wՄHP
'�-U��:}zy���r2p8�4�9fܤ�9�H�Q?�ft�p�Im�a�z�
)kc'i*���D��W�b!�<;� �x/��;y _[<�Y�lg���f�UK���{�Z��u"j�<�۲�� ���|��h�P�
_x���q˷a��`SV3�0��dq�ԩod��z�/5��3Q*�UI>zh�6�FA{�r�ҵHH�\�N�K�>�!lj��5�=&p�ؑ�������e�e}ho�$�0`�J�+���G=�.�ꤳi3ЂZ���$3$�!�W���}a0_�\�-�d����hJ�:1�%�d��ֶ�ȯ�cMtP�N�Z�60� n\����*��b��)���bC��y��l2�VT.�����UY��K`�&q�s��1|�l%��.BA�IB[@=D���$�!�3t�ˁ�i/{�%M�I�7���i
E���I�E�'\��!��\�����H�v?rWˍcV&ek'��o~j�y�"j'(7>�|r�N�^c|���`�	����mt�@�7{�3��o ��	�*'�wD��-ۦ[�s���CM�t�Y�d�#�W}�U42,�	d�o����:/���=�A��0P���a*hp���Nk��FX��%�,�����Cg�-Xi:��v��8ӾW�0s&������籰Y]^�ƃ~��8�6���%����@cJ� ��4�`"��.)�M~��̛����|�z_�?�B�#�P#[8�sp���w���c�TR}�PE��C8�L�cm��c���ʶ����68L�f�Oim�M��z O�����!9��;ѳ|�����޾5^GZ�L��vEP��RP[��V*��3ܰ'�3�j����2�|0�T�r�Q~ ��\�0ڳ{l��;ݡC�uvTE�"6�V��N�X$�2��D��������!�w��z�_.J���ֻ��xj@J��{e�vD�XОR�[�<�N>_u��c�^��:��
�0�H^R�-�&ph��D��[�6��t�ot�657��;���}��g�[*#W�S`n�y� &ݜ��3�Kp@�!�'��0�]���S���E]�k�Em�ɠt�DĕytJ�ZwfN٭�b���窶������/j�ـVd����C�'z!枽�.�E����l����y�Qe��?LH�]��{I�>���Bb��T�'c�����H��s)j�*b�[��i^F 7K�]˘���d�i9����c(~ ����[��(�.%��6X��8][A�ﴄ���,L��V7Ӵ�?�_efh֤[�9aSM��,��͔�
�Qk������e"n�*}��iY�q�x/�<�wB�J;a�T�c��SG��f�Ka��bMw�_�����_,�t&�aB� ��HغM�˂jOL՚�
���7�c�R�\�Sk�[��J�c"�Yև�x���Itl�����@NG#�i�\z
Z��53igI�^�����O��1UD�L{���KY�{���Q]d�s㼵�f�8�J��;RS���$����Ii�*�|�w`ڂ�VQrP�{��5�4�rH�DF�|v`a�u�����������z�K�YU_4���a�a�� �.9}�?+�E�J��[�f���`������|c����U�v� �`�e�#�$��祱�����6I����/�+�� l7�H�����ڝ;�������*0��>#�?l�"M�+�GtW�fz��2곙��K�-�hh�i�|x�y�r�S��quN�MH���@8�,*�ptY����?�Qu�qh��QK�Y�c�����<�`s����&U�
�s���1-56�pY}n�ݠ�~Uoi��I�9��.Z�e�.1�3�܎�i}���b�Ǝg۠ }LTR����
Md�6���k�J��+�E�Pt��	�z*�M4����ھ��SeԸyߗ�-F�H���E� !�����z�Ws?�!u�6;�F_F����k���a�RV�x ��gM:�+��C�@	e�o�������̬;�c�Ѕf+I�)�Q���P���A��Kus~�p��S~d<��.��HW�v�V'FT��][Q�8u��Xٖ�����z�e%.��Ff}�'�Ƙ��ս�3(�o�"����i����z0�-)"�Ǐ���R@c�iM�斡�@j`��j�A�{��f_�
����9 ���q��B�m�!����ц^k��\݈��|����04�ף/^��!�v�q=7��Ç���~Ux�
�XVb^nǐ���C�}��[�?��Y�+�Ib`sNgP)�]������ў���M5!��I4�<l�HiZN^����m�=�?��������gU���eU��-���}>e����i�V��a����M�'h����l��X,#H�I-d(��������]�K�N�Ĝ�Sx>hwR�[�g�2���տp!��҇Dw�K�*�&�4������PNq,�#y�|%�?O��4��Kp�e��'��܄ J�o�L|{{@i���oื*;�h�q�t��I>��寊fy56\����
��8�GE�h��!x���Ώ��Q����\=�0C�̲A�_,���~��z4��A�x����Cyْ���縒=/�8<4nR�n{M�:��
{�F; }�y';-�*��{^˗�(�-�	���bVJVV3L3 X��[=�Ra*'L���MϤ�]W����M���'�5�$�B�]X,as��|M��-��1R�����5-��	��b�����U��f"������6Ȇ���c�.�I��"�=q-�i�@ːS�tM��k*j|u��>�O�n÷-�gW����5����@��=��o����g難�)�������l�q;��1ƾq�nr��5R�n+��5c{�;`���bCϘ��`�p5��4:��������.�9�G_����TnRB�c2s��>ݾ�K�h�9���k�<�B��#1c��~J�1�0��~�"�`�2��1���i���}��뤯r�b�yJ��r�]��M
�_��獠��L^�{�ޘ)�S����"PƥV�\�d�8�YN���Ζ��賁� �:%��7��K��久v��C0c��0�Y���Z%� F"�6�m;S��U�O��A��Xf�U#�mn��CS��n�ټ:j�.œ�{�,�2j2(Z�R�ݬ84]�g������a�5�>T1���T��[q����/���R8�sN~/��e��&p�/�BR�r����`�ÉI�
�Uxb_I6�Ѩ��n=���{�v��f��l+1�ً��^gܝ�k����R"OQ�rX��<��c�6�L6{�Ė�Y 0�8(L-v�wA1ߓ��]�EW�/�󸄲�NGx\���2	�B�-#�W�q|q����op�/5�Tm�6�@�j��\�$<�J�5H�W]�+%(c2f�����?��u�n���0�;��G�Xf�F�$�f�SI��4�y{t�5���҃�O�аd�ȻOa��*���Of�Os�WY��T�j<c���	A�J��r(�^�8;N"i����&=��) Y�� �������65u,.Ct�(5/�������` �0m�+\ὃ����H�&^�<.f
�h�y����t�}:���E�uD��Nt�Uτ9G=Nw� Iܲ����n$}b�b1ə��@�{�+��_WC eR��0Y$��|���u�>�{�7.q?�ǯ�U����*��S�q{l����>��H�:�_��� 7�T4�@`�?�X/wh�K��ܛ��D�5��ŅM
qteϽ�¢Q�x�6c����w͑=S��fW]w�,Ii/+��FǺG�������c(�UY�<����P���a�\Ps���7�o>�]�<JE/O�T�V�C^%��d��Q�cp"���I!.eCW��1� �W�/��t���w�s�֟�������C�����,;�!�v{&	F�4�*b؈�g���)ۡ�)3�Ĉ��$����f]V��k� pl�4~$�@7D���O~tR�Ob���k��LpR�RL_��Q�Y~��_ˣI�x�D_��V[W� s���
l�����ZJO�o5�LK�, ��~4_��P6�n�E�	���t0�x�5%�7Ĺ��'1���dNM�#9�Лm�:Ee�{ �iA$��T!�4�|p�",�t��i�,1À���*�[���,.��tR��[>�b�
6��	����s�	�pp��Ĉ/	uU�3z���i_	�@9��|��{�$$�k��)�p[��)>�y��څh���5��% �&�@�Z��Xrm�S��_�H��'��o�:�pQ���>pyQ��e��m�Ұ	�02�H=��r�L�At�}���.W���&�m s��t3́�*ץ*�q=��	�� �I^Y�?FnH�>��.�^sq��W�?�Nu�4I�X��FĀb�pL�x�_�ʴ�Ef��=ӥ{%b4�Ȝ��s�U*�(�@����F&�ybF��#-<��=P=�&;��x��s�(E����ȯج]/�>n-�7}0�%��%r"wm�d��NM�V�c����ېu����%RyD�8��9<t���ª���4#1n �B�L��+!_~��N��~��\�PCS���
#Bf`ߞl�v;�ϱ���rC]$B��NpZ��DO��?��l\�Lrj�g�vJ���C��ǂN��eҙ��a@�|��l�ZC�nц֨��(ߒ�3�k��Ο���Ȱ���GN 
8�B��3��a����J�8!� �/S�b�d��!���s-Sy��M�J��s�'�f~�:G��XH�:��K�M!�!�q�� ��ӽ���B����&r�V��0<��m��rQSq?�F8�T�uh ���wn�H�RQ2��'Q�5����"VCsrvW�V��7蒀��H��Fͨ�dVy���>q�G�J�(]�mY���O�lȤx�Mwp��К��bjMRh䬜7�"C��#xF0��w=�N(.A���~�44<��KU�*:�e"5�mK�PyǓdF�
3*u�2l��ª�m����a'�i�ڿ"pj��JF��:]�n�/mj�oL��ka.��t�7A	�]�{������vZ���.ԓlDw+C'�ފ��)���>�#�p�apS#w�ְ�Q٫��ؤ� KEp��[�o���Z֮m6~��2&L:Y��l�E|s��h����V}c�;�3]NO6͒���l&N��J�}�40�]�$U���O���[7V�<J�  �&��+ïp�%�]�mO�ZF�����n��s��K�ӒGl�J^���`�*�2��˶���N�8���"�xxG�fZ�$�?L��<]}t��6�0�w��3Vqyo-�
M�tH�Q	�������U�M�C��a���$E��q\�4\�Qu�P15�]W=�b��8W�.�d޹���� �C��a�����PO9K�~��j�!�~�i�%��R e��M����
#D}��Nh���"�9X�+F�S������u�$V?��ȮxS�-Enh:��55�b�Nuqn�U�f=������C�#F�Ul�Il�&�F=֦�W���oR��o��*�0�xwv7��������C���0<6��N(�/.��M�p����"�k ��>z1�1��ZK%i��4�h�S?��%����m%�T�����]R­D�B���ү&&)�����&oܦSq�(�y�~O�j:^�M����VUQ��V��Z��g�}6^��6\��K�t��	v�����3���;�I��A�⪠�k���2�f,�Z��
�/U1W��8�W|]T��a�aT�zy�ߨ�A��/ˤPc�]$����V����yZ�fLqi�<Cn;�{Y<��2�26�%��88
�E�'#�r���U@ʘM�P�.��;K�V�rM�����P�t������Ćo5�cX��q3Ўv��H߷��+������G��V�1����zB�|Pd��7��%]��s\'�@s���yt��`�㝻�'@!'0���>�����Yv$i�'����m��b�r��N,8����汸�A{I���%�C�n��y�x�>q>��~��t@�2���Msg%2x �N��>���� ��M��oo�Ŷ���S��b�~�����u���{�K�8 X�?ٍ���=�j��r�Ꝝ����M70��
&#���Ko�Ο�������u���u�	�8���I�*Y�hS@����;���t4)�b[�/β1�fwX��o�M����2� �  ��6��I�j�~Y�𝃨F�I���5�M�D��(1�����G�m EsZK��^O,�	��Y��F���ܶz]7��1�,)����V���������p8���������Ғ~�ν������Vj]S���8�X$�>R���©���4`I�����bFE��_�ƴ��^}��s���ۀ�%��;�x1o�_3`�P2�O�D2���rT�*���ҷ��#�x��/��7�f���A_�����m6�G\W�ƆbB�֣�֥��]B�X8����A��-�T�[1�R�YBW�Y�f7Y�'	)����6�lu���[�]��s"G���ԍ*5ַ��1X� ��{�]�Um��[_V.3&+.,B���:��D|ӯ@���ff]��. �y��XU�~RQ���^M���n������|�P��"ٰ���I!�@�}���:̐R�D��X�,ʁ]P�4��z1+�A�{�%� �MF�:����sS����I��'􂤆O�F[o� w�k�eÐD5s%���Cf(�&�@ �A��Ɨt�<>��UPY��!�y?j.�*�ɦ�am����<m�!ct�6�a"���4,�u�pk�xӐ�[�uf_�;��3�P �n�~KKÒKh��m�lY�Ϫ��Ѿ��k4��A������q&$�_��Rʦ%�	d�V���M*���}I���#C�m�p�K�� 1�$��1��CY/{� �k0 �|<�CV��M�q^}WT큭e�nq̕qeq+b�Zc�Y7�۵�cg)�xi�WO[���x�%tn>Ep��?��Tg>��������aw�R*�V���w��_i+�4��#��3:�+?{�W���D3`P
5L���7_70�{�,"���1�{���$knq}Ȧ��ZVQ�b<��d�����0J[1��v��ʌc� �	����$װ���w�Ld�K �-Kv� �"�׿y4�%�L�`ϡ�ۮ�Z\y�p��� ��j�j�һ;���W�C��'Ǥ`�^x�?O5��"RA��;�Wt�X=�����{���$���F�6�<f���O�1۪a	OPI<��f9�NX���s�8��ܰ��������=��c�3Þ��6Ý6,DI���+*����[����w�̼���샼A���ù,�O:V�E1M#w(��2����H���,9�V�1.�lCo��4X��ӼǶ�Y�5���+x�e�}=%���#�������!p���WȆ�,-HS¬V�퇫(�^��l���X���9��r��RNs�X,�e�jK�n��o�v[���� *v�"�Ӂ����l� �M�/�H�k�}�eP3^L��ƣ�����.GƝwĘш-N�Rkފ��̹
��b|�e�#L�=�����C�a��br�]�O�^(Z#�?);��)��7�%�\2�덮,�M��
��g�BѠ�KӶy88��Art���d֭Y;�2�3vh�[S.��[Z����[����P��!�ɣq�_s�V��5h�J4)gMe�<oY9zi3����JR�!v�m�, �կj`����8T�cb	K��8����p�u��b�D!�@y����4,�s��V֦�����V>?M_e�{#�rY��
ݺ�1��K�)I8H+��c�)��m�M1�^���[�4�	}�;�_�`�S�8�D.�N�	L~Pu	�I؜�Ґ�����6�g@�	9kA��_�Ϯ�K�'+�ibL_��,�0�����?_'I��$IT�8�J�'hY��2�V~�9y���3)�����\by���y'�&D9��8t��$�����^��_6n��X�����G �����u�����z�k5�� -��g�Sϛ��e�՟=��rb�&�+��.kl�=x�a<
��!��J$#�WǀNy��`Z��13����Y��'럌���l����6� �!�c�##2��XVLo�mv��J
�]!40[���ԇ,�+��]ԍ��B�z���m,�jnj}�|Ϧ#�gy�H����4Ǣ{�^GV^Vn�Y{�8)!�y��':5J:(}�)H�8�b��,>����'�s�8�7�a|UA���sQ��N�b��t�X�&���_�kk����@D��z���̞˛[�?К��l�#�����C�`��3�t��x����{���\��m����@j�j>��yeK^Ex6��RZ��b�x��Y���^��}L>�M*F:zH��|�շ�U~ڑ��$�K@C"?�	)���jQ��n�W�s�0��KH7m���@��J��H��9e�K^մ� KJ��^�A �@Gd��	t����a�x���F�]2��(cT̓?$��Vp�P��ٌ� �h�G&�T�GB��>��9�;ɏD��Xf��'��Q�c� �)d��������%�j��I��j
ᜮsA�M1����݋Elz��8��c�Qh��MkF�ߢ����T��ZB^`X�~�zsr���9c��
R]}p�����u"��vDVH�z����n�@�!�Z7��v���$lx;���F�H���[�n��7>pz�YihW���iw�Z�c˥r��]���l�������$g�œ �A�=֜į�S�iU�ke�@2�97$ ���L쨗��,`�-�6�D�ňeXe�Xv[�%��@(�峰��s�d�)���N�F���������_`�J5O�tc+���jY�8��#��8�k(�|�-HZ�C�1���/,O�1s��!T!شK�L#��0η���5aK�i�AYE]��VVZ�9a��|�Z\����[\��\��ʘv�5� N6ʼ1F鸱���G=y!���i��bއE��!�����YT�,���4�)�ܦEIG'��B�y!��|�#��? �e�`�`V�gi�m�`����a���sc��J	g���}#�4��Ny��~�����Z~ �.y�ah��?d�\r�w 4s���ͧ��D��A�NUd��*�^S���U�2���i�b��?n#}�0'l��X���[�{\�H��b[��i����f���^�>H���K X����e�mLb<���pu�c�h�
ۏ=�6/��*����d$]XVy���W��}o�?8�،����r8����3,��$3p��ߓ_�B���m}��y���#]���m4+:u�հM�,�-
��I���zK�`)���P���^�0�y>��TD���G��Y���<�ƦK��x{'-]���g6�L��c�����o���-6� ��1�x}ik[�؉=�;��~2if&&(�XE^�^��N���������FxyJ/�.�U�'�H�v���؃��	�P�D#h�,�O�:l$R[�;Lp�=�>�v{��s5��)�/��N�z���A���݄��k��2��d kZ٣�e"� K����Tԁ������N�D�*i �g�2��/kxv-���x�%yc��Q���5��,����Ew(�#'���0AS��[�N��ObCK��M���d���t��q;�]3�86��:,UC!1�8��W��Y(�s@oeB��}~��6,�4Mߟ�"��kJ]8��6UFD`��LE-E��z�iŊO�?#����ñ�jX�p��1d��Ak���<:�������P#N�9n*$�0J����^�Qh"h3��E���[t9����L���O��M��ė`��ï�zX
M=�w��㧨U��ӃP� �A$�vW��S*�[w+��0��ev�R�ܙ��mT�V#[�2i	�~-|�ˮ��=�؂��_�_�/mZ������© ��e�8b�Gƚs�(2�aI�j�F�ci))eSRf|R�jƊY械����W�gS2�O�����oC�)��_p�~�N��U�n~V�",��	�]ngr�l����7Z����&Hw15D��E.[�=�Vi'�:3H qr��vt|k�+����eq��u�\.}��5f51�*�;	�^t���0�灠�aލ��ɉ�I����C`��E�qk�g�~ݹ�D�lT�蚁���R�ۂIv`遅�k�{�P��d?�D��nReP�u$�3`��I'��
0�����*	��[ I)# ����ޮO����|�VA��9�E3;k��r8P�o��Uq���{�{����1�6����Xɕ
�(��A���A�*����	]!kW�y'���@�E�aAO'����� ���n�74<J��T��DU�V*p�������/��p=����־^�q�/�w��{xl���ã��*��c����6p�<S6�}��֘�X q�Mv��ߎ��o�G��ҽ�%��T���m,������W-�$9H{k�Y��w=4k�>Q�`L-������ �j{ 1�v��V����_� t��2	�"Z{QN��z %�v��K�o�d �P`��rL�`.���+u������L�J�{�V�m�^	#/�O�׹�.��!X(N��KL-���_�� v<��i�#��e�@l/�_��J�Zv�O�sN;�t/NY��?ӄ�	���ۼn��W��|��ԡ��0!�0�Q�>��m���<����a�������'�4\��d���N3��&K���_�J�ψ컷��+��m@���uM�xYm����X�o;O�+�ȴa��Ѝ):�Z��F��r��k}~�$����0�J`��ŭ�n�fdV�DSh��čKL���v6�B������J�8xA!G���A��$C�W���=�1�����1jX���y̌� �j��j�S[C�r���GHa&�VO*�Xb���)����2�c�~����F��t�]m$}ʡ;�ŋ[J��	� ��{�cA�F�v騷l1��y�"}0�/˪�D�]V��g#�IB�u��ӵ]��g$��z��9v���C�t��ڟ�T���a�*��x�4R���
�R�
�E�/߽G��u��.���������Xn^/Y��wk�����GKM��J�^��K�Z���&u��6f`��Ϝ2���ƛtt:+���U�@�$^���B3vQe$��^.9��M6�}�U�#z'�_�u��]���\%M��xx⺽��3�"��*���$M�~�XG9�dz��5�B��$�\���uڀ�5���\�A���� ���q�$�+X&��������nw�͞W�f9�{��X�IՎZcИ8���xd��`����j29�zK�Q=���b�@�W+��`!�z��{quS�4��2��-U�p{0蠃	Abm�oH����}��첮n����AA'�e�LB���ZI�0�-�������t_�y�]��6Ѵ�g�\H��k���A�.1(V�$�[e�Q������Іn!Xo���=�#x�my�ͯW�^ٖP�6iv[����!^@�Ɖ�?uK$apMrwpİ�/�_E��_�w�P��2�PyQ�Kh��!���S��큰��7��~Tr�#m�]�8A�i!���U�n%�WЇ8�&Gޛ�X�P�]}.e�<h�,Y��\P�iӫ��c��f��P���N"9L3���N����n�o���5��v�2�ٝQ��,���T�-;Ѽ<��mI���!~C�uH��5�ͭ��UI]*���5����EN�*���\\^�vIc6�W�����Lec]Aھ�9h��k����m��Y�6�Ă�G0��+�Z�`v��Hj�N�n#}ҽ�Eװ�Ic� ����/(�����j�%�"FZu� �}�*@#�	=4ٍx+��՘�>�epr֘���0��m�"�@��wR�՗y��U�ΒHk�?��_g���uW�_R\��&���|.���8 ���Vw�Y��ͺG�*�����|�Q-�Q*�^�l��R�%�jĕ<��l=B�.3��T�~Qf�'I|�e!te��1eN�xy���=�0)mwS)q����ˍ,݋�w�t@��/S�X�C�q�����K	��*����b��vg��<���������r�d�;�_������]�V*��kT�1�����=!2'�2��^�_1Be,�g����j��>�3S�Q��[�t��j�cE���S�������Ca����4Ò�Zk�Q�GUV`b�3"��!�,���t{/����5 c���C�Ҷ��j�}�]���o�~5 �Z������B��-N�X�օ�0�A�"���6udzV>`,w.J#�2��@$p=��Z���A������<��8L=,X��v%��q��
#Msx^��v�y��7��N�6����<�{%���@k��s�A0��߁���{��}.�`H���ŵ�%Pץ	݆�9�awbqH���n'e��!Jw[,�3�j�g���TU:��=7p{� ��}\G[�)��'���^tG�ɦ���>='Ā�za(����d���i�k�C�~[���
)5"7��Ũ�w��ྲྀ[�� �����\���o ����L�G�WB�و�����n0p�?>��Jwݸ)����Evܘ��nj�ıک3
�#.P\�l+\��������Y��FYMw��^�2ɖg�[!�nC(�7�v9�p�E>�H�FZ7��R��EA�;���N�j�.��Lz�%;-D��z���Ş�����M�_��𾂋/�$�}��4ɓ�P�2���VF؎�u1 �$����S�w�Dʽ`����xO�@�*W!�\�P�2j��a�z��H5���� |�7~�+ϣ:>^a���8F]��pg�bhr�adHݾ��U΂(g�E8���??ܕ�Q��vA,ǵy'����V���c�OUi��`ذk����Iߣ#X�� ƣ�iqx��b�񝊫�m�����XO�o������Ĥ��ñ��q]���%H�$)\�-!�&����Ԑ�s��D��s����?���=����,�yXy�B�=o-�G���]�%��DF�x���!�1ĉW�B��5fH����cX��#d��~��N2�x������8Y3���g'�f�3��2�"K���UB�z�k:�֥)Z�ɇu��u��Q�f�,�">Vq�g��`���զw�<m��>KV�=�<�_�����KB�C�|�6v�8��{��[g1�a����V�� ���k8�$����m��O^п3����h+�/���_/k<q!��(�}���.�8�[]��x�w&+�٩��/���o����;�ڃ$�ׅ�K��ǰ{^�6�����B��Ȫ��,�s���p�'9�x� ���0r��f�)���[�Z� �К�)�!�U.�0�._�*��lٌ�ܮa��&[<5]�r�1ja&1#H�K���ф���z�G����j�K�v��B9�����g!�{��R�|����@��L�)3[�:ц�M8r|��G}�Z����
��kK�Y���i��=����Ndy�Zࠤ$��7�߇h;'_��Tx�����]�`�|�q�;!e�N�rH��韣��ԭ�5��=�W��%a�_Y��.'���9<p0w�)���L�;)��x�2-b�m���u��_|�6�N�P���i�2Gڑ��p��z����L8s?}A�`�v�!������Fg�5ۡ9��j���CI���'�D>��R��^x\�D�"��$�%�ą����ڑ�d��6)��IzW̧r���$$0���<�;苣��|�	:�ɷ�|������rb�E`�=5�`�:��''~=��y�E�ţ���5n���*/﫬$<JM�W��BL�<3Q�#Y���?X�;�u.��d�W�='�Ak�Y�����Ԯ@^0�o%ج1�cc�����w�����{�`4j�^�w����K��L���l�8�)�1���Y!b/*ow�N�q���w����ƹ�E|M�Z��Z����Đ��x�1hm���@]�\�����}_�������?7T�JeHi�a�&ٝ�Lx*��:b/f��{
f���A�s��r���卋�~G�xcd�o3��H3��#��*(!���h�P'����q�LJ��vPO6�]T���A�Ǔh�=��� ����'aLy5�@rs��W�9̖���=x;�����M����9+�h�.j������A�(%0�5н2×V��/����zN�6�E���j������X�R䓚UQ�f��s�SoGƷ�YԔ�<����.��ɒ%7�� ���R����~��=������b��N�-���=4��A�*f��L�%���& �U�yc�D�s����Z�Dx
t���['WO�i=C���5t$6��>|Y�$��������%�IX�~2?�''v��̟�%�g��4����NQ�p��~���g���?^(�yjƪ΃�j�5Ip��i/����;��u3rl��:���5�-3G[�XCi�H�'�Kf�4ᕡ�P����3��[?2��m�\v�c����uiHXTSH�����d)�p��H��.?;����a�(<�'�`LP���q�`oG2����W�6V���k�C�OU��-L	�dƆ0�q�����_�Uh1�qo.-�=��A���|���f�X��|���<	��1�c)����%�%0</�t�����h�]�bW�m�l�%��|��<�}[��+ז��&t�D��I�+�,b���];�y�M[�Կg��5�����gVLD��|��QE�5�Hl��d�S�쇏����ȭX���LO��X3>�O�b��ۯ�`bӊ�9�0���o5�9���o��n8����'A�Q�E����O�M���ў�lf��� ���B0��P�Px�#�i��oƋ6�`�Ql��ly�[	KXO�G&�0���w<�(	&s	tR>���}����_��%�Gjm�g:��?*�H�vI����1ބ���M��QX��	�ԡ�Ý�q�˪�Ac�aPC(�^��=~ߏ�^�vl,�āÿ�,�fo���blJL�M��z!Xi��؋XD����� ���>A��L��6��E�S����G��u8�NJ�.���)4AF$��
\ʮ5U�=��	� _��߈*!�̫������U�z����:�F96C1s<�l�5I��J����y?�u5����SS D�TZ`�����x+�����r�{���r�b�]��Q���n�|�r��t��v�ٗ\�$ I��;����,ה���`/�ogWb�aO�r@ �T-�5�o�o���R-��"K��"���h�H:��Đ��L$�C�tl����O��� N\����1��׿��ͧ��rLZ��^>��՜�p�ht�~�m���D��`p�����l�4���G�+ҵ����[�T�ڇ�r�Љ|���h�NU
�]W,��ڴ��z�ʃ�k#i0*Q�fD+�r�h��ӳ��7<�2C�~�yY�A��S�F�K�.�SlH�A�F�����ݙ�I�t�a&��OU -��>�m�g�Vo�h*�fQ�&Κ0XCI�.T����8�\�0u?
^�՟��=��R0JR�ó��5HF\�ȄT���uV��Qק���y���b�������o���-�L޸��𙯎��)7;s�%ҴJ+�*~�|��<E��u�e	*�vA���:;���k.��ƥ��c���Κ���u��ֵ��I2"/~��[���J�6��"�ϯg���c7�]��������Q���ZQ.N����	P��)~����yU�W4��	���>��|�!�i�ie���3�M﹅��� 3�X���g������{��k��%�P���e���/��	<�8Dw3߫���I���ߌ�`8^����E����tiu�^�z�/'���錡�)�L��b�V��~�+���Ԟ	�g�#�d �[�;n^xD�D)�¶�+W���΁�	Iu�UM�T��4?������ %wz楜����:�
ZUt�V����!�¯�O�]sd܄�S���3+�TwcAL���R��JͰ��QQ��(�c4��C��B�pt)G6� ���R't� `#]%��N���rk������Ղ�=��ˆ0�ܬh��~]�I��l�wh[*����:��	
=��,�]-d��sF�ݢ-�z'Rn�%m3�W�h�%e�ϱP+�r�wf��/�k\e�H$�@!!�G�ȳqA��n���ҭ�IӉ��&�D�MX���X��ȳ��jW�@7������H��u]��Tͯ�;�8�A�v�^t�W��!��cZUY�?2w�~�PYN�R���Jf��.�X8H%��~�S���`���Tp�a,�� ��[�����D����8�b�ʚ/\b{{�|���5AJ�V�Q8���MG�wJH��P��fՖ����*�wc"�e��ү�cC�|� �3��)�Z�7L����'y;����]���vW����Y���'�Mv\�<{�p��A%�x�'GMh�il0G�;t%c��r�ޅ���t��*@;��Q�-D��Mw�,I��^8�nj���l�Ű쌸�0m%�w6<D\���p����LԵ%r-> 츯C�$�.������Zo[����4�Y ��Պ-G��v�,��g�e���^>�P=Bd��8�v��4:��k�`�����,�K��+�׊�+ۚg��H�<��a�Wd9Eߑ�o�R���%]�~J��x��t���6b��o�*�B*���U@�/��շ��ƕF�c���6*�:dL T}v����a���02�q�V��e*~�I2��[��>� ^D�� -K׾�H98��J�>�K[eW��� ��u��fˆ��
�]nDf�����1��� D}�~cy�\�p�2^����>�g��o
���X���v
6I�>��#Yom�$`JُV����BGl�N�����!�\����<]�6�ϔ.�@l3q�6iHZ왛(�x���vNc���f����Rn���;ʆ��4OW�!����58�-�����8ס�T����aw�X�a��Qiab�<����̯�T��3�
cO�
@��HݖTK��DŧB���-�v��ܸ=V�m�<	�����_@Q����-���C��c��B��ƌ�[ZB���Q,�� ��%�V�����>�r�
k�J�n#XS�Y�	��K���	?���0)����;3gl�l��1�M�n'<�|:��M1�6E]xmsi��ٗO���n4"�Y���/��˶�W@�2:-�	$��l<g���:�
;�<u�oW Ϊd�R,}�;}2�m��U=��l>L#��r4@q$�.�\��+`�͘uZ!�Y)��9�!���6z���7�.o|��ePX����$�ͥ\���2�MTS�><3����,׃�^ێ�9���L��ij�C�ڞ��� �NH�[�Z���F3�Hh����&B�c/�K��vak$�Ѧ16��b���'zk�䈭-U�tV�"u��xfbҲ�n5:"�5���B���P�B���2��>aa�Wҝ���}��$9����6[�"Š�x|����-W?��Uo�ڞC�n�t�TǗť��1�9O��\��%��V8d��Z�����!1��bz˱g�q,�e�i#��o[�@<�I�g��X�)
g2p�6��˦�x�!��]�����6���ܙ� ��oz�!����^�Z���w�"�1!�q�(�� wu�w���:X�ۿ18�@
M��s���mk8:�������~����B߫�{��rV�(�N��X�_*'�b�n�Q��jo����h%����?�z]Q&�H{�-`�3���|Ȍ�uz�v�j~9�#��j��_8����G�S�n�a`��fJ��l�TW��S��{%P�u �P��Ȉ.�Yc���;I0/ȕ�g�OZ S��*��P�Kk+���xC�Q�G3�?��O�i/|�VZvH+�1QdL8��ʩ	�9gŋ"ki���_.�ܜ��⚎6�&�����`T����7nD��&�:|�2��+w���9Y�bq�mr�Ku�����<oh��M  P��	�`]-|��!�	u�܌�n��������K���F�K�h�N��}��^�����ժ����:����\�B
��d~���e�!�bY��׍�7	/?�P�g�Hb5���ĭj6_+�����-�C�y����&����
3�^�T}���=���L��q�^����� ��L!�!�N�L3�� <z��Uy#q�=�媪�85�ƐR��Σw�=�p״zvU������c����|��zZ�?������}c��Eo�x�E)=�[�q%SMz�pu\f�2X���D�&s��셐wU	>N�Aȳ�����Rv+�-;��QV=t��#!��xW�8�y<�|�T���i��]���ՖLa4>�Vqܞ=.�{Y����}�.�GQ��"G3��M����(��)�q}�G5kj�]�������3v��6��� ��/�Y����ʸCt2�·��RK8$T���r��3�D�p|Grb��kހIqt�Q�xr�7�.7�QߔN���.�i�D�ř1����&����,7{�����x$+3R��*���e���M�zzp��	�K���~j$�T>���]��
�=vx�Vu�-e4��@�w|����:'`��p���`6��G�E !#����BM�/D.���_��� ��*W��ꍪl�ד���6W�6�'?ل�굵��N���$>�v��5������ ��s��T>�7b����<%R��Ɖ���tol��ƺ����(��B��x�3;��0����aj���,[�h}c��M'�^����d {��:��o)�}�v�,�1��(8a�������V�,�3Қ19�A��6�X�u �@��`6<F�`�*���Պ��7y��@r�`őrtĸ�ݝ����RXDeaK��`��75�U&]c�s~ � ]ɀ������64/AQ����av��E�&�E�D;i�i���*�j��OH딠�s�_C��A^�1�Yc(1� �,�X�Ϸ��[z��}Y7P�����N����"=�m�L%!S�l�4^�� t��`ĳP/�I����߮M��/9/�#~��ͪ��{p����;en�B���7�7W�jf���~��b�֕�dM�ʳ���a� "�瀄��eHB�� IB����u���^�x�p�:�2վuMwR��2�/ʚ�ࡿ�:M��K�R�,!wOcՉ�;^�(�mS_�;��>pC�|nP�֚��)��h��|��w:�($p�$;e97	�;E+ �/�����8.3�,?>_(?|�)<���.�h]���ucc��6:�.	��7VuTG(��0"G��}�ynP�|�a��c&���A����� �e�8�'L�v��ׯd=���RS���ϴl!�(���ł*�e�]���d1�(�^X�Ȕ^A-�\������MTpR{��J���D��iK�&�Txʺ������	�la��*)������8m��M�C
ZHNs�V8ҟ'���v�6�]���Up��M�l��Ȏ�-+��ݚ�SѴQ!m�j-���z����,0�W�(��-�]�sG���?&�����1s��ol�u� K}�Z�Z��I������5�<�bx��������!�{w��c1���u�)/��~�f�=.����I;��]Hru�>�؊a�-���R}��e����ٝ�ڔ�ϸ��{�i�|_b|������e8����p1 AA����h5b���>\�n@B-$H��CXW�Kd��I�p2~�"��PsxZ�#$/C���iG��ԫ1\�W�.,�{ ���Z�`����$��2�s�hǜ?=F�F(n�w��$v$�4����Ht����o�NT�0孕6F]���Z�V�R�V���~Ё�6�e�B���u�=(&3!͜	����c��A��ϵ�[�B�n�G�'9�Ed�r�M5`�����A�Dz��\(Hg"
ε��\���vF�"�կM��D'B� �c��ٵ�iLxq���n�(�f'�g�%��}�}j�D.�`ߏ���,�{���e�L�[=f`X�mp2�5"�S�䒮d��fc>�|!�2�VwK�#���@�CO�o��)����z]k��Wo�k�7(�7 �[�2{�2��޺�[y�Sx�\3?�yW᥇4��y��{��Z��ۋ�P�=��SO�T�_�1	�'/@�0�I�P���<{}�":�O}aPt��[�QU�@�#�H���s���1?�7��qJhs�Q�Y���ٷȜu�Ł��R�B�R��U�/s�RZǭ�ׯ��<�ϔ<����(Q��	i�X���(u�P0㻖�3�N\cm!�u8R1/1�-�(���;bkC�hA:���*ߤ5] =C;��\mo�4�6D�ն�/�\���V���zZ=x�#�v��O��I��1�
�Ca1S]���� �D���F9��2tЬ�{͆�t@�{�Kד�R��������̊ޅp��'W��IQ�2����q�#���m���nfU�CC�_��F¦�y���-�h�I5�#��5������-Q���uV��A����E=v��\�n����X�ΎB�k1���8VK���ɂ)t�C9����K��T��88����tcŖ�~�;z�{�qk���k�tb@�Z�&�gKݼ�Ŀ�9U^�D�ëLcrb�A��k=���hi���Y�}դZ�c�pl���c��wW�O��R�3?^��
�oH���y�эb�8J��	�����@�����x�h)�0˽��n�Y=M�:K	QW�d�jJ����%�B�����2��dV��	�!��?�S|rx��d���T�V�����Tm���G*��W�
�GpF_觴�F"5ue@��t�a�X���+�j�f�)��n�p��B��R�>`V�S�%��:!�e ��$IQ�$Q��A1Ӎ¬�&'m҃��k�M�)Ż�9Z�c6杴��xf�U�mdyt^�PR��ƒ��s�i��e�E�u@?�8��*��f����"+*rG�A�}I��4��ٗP�~�D�� (�2�2�%��A�#-��/� �B�+��_��Oi���[Zj�HsZ!��@���� J�(�'�I-�:�������K�~:��TAW�jo;���JX��D�QMt.7����u	��}���u$�Ð�l�^��ZGPYF�K�I ?�#�/��u�E�O����%� ����Ah!�mM8qƗ�Xg`~*���m�I��mw�{ |�y�b�S,ڼJʐA�W[Ȣ��à'�||ac�nM+D"��(kyӟ���1�ܑk�)G	� ��V僀��A �0��NiϮ�9"c�2��v�F�\C+����yI�QB�Ɗ�1%](��"o�Z���aRS�hG�Z_ ��T�%b���
��2h�/U�d�*�6��~}�5:��Vc:��3sOFb٫2lҸ���Y��� /h�� ʅ�a�R��y��<��{�y�z�b�t�/�ot��:&�H�(�\�;��K ����|�7"6�rH�)x�Z9c��0�֪�2֛8���Ċ�n�)�n�e�a��cɧ@T=�mw6���u"�_�Y�(��`C��	=�xg 5~�ҧS$B�5I��\u��壬D���U��Q^7lSf}� ��\��VԱ�-m��6�$ޜ��t3�S���o��n�-�>��<��Ypݻ1��2���!�(mu[_	���jK��P䁛�ϡZ��2��͡�!���
X��� ns�>a)�ͷ����g�� ����t�r����f�� >z���587�S�j�kPiI�׽��)pp�1Ow�j7���\����|o����A<9W��n��Ztd� E����ք�b���O��T�]|�nS|m�_iz�wy�s��]D
�)/�'�D�ҜJ7�|~ظ��|����)^����H�)���ؤ�U��� y�Y�~zQ�����2>�l��3_��	�����	?I}dUǋge�B|j;8:���:�W�^�X@� 9�D�-ё��l����J�qSg�`�ULw�3{�I)R�^\O��Fo�\Q�z<H\�ˈ����om�� �
|�B���q|9��-���s�+ʸ�N.x*w1�R�x�(��c��&<h�!_�]�i6!B&���u"�����Ǹ�N�-D��V'�<�d�h������#a�)�	=����R�U����V$yу�AOo��x�ȇ�efY��:����g���؄�}ڭ�բ�b�9����e��N�[>�����}�<�j#<�w�b7(Yk���X�n�o4��;V�v��K�|�_!�T�A�/��h&Y�h�x�^��ȣ�W�l-R�`��[�ZA�X�;��鴸6�G_�}�󩜮�*����]�g��6��x)�N�x��n�$�	�/U �h�K��ZU-�s�u"�6�Vibky�� ɨ&7��JS�N7A;;���Ð��
��}�X���T3�^��
��6&d���%�	�ؿi-[�Yp��u���w,��
آ�{	�	m�;ku�蛇Rk"�-g�R��N�E\�l����	�0��"GI滂m��ݠ�^��f�z��U:*���b�b�����=d4��g��'��~��<�3E���Y�ϙ���S.x(�W��i_=U��,�j+�:��"I����8�n���`\lh��G�n�s
�m3&�Y@h+�!F�2��B��6��YQl6���RNLB(����7Ά֞��*��'6]�p�]�ɉ�q��}�RU����/��U ��}�J�7i6EY5��:"~�u"8mi���l��G,�����$��U������^�C~�M#�mwC�Y/�m�j�M��ˏ�힚G�W�O-��t 3��S*��z��E�Vށ�&����.zRw3������U>��mVO~�i����/��c��R;5ꏵ=t��{əL�X k��as$���Y�;�̝����?�)�)I���z����{�����S����A�Q�VzԿ/ܛĝ��~���55��6��)��DD�ɦG�x����8Њx�o�^�@[��݀7�H��`A��*�y�Mn�b�\�w?F�;�e�4����Po�{�+���	3v��4���l����'^v@
�b��0��|���"�y����h������\�@�3���q�� �	]q��;hX�;6`�
D��/��Q߻�OfDAr�R�RW�Ē�����O��t�$�@����8�!+z	_}&d��r�����ROm+	Z��`զk�1��v��K���Տ�'DXO���$�}ٍ&�%�Њ�R���:�31�x'�؀��i���z�:Y}�OwGI����V�N������C�\4\3�]e�W�I���F��߮��!X�|v���J!�, p�k!�u���cfs�Ҷ�ܤ~mw��>Fl7َS���Kp���t��ND�g|C�Cu'����>�f0�� 9��_6�]x1���yM�)�CC%�P�fd�}?�7m��5�ňU�۪-�N���jYZH՝Jǒ#ӍQ�r��{��ӑT�5W�l���R��V�D�۠򑶆_ �~�s{���N/'��}�׮v�$���5�����c�Q(E7Py!�`�;pK�����M5(.�D��G)3���KcT�AE*�i�"h)5Ð�hS�59��T U2t~�JK�J+%��ѽ���U�%穡�	Q�it��|͎WsDH�@o��"����y{�1���e蛮_�d�߁~�U9D�C'v=��>c��U-�2R���ڧ�.�9O�_o^�ۋ ;{����J���&����'�I�5ߧ,�Ɇr#[,W�c�m��aգy��L�G�H��Wu;��]{��ݚ�3�m���c9�'�;Î�-���!�޲s���!pA����L��"�s�N���3?���[=Bt�/;��q{6f���*�^��&e��� L=�U�����D��>,�M�o���h��#���b�ZϾ؃0)�ʖX�W�k�m�d��/�c�c�19�.'2�������
gN4K��7�a\b�}���'��X�n�8�L�ð�A�=|�r��WS(k�?�u?3�����|J 7� [l���;o,,�����4��<;��A�S��ޓ��MFaf�;�8�ݍ~�R5M�g�:ݹ>��F2s0'\Tz3�(���($p4Zɽ���!h��Vx*&O��M,w�au^}�5�Z��(ߦ��Fu�1]R������z^�4[?�U�����>7T�����4�/����/�.�;�<P����sY�r���q����	Ri
��������E<�Is�$�օ/b(�][d-�qzV��Gi�C՘�� ��zv�80H�v�/�JK��D[.S��s�Ɨ�6��O���;���/��h'q὇�N�$�c��3r޵�gȍ��R���[ A^|X�=�|�iu��zW���bH�zO�M?Lq�!��e��pd�b�fs4>�[��2X^qඡ7k&c���"c��Ĉ]���YV���z�G3(3ۂ��Zok�p���WJ��qq	/��{��ݷ!�2� [����k����G���G���x�7�;�&�y��p�(yb�2%ro9	s�e9����M�W�2A$��R��NA�d�G���c�`i�&�Q���iUvfKQ����X�x���%
�o>i^�)����t��w��V��~���=��D��Tǹ�U���`�#������},���Uo��7���r��<����,q���wz��L��������	���Z �%��H��ܒ �)0�&��lVATK�S.����(��}q�K�n(� ��|�Al�������_s]�C^吼"��B1Y7��E�܈H�&���Gj���	dGa~�[�6�Y	z��<(!	��N��ߍ����+�#z��h���B�
������V[Z=�J�(&�P��yz��mܛ�(!�4k�M���t �Éu�d�,�Pu^6
��Jh��;�?1I�����F��*�7��0֌+�t ;5U��(3�X�_闦�Tm����8���}�o.��/�P}8�5�i�8�F��L�$�և��T�/O��w���Q�������Kk��${��'0�*|+�E��;R� R���Vs;�J�&?���B@��8�ýC]��Vq[uw#-'�/���t"�H�l q�����0�6��x���wsT�/m�n}������|�ʙU� ��.�`^S��-ց�����"j�>ēНӂ���t����B�
�ե�
��Nex��)iYh����>z~��ԼCw���{�`ߟ�B�u�Do��Ӱ�_= G<w�ݖ׭��!:"��9�X=20p�Y�Ǥ�g�&�q�:�p�}��"R��f��!�H�˱�iE����u���uNF|H9g����s�6�to�?���|!���� ���HD?!d��<���Tx�6�P~#�;��������8k�e���ZÿJO|"���n�����It4��]��%@HK�f3DףN<xly��1��cSl�	b���r�4Ա+V���Y�~V9:F����J���A)��%�������[.�^��U���#�LNc��	��?��6���:蟇�Q�{(Α���B�!�е���A�G )�/2�fp��K@mm�M���4�3rŋ�=����+�Q3�<O�1�ڍ��В� �2!;����wTm���m?��/4֏��,20FKFIy�-�,�ӭ垵ѸTk����KP�:|}�9cF��უ�p$s�����ifP ���������j	�h�]�Z�H%�y�}t:��.
O
��ڃQ_
�#�@�D/g,b0*��t�L����c2&���:�+�M!>�:ۮ�16	~i݁�;�m����E�����Q��yQ��I+5�,��4�}2�`n��7~��mǻ4�:�m��S��c���}��l1��Y�@J�RI6�ⳑ\��L��/���)wÑ���aX���fś��1#?���	Q�p�g�Gd���inP��sr�~E����y-O�"d����)�a��K#��iƖ�{��D`8Tl����N�Eu�T�!�^�^�����M�\���Mu(�������f�i��l����J6i�8kY|�&�Q��\�ǈ�f*E:fJ_�u� '���Q�������jI0���0c��{R+�6����J���'���7\��,��tz���ٻ@�<L�A)T�n�ef������/p��m��wVRh�E�&�#B$"��^F��f�/W;D��Eעt�����2��@uq�x�+��F)��t�I��mVW��At��G�-�磝^)��^V�r�	~n=���=+�e�N���)�b��;���k��׊�E4�J�J4M��t�2����}>$���<���8 �A�%u��^�V#�:�lR����¸y=t�^m�g����D�^bǙ��Χ�%����P��S�$4!iF�+�����/-�.S�dO'4!�J��yfeSuA6�Ľ#�"���{w�I?¡� {��iX��m���������(X}�xW4x�8Z�f��L%�=o���Wl}�cU�4Ձ�Jmһu���X_�jp��)v��O򌹩��L{.�
k�7 ����s)�=:����(��Ki�u�q1�����_�� �+�E 	IR|��(�X��_��J��6����yXퟨd��b(�b�%W�2�{+ 3�_�%xN�$�ApV�Ǖ<}^-�f���k&�'c?����I�'����QŞ�X��1M)�П��ӬdY�C2��u�T���9���|�q����Z{�Z��&������(�M��x����O���)���'��N�$闯�����J���xx���v�G"~��g���<��G�(�^����6�8���w�R���~���db�d�)�!`DX�;��~�
�*p���#�������P\ɣ��5C��s"Y]xŝ������~�`�;.����������k�K������nqq��ϒ�qp:b~q�l�A֝���&[G?S�[
��ԙ��7P�r��$�C{yG����C�{���T�<�����������G!�����a��,�ˠF*�Ȩ��1��t����A�K<0%����$��t ��/��1%��+�ї�K�4,�f!n+��w��D�A�ŷ!Ϸ�T��N�I6xn�;)��R,:�ҙ!�����2�_@G���X3:"u��q��4,�$��}�θ$�4Ձ��m��8X4<l�?+��V��s�\���;Bg���n�B�����^Ȑr��vНL�0��l��ŕTسzjA��=�0W�ٷ���}P0ep^�ڔN!�l5�!�e<_�c1������I��q��[�(�q����2m�mZ�VP5Lӌ� �Q_�s�8x�T�Vlc�ɟ�0���z�8�T$%Z�pZ�4��6T8�eA�!���H�6l��B<�v'��G�{�����)��#ۮu�m'�%y9� \����Q'@�x��i�.^�|R�X�c,��Q���~��"ȀDk���L����qPF66G#��<Fכ���f�/�<�]�ͳ�2(�tgԩŏ��8�SKb	���(z4�gd������O��Xn�ץ�� b�+A�n�Uo����VY�
�N�����b\���2W����vai!ª���}��-���e.^�y��X�J0RT����|�p�`�Ă+��boX���@�u�c��ۅ�N]������8�A��ϮH��@d�ł6g�tTa���L��xۅ��/���Z�d�n5׬@�r]���ِ��4͗�U)�]iI��>���J�ɟ��N�:�ߎ�j@�΍�������s(Xޓ��DM�_]�C9����0��'f-�����O���+��SW��m�Ek�N���U�7g'9�������.�@z��8�ꑠ{.�������bO<$���؟	I�����_��O��e��\�}���hlG(��4��(��.�s�~c����l��V:`�3>�c��1o�BX L��sʛ�x5�h���wI[�Ɖ]���z6��$u����f}���^���XY��t!R@A���E�h�DOemv��D5 4k
:s<��{>��.�Ɨ"A�+/��(SĒ�Gˬ�]슆����.�Yh;%f<n�O�C9�^�a'��w�%)�>8��~��P�ro�U�eS�d��$�"���(X!v�Їz�
.L.��Ά��!7Wݟp��w?d�>�Q�:�#�s�4m̝���*3�_)�a�wt�a����*���&��럝Rĝ_1������z�{��h�x�ڱ�]BOD��bj<�{�TC��S��<O����oS @��T�s�24��:��T	�z���}�� s�����߸�`���&�~����3V�b�!Fl������h-^�#܀�]=�?b�P��,qu�Fu�I'cu�s��JXr����A���{�d�aQ����>�P�Ra�*��[��fd�E�aL�<|����}ə��x�>A��ע��|���c�wX+3.r�J���ո����z��z:��.J��5z�p@R��`�:<b]+�92y�S9�|1�E�;��> ��z���8--,��'x,=���9_�A/:g\�E�����1�X����O3�O�zOܥ��(�|�����F����ΧNS��-3��It�+�6��o��!�;�<�c$F�8�A��@+X�z~1O;3v(�TD)��CG@�]�k�S�J�͑:�pcOJM�D#�x�)���0���ܡ�|����f@�`?��O�+�m(�6Z� �`FK����R��@xo�@rI��:n���]ྑ�R�\�F�
lX9u��y�����\��Z�E &�G��E�J�R�R��G{��k�[�}-#��4�f�#��-#B��u{Ē(�Y�^����R�K�Z�7�bEΩ�A�i����n��kU��@�6q�^���]��?���SP�� ��\�Vs���/��aHks�9�ǟ�ANm�x-(�k�l}�$�e;]F�g惽j��(�yO��=�
�YP7ʗŬ���X��l�:mq:�$lGs�=�,' ��"�<���壜������K!���a4-���)�4���U-������)-�I�6_�-N�ˠ���6^�-9�e ?��EP����.�t�]wm�3�E|��Ⱒ�[�P�'$� A9��K�_�6\���pX�v# Ut�9bi�f�30�S�
A^�������]}�_7����Đ��6~$�v�14����G�7?$�!��I����}zI	��H)f$� ~qe5���ӓB'!#Ȭ�f9ҋT᤾*j&R��Y_�k4\nBD"J/(��6���Sr$Uf7RC��R|��"���� g�F��^��
�)�4��x�c���`S��.�.��/t<�C�2���y��L�R�q6{�D�g�rB^6s�� һeb��C�vz�<ub���.���JE-v��s)���z��NɅ{�-4xm5B��m����h��Fb���" -=�������~���m�1L�S��_���TN
�݄-�"�cm���Q)��l2�V��u`�$��J%��eL��4'D�D����Rv��Y�b�p����ϸ�2%�UO�L	RB"��},K≙99k�2����@���~�J�@3��n�����z�p��#�-�9�ҷ�>��<b���#m"WGR��b�d��K@r��������"�_���\g�/0�\�>)���:5?�#�L�lA�PK}����`-m^|���(U�@�a�%㉍����42;;Xi��ד��N��M�tr�La���*cOd6/�g�[�֭�Aw