-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
qq45bejbStVnFb0VZa0GWKuAtK7nBvcDaFkiNh0Dl9GXaAqmkw/Ze42k8ozihTpLZtm3qVVmzyMz
MITTx+QixyNYzE5r//sAEdRJVPKY1fwaxn3bD9VsEzOXtoAyM4cpFHC8zZ0R+gBRHmE6JsK+npk6
8yfhurLKYnb4NZUwgVJuBt0kAiLjY/GF2raX3g50nnCMeFNU69JyW/nIDdhjxaDo5P2D3AkwnTvQ
fbv3FYKUF8HsXLKsU3xguHO2uc9cGDgAry1hS+QfL8L8x1cy46W42KaSvAcjdCFJaFpkEi/H6o4T
aOBqvo/Wl83VvWefko9XgmJxi8wJ/n6WpKeZ7w==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 8544)
`protect data_block
jctzjxhn1tp0bRoZ6WJlITYxQtF5ybZYX9Y5niCL9A3YooUA/EmZykR4SMAg8IwQGzzaOKbhtf33
6aptvQV0Cp7XJsMs8VZSAgzwGOhc4qHvjYmHeP8L9CSrW7hsHHLzPo+IIghRPN/LdE4c1BPgxa6P
hVPAAwsIw0hU0iJaUSzED4L+fykdLHppMur5vXL84BfIeHE+HN8Jg7b2RomAo3HA5ZIxA8PtkFiu
kSUDPN4J6FMXncog5WliE4a50NFFoH5syg1/BR2o0xePd0Y55vhEHpZfLT2x+gK27B3aUaVEFDRr
jT575RD3Kt+7bzM3OuAgAtm0utXPrpG31n1WCJ7MIBIX6WDjtiYkjJqUa+gzaEPv8yrMndY8DaI3
4WfHV7rB2vJlwrMaC+tdsWX0pT81beUhwJHe3IiXewW+a3MWbpcDIRldNtaeQ2r+AgQGdMgxY68V
3HUMdregvQgihb2K5ZH7bljFNTSyOUVOJUktyqqbww+WrnVBDVoWhPfSRnDchSYR4dgDhg/OhPN7
yY+Pc1zWx9tKVtHNKZ4yToPVJ9CRA9AMZaqV5gHeOC3tUZdZZTKWn+5RSbD9l3Ystzct0rVYv4IO
JcyHi6kmyO/aHdRjd3hNughgNFMmFGk3+NBQ7BjSgwOjTFTc2jPShH3+Sx/Y1upMhbbp/MVwjNnS
V9Txcl16qzSknI8xN4jUYbzsgbtpZ5qw8dJB9HM0Y5nWVgGItTtL0OBJp6hYB+6AZKup5pjHfnUU
3VviWKuOmKINgXjRZyUDXQ0AxXBgbObnIMRlaIPW4f4bhIng8Yhr76xDHblE+Crn6jHOR2MTavYI
c3m9Q86lvqusl2+l5e5pRJ3rqu3xCCISDvC5vh8HALW9zC4INRfyx5UfbHuAn2CP7dpMLGt9mlMG
31irRO1wH5AVSREvq55jIX34aCLZXoEl2oFqYxP+VQl6fdrpgc3A64ZcC6+d72wd/qjtbh38Vtn8
yasfCq2lc2UwUzhI8IdmdPIpm+PFeTaW67FwbV0t3tmLDl4NUR8xItX9FWQvDzId8KT3+T447tuB
5J9DY6TqlcI+m0UCusI1CgK0iQYN2TvP2v87Ya6twLHS9q1C7MwUZGx5v9lXc1WqofFzqT/yHEPZ
cbueMiX+LBAgJwvHCj7riLypyjxzgpu2MzwT/aRfdhAQsAVXm5xgurRZKMaTD44hQXFMtUAUkuD6
P5rgAsOYwrRrXwXlBdXnejml86xxyfuWDyTqwVYxHXQylW6D8soahRfsmdOR5xXrkFeLupn8bSqn
G+usVjdVcRZMcaKVj3957m+CHZVHV5+7LiEzdfjNG3mvgTFKp9ONY0MgXt2ZWL+EivDZl419Ozw+
v8DjBYdKn2lmsE0ylO1s4b0w0udxCrVSIcyGXZyyOlX+fC/aCziFID3JiyL7vkPb6LilfVsMDufE
/OEtSwr8xGjpPtp6nQIc6jZ6Ix2uSPJnPvDy6cN7SkEpY5xHG097rtiWWFo6aC3LRxTgqb7sZjD8
f+dCd2cAKQ49e+O0l2r2rta2Z4srJi7GDIHAnO5Gh9j46nDAFfA5eC+zNJQcPyIduEEVFylyQwj2
VKr4oQ+AsidWaVdcnAv5qtxCp2Sz29sjd/cqOKeoVT4OYCHmyiFsAYtxjo8yhLYlLZrcORcJAnqc
X1zbJpFzY1KqL0F8XZOblULAzegnDMvX7rKsAndLQqvdB1LKWFXfroNVl0rpTyAhVwtDRmSl9bZs
gDj8yjrIqZnouhIhQANB2ftFhCezXUn6eR4PYyBtHdcmWdHUCSDicpdG320i8woRv7msLq0XYdbY
nixPQR2dS6NxSe7Drmu1X8aT4B3VzCLDTBh2hvA0/NzoU6lzblLCAZ3ez71DzJa/1XrNtXwJtoFN
hfTido6p658WyiiSn2GSmC0E60pVu5zyzORXeh1JpVJl34X9KsJKwnuC4erTf9uvxvL7nf/Q6Zq3
NFzhKAclCHdUxw93C2US9ErLM6mC+u+jJQ9Mmi38V1aK/cmGY0K6Ba3cQ/z1gkQglvnbPcM5xYW7
0OuD9VHIVt4KVLFG8rlhMQZnoELoQLxQObm3q5MFPTo2rmCNCvVDqyMpupTvDWgJxiNA4SREd+O7
UhOmwkAXoS35LWqaU0It4fopZcVsvYH9avl9p8PHPGSus45bIfAOEcQYYi1TB0PuBFI00f7U5/Wj
+SpyWWIKLru7DLYFTN+aF/5ZRHV+2wVnmiGJ7F7OeR12Eeor863hn+NWbAhaZUfnUe7Cb1/RNJwW
Zu1sAF8l/hTUy+iMHGol59rpIc2qLq/Jv1PqkpvaxkSe7KbzQRnPz0nY4jGeJucH+mQUYsm3gjiS
AbRONNAHSccleIpws5dHK4Ihs0SvMUMRYEV/eRNUb7WOBpvuZIPRunK7GF8+G7Y6vZy993YeG2M3
2OmSfsB0HRDJ24m+L8MLspU4/XqQuqW3kSnvntLN17isWiTa1mmPTQWpWr3bVCnknZbvLcB1Xmvl
geBv87ufTsPnf//l+HdfxrChQHtx44L6/CXZsJs9Anl64q7Rn/BDBLATxbHHJgCSi7S8CrjrQXpq
3zVVkes6CxyzUdNhp5HqTj5StEDwkHG+tzwfSMqM3uizfvqpw5PYSmDksHHVTgY3ySSfxJ2rEeOp
mWsCaNDZVd7Ye5xb4ukUWvK4uKYnU4WFluqpXeuSL1zYipcPCh6cmVq5KyVCPttMxDnxEKGidhEP
Z6Mul9IFCacmHTrRlgr7mAneySVwiHbWo248ilxxM+xb+lVuN1dU3PEGMo0lSOd06aPedICArq8c
hbIHSgD8XAm1GdQyqd2nip8U3WpZwXANPy29imE7XKHeidNbIb3Xp4NCUoJmI8wdDtKS0ihL09O1
Z3l3R2U2QzbE89Pbrnbp5+ObcUfCcx61keBUO5KFHhoouE87N7YuS4mV1eQiaZEX7L9z3+jFJd6S
uWmovzRxlhzXXjXZcBgTeloDpvRh90xi8+jiKnD27k0vDrdmQsdjeqtMMAiafYQr+Ej6MfiqQgcK
/XRMude6Rv5+1skc4m7JJGfhEFdxj59I7TOQxX0haPEQLV60hUfaaiZ+vmGcPlHrqjL4+oMIFbgh
y6mJBSqtJYic4xn5NDyB/S9VbNRIRsebsEHhWpR4a/9wjG/u7eMPir4rMO1l4Vgq4/APsVIKXofg
cLz/VvwhOrcfF9LVGnwOyMazw6M3k7BBeNpAtm0Vx16VufNCHsCDeQ5oLIBkvrMizMjIV4PSXdxu
6iNHcc+oqUSctLn3m/dFiZuIvPBb8nc2uttOZAVhfQtIRGnvItbkPmNt7TTSivfNh1nxy4u9QzDh
LGYe2eTW0eFJNuH7lNwtLwowSElEhKDj0tXza+1ZGiD57rgE+O8nLJhUez3lV9YmGslEubii9g8o
zN6c33lB6LsPlwMIqQAh+t/mcrgqYs2Sb6h1kO5nXbdfX29b+b976tuNsjEEc6GOVzM1RoN5mHTS
6nvVPm3be+ZeRCZIXqtGLLRxfcCqT8qzk+RM8p2NRF7zD0R293Zh03FfMoMRoEVZV7jW+5o9KkHm
iDRcDuBTbv2n2s6Sr0ph3kZIWACwdbSQFzbUFnlLFYo3RFYRWTuNXu0ekEj9ddTOcGIHSeOmk5sN
cz2NcZiwNUurXQaTPcZ1FhNJgMokXZIdqdQElLF0MV+FKw44kbTyz9lCUb1iMB+CTyw72b6ORVX4
y6vJWSVy6RxG++pqmVVRUSKMw0FdtVcy9k/Q+TeQU39wX7QR+YN1CzI8fPBp/viRTI84BeDDmRav
OdrPosD2LiRrhULuGdbE0kUCkxtE6wpdeiomxOgJePQ1sGIESZtGMtk7+c7GvPnnSbge1RtnGkGa
N1Pq7a5AFqfsIRc8XdaTtOIQ8eBowY01Ts/XtmDLXohp7pcR29zb2bMlSvpFKq90orw0lYSpkiio
KWeG+qlwIieCQSGhXhTmiOfcd7N4fHkb/I7lRzAR3RYiq0kbQNZAkRrM0ZnIlOWSy0oAh4xXJKcR
K7FzBFavHe7uv2F1YPTlOi/wvN4MDg9FIqEWCE/ThRjrbT9TUUEMSuADtbSXdWEqkId5aBgShUIW
QWp6OBPMlAHMTpzTNp7Gd5Ayrvg0Rx0aI3tmZJc+xoHh+Ckc5UyGzQpzTA8hrbSr1S+RYJ72MfHP
E91t3wzmAX3u0aADkLhNn67xZ/qXVIvJ8NJ5a2KegeVekJDlj7bUeXRtfs35Q/AAIEN11EvjGhU0
bWl381xwNzjyJ2GK3rtixASXs96X9J2o6gjUN+2XytQkOdGiB2c30WpuRf0YI+llpWco0zi9CQHF
pVa4MWbqX98OpdcsVJAO5AfmazFyRY4uQgyAlwh44WA4ldja4FWsHEiAEz1nfmYOQyUugS2Lt4AE
gBtEZW749vRYAKcbNqP704drZa3PhmQGi83ZFlRgLqDKyiMEDXEp+z3ujy0NrxY1nzWFEZMjBn8i
/h0vG6ck8c4tqAoO3ozbn0KmEWIC63/olupyhGGpC4+m2lZlSz9IwNnCSUZEH3PqhCUyMvyZzgDo
KIsKywW8Zmi8wTPsjj6RmSONUjPFU8V/L+5M5bsfjE9jOM8pVeaclMSIFw9rfBTb3rbnxTcRuhGY
9Nup/3MYMBHqg/rC5bPd9TzlcSBc2EukcJAj2pP/fK0qvTXaU8c+q/HcKIBaGmwW54iHLYJf9ABG
OnA4RhoUtnjcd++Tioh3gGarrN+pevUrqjgCDAiGou5lGXla6yYjm7PrNK0NoHZJe3O4PnG3HrcR
HC/xOCMOpcu5b3iQdbowARnE5eQIDac+BBmjoDcwAjRhfe4bR4tQLcatCum+a9uWU42GqG8WmISS
aipwIZuqp5xYilPLWis3rVtWT8h9/IkcUC3g1LKLLVVwGVC3rH1VmQtsFCcNfhkhHmpcbMfqmcHt
XMaXEl4cVTrefdGFtR6lGHbbj2E5SWKHm4GEmt2OCsuHkdFq43oXcwmKz0n6y/5nrIQe67a9gfrh
/0haHMPXMeckbcqLQTw6qXCKE7GeJvOn0z5Y+u8wmBvcPqdhd2m61/ikixVjffxfT+Ms59mOAfm+
MG61EMeT+HkzcsCk/SjzG1tyonzSR//6kprKXYU+4mu1LUz1+4VqmhEFWAEsmR0fbyrS9JIhWPtE
5TdvgbsyAx8BuMqiILHNUAsogi6BslTBwv2cQIj7w6LTVFmRSPp3o98FTNMos2zompkLfg6BAaND
oXmvsYLnP5ZD8dSHQz/S0HzmPCsYhjKUee/BCclEf/T26/8WqhvxI06Y1Ze7A2AZrfs2vPwDS/Da
BYDGjQeuy0kTzGBFI4IQxKH+V9R963Y3VkcasF0C8keyWrkTQKmS3C+MfjtcNXXA7OMYlkSdVpvk
DtKp6gW/4pat/ijhpt8c9HNqjyG4uNiiZEQjySbgVTRBsY7aZuSi+Hjp/9WG+2yLqgPpmT6myEoV
sway2zYxz0ok+fO4LJyq+B0j9kmZI+s3Vz4qSqqH4GzzTLHbxv0zhZ3gIwAdh2eR+8KM2g+iesie
WhKnKhvNGuM9qSWwyPLDqtQu6IXj75H9bwEWgfGyp50T06DrfBFGtLSSq3n7AY2aaaYVq2cDFXPS
xI012D1uN4OsJajfmF1oi3RYbDQxBJ1rGPcTL58N1LyqlgFQIW7x3Ugve+mh9qbeEP7utVBJdYgA
rdVsyEGk90L7y5cQwsLS7yphZNHUXO+ntm5sKMyqIUyAV8R4JMMm7bZAKAbdktMdFrdFIWgYKb1s
04dCKCRsu0WfmA057/zys3Pt6Vod7+IdfMpfO0kblA50lRwVHe5XQBAXjfDA+vSzBBN/ktAl0Duc
SIFfKt+mx5wc7wQyfCHQjeI7XnohSZQgW9rgcgJbsQuph3OUqtReAYjGsu+CYsdFyDSjRK9IkK3P
nFua/te2N+3XYm4M8ed/1efbGtE6v1ZyRHd4zEVX2daHNy/VUYkR3NIudd1XqSJdwYLEmCOxFDUq
aJMOmFwkyOVcoFLCp2/me1mhLXkltEOVDCG2SjJw2iGRDF0QULt1nBjz9qRDc92UDhFk6nH+3w36
ZM7O+12bk+CiikovEMhC0ehlqT4VHL0z6lKuEaAn6ztdNVKeCo8YMr6zNfABiWbvloA1aGT4GWu3
TKOahNn+HxQcjRpvVyk0Xlh71IDHBfN9K/akWZLdjCwtMSuGdmnqte5i4xWQt/uPWC+np9rEVLcK
bQALmTyFuWXZdLG6mVF8X8TdktmLXrqAEEzLfgPdiRFzepbOuqi4Kq+/xwXYMJ4gcNuUQ+5dcPBo
CzhPu2yCoWD83rUN+9QtOsRMXn5kpZK/ytUoIiAZd5HR5BsON7USKW4O4Hn9KeCfMb3s3+pwiXXA
po2JU1rGT1YlqnvorMMnr7B4/WEMSb22lP3kQ7aVURZRoVNxyOfRGMvNhS9xhbROczFWVUM62/mz
j/HaQoDiOQVxMj7njz9i58Mny2w6UQ27OUjd9D6h6iu55f/J5t5vF7F2ObXN3/AY+FzfnXoyE78c
068/6Skxj26lPgNxSg0WMPMeCXMRlKo8LZwjnb3ideChArryicNX6mjdTbaSMWGiPkZeQwex4IuR
/wGeZZr97hxtbCjSG/1xvbxmEExuRY6bRMHt4o1W02ZrZQrnsfJlFIfhYOKD87teNN+ljpzPBttH
dpdH0nuCs+PsjX/ocUqBOWDxAnSViYOK+FH8MujPGCEJddeaYqF2OEt73Bu5zLwD1Rcd4jhnjGVE
RG/I5prmhONB3tFeYQ8lSrGbT1Utr+AKyr/BvudxSrq5dF+ew+h21UAYxnKYI79xORYwilvUAMCj
H/mZjmHzA9vkoMr42nfHl4mcQu9SwYmsSbvuG7/kqNFguIQSdeG6Q6O6oT/GuJR3/eY4vyla7wwS
dMEuwLJwLQJZCGgL/1nZUwIrF/4J+6FOsZOlJ9rTj38iK4ixTtGJq2jqCca02NWVGZZf53bPGJ0p
0LUGiS07UKS+OyYmqdo42tMtejOfLVxwHPaSrXE9rMUZ8j1EwfSJfEUYlLc7NGtj2KsiLGu8HnwX
50P4aLiubtiHE1TquKWS5nacxcHw2MxYuWvt1ZI/0NXTxh3uSnxw5GhKBGe1EgWmxjIxVAy0JyWm
BGHqZ/avw5zeR68arkH1uoaPRDSPYGRFCYEQ6dagwGh14QXddOhW2M1R/mhhuVvAjn6zr9WssBj1
GgRdTSi9WX+I8WB207bGT8kJ5qRlXyBuDHNMKvADwhbN0ALi34kSQ5QapmzY6XYeISPRWvbuuMKJ
6gzhGzIiMk7Wq3jxM+B+v2ZRlt4iHKiLxx2PUh0KXEG39xRbxmXwtxEcWM0SEgVuogecmZjAujLH
ZtrP8rS1186kMFzj5D1Iw6pa8v3apXkShx7slnMvBgpNvvyl0cJOsMjd61RjUqsWqXFvdhydQbGG
uH9bK6BBQmUetv4lyzF8dL7uv7px8R66d9MlLYyQsMROyaUsctfbMtvVN+Ps1cJwGaYKfDoZuEf/
ocmuyIHdojMnGVQTU+SkSJzdsj7smlkI5V10Za38WEAPj1uXY2dn7Dc1l/bzNcO/TpkN3Ls73T1A
yyTQS2Gu0z69XPvS1hOfeH04jVsJecEiVwd5B2O0MTSLOSlVf7xVe5bRJsNE/r2bmchoSrVk1ggV
7UsWK2ZwcsQkckqt774p0Q9jwDHIZnTfPfpsOLQ0xkHUkt6netegn5y9JuSHLlCjp9FlHPgtKydl
3HYPHTtOCFNwyAJ/xmgcFfayq30/lPz77HIqzxhixW54X/PuTX3jNvsI3QLrWL/7YOghisueRs7r
+yn71VHI9yW8qfgIHKWuoVVo8ITiWiAv+7BzyThr4SLflflsqoqYK0SkeQyXKosmFPSg/rT3xUm2
QJmkeIhVjmfkFJEAzXBh0BSn9AD/sFq1sNt5kD2PHKLV7QYNTLzMbxuV2xUB1rhs+8MSEb4vgYcQ
pJzF9Ghe5Yg9aVa5SY3HObatCWVlVu4aezZ+axsHLAtK/3BVdXH+Jkl8rwhS0nbBI9DKn+fbjNjE
p5al0GeWdM60NY8S7LzIcynCsh6kjWo4wwM7KzfTiHklTl+H5DEMot0JGwSGkouavWH4f2QoRtPL
A1kT5Z+uT600visJY2O31bSclF/jbdJnZBq/4XRHhwG4SxABaYvjQbc3ALgdaC2zPJbXJwq5JiEG
1WJfoh1lCLcF7EmufhGWw/tEfmjNOV9rsJO2XIQWccldXeqnrY1BGViUi8AGNh01twCTQPv/Kp0F
lEchGC1HJBOgw+7t5QfBq8zfY5zVbCUV91TOcyxZVdwbYO3HUhTdVK05MFpsK68ulZ2sAt84WzMJ
BJf8QIwfgpwRpTc81AwimjoAZkT7w5/p34imw0+LJ0S0NK+xNqjFrO7AuR+r2xBkhqj6gqsHOjdt
k+zfAe/ujmtNQmEk8sxC/WEYvna3ZI6Ya0zytzRFWOdkQ1Dyf4gNT6V21XojgMg514Mxeym/Gth8
2RY07MIW8a+ZIn9vpsYOZNk6uskstDPpMAENP1FVchjdyqVOmoWwNFU8HN98zcUZcAocxEDh01nu
q//gwRwjiUGyrit8jSg3xQjfjL3UHs8mljDI++efu5tPFiqeJffkJ7XDTpFsq3D5esfkrzS1PcsT
dzuGpjG1AhPZt3dCaBl+/PRjCuqoKFVBLCXNbrYsduubnTa3Ly6VbEa6J5axPWGUipHIa21/8pnh
eg43PK0lj67K2jUZbjol7xFrrnb3ocbVIGwdLWmu0xND+MEfLtnHc4nDj938eqYCnr6dvvCsgpQh
7EQjUC3brKeWplAqY8phe6fstvUzNZRc3kQaGutME0FZiyqSKXPByAsyRZjTfqgMElMZXcO+Imec
B77FDhmJUWUtQF/A1ejyoUVL7nHPdkDBz52V0aQF7iylQ25DiM8e59NKxYZvbL21Jq/Rs8Xqgptt
o6VMYLTjtwgm6F6FgwuyWTcsyJNQLy8ZQ/SbCNEv75bSM4rOSXrBsiRXVn0Ov2ccEPp5cRaGeixF
UTy63mWLYqxnmiF4/l8RuZ9UwLloh9BMzfupf0bHAk35lbj0/2tAwvDc/zQ+12CImsZz6XSA3BAn
2YJ+wCnLYRUDfmmRovGMqPDkdUUEtjmMVLuzJr42AlazXJpEifQLTpX1fqxEaWGXKCr35SnR0Lh8
iBLyLHSejtTtYUDpP6BDgNZ0xVyW7v1T+O/kzwRpxxmzVaMm0Qt4CiuJATbIYD9SK7arcvnY+Dnj
55r1oE+DTlQKBWwgI1QVPVx0a+mpFInpp0sNpIDLD2uiMnGDN3K0qLFJEkZ8Ilj7s9eeYkdrFNn9
2pGELTA5+uj/ew2C1pYrHoOm29sYKtlHD/hKw1H1ELOpQ8/0j7WLkP5Wp0tME/Z848AvBEV5rqtU
BjvNIDRMGmOvj86SREvlXe2vqcMyX71mRQdYcFPmbmUYUz9ZhhgPbzZXHWoC4qmSu9PSeaFxwaOa
xLbKnuN0w3EyrknwYH4FI2lN/FJ23Er9qF7JSPAw0WScou+RbFrAQLN3abrLKiJM8FIFq/I8qXRN
DtLYBmBUNtQiJ1n+9dpLlUh/MqhRNp/JMSGVBAaay0Wru6uoZcJYphaC+VCSo80DuyC5TgdKEZW5
W2ZBwz15f9V4FIlvQCaeF8tbV1ETGzCYhG/hHUt0cRbGudr+0dA9T8F8QLZFWdLTjvsywF0jK4n/
t7omG1Q0xoJX3YRx7Np8tzSAhpFtMzRTItr0EbL3vZ2hBHhciOE5oD0pAU1g/8KqdgfHMoIYLTVE
LTWPYuRuH2y9fhSKySqyGzIq6R6eZPZBg0lQARsqPx9kl6TKafsBhReXfa56JuHthZf6Yud9VOBJ
JJiksd1iyJAaI+nJU+7ZcYOT4immuVGon9OGsquhxag5KiGOoagUL7Gy5sreyDnfD+hwwYCS7ByL
xOIO1Kv20o1pXPiwClQb0huw4p+ATUShEMFEQS13x0d6vl7jMeBeuvp2fnpFEi51xQyXDD87+ZC9
41uMS+yi63QEIZTmWYMO+iW5BAPCd5bZqpxm9r+x7akrPq4Icp7shZMHjiUXjM1D9U8Wu7l6ilYw
dH1kBzWuD/kPVt2xSQmSM+WiYLiIFXHEBnJw6LR2BV3dUdiIANlvzxFdQjzcF/GslfpapJWT+/Uu
FV1QbBV68iMqGObCpjLe7aSO6ummLf+Yn0VR4Tm6hb02e+roMCOORrtY+3+jf3eSDER3yviSQCrT
7+WcJh9lCU2emTc0Lb3yCOJRMRRlM5Sh4n5sv9HOmJmJDZ+EjGCA65trevy4b56tQ6ief9T6K+PX
eqR5ijLa+BT8EfnSVxhcNkuYqb3CXmn2rpAHSFvhWJlSZbIbTrwLNyTXaUKLIIhE43+SWQ7BQlGG
7l25l5rvIWSc+xIY7I25Is4kaie4w3yR8hZ1ggFmuTCB597V6IpqInLicxQmHwTwCP9jo2eHrUhl
N58nlLsmQu2QLan4RXOThcThyzSdlVAfLjkdRJf7vbtChGLXpAvWN4HY5mL2SVAAgp6kl/mqLB/u
uCZycQfWoS2nMNFnydBJ3adnZs/mOA/oG0IXfQm6jFw8Cd9ErUUSSTY9APbEvcwKvaLDb6ghZJ4M
3WlftZgRFc9ehihxvaONZnUzeeNglMdY97jrgDLz71PR5ONPYxP2PscE/VdUu0HPuQZGNfJZYhy5
OM8OJBi11Tp4V8VQsenhSiPslIPSJxKGyFb4Y/KzEtbK1kia96fC0WJavGztsRbQdcmXcDJ4aisV
leVEj14ZDebiubyIK2TzJcZH79GxUtd0bpyhxxW3C4QcFD2dY4reAj8zH8BEMgW17XaqnzjwxiYg
CJHH3Hr7+/e+Qv8cfZs6hLi3rSePhCLQbuk8s5qVi89pRT8hzpDt6tJvZN0BQeTsvOnAvlKHPsN7
tGewOnEWo5hUElydnSzEfhTCjMHRbiOE2plu/GPYZRZ+E2h5ROLoLtRBUKTzxoE9TeWg5Ci5aw/h
nvx/HFNKmFq+NWVRh5KJBth0rWeAJpi5kJ74sxB9RQ381ko+0IUzLKAUhnLsECXWcNMuLoDeUb4a
Un19BZwNaFMWum982fNF54keg+mMiES27zGxgY6XQZGpTQBxmFM+yag/yEeWgTQisuVruOS6ni5E
yLlWkw3LHdKPnSaN5MroHygsUYp0Ww8cokx+9azDhDf7UKst8xC4DjV/5kenb1aBzJ/hQux9iR4Q
Vdsh7FU0JKSkM2mAQYTZbZDJkM+9vngrOmcmE2lFqOEuyzsOkYKLsGbdsPsOM54JX5f6xw/eB7eO
K/Hsq2qJE2BvmbrpeP3WWWhGGF/AeeWI2inRYfbEmwJYVSLbAIgbM68EAkiHbBWD8qS7
`protect end_protected
