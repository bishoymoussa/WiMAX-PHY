��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$Rx�y�<��wA�*;�x���@�̦�W�X�fa�M-$u����n~�%���P�$��W��kYَ���P7�?UMfT��q�6�U��k�>����~�\N�(�����X�e���/6U|)�X2pF�]$h���d.���9E��WG��L�X"]�Ad����ľS���8od����e�GT?y	7�������ݵ�^��R�q^]�鍦�����s�ae���h��L��P_���ާ��YЭF���'\��68�b�[����w8�[X��V�F�0͘3����q諵�uW� �h�u\V�?@��_6G�_�*�G���B�絉�f������[�G��U&�����~�F��AׯK1�`c��[<��FY���4I� �#�G��x[X�=�Q1��`��R>(�w����R�O�?����7�,(�H\�#h(W�EH=�������yq��Ѿ��aF����:�U~m<|��.��0=�P/���4ǆ���T(���̬��A�Ɇ��0��$Bt�k�PM0L��Ev8g�.N��M^7w�eY(`t��M9��N?�r�/��yQ(XQ	���NP��Я���rV
�����2�U_�񃒟Koa����}�t�����cX1�Pr�*Cu�_��蔙mD��vG�3��BS�~>��2��e�@�,�_r�?�3���W^vȃ�H�(B�����G�}O\��i0�7�f�U���Gӽ�y�_�U���gzc�쥏�*�ʻ4`��и�â�&XƘ�0��S���9���R����>�\�Cl;��������h�&i�n���JH�N:���L쓘��
T{r����������������,���W�d={��ă�lQ�f��0eC���j��y�W$�6�#�c�p%US݋���iO�R�eĄ	.90z�^���Hlcƅ��=�I_�W��t�j�>Z����@O��p�\gÌ��|�4
�$ҵ�	�N�#&������-�=�	MA�ZE��Е�m��F藩p^~T[N1�@"�m�à��r�Mڞ[2)8w^C��}yj�N�͟}J�=�N7{���x�
�9x��K�~6���b�dQmH��;���P�5�Hh�o�U�Y/k��<5�*໔���F�g�
�F$���\�kaJM7���Gļe9��3Bצ���3
}r�	�A��^�+,�#�ȭ.[�J[�Q!��=�/.uK7R:�5k�+okW�kܫ!�����6+U�mD)���RuV�9���;4��P��sw�������Uƃ��d�\~
�]���_�Rg�Q#��g�/�I)����E�����%��3(ַ�-CQN<�WtC>0+�t�2�Vd�h�M��-��Ky*����jYqk�*a�M�^�v&��c�P_#��1Y��BP	F�	Z;�!��_kaiaO����ޗ=�so��b��#�+�\OYY2�#���t�$8)�O�,FSQ�<�;LD�|n������xS��fKZ��;P;/oc|���)�Wg,��Po[ {��]�8���'
�K�(}p⻊0q��ob�k'�W�o-a&	햕_�K���P�t��V�b>�<� q������`�<JLNS&����`ޝH���n;u�lx{8���n�i�5E��z&u}��sz;��rz�S��N�o�s�J0|
6�d�`ݫ���	�VE�$%B�B��(t�O��dÂPi��q�T�N�QUri��G5�������k�Xs\�萤�Ϋ�D��[r�74��A�Mɖu8������av�1�;�C�y��
�b��ʭw& r<����dѪ��j����EDO���f��F�����Ѝ@8��ˬ
Pa�Ccd�@I8C8��f�_䶎fr�*����m�EV���	���M�z�7��m��dr|3[˴��<��q�N2�]+c/
�f�a�h�8˧��d���ϴ�Ihm$��<�;l�/��H(V/7��{~��u�z�M���^���}�WVbI�%�Q]
BT;�Q��Kx1yh��E
baUŔ��AH��z��;�S9��~�v����2P�_n�J�`���J�e�V<���!CI�h�g��ǖ��\7�r�MN�O��)�r>P��G���ϲ�z���U;�2V8g4:�w���	�aK�hK�����M�������D=�
yB��<��4��kI񾙉�Z��d<?����v����#�֖^L�@k՜8�s`3�'1A�z>Vl+p����'L3�!����nW���\6ڠ�R&�+�{H�~�>�IxPcg?ý��b*W���� �^p� "�M�8�z��C���������d,�1h��XXT��N�h�5�Z
�	�)��0ٔ��H�4���v7r�SmY�F��R��g���d9a���\GZ�N�)ve�ʪE�c�X���%� �����(��Ci�v�w�/��u�ʇ|b/���������Q�Ң2T��?��fW�$&L��ǁ����T��(�Ӫ�ݣ.�����p򸢅���Һc�]��*N�4����V��ݵ`Hk㇥Å��Õļ���;�覉y>d��@+��%��= *�\��E.����،���fon��{���eFY�1��m��t�a�_��!���M�����,(������f����<�a�3tzr���ٯ��0q���{�>�S��U1o0M�'uM�5 ��/<Z>l/����̸^k�
^`!�Lٳ��``t��*�K,�z*����Γ���F5��+�Wy�VjiI~n�}� ���ş|e���x �>X���>��/)(�DT���d�f5��jJ���D ��Z`�6G��Ei+c0��W�H�j�;{v?�X�U����n+�4���O_�J&�[�0��A���Kf)J�%'+�s͜�v�"�L��ŞOZ$��Ŋ;�!���o��@lb�w����9�"Uɓ�JQ����01��(-�̫������]�s�q��O�O�#<as0����3u���u$n���ϐ�rz�W��l�?���ߡ@�qa� �s('����"m��2L�$�v��T0�?ꑕ�&ƺE���::
������4�-�E+�������X�9�Q���R(���,��lI��\��P�%��}?xJ��#��b�G�`F/Se���I,���vY��{���?+�����ђK]m�7�>�x�J����X,��\=3�fZ��-)��O��{)��%>�����R�ް�61gM6`2����׊:�{v'�ꆄ���ǀ&�e'�>�X�D/�؍�.��RpKۥ���Ez�$HYK��/�u��k=�ꕕ�܁=K�w�Z*2!�j̘f	ZJr^*t�ٷ̜��&��/�˰oǬx�K�'RM/84��j&�н��(���Թw"��Y����h�c ��^�/DBy�sH ͅ��X����/��	l<�[>�1^�D�����M�7Cj��-&�W���7�r?+�xpD��LcCK�iG� ��r�Z�j���������l{9�xqm�ǁ8}L�hs��v)�E!_���X{K�ˡ�����_�Uڿ�� �N����U��b"NA:b�{�^lȁ���C�N���X���V+����e!�rl񫴶��p��NXne��ywX=�����1}=�TJL8���;K��۝�dQ�@n1q�Ԯ�xS�`�d��t�j��_�4'��u�4ucMUD9!� hw�2�XH�L�WQ�q�M���WNO�3��=3����1U�S�8S�!H ��Tׅg7��RW`#a�l�8�s�`�9�}�/��P��o�A�����͊�V1�����b��b���)~4�B�� _�H����wY�֯��PF�^6�v00�.�WM&l��r*�'iDw��Bn�#��g'�G)�s,' ��94�k��1�}�q��hu�g���?�V�ʋ�/�g-q��ɢ�.~ƾ�hw{�E��%�-= �o���v����$	s݁J���u���$]�TY96Q��*K<f�U*x�hu gP�flZ���>� ��bXp�z�ZU����^���0����-@(f�D�&��px )�� �ڦ�㨈�C�4oU�&]mu.��<8D��|@Z�X��r,�Ч҇oe>է_�uy�\�k:��|'��]ՁN�E?�O��� ���$ɦ�73�Ї�cr�nc�m���	��MJ�������h�U)�o�� z�rI�\y��l礧R��t�6X�x{/�aŬ�� hQq_>&��XY\fiI���`Q�~w溧uϵ+AB�# �11���B}�dַ��/q�'�z>o�t����^K%h���\!�L؆75����n�h� ����J٥J�[s�]X%/���W� �Z�zX��nu�`��`�e����'�v�����'��+e���<p]�$��gHṧ��L�%�n�g+�]��8������#oG�(}�቏2��7}ϵ��x��7��J�<�N}m3�㾇)��|�5t#��D0���s�)����*q%i�f4�����U��q�q��ay�X\��9Z�;�EŐ˜CM��o��7�z$	pg���ZYh�)t��2tV��,�`�W��&�]	nϤZ~���w>�H��Ug���˗�܆���g ��ǭ��7��娳
u{!�����J�Ӯ�=��0���u1�eo� 	�!��G���H7ag�'@����.�4�yXA�`�)b�K�@1�m�A��������D�&��ƊS�c`�;���ag��U v�����P��G�(�%�|G�-%m�ǫ���cIF�X�5�Õ#��d ~%@�T=����h84�7(��ۓ�dFn�Ϩ��֬��ޘ�Ң�}���QXˢ�Ez�n~�פ*ߩ�S2�ON���[I�ѐ�h`�jޒu*X�Y��cE�1���^'������(@�C��f�r��	)_��w}��?Շ�Q�me�OY��v�	� ����@��u�Z:H�­�AB	���!���-�������Fu)�!����/IV�����
n�"�`?K�<_��j?�'����.K�"�o)����Q?F��P[�G-��!���	|�gE��n�~s��4M��;�8�%V�FA&-}8����R7�M(����Q�ĝ�VL_ ��N�V�(������| L���;��@��n��)��.�$���`?�~U-���uWQ��ٹ��I*_����/B��ެ�	 	���,��2��'E��8�w-����^ZX@���^΅���>�E��]��-��������-�ҏ�ngV��5�j�R}]�ר�a2r��]+��v�Vq�ȁ�������*���du���I/�(����f`5�I��!�DLk�5̽t@��L�0�ƉT�j�����G4	.y*f�TNr�Q��a����,Z_5uSJCǿp�v��+�p~թ6�D���:��[�jwfF�?��ʆ�2N8�঱�
�
�w*�w 
77n���~)�H�_s�xF� щc�G�-�#�M�����Ƿѭ��m$�в�������9��v8�����@N���Dɏ��Q䂨�f=Fdp-m�;Kp�S�*�f<���sG�8^�0��9��4`�e*����[⇭8+�����R�sP7���ɩeS[C�}����g݈�s���Iz���c?R�'�޾�����}\W^C^WD�`'��ά9C�V��,lѪ��b������ho�V�m��݇hl��Ͱ�9w��ȃە�#�X��.����	��+�WQF
�֮����ڛ��]߅9�󡑱e=Ɔ��b~��m!��k�VN@��o���d�Q'��-��X6F�ȵ�6(���C�{��D�)9�=W|�M�7��#�K��B��
8˄9=��7��S����"����n�^5n��>�Ťmf�Y��f,Ҳ�5��dm�ƀ谙��*�_��Q+����OXÎ�ǵckz�Y=���DBG�P�3��S!:t%�zu��^���>�E)�EJ�#�F��<$��~��w���X��*ӽg�5�� ���&$%@��[D}
z�Z]bY�T����TZ*�"�;��%o0��l�p-�v���ӥG/51(_�6���OK$��Ύ��\ܽP�"`�*AS'������E����i���.^�mދ����}��)!NH�m�����kRd9��A�,s��]$̢NrUHձ�LW��9��O��,+�/��왒�t�F�L�� �0Kۖ��f�U�������\�)�حU��$:@_R�':9ji��`[-���U���ΐ��Q��U�՗�vp=��).�vX����O�ߍ�F�
��w=;M��yw�����2�)s�(�Q��j�������k�PKrʋ&lX0�I�DVM�d{�Q����z�r(�
d�O3���^n���X�r����ߌ�ޣ۝7䱅6up��B��ٖ��_Y�]@v�M���Y�r�V���ck��(y�C �﫶�Do��(���5�,Q��p�+(ļ��u����GN^p戒�x'%if��i�5�  @5�{SD%į*(��'�^���Ц�X�ꭹ0~����c}�D��I��j�4�V��d��}eg�|Ş�F�U��J�U�L#�7L<v/T֝N��b\���,����i��9?�o+��n�����[V�njVyBC�v���ڠ"kF��f���J.�(H/Q�����N'��F��4��&i�.z�)�+��/�b�s?$��e�
�H�0x��Cn��96����\��l�xU1}�+���I`��M�H���� �a�h"���ȸ�MYwu��Dz�2�Sz�INh��^v�uT������ob��, ��pL���Y�)�򊲼p�K#nbX#y�z�nCww'o(9�֖U&���·���WT��]-u�'s����]C/EG�=N��k˻��C����H�֋��3��J�,N=Ia�퉏��ƴܙ�-ފ��?����ޣL�(�^ΤUKp���|<�'K{��W��dՏ���Q�>�r�z�Z�я��ɍd��Ȑ���4�[�j(wG��e�B$�YP��=ЧA��r���fAN'���eZ}��43<sg�~�Y	0��rg����X��n���7.�f�ª�f~��W�"fj�yӸ��j��ܤ��7��\�d0�@�~�[�ϕ��:ؾر.H\�ȝ��o�^�-~��x�G�`~�[�z;�N�n���c ����fG����$�O���jn��dCh+�Aufeo�¡Kk����H�6�`�ek����\���ȷ/Pyp�ʨDdI ��P�.��{�0�p7&9�9�����(���)@�_B�)�?������Mh��)�5bZA�^b4}Y3Ti�@�6y��f����	�hn��$�έc.���W@|�V�F��폽
���y��)��"/l�x	���+2��s�(�!d��#+���?�2t�v�yOV����c�~�/�;��7|�)~�͌���̈�͍s�}4q=u=^���E����v32Rt�%�;H�DZ�V�����=kY�0��	�50�.������Œd=NC���-b��f���Z�[��T���MPywՌ}��K70�.����2u��!���ءh��q��F�p�~C���n���e���r�AVD�R{���B=��{�T����d�î6�w�E�МLAa
�$�m|Ѷ	��^ʡv�p���%�zh����VEK�&�����nɴ<��g3�@'�Z��-r�9#8A�8.a��~�@���4[�̃�a��>n�L�$d�����/�y�lˇ��{�Q�\��z�B�y|dc�vxEڣF�,Nmh�9���ri���t�A)�`f[��u�u�F�5i�$�g�:�(̉W�T��ߚ�H��cj�$k8����vz���M�Uf�q	oN��ȭf(�|5�˗�Z��ʿ$������ �c�j�6��U��F���U�Kk�v��k����Dʑ�.�@t"��ou�c!1�����e�97<��"���}Y��>���(�-o �����VI����ط�(k��� #٭�o/���j�7�r�/��.Qa�Sݖ�c��3��E�Rz�?08��\-z�e׏:<��̦�}�A��3v���I�S��M����6�`g&+���O{���m��2�� 4��E���d���p��B�̓��ix# K�PP�G&v!	�S[<WLL�l4��p�i���`�� ����kCO���X9�,��2��u��3ݗ�z�|g�d@�EoB�wY�N���iW~zHt!<��<3�2U��og"��GÜ5v��ѵ�6��)�l��+W60�9�6}S���"�EE�"�5-�����ئj��)D�T�8�F��������̎�~�ˍsbSE�4��p=�G\W5�并lF�
*�nk �����^�n.����  ���]O�䛌9$m��[�B~s���z���@Xk�A!1`��(a�1�M�
��q��{����ʊ���v:3.��>Z%��kym�6������Z�I���"��'X`�>#���+��/�Җ������&8�x���:'�W+�ݨ�4� `�C{mȺ򚻘����+�̴;�G���<����_y�g���s���}�
+��*�|jZ��j�1rXb_u�&��,]�[m}}��)��Q���� d�Ǩ��_(j}S��%A,������W.�l��H5e<�#:c�k��R���X�x��
}ބn�s���z�(��^�2:R߈�ܤ<0^�f+g�8]�֋i�6�����Y���"z�yM?��PF����]�r��5Ԙ⥱�}��^O0D���-ߒ��X;
�T�I<�O�:6m�8z;� ˴�>ە�ZI`s
K6���������,����\IB̘Ԛ�x�=����߮�y���������@����m�+<6��cN�F��9Ɖ�ܠrrW���~4D��oU.����t�
�a�aF̦
�C�Ž��Mک�."ݑ�F6-�P�E��6��լ.T�Ɯ�G����ě@`�v���'� � �RX��^��):Ҍ��-T=� �	Ұٞ8����[Z�4��C��]�������}4�q;P,�8X��w;���#}�%�V6�/3�'�F���@^߅�`�۲�/��p.��z���zPZ-F+I>@øfS�=+]�$�%��������BG;��^CM5���&���>�#�Jͥ��0�9Fv������Jn,���<;�K��d0Xy��{��|��WZ�K�7 �����π��g�译�;�r��]FE'o��9$�|��O�M�Gl��׾K�O��,k�ػ_��[�_�Cy
G�X�߷\�#q{��9:��-itԭ��4��� ��l���h��P���,dQ��w=�T�zeDtta�J
�#ra3c�r�)t�-��mw��wr�~s�lF@�QB�W��˜d\E_V
�5����<�1
��9[�l����ķ2{d���E�~G���c�"D�d�f��3���6_^MB�=�q�1��`���"�c�@�C؄e�s�13������J�`
���l���Cq~B��`�9 e+���⌟q�m �X2n��"��;�Ô�O��ace!�����+gu�����=�ַ���U��x܇ ��-�;3���� .:��
(z\���U�xR G�Z���d�9��v6u�)H�#�D��,�u^��-_Z�X4�!Q����%����`�9<]V�g)��-�	�1�r��D}����	F5�'��<.�w��&v��>�s��Vf�q���9����ߐE��[���q���R5Q�	�.`��dg]h�ܣ�8�h�a��1v�x,��B�IID(����4���a��ɜj	���Zu�X��u�&�y>��QC��9jV	�r��7=E�����7'g�7�h¡+�{�:�^�"HԼ8��8pO��hL:O�F����[0�wǓ`���q��|��=Fc��F~a�6qe���:�[YǇJ�+���Y��ڷ�HiDSv������*���1��$��*��ZT�l�m��Oyu�O*ZOP��ɲ��ف�XX� ��B"#�"\�c��8��0me���F̓�=�v]�jw�o�vF��4y�iE�U�A?D�U�6�O�%�Y��\�c���f�yb��������[M�k�Y-��ATg��#��z��>\��{TC�֞�o�$Br���W��r�R������ƙB���3^5N�/�1�@��,O�|ƹ12�̪K��)�6���Dӆ�!Ƥ��auYѪ�__���Y^Jģ����5u#�H�F�T9�YQ}�X
:����|@9ye����Y>����ːS$.W�`�m?9�\��{��oA�������Ϲ�ځ(g��1' �&��,�ST
��8���ݗ9�x/Cٺ ���`ڟ}�Y>��_w0E�T"�e��`i6�YQ������}o�>�nu����:��w��@Y3;�I"�?U2��{�pc9��E�j7s�RM��Fq�����B"��ڐ7�?�3�2��گ���!�Mܹ����?� -��`��Y5�����k�?�`�&UC@_�`�t��½e"R�m"xW�r>��	��!��G���P&�c����v�CFƙ�u�E��Qb�8��~^7覕'O#L��u1��<h#E���E���X䘨f�SDZ�ߔl>����S�S�^��Bjv��<��h�RG1����E�4u�ݱ�����џ�l��Wc|o��s���5�����Vjc;�L�j�q�:2_ʭ:yc1���| ��bަ*a��i
�+~b}���u��0�}���[�"B�f��>	l�R���Q>ܗi-*�ƣ�g��
�SuU5Z6Au&����Vf0�Z��c�T�5s�{{n-B���W6�]�)��KͦL�ek(l��T�M���~V*���9ۄ�V�H1й7��M�<���}#t��+�$<�0�Җ��;l�N��S�W���t����iG�.W7��=w^.��ˤbc��;Զ��T�Ŷ�=�<�:9l�D ��Nq$�s�
�
Ke�0��K#,�+<:/@����qYG��ZPfZ�^bE )(u&�;����)j6�~��H0+�t/�@�~2�N0I���?X�sG�~�)J� ��,���2S��5����E{���{���̽h�.C�4��շC�͆���t�⼹)Ȥ��&�.=�N��3�f��l"�_�2��{���0٣�t�*g�f��{��l��w��^.xn <Mِ\\���#��"��t]~�@����~�{k�]���K�^��P����832ca���~-^A�v�eM5�JZ�Y�C-�v}�o���V�WǦ$���]���Yb�ٛk�NsF����y����: ������|�j�CLx�t��n�l:V?�P7y�+��~�E�RU��;�;��-% |�a�^���U�_Zc�t�F�u�*��3�����L��T;S���ϓB��T)��eE���&��u(��K���	dcoj�G~1�{�3LAA!�⺨����<�w;��X�N�^����@��P�,ע��-�WE��[d;l@/�ֱ}�8�>J77-'��.'��Oce�y��������Ð����5
��?�ͧ3Q��ɣd�gL�4�Sly#���"���QB����<�Ã�/*�/h���D�_�v�'r��(�c3,sȐc)�!��r�B�G�f��t�Y�ύ
9�=eR��jZ�%S�����H6q~OP=ot��ٴ_@>C1�;XL�N'�z��0��(����5�����z���|]��
�4�N[���~��)�k�_�T@ 9|9�E8R7�y���d2�-�ۯ��L�Ď��}Ҧ+FP��P�&4��;pTy�}�r���T���Ⱥ��z�;��tt��oR���Y���WR�����%�$1��n��-s���������^PgK�j�����������dx���
��9L�����tz�NT9/'���7Ѓ�]�;L���Ld{�M^\�g>���Fʕ�a�v��1��ile>p���Ϗ½�2)ͧ�h�M6#�ݪ�ڍ_��Y"���&�>�}��B�}^��e�&���=��
��KZ�p��^�	F���`��%rL�W?�ƼƉB-a�8ȼ\�#��g�m��|�4]9�;���m�d�N���PF%����¿�ne��K�a��Pk4B�x96�4<W<+��b�#�>@����V	MJ�0M��h�ݠ��`
A*	�ju�*+�j���vN���{H�q�޽h�xn;-�Ďm2%����1���)`��K=f�Wv��H��E��R)���Fh�%����� n+&w���so�M��ߚvV�s�/VEN=���^�oPnI^4gQ����nJ���n�P\SH�ǃb���]X�bȢ���f�k�s�IVv`��t7ŋY�4�$J�<�-XdQ�������20P���>� ځ���*y�^*ڜ�"���<�#WA	�w'���� 8���Dc[6�$�b�#L�_�ɮ%�d�aI*g׮�W�ZM�?< .�8�HC�yQi�'`��\��^�a$wf1}�d��f���������+���K�����5h�����4�6PD�P�u��rS�a��(�0��(rd�,���ί��ʑ�U���G	�$I�R3[��1���
�rP�Qmh��Or�Hm�T��}�\",�/7��[n��V{)hk�_�J%Z�BD�#�}�����L��p$�:S<Cj�l<����.��Tq���� ٷ�o��K��mn5�d����z�n�:�4qz>{��q�ջ6H�����+�	۞�+���I ������@��G�sq���~$X���l2�7+)ݻs�v�a���'���kI� x������t�y���7%|9���}E�c�Ε��n7��2�Į�u��{C�LTG5q�����!޻���zjۼ�����x=���Ay:<�A�+m�!̈́G�g�����1XJ�Q�H�����6�k�A�H�|��3�-���b��u�m�d��s��iB��q.mc�#Su�䲲�([isD��Y�Gn�?Kt'��I��p��R�]if��1�m��?�\�^�ަ� cH�V��r���l���C�Fڼ�q6)��ti<\DT�r�@�l q�]­dj�KF�r���F��.z�]�7���g��^Wb��#�e�&\�r`/�ʖ��q�7�ue�s�#��yCl��2wc٭���a!�g([�J���7�=z���Dx�.Z�$�w�4�Ĥ�ߢ�&�-q��?؎���õ���wE�Xwyh~��R7��\��©9w"g�W���x?�h�V����I�I"`��V�
[�E�٪63C�I���=gF����ǘdVQ�m�n�Y��"�Ÿ/{����
n,/+����򷒁4������8Ex�d���]��`-䋪��\U�狴�5/кG���|�JF"��Q�j�e|X��?� %#ABgH��,�*��%�D��N�����`���S��Z4�$/��4�=�tfd_I���g���q9�cuj�#�$��uT����enl�H�96y��<ThK��D��w*Tbw��H�týL�b������)����(�DGM=_3���!&qP>��Ҏ��R �)��u#�/V#'+���z�t�mz�D�}h�@��ʥi��Z��"ސ���A-�zO��@��[�s4�+Md�q�U0Ϗg
��>y�GI&\��t�>��*ɡ�z-؂%ϟ�5
_ԶmŲ�T����Qs���6M""m6���b�7t�v��삨�.w�5K�N��-"$����Oi�y�7�@2��)�1�O�*eܰ���p]���<{9�]fR觟e_+�&Q չ��p5�A�a�o�z���3���K�Ǳ�ER���U$S]xѧ��˜����A�H���jTt,[��z)�]�O�I�� ���������V��l*��pk|9���aMy�����q��A�P[vӃEL����A�db�p/Ö�2-9 ��޶b����7j�n�7��ڸ�JEZ���C����lkM�bKuG%�J���=�eo�G�b[�h�UM���Lu*s�d����>���Ek�6u�d��z2��!�I(�<�Л�����t7�S4V)��oE���{D�����)^Ї>F|�����
Mz���(�t��FSy��Ҵ1ܯrVt@
&��+q�9��3U�	=>�uNO&�ZDi	�b/]v�CF��k(�����DV��_��v�����Fw�v٠�'fm�dX֮+���bϤ|R�
�d���ڨ$y ���S}ȕq	ژ��c��7JkA����cs���PV6W����C����?������;v��4��2�����
��͎֕����S2KD�!������7�4���#�֊�t�����-@�b�#a�-�,��*�i{K�J��8�MMs��d��%�{MU���%�������o�nza̗�GRQب�_�,9
�SmI����o�q><�ƱI�������3�h�u Ȼ�@��Eo� �V(�����;p�j9���LO�6C2�g��-!�Mn������t=��I ���a�ާ;	&�wTrbtH��X�4�%�X�C�vCX�P�����s	]�BばtU'$��9���Nw�+�IX ̡��e���5��tMꤞ�v@z{�V+1�B�g�ũ�����+P�q�����}[Ѽ�j�� �����I&��9�'ꂭ늱���J�2��}/6oF)V�]0m^�B�i��/�!1��Uzk��#�ȳ!ĳx��`u+OC�����{�o� aB�I�s�)�`m-kA�����ի�W���4�r���Ʃ3�x�. #�ϊ��~���t�@�'���M��r>�`����9����a�Ŧ�%{�ãD�z��2?g����k�wc#�k�ء���ɸQ�caW����.$\�I
x�qBO�'�cZZ���ۍD..��q������L��+DT6�Or��ߖ�H�����}���umY��4�&�]������v?�*��T���s�ۑ>�}#m�?���*��4��@���JsĆ�>9���*�?���3��Ot���C��|ND���o����W��z�QN�FLܭ|��0�wܫ�G�4#Џ�}z�%���vx�>���'�~@`�9� @+U�}�~mxJ��d`UZc~$^�7�nTױ_��lFU�O#�Fg�E��ݕ'�H�^��Q���z�2������|�k�����4-�&b���υ%��5X�8"�y��$��&���Rq�}~,�M J�UG�d9��}V�a�ѿ٘�ς\3Ǜ�@��%.\՞��5�B1�e�^������a��8����Ĕڶ�O�c�u+���#�xp���s�+"CJ!f�x��"��@���x�)�^q�%B�sA��r���EٛDΣ�\�؇ԿO�(�.�r���1�E��&=ۋ<:wpKJ�q{��b����SJll߶����F����~M?���t�鄴O�N΃��1>F`��>a�ر78���b��%��;�9x��n���>~�jȂ��^P�zJ�vX�y�˂.�a�3��aT*��&�~No��ܻ���+�H�X���)��+.�z\PC�j���[� S��k;��\1ɓ$��ǰ)+�ܠ��op�(�g^K����Ψ��{�*yy���S�O�PTd�^���N�'"�n�$&��DĔ=d:��j�l�F^�+b!��c�E��qR����h�D ��>�����j�B�1���!*`��t�.	�C��KBj��cR��_4�`�xA$�w�.��Hj't�R���	�{[h+D����ܰ���i�[,!Pg&r*Z��30�q�o�T�~?�y����+�ᵬ�>�Z�o���Xi�pJQQ��7Vg�����YE���0�􁻘ƪf�����bv��u0k���3��u�&u����˜0Ȏ~(<"��dfT��Y�[�����:�����S�����B`����A�o��㟡�D����,+��)��±�6������ȁ���e���̈́TDC�� X��JKq4�����ݠ�O��+����9/G4�ʡ9��m���/���^���յ�nc�a����ِ�ٮY�x��˷R������+�E�ׅ7R���z�D���ohW���fg�Xބ}@L_4<e�o]S���l���.r#�`�C�Z?@Bm�`��'mT9��m�u�U�ǧh��|%(8k�+Dg�3ͷ.ڧ3�0uW�ӷ)ֺ�v)˟I�Up���j���j�!�Z�#i,v�!�?FT�.�`0Uf����m$����dUX���cqe��q{���#LS��e��0<�3�OmjgAi&�����2������D�5XAH*>h�<�+)��8��K�l �cL�� j�ձq=�����{i��e[�m#�%���6���%�����C�b�W��$�G�j\�H(Ŏ=�N^>w�g�	n?0�b2(ݙ!D�(^�i.�d}�DeIS8K-+���Mv�ݳV��˖h����h��"�3e�n�E"ᑋi�nG4>;��>�}�d$;��{	�lɷ�ǴB�6�?LQjO~�G�3���wCC�O�§�=sWc*z��O�����V��s���<����ԇ�*6}� �;��g�nظ��j2C˭�h�����3m��!��MuW���H��]�i��*:��;�G�N��6�GX��m�-?�q#TE�?�zm,]�DZ1<�hS&Q�՟�둬"����Eص�P�_�f�D��t�7P�������D�NY�>�zk+1�o��9*A�ͱք��<��؋���?{ÏݙY]�%?i����A�ݏ̛b�z��Mq�q�Wg;���憑
��P��W�e{� K��S�ҨCߜ0̝��,'-} Ŋ=a�D�� ���aT4x)�[�G���̽L-���>�@�g�K�Kܽ������Éz�Z�QJ18���`{�=aQ/���4�W�q�Fk�Ù�4v�?'X�dR�"�m���$�UW⾼�2�Z��?f�����#{�]IEf��_QB�Y`���鞺�Ȭ� k��*QD󯌏��+�&������0V,���e	}\�r�"��C�p��UqyGp��Ӭ�K��;�:�h��ƶKU��&��s�����&U�Z�T�ީ���7���N��+�hA������⃝ �N�'ǩ�*���g	Cjy�� ��,�o&Q̄xv�k��!l+ٰ�t��Oig�&��3ex	�yݫf����j?�k�y��#��s�gn�!{�hq���԰>h���wœ���{
�r�����v�z��ry�l�oe��H��k8p�2 ��_
b��5�y���B��=�8T�z�مF�D�4|J�߾Z�����Q�N���	���1^�nJ6����h�7�"���&��H��mL��F�o��d>�=^�3����l��n���	��V���H����"k�ِ��<���IZ��hF�7nxb��3E8�3�L���F���U�J"_����}b+Cz�F£Ư�h�,��jR@hغ8+�����qlԆ�v�����N���$�9���q!�i�+�_���a�׽�ڏ{o;h�m�4p�s�ŋ+R�t)Y��"� �*a�/)s�&��U��o���O�	��㫲��H@@\:���\e�\1a�a��\�� ���m��Q�1bF�I�z����F��n�����X�P��n�s�)�v�ILf���T���~�v�xM���@!c�hBݝ<F���8|�6�^5;}t(�¼���m�UZH�la�,~�x�����l����+ΫoH��~�g�ރ9�X��͐f����赡��3,]3ŦM%ś��@?���==w�2)�Y?�/��N�Y	. �����i���$��A�$M @�{Ɛ�-����-K���
��]�ų��:�]Ֆq(}Nz���N�IC��g��[,��R����V��������H州Q��L�{<ǂ�G��IF|g��Dc���G�!M��� vd\�Rx�kN� Q�3P ���r�	G�Nx��P���9W��@=�[���h�TB&��u^p��g�{�#A	1e��&��/����y�ڝ�s@���m}>�FA�k(�]��$w�MC�H���ZӺm�����|V�hK�QO;�\�m��/���[�`�AY�;4[c05�L�!:p��Z1'F���Yvx��븣M��	�B�﵇��ۣ+3��N;�D�eX���$Y��\��`���0K��
9�7�W���`��c�v&u%����Z��Iݦ������'�NС }7��-�
XE��?�-�N��'/���������6D4g���@�����~Ե��;�(�{�����v-&p���b��A����7�vE�ݡ�ޛJ��b�DJ7���K��B�`� �F�7���� x3��Q�#VU��r^d�����cq�!?{��psY)^���S�?lv��p@�v5Q�Z���՞�/qX��6����q�x0�u����ϑ��5��I�a�Qn��š�H���TR:�jl�A �4B��c��*Y;<Gii��X����pslu�\B�(���I��3v���F.�x�ۯ��?M������Urc�@�|<� W�p:�̎ $������?P5q������#� L#��=侑+S�|����v���.˟BS}�{�b��'Ř��y��}���i1�6p��x��0� *c�������e�ڀY�kR!�(\qp���h�vR���J���<�<�"#j�ZN`��;����F��hHv�"�r1^�J�Q����0��������6O����Ca�4���R3��Fv,���߇������.
�r8w�a�7�0�|vٳD�*=2�|��zm��ݶi���T���C0�S��,�aJo���?�S����� �*��4�E3�.�v��5Z@1�X}� �]>I%'�Xy�&��)�(��j��N���G�I�d^ �$�=�H[Y�Z�GHy�k(�u��Ɲ���+�%8��I��T
@�եrCb�a���>�����ܧ�Dx
�6�D�*A'�x^��_��T%b����N {������gڻ�.��t�z�n�&$)dt��ėÁ1�"������ �T#I�]��`yQ���|�1gz��2�zZ(-Ot����aa.]���͔��L��R�6\q��ؔtg�������{��
Y�����]<F�I�o�<�;�K_��\��_�����R� �U^4���R�x���`"�^w{��Y��ƅ����`��s��Ў����[�wLv��o���0���z:��gJX(��8��/�~\U�x�=&�����N�:�L~�3PO�S3��ȕW��p�l�H �鍷��aH��i1�ɥ2�����d?�Q�8��+��$�,8t�z%	{�m*�Z+�¶�L����@��0VtM���xP��4Oڵ��֌�߄��9�����K�غQ�9�@�ʶ	w�b��(�'
�Wu�1Z�M��5�n18��W��{��EI�g�&>��0���r1�G�P�^ɲL5���c���8�i����&)��k_�� NdNR�*�*��c�D��J��9���#�%����sX��2�͊MX���Լ
'�}�2��t��R��[b�l��ڑ�!�J%"�M6L����#��?f[U/��f�y+A��1�����p:ϟ��nN����窋𲎻M�9�7eOś ھ~"7պ�@ݪm����� �E5V�
�jѿ��6#cm���Z�C(��?\�_m3-l*�=�Y ���R�zaXrJ�YF��iq
��.��3Ϝ��Q�hS@���`�d���+y��� �S]q��ګ��GJv\����c��	�YY.����d��A�����M�]����q�|e٪�8��%��Q���uĎ��̑�	�����KF�Gti6����:l����OmM�#Vk�)�
�K��{�WuI�W�il�:�ƊF�ң|�����N�@o�d��s��O1M�� �?f"vn��ͯ�9y��˨�r�6;q�9"pA��c���Rgﱖ���j���2ٍ@z�M���g�b�55�
�7f�ZCM�u(��xR����I�)5,�F/`�)"�`�T�#R�L�9;�����/��W�[�y�٩���-Þ)U�Zv˸���(���8i{67T��s���2�䧘}}U���Y+Z�Io�R7�d��@�|7F�F5����R>���6#�]� �7�c��ϯ��ׄ� �������}�Ȣ����	�Ӿ�/��Ps�sT�oi�3;~�;���?���1_/��<v4�*,����	�>x9ȧ��B��cƪ}ɄC�v(B�9�-M�����U����q������t�h��J�a|�����T�|�S}�/�a�����cI8�����q=t��ɺ�m�`�S��`謁>�h�n¸��}�$���=B�k��̚+�t���	�f�����������6��
 P��p��֬�w�_[~23��ƫ���w��{�Op*�]A+�3�=�:[��h�^,��R�I6WʟL�Q+;8�f�4�iMh��Ʋ��p���xV����h��/���:���x4�7�ߺ����,���жՖ�u���o4��)u-d�Z�, �={�lE�j+UՑ���q�S�lFG�~G+2 7%�!�d~���r} {�E����>���?�Ч&��Sz���gU����Iy[tv�+�CDY��4FX�>��0�_/��'�S6/]��_��M:��ֱ<��@:��~r�����E�Éy	M����o|� ��J]���M��GR�a˱Y�l���/a�v�b�rk��?Z��P��Δt�EgXS��(�W�����<���$�*�#d	�[��F�%��HL��->,��Cw�%�z�AR��^l"mN��Nᾰ�v6�|=��2Xl���dAr�QFz��Q=�Pd歨�Y��?�ו��Vo5+�ų|Ԩ�ۥ!f#NUF���Z|TJ�s��!�����߄��I��w{G���k�y��B�=G��am����jB�4��rIx�!�s;��|.������_�/��yX�*P�h���"(*�.[���iC�}��qNH����p4���䭃2p��ߕ!�o9�uJ�Ƃ3w�H���_�P��ܰ0�iC�����7?:�i���3��*���'���%�ӂq��I���t�k\�km�ELk�f����^/e�-G�4me����/�����o2'\=�&��Y	��Bg�ƔF峲�qp��نg����&gᕂ��@��L�*~u(]�p�aԺ��=\�wT��$[���7V�/B��|$Y��T�Bf�_ ��Wa{�j��SF`"�Z�H4�(i(�8함��`��>�I_�g�R��H&�X@�"�Gz��ty(�[L&�3q��4�|!��#��9]�g2�[�/ T�@Z��.2�d%�}���T�V?H�C���,KZD<���EfI��E|��M��9e=�I�q�FMvÀ�lFn�F��_Y^ ��wJ���%!�F��#A�}r�{��؝�1y��E��8M'�n�p�Ŕq9+<^�����I#�����Q�~��|z���z��mF�u��r�S�{g��`
2�,����r�ތ���\�z�}hX��+��-� ��/��$
§���ڎ�8u�I�s�e���:�@�i��:լw"p��	�x�K?&�����`LtQ9<㌁<���Q�^7����P���[^��]����]��-�eˊ�e�#9�s���䶮�;\�CM��^rv�/�`m1P�{��j�8y`�E 5����#��I'�������Xʟ`$�-}i����%nhE6r�5���~�S�3��`Բ�ZC��>_���'�d�gFѶ�su
R��9}y�r;�y���u������ķi���@�ܼ�U�ilz�ҩ?2��G�}?C��r�������J�=�0��)��Y}�n#��VױGM�B�Ȩj�T���s$vƙX+(�=�ڝf*��T�$"�W�Id�~���O�wp�Q{��IS5�D=@Ӽ�V�Z��!&`��A�˓��������2y�W����%��~�P�N��@HG��fb���F(����*���p�g��k!P`�PY0�r�����-�(7��`���!Y1����RDvV���u����;�bW:("�LC�u1��A��.o�]�}{X��RI��b{��7���$E��i�N�L~)r��)M�	������5I-u���Usm���������_�h5$���?�Z�bh��Ҷ�l-�Vtc�YQt�G�O������V����.;[���8s��%�S ���!�$Ш���w�sY��HT6�iu����?����;�|�'�o'���ε`9,��;�#!J �U< �@���������t�K:�����{���܃�w')CО���CJq�Ʒ�)53��A�r�a�����1��_ۻ0�B��j�dXQZ����=��C��4<���o�������<�wq���� TW��@�n2̾󪢹��q��`�����C�<�I�MX�����˛"�%���x�f�%kgX亁9W�w�Yk�D��y���/KIA�Zԡ��_���_��Ǖ�A�%ǌ��*'px�vd��b�8�-�!�R!�@��Z��)�%Ұ&��&M����@^)���⛺>�d*	���Av�o{�~0:��<&��*rگE�=�I��(((q�a)f��Z$u��޻m@��$R���iM�ӆ )D�)ѕl�X+:����CB���걯�jۚv�;�NQ�&"����e�D�s���9��)61�4g��
�I����u)���.��+������ٟP�����c��oh	��A7/��:H�����$~������輺��G���bP���9�H��5��)�fy�(ҕ�ߚY��-�r=���,��L�θ�w�&u� �h�����(�������ʱ������qgXq�A��],{�7�?{v�E���,���u1`F^��-nO�yoé�1(hk����ӭ���̔��w�l��gq4���\����?v��萏sE�W���s��*�h��(�[����gPP�]���W�ɋ(o�,��P9J=sP��I��7>�G�����&R1���e��{���y�q�ӇNT�'ZW���7R,�ek~�i�c$V9!����U��{�kt�������t�N��aRМV]��r^��ՙK@kc��#F�8��j-���+C����'B���Y�Y�e�Dg���M,\V4)% �^SQF}R�o��/:4z���ؠҎDt��%�|�B�i> �(�p�0JH(p��`��_{��Ά���A0�'����ISD}�3��DV�B �檀i,Ŝ�i�uvVk+ĝ˻I��y����8���n��c��Qa���)w�����P�_�5��W؊+�W����ͩ�Y/AK��i�^�Zϳ��"I"�mε�s���a8fy��z�.�J�m��dHaMYb)b^X0�l0>/^����z2'Ou���.���ٗ�vng!ư�_"M2�x~�h�����_6xq�r���Z������v*���,��Zc�.*K���lJv�F�5�_=ӱ�h���krEB��Դ����N޷T�����&��LJ8��p	)���O�e=�C�:&d�aP�ԌI�;`�E��Ж���%j��\�3`��Ĕ�~�W�Ԝ�d��Y���[X0�N�p�����ea3�Co.p��ke�l��A��"���b�<�\���׉N?x��TYRza�M	;�����ǁF�#mE}U�������8�rbdb����j\&S��y�R�i*A�T�8<�)��"g~y} &l��Lo���.}� .��9��V�7{D�T�i6~���cey�sM�L���m������BgH}H8 �jfB@���i#$��[�Z����<�쨭��Q�iL#Dq�M��4���R��QȾ�׍���*M��������E`��"�Pv9v5��T�
5�f,nףM�_\���ҋLǆ��dK��G\�j-�{�A���! S���[�v��:��ְ	]C��.���Z�;�w�/�|���a�����׹��E�����֢r��Db}Y����o�/���ҫu'��l��4K=�,}��}v9��c���"�,���æ���dr�0���cưǵ����AaS�;o���\����C l)<��b~��&�}�Yˎ��,X�5,R��N�\��� ���X03�!�_�����^z��`��K�*��b�)(d+��U�C�"��ɶ���|K�'$6ƅ ����ı�2'�[2NJ��1rv�������KPZ�����{}�.AZ.��&ڤφa \��3L �|"�%��K�s���F�z�p�S�FڼfF�4R�d�% �,�۞seʛi'�n/�T\�P���T�hm�H��~J��"�nPa�PG��c�����[J��vc�:貁Q����i�lM�QBwV<���9B?N���N�."HM-�`�gc�޵Zu@Q�� �ӘSG���JO~2}V��6j!�-_l>��Z��!��h��ܠ�7(3<���f�"��:��]u��Np��4f$_c�K�K�'�Wu��ۓ G/ɚ��[�D���b9p��V�(4� k7C@�KZ|�b��qŜ�x
�i�g��C��
� 6�^Z�~��E��q���E%�>OH�"��%'�z�!�|�S���(?���p��Im�Ob�Z�(��5A���X��e'�:�ICy聸E=�����,v�Nx��O׍;uf1��\� ��>�=�EO#���P��}z�����6v�ʲ_��;!��|B��9�qqP
������jIu�g�pk}mdw�c��LgJ���p�1���4E5����c���/V��߼����4X�[ji��],<[�)���īq����n���W	��I��3S�d<����B�g�N��-*;=gix� >��,w��Li���4��g�a�������o��P[�v|i��b:�Q�����L-#H�F]�O�]���� @F��]�� ��@�c�`EzKzg�6CJ�A��`�3F/ރԮ�e�����3y������jτ8�����|бin����Sw�2fO�dh�t�,��&�y@�jZΗ'��8�]��'��~o����Ç�N2��m�X	7�R��u���֧L�5�����ؙw�A1�iaS�{f���4��7�iBǥ4!ǃe#	 I��&��3�.�����I*��;�X�N�d>����?�r�5J�Z�叺%��}�	�g�!�L����5��1'�i�2��Ӟ��U�E�`G`��j gP�_� @@�"�u�xTPӑ���]��ͨB�������.����Q�͔�M�,�`���_�,�i:�}V��n��q�>DD�n��=;٩��_-_�Qm	&�J�b�UK�L��t�#�iv���S��"�=�r�`����-�ovڡ&���r�|��7Dsa8(?��u�Våd�9�Ē�\�i��u>�	�외㳝�]�����g��� ���6�|�h�.8"���z�u�qxY����9֎����*F�)VI6m
ׁ0K�`O�[�^"�&r,�nc������X#{3�U�mrf"��<6�q#�'�M�{�_�#�U��f�Z�%�,�47�<�K�L�
Xm)�u�'O�1W�+��m;��h>��k�+�֛2�>NN�mYFU�2?j������(�O6��G�A��gjqs�J>Ug����E�M�2}1�M(S�<�N�� �!?�'���C�3_���]}��� ������6\�V��Ud��8�\���z[*,'/��v�7(�xې1j� ��F�
��d{�*c@�ϵ)�������ז'����E9���/�5�Q�T�#���	kC���U�m:�%�3���>�8:������6��/-pp����&���{,@�x[c.�cv����tW�לY˴ ����H�F=M�Ӝ���^��w�A�up�Z'��:1�6�K����ݠYX<@�Z��)̬d��ͨb4h����]ma�.�N*7h<��A46(�Ɋ� ���Dd���+�,LFZ�ث��b�@��l���{��%�/��F���6��v	a:&^W��L�%7=�>�#A��F)g8c�p�&�Yhq����6��i\���U���ކFt��h�*�?�bJD}ETX(�����F�e�ʠ6���q�j��^(j�"�
��hNs��K+8��,*�:��>)�ܨG|���=R�f��,��E׊	�(�2&���7� 4�溹�w`����U�T7�ݽ����P@蹲s  Jv\���/J\�����a�{���Y����.�kj�E����,�E��Û�����[���[.�	ݗ�j�K^�{f8�)�7���q�&��\Oo�q�EXz�4x0��c��n����Pc�V��� �
��3'M��У"�d��ȼ"G]��A��l��f1���X��,.�]��a�׉KT�H��@���	����;�ͳ�
1���D�|eG,�#O�W�D�[g���m���ؙ�v�zUø�����.{�s����L��TA�ܹ���O�H	��e�|�����Є�ʁ�p�/Z�� vU&��
#>UBN�.Z���T�?��r��-Q�,��6���b'@!,���y�ㅦx�b�L��� ��W_8u���1������1�1��C�� �D��sS���lL�JM���0h�
"���c<ݢH������'>���A�V�X���4.8�������ۺJb�b�Iep�o��n*\=���]�A�����x#nM\��̱><�MFŪ�s���f�D=f�|��Q�"�5/�={�K9�3�`Xy0�O��@�g�%&��y#��P��!b��C�𙸫K���(�RV�C��5ۜ�!�FG{�I��^�����-R�Vv9��6�I���f�[�{Û���"��DX�����1e�0q�ǌ"Q鹈4�~�9 <GZ�J\��9��}>'��g���"��G�\,���gm��6��Z_&=�#����(��D��t� �J���f��
�����TX�h*:(m���C����8	O�;��k�3��RL:{qi�W������=sS{�;h�=M���\�����]xSV�rͳ�A��[hE7��e�7tΖ�A�O��*�ٰ"y�]�o��Q��Û�Տ�}4�K���-�������U7b�B��1��%�aL��7�s�7`r��/����3�ޔ�M+��+,F��sy��ڃ�I���З?��CA�ePZ�-�,Wc��K���Ax&�+sLn\"��f�W(�V��jLzs~N<W�:���"Q�Oj!� �ZW�N��6v+b�S��*�w.�_.,m0��D��q'�(D�t�z��x�����6�&BW�;l��ކl�;S|�Z
�!�0R�=n��=ޡ&���Û�X/�wF{{6�*]�YM�&�@�|y(����D8�$h;��=�ʀ�[��K��JG�VT�Б-Ÿ8؏�.��'��X~|�X�-I��!Qr��v�2���d�>�}�"7���
��q�Sq�7T��'zo��1�s���:%`�6����˯!��k�eD�N6@�u>�M�} $�'���ʴω�� ���*����n[�S�O���a�3�Z�����?fF�1p��A�H:I�Ƴ�No��