��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$Rx�y�<��wA�*;�x���@�̦�W�X�fa�M-$u����n~�%���P�$��W��kYَ���P7�?UMfT��q�6�U��k�>����~�\N�(�����X�e���/6U|)�X2pF�]$h���d.���9E�g�����	bI�g��ȆDE<�篙qU��ٙ�����`�>��
p��Lż�u� �V�s�{E����E�E�wi��(���T�ǿt���܌����Wv��jՌJAI����6ã�I�A��0R=���Sg��CO���Q[ҬU��2eh)v�u�JL�P�;���0ڵ��}�{��� nYd�K3,��  ��m=?@ჵ`���XG5�w�?�p�y�u5�)�4�o�'� ��/�z���:1��p�o���:�]6^����c/!~����V De���@<I�mƮ؃�hj��t��7Q��N\�t������wG�O�W�x�U�����<|/`��b+�8�էr�c��~}�8�n �#�Z�I1�I��르�f�L<u)̅�Pg߅-���$k%c���؇���.Q��3Iq7#��ز�QM4�*ݜ�f��=;ǥ_y:�K������8�.'5D�lD|>�%��)S��h��s[�خ�8a��d��|����s=���X��]�&楺jL���1�З���
��}W�"A]�fF�ˬƛ�  '���4fÐ����u�-��XwC�M��L��DEP7�85G��2s�bpr�h�.�M�>��*�������E����8��E}�#�:!P	c5fKj�T`�Lxb��чB����O���\�*�[Ǥ�[� ���:%���Ё\� ����2Y��$���,�Y�ۗ�A�A�x`��#v����>��:ܥpȢ�XLMW�
��ʅ�&G}P3�w|mr�>v�� )�����%H��[0�A��֕O1�D�#��pnf�b���"4 {����&���\�?S��kU�8-����p�xHoޅ���.����LB�ۅ�}��إ��}���yO	9*G��8EυS�׌[k���~�yf@J������Aȑ��j�6�W��k�GeHxR���v(bxb���$�g�3 *1�F��;�Z�]I=�f��,j��{XC0�y��ps�z'C�}Ɖo��퍋�j��������kS �
_["�d����^�Ӿ7#����e�r�����)��Sf���T��>M�z�	���h.To;X�N��r)w[�
"���|0�+��+ �	`&� �l���دY�i�8 ���NP�S@���g�NTet�����G�PX���^3;�Ă5�ģE�0옡�Ҭ�ښ�XB�2NKn��D �0wh�|V�a ��'�-�l�c���7�ƫ%�Q ��4E DsJ�G&:0�`@�Ƭ�:�E�aӿ�y�@L"�c�-!Ξf`�L�	�z����s�7�&� ����փ���ga?��r��`��e�R6]��m!I�WE�b����C���r@Xir�Еð
�d
��a7�ǚ$�C�x�a��I�t�\�g~h�v1�h2=9O9�QE��ƺoũ��
|��Кݙ�u�%P��$:!��M���*f֪h*��E	_ S��ڒ{(��C�(5�J4jF����vR�.�E{�pxF�w��Un9ٳy�L+uAO0�Wh�:#����Ƶ��`��&��M� ��%4N�b���U?�R���n�����։9H�>�m	_�Zn�4'd� ��:a|�lW�R�=���;DJ�L��v��][��1:?fνR�����,WTj�ni��-���ɪ��֢!Dn �t�ocGw�!m���	�\��(�+LH��ҙ_���l���d�D��;�r�8mj�F�I���ս9@�!,��4��B�44���2�Ե�|ˁ�fw�?��:,�Z�l}�D�^��a�94��Ix$��4!�سo�>���+�Gǐ��7��i�ڪ$������D�q�TG�θdO�����6D�gD��-^q�i��sh�� ���*��A��� %�-��HǾ�-�.#�va)7~F��Ǧ;���J�ȁM2�.z���B:c��+�$��<U-&�n���64=�r�c

7�ׄ(��Ag�3���I� ܍OLa��8��6s�"�f&�Gj�Y+�L)����T6�ҡ�E��ׇ�߮���T	��|]`�85��{%�H�I�B�~���GØpJ���{W[��g�	枭�q��'�C���M��Y�VW^���`��X�@�R��:e��� ��8@�s�@k��)c���f=Aî�����NJN	B2�p�%�MؑZ[~3�HM�:Y�~�N�n��к��f��trRJ�<VS'it�.�� R�u.y���F6;��I��g�:S�Sґ[�R��C�U�� �qB�,���Yu0��P�B����P�8�vzSb�¾�N~tz��%Y����B?({=w��d���}ά��.}x�%�+���?���2�a���T��7�΅���c܊V��_מ23#g9��#�'m��ڊy�.Z��'�6�BOĽ��V8�[�r-ϪET�k��U�n���JI$�&���t��W
q����U߁�:X����>�=���_�9B{k*")�_]*��s����#��Z��t[�)���?���϶I(�LƎ����n������q�i��~�n�I�*ZM%��Ƀ�6�\#L!�1�p�&�V�x��;21$4@��/��d�����q�S�L��i�4x#jۭ�}tA(v6"$�G��9id� _چUT�W�/��b�+UL��Uq���I<	k:Q����/ ��K��U�����M��Vl�$�XQhEԟs)���.��V���ӝw�{�c����d�ɧ�@�������h�#{[�(}]Ęi��ʸ��˝�^q7��nw��쩭]���Bl��6t������Xt�,�Z�iFe~�y���	����B9��d����ߏ��z<���+���8�4�;�{��a��o�Z����5�_P�� �]S[F0�:���\X�V<���X�L�����H�2�@
]y��_�=�� �0� 5ܓ�%��g��ı��b�
�����jP�F.�|��.L�A|�7(r=vD<Q4Ǐ�f���d����dj�ʠ�>&Պ'r��0��� <g�*���F��Nn9A(M�(��)���ϧ)���6���ԭZ�g���2��2|�����se"�R�+��찡���r�ܥ����r$�y��OKJ�|f,m���3J��;cT\��I�z������@;|����aӶ��D`�0�[ʯ'���ۭ]�gp���a:��6G��J$�7��Z-/��\E�B�bR��e	8�P��+g�u�F�X�#�s���<>fh"���sJ�Or@�0�_\wB5bS��kg���YNv��o�6ʓ�˧'uq�k7FW��=�Ʃ�*�1�+�#h�c�Ds�q�M7�H�����<V��<Ȥ1��!h�i�XQqe({�"���V#�đEρ�s1���m�����YC`CQ Qvb�R*�����s;갚��G�M\�0dQݸ��Sq��9ܴ˞P�}���ۣ�<y�G:�*�uȌr~��籹��!��+tk�man�Z&����KD��v��el�M�n�N�j )�T75���?�Η<�t��b��B����J� Jx���5���9�x� ^�R\Bq��O�D���<�u	�
�b}����JD�/W��o�����-J���]��t�)ZAw���0U4��O끨0j;0���9t�_7"�
`�� ?�R��0-:1w�KՔ�e࿻$}#����'��쳓�����<jtuB]�<{�|��J�=�2ў2�
n�tѰ��u���9����UŅ��#�Ar�L({�������.��6���`)ʣ�C�9'��he���@hl����?�a��o�Sݼ�B4,6
���Q#{�Šn��r/&�х7���Kf���/�A�Zt[v��G�cJ�A�J$�\�9�h�hnBMy���"�25��g6�T�(�>A����S���C�U)G&�q޻G�`���r��D��ʀc,Or�.C�����{�� :3y�1�E��d9!�R�$J���)�b���i+�8������@_>����`���`z��y�Q8������?�9�θ謿*=�q���F��}��BR�*���9y���n��e �x����@�O�����
��k��Ty�#�<,N�s�"�a��!'��6��-�q\��6�B䫛 ���� _��Gǹ��E��O��lϠS�ټ��,���,
���F^O��[�_㉫q��z��ɩ�-�M��F��k��z9"�-K��O,d��RR�P�Bccr��t��ny���$;�����"!�
3_���N��花�����h8p�� hP��+�dWc:0 �<R�!І��{&��O�S����0���3�d)9kGZ�������	:�<��C�	�ю������;�ز�;,p�W��5b��=37���\u?�����Uľ�wzNmУ�D3PB#��,lw�TBjԔJO�3#��0%�L�V�th�?�M6Ȟ�n��rp�"���|���/�?�-2W��5�@7Q�����M��:���Z����J���Ͽ,�џ)�>��{�\�%D�w�ڳÑ& M�5�0R�J�*I5K�9ظ�6����x�o�V5��+�!Y�����L�J&j%�е��
EP$L-f�4��v!(����i����+Sk|x�\�wo�Z��Y��b��u��U���i>�RBq>���E�����zb�Fh��T��Z�QR/W_�+0Mj'�^���X�A>ji�@y{g [�l@��JWo�o��."�*�G��C�y���Ğ|���\5|o�<��<!���gMq�M�#��C�a�B=%�n��x!<�w�E�m�����1,���؀��uX`�`���L�p�`�DG���C��j���xYZ���h{��浩��j��0�v��j�8���[Nx��qS����:��$A�Bg�ٔ
"����9�(b�}�{����}�J9iP��ոY�z
8	���.�}��7<���6%�C�p"���:�i��>�b(M�_z�.]%6
�+#Y��˨j&�D���<q��#���V�W/Q�Q8F�j2�������/�77�(P]jҀ ��)���Þ��Qu�����q�f@u��`��6�]�Ҙ&�fQ��NK����C��_�y?b�J��ݭ�48y.�wd-dg���9�%�@x�H�t�O�����%gP܁�tk���Ҝ�6&�kJt1	-_��%�u��;k��"5-	AoG*�G3,�8�	�����B��T5�c��Jm�j�F���W&��|�T�cLw�-	����ё�������ͮi��4��@uBQ��Μ��*+s��Ԓ�6V��SʱP �c��_��l�A�5Ԟ�׸�,I�U��ZY��?�?f]�Y���Z	S�Vߝv]�4�1�U[� -$���7��S��%hz�`I�%M�G&�4�ڛ:�p,�?�
���P}+���g������ǒn��+U�b�ϥ�n���4.|�l��iО���!h5JK(�U?tx��.�k$�ʅe���[�Y�n�aQԥt�j	��oJ.�h����z��;��ֹ�e���f�)|�ʚnF:(�*��c�:�B�����ug�r��Ő�a����YH�l�cG���W9 .`�Kf	aHplfƋЯ/h�[�����"�������!`�+[����(���XkW��Qǒo>Qy���!�&�(6�ҩ�.W�m�j�~?OT�mi�'|�}���'�_���ن\Z�|țPv�`�]'ʚ�z�b�Vo�]��#s��&Єˤ�/_\�V,QJ<�0�_4�q�i�"�;���<�4���{D���ŢA��Y�]4� /DH/�/@������÷�G"ҳ��������'�<W�n}3��+��	�XS|`�{�qDB�6���O_�XL_�q �����4�+Z�ȹ�I�7`m	[�����6̗Ϫ��Z�F�!��q�k��*h��iqlܼ~��x?�c��5�I��#�)�>��5��P���Ia؊��{o]�m��S�s�zU��ˡGQO";��B��Y�u�QU�ܜfQ��`$�#9�1���a�T��V�EdH��z3v��b�EG�t���>5�՚�#�|"���Q�[@&d鴌��P�?ˢw
7�JBH�߭Ed��GԪ0����ډ5mҠ�3��.�V��"mץ;�k$v #!7(��k����/"4���B��>T���M���[ɔ+C���C9/�~�c�c7��r�>�A1�4����3�z�����c~d��풥�?�U�u��o�R?����enY�:����7���*�U*�^�\���P��І9�j�ۇ0��z2쵍�v��oO�݉%���%����e�Z����*e����wN2a'�P�a�J<�m�l�>��/1�!��8e�b�f��a(c���BX� �'D�\x�2l ���4��i��}��L�����?�K����9��vCЧ3���t�[h�r�|�����2���VD:�p�H��1��#�R�I/�m��V刈v'�һ+���Ԣ���L���҂]�,��5{� ����1����.9�m}E��8���p��Ғ��?H������U1��i���������y��'V�H �9��Hi�3�<���Z
�lQ/ �L���*���S����Kgoh7�YcpTA��l��4j�'.���j��P��}mryQ�x���8�u�w��\|)@��O���x5�pa�*����ZZE�ȋ�x��t3�,����	�'�4e�}��?숬bt-2��b�sz����)S�������lG��O�,*� w�Jau%w˕N���͔���:����	Z��������	���Cj�r�^V��O���u��^�q|%��%���i�oB�n��pH�S�ӨR�RZH��,��W��_�$��m�tW�rcy��ٺ����wGZb�|�H~��-��]�lj�+0��^$�'2"��y4*7�!R��f����tb��~u>s���6xe䳕I�D�����Rd��a��-/��j�/��"�>:HJ��xw%���	�#۴7��r����<>�)P:p�&�N��lb`�XMyvv�%���sB_O�f��3���ү�cm�W<�{N�����*�+3��ǙD���5��ާy#칇�{(�F���M��"�j�ś���i"d���C�Ɂ�ԛ���)yS�{�
+�ҭ�	�aF�5���./C�LIzJ�[�ӷ�N����ӝ&c��iݯ�L��"Ujb_{E��z7�#��'�p���7im�>"}<-+{Riփ��
���?C��X�~��e@�&�65�n�f|�������L�yʌ@5���h�Q=娀�(�y�&C'M�#Q�a4��6JQ���P��!�����h�}Y��rc����4#$N�i2n���P��K��VE�L\��UY����`�q� �j4;��E�ӺvD*�}=�.�:�O�쭘-�s�#����ӓ����H𔟝K=}f��n�I��8����Wa/�Ҭ*=h���st��X��ލ�o!�2�����3eKn8���[�G*}��f�g�	<7�]z(.T��O�
r��M�x2����*:6��)i͏��Fus3U:TX�ah�r�u{����̏�+qe*��c���
l������$�j(Rr��3����Z)�H�Y�$�>?��O�����ЪYY/,寬-�Tr냮�����6T�䌆�uE.��!��Q�S��eK�s�{a��^?�yB���l�o�BI���(&��ﱞ�� lo��HUtY�`�G
b$q<��ۙ�(z�-=XD ����&��rl�_?�n�O��j��TM�� �������v/�^��� |�C@�׸V���2�'Yr|)T��4��߱��d|�C�-T�B��"�9憽��U�pA>.Z^����)d'�|��8V}'J�p��kA�yߝ𡖆T� ��&���p�'!��>�IOd�c��󍖈���)���S$�"�F��(�~͝�e)�V2U�M�x���K{�8E�S$�tp��F�#�ضء��}7֠��z�����ڱU���[�/<�n�v�������<����b�ٴ{u��I�x���A��R֢J�+���>�{C�/������<yr�a�?�(�;Wf<�Lc��ӌ}��ӽ�4	*s�!�8O#��\�@���tP5��8R.k��)
tw�a�D⠶5��>�wY�� >���m��2���0h�t��k��?�k쇄����ؕ�.<�ŕ�}���&Ce6�y_n�����%4:�U�y����{�k����m�al��.k�؝�O���޵���ܻ�#��G�2'�ن����TEkl�q������^^��Y�r��cE��A���'xd?�&��9��ׄ{�-�mYz'��(�B-���{��̯��o@�S�}����ɝ�v2	���uF	�q8�'U��hCG��O��{7+CY냼�<!|N����N�9����4|�-q��(2�V39�=�<���Ц"��.J����[�n^��J[�D�Y��ߕ��3RF��F��7����t�y_�woa��_�J�kF���`�h��}P#���h?��X��B������g�/�����|�1L��Z���|��ź&�"���'3a
P�v�ԫ��ӧ�CJ,�#�r�Kv���M��(k�g��a��y����r!E��!�����<S6$ds\5U�S
U,� w��~����.��Õm`7�;tx���ؗL�\�?c�6���F�ʺܠHEd�"='}A��S����۪ؤ�bJ<�K��V$�#)޶W���]�E���s�����e���	}�Q����þΛ�����{�J{��H��Q@� �:e��ʰ嗁�E>�W�����������P�H��1�x���"x�x�N���������.�y9c�Ĭ2���Yg5���2=��ٗ��8/����韀F��Yey��x%�D��5M��3�W��<��z������+w�힅��L!�s#�HWź<���ɞ+}�c�jS���\�J���d���}2��#*�9#bQ��pu���W���
�[��� 8
J-Q��H�^���+��m���ud��D�4G��j.8ٵ�+k�t~k!`�W]��>�a�B����!��N��m�53��"�!��CV����K�a_���&a�������F��Z��׉X��أ��!�!��H���E�c�Y��%W�!���v������5�u�X �@k^�<s�B�#e�]��~����v��*|��*q#<r^��Ko��o��,|֘<V	oE�[�\|ojX���w���o�� .�~ F%�� ��{�$h���ט]�س�r��*�@Yr&�����%l<�C�lb�P/��,��lYݨr�A�U���C[#�ǳy�(�y�?�H@zT�%���E��9�GT�>����11a}v4�ۛ�|���Q���W���E��:��l/�X�J�R��+�e4�Q�R."���KАket,�ޗ��M}�j(����N'>��f�Bu$����ˁZ0�J�Njf'@�U����f��O������?ᅾ>�
cӬ8�1&�1bW�߰�"�� �D'C����K��МI���&(�@���A-�s��u��l������~�P���h��O��?��U���_�ՐBRMc�2B+��K�*vY�,�jz�U��$%"k��툨�E��n��.T�x��1��5N�Ǘ�j��@����K��B"�M��fJ�-�6a����iy2��)���'gd0�Whn�t󋗻Y9�%��BZy��Bw�1��	��i`"����:y˯�y �cMʨFhJ��E������
�K�����˷6�K��~��͙�~?�v��K1�hA"����5$�*B����eӼ	è��[H����B�S�ϫ ~��!Dd��鴑ဝ��6� �|�}��	��<v`�[�P7BNDb�bu�d=_l$�.Z�	{�ή��OC���N�i�-����AV��"�T�._�g%���#���`50���_���o_���{�:�F*�����@k�,$
���^=�Am�g�-%�S�\n�[�2RÐ._�\��H���e��y�L�*��Q-)Gns�d�=Ҋ���ɘ�S��ɲ�J��=E<�^I��Ͼ�*����?����s�:3���y�f�~�5��ʊsZA�a�ߔRr�\9v�9չZ$:|�iw���Y�d+7Q�$��0����vvo����&D2�m�sV�g��s[���Q��*Q�� ����4�.o�2c���6\ D2KA��l=���=4B`"2,[N����1����3'�v`�x�
��6�$��G��7,��$�0��|�`p,��GZ֕��>�e���0���m����7/�Y[;�0*`�v�@��	����-���"Y�����f�M�gi^�\a/�ƻ���I׈_n�P��i>�׹��8O�b������1�F���:�|@�f+�G:�Ô3iWkp6uƇ���^�s[��u��/��V��<]*;�&��[����*�Վ�=�G <���6����pU���0��&������
*�X�~�Yr���>D�o��%}헴��e������+0�6o[CHߝk!!ɾ��d� ��D�,�yJO<�
!:�>�>0��&W?�x0��p�^{��e��F/sjN���5 q�89é�I���7,u��=����&G{rw�.��ü&�dz,y�cQ?�?�$�ê�bɄ8[Q�6��4�$a��ie�|�Z�T_o����<�G���;�^�I`�\t�BF�CaOo�⽞��@N�]�b�zx=��WT��� ���И�=�gZn7޹�������ӌ~��;-]/"��Bg�9��p�'=�z߂r�-7h���ݷ]�g��� Ҷ��|w �Gz�Ď
\(�G??���/�z*���$7	�){�'x�N���U���S������%�Oka��d��6� �ʑ���69��0@�� -]�&rQz���ωCpK��VA���.B�x1p�����LRb��b"Y����N' �N7�i��d��Ə�j�[;�e�a*$!x��\I�Ht��&��-��lz^0^�$�Xm�?�����<:�O)(�̱N�aᒘ-<�nY�{���ʮ��L��k�j��@�8	~�Q�W���V$kǺ�=���fE��Fn�[�ҕ,�����c���7g~$��F>�%�	�t3�]&��"3�b�FB(
�<L��ROU�F��d6���d��F���d����{����V6	tH�fP�o�tWn�Y8���Et���{Q&��-Q55=n>$5�L �{��.��䰴?���m�-�`���G����)��ǳ���l-Ik�`6*#ye4��\f�@�0$A�����-�k�+����R��E�� V�ylˉ*w�xL_f�.S:<q0�t �0{�A�p�.��o�N����3z�s3�@lz�BKq�FZpd���/�C&�C�Ex��ȱ����N_Y�.���&9�kqJ�?C���ʜO@����pǪ��/��]Oow���O�$h�EWE�6,��1�������^���M+NuSV�J���#�k�L�䒽����t���SGm���2®���uɂ�ԟkT@0 E��*!C'�;����%�^��U�ᅤryޞ�WS9`�&jG���L��
�7�-9��C���=