-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
NdjvY3uHzii4wkO7O1oI67vZCracTttP4hVMW6U4fZ2uhTzyCxHD9msfwwRcMTkuAqUYIaU6bOID
l9+PE3cSCkQOn2IpvIsW0M4Ahk0u+WsWKKVjYN/ibbNH86O5l7QKpzkCAh6U4mQud8IZUGRu4n7N
0O3XI7b83pUTPSfqWYPyBfNrtpD+Qj/yX65NtJGvkLHQL+v37NaxSQkxsTv3UDgMTfUbHIV5KfWp
k+iseNc5A/58AMv6LUvrTJjxVJEl0gHaCrxfXFgTfdG2/EuK+h0q42R/MvGvCYXzv2H64x+ZAzEu
JuV0j8ILt0h1qxIZ1GMUr/7NpFZw/jPB8KFL/w==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 9424)
`protect data_block
BR95zhRJoDSpkAH2AtUQTRT64Vq5E96ofJXz0034pD/HcStOiBR63kQhI11OLia3L3nNDrmVPs90
AJBYmY3H0aeoNvir+NEPLNz9mcFnLZwD5mHrPgi0UIQBOVk4yp8NbBZvtQPDM1s8F1gZe5/OZffo
e1RAJPU0uOnflQOqqtiX6xwGaJVWa+gbtW3i6eOfEvYFZiIMXUkMBzYPPFvT7bd8GiLX7bvuRQkO
YiP95g+oI/ueY2Ry0DZj+z4wOwvCJgCHGAC898Jv/lo7Rko08+TUrueeVC/Z+NxeqVHoXGhV5IDd
zcaq94HfUP1Fm+snnp0G4WCKD6Uk3/2jvaHqn2sQ3KzFy86R4xFT19DhQiHmfg+qBQMJurnth7Yg
OsBZ41njc/meK32e7fVhiIXMrIaZRtQPAEg7lIcpVDgmAvdrsOm2YceFUs3cT1S51ron63gtw0wO
mYEdgwL3DnzQIz87m5FWlBMfgGKecRiqRg2ipW1VKKhTp0/vDTQ376W/OH8iQ5TFwe4myzMV8ckR
4Opx6UcNKmZfnKAU5zoEyJXraPgKgcHL0QPhhmJPdh+4RipwS9w/nJwYGc1hM+A/3za5xXNN5+8k
JfSlzACF1/IHox8zD1UxZ+OnSRxRQx68Y8suPl0C8beeyzoaXDKf1JjtqCw+dTioxExvjCm1q7QV
6NrXfBmNMK8nda/UJTXDwtpvEQVuc2tkibaMsdLjCsmbJOB2LF9Aw5dxruKwx5XT4VHb6Nb0eNx9
gxwkGwReMauI5ntRerjJkEKflfEfNNOEGBLJ3jMMz6sAlwoEApEt/Tu5FwVcnBfrTnXXWIbjqY9i
8YuD2rwz1IYTOqfcnd5M3eCIOAsDkEgpWW6fKI2qHWn8EVlYFLliqUfFVxoRC+yOGHE91846uINW
PdYUYJ58IxE+UhMt127WlyW50lJIRp5RmzsU8Uq3MkpoG/81xnk9t6d48oCFOMA5oqJIZ2BOEb+d
3Vh0uVv4kcW7bWm2RjsTENIMKXjq6QpyL83VkrJfviFcpulXjJWjheq16GzwAIDOLIsL3dfEF7rC
Rd0R/d8+lud5i9acvB7gOfX+3VsscInBLKZSfuSBccEuLGMlcZzplBpjEvIvwIz3LAuPYal05dA6
vVvev1qFZg+pfSO1brPw3Y0P5d0caXFBwM2bYu0RIT72t8nKKsTleoL0tQfspn8HVS3zxkovR/N1
LI1IXtV9vvlsQZ7ENVF5r3+un96pZtOaf/vUF9Snt98I3VsmTDHdQO1Qv9NtIlKhy0LN3eH99ezG
UQw3t7J4FkYV0UU9HfbThVgHmuJf5eHsDG+QnEsFwe5C7YezKN8Wm4yrxwtvApiHQC/p/uEvEHwO
Xj8mFfl9sTl4v/c+VfD/sB7K+YD3P4+iLCwS2mL2r8df08zwzcO7CD1iAHpuwDCSOfT9D+GWWIe7
L36rMaELMDMCoVgoj1Q4zRjAYn469CrRtK4XMc57/RR6uML536aeHB9ip2S/sSVEQpE5RtnbBwmT
FvwPGrakwNaCikgPMLzywtI92fapIDHbyZEXCNhJgjLnEHZJu5c//BMTcdJdsa78uFhoYSTHtg1j
1ror9vvgdoVqDhzeHy52VcRJrGt8/6xI7ZgK+c5v0Isk9ZCCc18vi3yA5/N/Ju3vP6Fn8/US88m2
OoBHGHxFPKj1e8xRz9jGiOJ6ntPUSILn38aK/ZZ65wsiT5GGkMLGUqBCmeXsZUOD/S1Ijkvbzv6F
YSZbCZMLoqi8qqF68kiWBb3vy46H6TX7v/dC2mwAxvZUJ9MBkzZHiKXSgJ10jv3fcS+OpOdikJn5
4awnAJEYSDr1de9/QLixbqLQCgdgMDX2GqDNRZ0iQHEj/vp4I/sBTBE+JAo1Uc7gsXXQYKnml6aU
ckI4ec3hhXcK9xCu2UmFuebF1uo/teVGwce9/GAtkD7qA/4WNIqNJDXHWa1jGmG+PP7qq9viSOP2
YNk9PAj9FqfcLF/wEq6Q+BLoMggmobrOloLYvRMNXxOOfRT7fLbJ0O5XfqmxbnmSWC/s69PUOntJ
P73OeyvXjSjuGmnaXCfpsmtL874d9uZ38kpP9Noj1jSlgLVScEjO8NZxZk7I30c4cuKnMKjCA2PA
XkAYDwdAyKMg2Tw3VTet35/Gm/RywNEHVcHTAHPW+6UoFOXgvkmBLuby5HVffBPHVEaqJsqkms2j
dSJTTXDXyde2D6Pe/AJX5ExgqH0uAoH0XF95SFHND5Gy1940hqY4wWnx56VfIfWqKl6LMCQcTl0R
KwQg6EdF/rjKqSrbexCwaSlPsK/RjFCGTEZWa6vvSV9VaWAANq8oNIBSjPpNVwUWtr3mmrnX3Y3I
3D7NgN9W42I8wNV8peGAUmbrZgdurgFka5WRvZEjyz61ss9yduyx2iaLsDeYpKKFDO/T3qKFVMla
PtU6Io961JddVANuSMBLPJMbUpFS7QByctjxOhRZ+wFXhAFKY7hCwAmBGz8F8qYfrsd2EmNGimlj
jO8ZkK7GI1DO8Qsmk61M0Afeo941hA0oI6m1mSL1fmXTHNbaV9i0g2lj++J5awtFHPgsAbAd0+ww
sUFonMJs+0iFWgre2PUK/0786Kp9A2Z/uzI7R2U2FckRtaLSbD6L+9TOQhnOtvdUJEEysRCmel6s
9MU1uhU6peDiNcPNsVbuPqm2pZPWQhR9plj07yDWbm5hbkmcDB9N0bCM/3P/G/VXJkr/8J0UE1Np
sNclUaGaRD8ujXZRKAUidGGNvd2lL2dwF6opy+qwRfX2eLXRwQDvGMVeG0h4VyNNxo9MEvAYcLsd
6X5/jNY/PzKgQiG1sOzhKbaA6Jpq+5ab1xM+6+56VsFnfZzCsGF/hZpMVTnBUjrOP1SPJUoKFphA
31y+xxeonAXZ5DWZTnOfbsOm9jWIt6E74fMiE3KuSr9N39lz7Skn++dKtUIYT/EA/HEpor2pRU71
gEelRYa35MEafrNeROqcRQpHHoBgDa/HKSABLamtXuhp26FYKXt7vk4XfwFduVdVTIbEFS7rlyvL
1HVkZ+uQJWO+QAsmIZNpIop0WlfCpwooEtV1U3UachNdb6wN6kSfx2guECYQI0RKJ1YV5umZBLb8
OJAYHJ3ZuS8tDLL/Y1K0rQF6UMLx7SCoJd591WcwlD0M3YS30w484cd3g1rkyIAlAOvbQuq63Gqy
MkHWZ4kEO7TKlKJVr9qvmmxNjDLfOKFApiqnKYq1IOAkONtCrCIaHJHxRqhfqlqMkQfWftXM7eUK
/+Yk+HCtSPVT/fGZ34ItLFthee0UYIV9X0e0vGIP1Y0Ja1W2MF9WdcPHxXkNxLhePbGS5Ksvz3sQ
1nUrVlUTpXTCR5j25DTEj/KCIL4lXAPZl4a04MU9N92zXjWexxd1CUESRnA0YgAxVasGys9lYADZ
FOdm/PaPqe21G2gZfgyXf5NZCttS603wzpLgvrSIDF52L9mtCIKdKtZKEzSTHO6VNvy86RNNSdiq
RPGdYhmDWVEg0pmVe3vAUmZW//4bRlYEdfI8qyr5T6thhk3HKsSr+aBww5v6hFXX0VXSarpdE0xz
BkqCon9wFuB0IIuzxzg87nAZiedKlZ3mnYaWXD80TOaZIpyLvsL9DTwGUTZ/7I6ofLsddTbzk6BB
m7fzRJsp6W1ObFNn6vzDdfbNkDuMZGKbLrcfZ8cUZJOabOjMbJyKWHQv8Bd677Jv61IicuEr7e9c
QsDk3cD1rmQlfLeNjhGwKiIU81F/gPzS1B0zhpRK6GAhLgXQS/7yDEuc9HDHuEbW/lzc6A6TE7aT
8Ph2/8xzCyz9/PmP3KULqKFp4QWO4TbolziiM9/vXAn6Yu6bn9kVVV0M/YjbUghoqp44zNjVaUIO
kWC/4Hw4WU4hS+eYhA9SvcgoDnJ280yOSgd27LDLORfK3MQHvBBgHtYIolV5/12EHvz0Bq/Qnc6p
OrkRek/2eroQ1egQ7YleIa8ujUb1JHQjXzcIWHUVt7KHH7bi46K68/z/YhqJFKSx+djXQo1sk9Lc
hK4gN20ESRBfOpx6LnlEdY3kxzrxee2ONNSa27VoHuWY3Mb9nzKn430DVEXtaNLTmxpmJ040DohD
N92vr1qekgqCU1TWWvgyZgPjZ0/C57MlJ5QE7UrLGuO7Q51cs2E08KLdV0UkKlj3qcH7RSlmS8SH
WvSBNQ4SadDN9yWQVeo4F6NGgye21yPXdBbMF0vo1QOGDA8D8NIzQUK/5/JdjueonK+WhAw3+jcd
AI+T/sL5/oSV0svBkiRN/Y0CDoaxRibAUGpARGkE4LfjqY6PJMfYhGLKptJo6ncHQXLk6ZZcBxM9
fGFtLr2uWi9DfBf9wjTGW73QN//xUO5uWgvQTAEgk9JaF45CxTO02qEoVNwDqTPPDWPRGjZyW15K
HrNDi7M2nKUxZsoeawYegB241PA6hybrRcWcdCabsSwnXtT1AS1ztvMV0Z0AQ0417ACNc/nq0XuL
hZuqw6yNKBuPFOXherp9/MW3qxbqxJ7LxuM3e8NSPtfkuABkrFkXPvU9QHSn7+Jo1fnCTv7KWPzb
Ti8wOcsLTIxrBumHhSLeng44m/KWJ6/Z4logxXP9WLzWr6DPboYSjDqFwfifIJh4RYAr4+CYA50i
Q0YvH70r9v1GxC4G3ePzPUYJ8SY2TnqmFvfVkrPKWkF0HRu1/zP1lSC5Z1Yw+5QGM3PzKhzU3gEy
OVfP3Mvw9VGRMvheyVhPkdVSWozfxEspOcYVlqFhhdfOHsQ4JhLEKBlx1somlOWs/HqtAUDfW3v+
es0GOJPqO4Fw422ORYhJQ1GuIxJIfS764utA/1Sbl8QlM7c5o3kK+NCxfig3qWrGf/9jSdbLd4cU
E5aVq3t0xQjIoSZAAZ/S6rb5ZMau3IAJ31DPwHLn0n0ciLSYOtAjQx/YA9/Gf9OI6AB84JF/vvuH
XG8Af4f+16ci5TTQNhLKJukcJJPquIjo+x9fYUWgqZDid8eiAJfZJR19ieTi4vitVdYV/wnFVDPG
WhHF3pOgjwXOefWPlaGhK3kOBCE13Q0PmGzJzf4UTDUuCLt/Ox7QjUMLJute78DT9VZNdr98tCBk
WFqhwdAfbONdbrCGSyRFTaiX8+aEthFhSdq+7uZyJ2fv4D51R1J0NZrbwMxhV7IkRUucjtUUeuA+
V0p4rjGgZCQPNhGwwTq8m5MHN5rdF7qRICVUinV0zMWj0S0xxgUMWp3HsxmrmibnkbLhOMKGgj8L
C8W/AppCqx0Ja5BqyTwsLi/3rYbzz7ZpqkIjOgLj9Gs15DjSQnAxxbQAxe2FvjgGpVC3IY3pitjh
XCL8iz8shAR4WCkOFFivsjE/YoJaDGp37uM4hIlB7L+x2QL5yrYbw1eynFP/yReRkv3s0NDKLv9d
6sCm5d18wiyBz0KKnPQqW4FvZGmKDo/0+7qWOnQPfafJAUcvS0lhLbMyWwd794NjAqlh7jtCUKzo
bgbUOMKpoT+m35m8p9Gpr7vPNK22UW0dia4FBoKuk6L+D03cxkjxYI8FdWcje8rDi0hEZlZLJqB1
VL1LJpBv0LgS7ypHs+ra6rd/3GIdf1sXDgSu0C3+W9DXtizJ3bTVVTaezKaCK0BPRQvVvXkfxHuv
AzD4PCOhcBMO5UuAH9qP6h1Jr9gvLRh1kfWTOiqSJ61MAau0YwdRGWGX1vbRMV0KczSOMMB0FsGT
5oJBv+13JwlcIZG9SvhXrt+8sUiA0b1Himo5GLgzQ517qfbFwkbMsJaZnowmn+tdXBTkiRSYGgbp
R/LvdqzhlMVmyL63pJDrF3W/5MnOcRVoq+2qdb1TxrK2l94MAb4ZJhe8i65ZiQDQPuBUlqa92av3
dXPHRBLQM+/5ScVdXXeUmbus6eNutr+w2b29N0BFkFliSZPWdpjcm0EgBn68yUgBPmFeAId9t324
YzamAO7e1JnVut3Yf8T0LOdcuhbmBMotMqUwSsuAnb6RQ/ct3ULoQCFMFDfuahkNXJUQhD59Idte
PocjZ2gYoegwD2aEuvzHl6c9FBXvjr9Tqz28LXDJ73yjKflieSePZM2bkngLM3GunQD8pj7PiqKV
kJKrKiGhEKbKerF2/hhoK/UKEXhnmeYe9gVYHWhS8w/IEpf6FN915S5RT7rTnKn+jp8Bi3cSIEpr
zofX35roJRmrBPokE+6T5Zp7XCB0V2EgyUAYUX7dsYycrTr0a3Pp2C43pal/L9gxABFHDUVd8GiH
E9gVEAX60fatxldkcFSG0kxp5D6ixKKKfYBdy2UvqORmwEu3mCbdw0P29gZbWobaC/IfeV8DbVOJ
y0Yq2bAJKjnGYSEXeaR9ztI96aEIkJldK//S7Olwkby34SJwp6BXFAIn6mGHxUcgDyaEReH0V/Uk
/MkscmmACJvK63GCtp/sr24fnMy6cbmxDnkO2cv0U4uoQ6XvoCt4yi86vsyPJw76Nqgbc33ksUI0
5nEbMaTmPS8VxHk1qdHDHE8OxJ91FbomsbmPirUOzfqM9b2XxhPV8+7r87LxQRDGJMlJMlKwf2NP
s9eKEpI1/xIq7ujcA3XDtmaNzFVfYGOQuHnRO7AoOR91+OjiuDOhGDunrf3GSQpadUfh4iqo4gx1
Cv0bMMfcqgL1sNY72gPNW6mfl9VUynsTEiXwQwcvlgZncVsLi9o53XTU5Ooozw4dgqWK0aqrhfoO
0B5mJ9bKohjY2nuaaFy4ucZbAxXIvXUY1EQ3Z5I7OCW0EqjyIo0EEIWNMNRxn/ZsS/1oyo9d8IzL
BA3CpODVYICWNBQvVTugF8ZL5xiJKa7mQx3Fy0n6fKTygZXKnBSG5b5ypg0D+LhnTlqbFBN/7vM8
CeoTAh6WSfi7EhPyewOakJFuKMzOTbDSLaOiJOL+fyCRfFLD0/g/5htPEVpcq1rLRNlGp77qCNe+
z9k35JHQhqeraJAPp3tZIZVxruURCdCLXntLqEsfsb+i3sZpSdOxWwDoDBLxMlOMxedpeIYhIzsc
5sLtBQVuqaUgLlqJa1KcAETxTeOQhY44PMhb47ksrzrSw4EWpgPindH72Byjgmm5kshm80Zz/mgG
f8ZlabHYreXcCLfxebC5tc5Kq0vHT2prkP9ZrKoskT01L0y/2x8k2gAbXEEwdelXI+ord0W78pmT
KXVCcxU2HiCEQS+Shddf6A5fO3izfMRQjOdV4bKXoDmLaZyMTOKnPzzWWUiZdmo+sQyCXdd5timp
NCd6Yh9HfvkkXlpAvVtuD+8FsH7ksM9qG9DDeqWTFiF4cayzoidwXYNDItO36StVtQLnkVLLVCAT
DvvGXQF2VcA8pC1svrU9xlXDZjM5KmueOKIJfHZwWDaUqPmXgzsQNMVmv9wPUOdTiTGjh4vFSgvP
EsLmhwddTAYTgCKTsLSsH3vaQpYqmVIuwb2Gl5tlM4blhTtxnTFJ6c5QdDe71XQahT4zzClSN3KF
YlMaSBQwkuVG+fdFFqgOnuybEYVmNXgtIlFJFMTm6+0EtyPE88u3QFF2XeqbLIEZ7FcNnDRvJbmM
RFNrnqvulDK9cUyh8diNYdlQhaUcB5gN6RWr4r8Mn0o9ns94HQl6/ud0ihRCr+n3JBvpwpVF7paU
chC2uH5jvCz/klYkoD4CrIIWtaLgzjAlpUN0MRqfWwIDKkuKi8f4cFsZuqxasnC+HvisVhu1Fuml
DXbTAbAD1n6jliYVmy0BWbSYmgZaGZmk2Vs7EbmuE0aBztVyJVsWnd+iqLdKykXCpCa3wN0d2Poq
3THXC3ek3QF7JcZBXI9EBgLhtfysSgMmRSzxMKEMFWRVnXdVkBEOpFr966W99PG7HO1lMnK/kunz
qFdxF8KHL1BB133QdYtGX5TwoDvh1ThQADgo6y1DfksjpINhwkdyLajGx66gv+5iEXiMYFyUEU4u
ovKipBjoaQFDfg0Lu46wXRUxPsWTDIWZfPzMxvw1pCvk8A59X8C+vHWtSDYke2pncaCM1tAGMKwZ
98AIQqN/bc551woPG5sGVa8JR1apAsItyVLX95dDrQblnyunSm2B0brkNjGCG4sBp3HUdxReDKTT
dq9mqTLIlWcmv0iEZKoWfo6XYUh+qcXgon6hCsPj/34SAzYTO725073Xw0kOFaTI3qXNTk7DGYr9
okVsHe/csErf206dN3zPdNzNJDdR6eQhUVVkJzm+qOGesy1XAfoz4KXfGVA1yx2iACO/J/B7cX9n
KtEyr9uXajTLx2a26MUr5z/ifB93FmgOVM/sf20IF6ilvscYLK56E0QLME2JKFAQPUQUZ2Za2Pnz
awfMvz0pWJZ1mEglN9j8IDZRTaQoxMzrkcZCu8mkdqSinGAmeTtXLIA6h2sYOkhTqqe88DqlvKJf
tWzUAvXT5LV+AL7iTlIWVKZTDZj7E6KAJXAVvWYWxIlwRjTmO1r1DbYD+8X9WODzC5O4/H7b+VPs
cwHiDvrY3C0uXz/OMUnuvfnShvRjW54fsG6zC2e/kUxwtAtGex32MM9J0QZBrXYjJH/ArYowAPm1
jLUdtXKcD6rIRZJBc54hYw0K6s4OBoszhHnvLN682PORSLa4uR8Ko+wiFJUzIk9y93KcOTEld801
WvOw7N9mr9U2cU3PjNgVq4HHtL2NQpOYIK4dXNP+kk8hOScVBPpD7hzjyeinHZqYyr1w50P6wksp
RmG636CvOyj0b32ZIAghVnFP7N1UUOlP/sLbaONgDOJSMPVcV21uWi61c7h6UBmlcMKx7c7hNM1r
+tUZvF/UGw2MPvZKGDbLGvI1AEVgHxcbNCSjSE6H43TUo7BffqSxzLDL2Ga0gRT/unGd8VPgnHvT
PNfX4Cw7KvMDBG4p7NgPD679pzN0222PtqnCPlO/wGYfMzE4Ind6I1XAdcrWmFJUvi+ZwR8OELXI
VbQqo0DdPWaOiiqqbWl2qGfEZi+lzOnWwKJBEA8SREhobyQdPuvZAfT9lZWe4TlKBq7Li19bXxbN
tGSN2mlTVk1tG6Fy9VcZyxmF1Dy+h8lpfcVnYKRgFFiUxxH+Z7NBzY/lMwaK3LKOQ8MHJK1oiYTh
5WxhAGmvIqI07eUaRmhgVwraF33D19+tn7u/+Xf2jrPDJj89GgI71J2kUJth7DUp0EWyzAXwKyVu
4nIZrvrNAezq+CjSCO1NAAOvejyobnyJKvy+o5W8m3IJBaeDIGWRV3dqVGG2mVyTWCLYSPH3gS/F
pezJNcjOTkpVsiePcxdbi+spg5y2J/PLQpkr5WaaM2K9vi8O5ngwTShJ5rMXsc+lxmqwgHi2Wvjh
KcOaALf5oqXlZPnEZWfkSPogSxslDw7bxcU3ZjoWfwHakJZv7GgXO7b3Ag9e8f4K6IUdGJSsDTpm
rIhKraxqz9ReG+V+FU3dT4istwFkfKu3ZHKJAlk1bkFUW0vwyaCJAPJezdBJ+qeUokHEdDRTgVIp
0UeQVwtpLuN4+04N8uARiN3eozl19Guilf+Ukv9NK8kLtQSXF7Urc1T3KryBdtjNIdvU1VbjDGZn
suZZyT6eQJsV5rTAWZN+0khFr1hkAstccaBPxCJ/hZrQH3wzSjopgqz5gweCwOgWuz5q1VD/faJ7
jkPK4L+9J7SMhSRRG8ACws5zAk+s3fGyYr8L54I1LSGKxpdBOTo5ryJNOg2LoO7a5GOdOBfdZrRx
CUY1ISNWzBAkOFFsPu3vL816Sshi/wMjmQZCL5qQ8huH3yaibshqqeomPuQO1hgFC8swOJKHqFAW
beKkauZ0kCyr/O76KRl1qY/oT+scJMxlNq6cK1fO6L26NzKpgBK2VfQn929VC7Mp44Z3l7O/U+BD
3tNSaUiG3f+8Ofq3L2o4zRrpNYW32aKVNr0yVYDk4l6RuRo8IjwyRyDh7lZ2/+OqIUWegJduiY60
Wb38wZ+VMUT8Fs7E2mhPGEb2xxcXt68HHAocB4IT4mhsUqM3RCeRWeC8jesYmK3aB/fgcFhvkDp5
Qms8XQr/jUk7DYV5VfVBADOPIsgYyVEl+eFdSG6g/yqwzto3MPKjUdTfPMTk8N28lly8z7BoZkfe
beNO+UReI5fSmcgSIty22MBRAnUpyFupob1saUtq1DbkHq0v9KwGECkekYzLpZA26V5jA2icvh+E
XrilE31cji+K5T4jaqE8K230c6/5WD8wLdXASmkbpORrA/qF4O3sUQt0r9inKh7AjOWKqGVw7qHf
FzSFPjIEPlLQBJZjJy0Yl5ThupDjFgFG0c1GiPb9Khhdp80cfnr3bDgRDIJLbQZuYQEQyeErjIiz
+xUQ4VmrOqPRlQzhRO2SwD/phasUzBEByeVvyrES6XXdIgL2xXnSBeCzuAV1xqvPctxrG29tLcKo
FUzOGAl7H9pQdypNyhRupyp1lEjG7FcrlOhkU4Q3dO5fZSXfZdpgTmnjLV8e2nqvDVr94QD7uA0z
f1DMJ15z/hPHWkRjcN3ObKQHsZZ8wL0KxFQRrgTLm5n5aeGo+4Sx6WI8dGjnfLtaWDRzVm1R4jP6
npuOpNVWEByobVdaiTHgGPvMme0b/fJ+NrLg+33lxOuh5Q+XbZt533UVrbB2HbQc/Hho5zHv/WGp
67jmzWj0JdRoZw7Ex3sieI4URpQbJb+OCrMqRTM9oGFg1dgSCe6nkta2fOWnNp4gOUWtA5XIxjdW
rOpqcgXsM8POuTkKtFN93HPKKCtwzv1lqxXVQFU/m0HT8ZDiQVCqJ4Z5eXsAeRCVVYotBbqnZhZB
h9cLlciG/quQmsbsy9eabjGlPChfiPnEWlgbsrAkIhnSKDLVu0T9WgpwV5xQ9gFOqveMtnZ0MMOB
zP/NQfH8i2E2xZtwaHOc1zX1jNtcYl/8bIZJMuqDF5iIUCPLzdUPxhpKi7V647wb6Dea/m8FYRwu
zGaAlUhOSt6zlCdyCuxE1eNGcYZUU+MXxQSp3Auy1rwu/cUSVlN6F32NhtwDSN76woGAwil5Bqjb
WDLoM9ArHQ4HXG+bqREIXjGOheeaVFLwNqQGJHPZH7qBWlfJkB5McLwVKdkCCvrlzPbxkbdJJHzk
RRmKJh0MFXtlDDm+ScIurjLa2jbvlFB/4JcuU8KpQTFrfYtxa9HhsSzR8filAq+4jtGzaYLGhyIz
IcowDt2MZHK/on99pcrjV0gwc+ro5AJXJ9jg47ZpiH0XArWDXO5KCiYTP3h2Naq2pSPy5A2/n0Je
+5TRKtw8oBh/ZMhoSJBJX2l9YGbdXF4fzr66kMSArojlMn4Gu8SC4G4Jm9R0Z9nbXQV5N/EwE4Rm
maTAlOrb82YR9l1jDwWiioBVvB+cceO33DlkpjpBsOeG7mHrxoJRSFk+9LgLO4933XjlscR/84aB
lkaTPvPSJJXx08g3FN+Iwn4ioYu7tHveUZMRqoVJDSfSWrdeyAwlbvuEczWeSEqXehWz+6FWkzVA
g/qLDHR2WrXd+3tqdKGofkmQux36n9slpaievwJvvHc6MMDnNOIiT8u+pAQp4QviAWP1ehAsztbS
l+T6aUX2g1im8TniTKGNCMIYWiyJpPzmJaOouqLT97Rx4w2X5gh4rIm3ZTbTVGOtYWx0zuNYJPqd
dwNDBn06mthG33JNTZ28SS6KEiKvLEe7al7DKsK/dNC+QZK8TGAqK+RD94cQSk2Yx74e+FmPn27D
TBBE++3sl5e51Nm161PscK5Iru7cM9bLcFOLli2JL8mHVp65X/qRRuxhCozEGnv4zHb8JcQylmEE
xk+wM5ssnwlTLjgIS1auCXoF6atmqie/UlP73QbSatGRirwIysJHoc6W1IIaZirdweLaDR73evGK
oZjWqhVnDG98Hapxsc7l1iROLZo5NiVy+qRuLX4nAsRY+DV6gFruUVzTKxnlfXLLJgaMjd6EF+P1
bmEZUh+hNhADrXvUnTfVMBiSLFj0FM2wTbcFgw2ArA0DUCBeXyuOrTzUeAXNW3tMSGbN88/6Xg8F
uKZbRGJSJQibYxHxWSzcPXfYqkyDijyqZ8SeCAyDoiCtp76nzQksBLKQnms3H7JLmF0X71M61qaI
Jh9prKJNKQdkQAx3+ocAG2h50cfpavZlrrdMAGeGhn0KoJBqJdg5Siy5zRJRcIt4g6Eu6H/utXOH
BusIjsf53pi3rwEkgk0G8iwPsL7K3KtD8rEfBpbUxZkNTY8YtEIkBeDBN0Q0DlRnE8KXkLq8aC/c
w/33Vwg7+0UlwLNf2HLw1MmlRKHfDcgPBqp4dS/Jvpm0nynHTfYpxFKMxxSFVmvqTSHEp64DwYey
ATL9em8XF9taXphfIqAq//MTJ3KT2W7SD+6poTdPjfAL/u0CQuEVe9phdSB5kMI4g3wOVQGNjckZ
BgCns3e9VHILsdYyN9T+VpeXO4bSZQcybIUjcIu4gWTF7MaWwlUSapCobtHzukb7ZUYckZRWNjb2
9vux8mtFYbvF41DJFIFZXIlvGzdUDDuuI5s7hiKPK2Cj1eZObvY82/8kVy5FK3WFWcfprwVXnw8u
5iBLOHfk7BSetTh7WNxxSfRomsp3Atj/2Y652ix0Zx2jQ9pKLxgohA63AihcESBSvlBuvzA6hU4t
sqKGMDVoeR4ghcWOzs7n4tfIxg==
`protect end_protected
