��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$Rx�y�<��wA�*;�x���@�̦�W�X�fa�M-$u����n~�%���P�$��W��kYَ���P7�?UMfT��q�6�U��k�>����~�\N�(�����X�e���/6U|)�X2pF�]$h���d.���9E��WG��L�X"]�Ad����ľS���8od����e�GT?y	7�������ݵ�^��R�q^]�鍦�����s�ae���h��L��P_���ާ��YЭF���'\��68�b�[����w8�[X��V�F�0͘3����q諵�uW� �h�u\V�?@��_6G�_�*�G���B�絉�f������[�G��U&�����~�F��AׯK1�`c��[<��FY���4I� �#�G��x[X�=�Q1��`��R>(�w����R�O�?����7�,(�H\�#h(W�EH=�������yq��Ѿ��aF����:�U~m<|��.��0=�P/���4ǆ���T(���=�ըTW�z���BHMU�+| �ڋ�݆ݜ,ü����(��pa!��� xR�'�L�wC�ʂ:�(FX! 9naq\Z�>m���)2��CE�* �.��*P��"h(h2���f��k��`E��Ⱦ�7Բk���_��f'�6��2�1]I!�d��*g�Ɩ:{�3ǚ}0ߔ��քs��$�����V���7<��%%�v���4Ȟ֌�����?�Ak	n�~V���'Ņx��E[�(������m�T>�ȇt|"� Jl��	�G���U�o�Rc��;u�/�C}�p�������?҆�'�����A|���)+����2'�T?����Op�c��-��.�eFdX���Č">ā�΀X��ј�$�$�S�
�a��e$�o?գ�\9H�?ފ����Qߴ!k�`G�L�mb��s)�1M�),a���]Jb�xy��Ӯ�l��}76�j���!�wL3AA�= y���~�XG<M)&HE��`\��Ʃ4�t�t.ʃf�~4x�H������(��Bhʑ1��>�v4�:��p�i��N�K�hl�v�XM��m灲k�k����}K?�h�ϾW�jpi�iy��7���N�ŵV���~\����$5�')b��� '-a����Rrᗭ��`�������d��S���/�=��^8�<S��+gg?����o���,�95,��*���D|�s�$4���3y2X��ч�R�|�Zr������t�f�~��Q�R@F��?�5 W�tmY>�=J�똈���ܚ֗!i��El?�M�҉���}�#��:L���Q�����/Ǵ�&#� P����\�;&:`����Dxh�{"�ã�hC4�=��6&;XU��3"2=a��H��d�o��D��S�x�-*l~���
�w��	��i�^�X	L��ĦD�%���x(�O����U��k=TH�c���uF�Ncѡ�����Y���>B0:`:_[�k�0��2ߞ^�Z}X������P����ߍ>��@�O.8ȫ�w.�JO��1=t��!��39�􊲼=l��������&���	�v�/�jwa!F���NT;��L��[�����nv�'�
�2G.{Qʰ�h�zE���N��W�R��	�9lͩ������]vi�pT?�����1��De����,�w^����X�ޙU������}�)�Ty$LeZ��s=�|J�gKݖ��&9�/�<@(|�H����� 5��7h)l��k0��Ga@#��<9�p��+n)�Y�h��fI)�!Ϥ8�$��ce��Eۈ���)�ˌjΪ�J��&VP�P�j�!5���@)�vn��/'6�m*�I�}�B6J�m���J�`�>���v����;�}����&X�R�eN������>�{c��>^��'�:|���˚'�Gb���:�Z5�M����c�[E\�̭���09�ks���߲����b*J� X�T!�2t^�2t�R����~W*��C*�)�Y!��UzE��}B���4�����%^xB���t^¬��DU���A�/��6�7�Ǚn�+,=�?�`:�#i�p) 
x��a�4T0r�^�(����#�$+=X�@�}��[�lͫ�D��8���@�r�k�N(�z��Sנ��{�!��ѱyf񕐗������X�ҍ��
��G-���Ha�3���q#ֻM�TtGH��$C���R�� ���<�|pÊʰ�'r�8��\����/����
��s� ��k��᧕��Wh�Hc����r��q�db&�����gZdj:MX?+6Hx�n'cg�pRf$�ka��\�E����n�$����S���g�W!�x���m�h�Aag���2q�.#HG��{·��_��Q�O�ޥ�K֋�MǑ��Gzg�j��C������fK�<������u���f�.mWu*9�q����N�5<�Q�<�<K��s%��o�4��?ס�x�#�!)bQ���뗼Dd��AaaL!E�Z��Bp�0J��P����x��'�\���Hs���]���wJ<��m���^9���`t��R�>�y(W&)��TԀ�ӻ���!癐�l��&��Xߑ���%Og�'60��<fcX�<Hj���***Aʢ#�v�����_+��6�=#��yk$,@�/%�쑧h�5
'rs�~�|V�$.�$!0��@xE@�;�ڢ���[������ä�ۼM�$UB�Y�Qi�aƁ�c%�H�:nw��y�����>��&^&�u_�R���y�RA:���W��&�:Q2��"��~�T	m�d�b�6-�E4��i�T�"�g|T�F^�\�u�*n���"P _�>$?����X��h?se��ZaGI[�R@u���C!Rw$}+G����c1_���/�{�V	����Zr6`�?bW
X{Jd�M �F" ��M��k{��Fٞ^>.G�kV������R{(�����V�ϑaN�����Ҋt}v-�>W2~t���D��~G�h���Db��f+n��sH�T��z��Z�1yd^gd8,4SSk��e	�׹t��-��L�d���߷w�����/Q���03N+����٣������y�Ƞ4-V�PVa�:L����:M-ш��L2�v��k��,�z����(�nVwӾYA���A�QP�ǃ�6N�Z���mk�9Qfq�+��?��0�����l�N�E�@�C�W�%�uMtA�%YX�E����&T�1\��ߜ=��z*��_�k{�Fo,�<���%�%w0�֦(�5�Q�ヅn�>��p��[ �_��:�5=�d�=�}��`(,��:���_�x(1(�Z���%��v��j�>�>�b������G_��@����cE���D��|i��}1M����ILj�̯�$����v�n��S�,X��9W2G��V^j�{���q��3,�5�͝.�Eyc��Y
_8���"D��މ��p��p�Ӣhг���^/�2���*U�$���m�7�Ë�&��`����)x����z�'.�3���@i���1:Rql)��p�C�y�I�~���p����0�-Ĳv[)���k<+d��S��� U�U$Vq�Ů^��)�C���׍#jt�-��7l�������P��c��Ý|�{q3�-DC�<��|�"[W��<YZ�q%�$-
̈<���i��*ICN�f��� Z����\���?����TV����^Nu{��f5$��P���j�8���}�?;�/V��w�������ln�]#"�{�:�G�$%ȃ�f�!�\�Ƿ�ch�&.M`�Z�B�{�J�QmUN�n���S?�4�%V����0�ذ��T�6��kz.:2��SI@~�cWT$9�cR��3����X@�'2o�l��:(�m�J�;!�������5��A��M�| ��0 �S@��@�^-��`9�D�5@��"&.�.�_	j��łܧZ���y�L5��T @kW����F�b�Eٯ���^��>1mf22I��)�l������2�E�3tkN�`[ѥ�iJ+�a���>+�GZK��.�����%S��tɊ�cWCÝ��Q���\�`TkS�l�?機�-$�8��k�_IH�~�c���K���L��p��=�ހ�"��{���Y�5����B�,M�D�pJ�ǒ�����@��~f�ˀ�D�_��v�/����'�rO���\�{K��͛�[<��w�Z�@��!����������Ұc���J�[����P%����F��kW-�3xF�o��s����K݇�-�̍#����F�v�a�[��y��(J����~Uv��ʦSs��կE�˥��d(M���x���V�"���jj��b�x��t��d FК-Z�a����",�2F6	Dv�,X1���&9�I$0$#1�B� ��l]����dUp���O�>;pS2�SXY-�]��	PYl�b� o_xfBp����U��:.ʩ�%�3I���]'��&D>c!�����1����W�M�A�4��v����<��}�,%ʗL��`�TO���a�V[���zc5�Kz��	�K���qύx��xi��b�ʧ�l �*����MC�n�4��ܣ��'UF��l`�u"���#e۵��n���#6 �W@x|��!�N��o�2t�~A"5��Ƀ�_Av{a�h���1I3�6w����!w�,����4���l�p[�f@g����6U9�	`B�ߚ�Th+�QD�Ɂ�٭��A�ɨ�b(NJ���#�+V�m�RC�J����E���<��/ʸ�-Ԥ\+���A<)s:��^�Xe�q.�ǘ�-9;��,��"2�tj����v�'C���u~s  ��V/}{��-���E��6�g�J5�<���6�B��"b�]F�D��ܵ���"P��{]:V-��Y�_30�ɼ=���b� (gU�J$	k݋��o�K�~����s�B�-�7*&�g7�]N�m;�hA��].���em��0iqP5���*���%+H����C2��nܺ&t	wAؑ����� G�WtrpL�Ɔ�9����48xU�F�%�5.��q�܀J#H����{Ó!��v��D��&t�.��)�ܶ�q�}�uGKkbu����� �1DCM�j㓟8�r�YhZ�%�*��3�C|�R��+��lv5
�w�6��њ����0[�W�^YISd�i_����<"�F-3�ݻv6��!O��n�δt�'�� \3���6ۧ[YV�H�4�FM+�{`"19�����Iir�;�R�ctERj���`B�[�!��c�8V��k p7�Z�|Í�ZY
zl�L����T����T�����r��R9M�w���1��B����X�D�F�I`
�e�86/aX��@���턞}�/'�h��͚�=ЯS�ؖx;4<���H��\���b5$� �)0��~� ��dn�����6�^�D�i�1;�_Ցr�<߬�ވQ���t���w�[���7U#Y����e�M� ���gkq�=�]z�����O�t)I��;Ֆ~����Ek�J�d����CI��R�<!�16��`�����
�06��y�g���ʴ�Q�L�ϖ�����i1�lJ�'�E�&���l��G�ʅf�Nd�ƥ�2�B�B-��f��/��	�G��������.b��9H �����OVԂ��Y��yt�4��%�r�?3����bNfQ��n>�h� ����Ʉ�$Mݕ�k>:p!I>,�;r�L����l[�-\�����Zx�.0��ٓ�I��͛k�:+E�lF�[�X��A1G)!)9˕L8�p�B�:�D�A4Bݗ��վ�[��
xɨ��gy�HA`�͓pΌ/~���]O��L����奎��&,��N�E��K�Z�̛
��PK+�s]+ȸ/iiV��b\�<��e"��#�����	�������Q؁�c�S-�~���%��f�+��9(� е�3��^�&�W�p���<*�����|��P��m�0`�<ݐQ����~C��Ε��給k�U�*2�bd	�}pd�TTr��S����+I8�%�\!����.�IO<Ùc��$�u�>���Q_o~��!�h���Ш�r�S#3F�hxYE\."a�t��[[4�XJ{����T���'W 0$,>��{�l�@;����n��}�4��[�"�#��3��X%t�c��c%�u2���%�s7a�!�ܮӋ;��59�դ�6���ȍ#j��H:wyގL.�����s����K�<��OߥH�A_
墍ּ�S��"@\�R0˿���C�u�K��G��^PK��l��8d�4ĥ�a��H�0	��0�~��o�����_��q��wv���������B�I1x(����
-X;A>k�Ӿ6��`�i�u��EMxa�d�?w*	bÓ?�a���N��r
��]-�4Q󖧹���U ʦ����+ޫ�}>@��=�J-y�jX�c�ʆ�T��fm}��?��HV�Q
�/;�R��9�S�$ �ia׏��	��R��9K�?)�h��꙼����Z��Z�A�F���~�G�F9��L@�H�x��B���YU������{�l��ۋ[��(��N�縉���k��D��R$����Xt"$#eB�����A��i���p�މ�>�������g��o^�[��;C�g��:�ή��l�qߛ!���@Q7'?j��~��_���&����+뮽(�L%FP?�m�r�R#�F���e�<0�D��(�5n�| �#�m��f!�Y\{��)]�M]Y�괅����֥Ť�o���@(a��N��N�E_�z?���4�Hk�;e�K���=EƊ�h��0g!#[��Ų��^&qvܖKGYz|����R�Ҵ\R�'�zAs�nƿ��ܹ$�3w�s��N����"��Ӽ�?+�|�X��AT�om�P���rR��I��+9i0�,ް������7�S�^���{0|�U��&�}d�O�T��';��z.�h[�<��b���:�n�#���(���*��hs	�r=��A�����[�����w������^sVajضX�"�%S����1�=/y���� ^?�^�e��IҰ|'	@D�$����Ƃ�\P"q�A�2\�g�
�_��G`B�|����?��*� �&o�"�e�3�ќs�=�T��"�ئ��`��id�N�g���G�zS�LN37l/�����[�(hO�bm
Z{��ڀ-�p��GB��p �Cr����D��|}<ٲ��AH�N�M�h�M��ު�L�RO��іih& ������G��a�aP���琒�������%3�P�%��ĭ���M%('$;��L�4���e�|K+�Y3�!P����V9-l���^X���~�<���n!y��4M�],j5ӣ+���GF_����M��d*�䠉��eDk���ճ��٬�c�~�j4��	��ZP<���0��s�(��s��ὃ��ѵ���>rBK:��>.�^�4ޣZ�� щ������ݫ�c�o�x7�6d���gc��ǂ���������de8?X@O���5i���������Ĥbc]YA
����D�̧�5_��h����_��a8���a/6&�}�RX�>�2��)��K�4��~W��MQJ�¯���9�cȟ��A�8��!�K��u������j/j0��b���ZBE#褑Un�z�3�`:��me�4�P�3�n�Z��LdQ�:�&��!��J�';�c��q������^�{�u�B�\�6�eؚ�&O��}R]>�Y<��<?�jD��]�2�t��ʠ���$��ś> g�Zn��?~��V�`2�N$�D��� _x�G��-�*��C�?�j�h�ZI��^h&|�A�Y������3�̯��'��Z�_0���%e�Ty	h�]/�x#�����_�ZR�\.���Y�v<�O���/<LT?9�w,�g����憕9�\C�����po.B�^T�[�-�7E��>%dz��vh����|��Mo2ˤ��P;�@�Oۂ��o�Y^@b^��{��C_㠙�A�?�7�{��>1U4��=�ct_4�gד��1gh�et�A��rdl5M�E�"���QsܻJ�iP���g��d�`��ν��4:95-�>s���q��l���a	�)Y54�B��a�L�i�����s���Nپ[Q�/$�3,�B�jmM�����ҩ�g7�m�Cc�L��{�k
�t.�--�2��b<�����{�Sv�}���щ$)���距9j���t��+X:������k9�����|�QSۨ�䦑��A��w
[!͌�2�q���^�&�O/�L���=%/$w���G1�~��.�|:�V����M�5����=���=�6�6U������(T���/Z+9��b�N�l�0�q�/�( ����O��D;Hl��x���5��kd4��0[(��!�-3����@����C����z}Jɡw���6�@�ĸ�Q��G%��b��
jˆ���a���m����Wb�}��ʙ�$	�vN�'T^~4O��	X���&�#�wй�c��/N�bHw4:�<S��lL����B����'�}�����R���̄���ֽ�-����>5�rBWE���ȄX_��i�����>3���lI!�������V��r�XQM��%�2t]&x�?] _�	z5�D-���Ut���h�EL	��*{���=��@��I���D����J�o�,�ɒQ�*�����f76Ǭ�,�y�
�F1�7�����x��֐z"�z��mU�O�d���ü*�F	�`Ә
�՘A�>L�P����?�u}-�e���/��ź�k�(M�rT��i����h����)�Fy�D7b���Za������7g����@��� 0��q�[���w��U�n��DʹEň��.���U��o~��Y�V-���+�b�~�<GcK�:3�zf�Q��Sm|C��_�	)\�X�eŨ ?l^se&�Fo��2����4�?&��N��V��#����ȯ���� �XoH$��lC�F~�zw�ܵ7�z`ňO��� �� ��C��vx�J��f)Jv����zh@H�?������N����";�{�4O��N}��X�q$G�,N)}`B�Ӗ���ի��n�][���}U,�5'dJ<�g�����r zE�H�p fh�o�B]5���̲��I��r��Ҵ��^���z������sM����.����n����U�GV�*tZggY�a.�`���	w�[�D�'n�F���F�φ�t�$�0��+1�^�����^��qe/i���JO�@U;�k�E��_������rB��7_��K���#�A��3#�[� l�	��=|m���C���v�@/�f9hx
�7�ab���θ�)����o�EE"�U1~�`��n��x�i���R|X����1�^�'���Dwl�a���<�}K��s@��ư@mWAq����C�K�gN��I�7��l����T��I�� ��n�gק����1�J61D����8� i��M��Gqd�B�S�c2�V+,ƟJ0�
?۠�����P���ip�:�� � ��տ��&�m� ��PccV6y숕�i������S.��l4W�����:Q�;����fu(=�¸Gӿ(��r&�]��P����nV+�Ol``������|�wm�������$x��>1Lk4J8WW���\;��)@4���/� 8�(-������%�'��t�h�*JY�����7�8���� e0U��Ss ���i�t�Xِt,Qq��ao�ek	4<�}��i��m�1ZQ�\�9�駳�{�э�N����z��:ۨ@)�xa`>b���/��7��w$�a8N��&4���a-f3� �jjN^!����jj�BJ�6��"۬��Y'�sIhZ��M8���t-z;���Z������Y.�
'�4���8: vy�8��x��T��9��,H�h*i��NSE�z�Q��GH�\��?��m�܁��.�=�f��[���� ?�c��]�S�/A�Xm�J��s3k5 .����a��4{֗�n[O��Ve&���h.E��y�ɲ���s��KuA��>-�9KEӒr�����-vEH
ا|�����R?؁�ڈ2R�t�i�F�� &����l�f�v��|I�wj��f� �!X�܀umM��<_��Ic��g�c8D n����U�)���q-˻��׍�@}-�k7�Z�*A�=@����|8X�+�3��h^f�#f��Hߎ�]�҄�Xr�jZ9yh80/�O��:�ޓ�t�����9>�W�q���c�`�������6j�[�{h��iӶ�.�F�v��S�M�v|�;ia{B�Ub��u�ȻK%�|�����:`G��r<LVL<a�'� 4V�f���4;)b)j�߇tg� �8���Pk}V>{t��i�Х��kI$�r}#U����G*��"|3W���ɜv4�j�` �!��}aJoQ>t%t��g%,n����L�L�h���B�a̼ZeKJ[�$�1���23�
����^$�a��]-D�Ɓ�Z����Y\l����c��φy��d�PJ0U�j���N�Cȍ�r:0]���QISA+�b���q�8��R)��� � �a.���ԣʏ|jC�Y�F�!6}���o�����FJ���Y;��5='��a뎇B7<<�M�;P�ZP�h!\�u[� ���i[Uc?��G&-�~$�U�g|��T�6�,oi
!kt4�N�w��d�[_����ψ
���s��~�3Ee�ݽ2��U�/���j���,x���;4�-Π��~��2��HȲ(����R,�5��񪖪�����5Rnr3U���{��e_��:�U{yp�GQn��%�g/_Ɖ�¬���,D��ºE]��ۈ7YEŕ|���"��a9t���\{�A�,��@Ay��'��_G�χ�A�C��|��bl^���S**-�sc����6�7{;̄T�쪬�8�=w��K��P=���{�^m�(�r��Lz�v���鸪��ct݀=uP(޶�:tg!�o*�߈F���I�G�`?jM�6C�H�fH:�����J��WǠ����ݬՈ���M{���$o�7 b~��D�5*N�Oe��g%�i{v^kr���2�  �`���P���� X����a�*p�Xc�3��rqh|`��^�a.����u��I�������9�}����d'�n�.���7..R�Pc���XF@�)�7ok$�V�(;U����D��Lݍ5d��3���*g1k�;p�&"_FZԲ���*�����4���
ǭ�6���t�\�tP/q���	����"'����l���Ҙ���ҏ&|-*~*G�}P��d�'�� ��Υ�����[ګ�.�"�ك7W>k��G5�)�
5��>aQllܠ�7�	=/v�f���3ȩ1��D�5�儍�?�Z�Y��Љ��ٯ��^�I3;c��7o��ЍV	�.���%1.�L�l-�K,���D�P�c\TL�z��J����nN�E�߱r���U�;es��p��Xd]c���T�M밳	A�(���[��zl�t�,��fm�a����SOJ�Wak+m���-��<G�O��w��D؋7�TD��Hɽ���+��B8�t9/iJq%j�
8��zD�Y������F���H
�]u�>f>5䔩��CSE����!4�������ΏU�0�Շ:�-�5����vU�k&yR�2�Fb��\b�"S��-d�������V}A4B?�x��v�ؚgW�W`�gw��;8�`�nV����ƭhFo��VIx��w��B�47����u�̯%�h��V�VE��z*�)�G��U�ȽA'�%܊������-4n"��F�ܙK��5�-`a�?�
���u������cB�b��<�����D�Z������t�4�<P�%d+�XPՓ�|�G}m~�R6�@��/�l���o4�uL$_��H75j׉uv24�A?t�7�����#�@����9'�.R����Be�g('����\�� ��6E 3fh���da11�&�]Z�OV�r�k������-#����`Q��\�� �0�M��?���4WV#�z�M�j,��d_�T���T�T�w Ī{5>/v�&���(n���v���l7n�4z�\B�/���Bb�Kt���	ѳ1�4����`�=�T���l*�T<�����{�#d@���g�	��7ŽQ�M�tW� � ���ǅf;c�����_�TV)|�g��y	<Rc�����������V��Q�^@\�
4�=���ҒP���&z]Z�j�8��9Yܭ2�z��~|O�:7>բ���������4lp!����d�6�U�x�DiG�zN���#���O0]�ol�w�E�>j~���'D$���\�4�]�p��?_�&/܄!>IfDz�6�v����*;4�k	׷�E䎶Xd�������*��2�v��Sv���e����Jӈ�U[�Nc��8'@(�m��`>!�t�\l|����):�Q�a���l��!Sl�4����k��w�E�K+r�ݢ����>6��oV�W�M�ˊ����	\��N�l���1�����o�u�o��X�z�DH�ڭ�_nj. �O1��6���k�u����%�	(����g��lk	ۻ��^�@4zGx$��.Rhլh���d2_��˕e���v�Z�L�I�(@��B��r��'��Ϩ�`�?���i��B@���3ez~��t_]��tSۏbl��^;��\��$�D"`eة��Y��\e�����v[b���O�a�-?������9BA'�Xsy�Ty$�5_1��%Υj�.���k����~Z3�|8*I�X����r4�S�q�X�����y��Np
��׳�w���G%�R�Fxx��	T���à��H��'� ����Of��p�>_�����a"{��'��9�:ʽ��^��).i�^�s{皧� /�Oh����[G+��]t߇����@)UˁSb��i�7���6�"��?�y4�>\��	X̄�r�����f��z��s+�j*���?m,x��;�j��yv�O�i	��\�d-VIR�+�<)3
�~![S�Ya5�cL̈82�r#;�� �`�-���>A-m�Ig:�Bb\U���e���`��n��m���$��Ъf*��_10S6O��'��g9R89(��3�
�S��)�}E��g�Lm7kl��Je�>�$ۏ(cbK�ZʒM�l��9��sR�B��T�ξJ[)�V1E�J�k���Yh��s�:�{c9 �|H�Q��Gd����{h�o-B�ϋ
�F8�[�<�'�0�8�L�wڹ�p6Ck�	�Wt	i
��l��O쌸F|� ��I�E����	�~�A(�;'#@�UKLs$�ԇ'��-Ԭ�k'h��	�{����h�R��N�a�9�U��cr���_dmD�����@h~�0��=r�y1��0X�qw~9t-� �/�:�pq.�'n�F�����q劙um���w}`.������������j��Gm�	���:
��ξ&� �U�Rw.��I��5e�Y�2cD%�t�R��
�Ȣӥ9�KM���v��A5k	WB�?b.��K��(�S��	]�Y�}�p�<����P`Gn\]L!��:(�^��|�ϲ�b���U��W6V���L�������]	�NP�AK�2��.���-%�k��z�de���͎��a�G\b��'� �42ѱ��NB����P�?6z����]m��P�,(�
���n��|hP�{:E:AF�j�&�Q��,�E&��K�&��a��qz��tT;�䅣�2u�5S'���L�d`gf:��^��Iq�6>u�Y��~C��VX����:����I�WIs�%��ͯ���mN����jY^�
�
�␆���1��]$o�����C�J��Vh��~8�q�k�������ڂ�]x�b%Zie�V*ع����\�R�r�KP�9�ݸTI�`^����W�Z�}�/03���������F�v0fD/u��I;�����*YÄ�Ka#��=GBG��W� �ޏ$)��Ύ"ၠ*!�x��_�&k�9�A}�u�H ������*���k�j�1��(=�-�������xR���BS�r]! ͠�5(��j���\Հ�:6b�%�����F��X,���6UM�D���=;��� �s"�,����ǳy�kC7��1�
=�J`(�)���d혶m�EJL�ZM%��`�T-Af�%
Nd�I���&��Q�����*]��1���ϝ�HJ[v��6ڱ,�$7S�#�`�����A���y+��BX��YG�>nt���k��O�/�:h��)���kq�̎d��$U����g�#�:�]���%��\�J;B�T���\&v	��}�aŞ�c}��L�}J�d�6�ï�?T���/ ��̾�-�'��p|�-A�5�� BS�m5�=^��:A���`�������K���7Q��(�������������˺&P>S ��)&��'�؍�(�W��R��/�_RC��#���ʴ¡!ȅaMެxww�A�w)�⑕(���srZ��o����n�g��^��2�{�����ng�O��RB~õC.�g.N�/�s�L��sU��c*5��5��o���˥��t3J�\D�φҸ�l�ۂڌ��'�G�&t<�{��tj�ƕSg҉vSQ���.6u�7~��xH�?���V���*��9��	�����S���{ի�'�i�>�vsI�Z�i����Ln�n�+sB��B�ˠ�GP�FȊ�r��F�S���F"y���`�d���^�����Њda����(��l.0C\���xV���|�"�hI��[��dl� z5�)*�����]��;�#����q�/�eяܯ�R҉d�oŷ�a3BNw?c�{���΍@H�j����ݑ7~���fQY%Zǧ�ȝ�m^\�j_$3���:�T�R�r^�A8'���#��}x�?��̔J1�M��p^��T��#�l�Ii���`V/�ѯ��"�B��ꙫ�`]{gx_��^f�����u_��a�K_(�c
	C�_0{s�CƯ�J�ĕ����|/x�Ѱ9�t�b�bŷƢ�Z���N�ţ�G�$���Ys��{*����q���BEC��vp#�{h��9Y\4�T�psҶ��%���p�y�L|�EH�
�V�3�b�`�h�E�z��D���S�j�������-�~�n(�GQ�)f�T�f�8�U���Asv����د[-eMQ�"��3zݕd�d�K��K	m�W#��b<-���9vJrE�J����!+����G��� ��mQ�[w� bW��GR�6��No��b�%CVuc�Ș>���bЊ	oYɇ�?�
>L칑h~~jSv����'��$�to�0}i�`���q�<�gi8+(��l�4N�e��iV'�#��Ơ������dq[�xQ��(W&�A�IS@�ܡ���is�󏈮`ooݝ��# �#h���}�4���*�Z<����}�yEf�zw'���[� ��D_�+I���7w�N�]���vϔC�"���R1㜽)3����a;�mп��_˲��K��u~�.��smdO�I��JD�\��j�=yP�ˀ�m�n̿:7��0!)	.��q�\������X����^�<��,[�_�@�[=TR�:�[���=t3��i�^�ڐ/��
lD豉g|�:�h��$_9Nn-��ޞ�=(��n��9ؤ���c�6+t�k����:>I������UoJ�_L�@��C5�E0��a�{�f�1Eg�����y��j�s�6���A��!����z�� �)!�b�G�un�3��!��2�v_��7���=b
�иL�4�sk��]a�:�P���%�I��%�oU�kr�]���lu�_�喎�D,���/�)���Q���P���]V����2<�Ti�s_�����A�]\��q���(k���=%4�f
�/���Ѯ���z!�V��@�w@ �&�1MU�Z�:wni�P���c��7�Wr��~����*QŹo�U[E,q��>��8Ee�6�ѪDi��a"#U𮓉�۔����,�%J���+"���a\��,�\r��~�
˜� �7��<�j��z�T$)V�Kr��W~|�h.��-�'~|#�����`!�z��Q5 ����E��ڑ.��[��|�)�AR�\L?���CP�ł�}����y��ɏ7x��JS:�y�;:5К���/sV#�X������ �6ȥOn�/�dt��(���gFi&�撚�=_��i�"M���4��``5�O�Z��HYOv��MQ����L�@{��?}*ˆq�0[է�\����Hֹa�b�j.�9yQ{���d������K�`��Y詉�#b��@�����E�� *�tXP`@���	��o�^~�і}�?�)V$�c�>l�����ģ��^a�JU�ez3��BL��Ih�	žL��xц�ןx �@�J���UVPS'k[��T��L�;#&^���GM��vnBi!G��iE`1���q�����o7i~?�B]��H"~`��O�,��9VSkM�9���4������l�0R]�q>ؖ/�]k-�~���7��
KA���Ho' FB����U:�7)��!�=�����X�ؖ{΢��} �_�"�]$��ʅB�_�2E���ɯ��X�A�!��+��N��@`�u�%U̾�ff�"ȣ��R5�H�Eﾉz�I��E5V4e��a#Dc�A��y�D�;�`�[�`����af5���o�c�,W�ʙR��p��'��Dt�}��>�T��������l$y0�=m�F���f�VXE�+��'&8u��|	P�~
�D��ֲ88U��R�vȓ��F��R�a��w�R�S�!CT��w��Ur��Ga��'%�����e�	��XЃ�p�:WA	���Do�&q�5Uլ�n��n�~�T,�.Ei���Y:��ġY�N8���x��?��/��9cd�'q��s
��߽6�$���LX�Kw����>B�Z:-��q��ʺ3��^���]Pl���n*n�����s5S�w�֓�}��Z�~<��q�ǹ#4�ދ�x�EU���������$k-�s�� ��#}���.��}�7j ��k�A�����!^1�/�[�I�c$ˠ�"�&���t�ڽ�,��<��8ə}�;���U���1�����拥X/��M�w�y����Q^()@���P$�t�u:��⋽Z�J��H!r`ԁuS&�}.��U�X}�J㴏���Q�n����uƵ1\Q��� OsJy ��$�8��JU@[C�!���i��nH�Eo���jc1Ty����m�ڴ"Qar<���N|RaLmd �<OI��#�2���-��;�}>�z*�k��R�~tIkK������1K`�Y*�R�^�R��!ۍ��Y�Dm9�ڃ�+̇<a`z"�7��3'�E��CvI�8A���n-�9A�Fj1Y�y'�đ5���|C�p<��+C�Gj�&��l1��C}ywRj�����l'�v	�7�I�z����בC �Y|���s��3�\6 .]����V�"�M��٩"��j4l&95w���"%w�T�M(M����qd�Q?Zy�*�2`Iyz̶�TB������}���npE�@�U$F�2�f-���˪�nf�A]|1&,;�3�g����L����w��$|5�&Xu�+�AN�N9|�s�OY�Zx�L*㝚��a���"��\w�w�p��s��߫Q�t�;1b�-u�Xy��B�c�MVj���Z{Ӎ��y���!,xh�B�2Wn��3�x�K�]ca�Lp���J��@g����ۮ���t�"Q^���IF�mõ� �De=g����r8$��2��yZ��<2�A]R�&22��`Q\�v��;Tj?,jVAm�@��2�Rqb��+�V ^�ݸ�V�	��&
����$��JAj����Jz�^u|ܐ��A��]�������:p'� ��,�EI���G�����$�jY_��찣eQME�\CRh�y>�/U�s���Я8�&��z��SoO#�	_T��k4�����t,;�ఢ�<Q"Tȧ�"���UDͻBȧ�������rO�����@]�*�߇��\��
%g�+��eF4��j�o�~��}�IW����1� ]�K��3�]B������b�Q�*��V���@�;�x^D��N����f��2/��=�D�8�e�A �^�z�k���#��;�Dlѣ����ˊ�+��/tE��R�;��4�v2�=���lM�@��=���;���isn삱uZ�*@��H���~��ԣM� ��a�/�������<�X�j�
ty��с�vT����\U��v��Zv-�;��c'���0+��n�T���#�h��lmW|�_�[�v��uG�~�P��"F�5!�A�R�Xfq��H�_f�E��!�U�W�Q�&�4��iׂܹ?���w���S]��4u����-B��|6�_�ġ��_�; i����sX �&�q�&R(��F~	èK��}Ț51�z������ ��!{�xӡf�B�b�����g�k7r�QЉ��\�Ss�u�r��)�	�Z,�VxR�B(�R���foh��i��̏���j�sM���f��CDx�1q���bܱs����C��]WH ��Đ�X8�R��e��Y��嚩�V�rL�n���F� ���-��S�&�xw^�a\��y�֢q2�_��?���6읎�l��h����e*P��%�'��<4.�v�W���Ջ�v����P��x��^M���(>��״A�Yra϶Z�M�O�.���B��,���ގ{7Q�����*ʛ�~|�p�%��l�/���|"���I�|`��	����I���,�Ǟ6�w�!�i[u֧X,�D^;��^c$L�z��X�0�S`o\�wFY77��XUC�ɶ��,���Y��p�� p��>����!����)}h��x���5q�s(/]��h����[�8��q��J�9���	==ehU�>{�!�0�A*��h������n�]���pr[��4��~SN��r�0��yŁ����nM*�Ar^�>�e�8Ux�8�,��D�c�ݚ>��5�U��1�<aU%��0���k�T�Xohzs�jbM�8AC!��Ւdǐru��H��E��7h��c}��<4r���u� D���_;'����B��s^�@o��r�h7��I��V�0يv�ݮ;�"�����E(�����^�$��뻷�7�T�sj%S��RD�G��Y1/�P��U�Om_�yzL�m��xx�=���g0�JjFGN4���C ����F�`�ݣ�!l���
�G
$�X����c��J��`�I�P��f)P�zޜ���,:j�ң�����p��N�c�,�\�0Qv�s���>�'�hf�ﱦٸ�`��>���ڬ��T_�#�p���a�P��!��v��k����K�]��R:���xt�b�2�vrJ�����B��ğ��O�>Y�S������n���p��w�)��G��P����A��wg��+1+2���Y�ﾜYO˟�C�A�~�;>I�1��u؆O�������n6ˌ����)�&Tc8�Χ��O��W[���sp,�;�TT�ɪ2��:��8�!���:R�vFJ�R�;)l��z:v?Z"q��Nd���,S;��4mPR�_Y.� 5���"'2&#�sΤ�O�!L��
��Q}�0�v2=��"�7g���VQ;��� ��1�������<Ĵgi�C�8�A�t]W5X�l�Ǝ���%d^�����ϒθ������jU[�M�����]"'f�Х��\��G
�@'�܄'�h�[��B�L��F�P9�Î @v*{����Q�->�c��?�ϷHm-٫Od�Sg�7S��-F��uQ�+
G�*�� �/���emay���[(L�]��śp7�F;�ҍ���宠�;�����EZC_OE����?ʵ�1�>���J  ��>�Ƥ���YXb���
C�ٴ�*�jj���3��)c�|1����gB^�_�l�VCn��}�+*�3,�de��y�N� 
�/pmk�n��ᙅ,w��vo�2��(F��ts��ꘐw�n#4����9�7�B�K��@z���ݫ�~z�D]մ���~M�沈݅Y����q�S3]����U/�iv{4��M���]��&|��+T�n(ǐRom�}q�F�@/3�1ɭJ�qm�@4`�ǒ�"�1���5}���s���,P2�a�E�S����s��o;;8'�	\�o��H�9w2��#,�VK��9�	b���p�i�' ����U}��q��?��_���$PUSO�)��<KKM���*DH�x�И���;��CQ�.)č�]�2%���
:bd���w��֕��R%9�7��	�R[a�/�=�\���c����4��;��vQ B8��������!�f�1�-����
CF�;�V�*!aQ^~�"�v`�u�~��*�G?shȠ[���m��S��o�?���ʀv�?	^`�����C���7�7I�- �i�����>?a�g�2�#�ܰ��3L��_�v�N�qj`<Z$�>���Hd͗�O���Q*�-f'��M����z����χ�(�a0�z��&5����|�M�Л[��(��#���;9�ٖ�h�+_�W��Q����� ?=�y2P)���\эJ��vT�����w^>�N���1	����uwy7뱗�C��V�0��Dh� ���X���ϣ��mL�
�����\wSԤ��/�OX����\�aˇ22񁊨9�%��'��ݐR�5�W����K��Tv����#�5.Ryf�@�O�!?]������U�����ȴ��řt¥��P����nRT��ӽC]�'mChG� �9�i�:��5:���,��س�w�ؠ'�� ���N��1��_�:B��l~�Q��9��l6�@�d���
�nz�'$A�q�(;���R�`�U�u�(h���ƚ3��tT]��vwl?X�1.n�Ѯ$ǧ"]����:�4s�Y �^�;K�.VfБ!� �����m����!]>1�gDFϓ*v؈ӏ%c��X!��÷=MG.�H����d��lJ�ִ[NF�dG{�k/n��$ߖ*MEvO*{/�#��x�����}�EG��~�*2a���B�A������~�2~�T?_y#ߙߤB�n��2aJ��.o�!���i<m�`%�)
5�RK;�0�X�$6!�{����z������)n�KK�4�]R�e"M!m�g�O�I�7p~bt�v���b����#��]�:��T],һ�uUKT���9u�	t
JZ���w����(�������8fHR��}�Dњ���^�Z����w|��3� ��e&�H��ގ��
��6u���]�Jn�O��|�|P�d���LNb\�	�t��j�����Q%�<vS�� ��h��'ܳ%9*+�t�}����i�<��`騤M���t�mR��^�U4ƣ�e�8�6�f��� ,@�'$A1���X/D�o�&plQX�ѷe��hU�-��O��>���-�ai؊�Ϸ�,a:Àv*AFdLn��*1�3�DtQ�U��i?b�>L��a^kif�Mc�j�gRe&m��Qf@�p�l8�-��S�,yZ �5�0��p��P��)���	��U�������k��ݣ�{�����E������/F@jUv΃x�vq�eЖ�I� ��6ixջ�i��?�Y�F�� �n^�_�^0�k��i��V0��HB��p�����Zþ��3m�!�C]Y����{>���5��	H�#뵘�Ȏ��ɉz�Ҿ�d����ƥ0�;l��#���7�Z�AF������4�HY���� @�^/ ����f-�ڕ�S�&����m������ Ak^hgH�v�FeM���Z5���bt�cs�v|dd#��2���ǁ$ۻ�������9�[;�i��"A���I�r�uJ��2��3��w��q�Y�D��*T�p�(�4��p]TF9�Q�ͮ�b�5�iP���E5:��0u����=�R�;L&�'�S�gx}a�b����ٹNO��$��+m`g IՌLg%?n�K0I%ݿ~w$�c#2�����ĄIC�&`�H����V�1,:,G�IBDw<^��B�dDf)EqjKqt�a�K=Km�ǵu& ��t��O|�-�u�B���?_\?A���J��aܓk�X�J�������*�4m����4�'uN%���B�`�~bu5v]W��7�fW�#	;�z�Z��:s���Om1K�0j���#�/J���8,+�G�J�w�O�_G�K��Q��Y����'Lʹ�ƒ��p��]��MhϾ���=�B.����}b&\�ք��ޱ���0잕A��]Z;�)�5�4�4�!NػM�iع}�q�R�=�`�P�Z� ��N��9%~�M]���oC�ʳm�R��[�jl�E� ۠R�Y�v$���Ү�4*��g��]F9��T,B 4�rߏS��b�g��N#cF"��GZ���wiW9y�⹰x���³�8CW�^�0sC��S����2�aʯ����@RRd���F���!�bW������fF�10�����}Q���L�턱:0��#��i�8"�6�#v���R�X�p������l�0�9|.������W����`hUWi*���\�����k\8��l��(w�����mp^k�^���]}��O��J�
4V`�Ԇ�K���Mx�3��& r^e�ۼ %b,N'6l�VFo�5�˚?�
{Sel���H�U�D]4�f�4T���i�,��h��m�������­�-G���ŋg>�YL�F%��j-��2T8��t�M�8���׆,h�G�N?�Bt�O�6���1����X=���$8���k�I
B�ͽa���:P�X�û�(���I�_'/o�
�V�Z)5�e��:������C���A��e��c��H�U�`�(>�jf�#D�i��O-뵕�*Y�S�z�>(_���s9���
��BG��g�_�L�"�e��'r<_��m���{t�] I��I<�޼.~�Ƈ���r���0��g%_qH�H�	F(�Gw{��)a� 
D��5>�tN�`�E:^A���G;���>9r�E�t�/�n��[N?b���-���f�Cl�m#ܝ����H��h��Ҧ���?���h1(�9aU��Ǧ�u�����~�琽r�gT,�(��.��3��եSFZ��P~�(���7���Ϻ��+�HM g9߾���Ȣ/+�(��^�wD�9����4ĕ��nb������`^�����x޾�a�C&��{�.I�u ]~�v
ۍPvko����zlz�Ł�<-�h��E0臲���S�$�*�!�4;4s&��!j�{��~�<��\�dk��O��A�¬߹!y�8�0�!�יִ�:+/)&E�̭?u��>S�&;?���b�) #�z�U`����"�@XB�m�}�6�An��nŨB��'t�FˇEAG}j��c�s0r6ߔ�F�p)����m�v�S�U�p�)��!�}��w]��gf"�)n��Y���/[�s��)��-��=C�5`�Nl�k|h�E��r.�����9�f�6����S����f(aS�����1�_ j�u:��Q�_r��u��l��hk�S��3�������u�VH�"���G��j�r����	ee�p>�
��e]	�:��2,
�Bƅ� x��m�ۣ�Wcrp�N(���H&�m_���yj�X��(�� ���^!�zU��Z�f�7�(��5@����~�2v�b'#��=�"�|L.�/��	�7Z���Ͱ����&�F�b��`qnP	��Vb�M@Y�6�UO��?ΥE������7��,;��C-����}d����)7c�AȓB��P[���p��âPе�V��j����r����d���1A�����p�Ļ�yى�R���r-(�+A�6;��,1]>��������PB8��K��+���X���΍���zW�a��6S�+�IGp��p���)�0N9aI9+:��0HÀ�wm� ��P1��"�0�_҅�)�� �����p���H7io��U»����r�Z_�	��Tc�E���	H�@B� �9���K��������m�0q<�\���W��h����:O���+m��-��
R�\��	�::&� G2S�[�I(�6�"hޢ���/��ڍ�%�-��/��!a��ړ������mM��d��12Ydl�K[��2j���l	���GlVi�A���+�䱧z��m��kK]Z*��	� ˇ�!�&h]9�tY2���d�� ��s�Q���{�$�2�6��񏌒9��qŁ�K���CL��Q	[�q�B�A*��l�5��U�J�(q��i�Iz"6&E�*�˽����VP���Y�+"�n�J���:
����BX!烩����n����(�Ꜿ{UӜ���׮�� ��s������'�3�{u�k��3`�����մQ������/w�X��f���rw����:[�Z;�x�{ 7��n�yI8F�C/���������>_>�y|�y�}�Y���j�ke�؋`��ǵ���
F���G���̨�`j���~����%{��ݚ?��sg[~V�w��B̪!
Qb�.��y�ES��Q\J �rtۏ��mv��@��n�rL?�*�2F'�D������Wz1�T��2�m�<i-��p҃,.�@���:g%�c��j�J�⣼�q[V?��zV�cm�^a�#����f������V�R �R&u�IG�kE���/\fP��զ;�;K;�1j�(�$C+��a��y��I�H@;4l��C(��$�;���?��������|^/�,T<�5,��Y8��b߶\=���Df�㠟Rd8�hIZ��F�;���̀q�Q]���_�qS
�9j㷍R�3LW��c�����
o�%K�T���t���ݚO�֓��!Rݓ������ B�0*=���ar.h���1x��,���VUA\���t����t��bw-K�7�����P�Z�
����Y��lɲ��[avZ�ܩs�ĸ�^9�Zhf	.���sb�Έ_�V?�RIT�G�HJ/������-����t,��-A4��H`�"]%��>ݴ69(�o��NP^���p|�8�3Tv6B��;)^�/�aڀlaݷ~�������ȉU5,mL����/�6t"5
H��e1��7U�V�n�d���_̊�������'�&�,S��;��+��9��/'3���#���,���e]
�c��.�����`�_+��R��WUBk>Zd�����U�/���D�K}]�M%����?�����Vo{�w+�/qσo��h�/1you''�6)6���dl]����YZ��NU�4=�����Rg�y- =c�f} ����˷YQ�첲TI�w����}.�C��Q�My`5���W��)��������`o:!3\h)!-���]��{���$>QH :�ya|���D��N���%�0G�^W9j2HL��)����EⵗaFݏ��ò����}Aa�����H���Or�<v�c2Ε#4�����,t���U����gbE��2?jr����A{�M��jE���$3?�`)1�d�Ugr�N���[fr���ZOE�����6Mlg��wѾHZ��=f��U�I�d�,���A��E��ovd�|hHム�,�����:�o1h�*i�L7e���]+�^�S蹰�5s:���#\623����x���+�C	�H��82�C�x֍�J�r��=e9��M".�m?��*�e/
�_Z_�dB�X4_Y�l0Z�"�صG��+�!�b�gMr�ɀ�^�p�ȖB	��kї�b�w,��so����jK�́�������Ԝ�/:�O����IV��"x�f^�<^�-H�N��p��g�}�-R��(���M��E7>��h����3����9̈́;C�!\�����	ɈOec˗Gl��:�0mDaUB*(uuwA��n�Mm��ȫ"Z+�4B����i��H��R��>��Գ�*�����q��EZΛ�ޚ�����&��b �J�@�$wʶ;zv��]� ��u42y��G��3%+N��]t�Q,A�L����R����ʭKm��Y��:�O�x�01Z�94���H<��$��|�c�]4M�;�VwPv�h7�X:�g��y\Ϧ�}���.^Q�ma;�����,���cb��c���*�FU\�R�D���Xi6��x=�п��Ru_cwC���p[fѷ ��ZM�2	�!�t�rAB���|�:��J�ʘ�xX��{0�bZ�����v���-�>����D�Eg%��.��6��z��#H�T��>��*��QS�����>��4wGseA���"�:Z��Xa�lΧG7��^�KQ���Ǯź��U�K��o�p!����Ȗ'��E$Ċ�	�,�6�g��<~��[x�)��%�t�o��Q�'�ǃ��>�xeu�f���&�`g�B��J�9U�۶�عx���U�������ũ�����F���+~�o��"q��.��JA�x�ځN�HKv�3��P.�$/r W�f��4e�}�7����^�sI�#���X*�������UW��HMp���";��߳{#��	ѕ,/x��"_Y�N�s���ƶ3�Q�\Y&�{�2TN������+#ӫ�	��8Le��!��I���mbx�|��)JN�Wi��L!%���ڷ�"i���z���8� �O(,��3�P�;��8+�^\�?�S@+&6��g�qfl��P߱������v?dq�5FjaNNPG���Q���n���Ҡ�Pԉ��v����L�mu���\�:y|�w�*j1���%��^�;��"���6˘?�nbv�X�J��>���m�TVH�E;
�̓�mW�K��z�~L����
5��񱃑���~zwG������W��OQ;���@��X
�Y��-��Q4G���gi��y�����nqĜ˦�>�h �r��T�����埮�F��ш^�Y-�=��U�a�P��!Kn0�w����F�D�۟�N����V��Y����D�v��E�B?�u��Xÿw}Pl�*OM4�B�v(�X=p��'�>	It����֡4Q�Ny>�@
V�T��2�؆<��e
Ѷ��S��48�t3#�3I5�z<� � 5�:��5���	����`_��x)���`y֨�G@=�dcin�c�V���v���ˤ���Go��X;�B�0��%�����0ܷ���
zve��NN��蹃�~������;�a���hRq
�.\����~bT^ d�o[fT���g���ꯩ�x_��|Zo0���d����'��B��̸Cwk�0��`�ӌNmd�ْ���$e~���5݇��QG�Ӭ�P�I|9��=����I�+N�Z�����[�����q�f�+Pq�g�>�s6t�U�O�^P	r.ى����������h���E��`���n���iͮC2F�\x���p��m��,>����M&���Y)������r)�?Y�I�'��B�dW26�Q�:�����!{���-�.�ǒ��6��Zv��(3!����̆M-aW���L.�_͝����|�R��@�g��*f��`�9��Z`$q�bբC�H�LL��L��qKB�4��iiSfow�O�m�ʡɉ^�����Gs���ɉ5���f��%���ι�E��l`��1��7�<r	-ۂ�9�]��|�����^�]�D+|�	A�l	L������4'�Mg�O%��,�qj(ay��BS��땺�;�!�.�a��Uv�����=��7ŏ3bZH5A�dǛ�^�ࡲ	!�zu��h�}:8	.Ɵn=��r!#��c=뙤X *�-�D��y�*Kc�=����Zʮ l�Gk%��7R�K�5o���v/��t�__�2�A>��(jsX$3
�(�ۣ�N�Ð�	�|Y6@!�7Sܻ:c^m��I�v�A9�jE�0�;�� 6��!���N/�n~��6�	��O	:x���J��D8�Sb8�������%L[�PE�����<�G�'cAf�^? �12�uiw48���
�[˸��Qb�\O�{W�����SVQaϝ�����ߋU�<}�[[ԉ4輝Lx�]`�x:ܾ*Ua����>TR�Ȕ��j`T�ÅS�4��Yv։(��-˳!5ؼฟ܌�4�y�{i���l��?LU�� ���s�>V\#���Z)��0:v�P��g��.��jy�o��%&#Ƣ)K����3)�Z<��)���*��K:�ě+�ҋ�/J͂�R~xa^Ń���7�7��ҿǅ���,�$~��U�����J錋Q�_�)�"K��y,˻cv"œ6@Ç�_f�F�w��ckcS꯫h���&/�̱"�|���|����K߿��s��D5En8��<|c�p,﹖M���@���l;�ו�NS��{� ڑ�(�d��@k�M�S^��!��E���4mx�4�����YA=[mc�ς�wPZ�=��w0j��"����n�"�0ι��� �:��y1����⯧]��m.���!��zB���Y3�W
�/W�z�Ʒ��q�@k��w*.�Ȏ�|k�Z�W�T��?�e�˓Nژ��ե)
�5���d��XN]�i�� �,���|:�%Z:u��~i�k�wN(	��}w������o���g�ȹ��e��_�2ܘ�M5gǋv�w?O��r,���G��\�շ��&�!��e`�O?uk�"�9I�z�l��+�F��F�V��nl���,>�����RlP��*��~�)d���D<5k���9�m����nk�O�N�%�@����_�P0�Ӯ��;S���[�R���_�rG�����ه`?�6�*4�r�e����s��uT��@�ص�.�.6Ơu!R���Mq��%�2�5��>)`�3�}�51��'���ӌ�F]㎫������"��Ŝ�}Q���ΰ���������^�h���.�U�Z����<)9��`ba?%�h�g�!G�y{�~��$�m	�G�������;1�\�~��P�G(���k�^*���D��0���u:���B9�i���ME�5��2�\���s1����-�����;�+���U�$[E���ZLBI��}?Y��0J�^!��k��¶�CiV&�^te Qx�&�}�����VAKc{�jІK�X~n[8�3;�-uJ��1�Qxw���L��a��bHZ�a�>�~�`���E�Uy�&�2�|��a5-@''2~*8A[�D��J�FX~[�D��$G���,<P�Q����K<~Tc���5�b�`�:��퇴۠�43�݊�b+R�~3�p������]�g�a��f�t���G�qV�ag�L�����8����l�&Tx��#P�H�Pc�qb����Al�����>OsX#���P�7 A�1�y�F�^q�q2=?QK:"(���Ig�}��G=D+fm��0yy_⥋����t��`B
�3��y)�o��
Zn���ٱ	H  �E�z낉E�¼(m��iV���	�b�y�W!�%2O˪����6K����2�Z�e�xa)�#&%�>+B��]�����r����1mD�7% �jb�7h����%���ȔWՒ){	�| ����V���e����@���~3S�>�N0c.�nj�'�������h�E�k0��*+��
t��� \�Ka�g��jS��ԏ����*��|bu����_�H_������j������O�I(�hj�:ǜ'H��|�d<8����w�x�<G��o�Q���VO7��s��ddmv.������-���f���s����p׾����G���F�9���
��lj�H�4i�#����������u*k!w:�-喱�[�(�*������ȶ6�_�o�SLJE��6k��\��^�.�_h�j����h�������8.m.�A-$ްҐ�m\(2ʓ��̓���(� ����i}����x;����s���z)^�qZ��1m���Yݧ�h�$�0��t�&x6S�.2kY�	���@��G���=gw��{���`��;�l*e��A�/�����������O�[c��J@��$X�nU&Ujt��Z�(���^b�Y?"�#�njk�
"6��]C��Iw���h�^�^_�eCK��\��i0̠�h�hA�^��A�N����{$����Rj���F��Z����hPh�9�z��U��I�����O ����u���ă�WՇ���*Q� �Ev�1J��|:__|��X��)�1�|��x��6��:��BP���惓��&)N����3h���k~�9s�`_^������L��.�E���
FL�Qr�Q���Lԥ$)w�/f;_�?eru��3F��K���^m�H$��׀�!�o_�6���X���<���}X�4x����1�����a���.) �,�ru^˹�K+�Tl��a�#Ί?���Z��A�k��!��m&�Hd�Ӆ�~ZB�Mƙ��7/I7���6X����V�.V���_�-�.�����g�x�\�I��/�"U��n����s����4�6~ߤ�9�������������4Y1�!��2泉�p����B�	�ejQ���N%��?��ga�2��^9qO$�>$��<��Ѐr�{�ȵ�խ&���w�+�mu�<ir21�-k ��(`�UH����q�JP����a9-�~榲�di��	e�Gl���'�$��L���
/��a���dSfͷ�oZ��x$	{�|&w�7���tc�F�.:���n�֟�JPg�܈�;�Nd��Q�%�g7�q[�d4�(w��ࡗ��W�@΁���q7�� �/	0e�/�ɻ��}M!~�a�ŷu�ʶ�R,��OȀ���bb��0c�O�ȿ����4�˗d�W`�L;���J�$;�Eb/�Ԟ�\��B/��}d����WSE���y�<G�9�O�TB��*)�t�R��.�WdG��{�(�f�A�Jc�qD�k�aU7���]=�@�z�qE,�h!��Bl蒩*��[R��V%2��
����<A���p5}rAĕ=Ya��"((�iS.�m�:r�\˶��tW����I�l�N�sÃ�}��8!�kO��;3mԈd4X�ZԔ�+��e��f?5V<��V`^ZL@���z;?㢊�~+(?�x��}����"�~,�4�F��QfAT��Ad���T��"[r�:Yҕi��G*�n�����W�w�D��r�fV�s.l|8j�aʪ��cyyG6�R���2nNsrŪ��@lؙ�����)Jm��Yݴ?�C֎��Ɔ���C|\<�ݹ�Hp�J��^���)S@.T�R$�X/O�}Q���17P;���`�ޭ%?������h��"R}p UU �<#���'#�_����hN��������-P���A�Oq�9��,ʐ#%�:e�G�஍��,�P��v+.xqahie%:��7`������1AO��_UBI�b�m�2�����	�;�4��� �w����,�B�D&�Si�b~�3K�d�2���߸F��g��C3�4R�Ҡ덜���D��|N�-�IE�����E~��,��� %OP���&�v�{-�� y�̀��5���>#/S�7r��ʗT��mݟT����>�����'�8� � iz�h��%��A��^y�!1Y6e#A^��JpT���ܶ[�A�2����E�H.|����d��� b�*�L�����-���"i\X��It2Ξ�B��|ӳu(�-��x�S6"�L�zX�8h���Z%$�Ő�i��ObnM	�d(��P��n�  ���P�-��dy.�P�ϕx>�f@CTumǸ�{ �J�a��[o���������~p8إ���V�-:��ב��Q��Y�Vˎ����]����WaT�3Q�!�DY���T6�*�,Y>^ع�O��r�Zz�
N�-7z+&�D�R=��u��q����k�>��ȜC���j6s7�S�A��В%�PU'�,:�m7���MM-�k饷?|��#� JY��/�`��7�h��w�6E��Yt���t�'������(�m�S����	H�\��XS����W=K�����v��1;P��6��̽��{�w^Ǣ���͓,�2 ����4�������0/.N����³�砓�r��/��,��D/��@Û�Y�Z'��ʅ6���G\�2�s�sj5<&_�7��~;��"ث��t=��Q�g�4�w�oX�+��:0?�Z}s�5P0s��D�AQ�r��궲�XF��&�B����-}�*:5[�`�����3V�T��=ML�ه\Fn
"������'AF��D4���E)��t�q��"W{. �&���r1c��y�.�)��B����j��'������b�sf�r8��u%>���t~צ��	ѐv@��>�E�xs�� ��+&0F���i�M霮��e�Tf�sbЛ��ڨ�z��d�ߤ:@^�K���\��J^/�l��N���3����o�M��y�����}R���s&M�L��H�9x���d�UeD����V�SH�=���#j�cI_A䵢�ZSN fߚ�N&�\�;�AT:XW5���D���AQ!g�իN/��/������ǱG����n�+�����I�A�U��l+�ͮp-�!��N�׽rs�}A��<�n�k䕑3�Q�碟�`5Op6����Ŕ}�f����o�++���\S��9Ʃ�I��P3@�\Q(�K\������|�@B���KR���!G`�ܖD�|?T?�w t��ѾA����U�⢝9Q�c�r�=(zk|3�����n