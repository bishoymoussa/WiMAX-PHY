-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
wp03Wnr9QQObYmNIe89wxenBPJOAP3KLxodPeYEZb5f5K7wT79mKFXDQXgiLZSKMHfk/LTcy+/8K
2foo2nmQBZ4T6Nb6SVYfQvfQ7viwXFuxomJASpQJyBQHPWHAICEfMHAaRqS79jYnlIFRIYd1o/Tr
U7Xu/ViM+nquSVcL6hnW0yEJO8WFzi94vkfz3uY1H//6DEoJD/Waa+eDLuAdO0ep51KLLZQj7jJx
0n0t4g6tT2N3yQQXcHU6rRZZ65QHT2ndNGRP5K0yMEbUNSainSCI2DrqUsc3fuZgUvMBS02otwDA
Q+nutAMSSNQ3OQXeS8MsDTIRfkWhL12KK6yHrw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 3008)
`protect data_block
SzmLaBn774AllJRj1/GOk17edd0F8MZziHDPqSsw2LfbFP4ZPFABbsxyyYcmB5cVj4FyXdIidSIn
BGkOwStCaO21kcIPapquopnsCXY2MnhryE2+3oeHg6jQYd8hWe5J3niSJmfzxnKRhp1Pwdae483W
3vCllc035SXgZC3eRHNbeSKBHrI+Y68ciFtzFZ6+tEgf4G0C+ZkE+bJ3/LwcCVct5L1XSEvzfB8C
YLj+gskvXZevmJakhuGPt9yN2tlqGg87iPdd7fKj0yz/UUCjvpGzTKUdwdExiS81dfvwHudhv8eT
EYrcuI3f4NVUJ9QEwud80Kgv/u2JClqK+5xWFGNmIUroUkMY5R0G+xptrUPFQgdJSsR1PcHJBGj+
MbVIjwE18427KmR2RbL9UWkacvom/gvlTdL02UQsH7JEJphi3fAGozrUdsc+UK9/dDHHaRwvj6mr
FnYs90DaqeU3i4dSTEKeRJjRRhlu6gcjgmHistXOzTQMN1sKgAA1yhli/3NvbO56sMTphJYzMKAL
NMEB84jQABgAMXERBaDo+JNHYzOzjPTGJN7X+V5mHlymJQ7qAcO4368e5DGoQPOSj871x82cFKR/
SWA22yI1UmeYmpkphJbGBuNz7MW3mwuche7l6fu1cbf+RGTAO0v+HVJ6S151Kh7C3BgzyqS4UBAL
mgEx3+jXFOHDq6v98RD4xazE7t1MatP9Y7/UPqXmAgjb8f8bHmaEZfvaAFZxHHH9WhTFsi62fbTk
Hv0IOcmPHNbh6VcGei0JxoHdMy1YGvROJAsJ5ttT/euqama4eubLIjg14zDfRqYFDxFsWIw8Oi7D
27QaFrVEooyMp7bbO94Yt2eTnXc103C/IHn6XJC8iI/dNr2olqkUonS0JErViGP7tnjohiEKaMpd
uCBisFztY3VTGoBHCKLwWDGDsIhbtDLzzlI7427riR88jM0xycqC9cLnOzKAC1ImUcie5hgRSPoY
NE4EkFwRKeaXDjLcFLW4xKjXESAQn+6L4UpUJuZjxe5A+hDEC0Rn26MaCX+bjL/TqeKXX+sAD3I8
ir8KyGKoTlrRE3X0Qkiq3AfpxcPTZAkUy0SmY0XbUX6nL7bci0UtKokjfFYGSGpS7Mn24s2oEjrA
9TlWtMwDHU/w2vrJn+UNkB0LJ7+rpS789nz1ho7HRFxxITyNXZm1RTqzLicO5qLJaatKqt14X1d7
2800F4367zzk94dXPdNZdkMSxyBx6KPXwfb3gRKk0GiKIcLfwbYbMbe/OlFEtnTT9Z777CoJurFa
rwsTfURscX8QO+RTkRcs0jq+4NJSRnybQlJVgYfqCi2j5Qh7MpPDCEmTNoWwgSDLturCLXkD4ym9
skl2L+iMJaffCS4EfNCzTFUu1AlCRzdNIp5oNAW5VgjtTnkYUU2xlEzTQ/JGQLmjl/BEbVfnjEhR
GfJMvenW+Jcatf1VMGxeVp/evyEpz4HP+HqKwbTLAZcwKLFtUN5IUXK3smXQLOTHPK1ksHB0ebBb
AusPjRtuR+BiW3cX8NUqH21I8Fdho0GSpTZ6o1HtoM8ZdSb/1bmQ+hGT+MyhoifJSXPBa0MEW5pz
BpEKPAJyTrRtW/YDmTRTwD3voJarWIt/RMylPbqt3HoaaH5nsAOkyVl0+WVL7zgBdk//B5gnOHcc
l4zevT2MvikkqqaHORsQkp9TeaHnHUJnNLz3LOSt3dhwGeY1bb8DGP6GeTQDdebCFus3EQxdCml4
Shh9crcldhJTjecyzoYDvEAafA+WPbBPNXzTPprU44ojB0u11KKpIKhQYyFjcQxavEUfnxsn4haz
IQ/u78dIEYHpCxLubc7FrPI08A34zxEFu1Mq7pTzjt7jBWG0lNiYGJwRBqXRUh9dZxew1wNn2b6Y
C/KAm9A+MYbZ+H0X3/tWO6NgnDUPo84QpqCjIktPjNd2yCX2PDMdbyl7iRHcBShC/YcmrcejRIn7
BL+XRUaAJc06ZIWexdkc4eHoQOngDf56JRYgHXR8Zu6g1O+LIcjI/h46eGuLLqdznOoieJBAeWWV
fo0hfbBxCq/8wQ178ys4nIJWoAuBgTosfolZJDBHxcZ6+JLL21Y42I+EuZk3KfEcFwco9luXPlKu
o4DVRPzcNgwtsoS9K10Nha+KJXnXbcVxpn1Mb7Nrx6tUic4S9NAXgGdq+n9o4SPxTMPCiWy5LVBf
7emaBmlJRAho8wHZRoinl1qzesGLMbi1wURziFWgzWJhlLP5dZosZL4KaKDoX4NTMEKDauq440XX
+dmgbzH57FCzwNXVnO0Jvlpy0SLxa9VSCPQkHdtmjg3GU2vHHrh5Bolt0D6d1b3xns+2aTYvfmbw
n21ui4K9PH+tAD6ZRXSSlPXYlC4SylP4j5zj7R0COhFx+KgGHSVnzNegdSMqC2vYV4QydJNG5bJX
yplOZR0wNCb3YF3Y/rPeXl4/hD8oM737XbH/FMaOT0csCRr+klIF6tZE0NooI4/PhNbC0bTcTGvh
Ab8m49B9A30uwUb0rbR/kO49M7pX7sEBRp6Jxuv392DeHIdxKBnOOchwCNoP57xkINsJFrv2+15W
ZNetX/PIGeMA1c+29uX6INGAVdzTGd0/U13hakJPMlW6NfQdWyEvOwI6GyyP1gpWr6x4aVp5AGCX
FHSRDkLw+lJlJhC9/SaqDlvKk7OkgCAmNMxDY0UQq/fLGfXLfdm2X8ZIXyBtokRNhyXMgbWvH4Lb
z5E003oHrYfo/Cq3cBPdJ09I4l/oMz/u1bTvjiCLAsK/EFdBSzGPlJkgS38rVWMdQeS/jt57TB7c
lkTdPufWsrD36CsomZlVajQgQBBCiUKGILMYTfo3C2a8davKluLVm7tQG6ZQbNFrG9zOhb6no2oH
ORtHvro6he3J0z8F1ttTQxGEmmBfWxFQ2bnx1AuvvTg9gF17Q9NqT6VtPcW02VYIv9PCgt7jb+xB
rrCUJ1LIHvMI7WWlLcxPyjEKtnZAh16mxLx5BcZG3RWWCOFswH64kbxOrBYbobaMPDnweRCDhy/N
fE7yWvCNRymwb6MwwLPopXwMcKoysjHTiNc1zeZHApvOfQ7gAfLYa6PlxZSvEme3Hp+d/cRcBAzn
ryvVCBRSnyq96Omf7XA1J8rMcIXhQ4xY2o0zj5bcxWnnKegJUql7Q1sq+dPmxibjJd+AX8lHEY02
S9BjISFQS+YfodiuM5n6+iC9rXClRNKZI7q3e1wWiNVd+jz0gDr8XyMZ0BtPykz9k07IRcx6QX9j
AM2kKdSJcXT3gtAkl9/ryEP121qOORHaoYCPofr5hO0kXI8625RDOWLywVoE6yz0RMm3V2QBKWGD
k15kNVdR1qTaAD0T/iDyyHktlZPX8u+7yTLtOX6drec7qngovNQU6Ftnnt10WdY5tRTnVjYffxIX
huNwHYG+p6Busym7oUFxLK85Hshinp+mLRWrYoHUBxTYo5gkqdgBpm+bFjzfm1jREUp0mcVnjydL
JUx1X9SgJhJSgznV2ltaZHwbOrXTouvsmkS7+iCN7p5te/HKlwS7nDupqq5ifJZJTrlezdyRCloJ
EYUvr4GH/UJs9AJKff/ygxckppR07BfioZS08tHeg2HFS1KsS3qTsguOM7atYu4C/isF3iXyRYZR
8vyxwCuX2DvSJjrD0WQQ6Vw1OIoIaEnUNEl46tgEzLIYsfGiqvoSwIBZOcSqsXjt0Z5NKXIyXgKM
RDLS5DDNsiuE3n8WHj1SUF8dLtEjjYTtHaNg6flOJIgFY691uD+FJc6fQf/DFrwhavKe3nOIweyB
v7tTfhOJWF7/CUDs3rn4bsQ7yfc5AOGw7UznokBbzawc/EVjiSWxsnPh8d58C8jS9aiCWPNHYCRd
DwX/oJ4LVtCEmQnPNLTcZF+StWPYhQ/tUlpW2xJt/Z4th1LcsSk2l/hzAxorZRdCzWk/Ra1tPmt/
44rnujvjgDm+AbdqrV2LEiY5zveNyn8pFQ39Dzvg4LJuovxvxoM2sfE1NHY=
`protect end_protected
