-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Wa8nHQp07mS8iK0XDY2SWufuLofW5azpqZ3wqqvMSy1lCzwyILKLFA7BEbJn5PQam7YHxoZJpezG
HWuQC3X75wRdq6a0BhBMSXIuO8zOe2hJQpMUb9A5rR6IKjtlT4ZDbpT8HOt9aMKN8aa94V9DWuQ1
D+NLq82r+LyocoIqumBB1F9d+Gk7eAWB7tjg+UjjVYL2bMSQMh6th8TmzkzRs0H6m3ZKvDNMSa2J
9m9E0dfM8RSYjvXMvaa/pDlzpr6h3oi252dPDI2jhXmJJRyzQXD3a/p9Gw0MWMD+NNjm1K9yJPbD
13UiOcj/vd3q6b2Nf0R27DX4XB6XVbI3XtMTGA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 30288)
`protect data_block
9tF00+zamNIFpkHWHB2i72kmeovKc0Ezb9ImuMrRIByrnOluu1LmjxkmNKtmYzKwjxKGNVsZJaqH
hjEPnjJvvbdxdeQyeKJp/gb1Iv/IK867kuwrZmGoBXodnK+KWZ+qlaPrUXmGsi15ODqTZvzDAv1V
hUpVrX4P4rjAvcoZac3jf2mJjYMQeG9tQeyoLfj+mFaG6o0D6THQ3Dersw523RWyS3o/CAj+UYNC
qPAQrC7VkY3rg1M3UbIbRb04JHgKXjvH8xw6dghaMBYANuHl3uORijW6n0BFccjBwT1FyQBBp7Xl
wcDoYr7/Ip3K5AkFFXRKYTEzguzeqXbzvJuG0Wba00KKVt5DXKrECHAwDSKS/lYbS5KFsyC5iv4Q
+b8cNju4IRbN37fnInpIfdkWU3zboGw0Ex+trVhEPVKxjPOJqmDHQd6OuIS8lDxCKFoiQUDadY9F
jH8Y6Xk+XiutS8eRm2YtTFhGBoWjGHQi5lqKNPG2e4VeJlHWzoNS693j3gHLlHZFoQd1YL1AqTTE
SCJvB5DJLFpnbH3Yjb5PZ67N+76/Ph1Ao1pcD1l/r2W1pZb7xcBgTtABEvp6vQcNzdFncKNCgHTB
kGUPutB/+f9bswNe63DygtlV0H/bET821OKAm+9x7R+Sgdr5C/HJMIr6frPacPu4iLFhpLAjQKYK
77H9fUftabDSs6MfGWgfWbUtODYqxPHfsI/NoHd7DMQOhhFTed9nzryZfzusAxWxmK3fEdnl0T07
RAfM7I1h5nw4sW52zGtVgULxC5NW/AHqtY91irSYmNP18z+OWGI2+88NJ23roZajXL0G3UWQ1C6V
fiim1kJff1a1niKejP7itqJ+P+dMEFSo7YLZUB+/OcvqjAdfOuXzz+kgkp5MG6KuRfQpSiIqT1Gy
+PxwL0Cag7ka/8Ac8Pu5ssYsLE41yxcP6Sh5kRGZr9JEq+EbuceC2UJcBHSELdwUGk8xsG2HnKqC
PiiHvuT0roKdxfEG0bLLrOdfQcG8UV5Cdd3DsxMpwCVR3qSpIbZToI0q1LKkZ/VhSg3oItoW7f/p
59EFMaDHKdpl0BSIF2MNXyF9nmaMEEfsng/kBIcFrI/dG+CUP9eBoagAj/l9RAkgoneOncoeG6Kh
O26WHyR05CDGJ7+xP/e+25WoORo1o+TyJIRSMADGJe0sbwZT8Tcxo46PuJJesjCZ55kG9c1CLvcK
ims6Ty8tnU6hgjDaRtqU/pqT+DV/eBjm3Q6y+709R1rUDkQZIN7QfJGBVUJOE14S4KQR+i/lXKUf
GHhY97HzVldboXBo0YlUDC1SX6xQKeoW0hUDq/NYQWoIccUaGTy+hX9V/3xmicOq21V482uCsgaw
QfankPPYy0NgEhJekcX4ziM+P31LfwKHMwMxWEQrFrPirgBZt62AqzsE8bPBXSsz/xkajKcbbXQu
wUnAdCaOZxhU+gfymWow15oRPaCyTZ03G4uYGHli3UXvp77rd9DdvE8gs4eRYs1hnatUmSYgN3Pe
QVUU/n738p3AqNvnQNcZKMv1nouzJ3UN5P3NjjD910SJl0cxD1G8OFqvvlvUGLBu4NdCSWhURB1K
9Nkb/EV0iuxxrMvylKBpMJaq2k/4ZacnWCQo3yh2p7qHPPMye0l5J5qMA7BIcliQE2d1bHpFdLBZ
xLo3+awVDzgoYp10Ma5tmLcdbyHGmnNILWEeWMx2T8YUQmfNIXYc0wWuboJkzh/0RpLpg4iYLW0q
ZFNqikoC6Pgq4Arf3eqQcUHaFL3RQURAXViWYxcoFimh6ZlHe/KnnSkekc2cLb3HEngN9jRe7ULt
jwCG17aXc5vsYc59TonjrM11EvqB6g60w0OKJAYTJIw3FlfVO/v34rHtnVA9vCMk3D5VuOzw3nOE
Q6a1kUNN4jEdnwn1dGofdzVI4789A8GgRwLfPY6YRnnlFcp6qvopNRuct4c+5PWym6XwINmyFDVY
VJBEgGhVNQmWFcJqoORSiX4S46QCzwe6uXgKtTYlEXnwEqMkXBa+9tObpUYJ0fz6pnWqJ/yvVtsC
MUW9Z5W/QTsRJtuT9Zb3To+nM6rHSqsBoRcMCaYdnzzo/DYEMXep2za2oL1IV4NYRvwL9viK1bf3
lXYgdedlpmrF2XKf5jd9uMGgFL8c3Pkc2L7hoixMGgb3BnNH0CmtUVdF3a/5IYiSrY6SzuwF+/u+
7Ffbn+b1R/RFOG44aYipBgW93HZuASvSjbQk1CdMIMUuN3SqF+0Q7ZhaKPo9NkZwy93GxCcF2xtV
Yd5Uq3kZTBUOV8ZPeJJWdeOZlTHOh/mAovHGkimySl2KKp9mzQsscz6Qu+EEpi5YXOSxE6xibwOF
xbQ9NyZwdQ4Mq3YpmFnG81z/Q2Dx2or2M+MXwACeikBhvJ5YBBmunkZYXnlNnXoZQdEwyOLPhuHh
krzvlkRP+nNlvdriiqzKZd8Yu6e75+IQ3biLwV+z+JSyS5hNs1uk0Me3y5HQIwK38KMmJO6emO8L
JUXzlZcxN/H6dQc7934Tvg7WJPiJh6/XG3z0H0Af7iliBvqOjfPBSdfuNiQrKO6OInDIrzASqCAO
UK8Ws/UxNXhvyBDuggafFtetgckcAh3JfG+ZywMmy82woWud981dxZS68U1LBG+4c2z6u0uVPPdb
c+NZxMiR2/C8K9sFF8FbtCyy/F1s6AmaD0tE5rDP42xvirlIBvCiMxkEhYdhSTXvK/1kOaJKhgdp
9dQOYMbb6pvliM/hHsIBX3rLgj+pVAWAGXqUfYf4M8tnyMkRFJrgnlLvJ5lhKjKjcNcGjxMF905M
P3teejiVRK6/b0XEw0Ixb5IH8l6F6p7pVUJXXOUUdTG/yYmj7E9wmxd80hbHP9CQjPt3ogL+Hpju
Zuo8B/EypLAW6JNgwt7NDr/M2/dW/6fZO8gbGbMANdvezUDsE5pbzb+hrz8WWAAbqyHZ7ulLgH29
3zpTQWMMILdWBmZntPZTEfSgoS3R2eBfyXMJdfq4bVOD/BrIlTvGjaGDm0q6dsvNLnZtHZITeRQ6
BYNMPJxp3ls4asTPHdWPxJls0SWprf6Y+c92JKDyLaH0yTUYRi8kvFIw36UzrwW0T1Tj9TlyCE1h
7FvaN8hNuB9jMY2E+UiAgK3GP+ADm/zVKQ/Lt192rHF45yoKJ6PjEgtsBtg4UZfjv741B2c/Cp2E
x9agljga3Zz+iHWulpWXE2QuIj/AWlpIyUNEAdb5wMfZHkyZXBC/VlHC4v+Wl7LXIxUYnO/0PH8e
deZRAR1eBx5o5TpYiDI4KPfBIdGhv4c+9ukPANgdxVO4sBb4tVFYw0Fp8CDwV0eJ3j1gKvmvaoZm
wrqBUXgu+SSh0uuc8SN65BUwOhl8Dwnb8JIS6GRhcjrnjltmINW9c8Gf2VJCW2X4IW4Muuvg3A0v
bfFSTxa9f3SwaWCuRhUm7eYBhbduGfT4rseXOuCXQ0+UDaWQ9FosXNwf1hG2r90u73p6A+Z7u50J
xKeOfs+OttzHlRKximBOK6HD+N9h4+SV7lwOqwOf0cZkTcg5iShj3bZIx78PVhz4cJCm/Ux+VdzN
Pgf/eG0yU4vqCW4wfZb6YzkwgAYMvm/3M+DtXxyOmOX8XKNfs75a5LkD0OtlYDKp/qYmnsn+3Vy+
K40sbGiTYHoNNmIr/EX+Hl24Z+jgRrH07XdF1Nt65WTIoYrSDcCN07wx08fmBDGcbacraXlTxazK
3cIO/mcKTIGxDqewYZc5otRXxO4NzTjLSpRsS5E6i9opa9Cr7GhXd0oMyyQGDHuKFwR9Nv6SydL2
9GzlTfyoWT6/ukdvCuHmMLJcmL5NwV9AhdxNCnjaStwxCzAVZOgPlqWDdvZSTNFtqT7HZEA2wYZB
w2hmGpU+cVU1pLyFr+zUDxJPvjyoZyFT/joHWiXE+k3LK0f37MQA+mjj4mrzGoAApCrKXAD0pz2U
BZEtCHETNfa/2zc6rB/6ea2VKu90IPW6kaur9KTgbncl9gd82XoLLqD2bRlyWfqN0/A+UodnZCxy
+21mOEJKtpTT0pDgnYHinjnbu3NmxcEw27QvyZtS+0k1CrE3LFqMs5fAGuCcdUClB/xqmiA9gnzN
H43vKgphehmglk7lVLxL2+4Gw0JtAFRxlUu9xiYdRGM6gu5cfN1v1qd6VIdeQCQ20Hon5d6t2adX
d22QJgFNTjtPS4hXOCBsF7lNZqL6ugnvUPh4ZFo21vg0lwl/e/SOhjK2EFBGXsFxfnYFlWc77uy8
V2RHqlLcF73AlZ119gzPv8sTRYdbi5GXrCLxbHzjwRnsYVHUwYi7Be/jwEjCBgb1VSFWqVd6Rn53
YROlq8/8prehcXR+4t3GJ0IXFKdHcuPKlfBJbqQn71z0ceGQYNstZB9tdDWBe27TTUXDuLs5O2iA
pcX9G5hN6Wg9qngbOZtSWJyWx0BX2k5x6Iall39Lvval5shZKm5o3C95jd060KNWri9uFWqWWvHN
JXfsRxxOcLJ+GjiqO0XzxMhHnrtUvCCJCXc2xoqRotv/EF8COd1NX7F09h4oSzOe9gpqlObCQBfK
NM9cmtVH6MccpFh30CaYJAH6nN68Bf8OK/tf6A7KopqHuZj7DGc5dYl0//vw/0zMaZEDwpnqItAw
i2biNKWISIMPQby2xhZpNNSwRQ55i2z3TWgZR55a8BXQYv/5ael+rc9HN6duXCbuMLwX2TiWV0TH
jmYAo5HcFFOTR6IStRyMYX+CQ6RQskNtJjOx+OIG5vMmQ5DBYpXY6tUaTA038K9gwQlsxxtY9lb6
ccd/2xZpC9fu+mCB85ZIdXRs2EU3RnFuKvBLreVCemP2W05hB4OaVE2PovokR25PNDQ8HEpNbBT2
JYJcmPE2+CZe5CzmDCwkVZjClrUq99RwwNUdeIUqbXK9tBE7yVelQysh7EiyIO4qTErTm6lUyyRJ
OcZqVznppkwttCeppaU23x2dtBWBOPAET3rcHhNLGGHdTwDLJpL8RxrHn/M+lZd4MTUHpr4FlVxi
QPwb0bA2oBKR8AyVenp49MIlg+r1ukzUteU8F/hTnrrGrxSgrwmdcxqvGTgVH28ktzT14jiKjioq
n4utI5vuyXxuaaRSpJXlgKbXrfFzusGMvU1wzB90DnGr9Rfm1xqZStV1LSFiMe7pD7H+Pr6xSyR8
KPbMGih1cleDvgCw2LBD4AvChyrjTXv2DmVZIBUXm5RExvLji2RJ6wVcWcGQ5EZY09ROKz1wOY8L
V30cXWfw+zMskOKZROwj5+LIUEWelcPd9W699BOTSTRI4WnXYEFDIIWTUun+vYJ3rYNWlfl2BR4E
nmFTKnJi678cQfvstbIsDklOrTFMOlP6G3I23EWGG2neXNBRc+cJMhuaGUJ89mjnBy8r9J6ABjnP
5s4/Cz5U3OqZa2eliT6bss/ZZaO7fzhHiifTuKUEPTLCTMOl0T6d2sYvrlBu85gsKtGCUpaodo0U
X5YdwxQovmL10VBN93ivZHA+K7kdhS3594gHy8QJHYxa2NSL05d4RES6YetSRWHwv7RfWZMFJ51z
7OazfxyO9wKe8oQ9Nji2j+iSWXoSrF+Krb9alGWqoWKd0aVxI6YkfQDfHDiYoYSBPdiPO+JTSZDB
Wem8jBqxXZu2sbv+K8TJ5HEpwBDan/ekvXSVe2VrzCGaDelw0X9Dm2qqn8xCuPfJiDejwiETZUH+
Yl+feCB8zQlRq8QqxtHh6K95t/Plg+ANPOG56FTF3aQgqUtLEklTn3z06lgQ5sT0/ECT5RUlsDmy
HFifcVk0gW+YxgXmWKS/mHz4bWrd1mmXhrY+sEKIi0QaXWIJh+A3sxj5cNP6GaDIvdrjLMH7aSzM
4Ki0BIVPiBD9k3buLNGc1qEWUwxC8Ar8kd786WcHW1OtLsn2YkygxBixF9BwN28ZzPR6d7cMy9NB
K+8bmmGFdy2WOr70rFhMcrEaKZvRLDymhUcAqBKhffUsKYD8erDsUfCDaXXH1OiXWFy/+it09TyJ
uCZdW/gZBecbsWC0EFGCaM2FF8Vbj1b1IrMGQCCtguUc7pdeiTGFp/j5pJ0ejqmQsc6a6yNJfatd
kWwtsyWpKVVyshjq1JZSp+oSA9dtCqY3iRr3vNWnPbE/JEBSDZWNuUS3+FkE5fEpCA8wnZECiVSO
/gPH1wE2m4f42VruMJVZRhaoyhamh7MG8sgcJxmKn4t1i/kFcQNIW++iV9HadUeo+D/YgSLAvmDi
xxGz6I/65ZmtGfDB1QdFZ5dDK2pKpGopXDInEIwqxX97R2sYAThlQM40dxradpPV62eKUyV/Vl3S
TMPrj/W00ONhtzRXnOiKEt3GdlxPtpdMvmMKnpR0jfK3/Rglz47PQFrweBWUTjknaIx7lcbyyecb
NNpHgJzXal1SYhdgKqgizvFOXEMzI67z1zCzD19OJXbXPIBjUG/UTQW0yxkEkyBswuI2ccjfcOAx
iqNs6R8UGCwMYQiUfAkjUznqA4HaTBcErsauLv+1kS0YNQrKPF2KdmFsIMYsG6xUBgRYVyHxPIHR
0YWSV5FYagTEBjYKBRhUkceACUEXqLWR/aRykzwcviRw+BrVyIgSc/Ww1m+6zXKBVnI36N1yOOB/
vQNZRKohGD3heIMIQZ3xSZ4W2stFWCJIB5DYl2261g+PYXdgegSlODpR6sTfkhWwxCpZHMRTVAEO
8DCxC9n/AxFPEc21W1zi13oRH0tCx8qUowQrOWc8wwsdTtS6HAsuhWmlpCydzvJZ3yVBiZz3P6O0
bLV+VZI6YACDtfmyWUmFPb3nT/g1dtdngp68qhJGd8kzLqJLIZ1eb0udv9HVy6lXmieLziuhds8s
hTMqhgii3kaMKg6OiwlsQoXH16MY8TcpGBjOYzg/eKbk/DZjCEy0bffJEXPb8z9cNh9qMEgYPiaA
rU2jG8/yZdN3uYWb+ZS7XPTip9/jlE0NZfWCNtFFZxGUXH/zbyn5dnM5UEjLo6USX15R2VtVcnJA
xtiPsQKHa8WtqGYGa72bUjNmZGcUCBfDSQXj6NNg/YZuLg7XgZYnju+NabdDUZeTbYrMyMHwJIdr
BfiHDnPw+lHpJrziDpcaIBt2BDvOscx2DcVGEXuvz71zTlnIRIX40Z/xvoxzRsRnS5SLaXpKyqRx
HbHgPFfmPww1ofPDIse4Kyg5La1U7y/YHilUZ+Go0IdJGFTh5IgrZNsArtm3KooXKoP6EJTJ4eor
VnE8wrT5ou6fM3dFLbYkOASt0DCgmkPYXLVrZf3scUvyHfOb7P5z7nOARGqsUtDhiHxGYQeQxqRR
D5kqRFygNMnug76qJl8k3UwDceyXsE4PphmxBWGVAYxncMXyAnMWrqvuxhHTmA7ZJTpstliu2/Tg
HRuA1vMkS6iJx8khLLgj90mAAYj+OPzPzs9xkv6LaBlvy9r0nmxMdpPv3GAyob0lkV0aq1K9MT/B
skO0xXK8zGq3IIu5fDJWAh5jAxyKxpSAxN9gq3OzWYYd6DVr0catXJJNtCEqqNpGTitq1IPS1IRw
O7MiFWVNY16aAfRnFjySevKRVBGxakWRVufvkFRqS+envOq0bs6ZiuQkOURgaOTMxpwIVM+cix/n
1MxemsUrzJEXDg7Ku1jGVVz5j46qnzISyMUEal5P6544nrRNMvG5AnTNFv4JWw+4+08Ohy/H8TqZ
3jty57gem6NB3AB/2w8ylDaP8ywK7sp8ktoTp2wM2rF3yGlx5Ryz0yh5qtgsKVHPsZLkcD62rPVy
3cQifoqDOpzxuLG0PsZ/8HGgFdbtuvEJ6F39D1POEKsbYofT4csqcra8nUnPPqjwpFsJ5m4TqaRl
TlloQdHUogyawNPKX/RZUkJ8ggjFv+mZfkof7aWA74hlrfaEMqZ09piPxD0jI6W4RAzuunBYfQzT
LJGAWS2IRLhrgomV4JYnXoRm83Guc4yn9Udmg5BGnTDRHm3cfgdyQ8ndOu1GYbQLxVei9HDTFMGg
vwBRAYoPYcJeBN+HoBSEpnX5C6WWFtk9ouzpaMCXrYEFxONWPxERYYBArVBSN1tqaoS/suyraSrV
WZiREtZNCNgl4ej0MiDg+5PtMpCeX5p0Au1Zc4WgC4ua2GT2cTJ2hFUjkGwV1IOBH2usDimnJZtZ
mXNHcOUIWMpW6Sgq4F7Df4lIPUNFROEAuUHi3H1f63Km1pFySjhigfd62zh9y9SfSRRB+ZKx90YI
VUcM2M2XTHx6ij2qbC/XbdBYiqM1C1g/1Uww9OVIVotCzFiT96wzaw6egsu1Mc5W+Zkd/kyoytBA
lTCKjNCRpWKR3m4JRO1UaDwjfiAK4t1O4vrBcE8Tp1LfoB5OaA7VJOCQgZaPab0LRHKKOHfKpXQv
3at5SOKwR6MKRKYuTDglxVORIUhX3rg0Na9h/2Ngledbzqbiflqnm3GMx3sKM9am/kREisofGIhS
03kvrZM0jnEhK/s4syDBOk+nzbBZctgNqjf7VaAo/XFUBQIOcwn1ecfwwwH3NRquDp8VP6kqhhLA
4g92A2L4rVnPnyH4ZiTdwpQUM4dDS6xBfbEwFr1q6H7rJlWyFem0euEMP9qg0hOw/EieZlCwAItk
Tt2jaWnVOG+5DpVlqJdmWJF4e/DbbXcVslZ+kPA4bAYADlhtbHMLuyjN1l67PK4Z8ZSng7G4V31z
zPupz4Ks+DRRUfJ+ucceNgPvrApEwKsWkrkbCrp4G8CymP3rzDy0bNvvTM8lfOTv18iCT7KiMe7q
l975rwlcc3CGfmi+m3hHt43WCJEerUvt60CHKVaL8somiWaJN00BtV9G18+eoSSSKMSM9NDD3uz9
kY9H3NPfvITnWfztRpUViMM5YqvG5Oo7aY2KT6Q2+W6C4QIolSzUYL+5tJQt0Y6bqVo7AUGxqSED
crw9w8hD/Lbg02e41q+SjyWlCFsLAObW2dPWEptNY8xjzCASYGst9s6lvP65UcKEO2UTYfTScg+k
tDqn7NeQwb8SnkcypX7i6QE3mtEHc1zhI1vK6zflTiEMGT3DkiYf2hAp42CrFOYyUpCgzWifSFSe
sCZonY3kynvnG3rvlJ7uVqYIclg4ML1HKWG5rXXWTtu3RYov5+37YDferIE1oXpY95pBgWBH/tpN
DuEk5FuL1xdW2LXAnkW32CzXGUzQSxngo6TUdSCVyVLZmiDzjogNU/xXzdFlgivYHGNMRXvCfC2h
ekLOYBLvRp+6V6XIVE/vBQp0LPgUKXXsUVaCyUVJTxGK9u6xcQ2c/ln6qpIPf7hriBpaorCszGcC
poO/wwo3gltNIQHaf59AC2gruN4t6JUoLhxV12YYeA1hxJFfPDMsGXJrcYf8R4MPD2HroBw7XWqc
RUw/oeZ7VuusESM6C3knp275nZlY/LZ3fWN5xQmSadWAVyn5tmeXCOVfTk0KN0hpPsnOlas+9uve
iq+sPA3YLt/VbP4QaVLqT0OBZKxDn0A+3LDyWYHqHaHE1ndRJiW2LdWIeSN1tkdSJNm69YbxiHyA
YExSqWHkZBum88hk0mk/iFG1FJvgLx3pNBMQU/mg0UUaNL6GM6ytf2Q2veq4lFyrrGaU/pHgqaOR
mBhVNiXABOb37c3RrMEGp6J2mos/7woIOwGKcDrHz3dmE9/+DNO/UHsRZRMj1jAkSQuI3gJe5qR5
7ov13xcvnlN7v3Zcq7n+8h5NTxUCeW2LgF3OJUB6d6NeI27tc6v3mLDtMKIu2auohyJN7GCLU2jF
/AUQyFVcv0ybgVvldLfOdfHsPsdYAOHB4ftVKdoOuJC2l2UG7Nxwm7PU6vrHk2W6syCGazTeKPdX
LOczxc/N43qr0C1YcP9HyAai8qHDIttyQc8VprwjctQhCdGnJEFAo81LhdTfJLyVxvT7A4gUfJMc
OXbmSHMjZJJTfV+O8Ztjaz8viYXBK+RGgb2dc8vbLl6/WSngEBVvR9TsXwT6oY+TDInQL2VMo49U
zCFtCrqAjhzujfkKr91nE18TrCsUcKr4xuiXHVh2QBX5r6Og/T128nt99o6SI1aVbTQt5iav93rJ
k1eu/x8oFnrnO4WDre9gTopg4ZWHsPZM+K8at7yk0fO7Uw165dn+v00urEgIC0YsEWNcE+74sqAS
8mph37de5Ou9S6RJdATZSSChF57RCFp7WBHw6Qb7AFwGDwdeV/fDIqmMND72LaAtDIjc9/vsZTi2
C6HLBvadr2uIW0S1DV6/eI4lVQePkS0z7CjHoinhGgYvRtgLDRUpgs9SiQJuG3x/qs+t8r+t5hRN
1DG5GtWJWrrY9qbYONFZPqkyahlhT7PW87gZEhvNGDtDFzY9BhG7V14FTeRdWPL517bGrLEIitGb
7GlwW5AnhwatjGqkCJXZKCdPjyztGF99FvYhOm4ZhXse3NIuVuFZZhFKP5XPTkupPSe8KIHT3J+O
IICuCnyV+PQQTIElx8RheeceIdmNa8EZCGvK9CJWCjael86kUpR3DffyssxMTzvQKvtZuKRm5w2A
fba1VsEgsWa60AFWwsfDuZfpWpBMaR87XTnylAjFGUBU3eFYw8y00bj9zMMljITNb5awO3Z8I7yP
fcU3w9P4elUh9c0TrusXqxIg4j7dpa1ePec+hi8Kji8NNoHF5b6ypEuKzDi5v/tY5vxS+OK7WRIE
BF79NBG9dkRDBuhGo9zFZ8TUbRl9WRnGVdEdHKqe9CZsOOQ/RvXm2MGdVB6412R80tdarD9SMFZv
QzEx+qCRkJ3UZB0VKG8hgmDWi4d8U3zM2w2g2Uvw6WOBtpQGVosXH08popef/nbN+Y1xtY3Y2t3j
Hec1mwR4wzjrSPVvw016yVk01Gr1iY3M7oSX8meC7XKOHUWbSMLG5zDD0JAKEufh6fy+bfykVliY
HzqVAgqnTpB2xhREe6IIEdzj4hiXbldH2d0Q4H2UyuAJSXh4rt1UQiqk5+zFMFmjuqQsVyuaNJqv
AKFAFldmCw8GadYRCBYY3YjQ5NRLAnV41RBCm8UcAIjwqH67w23/TsGyvur+4ulVJZ7KCAkWLBL3
5p+cdFlIJUErHDZ3zJm/QgApmfTxIc3r9FUlvXiU9ytJK5aGy4QIl38fWJnDJDdRyIC5tU3nZ3TR
x8oiF/EyRpTV6KuQLQhQqZFTz0iuVMVZCiMCBOWYYz0HRigAQrizyrNqhli3yaSMJe7PsyF4qX5T
YzMnvMHnSkDa8EugcXhxxKNDUkQYGeKbvJUi5KK47ZjIiX0FKZRgene1Pmh3T/4Khvj0fg/JS8rN
40zp++QmIPf4WzfxELDpAAzAjhCsX/42hwgdsUGgHi2plmUCcPP9PWuCSDbBdrxQTU2WMa8FngZU
h8oHDjdFr8cOEoqaQToOZv54I55UhGjXrz0mXxJxhF+bs7roQux/yW0dwAQy1sItxxHdnkOU9lq3
K7WYp5m2gLvo8qLSkCNbS4wQa6fPIIFkYul56u9EOFTjmKEgADl5Z9tYQ30S00MIp/omYu80rmI4
LJ2O/zx0Ns9GzuK6gGRWXb7GTClCq+WQ58kq5E289E0hMQJG+F8NMkAm4cbcGHRZbugQytqyZROE
0f3Co8wCNSpp6InwB1Q2wxHJ6I7wuLwGAZyHbsaLCi1FlbFSfN5BLZKSpAqHGPVsmzSee7wIJcUM
FSe/m9ePiz1bwdX+FNrSCMxkMC5kkRHKfu4BAGTmAGxEh8O3wkMObuDCgZ8aN8WogGLRZyLki4je
36T6JyEa/g7+WVXBBCmhXkMHktANjp9uQpLx1I9GG4uf5xHOM9NbxHJfEMvtMZK1Z0twHbcsU1t8
zujctQ/RwfkymHhn5ZR4spuBHDf0tjZeUKxTwGfaV4S49RTlXsfksXJNyZt1OJ8ory2HCbt3duaD
KeptQ+iO6fb76y4chP4p+CFpigVA2aAPFDTllHhHow43cenvcye77bkNgyM8pMVkcIHqMCRZctE9
u5zZ5yMF3/guQJqye2QWui54ik03wJI/vmT0UuPkAGfSOOCXS6nXZ6ISP9wYBHk3MaoSKN6DTSAP
U+39i+ullmUy05ghLfvk33QeKwvAYo2QxDOe2ERFfqCWGYtaWVpqUuiQZekfcWQUhptMdnHMBc3w
PBWlxz/hsYPWXZulL0Cc2uvFB6DSo90SNFbeALT3glxdd1wQbLFAKztTxdTykeXW2yawyxiafZid
vsJ2QvoekIsFMxPFrsEMT2DiiELGcG/iKKBt+fwDYEbKNdDfTGJ3ovBKiHtRqBS0qeCdLeggdogE
fyQBIIimdqSnvk9Lv4H4zoQwHjF1mKiFKesaH2wIn0/MfeWrpiH9/Xu/YBlECvakq3XqR1GP7rKL
YOLL9zFB74DINJw/FWHuhER1H6iiyEw2ly0f8JQzgN1EP17paMYapsBNlt9v8YlXEf5TO+tcS8E8
8aZFQ5TSq54BxXmREOtOfyoYUKrkF7J/j+b0bbIxENhqEusfO3NHsMWBTVsF30ax3sGGDOnG2+d6
2jTrQFxHLhOq/o0oQhx+QO9VsecUij5gWk+JA1AnIIQa3Lck8y01UwbArL+46BPk/DlhTawznyWV
NrZus2me4F58lxxEEeFenhRypL8di6Y0YEfHFA5QjBVUT+UBoVQPKSgqch5oJNrycTCMSgv1+TCV
3yZRI4STmB97ebsVFH3HEHJPCulJKjMGqd99aHr5QZea7RzQYUj8fqJ8FK2agZTdI10Fd/VKUI8O
H+LA1Knbz+694C5vc9oFquDXzWTt3fXmQwqjxEj/5oJ5Nf0/H54dHZh8KkSR8GmS6BC/JIB4wO0i
OzORmUaINZ+JX27pAo97iaP2GzryWqKfQt3E7+yjg7opHiVnjR0W6hpKXMUba4fMiIYOUNlfxeFQ
XfE0g1a/XwBzt5FQAaoY3LrR9tFYQGdEAiG0OTObLHOXxbHGHwU9Q7Rw1swDQe7p8k8PaOk3ZALo
U0EakHHYGzYKuzhDujqdK+kVYRIJPaGS7L9iSIx/8EdYgfmOOgsc8MKeyrlS2WO5YYeDlowuTrxt
ZPUD4CpFi2rGuCrpotjecw0Aypw+i8eY5rVIOBgPrIMRA313ZBZYEd4D0kiOKBfG/P3vPl6U3ZQl
PR/XGje651LBuE7ENOeH26d7h7gJWwx0AaKLhecSHvGKaupbljDZfTkhlLVJvD7GXDAZp23u6/va
4iBrn0aeyvHiJic0jZKPqPXop8CUdpb5Nj4hkv8nSZPaxOYwtN9RC4XWE8CfjPUfc5PFo1Ev7WIn
G1+r/FuVKL5LhZbcxDYropCP6qK6Tgb0gKSnU4ZEIS/hteT9ebrXlqBQDbWdLZazH3eh67iO4A08
qh+Aj1aK/zA2sHJ1Cfnp5JFWTDpR/+9p9snkf5K8077KScuKm8bL69NY8gfiWUJ3vJk24YTyQfkQ
k1Fh8040nuJt7AYXr+XsJV/d4NPvO9E15YCsloiWJ+h9H8jONckgVvK4tsuvIuEY/W/DV5mB0Cp6
0nzFkuJu/yi6GXkKlZfXAKQ9Oicjqu3PaFdaJqy37iWjc2fuZ5VndGxMT+ojoDXAwGAUXAGXEWa2
dFabJtc2sbEOjFnCOM2NGqxU7zH9f5RddHJM4pnNv9DIGM0bDK6UcUQoe2qMBykUNAqT8/eNiMDu
/pYxOqJYkEfEb7BKhjbgKf0KpWyzAt3e0OhgrWbmrx+sOtg0/aDF+MXlKQ9qb3k6cd4upuXxw1CF
/29BCnl3MohFvLBQ1BAWHYZYuXCkURkcItSFv9+ag0wAas6pvT+M6m9Iki2UiXU+NQvoAmpiTHv6
rBvsOJi0G8qgr5gC6F+7gQmXJvx3cVrpjyL+hSVQxBhjrXMAlg8EebT8Xl7nlegRisvxa++UgCGi
8BYULWe/8Y8vNRYAGE5hs6N2iBLlgowMaRMS1beA5J4bsVL81GF+QpBBEw2YXE9gtHnqOjPin7QG
YmmBvlWcmv8I2GgtvrEsQF/sgZ9h2EBO5ZMkswG5pIGflIQU4k8NrGv5YOkBWqOew29a109l4qCG
lPLSZNhVKYT1L8P+ulY1aX15olrSmX2Qh0jKjd6Mwt8hLoZxMDuIBqW0UoM41czxfb1Zeqjt/t4J
OFwIb2d+tXB3ZhYpbWDT42uKlC0ZpOKjgoVuMYkttC2KDlZJHoT7n3zPg6om6ZXlsM4/ximimh7f
qoQcss7xeWkuZQJ9uBWWq4nc1BgVVk8Do2VXfrK17hQYfdPtB5tLuYqWlvq1Y3vA3wa6fQdz/2zv
sRCmU6sBAvTr5GNPZeg13EbVLGFnIuIi9XJJEfX5tzcsft2u2/0wGkUTQhrbHVwaY9y2g50UMPoe
CeRJg/qDq10ifldWRc6+uQOHk1dvKXapOi8DYXB5Y4OBkpA089yS5ejvD/TOoxu2hSC/gLxPC/cY
gs8VS/jPsGVXFVAfJrtWNhv9BvTCO3TWJFXhEOCnJkrvyI4LbSd+QDDblAbGuA8XzUi2Imlxg/0k
jOpnh1YQsiZltLsGjQE3/CgBPot7k0V3qGkGmhS4GnpRvv+FDBSwHYdmgDe9RJG96JGuO9aHgpRy
QfWieGgfWAVb21FfO3QF30Kxd+bjyH5kxljjI/NMYiALQ4BQ3Enn6GJ1HcjoMTiKdREsuzDhoWMT
ki5uBcPX8BryfD+eMIJQnfgUy1iHW5XwAlc66G8oC6pveR6o9kcqHlzjOv8UR6fU2s+2rv2WW2s6
NpxxCYXTg7Zd9h+sqH4AK3Lk0lw/mauih7lnyGRaRzLgqjQR3VeytCJRb2CtKyKilUshyeRT2CDC
snrvbqFy7Xo0yXEqAMzoO507azvN79iXRZJuHPZBPRmMX7eI1smsyqYTLmsl4KxnmGLYCfJipyjN
dr+s1Kcj1OEoK5xhMXuX9AVf9mPBKSdoX3gqheZxd56pLej/WuQ/7KWTJs95KfxOoST+wozXWuIa
+GI+/0xSrw1LN/8YvNGF91p4few0GnfooMzLBBgd9U1cng5Zoy5j1QT8Asz7sSMHLszN4S2IFxUA
6qaelUjrzoLSvigE8osWqZNtuVrf2qh10cwCnix2MLycKs9ga7a2l2Y+tpxylZlqCSX3BPaZmMAy
2/9btKfylwyS1phVJ1YDdcJHXv0xwRm9gxDtx/BbK8qcC+th9D8/jtdAYFzCcc5zbh+ontQHIP6i
N0sAfvZcrL3zXicsP7kRwNLIJe1yuoIIc/g/vLrBE8ZPpaRHgFEPsK3OV6fC7U232r1xPnILzwse
nMjUpSALWiR3m434HTkPXSRUIMAK8z5573/0ejUxVqY1CKW3sGkkTcvocDoVT4ekl1pDVSH6pWI7
hidxMpr8zI8IueDkxTOsuWT59Omy5zy8qmwKBB3ZPpKlsSckxGjytzXzzOkffDkBLQhopq+4L5gR
IH/nMk8xdihQt7fXckO/jcrTMHkJ3Jx4P4Lm1QBDp5UOSMOFySfusPFksL7Uk8fhP0SAUf8j7Ivh
r+CxsOes5jU2aFwnBMqcR6ZFl06MC0fwv7iupG27Xll9XJqr/8ar7WOxCa/lDORK/5fntmlYTRMA
08L66WEW4yBRlxCRXmWeGbiPJiQB8NakpE0V+gSL+zExWE1nQGHOxGRUiV/hz+grDblIkI3XYpFW
a3tRmeMKgVkOALLDQrdavmGHQR2uA43GyYEagWJ8fHsGIppOX+XCpCQfTr55tqkwSAtQFWlLu/r6
ksBi55k4oz+mv2A7yTKMN1bIEfik742ZTE3oFHc3cxGQV1Fb06WZAZAXohpbIw7kWWezE+wjLxEx
bqyypqwQ482AGXA5VWqVFaZZSQgy1zwFDbRIywRBrsJOhbDMUXp7yBq6VUKrJDktvkOo1TEjRU0u
mWB+mqangmITkjxGhSfxm/ujAbn/D7yUkC1wvpzx4PrmzQECdQkGkFRAmmu/mp/LzRE1GBWh/kAt
hBIg5mgKmLY7tZVNfdOIjVJa4JpyEC9DjHS6L3U7X9CzrW7eJEsRqeWihHBnIdrAWHwzgM7ZlOL8
yfgPUNySxarn5+0GtCXwdl+WHdo00x63RDLUhA4rwX4367+S5umKLXihPQElOdlJbxfFUuJn9PcH
Rn4fJomPy6vKX/k0uq3TgY7K34KmSPgWtzL6q7zgnlbdQ2ozGqEf7uTpJ9CMx4B029UoGvPrNa/d
lffmR8eljaSAONlEr/fKYxvPBIW2XY6QNuj0YvFdap+IUGSBEjuljONzeTNb2wkLCaTqHOp8lF4i
+OJ5svq7vEk8Gp8ZQZHqqRUI4OUrJUKKvWJIrPTSCbapRnPUkxeJXPZHEk9e1mLAmA62PNuqktAg
Gi1LxSJ5AjYSwWmDQCPQ6qxJ7zTAC6V1nvXK/+hWgBrXdwGlhEEo7X5sNPu6js1mSB8aVpYKKLt/
cQ3o08fuhbe7xKAsc+HG2m8dzRPntIHkgekx7AC3jgbj2GKbpmcOkvoyl42nQMgZDPps2zO0mlDc
9MT9hxvlJbSk65b7yXXhwppxo9yD+hgpR/muvi7MnBi49KGYKTL+T7QWDWpHbD2PSbSSgRED3M/m
YgQc340+zP7kTT3D5WCV+JJhJQ78APS8tliF+N0Z5qT5Wkok6iBXfTk+NCrYCUhJS71fLg7Ml7Lk
el9K1Ya+EyvMV7eWWxlzJVSw8Dely68mcYSL0939RbA1awDQpDFskA7GcPQtUxY2wr+E5gt4RfwS
sAiL9wHhUbucPwWVjgDajDyer7NlYrmTJkXwHhjH3ChDmHrHZ4FSEpqP3g9mpQJoTf9mXZYIYeqy
+tDrzCSthSMkxVV9gLciaxSoPNRfXeM5K53E1tsXf7YGNnoLcbhBHe38w2akihl08oXGpqHYEvdo
gA+SZGwgqaJz4Btpm+7C/Ssc8gfRKkNHtdI47NM0wN6d28MEVRT0pxC5Rmfa0MmCsrZv9pGloXo2
mJn1YpJKBS/6gZ/0OCtWqM1i/SM9W0w91RM3PBUnmYU9uFwRZdMBjODRQIBVK96HtxXHOkgKpwAH
2YkvTVi3U6Xec1b+ogZsCJyFPbs2ESYTYx6o6WnJD4BI5mCD7Ack+mQV1sFKEuZziLQAFeYl3msm
0rHs+Bc9G4nrbLMZx5WqugqSUjdvX0zE0pKFYu4UgN3xWST1s8sFPE3s6yw+I/mGUeb74p7tPjZm
bUKcY57kHcBY/dvGpxD98vlOqt414SNdXA1l7Cf5wA100uH1CqplL0aoNSQxJtxUV13dZr6tqUml
lzEI7uXIfXupEuSY77Msxu6Y86XtJ+RkaWaSb7uXUpGabxmz1RcMxeFQcc4ur6vw6BoesZ1zKfYM
w5WIIeduLfa/p0Lhl4Qr/N2YUbguTB8eQTclnohLW8oIkWUNyWVrHRJAa7yabGFz8Rrt6Qe1ddxz
NM5bUT4t9WVVURE/hDsi09prVYIMiDB/JzHQ0WiJIEWYQCUzWnXQOnMRiM2z7znYtOGfy4lXpyz7
/WRx2TYUUE2x7kaOXX/uzB0UDAXqKCQL/ddnR83MUdomQY6sXw0mAVAtOTYJOMxyLl1NrIAt6Ayu
oSAUxsnikPV5WHzkbpc5245zc5qhbsLfNlZcOP+tgJe/LiwQDtbKeGl0P7zWkOYVWl7ads3lP6Zg
Dqv6wMq7AGsJytvhKwPC5BCbeMxEEvgD/dp1QknkXUYsMcfn4YLPEOjUkd3mfSzhOEArv35gNPRm
1IGGyni0VJ9j0TVG5F9/OI6kB998kU8ZKCOntUkp4ZKyMrBYU5/rSblZFKhgN/qSJ1hMdYx/JP82
piB7V4yEfY8nDjUrtJ2ApEkZcDXIDy8FlSHv1LuxZ4hToayhR4vyx333huC2x8TX67U9HfFU7qLS
Md07N4ewvZfX0K1ZKjOCk773dcotoib37dq70wvEa+518lpb6RwTD6WTGs0ZYygjDfKMOIgiWy96
wnuDCCSLBmEVP2U464s/NOu2aNMHR1NjgE6k+QmovsK3VXpy0Szn6NQJRUPnxjgfMnUO2qRIBdLt
JCUswp4LY2W6pz/PPlcrG++JA/+F26rdNUMauzgrZqX0KnqjQ2Bp9BmgQAXX1kvWuRSarSCzwl2a
Ae1DWdlSQ01cDdSRsFAuzdkiU3XW04Xj8ycdtt8SeDDRzm8SYN+aY9OMP1/uLvWC+NemwMCi66LQ
HnSNjD01kKh/bYyHsyMwXlslUThaMOj/zRUT5Tc9H0l9HrBMzyQdPEN7TmVYOQib9lsr/2NGHWYf
Y7Pa4gNwWEmNjr+Q5q2xMi995MlTqq7GhQf71YrK/2WF6UKiMHy89AF6BYb6A8Q/QGFXa1eSqyQR
OcqH9+S964moW+QSR0RNhHVMXBEeqq3iBsP36RqWjWogm6DB28PCr8TWc4yhE+lz6mUYWsEsmIPm
WD8t3Gxx+Tr6RRoFa4pHPyNU+6NeBo+9oMrTrHzPrAhn3wNgRKd5hkpLbw7PMFFmWGKK4TM5YZMO
aYF1gMQmAeYoQcIJVUqDZpfOpv8485MGZltXEoFLN+IXNX5bqZO922XnHzHZTHEcVfus2Aj4rsSX
8+gmWNI9zaYYyK//jngOtMwSxruxD1d2oV3jKphTmvl4UduN6JYewdsnFQsOd0AABrTW1ynzeEuU
fUhWwj6FYfqMqtTOZEHckB/dGHF/TApRLCkuB6K5wbqbCUyQZDTLo/czx8UNJ+7ElKh4y/wSR6Mf
8u4eFGl8w3JFfjPx1mNyih5SzLVuIam2hZtWDh+MllmUDMIgXw/iEhFTsiS4b2RZicS7mOng3GEC
Y/hLdNlbEyqbHp9boGRlQW/CDkCE2nRgGMsdKGusaEc43inp/Zq+pWHwrBc3vkbnCv849+n3av+e
M/BcFr0AweVi3BvV0+8iSYddCIgg3aJii4I1vvGJsXqowrwuCBXFBbW3JuAfVRMz44lp6LyToaa8
TC/IQnmanL0C4FuC4OJ0s9HXezCmN60JkmqtHhQgF5AqJ44XnNtQojJUNO/Uqip4744gmUsykN4Y
PEL1rn8fJHcXh6omWVta1Tscsyf7hSffEqv2DxPRrhYaOjI6ItKfARyZgSwsVUfyVPWIkTs0WeuE
UgU2MjLAyxxReyACxxnQvgt5INc7CMn2J1lqGsq6xYoJVcT34B/3ebYQ+t0+rwq5tg1usLlD52Fy
hfaMPMa5UGRl065a2gWF4jnc6ept35SYqoS5ftWaGUkx4DEoGcXUyLy7LG6qa32bznn+V1reFZ+N
PAbxm3XP9fY/jSF7KEvpkgyBvOym3UYXZMek0s0qv3wNFi+JNi+547M7+KswDa5IparKgSzP62ph
oRPrdXcioCE2hQmBV6dGERLGEMxo3IHJGyqaVg6VWbGqrn7VX3f3RebllYbPz6EI9N24KrcdblEh
EEAV+cAPhSF4nxw2h2dfgsCo5hxI9I5Bttyh3VCJWoLYUnBy2+BY5BNWUDEJSTfpDXHkCjj+d52X
dIeqEERzV1+scEwyMFwN5rB2Yu+7nkyiy7oACkmiwfe1nkucoDlpZDVEmdUfrxiBKmyFr5exrH4J
wOA2HJVtxIotttYO81WPAWc+Tv9a48ScNQTMio564TrQIYKmFBAsdhT7E3j7pMhse5GsGUDN3KF5
S+GDoQS3GR7uqjeb5i7/SfVeT4JgEO5FUy77j0llEn5OWeQvSTSCfmu3/XayGEIUEgKrDnDxKXqA
J7eDmYpLKBEjgk4HH7en/FHBvCW+Z5dL7ZXokVuW1N8hlS91SAX/KqWtEUqZTWDGnWeDfTeKyG6U
BAJ0CfpWP6gVY020yLFwJOTALFVXgM4GL+D3pqV3eMeSRqarvjP+bY/eCkIyjDvaPri149XeHgm8
aQDDKKdXBR6jLulZu5ayCebYPglvUBplalDaPbwHBXZ6vIPAoN0M8mrdm15mDAz111ZPeeKOfXWa
88BJh8FI/aRVh3JrGjM7zRsTpLEyAw3URt9YXUNT3lJkTUbbOmP9U9sbInInBvOvs6wS14kAIEGI
DA4J7ILBv85j23tob9Of6U3/+CDdm4sD0r3bKjRm1tTkhuZqiaY/Nk+j+q/5PxhJSQ2UjoPa359b
slBnQrJTAjQIcS/wO3VaglGuCLCgCsV5HTAgpRKx/w7JtuIGtbgO/H7VenzzWRNKDw+G6WUZimfY
PN4pe0C7bojk/n8Etn79BNuuVX31LpO85d2Ugr0fJ5mysHm68kqccywnBQC6uWuaCmuA5vqexA73
BtP/Yi050rZPtIzG/g15SYphG3RwNuG9aXNw99iFwrDoikN6HaQaZQA085qx2w4vm/jawqwigyPA
8/Z2wHGvq3lEQCFVgxH2PDZYg2OdQ9u5DyLS2uDJIAwLZ8MuHJREp1dFJ64rc3/cI/kZyThmf6uH
J/43jHIetRrHJWo2+DEGMnSwzAHyBPWv2SeFUK9fzM/bIZm51oEO1YsfQTrCh+0uVVHESl3CxCUX
Jrn224vsh+YJF/H0029eQGMvX0YEANinX6HW3nu7CnDT8rMeGd+2UTR0TeClfrGkrU58w3WL86PB
HcKGOh5A2OR8280Zvkc4TBJfd9mK4ztT8w1UVVpQgPvVy6nryt5BKLvHytyn6Tn7pTN/DBcq+Qod
JLO9cOU3w/QT9M8hjsueyBAIkI8WtsTVIMxmAhoMEgrnoKO0W1wJ+wcQvGlyvUdNPS6JBQRa0rXX
pp9B0BVE18Ct/pX/TMhKplDTRXlUzqerX89kuaYJZB0zy595X+6KGKwvHZnBz6IYcD/KLztQ9lGJ
Aaz1wY1w0ovaT+kj9eZVgmXSTsMrABylkCyjGvx+7/r8Gnk3M/UoWgUAj21qlFWJP//TYEVeuvQk
48PFYhq8pX0iASErHpL1V4BSSS5tbPotNNHgGCVYzBmOZs5HbcpgGYkAs5+hypzLYPEadqJpNScI
54QGfjaUEf0AC2PQMTmfZ/tYwsHdZV7zSw2gHwfh7vjaJHIsJuT2f2+0nvd2shQ28z/i7mUt/ZQU
sZE7xQyiZK2i+smp1+IntrqDKG3kL172LjTzMLhl3+1yRun420Co+dEwAhQAqbWn3s2SdZq5/nWQ
i2JTz5hnuTp81YCM21loFz7R6rIBxX2eCFe7NdCJyibRTOpeNBGMkdUKNodBP2UT0et7dBr2P+bc
nPudCwolZ3umImebvgdKHTNmCfJXyZyuBLfF/MEcLjPAegBnU3gGvLmkgWuibahXqxCj5MgnEYVq
mfVyp9stlcplKyEKYgvfxetoIQfAG2lDYFu+VWuYo5ttHxJ+O9yphBBnA5Vl8+HDZq4EV8EoCrTx
ICJ8w0bm6z6GGqwm/YbxnBU5vFJSjuUDhvHDuMgptmwcgQ194F/zLkF/bezR1GfpsV5FEDc6QF2M
eUO3RIIegQ5NQe2i7wG0DRT/sMWzQNsJubAl1gAUetxSk1SOF8Q6O+BQJx4TjoAeL0leZbPaVrMm
956K2CtNhDPxHtnG9RErIARCI25J2mZkRXNiHJewz3T/uxAsGIxQc/aNS8xDuOVkCj8VKoo2tjLY
ZMxNku3nCfZUQJtsIGn4Wj6FhZf1yfjM7u98VnxlLq99wSrtLb2muNyp87kzR0gMeH4TCcEeThpl
DQSOCGEK7K+inxVW5Rsicjt+Pyl/JUAQnAN1YI2biB2sB/tS+dkX45trWs2vp+1j1nYYU+CxIWXa
35CXnLYIpUfmRf0O847NpyzhIgVGn8ZvbBxvhCXtfI4fAPqRg2d33CQSOi5humM+Ys5dJ0HvqDNR
VyQGifKAupxio49ALXH1nz82cx/W8l/nE12EKEnxoz/Xxuv0sAWfXJRCzd0qnpK53StAghHRK3Pj
8UelLSYDmZT2Jp7pjJJ4PdYGCKHNiWQDpKxGyHxcgFrgcP/FhZjdv77zsMKb2SoUIWrI1ZNvvhif
0UpEajSlOExak7/NWdoyVP12cs1OczCDMmOUgxKR6Rmkv5CiE7b4VhZ/mfO3dW7+HmAdjdHHJfsJ
178EmO7rw/HeXIvG/Dmm41OzVB0c4yiHSa9S6Htb2aWUougfDfraRv7jB6mlJ1v+xunODFC6+NB3
4za8A4fjXHtLlM8ChsZ9tLnSCKybD3BXeQZF/10LlsJ6LtLB4b1Zqy/B3kbkUdOi1iQb04+FFooP
x+GxCRLzzLrN78Q3SaLuHaVqgEWKCrcKnnE61RROm9eWT8dHCKOqMd3XoAXVFWoKXHGEZwl9wyUU
bp5YjfwjchAm/hy8Qoo2xNVMUujx4KakgoqQutsr3PbpA6eZdVJUU6GvcF2/FCqbLJyM4hTqiq1O
YK1s+RzoMUDfNAZ9+/+n/DsSk8737NcVnWrTfk0sC8FKHWViArkbbOzwWxUYPQA2z/K6vs2pkSlG
xDGCk5gKK8PxVoaxbF6BoG4RBmVpW8GCD3wyyKiiRNVM1nGS6u5YtW5w6B8HKWF1GArPa/zudQqJ
6I/Z/kH6aIwVkdfVlW1D3g3rvAK0qIIjd9vrKcquOwdH1q1TTQnve/xLeuuQOsLICqwfipsWprMG
OEUdQuDMU/7P7+0Oitfkp4PePex8NWa2rUL3qMNqCuvzehrq7/hSCO5F6NRoblONmNISzIfT9CqU
1Y45lQc8ZH0NUDXTHPScg99nEMSTiIqH1pPnk1RQJSfvlVwbXVILuecER3VKNhIZ8dbNBR8a4U6/
zOxBWi/u6V4UMnE/mCx9kH1o8zwwsS1RyMjU4hoGt+uoml/NPhF6tDin+uHQBPrl+pgL3Ynx9lgV
3gBcDDS4hRMP4l0rNMwwBKx8bEmdNh3XDKFu6ov5R6EyFkpyHeh7SkyRvKHeCB7RckSivEVIjKJh
XIEBh6M4J9kGG6JfJR2iOmhRwh92wv6VyTxn8xdgChi6eXmsERkKD+qjYV9MVEZ66JMn5UdKovYq
EAm3qOYHllJfmViTDIphA4rThz95PSH09rmfQo17KKliUWkn1P2pMl3+ZTcg97DhFYpgK8H4U2W/
j61f/dviHRYZCs4rQasJ610PZ6rZDPJrGqcVqTlC6yPJ4RCM93K+oqsZZxcdjMUI9QMCuF4QS22d
jIkveDqESs0qRvLKPX+d5O7SOgeGAnwZe2sCbj4smceoaXw9QMWSL/zxqdpfCgG+2Y0Dwt1OrSWS
U/9/Jt/PS15RBtDVSTV0L/wd6KMN6Ug9ODYW3AB4E+aY8y+PkA13TtMchtZpzijeU0jJx8pmF4+S
2ECctpzLxDS8P9RPIFxM8DXNy1jorAuW2q8oYWx6fQhHhvy7W1YaxfZCjshtTzWK4FqFmu3aC/1G
MlPfUgUrBWeyAtrtQ7jPuAjxuJiUM4PzcK6rAAXzDZFP4gCIVxnoR1RZ9FlsP5zCjXZKVlB3CbrX
6fdiu4tjhIPPlyjyPZLkq7pck2g//4Qf6m/Lo1yNzyDYFmeaOfZO1rjR8+yRqfnoG8w5LF6R7DCD
2mI+5V26UDD/xYB+Zlehh2zifdEGDtr1b+W3otFE4X8VSNY2OUdYooZD3QbUpzygfGCWNxM1Ye4d
h9AHfKofGvRhFNZQ1e2yRa62WFgzYAOan1Pr1ipEY0g7PBlw92skUElrWr/Ypyv4kfRg+dwETQBi
h0w6UmxGxDhWLHn2LmZKamqteApvtmSfj9b4rv4S4wyiSLTg/jOIb/qutwt7ulRXSct6zxzgP5Qs
dhujSDjvkfwhEDa7cuuHw2qTFlQK4DGVq0Iekxzj/jjGKsEuuhl7EhkzuAyWL+G3+fbx8VGHCJrq
FQkMwwymxoxLuJ+wLnCmLKdlQsoTeUa2a74QjzDtYD0OBdVDFLNOSbUPI4oWCve1X3TJ8lB8KxPR
ORwcwC9dTh2BNoUFPpsmzdDFr1Z/sWkpztnPLyOLHONy7yhqNy/m+vC0OVDYBd0UzUrH2QstGKiA
2v5dAHnwhkdKsaWDzjgS/7798NVMjW/3zZ1pWDZxxufzegstB7TlAJO91GrhY7NbtnQYdz70ZUZk
ssEvLmhw/j3xDwFYPXcdZZhTCiqC/z/s609uK5Wqn3ZK+gPU668RulVtq7zCGjuad5xu1JLHDai5
6wVEns48dAiUb86kLeaW4gcvN4REotz5W243d8iicVnuzC+PXZDR1uAGSp0Z+6yI910Efk9/4ZBh
r12lGOVxxiZCcTrtpyCMbc31gMFtLb6sfLIkjZVvx7ovKzccfJFY+9WsgD5GmZpEG7Buas5ipPhS
w04ovBNkoNK8wUhY1ShqUEZfKNyL+1HY61D7/deX03E0nS/ACMA1t/XFitVLbLEZ1fCO9x+hAE7V
LGanb6nZGDHn6ol7BGZVvPNe28MSjv9GfPwzrBqjryNJKoaYqPOUwlmxhXfQM3YX0iB+LRv0nRxg
LaMr7lN+Sy6pJ1Lw5AY4w0blxlvzkjPM5L9XcRmhroN8DfB1DUYlSnp31K6UWg48fDIX4KzE08bH
AP5ZUPqGpzd5SMrJxdiyLoDgX4hGaypjf0mrnqfvDeyNojFt28GcF3iGtNCyKCcJcjx6bxPbwqCb
2aWCVMuHFAM/YShPn3fTq0eOrqQ/u9Jl4YspCFbxYHi1C/stRPWCz+lWKGqy0yC8dTr5r/pQXafG
imoYqNPeWIr1kjTcnv2pXE0f9cV7dh9Fg7I/FzRPJ8NbDmCcy73yUruUGXGMlewQspVrepmygVZM
OkwgUrFC4GTnbxoqw6TTeQJHpdqCwgUGNUQWRzByj5XtZ/FzAPr23a3OCEbuqWVSkPSTXq2YCO8U
qq1AFJxbcDjxGVLIojTOVuwMFkCQayJ0jmSmu+4y/9+BE4g20T7wH048eoCqDlPJperGhe2QoAXJ
4LOcWrsgsQlmEh3PGSKTL9bBQ/ucM0M0gh6BgjuuObbcXAqQ79hzI6PPI6OS5gyenoyWSOsUBWi+
0v/baq4UnVHZPQlelVxi/xdVvM3EeWpyvI9IM39rTjnk7QaXtNSAkgvvSSoRf4sReikJXQJBMsyl
wXPsOb1PnnhF2rpfDZtW/jVoPXL0qr/JUWLeA8vEKiC5MMfRAhDaAzf9aE2IfqzKw2A5cTKgKSTE
01/yrysLQm2MH94m37rdDCg15Ja8s4qukewpBnd4TQ5EB0sMdO3162k1aJv/ZJ/DnhA/+kkx5wPO
KgjF1mF/U37K2UxsUAPoo9k5fgVCXZz8UQFmvE5XSf8L+HG45+VcRUbXGJzc/c44y/vbJRr9uNlQ
/bJNPROI0caDjNVfEY+V6OetZPzIUwsEbjySrp+09JqO8g2MpR/p3k9Rgr9fTdcx0gj8KWRUp/ey
BhVjN7npKN9LV9fz7XBT73C2Aa0B/0ZVadJdpMPx/nSDlatgC5i+I1eKvlqJ7GZknVjsepHkUzTW
YT3uubfKgQwNP/d8yExXcV7KZGtOKyKvuo3p1ty4nk2c+LLgFSfOLgeCKWlB0VTRzn7lXggBPSrx
jGZ+4CK1T++68lwSJ3b5vGHhz2X+MnqyrOIBjL2JOwIQAA1xjp+ncnloej+kkNurR/Z7XWOalICb
clyXyv+yxZ0VRSJ+qAICapGxQf2y+MUIG1m1lYBtmki3hk1CZsCmkc54tPRDkaHgqmV4U5sF5Nl+
LqA4LS5ouo0EvJLOa1H+HX+uoo5R5muLs0sVYATN4P2UFjjGhUQRcec8uHGiS2X+P8ueJ6Z7QfZx
VbMopDGzkF/0HlgGhGsVFmf4QNYX6gvk9AyU1eR/HkADh0EgeKdgNsEHSaojNtoAIOW1E6GOJj1H
Qi30gpu80P85G1o9AaPKLSUmpQR2m0nk/qHxKiZm1M5a7tCLfwC9Sbsa1cDYyN8dT5LsCsn1QMqA
k4II8E0klfU7owcgE8mG4FaxJYpa+qnh/Rd2X9PjYWYZo6xxuQowGnPNFy503p9rlKl3bavE5Ivx
CBn5S0/9M6GCsMKfPI9lQOoXEbihM6NQ7N4FaOMBFMKW23MqFZwC91L1LphL7yzT9lsuFKM5ixz2
o+XYFRcRxfwy10m2ZLEG2GGpefKsyXlEmcJpBlPyTcX4Le5V84xNq+Sgw5y/FNs6ltHZgGumb7Uv
o+VbIIlU4TJd0GIUuw/VSvy2wAw6zZSM3Ahlp9LSLOx2Ot1v9o3vs8gJt5REV93Qa3cBNOwPHOJB
g/nNfaWLBxsAetJjn4OOziJZZnVO8Mboyj/AWQ2nUdKZ6qsDYAhzbzFdJlv7nnpni44zi4zMyUbZ
3Ahv6vFc+sqvc5035m0cWl+hT2XE68j5CA3HqsdfSrkBOP/ekTf+ltPvDkHtytal/vrCVH3D13qZ
QrxWY1YHn0h2nrH4cFoInApWw90cf41s/kIFjQU14Pa6DKm7NDztPEng+z1Kmt0kziE6yAvWmf37
AZcWfSyIkx0uRsZ5Jm6eaK7p4BLJmdp6rXutijjnMavjg+f698x5OhQ5L+Y8zc2/7ptGVGLG7mKA
OFsUhhmoQIJmBLYmGg5xQUF+vSrfwdFEEMSijYJzCovQyB+eJEJEJ/54ID2OH6zzWInGaULsUHv7
bEv7931NwjxRO5NARBy0tWo+pUPJw+sbiEUiCKF1TXolYrpLMxcT4/r8iTIQEiCPk6G5vPPeDSQK
emVwaxzAK05JZw8Tf2j0uNQcEdd1OD2+6vaAr1kZ/NglCbKCJJHaBTBrYnVT+VGR6sHVcFbc41vu
6zGZ4fWOrIHgdO6DzXSywXIeKpBSoNRescde7Qe66ah8OnF9hWcytikiKJ/xCUE/XfAhPYvX6UYf
GotSBwDXG89nkFaadopj7k+ish4KewtlcHQpjfgY/IAwvgthoBP/bPcZ9kkRW5mCYPHgP1s/Cwvp
yIq6tQIo7Wf1xinBqcPJADdDbWPadpLz3sV+sQTznyWg4n+LCJsgAmJiV9YXH4R30w7hPF9dnuNh
PfgxkBXBwmls29qzE7gvx12vf40IzjNq63Qz9C1HL7Yymvfub+T+FETxhjHtZQkZbq+bPve7HMbe
6qplDJxmeMheLLj7GSHnYFMyHqX3lLb8BS9S5T0yyc4P+Uh1/iH5D1oCqpuncqG9FK1GNu97FyPP
2fYdMCTgwuAGyOIeIJ5OExkaM0QbthFjMErI/GZfy5ACbrZ0bGQU6QscVm+KaLWAFBpuFNrHraSj
wkMoZAqSbH6us6m324E1i0jvKC87AyFKLGvFrfrqOSLy4h8FgrflqaE9ARdz7boq+PfyOysE3/xo
oINtUp53p2esigG1tn6crg/JwdB7hbhyBUlGXisQ6cMMOCThbm6TON+KXOuv5EtRSutmsx9LeZDB
UoYcQSepScyP+s0hC2rNLQtjbFOB8cpxa7c8YG2uksgL8Zj3uCeIeqhf0XUrOwW7CaRgMc87sXLS
P6X+jbMSr4BNnHR+Ne1aMMEsyIHKsBm4OZeq8QSF/fhiSiNzRv0HuGMM8bMm0dvzKyUcnRA2UQsK
f8Hj5W9s/SilINqWwRJDGVIWxUaVGiidD+zeT3O6hEFFnSDP/y2Qy5rpP0mG7+nP+wvNNGFmrp68
vGns7iv5/8gi9oz4HCgu9FfzbQE2OJMGdbzwgwg10hzy6z0PJY3NVsCKoHEmI8iIC3q8255QRWha
B/CpEDVuDpTnpI0UtY6p1u7wPK9Arcz6NfknC9+MbwgofSI3Df1Ho06v3T3Fnc4lU9tvSY48hE1p
DLpAtSag6AOX9muMwv61w7l0US7cnIXqNAIpiQeuXhxfEpShQ06ceTWVuilMD0uqFXwia8QR9RJY
FdTFAeR4Q9pdZFL+mMbi7cpLUfDeuEk9ELZWW2h27UOmt64hqWtN7CIyvQ3LOJoYKQvqk99iNflJ
6uIBOZ9DzMi4g/iiGdNV99h/SP/hv/cjiUhVBnzaFI1uKWLe1w621OrechRE3dCubiMOWe+JCbGT
olAxjk8AbmBLkub1DFvOZhart9NfGGu3WtALGFcLaK8KVdvgSBbP/Wd/imhyzhTGyPB4u2X3wu/g
TaAeGa0BmLLE5shmktCsjVs90QzWlM43GNmc0jKFA6IwuBQ/frE7kASLW1cvVP3WxNjxM4lna6Y6
8mc+lXVJ/80KalIXWI2SG5pKs9NzoSgQIbNJb9RehHQMFE9AGE8F8w4ZhrxbqeiaZxtgkL1Zc1WW
H3HzhEk/j+eFE0VZhI7/X5R5zLg7fcri1Q0V6uX1uYEp3gD73B3QJFd8GsClJbfAPDivFCmJnMuN
dRv5QXVnZue0B10u60uHadK0a49GpwIQNQoT8X7R0ULdDF17FsfrBBSSzGhLzpmttX2vVflzYrn6
m1Dahaac5b1MKYfT8TjBEy21eWQYt5zsrreVm+M7ykvXrPms90KvU13Sahm6i36JXVJAfubnhzti
Zvc/NI4UURDffFW84c+3DF5xbZs3gq3nBmx6d3sasYjjgaFVpSwn19YC8bitGx5kSGOY5Qky/B6S
KNvZ+JPFuKWxbK9fUcuXyHvo+IIYd+Mb9g6xO8Y9m6WlCuTgKz2ZFCf+hhhYdICjKQlGo+ENIqbA
PYac2WGGGLg9H2DpkJMlZJHPDpFv7Kli+wujrFg6cfPK/Ov0k/YABHHGli5H0RqJRxJVugwv89Wa
T2Jq9rBUPDZ8c2hCmjXDkInpBd8eGJDoZL84enXySiZ1mxBtjXVvrzQxZSSjoVu7qskD/s9HDqJ8
GCTNdVKO0jK+OHFwz0wZcFMMP5Qu2BRw+Cead4zzruCseKxw3TPLD4VCsyq22Pbkxk4LbEmLpFE3
rW/9xS5aSirD8A7Nd4VyHTqdnZeC2C78xm7EI98YRX3ZlbxaTGpSn+WnYlZvL8QY3Ebb2fiWK8WH
PLctb0UdoFONIGlHEVafazLT1xOIpHkF5LrA+cdiB0f7bE+zvBsF3YZMIirz/qTM6fXBKTgjoi81
7R1EbrcupG7pZdhtuRHxaa51UWm+DrcIguapo0UXueqHwzMIiOA3KRR4fZVx5sVWr0prYZXJCaxh
BkS7YjIapJe61R7K7dvkDZh4a6dwpotW7vyTF55s2iPS9txDBnxbKj8oSJXD2CA6ChXGL0uRxM/x
6dOEE5MnopSVdlUHTdO5R+ohl0AYxPuj+rP5aeuY/r7wcS+xbLk+NDWKwIagxFn+qfRuh7qI+ii+
aM3yEuF1tNG1krVyKUtkieP+IfsQcx0wMnNjkonrP3AuAlEXUBtcVGrLZq83jk42xkGfhFLfHFxy
BV1biNcKJMKjZ5+edaHK7q7MTiUn7pQospUmUDEVKp54+EXG1izl5KFjGBkz5c0CzvnaecJyKV0z
/TebdD+EKxUXPGEJVJGIZdD2+ypH5/kwk7bn9h3YU32UXjY4sUllZ8SlDyaRBcfBud3NwCVCgQzI
ZqOMfdP4olw8yhUUuBBOm21AkkN06wmdWM/WyONLLf+OPIQb0LeAmj716sIh1Cg+LyHoa+ONqOCP
4/FrN8tPpMqJ+Z5lYr5f7taCqykf/CMVkmhsbcF3/rkckqZ8Q5ooq0sXguVCjDzjcHqzQGgKBOZ7
u+lq8ZaSdAi4iQxE5rPSBavvU2UaokTCSCehxlEr0/xgKUlGWZUiQUSDUZkmGFtXG3Qo4nmJHokC
nsRWbg83dwMTSxjC/spazOp3WTO+6EeBPj/IgFAo+nizIrcmUrDeB8Hj0Xe9NZonBBhKMPhzo+5d
rNhdj8HMy97REYp9vGtazdSmrpwe5yiLB4bVGNFSzTjNs4dEWew8w+E8OTkKxo7yDzyy0NU0ZGLj
7nAwRYHLtQsinznShpF0apNuG6d4xbsaQdRkp3nzCzBqIAfUhriQKMVq53xXy2Uaw6zn78pRKLLQ
EEMrRAaEJhPQj74/HOjxhYAto9r4CxXJKTxykGBeEYly3RQFLbs5SDdvws/ky6ky3KTuiV4Z3/iY
ALPA4NNC0sQkGKOPso2qGsjsAQ6Ewsnwpsg4graHva8DGnN8gQbsb9cZ+qCERrrKI7LjjgY7YLAP
+PqXqRkaLU6BSVhJzymkNCxtbzKvX+IcmtDNLJa41uvD72/2v83dpQ3rAmpzeLbo0C53etqc1PUh
vZN06Oqh+x3QAT+K1vxBALaCTEF54KMXjb8CfzBiqSSTDKNvVytkR5uU3MIDQ3uVJ43LXK1JtIAL
O9tkumeF+t6lAjEApmnXKFqdEGyy214tPI6moxKXpGTksXZKU87ICigDHRybsPj5954dqxt8aoA9
hYFe3xGCY19Hp+EPTwe3M4uWmiGVyrYXwOWrZy9Cyb8064/iaLqSHUSl0FMjpth3u9rrTfQvPN1M
lEgE4UvA+wHSp7S7Cy0ZbC5T+3GN7uMx5teFds1fIa+DNw1kjy4PDjYr8uCMiTH45oW3vo22jq17
6YIlUJ+N+IT+MQs7YclCeFlSAqJEwqhNr7BhpvQbJAwBVHirSFKDtr6R9c09SwBkrHxqY7nkcL+p
YNLc3o9Nmk/Pki+7syxOrjaneSDI6khWniM8WFTz8X0Ql38LfIvQifrE9dBZFptdqTMMB9QcQQX0
Y+In81QNV9646a+z2QYOO+xmvhLdLYxPySwpo2dFfIYw+Qrg29kTJA1nSwgjsD7PqOT/D5dpB4mS
eqYiadU6eGYxDKE0j+x6TtHNJpnUGX6Cv13dDky9geWj5MvMZKmcHwhElJqNzTTQJtXvSEhrWO8N
JhKPBZFxnIXkbI9coY5QANYOrHGiQ3EYfmh3/14vq6+hvGavvfEr5Gx0g5djIHAWMgxdktckEgSG
a9soUwespcjZm7kxJRZ5W76fXEAI7VACSCYDnqfON8tJ2KeF9VWY9G1rFCGYqo1AOdZJmmBHznUg
o1YFQM4MZTF7bFiTug6LuzUkBvO3YFC7KQg4o6KEKzf6hc9zB8MD6eFntf3q6RQsTyXxTjj8BSbg
p1lhgYGk4Qb3zgtx4uvBrEqDALZbD8sbv3O8ThkNPPXd995MrXZ/ptBZLHRUuwFErCndL0UQzqLH
rJo542JEJ6HVckWyroOxMMIcBmwP0+afXcuJQjjZFiDlSyscZFlFiscpcmEfJij+cF+4xX1V+alZ
k9BHOq2zhIhU3bamtAv2xOYiOxChAANDHQUZBh71IeYF5XomdmDn8Ts97ys+jCMX0+33Lkej/4+j
53vmmeZ47k3IefzWGabYcmVX8aaF/QExoiBJFYC0DUFjbaZpEGjlr1xhO+Sv9a4djzHD23elv02K
KtnjbKf8+pUPOXN5YAS8GBNzooZDnXlkEMAZoZnF2Z8e2zngRaeK0gnOZ2gXQ4apV+559mELOMoN
WxL2jM+sKLqkpUBLM85Gi0TbWPksdOUSvsVYrkPnsUUOTGi6+euzoZ9/fq2AmAgiyKucwdir34W9
NdhChdhNtP0z+A+bElmFA+Sft4QnI1Hxc6QFIpKuK+g45dat3hayMrYdbAhTlOQ6++29JCEJbGjG
8zNfJLK7E3ppgdlQYMFI7UwryRBCGa6/471xvrd8W/LFuA0SQGFs/yoVwtvwc3FiuSVdF5QKJQoc
9PSWlMu3skTZTE7qF/acyCdoihBGw7QtjH1RtqB25RbSnL6Drh+7YFw8U7O1JiNOCb34syjdPIwg
ECOSGaxyoaGoHGLx72NpKHfXzWY2mbjt/jwN8luV+B7hdcNJr1AT39V4kj6HbaWDThSkfbdMSXQj
vDxUIxwhImqX0otcmL24tluvr1Wj3x/Q5PUknMHsZPrDLQi7/Ry23hrXFaoPBZj6/GSTTvR+wQxT
6STsMNJ4DsBO8PNVhqA8OcO9TQVVdnD4MnhoQgtJN1YkWQJuyFMec/VWnVKiSTphKVehdbawx7xk
unH4PI8QvGWb7lHwmmtd/xsEU3y9W+2vRxKWAodJD1NhNmyPB0IRLFVyH0LePyUvEgmmhJHPp2Qx
r1Ls+N9J2EJiBUYXKUZjMkS6g+8WadjaF/S/zgyCml8T0iuF6K5sE93PanrxnkSvD4UST1KynfZj
6K/aY/RVLDdUhyt+nUCJDVkbVoUlO46aQMKIdZAMW2RPX2GHQQ9uc9WSnW+t5ZjA+AJ68nxTgbV8
xk2nYbOmtoJHnPdeGEslvZcZAN+gwiT5+K2PC1/80PsRsAE/EsTxEHYwE6+dxgi2E7nWAqKE/KdE
VzY3AwYmb2/AjzcRLhSRx21rsUQsk2+/b2gqxhMFNaRgVrVXtjS0ej0EaGFWzoi83HdHM7GFdQiD
iQsxstlKitaBKeU/JrOcYAYZeb7aYtXxpCXRC5sr5c/y0M34oPJHLHxu/5RonKHLrCg/hsXzdkT7
+jhkUwVGV5cvTYTjQLgl7lQjY6Jt4jW/OQP/WDhH1C6g79oWjZFtUjbgbfaPrJTgpKbONKctaA6A
NT31/92PHbw3tb3w9aRucn28HCfmjj4/TNhHhyEP3i1KoUjqXgorgcBSfMJXFIZJCryyzM+wCLGB
rls7HBJRw9HEhzifuSPs1dqV3hq+Hfcuu9DoNviCT7s7kS8v3lKn+L9QdY9/DerV0vFeGAj2dlGe
y4+03wYWz1ORLpjqU+7yoRG6tN76GykzrjhxLo5zaa178LGhH+atNo3bbhmAq6sTuSzZX1LW77/A
2aeiJiPMSDPOHHkGkD8t5asJMPdf9Aw7cyDeFOcNc1j1Dre3P8IlOOQivlNrXC1PtszHbjFV5ZFC
P0F1blWWjP+d8PfDppUNucviy0H0AfBb6MolB5V7kivGvZD/+l1DmgCJ4UrvQdwZ2ZbOGbKw/yso
mNHouzDAuIAVJUDVzyusIQpZ2DkTWZBpjPsm9AqV7tKGB6WQrkfuoFf0/Syg4ajYXeEIqyAzjKj2
roOP++SKNVtBcSKHnIFQoWAEiZNmmD2P9vQCrBFhGk95UTURNM9fdEYRfFQKV1Ivhfmmvuno+n6A
omPAQKEHmTDpPHTfIJvW7FPeFDSzmwPNOSXf7hmj01mlk/U5ADUJsUb6tB5JqG3HIBYgzyDiMXT/
cD7zQsVo6OCsTbid8HpPizS6AMJ+O2h8SfLDmqa0SvyJjot9E9Mx5RsXphIQMTDDWiC036l8HN/n
33N/GMYt2YxfsOOQ0YENHXREP5XqUZujyzHBancCeOvqVCOG+dXRnQWKFEwDu+n5AYjw+ALcV9ga
NPdqTibyLkZKMVdMsfqa9Sg0br6ABVBVEHzOAm1jA0r1bs3lnQbTOKb5MtoJpKB4Pn4TggATYYAm
WxG/N2UMs6E0myaFllDpipilJIB2OpEoag3DJILDw770KXBySxkX6hTiOg+i+Aj226VoIbUTvDrk
ZDtXzf1+zFLHg38cNTi8K+uQHRQwy0EJk7NPbxs2JN1E3BC6mOMCFUutiZ/X3YhMQqyXeZknYF1s
fMknAZhjc/qo4Yw9KBgP+dVmyq9/4Sw/MLIwXwJC6T0pMYY9ilN/6BhJM6mnu193OEopodJ5oRyi
fBtbXRxNDkqPEwUkdxRji8Io+q2PhtU+VpJPP4s7z5ynJMumjm+Kb2DyaAeCcafMtJXdsT2/E3h1
NqqEc+cw0dI4vdvgHBDzfz+JWkplEn7V8BYXVWjjUl17vVtfVru7KKpGdFmq5xQCYV992uEYL4u4
PAyZWc08IG50rZ7v83SOyEI9NiW4lG6aeSKy3/YNDSqqOKvlAf3CA4yB11crYYo0eRyHbxXUlBRa
/v19YqbLaoe5BLXtqlOOn54bqg8V0aiKZmnef18HyCdFr7Vi3+58Nmg9ePIZ4gXX8GgtEaK+5/gk
eprRrvmZaEkoTBrUxc9RL9YYTtn+vTiqxCOhhtMd5PGLPfr6KUaySJiBLWjuuMUxXuRD8VrdSjPH
ZhM9I9kyueP5myYmuJMDmk0wzJE2q59YI4AJeUgmFitq4kiMAywk5M2+99/aX0aQeaQTovB9LdIn
j0Wh+zWSRdUzCXW94VVx8CoaM3wruSI0/iuovQgoXyE0eCH63qt8gmG6myIdL+VDKz1GEuZpW+3y
TuxsqCuLm2CGIfVLhQKwcYvrT1gMxi3RAO/GQXXfocy4wk39x9fUpKwMPxiBiaSR+oPzFe+gN44K
7j4dpzT/Mc3sVzUMW2wKDb8Yqu/SFxqNa0QBYJJsW1YHkRBz9NNRL5c2PCE8L7oMaZkpieProntb
lUq5kcUEK5OXnk80TQvJfxG/ocDANmjlrgAxMUC4mGpmvy81UnZ2BNbP8uXV5ru6eN2PZV7zvEUX
CX/nT17/nerlbOppzklcrbLAl+37XB7CZiW8rBX61ZwIwYzw/HERJlQIWvx2TErD+qZPbmvA/+6T
VP/f7NcFxohRQOZlrc2EyUg63gBb0iGshdKhcga9i91pcesEPT36EBhxfSSrO1NJCWnOPKOfc7bd
T9F5VRk06f/rSD8Lksyc0XWDuQmvEL78EXZ+e8oxGYl6gU3Jg3fivZXaDOQzhuXcIK9so+9Exgpl
F1jiAq2jDeWrGfIddcIcImbae+CTJu1Y+u1YjBygxmL5HqVaI2iGASKSSv+TyAuFp9kvyk2umajC
LVEJDwCWanoxhUamW70YcJwQ2O2tpiILRVt9Rn+zWfFVcWBaOfDav8OdJCDPF4U2TLvCZplh2I2k
b12DU523c0/ImiiJde5ADmUbbBDAImULroX4bVceec0aAMyhWsmGS0GwcmpX7QRiFHi004Oh6R5C
wrPiogowH5PaVyNas29HEbgxtcS3Ep9A7CFHrqFfaKp8EA8oNyLUPMrxqnQ6wg/1a05B95g1+yRy
0yKwdNU5jHdS1GysOWGFEa05JkI1pG8O4H+Laz4BInRMUpDMng8P2+1O1+Kv4tkjBSizt2+iaaPF
nj+E2VrJW3VMDZVZ/anET7S/5EPHq8NY3p8xFLXhrFlFhk+IPIBMEnh0JKlfGQbvXsnQygVK9m6a
cR7RKY1aBDWfcvIUCFYJpCCE+T4SxFdXlCiR9kj8EA1wDkuXbqySPGmHpJK63TNw/CEkjXARHaCP
Bda6rc78vaweIzo2pZb8icwOO40CNb8tTGniknb+RIJeVXS8T5ICkQmOvqdWJh3f2Jtn1z5a+TM8
WbNMO4rH49auEelW0NaKrGww8S0MSFzSE02Yp8V1r+cClpe29SahLoXPzwymghj57dACL9nUuthF
QHsXTy1+nKC9O6KeQNzdppTzvF+t1kBzbO/oPiJYuKNFPiQZGHlQ3eH6H/XPIkix7ugAeq3xwTMd
J4a5uT0VKv24TuI2BTkZHeF2lAkok+M/yhsTl1XFBzX0Bx1W0ESitPkDtlY+1LJJ7KCc+ZUpmaSe
YpYhSEiTjO2myF40HVQAnx84nTXRlFYkj5rmkrUQf8/eB7xOkrWAV/IeCA46RusJt0kfNzEKmiKM
Mfc31Mw51HM+bgYkfsi9+mN2JHgOE3vBNXcVXGvbXJbOT9jj4M/2ycr7j8Unln9JFUME6khpbYxC
vzwxwlAjoXMZnaoPOQgOIkm32X2/KoeaZbgBAzcbYs54002gdyNJQq4pL+1+md/GMunqaEMk1yi1
9rLMBKERyfEpKTEDU6q7W0Un3D+WYnH1OQTlDKyuwiwBnognNfimAwtLC8CtNWulRT2LCFxx5eNq
aPqFgDtS+PSnWusEwPW5bhaZq6xoN16h9QgUhMDNhK/WutXmzY4PIqW91Bw+9RdeANgZCdFVMZR/
2f8+3DT1jzni7YLF1aRebZ7RlCmTScMzIQlQ1cGf73rqFrVXm8VqKlbttKIhF0kySGDl98ucRVcf
GYlrCKN3/wxBHyRrJez6FVER2BY7AybtCW1YEDyi0KH09lec5/fHENkZrjfkMhTol3lNM6vof+94
qVufK0pionMRxbYikSyDilFp0iZI0rDLCa4VPfmFwcNVj/+ivXrDwKI4VIbsIwYJhkI+MOCHJ3E0
XxAY5d/RjwTFDtXea4Y0b6Fns+0FkssQQKmNG+Gm3MCW+GNUyctRJhPDtr/hbgMe8E4ZfZYz945N
SQ87axJ6tAK1tId/eTpVbHJ465d356dSTqLpnD2tNB7DEnT6/+0Ee9DfFcw3ECoqNhOURFVUYHrk
mVRJuxx4957dThQEKrraBatyNwDXNbmG+SHTT0sjY81P0ek9w+AbTl6rj+t6sO8WYunnXCJR8fVx
uQrec+PS0sw6eLm5NrFgl9TWprEm4lIf6bNQx9MmRJcAH1rCCsAD6yDTGcG75KrRXY01HoyjK51w
3x1Xn424kPUtjTf4atO6WEIVI+KQbDRbRdMzb8/Gt7Lz0dTFcbXjD/7UUewD6rPbkGU28CLawkNu
0y0o2XyUJSPED3JQdDiS5P9CthAskXEi5mv8sbzL5iH3IyH2dmPMw0Yfm3ioN5vk36yPB+iSFo6L
8nloMbz5Y3htmD+zkyLRC0SUFzG2zEFFgvKjXEqdtwLV12AzOim3lDql43qLU9LGCDsoIO2cH1o5
9Pw3D5ShQVU/436J5pbFi5BoJy+JAYZmtik21pRPIQZi600mLMBkO1LPGKiYtaZ50xtxKdhhVyx5
3FKoeM+jY+G3L//LbGI2OLFp0qg0pab/KgMVPiJKxaqChyB1Wis8Esg2C+k/kF5Px4gR1KzR3By0
mi5vJNhGGgXtvWfWbBVUCNKPHNn9LTU1W5WeIoJ/nuE4O2FbVUYG3oEzTFkGKC3+XBaW8WproS+Z
Y021LTdgJ6kj97ofsNkAIvYHtU3XtTKt9Vly+VB2xAHQC4SNSk9NEWdDhMxWfgAuny1bYhVf+sTH
mEcqdsC0sCRw+wEU5AUXBtDlgwevlA1vaEy4BYBXaDIDBfOmxSbTjCX77LCffNhFKYRkOpwAwFnh
dWMNH/9aulNLwUo9iKvLo+wJyrwJJtMU0B0vLwqNDQwFcoJcAEPw1a3VV0+MOxo0XyR3tnBp9vXy
PjztfLyGsZSEXvdontA4yDFQjPw0uvctvAEUxxcBIcD4QCBGmtznJDBNpmZFjAiFnOBs7CdqY2Uc
schvuKY48Xsy/BJS+bV3D+z8pIDf6dUKvSXWmUiwQLonOe7L7HwSuZgiKpyUrgtFpDVHUTCwAX2l
HzGiKzfBcJPCtPlan1t+0/jQ5EalP2A9t3wZHwXKx84ZB8M+6sJidqYfdVjZTbJz11YpD9Vm0NzE
6xK6og31HxItKT4FRIx/JI4BZbk0QbkJyiq9IJrt9WJ3JaH3c7sLp6za3C2/NoXeYQhw/Hwf4bJ9
I2fuq9/CQ81BiHG4WU2I3bnjlyggtf5FOmTMAmEGuRe3KEQhzbdnBePzCYd3RDdQhw0hf0rTcCyc
8RM4a1M2X8l08XUrNIlmJEluqebdAOLpe0yp12ErOG8rHHn95JRFNLNh3/l1bslC1IR5YMibSHSE
rwSPX6H/cx70zwAbzbFa0MzGgzjmDZuoHpkYfnkbYGpqFIrWzcH/Qc3JecaMqlVCOaaAzXPjz6U6
bBWR1SKJbpdUqqrYyCYYjkAaNeX1O88iEvJCue9LRK1ooCBrjrAjaeDnFaTky/l2n45HPH9pDu1w
ASdl9DI2PV7JMl9Ti+OUwLkhVzJh5vbWsbuSDIqGo9kzo8EttU+653S84yl4BOxltScSd/ME/BLC
Mdmj9egjNMtmaQzqJF7IxpkB8xnimGOxHYsQaiZz4D9GFe9jy+/lSq6Rm3HlAkUx+GwXG0J4lsK+
Dath3aH8OwRXdczAqliN0LhvCfro5gnNY8tihqY4PUEcZjvmH82jlOoRNsJgfJW82bzguQakE1KW
SQImj1BTdbmAY1l0NWwc6DNJ6+YDEQbgqYpZiDENVIe+VQJ7vDHYfLyLaVkcaCLHtvUvDRbIaZZo
DYF6PcHGy+ChUgHIooMR40smV/dvOyKf36ohl8K3K93x3RWzs2ukYt+SLZT3+CdLzNfPwFT8PAnc
3MV7UyB2sDkRek3tpowCtFjohTX9LIfEP+UXj/NTvbFYEIC5DQnyKCK812wIDya8xstP9ZDurlOJ
0RWn/l+6MB5LBN3KM2ZeEoM08/V+7+zerijOLVi86PkwZC0/AtwRF3Qhg4QQznz4pcR6I/8IscR+
GlJrf927UlQoi03J0IUaxTaIf7Qtz3xCpQFn4B3Rl3QXqAWISdjdMZnmJIU9y6In5i5fxlKq+F9E
XKXT/OfU7JCgVYQGlRc6EoaSp+3Lr8HCCX0tgaqx/IX6cchiBZ7EmICJ93e/p7YybU9PaZxZPMlV
EJQTnKcFEQCz5VGvLWPi8QyqlIzX0P/l/G+6mX27UD/37TAxCIWjGJGw6fFcqdYquVy1Lci+Cbwx
Zmv0NmFzpqQ5t1mzUs1iqIHITBD60gjH8tXCEuZcIhIs9UetU6gyUp9r9OA5we78cjFDggjjygOi
406buik1sV3HNKQWcaJUt3pvnz+pV1SPf8ZEhZlxn0QENxbwhItRKYjpy7p3nCtSYnTsjDBQuAqG
+Hic1XYXscJWrR3mELio6HrC4vOr1qmESjn0mdoUg4UttWnYgJcmp1pKUo5TnNqMfuuJdiOQ4Sr2
jo+W2bOMB/ejIiAFnCv5fIyQSoKRv9X5GnX9I9GwMvQhdEWJcC4Gk1nevYxl35bW3GhvrLKYD23n
ETQdHPiUbqyZvRx1sihlHKWmGl2+WShNOBgHQkZG9ukttaxjsfqpw+CeO6HpxfK6ZPV2rF7YSgfP
Ny7nROjj/FylY1BeP/2ZPyQMvwyJN0RiibqplHpn+uMMtvWF4tllBLWFZrwrftVYvlz3pMYNqybF
H+Sfx7q2APjsXDpFaSf6DJ46Bt2+cF/wFKKyVJOJrdRBFsHWw7Ane2NXR6Bjf7UFkua3OpEUVXfB
Jj3Fr5N8uV2gnbLTEFVBQCHN5s/1ir1G6da3moIS7o7DNrihn9aPK2YK+CzeYgFArxjm4XvCVry0
hVYtgmJ8BuvirlI03Wqv5CDys544RzrfUPJtNp0gBNPkcmgn3m03arXNyqtQ66vOVKRUgzLNETw/
QkFXGBSyoWocht8ryfALB1y7xGAAws8oeaWmu8pkENz8jGq2bxnxlYdJyVQGJc2nFB5zF+jmBXZy
J3kWhIyznPooqT0+11l2MMFwwS+pd+qH4UTSWI0Lki8RjlVf5YolYofKDOpKuO+AOL8XPmwn3j/Z
6qYVnHgUhkkTYlH8Lyot7P6pHreDZYgrbyr5MqDf/5276HKngcPKTxiJiO4fDkjLae+CQl0Wb7XX
NFTJ82YLJiDz2K5YHGguqt7o/ZPPOtGAofm2O7n3DIogFw2l1noP53lQEVtqmcECujaDL3xcDwjO
+OzyhR879pSL79ZxCXjRgm1s73fAMxPxlEPsM7bxQiLAI0NFYlebXaAq+7kuIrIGE5GwCBC0d4du
W2kIqC1ZVquROQxmZuGenBtlK7Q02lfporXkD2/3aN3c+pxiOp9e25ejt4pVYb4jnCyo6JljwZrq
OQmgJD427DHcUOgJUHSTdSq6s/SG5tO3JHkclrxjyrn57WiR74+/JO9NvaV/afCf6qT9/g6mACTK
PEwFLGL0fJwmtsI6tBKsEVarQPQ/QrkdsQrATc/nG5V+k5xMmi2t2RBuUkoyfFO67z9Dv4hBh0sV
xa1lo9MCjsQmbxyAif/GBl98j7XCYy92TTvD3QqIxroviz7rIpsGxnwR0eQXEeYsyMOAUohqvE6m
2jf02ksWDuJVpQ4xEZnLruhdU3cLZKJb/iVmGhr7WszPtmPh4/SFIazLHvaYR7rZIGiS7nVyZ11q
4p5OLnvjAEZxcwa95aA2a2ghbMgJvRgjAwOKyENcviAZ9icdbKtivgQV28JGaeCZb+hCjL1gii3b
QXFYNNn6mOAcfCTfqFSDzEIXO0nulFWllZonCqCpPdSLC7YGWheqU9TBkZBCKsT7lWwy18juN8VI
A1fhNEkIJecBgBOa0pwuNvezzpBfbGoGSNgm4h2P6e0C9JVQpJ1+K836a/OX5ssvrQ98VmzI81YF
jgXyo4/qNqAhoIup2OhtS8Ek38XnWM7qX104x0G+E+aFt5HzI796Rkj/KTHhKPhNvkaq6Mvo0OFj
jzSQN1FOK35Rack2Ky/8ey6MV0WyaB7fi+PAwhasiyEQhPE8BFPufgRJBW71h3p6THGCiDvTS8Jh
Z7q1pfQJauuL52afsansS0XU/rzwMBnlt6rKqi2kmT9FR91ujrTEV09E2eZqLStfvrJLX2gZB5WK
fHCzjVW/pyoJ2uuZUZl8Zm2ZfuICuxmn4uReEiCFsM/WEKSLlBOWrF84K+QGwoBC9E2zEi/SYAi3
F96sQQBwfrXhUq09i0yFZWB9o1aDKsQs1bdgaArgmU1osAOwIlp96MEpic2b+n/TgxzuAieP09Cy
r4qytnmAXDcQ36eTFZeZwpMfX4JCGyC8gzCqtrN6CI2dPCp/aRxZskZLVEWaqMLp7FhX5FreJjxm
wt68v561WrXfQtcgtu1n+mOwjQWEpO8iuwEuzWtvJCDGFwZAj1L6lu8a1MqUDPbW2yTNcJ8uU/qU
ogjO212VHm7ws28QX0q2y+sE0y5M7NtyvydxA4b0j+R8pHe52PfpVwaETS84/Y41be9flvaDlWfD
Wqy35XfAOR/XHZAWUBIDu08p0yx/LzGallhwuW49xXUr9NdJikq3hDGt5W0740pFunRQemz0XWXz
VLQLTYJxCcmqSmofqhDt6jMgMBAU
`protect end_protected
