��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$Rx�y�<��wA�*;�x���@�̦�W�X�fa�M-$u����n~�%���P�$��W��kYَ���P7�?UMfT��q�6�U��k�>����~�\N�(�����X�e���/6U|)�X2pF�]$h���d.���9E�	�IN�f"�\��e�z�y�b�����Oo2�?�qˁ'�͜k-�K�P|����y:����3�l�d���bl��ˢ_�d���kx�rq�mh�MذM�`aS�.�DW�mS�9���Y��+�>��!��!�T�uOB���,��\L�7m�O��W���6����'���j)n_�I����2:��$�K�2�Sʫ��l ��!���{�l����.�j4�	��很�̢=�����N��s���s5���_�R�>����ТP .W;������	�"�מԫ�����]�#7@O+?�⡾�Ԫ���e�O�\A�	�ͼ���ƹ�d�	@�nQ˰��E؁Bf���|D_�%au�-�'���w�*%��"AM$w�*4���J*!﹦�2�N؞m�����Y�#����^�K]g�y�b���8����/�~ ��!�^�:3w�P�@T�Ea0�!�x��9[��y_�t��>9c��Dz�>�XR*<�	A��']�T@�mj�\�)�bU��@�?��E0� ������LԒ����35�(��R�dj �*����q��S�G��)�r�&ƙ�ɹ� �6QB�b�բI��d>���(*H�Ul8�%�o��aK��Hi�k1ތ�5Pӭ��/�i���<ɡ\I�n��*����:����W� &4�b�GK�Uh%�?*Mp�#��<c_�w��#I^��r�i�/:!�贸�D}�~��n��)��� �|M����t�4��v��H�G�Y��uQ��K��V���g,Ͽ�#̓�����r� bi��W�=��<��-�,��B����FL��CE,1J�7$���e�� ���ojX�d��:\��)�b~��ߠK��8�L�Y�듄��� ϰ�d��z��ٸڪJO#�9�.��S5~0�mQxW����#�T+Cr,�)���&�x��������[��=���J��h}<��-)u%f<M��bM�_���0b\⽺z�Ͳ�� �u�R,�s�Ad�^%�u�]�Kt��>�:�76�CZg�ɠa��$�G��}�(�K�|��P/w���kx�@VO-V�cڲ�W�g��:��-J��8��F��O�41�.�,�f�Z�����j�JKM��!#b�*�y�dA��D�p�B�����߳��"����p����z�v^�k��l���|G�C����x�� rF�\g�o)8p����h,@QL�-M�=7�|��G��<�G3ɒ����q1��sf�k%G��c"9jt���@��b*oV��#(ty�2w0p�?s��M��[\r�+5X`�.�?�9��7��H@׍ӰGd�O,DSn�O�*�Ӫ����Tw�[;�tb1l����8ĝ�SN�X@�N|��lN:ַ�_w�Xo�=���L�z	)�3%��N���5�/.��, B�w�܍����6W1 �Z�������۵7#"�6Q��Đ�;|վ�e�5r48e��p�w�LӮ��tz��R_���H�����7���n�l�ʒ�m&-XᏢ��Q��{���9�q1�T��5ȚγN5(�1�u�PFN]3�R�d4ȴG欇d�\��Pu�0�҂FT��)*h@VYcGRx�Dhw�+*X�d7#~��Z�����e8�����H翞dP�k�8G9B�͡-�ғjF�4g�IF ��+*@`������xQ���\�`�ű���$$6����B��ȇ@� ����뤋��w?�%�O���x�A�4��	* �N ��$�����{�K���徏~�v���]5�8������{�{I/� /�!���!��_ڝ�����%�d���{��ԃ��S^����M�*�-gW6O�[He��	��=:\��
WY�\>����?П0�+2��ᙠr��,a�p����Bo �J�'�:,�*{�1�_寺�R���9p{^T���(��4�8EP2�?��t?����������~���cÄ;��#W�w����H��UGV7r���i 2b ��5�ڀT�{b�G���4��Jy��ԽFu��sy;>4gi��� ����6��D��!.-\�e�=ǉ{28�<R:ɢH!Q���d3>e^f@�x�g����7sH�0��x���Š��3gL6��2���$�
 mjO w���Yv2z����f?�-\���^����|�u.[\��	o�Mf5C߀
�\�K���K�*���O�������	\�.)��|�P	w��}"C:��2B���t*`������8����A}eB%���ݙV���1HCG;�{r�����a��E
F��.��I/��|�]n�V��`��j�kaZ�	3�ؽ������^l��W��&�|02$���W,�Gk�[vG~M'����N
�?:'$M��(d�T�?B4a�[_���J�v�.�NƑ�� ��Vt������}8��}�b[
�	�������<U�W˪�딲�ҙ���M4�>�v��K�۾�s��yi���ArL�W�K\V��t�q/
�,�WW�g�B�kg
�x�*�j�˶�m��nȽ4+�B��]���ZZ����Ȼv��\�m�d�m`����/�.�}�3�����[��6�;���rC�4�(u�d<XmQ�3�����8��<��'�FyΛA�[mV<p<7��`����B:q��F���{hHd[I��'�dX?uL����}�X��;<wZ�rd)�/;�[`��S^"��N�殨'�xMU_{�	�ơ����3���t��#/��|C�Œ����p��`Y@�L9�K��Gfwm��V��X]�7�|I8���͵�h�!5�΃.��f���8�F�D��z'�NI���p�v,�N}3\��M������F(B6�����Cń�L�ZR_dO#;�%d����m��Qk[�i'>���\ߖP��w[.����r�:	Կ�8y�K�t�������1�o��U���fk_�ZUifܐ�Ҳgf@hoMH�#�3x�d;Z�V�=w��8�Pˏ@�bc��J/3�?�,s/`lx,�*�M0��X�џ��I�/�����29��ٳ�p`����5�gi`F�e�ݺ�8ȠOўB(�g>��u�(劘9�Z��(|��n֕����a�w�Ȅۭ�5\�G�&p�pW�G�4���掫/@S�Z��HΥ�L�>Ζ,/�=�?��]	Z-�tˑ/������鷟��N�㕙�gPDq�ɟ^9��D'�V��E��O��>C{p��K�`�IP�6�cDZ��y��|FϤ�Ky??��	�#���������.쟅�* �ӥb�ƥ����a���d>�[ߠ��Q�7�Cצ���FMq��/��k�)�K�J'؝R[?T�&������ՠC����k�w�?�����{4|�M���_�9�5nΎ�ڢ�^E��.��Q�����h��j7Ae@���E�<�ȥ\�������t��B�}R����΢�905zd��j�lu5���%"������bW��IJ��˸�����
.��D��ui���I��O/b��@�eu���dSVw��A�S	�}�8FV����I��� ����ӟ�2�Iz�i|�\Ih:�^/l��`��q�d��[uW�b����"�9f�Ɂ��j�m>Իoꕡ����͸�Ĕ�l�M5Sa�-#}��j
_	��ƙ�
�L&qR_R���@�X��c֗?l�ƪ��A�HE!�#C�m��}�V��q0�|u��?}�w��Pq�+ʿ5����R�ӽ}�tbP2>Wp,�uԏ�W��˺5Hܪ��?�B���Q�<L8��(��n�e����
N�Ϛj	��z���"kb�o����F���*����D?~�Q����x �G3���4y�@�;*��p��0gR�P���/���@a!�"G���
7Zl�V�����H��%�5���[\�&�/յ!n��/���'%�?��̣,7�����2/�o��gJ@�!ݜ_RYU���V˨v�Q�W�"m�����O���
��P���z��+�xV�?�B���aP�
�
�Z�e��>7pEhr��3�RS�׆Ef��
����)���d��x�!�B��K��{�|BR��B)l��a���Vͅ�
�^�E���6SĹwV��Զ��yh`�~� �)4�tb�]�WFЊ��u�z�t�vSτ?���L�k߫�0'a��ʯ�d�@ Ζ���Є-��
�/M�yק+�h'�C'�Y�p�b��'��(R�:�C�����H�j�~��R���:��G b��3��5t<ꔃȵՖQ6(���Лy-���q�J~��j�< �vΎ@��Q����{f�����n�n���|NQ����}� ��\ͱaU}���h߮���9�s+
3ҡ���i��������zL�^B��t��u8�p�D��-#�*'C�Ɛ{��X��^�5d/�E���7�(�D~�=��qj�d#�ܕR��<n����Vd��mTb��H'h}���5�D=ԊXW�B|�"��>��G��E|��h'���IE���=�ғ��g���ԏ+C�u�V�K ȣ��Q��x���#s�v�u� ��M~O�*a*��(V޹�[�GBʝ�Fc�.�����w���ZMnHG-�n�X[�!�|4�#-Fk@�_�$�`�u�]�2���1K�O�p)ו^��ͷP7��&ar���x�f
Fe�o�0N�ጭh��;Ӽ�|z��QE�M̌āJ
'�Q�[�
n�	R�Y�b�a~ZX�Z-��;��C-�䈛p�T.�����^�l��Vʞ�� _)�,}���G��G���7ɧV~]�D/L(�ML�M�"�L��:�gR)I������A�.�.V��ii�c��C�iA�lP�Jv�"�o)^��/ͨ�P��+����ɓ�����ˉ�@��(�ȁ��ւ�G�m��#��Е�Ǣ�=�D��ת�MZ���{� F�uC=r�o���%����/���}��± ����9���i��,�F�߽�]�IS�&���6~�e�Ƅ�`	f�;:��3��h�4^gY/j�	����X���M°,掘%ʴ�=	�y�Kd��i�U�3��`�ܨ֘����e}R��;���M���5z���A&g'.��9t�פ��`�,�<���6ΓY�^+h�+��p"tOĀ��>v�F�%�.�
�F-�a��F	�tu���A�2L���d?b��oa����<�3I�Zv���ԃ堗eU_�=��M��'�m)��6���%�	t�B��k�������˰P��	
[	-/�
�c��D�]�60v"�<q�q����ʃG�O�E�/��L����kq��V�N,/����·.!�Ek����Ƚ`h���f��=ذ�r�Zx�D���L�c��tzF�m��E��ilw�7�6�`?60�r뉥�#�,�Y��Bm�&k<Gr�T��@pR�p�)�b��(3D@�q��ʜI���d� ���f��B��e	)�g��*b�,�h�=��zX�= �l�	��q-�ϥæ�k�O�1rBt����mN.=�k�B9��e�b�r  ?J�n,�VЦ�4������A�:8��B!F�o��D�A�dT��=����b�#��-���*�%Ḕ|/�3;b��ɐ�,�|��r���!��9Ѳ�nY�+��$f�w���m#�9G�A��&�>L
sD�^�]��G�z�\m���;�v���_�XtB5��\�B�&UB�F��?��F���;�{��Q3��F�_%Z�q��7�%�m�[�R� u��,���^�;� �a���j�B�i��$a��f�-��?�C�Z�2�!��LÍ:�ϧ'�d�y��m`���ǃ[Ժ?�q��Rvlx՞E��Hߘ�n�z�]�j:�X{��n�I�{w՜�K�-��C����?�*zd �\Z7�,�3���W��w���Kᆙ�Yoq��"\��]�zk:\bƴ���'�c�z|Z'hQ���,�%�D�8�饌��a��<�~M������5���Vt.ħ��(	-��Y&��������M�M	 M �U4�4U��m��W��0�'��g��ľ��1ϲ��k���ۼJ��Y{Ùw�v6M!� �[]��چ|@�sx�M�1Ҝ&͝^Q�>]��z��W_��	�؇S:��%���c���قs>�6�Ӧ�R͛R���ia�v5i�T6�5F/n_���#K����G�h��T�Y1h�wk5{�o�*��)�0@<�Rf� ��9<��F-�cB�4��qa����4W��Bx	��������g��-���Y3�qФUbɡާO�͗}06XG��Y�.(B0*��V-?}Eb�截�vA1�����j8���0s��$I���[�O#p����P7�!����b���]n�Վ���;J,9s�n+���Riˀt�`sd_Si[b[���c��Vp�_��KO�_��Z��
��<%h#�� �QW����*s�
ʄ��h��K�Eh����i�裳�4�^-�)�S��@�z�^�V�5py�y.���4>�3 /~>��%@�8}f��¾'�$5ؼ�hr��	̨�/9��[��N�g�S�%�Zs�t�#�J�n�c!k[��J(�Dҙ6�Wz�-Sqf�ɲY�zγ8��2���3P��G�,��%OF��8J����):L��S"�K����3�n���@�/��2VXr��ȜXmN�e>{��������3���TC]M��M踒��moՓ�m�?ūS�1����$�K��I{�D��Azh�}��,p��k�����K����XBSև�fEr�q֫OI2�5Y� 2Z^�]U`�[��cv��|�t�p���6l:�;�r�<�2VM�V�����2�����$�Z2��[�H4�	��'T/ȍ�󚖇:�vz3=Ӗ'/oރy1���#f�
��Wt�v�R,�y���������"���1v��@:���&'���L�ه^�,gF^4xd��Qw�\�D�� y3��hT&�я;��T4lG�^Ϫi���N5|=AB�ґ��;s���'�ޟ�b6��j�C���h�%R�_�˭Ԫ:��6��\:�m�a��W|畭e��_���c���7ټ ��_�]�dH�V��;�2a����ya
lɇ���g��i���2gH��r ������ֶ�)CHW�%��p�"w�7A|�`���U�����mS�Rc�w[ya�v��W"�K&y��gZ�vCH�R �?㯻�B��Ab����V&`�,�tE�'+%|���Q�<3�e#��dV7���ZD�&2��u�l�{�ҽ�Ew��_�&5�)䲳���Ԏ?���WD�;����'6��^v'd����-~��_K���,0�I�e�y��c��8�,�\Gc�	'��G]$eA	�%�����0s������9����]z��e8A;�6�i=�G9=@���U�C�]KQ����� �qp��P�ކ������3��$�0[�C-���jk����=��N�Ҝ���d��@}gxp,�uױc	 ���9Ţ�R�{�����kku�۩�B�ng^ɳ'�*%� -�U=�@bh�U[�yQg����uV|�iY[z�eC�H�T�����~�!�z�W���������ĭ�c]�r���\_{���-�΄V4|�L��l���' V;b.JI7�Q��� ������9ah@�'��$��/���]��u�FM4�p�Q���D���Au�:h)"LVR�Cɱ��C����`�vp�"�v��@�Ӕ,��Ր!��)���F��&]�k���q�oڏM��`P��OlJ�e�ӑ�H�]��;���Is�~��3R����A���:�W]����Eq#i ��R�d��c����e$P֏��5MS
��h^c��J��X��g?b������\<�j��=5�E$�p0��^�ߣ��a�Ø������ ��+�~�5P�i@�i|��5x���7&�d1����
�S��H ~�k�M���Y!�(E%y�7N�Q�Y_>YxV� �Ԛk��Vh�D��wWD{9&�yjg�F)J���k$g^8�(7��V�'~gX<<(r��rS�Lݑ�F������Gp�c��,�����I�C���0����"��h�Ubu�ֵ�Փ/� �%�[�.^�E;��3����f%����9�k���m<f|Oo@�zw_�`�4ك7�3��0N4O�ז�S��[5k��Ek�\�{�N��Ǧ��?}��?�v�l�LgR5VF��^ȴ�&�*^)FU]��͉�I��b��۸��̄��/U+����a�41� ��/eU�"���N&���(�n��O�yΒo,� ׮J�TΠ�M3��ϔ[ t�|���Ǽ�oQ:W3[���[%9J.�}(G�����LS"���8��1�F�^��%����(����IX���~S���[��a�����Z�&����C����Q��F�x��d;~�g������15פ<�K� �rt��@�*�y���c�p����3M�4���'4�d�z��C�����`?͖g��M��޲H�]��鋝aZ݊b4���_j����ZwG�O��8�o��(��;��|�,ź{�$��4��搊Bn$���}��6��K�%���6ɀ��~>N���z+���@_�f�J����vri��l��W��D.�?JW���h<,զ�~��}ƴӟ<-�����]���d��omvU�<zhW�����n���.�}�M(��CR�ۘ����~�)��|>���r���|J8ֵ6:���Tj<е)
�{\�{���dS:�*]���I���C��hL��,�k�T�YT���`�7��L��/�E\�<7����WA����'s�E�"���!��Qj�A�'��H<�&��
e��]�����a�c5`/��)��v��<�cAh��=�Ԩ��=�Q^��uʞ�dy,�v����4$?9�}�����g�	<����k�(x囤�B������>J����+�\�vhY�4fػ�lͭ��G2XU*���D&J��a�4c�^�`��{:3ɿ��S�o#�S�shV������+G�2��SM��8 {��ˀ�Z'x�[A.�-��,��]�~�8^��V��4��+��}��|A������\e`�luY~�CĬVͣ��,����ת�����'���fSy����t+0c����M�6�!��I�'+����ف4kyI� �,ѱ�K�k��@O
�U��~�5����q�mӀ+�a�����"��`�z[��w���c��?�2�����ى����O��4p.P��N��
R�4b2�33r:߿6�@c�O�ԧ��"מsKa�����bg��ǋpS�T9p9ہ�jIXE�@�T��� b\�������ޢ(�㔋`�y<5��)p�ѝ�>V�8�Dw��c�ݗ��f��HTaC?�h͑��9L�6����Dx�k�r�{M��-g��&�ŭK��7Y*$N�]Fl�㐻Ed�|�#�4{`�_o�L�b����a?�����m����:R�2"�C������֍��+��h,6�;?g�P��:Q�st�D��֯�o�u��w'v.ЇX*G�R������~܋у�N�'�|t�m~{懑��R.3������'U�N4r42(z!Y;�9�,*��n')����"S���}a8��Ҿ���>&t.q�ϳ�;0V�=�&N>*�jJ=��܀�˔���	���H���`��w��_q������5F:��e���"Xې̈́K���I�Դ��fTM�k�hM�_>�wgYu�Ҍ���}����y�����y���1a�02$�i\$w�N�S��sxF�8Y�m"�&Q�6�2w�N�m~�^��v ������Q8���:�t��
�[�D w<������Y(���V�3=�`n��`�dn.������AZn���,J�k�1�Z���1.-��&���)h���f��a�W�-XlG}�ϟ�J냆��������%����<���� �O����x2�B$�7�P�7�)�t�k����|$���7~���	@[R�U���~���cO��jl����-�IA\ɋ#MdG�]���^+�~�O��}4�xg���-�`!��@���حq�Ͻ2$��w:��6�G��uq����=z��JVcQ���xnb�U BC�O�����c�lGIAgp�p�DXa)�$c �
]H ��O"/���5��2E
] ����,7����|wj��S�Z�-�Ԧ*�&q����+�S�����E�d��.�wU�[ꆦκb��*�O�ؘ����d���5�7����d��'@є�4Z}fE_��K����C����S��n��L�W�F��Jk힐0���}rS��ج�8�38�&Y�ɡĲm�gsa�{#��9N }.�<�y�lf����W�gL�A��eÍ�b��P�Y�!�_��ܤ�t��&�Z���x�N�&
�����0��,�uD8�T�o�����Z�O�|R�~h���� �6RY�_v�JC�Qi��%��-cVY� �B��������jC�P�sqY�Xʇm�35�%�h}�ʾ�a8　�{n�1@,����/h��+�rކ.Y�$y��u�~��(f���by�%.v+����4�9�
��?����u�w:z��.�� "�����j���n!"�����}X�3O��DJY�gJ�~���,��b�w��Y�pB���W�$���Vl�sH&41���C�"_8��A��f�G1�4�`�K 锪@zn�*���/��%a���W�q�!���c����j�p;��p���%�'x�%�1K!>��i�]�� �)��J����16$�����ًiLM]��.��9$��5���������~c�JW��d�'W
*�w��[����}�w{���#9��n� ���kXE�b�on��� Z�p�9RH���� �j��s�R��#��bE�{�TQ��Ʒ�T�+0��#T��	Xҏw�@���m���)�y��i�&"W-�>�/�e�OW���1����vx�.H�r���s3���H1�?$�@Cad2Y`��һ>[5�����R!ˣ����j����dC��Ȼe��бgڈHBPMi������E��r9�/��p�?�SԵ��>~���q(%;�O�iI?�4D{��^��+���Ed���ȞH�t@�.��!�~E�Q+% .�j�_>�r�۸i��y�/. ������Y� |"���'eЗpW�L�5����y����b�)8��g��\V�Hhi�����zl���aMW���ggb۳�V~�-ee�v���(%��.ү�_Uz�6d�G3V��6�q;�+W�ȿ��w�@6�ŕ?2O���;���&yā�~�BX6<�Ύ�=������赊y�-^�1(#)b�cO� ��u27ĩ/�
Ŋ�b��$hXg�e��֨�m��L��5G�+߾f�5�fsIx��y{D���8)��%/֦$釾�F�NB���t����
gi�Ș�9yN$�>����� y^a�̰'�߼Y�����3m�f��ړ>�����)U��4�7�:�/�`g��Ƿ�V�@����tn�_�BO�W���[ݰ_X��+�A���^���(%y�$<�FX���7�7BHD=<7_��*Emß�0�}]��e�(�=�:�x��-�?׾���$�pj\z^�t����5<���%[. ��H�hT��t��Kt|��h�')��E�K�6����[�_��|�Sߎ�HNv�P�$W��d��'��}�Zթ7��u'�	��`�K3W����+���~.���F􉻿�q���Lȧ�C������ix����OX�f�U�� ��kK�*��y|8I`���������~D)�o	Y%v�l~�\��*J�i���P�cY����f"��˛!Ԅ�Q�{�{k��Z�/�a�������9�� �V�p��<-���c�AD��p4<�2hD?��o��X��5����-`�q�i(+T~LCo�<�J;��6���k�jY�/��8*D�Y�bG��= �#�_�E���qڋ�0ÈӺ�o�݄�|��˯Ys2F�4�:����`V~B�j&�S��h��9����z7�N��b�k{�U���������*6I��LǭL��S^?�44��)9?D� �!2��C�w�APJ�I��Z��5�(��c���Da��ʽ�Q^a��+�uL�?u �L��n��J�!;)� ��=�T\4A������#�;��y�v2��XlF����X*�~�X��~u��Sǣ?�8�F�[���@P�5���Y*�"�ÿidj�JI[��p����V����ƽ��]�]o�:����7���mAׯ��M��C���p����Y�؉A��X����$��s)d�vO٦<h���Y������pP'�Ё�5�7�nk��ݳD��������K�*�UZ��L�,����:2}���-�Jѯ�s ��B* �$>�Z����:����eC)���򬷮-�6ֳ��r���.͏���Q �8D�,�N��x;�r�b�@���Q`�P�0����*������������u��ւeA��f��qiD̚e0<�O� M�Dg�	ԋ�u���-E���q#4���$�d���Pv5�����Ï�o��8�A�X��?��<~��v��Uk43X�\6*͎T��n����C>u qh�mf�~�8 N4�'טz=��D�)R�V;+X" 'E9�$��Mڱ�r+�AR4~��:bJ�j^����i(G)$����-�jT����޹�o�����7S��=�9� ��;@1Z}A�y�K�o��_NLc��Tk?���F�`�
3�O���e��Αd� �u�<00w\h7-�0g�����i��U:�IMT�-����� i�n�1���4$��}s��b��)-Kf
�}5,�kg*�a� O��-�*^	!���� ��N�= l��,SH�BdU�����P���d�Ќ{A����	K4�#�_5����@3K�m��@��nl�`��N�ϴ��мLj��Z����츃~'΁{[��z�Gݖ֖1��F6y�O�1�M{���:j�hD�Eqɦ�S����`<2s{��]×���g�q I�9�R�A#���2��M9�l�fNL�u~z"4k�[�E���4)tX��I"��<�o��8�]>��Q7�Hb�l�K=�ǚ�$��#�7E}���<�= ��f�� M߲y;/�
	���fɾFy���c� ]��&�̃��Q6��O_4�e*��J�pr���	�S���B�d�o����+�����i��7��QbD{�\˵K��Zl?����j���n3]2L=���܋K����3���ݠ��n�k�y<��v��`\�P �4R����\�����7:����|�(���%T# $��f�����?���E������ ��"�I����3�񡁡��v�@�	��[�����:lg؏��������>٢�r�Z��z��il3��
e��J�����^�%kw�D�_�-Y`��޽�U!�� e�1���`tE
���Ρ&��egbw�[��.��Ai�i��u�����^;�@g�]����6���L�(�{O
=�N�c���Ez���R�|L./N��q����I	x)���$"�_H��=�a��m^4���~bAy����Hʏ-� �Ne�]��n5dj�r�zέ��ރ��+�)?u昦� s��ڀ볓�9�Tt��!T]Sv^!��<�	���Y��>d`��O�=���}3���:pܲe\I*��<�#�Po�w�T�Z�%��
�D�#���|߮���Is���l_���mӕ���On�O��������ѽ@�9��eIlmP)�}�jG��j�@U��:{�X�u�&�<�M/��ߝ��t�\l�蜐[,VNKsrM���B(�^��{���!�ةa�"�ФflۏP�4s.L�L�y�T�`�8��8�9j���KO?�KVz,p�z��!w����Ԕ S{�Ty���)H�ouIqF7dI��
��-|��Q��X�M+�N���5�egt�΍Df۞���/;�Cp,�g5?!��NZ�D5cY�g��	i3�B	�?iLQ)�!�9��Il��8#�O���[��
���~�y��㘭4Ybd�UɅ�ZaJՔ*]�&��f�6c?bX��#Z��~�\���C�1����Ö`�}���">Jd�C��J�2�U�?�ҡ_)M ���cŗ`
〸`�Z�b�p�8u�Z�^���p��3���u^r҉W��_2�x�\��HD->C@�����;�����R�.�eVA;+()��:�g�/�VZwq��{��Ą`�~eh��'���b�/�p��P"���D��s0<4ʹ�=�UY�xw�N_���6�RV�K���eN��1D\�uG ����~�}A �k�4nj� ��>վv�
E'����I�豭�m:�5����7>V�o\���:�o�9���?T�Uj��7�*�,�6���!�F`|�d��\{/�n¦��� � =���(*d���Hl&�Ő�P=4��h��3���5Pq�%j,�����(p

�kzV9�-<�ruè��J8�!���"����F �����[={�Sy�]ω��f�/z�qӖq�,�-�i�ƫ ���N��j&�L��x}EE������ jȋ,�/r�?K�����b���7Fj�,�y�'��5ZZ�	�m@��W���x�*��.���}���=jZ�m�fF��>eI�����E���s�+�5�}��?Q��~ AI�j�i�K��{�+�T��F�� �P%��0��(T F�
=Í�ԆZ87���M�hy�Y3�̭&e�����u�T�M@_���76����
z�x�C��t-j�5��v̏^�Ґ���'�[\ҳJa�PA�qUQ���Or��f��Tft���=�jj�Ԉ�qJ�B�g(`tQ=iR,Jٟ�rI�l9q���Pl��=�$��S�B��EXSnZ�zD���U�ɯa�hFZb^!�I�-��d��Y�6!af8IƖM�D��w��ت��3LYj=^B�k���t'����b�k�;x/AĤm��yK��>��?�"� {��x~�W��=�.��7� ���:�`��4�0Γ�_j��G�b���gL�vǽ��G�+��B�v78���[k������տ�q��v�≟�]ȵ�a��FGtkC��-UJ�*DPW`��n���h$A�C���(��c�<���[Rr[��M8���OJ�jl,0�
W(LW�8u �k0=���|�n!*�S,9Br!V�����N���;޸Ú'<`�$˛��þ���37���8������p�7 �
pI+@�����o
g\��מ�F[�UK���w�XXߐ!�[̽���*���5ud��`�~U&�4���cR-א�+�%��Z�o��~D��bǎh�3&�!�=	��� ��l,��Ư�P�\a�0�V����{8�e�Pȹ}f*��
�K["�@i̟j:\�9��q�[L�i������l��8z��!i�w����O,r;"[�X��B�ρZ,�	Ż�&�R�JC	�)+L��/�1vE'-D�HʏM�k`B�}w�<�O
9+b�4��c����@���:���̗�_�1����	ݟn����p[����f��~r�A��-�fTn����Ms�*{�X�17=��%^�#�.=`�jP���Kr���3NC����h�y*m�S:�n�v{�/�h�А1��ky�vx,`}>�nH$S�U�r�"��-v*s\�ëY�7fÄ��#	�,a`��$������C��
,����<��g#��]���H���-tP4aɹ�ı�a�&>@ʉh��V��
K�� ��O�d�����(C�R8�ޣ6���Zu�S+;���kvY��~����-z�N��
��5�Y��?�_���N]%C�w�d�j����4�뵌Xy{��pc�Ϻ��U��\oN�BG�+��jm\�z��tx��Ii����V�C�ʝSICp��jp��~��2k�G�<Idi�����A�{e�=�(*�X�Q6�T}�1����>�R�pa	Wh�sj�1K�#$��}��-�F�wʧ$���(-��όӈ��/?�F4�=�fC��>��=f��9kU��ʧ�زo�s/ނ��諚c$Ĉ~m�*��p��]P���+���Qm�J�'FX�?b����:ɡ�eo�e��*����|�9�b�N�v]'|-W����VI�����������Q���=��@ĎX�����G9L��#�z3�qǉ��������~P����GAH[�-��Ny@f���6"���F�l�z�IR�p���qM�?�0��.�HU�T�,X�i@z�tȅ�.��Ji^Q懲
_�����c/W] �H��>�`@=	:-h>�4�'����)�(K������"�GG��\}���z���R-��ѼgO��G��G/{Ȗiȳ
�}����*_	RĹ��b��j��7y�9%�o*�plw��@����*���:��6�	��e�Zɜ��9�����3|����Ǣ��/��q-�o���#^k��#� z���k&���m�����"�*�;�HN6f��d#��q[\_N�t9(�0%ڍ������隻[	���7ٶ7���2*h���G-B�'�����U��r>G���гφ$��*��x��z!�'��� �;�Gf�a�L�e�SZCk�ψ*�*k��xS�Uݕ�B�s���a��W2��(�Y��>"7�� 踫��O8�&
����5�]h�{�[�ίwA2�s����^����F隩9�$�_�k!i�@�WU=��L2����௟ы�Ɨi0�C���"����HKF��t�גv7S3�pڤ7y~!D��ꯈ$�����㑉E�� ��N�G ��_[ֳo	�uS���fs�UApz��:
�`m�_�$a\�4�������咙&���+P�k�}�)��m��	���m��6�UT��}8��*�`}Ѹ':�4g�T=?e����s��h����_�,Q���8Q>�->s_�R�[|;ZU�W�.��W�D&��?&�_�<�3��I�a��k`!C�)J��eN�"1����=Q��wY���e�*�jA��::+9��#�-�cI�UՖ��޾8u���H�)ۅ�Ϗ���5�
l.�Q�)��y��Q{�*�p;\����A<�!b�S��-��Yv�=�I?��c�^|�O@\���f�lO���h�X`|&�&��1H�Y�(�������ٸ��J=�#�e�~�ǆ̿���}�J���,O;:�xL{��:qC�H�����%���O���t�xC9�ʉL�AH�F�8�Лyj�n�����'.�d~^F��:��L�'�!WD��S�4��� �WuP�Wڭ9��+��#]���'?6'#d�=1x��njb���A�1 W���{��)�cAƾ]M�\/�tpC���>�C!����- \��C��E�����R��."�:���ߓ�rG�T~�KI�4�5�!yD�-#
mz�z��R:Ѭ�"c8��&�+����"P@�ej��=OƊe�c�O�o���#�$H�[�.�M�N���d��-FBg$���`q�m��-���<c���}����GmZa��a�5Fu���#*,�&$"�7���!Ā�����[�j��{�Ó���5�����x<�+8�nwT�u����y�/�"v���
�.�Vi��z>���	�l�3r�$�yRE���z�0[�k���T.s�Ф���:d݁�xit��Yi���n���E���J����V=&k���*��S��E|B�� �Um�g��@� �Z%4���"��^'/�VnF���I	�&p�۶��[��ݧh��xX�o�AH��%B�ʡ�Ğ@bⲅM��2��y��p�#^��+�8E�H�'oV�Ϲ���L��ԗȑ�U�N'�@L��N���L���`e;���bL���k�5�	D$�ɻ�])O����BM�m"��9u����=�~�?��-��r4�盗��#�r�T���1ϱa���V��p��RѨ9G��3eZ,����*�rw�Y����p7��Dޞ��x[(�Mў�vaeJyHr4�c��4�.^^gw���l�(o9����E�Yz
���ݳK�DO�R�\�H�����x�f_QF�������M�
�1?��I�A�?y1�_�L��'�3�W]NTç����C��yq�x�ܥ�If�'��|�2�(;�@�θ��Cz{�� ��g�a�c�9�2�� ��nժ�����U��'aF��L]!���V��S�T��8��c�s7�	mcǁF"�(?*N��4N��'���2������H��]2�`�YKȫ3�m�
�E|V��]�e�%���s���9y�����گ{I��<yG~4�kMm�2_�l�r)j�`����ޣ��,}Yz����~MJ�R��w3�����a�(�j�.�z��lY��$}��0���sdX���0S=R8��q�}��*���10&���B��,]s���6&��%�[p���w��n���ԨNex��B�$���N�Gs#*6���q=�{�W�w��P+>�	�pA+�$?������Bh�
f��N��y�.u e������30�n&ջVPKB%m|�����j�sUk[}]@e�h<����?���
�C�3[{��n�C�WX:_�/S����F��{��;�So]� e�+�\�V�&�X��G�2��7!��U"8��cP��8�U ��
]���=^����is�~��a٣�-�L�5���d�T��6��r�>,ŧ���� ���J�k�$�{磊�I&��.׫ft��F����ȫc	/���jM����N�tr���P/m�gL+_���ָ����fM��ZDMn�淟6�o'�����ʔ�f��19x��}G���++�q�E�Z䰜Wjв��6���
*,M,���`?�Y=��ⵢq�_{�I>ZDG|MP�zJ{Hjhۄ�j3�����Y�j�^E��'w�wf8s�E���+������zJ�
���|4��I�kB6��jz�.�C/�{��(�B��G���A�a""�������*�s� ��:h�|�n�^�\nm{��R~Y*�~%��B�:u�ؒ�q~�Aڳ4��7��O��rV]�| %M��;���3�4r��;�H� :y��A�����ym������Y>�Y�/9��a�<�3�9�M(�U��P�Jw��&w���o�r�*QtR���*�����2��9�(�z��@�{|�R�}�w` 
�F��������B����Q��U�70�ϾH^�A��U��"����P���p���h+����l'E�����듡%�Ȝ3��Dh^%����%x��ő
Wz�f(Zo���x��|glVt�1}!C����+R��1�#�<d����_�۽�q$���Fխ|���^���OH�JC�/
�8�R�Ԥ�.ƅ֊k���^#�ul�/���ݍ��`��%�X�ϡK45l�\2X��Le�/l�n�/�*P�8��1U��(_}Co�X�F�S��@nw3��Ep=9ؐ��6e��<�+zQ�c����򛖘mtx��.��>p8�k�Qx3��u���iIv9pz��Cp'�=0}ǆ��$����v�$�*��M�t�W�}�r�h�ՠ�Lq
�8�7)�W&��:a)M���wl��@o'l��ɖ�F3�_:+���x�P�0d�&����Ͳ	�����Sɥ,]�Y5���/c��21�̠�Ђ�E�%ɪe��T�D7(��%u4{]ؠ�f�����mr��F���i�=��G<>څ��L��F���[�������ҞQJ��%�t����b]�0a��Q)���[�%9I�~0*���{
H�Υr�8��JMC1m�\��	��J�5��q��5��M��s�d���o�B�~�΁f�-n��<�زB"�$SoA�������T��1���U������z�Z��S�����aG�{i~}�2]qz�� Z����	��8�b����A�]<�~5A#�"�v�k�$���ɴ�^�j���m��߰ݖ��|y��J��8��ℹ
P�&�c���2�y�lAJ.Y�5��nrP�jS��|��9�$�f���&⑲�S�q�iHp��̰����8�̨����U.e�����X�Z�P/�7�.6�:ulA����s	�ʄ,E&.x�g
.�.�>l�����������t�1��->,N7��!�v�<0}١�C�� b��X?/��4,E�mk(���ƴ6�9�����l۝(f	oN�st��|��[GP�^hם_II2|<͡����N�w$��@tj�E;���ӡ:�zA�G��I-!��8�	~b��-���l��?�T�q_��LǍq��i ��~܅�`�"n.��D��b�5	��cf+������mZ]� cP����x-�I7笇�~8��d8�f�	r>�c�#��-@S��ܒ��T��jޭ����JJe�|r7�!{
1�p���wϴ�9j8�uQa�q�]GV7�]L"�R���y�5K,���ҩ�ʤ��N)��|��G�r�[�$1�Dz6�2v�ˏ�UQ#�q����=e�E�L9����8ZC�1n�H� �ZTa�ݦ�$���
j�/��
J	ԛa	��K�9��z&�$K�ʦlQ�<�v��IP�*O[�]�r<)��W�iw<�9˓�Y]��gjE&K��� �{:h�%q����?]�c�ksŭ��E}�]r^J�!�߳t.�jܶCJ�k���m�<EI�T];���'8����F�F��&*�3N��]�����	�2`G��j�Z��4u*3�eH�0��`)J��^ ���9z�_j@l��4̽Q�c�\�� ��������rް�4A�n=��6=����G�	d�*��L�eC*<o%/�ˑXzv;�԰��Y��:�q����Ȱ��<C�:�~9�v�y0��x��9��,_Fh�t���	���bJ�/��5��RC��AN&/�A�df3..g�� 2B���H9�hc"�+��W��/��8����Uc2+��Mc���KOU���Ԙm���3�YG����
C��l� (�ً��.�o W�ೢ�_Gi (x���:>u�:W��+V��C�Yʔ1�c>��Ϛ��
�H�9Ke+�oh����4��6�܂/���[����[��An��:O�z�M�P|$����/dG�u�<�^qA�TZ���	����#Nϙʇ��>������]D��B�M^�6���}P��+�a�P/w^t�}��8�tŶ����ӢZf�#{	�i����ˊ	��˦x����dG�P��Ͷ(��s�s�Ok'D1E��i��	}�"�7v�?��}���Z�������̟9J����@E���N��Hi���0�?�W<�5%��U=��'|p$.k��ٯ���Ռ ��?^����;���}���-B�w_w�R;�\�x����--�g7���,G�H����we_��[�jہ)6u���T#�lf���Ȣ.9����  |]Ɏ��Y3t��Ҷ@eZ)d`$�*�id��	u�{f���j����������F�7i(Fn���N���{%�ʒZ�DѲf��
�T$���#����N���Dy���я���"�j�`fI�U%9]�<A����Kg�H�Ĥ�.�\����8C>�i=�i]����4�#Z���]B1�F��M�C�I���F�Vf��r�k�d�O�[ ½��7���}� s�N�)��O�i�a�ҡ�w13f":���i����4I�x������jG����*�?�di�;��e����8ۦ% P�������
�o��Z��Z�?|��hv�y��2eb�{&�O4����|`<� s�µ0�\N�p�t���}��>�E�o1v&�[w����E̤���#��dhl�lm�j ����Zr��d�5�.֦�>9�;xZ�t�I!{.P�;��Q���!��.����.�s'�v����=��ሔ�qQ�������q�L�<�N�=ʴ���(.�<�וQ[!\ڃ<�F��Y/i)n��Onu��4H����.6�;���� 1G�!y*�+��>�T�Zz�Զy�����~1�<� �չu���c�bo7�M�(��%ܧ��f�w�%�>��H��,s�k��%&�2�A� K��zߐt��r�������ɉ��F��R�d�lT�cR�D9�h	݅�R3e<8s�˞;
%c�ߪ���+@+bƊ�z C���	[��;T3`MeZ��g����8ۧQ��#�-@����(���&aȴ��ʾ�t�����g����ޘ���L֓A\�~⩻ü`D�w�&�\���9�M���o���6�i>��L�L!7*=�JU�0�l�B�I6b�j(G{"$� �!��޴J�|5A�ꕞ�� ��<�eK8� �y*���&ێ�J��5����ӔhH/�$��*o��k�2�ץ
���i���B8�����D�:�5�x�H�J:a�-�>K��ŗ�m~�wo�.���S�nƖ*ACI�Rؙ���d��,%��Ro�����es�����"����%��4T�^`������9����c�\���1[`e2���RVq�Y����/�z"M�ttP,��Ԕ��:q��pѦ�3�k��6��$�DE	2/;�ڼ ���ԗ��ν���Q��	���6^�F��y�K���[��U.����B�*�#O�j}���t���S\������"�:��W7��@=��g��5K-t8#��9�}�>���S|����|X�QN�����B+c�0䞲8r�h&\Y ��Hà�AH�7�f��Y<�r7��2����4k=����1��4Am9;+�����F�v�x8=fuVM�߹�%�輅���9�a<�4!}:�lR( ���Ny����0h�'�����'2Ý$F#߫[��[.e��f1��F�QI�hX��on�^h�/�F^���C��2I�;ߣ�;�;�xl1�7!j�Ϲ%��{������Gs�����z�J"uv\�VPn�s��<�P�~(j��숭�����dsfGe�h��'�G�=����^^����&���Q���g9�$�!5�\��h�qI�P+�7�ڂ�D8�7o}:r�7��!Y���Kd8f��~�*(B��jf�̋�*��k\�$։��_��r�ʐ�4��v(�Gr�b�<��� ��
\I�Úb����W�F:�Y���ι�h�t���, �r��V2dY�ѐ(�e�`��W`�s�Th���0/�4,+���2ȝ��5í��d��L;��g.�����W j�)����C���J%��dX::�`}iO�w{\0�Į�2��ɪ���~I�@*�k���	|<�5�3Qcޝ7��gc��|�f�ƨr\ML����K � ^�-�����d�I��=�4R2TK6;�I�i��L����L��� PU�GXT�h1���l���F���3������(8��\MT��~4���(B����k��p�qO^ÿ�ߍh���n|R��qǈ��&O@�Kxy�����y@�S���BeC�yF	w��>uƏ�\�����C�g%s	t,�[�Qd��%i#�\��L1���(:�97�$��4/{'��IZ���em$����kGͼ�>~��C�C�G�*��(���1:�P�W�G��P�e�O�ڍ�t����L߷���s�xm:�i`g�${X'"9�(���F\�5��
OZ�V�_r������{�]t��r���U_��,<|)S�iy�Fsp����?ĝ[\A���I3c�4���&.�JO�i����!�y`����'n�6�R<^�.s@t����_J:��#����lEj4���W�v2�������y��s.b�N�T<�\�IR�iง*C��h��ւj����A���dz�f�pl�Ώw )�7&����M�O� uXZ�D7x�vX�`(��d���x���"sѭ�/�-�u�6'����	9��y9�_ѭ�C���W������T�kf*F��)ɖ��?�i%+ɒ�g,�(�.g�O�;��R��M/ݸs�%����i�[1+K�{�f��Q���4��9Qݶ�TX@^�{c|o�8E��NY4�;.���S����[�d����$�G�E��D�-P�j�]$�6+��~}!�\���b�a�b!.��Le�7�pz�� |��r��Tsb�!r�2縟��T�qC������
o�O�z`���6JM�P0Z�����w��y
$��-,��g�Q��`)�4T�&*�q�-}X���4�I�T��x&$,��N`�J�bX˻�
�*]��-���,��+��U�⢍�$��N��<����p�+_��'�T�F�"?���kZ���~œ��V"֑$�_>��O�	C�5�z�G�b���43*��hWS��LǏ2A����4-���6����!x$tA��UU1eA��Y����b�C�] �V�6�H^Ge��w�1w�ĿO��u�w1x?�H��H%�t6h�g�Z�s�ig+91�����~3�FVs����a/3 ��h�ی:g%��&�6=�24g�|�z�� �@�{���^ř�����d\�/���a��/-���*�.�XW�]2��v~V��"�Lrp5D:?,��@r`���n�R
��k}�W��]��X��ϟ��m�7P��P��[ur�jD���J�	ι��QJ[���6co���������c�g�/՛�x��8�K5~�)3������=5X�NK�E%�ʷ����=�[�{��e��(�ɀ��j�S�A�W��G��Q�w�(�	��M�;��MYBh�k	 ����r��H�ܦ�;��T�ި�A͘E�Q����[��7�Z�i[b����!I!�·�w����ɇ5��j-�������>���J1�J�/C���>�i2Q��˨<��r�������Rqּd	�V����`n$D�hP��hDm��FYfc\�4٢�*E[I8��,p���u���s'e����mQT�ҁ�������]QjR�g_�0*�:i�f���dM6�+����A$oŒ
A��kx����ZC��y4�*��x��[Lb/,S�����S���e�b�i��h��I��k'4�C���ut����!�	�p�ޟ�H���W�g� yZ0���3�p�;����Ĕ�Z����s���K����b�a����nyQQe���4��d}\�-q�7en�TT^9 AN0*�3/�h��4Y�M�T��I#�.H�i%YÅ��7�glV:��lо�Ad���)�G��FC����x��B�Kl?�g��Y���m4L?j
�e�h2�`0o�p�)�����b�Я�!�
�E�!�b��/�U�9��:{��UY^ ;�5���Kwu���$�6��e�z@iP�a���C� �X���t��4<��\~]�w�abh3��.4q��bH�抴�2jik�XC��{����]���V�]��M{Y�X���8�fcq8+:_t�hy9LOt�F��ۥ����-����{7����(�"�[-p`qn'��[�b�:�1�8�}!H��	��g!ӉQY�/�}L{��w1��c�e�8E��e��z��&5���}��"z1p��g�3�9�m�/&��e���\�h��im��Q�jM5-)*�zޓ��%��>F@c~�B!<DjW�0���=�s���;��=��g�_�+���^�;Ls��_�7�9D������W��E��(��2'���b砾��[fE�L�h�e��$՘�,I��(��|�� ���p�������H��a��c Ǆ�y��h�(]�dF��O�22&|��äH3<�����`̑�L�1K���~ך����_�������CC�F� �bUԹ��X,��P1�ű�e��y����z)�`�ȦS�M�L��j���t�~z�Sd�������<��a?Ғw3�����X_[[��`���Ӈwl6t�e�$���߭�r�-��F����|L���B㷝p4�2�d����f[\Bkc[�d��/6�H@�	C-p���u���&#�Ut��1R�m�6�+S��J�a�л#s���l�,�e%lt"�G���
L�����1>+�~�6�2ϐ� �\�W!?c�]�.��2l��\c�.5G������_�\���R�ƁOe���a������K��/2����8����Ŷpz�+�w����q�rud�R/�ю�}P�����w��f�V"�,�(X!��{?�`af6���AH�c��W�P�A�v?QU�����YB����iNgc]6g���6���{%mx�!e�8��խUJٟ���!���K�U�$��ϩ��t��*c	�A�&�`G1,b�:�-�p�L�Ȕk���`�p(��Q�"��]ކz@�<c�GA[l�B������.�8e�?�d��N����̶k���=��}�A����,A�t\vC_���F��ؑR���&�<s6x����,��Jf�#�������,Ú��y��SN���0�G�s�Jx&����S�)�b�����Q���55��Vn!�uĨU����tް��1,�i���U �,�:�R�d\A��q�!4�=��O���uF�Y���Al�L�N�Zn��8�e��Q��bB�9�lēe:M}�H�|�@�PH�̘QE�5��������R�me�l��+>�����[�����e0p�/����2��|���cߨr)-�i>O�R��<-�9�����:����f�1��双�=�Oea�a%�\C!eb��K C3�_+������jl��]E��¿�v��5wAH��3�� O~�˚��]�I��Ъ���o���C,Cm��\��N���\&�b��[@N��~�+d��ya9J�l��[���K/�yA�HzQo/r���B�'�o�Q���2�B8<KƂ�'H��X���-v��XD�N����Qr�8�Kng��r�n��9��2�K��)�mG��tQt��A�8^�)h�k��(�z/��_�U�Vg�:��U.����s/�8078�v�Gt5k�]$ �0�����+���Y"�W���� >7�5�d��k&��	�8�>$�ôE@��-j�R)����,������{1!o��ߤ����"�xQ��z���u�T�Dk�7�����56"{�}�Q��'X�^� �A7;�Mџ4,�����̡��T.n��k�8�R\>G�/L��
����,�j�k�vI�G�j�~d��o�j1C�F�� ���&�rs
��R�vKJ�����N��:T������)8i����Av*{��7���/V�\���Btq0�F=�9J�4� �5p�∤�댡)���Q�Z�f��2��VZ���3��+�p�R������F�b�a��	~]�=� <_
�=�o%EO������%�,}���oI��<K�J�/��ȋ�����3���CP��V"���-wJ6܂ٻ0��5�?�K��	5Y��>y��]�v�D�@F7�Շ�x�ݍ�3�:�M?a|���@��+2dǉ~Gsܞb���Zp�j<" <=�|��A�'�%Y�b3诐��v���r�ia�RޟB��ۗ��d�-���˨:���Ow�PNg#�VY��^"�-rN:>��  �m*�pk�d��v- �`D��G��b=�5~p����%'��/��m���ҽ��9R�M�M�������jQ�Al]f�R���u�C/�$ʮ�׾W�UdUN�`�������n�ݍ�n�L� ����"L�]d��u�j�G�'���#!��d�<�����Q�T����2_��<�*����][K�L3G�;}�T4��|��ykE�Y%r��R��F	Qu�Z2���$M�S��M��dK������{��c!Eg�F�zo5��M��JoồSn���z�b!:�͒b���]J���5U����� �;��͡`� ry�k]V���r��
�\=D�P%,Wԣ��m�6������ul!�-�@@揣a�ݡEdْ��td�v]���lDZ�ƨ��^����f�ŕh��ef�{���Q����5A}L9�Y�b�� �Y,�hzfYK�ݳrEMp��Lr�7r1��.�]� ��4�+9��p�-H;_��~�)d�8{��4?��/=zj���Ĥ0���A��?#E�'8��}����0��FL�>t;s��\���c� ڷ�]�'��}��v���%f���8P`�m����Z9=�����sP#���r�&�m3s�_l��}�eZ�k�k�U���$��������p�k�w��5�~T�D/��k:rմk�`��G��2���xiIȔ�
���e�>	g/:H8��\�+���!g{�z�֌��[Z��ڟiD���*�.;�ÿ�����l���A�>�!l�j��@p����yY��X�|ҙ2�*ݨ��{�|�Q<�Ϟe�^Z�r�\��|���a>��Z�Ў��zM5,
�fE��"d��6���%�1Sy5�^+�Y��C?��&9�����.ļUM+y��s�\��o�2��t����2[g 䇶�8i�)��H:�5%�\���� R歩���Gt�g�ِ���#d�u8渵��W��B�[��˃;΢8�/��"$�es����e���t%e+����8��n��)����[�cH⽮ءY$}���͌�����SN�U�e�?P�oI���%�>e��.�/K��m-�Y��"
W�?%�?�"��D("m�'p̵Ω���A���h�����ә�׋�?V�+����p���Ջ�Ƭ����3��X�}�\������<�%��e)<���ژ�]���v��=��kx��nY;��j�S5���r���V�:Do.�5Ġ?����vV�=�S`<<^�0� r(,k��@��q��Hk� �@��r�V�A��n)Eh���Zh���$;�K������O
�Y~�� a尨?0���
z�Ok/4�N��&������P��$�gF-W^�cGT��Q������M���M2�rE!/]C�q ����d�*	�m �Kl �۷��ދ-*���b�"�Y$��
۾6�� FP0����<=�M��c^�z�u�
�dL`�z:�#q��С� ����X���t2w�y��3U7i��n#4>����ܕ������|�����TW��~����Zۭ)�|F�eިMZ�S�j�O>��ZO�c����J��EvJ2�\aҐ�r�HlRQ\o�0�W��a
���h�a���^�csL��,��zF@z��s`:�N5�n�К1�_�pC�ū�����+����`=��䃞D�̘��ьx�XX�-�&1j����ӻ�'��W��?,怒�K�j~��Z%�{H����\x��|>����No�����Z�����+��6�.a�"��)�<e46/ �Y��G�̈́�2�Es^P+A�ސ�VX J(EG\��ܱk�sO���%F�5�*Z�WߞֺX�QU}�*�<e$a�7��Y�(��F|U)��r�j�������Z��ă�Foy�m:��b�*�{L��Kf���Q�Ǥ�	ݣ�*j4?\�Bq�:B��S��Z��.�aҢ�_�ȿ��������e��>��>�by�/H�tHlpg�	�4����Q�p���h�j��r^y&��Z�:��Ԟee�#rǢL�~uw����Q��^� ��æ�ʺ���{������ �)L������	=�R��'-��Nd�ӹ�A�$���T�L�N�}�:�Z �#@x���e�Ǐ�+���1�k.7Ј�Uj�چM�������/��r��G�t��:8nvU��T��V!.�8�`��X�Α5��8�,Q
(�X5+f"��\���JWܜ�^p2`3�Ѳ��w���)Qٿ���s	���F���n|��P�X�`*2�=��*��Ԕ�[bt
E�;y�x�/qz�{~)R>���~E�
4������r�GK���s:v���6A�I��� �9�˅��S(C��t,�dk1�����c܅�jH�RԮ�,�>�س�8���:�2{��� d�E�=�e�/�o����?���������q�(�OQ2�ei��`�}n���v�pB�=_�mLp{aw��1S����k�cT2��
�^m���7�
"�?ZIl��ﴌ����{N�B+<=��C�e��#���Ft&��ڽ��ŀ5�M���^��Y2�H�8�[D���(U�F|EF��{�1�Cp��-��_M�o��M��e�Kda��REcş
�!D �,{vrש	����'iO
3�ċ��8�TJɸHD!�'�}R��R��˹\d��
җR�h�AE��7W��#��m�`:i��1so��rb�l�#3F�����ܰ"Y=X��Ncz�?�A��ʻ��~���L Gʢ�kB
���Q��S�/R��A���G�!M����Ԑq&�{%Q�X�iݣD��V6�Cn�=���o��ɼ�L���Q�����2:���)8LHČ�S!] C���CɩK�J}�,�X:1!3.#���\\F[��o\�W14H)�C�u��^�n|FII�gCD��4vkn>$�|K� +�E�uG�&b���i�Y�C$�E��Y���z��k���� _�<��w�YQC�,�XDO�L>�`���1ԇ](r ��j1@f�M{	־�Ma7��aɫZ��X��`��I����N�/���u$�&����c+O&1)2()��OR�N�͋�6Hf�4 $�&�I�c�}P��:SG�+��v'U���C��~*(�qv���%A�(�?��p��5�s�jؒ��C��%�X:=3;2�<�p�̨x��^4O��k���8�$l�=|��K�1�қ��2޼�;��	1/>��u��ŷϛ��&�v:�P��^�,�W52>�g��_�N�1#	y�A��Smv���u7���{A�w���W����\9����-TΒ�q|_���@D$��f���T�U�>n��*����?;Y�O��؉�� ޗq�Eq��'6!VU���]��� S�7����R�5�WY�풮
�;Fw� _V��~'�kFu���������r����W�:�/���hg�'�*��8M�>���������V18�:P4��	�g�.H=���ƌ1���� |�8B���!h��!?� d&�5|P��w���w_qp�;U�$O�I�M7��Á=��x4F�E�NYy�ҿ���R]$*!I���)�pG��z_p�����C!&[��Yݽ��7� ����>��]`*���怒�daAH�.(�N�Q��_���VwN#c�F�ײ��_�����&S���
����.���%�F�ڸz�!ؑ%ʃ�'���.e4��|;��X봿Y��H�
���ş������Eh{��v'�ܲo#�5*�;���0'gc�V��B�OEq��q������Y㣆���Ȝ��A�PJ���_�Q�+�p϶�6˲��>��J��8=h�;���#f�%��e���i�я>�#�F�EN�<�ٯ�h�-O#Q���:
�6U7�LhFWiUA�~�Yd���;���l*�����tKK6�Εd���C��¥U�/�t�[㿷s�'�d�Ӳ�*ƅ���F_�����k��A��Pt�ˎW�֑Ȇ5��{����.��1��"��ѻ�)�$�,B r��r'����R�ÑJ�#������~-�w�h�k�g��"=Cb���xYz)W�58��Z ���u��?6���ӆ�B�wE#�	�8cL����~�<K�Ct�,��h��H^�~2�7�^���L���O�g&0F�}��IndsW~|Z�c����o�s�v+��5�-vE.J32�,�Tf~��n�(���9b 1U���+��5\C����|W�Mk�c� ��{��j|�Z^L���7 ���(�˱�����ph!�m y�
�r�6������_�g+����|�o!�������o��� y�2�/�U�ы7!c+���M�Aa8>�dʗR*:a,�1K��l mK��LS�Q����;��V�%��6�$B+���l��n�	�Z��{�d��3��n�G&����2��c�f��4��U5����`��^�;*ʇ<�}�R��C${�t8�[|��k��bO������"(A������d�am��ձ	"L��хe�*����8!�TR%(��at�[Àٯ�P���b���Y�n�%IC��u�z��� 2=�[��QA�4΀M�+Q�
��Y�9��&�^!�*H+W��N7�D�5�4�)�2s��q�w��X1�_���� ���͓��K�)n(�|�6`q�N������y+�YZ��S��͍[�I�$�)jekh\�æ���ĭ�z�x܉t;f4�;�fJ�2��ҿ �� t�P$ΗB��	ߊ�?[��m�Ӑ�,z��I���EN�Բ��EVS��y��;s�>�+P���
s���uDz�����;��DKxD��-��=f]�v]�#��(����AUx�y�S*�S�gǶ��MK?�u���]�Z�N'+�6�ϬEwaYW��~��C��������zԬ�V@�.���w�,&���A�����<Ow�5�=�����Զ�.dz���ThX�B-����a��!��׫�����<�t};~#M��~�8f�� |_�<�T�����8hX>�^?�!�N����'J ���`b�b��0��������f�sWm���i�iEq�3�sz\E�e��b\fVXzqĒ�����~=�0j/Ѣ��9y�'�K������X·�)�WהrK���+�1.	��ٶ����K�El)*Fx/���x�>�*�D?�{����_��z��,A��*-�����e�i^�rUa�Lh��6�w�_R���f IS:�����S�C��n�(����8ES������}7�\���t��	���1ڲj���r���M�=��sZf���͢�I�~#@�h���_�#��I�����q\�SgP��ʖm閷e:X��ھ�p�>;��oQSӫ=�c�.�I�E���y�L���E����$t:��麚�ȸ-d�?Yu��	��͊���r*�6�4�r� zNU���S�3gl�N�ZX�O�41f)���dP��x9B+���u��\�uS�ܩ���d��������H���vyi��KO��2QU0���f��i�ET��)\�EQx arsB�M��0�^�d�#.e�_	r���
vb��f6���|�����l�6"���}��y�<s����|��ϼ
�2����˶Gڴa�ؽL�|J��ۈ�Z��
�|�ZF�ª�o!؈V4ԍ+���j(��O�.T��X��7�uQ��}�ѵ����p��,2�Sи;��w>�-���JF�I;��>3ほ�~R��
	�8�����&+�ZYn��_
����h�غ� ��Ԧ}�MA�N�ovOx�@�ب?�I@Q���K�'��	 ��v���b�z˘|ie�������(�x&Z����i�6�h1����M���'������?�U���a�Ou�!B�6sb#X� �h2�7�`V��p�B��,1�*�K��ר��j�X�5�~��K��x�Q�|��%�<���z��9x�<Q�v��^չ�>�/�^6�S���z�q:�[���"�^6�ߑ�s� �yw:�S��&��� �ˊ�E__���V	`*�9h!H�������J�������m���'b_Pq?�0�V���I�_��Ɩ����r|L��S�OvJ�>�!"����%Pb�oK���6R?�59�.�� r>�o�G��k�i���̶���"�_�9P�u��mOgF��ysEz�n�{���p�<�tG���y�-�oc�w�	&w`���ӥ�W�3�y:Q/]��m_��fP��<��yN?�)����jP�x���A֯0Jd�h�G�zAc�N��x54.�02y��������u�P`��"d�����ɸ���q���5ɹ��m���Ɯ	�����#S��ӱ���{��Q���rW]�S:����O$���=��e�s��B ��wl�"�P!����Q�iwN.KNu��^����D���}�H��E���y���hogtR��s�g�`���mp{�Wjo#��p�]�ȹubf�`�F��~��
a	\���������6Q�� �
�ah�OM��2�Ɲ�xg�&TO�in��^�L��C��6��b��.��Y�myk�ь�����ٸ�����豐���r?�hI�7���D��[���u�(Q`'�->X���t4��P0`��e߳epT�m
��p�����I3=��MM2P�CJ`��f�u�C��e��HQ3�T���8�ܠE�u��^jqj6����d�Р�8�S850�!Mw>��-¡�0��Z���u�-b�d�n�`�gA����*E���n��m��(�A�\�6|(h 0)����X��ֈ�� ���1 Y�wY;c6�tV�J��iujwÚ���5�
*<q��MZE�P�X'��բx�%�B4I� �1%�R�{��k�Yi!]ZkA~P�Ђ��w+�2�2ǟ�Y�-o� fO�ro?�1�%+m�DI���F��w�LȨ`���/o^�D���gR�h'�by'4�c�̣\y�PXB�C�������� l0� h���� ��d�
>���%P^z�v�ΐ�l�[mG��g.B(�\n��"(�����F�.���=V�	��5I����n�����Z�e���_1�_3��!$ζ�����m��/M~Ε�-g����@r9��!.��V�סO�sd��&aH�>vV�V�d�H+y�D��:ơ��Фn��e�
>}����#4+9�Y��`^��/X��=�ɵ7����>@:���`�Rg�0Vy��ݣF����l�*c0�01:�P@;+��K:��%�E#�G�fx.'�k�85�Fx
$ Mi�k���~:Dj�4%�r�9S�T"�Mi��!*�ED}��&�#?\��],-��;�����IFa�RX��pXq1t�-���LE�	e�d�j��p�Y-z�O� �4ش�C�܈D��r�T~��_�K���2 =�2���+�Bl�����1k<�g�m���us	"����0��F[k!	�Z#Uh�b���PҎs��eR�̞�&���Ȋ�5�9j�����h�:�ѣd��Y����������5�͊���&gzR5/���)2F�����	*�!�%h]�ew�a��#k��Y��Z�� �0W��Mo#}	�;_��x���A[�ӈ�
��sW�l�w
�~�	?R��m���!T�z�|�*[]�,L!n�������~����C���jS9>�]���\�������݂�������TDujM3Ti�_��ܬ�w����X
?�pi�j���&�
��W�l_���}8��!�z�[���q�#Ǽ޹SU|<�b��!�ΔKo*�V��[�P�W�Ǆ)H)g��ca�ܛn]L��%�{x껧�#�FIb�69g��؝0o`�*��Z�^�v`�A-u�dZ��yT���,?D���4���Lc����Sa���=^Ha�)�&~]��@�0o2�>D]ؙ���Ų3�����3��8n�y;%�_�`����޸~<�m7�ǳ>�[s\C��P��ف,)`��Q[��
��z)<6�p�#��H�;��O'du��!��j ���������^n���%�ZD5�Ts�����&�Hv/�B���3�o�i{*�\�q��M�Ϯt�l��+:W�H^
���N{;>C��g�69���}�o��j2U�/�w��X�9���Q�`��:�,�����<���w�A�+�i�b&0R E:�u���JX!��"d���\��O?�&�[�߰//׹����y�3 )��9�Ca�~��yXE��{�rP�Q�+��X�V����Ew]�$x�'�ןm����i���=l�
�i���x��o��:kܖ=%guW��\��C��U�S!]����[~#0�wxF{R6�9�/
��F�_�����8By?BD<���g�GS�3l��e��oꛅMx�}d�&��Y�G[d���_�
u��i>}nLuGx��mⵁ��b &��>���"L&`z��yՋ�ySf��
��<�xѻG��N��\��Ucw��H�>��;�J�}�&��a昌(�J:����pu���χB�����M ��@o�TO�WIO{�%L� n4��J�����2��rz �:V��#P��\l���z�@.�c@|�~������	`�i��r����-1��R穙	s�Qc�dh�EU(��d��XV'S���i�Mc�Yu̼TJT��;%sV��+J�r���뼲�W�Yn�5����b����A3��Rk5I�[
1y�5�5�pkm��F�xE��X�L���JwY3�gV�p�JY^�)��ݟ~G8xx*��ܟ�ne��h,�"�fh&�H*�V����[zD�}m�Y����N�jx�z���8�g�����f�<������wi��~��}vr'��N�m�d7���E&"%3��f�j8�#2_^5�Ʊ��l#qՏ������q��+��k��D��6���A꯫�S	Ao���kO��[�Ky����Kփ�f����
A-��p�JK�C�7�3a��̮X�p.,os�CÌ���	
uz��Ğ� K-�������#w�B�	I��RSۦ��b��݂}���I
�DjI��XWC��=�ݐ��"-�����p�~��ڿ6&*���Cv;�f! _{�����v[��²�U�f�}w��\�nC|�k��z�����e|a ��[vq�˼����>p�3ތ2m��t��(R���M�W����Ԑ��6H�Su�篞d�K�]�E�k����C^�u��\�r%�n'<�`�7+\�t$���_�F��+w,Q?q��
�S�;S�@�v�?�*z_\ !����
x�JA>em'p�{�4U�nӝ���푹�q����+���~�rM���O}k�sȌ�4�<sU�,���W���ŭ�����G�Z"*]	�-9��Kt˟���	��7��Sv��<�a񧅩��,�t}{3V�a��c�Wh% �,�蚚�1-����
2M��q�c�V� �5�K���-��۸|�C������G ��r�g�@�6NcW���9zU�_O���C:ˉ�q��ƞx��o]��R�	g��@Y\̮�
3m	Yd�mĥ�[c�����U��54*]�Ls$�t��}8*��K�A"�t���[�GB˵c(eJ���i�Tŭ HmP��'L����qHg����Y�W��'+:n��퉙h��0��~��3����4�I�0	th��<������)IF��j��Πr3[�Ǌ;���] ��	����/���mqci�Ơ,�����ibӌ͜��p�r;�u�=�*�E~P��ԡɐ�4D�඿7ƛ ��c���(-��0�{}�n�_��4����$3���$$�݊ R%F%Ύ�����6������t�r��1D9@��p�
�fT�Z
��#�����y썌�%���v��2�������NB�rɧ���K5��t<��f����k���#��D��/��t�t���b|"���
ג�2��c�����;��T�IႩ��O��Q��!��S��1�)��l˭������a�ץp\� G^5�!�Q�����7g�ַ4i��h�[�BЗ�ͪ0.�^�?���%QT�nJ��y�$]F}vb��0_��tz ��_�tN99'�&���|�X�T�ȩR����h�h��f�����zۙT���Д��Q����@�kwx�g5RHt�n���Y�Ȁ(�Z��r�q^���>A�u�T ��n8���!1���%�����2*�N�Lg�Ϧ�uR_5��*�����ש5��qj~��v�'��Q���M��/�#5y��aEk)�#<�?���m?	Z�%���F����1xc�˙�����x|�cc�Q�eQ_ܤ�:g�:d3�mԣ�2�
��3dkҺ
[T_Wr:>U�zU��s����ԌF�����7���]��Z
ݻ�#�vc!Z99�~��M��"���<�)���P�t�ގ&�M����*{��v;���=d3��YJ4�j�AZMU #d���g��`K�6�6�1t�l��8�Y�8�9����vq%����V�@.����4)��� h�<q<Z� ރ��8
��n�ۛ�B�B	�⣬��^J��VHFH.���4����6qV5d�(T���3C����:%��ϺJ1��üpFl$h���β�v�{�t���Z,��8R �4v�6�C6W]7X� -��}a]��}B+3t/^�+��?�u���2Zov*Kdl�)K_,)@w'��4y²P'~��%p���*���}� 8c� �`~�ظ�y9�t�*���Z�-�e�pQ�R!�TM�ߎqC�6�� ���܋L&�?�[�4�/n�2�5�|C���J�����y��~X��RP2��K�>�
)0��3*\�oI6䛌�}�4�EǏU���6x1���i��Q�:JC4�K�(��=�⅄A�)�#��(�qD��j�-|N��mv��#���n���!&	���x��|>d�D�Y����m����@�����<��(����W�J ��*\����en���1g��5"F�|UJy ��1
1��ER�c��5|S�-��m���I~֢��|�?�6�~E��V�����M�$���)�m���Rl��&r��$����"e�b���*͂�z�����7A�-m�쉟*�έ�'�>|�6zC9i+,��NB�͢O���{�+ƅ�����Zi\{��.�B�B.2�mj9�9���U��� :�<���g;}�\�6m�-�̹�-l՘E�m�:�ʍ�wL;
��Z��]�����Sf��8@�O��I��&��ƭ�!2R|���SϿ�n ��=Y���Sy��G��3CB��0��0���|1��\�̩F�ZɃ(w5�:�!��i0+�z-?���B�>RǑG�U(���s 
��2�6�M-���������6�[=��t���6�5���B���_L�Ώ�C�F,��n�!�5�Z���. �#ޓޠ��m���)C��,�l����_��ҩ��v#�P�o>t"�3S��3���w���B�S��FLγ	�+�_�~֤��L
�,�Z:O
�M��*��H�B�{L�!�hl���
H��v��82$���0�� ��
�t���{G ,W�̅\���!̻W
����z`~��c��n<Gw�tٟ׀�f��ݪCt򡱮hɿ9X�ٝ�ߡ�I}�АF䇺V7\�%E�"r��c^�%��/��'���'� x��AF����c
��~OP��P1Ծ�эD�z��kop�v?�~«��f�����::W*���,t���[C����P.�=�{��󗁞X����\k��.P�4�?4�=��<�g~�6����5��O�~��U��eL߳�u�W�AuY�U��f޻��Yh��B�6�S�⑀6�,|�g|,Vb�%~k�c]B��k���]毱�8|,�.�̪6������$3\v�[Ɓ�J����_��/1��1盤������an^ѐ���޹�����F�zpk��Q��Q�.�䷼�0?�kFr}T�,=�ǒx��$Ua4�7��{��� o���wf-��qO��!�I�*�'a��9o�]��<w�t6XD�?L�Q+�1�|��?O�ib�~��	�ɔ��~x�#��x}gM�'u�2O���S��������,��7.�������R��ۤ0�{���WL��]:Cb�p>#{���9}�ē�:��世]���Io�J�ڬ�h��j y�m����¥�f�%���u�I˽u�!��+�4O�����|�1n�ê���6Aj7�}�ì��������
��r;�c�8��ca�&�c
���P>y\{q��ڝXR
(�����y&�?����H�L.o5qg9��vv̭����9t\Bď���^��"t5�\�H��X�>�*[Q0�ώ��1�G=�[S6"T�7C��$�d�"�CsLC�dE��w|F._DG�����GzgZOq+��D�z��D���<}���CA��ė�Tƪin`�aI�_iqP�*�y�;�����l����jC�W���Qkc6��kjdk�g�y�)t��Q|X�/���v�Ϭ�UX�_iɈ|���z��z8�-��C�zy���	���ij����ih�����w�o.�o|�
���_^��f	e�5�+C���~�h&�A���E=�&:c�ޔx��H�M�/��4ZI@с�0��]Шh(�t�ҍ�ЀX�����2�j���3��Q?y�,�2CC�q�H2f̎�f�����$�	�\�A�>$҄��ggN{)G����IXi����2�N���V�%,�K�ҿ�<ڝ;��!y�(]EtY��X����;� V�ڇ�JivT��7���0�ՙrd��a�O�̯�$Dx�R=��KA�ޡ|�h9�2,�CTf��G�bz��-�T�b׭$�F�����>R��Is���7�0`Q ���DQnW����2K��Fܞ��Ք2ҋ'H�[ �����te�N�q8|��>��&���1Hé�k�a���&�w?����'��Q�(�{�э���ѯ�V
c�F�R�"ENsy`��������[)$>��,���@$�u<���吭y���!U�Y��H<�<�V�ן#�%�|_�ɇM(@����|�1ux��χɃ��d_<�{�3҉^S��ʠ�i�JU��Kf���Y��O$�.^�O �2��S/Έ�2-���m�@�
�;.�.�8���(�1��N��0X
�0�ھ2��"����o<^�Bo���9�`f��N��H�Kl+\���X%�e���RSR��>^�w��	3TM_���=�to����mL�jR�xխȏmC�1����+�&D�(�zU�\C�Й]�aq��\Й沚��������O��	���ͺ<����ہ��]���Mr[Y�Թ��-/*�@D�R݋]F��o�a�y��{���I��Y���������vW����A%Xc��h0��5�D�!<��߫::ɶ�~��+%�S-f���I��HϹ�L��5�W=ޑw�9�����-��wl��PSƝ������s�Y��n]�C��Ź������F�zt�9"�1���x<ejg3/XS�/. �
|�6��6�(�L�l@��sEǫ����ި�&8�F�(����i�1_��a��x�څ,����#�j��3�������.W��NԦ�pBW"~���P��$3��#P�a�!�[<cN���r/������h��S]�<��v�'�8B3�u�����.�[~J��� /l	X_�n�/�;F���ڹ5n��"vk�`�D�s��K�׃K����&9�s9ol@�vW����-u5��<Eor�j#�����Ȳ��;#��|/f)#d�#�o�E���p�[&S�e���h��mm�
�	�'÷�O�<ȤJ+�;��R��Ň���Kz\���q�
�`�9ӯ������w�2N�9����G��1U�����;_�=�|���%tŀ	�H��ͫn���_������}��_�d���r�K���>�2�X�7�3��@�L7[{0@�}�N5�ݼ���"w	�^�sW�"���g�Yhg֓�r굟�e���r�����9�QY���_4ۛT1��p
�Q��C�s����'S_;�R�����ս�T)�o�����~M�ho�<��0Y��d��g5��O���F��v)��M�4[M�>�^Ȉ���2�%�SR[����QW�RK_����7�)b�-��T��cFK�i��Q,	������xI�4#��_���|��˟�˱t/K*�@CEcw�z��`�[L����pt�J���ي��N]���Cy��$�]
Б���ǟ���Q2�-%EF���Z!žH��nHg{V��af��Fn_Z�@i����������V�[�|'���Z����^c����a%��j�(ۅ'a�_u2"�	wq漏��-z}Ќ�\����q똵*��xZ�E�h�"'���Wh�^	�.,��(QF'N�t��J{�9/��F	�V$��x�Ӧ��&�Ι�e�)ߛ;ڌ���M���hp*�l}Ι6۾���a_+�8�=��:9�ґ�Tܛ|ͷ��AG���+V�~ܭ�X�6��V�j	w!Y������`s�}��08����U��\�������Z��N�_�)*�����?���d�G�o ������i��L����ҭ�`l���[�S��%y	���,7���*�L^ss�)�����tz�W��w2����ڢP܌�A��⮃�Ȩs�����}G4Ts����?Ge��O%3���#�q���"�2N�a+�O~�!�1�d��m(����6Ϫ7;�;��Z�B�����QEi��h��M�~+� Uח�*y,�ɷ��C?/����0_PPoT%�������W�m���ڒ�LL9ҋ��
:ӓ��Fu���zɱ��fa?5���B�(���9>�\*a{�}5V9ܩ��+���w��id����q�`�xaܣ��U�<��B���>�^*�9�A�hs2�#v� qa�Jl�D���P����+%z���^Y0*���6�y8�����VO�E����h����09
��(j��v�Ywp��a0���mD(��h�*��@�V�I[��4����D;� �8��I��I0�o��©��S(�t����)�_���צ1g�����x�Z���L(�)c$�]ÒY�P_XT�h�������wY*�p�"ۼ0xHKʆ�	c���_�E��N��)d���v'�����&����s,-��'M��}B����� H��,T���É4�}�r�>���$�����o��pV�G�e�-���ε��#�[��$]�<��A3��d*�>Ź~3E�;�M��	<��R��+�(4��'N<��-J㞂)'-���Z1�;�"��i|�(�����U�X>\��Xj:��X�R����.�r�R\ �[�i#�S�&��o8CS̤R��Zwj�Wn��Ґ��@3;�7�?{��R�%~�AyO�[f�`"��`/�c��\+����
�4R��t�ZJCc2�&;;�1��? �￵������Ȍ�x��↦C���yޜ&c�9���b|�(�8z��y9A��	Twbݣ�^+g�Fz,O�V_ʉ��>&=�s�O����IN�sc�$0��O$��8��d�P#���C�kRe�� �Qp����K1"d�ђGY*��R�b���I���S�����}A<z,�a��W���^��J#ʹ��&�sY�;��I�I��L���!ƊhY\�b�d7�Ǖ����L��ng��]��~Zƞ�1+�Fց�Ӭ�s|u�p��_*XT���&�����=�ZS��b>��B�S� <X҄R@^ؘ��q�~\U}uw�
;H�Lzx�wʬ6o�������H[�uRl]0�x��ܫ�E셵�qZd)����\Q�h�\�v^�EӨ�1�v$�jY��Ug�<�R���JԼ�
� ��M*R�x���@0k����W��G1qG�zU�9rKd���� ����s���:�r/���?������L0�NQO��Hlt�~�%[s���O�(wQbWT�I!O��zC�$buc
���b0�aR���R���'�ύ�V��vWD���37g0!0J{,�!d8U{����y^=T2�kS�'�r���rn6��x��|�]6�~K�	���u�F�V�i�o�>g�'�����i��^��AG�`_�0C�~��;��|�h�z�p��cl}��$@���mM�� k�1̤��VM��W'�*�"�_�q��CW��|_#v��H����5�冟�x�&~���y(�ɻ�ͣ�7aCJ���ݕ�I��Xk�����y��Y;��U��g�����#e]�ȓ����?"{��A�$�a�T�I18����S���X��b6�2��L_r�Ov�)`\5�x&L��v�.�3��iu��\C�T��(���j�6!�O=>������sHj�;����my;M��bk��]۰��Z�IB��f3֫�=aGc���&�9'�f�En+R�*�ѦG�SS7O.ϱ^C!��I	Xs���S>�Q�ގ�l&�'����׶|�/���� د�p������ߌ�� I�x�Ffl�"���I{$n�Eᰐ 3���\ˌ��R��;�n����RXH�Mg���	Eٕ �!�{�����~���P�N�%`>kZ��cUʷ��niKT��V>�~O����#�L�t��J.t��9�պ��܋���h��w
[A���@�M!��k}� ��f�#-�lW�!ƅ��*�@�Nx1�V����&�!�y��$4����}���F9��a������S�{9��T��u����U)�ś s�Ƭ����0W���͹a>�@�%A?��S����[D�����;�^Q)1�զ�$S��!�ѝ��P����Nk#x6�o�X���n����8�%�VA.���"�2���7��F�#�ms�c.�ۚ�2c黪R% )�b
���.��)��3�V�
�w�<��k�y�0��iI�WTѓ�,���0&�]��-�u���,S7�*@��s���2?M���*\8�^�
�X� s���r����p�m��s|;cT�� � ��[8t �%��G
)`R��&A�Иl��%��3J$[�O]U*"]j5Z9�f(�� !3Ϣ�uC���=��ޔ�oߓ,�޵�7�o5�L
��>P ��F8����y(����[�(����9@k��y/nZ`���=�j�Zؑ�rî��*&ݢI�x����2�,dL;;D��_JB��G���c�v�d?������B�A*���*n���Y�����S"���8j	��/��uӷ���xcD��J Ϝ��
b���3>$pI�ӓ������X�9����`m�ܪ3��?�q9������fw,�HBE���\RR�}n?}S/���]�_P𶏪Ed
]��I!��m�h,rYN
���T��(���6�޲��o/�%�7~K����n�%#|�._z7a��魁���u�ȏε��p�5 H�=o��%5���PτX(�Ӌ��'�i��k���Q�i� �H}3��H������vc��Q�F���,���U�"S��y�.�b֬>G�6�a�G�j$^e,��:��JA����9A����1��A�˙4 �_��-�,���
���z�_H���\Z9PKE��m|��@7ŵ	��N�v����<�!ez���u�|�P��sQ���W/��a���[���j� ��nc���J�����%m�͕.Y���P�j�G��
w��!�J�v��4ߌN6E�5���ckH�|7歇��ɔ��{5�k�l���tP�8XKA�b��'�jj���d%�B�?l��ҠI4���^��2h��+9��T�/i)oKla�B�`ZNN�w����I�H1���֋PRCd�gwqD{qZsV�T�Ŵ�N��v&q�[wBg�2w�</��kEw;����ԼWQ�p+YxZ�>�=3g4�V�CX?P�u�Z�c���٭P@`�y�+A�2qX��Έ��T�iQ6��ay|��]#Ţ����)��p�	�8<i�%f62Z��DJH� ��@�)�����*�&����2M,��]Z��\ՔƟ�TوrN��=�5�
�Ǵ��.a� 5��I}3Ө#D�.{LF�d�P�RT�S�8E@�Nc��y�R�о����_n����}:C�-H5��3X�MH�]Ʊ��Mut�!�� c�r�=��d{N��>,�u�2�>7,آ�e�|�x�l�"��s�e�bhK.#�s��U�zZ��Mq�к��� <V1x4K(9�Ad������)	J���1�!䑀�v���r���6	��@3�,e&xkx]���o�������ON)��B����f^���>���yX5���q�}DY�!����-�Fچ_]-P�ɫɎ_Qʮ\�5������W�(^�	/y|�{Y�^��I�(�BR�7(�| �j�u*��]�8���g
9���Y=�s��=4 Գ��V ��������
*���sB6�2!���F�����B��M]	]#��/��&w(�D���}�CӮ\����|��.PjrbI��W0�>�\fz����A$��4���Uˬym�2:���ޜ@��lb�s�/�/�.��`�@��ͫF��E1�4zxXCK�B7;.,s������я��kYћc͝�8!y��P�����$���I�8JC�^�?�]V��e8�ڬ��(�dJCP��64,��F��$��O@��	�A��
=�0k�«�t�$��uf[[l��� /�y/�:�kv��2�ϕb.@X������4��Ã��0���И!�.�J/�`��Zj)a&#�t�������q�:� �y߻�ď�PG�.4m�V?df��U=��N�_��}��@���W( lh'��鬇�W]�yD@�:�)B�E���4בX��6id�h
��gp�2�g��vWv��D	� "J�ު��ʤc���}���1~�_N\��pW�n���8q�U��������?�<��<�|a���5z��Ԧf%����I�֘Z`�t�4�ɵON��; �����#c4ٮ2P�U��#�ٞ�#O{��э�P"o�yB	���>j��m�S1�(�M��_�cKr��/�%��G1�̟�~�W�d��Zg?���ѿ�+T���2�6�1c2���h��b.�v�UeƓ;)����9��� �)��*�8}��h ���K�"�mޝ�l%M�v�T.�fqQ�� ��x�X�"��=Y�-�:���{�罘�����t���=g��
����Wj��T�L��-ˍ=ֈ�ה�P�^&?�����J%t����I�^.A���8T���J=��5�L�)��ӏ[5��h?(i�١�)\�=�
-��-���a�eS{?�Ț��b�(gv�v<C�M]�'���AJ�C�4��u�ɨ����'�?���3�Qi{��C�H̟h̳�#R�`�N����s�TK����q}�j���w۱b�&���@	&�=Y����dik�%�VBk�ے�?�p<r�'	6ea9���[w���.�Y�	
��ֹs5@�"�C�5N��#�7!�hy�9qF�,��ɢ�1"~{�]������xm5����T�v�։��s1�Z�(����l#l��8��Ca�)4�ԕbux���L}���9��Ѝ��D�F��b)�*��)|C�|��7����A�Ŕ#I��!A���ױ�v����P���(�rz�.S�Pʩ�e��\xb�w����?��5I����S�D�>,c�d[q�`�w�\�7�'还ʿ���_9lCd,�j��j'�#?~��ڛ�k�Ϩ���DE[��Cli�j%�*}J�@�n+��K�!}�w)F:=χ�%�g��ڐ�g�(NM-r.M�Kp�4O'w���yjx�}�<vr5��(Dp���)#m�2B#�"�@�U�����7�z�ח����ܶ�L������,�]��F�J�$?��a��
k�@�$_��	(������/�B,a��m�띨&��6g ���o�֚iI;��%��g�;{-����po@L���Q��KaG�N$\+�j��ivs�H.�嫞oY��y������X�'���ȿTȪrSh=ϻi4�&K��((�qc_@��Gb$?�̅���0Yț��٢|��y��#�K��H/�U�?4k
%����P�IHG�IO�	bpϢ(ǻ��Z�\�h#�k�.�ݳ�JO15'�n�q��Q}��8���0����h��8�ҹ1�R��?E���j��rxZ�0I���xj�iM����,��m����~kr��>�X/��o$����"[�H;^o��D+F�!�=�D�,Aˬ6VLb\�|�o�*%TlR(D�����QV���u������\���JB��
�ې6X��E$7�5��y)���I�g��u�ك�>_���g�v������L�vZ�ߥ�ES�S����,l��"v�e7�y�t�"B�����ttm����2��hk���E���B��PoQM�＃X^X�8#/�Ɓ�km� Kn^��e�6SA�y~B� �c��:��C�B�Vw��[|_�m�mD-�1� .(mbT��?�j����%�P���H��K&
V:�p��6�u���$T��"�χ�RԺUR�+a|m��@�bE�֘� C�C{!f�b�r󷙝#�e��Y�D(����A�h�,z�&�w_9���$���������D'��U R$+�;9~�jX�wZ;׃g�R��H�w�Q�ʈU�2���Xru"�t�2|r�D�	����?�!ף�	zAٳ�8�vx>��{���?����j�ƹ��[����Cډ~�LNB�o���<
�ۊ��M;N3�Оi+n�
��,�9ኞn�L��Y��f֧�8}���ٽ�0��Vi�HK���N�VnCDT��t-�~��L?�V�����>��)�}<�f
	�[#"�3��a��WZ��bU~e���\k�=���nmy�?�y������8�a_$�^��ԟ�� 0��G3���<��v��'�.��I�P��-�y��OPa;]
���ׁ���ù�ΡiF�����G���������@���.�ݢʡW	����zK5TC�7�_}�m�h�X�=a����ţ��P,Y4rW�XhVS	rj⦖_N���[�@�-�y}2n7G�r��������W^��P��oBP�ڵڶ�vv7q�~�؎J�샮�EϢcl�u��I3����HÁ��ݠ��i�
W�nd1ʿ������2����1LM]����rP����RŨ%�z�CX�S ?.%�����SKU��Q⥆6�C�A�SY �)' Пi�ڀ��\Gy3��5���,_i��堗s �����=��p������楩a�"y�e�֊�3(��`�?�R��Ӿ.d��7��mE�$X B8��ʭ�@P/�-z<��1H�ҵduǯ�z[�������1'%��K��^����>,(�;��b5'�Q��6���}���>�j�OQ�*ō9�z���c��t"#:H��Bv`޹��Z���ھ�q";���������>����@�5��fPZLF�*� ��6�!������K�5���3��V�ݞ�؂L�o�)b%�*T�h�����o͜���<���أ�:��l&��l�:�������=��r�)��0P�w �}��~`I�
�X�Yo{�e`�)ٮr�E�<
đ�')� ��]�,]���f�j_vP��*�1�� ��G=B
����3���%�߭&�r��1��d�³c�ͪf�|(��=b�vT"������H��t���	���{)��1Y��͘C�e��Zb ��h���܆�$n��O��\&Ճ��ݐ�X���5��Ȇ9�1�tPi��h���h�g �_66Mf_Iq�|m�x��<a�{���԰�v��40�KchP4R���|����-�7�2*a�B�	QL`{�������Q��R՜{M��y�`�;duy�O\w�[��V���7k���9%D��8 ԑ���r�LТ����Jvc@G9e�(��j�!9~.�$�)/�4LN�Y���ڳ����FbY�8��C���=u�;�7�1�>rc��i.�
S+�4BE��k�]$�2K���놀�$@���68MԸD��Jw/���-k�r:h�st�〴��x'Ӌy�!%�3��8��I�b��3��#���DH���j2!��;��'��(��{$�]&�x]s� {|���N1���H��7���=���-�~� �%ONj鵴�auK�(]��+��NS�qbi-�?h���>3��]�p)�h����[ H�O
)=Yzo�B���)���(�8bs$��чP��V�U�_�%0���"�Ynk8+i΅�2sw���K,6�m�+��?f]Q��/�l�amj@w�t�Upei ��xκ�z�Ĥc�mR\G��Ⱥ<����ة|z�Z���~/v�W���J����l�`�ҾM0=�Ʊ��Y���:F4-c��B�q7ژ�舖<��`0�2R�)��#�C�B��.`�<R�X/-�@GXu�\ˊ򲕶�"��V��>`���E@LKŒL#������)wB9��p��:�t?8b�$�e瀯�b�=�v�d���p��V�M�Mt�K��/h>�ƯM;SY8����\�����Z�E�yz�O�Z���V[8���Os1.|NȅA�HPH��p���K�-Z��U�bf�y�?QP� ��x�A[VE��HX5�u������sUsz ��s���4�z�5'� ��H�ؘ�z�8�=h�����O�� m����7�d�ؼ�%�SD��k}}���9݊X���L�������
p�Ƙ�0����7w�b&�_+�����+g�_ל���Cd'j����x��+�8	f>�?���_w<ʟk&�i�ZX���0���%��BB"@%�f�f�\�"�&$n9lz�~ֈ1߶߉���G�(�)w�3qm�F/�CtC�Qp!�-�H����C�%f�+�P��34�L���qM���`�xU�M�&ŋ�TrЄ&�:��G?֊]0�eUK��6rZ�>��w�H�� UcH-ڛ��S��[���T�\NPSp�"��~e��	hM�_t"GM� �=#܋j^=�̨D�B�Թӊ�s�Mm��2���`F1s2R��0�������ط:m& ֺ7���'�OYձ}I�J�d)m�o��������R$z�(�F��o�fK<�Ȭה�Ŏ�N�9p�J���Z.zs���ңv��2�� f�)����q_�mj4����+�_�B!��r���LN�
eu!����8�%��|�|��0<��⁍&�D7�g)��!�
�]�ǒs�.#�}B�,�OD�)�})����гԡ�4c��"�Q5y�n#�23E�?\�j 8j���4#��)lU��]���5��*�)Oi+C���A�t�h(��eאN�L�O��/���O�)+��x�K`'�\��m%��e������r��*�f	�Uɦ�Y���5�s���6�#���U�q!����B�N���BrV�w�qPǟ��2�U�!a-�?_�vΖ�'Ss��t9���4L`��3+�af���^SVO�xi�i_�x��& M�i�n�E͏ah�����#{)jE�.K�ϭ��0�Nw�$+ڊ�������+َ��a>����%��'��3T#[A�H����+�8�՞<�	M�a��{m����7q]������7J4_Q{U� f�s� 9b����'�����.�p{t�eW59��P�`ں
"���ݾ�0�Qp��\Z��H�83y���E�.%�Q�f?g���P��=
��:C�O�����&�@�2��F,f��N�;�d�T���h�с�6�Ķ?����vT���\���e�Gt���F�˚J�ʋ�}�%��J[۶V-)f?��<8����$yG?튿s�p��W�����&pi�m�	W�O4���:oxMެ����-���ܻB�L���jw�*�c�?��D�E����py�~�t���B��-�,��h���}��itI��oxyy9��&�H��S����R�ə�yQ s9���O���K$+�e�|�]���[�jZ#/��+<b�}c\0�<�K[��wʥ���4�	tq�=gNt�A�L�F�k �tJ���˄����f�G�Ϗ�8?R�����{��]��I�4�	͋#x���*�\��_��\#��>�EH�E���� t�Y�^��v�PQ]b$X�8�i�<v2��3���{��$m2��q�.���׺ �����%>M�K�-(�lJu�O�]����i��B+��yg�U(~���X�
�v�&j	u��1��Y��ʘ�~���w��|'�sN �k��5�t��.�����"�]K���W�;�(�����k��j|"�7kt�`�S�m���C㫢?�3Ua����aZ{1f�=u!9讐��c�S���Kq.SL�x^'$����q���J��S�ܽ��:�jn�_�p�2�i�w��5i�o�A����;G����v��,8_��h����T��������ؑ4�xZ��z���%$�!G�|Gx��ϣǫ��1��� y'�U��8.q��W�ŵ�ڌ&v�s"��B9���s/�d�Uhra�J׾I`��5����ޞ��U�|��|�;��Ė�'�`ջ�ǫ�X�x���\ji�9� 輰	1�@�)��~������R�1bIQd4�a�/��Yǔ����;7MUw�,�!����r���[K@�ջ��)��_����){�u�Q�x�㞊٭s���:��w-!`wUyp"�������IG«X&ǌUe35ꦋs�ǀ��-�0j���R�f�~s�%G�e>�26K��-��`(�b��=�=!�ʕB&Wy��6�A�����+lPy����RJ�b�c���ǥ�E���g�u���-���O�dd�M�>���ym�a@Vl���Ї�[ �tW�9��/Kȭ7|&�HoU��OП$�I���&&���t�x�r�S���ũ�t�(� ��B���>0��6�{�
��xէA��|̴���>@s	�H'	9�N93�VY?�� ���ݜ3��IR����? }�*�H%r�Xn��B�\"r��0�&� A�צ��~�\&XG�X�J1���r�s��ٖ��5�|�d]��&����"��JG	�B �	sx�#`mt�rإ�fd���@��))�U返�~��$w�;�m>�3y��	SY,�#{R�9uq"\�W�rT4V;@�"G�}�v�����އw�ǎ&9w�"܍������q�i�l�c�f�蚎�,��.�/��ݬ���c�ҫ��6y3��$���o�߻����aaݕ���5���spok`����<OC?��_����{Ǒ���wQ-�����P�r!`i'��v�p���Uy��n�ོWr B%�O�C�:B�88*Vm������ʉ����1���^�C�hX�en�*�8�iޯ�[���]$���m2�cX�[z{~�C�x	��?�b��É��5�₧��	D����wj�ӌN?�����^�ׇ=�Mq�>�sf���YA��Є �5I�څE�}X����C���]E��3U%�#��k���.w���2�:鰆HD�K�t�8�uw��u�G� �Z�ۻ��r��+�я�j�oZw�0�����vNx񿠔����@�лG�C�05���X@gv������Hk=p#�3I�jz�!Rkɮ	gd�~@t�̶i��M�I��{�t6���K߾��_C�"�@�z]��2r��K�C���PݨVVZ�ո�~4D��e>�|����E��.Z;F��#�ͫ��$C� ��CS��+ȉ}<��V߿b����>,��5�����89�VL�C�um�x,�o��V�LA��ʷ�_[?����S� �D�f	�{���EN��7G�����3gN0�T.�d"�Ua2���M�Z��(����26�Z�P��WP8��^�q��a7>Ž��*�՝�#����k�{П?� )���k!^,K,�pC�K� G��*��w��
���	�%�{l?�1��FH�r���C�ߧ�l݊��pP\�)��N2�/i<�c� �ÈՇs�¢�Z����B�/����<��@�{9�T�g`��v��BG�B�����?O���-?��G�
�)Q��MC��F���
����(�Q�1ӭ��Ѿ��7��\~�Sm���%�$���]O�O�q-az朥c���"g�n��n�J��Zԭ��&ty��ˀ��A�Fb!�U-k����W� ͕�Zv=����o;k��G�"�$��B�J�|�Ǳ�e��ҡ�_��d+����$��͹8�6�̓���쫰��n:ֈ�%�[+���=�T��_�_h!�U)�~& ��m��n�ӏ.Uļr��Fr��%;?PH�E}^Z�	������iN'<@�����o�J��_.VH�ȅ��H���\���g���l�>��"��h��U��Ŏ-��~w����el�Up�cNe�PCu˒�B�i)FаH~���MF��`��0��}�v��i*�ԩއ�u�!�����,+c�2�;#J�@�s��"0."�e�׆�8 M�7d����Q֍�ę���<O@[�C�� �Z�O��Z򣛝������M�/u�~��b��QZ�YEA��^�<ݿ<���� �� �t�"ZT<6�h�[��!VR%ol߅�_a3u�
���/�nO�ߗf�[�����_�R�b��`K�Y�}���-ah�8�pD�u�Q��t�lbjtO~9���N��*{�ڈ���!��bÓ	�����:�lZ�c
�"c(��^Czxs�]	�݃V�u~���<Fս��r��L��^�z|�:01�/���1`��R ��9�ê1n����^{�eɜ:�(�MSm<�ue:���!��r,�c53���9ES��$l����"p}�,@@�P�+d8
�$��R��3E7g���h�5~�Y���F%�L��Mp+NʎC��c	A��r��������|�C�I�v�[b5��� X�1����D��2�H�HW���2L�W��qWw���w�FK�Oi���Y�a��m��z���~�"���l�1V�0�N� w��sJG����X�2���T��-=�!�����������G�����ߝa���-�������x䜄�B{߇�fz�:Y�+�u���~�Ģ���?�-�
��
p�M+�`����Ċs�*3�Ve)^�J������1W�
����e���bhgKj�,��V^��N+B�!Sk�n����׹���a-[�6�{��M�𯭸��D�%<$��|70��%Ҹ%�Q��P��R��o�հ� �Ѳ�z�<�v�/u��3��q������V��|O����oS�����"�v4F�W_�٩�k�Dz��|� s��� �>���������j<����l`��I�y�/�q��`��c-��茴=_LchN���Sv���:3QE���*��I �%�?�-=PuE�¹f��jw+���	Q���r#�$�"<��о�H�z��^ۋ�p����Cv���vVB Hb�æD�\@)��h����O�{`��8��ORc�&{��KnnfЌ�	H��o�  Q��r��8���G��r[�sLl�f�?GC�����ʡ�59Ʌ"Q����X�"7�T����
��5�Ox��6^
eB�j?m�{�@���C$~o�.�A�ЄO��!�cYZY��~��/�.���7�t/��uY_�JKH0UY���ɇ�:@���>�q��6��/	��7q�L��o�%}M���Qx�s&�+��5z�[��NS��p3+��Y���h�E��� ��5�k*�y���4�as�O�hة/4��cUA.��t��ȺO��d`�ڿ#�*#��Fi�ѷ� �-����谛zaN���"pU�3E�+��0}s4RRK��nq~�h
�U�	��b�u@�a�Yp��:����.��n���m�k��4)c�@}�ϮW-���>�|D�5��`�Op�@'����1�'bI�m\�1u��|�^>}��}�VP�=� l�q���!��/E�'sF�pus��[Q	i(AjZs/�UlJywZ��� �~��uyNh. L��r��	o�N�FXK�z��Fب�'�(J#)�e���������P�3���b]7�/"{`YD���9���+G�-�~JAAK���v����q\�.m@�hE&�h�pU�O19�{����pt̄�� ��⻮�^w�%uc ����(�6Ycj����XĠ�v$;AY]��N�e���q�'�+m�E$�o2eo0��y;$�kل�c,���?��;l���+h��<XU7:����s�/�/HrU�JV�j��r���Y�hm:��
2^��4��H�Dq�xB�<p�*y��C-�X!��^��NV��1֙=�>N
��pRH�W>@�1b��k��y�q�����D�=.w4�[x���+	���5���v)���/f�&ͧ7���@���ˬߋ0�_��`�ͷ�X\��D�v�R�G�&�H�&��t��b���-T)]A4��䃂cd��S؋��8q:�&ڜ�w�������|_�G7�dCWN�r�4��~�3��60���6p��Q��v�{ oY/#�>g��>��n�����	3��L�}'����`=�~I+H_.�������
�������bv�TE�CWn���o$jc���&�#����O=��W3���m�C,0[��	O�*��9��Mծ3xѽ�R�v���<�� ��NBVCC�Ɲ��پL z���W�}>���aE� ���3���|�'��v�l�T�,�^�n���$j�'s�!��z��d�adAv���{�=����<��̍@G*T�L<���4�'�����vܔ{-|b)s��Z�	yr��A��弝��ƀr�_H��[�Yk�UԣL��bw(����$	��e�En����U���ш���6���uz�@�]�CbϣR����on���\lG����b�#����7���K�(�3�
����7�����3K���a����w�GT\$��,����8��|%1�O�.BPwe�.y��@�f�tuvW�1|���7�>���j���ဈ�ДgGe��l�á"�tL�Z�� )wUz�z�������9LZ19�($��� 5���N2�:�~~�5�-4/4��cL�^�I��{���gZ���]xq{���e�-[�פ~ym���-7k�����P��� �C��A)#��������6�ѐZF���� 𴞔�ZA�)ik���_�*�*�g6�$� U��EvHy>��jn�6Uj�mSF2���\u$��Zl8T~��^U2�S�H|Z�m�*�Y��!����1N�Y$������ʣ[������x�0�g�8~������p#��#+�q�i���_2�C���������X�����4�@E�*a�<��;��2�b܎2:+�?͍��V�f��ǹ�p��>��M,H��7i>M��,����Sq�wx!$x��e�)W��7כ�Ӟ-�g�ę
ڹ���z�m�Sw�X>��Z�`י`�G��f_ ݶ�+�O�hO�V	G�D��]�[`���>���|���C)܌Z��}'����tDM�=��e^�w?I���\�V(P��L�I;�+�h4 R?��	Y�W��s"�+9��m���C�j5s�:�K���S̉鋩��Ql$x�W�޷�"�C]t��3Ihzw�y9��[�����:��� �b�X������g����Nc�s�S����D��m����~n�����&1���|���Ήf%��Q)s��K����qǦ�w��A8,�-g1��(�Z��A�%Q��ͨ������~��b�J�堺F��~#A�O��e�EXCk��8�����ᕪ�7������j
��������I������P��2ߖ�ΰdT $=�
�{v������ht���M�Z ��7RH�G������G����9m�ƚL2��N/6����h��9��/A�юԴp�\�e�ϼ�ޤ�������95'P�>��@� ���ܙ��d���Jԛ��ʮk"2��b;�cY�M�f�� �3S椨<�M����X��\ʜ�p�$v�V�ÍA9t}�6����x�zu�������%����>FVr��߹���"�\��p�J5�P#�ޡ���4o�����f����J=�����x��>�?�r�{���)���vfd�=�}���_�!
�1�z7O�9$Z{2F�����>�0��iv��7)η�*dҁN2R�����s3����bZTZ�<����N)uڞP�C���r��L�-���Hg�2�j�Uª([��|t@qU��l�⮳F ���h����[�$�����V���T�o����Ĝ���L��
�֢���ݺ����B{gW�2.�>3nצIC������,2��#Z�?���Og��U\{?,	��t^���\:��׳f���	���Dwt�o�<�^D�ݬ'�m�^�yT�'<�����:��I�>x�){�D���A�`}�0t�ET9��s���I��k=�������nQ�ː�|�8���Q�s���L� �aH�@�3,=>�;��� ƤZ�U�Z�����AoG�;�v��`���R��h+�(�k`M��@V��9��lƹq�,"y41Fjn�w��Zi�x{Ywg�-8K�A�x �#�铓G�%�S��UV�W��-���2�$����?��Р�fP���=�Р\���M���2
�ŻJ�����<RZ��L��f���{��e���}��5@� ��IHE�wz�^�jV��GVT�B�Pjy�#1c�'�v	S˼��^ą;�_t���b#��/qء�1�~��Sq9d��B =_�\�UP�]�a�0M|#Q�
͟\�&�C?]򉧹k�Js���)yĲ#�TO��FW�t��s���%�٥��ʰ��eb�m�T��d���{�+���S�Ŀؘ��m" �N<�>۹��&T�����L���"�IK���J�щ5��Y���W�yR�AKfR�䢫O/�g��6��X�����!	��!۸��`��J;�*�:S�+	���'�񥚀���[Z`�b�����' ���$��o�F2�c��F*]).��$�NUf���8��a�oH���ٳ�]>���s�yL�s�R�{ѧ'�~b��uͺ�%���Y�p�/������Y!O~��D�%�ʀ�iX�4لf���"�z۷�If/�C���7`Ɣ2�y��O��bD�� ��&{�s��/�t ��_���70V��B�|�8}�D�c*��,�t����]��[�x 7��f���ADLf=B�� :�ryȁ&�xk�Q����8���n�ܰ���x6�k�<�-]�*:�`�����]�ɧ�o-C}�y��C�BR�4X���񼁗����e��ِ����5rXӆ�oV���9�L�j��V��a���X#Ѧ�ܿ
�^��5Pf��&�!�ǝ$���;�i å�	�pO�o�;Mz���4�h7��b�u1\���3(@ё��|+�!=�X.���T�5�t��Z?E�f���CM�q1{�9>��U�r=N0��V������@T�d��6:���暃p���Z��������8:�� 0��^�w�|��i���p#�u���
�������P aWt�$���u�$�>L�Z4��M�`b�+�Ϻ����7en��D�vN:s���I��<�'�j]/J�h,�n�hI��ٛ�ZU�	T<ת��m�}�}.n�5Qw*�B k��#�I5*��&r�'�A�"[ŗ��� b�5䫈���4�"=�Qt�'w]�3�b�|�AXc�����Ƥ��D�%�>�_[��G#�ք�]����=���'�B.T����y����%h��T7ֲy�����qX��b�ڕy��u�
���pAQ���C*�O��x�Q��ʇ�pt�i����E^�O��%��`�^��'��X4���N�c�d�/�$�`S��_�@!8���v� �����F�����s4�e.���ԇ(�p��k�o�����R�"��1�>=� T'��'����ǍD��)��?�ι�\�߳��zlVcq��zb!�G�L�wB�w�ƕ]N.r�3�@���^�����od�z=�ߌ�QX ��ߛ��5��&�!���a�QwqY�-��8%�������\���/�;1��h����(�6���4S��p���<�?���PU��w�ݫ/j�w%EAQ��|���=,wAxtf0�ʵ�\�o��y�y��Q~���5r_�f�U����
(`��pLj �d�2ȇ+��?��
�J��"T0�bV���i��[��c胑��� D�_*��W:���6Hs_e�H��
�v!��x��»؁c5�u"89C�8�cqeY�y�W��8������i��L����?������Ꜻa�^��k�V�;*�K��X����B��W]��CM�]�=�.<�Aʻ��Z����	;v�=P�`�1�PvfBV�e8s���S�@ڠ��]F����*��0$,�ٮ^����{0Iq� C�>>��J�T`k�ŵ��U֠��J���r��D�f��_*-�Y)�G�4��9Lm��w����������MM�=���Er�)�~&�f+9�jDTD���@����5�]TbI�ڑb���3p�Ij� ��(��;��	F�2���؞�b�?�lhuҠ#h���&�dw�� b���⁶,�w[��ҽF���Jt�|�)vNTPb_��"1��Lt��iע2�i��[5�}�#�/5�4�p�.�NMx��,�|б�0)iz� �oO�hwf'j���?0�:�N<+/��jQL�-X��BUT��φ>���8�t|�W�0z�ʗ�Zc�ȅ��#����?�pe���},�UO�U-٩���F6��<�L¯6��;�d}�I�k��S�5�f\>�+^S�sld�G���yb$.�~.�(tGψ�F���~�,E�>�1*��t���=���tr+f�vX��M�m�-,��z�-�"6����l��@3�^rN_J'�2�����w覊���x�u�
KS��2�D'�~i T�=��~l| o�_	�4��������n��=�do��ۖ{zL(��ϻ�#�
�֕�2h��쟵�bP��v�gĺpuA�cj�p�t�#T��M��?����ˡ�U���]o���\�`�2o�ejW�g���g��xg�/�OI��tA�J6�3��;��*d0w�$|D��]��;s�{3�xUCڪ*��d7/sB22��K}pd6�%9��\�+�_�]N��I�B�XV~9;f�ڗÿZ�.RA+}p��p_��s6'ā�n����
��
'Y'�Ug47�gS��f��ge��3�t^�3c�9(��n�
�s�]������̑}'~?��=؀���zL|�ޝ{Dê_�Y�ĕV70��h���ZѬ�Q�`�Xx�b
�ChJ��.�zD1�-b:��^c��{�rۡ�I�2ֹ#�u*��y~̯�Hm�`��{�Q�f����fS��!��Z���U��q��2��m�l�9#x���v7�8�[kh�hs����0<�B���f#��{!	����%�b�s��s �o�~�]�a+�[lz�*� d�?�jz���b��X���x�����
�����%�������sl���bʔ��$�uRlQ��yt�F̓m�;�y���Q[?�y����ꟛ�|��y����CV�b��3iD��;�1<��C��PW��4k�z�J��`i���m�Îb�P�3�/�~����j�� ��g#R�2�����D����\�m�}#�b���S�9zw�&�a�r!T�/L/a�_:�m<6M;ZeE��;tc���Q�^gч�$+ ��N��_�@,��҂��6+�Ù<��~*��L@�D���0A�F��+T8yFz
��L�R����]ү�c��
bpG�A���^�s�(��)���W���o��7r�XE�)�_�SC�-�����C��-4���=:�hZo���f�J��Qpro%���Gb�'�cA�oL��=<�xwt'U_H$��3U�8 ͊u�y�ķ�6�D��t���58�������yUe�z�ϙ�5`�$.[1`�U�g�Z �{!,���Uds�E2�0�}��HQ�"��MUp��r��^�h7K�Ǖ��dg������DT˵�� ���v�[ߛn�m>�x� d����Ù-�{~ӣ�_+��v����s,;�
���O�g�-r�StD��e��=Q4�BC}#zu/%�P�A�p�dk~�g�Qwor
h�g� kՐ�y��K ���l�Ʈ�a8��24�'-�����>;��҂*�=nu����Q��
D�|��l�@����|X�]�\�	ƈ������Kv�6�mw�7���pñ���]Ģ�<�ؖ���c ]�Ĥ��bWJ!��)��x�&P���A�0�x�����dF���s�Y������.4��I�B'R�'#X}2yd���2��mW��}P���#w�69u�sN�sR�3�z�r��h:� �`9P�M��>�@�3�<�%֣����w�	�a�o���͹��qB�Z���s��d+a䚂����h-vL��M���g���g``* Mt"�7��WP;`�NG�҂��
�D�����8(2y��X�Z�<�z��Di��=�Qvit��=���pMY�kA��+6�@��pd������0:���#�΢��ơ���Ey��byjsQK�iY(��_A�D14���M{4e~;׆��mz��o8j�e!M������? ���?�[�>Gd��F���4 �*�)ϫ�����,�`-}�!�gޭL�ߦ�3`�ZE%Z���i��Q�i�ផۋ�G��+��f��2rX�zd�M?>��nM4]�>�d~e�\�u��z��5�g�<_���j�w�/�������Y�Bg��%��m؉�T�5R_"����q=¤G��͐"�T;Z��"��Y-b<�*�֡6��Tj�rr/��� |�*�!1�)0�9#u��AP:҈/]�	��x?n=�@Ů��<� ?�q=�&��8B"(t@�����T*=T{{rg{�D%�e,,�6��Q����4������7��2K�n_@�beb��}}�D�KAE�Ry8������D��K&n�����/�ͺG����[�I�h�L��s#��zf= ����w���z����Xe�F
NڃP��Ҳ!G.�0�/b�P5E����vT��W����� ������MY�_c!�ӌ��=c�a����)\GT����xc�����E��N�܎�z< �t��Az�ۛ�j쓾�T���B����(%$���9��l�T!%P�E�]��DB�
�~sXݱ�I�|��sӓ5.)��&���˝ܟ��@Je�:V�#�H�/�z�uW�Fղ�/M�3(����p��|�ՇFڽ.��ow�1
���$oBO>q[?��v��Ēj��|X��?J0�{#���p0��I�e�&�ے�
�n{�#����n���@J��WX�5���# ��	9�&qq��_�>L��ۻzZ��O���]q�,]�`lR"p^O��|S�{�iS�7T�
����O��\�ɛ|�����ˠ;���S��!�~�+F띛��[�鞍�'�ѵ',]���ZcT�S��a`7g�{����\���w1˕Q�E����.���my�P�U�����_��������΅$|�¤V��������^ƥ�B	�2Lȇ�S�m��#8�|��@&�Q���+�[����M��Ꮢ�M�l���J��G���	�a8�z�E��v�5�YM��F@�	߿��߉
�ƃJ*�vu2Tw�m<D�FA��L��?�X<h�����a�E�9V�e緟�У�F6M�oc�wu�ڈpfc�og���07�#"|;�z�$YaK�����>Xo�������Ls��`QKiշ���SLU��D{pa����������y�X���3�� �f?&n��l����1���s��q[�%
��v/��؝Q�Th#��!�m��y���\�ڮ9��ꋽDp�:���L!����5�݃c�Kn��27�T�&_���Ha��d�;(�������TLg��	(i�-�i'U�0��z�n�1�뵬�r*��U��a���0+�#���<���ksL�g� � ��G;�+q���w|��y�}&�����*UAEA�VB�PL,�8QF[=�[6@�ƣm;p�O�̪�j}�t;�-ű���6����p��ݽ���fav�MѪ�|>����5.�@AF���G��a9�V͜G�"�ٷ
�^X�6�
�Ϣ<�v�}:HI�bʟ߄�}�x#�+A��.2`�#��6(�Ф��)հ�u�Lk3��T3E�]xGVV}��*�t
����ϋ��[(&��6z��ư}�t'؈�����%,Ԃ�ַ6����Z�{��33�L���|��f�w^�y���K�� as�HX�^�w�y%u����Z}�t�~(��a@�S�Oy?��@�S�6�I�:ϒ�?�n� �kJrll��Ѐ	w�"�w'�j��V��[Gꎁ
��s�LP��Z�hk`wcA^��IL��̜t�~!	�)��;)�!~ܗ��|/�H�0@����l��T�`�#�)��#C����ܚ��#a�ȇDV7�'��7�j)�=����h6�@]><�ލr��ZBQ�*5H�-m�^�����I��(�)�ƨ�������|ı�����c�ea��j�@�O���_@�x e'�0J��,y�R��Ry���7���C�Z&۰E�6큂�y�}h����� j7ޥ���
LY�7sՌ�Y��	$R;�mF�B��R�Ӧ�]�(1�`Anֵ;�JO��KBco�X�ߪ��}�T���^�)idV��U�e���'%X�S��>���v����r�%"�-��O)J���i����="�k���A�� &T�_��~�J���Y9֗�RЫ�2C�C(�~���#�W�GU���8�v������N%x*����2�>��ݲj�2- w�\G)��7 F���]�H�k��|��DW%8a.��Uj��η�aY�㼥M�p�Rb������>>�=��)݈�f�
!�(`�d&o�>U�阻o໠Ծ!��e�rK��\���S�����g�ų��U��^V�,8A~�&dfK5cNY5��c/�����+���F�LM��{�LM�U1��5)�����+��#q+���n'%^�s.S��N�W�W�R�5��/��4��͙��%lj��::�O�*���?���_�����d"!�5��[>��O�i��t	B�-&[!I��km<.�h��X�tU��5�.�8W{�qjB�W��d����� ��S�j�+�L��D"�/,����X�u�/Zқ���N�ȋ��1��^�̏��<��"�lF%�^�`����;+삏�sܶ�-痾�L����aj{
���B�����L��%�?���AJ!���Xf,"�����iW8잓�¬�כ�]�D/ZP²��J���� �KN|TA9��.pfӦ�ӟ%�&�[H��Ĩ�l�$�Øܾ��	'�1e>y������>�h"�"��u����kJ�~ޜ�a�85�Sl�m�}�E	���X�!]5�&�c�D\Lى\ڏ��Sx�C��i:�`�w��R�`����73@��Z�>P	�sIF���'g��tHp$�{���ڙ���ω&	v�1�OE�9�+
$ԫ���փ862����w�:�Q.���,$b?Z�YB�)a�!�������)�
(�<�;~�<k��%�y�D�]�6w��|s��Q�r�Vy83X��~�_����(��5T��VWП��$U��r&eN�� �b|#x�����2���E:��qk���^��\Ґ3�(��Xf_�EØ طB���~z��X����t�S-�F���xa3��@��@��X�0|z�<�����|���2����� �$Sm-7�a�op��:�9��)Aj�i��5�2G�B��I͟�*B���P��o����ܣ�(��RV�b(�ؗ��[p���-���Q_Sܢ�}8����Z�:g�'C��w�E�G�}Q7v�2�dI:��^Q��'��&*�ƥ��  �����p�o���9ŌQz�R�Ć����ۻ��ި��8�Wƾy[0���7;� ��)i�S�߉jMS���n������pw*��P��I2F�)�v�&��U'/ac}��얥�A}6���ZRM�J`x���������(3ݹ�������y�;�T~�]���9����㎊\�(�+p��3��l?���a��	�� V�����^Fj^t60��M�5���㐈��w-�g�Dt��0����dFj��q�se(��*T����+�C!zUU�9�%�1h�t�X������r.�eY喋�}+O=5^B��F|?�����&RH����k���8ܚ��o�|�Æ67� U�`��UU��i~�xԷՅ71Q�'�7?�J���ڇ���2�ށψR������P���J�-��k+Gp�
�J����U�:�q�@�e�vy���w=l�Ck ��V+4��s~"����G��@�=� �:�p;o��T�Ǥ���g`K��
�ޏX� �#ǭ̠Q7/�z����&���p�B}�k��r���(	�	��!�bdӻ\�&vW�t�����6u�'�P����Q%.)����R�Jh{��>W������s�J�r5���y1Ui���#r�X*oͬ#��A$N_��
09$&�&�����q�!������ �Op���8�(C��b�]+Oט����/	Dۺxl�ЦTQ�h�ur��.�W��P�ț�h
q9� LL,+� Ły�J��IG�r,�L��K߻�Ay�%����� �g�s�V�H���p��ph���4gӄ'Vg���p]���(��&�X�a/=	�ɬ��-��n[�]0��H�7�ǵ��:�aAb��oV���!�l���,�Zv�j��Ϟ�%��n�B�'��$��N��!1u���o53�P�F���l�]�bÐ@�T
ۃ��>p����x*u�A4�x]](�W�1a��+��=pz�kcYg�//�:9�:�}�,%��ݘ�0�O���bȲͺ{�{rO����F^�#��Hh��K����)*�z|�ׄq��]�쎠�ȝ̢Qc4�k?�s'�h�{}�.����1mfzf�U�bP��e���¼��a��U,N;������f���b]�F�B@���݃Ҍn�l���+�"ZJ���]�Aa��_�]�oW[ܑ@Q����U���r��/ZS��3,�9���� r)�����1Ǡ����vC��N�݈�y�m�`35`u��cGd�sz��آ�);cJ��P[��9���Ҫ�~"	�
�u]�ʚ�����]Q^�D�E������G h��BkF53�ZtW��믜�H�Ie�y�]�;#����YP�+�F�3n$}��8>�9$��\kw�����{X���+��n�hI��Gn�C���h<�3�QJ����%�,�˖�8$��&Ȳ����;�Z)i��<r��!�1��1從:B+�dH|K��(�!v�\`~���P�:00�,c\V��"{3R�3 O B؛��z3���gr(����ɠ:�m�ydx��z_���X=�U�k��ގ���b����6V �ن�B5�z��j�ܾ�Q��\����_/����;Y�/�u��l-��rV�̓�M��(QZ���+�
��8��5���1����i���2 &:R����~Z�.@�^ ���Tٓ��I�埮��	)ύ�2��b2a�$�\9�*4\�����x`�됔C��_sӞ4�5Ν�W�<2l"�RM+ ]����uΫ�*Qa"*��#>�Y�Φ�}��	f�M���Ţ��F�@BS��e�l����fqf/�<Ϊ~�QU�-� ���=��+[��r�sf`�֔��ݞ���AVHA��� v>��#ü|c���J���d]��Y�ɘ���dDm*���Yw�ʤ�O��v��~�*˫��	�7�ν�E���듓�����<��7{?�ζ�������:��~"������c�.�E������|�ք�W|�a8���s3�A(J�VO&�pf�*Ԥ^Ї�9Bv��O@�a�h����"�L���Z� q#;r��pIi�MP3�}F�Gc�Q�k��6��L���ZZ�\����qbf*/�X��vR����$��kj�D2�[�cc�Q�g8��� m����G_�!�"g��TU����e��b ���7�� ��ś�Kg�C'��3옋>�6Xk	q{��_��*���,�������g@�q%�T2��k�=��c�a������_~8W ����K�v�7u��a���.��2���D�V�D��ũ�4y�w��$�V����B�<��9F���cv$>�Ym>���@6ݻ�|[��^�KR�͈k�wO^�xL��+9���<m�T1��Z�hO��������#��v�s�_4g[��̪R
��f��aL�_�L
~�A�~g ���N���H.��b�N�n�#�������j�;H��2G뫜����T�� I]�.l�gݥ"�	�,�5e����Z����1`�GA)�D��1�F�8�	�t���HIu�;����Q .}�s�����AD٠�͗���[�|��B�oSMTn$�}Q$�J���ƪ!�\�K�����-�۟M9�b�+�p"��nB�	���R�T���#���6�͆������5��#�.vy-��E�����7Ӵw�2�g'4F�*l-�wt��"���evr�[��$)g�9�>�ϲ����q�,�ѩI�5n�\V���Gr�q���C'7۵�`�I��o+Fch�������V�W�g4`e�c�lJ�o�J �Qq�m�c�2�:�!�?/��LGƾ��4kXAP��\���T��dF~O�9�kK�h�27$D-"�:��w=�U�S������� ?�,��.�-��(�h���E3�d%*���I,�%w�G��l�G���η�`9Г�Պŷ;Fm��\Ne{>��El9����k�M@���'N�t��o�&��y��y�LK}i��os�����r�F����E�� $(�FB�O��ݐ&�
��B������SӚS~p%]�X,TExD&�XŁ���l2��Gc+�pi��� ���J�0좁h��(�v.���$}c�IR��ٲ�zW��|,�盗��v���_F�~e1�La�����2���I�j�:��j��}���̹���P1&v-n^�>���
XyZ��T�	Lv�ֆ�v�R<t�n��ݎ���,��g �;�w��0���U�Kdw Jq~F�h-�����T<G`��Gk����&���]�@?,֮���̅��wSizn�Z��;a��y�#�(�;x�Q�hPD������ߪ���*��Ѽ������g�4Ĭ{�� j���.�\��m����}Ǻ�1;f�^�j��ٞT�Xgp��دG��K�p.ȴ����Y�C�,Z�X;zs���x�[K��*9���v�˘L�_�G6��
9�s�]����I�$v�9U�����k���C{ǑZ��Y���{3�J׳PR���v���$��Òdܠ}F!^|�5����o�Xz�-ZҰy0 ��VU;i��a@^��s�d���������ʇ6�'_��O:�1%�j���w}z����p�}`q�F���ޒ�<�66`&+"���׷�IRk�(��|���x8��@�y���f�A��?�J\� ��_/�� �����`Q�:=�n��>��O��6��� ��
>f��d����
��jL0?͠^{+誥z�ɟ��*UH_=��;b�i��.�
�G]`~,t9M���� ��ӹU� ������
�J�6S���m���R�v�!gx�u�'��
�`�^1�4ֹ��om��ӄTW&����u&�Yֲ�s-�0ЄqdZ6�K/-��{�˨0VT-����N�ҩv9�|\\��̟������;�A?�5)Y5��,eqhNG���T�Y�Ի��~��F{Z'+[���p�o�����]�����=�#��#�:ȡ��Xt��M䇯�[-���_E�j��&B�5u��] ���]o��� p��̦w���g</�m����5��y#�o��`?b2 ��fpn��[NR	�A�O�s*����MA1�����M���!x󹉄<F��.��i]���!��d��8���ƁSx`�Q6��CkY�$$��ie�3Yѫ\��/���
�ň�lm��v"n���R�w%�A��l�h$]���j' *���t����*��՛L�K������������u�˔o��������o�t���3�S��O'�}�(م
p: :"����{��su���^^s�%�\`1+��q�S:��RyB���ʵ� ��9L�U��G[��l�X� �fHDU�>�n$�2�������{�Y�i��v�Y<H|� �]Y���E5�@�g����҃��m�z2!�6b5&[��)���ω��C4t�#���Kj۲d��~]���G),�{:��7��� �/n��~9�����+��(J/�.�Y�r��l��oR�	��װ߻❚"�
Ѿ����V��X����Z���X�3�v�<�(���R�Ùd�؈\���H��"_��j�p��Xܴޭ<�eJK�ϠM�=�dE���*o����-�����
ũ.�}���1��K&�DL�H�A�8_�|��c�>�b��&#�Ճ#�I��MQJ�jH7�v+�]C�HJTV�m�&���X�!��d "����T��	����;?�
#�f�ɩ�٩S�I��:���V�y%L�O�w�0�^:f��kۃݢ�9[���v�a-�1A���p�C�r0�b/G�鿙fJ���-j7���r�(�q����������� �$fu?��\.1Q��O���4`��j��s������uiKyT����-�m�����plG�a7ԋ�d���Slt��e�acU%伅t�Ŷ�� �?�+Q[Z��cg��(��U��T���5X!"ſ����$|>�C}MV$�[�Qms1��uj&���kE�<D6;8Β� �B>�H�ɨ5���\2�m4A�,��0kW���((�:�<�øjL����`:{*#Q���`[�������-���_�j�c�@|�Dj��fԟUG�����a>����>%4��c��]���(�ɝ2Ɗ+�A�w4�����ߨ���z�|�N쩘�`�&p����K�l�#E�l��#��-��B$p�?�/SX�M��'^�R0��4��]�#y��%��4C��b-������{�,��E��yB�s�rk;��!�G
WT��y��#1�ݟ�)1j��4	�lzE�V�b�g�;���t�E��M�V�:oԘ2W;g��r��QV��n���R���g)qI3��-S�/� �h }�P��	#��ה�����Vy�
��mZ@ 9�R`�>w�㭱��	���N�\�LLvA6oz�] TGe���lN(@qs�lN�	Ĕ��"��Jn�1Eܫ�����-����ف<m%�ˤ߾���;)���}��dg�8�H��ǽ�[Mn��/\Zi�9�E�i�9vtM�x�ʝ�I�Є�N�Kx���B%.#�!�X��V�ӈ���`�J�@Mk����1TA�]�|�3�5��V;�x�sQ�.q�>q���I)XJ���������X�R�t�o�|���#Aws��K>��f����]��G�h0��`Α�E���������ɗ�>��U����B
�.`G.Ҁt�����SxW �T�<�g�+�����h6�2v�3.P��y����"�j���w�N��� �U� �/ٗLvZI9�ǲE�-eA6�av]+�@���+q	P&qE}��_�~>�g�<	�=c��̵|�?���v�G��p��aG�6ڦ��DD�i�_���dh�a�N�kq�m��SS���m���JmF�67A-RGreBKs�c�`�-��Г���^h(�l0NI������0J��t�?��������2��fj�<|��w�O�t9¢��TG[r#Y���p������8�S%�2��1�	��"�e1F�F�I���Tiﹹ���]٥��!�2�0�V�1Iwf�4^���9M��^�'c=���w�ț�Λ&�x���ƅ+6"ы���1�+iܟ��v4��/Q�	m�Bq���E�L��Ǜ�o?�� �T��&k��+�9G���yCz�����M�0�O�j�"�S�Zʥ���X�}��cb��l
M�-��X���fd+�2��Qf��,�D���=��z.e"��iWB¥!(��\�������C�3���U`���,��:�7����Kp��$�����v����j#Hk ���M�+��h��L8>���vus�J��luۍ�v
eiZ>Wd�߃A�z
��.1:m�~�>�b6���vyǪ��U�S|�+�T N4���#y{.=��L��r�ZSPZ�U����siQ��
F�v��9���z�����F�S`	������udB������5=���3Qw���2&������qr1-�i�LEwm�@E���w�Kt\�L0�#.���l�@x)��RfD�� �Ͷ���.5��tV�<�v����j��/��|���5u*�?����ӓX��:���o�d���
+�kE8��fȏ���OɈZػ�aH~a��	�d��7H�Aa]�<j_Ʊ�@h�{]ʷ��h^�
�!`�Mݢ�<h��R:t��B��F�a��7��A�^5��/�2���J�b��IC��?w�LAШ�K�Zk���r���.�g�C�{�5�6�;�Tb���E�Z��7o��ժs�+6}CɃq��ڸ�ެS���Nu�7O�D��s�����+�D��# +Y���e�3�2`��aUoVl}�b4��-�mQ=Shk��Sw㹭bM)N�iwhx��,I��i ?�,���/|����W�i�g<E����,46/�!���8�t��<]����w�T��jv���.1t��P�l��ް>��7{�����+ֶs�F���]@�Q,1v�a�"0��M�nIfAp��s��$�uj�tI�í�0V}@;棟�[��O�_SN4Oc���	ζډ%�.��5�.��A�~�������ogiĳY&����rv�op�.�jS�U@��m�u����}��h銤���ds�H��L� /&( f� B�*���K\Ƽ��nSC*���0<��v�k��`xuqގ(���"*��C�Ç��=} B���]na�~��,�,�_���[5����j �$��r�<��7��\�����Y0'ƺ�����#��4`+r@+�A�Y�J��-}�E8Rg�m;�m��&� ��)Nc�����	d_�d!����`h����`���L��65��fpޠ4�Km� x%8F�t@mx(�[��ֹ��K9�^�;!��;�2-��P����_g3�ߒ0&�:�	�Sr�)Gc����<����v<v@q���~� =�ӟ`Y��D�,�����^MLd�L&�Eg0g��������B�[\�B���=�f��^����:6����Q �a��Sn��I9�ϧ�l�W�1��G d�����@([�l���P��3��������v{��B�{Dĸ:�y�����I�^N.���B�(���5�")�����qt �zS�oT�Qm����
k�7������F���2��=IJ���0�C������z7�����<#O�¦1|v����G@�*��&��0t.���WQh��u9Q���gV4�D��4r$�Z�+�����F�K�<B���ˋ0��Č1�s��/�^�ZGX����ǃm��|U�'���ۮ���	�Nz���,*����&�e�veb�,�ĭ+��p�:��Lo���K7+�Ű>u��X���c���-���{��*;2;�A��y��!�0��?�B ���k��%�h=̖��U H���T��L� 3�ь���V48$<�u$U�+�]$Q۳X�Z�5����?�ɚ+����sA��������� Ä4% ��<�����N�ؾ�0�i�K�
&sO�������[��~�*B5P����u���q&��|����$aRќ|��N%���.��)�=g�A�� ��=;ؑW�ZR�c2l��b���c�2�}hc(D�ĩ|�����F~G��'k��ޞ�Sٓ/
PuP�GY�v������}{Yj�xm�VW���}s�#\��0� Q�dMt=4���8mx�=�vp;g�<P#	��<��*m�`5?^����l;A]5h�w�|U�!�,B�9[���"��TZ.���qǙ	A7���j����q��;�b�\��iQ����r�{M���ƪ�aVj�)��͟����N*�I5���x"n-��>k�c��3"q��۝I�2�D�(��ߎ���t9ό���xz	����h�O�q�z��S��?8-T����T�r:��Q�,��y��re�ڛ��IΙ������`I��q�w��H��V�*O��'r��N�F
��$���X���|�(��|?�J�s�MQ�"�9�{`�ܤy<~GQA��������M�nf���HC`���+��C=
7���T@�l��ԿYkz�����W�y�������r�H '������/�Fi��Bj�Uj��g�]�;��y7�������wV�C�K�ɺ+|.1��!R��u��uz怔���>W��NB7��D s#�-��n�H���jڤm$���&�y̢Oh��2�P8��`lը�'$7sw�R�-�M����[X��������T�w.<-��FD9XC��)�Qc�@0��`�L��Ƥ.���>�@"�Z�V8�����H˩��T�C+bVX�mƩBm�[�9�?7�X�I�Dy��Λ��ҏ�èS�.5v�]:��LDfݔ8R5�k���{�W��d��5����ʳ�� x�krrR[�fRh���1!\�:O	�C���Y�����������@��֧���O�R��[����rx����z�}���P�W����J�� }p!B�)
�%"��
E6Rs���]���翤^�Cf������JDa+�*d]o��\'���w�Z��r�N������Ҩ��v�YK$؜xS�C����z�5��4W/1����4�����=Zpx�ˤ������p�$��*�gy�dAS��֧Cv���������c��L�+RIx*\9�g>�����M��UB�N�7��тAܣ�e�y���*��ײ:�i0���	9W����S$fh\��U�Q�0Q�Z�8
J6oY
�E�)l�T;��u@�R�5ݴ7�ú�E���˶#<��H��"�z�J�> � ��
�D	�$e4L�:i��8ƒA�)͒(_�@fd���'|�J-�j�������nFq�7P���X�i\�j��8ަ��������)�_R�#��N5;խ�/���*]�M��o�u�%\�n�(�BVJ��C����&�{$0���!�Й[��P�Y>���I������C/�+<��,�L�i�<�����nt���VB����A��{�6����:`��R���) ���K�oO`��;�N�2�0qM�5��HB�`����T�J���gS��
��h\R;��<3�����f��j�e�v ��A��e�nP�ˊ<O�&���V�2/����Fa6���|������1b���e�BMD�=n2�x;���EO�^ZT��<��~��?sI`��O�T	�ʵx�Be9'S$Nf�O_�L����.��"�U3h����j����]��3x$�Jc�T���543����y��}�dS��Ꞇڷ�ˌ�^R��6?>̂�'�z�=J&��h��
$f�((��q7j_=�N�����P�n+�|/�g�#O@������9�M7���pK/�T�Y,S�U�"�����)�9�q%�__\�GC���������m��*g������!�a�d��A����_zrhS���b�:w�R�Oj��0L��sp��٪I�v	Gn�C� ?�����Ȍ׀H)��.]�g��t����(7����Z?(v����lu��a,!`f�Hyo18�.��[���c�{���wi�h�5M<�0��T��u��~	t��2�X�x�و�O=�����i���5�Y���:�
A��x��ӚCy̑4Z��z�"���^��6Vs�Q8P��<@�KSb����o��vR�l�?z&�G�2���{����\�sO3Z4T-��&�)���{�JǇ�c��U[�V'6��j۹�Uu?��������xC�5V@�y6:6"S`�a:���/Ljp�@8e,��p@Z�C�'�x�{򴘒�@<7�-.��A�>�Қ��m����1��K��$+avS���F����BF�@�1
$��͑�B���$�y�?��/eZt;��� �أp��ܣ�9
�I(L�wE�v���#��G��2�W��	<����0_�a5���'������z��S�3�B�'�����̞ L��$�
��O�ձ�%�6�����[���ˉ8�tD�6�Aj�YF���h	)|XK���'xk!�&p!����K@}1����0&v�Y:V�!� b+��-�=	b{x���n���=K5�	Q������ u�y���[N�÷J�i��>1?s���Bzx��m6�Z�^�����˞J�\Ɏ��0����6������+������x��ߎ�j�5���ӆe.�ߣ/������k�7M-����P �层ϸBWj��̅^ ��,Ħ^�?F�i/�+h�+��	;���r��a�W�b���#np=�=ku�Ps5�|Tpp��ƤO���5���\���?9a�6 ��W��p�ݍ�,� j���9r�1&�5\�YA�~�kt/���������g譁%Q��n����� &�D����ۣ�Xyy�y6�2@ק[����raEK�	Z��[)K�"���o0��cX>��	�ϽB �ԡ.o�_�#�{���GٓZ�>m�؟ߺC��L�7B�e��'�-$���p6���̭��u�O>P�^�{DS,��������Z�ӿ0ᕷR@�e����D	4�o]epɘ����$������La*��c������YޕI1����uK�CVW �)�fCI�&֓Ur�%��Ll���%܅`uK��L��l!2]�A��F�F���!p9V�SM�X|�v̠!�vJң�R	ٹOI�2�����M��Ϯ�x=I�r�AR�2(�� �S2�k��F���
ϒ�g-S#kzX*6G��F�a݂�T�"P�m�c�K�9^�g<?�_aW�/� �1Glht����'�ϊ�n���dC�:�ID����HK�`лtJ����̄E(�9��|������6l��V���c�(ߧD����� l�v�bI�7�%��ӆ��"�����\'��˛F-2��C�n� �DmQ��ǝ)�13]sn�k=C_Y�C�mU�_�KX�g/ӌLj�W���W�J�JRTeY;�$�噆���c�η�.%Vb��}!f@� �Bp�b	�0g�v�,�.�y���nꆟ��6l͝tŬ 8;��P<���nL#h��U?�L���$���)3;�;���q�M
�7
d��R�;,՟1̃q��-+�E��T><�)~���j�2�W����:15�L�"d���i�A]e����C����Ñ���~���k5[!8��� �3��n]���\�q^9�H�o��o�#����vaZ�cAH�O�Fr�c��_(��7W��_��E���Uݵ�P㚥J�*�P�aR�����^�$9����ɋ�BG>�9�&n'i(콦d�K��)e�e[`��M.�h��%[��7:��GtҲ�'���k6���s�3N���qU�E!����w�CH*AI(G�8S�	d�M��[|�/vD&U`���D�J�h�Hʇ��t��M"N.�@�_&�����T�ư��.�?ɒ�G��w�F���V�Ǝw��T�ۼ���7�L	fC)-�'���iy DB��c��nS �u�+����,4#�;��C��&Kwu�!�e�w$�ɚ��427���'܆>�-ɴ�\lF-m͈��~���/��Z��V�?;#	D�l�7��dhV��D�Ӝsl�He��0H��4�Q���ػ�B�l �0<@��b�dK�Pp�Ͳ�F��юYj͠=���C��w:s��9������<62�mY)�=`�n�
��39�}_���e�M9���,cRK �͞�%��vfU:A�_F���-�T�ֻS.��o���k�i� ����KQ��pSg���df����a��nz�@��`�f�Ԟw8y�8�_n��<B���b����4c�Up�/�V���)�ͫ�
��u䒩�B��#��Fc�+4I���_�bDS��L�۵з��S��IN�8�M�[�8�3v���)�Q��P�Q��ՙ]	�?4���p@@^ӥ����jc���t���v�.Q���b�~|���(a�Ӱ���r��h/qsND^����%k�g��4�a�S������L}-�: -[f��r?���V�T@�X��[�A��G��&n�	%tf��x���܇K���p����1j��okb��Ϭ�u���s��=�.v�$B�SsAqv�bS�<��_��۟�0JP�<�M�ϚS��٭d$c9��ɝ*B������eXk8����j�
{!�����=�b
4��9�)�?o�:�Oq�$����`�c���W�&�%�ƙ��G���e�$!'���3/�z���W~#��!0�O�Қ6$�4Fu!J�s)�h��-U��d�T��Qs݈�
�Rrތݺ�Jò�c}V�pm/��MΑ��?��^s+�׌�s8Yg�=ݻ����+�a���?��g>1��w�a�����N�y�`������D��)O�d������"�֋{1�,`[Ç�Ä5p��R���/l���M2Җ�f�b��,7�i+<�J��y�=�v�]��[�м��,[��k�7Y&�,�q�of՛��H�Y5�?�����������Q��:JO��J��'=i�!ߣ�l����'�򹋆YY(z[z��)ɼQ�[�\��N��.qB)��p'	`��S ���d3Y����/x����):pTf��p�d�	2AF;l��RS��0�XU�H���j����&��e�Ĳ|���4��Da|������#��@�J(ʨ	�d��Z�_����} �?�0Qُ�~~���f|?K�����ƪ�pOm��TL|�
�In
"-{�I���C�r�˺h׎[�\.���#���S��7�=�e�7���1鿛]hv�7_�*v��%��av+a`flV��O�K�B�{~3��M�}�q8����;�K�H���O�<b�����m}����
i1ǯsF�4���{e���h��=��P�@�A�]�����&6
]^����/�Ӵ��|���jƟ�gk��=�� 4��x���OB��"�e�F8Z6�Xz*���(�U��^�� ��M4��  F��N�"c&8��9�VWH��D�v���b�I��)U�"��7{a�f튋��[�JOe�?����+l>��	��N�![�ؼUBP�H�w(S�e��P��d�Bz���5+���y����9��L���D�C���ͣK����P��6�"�6�vL-{2i����7��x���T���4��Zo�W��׬#�����������^�=�
��[��U�S�;��e�(�i��aߌ��=���5��k�m�x�\��K�3'Z�Ic}���ps�Y�5U���h����=��R�1��XR���y����E��!"s��Pn#�,��{�dڜ��?.o��|z�]d+�^d������!�H<e��~i6�nB\�NPH�V�\$��dp�ܵ�w�
ŭ}���v�q��Q5^`!�,q}�7ꊉ�%��9~�{�
��q����'##�󽻕���p�����j�ez�냇.�O��T�i��C�-�i�Y�ggi�/����moNďdq����ȭ?=P	YU�8Ćm��a�h�K���9	4��(і<a��<�6�Rg�
O�dz*�y�X�y��	�м+�/GӬr�J��J�uf>�:�eI���)�7!�D�5�3���K�&5{>���|jr#��fv|����@SJ3�h���H����j�ʮ	��+�DJtj.�Ol�j^.��F�1)����G$g�&x�G^T���O��d�Qj�&�'̀��%$�P�~[7���t���`�r�Z����~Y�e�JGS��*r�C>�'�%Tλ3�e,sXL���*��Lac�0�@�3寬eH!U"�h��wer��wP��o���x��2#�2�����&Cv���0D/{�a{����+��J����+�A��KC��RB���5s��k?�o���XGC��{�M�43?8쵾��G�����Bι:��_N�̀2$�/O	���|��7p�B-���$5y
� �A8BFz��,7��/5�cd'8	�ny��%O���PC(c�܂�FF��������� CR�����>D������^�c=���C���e���v���a�6o}A��Ai��~u��Ӷ�ģ��|��`[��.��b�M��hƝ��WY�+b΋�s2�g.E�5V�4�O%��F8mTW�`FGO�d;��w�b�����<դm��N�M�T\�F8��؜���X%T�
U+e77t�r.Z\�^�Z��=Ďࡓ����3� �,���_3]q쿊B[wR�c����z�B{� f�!.�(l�N�	��@�\���)��E�M��F�Yb���N���(��%�������x���e���ޓ�-.|�6xL:�7�1���B���񫄭��+y�q�@OO�⺧��!Q!h������O3I�!�h��y����Q �#l��r���~ң3:���q:�z|IxjH0^l��4N��ӻ��KR�p5`������6D@�����Þ=�)��� �di*wLޓZr�5�,=���a��Q4M0v��8u��u��=)��6-��#�YF[>>���ү�5:�m�����eE��@~ȩ�p� 0从�O�9�bq
Q-?= %���t�d��F�׽T/L2��q���z{o�'�g}���K���i��*������p�JYYu|O��Jt��F���I�NgSu�������P`K�"�E��XR���1[���OG�N F�$��J���C$���U�,ez�&Os~.�Z�=h�>xo���Q$��&l�T�[ߞA�l%���tg��9d~ݔ��34�H���XH������"Y}�R僫�{���i���f��7
�y�׿��,�&v��^:��a��}����Jz��z:���ߗ#��;^]��r̷�ʝS������ڢ�0�j�bF�4�3L6��r��@Y�)a�:�x]YX���>M{�� �o�@�^�ߪ�x�dd�hV(�1,�r�q.G��·AtR(W�+�un�P��Q_w1(kC),����@~��c�`���41u$x�����,�G<�#~X\Ї�|����B�G��%Pt�w!��C�c��4v�=妍PW��K$��T�m�����!�8JJ ��t�Á��
����$��a��������Wp7��7R�<���m�:+La[�$S�f��Л�Ȏ%�Cg8�A��!�r8��qp����_�g4Ar� �d����/�4̾��md����a�!mb=ʷ�I�4����2"��q��i�Xd����˺"�鵏f������;��wa�0��$=�g��@ i�SJ�Rv{�a�%�&��b1:�6�R�������/��l0P�L�a��Su��u���&]�MwH�3ikT��fqO��sH��̚�Nrm��h�x�P�!a�0�\$��lY64�<����-G�$��~)rⷀ�m��k���Xm���O�֦ங��_���Ư��J�~��<'�CĠjX8� Nq��`��dB�p���6�[520E&R& ?�fA�R9�t��v���X�������)�:��r��c �֗:��3��L��b��i}�C�η	�lo�b�F
"���h���=�l籈��zgUCyy����=a锤N�1�����w'd��V-���,`�V�a���Ι�x[D��;�Q"�x��8����It�b7�R
n#��Y�=��L�OL���w�}۳c�H��z�}�]X҈Jލw{�ʆ�6`�D���o�N!�d� �ҩ�޷,W��F�)i���9Q�x��@?��L�8^���`7�Omq��|�t����y���]��YS��ج���, �R2�����V6��Ci<K<tǡ�0ž��)ު2���ic�p�����s	�Ymс�Ǡl���Z�N�
�M�'g'Q��3�k"� � @F^�m?����>q̳�3�yʚP�R�W'���C˄�x�I����M0��H�{XmԼ!�*��
�ބW�u���&�!�h��c�;-
�n�J��ܯ���Q<���Fq[%3�a�������n���T����*!�
��E}��{�+�"�@j(2���c��/���P��[����z�ǆ#װĺO@{.z|�x4��8W��>���C�S�"�Pĥ0́�^�q�6yX,%��%/ځ�a�B�b�����2D���"��W,�"��9@�S��G4G���r�`}���x�B�VLg�b�,K>�a��&��ܿ�[�3��N�N�����c���^A��$�q6<U}����N�Xh�5̄���m��@޿�x�Y�'hp=�o���?g->���A[f�`l�ҍ;�m���O4�Jw�?U���H��'ǅ�V��j!�3�xb̯`4ƶ�������ؘ/�w�i�CV��0;\�WSX��U��N{"�9^N� +�f �l6� -g>0��
B�,���;w�p1Y�h:����
��Lb���I³����n�Z��-l���J�ޝ��� ��ŐW޻(��j����B,x����eTڟ3_b�H��	\x�֤�H��l��1-/�	����� ���Q �BfW�C��8C�qw��RUſ�+�֦ǖw!X!{�Q�].�5F�7��#])��'�$��=T��%���g���5��%0�bZ/���%��m�K��`_D�����LQ��Kw֥|8h!��j�G����~r�z#]M���x�=���'���:¯��$/��	�����w���Po���$�����|�摟Izݾ8ZC5J�����vƣ���[�/&U6�*���� 8\�Mq2NB�a�?��T�!��9�R���G�i=��R- �0���	5�e+�S$��
��lg�3Y��]<q����O����G(�4o<?	�R:e�N���e� +�)X?To�m��H�W���~d*6���*�����]����<*�?��W��IR���C�/��u���L��.��
�nٚ�"Jw���t�G�4O�y���Î�>l��im�dӫ�)���Y������B=��9O%����dq�ޑ�y�ߞ7��-E���o���3�d�qj�"��̤����,Ӎ�� S�Ր!��D}b��F���W�r�����p���C�1����C��j�����֊?�����_��4����w�b�uz���M΢��wp���$��`5�o ��������Iu���{J�Qt22�΀�_l3�p�k "1��4������0��h��lwF��JQ���]��.���/L8��-�����V�P%�H,�=�����x�cѢ�" L��:�a�����E*����U���!G��Yfe%�~��$'�+��|1��<
Ҩ���Ri�@lS����*�"�Ý���@��m�wƓ�*ӯˢ
�O��2O����t�ɝ�k%�w�|F�3��\�	�q�e�ɚ��=��k����Ԝ��ѺW�$��yxQ�2�u�b�p�Yz�ֿ	.#�ǐ)KJ;�1(�x��T�~A��XI���ڌ�O��]�%��ʝ"1��wҺd���#N��!eC�OO�}�ε4ii��,2�[zq�)��	?P.]���G�N?�"��I�d�]0��@�a�2X���[t�I�L֝я��3@�r��Ub��wft�'�&nL�B~�6�D�P��I?O7p';�rKz�����=fe�$���z��;������9���!I�p�n�T��K�\%V%2��1K({��F���	��W�hSl����������c���ݼT/�2����F��ͫ��Q����2`�5�bvl��8���Z	��1h��"�ML���iK3=��v �+�^����geYr4v ��[�NǞ�0��xh�+�Th��g��,%o����V�E���b�q_����bd��: �=���`8D-3��wߏJ�/_�/�tB�W��΃�<��͐�k�nT�\��\Fj����� ��Y�or�8䐙P/lK��'s��=��ll0]�!ދY�E�yn �}�̊�Y@�+������Γ�ue�^��l m��ʒJ``T�J�]nI�f��ef�f��	 ���c�s��(\!�9.���QL �0�?��;�a2϶��,�;��7I�OA�d�cF�H��P�����[�nZ�7<j-|H����<�N�Ƚ�'��N��q� 5�H ���Gu,�l�lu��K�k	�	����aM��!ELzH&���#����{F��؛h��f��	�=%��}������26u�5�R&�̟̗�>�Z�.�c�1v�f.Q�� �G���N{ƖW���k6��C�QR���T�Q|-���N���m���%s�;D�㄂��z�\���6���6�>��ޓ��j̟l|��E?�������AC�Ê�f�c̸����'�-�������פ��Y��4lɯV�:r�V�ѳ^�DB)H��r�qzo7F��66d�0�S|�����%T�
����^�����Y���c�R$Dy.%�z�yu��7��˾��4����uj`M�����n�>榛S�e^2��],��NJ�����en ,��)W�8�(��"��q��(	� ]��W�wR��+�Tj$V�+�\�F"�����l�?i12�=h9֙��Vk�ގ��k9n4u�OE�u	UD�}�B�>A�g4\��b�����B�9�x&��&�f[�wʾ�xl�$1q��s�v��{��X)�--a��xQ����s��/!H�9�nw5K�,�����T���\�NzF9 �������;s��0������U4��^]�& 	�l�}�TX��Y�=�W|��nu���+�Yv�[v�/Z��(&|hh80ִ�!�Z����H)eͽ�>���u{희H5e7�$֠S��B-Fhw;��X����򯨴Q��'�!<0�5��&�f3U���n���o;o׷�b���)��ډ�J�{y(S}jD�+u)��޳���d��W ��,*g�Z��C.��'�w�8���УZ��Q���__��&Af�� �9���]�(�H���yd�/M8?���nl��:��9�,��^U���F<}hb�p�n���1�aϴ[|�ţ�԰��.�H� �����