��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$Rx�y�<��wA�*;�x���@�̦�W�X�fa�M-$u����n~�%���P�$��W��kYَ���P7�?UMfT��q�6�U��k�>����~�\N�(�����X�e���/6U|)�X2pF�]$h���d.���9E��WG��L�X"]�Ad����ľS���8od����e�GT?y	7�������ݵ�^��R�q^]�鍦�����s�ae���h��L��P_���ާ��YЭF���'\��68�b�[����w8�[X��V�F�0͘3����q諵�uW� �h�u\V�?@��_6G�_�*�G���B�絉�f������[�G��U&�����~�F��AׯK1�`c��[<��FY���4I� �#�G��x[X�=�Q1��`��R>(�w����R�O�?����7�,(�H\�#h(W�EH=�������yq��Ѿ��aF����:�U~m<|��.��0=�P/���4ǆ���T(���%Y�����3n�&d��֑��R�F?�;.!oiOZ���c'-2��.q��m�s��n�#�M;[��4�;����"�$�O�ЗǅKq�"�	�>ȲJsb�u�F�u@�({�X�\���z��'�űJ�҅Z4v�+�2�V�Ľu��kyF�t��#��U��H��t׺�|�a����%h�>W:b9oK	Sp�_�(�)�40LQ�:��wu�Ƚ�G�w%j��N-�a��J*K5�o�ٲ*T�0��+vƘu��(q�DkS�+d��S"5j�8��9�G�?�-���R���C�d�딂-�(.�y2ADq�_9�k宕���]Q�I�\u~,!�8JN�b�}5&5�R�H0@�3�"����r�!C�H#
�&H�J���=����d�d!u b�����-<Lo�.VU��vD8�5#�7��U<ؤ�?2T�~����P�:}�^z��f}�RH�{�t��� >8wv�_��^�,;e�U�\L\���l���$�(�ܹ�J�B.`\7R�q6W/�����<vi�P�l>%3�d���3�}����7�G��w2����I]���K��7L�6I��f�'K�/P���F�yX�~�2c�<l�)9�[��ŒS{ȤK��
H��d��m�� ���Nn�O��=➆���7��t�no�P»�w�d�j,?���h�
�	n��jx��\����`�����䊳C'�@J�d(�c��?��@ߗ=�hl�j���[�~�V��8\�6��^�=��"1)��,�A�6��F{x���T))/���frv&y�9ǒߊ|Vv���l^ L��˝>D�:OϱE%����UϜ��O "����q�֠�q�����݌��N���C����HB	�/�q���Y-�|�HC�y�t���Fߴ%:.�r5�a;r�����oO����z��naȤ#���6����1Dߊ���Nk��.�I��>�<�9��	�"�Q���UK[ ���t�-�<g�Q��N��엑��\4���B��A�ܷ��y��9Ls��z�7��^�qP��Q��#�X�	/��m�ūV�K₡>
َv,��ӯL�8KMʋ,/�E?�=0�у�m��u�4�D����φ�g��5��t���va$��[��|z]���)��F����GnL3�W�M�~�ȵ迿��VL�x{��u9g�h ��掫�/(Z�pQ�pd���<�8� �����nm�@���9��O9ȉ{͆��nDrś!R�ıg�0ld<���w��զr����E^��� �ɯr��<��#�)�.��2�B��\�^(f�e�k��?a�hx5Z�`hhf7=m�ϖ��'���&������J����('S��R'�g]��C�L�9���^�=�/k�2�P<��d�؛�FO���p2�ҹ��N����D�����Ʊ��=�2-g�Ӣ
�6��r�{Qy�=�9���t�X�;��q����L�qa��R�6�wF ��_䷓�$4#��:5�|�hj�Ѡ���� G#��vD������{��{j�d�d�fyW*؏{uA55_m��Xfa���k�.5�:�$���U|���l𪶹r4OmR��<�����ހ��>B�VF�)�5�9�UԦ���NG`���1V�N�yBK�Gfk������x	W�|�-�Uf�W��񙻢�Q*���ŧu�����ȡ�ץo��Mn��5ڹ�]Y}�"[q�&��N���e_^��JHw����7,#�T*{�ܞ_20������S�f����9d`�a.��{:3	ԓC��ȋ���X�lK��=)0tܕ.��z�$l��or[�G_ﾍ���(9�(!�a$Qb�Z8��k�V)n��.ً���Z�����'4����Nq)��Yў��h��?���v�}Ax������yE��-R�j�����"�'ɌA�G'���-)��Y��X�=�GrѼL�����t��hW���P+0aP��qQ	#䪂as1�x�h��_;�DR-a��Ҙ�c�b8�i�JT���(ԩ:����P����n`vO{yUD"�p��&��V��<� ߿�b0($�c���(�ƈ��I�%\��%)�j���Q�1I�$nV����L�������Z'ұ�յW[�}	�w�G����CB��L\��}V�g�����[��J��U�+5N��CNe����)�Y9�'�TD{X���������+�*J���}/������a���a�f�O9��;�͠.����ŵ�֌�OG.�w5�`cuOR�g��?�r��y��E�pԨ�V�E�m9��=-�{���e?���cy�ñ�4ˋ�'r����`��nwGp�c�� u��8���H||wy��<��Q��wD�`��

��xQ!`�+S�y�Հf�h��񬯢��vRQ�q��AS�)ʳ�[���5_���Y>������؍ӈ��|[��#u��KD��|��Swt�_�3���`�2&�CU�m9i۰���ъ�<�ț�T+3��=P�Ъ9��'pk��(g�P�G%�\�MS����Íg	���<�>��b�8,���V�+��J�z��W㹷���6`@��"��~�DǦ�?_�����R��'n��2Tf(8�1���"�2�V���G;pD��'FЊ�1{�g���c$��c�.��..�S���!�5�V����(�+ϐ�6�F�/��!0w}� �5��1Љ^�A)��n��u�L9T��κۋ�u�
X&���'��w�f%�Ĥ�q�Ń=�5=jR�p�R/��~��1�ŕܰy����5�$�f*
QyZ+Q.^k����;��|g��������M�ٖ7��79t~O�O\����gK���,��r�Y#�!T�;�R���a�_����9��� [:�
���<�՟N�����T��p<�X@�{�n7�~��o�`e��~�C���+��	���&@|�2��H�b�Y��DA�'�h���``�tC������~2 a�o#	�����-���f�!�S�i�(K<C:����z��@�G�@Dʆ	o��%�Z�9�.>�݂O�)���QgB��W�zӎ{�tj:�(�M���n�6P � �&C��-vM����p7�KT
�k�ϫ��B*G�#|���j��d" ��mԙ=Z�T9§(�6[�zl��{`@���0�4{�fP�uYבAJ��� �ʷt�jq���P�W�y���C#(�Q�L��MB����F�YZ�z~�p��P�&q	�p��7�t�kS2Fhh�
<g��'qlǎoIJEH�p��Ƒ��jF����t	�����f��j.����W�Tyon�q�#� u2�[
�l�*W�ksl떫����kͽáV v�+Mf�P�Ei���GV�q�De,��J���"=����	4�;�A{Ŋ�Z�ͬW ���r6��_�!���a<_�;6�Cޒ�-� NPF�4fV�-4�\���^ƴ#BCr����+��2��fj/�M�s���q���ͳc�zp�2pBD��!�<~�u��2}������e���$��Y86`Q@ _��e�Grm{�T?�-��G���P2g)	���z�"oq�4ۮ�6�?h��7���K�Z~�e([��_������:��d��`�Jڤ��*WJ\83B���!b�����ƞ�d�:t���{��x�z#�e��\:s�Z�n�(���U��洇����>��+F�m���Y��R�$�;�I`zCQT����mg�fe���ZpU��",I�*����;q綤:�\�0֫�-��s�HtZMC�]�I )�������0�i��!�v���-�Q�,.숍\, ���G����x�sy���=C���u7nn&�i��I?�@����l�����:e��?Z����|��d�J�eA�(�/�#�+���e���hl`�7Z����eoJ��H���������fQ�/2�����YN��	�Ko
ߊ ���~���ތ�\���w�0^_��-�bK��<�'�u4L�V����Q��FK'-�EK^��W5�O令��~4��8>+�<����3�3����j��<B�nsY`X��#^�P��J,Ae�U.��
����PG�x��HX�j�nZ݅~��Բ:&2��A	�^�|�;���p����'�{kgc�[��@C���$��~a�.b8���!x���˹��dǫ$��1E�W�����Z���}�_��yű�����4�jw�.�Xv���Z�3�C�y�ؙ̇N��&tz��������S�����W:ɩ��3�n�
BC�1�uŃ/@N��$��<~p�`ut&�>"j'�=�[7�k�]�a���hަQ��W<��!��tp�h��1��e��r��/�.5R�
�����9���Óﲘ��YET�/�fco��Cs&�Pb%4f�l��逭�"�R}�5>��� � �!�4�������bp��R���6�oI!�� ki뛖͠�DӁ*�n����Ta��Q�����Hf��$�/��L^��Z ��2��G|�Ѫ�ZG�u
V�|�V�d;	���=�VvXgG�vW��l,SA�� �򺪡cg�`�U��ڹ]b�٧|V�t~�wz�+�@F2��J�**Ċ#u��h	Q�,��hAXY�#X`a�.�EE�(-��7�i��fH�ZX��?ş�; sF�b!�ʥ	��'}P8�ǿ	��)�7��h�b|��B�V���q뢇0���:�����p),dQ�5��\gyF���x�+����*&q2�C�Wg��;O�z�͈a��~2��I��� �5�,@ʓdd!�V�I<�7ML�)���B�+�e���9�p5�lϷ NV"ƃR�˵sK�^=S��7��Z9y�Ȁ��n��P���ʄ�z�8��Yz�� �jkgt��m��d�',�2���� �)u�7��?x�@�		�Æb8�ɢ@'P�89����X;��[�ߖ��[i��R���&W��W0��!������=���ۤ���p��~�,��HW�ԝ_�?�
JJ�s�.3�1Gێ(Ԗ�;�k]S�O2��8��;�PUN+�U3J��T尿�"�L�{��1���
a�����9�"#�#�~>k���ع��8̫��r�����Q��t1#.�VD_*2��������O��9��	ZfO �z\���F��1��R���4�����\�&!��4�ORއ���n�Y`�t>������v�3g<��^���ewI�ŚW���0C�A�ӐW�`�+�%52��@�	�_�(���������}֠>z\�|vgb�ʽp��9u��K�gY}p隍���O��u�h�*1O�3�	��M?����*��]|W~��P��1��(&ά��6Xt]7!�G����KP�)F�l��Y1���^�z�� �`z��qoI�k����_�M��~o1��&��=u(k�;��"/��m��L6/�ioy]	|�	yzr1�H�L[��0\Jx[�� o�]Y����	�-�G����ͪxs����}�ڱ�b�٣PڻicC}Ԕ�G�
/���-❘'�%@ֶT!�wH��͑s=�P��z@��Q�%^��"j�=&���T,f���uS��5��\Bш-إL��|���m�|fU�TsLS�jԲ�J����fi�:V*bG��?��p�ф�^nZD����|�Zޏ1!��\�!����T�Hh[v����G#Q���4!m+�~��d�7��T^�T�,�6�t}�wC�`'�J��z=�)Fs��l�73Y
yZ�$ s2�*�6�i.\�������߭Gap��N>[�^x�tP��V�8� �K�#��ֈ���F���f�s'/K����iNk��qN�o�� Ֆ��^�fs�"�!B��2L�)E�[���]\Ѕ�]�A�rY�x�������ӳG&k�.���}��JZ�!u�D|�]�D�`*���ᤓ����ʋ�N�rQy#�5Ϲ�ԃ_p�^���>l�!��R��ବ�B׫����󐔁2~E�����'��&��W�P��p�m�6j_J>��$���A��,XI�|��<Eef��$}Yov��M륧jN9��e�~�K�@2`�`X����Wu`؎���$�J6!�D�*�в���=�.�I�q֐�X������,�٤��͞�[-�����Z�7�Wy�c:'4�𑇑��9��p�>�4:X��l'�9�b?7%S_b<�r/�H}����m�Ȇ
E����*>�Agn�VL���A��5l�{M�@������f޴�.\t�~����C�񒳙��Ͽ='�l=E}��?uh⓪�@fn�S�%��;�up)�ۉm�k�M�^�BG�cr#��U@���ņ����^e��&�B��k˄��8�A?��wO5���@��:p6��}�r�C|M
��L���l���F�	��Ġ��߬��c�ƺ쾤�<l ��z�Cp5])�1��Lh�C����m��'��媽"i�w�>[(��W��R'�T��i���*#���p�e�� �����;C�j�_w�5��r{f��b����F������<\g�I���+��xax2|���m�~+��ʖ'�����!ĥ� ��:܄��\>���+�J�hQ��¶+�[�y�F���b
��?W�9<n���M�'�/�����9�T�$!:�Ey�&СƝ�����F����p�O�e�7捋k���͎Q$���<W�9�~k7��j��iQWi�mϣ	܊�#�<��L�8�	�Mڿ<K/����{w�̞/R��ȓ��V��|�e!ǟ^�����L�7�襙|�Q�OS�*M�i#��Q��8�J����P�<�\���d�gF���xC�����	�P��8���9��X ^�>, �����=2ݷ���l7�90D<�����B�$��^]�;j�P���OX��+}xŹLFA�޳�����i)�-W~;��F�����\�Q7�Y�r#���?�:������0�u�ә�
��d>���,��C�w%��r;�4����G���{jr���P/"v��*�XpG/��/Ռ�����~�?��x�<�C�.[�a�z��E�߼_�b�d׭��n��4��5σ������@[��9g��C:pM>��e|Ҳ�-�:��&�oK���(�\��ϷO��KN��sz�!έ��5j[���b-��XGyO�C�����P�X.�:�ڢ�� �Y�[���MP�\�%Rh�:��=�C�SN���CҴI�|�if�	.)Es�볃��A���$?k���Q '��L��@?m��xS�a���N�ߥ>��[���cK��fh<)	��)�ozC֓��q�I��,���1B�e�h7t��R�NV�Ln�+-�i�$��?�v"2IA������i��c���-_Z����e߭[��%��l_�L�����#���?d��O �m��k���}Z(�i;���	�+-0����Ơ˪VR̷fp���ur�Y�̶4"`cCP�:0�=��nC2�J��]=��D�칍%�_F��(�!q�6�g%�G�(6Mk�FA�
�Dꀭ;U;�rq�c��4`�og-F�La���&YW�����$<�s������k�5$�7�����Ԙf����ǀ�Cϓ/^Q�>�VC�T��H�ӟ��[��d�'�׿G=���U�>@3E���l��[uUX��&?WX��Ƕj5"I�����I��[%�2��RU�t���Cܰm�k	��٩��{����(u>�2�-��xb����wɮ�X�(��4OcŐ�p�4@GS
b��d&}��&a��-ƚ|,����F4?�T������창i3>�#�z�/�e��X�� Ҋ4B_��5�%Ec�k�'�8^��.H�'�e���z]b�(o��l�Ⱥ��A+�0��ܿu��P@1��+��2���
���ɨ��S݄G@�Q�7��b�M��J�p'Ur$�;�P �]������pK�����8���!��Lyq�G*���Z�{&K�>�/������0��y`����p��j����D�PC����q��ԯ�y?�r�nJ/��Ez������T%��n�k1�h0c��	�vP��,��K�4uH���B(�M�~�*��$ �2Nx��.�aK�0��M�W|����j�ut�����wVƳ�[Jyɔ
/�	��z$'�/���;c(�u;Ӹ$���y�z�9NXc�/���W�e\[��i^�c��{���+�F�́h&����'��O���Tz�ꤺ�5�QLX�C:�m��;���6ou̗�>
����:G<i4#�L��y'�\����J���ki�	8vpw�si�C!���g3��R轜�BsC�#������MzP�qRp�Ӏ�Y���.K���̇m��\�:P
�]!��et�[�u}��7Bi�+�d$�:}4�8l������,<���6�Z��j���\썋UH��=�����z�\�ͺ���+[P�noZ�FfB������B,4B�"��5C��J:HL_�1���$B�j�ަq{"���t�7�NqAXzE�,�$����ɛ;���~��
�����K�tK�i��Ma����ȶ#�d�I�H0)�Ձ�#��=���ef�p�J�;F�m�=�|9>����,�%����e�B�H��^� �?��L�eM��x5 �:".Ɋ>����&u�#��Wv��n���I��N&��<����\\qٖdf������&�� ��-�Åh����';tYL�>�
9Or��W�;�A=#��0�H�PrX�f��ш.,}R�j��Yl ��Q%�����k{8K��9����a��\2�)V&���e�u�9-����<������J�.�$6�pR�}�R��'L%U��[��i�s��p�jI+���R	���N�,�TqG ����� L<�T��NK|��$G�V�>Q_a����6����0٩4�_[ze��֝��, V` lɤBr�rc��|a�����k�{Wl�/O�l��XrMG˩]�F4�~�2E0���+?���F��Aя������ٷ��L��`eY2�ZtUG�ѕ�q��^$�@��ǫ�CB���K'ih��2���4{���2��!6�o�lavf��h�#+��iq9Cy�~�HwP��/�zٴ�W\��j?�%�h�7�8�T�4"y���O���dK��9��U�@�Y��ݝ@(�:\g��,Y��
!�yG�=�@�S�@����/��$w�����uB9�����G�1�v��b�e�:&h&���+�'�PlZ��9P�x��L�v~���S�Т�]~��_3��6��7���e:���^���D�˙�~;?�5����l]�'M�T�g�!(B)�/+\��3�0��H��|lq*s���)�x�a=tr]�d]kj�y��B��>q�!����w4���z����ė��(A]*�>YHh�ܠ�(���!��rt���-?��PQ��R���Y�4�(���2�/��KkZ�x�k���y��,��Q1���gW�OH���(�2{�U1�����\7d�!����X��r 6b�ބƁzs�-o�=
juq@�C3B�G/�s�@����,���1�I�sav/�	b�нA�mlr�O�s.]��B��U��〰񺊙y).���QG��٠�$na���1��ؾ$D,��w���F���������	�����8y��10�)�t�V�*R���T���A
=��]vC
��c�)H�>�_��g���q��zWӛpɓ-�\uL3'���#5���^�]�w�F �!:��{^<�T?��\��R��lv�{S�\��*���x7��u=��1����J���� ��c�_��~���
-\�f�J;>��P��8t��!�C������+[�c�s9Dר�J	7�Q紦HGp�r�#������:�ڀ����7թ� �G�P���d����2{�E�[�"��u}MLoq`VJ�դ/�:+������E�~�h�+-
��Ɏ&w�aY�t�	�̛e#NM���w��𽈓���ۚ���'�P�Ow>ٷ�Ԅ��$Kж�EӼة��bp�T�|���>����p�^��g�+�1 ΔFX����8��^�Q��Tk��S�J4χ��0�k<��]$�+�չ�Jfx�|Twq���9A�7~��5���.�|_��>�7x�
�G��ŵ�;t�a?�q-�.Q�Im�DPգ�C�L�������8�J㙹�Ҳ�p���K�S�e�����p��a���;�rB>��Z�$<�f�aˌآ��a�ܥQ
��j¥���T>7���<T|����q迅�������y��2��������!C���M��Wݼ�Qt#s���>�w��Dp�F}���?N]Ƃ��[���ſ�-W�/a�vf;�Aj�g�JӘE�*|������|o���B�[�^>J�OSC��kew�o��g@훤���}�P���C}�F�+w.��X���B/�a:ei���B!p��-�Y������%i�~Aܚ/�|V�U�55ͧ�!c��M�-�tk?�LX��YA{�MA�!K��AOY
�����oK���-6ҕk�_p0	�
��&�gc $$C���2 0=�O鹧�QQ�
��o��cX�)G��H�v+߻�n�fj)3�v-��<A� Q��_p/#����^��Ɔ��M�dW<y(�q��3����O9�k4����f����=-������+W�,�A���S}��4|����J5�VU$�(�&=<�|���eݱ� �E�D�x*�Az��5�ڍ�����&�'��;̯�x�yΚ��D��{D�ي��$�pnx�(�$�D�$Y�$#y^h��0��<�t�(t�-Ir�����*f�|�Aъ D�>�ea;��?�p������#�]k'��	�d滜@n��*����5�c��E�!���0��pX�T�\�Z(T��N�����C����Io
B�Ǝk�8.�!I�IY��~,w�]�ţ\��=U_4?9<#zl�������孟��9
�zb@ �!l���U'�6~�y�L��{;��mr��+���:��+�g��~�˽�����ȷ�q��g�{��cx����(��)�k_#���i�=K}������{{�l�V��?&����^�1�#O�J  R�d��{~)�Cz���y �Mg�[&����81M�H
1���BDR�K\������g-C9�-J!?�����*3lp�A'J��M�V.�z��y���0����BW�#�W�xj	Z�@���7�g�
u��R/ͫ��ɬ
��3�C���� ���6�A�|7����;�)�v��-`�u1�ǉZ��	Si�W?_R!���C�d����+�h.�09�G����xC���hd����ax<��H^�}/�A�R� ���r�Y�����4����yL�i�B��v6�s���g`�ǳ5��7�~֔mT[�+ �{�� ha���ڒ�a �ģ�^Tޗ>��"Kq�@ScZz�z�v�O�9�1?�a瘰xHҥ�q�@�4��O���
ruK ы"J��~\;g͙Zk2Y8P���t\(P�bc6�Uc��47@O��������p�ӑr1��g ��wa:��9k$CPr��`�D�8�8b��f۔��~�ݲ%��)��G'�a%����Q���
���x�M%�����L ��������{L���?�e����$�Y+�+A��0�Y�I�o�*�J�aYz
r�z�����T0�\.ʘ}I���.��6���hDK�ҷa�Y4���'����7Pk���I��1���.Kcn
��)������cp)$���1����2���/c���C;v~�e�&�Z~���t_��"����WT���(�n�5��΍��O�Q���W�G~�7�6I���'�
p�;��e���<j��gRcd$`��۲\GGb�H�1uz5��OoɄ���ԡ2s��٨���$�Wa��ԭ�_v��"π�[�c6���#o�5%Ih����-��J�Fz���#��_��j�U�ט�ւ��y�D��qK�+�����|�L|��_o������f��w/�1�q����b5a��O�Ő1�<�u�9���'t)�����Cˌ�t ��Ȱ+>NyO�T%�r;,���w#;�۠X��vN�r�e�Y�@J�#]�D�p�-�. �3�T�/r6{�Zu���u"�}TR��ے�gK0P;]β���H����c��U61_�E���Z���]�@"��wD��4��2K��;����������F2^���y�w멊���Nt6sw~H��'0��~�.�R��uRM���(�k��H'����	�۹��|��Ķ�s��5Y��2#T��p�D	���r�kg�w�;���,�&z��"EFkM�##�m7n�^i��u�_Ƅ2ɪsؿ
S�#�����8	?Bk�t�<j�vj�$(�c<�u�Y�HD���]}�92�`;�&�m;vD"�t耦����8��c�(by�Ab+t��h8���D��:��u*,��5��N��,f o�a��i��Tr��{N�/��On3$�~�?Y"1�/^Ư��a;�bO��;{T%:Ʊ/]�l1�؂�JS�`�RF(��2�u���J��ґ��L��ͧeD�����^H?������C�q�0��k�|�ޥ��,�Yt�G_��u;�P ���X:��рA��K	Gf�G8��Md�f�t}3�~�j*����h.�\L*�{]M��"A���ARH��<h5�|���W7� �1�\�ԟ-�JA=���-�����а�;f����u����D�q���иZ�)�
g	�%�q=y�"�o��[�����6A5a���#��� m��vԬ��I�4�*�0�8:�jE߀V=����Y��  �3 �}��1�C�	%ߺ�ɂ�YLA߳e���	��o
+b�)b���7pSt����2Ԫ�����=@�	�����/�$o���(��<@Z��2D�m��w�u��Ӷ�>�3Ro�?��z�zP#���x��Yo�P���������#\�2�yy�\H���ӆ�,I��� 84;o�[�!��9��k� �iM����6ô���#�>2��aʹS��a�^�)��!9�U�.�{�sIPT��v�߮��(�^�K�J�F>�݅�İk,�.�M��N0�xUz2�*�g����D5���Q��T�0
.cS��;�1��F&՗�8�_��oO�S���(�tp������ ���|e}�s���������^r�O���g����s3�8)�6:q�M
yD�4Zz�$`"ǥ��'b�R�p�hk�q�f�/��0���������z�j9 Jm@��Q:CY
�/b�ҁN-��
W��d�Y�"ݍ�]�SSS�?<�}�w�ef�=�x��\���h�;UR(�d�J%�'��L�ʭ�i��%�<�w��)����T8R,y�`�^�0�4=7⿦.5FdJ�H";��|fI8Ax�rQ2
)�����0bx8�����rX���l��Q�x�E!us��S/��-��q+Ԭ;�j��Kފ�@=�͜?7��p�����k��y���LZ倆��Dm� C����z/'��%�k�;<�,�(���uk��%���w*����>�D0��':@�����;�>���,�i#v�s�����ߞ������RpZYcn�g�J�b>�����U�h��;�f�X\?E�X�k�'��}�Y��,�;�8���23�w�n�9�e%�͚�I�����#��q�@�ϩm=�{wa5�����a0G3�Hn��-@p��6 ")M8hPӔ��:� ���ģ08o�ynm`	/=�U(6j ��o�H���nC)�޻uzf�[7�,�a0���Hym?}eYL!F�؍���u�����e�e��s����q������*".h��l��
���$)���Gb:�q�&\��.`�8t��FrH�;����1�/���.)?U��2� Uuq�$���|g�/E?P�%��v��ɥy%�%.�	����&Rߍ�g��$!�Oa���u4����7)�pr�4�1�o��9������ۍ�4ʘ7ԓ���z6�q?'Yg��i��(2���a}����uK?�3�r��vo�^deX}��&��{T�x1�GA��s�a�)s��Ж� ��
*�Cp����S�{�O��#����r%`B�0�}�+R����#\�$����_�Zt��2`��Fz�G̭H���-�Ϳ䣲4�(�8�"�VOu #��ZjE@�վM�֐�$��W<���9ы�"j&%e�{�LZZ2K�:���z(�Y]���X��� �ۼ��?K��:=��}��HУm���Qi~�"n�[�~�K��|�;^o�ib��ѹr0��r]�t:�`C��2�{�U����d�5��h�A����M�y�n�Փ�m�9�),}\X)g-&=Wv��_8p�6?v���C�Vš8Fw~��)�~�4�ޱ���k?��-s�X�:�՗�ӣ�v�-��ڐo�;{z_g���G�-*v�YcRƽ�:W�3�����{7@��\i��e~��ZZ��|D��Zpj�?�ϸ��Ӝ
�b(�̙���bMm���w7}G�>�#����[k,]�*1���[��E�-N[�r�����\P���Z�`���#���n��(���U�"<���&���J����&3��I�Id�>��ڦH�T�O�~���no�udЂ�F�mv'��Ѽ�fa���r?؞����>J�_S�]ǃm�$��G�M�4-��#�6���4S&]Tl_\{�~��8,��7z|7�\�d�\=�#��Q˽�c
ca[p����m2��Z<�@�+���IJ (�P4��*C�<E�bd^����:�'�"��vk�eq����0����0�xo-z}C����<]��!���!{��"���	dS �F>k��Cʕ�?&-�#:�����67�:��m�[|��E�KǢ��.�U�;�:�I,hϧ�}�u��sy	��������D7�M���]ʼ�2B�Ĳ�'o�3K�r��pb��K*	˾݇�綜0Xc'�����W��4)��W�q���3/�K�-7>y�Im=왃��@�|�[�x�&{_��oaH"�_�.C�|欧'f��X�g���d����������ln6�ރ��D�i(�k ��ɠWv<L!mo��*�\"!] ��3��<�R�>`� ��N��KǻLj�T��O%Zٵ�AEX���:�Y��֌�b��Q���m�,�/�Ս�f,ҳ�s�rٴq�5Ê���M�K�]kX�F�XF�	��^b�q`��ve�h����OX?]9LԾ�v�������o�9��'���ܗڸB{+�>�au�"rgRGU�q��h�l:�__Nj���D^"Du��`q���.5�bه��rLTJ��!��K��Y=�1e���'�֥۰N���t#*uP3/Έ�\�	�T������� (�Nc�*��r>k8O`]&�Ӿs��3�9���^x���:��)��%Yʵȡ��;ιC���F���g�X/�$�
��x�wS�T����;��>���`��3)p��d��(-o+��"��e�<�E���x}��B�_��d��2�����"x��i���k`L^���,�!�N7�Q��G��8o����~U#�D��?��>��ao�t�(�\��VȆ|��>��0<���$��Z�F��V��ϐ�� p�G���tP������YE2���w�~C�� }K3�7�7��%�Ɛ��^���:Ȼ/Bl	BZ��m�*�Ә>՞Kf�t߼8f�׭{�"-@�K�jr�L[�l��>��5�q�|�Wt$�U6�������~�7$%��#|���mrx�����@{��U�vH�i1l��a��C�v� Ow�}��QW��C�CC��KfFo�Ȋ;��-ܞ67����;�L��p�}9r��v0{�Jr���$D�WU��E����V,�X�޽Yu�V�|�1LpK�]z�.��p?��������]$ǵ�����k	"Hr�6nq`_���է������s�p-���������@a�x��^�ȵ7�{��R�`@�}�r/8^.�C���8�C��]�H	�F�kiA\A�<����&Z��h�P9�m*МK�׏�6��RS�ӕ��b��+��Z=�tEU gl�o�,uw�NL���o��j�>�DU�aQ���P���ƅ�埶�T�{<rR�ݒ���;x0,������Ƈ���#����y�mr��e!D���I����O��p�x�����,��$?�i̱�T\Ĩ�_%[(&�n���L5p�zL rH�����Uw�-%Y/�ҮVc�JYmCP�;�А	ve�؝:ÿk��|�'>� .��PPQ�vT�V2�n�c�B�f�Ƹ9M	�8��N@��A-L�1i��y�IX��O��˜.�����,���P��N������ҀrQ	%N��-����BԴ"��\�2Ky��� *@`0��]F�5 e+x}�P�[�ѣ��z����/~�F���"I�$"vE�D���(���V�}�CJ>!8�w��I�W4F���@�mwJi��K�lg��~qu�o�X}��nNL�I�
���J8� ��7C�oV�>�����I��.�9�u�`<p�w� dI������^8?��4�e�������@��{�[���H�n��ǣ�ڷW/m!XC��8��6�]i]5�AҮ���%�4J �[�'����$yVkNm)4_�r�����!�T�!��f���x���~2��%Y�8���T��X��"A|���(Yrϝ%�)�9���%�I�5w'����A�qg��.q�+ �(�?�KG��{9����J��z5�xc�/)���G��Z���)��q\��1�"�'�'M?;7)SI*:1�ᣭ�*U�Hڂ�2go����ٳS�z�M>�S��2��O������p�����90F\H3�a�"��,F`*-�`�(C�YY�@��$"b0�9?bZ�{� k:�����xuy@�z��A2$�b=�qV!�g�3�$y^����%&�uIv��A��oT�D<CIG�`]v��@^#}{Jt�w���Q?>�D��B�lKY�
7T��i��b$ˤ���0���jqt���}fM�u�,��ĵ�wKH׊�	(՟s�z�#0��/Sf���3���F$��X�"	uT��p���D,P˕���,�zkxէ� ���y� /�Y)�F�����cߓ���0�ʤ�L���ղ��l�=�e��H���!y>v�Q�Zg>G��Vr�yUڰ_��݃��G8�8ȗ����F�<rA�j�H?�L�bpP��6�����b�T�!r��o��<��b�W��&����H��-��t��\�!�<�5�r���r�c�[[�ф�BBݳʏ�����)�؋gڻ�QI}o�s��A�PH2�Աq]�	$P�P�9/b�,^�F�dCEZ��|eN&e���,=���,�{���g��N��ӫw�C� JJ��_��k70�Js��H�/m���7�<����4�>Y�r[���=�k?~�p����0h����u����i;L����Q�n�h4��2�P,B�e1^M�v֧^�O�"�� ?$y5���9���z���Q�ь���V�B�S��R�J_�:�;�3�O<���}]O���jb��@Z+��� �;-�WhA�@{-R:(Bm�=�.A�M�R�I��� {DoB��t'�Qb�b_Ơ�����v���O��'��!i�ɇ��}��&���t4�DL���ka8�qk��)�c��T�-�A���X�BZ��>T����Nl�u������z=VA6�W�'j�q��-��0�@��n8�G�|�(�GOj��Ģ�i��̨��VY�|\�ŉ<�t/���洄u-��	�ث�BE���=LAY��(�qz{)?�R-����M��2���q*���*�	�/�>�ZJ���1G�2B�l��=Y������>l���&��`~��v�a���x�{��#��oK��g����5��V�(����G�{�ny>���ctu��	�����,���9F@�~���ݐ����R�!��,-~���PN#�s�hzZ$:}�92S?�s"b|[�a�0��4�GOU���]�?�!���?��EgC0�/郋��KA���9�t�x�_R����$��k�즪[7���u���H詍"����[ɖ�>�,���������@�ⰷ+�2��5qk�$I&����|��H 9}�su�"��d��w��k|"E!n�>/�
�[p͋�ЖV�	c*���{H#{�X��~ƽ)- Ǣ`��>w�m��D*��^���)��>���>�)�v�s�L���7���r}��E�:G���2��,z�v����6���`�9,bz�N��3"p<DH羳����ŇSs�)�cqA�ӷ���	H���ɀ]1z�gb�s!Cl=Ơ��Tn�H�[�Q����ʂ��+�3����y�V v��l����|�:��.��m���<�|�
����^P߆��8,�����m0;dR���x�=���+F�}E��	��h���1��� i���%�6Ų�1�N��5�����%�i�c@��?6�K �D��,'�(h��E�U���V�{=�OPΟ����(�;�Z�Z��5��@Pw��^����N��N |�+�!��fBt�9��܄�m��hQg�+Ȓ)��MH��o�^�_O,��^��+t�Yn�k�Ix�%�xk���6�>�[]���WM]!r����j�#B�3�}�ÀE
�}5�� �ȴj5=;3X��ѯ´���À�l=]!��I	\9��a5�=�)����04�U���j���Ux+�w$�6��%��pt�0-��d&����$�>�c��������;��T��d��q�mn0����RM���\٢����[4�>/QD���znO�e��{U���8gX.��������^�KV�^E�����M���[!�Oz5t;�q���1@�n�qX3J���v�z=���)Z@�J��f��jCk�4�cq��ދ�>~�i7�l���u%7���U��D�\�~��:�ݴ���>g���M�a]3�VP���	�p{��˂��T�d�����8Ƚp! 'I�/gH�a��<?�o�P�i�]�
`"�{��.�|�=`dq�?&���}w���#M�|kn�m�k�,�(���.ԝ�Ÿ������C+.e��x ��P-=��|C>�-��a��NC�K�q?�����V�2����<�'��Z^�����t ݈T�FfR��J&���P�)0����O�5vʩLS��xt�����HAn�2k�i��С�D�iH�ɂ��QG�g�?ɏ�z%�s��g���~Y�8b«���y����F�� ��;xҜ��;>պ�)�@Z��������<�p����B�߰�y�ט��Ƨ�Z �d��2���`YD0K�p�O�p�����R�R7���V瓬�\�����$A-�iĸڐ[1��d�1=8J�V�K�ԇ�h�����G@��B:|9D�u�`�X��KT��(#�(�I��m��3A����S��Xj����������85h���&7Ux$U����/-x���a�F~�����cHyIpC����w�suZ�D����B�����y�M(��ղ�6*|��F�B�/�i�M�d:��c�r	%(��s{{cōE�� ��>*M��D�� t�p5V*��׌���U����M/)���̗S���x�'�iQ؝x��￝_�'x���.�D�F8s��h��P+5�_tO���F�Q��2�F�CU���r��}HbQ��
�����-m�	d��y;r��g�T�b,�**ʏݕ[��!��!v�5�V [:]-qb��[}%b��tܹ��g�?ɟ��>���3P�gb|���}��O��*��^Eon�m�l�	8�����?��0��0��yg��[h�=r���rF�Rݕf���#�A}4���E���/~"`�v������ē�� �˗}�,�oK��p��i��y���n�GP��2:�=>e��;������lk����@���J�G�]���u���&�4��o�s��S_3�H�2�jwh�1D9�}���Tԇ�k�Y���`we�(���P�Lz�-F\΍�f�TS��`��$D��SXqm9�cj� +��0l��_�PZ��Ko�-��a���j�;����$�ɽ��4�Wt��.~5y����t|�>$�3$9��C3}O��_�Pb�Br-�kd�H�q�Y�%�h� �����S�	�o�.�M�gD� ƍ����ԏ^������X!����X�h�VgK�wo��b�B\��5.����I}UG�4��\2q�2�k��~8@����sw�LB‬^���{]^� o�=�� ���Ε�|K�k?�F?kɄ�:�،o��dc|���#K�t�cИ�����_c|!���z��	�����k�Y+w�%  x�\]��ʲ���� �vT�p*�5,�c-x�wK�]�f�KR��I` ��%Ó(��9n�E![!&@T����*���3�/�0�3��R����f��yw��ee�)P~���*�vf�g���6`v�R�v�/�qB8���wΣ�'�6i=U���@ݑ��ͽ+��`��qF(a~C���Zj_n�����ب�&�CU3�wz���.JUgV� �֮Ay[?Գ�3���n��*�E��E.ۇ�f��p��Y�UC<��l}i�DR����]���ߙ��[��tC�%�4P�'F3Ut���lbzYJ+�&(�5�j��/���*�jI������k	���L�!�T�Q�1�r!TO1��U���[�a�_k�O�dH<ٮe:S�#�G���"#����c�(8:ʤ���x9<�K3��L��>\CL���ĮGݥ����,q�[;�Z��+t�s�Ke�'��X����ul���Or.����?r�=����;��>�!2 |������_��Ь���x����R�s���$�f}��n:dN���
�ctkG;��앉����-�
�Ǥ�I � s�"fz>K���X[L��q�R��vzl���	%5�ų+� o9�"����~$`��߅kJ��OR���O���\֙��	�F���l�ţM@�|6J��.�Y;��lD����wj��Ν{��JND�B�@��u��{T��l�
 I��6��e�qS��P:h���Tҵ;1�o�:Um*�َ�yD��l�-���s���3r�+�@Z
z�M��~l�KOn[���*��	�cXj�r�ޘ2��v��AxJ�O`��Ϻ���Hw�1b�~���^X�AǬ��	81)� }O�쪴�'�d�2��8���T���tꡩ��ї�s%�
����a�h[9�6����I!�璻�L�ʤ��#��F#��u嶊��׫NFsDl4��
J㱆� ] ~�� =�Eigt�w�Y���:	�OL�3���4<�1{,��O�E�jC��Dܟ�GNt�����g��n���V�o��d��՝ �GE�
>�Ֆ��Ǣ���D�nhH6��X�U  G�����1���'��}����[����A��ADȵ��./{2o.J9�?��\�_ ������i{LO_�vY�ۚ����|��4�z���R�F����t��Ş���z�+�&H��+��I��ÑK��g�<�>E|�U^v��FebIü.@�vF��M�{]��]88�*�*�U��q�2e��ywY^t�+�b�#ŗ����'��<A���՚���^4w4mв ]˘ 2Ř�e�@��jK�OO�%Ud�y��;m��Ђ���j,J�����_��k�!~<���\�PpV���؏w�z�mf����:ܢ��̡�Zd��X>��ޠ���W�@�q�"��r�����:�}}Q+1���X,n���n��LU�Fns T�dJG�?4�}�ɶ�~��"�Z����Շ/�}X�[!-�ʤ͈�!!)��� ���F��cyYs�u�>��?���>F15�ˉ<Q��B\�#�@��<�|n.s��*Q��JL��8���(<��A�~+E�0r�v^~�HB�ˠFz����j�"�e���'�#�	��K�>�QG��oA8��>�2'9$�Uٳ���8&a���"�L� :!�B�����,~-2�m���6�Nj6�i��鉰�~�L?䙶�%����az�]�0��BӰ � I.��]��e VT���\L�'����q�">2<�̔�j3)�)�wو�a��H�/	i��0L���P�F�� �	�\x�$��bn��e�t�����# �V��"���t����c��Q'���qC�����m�6d@�Q������m����!��{<��7�~�E%��Uu<��M<l�'���.6����r�e�/����M>br��Q[�x���A�Dz�v�W�9��P4Ekw��K���W�3��h��FR2���M�6Pm\μȐRX��Ԏ~��{�3��7��@�q*'x9A�IU�N0!��?�d6�x��` �G�q�����Zju�س-����%w�b�9�<ɋYa�ϠRCqsq��4�I`o�����;��7�9�������j��������+��;O����|�wgΪ������@b8�n�k�P�ѸN�x��R��e?&j�o���D��&L;u�P���xܸ��z��'j�ܙ���V3U��3��"!��;H��G۽�*�F�lWeQCܨQ��s\~��iQ���р��a(e!�Н��[�c��DTY
������[�6��|)%��Ϲj�=�w"�m�}�jU-��(���Sݏp��r�^�M�>g��ڰ�{��f�cŹ�6��MeFjܬ�KxƱL� �l�4m�'sYa�BE8V������r_��G�����px@�������
]u����]���p�xX�b|`8������S�n�Vii��^�)e}/���z�`�ԊFc�6n�_��)�-�P��C��AЖ)	t�X
��w�V$|����������
�z�������#.`��-j�h��N/7����	>Y��/DH�'���]7>i��^m�ܽ"��{|��X㶻B�: 	�`9���]Ve�z���t#'�悟��J8F~��؆b��� i����J���,�,�	�wy���z��T�&&���u��Q;�<m���6a���ĊK8�~0�蚪"��#�6k��*�Q�X�̼�o���=[��7� X�Az��,���Ӻ�:��U%�%�.��r�8������F`�:5t`������A�PNֱK�>��h���%���LD��	�&�Y�Z��7�k�c���C�|ʻ������B�0Jg��ax��`T�v!�y�Q����=�z���X%�^�}m]Pp����=�N�˝�b{Bo/�b4�sE�=D�<y���p��,�o8	����?�Bl~m���0b�/��{ۄ���] 4���a�Z�
'���טs,o-���;�8�.�xќ���3݌�I��լ�'�s�)�������G,��]ގO�׻4V��bm+)���B+�u9�&��OU�v+�~�+�)S�(�a�
l:���Sf�׾��1��{מ[�hz�{JC��l�_�s�u�?�b���~�8����En���վ� ۭlQ��d��	�-{��_��f�#
_([��f�H��Һ����(V�2���/nkv��ʧs�┷�B��9���~30'�����<?��]�T�<*[����aa����}�֤�0���׳���<���w?����6���
S�ywA!y@@��� Z����T�FT�����I�a�'�B=e�1 P�C�ܸ��DF�XT!tV�?����D��Rތ/���ڗć�-�xn��v�uPJ��0��|�#��ylK:��
5��~.G��蠹ry@�I}�8�^��)�Ə	[p�_Z�������]�%;�;��8��f�
��:�XZ�H�!c�x~Z\p��v�o�l�t�)/�Aa�dY�}2:s�W!����'���r�����q�D���v��|����2��0����1��J��l��`0��ƮE��t6U_���~&�Y.��Gk�~�=Sn���oOԥ!����|VY���+&���2�k2������Η�h1��S�aB��%m�j�J��j{�b�l�F1�י������)�!�G�eZ�x�!��yۺĭ�C�s�߱�~'[np�a,��^b�"΀��H�Y��v?wr�r��TQ/!��l3Y@|�����,�HA�s��!�~ %*z*���9L<�K�`�*Em���୆���"��#�^�P�h�H�0Ұ�_�<��@;����i�@]�F�A�G�7X��0�x�纾��a���.��'�T�@%:Z��!���st�6�J�c��@�]55����^� ˙��V�X�<N����I�kf�����ҁ�޻d��&ߣ�)Hp�<*�F-�7�������{�݈�Ђ�!�� Q�L���=�FT}jp�����:�D�3:�.�N����L3��fS��D8�U%��*mK�/��p6�@)�Wʈ]v4!縭a����^��MF��U�M��$Ë�O�C�bZ��~d�ny9틥����n&�w�\�9i"I6<���<�Z�㛱����6,�P�^>���q�=���g@
��.v,P ��S��q�Y2ɟsKD8����Jo�V�H�)٩Q�u���5���4r�僲e�4�F��l��~�j�5��C=0�;h��?r�ȧ<"�_
�0�Tke����!����It
4�e��ʠ�K�Z��POI(&��P������ؒ'�]��C_B,���0K��?�^��ѣ��&�]�3)���� ]~D�L�D��6C���$,�U����T��DܥvW��	P��]�fv�T�.�pO�:#��"]�2Z����D��e'5��v�G�2s��X��P0-u�xOu���r薟���~K0F�P�%>*k�0��g͓!g[M��(�H����1�J�ˤ��/=�N���S_�SN��{yW��U��P!��_QL�pVY���N�-�Fc�(@��|r�)�r;;S�%��	7�+�!�J[g�Q����QZ�����h0g����<��b�irT��A.�w+?����X�^V5]��d�|���Nf�~`�}L����~�����@4���T�+���	PW]aM�>�L$�W�	�kS>V�d���W_)ib������U�׉��#S���T#�����0�"B`DA��a=�S�@��C9}?�|3.��m'>EU�.��}���`�%d骺	3�[\��pG�L�US��o�Im�O�z�;���hW��W�9B�fG�	�YZ]_1;�{��4�<?Z���r�D��>|g�7�c31�*�ނ��ۖ��"FFѼ9j_$^��~jӦK$1�P����	�R21	c��)Z6�;�o&�Z_��(�[�ã�<�9��G
/����}S��_)��ꂰ�K��P;U��A��s����LkUV��U��J�X�tZb����W�G��C�"��W�t\+��>����
���̴N̆u�7��u��C��<���OP#1)5+�5�F���F*dê��9�H.�s�;r�VTKa�⅂@'Ϯ�����]�
��,B<H����]�Rr L��@�ڐ7oLW��7Q��E5m��Z�bi�`�����������"��{A��'$�H�Lp~�CI�-�(����~�I)N��FP�F�I��]`}�z���h.ݿu_p�š��_�u��Y���cS��/�����,v)ʥo$o���� ���FXͳ�����M����x�8)��犃�[ڇL��-�n+��CVL0��������`H�q����;B�b!�����N���缸�G�H�{�t�8���L�*��3v�q��M�f��0�yu�IL$��%�� �Uc�D�!t�&�)/�-�6oY
�<o��<����:x 37��62�kxY��6'�hD�� ���T#Mjg��|M�%���VF�8|m�ְ����$)�г(�;�����"A���_����v��#���fZ��s�L"vO(���Y�CU�l��N3�k��n#��d:fuD�`ˉX������X[���CfT�'��l ~�̲tbL�x�م�x;��`�wo˲�Z� ����J�{�AM@<e�%������_�	[7'����R�pa(&��x���4���y˺�J���#��<\6l�V	��0������Y��b ���C�� ��l!E�]i\7�r���"���`F�v�B�y�SН�W�I5o�J�O���_�%�z������]�?��u4��]>�z�/A��+�XD�+�g�׭��ݒ�.�;����,t�D	���>�I�4z��)�J�����������<�ؐ������η@��*;���2����w0ʲ)K�ǘ�5�uA�*L�SNq��������{�\i���{�5��$Ǝs����"P�A�&:�D�^�^���@4[x�zV�����"?��/l	:8�L׾9F�T��p�O�r9T�d���w	$����搐 ���`煆�&}iW����3��$�+���'e���i���Y*�%�Ѓ�yu�o��#? �G]��஀�!��,r(���@	g��C��� 8Ze�	�|�� �(�~��Ba�r��H���*h&$g�F�a���!$~��
�DG��5�T�I��;�X���J�lЄ�!{���ݛ�7$w
�b�F�)��I��H�Ú�MZ֖�)���k#K��p?��?E�Y�IY�]ս: ����;"<�J�y����Z#��VD���wD}KT��$fyY�������{J6�3�#i���^��]�mX���.�&?�]�c�ˠˮY��!�{N
��e�
�0�n��8dW��,�a�\a�u�/E�ƴy�R����(1�|�<�C�P�$#� �k�{uV�N���T'j�a�p�MM���AD�tf�x�(޿uN情�e��̃�g�p�b_@��*�"(MCH7���O�Y%_Uj$-�ż&�B/]�iN]�z5�m>���x�����K(
�������c?�Z�0E��
�d���@�hU��^��)�~+����W��k���Mԟ5t��Bk"���P~V��*c�|�����v�;\
�B�J���Zw�[��@��!��������nv�<~�ȯ̘�]�O�XA"{~m�o�ؖ 	�hbDi����Ms�8 e�;p,�K)Q�d/�Lo�Z�$�l�q� ~N�W��Dd҈�ER�~!Ċ� ի�o7[��4$�N�t��~g��}\��|����<�xҒ�)�h��:�B�B �F�sK %�G� I[����0�z�q�|y���xmT^[Y�n�P���TDkѝs�p�mA�+�K��d>�n��)O�i1��Z&#�݀�.�zYė:SK�-��V�g7�B�8W��	5�L�b��qW�S�=V��|H瓐:AO��80D�<��H}f@=���`�`Q@�9�HH
?�@�q6��xy�� �Y+F� `%���}+&"�PN ��+S �{>E��mͿ�ua�*��;�i�`���mZ��,�ւ�28�=�#PY�*+b: � �3;d-�uW�$_���W�M����-���c9�/���(ղ%<��5#�'w6��~^Tِe�M XƩ��8^���E������_�ㇸfY���ϰSGo���o	�挵�+l4��4��v��,~���?`}o
��2��� љc�K��r$8�ZN[���8�4z`mL�hO��<�ߕ��/crc��[�{�-�s��8p���W���d�s�E�	1*�8��smwOM6���֕ (\��	- w���<6��|8����'#Zܮ��o��{R���dLpc��̉-n �7��4� q��"�AI(ֽ�Uu���܂g��;�R�\� ,j�eg'\I�#=�r��k�3j��B���� �\ޱ��Y�C ��
�G��x㇭
Z Um��%�A�c馱#�{	��n8���`��P�Ќ�:dʢ�N��OOm:\�m/4`�S�~�ގ����a�`=�u8 N2�[Ǽ����2�(u1;���Ju�2-43��7eg�`�EL�4���krT��B��=���pN����q#/iB���Jw�s�4��.M+Ayڀin����"��GV�����_ �����v��;Lu�_��!U#��,Eً�=�;��יpN��������������h�ժ�]Ox�m%P�g���{�	�%Ol��M��u�sv��@<���[�^����M���JG�"���ױ�vy�V@�P�!�0��	8sw�N
I�;�퓆��]���5J�E �k���w����d��F�ڮZu�����]n�h���5��ߗ������o���9#��ן�[_�_�!��FμH���	,]G�f���AG�o&�G�[<o<����c� �K��F�*�Jg���y�X�>!�t"+3u
t��k���:o�@����c>��7 ��Y�N�L�ð��|��
*BZC�Л�+���VN����;�����cɧ���n�m�;�Ӄ��"<�؀?cַ��������b�}+̼����j�&Ƣ�Py�Nud��1�� ��&�֫�,�K? xL����3U�<q)(˙�Z���{�������'{�@��k�S]�zז}���\O��)��Up]��llw��"����xu��d!�����9��L�)�朽��4�IVl���M�_d�[z�����X�[3���~�J�MP|�:�薠�D�r�YpQ�y[r��V�Y�G���7$��1 G��|�R��ܦb��/��#���6׵~�};B:��=��i`!*�|E)��W��2`�Y 8ݺD���I���Re�Xg��Ѧ��R�@���KP��YT�m���:A	7ސ�uBt=�rZa�vì�q>�P c�7BbԐB_�Y\�\�j>`/W��l���&�*�۝��/q���}��E=��3HŒ;C5�N24\&ґ&{Ӛ��{��	V����V.�^���$R� �R�t��q~$N��=i�Q{p}�
uLT��b����[�8a���7r��y�L�����54-�i�Te���І�ws3*���(�����BS���E�%��[i�$-��z���k!c��D����"����dN�7/$bZ<Bylj�k2e�}_�^���6E;�o�hN�����������X���}�x�����s�8b?kmW��Fχ�/)�e��9�n�u����j��l���Eƀ7�@��3I�!*�N�d��c�ޘ"���X
c�dO �K�ħW�k|iHF.n�^�!4��H�d��r�ɪ����%�b�n7�.9ʎhA�S)Ꝗ00��K&�uzM�o�wga)���i�@�ј�X:�آ�w�z�R�9�&!���=]ݯ�Qc�CY�<�B�R�H����W�)NPn;�wЊ�lU�Tx��B��=�`�%f����#.l������ ���	�i�_�|5���H�����[ͺjZ�X:�|�̀8+�	���n`�+���'j���L�-=AWp����:�j~��Df��)��%�N�L;�Z@J%��"(��B��Xݳ���@Y��A�q���~6�!N�ى܋���b9��')��/��7�N�ё�(�]F5�7F�7<w��f��r�~��I*�f0q����A0��__���b`��j��*��%+Iw��b�6�^�"D/6�Z��XM�E�!!�ɲ� ����ux�TM������r��9=|�r$��_#V�1G��=���:p�a&n)�8�
���N��֤V��#��A���5>��0��Q��#��[�f(jk�s���2�NbLJAE�{���i�������ذ��N:��k��A���M����Rǀ���r�	Qot�
�bn�ȹ�����Dn>�e�c5
b�X�&�מw����F:pR�=���uh<��A�^�u�me���ΚÄ�7���	���a��[Nğ{ ��D�
|����?Hn<�blWg����(d����B��a+�8��~X�$�r�;���'�&��8���x�`��Ё�����=kƮ�Z	c�bZ�o'�R�UCaN��LL;��8	e5�ԇTܺ����B^$��Uca�E�6h����<T$�!��˟�!MnA�雳N��v���U����kׇ���c�,E��AVf�|�nïjyC������쒕.�f�K|prȲ4I�z��%/:���B�N�fC����+�Td����z÷{)��Z�X���=�%��$�"7���2H�p ��[�uQd�����D�}5��X��C�O=7q�M���׬��O��}��9GF��^ݨ��=����ٟ �K0�[��k�O+4��Z��R\&����>DPu��������"�d!wH7��I{�j뺚܌7�,��T| �����*i �1�e��Ծ�Йk�����̩�[���:I&b��q��Tea �	�G���jx ���[��9��;Fdy��M-��P.2/}0\ȷU$���s� ���c��y�K!�Bv���g5�c|�,�Lcl1VH��<6|�׍��m�t��`!� v�Q����C=<jЎ�9�R�r֙?k]��F4���\�q�D��ʰ ����`��>����]	޳����c�C��j\�j��=��& 0�7#��G]t湸7�iA�Ur�����ѐ�P�S7_hlJ��ʋ���v��fh�ź}@�ˢ�h�x�^�Dv�@��x�'�ڂ�Ӟ/l�B�<���萧��t$&���~�?�Cؿ9����܋�U\�|��X	'2%r[�x}7� 
�П��4�9:��̧=�%��+�+�</��b�"OF����X?Ʃo*�=�w��M���^(�TZ^��J�"���'qka���E�n
�3�ԇ�];���n�� ��p�T��aT`Y����e�=y��M�ik��d��;�m;��F��8��0%��$��_�W{$��1�iE�!�%� &	ޢa]x�(�[���E�s��<�<̷��$~j*����<�B���6D�u
�&-sEU�
9b˭cM����׃no_D�h`<W��a5�6���TUS����D����;c��sl�uk���t:�x�i����ڴ(sd�B����(Y�V�� ���M�W�=�@�U2�^s���i��	 a������h
�f�h��E����#��i+��qD������R��A�$~@5�¢��<ؿz�1��O��	l��R�c)��((�9³�Ls՝KF���
H^)b͌�'K��+{h�Q-�o<*؏�<<�FT��YA7�ʯ�H�Г��y�H�鳋L�S3�fݓ���ʐ��,��	�tr8�
=*T��f�d�M>�`Y&u��}��߰Q|AnN�zS��_:-�<�FH.A��\��B��Yx;��?� qq,J��$��;Dຊ�Rs|���~��#����N�~1���l��z�b���;鹎�[�,f��%�b��B��܈�����+��*6"�ý8�\u@T�%L��r�,�X]�n>�+;�����9`, )~d؎>	e�A�+��'��R�n܈sV`�}�� Vf�?Gxh�(tz3Ϲ7��_)�>��T_�YR��B�Jb�� *p�i�m��S@Vf��b'��U5q�c_���,;���5��V{|h�����B2���$�S���'Yr�5w�� �i`�Ă=H.֟���r#�O6�u�#�T�e!�M8%��6�Rb�б����Jo������&{6Յ�� �����0tc�[�C z�^�Qq9$��|�C)�tYd�C8V�Չ��Rtq�J��@ˈ�X���zQ�������hْb�N�G�I�(������l��(eÒㅫb�YФ�Ϗ�{d
0X��$}��:������������[m��sŻ��.��ɑ�8����)�����ˏѷ'NdT4/�˫�J�7�x��$��قhB��P+:�7���
ғ��ǂv=%��ɲ�F�!d��HfE��imT�
.��#<��.K�)�jw�E?e�g��e�� )�=���)���<���6�}i�� �"D/'��f��d�ji��7�ZΚ�����2�ߦ�j����ܭY;j_{�0��U�8�=S:�Z��a;�p�+dA�ƃj���tL@\)`~C}�nO�H[w 1�� 11c(�=2�qͱ<��hMQ?
n�#emm������a=����(؂M���*������`��%ӰQ��dZ��M�}"��$i�<G��ID��y	J"����U��x�p���%��y/i0�ѩ��5j�	�_����GKWH��*��d�!B:Gej�C�T�ۮ��.���e�����OSP���k���p��	Ӡ%n!�D<�l���Ř#\�w4C
K��j8hշ;/(r1��v�#P~����,��|�x�3yCu�Z�sQ?�<���^H8�*��¤�U"~?��8ie%;�;����#f� u��9:(L�am�q0�,������9��LY�� **beM�����ǵ���l��4 UA^:�����4�K�}��dcO���&�L}Gq ט�����O�� ��Çl�ل�<��L��	��K�oo�[�d�؀p�����7�S���a�j���S��(��yV�l����L�M��D���y?sg��'��$�`Yc��+�)�-!��ͨ���K��+�Ϊĸ�e!��Z��m��sL�6ާ�Ϛ�*���E�b���S���^/�X�q�n��ǟ�E1R�OrQ��W��<!��U��H9!��#�B�H�U��}(F��� ����ȕӮo8��a��O����ř=���e��.�q�1��S: ���R&�g��G���ֶU�օ��OkDAs�7o�Ƃ(*�}R��kX�S:�0�X���~j�LpP��L�P��tmH�0��K����d�ЯF!Ƌ�#�rV�}��P��chSd�������/p�Q����dx�F�%�`nj�"��N���0`���7����̈́#��*�|�$.�p�1�2g`��B�[�~���~�[xc�	��<�/𛓢.��	�w0n� ZR
v�h���wa7�g���
�kiƆ�ֿX��!�B��~gVIl!�I�_nD� ��½hM*��5�a��Z��3IX�+®�[�b���bq�e�� *=��_�7$j��w���b�]j�.+�Dl-��Rs$H����}�;^$�� �+��ʅ���J�QR}��i�C�	W,���߂1� ��O����e�0��.��=��񀶷����J��?N�ƾj��h�t��a�#��LTȗH�u���b2z�
`{������<�Ȧj��"���g�kUw�����G�)z����c�Z4�R�?�����gvg���DH9��U\9@3c*�}���Y~�����ᵸ�Z^A�|?:�Q�)�[{�J�/Ӷ�L�*G3,�
�eh]�ɥ�?R�$��'}��� �<�ON�=@�Z{�����ҍQ+�2Zإ��)$k7'�(Fh{$�;ED�^�QiO�[��W7�%��7!z�0<P�w��a��D����:�QT�W��R���]ڢ0��U�����6ڕ>~�A启���^��&#����o@���킯�ڎ�j��LMҢj\�ń�i�K�b�5�z˨����ȕ��Yj�x�sn\(s��ږ�:���J.[�{:!W	m��t�⸘���3�?A(�r�MJ�-s��[mu����ut��&�St\��l���5o�����`s�	E�@
�YQ97	�4��y���2H�(��f���=�
g�{B�%~�:�i,�Ev>q����zl�b\���P��סa9i�)�5��.��.&y��ʓ�R��N-l�G��	��vcr5/s�X~���k@�E!Oe$p�Y���pA7%B�=Ĵ���[���k��VP9���ټ�����d@O{��"�4��5�8S�)d�:��g��[�����>aXH���t����������9��#W_�`�R��ٱJ�#"�Ԇ �4����v�r������̾ty�I5�Q�j
@z�UJ�@u��GbS�A�3�SW)���w.�A�c:d�8��/_�2_ӌ��u�����=3�Gs��T������t���Ql��t������* �%���^����4�.����X8k��{0��g(I�
�(�S���CR��g�#m�^,���m���}�����a�*Zj+��B�0�, آ�%t���@'X�lO���A������ߑ�	���ud1C�b��5ʣ�K8{c�i�>���Z��QTfg�E�C��y�ǜ�r�+�Y`��<ѩU�uC7y�y��G��ڈo�OCd"���4����p�9dbԴA�.|�S1� ���p�h�m,!f<�ߖZ#��0�3ϣ��������,�\�ʸe��Ŏ�VY�;%� Wm�2|���L������8uN�F���UNC����H@�>�kX���Qt���M�Fs�m��ŭ���#����Q����h�l���7�M����3�]�5�A:!cv;�tw��_*"HD�ۀ�������Y�C�{�b�ŶGfE��Wq���O^��u�$򈛂2�⁲fƐ� �f��r�'R;3B8`���
�jMޡ춸�}�����qD�6��°wi�I��҅}���k��Q�+��D�y����f��[r�����:;l-P����T�$p��Cv���.��#jg=�������K�t��	����?vӭ�vÒa��͙�9�_�*����ݻnx��'7�G�i�N�~⒀���B���'I7��
����A �n�N��|�8t����$�2)�C>Ї=6�4mxr�$T��dӼ����p;*n�H���J�dtR'x������je��^Sd��
f;6
��Ӥ�R̕|J��'k�8 ������P�s'��5l��(hƼ�|�2,�'���(�^NT�d)Fif7�3	��Z�����1^�X'��l����օ��ksElDz%�km�ɻ��-��Xq �3��{�(?,vͼ�O�r|�O��6Ңd=���M�#n�=Y��K�ᷝ:L�W����fS��a":�������"S��
���2tX���f��]oi6������q��ڤ$��G��Aj�q$�脌�os&+9]�\�A���	����H�C�d��^̰#+�JI:�K�_�Łxi��~9�#E��x��`3_���K�7��d��j��E�"I�f;[�}�;��S���@���T`Ψ�	��X��e	�F
M��I�f�W��&US�a���N@qڿckZ�X��L"�`P�)�:$
��X���p��/���D�FnTR
%�Z����op �������/=��Y���H�lأ��=�h�~.��<Q`�gc#V���Cw/u�M��
H</�`A4Ʉ�/>����8@4��ֲ;�t'GB����NK2���t:�Y�2�(�3�K3���AS��"l�Q��-P�
�^|�d�l4�������L�+u���[��kPG�O�ܚ�;�x���x,�HXX<]�Ϫ�m�AKGEL�PWE��\F��ۖEy�P��C�j��^Zc�bB<Q1� ������(� �Mx�B��(L���R�^�Ջ�YgW���/ң�q�6�O�)��u�,��� �>�㔤.���W+k�cÞZ���W���L�N���Qw�u����A��D��'�S�ߙ5G%J�o�7��[V�<?����!�=
f0.'������D��F���Sej�T�og�X�>�ˏcNB"!%V�7�*[A��~W��(o'���y�)�6i�:=U#LSM:���壮��P�MoA9C��� ��fR?N&^�S�/'��4V�N�pګT�P4y �ZGr��.2y�O��Ʊv��nᇴ1��y��F�ߵ�JzUٺ��h�&�S��9�5R �=��{[��"eN��w������v�$4�P�|�(�kv���/L����됓Jz�Q��O�#���[�����e)r�뭪�r�~zX�LW3?�|�OMͫ�����(��(�cHsdt�P�Z�^ʕ�m��K�,Haw���L1�Ḡ�W��[��źއ����U�z���W�G]vv)a]3�߆V����y��_� ����P�@������5��W#�58 ��LV�i�qL=�̳(��j��͑am@�f�LȺ�~��kL�U�z��C�;�fm{N���FJ/u�8��%�G�r:��8���!�z��OT����:N(W�En�u�];�[W�$�G�J�6�W�M�qF�U}8�P� "	��\��@�����Ȋ���
Z�R��M"�n].���NU��g��ܯb�6�"��	M�l���˷8B!"�O��Nt,��ݼVj�ss�Ǌ�_)��(�Q򤽤q��X,��4w!�x4�4�?��_��_�������b� =�����wb��FՍ耭=�k̾�&P��X�r~����&41A����<�)�[M*�V�(3	e;,�Auu�5�l��3�O"�wݚ�?�Y&?�<�)G��y/1�@��+0r�
Z��rM?1O�� Uw`}%Frb�`�Լ "�fҭvx%���w�B���9-:�X�@�_UIt�L�X}�1��#�G���^HI�b9��[Kca�{)��8�NHVD�jl��|%d�i�-����Vʛ��'��o���q���+4f�[�b׊���Vt�}᳏��Q@��th���J�(����&E�<������rQ.6G �~��G-���YƤ�j�'�-K�d������2����n�M� 6O(��"���0a�RY��vw��+�4cb6M��L��:�N��#!��܃_��==��z�D#�=H!PNC��2���<<b)Ǖjg�F�!-�<}�,�k\,�Bk֬(��(S�����N9����A�@���K�eC��b/��*���)�7��d�zί��B�Y*A�ܸ���D�i
���Q�u&��a����q���h�d�y,zz�B�X���ϙ/	�f���m�%�ُk�y�z爱M=��Bh�w⑲���p@)���Ka��"�T�]��֜�����O/N���/�ȅ����W5El6�3T�F4���T�sN�!l���=���j;�:�f���YRC�0�D�W&�@1�Һi'{��|���4#��0Q���?�F)!*��\���>���9YBݧ �&S����v&G�Qm#���(u��]��/��ƨ���qd�K0v淊�p�}F�-~����)Q�X��$�³�$]{��N}��e�ղ����Y�v��:�य�:Jm�G����眊䈆�v��jfgj���Şh3>��S���`x��T�)�ҹ�?��C��S���N@?4���;�"#I>GM�������Rq4SGK2J]�Z�Zև��̨���}��{&lZ_�s�|�+�>m��Ѝ,Zr�0�����]2R�QC��%>(������x�>{�A4�<D��!)s$�T7C�w�Ț��1s��;q*H�M317̙���)q��n��Ά ��,!���[iO�a��;h9������m��j�v���%��W:@(����2S9�ԃ6�`ƃ����n�Ĵd.	Ѝ��V=¾��Y����Z�^5涛g��J,�x���?��p�~3њ���)۝Z��dH�f�ט:�˶G�+�
w�"?M�h�t����|��Ru�>f�K��@C-�Ϩxa�Eg��$R����zEԦn�+vY�^C7�V�|9�"V�Z:� ��8-g�]��Τ�>�B a�oi{uOX���!�ܪ(K$�2A\�*dL0V!D&�R�[Z�t�=��Ġb�HT��6�~�٪��'{x�	���CP�,��0<���/�J筷��H��y��ʘ�J֓4���2U��$�{��������ϴ���n:��|]��.�5p:*sOfu�X���7}�.r���r���>�#�h1p�n �8���-('+�:�ᖐo��?h�-w������;��Ԩ3�L#c �u�S�@F��%ģ+��c��0XvW�Q$�1I�8�=�`���#�?�,�x.�9�.�[��'ݫ��� O,�$.�l���S�����Cx�\��Fӧ��4�2sM�dLi�/W���o��y���I�4�p&�]�0Kb�?^L�� �n� �wS�+=�e�V#ԧ�qs�tV9�g��L�}|�̚�L�$ex���j��Lxm�|���p)�T6s(	2���[�V�A�f�%�㏛��(��Ck���y��f]>��� �&a���P>�!W�)�~ۑ*6sJ�W��Xb�ы�4u��ܩ��9���!��H4z4V��T�4]٦F������Btc!#�9?�W�@�f�2w��`"c�۝�kg��U� ��@�]vs6�_�Ђ����gb@(wW���a�׊`I �$`�0���?2P�"S�u��h��WW](�@�p֓��V�I�����,�)��7�"���̙�.�`()=d>�5<��OZ+��%�#T���dº�23��;֔[d)9dw��_�8��:�3f����t��=�^:����,�73x�U� uH�I��2�C�^�W�F�a|����_�)n���/X1�J$�i eo^��
"�n��1r ����А���]�/�{HQ��u����6iF����K����R��?�(V���!�i�H�O<bzos�.O���7��ƛs�tU2�9Y~�FRZ�������l��U2	������7ܭnJ��1|>s�cڦ��=����:KA�T��d��\������q�ȋA;Ӭ��#��-T���-��*�<?�:X�o������p��J��S�1ٶ��u���iF��H�`x�PH�i.����[������L�����c�9}���V_�w��ʇ(N���䶮 *�����Y�ի���	D�r���o�;<�t��ق��< f��ο���t��r1W���r��G.n ��X:�aa��'e�ǘN�`�T�A*@n]�2��w�r��Fa˪&U�`m/�F*���o~��HԲ�ez6�@�mE{R�턡�$��?t���Ph�;4oo;
�i��W�*�)���@�1w���W烽���M�Q�ة�}�|�+wk��Ь�.�Q��m��{�)J"���~���f�` {��`t(r� �
��;bP��đ�@�s�rV�Y`9��%�9Lxc�o���9�w���ICv���`��:�W&�-��������uWP����)B8�sI�3yk��1%��V�04����"��d�R��g8��{E��Jk��IF�|c)`R �F�a���Zk���ɳr>x,����U�b�zB��|�K�)���n-���'}
��,�}�T����6wH�%E7�0<gk@zC�K�t9VB�!R��р��cw�3�Պ򏔲�_s�X�'5�س���)ZE���E�;|vƽ+�#�-��;��|1b;ؕ�:��u�XY;�B@�)�����_i{�5��D�M�FU�C�,1�K����Bu%�Ě$���kM��[ |���I7�ʏ+~ �=*`1�	/�?d;c5պ��yP�@1D�Qjذ]��C��}�d�qm��{���,�>8 �iS��Vh#���q�5���F�y(���؋��yoG=6V	�P�(~`�#���P%��]^�r�H@�A��Nߊ���;��pf�8�n�n��S"S��J�����ñ����J�Z�h��y��hF��e��\ѯBJ��Q�_H�k�j��nN?��}H�����M��5��S$uC�Q�$1��du��~���X���:ҭO�x�L?R���t��mKg�Y_(`��|s@�]�L9�4�~'�gw��g�y,[�aȚ,�	n�u��?>}�*�y���;~9�!_W��4�)G��\���V�ʖ����pS,�����������/�M��=R.�v�`>�s~�~㱘���z���*pۓ"A� Bm��&�)�M�->��T��%��2k���1�i4 �&/�U��R\�,+UH!�s���T;�.5Ҷ�)�I��t�\\�����F�佷������-�U��v�wӒ�p��?WJ1z$���J�a��X	s�5=��H���gq��!h0��"��P�hCX�}rչ'������H-��ɯb�b�~��v���Z��l��V7�ۑl{��-MDl'�y��1�w�PY����kզk��h���-��Z�8%v]��|�>ge�ΜCA|Q5�nEk�f�R\���0�il=���W&�7/��.Ou.!VC������.��⩖u��Z�F8<�ir�9�baDS��9h4�cr4�U�P'[M��)��_'��{��-=��UR�ޡVggo�/�z�Va3�f`�frr,j��~�94E���^�Q�t5���r���w<?�4j r���NS�JӀ4M���2�U���L��HF����@��ڛ���6*n@�P@�a��$@,�z��)�pd����T�J=.�&�o ��/-|k��'��p3�;A)�5��ejg=i�#��%�(�=��mQ�I&2y��X%�aǓ �"/1n�	>�sT�"�H�H,��g��-l���"��0u���pr�sxf��m�B0�cSw�.��$����{Q�>@�]�3��ӈ�j�z�.fF6֍�&�n�J�Q0ad��ImK�' ��e���\���{[�PL]ơ5l���>@��,��b�������DH�?�k�='��笒�t��K0l8?�T���Γ1���������o �a�%ٙ�R.���%̈́8��3hL�J���y@�����Y���=~[�[�b�08?r�(!8��\5�z���x�Xa�3��;c�u��M�ƃ��s���N����+�\(���k 5�'Uۼ_��[�#�|]�6�|��w����N���RǓ� P�7�,�{��oǡ&.�
�6�8�}2�/��_���Dp��G�A�dT�̏i�Ɓ���ðQ�{��N�n:����vE\�`�*�{Q�L��K��W6H�y��~�%:&Rf۪�ĜTܟ�Օ����� |$��
v')3��wV���qɬK0@Jo��q���h7��_��������9�����Bʏ6o�M�Ļ�:]�p/�mQo��y��e眾�Q߈�F��<(�}�q| ,o���.n�<Ż|\|	t���ؤ�!�m)�0��mE�Co���#�����N��Y�u�L�O�i�DT��A|��l��j)����t���������Q3y��f2�R<�R���.��y�o�ا�oEɎ�)�9�� ����ڛ�"Тt�
z��~�tՄ��&כ�9��ڀ��2@Bq5�����P/)u����A
������.�ܱ,��8�WS��X�o��A�̓�52���:��=�k�5I���Yd*���L1�d��7O���~�1���D�s�J����<?܆��r i~:���Ck���?k�xϿ�ѷ*�V\(��� 6v>�ثG�b��}#i�1!^y��]��U�f�B�&�,�̭�L/u�x��8U:���f�j���C�2�=*g���g�^�76�'Je�*d����☤�Z�e�x���,�Uf�]���f������䎳�J7C�a�j&w	�@L�vM���RLV�k6��Q���ЮKl��Y��H�F5v�J��a��3A.�0�	a�453l�������ty�D����J��&�U��N�N�bl���B�k;ZĔ�YE��%�T=s�N��B�=�H[��uǊH��@�6Md#��5�ԧ(&�ꑉ��o�_U۹LD�>I�e��2�Z���{э�;��۸��������y�ܗ(�LA{�J)������Z�G�78ݮd�����;R�+���d^b{�\��U\��6o��;��K�<Q�^��px����p
����ٓل��p@��\����K ���L��Z4v��O\����1ᔝ,1��"L"/
��}��C'Fk/���|{7 50�my��E����J#Ě�����e�Sp)��fƛU�����B��@�����/�2|���°��X���&��v>�0f2c��9�,����zZ+_�eE�V�8��i�����R��N^/�[�k������R�n�6�i"u	UbC��r�K���7�q��'O���W�JD?�$�O���E,�]��=�-�����^���}!����/�H\&��b�1���	9�G���v�C���+"�]T��$�Rg��z�x�?j퉼
�2�\zK�I��b;����M��ĩ��?t�u�/?�v|~�~I�x�- ��Y�>|"k2v���W"\/���m^.H��?ѝ%K�����N�2H��C��9��ړk����0����Y�-4c�;���/�g1��m��y6](�f{f�#�����uz�U-�W����8�T(Sz�r;)6�*ɣ��v8�s�1���h�)���WM�n�V�r�x�w$�tC�uV�lG��p�HD{�{T	ϖj�c�NeϽ$���s�#B8��jo�Nǎ�Kmk�MV�G��|�Ā�;�L �yj6�_ +��AV�����S��P�H|��4	��Dy�g
�;ί�΂�����\�U�MPKS�o��\ �愇YĢ����t�u��"���˲����Px�]Hj����{���uӺ���Qń��vn�Ģ�Eva������W�~]!o6U&b�"��5O��7�嵘b��jaB�Oղ����B��L$�ḱ7�4X���z*�hşk
��i���U�Q��@���$ThS��������Fi�j��Ⱥ1����reV���8���	���2��
��a�=FiC�Ud`0���q[�E�QH�5D��ZΩ���	�E�j�86O��@�{s��a%#0�?_i�/��p�5����ս�>I�r�����v��`h���u�T|�mx�kL�������zu3�аx'�'x�R�,
��Ѽ�v��>2��>�/�G�7���%Ή�W�M�!�TP��������o��L�}.��Шd�����;����6�����K�`��"[-�]|r��+�&���w�L�@bRȽn� ��d���F6m��df�"�jJq�c�rr� T�Z������?t��X��ـ�8޻	G��WT3[��ի�m�Kl˺�1�[���A��6��7͎>^O�W����3���%��O4�Ӯ �T�ie�O��`WW=�A��3��%k�쯼Y�1I�z
� �c8ZF��I��A�0�'�v�c�\Z8����#�ή���5���0��sڷ?�ф�Ś�C�2�R��X���Σ)/���G]�w���H�/Q�PT����R �?�Y�a�U�3T�~���!��~�Uvf[Bͯɚ��5s��\ ���ƍk��ѵɭk��*8�a#�=��wm6!c�h�� Օ
r��o\�^)b}Y�6+����~�Y~�0���wwd,�*�xI��do_qݮtt|�9���,�W%D��TvZ�����MF$�hl��)���,�ED��i5T�:����O���,6�kF�%�A�b���x�'؅5��䂊ZM��c[�=�M���;�����6;�M��K�����i�Xh�C)jb�\O����1PFmI��H��!|�Ax�M��N����`9�u5r�K�B�����5ʯ`�,�7Ίis�tzj��P\* ��)α�WP٤�c�1|�����N?g_����;+uξ5*�"��'
4�_v��c��ђ�D��IW��q#w8Z��;�b��z���
ț��[��v��Ԅ�q����2d������']��i'.��>ȱ3�ӄ��~�!�*�6���D��?���y��T���a�eKq����U�E�bdO}ـ��X6�O���K"ЅH�rP:��ܥ�ΎU$ݺ1|�!wh�w����,�B�/���]	]]���k�}idж���"}�_�gT�>,��a��r���L��ql��B޾�����~��=�����o��%L���o��K�Î�ub<G�J
a��6{�o/��� �#�,ۡ�=�L�vW}kD�~nHw��Ykd���!��OO�*Z�Ec�T��mZ�W����7&xC������� �}�0@�~|��R�"�Q��@=nɘ�]E���|a�L���|��6d�(`ҵ�O2�����YT������Z�ϱ�x�f�~���Α�<�5��>aے�����qSg����k����ؼ�'���<��B�d�S�K��DU��yy���I�|�pXJ�@g�I�8?}�'�����������9k�/�d�+'�C��K�2j��gK�o�c,�Iޫ�!�'�^}ZR Q��������(UQ��)����B(�\_�J�wa�h���rp�ϋբ8p.������xq$�^�Iy��u�J�B��_�|V�տ��B�8~qCXf��:)���o�O��`�����<��W�gM3k��r��7�b�ĩp1��M% o�:�9����\�� �ێ�~�z};�=�<���n���@��~�����?z�s��n�o`�|��^%�\nQ�O���vHw����(F2lZg�:&њH��҄��YE
lKa`���p�8m�n�B����۲a��j�6T���.�CXv������Q���j�������2˺��{��>�'�3gu��*�>8����������]��<����[Y(Hl�'���D�h׽VQ��շ[��#�?�M�I���xkm\�x9� �2���+�rY#�i��[�B�l*8%А/��/��{#��"W��pod��n"�Yu���R������)�z�ƫ.BS��$�u�0X��+ZX;D�R�gw�����on�M�/�o1}q�Zu�苤�S,�M�&#+�����U�4K��0���7LZ��%?����yN�F�y��oU���h���J핶�!�H'�-��f��jޟ)v�l�����c��=ʉ�ʖ�O��һ����x|Б�=�����Ϧ/�g�o�upSM�<��"�� #�a�ss��;�ځ�-Liá��]�|:���?b�H�~j�o��V���U�uu�U�@ޗ�贅�����a]4ύ��w���#Äo�}���1*������{'��3��dD�a�4� ���&�3���+��B���I��8��o��tz
C�e�U����2� 1��+�;�e�mA����}�3"&�4��ѯn�����t�k�0F�k��뀠��85��a�0dc������ӫJ�g�w�7R��(cU���n�V&�f�1��Ȁ1M)0������������u�6��r�'�O�}��U|Y(�',�p���E#3_�G����������0�~o�z�B�|���M/$z���
DU�kb��sc&
<�������ҕ��Լ���Vց��=i@M5��pR(VگE:^������B�{�VȭK*ݐcV�%�A?=ݯ/g��I}L�陜
�#R�txΛ�<��)�]`�v�'I�&���,&�������O�u��I�@�-Z��u>���!�`X�x�/�|��4��SS.
� m�;i@�᤹|���W~.Z2��9��J�*K]��!�{j���1@�٩�L��R�c��J����!Q��	x_����]-޶��I�[�j]�VA����_� 1s�l����@c�x��䆞�Có?F���־�p�:��ɷb�^�:#�.�\�~~ �g.D��E�y����6�xW����wuLo|�����w`D�{��S�lվ�^����BӀ����7p�/>!_�2�F���_�x�z���:k�b+��
�l�!�6���~�A{��`i����:d���[��%SQ��/��K�����H�Щ0�C�>�0r��b0��n\A-����b��y���N� / � �ä�V�ɏ�z����Q��Χe;�IC�G����P�9���G�mc��l��b�`=F]�ծk��պ!�k�:���̝���+�V�[zԆSܩ���&�[Ɋ�U�p`���;�`�-�V<�|~�7�=�=��Q&$<�ՔB��7Y��a�a���֍�����b{(���� 00�6
�O�;���䗧bԆ}��"�������c�:�3�juޱ�I'�.���𺎀립�A.;���D�E�O,�I^ T��3��������;�r>������	�eՏ�!+�E��'��kd����ăC1ֺ��L��iš{k���{�ef86jl:`f�H �طP'G>�X�h��t',g��D�8��!���< ��}C���w�?��NI��M�g��8�?:�u{��U2�"=@2�ܔІ%8���`�73��#	�U�1�x��}�#İ�"��K�C��7�,�����w)p���Y�� �j���	ľ�&������5j���[�P�|��Fy:�ǜ!-۶I��� =]�
f�05�&i�'F_Ar�jմ̆6��"�:Rm	i�()1ݺl��K������MRp��M��k[ֹ�$� �`��m�t��ʽ�R���1�%s�)d�Y yȦ]�_����B��67;v
�0����E_�P�(�ZW��@d.��7t��ۋ�[b[6.���Y�	8n{z�Up�y}�'Rf�maJә��B ��}{+� =y"B�O�Y|��
J���m.e�̐)!A�Y������C�f�Sb�!_��p�3ӑĔv]�Z�2��lTgh������*�5؄�`���a+&���^�eQ�=�wf���Uf����]���{:^y(�%�wvM5��SY7�S�f)���HfF��Z=��-p:�u����c�ߌvBo��e������=���n�y7��型r?l��o��!�N�9���-��P���0���M}�;��CI�n
���0<B6�/��B
!٢��G�rW1��#��R.��6&WJ����&�}o6���BŰ��A/�x�9�Ǡ���fF����B�+��<�Q`�k=@u}�N&�~P,�vCu�EH�ݍR3�i0<�q�2�u�{S/JIn2U���i�z��s��lH�U5/kU�Â�'�U��Dr��h0|���f�N3����s.��:���9�O��P�'�
RA��6��ݬJ$[{T��Ϟ�Y
�q�[6�ԲJ��=S�N�Y�>i�еY�Q������a����b��Ei����ǡa&[��5.�$.��&S0I��&�p� �t�;��L�qaq.�V�׈V�]$�5~��_�]ً��1��-����}3��|�0�m��|���g��C�0Iuw�r��a��*ء�	����=@�x��sZ&�9�h�E}���3X��q����)e����uLm�1�o�v
ylN� u�w��zR���S���%��E���#d�Q#lo,ݹ�<���R�Pv���^Ҵ��jp�]M��#����Bcc��m�������X��okǹ
q�p�[;Qa%���� �$�L�;�S	,��9�K��G1��r"��!������Y��%.ۇYL�kyd��M��އ���e�m9}~���H�2�@��ٲ���'A݇���4�E��IQ<����Ǖw�&�ӫ�:���O]�d�����VY����n���V�U�9�,��
\ʤf-{�+?1H�q-\�Fͮ"�Kʁ�3�\��8������D�Ju�9n��":>V��M��|g�MZ�TBy ?�5#�D���=j�b�Ѿd(/��E6�j���eG�� ���j���w�"�<��'V�M���K��Iz\��U.hp�ᮺ)��9R��V\>�X�٢��-(8��@�'�^Um>��0��F]�\oUtM��lI������=�$��� B F�lm�˪v���8y�bK��jc���C�(��X�`rB�<��}��d���"�"���"���ʣ�3�%�H:���dek�ޟ���*��n���b��-��)���0��@`�?�`�;B>�ɘ��l]ݶ��`�t���(���Y6j�7؁4cj��F^l�^3m{'`��g���S�Ѽ�	~-���G�u�*f�z�4bl��>#I��+gVܣ��&�e�	W�.��pɐ~�i�����<��K���ˆ�0fg��YP�U��O����y� �h�a�[�{Xǝ�eܿ���A�9�܃�@�	�io�j���B��!;��1'�_��� �N|�
�)ծ�D ������67��͖� ^i�������w[��� �A��2��C��c�)��30��C� _Jx/M�U�@�<K�c��?�Ɇ!���)^nRb�a&�0w�"��C�)��t��G��mR�}�@_J�+���R9�V�byV7KKe^RG�H�.$y�����#��%�*�*����&�BU�Z(_�u��őM�W���:�t L�z��0&��deO������������N�wI^�����+�B]>hY�8�{ �j˼�����MĚ���=s�ُ��00ή��w����7B�����Q샿%��˩I;����u�s�µ��2lj��t`���ν᧷���#zb�����>u��R=��yNe��`S�S�㝛�\ʹ������v+�e˖�A��l�H���\����] ��Z=#�W�J�TZK'��̯��f��5��ᙼ-����	����N��<����	�C�*6;O�o�Z����M#����^���]o�%۝�bf��ǽ�t84�%>�;t?����$ �/��[<7��W<��� ���j�`|U�	�Nx�L�`X� �<�׻5�ld�3n,�4�R�&y�/���>��#���v��LҚd��qO�%e��3ڧ�j���m����������PB�9�'ߜ��F�c9hM�%ߚX��BiΗl6�wyd5���z���k =%+�	�a1�B�B]����ێ.�N���(e��mݥfT��ʯscu���3����ش�T����Lz��[ޱ�r|&0��YGk�0L��>\߇$B�Z���=(1e����K�E���m���N yB>��V��J�\�/յn��V��߫�+���U>��1�LY[6S*���i��~��~jU�Vņx���9�I�.��A8�ҡ����Z��l��%�*5[���1W�� }��a�h��`��̔�_d�J'�L-�n�����2�]Ԁk?`�F���l��~��WZΥM>9�9�шc��Tt�ۃ^&�硹M�Z��i��=�62qf{�nx�$�[��N}쉬�et�X��i���!�0B_c�k����+r�-;S{�[y��D{�1����b�x�f��NW8��u���EW�?�dCHg&� ��m-j��_�րQ ��1\o��&�B�^gt!P����r�����Q�x�eM��-G��˫��O\X8%ɲ���h�sE-D�Ї[>eN>Ü��@r�U����j�`�a��B�0Af�Ȍ����$,��sq"U�-	���|�
7��ܛ����z-�����XZ�B^�;:,֨����a�x��-�!��a��������?���=�2� �N��Qj���G]���ȶw��l92ޫ\5f��^��";����gS��M�qT���7��ӝ�B�;֝r@��}x��sP�ĝ7�q�eB�6�/D���ے��|O�%�TC�)��~_#�#��rj�O�s����!V(�G��VhtT��E�ꌡ��y������>���J(!��<�n��0�q�ޤO�K�fON�m���j�n�	��/�b�^�.�w�yh���������j����a{j�V�nO1���~�%�^I�����<�j��t%�a
L�,�*om=�7���z�H�����Ԧуў�d���Xw��q}סgp/V�l���|�����A%o6��J2���n#���L��6���^d�q`��C	mo>��]	�i[p��.LŌ����N����A��/���������6�qh�0~�T���r�����f�
A��ا;MR��+P��k���r�E�M�^ ��N���_��X�$}�sD�/���]'}$��"�e���kAE���e0���~
 x9��?�Q�˸�_� _�c�l?@�㯽|��k��H�V�=����؞z��k\`��;&/����~wy� v�^���Y1\��Ir��H�ښ9���T��W��raD`��#PĚS���1�?�]��KR�ٿzX�N�ڢ6	��6ڐŞ��N�����J!,c�ij����G܊��"���gZ�mh~�0ݤZ!�>4J��^o)�-g(@�`g���bB�(�M�9ㅾ4�M��e+Dm��x�uݓ���^�O�-|�a�va�,VN���_E��V�5�D�3)�� �ff(�֖��g"�4}������bC�k8\K�g7���I�����~�&�*�SG��F��J��;�ַ Uw��V����9��X��*(�/��M��B���UC�����IĲ,	<����~�ԣ�qdOms����������!�,q��1f_P����QWojhsU
�ڰ�S#���aJ8P�W��[��o�0D����Ҷ�z���[uw	hv])]�R�r�<iëu��R,-;�������� �Dյ����i ,�+#=�������6��4?�K~���E;Щ<8l��� �J�"�d4���f��)\��rsD�F(O�;-ɿKP]�D6bq���)�X�%�y���]~��=�G��!���9+K��ڪ�����,�GGm
��B��Fь��)���7��r6�hzҎ�T��1#�8J$,�g�C��\�I$!���k���c�\��|���*��A�_He��0��J�D�iJ��;���>�\`M��޾o��$VV�,3�uT�ĥ�Ԉ?Q=Oar�M�����b��k{�Yŀ?���y[�����9?��4�r����]ӥ��Di��p�\��끝i=+�|@f�W��V��r��R��0�w�Щ��#s��6����ZԱ��>0h}(h`+���B-_�M����S���XC���ѯ���]J�Ex� fM�.����RSl��H*R��;Y���D)�Z{A�Lu�f�����|��\
�,���g�K�q��_N���i	��Kد�����5���'�C�w��m����Q��=��� ���@�.���Y�#L��3�B۫;�/��*���U:Ղ�A�Mi�������@��<[���qj�&JO����Ҟ9�3!, Fd#^�X����
%�t�W����?)/�Oc��m'�("��9"��12����]�_4����Ky�A�dI���� �}�>���mX�-��T��a/��)ҵ������"c�wb���ۅ%�@{��8;����$7�`��s�W���RZz,��n����pSs��U7y��7:���?�+��+�x�>y3���DewB<`��?p	!�y�V	�^��a�W���������̩���㶓A@^��D{�+�2��L��gKNGL�=k,{�Ȋ?����GRA��j��eٶ���%KA�Rd�:����!�4G���z���+�F*ւ[6(+� ������TC��h�y	���>��MP�<rf�-8��TxN�ǎ�-���H�J�r\�=�)�J��kC�u8ɥ[�Jٕ\�*��ƻ���+`���}��)�Sǖ�衤���X���%{��ߥ*)Sej;0	ac�8^i`o6��=���R�������(�ǐ�two�����j�Pn��L��@���&<&�a��%����)�SW}ך���Ɍ����I%5�V��3�`Ĵ�.�QT�B�kM��m=N
��vr���S�k��|�k �Kn,�qnp.���%�m�6N�h�`����m�:���F��P�м"�����*�pÁ���;�:�7�A��>?�?�3�{���SzjO������=n; ���v���j�C��T�+E�����ɜMA��pk �a��5��u���c�r���V;��7�?An����k���n���ֆ�ǧ����B�%\�0������^�P1�)L>-�6-�f�]io2:�{|���Ϙ�7����6\��-�:��C�^u.��qٸ��\�f��s���Eky87~�n��b d.a�(�C�U
�"އ=$�`�74�7�,re,EcWp��K�W6���3�}�����u�������2e.�[/O��V8��fm�(^?��sh���+�T07cq95,��:���_wㆡ\Y9C���31�H��;�Wȓ�&g�o��d-��`��sց�W^����kC=ե�����Z��y��o������03I���{լ}C���R����0�x8i�����S�0 $�
ɽ��d����o���8;�c��*�B9l9�>�{K�eD�Zygu��=��Z�qd�G,���q�=3�P����P��u��MF%0��$�r	��)4\��i�?�ھ%�M:�e���1G[�GWw���EH+n���n�Y5ب�	�m U�o)~�H�g���(C"���H)Y��/�1�,�l��<Q4�������+����{�i`�H�u˾\�bj�(��K� U=���aO�O������2�SF�o�2)��3�� �,(8�����鷰��{Yq�c@�C8h/�������1͓�������VZ�_��-A @�	�2�Z��N��/���͒�A��O�H� @��Λ��p�������]�����B� <�W��B48v��]�M�h�?��v���r"������C+��нU��<����a��͝��*]"��6GS��ʭ�nF�+qMl84e���߫�z�Z �
O��t�_S��]����ez�=�#�8NzC��b�����v�x�� ZLҨ^X��¥o)B�^��DwI��P��z�@�)'�����6��y�v�$K�6�˥!��fm/�l.Qg�S�Ƥ�3}�t�@�N^	N}��ɋʳ��O�e����ɟ�Ь0ѫ�\���M�lzzN�$n��>jJ��)��4�፰a��(�n*
��~-�vᰐ�t��?F�{u��)����{��T�}�ꋮU��U�܏�S��/�G�[-���B�&���$�F�پ|1���N��\bK;�?���֝�Cv�Rq�5d�c��X�v�FK��~i~���!b_W,V�[q�OnBew_=g@�
^O�b<�|�\Re�vI70�@�̧��I�H���+:�p�x:hP�JI �,�i+J╴�'n~����_A��K��
τ5#����'C7�|q@*�i��3hR�n~i@�)��7srY�@�}�?�7b��C��"�N�
^��]s ��t��&^ �.	0�	�0� �]{�(���+2�$��Ss�	�س�}���j�W�)�����b$�f܀D�h�H��%��YI������H�W��J����j�5�NN�L���^y�S�-c�����YO���+L9_ ���9�����mc�W�F\�z=Ɲ���͗-�HT5A�.���,H���~
�U��S���̚�a���1ɻw�mLF����gP*/[]��z�4��~!o�n;���Z1\��Q�*oZ��{7�ZB��px�-Yto���z�^o4m��.��?���}�vX*��������'X��g��Z���g !F�gw����m
9�m��#p�y3�<D ���Y�f��%�9˵9)��(iu�Dd#3\AG^���Q5��I��)63�)���|,}-a��P�ݑ���r��(V�X�������/g�\��\��[a�0�@.-��GuL�$�N:G��UTd�gK��w�9:{�":��ϥ� GG��Ȉ�"	���AUb:`#P���Bm�Q�e�\t)8J(o�ğ��5jf,G6�40I���wj���<i׮��Y��Ҟ�f�?����1̂w`��@��[-s���R��R�͛�,/y#/@N�'��w����׬8��Gkg0�C�p�O����_[�~�Ń�Z��n�- nR۪����1<��Ȉ��ѕΐ���u����e#�یMN��E�-`�;���z�yć�E�J!�?Y_���GCy6ǖ�#�jj~��_�"Lh�5?9�~�B
D�9J�*���p�l��O,�P{.���P��%@��,�[��?�.w����)�����en&$���B��fXX� �����|m��Ҙ0m+���HX=�&��I��AF2����Bʅ�,i� ;�&@$�"���hO�IH��{�03O�z��P���H��nˣc6�p�Uߒ��Z@,r�.����Ã�(Ԗ�[��u��M�6r�*�	�T+�#D�#^^����y"d2E����<��^�7���#b�!�s2�����Q��3�a�S�����'<�G�"Q���T���ɬ'EM�U�=�.�#�=A��mԃ?7�xx��	`Rv�{�Ο2c�pr��˯��&'�mu�6�8#1�Ti9}�|D��=ӊ�0sj(*~ƨ0��G^�TzP�jG"s��-��V\bp.�	��^���<Hٜ�K�*��A�&sN��5_��D�bP5��,W��V{�T�L��,v��Ȗ���cZZ]\�}����F^��01�'�zDk8�;WZpñ�.�ޕq5xI!����˗�MT�w���W�6��(��V�m�kAYt��v�  �g��Jg����I�B�#Ŗ��A�C���*���l�j�t�;��/�NJ:s�#��o-�~y�9p|��
����ωy�W�l=�}�����*���*���	�t�B�x�����������)Q����_)��q�f8&����d~����K��%�6S����e@@7�������\( ����x�K���hxg��I�2!�Ϗ�"u԰*}��,mk2�J률O�LK���L��Qˎ��eX� I���	����$8<���Uf�G� p�"�����IȾ�Wͷ��B�u�܂�q�4�_|�C�4�1�p��İً��<Y*8��_��}k�N�W&�.t:�P�����.Jh��N��f�.�!U��M�4�h���� �f� ����6�R�ڤ��)B���u'~�6��
Oɯ6��Ag��!q/���H̻�|&�Z(�������4��[�l�
|�g#�-_�ZD3����g-�˛����GqH
��W;'���@����X����\�N�	��P=����ߵ��	>��0�M�W_爙�t8��uv��_"��v�e#��,a~��F�^�P���#�VQѴw(�&�s�S'xݴ0��߄�
�$7��n#�1/����W���c�R���q�J���y�m��|�ט{�3�r�+h����(�`��������<�Y��%��$jY�2;\%�h�c��4�6�ڏ~l�H�O)+ٓ}�+w�p�ju?a��J^o[k��~Fv�%�)�fI-��+ �_�I�L�Ļ���W�s�*�+�ܐCݨ����� ��K�E@���)�2
~s]�1x���Jd���BO�f���E�.CR��;s5�@��B4
��T�k�膨�[�v�V���ޢƔ3ގ7K�t2��3[��a�Fz��ױ���4Ch�%��&,q�=R�8nO��x�����J�*h�Ή�T0\��6^��J��8�N���&L/1~<h�CY.��X�x[Y���##K��^鼏��������<�Xe�I'�#4/〱�A�i�����Z�{�a,�KM���>�'��� '��\5��A�i?�fJ�G����(�;�]sՠ�i�'/��;����;���ar����A�%�}}(oh���r������Mh���	���>2v���l$�tdoPXt�:^��m��v$}Fi���)�9>�g�t�Z۱yQaEF3�|��q�ݎ�c?�����w�7�B�.��/�!���ݹ��-rH�W ���c��_?M��Ǌ�i4�jB}5�������(�ʐ8��,��y���ˈ�*�ő$����|�����8�JCRY��w��D!�oV]`�vH2�<fQK�+���Z!��P��9԰�����ڴt�1V�F�b��-2�[����atCf��$���m�o�E˷�ٝ/吟kK�J��a����m���+�X��a�0���E�.��nA$Ə�f|:7Q+Ă/�T���Q'D}�l��?�Z�>P�����q�&q���#��ɠ�+�F�;�������Tr~���.-H,����vgμ_Շ ���^Z��z�k��	 ���5o?�^�!qV��y�<�2՛��	�ҦjHi� ���=��UE��i�Р��O��g���J�_%?Ӱ\ՠ�������Er����bA+�:P�c_�] K��!���=��o�`���7՗U�����u�꽵�{s�����đ2�Qgs�����%��C�}�|�YD�+�=h�M�̈�S_f�L7�!)F���,*P�x����`/O@k�rSC��S^DY�M���mhZP���=����d��w�r���Йr"��T�c�p	�濗���;_"�}s��������q���澾j ��p\h\L�M^C�1�78��͡x��`� ���r�-�xyrނ��)U����r�a�	�<^���f�T��q�Y����'v/�aVm�P�4���N��*U�e��+8��S1��?����:�>:�d��KL9�%� >s�d�ë_+*�P~�^јV����� �Ir���e�±�R�)@B����Z�nu1��5\�j�X�o�M�ADB )r�����i!n8n����3W8Dj<��-�H(}ڂ"̽�ܲ{-����}������5U��'��?�y��5��t�`����d�� ���}.�k��Kؐ9�8���ه5ܳ�.��������T���%������.ɖn- :��5���j�F;�"¶�S�)�<j��P�W������N�T7c�3|����=�bM�Q�\�Gڃ�K�����;:����_��0��Hsuݓ�ӈ;��u��]�v?�'b\m�^+>Yx&Mj��R�CD�?V�0�d�c?�x̼�ZfHL�-L���BP��$��w�E�ku���}GB��w�I���{I]�(i��Qa��Nϣ��SUeZ���6}$��D�iu�+�ꀁf�MM,a�8�X�������+9g��<"B�aX��3��а{�G�w��9�m�A;7
Fe��������)�v�n�9'W� ���u��.�%�]���c0ݯrwq��X"B�K9�	��{3���;3Mv�����o����?]�;ߜ�E�	@	W�c�K�%V{r\���M��ݜD���$�[��6r�v#�L�V��F�:O ,P��?ш�� yzRJ:	t��^/�q�)�w���s��"�ykp�/�
$rj:>2f�����U�n�kg�g��w~]�B����A=��K;WT�d�gI1�=w^��餔G��8Iu��h�����&��kJ�\�aڍ�
�p�`3=�H�&vz$͸l`x؞:p�@E*�:�)΁a ;f֟rE�_�W�֤��\pz3X9���-�hp+�G��N=�*���<X�ք~�R�j�� ;tǂ���C�MĢ]��
�%�b���@�_����u�	���qM�)��a����,ȑ�L�Y�$��MU���/{�'	9�A$�PUU�?���sԅ�πP�j�{Sh~�ex�Oc"Ƈ�Xs��~G�h�rC�<�t|x��9��z�q֓��C�"�i�=s�u���I&0#�<�696��S�
.m�jO�����f?�R�i�7�0��tc�v�!;�����p������	~�LB�-׸Qp�h}{@�:}-�D'Ł )-`sYVq-#y��Ա�!�_�z�p����S��3��������P�O�qS*����eb[*Kfu��J��<M.��ev�����NIsA���U��D�0X$̔���ծi�`�����T�H �85��p��~a;&ل�z�nϚ��į���y�;Ui�+�7�J9i�ߣU�*��|G%w�l�F���BD�+� �S���za���:{.�NR@3�@�z�&2b0�!K��ɨ4�/B>�/����-��q������?M�ר�x��O�M�5vZ���͔5�&RB.@���扣�n4��5�6^��X�����u�<0t��/�>�$��u�E�OzT-��'�f�pm�#;����B�SG8������Gί�.4��~ҍ��uҢt�]Zk�hk�$=��ꕖ��/C�W_��(��sD�"��A��jx����bTi��/P�[.�I�����U]��b7^��������
&�W1N�	>Ä!"o� ���C�Sp�x�^o��I��p+���y��U����vm���=�e$?�f��
a��� Vi%O���(U۟��ݿ�w�.�e35����de7�ew�'.�}�ݦIG�����T�|��Aţ4��(ğ���`��bF設r;��ZV`�	F�h]� �rE\9N�;'�B��˪
v��ϩi�iw*��о�ܽNw�� ��VQď���U$�uB�s�HZ wFo�8��X�N��N��0��W>/R��?����0���f�.��^���2��7<�6��
�ے�u��@4��/�zDB;uX� ����S.�]�� v!#hs��76k��'J�Ʊ`'U�S)����N��I�p��h�M�|����.�S���{�SN<8mP.[����ՈΛf&8q��7g�y_�����;nd���"����
�Ҡ�K<%�f�s���k��3I:+�J����p������<rY}�c��:���� `�ek"�G+y?��p�c�_G��;�t��"]{�Q���Yrl�fIֻ�b�Cd~BU�ҼḞQ��{���sC�ܝ%���3f)����"���&�ф�i��6�z� �B��}��4z�Y7ɼ�\`ڄ@U�����v�	�Ʊ�B��a��ݤn*�a�����\��yXuw�*D��oY��X����8��hF�)�3R/�s�������7HW�yjn~Ž6��H���;�k��q���$V�<C5��چ�2��~(��'YfP�`��V��^
<��Z�"�^A�:���r��ʁ�8��z���K��%�(k�����L�G4��m-<�H������z$ٴ�|؄��&Y���Β�����J��j��p�9��@�!��<��E���Wc4D܋ࡂquW�[�⟆.�2��u9���o�M�i�35��ƔBBbr��x0�<J�x5%�@�_�Rf�����Ǧ� ��^�c�@�eVd�����gB����¼"�����[�s�����0�1*������*٥�=|�QK�<�
&���֮��B�.։��)�N-Հ���9֩��2֫�ճ����|"�+ �x�`��#��?�}���x�Y���Q�X��v��V�o�����U����w*���l�tQ �|��lۃ����{�I�a��5Ya�/�y���Ҏ�hn����T�$44q��J�H�<n΅�7=�w���e3�~�<��2OC(o�VA\'BKs���|n�&����tm��zņ�ƍvƕ���Y5�,�#�J����@���͉}j�3�e*kA��V��*����m�� 'r������ق���yX�&��.�!��g	�|��[�����]�VX@�O)�������]��6�ꪅ��Y�k�4Tw����!@��~
o��-��1P5e��6��v�s��Ic�֑lhе6W�d[�2`����`*8��ׯ�f�X�rC�'G�`o�7�4vՏv�]�7}O#A�|�i�D�׃��ȟ�4�^�T�C��<_Y���1"ȳ���vu�sؕ�=��⛍���q�z����ԮeNA���&�ه���l��5�̝j�=�M�����gq0�<�xc�}��w{�[D=Kb�-�������U�w�%pBTO�ȒO�52�/��bx����@'ۘI �:���ޏ��2���̿\����`�)�&W�n�ok�0e���Æ�<��=�y�\����|'}����6w��h=�޿Y1`
2ջ6Q?K7K�۽}��ӽ&�k��K�I�i�</*ވ�������<�ћ�-���g��_ՕH�cCI�d��[������47D��?�w+;�*[.��F*�ӥ��2�zcG�UU"�%Pȯ֕7[H��}�@0�W���`�#~Og���+�#u[�f��JpL��@U���hߪ���M�����,���%�*�}r���B��U��47Y/)k�g�e�I�Nfem�oŰ3�W��ܰD���'����!�B�p"(�"vp�ND劶�%��# 5�Qj%��+0 6s+@=�L4�M�B+�h���V9��j8$��.0�I��!g.:�x�n��e���Dp�����H.c�U���_����d��.h虃r��ו��mJ	ڌ5����Ɏf�Ŋŝ��	����_�48��iC����G�<�aYt$A�e�Z���D!�a>�5(�~C�U��Ք�ɮ%j�;�m�gI���3qo��,$���ݽN����LLA���qSi�?�tO��B�J�{(|��))�̺�F�_�w_����5��v���� �>щ;N�W���x����F�r
&��q�*9�ˉ�<)�����z�b6��k�2&H�	�j�	h�T��庿W���	촺�<u��zM�K��
,���1X�~��Q�9>aIA,�[A��^���R�2�t�f�Z���N�J�RZ��۴HG�L�E���B.�����v,��ppʯ��+}�N�)��n�Lj���υ�ᇓ5��ߴ�)���r��u-A�^�d:eN($@�a����*�.ߡ,��Lھ�����4���y͜Z�=#N�$X+�������|��,�؅�e�8�Ly�z��aC�P܄ǔ
�v%�sL���<�H68j�:)IJ�T���O�������P<��L,(6�SL'���*k�oh��B����D������`I�q��l=:��e -��{��<�^��]�U�W(��KJ���d����R���)���T9,s�Y�O�b�w �p�~��'�5���`�E�������Rr}�Y��(��ڪ�֙��$(��~��p�������+�=Dھ�>.��M���Y�w�F�1d'Dn�N{��u��H5G<�թ��(F|�l>j�%��+��R�&S��&�&k��-�jř�M��	�O$���s+���	��ִ0ӊ|-N0<ʋ̣s���S���[��ى�&#��sa�=D�����>	��e�>��o��� >ejlr���n�<%n���b`S�0C���A59���d*Vc]h�Vu���J����lT�]<DS{�֋>��5#��N� G�Q���E�N��<I��f�����ߣ���?:�Lz�lM��8��\�lMJO��)/���H������؄�Q�8��׊h܎吵�B�6��hhbŘJqo�I[������1�c�\��}>vc��&��lO�i�R���K=1ݳ��#u�KC�M�� �H����É��	���v�����\\FJ �0]b>�{>�7�I�sª���4AN��J��V���D�Bt�JN�� �:����۳m6�L������h�Q��X�Ȏ���[�m�b�=��^�tT��?zd��h^�hi�<*��}���۲����/[%V:yw�Ljb!�D�f)å+l�&�՝U���l�ѓx���^||�Ho*X�/�Ҿ��;h�_&�8$� ����M	��C�1vdz��oF9\��]W�j��Ƥ��^6��Vi�~*[�u[WY.m�����ˉH~�+c	R��ʟ�����S�1�D�Z�����pxY����OjQ �����ĺt��\f};����Pi�JHyc�\6b���Lx/�ĵj�s��(r�b�=[F2ݺ�4|?q�L_��|���,FqZ5�t)oʰ�s�;�\�MqD
��殪 .�GL98�#CK0f��HCH�*tb�T���j�����<�#:��xچ�^���O�xj^��JB��_�d�cC�،�l����C1f�Dd`�q�&�$���y��k�k����d��7�'��O��&@��@��v���뚰ֳn��m�<���F���`�I�p������?��z�D��N<�$��87��,P�g�?�@����(��џ��AI�����&X�g!� 9X��5�8�⦱��B�ip��+9iA9�S=�.��ȵk�『Q�o�%�b_ytAI�;�uc��e�!��i_�������V�ں�o����K����3�^��е90թ�J�+�o;��\d�hq��IQ�:���~(V��� �yڮ6�lү�.3��10^��.�jl�՟v��7W9�b=������j���m>���gA����8�rt<��l��V�^FѯM|wHS}�*9O�P���*�uč*|���V%�θts�
�ֱQ�.��yf)�� 8�乻w_� �Ok�4�������X��7����G=Hx<�r�Zo���Q7ŭd��!��ǂKX�Ro�W�{{��H�L�F��7V��	���K�\�Qwߡ�
V`TK�k:�)�����3n�Zl++�D,�[�����pв��@	o� "�P����ҙ؇@�/��1�}���U<� �f�݉��y�J������|��6��:f�Y�@Wᡝ�_@��G������5C�lM]І���?���
�o�W�0�6���au+d��<��'��,�Z���u���{^�-��-;����;	�և:w����ag(����t̎�.�KҌ ߦ� y�����(���e.Xӻ=�����,�~1[@��3��)���ے�/S����*6�ړ�ݪWh���3�g�ꦺ���8�"p���2(S6�G��G��_�\4�78�>���z��`T�$�X�D�ˊ��k�yn����(�/��|@{�\��']o�l�w���㛯�"����"�Qwf��p�� "0_e[���b���-����b3�+qȻ��f.�L��H�z=�rn,�CX-n\:�'3�e땜%?�d��������W���{�~�8�7}�qG�\l�P�s�������T�V���2	�Хë2]�ʄՔ��]@;XRsA�]�Ds�;���S���7$�BY�ނU|{:����ee@P[>�1�n_�(F��d��Z�	��%x{OF�.W���p���f�C��	8��{>:#O������5��)0�٢���<����T���%Ș'P.'S��|@�WKf=����N*��Y�ź/0fFo=^� ���y^�4Ǎ�C�l�?���Ш!S���ǩzxt�Y5n�ج�1AiX�Oo$0@�)�����*��>�	�9��-<g�N���߹�,#}��_h&TČ��������u=] ��,���� ~�\�j1�)�a�K\AA�ԵPF0qs�[��#��j ��
.�v���:Y���I��k�~���{yZ��`A���mWO��K�v�2��.[s!H�/1J��n�eT��";X	˴x�����k_@���:���$#��
2���r:�NB͞�ò~ �7���.�H�;|5-�7c �P~f
E�l7�����璯Y��]�� M�3�-Q,6a�'�=R&w��K(d:N�
C2���k��$4�?j��/���ansC�셓�� � ��E�aD�/ Ӱr��&G:M�������5���6�F3:��*ڛFߺ�
~HTA ��(s�i$�'��r��Ћd�>
l�x�9��&�� ��G�+�dɖ���2r�> �o�Wk"|w��b�͹�{��Ѥ�>[���=��
�ц��/,Y��U�JX����(4���@�v�д����[c:��"~Py�-C��!* M���p������W�7w�C�*���	�yjP���`pp�����O�8WW9���7�=�E�pɞ���a*3�:�,T��qsw��#����o㌚�)�z��F,�1�	�͓{��5d��U2����4��s��Mh�fs�"�pZ�r���?��_	�ͱ��0Q(Z�2�5C;��<���G�Y g��@�d4"�]zjA+�����xg�Gqq�,,��>�Tg�_Ot5du�tQ�F\S�Gm���D����Bm(z�v� �E[4�a���j('��� yB	��0�[�B1R��yDb��j���N�%��H�o�͊��Ҋ��ĖC���\��'�%�a5��{��k����<��М��>#�o�`��`Yg�ؐ.�[/5��L���i�3�Ae������7K2� }���E?�"�ƱY�f�󾀄HAT�ht�Tdu=4�����8�wgح:YUQ	������6�ԉ�p�靼��'���+�N����NQ���s���1{µ)�~�p��-$QA�}�R���m'� ��P�Tw�@�gi0X#� ͑f�BR�ӱ��T߲��x	+�O��7d����Gh��:4Y� *b6���[�`�R}�Y���.�+p`�m��n����X7,E��N
 ��]��4�_,��%�Nc=�>���$ƀ��=�t�'�f����%���.d�PVק�`�&E����^��.�(l�?_d�Q����=''�^l��N�+�����Ke������f<þ��s/��G�C'�#���io��8a�F1���z��R��m�F����Žog^s�H�m���KRT �-�;CӪK���|�r	�{�CA��Ӗ��*��O�E֑^���X�7gt"���	���Aw�atm�Ę�w�Uf��X�
{eh�l�%af�	+Q���W��}Kw�����i�au����@,��#�"�=����3wm5)�!d`9�k���B�Jb���C93Ğ��<�mP=eE�|���(@��AZ�XOI�5K��B���^�'l*�\��F��QVA��q|�ڜ������E�.���{���*q~,Ğ}X�K�M������3�E���8�c��t6�C,Ц�e�gq�G{�L�S��e���7g���d�~y�2|D���?�]�I{p�
QY�m����C�v��d�![�>%@���=�^B�؉�9����}px� ��* �s��7�u��:G=Y��j)CY)���aO�|�1�<�	��8�6���L��ޒ�^&A�_P���q�>��^�zF��$���*a1�^!�D��{�$Q-�� ��A�>/�A ˤ����IC}f���e��2%��и�ѵ���[/��jls��oa���W�o����[��h5�����cb#�T��ƹ�D����2��؊߳]谒�'��#o��g���d�O|N�TE�c���Z���>#k|��ȃ'�=�����|gO� �	;�?�9�CH_�f�xo���}�Jr3lK��>B��nV{���R �A��/{A�-�����Yl��Q�9�ؑƨf���JDu�`!�ɱ-�W�v�p�����6C���:T��75��)�`�-l}��1j��+��&��|�ӛá�k<���}KT+X�ެ�/<P�,�e������Yyh�4����$ߎ�!k͟�@[9��#���H�e�<oy�"�%\" ]!�=�j��c9�t=��EK=�LZ��@�flTWal1+>��+se���1��R G�d��4�A��^�T��6���ۈ#��&�@Χ(�<)mET�3�<0 ����"j�`���I���X��}M�GF�:�t �P�5i�}-�/�� cuU64�<85�:w����A�D 2���ж��QӰ���?����m�F��ӝ�FI[*�{ɑ�*�n��f��m@�$o�o��Zؼ�J> � V�M�`X�� A�0���_B�y	$Ƿ�S�G��㦮���kDy����Wi���*#@K��	k��������X4w�P-��pd�GIaB�3h�m�?�p�k�BZ7���)�Mn%�%X[���%�XoC��]A�1;��xR�}F�+u7�cI�C��py�� ɭDv\J���3L7r�.����ߑ)઻��c;���g�n2"9�@;	���p�j��Q8B�osgk��S
��Y��W�B�X�1�s�'J�@^BKSJ)ۺ#B�:�3&;磵��L��\�v�INQ���6f>Y h4\Ӡ��;�۽"��EƤ���҅C�5�R��HJ�;:��,���/�\��_���(f|6�D��$$����,���t�ߚ���hxf���xa� @��R�ֿ��i���q�,nuA2�I�U�v7��pY���:�Z���G��8e�Þ-O�{���)�[���P�;��j����7`,)޹V)wW(a��tp�g�wm���o��F����~H<�h�EdAX���&��D��^�٩֣�8�ߊ�U��D�����jKz˲Y�8�p����[0o`���rq������O���R �ɾ�VI�Z@��p�p�6:�;�J�z$�������{��6����0���n�E���n)?����y4�㉗zGw�s�u�@�b��y�xg#�.����<7W��lnE�O.�*Z�!}�/s�t��k.IOx1E�|��o"y��݅�H,(���xQ����a��%<���66T҆�ƒ����:��jh�n"5#]�O��[�M*�PA�<Ç=��ӎQ{H���>F"߳��~��]�r��UR �rf�Sl�;�������5FOгktG��bs�ɪ!.f��Fh�*��a-Mw�^u��}�X�M��6�+�l���1����n{%�����xڍ���i)��1n5�o(A��KHC����|����ƈ���à��Ieޜ�{�����~"�O=�_�
�5�U45���Tf(�h�\���0�.Ǟ�'.�U��&Nc���#v��ј�:nE8�ќ��s~-AK�vɕ���̬w[-%��C�/i��V\���:Dl�5EJ��7���V?�W��>�i��ٌb��w�!빕���4}k�G�9ꯗK<���@���,�@D�T���:��'��?��<��?.`��j�0�tqߚ�wV�s��44j��邤�6���j�%2l4�{���9d�W\�T��lnY'uٔ��߆ޱ�;	@�	�$�g\ht|q����t��\o&B`�1YX�X����X['!7c?���9�L(�vVFZNvm*��r(ð��g��N���NX�cb�yB�%t�����,Z5G]�=�u�Zob`�5�1�c��6冧Zt�)�F��c�G�v�gl9M���Z�Qg�.�i� ���Pg^���GB��ue@�S  �0{��P���8:<����\�D���׫���*�j�!E�	V�0L}n�R]#��8'?�D@	yY{\n����%nB��V�s��Gn)���w߆4x��B�DH�4�mX��J�&�5�����.\��ڟ��8��X3�3�k�ݖ�����j��4ea��Q��rL�A�Xo�jr��y �0�k��I�Z���U� ����ÑP�$YX�0��qF=��LI��<�Iw>��&A�RY����+�)<T{V����L�m�[C� :�)'7L(!{`(�C�/��̺�[�yP:��n*�ũ.�'G���H	��a�<(a]���n:'��l<f*��'���J�9�N�ۡ�a9���
~�
~�(�xt��ۯW$����	�I�����^L]�QIPq3�u��W������x�ǌÁޤL�e-!ō���RM�x���y�I�Oe~�ן�#�,�N�4��Ւĉ�x�3v��t��
����[�<zɊ{d%�1�������B��ǿ�DGw��[ݡ�YT�!3����2��JW��]��h����gy�%S��i�c>��W��a�����"��S���ϧOЫ�B���F)HxXĐĩdo��7э�_�ԧD᤿r`�WN��E�V$ɁE�մ
B�U(����P�D���uY�cIU��%r�Eh/��&�c��n�	@���C��Tط��I�{9�|��uG�� �g�e�,�'���s�� �2Qs>�^��Y���	̎ɹ×��n�YX�@)�ʀ�p�	���z\�w # ^�ݞ6�Hb��1�QOƍ��A^�OgRh��g"����KD�m6�����V����V1�*�c��Ѣ;3��+�1/�/�ꙫ�q�=X��4	9z�R�>Ԟ�6䆻x3"T��e�����m�:y�����N^���M=���/b���NL� �D�&�H��֒����}��0�q��=�K�P)YV�Rs1�!�����Tō,}�S��k؁ ��35	- =��EHF����8� ��=��e���qބ��/�M��J�,[�\������>,�o�����J�Ջiށn�V���o���ӛ��%�ºN3A� Ȟ�b*�_����~3���T��i��g�.��C�۔^���Iˎ\D5��I���^~��b�6�ojeo3������w�����ˌZ��G�Ġ��?gtLšJ���s継�V�7.p���Pk��>�9M�~��������WJI:�E���m��ݫ3�b�
2U��Bϝ��堸��,�nr��d��J�q�(p����@m�dn�+�#8	qd �gk濖�I7�����ln5~/���<i����3�0g��'hzab�.;�"\�"��m#���-�v,�K@m���o�
��Y�n�;Se���͖�,����tV
v^e���=��1��k;��w���,�s|����ZO�d*j���l}�x���Z�3�S7it �����ך�$ޣ> d�y�����U]���:������ϋS��\x��.#������2u�5�Xڕ� �ɫd��f1A�f1-S7����O)&�0y��+W;��܏5!�g�0q�_+�s��׻\���e��Dص[���H,�]��In�ro7�~�+�A��'\]&��Uq�J|-#��Sr���zÝ�w�,̀p*�v��u���Uh�\��;�~Ċ�ej�-���m7:��·�L)�~}�1�4�$R�FI��de1��տ���6�]���_v����ԁ���ޡ!���X^P�����x!��4g*"�&��U�|�H���=U�_Qr(2�w<��n�}�@��q�n�#���릎1�q�ڧ=�M��� �N�Q�쫎�%B�[�]�`f��]��:
�W8�>ҌCr�K<s=����� ����~O�V�A,��+�0­)���Ύ*��)yk�CUB�c�n�n?ֵ���=�A#}D�k��
U����10��U�!�!��]ϣߥ��#��2��ͥtZL�#���a�}���y�Y�)����]���h&�m�Y3���nv�}�X�8*e4���4�P��Tˬ�0�����ƹ�Q��Yl�+P�$����^���1���;�fg�ܲ��k~ !����	��nF4r@<y�K�r��v��p�ke�;�������n� NY�H:��NRvBQ)�U�e �Qo>n^�#��r ���3�퍪���[�"��2-��BG-+���Y��<)[�̿�0n5���眘c���� `bӛ" ee��U����%��� ��Q�W|��E_`�Z��`�]>��aj�8��A�ͥYc�ͥ~R<��kF�OU3F`1��?I�_��y��q.T���U1��5�*�[|`�i�y��dt��`�ki�{���Ҷ(O�`>	5W���Q�١���Q����L�և�4��FV�O�K����Q��R;n,ˉ�6��[4l/��ǝ~���X�I^g�e[���+���@�Z.x��� O���3;��)V��|j�(����޵�4�ʈ@u�KB��N|�P�'U���*������n��u�5�)����0�$^]����C��k�� �� qF�?`��a��r��P�^�#�@ֶ��a.i�k~��3���K"LvsmcܢƏg�6I�颺�Su���O�����es�+VlqO���sP���eyL�-;Ԡ�sޗ���\	V۱s/�հ�3�#e�A�a�+1�j�JC������M��Y��j[��!ixh��ߨ�������a��9��f!�i�xl���rL�T�a}k���Pv�Z%��;L�0����ucytg�������*�`-��YT%�O��v%c�:50.Tbw¹n��uW�[ϛ^�Z�i�y��c���·�f|�oZ����8������{j=����(�H�%,�>�S�����\3E�^a�E�7¹1�����b���`/�},��?�ݖ��1]\�U�6�3ZZX��ӗ�B"^%�C��	h���#<����,љT�\��M���-R��m������0l��ܒ�!d��)��7�z���7>���%�0C� #�oR�y"ΰ$����);w�S�K���j��/Ul�4>��{}�DB[+��-5oƫ�!@� ߤZ����sI�Y�(����G�M���`�Y_N-ǐ��:ꆩ�A�L���쌌�����C�	M��t�Yv��ĖpQJl޾V��򭬢�V��?�!����\�P3��)�O���f�ՙ��j�]�̛*؍h��<SƨY���RN�w�Ixe
]�	"�}2ב�8���Ha��5:�+"!�H<��.Ec9�}Z�ڮ�mq��i�z���a�DC_��ړ��P���'����������"F�"�16�\�*^�X���Z�ͤ;��N{�٩)U�5�ޒ�q�Z�,��F=��@�H[ξ���h:.yrP�w��>f4�1)8�\�6A�g*��\�B�Ȗ�w�)$|�7��y�n��&�eY�:�S�p�}J���g���$$iCn��c!/Ӵ5��Q �[&"6�c&�(=L�����aG�e�]ܡt����}�ž̠{Ҙ�BD���k���^�L=�4�nsz}R@�y���.��3��6���6P�Ci��y�9�Yn�-@��-YjL҈`De5�OxK4L1�=�I�/���N��_���Uxw�7�����t�]F�Q$�f�V\���	��L���t�n�2��%^�y(=) 3"[B^��m&�a)�Ҫ�!��FS��\h�O�($Y�&�C�k��(�--���I��t�_�X�7�G�f�����a�$�Tʑ vqS9�@�~Ni�����weSM�S�=Tv�������v��b?!87�(�&�1���+��P�2U�$��[�dH>�Y+��9	
��K��+�!;X�ũ���S)1�hm��
	gpRgP�8,�)tWh&���y��{='T���(����:�N��|����c�����O�*ڞ̅��q�tMA�Ʊ����d 5J�ע�)������~��f�u��&������� ��b���=Q��q_�ⶱq��S�C�7��u�N/c��s��|�!�.���]��\zn��/��3����噢�|,�������$������ C�O���&tś8GCnV�h�v.��"�i�հ�v��X��L�Ѡ
�G{�m1�7�MA{��o�p�(W���y�M�>����=��P
���@�zM�/m��A(؇h�*��W��;���ylS۸�� ��}nU�8LvP�������A���Z���2� ����;)����21 &��tc�̈́�u����hYW�\�#-�/�<WoA�s�3��Kx���Y�ȟߣܳM����xn:�I[�
{p�U��s�5A��cҐ��M-��d6A4ς��}	KY�jYX�hk�7�m�+�t����Ƙ�Y�X��Y����5F�˷�����XJ
�����W�b�g�-3k��s�R|;j�0h�
�J����r��j�x�����{��8�[�n�>Yæ�g%�|��䡘��Q����J�!vۙ��{f�YEe�alZ�*Ms�^�Èօ@\��j�K�Q�B&��i�ֿ�!��}	ǁhS�8 e�눒�:�~�6��~�h75�Ĺ��z�썯]�����_��Z.C�Tŧ.���ŕ��?JC5u�r�-��쵲r1�n�_�)�,�����0:9�X	I����Z�V��Ъ�9�a��%��9�W��#��9�mS��J8sSza�ݳ�����Y�bs��$YG��]޲��{zu�`'�(#j��@zD;c[k����VS���o� P��%�j�R���p
��4I,f�r���(>Y��J�7�Q����'�	Rj�m"�s�}�O%����X��G��Y΄2�s�+��~����eg�i�啃�	w>��,�GU�-D�nۭ6���?�q)�-.�쓫�Ny��*Uz��b�;o���V$���-��!K�~}���h$d�����jϹ/=\5�����R7�< n�`�Qwɼ�����az�6�uŚ_��j�8RV�l>}%u��{ZSC�]'\���>�du�^rr��
��R;��P�?D���ծp�y�|���ʌ:�rZ0����@9�`.? ���/N��VdjT���)��_H�a���ɩ`����@�ѫ)�M~K�1��w�4��뷉��|?��)�	�	�܀Y��Pf;6�jg�ZƯ����:U��x8<x�-��!Ϗ���(����4�\�ql�".7�S<�9[��q��`ĕ�V�m[?��<����mwg���y��6�樊�������\/56ǯ������g�̽�ua�r��"���b��/�2���}��r�&��l+%�#� ����>��8yY��A��c��#Ʉ���2�׌��N;����\s�4�������c>��)�x��{S������D<h�L�}���q��?ۓv���vD�~�"bU�R���h����*�2�{k�ʹ�`�'�?$�n�Nک���J7�=��x���NK�w��a���	��v1�TK���O7���,��g���-w�H��5�����_�c��
�L��8��"�V����T@,;VZ��a*=�����P��G=ဢ}J0��X?F�mg��c2)��cW�ܔ�����+aT+P�pHWz�uS��J�4N�Ή*s*�	�k]=*�*�A ��=����-�S�c��c��o[=�l�!��tg�E.�#�K���C2d���.ԋ���pgbK>�U���8IWJ��=)�W���l��w] Ϛcٸ,۬I�B]���9���nk:&S���!pƀ��2`=��kJze���gB'@���?�jW����pAI�\)��ʡ�Xsug-�",�N7{�Ҡ�]�HnU�Bc�$�U���&�������.�I�:aM��wK��!V0�o,����!���G����d4�C#ZPk�YP�`��!�C	���z|i���^짘M�z�(N����l$�E��w�G���h����Jh taT��'�U��G��<5���dxf�mD��M�&�~/��:�m����(S:����x� ͧ4�.����_#Ύ?g�Ȉ�VˈcO��^|#����|oX���F��#�B���̯^�h5NN�d�ǿ?��$A_���L#'�8��	i*������=���Xu�}y[��M��N�d�ᜢ����2���b�Q{���a�Ν�$zy�NrMcw�7la̓@GG�T�|�(q�m��o�$a��m�b��ȏ¤�{u�&�"*�<@f��N�B���1�|���p冺��"�-��֐v�gzko�.L���TA6�Ԍ�T���/�8��o�u&��Q����K尛w�eՁL@��~�/�wȒ�M��{�C��a �IõU���ې�٢�*����o՘E х��p\�7\�:rw�	^7L�r̂�����e*�E����f���J'K���� �'A6�����y�Ֆ��ڸ�y��{�����X���E��Þľ�g�[?!���'�p)T����o��"	�U[�Ҳ�ȕn��|��5�Z����酹��7qn'��d�S�ݷ�8��a�` /�� �N$!�\��5Wc���˔�#J�k���.�ڴ�L��r�z���Q�4v�7w{uJwԽ3`OcW��ߧձ��G��M��y�vNp����|�񦑹w�8S����}p�6�A(:�`$l�@[�U��d*��d+Y�+������)%t�_�	��4�z�a('�v�P�,C �&g����R�� ��߬dP������b���6@�6�|)��q�u��(��s"en�#��r�V��������s�������C=7��̶s�>�YA3;��6o�XNV��H�Ã����r�P���&RO����Y�?��^^G��L/���UZ����}b/�t I���~f�qu��;���+�F:;�,a{_�N��'>'���*�xo@�/a�Z�5��HҶw�T9�`�ƭ�295aBA��	���|�9^�I�
����R��E���|��<����]O/ZZ���|ss<>:�	�)�ۊ��$�{�q֩j�o��*�Է�sJ��,�ua�i��'�V
9g�r�=N���)�]H�U�c�=U��H0����G{t:j��i��W�m+f��X5d��i��j�s�?#���~J�~C���Ûiݼ?8є\1,-o@<�<�"�K5"kƘ�H���2Gc�
f�>~1ḅQ���˿uq���ֈ\�z`��>SI��i�!5���o{���^��H����}��yi�h��>�7�]�����\�{;_D �&8����f�#N��$�J��g��I�m�V-9@;J������h�xx�5w��Q�S��q\� "��m�H2S��s�ø�_	Uq��i��4bā�%E��":�8?�}�8A�C�_��3y�1�R�l�b���iל�B���=�w&�A�j�|�ޚ/�<BB\S?H��uL�*�£�,}��Pm�w+����h��1O3�����f��U��){�P�0� r\]���� �I�RF"+
=O u����դo���?	4�2)��)k+�MP����<HU_}�s~�^8~f	����Ζ�o�
+��w6�paC�LG�נH啧V"!$�ĺ�7�^ۭ̬��I�a�,]��1W6u���P��=�oa�bt�=mZ��J���XԦ"@�\S���	h�KLv�$h��	K�(%)M�'�G�������I��ùB�i�����j�A��9�Nk>�#7Iv"�}2et`���-'��ɦ��2���H�9�Ќ�����>�㻟^-��h9tOxQ�kb��������S� �?1�_.X����R�˩��&�?K���D*�[�w�p�"5��"ݿ_��A�=lc������?����劄g2Ki�X%�"��PX7���U����2�z09���1�W��~�ڬ� �׊HP�d��D�Jk��D ��w�{Q}$�d'�?Y���c�̾������S���;�wCwgx-\���KCHH#�:o}�x�󕕣?���:�!��s��?1uF�^�{��^~���k��*�_ �G�<�����v15=��F	��v^P��p����4�:bZ-hQ�mpo�=��3k��T����2Z�&�\��z�v���e�g5WsF��[I���B�e���E�MA���U:4�}�^�?�$�Ds���q�H�\�~6�$����L���")M��
͞�r�=A E˶�L�����[�xQ��
���i�2�Æ2X9����o?ޝ��;��o����3�ʘ��@�U���QZ���́��)$�����!�t�Q
ۮg�L���4�M��O~i���5!p,�Yܹ��nln�XT�V��7����s�b�s�Ъ��ㇾ#T����^K�ĺ��%l���y7�{�E�(���r=>���Qu\��@����-.7��Ix�Ǖ��`�A���߲�&�����}���^z�r��i�r���U��jxx�����@Ɖ!�$AƱ{�`��� ��mn@(|�0N��{0m��o9���T�}�7��n� c��G�\Jθ> G���p���v�|�3��xf�Q�찳0���}K�k�6+d�&@r&��7�S�<��x��n#��5т�Ƿ,�{���k���w���px�Z��.���Q��ME�&ᶢ�d�����ô;��T��2wT��&@Y�ȷ[:וɣ�� [NT�&F���-q��9 @@kx�(.J%���I��ր�����t��<U�X׼��R�u��$SsWm���.��L9ƭO%��������������5��Jq
13��m��|�+;�4_���01e 
ÍsD��@��K�T� �X�l�_槳���U�y��)��x�r*-�vP
���I2EI[�QoD��p�E��t�Q������-/�;\������܍D���/25ȵ!��l��r�ꎄ���!zF<��j��	q��A�Y7(�D��Ѯ���,L��w���Y��Nc�xQ�v�﨣���|M��
�Y7���$B�E�J�J۪=�(��o}�*H`>)��&|W���{.���}d��/k���L(��%�h�(t)���"�v,5�z9���/`�Km�]i�f;��E��&1�|����7���bW���E
0��~%�?��K�6d�X;#���([ɫ;W~��.I%E>��H��J5->V�g��P�ٚ덤\��Q��8ƳM>��O�X�(�;/1N��Z�!�cqӸ�N�f�d{A��C��N0���� � �o� ^�:k,u�kW'�d�!��ߧ���Oó;�~A{�}X2F�d�$VoH,ݾ2�5 [앲H��U�j�=/T��ɟ����|fQ*�7�Ώ������r#[�H�N�Y=Y%.N���,Zq���i9?���X���ހ�C4��,U�}o'�?�7���[O�G��'���J��޳;�j���"y�����)(o-�Ih�C"���h���2�e���E,de�J�SۭnV�-�Mt2�}�q(�⩂�{�0��(�Hff�����d���P÷UVG���s>.ZV�����#�9(mZH4�/U-ى�N�	G�F&;�6kN{�.��5Hg �R#/&��,��z���u߿�kɀp�o݄���G�f�RlT��O`c�˄�h��r�_/��n�3	2\��*+73]��i6!Hܭ���[��4�7%����F��P�<���Y0�mz sFY�>�lK?�P��3�`�mT�S`2��#^E[���(�jr�,V!Z^�2���7<y	��@˸�qV}���cO��o3|�J$+6�o �ۣ��	x��Ϗ�u��ŠsM�u�����{�o>CQ��ofRB����M��[�&��Χ3�_'䚅��~��U^E� z��|�Q�ƀ�/'Y~a�?����͠���n��g����/��E�I]����\�����L�y�0��E7�:�c��@��ʙsp����	r]���y��ͣk�� )!�+-�3 �i,�	s"Ф>�&�vȑ�	lM$���^����0���E\���8�x��1'�R@V�L�����)([�~sLQ�Ecu��~��%��ŏ�.d߰2ޖ��Mn$W�m�;� cߚ��Yn�(p˟�I�V��g)�l�3����}ެV��\����
jɍ�O��z?�>_@��(���w�ъ��{g*���z��>Sx��\DILJ�l>�c�tfԬ�}�`��bJ�{��ǊbWAÍzp2U��	h[�8nم��U���ˬ��|8U��:�����3A[6M(�鿚rA��ƪ�#��l�B!�V�t!�¦)?�d�������h��j�h�:��;MX�&KdW�� d��L�B ��/L�nQ����2����ɆG�A��f�rOo���Kf��}N��N���
�q�n�Uv��_�� W5��rߴ�[�? �v��>�H}���cU�|��-�M66͞o�B@�F��<C�c$9�=l�'^����殪�(1�˝����� P�' '��n}v�8sEu5x#��1��ez��n�C���\S[g�k�X  ����i��k��q�q���5�SE�@��@�m��}YogAfB���$
 -u^E���Ԗ���713�Ų��G!g$@�ZB�3�'�pz�vG�T�`s&|�Q��;�6��2�d/���|
<���~��ŷ@�� [�~��ա��xWK@���=��O�����>�ƹ���fɁ(�j����Fv������gSn�S��)���l�ai����H�K|��޺_U����R�2o�`	k�c�r7>+;�ĺ��B׳�W�{M�?���"+_$>�@L�$%�Ɓ�m�:�8��t��H�`�Z���'l�Tyᜢ9�Xv> -P5�$���B�L&�<���
+�A�
�bp��93��T���v�P0�i��fwؑ����P�¡�di�����H;����p*��b=�p�m*˖Ro���g>�c��0�$K�	ؙ��+��i�8(:��Y�#X�k��O���Y"8e��D6�B��!#�,��°WO}E�8���ro��a��8".�&
�̲�ŭ��t���,id��Z���q�������r��4���}<w<��I��f��"=Il���-����,���RV:����N�`��W̃Ʀ�Bb��6i��u��
������a�� ��ET��h��0���cK�*&��!�Y����M�,rdh���r�̺�bBf���J��~A���藔����{D�y�+q�������*\�^$��ɰ�'G��������P@U�������Up �kv����X4�Q�>\V���uF��W#�#{
>h�79Z�L�d�h�C�¼�!�R`}E�ل��t�Ps^)�Tw��&���Ĝ����X1�X3`��Mr��{�+F[�7��K�n]��P�����R��5:D��'��;],�z���E������<~��Ye��z#��@�?oO\���  �w���Qoh��\����|$7�=c�'i����|[�ѧ�1�vu��I�^u ~�)3Q>�ܿ��R�� 4R�m�)�g"�x ���0	{�vf�>�lU���`�����X�.�&O�
�Z"#!��$N�~ڲ�g�O�Q+�}��^R�������fΜ�(��;D�靵"��:��U��<H���B�c�d�`�S�$��"��Я�	T�3HW!1HH���Û[�Z�HI�E�����&�6��9:p'|9J�	_=gy'�7[�9���W ���$?�V�t�Q�vڶ�t}�'T]r4ƾ������R:�{½��)�/�;�'H�u��N�!^yn�.��qۯ��2��e�pk��E�t������OSz�-���FT}�Xw���3Vv���Mcn�ߒ�+�:�I#���c~f5��°h�+�5�0)�+J�B�cA�JB�U%�'�`�л��5L���D w?� ۖq���^��+��jU�s�*�� �w�	$\�g�����U��p)���g����5PQ��\,�0ϴϩ�%E̲�`�]� �+*��m���}��9���Z00���S,#����0�)T�2֩JZB�M1���Ďj�c�|%��|p��9�m6�-�s�w�5r�6Au���7� ;1P�$r��h��G�
�Z`kߙK
�=i3�l��-b�|.�P!�!o�Q��� 힚w+��2Q��AK��1�P���97���D�6	-J�0�1�)q.-w�T�BO���xCo�{;��W��S�
ѕ��� ��F�'�B)���L�G�z�!]���~X2�Z/�&'xU�P���ns��"�f ?Yf�.d"Njq����J���V�eJ>e��@
"��;z���O��Z���t`����f�"���rC�}4I�d��� N��*���p��=(g�[@�O=����~�a�um�f�X,����C�X�$��T��&�?���ɺ�����S�[�1���c)�o�<��!�p�3H��N����]Y�4K!�}D^�׌Q���X9v������f�HVj�,3 T�f���T��V3�?�_jD{��7[��o}08:���?(��Hϔ9T]לW��<��H���L_㚔���B�@r�)���HT1��p�8:��LXð'�m��O���s]b�%�u\�	�F���y���X1��c���y�d�Y:Q1>f+O��q�����3�r��b؃|�;�u�c{��m�F"D����q���ůY�(Axl�U��ݿ~�i��JV~�^G`��2jg|�'���%�u��\��uO>uz���aT��u��"z�6�yх-�{�Ds�����;!V�i�S�l���j2�vJ.Z�)9��{�ð6;��� rc���r|0#��NH���v��x�m���f���&���uSt.N�3���s/���Rܨ)6��1Av�}��шUL%�ӌ�A���U��ԥ��0�t'W��L�¯�>�ۄT�3 ����M�>@�-(�����jr$ �Y3��tE�����E>@�Qb�qQ]��A�/���U��a��@
���c.�Щ�X��&����WڡEJ�Pv�L�v��#�ɏ7M�B�jR�Zg۽7(��N�a0���������>���)}��7r��7n7*�,��S>O�D�'����(_�Z�j��4�44� �"�3lG�LꮵF$
Y
,j�"^�P�	a�Mȑ��8L�-�s5Z=P�6W/�4��RW�%��Ss��k�5�
drQ��L�Hh�pĨ��W��$�q"��f&�HR�Lٷ�[l�-V����lB[c�OK[�G�Mu�2�q:�8�X�og�Ό��:���9�TW}'��3�K���Ê����-x<����
.��PwP���9�/k��������%�{}�'g$�G��B��>�ݐj��tqӥ�Ꮲ�k_ė�d85b>|��Y�����0�lyG�C��U<�d%�p�1���9��i����ʤƧ�v��,MT�3k.&e��5�cB�5�D��2��6x`��G8DQ;�q�s!��5dO�^
a���/	 E��;��v|�}gV�j|�M;����d(ʌ����*����N	�
����l_K'�Ռ�4�Z�c6�%��4퉾A�ID�v:ȩ�۫���W�+r��%���D䜪�]ÙG����ٖ	$>F�T������������&��� �n����pHyxܐ��%��!p��\D6�y���Y�H�NJ�Vs6�񱾛q����0��S"���(l�+^�����=�G��*_
<�M>�E�U�g+ih��4e�;����O�tgUG�[c?��w>+�<-�v�l�M9������Et���
�Њ�7��Jk�˦�J�q"Gt���^�~����r����X_�P����>lff��)y*E1�ּ�dp�Bn�D�E;�j��Ԃ@����~���G�*�0�Y�I��uoH�"��(�*U'w ���������*w6�k�v���Κ_
������M�Au$�ZG��%��s�?��"��
0��:��_��~���o��CV8�ڤG������Ah�\��Zb'4\�,��~�/x�;"�JToS9J����^��/!��N�6�'��{���z�g;�hFH��x���ʬyTK|��ޱ�N�z�y���T���K�idO�D�w��/e�G�h}��ڨ�~n{d�K��Ӭ��ܳ1����[I�V
Rj9�X���\E�����"^k��uu@h�� �� G$��u�s�E�|\"�P��I��bKI;��
�Y�Q�qք P�sm��(ԙK|����
1��/�E��?jZ�sC�=�xH7�fkVC���W���ώ�VF�q8	�qC�I�L����:=�D��)�sZt\��|G�*2����W��Ù�D�I)�n���U��`�ȸ�O�)��6�w���ި��Yٮ�X�o�� o�OT�ˊ.>�ˣs��]A`��[�ܗǽ�]l�$K�����O�80vQ�-�7��p���$��!c� ��UCW���u��t5�Y��IF��b��pE)�	���M7G��@&P�h��ι�x1�'���L5 ��j�׆G���vN��8`4/�m��Ű��7�@'$��5g0{3�w����	���4%)K�������WJC���7,d����%Yz�ӷ��_����p���2���[�>}�0a?�{4�0q�QLaW�����RWt�6���3����J�Q����#U^^�b)ؾ�f�<<K�69��m����^,JV��vH},Z�ZL<�-�s�F�l�e�qe�(Wgo�Ц�fZ;\�xg����E۵��ճ	5q/7�*�����u�1|�8|8�4�I�I8��S�_�,����Q�?��9���\\�@(�ȢW�����Ϩ�C�%2X���2�;M����MK�oJ����<�Ú�V3񋾌=@ �r$^�)�"�(5��X�l�tA��c�����m��͛)�n�i;ӿ��;��@Q�bʐ荘L�N0�U�q`j�v"} 0��z���ڰ���Y�$Ȉ�����R�Y�R�󇴕!��+$��DI%���#�7��8\��$��E��TF�K����I�qT�[���5#��,��ɳ�T(���7$�����*ɘB����z����-ޫY;�cH����2��과�/36LL�}#�wNS�(Ԇ �͢�'j�I۷�l��J��5b��!Q蛵��|�O7�:�}~v�\'74�g�-1L�o��z'6�-M�\���gX	%L��0�-�.�|�{yհ�xS�(ē{R��>	x�h��\���m9���w��.�Ҥ*%2���j(|r`̣��}��6�}V��ۇ�2�[��d�zg�=Q�+
}'r��nLꣵ��(�*.�s����Q�gI�6TA���Wr����W�):y?��JYi0�	[)Uy\a,��\����-��}�	hR��]S�X���3vH wof�v܃m�ѽ+���7��;������TU��`|�(j�� >k�>L�~ ��]-;A>��&^�ʲ?�vь~CY�g�r2U��g��W
c�@�!��q�*ȩ�RO�a%�X��N���)U�*��NS��Μ�	�٣��VB�L��Y�nf��g��R�ЖA�v-kf1�̍����E����x�N�H8g��-Tq�̍����X"߄[� ��f�RS�Z0^;�#����k�4�Z�64b3��S��[��63�M���WEW
��n�S�8�ς����~�v8�i�W��F��F�̌�_[:��Z�G?���1�QA 2����k��nLYN����Y�5�� pi�Zyތ�0)Gz���y�!���=��WA���X�c��`vO�y�]#���Y�謏�`���D�r
>��i8�_���%\���x���zG���¸��d��S�>��I�L���s(�ی�����n�ʧ�|]Q�r�U���L+�BF�;gU�Z����������R��P�5]�Ĭ�"�z�����/�|56�כ���E�S���\EvlxK8�4�Ř���;m_5jByN�#��	�l%��	~+$@����C�S �h�x$�2���R�$s֢)��a�&�R�� -;���݀l��X�8�=�μ���G)ˎ珰n���<���8F,Yb�8c�ky�_�T=ފ�� ��"��5%P�x�_\4qϭ�O��>�E>6E�Sz��{b��[롪f����|M�i����ƿ�z˚�У(	q@�л���U���2M^1�ZUMq:�Wx9J��_�D��o��TJrI�D����H��vǢ4��Ө�>*��R�$Eagh�l�Ƥ����+�`����W����X[��E�)�W0¬�%�aiY�$;�攗Cn�\�|�.#��Rڍ��;����J�&����XF�������R�[�ߵ�������j�	�iґ��oN�xj~�I��eQ�{�D�f���o��N@�L �p��*W=����Y��w�s���)=ghӢ:�2ED�pSY��1J �F:t>��F������N0�A��ot^4Y%��Eo�D�ĴA[���昋����x`sUW�$vkn5�칍R٩t��4b�f�'��`Ū�������&"��Ěwzm �8�B���T��f�& ��$��E 1�h�jф)���s��Ƹ{�0e��PG�`�@@bX��r���+� vh��d\W�H+���5��6y6%<In-���_����!��͘JUy�~���M�0�̘E�^��e�X�x8����S�	us����g7�]�.��GL4�_������2q��$�e\�-����]����3��&Ʒ�Mu�X�|dZ�S��yN_���]�����JW����h���)�h�MqK��Z����3����2�/����1�ÆQ�r�v3dCdep��aT�	Xτ}&9�|ɺ�&[�?�<Ү&[E��|Mm���/�o_�t]u��K�#h���(�LH�:VT�����P�j�dw,uܨ!Ծ<�$)����W2?���߱=���J-{��L<��k��prŞ��aߠMhB7���1w�|S\$RR`�k�������+->��T)���-�F�O��mॅ*C��R�X���}��p��~�M=���W�]6Da.2���a?�����4�(��ǅ����;������pɣ��L��[���5��]z-������{|�ru���E�e�TA��r�ѯ�a=}���4ѽ�z���P��>��rV�P��gc_��I:m�?UH��Ut��c��|*;.���K�&�d(W��g.���X�%tA���۳Z>b��#��(��=���+��c-�����Y<b�R�҄yc�"��-}�U�$;F.%�)u�Q�.Q�}�|UV�xB�o��5����7-�mN9�6ŝ�n !8�΄8���e���_ 
�0��?�(T��<li�P��]�ez�Y��j}�|�$9͔��
�X`��=�ϪcY��p\*��bܚ&��ù7��Hw�?�
O�OO}]v
՟��mw�G�2��(8h�'�Aף��2�a�x���|�U�Ez�)O�8�p��|�Q�vy��M��P�I�V�qB�&�2��|>	�B^�4}��dKS�0y!��N<=�i6W��&4�|�1/�R��|��J�yt��B�ر�s6SC;T�l��I�X�%M����'�}��^�[��c��ٜ­��x��)҇�yD0�1s��m:�Ѻ���:G��E�8�L����B��r';EٶM��4��IiKs��z��vI�v��7K�g\����מ�	34��Ɗ��_U�9Q�c0�k�9���%�TM�뵴�����׍g)���E�-N��=���W\����]3���]F�1wd��Ku�SV�)�#�F�r7��#O��6�h��}���r��X�2�~�n�A�j yT�Z�R��a*�;6��0P�� �a̙�"0�=�l�z�����Ӡ�V]����i=��o�@=�5+Y�D�� g�]�C%d��Y��)&�Ok����U����Q�N�J�@��6-�$��F��;0���<�-j�zAi�"4<n8�s��+
9u��a�PJ��dڭ���Tk�"=���~f�%6�H��҆É\��K=f[1��_�WE;J�/(�^G�����w|�;X�e�Y���-<UqW���pM0wB�ѩ%��r�4�*;�z%Hl�W�I�δ{�L�n�uy�.ɺ��#�1k�G��jT��EӍ���l	�
�2
���9c�P�]Ք�ɍ�F�1�9���\�}��!��V�䶛�jM.q:.�}��PB�
��j����Uft���|�R/p�X�s4,rHa�/K�y�K��}�5;����G������
����T%�q�^D�3R�_��bVϕ�d9�  �k��ᘕ6+g�P�>��嗲|�pg���Fz�'�v�mb3�����Z�l�_
�xH�m%p�Ϥ V�[G�w�2}�*T(t�9=H�����ח�1��Y���oC���.�8��< "�ˮ��
���)qh��'Qk���։�0j�t��2	�$Y�P+"�s6B�#����ne�pt���-L���B(�_Z�rw�.�Ϊk1��`.�x��6ET��jѸ�J��׵����c��U����v�����I��>�LhF��չöc�M(��l���u������B ���$�,M�q��eʧY��������t�.��$H������g�x�a�Oo��%�RHJd��V;�!��4�^������yRAcDn�ؘiO¾T�&�)1��3�#�^+Va��ʍ�_JP�Z��Zl;Z=��A��t�2άd���_��]m|�.���̒��u_t��@�V�NLR�,s�(Qr��uW���1�I����MBA�x6�k����"�W�Y��o���PJ\�}��Q'��������z�=��kɽ��k~@�I��+��\�3��L҄d�jJd�㞂���ywS螂�&L���loT�Y�-3���~��F�s�lSgF�R�4�a�j�D��'�ns�6��e��{`0Fj��>�uU_P���+�����]$�K�9�kS�@�X�y��H�GA� 
�u��o��ݔ�>��j��F %��}�K�eq��T|�h�5�u�7\�>j�������ً�܆�B{����l-����#�͞��Z��:/4Z뛢�.R5��O!Y�B�n�[�������6FBi�Ꮶԭ�xX��bw���J%����+�b]5U";��0]��x ���5�[�@�hE�X��#����Y���fمl	U�y�uLJ��P��|!�X�-o�.A�dAf_қ�S��N��e�67�AG�T�d�];nx���&	�g�P�5�ޤIW
:������A昇��p��4��לNYh�S9�(��O�2��P���j��H����9�8���yF叅������{m_�S���V�9u(Wg�d�sVQ�Ӡ�6�h�t6�,\��DA�9Ú�`����WZ>�$aOtp$f��z��5��W@�sƉЮ�	�H��ds�M��GS��b�p��k�G�o� ��M������p�cP�'f	~�}��� ߻����E�a�!l�����������)�&:����r�/��Α[�~#���v	�m�������ϭk�<�дf����>Q�Z�����r>KYuQ7OR��[��&7����q�[ h�����)��0�3��k���I�5x��c2��c_SR��qi�B#�X����c�}� &9�m�8��3$=�u/6����A�lhA�Vi|��2�)k6�����2q��$ҽY�92��QS�,w���}�]^|�5��E� ����~?��w�C	}�(\F��I
��5GX�+�����芖��T��
�I��e�!�`���$�>�Q!�nƲ����l-�B�����=z��_dK�$�/)��; +��Y7偢�	4$Ķ��f��:j.�o�������Q��v�>�0��_P�a�]��b�ms�w���uݠ��K�g�C:�LYYO�G]�|�j����G�)���#���9�
"�����},̆��n؂{��VJ���CC�%�#fWt����P��3+�L߰$��m��Wn
�?�^F-���v��S3R��hX��Gγjq�P�95hb�x����C�hOO���N@�U�M{�Y���[?5f�ժ�R��������� (L�(]P)̾�`���j��Q���kM�X/�Xn�"�Hb�@�%{�j!�,�����a�8�S$f���N0����G	f�Q�0�n�,-7��jp/B]w�I,z~j��m i�c_��|�g��y(:�q�5����2W-�5����n��#�7���H	ډ�ȉ�_�ȇ���3�=A��U�������cn4K8�5�3�����`�$��y-��/�s��;]��];Ay������1�mNC¸/6LA[�g��ݖ&�>�6��C/�q�(\K�j��,�ͪ��q��d4�t���68���tk�e��r��6�v	�*����(p�\�y"�=��[�_/D��X�~{��7Č65���#����݅�Y)f�Q�>���@:�U�b��l�+�e�JX�9�l��,�e%^n�fK{8�,=�[H�&��Ƨ57�_�wAONMdH����ԍї_G�@�����B�=Ex�oZ_g6���s�jФ帉���#��u2�3��b��ݢ��Do��E��3i����|H؏���+�d/S�kB��Z�������q15���Q�h�7i�UZ��1ӿ\����%?W��Ux~�'�|�E=tgR���m��FCؾW�s�@e��Z��%�+!�f@3R���!&�|H��a�"� �"�����G��$�7emL�!��7�C�.�s&+. �;��2EG�r�
�H�����6+��b����!d��=��֦݌�K$��0�L$iz�~���'���>S���d�/�N�kl�4��U���N���狣���eA�;��AKi�sC�r��Gmf��z���&2P0���������R�Y*(�-�����U#�*	{j���"Ya;����XzЅvrR>�L��V�R��%�u�@����h9Ȧ(Xr����I�{��&��ǹ��S
�}�l��@� ��m�$P�)��^m��w�&*�W��$V�Ft��bs	��OpՍ�P�NC�i/���ra���2	�E��ҸJG��h��&9ٚ��]ƞz����9ZՆ��ۢh��,��fK	a�N@���D�J3�x���+��E5Bx�|�B��%j�֪��I,8�,r��\V��l�x�J�˄����V3�;7�U��=��&�֗u��'�ƣ˘���T������Q$�q���Mۏi*�C4�|OF)���٪�^�]D팄��U����_�̩d5Ć�pP\��k��3$���]�dK��'V�
�oPB���!����E,�Z*:�$�3�xQ 
�KqcQh���}�f�ݣ��#����d���A�/M���A[
BO�hn�3I/����o�#A��"�Sf��)���<�z�F� 8o�i���j�x�H�KUZ`����>�HKXE"M�[Z�~iPH��#R嫸��K�?���\����OQ�Q��� j�ް[>CaHQ�Өi�4���=�A�xQ80P��9Ѧ��Gz���d	��������Ё6&}8Q������:�`U$���z�c\U�{�XWnyY�_�:Bf3������Ţ���z� �j������>a�/&�p$w]��{�����T�������e%���Կ��g'V��Y�+m�^dύ�������?�K��6ͭ��8R�#+'��C�NQ��j�_��#���#��6�M߭'�n��j��D9���f��|�<I�#%ṥbd�����6E��clS��NU[a=�դ�i��V�\����R?S$��y��~�M�^I �G]�o&5~l�wz�n��%��Z�m���̃#��쉧�{���ʖ�xMuu�Z��FA��
E�����@�J�����j�)=���Z�#�_�!q�F�y$�l��e8�&<a�ś'����+7<��`���}�5�Lav�$ù�pj�31�1�-P�1e�8�Z�<���^�y��LS��ʀy�c�Z�x��1���+EF57n
^-�l o����g�E,��g��<��B�Bd,���F�䃲Ei=�G���`�vp����X[X��l䟡�R$��z�i��;ʋ8w#;?~��H�Ozέ(�R���� Ã視�q��Y!E�}��/���b_�\Ӡw��o}�I9quu$-�?M��MR# �������6]m|3m�Uӫ�Zt8�2�����W[Πi�`�
�a���%�X�4�}�O︣0�g�> K�B�ȏ,�[!�MuU���a�tUv*�y.s#G�}�oj�~̵\}��ŀ��6s"f�ޞQ9k��U�هn�� X[��$ќx#T��aER8w ��J��In@>;ѿ*�@�az�wO 笤'�,i\�Hb
���y��b�6��wB�k�*�A���9���)�bN9���q�2���Aï5�S�hPٙ�u����!�aKU�이�6p���J$3����������*�E.z7Dk��c.�pϿI*I&H0bh↟y;��5L[?���J���=����*X�r��Z>�=}�-�y=ւO!^���y��:R3����j싣��I��n!:R��0-x֩.��>N���݄�!�OfD��en�Q�2)I�/-�W���ë́�[��\;a\	���Ц"�*�F�yA�3\�+�u��l��^W�����Eb���3�{���<J�A��I���c�)����W�좺Qp1�"ۿ�As{"��Á�4y�)�����[�P���w8�����T�| �R	��L�9ThQ�C��3m�'��P����hYBHe��<�o��	��C���*��~u��P��nr׿n�`a3����N��e�/Q�P_��L��+ܔq/T?o3��D�bA�I%M����D��8�z'V�����]�#WI c�b��Q��.��t�g�)&�nN�b]�3�-��^k�c�"���%�n�⼅��E���G��]MG@@�-
�u��R]��A[�}����~�B
Xɟ��ǯ������?�r��H���T���Y��?�T�z�э��
BP '|�z��*o#�U�ΑuC�P��άL����dҵ6I>�jF�Of�
7�kn�'JI�3OF�w>J� ��̖";��ƽ:����c4�d����L��~�U>
9�"�V���y������6�������(�esy�1�O���.�g�?)]���xm9Ji��<�G�#j��g�-�W?]8�-U$9��c
7�X����!';�,;<\����b;�п�z}o}�{w�����%<�d��?3���R���Wq���e��Մ��.�����x�V�k�)K�T�X*�787�x�sK`��8X��f�3U����>�T�[Z�!�`Ƨ.o�aI��1o��Y�`��K�i��:���ƌ�vsxe�t�#zU��,:�_��7v �"(]�B����EQ�r��m9P�,���)g@@��q���4�ޅS��ߑV'<.Z ��j�\c�|H�Y<���.`�o���kP���I�
Q����PUK�H�7�l��+�u��r!ӌUȃU{�x�f
�ܟ�C\a�4��֝�J�o�Y� t���j����W����$�̥ ���t�Th'�;��OM�".t<(۽r9���i��Z`�;H�(�݁܄ X� �y"a�?& �*��+�wEAG;��GF(�e��}v�ƽ�)��҆�oJ�{'i�]X0�e�Ԓβ�qoD�r�$p��z}� ��:C��w�4�t�4�*��L�A�o<�E�V����&�����HU��"���H��P߰��O�+�kb1K2?r��GU��.�����.�r�f��[��`��7Q�J��9L�G��vb��C�,
��+�j�c+��D.>��<|����2��`c� Qf�tG�=@wQ%~Q5���q����#� L#'!�R�bFS#A��$6{uQ�O�2m�R�C)�L& �GXһQ(|$�Q��0#$�Cfx<X(0��,e�4�1����0�[�W���7�3M\ɸH�I��DV��'[���|�b�g3^�x;�sQR��F�0���ċ����2l�zm^
P��F��6EYpt�>&E��7E����9�IiDc8���3�k.����t��#�+�6�]A*.t;��-RU.!)��]?R���������q�r$��zH*/b�ve<�pM�Y�Uht$h������\���iwF��}�|�)�E����:��o�8fW�:��)P�*�x��¤U�!�ۤw�Fs:��7���z�)
aa�&���w�ߝ
ħZ��s�fI�?�r�u�V+f�X���d�PQ^���(==v�g�yU->j2�va�E��T�>�PHU��@��*�D��Al�V�},�ku�U�Wҋ�&@��wD�]GZ��KrMά� !� �R�V G�����eb��'-1�8z��h//s� i�,�1��NzQJ�M`h�_���_�kp�`����
8ׄZ]?��<�i���+aR)F_�B�Qƅ4�`*���Y(v<8�+ ���0dP9-��CJ(�/\���8�O�u��bZ�簪/X�,�(#e�'8�h2+@���@���ˏ
��dW�\�.�;w��J�Ő�`"*~��Q\�E�ZTF	�mܘ"�S?�gԓҸcB�^�;ćӰ�2N<9Fx���U@R�Úah��Y���(!4�pʚ -�| �s#U�\���a��wf��$L��&7{BS)-$�<nh"^Os^I���7!x��2���G3Դ?v��Č�m�#Rv�z>��,�bh_��,+Y-{�t$Pc;o���?.���KM ��2/\� �bj����0��b��A �=���n
��#���M�]ٱ+�CM3r�o��hң��kF)!���ǹ��f�_L�n�̽��;`���lPI��(;�������?�<Q{�K���v���Ӫ%,�Ԗ��
i�4�B�d�=6��I��?w4���DD������&��C����E����	E��@*��	XaL����/�+M*�~�Elۢ�"uo�I������M�vm&ǹ��޼��-k/��S$[��Œ�f������#�nӚ��l%v~��I�`W֖K2�*"��n%\i���-bZ��'l>r��_�WE3��nz@�d�u}�	�4w�	���{'�H�I���Tv�6�����l���!W����^D��e�|�?59�މ���K�����FM5�L^�i�b&��C�}�S'�-ΎKe���۾�Y!'�5���s�ʓ�5��m[y~E�P73"����Ds�YÏ'rX̓g��mKs�5�h�oЫ`%��`Z�[:Xh�p�e�*&�Z�ĕ�w�|�*�5��X�M7�"�s-���!z������T]Z����Lt���]4�XH\��`nV�P�ǣ�Op��)g�7�k?v�H�љ�Wff�7��1�(=S�@���U)�ڄ
��/�qHg���*wr���O ��I���[0:!��P!�Wo�qVp����q���U��h�Z
��+�>L�:x�"��`��H�HK�l+'71�p�X� y�{�r�,u%_�(Œ�J��C�ZV�gɦ���j�X&v�|k�=s�g�1?9Fn�n��Q� Xv6��B���"Z�Ǉ��Ja����(��k����?O+v )?��`�}�)kd�%Nd'�0����&�]B���s��K�f�+�������LEԴv�y��C������,C���%�-g��঺��#�SY�|�n:�T�Em�F�q'���ck��>��I)��Ꮬo)�^��[�?xe����mFq%�ӉNM9�2�,<��ā��XUM�Zds�5�bi�"W- ��ɐbf�k�8�������+
�𓏥��S��ǡŉ�i���r��"���Dɧb���O	�e;OۆL��V7o���:���#�`��;u��n0Źf�2�p���Z^w���c��F�B���K��_m�����	or�7��BZ4�F�(��I� (�؋ Ѵ��'B�G@�y�d�2PC,	������EMCP�>CX�.!�䒼��SE�Ƿ�
�4&v�|��sT������p������,�INTDKM�U'dLl1�4�C�"n3�Y��]�N/�=���P8�f+f�A�Ķܲ��ʎXs�0m\R�:���^�iJ
�H���%�f4l� L��S��|9�.|B����N� Bn��g�k����S�ZaP��̽��)�?���Ņ�Y{�ˤx�$�~�O4��S|b<Am;,6���LGr�̀𱊆{����%�Ɖ<z�ŗ:�;٫c��6��)�8���!T���]����Ye�IS��珤)��|��2��-�
z��`�n��d�,_�k�Ծa�s��'%| Co��;�ƥ�e�g�w�-h�$��1Gq���A#������&?�����/�I'�@4&,��5�ߖ�qdW��\��%KA_Ǹ�u�3܈�)���£7t]F� �p��\%���>ؐ�	ѫ�ڜ��e�I���N�6��ck�Ɣu�Q��hۜ�{2q�X�����xժ����f����;C�5R���˿A�)k����_e�8+�*<�+�S�s���Vn���GUS�6��%p� �WG�Mg]�+c��@� �b5@�h�Y�:�*R�v����p������$'5��^��|��xwϪL+7��M��<kh�=�E��u�z���<�#-��6��]���ٜ>�J�Zx?¯[�S�Y�m	+�A� 慙;��|5Y�Q��9�&�с�#-����,��l��Sd��
�O|F.}�	�8�:�8��07BD�f�ީ������&�2�(ڸWi��5�hF���g�#�j���FF��@P����r7��D���z�|����\�i�n��vBD^ݍ��\��C×��BpR�����*��?�����E��7����}��r��O<E��Oי7A�=�a����'o�T����"��Gc���~Y��)�p����ہ�2�0��Q�+W�P���8�s|evF�����Ɔ��=����A��~���Md���N�z��������J��{��XB���@Gh�.���yo����R{�L�#�!'m9���Pßz�k���X��H�M2R��[)�)��+�(�2�C��Wv��	��g��tƤy���������G���;�8<�C�?��N���I�#,���te]��ʞ�gٵ�-�#�^P����� >���d��q)��1T��@���T��P}Y�¢x�< c�:��B�"���(�<�߿�:f2i�P��3}B,=�J~��^]�&�����g �\����}]��k��Y��Js*�r�e��z	B�2��g��J��am~ч���g ��fY;���<��3ϗkm��E���]�[�G��%�e�L����{W+1��08z�Z9F��;4 |-2y�t�Gc�0^�����d/%*<-2��L�OȬ)���?�s]���''���NS|Ѝ�$��쮮����k����_eW�ʝ/)���'']v��ѦÅ��5S���kQV<��a\6\��%6�c C��;_����*���ָ����l��&�Z1�4Z��h�����Dy
��4�@�����\��]s;��ܽ��*���{"Yï�َ"��*�C�-tyeG-W$��M������r���1��it:Mb>�� ��4���FRO��q���?E��ď0����%4R{�#��!�v�?B_����Y6iِy���b��U�nz9���Ȑs*t�L���F H-[f�J6�*�3�E�)���+m�fX�i,"��V���"���}���tF��JC����*�t����_)\n�@�)��$������͓�\e
Q(NH��U>?���lt�U�"`Fa�"��|&7z��8Z�Pݠh#'Y�&,|�����q�g��sɨVX��	&���c׊�F�p䂍��S�\��b	Ea�����|K��^9�\���FШ���2aor�@u�]4�9�hW�U�Ƀ/�F���	���h<�|.5g)f��)0�*��P���X���n��s�I;�Z�'Q�b�{��%f��iLwLKS�4�PE�R�8lŮ�1\H��L&�f�mcVl�o�2R��˸1!%R��i�N%�E�j��n
���1��r&��GҼ��ǛA�ʤ�g�Y�bҤr��N7����1������Ѭ�2F�Bx��&B+�6*v���#P�/2��|7�|�h���W8��s��_��n���^N���B�z9���Q�$�
=`�ʳ�8�g��3�=l�JZ�i�?�
C'v'
��<�9L0�fc��w���@>�Һ�^���G��AR�aߌ��֏Ф�o@��jL8G�@�\4e�(&Z�|����0���D�˱���}���PJ�'*�f����!x���z|DF�rko�����a'����C��
�i�t����
��!��#,�W�jɶQ�}\$�j�"��4��ر�Q�Vz�\Șz��!o��|K{��-{3�.W��х(al�^���ֻ�K�xby�
	$��P<S-�����MC�,��;��aV��{W�$CM�mV'����~���h�����*iΝ��P�#螌�7���l�`��ϯ�%��@��K�k-k�d�A'�IQ��g��g�yY, =�#�y��}zXld���[}�����t������LO����P�..Eh����&\A޽��qi����+ְI���&N�٨�l.KֲY��f+o�\M�<�J��8j���|3�r��������r�  +�T>ļ��T8���Xq�C��CJ����x����p�͒�D�F� 0��=R;�8ʔ�y[|i�=�r�pEm��9[<h�:N��x� �cA���N�� .g6J�jϰ+�k�@����ɥWC�~v�!;5mj��<&k���m���"?Xk��!�08�mx,��B6w�50LGJ��mM�������K��LJ�Ļ�B�`,�L@܎�_�UM*4<ђ�N���.t"�E�&)y�"2�J+���H�`�y7���C�3�r����6��ߑ�ۄ2�=,>��<u�i��&/}�M���o�������vٷY�.�h���n	&]72p����*��b� ��$��!�%�13�o�)�҈��Я+A� �hҥӊ�~K���=������`�a��I��zu�?t��nY��WVN�=��(*�̓��eǱf�ʔD"�T�m�րҪk[[���D�K��;��ރ���������q�s F��d�2/��?�}Gp�A3��F
��I���&��c��ch߃��Q���y�3��6��Yb�TeH�G�@��'��ٲʙ�H9�Ϡ�lS�ȓ�DJA2�q�������C���6��Hn3��@7mX�Z�H�_=�������溵R���n�"Vp"=�-��˜� �}�n� m�]�ɾ���+����κ�>��L��q`��_��ݣ��ZN��/���Z9x���y;tK���v�m�����6ur�68���̏�I'{��Q�ݓ�c8y���G��M�~����E%��Iz�&!_\J/+�B����zm�7��0���$��8�7���^
����.t�&�!�kF� .j'�>�e��(�n��"_BF��G��\�Z�C;Y��⼊�.�!c��ȼ���Q~d�w`# i�x��.Hl�@����r-S
F�7��NW�@��/������s��{&"��;�s
{v8�2�%!Ѡ�+�T����kL�4�VB��*�D�H�k(�����0U��v�VB肍z���ה�������ꑤB/�6�$��; ��n���G�S i����N�)s�n
;q��͌6p��P!�#*@]�5K�@%��Z��b��ջ@���/��H�!�ݠ"R���9�6!#��NЃ=�Şg�+B����Fx__t}kҩd�넩 F蒝��$B����#?�B�n��c2����q��������A��uQ�:�)�+��I�r��٣�X���H�����YU�!7�@e�r�K��#�R�4_�/�D�@a�����>\�eS����!豸�j��X$cXXܾL�V�N��z���j<�.W�Z�P�7[i�ܣ�=��M��Q�$X�Α(���I>�H�h`1�� �o*G�9��1��"��{|ѿe���6�5����R�2�$&����G�*�$er齤fw3�V&<�&�Zt��8�jpϖ	wk����|�_�H 6�I����_��]��4 FN޳;��A���+�|��P�[�>�y�����b+;��A w"��h�A�/�S\v)Sȃn���t�G��T�;�!�r+B*H�{���%N�dk��2s� (Þ]|���E����w7�պ�W����/
uS�0e�����׽
aVk:3�-��dc�i�VEԇjN5���m���4B<v�_{LsA��ƃGO���Ũ��T����H��l�*ND�C�O#�Ћ�<u'�2�{�`�B���"�ȩ�XlyWY��藈m}���{�e=
�>@�ff�O�b�ɴ���rQ���C{�%�q�P�,�!8�*Gm�fZ�w`�FUY3E�fD�l?z�^��^�g6��5`Pq]=R��Q}�K'���`��) F^M��1�^ݩ!Uyd:��+�k����֕u���_�9ة)q!<�e�<��}�}�'��5�M���L��X�6ՀL}t��/"�^��eP�U�͑k��k�d��84�S�?����^�G�,��������Ni�S��Ue��z�k*��:��	EEyM�sY��x�q6"6��o���=�XD<Q1�k����w4������nj�E��b�YmZ`\�K��0�K�l.0�����G-�����˄�4���)�+�Q��������p��-�0����aQ5) ����<�ª)��h$�×�Uo�f%�eU��\/�4!k&�_S�碊� �^ Q��N�	�����;X��L�NY�!��%v����q����N��].C��y )Eb=ō/ ot߹����v{]���-BC���#�G����$��W��Iϲ�,Y(Č��޲ye��}�;�P�Kr��G�P喼�IV����7�2um��õM��M�nt�3M���j�H�7������/�^~�J�:�S�&�w�iY9�w�R��ּJ���D|�y��`,_ \���ന�s!�1ݟ��~�Pj�:_;��X�'���-�6��S��)W��II)��p������v�Rkc~L��,��߻Ó>q��͞)�(|g�/$���}h�5*�M�u�F���GZ�	���tl&Ke�d������ ֎��UoY`t����tW�l�26|�����eſ�dG��r(����wW���So[jC��L�1����>����ѹ?n^�V1\�CF�}t�]�T#�"�2�}*�R���R��vm�N� L�A�2��q��B0��U+�c(�%8�;&W�,��8������Z�G�ݒt �d>�U0�L��b[�������ڻx&�9�UMD'�
߰�ʟ� �b��F�A�Kj,(j�Q1���m6&�/��5+���,3��f��w<N�� u6���m�
��ʽ�5a4T��۳�ܱ�=����9`��Mn�X �b��^F�F�~f	��Er�>^�c��)'�d��m�;��2B����s�?(2J�J��׉�<`�>c�
^��j���D��.��n2OdGG�����M>�F@-��1U���z�y�6�s���g��{�aǌ���蚞eC"���1�2��\�ъ��ͳ��D
�ԁ�<�Z.7-s�c;�` ��q�T�pg-�,9�|��Fo*/5��,�z�wI�Pg͢��Js(�IpD�}�r��"P4�E�5���jp�_%��5�h��X�#j\��O_h��W��b����ڕ�@H�ZA5}W�\�r`F�1�!�;98��LK����i�9;�wЖ>,b�wC}E��!��t��#�d��� �6���8 ��	�z�������u����f�||'��UX�M����ڲ�͑B�� ��7�ԙ�a�~h�o�U�ZZ( Y���Gu!i���	��Q��1	�X���J����k��`4��G$�NgFǿf�9��Xy�X��v�� ��}ah���춹Nli���z;2�4��[5�,�(���c�Wt<��sȺ,�*���1���ɾX�0;�(�	��"�(yF ��i�:%�+za3�E�޷>eƎ+�b%�-\*�Wbf�,[H�w�y�1>�:���JSAxxΡ���|J�|IZ(���YL���GV�F�俫�D���\e���f�	�i�>^#D�j���V�U�����z�sD����)6Z���ܾK*�/�o�!�(�:�D��A��7��k�]8r�d�L%�%e�6��.9�J����c��r� �����Q�t ��F�d�yB�/��1̴�����x����C������J���e��I?v���{��0x�������5���a,*�9&>`^�Ƨ�Dz������'�>|l"g�l�ω;"��:��ψė�4\o!�t�J �*1d�2��;���DGIG~4��:-0M�+�P1��`�R��o ݶ�p�����S���dI/�6�t��J��������-���ħ�ė�УܗԔ�ȥ�����̜W*ooAa3`�s����K�[?q^h(�3IQF]���pԆEyz�4Jnz�kp�j��<v+�vޅ^Q�Qq�9g����מ��\�I͝[T�Jw��t�,P%��4�	j63}�臃�>��6H�^�m�G���\>��t����֋�	�?�+b5G� ��FlO�U��8��4r��>�dPLdkv��'RBn�%)Th4��»���85H���,���\��6�X�\C-����h����MWT\lǷ��3��0V���M�y�<�<��AQ¾GJ��/q^�u�<f�B��Z������ݙt���s����@�B<L�I�ߚt���꫏t��4_vGn%���@�HP�d�"�T�֚աNXڬ����):��3{2�,��FT����yXQ��;'��4����<���FJ��k�*_�/�Z3�$^:z��6g�+b����G*:��s�;.�j����
�9�坏�������B�1��X[JU�,�m+Uew)B?�k�<7�2��-lЂ?�����[h�rpi���T�*pքbj]_݈��t+\�CC�-�*�,�� Rc(�s�A���ݣk-?T)�%OE�6
Tv<W��Yj��������7sכ���O�3��R�~a�5L�1_6�ʳra�KΠՉ�$�-J�V��8�}�(��Υ�JM�գ�
���KL�^��bJ�b.�<�1��Ϥު��t�Xe��<��Y%���WW�O��_�
A�� |�D�{�m�dG)i�PB��v����z��-�,�l׼�t���VӆI�C9 �ϩ����z�߼���\1P�_���q
�P����/:��sAZ�|H!�`R޲�_�mv�@:�g�;�V�M�m�r��y�tC�&�A]А5�/R{t=g��_��^�?p���)��G���J�־��� ����kB�R�^P�k��?^��Z����V��-H�G3�h"hS;�r���`c0�S��}�q���7;h��g�x��(�g�u�?;�1��l=�U|�`���Њ���b%0_�1W[��%S�AA����o�7uiS$nym;������-\��[ ��d`���!r��&�%�qE����-� ���:�Yښ�Hq�3Ը��� ��+��������3���b�h b��Z-�j�d���
�j��(��s:�:%����Q|��g�
7��:�]�~+씱8�B�C�4�4����FL��=E�}Lq��m'p�� �Rnr+�D�k�����[V�� ͸�h�3���gᇏ�e��}~JA�;��l�,T<��L�`S(CW����B�PNP{�F���1ܥ�� ��L'����wu
?�Z4�*s���^�����9�$�ܻ��T����F��'e���l�F�KIWI�o>�?A���*T�UB@>��Z���q��dC�/4���. ��!3S���kX-���ќ��/"
s����G�@��.#�~����Q_6�6�u.dhIh��;A?첕���g�RRU�K�oū�|)�!���n�P�r�b�!�p������wC3���P�9�/��x�F�-�@�cg��NwYB�rƠ��>��� ���
�rJ�5��ʿ�Ȧ��D]�5�@�	�k+�����h�z8̙ᨶ��O��s��4��&�^��V�P��%�FkPJ<��N8��ƻz�
k��r�L6t�����0��^̷)W9���!���K������'�,������ !��C>���GB�� ��OՉK}O&R�)Y��ւ��)��5���w� �x;j�?����p�R���e��\?��\?>�D�����B�KL��W$���1�}v�C�),�e.7|����K��	�L���j�X�_�>�K�C���/:\"���/����V}i%�Qu6�8bz"e��5�O�eÈW�Q�|����~�R�%�&s1���Y��L��v�M��ی��Bh��o�q�%孶/%��x~"���*�gIFʶ���|HDܮp��}��J��oH�H�ʒū�P>�
(4��}�O@��r,5���]��_�[�C�h�F-�q��>oM�HӪ+1��Xa�#��p
��nӁ=�p��=�^�4 ��Xi�b�U���7����;k$h�����c{�2n����	�]
��Y�,{6XA��56���A��iNSI5C�IM����F�M8�L�������k��T�jh���.��z#ttxۑY^��z���>����Y��xs����@�F$Q��ڕ����zL��u9�x;8���e��G¸#&�OX�꜃#E�fv��^�[H�hW��ĊP�PJ!��u���	e�tľ`|��¨�}���[����h����� /S�����z�&w�����j���v�����_�L����Iq��Wlq� 9�%�bJ���A��X�3c�]�?�0b!T�7��<���TN5�Tн_oI�����Q� �8u̀���j�`uW�RN=3�#r|�K��������<�B3]p?! Vj�'erL�^<�����+�C���D部j�g���C[s�] _�e���7'��;X��fߣߓ~�8R��n8��؜���Z�9��צb�l#��
�T��u� @֍���Gj�z-�b�~ �J&}r���?X�K�XN���;A�9��Ɨ-�	�`'~�9�Y(S����Jhm��d�@��3$��7��Ͳ^�)z?�~��d EJp3���=dʊ��Q.NQO��J
���Nm����,�]����g�"�qD\���a���B�á�&���[�||�����_�R�4d�/0��ԅl��ѾHuQ ��>������[���?�81y��;�z)�h����O�"�
�����x��3VN}�~�_����TQ�P�e��,�q�r�#7�2t]����Dn�-O{p��Y��y~6���e�~�%��e�� �q ��Rg۳��.o�Yĭ�TM,�`<�I��"i���õ����ubJ�����\������_}|Y�� �Ng}Z��V>����0��C2n��wbl�WTI:g���OT���n�rI豭)���җ;�:B��y����O��������%5]R�ClM�)��:Di�}o(��S���"=)��X�a3������m+OYp�0����g��V��a<�(*JeSO��P��!�Q���8FY����}���U�/�?���,�����&z>4���[�h���hI����H�)1�Χ��o)��@r, k�;u#�5N+1~��d���FUaM^3n��=5�!m�{�-sf4�5��߭ޟs�c��&��;��욤:��H�����,�+>����p9x6��p���.��L۰�����<A����S#f�\'f��Σ����/�PO�����&wu8��~�e�e��'߻@�"�!����3Y/3�r}Vf��H��N���n%[B��|'��VXfa�T~']����� ^��Dh*�tS>c���~��G�}T��L+��P�/��j�
�m�R�%B�Q��
Vv�D%wŢ[����]W���x�?@vn+����ֳۃ�[���
[fQ��&Yb�oSs/[2u��^��I._����_��AjĨأ�˖TCvɑ�F�	�OI�@X�)sq�:�{ �k����d5=;���E���T��f�jal>;�t ���HwP;�Vo���-D��-]�����>ٲ�"����oJq%�d˕��B���(c�����=�L��~\�1L���]1��j�M ^4��8>:I�Y��hoè���b��V�/;�6C��£���RE���r���Z�>�r��IWiS��3'������/x(z���m|�)�H,67jջ[�O��ܼN�n.#ЭO�����R��	�W%l���B0���c��m��[X(�S���V�����dT_(���ѣη������V0��Q�۝� ����{���,ܭ������Ml�O�1+H	��E�N���M����c�HYp�~�2�4Ċ+?�Rz�ezp{����u�,���M�_������]�Q��]CkF	� ��H�����`��F�����%i�0ҚH��sp�S媯w�B#+Y&L�Uƣ���������?m���*C,��?��TP�h��C�?�u�}"쉸��(6^n�h�%]�t�Q�NF]�tD�*�J�����tq|���,��`Ѵ��� �J7��(?9��w��f�Ʀd��s�b� 8��hM�xD�8�A6¯�����V�^��l3[i�zz�����7(�- W;��8^ ֶ[��fա�W��Rw��i���,���[����&?�p7��DKw��"����g}w|~w�înR$�b���SD�b��Y�G�"�Cd�����TV"s`R�KQn�Yc9�`)����1
�\,�h]��<L}��)fG������Y���V�Jh�����ٗk��)R"���:pP1_�V����Bc��2;Q���n�lC�����]Rx�c�������Ys4�s_L�J/!�n4��*�4�a�v�����􎞹> ��)��&ז��Jd������ԷЖޥ��̌c�3���t8.���X4Bu�Bj�<q7&q�[��m���4.Ąu�ڥ�V�$(�@5�A~H}Ln"��[������7g���;WU����Ef�?�p����v�^��^��X�^��63y!un��x��3\���"؜y��N�\;$�A��/�8���8b���l�f,����*{����kPTgK69�_��:�q޽&�����MWf�%t�g�GO��	vH�v |ߤ�	͵��H��ӥ\���3�K��+:�Q���k�f��#^�����{ȴx��[bL_gꚯ.lz � q��b²�2��8L+�~��-����Ok�V]�\W��A�z'ʶ	(����]�4�u1c��q���;��� MJ���U*�q�>a/��]E(/����?�uԜ�ڶ.!&?����1�����U��f�k�f#�h�� �Q���֫4���u
�/vr XA���{��,��Mm&ٟ����|��ec��ԋ��� v��BS�ן(�+�(���a����=�	t�>#�'=����ABf6yE�<��Xη�'0�W���8�p�����n�:�����ˉ1��pVϪN�����u� <p���O�4e[8��ە�*nŖt.R��`=rl�z�
� ifݮ͇s0��̼�������b�$J�8Yq��í��1MJ��o!9�������Tx�r�^H=�^�`�<�M8P�f�����W]2��($Imlj��4��DJ��	�K��NN��X�Im����hm�<��S�ȭ��B�@5�Ƿ�����Ħ��L�2I+1���+��k\�c6���ڋ2?@�p�����ˤ�}��*&cC'I:H�E�B	��gL�YF��͙lNC<<���G�i����0�@���Ī�3M�nh�CVmT~�lm�`����,�H���V�#/cR�wl�a������h�9uc�eE(��K�%{�]!���K&�xf`_������ X��%��H\���q�V
��	'P��N:t�������������U(�������u�.Mr�\�U��%�q���|����"mce�swmr�v!��_�`~�(�Z�|�űP���� �Dc�t��mn`f8�3��7{Z�lz]q�?�x4�	2��+��ն�_Pn��-:P_�5��քe -��"����+0*T���
�V�:h<7:4�>}�҈�Xu�����<��#��2��2{¼�L�x��03�;mȄ!�D��C�Ť"��j`jL*� �w�T8T�&��蹮�dr��:�P��^��_�5鐹��k
 ?�]pۉl�k���6�����G�Ao�j�2^���]��d ���^��p���	�p�-�˫�$�H���XI�󚇃�OE4�c�f7����mLɪ��)C�� ������b��k%��*����*Q�Hv���Hxv�h����˹��FDcIc�OhK�l��/Im:V0>�4�k���FZ����6�7ت�CC�Y��*@Cw®��[� ��]w^<���8�.�=��^���ѐ�z���J�3���w�9��Z\]�-Ҹ ';�� ̧�^�ʏh�IȤ���6��X��WW��+��_ *#U܈�K[���ÿ� �9�J�Ym~~S�%L�w���~#j�Ϳ��n��$h����!���Rߊ�{�݈M{+�𰅎�{K��T6��䲃�P�������ێ��)��{����L��Jܒ����A�X���Ww�;��cP; �Y3(_���o���h�'�%=.�ԝYߎ<��rR$b)�'�֩��N��3��Z�<W2dB��E�Q� �x-�:�L��^���
�� UF=�>���ZF�,������F1倏��<�o�s��m�5 ƒ�dwZ���%I��W|��v��5'|\�����^���@���ָA�v	_i�M%���)L(7^$��9��7����?�&��>ľ4q�r�9������I)��ߡ�J�������nZ1u�C���z��u|��uu�q)��رԟ2�LR���r=�"�XÕ�2Cr�wp0ŝ~E����8ʒ|�W�VV�i@<��R���SBf��lo�지���,P��nՕ=�]f�9�n�$A�b�+�x{q�.�N����M���	�����U���Ua�s�Q^=�!����o���;̿�Rk26�N��.=��q.At����͓�V�eIf�S��ChuPЫ
�Pf5ê�R���S�T>L��EX*-t+6-|�f�|UK���IO�-��(E��%2��I3��Um�y�~�9V}��i��c����Z$�H�	�ah1-�å�����u�e���L��k��.�l$n��2��m��1*�GA%S��,L����N�5���w
�EIPa����
�%�0�ME�}+��b�d4���x�`�iEx�1P�ı}\k��P���=p�Vԭ�S���O�\�Lק-V=��ʶ�ʃ)��N�����%_N�?�%�0�w��Z�$`��RRm�� ���9���4��SA�����lo6'�K�E�(�_[�^�$����G�ɳ�_[�E�F܍��ۮha��_o���K>��W/+K�&�M���R��+�h\��#iG���W�|O`o>b�`�:�y�Bm�7v;GTFN�`���o�|U���A�^S�RMx�Z�]A���b!�����D"�u!�d ӶG��(jk��5� K��s�t%;f&���r�r�X���S%�冮�I�����3,�u���Dkv�}.}��
� Y���)�� �k��L�F����@*����52������tJ��W�u�����7LI�#�1_�'��:�JSz��|{x�q�m���_S�:-'&Z�>�^��/��CQ���l���T.��(�������}�S��J�`C�ط�I���*�hD��q��H�iڍ���TlIJ��e,���X�*0��?�H!W���L��MP��%̷�K0(``��$�:*��J���N�����胀R��F
��kq�L�6� �ߪ��N�W�Xη�d�F	z����p"��7E�m���[�S�7_U��L&�亡R�j�{-*)�cz��ZF�Nu�An�/?��2�JŨ���҃qwt+Y�*� ��e�7I]���5�j�����*�@7���)�ڵ�����~�א~9q�*�������1�ܑ`�"977"��y���J?=Ħ��E�ڪ�e׎�0ݙ?�eݍuۦ��f8��JQu\��9���5����f�ŷ� e�,��a[�X��Z<X}t�׮���F�p����g���t�'Dmb����'��%��9�a��4 �X
0��8��b��8��D��MT���+z���5���Zx��k��i�;|��A�qt�W�F~3��r��,��D9'�d�eC�&x[��1m�7f�y�#B��k� .�;و��͘����&�
Z��Mճ�o+B�|���%��k��W� ��r�9��N�$z͕գ�JϞKi���է��F�mP6cs�?!P@�h2h�U�q<=7�-�'�G�wyd��:��B����_�Iw���C;=ti.2_}�;���.�Ք�)*+���!08;i��Z���rTL���Hӱ5�A�[�$!P�q^k�܎�o��s��q�F>�&2�Sy�]A���n�q�X��'�v�4�l�ggL��m�оw�|>����04B���T����ڕ��E�C��0$�^���3MpV�_�:��@оss��2Z\:4C3hF{IQ�wo��.Z��z�7k�8<��Lm��;b�]���lnr��sNyQ���)"ϫ}wٺ�(i����f.l�&�q��ҏǂ��j� p�tl<�9�M�����/ �I��U�E�|�t������Y�2��
"��F��X�I,�/���ǋv���%e�ϗϷ>�s=��~sؕᮮ ����z;!'��	����9ڬ��ۿ>���us=�O�'~�,����'|��f���_��eYӗ`L�(t�>�����cc9��>x�K�����Y�ZK{�|� �iX�թhSND�7�ѹWQw�w�橾��?����E�b��n�hOu$�� �C�I�	Dh���礌����,��5ON:�f��}�G]&^.$���mZ!���z��A�6�
�&P�-l����\E�����԰�T婸m�F��o�$�Z�	`�������1d�;��p	V�vw#Q��T��yZ:8Q�%�Z�g�MϛVZ�F[��s,�����b$p��]H�F���HE�g�u�Hx��hϣ����)��6�ʁ��f7_ZS<9��P�zƽ���+3Omă��QT�Ắ�xT��p�[C�}}1&�g���&Uy��:�sN��x�|ħ̑DNݦE��{���|��ȶY���a�\Rd��}�
�叞15r�1�����I�����Y������{��,�귚O��$���h� ~�m�U2 T���-0Wt|��.�&���I_	���f���+����)�6e�3Xw��@I�G8�$3�GX?��sֲm�MK; ��_m�@�a�#j�$�(g�ǻ��RB�P4p��?�^BCi��T�3�`q_[��8O�����@H��}z:�fl�b�;�����ʄ
 ��y���:$	���R�W�#�-G�ݕ��^���ggt����/�V��~��h��+�i��cև{�tN��Z�w{P籯���&Q`쳚֕�h?8�����~�1!�C�`途k��i�փ�@�Ub#Ғ鶫���L�Gh�B�s@ߩw_�ÉG�y�s`��D����V���X���	\'"U�����a�>�Z���ŵ�d�_�0�7Ql��2!���6>(�g9�u��0���,��%����6 ��^p�1KI�"#\gig�tސe�3���5���8mY�5<#)��N��	E�wl$��^��9~��+�nN�B2����6=G�논Q����?NF�H�?�#��NJ�Y)��炋�U`;N��9�R�ZN�ld^�[-~a(=y��1V��J!P�:�������7Vӗ��:�k�%�!_ٓ�B\�9:�³�+��s����MԪ[l���	-q�j��E�ϵ��^ln烃P�G729j$ח�`��^#���f_�M��w�H��1���e6=}���4!Pm���5���W3�UeRxN���pn���j!�Ԋ󣍉���"��ߨrY�(GFƕ�h}�ēf̉����& lg���L`>��K���<�I�����hP�&�>��r���Hn��W
_�#zmD��(�����_��5ݥ����r�kV]Ӫ����%t�0�[���B��K���X�`����oIw#`~��P�y���iw�)�+Y�QUeё�p�(G$՝�BQ<�B�;֙��%�#�8.7Yu���;;������.�M�K%��O��i��5�/�cE�+�V��+�7|i�#	>��gݯ	�H���TZviU�߰���(}r�/N�J.��B'��«��y���L�K�a5��-����{�j�2eQi���/XIS�w�f3K��fI2MrsQ���Tf�X����#�FU����Xs�u��L�֋�_�RY�Cp���LJ&��M��;)\�� �)��]�>Ҋobl]�Ҫ��E��~�P&��G��#�}����S-��NJ��@�"'Nh��2��˝$�x�x���D�3�>�������pk����h<����p(��;`No�q{Z���ڳ:f�
�<�'	B+����F#����d�bo[ɀ���B���#�:��^�#�X���5���*���D���ݾ63�~x'��~ͣR=�0�X����cjJ�5ύ�,9����j�&�5A B=Ɍ1�86������Aw��y�T ^�-�eH-���1�:�(8ݵ�8�����Hd|p�kζ��a�J���:=W�
��,70��e�8��a� ��,Չ\�`kL��n�巶��_|E�|��q�m�	U��s�/�Tb�'��g�e�����e
S�r+��T:[��\�D*��v�!��%˭�&�TG��F�.s������`�	x������]Ŏ���,;,��$�L�^Y���ܻU��g&�e�.��/E�j�����z��ͺoO�֡���!N��+J\�*0�j�!;Q��՝�+��H��/p`ۣ�#ZW;o�7!U�-W�뽡�����|��3lAl�D�������5);7�AQIÍ �w\���(O�M�F=�q��=���rQ�y n&�NS�G�;x`Ju����݇$d��o�=vyL�]Uzg�j�]�1�j�45�*M3�0�Bt\�JUN��I�Z.n�I���$L�������$�8SMBž�)�4�0!�Pԯ/iB{З$S/�	�˯ �_��V���VL-I��o!Ô�[�|q����9�oa��Lmq~�/^�����I��*�G���bu�g0���m��)>>P���A�ժ�˘�k�D4�LkUn��ɰ$-��6�g�/L�̧&�9��8U�[��ޘ�q�B^v�R6��W�������-���L�+�Gs�\/��P�ͥ�_p�*��*�F�I�
�AC.����+�\hD�Q-�֍��<g��k���@��fJ�a���5-a�2)�����>(�S6V��&bM*�{q)#�D3�����}�j�I�7���u˿i

KV�ȝ$tw����m2��^'�_H�E1�XRs�ݷ�f�,����}��uL~��͚����0���f7�|��?^.��B�R񳴕м<]%�f��Z�2�l�0&^���Dś�竷����{�(� ˊ��#�[�@5���Cl��y�:�(\n�=uv�(���g�U�f����U���NQ��7D�'����Ў]Q����D7�z� �W��G�#8�-߱���<Ͽ��\eGz���f�*�����@he��^p$t�5�Xc}M 9���q2V�c����D�j��0����E��'b�t2n�gx��%�T�!��D^����v��թ�'E��U]ʣ�>/A����!5>!�`�%$�qV��[g��dn��V<5PK-��b�I�%3�����F�f�`��ك�l�E�&;j����i{E����i��5m9��Ud�����\�i��!X$�=����gv|-45�P�Q@>uY�
x\*�զ\DE\|���Y)���#�@�yƎA�j���B�� o������,F�����[��h$�g�4pmk��k	����-u�=8x2����?�w��C��59|I4�\p�c埚0�*|>�-O.	�E{+˙g�S�1�(� f�C��:^�����
'Yp�h��0��UY�
���.�4;yh`H�0Eߤ���kSJ����$'�{�z�0��%�B���������4��\REsJ�q��E���z�ŧxQL�r
�{	���ZN_~�a,ݦ�)�5@&s����"�s�7ڭ,����j�d��RY���D�������w9g�ٳKVE�Z<���sPK˱��B��J�1f�)x���\�*�"~B�����|�W�v�`j`���:�9�EC����|}W�l�=Y>I�����CL�P��>١d͟>�h�a�»8Y��ӹ��ļԙ�.�K�o���O�����ǃ���[1��Z��<�;��&��pjZ��C����p��Z]��ҡhX=�ۇtbL�����gN��4���}�FwR��Ϥ���8���$���|Sz��ԓ>f|�'�L��ޡ�C��u��F�I%!n��v���1e��RV}����$��[Tl��̭��j�H��X��f_�-���x8�Ժ��&<��'&�\�ᰎ�ʆ��4��c����k���zi��nu7J���9�&��}���ϐ#د����R�n2�ob�D��G\,V����/�cxG�x![ed�M��`Y�����k���m
�Sh���QԦ�o�1��K?w{
��&.�kO���[��rnW1f�l͸�K"o�5����t�2�r��"�|/��06�#��~��W����sq�����/�?%�,@�µ����B�zƭD�����d�h͉@��l1���א�*~���vw��S#ሌN[}�^z�_p���gH�M����4ws�KmC'����h����Jv��}b㇤,o���W�Ҟv%C����S����N����Zr��0�����^�]|ǲoc�R�ni��]ˉLbwG=�j�ާ���v���ߕ��� �)���:%@��;�5<3�^ҎU�,p���m�i@��gɧQ�B�H|	���Gӣ��������1�ѻ��܈=EH�°!)�
$�*.Ъi�$�P7�(��k�X�7��e��1U��E_�] �� �l����%�̘-ь'Y��USY�lD-������6ᰰ���BMƁ�[g(}�O|�3�U�#�)ڗ<u�՛����3 �(r��܅Q�5�~����7#�,��6?;2#��g"#1�t�<�,�S#eq��G
�j��&Y���� �C�{���� 4e�-ۈgr��M7�\Z�L�["���g�K��Z�v\^ޏuS���[îO���0q�z�k4b#�O�#�a�x�]T�m����ħ-�Wk��m׆�!�P��DT�SyI�V�zCi5Y�$�h�8�X�0Ŝl�7��VZQ�'���Q�i��Nx^!n7x��B��4�����u�����3ۃ�a��_T!��z��(��!:�91�*"jq�/� � kӪ���ŴkNh�9��t֣�QM���$wj�@ ��(��#���{$$o�|�_�,��(_���0o:u!��6z���k�q�c�]��g��c�b'�k����hџX��Q��[VX�� 7��\?d6�O���J2}LtP���������<[�����O̜��I5[�\4IV`9�9��r֗}Z�����/ �XO,_sC@�W�I����@_7Z��S���'�L���wZX�J�r�<�Q��x5fe)�k�7Ow1~̬��W��:�P:�R����{Zय����q��݀�0a�]<D��K���i�v��50�@l�00�ilKt���	jb�)�lh���=w�{� �!�-3��vZ9�,����o˝@��=yw%�k� 
�1s�Z���~���c��Wu5�n~\���A�Ǜ�ׁE��O�� %�55cXMk�B�_�v�!��&:3/��+,J��L�C^#f�@�h�E�q��(�m�+���K[�U�P���X��<���q#5�&�b[c>Z��z/�c��n7&� j��F��C3{�^��g<Wq��I�Z�����U���YKXր��<Z���.��>�:KH��x�x�����?J���=�)�8Q���c�w!��ca��kڞ�;0��R7wb��߷�zC���*���G��8�g��y<�DќM�Y�Dܺ�_>Js��S���E�K��ՙ���o�ՠe?S���������jթ��Y���9i������LEp"*�7n!�3Ò=ܐM��[T,�3��������#�=[�x��Y1�n��!� �sd�ۘ��k:��U�*�T����NDZ3���;C}�#�7��,�Ӊ:�S�v�_�j
$з�9�D�\��vYhE��
u�$XKUnC�X�x�ם�����+ �m���F���*�Γ�s��RXb�M�������l��w�!G)A������|j�����A��4BP�؂��vk��J/Ua�X�/�|�!�� �9��7�����r�J���?�0��5 q��E�{��F���S�Ic��|V�����9�
����a3_�ve�Af�nu�����@�h�#��3�>-L(h��:ۯ%O��]QH�*��V���w{WI�"7�d�c9;�p!�t�\�k�u"�Q�0�g��ӧn�]�/�2��&A&��91[�[z8	(^FGO����]�1WL+<2���Hy"�Qǖo�i�6�h{�m��G���2
�ܭ�7Hwp]�z�)��\�����z2���������v��ĝ����X���Ub�n&��SMֺ�Gn���G�T�c�E��|���:?@�A�WS���q(��b��/ְ2�׭�  ~�C��1�|lt����' ^��E!+A�
u
�P����%� �!�4j�PLы�#�| M�H���)�C�� 9{�uKҀ�^�8��f�����U~c�'���J�����d~Ц�vUY��tQi��~#ؘ��Mb��e_��-�����z.����?k`�ӫ3� �୥����q	�L�;�^d�
��X�W��r��ձ�)�y��Aܯ��Sfi��]��;G9S�#I	O�
vȨwf�����1�|m����&ġ���r��v�������"�C�F�6���^=V-&<��Cr��,>`7ZF��k��V��� 
<.G��mA��#ؑ�K-��.�����z��Z�k@\�3�n�,n���Wc)�d&v����̉y���#",����#s�v(P��O��#q��/�QD��m+�x29�s�ٙ�ܻ>D��#��QhE=�_�t�H����\ΰ����x�b��xA�*��t�m"��^��F��v��أ��e&�M-*����H�8��������|qG���mF�^�'��wd[���֧�4�r�"�9�o�[!g��k�_�GP�Jm�gc@X���E���j>���a~��C�
T�ɧN�?M�̮:a$�b�B����8	�� �Q��_nC�7_b,\�ݬ�ި���%Oi�̮;�_k a_T��L|�ɇ'iB��2��d-�%�(]�;ڝ��تʾ�y$�)�+�#W_�5����'������d -iЖ: �{z�}� S�-���0#�1�Gq�l��0h�v���j��8��)j��}L����u�Fq	������C�c�����N,<u�C#�� *�3;��p����.�:	TTF�<�^�st*{`8=e^��=�L��^����ñ���'�h$��͏1|�����IEl����:t%��W��BiN����XW�{1�?Z�IJX�R������{Fm���225zf;�+�#�| ���|3dq���R�_)Cgk7�/���c��`�\*T@5Fr=R�D�x��h�/e<�e&1�P�.q\v�A�j�Ĩ�)\Tƍ��[�%%�<c�j1%j�>�0+����.��@h�W&P��V�h�H�4lN�1�#�E)/��ߘ)�SC�W�)���E%�"�8R{��1����.�-���V�tE������MX�]��/q�*�6?m5��84��D�Y ("Q��nEa}��)!�T,:ޣa%�'��W��b��V�)6K���Q�f��qE?�cu�m���6;n�����CK�����ie�wW�>C���U��,x`�_7���y'�{i�:�O�hf�+Y�� �s6Px'�>}�DؐV��J�w_u�Hw�=Jj�K��@.l"�[�_wr�25��nQ>;E��|�`$�my׽b�ɣx��6����z���z�y���j�|o��
&
'.�ALd,�� t[ d��(رqS�R��"7��-��:��٥���;��~P�[hqIh��z�:j����h�7�՜�jV�B�5~{��I�W����$U޻b�%Y
�G��hc�,��߱|t�K���񄩝r/W$���4���w��_��>��Sܕ�Tϗt�U��E=q�d(y�VrJ�J>��-�� �7������CiΊ�?ڒۯ�:�ZiUQPek��3c�k��v���6 ��@���\���a%g�>�r�w
����k��$gF	Bo\��4�;|$�Kc��nw����]w��������\D6��r)S ^p�
�>�8�;m�T�Y�6�y�2�A��O�^;�jV_��J�~�����C�U^̿���,�+��^�VG��_�?q(.�<͹_���P���tG]'6
�_�>����1`�5�i�y�	�ӗF6���hE�GJ�k���g����^p���bR�kt����so�-�Ja�������끝1&!�pp�d2/���[�Ⳟ��r ��[�.Or*�h���oy`!N�-�����쪆����%}n�d`�r�o!�b̷�^Q���ghњ8�;�ES�nl%ښ	�rTi�@)��yZ����1^��P!�^OZh3�|| ��`9���ǎ�_�`�@p��m����-�}���0�ւ.3�	�0��=�Yb��q,;';@e��*�ul�5�.��R��� nFڻ
�������Ӗ�ӱ�+b7<��ѳ�0ǆ���38�N��%Ӽb:�B3L�O��3�+�����>t�RX|��muY6�m�(j�#�l��5(�7n�Fe����t��dg�l�3� ^,[�_3~.���~o9!<&�L�iDC����Us�Y_�����C��r��`K�Ě��|R�gn�ru!'=*��D�E�3��?�k;Z�Z7\Xu	ž-`j`�[o���$�ym�A>��O٫�Y	�s��g�,t&{j������أ�v5G5qWKsZ�Ա�L����蚊҃}�J��ȭܓ���5QM�ȢG�P&��a�ja�W�Ն��+w��w��)���Q܆�f}��xRvN�L�l�m�mMHx���R�2Լ�{0K�8�����]�6N.�K
�V�c��=$�/E��~&<4E)�A�7~�t�mw��29y���z@+��yRA��eW(�-f���&Z��V���s�G7��G��
x���J�X�>�TN��Yd:j�ƙ")c�Эn�(�E)�;v�\�����3�6��P_H4��qm��&ߤ��.�ƾ�H`@t��>|_<�'������j�����wӪ�yS��m}�L$���	b��'�1�{T��\���'��H*�}m��O�|�X��&�0&����1�p�)����U�H�r��_m9�9r��Q[��x�|g#�-�a��˗|��E�~=�/�9<�z�|�Ib��f�^5�3ݓY�_,�W�Q�U��6��Ǒ_v_��?�9�r@�x�&�1�5���K�"*f�r������E���%;:|�~F�0�����LТ��a�i�6�}���XJ�ht.	j���V�ӧ^)<��O�3($W=�jK����49}|-K�6v4�&7h�����\gc��Bp�����:'is�!�P�!s��E�����JF�Yp\��:��Q}i�˧�4�&�u��0'ofD�f��=��Z�kc8zt:�ώ�:��7����]�U�̏�:ۻ���^o�3"�p���2�B�l��@E�����>�G��������[��x]����ċ[0fQv`M3}�u]��WGh��8�i��Y�	����kՉ���d}+0���G<H>�Y彧�YԦ|��3�*�}�,$o�� ������0n��%8]/�\�)=`���3 {_���=�xF(�f��uz۹ߣy��8U����#crU���N�7ԟ�|3�L^��*�--�"�5�I6:�g~��NZ
�q1��������G���!%e�~=~ko8[��5e�3��Х�۟a�,�[d��9��Ɩ按A!��$v�����b�</�X։�c�<6xl`�����џ�}SP���ڳ�J9���m 1��桐�����+hwu*��~w�j��@ÃIౌ��2����$?j��b��<���-�ʝ_:顥@�?1��8��G7M~3��f�fWz��Ĭ�A�2�����-��{��ַjq�}���)�Y3Ru �c{�*�o�*�+P�0�,�v��~C-�N2�8$p�d������@V˪��v�/R7�d�D�#lU����;��iRh`Ě�ghEu�����_�F����DEX�M!��^[~��%f�0����p�)�tZ����f*��z�:~[�#9g����cBP���HVt��`�h-qZ�8�!�����B�-�1d���(.���̖�΀��U���7��(�~����2f�U�Ϋ6		~���Q{�X�("mI���>�0OvW�i���]4#��R؊�0��9�(jtm�J^�7ജ���)��+9^�P���杧�r�˨�ز�����0<P�-%�rj�'�.���ҿ��̦tWINZl��p�\Lx,�o�+썷�-�W����S��Lp|���K��y�Y�����y��6x="��aӰ���C���`7RTmH����=��ԫ��炵	��>����,a��[��?C���
4��Ӂ���<7@
q8�nȧ@;�T.�����ֿהH��YK�Ӡn~5^c��Ivq�VX�i�k�����j��D���	��r��I�M
�Z��#!g��r��$��na\~����'�J.#+���u�h�@fR=4ig���
�����AE�^�c�a'ʐ_�Y�̰���Lձ��ܷ�p��A��H����W=��LM��ȿ��R�.�Gn�qy"D"C t �L5��/$���˩�q��XDŹG�B�ƀ�<�ѽ�.@���)K��Sd4iвҹ�I�ɖ�&�}���Հ<~�?Ef��y
�j���ѴrW�o�,�_K�K۾ev.O#�;�M�O%XY��D�\�ٳ1�Ԅ2�dC��,�ܮ׍����0�8�ѵa�B��j�������ʨ-�.��/2ϣ��l%�]���W����pB������Zc��� d�>��
!��,G�ŕG%�w!1�x��p��^<���9�>O���\Q��hb��/�<n�vT��);_3��ph����S�aoI�)�m/�8��-V�K^>l�Iטم����>nN���8�;%�!2)���.��<T���ݕ?���dW�f(�g��I�����h�م�����Ѻu�&��Kg�8�x�`�5�T(Q^,���䀣�'q&
~j'�̰�ϯ ͏�G[�.�d������x�6ӕF�����g�&Y�8`�����Bou�
��Sd~�+I��Dc���#�Q9�n������ʼ�������ޘ���<V�y��i�2�Gy���:�c&�q��"8.Yr����શ*�(����bՇ��)������h6���lN�������%+ 鷾��~-wl�xd0xW��� �B[s��\��d6��h���|Vb���-Q�s������>�����Ղ3�^����\�?lzt^�,�8/}fJ�"/�a�nM9�@�r���T��q��=��k{*nYO�ݕ������ǿ�?{�l��"daϺP��>z	��)-S���< ����-�eB�n�Fk�G�lJk$�K��u4_o���c�i�9��,�e�ѯ�Ib������I2��W���
����K���X��4��M�wM͗Sߦ�����K��.�O���8���κ�_x�0dG��Ɍ��`���8��ر�"����dH��g��بWڌ,Y�]�S.>�4K��AT�jA�W�5��',Vh�����Zʛ�����:�@r�V_�.�v��ܾ�6z֓�f�5��`6���M&����m�$RB�q�ko�=?TYO���=����!��z�~mWs�|�O��{2� G��������]�pV
$q���
;��v�9ެh��Kp<X�v��cr�1Y�N�\�Cs�0pǦ���D'r�TQ�B^�������<q�C�W�U	.����:S��a��wi��<l|���ZU,������B����f�x�9s3�Q�$�*P����
ӊ�E�Z�3_i/��w�)��v�}���ƳF彀(����3��
����%��s��u2HW��$�ٰ|+�`�'�=W��uM#�t�
���l�x%�w�t�
f�L�C+]Ò)�P����L��ݻ]	.&	�z��s�T�Ol#�����z��Qԡ�m�8h(b2W��D��I�&6����<����$�=��6�o��e�Lǲ ����3�7J���F�h�g45"7�C��-������N`� ��8`y,���򆘃5�pŰ,��w�4P,�s�x�zIL��l�R�:C{�Ē��	u�Ĩjj�-?��K�$Q��+y(�R���mȲ-��)�� YYBJ�����h�z �,��&�ʑ�����`��u��V���p��G�?��G~H���ϰR�6�fP&�|��_���|f�>nN�nrc}T�ڙ��+T��'m����Q�݆˂��#���zghU��@�Bt�s�$-��L�>�q�n���8�,@���}!C�d[d�[�}��vFM cT\(]EjYhQA��s�K4/���@�ғ����x��3��=�����s�}iK�C�~b(ȧ+y��y����{ވ����`׉��bm��f(�-��uss��Z��b���"�9?��:dF��*Y�
B�Z��|eTb�� �8F�9��A�7R��C �Ju��oR�!��<�3���
8�HE������Τ�j���Ě��*4	���܊�ǽ8�S1aی�/-M�&�Sz)�����|i֯��cind�6gÜ�vg�Ќ �S�Վ*��$��c:iR�1T���؝�U��Ғra1`I�B�{}jK���)��k�j�@8�zZ��M�M�]BmC�3PR���\�l]�B�=��.��eĆ��]�d�Ì`�^�93b�f��7�ؕQS}nЋ�\K��
�-v��6`KS͍��eH2��L֮���)���vk������1�J�aae����apFC�o�z��-�BǼj>�lV�smϤ�2G�E���xeb�o�9K�͉�k�E�����ӂ��b}�����r���%���Ώ>#8�vd$b�����l�Ay�Yj' ��������l 0�i�n�����w��Kb<t��{y=�������#��KeK>�V&54��X���U�
3^��Ç ".��Ps���^HU����VA"3�#6�ķX�)(��vO��Wy�U�p��u��BݦGw�/���N�3c��J���:��ݠ,c��4C��0��:��Xk��/���v[hoK�R �����-K�x�D���[�P������=׮����w �e�}y�P�=���+\���D%VAm�CC"�ͺC��g'�q���!+b)4v�@���ꯂ«���4
����0�+����fu���z� Ə�̪��Ens��Qw_)�	���eMg��Ƴ�s�C篺��td�!���
�Ή�>��_�4��dd)W�pT���5b�f2�H�'���usȼ�!̇m���T,�갗����}�f�',$�tP���1�{������T]�$��'�#�g���&��V��ΰ���L���m�Q�}yeS��3�?�6:�x�;��a�U�W WÑ���juB����6f�~�ruTOfL�h������!'9p���M����� �co�M":�0S��p�6D����1XE��O�A�QIE$��ia�ڐ�4d�;d������z���i��(h�T�x|����G��D�����##�':0*��ɯ�12Gx4�H!�Pը
yL����I;��!8�c)�pB�9[�������	2��N���c��������!�;G��V�N%7Sq&�k5�.A�� �'8�a9�u�����*�X�%Ĭ�1������˟�j�n9!�/ğ|�\��N�����u=+���k��1+�Vw䶈$`2u_� N�E����Y��d|��B����;;\Ӽ:nr�ˍI�0��$n��(2:��Z<���@^���CƐc�ʴS��YZ��:q3���˸�����_�Ԇ&p5�%��iA���_�][R��:f-��'<;<p����8w:�[�/{bw�9����� ��j�A+)��+�U4{���,	�ډ�#���G�?���l�h��@��M��!Nkh�q�˟�0��^�	�U�����j�O�է�#��̲��]�?S#���t���<�����3:�WEv���+��(6�����9�1޶6\>�.����ܜ�> B���OȮ��i�����5���y��7���Jl�*�ʓ�#��Hn�����K��E������@�F���0� r7���ڗ�N���Q�zA��APg}���P1F�
x�����¯����)E	�p����Bn��~vj�a���`qY�0B�\�G�D"C(K���m<Ш�V}��t�����W��ו����^��9�"�涸t��z���?-`�}6����"����;)g8�Y��3~�W��`�F���}�d4S@�1���,�~tbs�qC=$$}��� �L�j�g[S����-��yey.ݒ��C��}JT/*+���|7��R�~B^�>���V�`:<Z��܏�b�!��|�NXܕ���s�<ͯ!���0I/��n{*"x��޽Mq��$�l�Î�<U�ZX9s���!�������� bt�X���̖�����a� �yJ�>np�@ �bx;�eh|�K��LD7�����[&.RԅE�~o�	/��^�9M�9yDTɥ����fz�|�L
l��re��������9�;��ԍ����J����W���5ҏ��e6�+�
5m!7�HY�k��򕛧��7Fg��~C�#m��' u��\�/�U�e��M��d���eZ6�8�eq��a�"�K�Ƶ�6��[&f�6�~��eFie���A�������u$�d=A����2vQ���zN�v�#/�A�F{��4 �{(Ga<p���֡ֆ�2I��&3�����-R]�LY�RTa��Y�+d��U�s��q���Y����h!R���f���m��=/���
�����T���+��=To��D r����ɣ��|9����v�����W{�H[B�������?����6��j�i1��i�Yno��j�$�r]v�Wʓ�!m��K_�,��iQz �^��~�Uo~����v�����2�m�����!׸���y�}��+��'zP��X�/��3?�o�|�yUe��rY�[O��$��4�FB[8����SA�׻3�Mr3��K��i	��͋����;}t�y(X�k$�|Mf��ꄹ��L%�p
0"xq��=Z5�;���sp@����X��
�48�Pp�f�/ӌJ�²'��DVV܊�y\7w�f�s$Ϩ�8�b0�'��+�q��&��w��6�g>���Eh[7����%���
Ϲc��D��*z,'G���kU��^����}ZE+ѥH�孧>[���lOYs��_Rͣ��`���Q
�9�h>��}���h���o�[���|Dwfs�f_�N4�Gxfj��8��Ϳ��H�Zqzj���b�gHU:�	{�IDS[�s�r�y�+��:^�|^s��1�����YQ*�ВUV���Bl���4�������o�.�k���sT�UGOU�ͼ��H�Ӛ��	�/+X���YB�Z�1�ʖ��������h��n{��)�0��j5�G�����c����/������N|�Jcu����2D�DK��9�wӉ�ocm	�U&II[y�< �	����x9K��v�����:��W����Ҙ�"�� ��~ɒ��{ܫfB�)G�5Ua�~ʾ�9�Y�M%e?=k���X&�Xe.���BZ<�(S���xm��\��������1c#�ny�Xt�	ع2-�vT�k��VZ5�̀�o�V��N�w.ğ,��Z��p��;�=r��Z���]7E伍j���)�^���G> Eђѭ�FF�G_�\�B��${��踕�)l�|�H�O�WP��W����%�lJGo���߁�+=q6�%-��}{�^a7\�ļI���ب'y�ѵ����wY���Ҙ��f�?��U���N��s�gHH�ʁ��ż�_3�Օ��C�C᠃MAq��fm�3*J���o#�4ۨ�RU�J	���)<���<�0��'�-��w`2u\�흫�T�ݴ��+5e|j�S@�/҆+�F��~�T�����x����V�G�X���<������u�������WG�{�1�2�NA�|'��Lԥ䀴3�����"�a�L���g���#�L}�WG��$�]���f�J�! $��m��p-0�p\�t���+��Snpѻ�v_�/��ẅ�i��E��|�V�k-�Йx�47:N$�2Lx�%Ǉ58���I.dYZq'U��ѡM�U��?�jʫY��(�3
,����Yr��\D���όN�v`w�ꫛzȢ���&��3��SrJ:��迅T��:y�6M���XR�����4�:X��6��>�_�y�{�Jyi�yh%�B�E�[������MӒ�]z�� 1���j�j�̩xx��.կ*���0j�$��D��{;�%~�Q��0�u=����؟�����hLx�ʒhg�ǽ[��;k��sA���Ek�~�"�z�����x��Uz���?m���G6�����ŋ������Ľ�֬�H9���I��M����d[����� b���Z����|��e����������?�<>*��?�o�B�!�_�#��@����fMꋻ	���_��D� v�'��1ﯛ���&�E���W�:�rx\7��۱c�c���LDԞS!hsyP�	�����X[d�h M�8��T�|\;�y��9�����o��L��*۔�o��4��zr�kD��Ǔ�R8���f����h���b�]�D�K�34=,��Js�{��5�`����F>tɷܐX�,0IDN��Q)^�Y�wi�����GX�;���l��'���O����
Cw�ݵ*�-�biJ㮟�4���^b�@
�8svV�x���Q���o:��:&��OBŵ{V� +M�n�>�M��_�tb)s�=��һS3�Q��4΢�Kt��k]�,�Ro�R�?t�N��=��Sw�t�)�TԂ�/Έo: Zon`��m��%z�3��X��+/����iϗ�ePNo^�KPC�!�����!�];�k�M�Q��d�������J��#ʚDv憎���mw������W�
�~�Y���rϺj����ufV�chr��F�"����4���#7Ҳ�!��o���P���j�9�G[o��j��A��ȬJ�N#����Ŧi%�>1����ƒ j26�,.��}my��@a��m�}�^ɫ��WZ�֯�F�j����1W��(��\Ois�r���]vr�,�A,~��z���-�! �nn�Qu���3� 3mKF`�;� xpU�ñ��ȗn%J�|@��瞒y+�7[��ĉ������g���ʹ�.+z���ұ�[��)S(ʑ�}ثΧ,TZ\�{��|X!7�5Z" 0Q��")���#�c��j�+�vz�&���勳P��"�������������f�Æ!+g�֟3��9c!��ܰ����sT��F"��H�2�p�	�1L�R��?�l�����-�\K�_�0�npz:���J���G�+u ��	1�%�Z��eŪ7�=(�5�Q�Q9��҈��֩WZ�ch)-��YBU���!_�W����hPk�m�Iz���<������H���ZAS��g?�Ws6����~9�O��#��	����"��L
#�k,d�˲���cR�5��y�����5��V�P�*(�2q2U�#C�1�A&s""���k0aM�J��-�+n�Z�懤C��܃�D(=���2�-
�I;ͪ,�^�bg)�T���0�:n�x-,�0P�����s3� ��gԀb��
�B��C����0�H�j5�L���/���ѧ�)̣�s߱�gl�5\�R���i~K�R�4�Jgd1GtM�U��L��3���Y�kմy��@�(�W@#��^��HHnDZ�u��'��DvI�V���7���z��|h�p��)]�Om��ݦa�� ���,W�� ����x��a\N6�B?��HB.��"��`�8����=�{+�
��� ?n�42�\��s'�SkÂE)oD��:wf��2�>�H�mY�c�yE.��^~��a���\��SF�C8P��,_ h�:�}�e7���%��'u�dUo���x�`��ԟ\�pTHdX�Oo�|w�y�0b��qп8�s�O�M\R���m�����Z�W �.D��?Gz��� 	�(�^�q�5(�W|��ʣ�u�ל����Ǯ)�v��b�S`.�t��|�����~R�+�[FL�����$<�jxI���蝘�mNR'��� ��Ɔ��X�odf��xӵ�_�6/�n)_���`�
[�hVLĸ�kR�����缹�F�ŉcJK;���(��wڼt���Ñ�)4������o�*���/�A��Xo��,UC�Kn x2�>B�/4�=�q��F��w���=#����� ��jR��$��V�����J�?ن�x��Kj��\	��ٖW���EN�q�-���$>�L�7>��Z��>�Q��3BN/�,I��R�'�'dқd�D ��ZnF��	��\aY0=,�ґ��?�:�����d�	��%���u쓇@��mc�Qe3@�0��~yW�u�'I�z���l���n n!ƻl�೚��6���]׷Q���s$,7a���Ch>_����v#���O|��$�4��F�K��_���5zq�,�F�����zj��	��a��|`}/�$6Dp%4�%]د�x:x�~��ꉁ֫��xHW+Ҥ	͊�������;���R$|�p���r��S��a�0Ġ�M�*ݥ�c�q�IR��耄ٍ5�-!W�]ճ붼4��))�(�i�S[T׿M;/t1&�����nL�>oekmwG��%d���fv����"�R�N���M���Bď����4ܮ���cIl
���s�n�� �J��فn�U�E�0UE˟G���2����6{�X�1�=VEu�){��]D1ɧ�������U�9[��Q����/K���L2薖�XU�1N�&Gk݊OwG�nv1{:`�
e�ܴc�"� ]B �〿�%��\tͳ��[1,���w��3w �� �Ln;�����[�>$67x���j�c�?�תٿ%�����eф�.�|9����tx�)��K�'�sH��<�de	 ]]�(`����#�;qK,�,�Z��&o���R�oEr�G�+�>��wF������#�ϿS�#�B�p/���H��	 V����+y4���|�� ���*s@!U�)E�}��Se��t���H8#����3��x����*���2�@>g�Hpƒm�?��|��������u�@�&��H����/�%*/Kch{��6ʗ��������I��]F�#�N�ąfJ�KH�!Y⅗�C�w,"�KRY+#ֺUd������1�}�m����[��+�u�6�@���ǯ���Z�K�7n�y��>�$5)�0A�a߼���ɷ9[��AVE��݌�Y7$J�����IFto�%��7��ur�����:�S�4������������	5[�T���Y��N璪�x�:c$�6vu�{"��'��zù����-���h�1�B#����2��e���m�zS�t6�-��(�'�֑6��(^��:?�6�����F��g(7�"#K��c�u#o؁��ޠ�W�l+yR�lU��4�x#P���ف+w��2���|������qQ�a�c������ό�m�U+���`��B�9���Ob����gZ�y<���!P��X�G������(v2����[�SY���2%�¥�R��24��۞>�R^7ۚ��u��z>a���T6�����y���n#�ےg�������*v��;u��E�w�t+݂93��L��i������B�B�HO��������^����;jE�Bd��[��4U�k2
`�ig�ݒ��d�%N�!:�u{j�����rw��kIc��k*; ��$�2|������9�7Otp���m]��g���Ѐe]�M�2�4H�H�_[�ZV3vǰ����>����}v
2�pVB�]�n�_x���J��Z��Tq�P�����-�b���U^eRL��4���|�Kւ�V��^}8Eʃ��	�4��ґ�=W�6��y�NLXl98I��(\�f����k\��YNe}��4T*�+������L� ]�r���\��?�T�n�9������N�/s_�v��`j��$��մ����Z7D��x��[WJ���\-��ȕ%�i\�e�N�PI��_az����L�6���(�#��df	� tzщ��9�T�%M�~�ğXSro?q~�~bE�F��vK�aZ�q�][S]h�Adٱ!���;�mLZ7,0?��V��R�K�xI2E�/�n��$9�wF#ǒ/^%�}�D�(ZWn�v���AZ��FU�٬��0ZO>�_El�~�B[i$��ÑJ�z+��ө�RC� |g�2攲g �'������XF�_(��0��W�b���V�Z��f������"�$`��b~|��R)x�	�\6^I�ҟ�3��q)~�b��~�=u���O)��0\d��e�&yyKy�HLr���:�Md�Vz�w0㶻L[�RN2(���U�N�ԇlY�`��l�縩\�ٖ��Pu�Pf���]�=�� `�]���j��o�Ɓ���z.��cG��[��K��Uy��Ĩ��q5ꪬ �㏾���#~?�̷D2v2�T�1e�9�W�r��N�H��喲�f�Q�����t�M��|�(��V̲S�X<��?�/)��*�����_��A^258u�rX�`�Mm<�݋�EF<�ԝ��TL*th��GT<E�$�H
��p/���U�f�s5aƶv�襡^9WЈ��Y���N�F��	 q}�ޖٱ��ڝ�����9?�c+��m�M��lFĸ���D����&gv�hw2q��t $�7�y�}��ۋ`��w2{_%�Y�O���N]�E<�y��i����@��,����Z�}�k�S���8UF07ʖ�G�-'�u^��>�g��)"�O�3�z �~2�ʖ�5�~�usS<�N��J$<6:=0AI�|���H�; ��$�jUu�I��߃c&f�)sǒ�k�|�@��4&��*�RZ���D,(�M�	�]p�-K+8�Y��}6zț*	��Yܴ�hT+��ºVi5�5�1@S�S\�%�>���M��驄���K�-�%�F��Q*�(�������P��sӌ�7���"��	�]'��)rob���+.],�,���3�=�VY�e��b����N+z%��uԶߢ?��	M��*c��R�*I���Ȩ��6"䊎^�&�&ǥ>�z0T�)�x��D�Rݣ�f�#�����@�(�^}��a���i*(
�yA�>5�K�`����lɓ0�d4Z������10�Ug��]x��8~�a��*l�Bz� C�΄�w/�v��>?�;^��K�pr��*K��AXU�ޜ�Jd��f��Z���N�0������OE^��,_��K�x��i��_|?����+��k,���txh�Z�>��M�M���>�ƙ!
����
�U���\뇃�������t��H�w��QL��ฯ ��mŹ�(z.��Ms����h�+<椖^������Pp�`/�t@�g��ȃd#�?<Io��j�<2o�Kt�7k�6a����5b�$-y�ț'���7�6K�f�H��5]�V��!�a����ڡߝq��-B7����Q�1ru�o���;�m�6�8��Q���E�m��E��֨���6qj�a�8Lb�N�]��w��7c�d�g��m�( �d��N���^��;����3+A�Y�؄�ܗ�d�Wp��f[����F��D��g{5���l%�6�<��D���Y�JP��.u�i
�F�O�#+��<�m�n��]�'�{^r����a
}.��ѕ_9GĂ�ҿ��	|<`�����?R����h��?yK�z��{��0v�똩͗z����~�MU���g��J���Oӊ�[�q췏��Y*,gia�/�%p�ÔY��W�1��EnhW��ohޑM�5�%���q\�&9Ro���Y��(�1ˁ�M�a��ߡ|¨�iXڽy��R���:�I���4����������[����������>��j�f,�O|���81N.�I��@���Gx�����!e��*�ަE�W \K����YE�MRs�1��ڥC~��G����ՀIF�g���; ����-6{���}��K8c���FS6�2yA�,;���M���k�RUBB`.L�O|�~t@l�EX�N@��E�϶���b��{t��XF�HG��/�ߵ�� ��nt���@�6#�q�"�\��n�:���i��=��6H���9)�#��ե^DxI��K�8b�� ��|��n�}��SjN����>�  �__M�
�.r`ܹ�C�o�ԸB����u�U�Ae�5�����߼�rz��~Ԟꃯ8�t\b�ؗ)�#  ���j��fhnj�r��Y;�����~V�o�����Vӥ0��O8����a(`��h�h�/�z\�j�Ѩ�D�Y�v_�$CN����~��"�4c�g]��( ��� $��f18�M3?+yy�u����x��ꉖuʈK�' �y�ܛ�P�fAN]/�,;�:\S	C>*/t��r3b�#�I��
V(}��iձC�RYRݰLsv�j��U��G�y�K��ј����h[�̾R�&�jN;vd�<�}��5'X�$
s�i3�~��=�������~�>���H7 �H���q�E ���`�5����Q���Tt$�Y}u�n�7�S���&(��m�y#j��5d�N$p;�#�K��acn��G�@_��{&��6ȸJ#
���L�c�wnpa�0�k�.G�+u���oa�ҷ�g�)�T�"�Gh�3!B)H-�zãM ���Pޞk
}��<�6�8���k&�X���lYTj���dts��Ʀ|Y����Y׼Ez;k�|kU���n}j��4r�n�(��A������4��z�3>%�H�Z�	������oj�#~�r�K�>��)�.�H�S�B�g�p&��o��$��&5�ݖ�ț҉� ��"H���k�B5EQ��1f�/�q�$S�m��Z���:��`�E�gaG
3!��y�[�90`����{�U�߁^���nS�����0�E�������/�r�_���@��B`+�!G�J#w죓���[�I��.q�sd���d-Q<H��#l.U$�).�y��U3�c��X�����uK��UXL��b޷g7e��R���笯Ro!IB|�%~�5p�`����Q�(W1:�D�CC�E	� �WI��oL{?}�.�]�]�J�n�Ϡ��M�}x��(ke�ߙ�U�׽<Oz����%9�!��l��ꤪ`A��G��Aܠ��r�o1��L����uU��R��]x�a�ƨ������#��'B�
�H��7=�.�I�H�~�`� ���I����v��~R3+�:�d�Ԗ�ۿB���>�S
��|o�O&��z�UXL���TY�{ۜ���qǀ���MU"��D�0h&}D��
���i�Ά'�;߭����پ@�޿F����Wr�5�k�ES<8S��1%ͣ�U�]�H9�C� ��Z�,���az+�%�.I�7-�9/I:�)V[�n
�g�g�3�E��X���
��(�Z��Ʋ���M�	]�2d���׷}c�H>�M+�?_$��#�W�H�#���m�>�����Y����	>��3���v�n['+qݽ�m�����_CE���Qu����ƭ�Qf��uZ��g��/L�[�x.@�dc�%;�ƥ�m��-�����`݌��o����T(�����y�n��7
C5V��� �0AA�%>��?�� �� n<�S^$d;��m�u��1����i#�
b��7�Mq���I���H[>���q���a߳�����Օ^K����kIL�[p�YkN�շ��jS��JT[�<S�ҡ7di\�!�Qy��4P1QDS#����l���[G.NN�v�dnh~���0�	����Ɗ��7���Ď���Ʉ��[�a+ ���:��z��azdZLx��O2�mT����T'����1mG�b��q�i��C�4��vjQ2�ͤ�j���Ħ������-��+���a_�u�����!�S\�-�ZB)X��C"k�^dP��J�A�bF��/��y��vAw䝰hj���T�.�`\BZ����3�U�l�$�dPw��[���ϰ1U8C�O�������_�slk�AN �,�a�yd�.��y��ٛ��l8",6�Ϣ�W�L��{��ir�1�5��G��C;Dzyt'fl�#�OE6�'S��ԡ��\R��$L��.����DZp0=EK��y-��*G2�X�R+^q%�@3�DjK�R�O�<n���V�q�{��)�� KĴ���z��-�J���*����<���-����~+��M��d����5���{�8�_WY��J(��;k�[�w�`%�=�i��{�[�as^JϦ�ݓ/�}z�<�O�K4yF�!w�P'xf���	���Ҁ^跫��g>����2\oبb
}��k�P��4� ��T�^W	�O��m��c�I�Z.��p6mU�,B�M�2�� ���jPݱ����X5� % <�y	�^�>��BM�_hfx�xz�)�Ɠ�@�~��b�yd��ާR���gL�,1e�i�֝�K�����#.��20K9� ����p�WFƕ��(���IY6�%fA细�z����o��qV��ME�6�
�%#m�jp��f�y�c.�+�ސ���ݓ
���e6΋e�,N�dk��}m�)��.�e+���%�ej~���������T��Bg�)�;U܊��̭N�5��f2�1R>�o��Do1 wMy�����PΜ�tC�:��wƝV�΍��]��m��0*��==���_��EM�'GTJ(�4s��z��ɳ2��:*����/�dF8�^�_��s>J��k�4X���yK��Ӓ�8��?��T�����#�����}+@|hְ`3�� .]���=�#/�fc��R�`ᩞ����cV�`�y�e~�cu�x>M�K�p.c���9�|T4���Q��B|��y�<y^-jP"mfί^e��}�0���U��IڂI��0[i7�؊�A~�4�+�L����ں��pŅs.�����jJ��u89�W�<. H���0���/Z�$�]��.}�0�EѢu�V� Å�F�X�(,��ĳaE��8����qC���)���S�ڑ"���jw^��#8v��\��^}����ӵ��Lhl�Q��/B[�%��ufE��k��%KcD���a��Ԇ3,�Vn07s5�Ǿ��E&d�e:�@h�X������BR/R��Fj*�{NsR��
F�}9���a��܈�tC<u�Z���8jXGϥ���vP&y���qB���c���)�߽��PP��h��Wx���W��K�~���_>�.70O�jFrxF��;�t}f�A��-��G�Kh���J�F���E7W *�s<�|�h.o���f�;s����%�Ѯ�����&hWFMQ%X���0d��\��A�&��z�S؃�klLǩT�zN!���X��]�`�(i��T"�������o�W��;�RV,x�^~"��V���$Lo�����!�*!Z�k�с+LU�]����r��{~�J�o~���-��+пq��"�� �h�J_v�Eĵ�A��з�v
�*LD�Ӊ�sk|��O7����G\W�k[PQ`�5�������>Py��\Kw�[�C�識�L)F�<(Ӹ�;դ�F^�|G����q����FA���G�59=@^�M^\�T^8{�2Z��ض�J��Q�!�Yz�8�W��컪��gvRp�?� �/:%�s�dG/�V�jB�9<�u��0�I�hQ��;���1晒:��*���Bk}�����-�u�[qy��/E�F�y/(�QSe&�&�;��U��Y,W���:izU����IJ���S;�.�0˓ӣ9�k�S'�<rӤ��w�i�$
�Q+��eW7\�:�=I��C6�:V��~�,9�n�R���������k��O��*C�h@�P}Գ�p���Z^�~��:`n�h�{�y�|Ŕt'��g+����#�o�f݊�?�����ƌE���1>��h�>�}������^�Ǆ��U��ͤ�ц�1=g�ǧ��	��RR�k�|��c��%/� ���ZǍ	���`M��x��K9ȝPJ�&�g"bݲX����M��c^���׭ [m��u���T�NI�Ԅl��s@�0�e��t<���2��D�ǄC��S�v`;3!><��H6c�ԕ�0ٌ��v6e #5�.VG�4�ǈ�*����f�
5���tq9�w)�c7��ek��G�<�j� ��é��=�b�e��/�j�	�'�<��zдS�<gz?e�׼�d�
����(��"n����hʄ �PS8�I�L��W��g��ѕڭ���C�?�x�I���P�W��'b�t�@?��<�B��- .B�9�G��Էf�E�˪,���u^Ьz+zJAȢD"�u,n%
D�d,N�D4���T'!w�"ܦu�l��d(���Glq��1Yi��F۟"{v7����_�z�F?.�����}�֍D���S�d��~��l�	��#]&k��':�E#��9�`ס��_��}uZ���{O��.҂m�����.1;�#6�k2�����9P������q$J�ǳb�nw;@qm�v����%J|q��)l���ZU����E�HL
���D�G�0�[��Z�hs���~�*;Uzə^��@����q�6�%+!ؔ�`B����G�J�h��e{J�q_��~�
c'	*�Fݡ��k����=l雙�c��T�����g��wjk���*D�a�x�<M#���{�4�P��ge�f�Ե�S����0_�\@Te��F�����B�9!\Bg�_o
��:r�rO��[��]D�����zfx^ d{#��4�0���E���-MZ�6k�d#���@p�y5�\4�� 6�8E��mb�:�{�k��?�s�����xL�a D���n��K��I�����F$�@?5�T&�%�h�}��4KE��^@�q��"�)�L��%����&�nI���B8���XUSML^�_f6F�۝+���diW��G��<&&�kt�)���L���3�tbj���>LҐ�b���5S��j]�p�u0ui/YTt�n�d��:�Δ��G��O�j#�
�NI�K��>�q�N
|H���]�"��kVs�<\L���'�Fh��H!�b}�X3��ӈ�W������Ѝ�
tu��?d��:�1��ͪ_��F/S%P�q��c$�B�f(�7���(jɀ��)���Ӓ�_�X:��@Ϯs�;&�u��G�.c8�����lnu��Og��_�	�PݯY	Y�E�@��,|oda�
�2�l�L��f�5�l�z��ק�9��2l��O~rO8�^U\�ꦷ�� h��m�s�m6�Y�ᕠju]?����Q�n���j�բ�F���u{(��$u[Ej���r*��)��i��c���;���>޶ˍ�r��M�s���v�X�!��ǆ�5*�$>�lЮ>P��d�_����3\�rgf�S��yh'�:Ʒ3����[�A�6�sK�	��|��WV_�&[�vTb�~�/I����,R6���B?eHUF��\��?����I�CH���?.����.ޛ������;�6��_-N5�y��<���)<D&����9��묶����b�~�K�E�	��� �*��c�I�O&/���� 5��]����8�4����}���)��m^p�W\%��\?J-����sp�<RBe�_ Tݟ�;�q �J��HГ���\�:�-2߶g�:[��me԰�u��S�)�rڒ򃫥(��a�����f���B2v�〒��	_�����,��Y�P����Dx f����~K��3+x��	�s�/'� RN��Z:�}m��6��:���r7�<j���Ă��v��7y�/cFe��"[4(���A���R��W2 B�XoGy��iM��K�ߋ�O��pG�S�^;ahN.�A�U�d��2���1A�� ���q#u����)��TA��˽d6��G�n=�����cqIrr��Z��DV�P@x�[@&��l�� ���X����ē�x��/aI�=�w�\���WomŮH�� -���1QB��ҡu3Ŏ�-�m��B�������%�TK»<(��9�u��e�܌W�?Ե=[|��aY0�/�����PL���Ԑh�@��+�M�}h%�w0	�Ef�v��6!t%�S�r�+�yt��Š�w۴1;�Y��M*�?���R��Hr��S��A�G�"͏5���.#zb�5�J��,����
�r���
�X�Q�%�����'.:��� �S�E��<D7�_X��ؕ�8�A����%b�1����N�)/^m��(s�Xh�M�N�Oa��"k��b2��E11_�	R�/����|48�Qb���A�wo�e���냡D�'_�.q����6��
��T�ʥ-~L|\W;��__2��[zX�C�W|�\Ʈ�IK���F�F7n��Qx������Z/����rU�^"v5	��R�:S
(g^K����ڨA�aR[��w�.�]�'�]ٟI��R��]�&�2F9$[�N�%�?�s|<�#~�����n�3�:��ʕ`�UjV�ؑ��6�1q|%'Gx$��mJ"
T�K?��ɵ���>+BHNf��vo�j�hT��>3�%؃..N'y�t7��޳��Ϯ�d�m����Ue��w;�STs$����Ն�7 轶s�H�a�lD�S�ʹ{L*^y��V'�P#'�@��Ҷ��@=s�x]5����F֒f���B�{�|�o�_����\�|?������5m���{�4�u�Ó7��t@p�ʠ���Q��_�g�khpE\o����QN���"J�G)c��%Ѐ/s����}ZL�[ؾ���k)v4�cvXG�� ��C��Cg�r"G<�.����K�?V����g������[�;Ukڡ?h)
 ��V���Tۇ�������{<~:�?�Z��^��ɧ��/5>H;��o�ߙ�����	���_�,E����4���P��ҥ��)q�}��$��F�]$M.�?s��@B�p%;��^d��h�k�b[��o��d�^�DB�S����3RF����������;���Fњ_S���7�yh艠G���V���DX�|���	5۞2��S�	�b�!+��vf��|�ࡖgh��iծв#}TQ`��z9��1�/�1��;�ߺ[b"����r���^�5��?�ϲz���3�hĕj6�,`U����}�3Y��䆎��)�����S��+£���I�2m3F�(l�	�����P�׽�Ƥ �&+�"&v39ޢ�=��-�AM.4��";1˯����1�Zq�
��^�A�\s��ϡ�L�k�܈q����v�Gb��� �C�]��ѥ/�Ff��U�Ʃ,�"ʇG��o�i��<g��/9�&l���`8x�o�2 &<J^�ōE*Ib]Q4��Y�ٶZ����U��"�7Qwv Ĺh���&A�E��˕$��g�K�/z�.�"�����5��Z,C�.=�7<��UfQ�m^��1o���개YP`ɗ���l<����EHnnR�	3e�)�7)Hzō����|�]����&D��;����h��Ƭ�lor��ص�0�L�O�.�2G�ε�?�~pq���w=�3��@��O�PT�׎o-Db����y"�W�A��y�����!�O}	��d������'ßR����G�����&3.	}��bh�Q"�&x�e��4TI�y�R������{�Ǵ�:�}����Z��ĺ0�˱�:8��~^|N��z�R��{s�ԋ�h��=ûPp�`K�^�L,
���ul!��J��H�5K�#U��4�(lSb�i@��O췉4��5͏�)Id`x�j���6�j�$dI�r�bվ?N�	eQE�=hOW��ٵA���A�z�~a��A:�w�Ż=��<���X��v�LqN��xL����� ��q��U� �Pҋ�[���)�Bi��0��T�.'�o^�u��R�e-�{�&us*)��޵����џ���Y4�8�hio�jm����0����F<���W���eR�m^r�.t�F���M^!*�D�&-G��p�k���fj���e����ru.��LM|U*R�B$��@�*WIhD7��i�pI_��f
����U���c[�P�"��0�⪢ΎkR>�qB�6_9j��)Cu�� X�ȷv��T�ֶP�H<75�LW��:��e�E� u��V c��L�{�&s)�2]��uAGZ"�}�o���d����C
����l�V�tٍ�����c󖶱����������:�h|�ޖ��/i���zR�S�˻U�p_C�6�N�1vV��-�ٰ���(�l�?�H}�i�;��<gmӭ3��p�%������@�Lc��D�Μ}��i�`;��h+�D9�h��M���p�f��HX�{����A�ߧXw�F8��KE'$p���n-�s�>�BD�>�7��M> �ϱ��tO���_���'}?���Ze8�"GI�R���|�L�tn3�͚��S�*b�Ǒ�U��Ey\��%%"G�!�m�"0���|�����8���I���t�F���l%DT=�l����u�1��b�2�v]9��q������x�?20�%�{?U�� ���&�IIv�U{s�x3:^��2ۢ��������� ���E�9�eBc�H�cp��w�d!�M��E֦����[��f� {ps��P=�%�u���}�{�t~���L��쏒�u���<vK��V��w��m�Qt���-�-1�1&d���d�[/,"bm��x��MiKR��ѯ����G��75�Z7;$T$-k�"�@�Sp��|D���uz :�܎���N
W��`�]��	e�M`�3��r��C�"p3j���f�~��S���Z�!.Ɂ�1�}`��p��N�����"��O�	d��	��Agv�e�y�K��݇�X��[���Bp�^̯:r���jA��c�;����}�����1lw��w���:�HR@Vl����b���
�+�dσw��hD�ʳ�x���j3�u��z���DjU��O|z�'�H�(khsv�n���A�?����'�'+�:��,����)�q �B�����>4`�W���%߹n��D���c���g��K!a~����w��5
%JT�D�T�f���6�#Dy��r�`Վ�>s�%�5�&ζ�bȣ�ȿ'yX5%LO@��*z ջׄ�������Aҁ^��M�|b�3���j-�U��h���4b��l[э�J\>C�>��|Y�A*�Y�[�������o�%�{y�/�?�۾7ٙ`ng����f�'�龶B�K��%R�S\h���M�����-@��@��t\�߿{	k�`$(~�TT�/틄S��ǜK�����ҁNXUiX;k"�Nc��N�p����i)����y�g���i3��$z�2���VH�x�����n^~�{�r5볊��&�b��h�
���o0̆-�l^J�Ձ�f��gA{��ϵ�s���3gS����'�Y��4bs��r�E%:>�9���R� x�����C��[�kC7�GFP�� (�Bk?�N$�bam��,��va>�q%����+��8o�p#ƒ������idO�j�U
�i[]���[)�-��M���P� �<�y
[�7\��o,��z-���Pكd�6���F�7W�f؏��H�\/1�9xz��4 �W�)��&�g�\z.���}$��cv�5,X�Mj�C�P�R.S��lo��ʽ�"Q�Q�5M���߮��XL�ж��.�\n��k�`
�2؍=٢I�q��4�(��s�H��f+EYTB�)�0\QS��zɈb�{�@)���i9��J�9���\4L�يIF?���&x`+0��Q�IxR)2�&��,1J��U�\F�I���h�j�@X��=c��܊߶��]˱��.��]e ZG�
ޕu�S�: 
�n��w`iSɅ_�����+���o&��0�5����ӄ����:'���ԣ�
(K6p�}z�\秊øW�h^%އ)�L���=U��~�OX�d�x	�Ӣ��ǖk��<{�H�p�]��2cB)�jE�} (1��Kh>]V�-��%	��h�|��R��X�:闎Y���F����(�V����cJy�߾�#�ǟ��[��!��Fl��HmYԃZ,U�U�d�(�4��,k�R׽�kA�D&�c@�i��_�~
��rJ��Vz�B�EI�S���1L���?��%�X���o8���s�
����k�@�!�S{H/A�9�6�cgS��������|tWT��哃����A�W��4��(#��yC�uvh$�x����,d����0��.]��L"B�fS�cD�K��}y���q��I8� �i� b'��Yv !%��{�|�t��TAeC�+#Y�6~���=!q�/[��#-)��8�ɽJ�C��PraL9�2y�@%\qi���>���~CZ7���v�Md�ɻz�qEI�ˆ?R[�i�U�t�S�Z��S֕�e�92���������I�t*$�D���/�\,� ��I�M��o�#c[o��[SK �5c���+%_�$H�p����Q,�D+4��_��}	����Rj�^"J�Nt)Qc�����Y+MN�/�2��+����/���@yNIU����9Eƀ�����5�WxzbVi�tV/D�V��b+�TNUk���0P^�jkU�3�,]�3ͮ���.����r���>���-]���lE�;AM�J�I�h��0��C4���4S.x�����.L_�5ls�FN�׳�p�P�+�w؍q�ק_O�R�}?*�q�?jX1j���Q��A9���>LZ�x~��8*�׼����O�s�Y��'�"���,qď݀�ͤR��7��L�x.J�`Y7�A��T�'�4�/D~�l_��.�����hs()W�T�p��~F��"��K�����0��Ȝg�9�[�Z!�x"�~AS��(vh�.�d	�.�� �`�c������	t�"��g9���M4�� ��u��Z �$�~vA���FH5M��@�
�o	�0l���)Z-�+ve���*e��S�y�QW�F@ѕg�Š>D�Ok�&�f�_ l�%BE7���q�D�sx-�Re� �WoxB����5f�?T�s�ȧ��ԝ�(7g=F�{Z���/f�8 k����&�E{Y�56s�&���.}o,�EZ��W~��E���х��1�'����]��;ẉrwj� |)�
 8xN�]Qf�5u(��իKE"U�g����wU�^dt�v�PGYOV $�﫿	���*�l��Y�0�%��ީ�9)`�X�@K�3zf�h':�9x6,m��N��>Ҥ��n�x���J���1��R5�D�"/>�W��+���g��P[GN��6��=Id?iY*O�Х�W�D11.� l�j�'<^y����,�yau7�v�a�ٸ������$��H���VI7�X���"Z��@������)�V����~�	��)u� ���+є��8R�X"�KNa��L��Ȯ߈B���U�@{o���տ%��/��Y�Hy4������m�`�O'��UTX�=�͎a�>������P'9�a��Q����ŉ�J5�����`�ZG�¶s���n:��{�:�NBog���Y�CKC��G� k�2�L�MC�]b����Y�e��R��q�&��P��lCQ���901�$���ϣV����x�Ԭķ�&�16Ȝ��W�{yE��h6ɨm��Q�
������`ڿ�1{QMf�2 ���_��Jl��!8[�i�F�W�C.����51}K���6�f�����:5b�}��=���0p���ҿ��:��&�c[V"5� �s�O�� �������fjo����
ڗ@���'����Lw#ȱI4�ְ��5�5�d��"�KA2=��VC�{�b�O��
���/��I�Z�����9�ƹ7jT�.&�@���K�Xk�E�[,�`�x�i����J�ۃPܮ�W?�F���vs�҃-���'���n\�������,C91��9!���ޟm��mj�������|��e1iDK��0�dqK���ꑍ���gƎ���AN8�������Ze�s����eN�Yk���K�u�?��xU�n�sJ�
0�_V\ѣB1���Z���|�~��M��H[�����K/�Olnk�p��a��GSl�D��?�Ǣd��-4�D1�
�j�E���t�g��2}i�޼�	�H~u�5��� �P�v�IU��f�
[�#Y*&?��M�$5Ոn1sd��:�]���b�!a���B	¸����s���	��^�<M�V(�š5�3��
�fէ
7B��ͷ���Icc�ȇ���*g����5�G*���o����p�����)��7pz�U����:E�h^�a�8�v�	�����j�U�n^,��mTS�\�_cRM��.� .O�q 0 i���ٺ⮐Az\C��XR�B]����˵LA-� ��(�3��ш����������:��%��n� b�PV/λ����n�#w�%\��}�����>�'o���m}�êpF��6�Ytj*�G���⿟n*H�t�z-ûc�S��F�Dw}��F�>K9�����)Dobr�J�I��om�hQ���5ǃ»��Ò��ᥰ�\dߌ�ͽܡ�OەZΠ4X���^ڟ*(lN��\1�h��-��*�J~ID{�4T���7��o[*���Ye���71�����I���l���Y�	�m9|,�<.[S��Zl��mw��O�E[���K��"����2~H[R�B�R7f�3�>����07@nҏ�vZ���X��)f���Nܣ4c\C}�3�x:ƭeF�Q`��Y�c��	[3"�\�~�.��,Z�]�G��~�_9桦�TuiLa�%�}�2�;�r�B�X�֟����D:G��H8���ot��<ѿ�+p/ܸ���Ӛ0!���JC��r�WU%��C2U�����2_V;����3����|��N%J���{7�H���!�UH�(��ݧC������5�zP�fSoc���6H�P���S��)�V�ѱ̨@{���s��rG{�~�1_��:�S�)V���7o�w������aa�<s]�~B�E��Og^d��'�b
u&z(w0�6|{Ֆӹ����]}���o[���H���R*�.��ڊ[�q�W��!����Z�3��{rO�Ӛ���mҐ�!�q��D�>���28��"��jk{y�h�]�*��ܗK�+F%�Ը�T�z�+m�����^���a�^WalG0�
��j��NP����=J�.4�g3oN��.�����->ɣ��)�u���X'VCr������
j��c�yuZP�F�T3��J��!MW��BƑ\ĢEQ���܊�||�l��8\ �|�`�����hi�[g!q(�k�[��B̎MFm������+F��kԝl �[��zc�O�5GF�	�49�ASe̐��;Uˌ%���h��o�������0R`�{L�����M�U��>��C�!��./aۚW�����
BKt�?�d�fّ�$�5��8-Pǽ&��
vf��U�lc��e��F�G���G�M�@!����B�-"�:1����
ЦE�]J�ߓ���k/%����ml���k,���ƕ&��1H�U��-��L�hC�2K���������5:��7�+��2F�)�-������_�}� -D%X�W*���vp�TǸv!�z���5n�cB��=�|�޼ʻ���_�JRdf�@����h*��p9,�k=p_o-�k�%���̃w2���!U���Dz��{\��J=i�z%Dk��Û��x����	$е1O]�����Q� ��.4(d;/k����p�g���"��\�����u�1Ѓ�0ᚥ6���z��2�$�i6�r]E�v���4�Q�}:k)b�)]��{$���l(�����*��y7D�jx��>�w�c��S���;JS�e̅n�?��6\n��`&H�����Q������3t��s���]�UK��`a9���'�;��l��5�xbY������aq���uTY�I�F��"������\���ɞá�L���[0���7w�B-?�������nR��i蒭Bݾj�$?\!�i��zE�ѯ���9>LPU�{e:y��y���=�cƒwO�Q:J ��f>���>�^~N�c��5Q7��F:d3�S�� 񗿀.%C5�+q�N�����������kWU���`�w~Ȍ��4�cA}�Ә��|�n�Y͈�@
��I�t̜&��'
e=M�ިOG�"��rBψP�:��H�T>�o���#Ч��Dy�:%dpr
r:Yg��';CV9"�i,Ҭ����0���?�w*�*�Zi�]7�⇾vBL�>�Ǥ���Wm@r�$��Dm�5��l�06l�c�'d+o*h��2/|�
�L��|��f�]�l'5f��*.��\o!#-���+��_�A/���m�����?����u�@T#C���?s���|Ό�W\�m��9�:Vdm�`�^��e����.p�g�6/��-K�.g)~e`��`���1[�G���{�-P��$[���0��%��f�f^pfQp3@����xS¼���F�iq�8�3C�n�usc�C����0v�
�2%,e��*�M���5V�T�<��_�?L�$�5|�s������뱿e��эCj��?%M����s��.7�aẝV�S��0 �ݼ,G�L会��"�O��44�&��y�Yl@�m?uC:�\ծ/)3��qo�_y�ұ�]��-:��?�8�#`D�[��J�! 6&_̻����Pc�h_�F�OϢ��nP�ʌ���z����F�R���#(2�3��6�Ur�b�I��I�X/(��~\�4]]_JX:�����@��U���fM���%�h3�}�ƊM�x�BX�.kt�x;�~KA��e��6�ZvR'M��{��W>�s2[,����^#+a��v���߽��z�b葝ch����g��.2���t���� �;�4)H.�g��/�2�7���&t`�����Ǳ�x�'�Tk�%⎖p,`��pi�:.\�^߱��ҦSϏC,��h�=�,�<�ty�d���Y������8��3X����Y��p�X�c�jGw��8��PDc�.�x��A�󫾜D�J:e�?~���?�?���g/ì�v'�̽'
�n�9�,�S�ݮ\k���a �k�z�����z�N��"a�\��=)t��$+Y�!%k�{��,����1�k��p0i�j�$~��}��a���pчDE���k��ﳑ^�P��4k�Y��=S<���+o�|s��re�R��h��t�0>綻������߅`6�PR�,\���z�:�U�&�a0�g�6ا�����	�G�b
�1;m�%���Lp6����j�:e.�1ĉO�e�&
�̾ٻn:�ٴ�RC���\ϓ<�R�Z��V`ݐ]ˏV�E+��%�������n]���#"8+�Vl��M��P��z*�����]R'���s��x>��(V�Z+11H����8��yz� <H����Y����d��[�x.aӵ�YL�	�� �����Pa}Bt h��x�
Q���bk���mN-o��U=���ê�S��X�D^�2"��E�^2f	��? B���^�(]��Hkm�Z�أN�v޽�b�,f�W�����=*Yi~r�qqz1\[��L�*��Dd�1��1p�#rB�C�*'�$qOO�g���t��il峈�L��q[P�a���ׯr�m/�M������B��DOl��&�-�?1a���O��L�ߘ/�S3���w�h����)�	��:�_^��t��?��<|[)r�־i�G�yK9���*����m�zq]-27iGϬL�]�/:�!���, �'�x?+ʛg=%+9�)�3l�P�L����y3�G�y�<�b�-�ƾ��S�%��Iu���3��S@��Ŵy�e�4��d�uG��Y?z�ž��=gn-z���~xE���c����g���Å���}�C������]YR�֠�1��,�}��AP��#��V0��	�sN����*�<�j�2!��b�4�M��y:Q^q�(U�sf�7�.����)�W:!И�X��+O��C_�<#��+���i)�*��،l>٩�u�ܒ�jW܃PP������x������K�w %!L�?��F�x��B�(�^�a�c@��Y��!ϋ�+��Ҕ�:<�f ]�hL�2ڬP'e\GD�X���J���!���&c�՚��U5��h�O~�t<߀���,���,�.Y������7�B��k�a�ky1��R�0:0�O�Ei �P�I�#W�3�EM��f���}�����,�c]�+��[+��6z��gB;����}zC%Ceac��1	S"�A��bv"r`�]�o���C��ȫ?��\���j�_�*�]ʍ�B����K ��q
��S�m�/��@����j���>(@��UJO�S�W��@bX�E�P�5��{9	��~� \_��{ ˌ\�f2t{�$����#D���P��á�O~,*	y��ţ�]z*�M�2#�݆�5�(� ��"[[��*Y��ȍ��FJ'�1�"*�^s�ʼ�M�cj�R�GNj�l�YR?�I&z�H8� T@.!�W�0$�ʞ����Qj��KT4��*�y��o�!�t�����g;���{{:���'�M�W���R8o���Ş���[K�f���|Q��Vk��Ga�f֔p�w.�� ��Eω+��R!��\d�]��a$���&")��-�C8(�f�+V��C����z��"�봏���o�ɪ�'�(�l[7�������A���i��)�g�H��EO�A!��B�_V1J��G֯U���gr�
�)�j��pQ�Eˢ� �@f����ˎ�3N�P��}�9��셔��b?��f�Ԩ�i�)�i<�UQx�ة����[�V�>v��~�iT�.�L��[����f}'1?��%�e�./lY��)�p�G���#��yc�S���h�M��E�{�OH�8
i��6&~�`�X_|�! ���d���9��b-��᪲?[`Yd�B��z�����eE�6\���Ymb�;��[��*���dI�*�������;���.�U�\�6
n¾��;-o?M$�85�
 ���& ����}r��Q��;3²Ǧ�Z&�WE�kS&)F�3o@t�]��Ç���­x�6LSV�_��kDC�7ֆ�h�A�ƿk�84 ���(�)s���:�m�G�PND��/���B��Y�ϰ ;9��ޗ�b��g��0Ѧ�&N"[q*�1-��e*$�KAd<K�AX�2���Elp�d�"����w�o�����8��D�A�i�I��j�����ͅ�_�� 1V�}��]XD����7�_:,�Bv��R-D(�)�fa`���LA�-�ZbQ��X2 �8�2{�l�B���Nj��-D6H����՚��'����v1��[��ǐl~�Z�Gj�hbǷ��F[ү&�f�~��.�2hF1e�@_ҜJx5L.,�b��Sz�W��i�܅��|�e�|�C�O�Ȣʘ~�`��l�����
�(� �gK�1Tξ�7��G�)���p��A� W�bM�q6�X�`���fj�]�#��;ȷ$���~E�-\��&~U�T��Rk�%�8�s^�[8Hm��rs.��ڡ$�I�1slb��W�v�'A��:����Z}0�K ���3�"�NԠ�xF���~�+;��L�fy���R�f|�.��u�X����H(�����)���}���O/�rǅ^r)*��<�}�{b���d�<�uQRGJG�V��\�$��x]�ܜ�\�l���1��P��ڝ<݇��>�������z:N8����d�!}�Wՙ���6���� ̺�%���|��J�J�|�c�tSM���	����_�y��#����s�e��>G
::����:�������7}k~�4� �K;!�Z1�쑤��v}^�D+�����6żL��d4w,	L7��PDJ~�٬��f c,|�N��J�w���FR-2�%�UfLM�x[p#����2�-�]g�d�PeA�`J�R%.�l��{��G|�,fͰ`��ie�%�'���f�f" ����\��o#����R`�uJht�����5�!+`q�81��}(�>�Fx5ff3���x��2 L��l6;ҝ5�-b.�Yx��!_��3��2��4S~�6�v���Sr�]��z5D�j3�%�VԽֲ���Mi��5Q���}��@��]��|^�F���/Ϳ?aQ���-d#�� ���9���u�����c���x��v��s���3����)���\⬨N�OϏJ�^��kR�����"G	���K��F�`J��m�ӅI��ḋ#��T�M$��13{E�>�у�Ex3����yڂ5B�W�9�D��~%��A��p�,?�w������ȑ��c���3�7~~�u��6����Y��ý��M���L���7�6ܚ�+�s`� ~F{
ϫ��Y4�gq��W�PoT�)���U(�觧��da�}0�� IJ-�+�Q �7ţ���)��<��mE0<';֧��d Nŗ2�c���^��&�a�Y�1��̈́mາ�9��D�L]܁1�~��|�z�c��J'��U�?;T��!?���^,��7{L�v|Դ�v6K��"�1`��z��j#�V�u��݆)�U�Tň��de���b؀s0(�w�wي�k�ɂY
U�@$s���f3��L�K�iC���Cp^"$~,��,�H��|s}������F�ح��?�� ������V�tl�赨\�a�j�ַoc=?+�: cv	��L"Ӥm���t�ˁ٩�Ȑ�T�� 	����h�ݑ���#&)�Y|`�k��t'v=��鉆	]�F-�a	v�Mk�=j���6���>���&#Ǘ�rF�+:������n�Ȃ���Q�ڊ8<�fīk�o�����/^$H�@���}`�N����h����/���_p�\���$���%���z�ey��p�/��z/E���d��"�'vwv�l~���D	w*<p)ƍ�&6\��@yT%.8[�v��=*����Am�)��Q�k?���e1�c���ҪŸ.π��M�|8�ʕ�JP2��~(�1���~νj��oR0�3F�_�B0�l�#�![x�}�
}UKV�v��@��H4���� ¤�'j����(��y̱h���� ��3�A$�Y��$Eɱ�F�2�y�!����4������;4�ǽa�����>��h�(�c.��ζ��'�-��gK9n9:�y�Ab�ɂ�,�3�p�%���[��[MR 2�X��Ċ&��s1�ƪ��ӿz�b�*�	#�(��>��j�lJ���{��Uk�SC��7F1����A!5�Z�|xL�@ ��C�����}��"ƍ]sF�Oŕ�H~�T��2+�ǲ�ٞ�x�i)�o3uP�L���X���Il�f£�Z��³~�+���4��2⧘��=�@�����p�(�|��=�$�p=�:�����0G�ѹ	o�X��"�[)c얥���";���}6�(>c��bw|�	�H��
����R�������W�
�ص���]�fq�/��D�{iIt>}=�� �e&ϒ��TG�-(��I�KSQl �i�tE�s���U�OX��w1�aw�LL�'����_����X�[�N�G'��6���O@KmܸAh�R���&�=��<���BURt����6���C/�x�E�h��녴�U�K�����%���J!ӛ�\��ۨ��.ц~.� ��!�-��>�(�@�j��#|��%�@DBn�u�ٷ��J4K�w]jFZ�H����7����$y�YH=T%�1�h2w�,z��$i�5;������b:��G��ޙ����lc`���Ols{:�(�rN��~ץ��g�`����Z���S��d�!��*w��D�G��2�\�����ڷ�"�Y���$��X�Q{hc��ٵ �OI$g�5��c����mk�D������"څt�w`���07��`�~��	�T�+��_��H=���ţ��FM��?7z��`g� rx�>�2G��H\a�wp/f)�.6��D.T�RZI�h�E^�!�f�\���"�y� �㺵��&ѣHo����zq�y��c ���L5�yhP��&�ώ�L�7�i=ŃiLؼW�rU1.���߉��`�'Q��ߴ�:
A�@" �:�>��4枪^"o�������퀳�qt #Da��]��!��A�Qʨ*�����}����	:v�h��S<�U������[�R<5p�K�'�����r��Z͌��� ���6y�<��BO�ć����� 5��ck�m'X ���Tp�xGĳ.���Z����Ѯ)��8J���O�m�e��m�_�5B'����� 5�ۼ0�ї�2W��\��40�1�����R5A<2r�,o�l���z̘_)�cP���i���a�� &�����̡W1{�q�324���� E�bf�ߵ����pI�q@����:�x;�H���3��:�j������V@}��]Ԧ�����s�~�25�M�7��p��D�-�#�aλն�uQO>3@v���R������ךJz'9�8o�G�5}d�Y1�4V>��8���������9��~	L���u� $�.��b�'�>h�ߛO��0����ꄑ���N὇�p#��78X�X(��"Tc��}j��C1|����W)��i�E�v	_������^]�8��H���������
$�9�`���.o_�i�ٔ���D���=�9�z� ��9ͩ�%���W-89��+�H{P�i��7?^-q����ԎџB�ص� ��My��=鿮)��,l��D �&'?�Y.�I�?���|"NYU��%�;�iMչ��D�pT��:��'G3�Hd]ks;�z�gf˱2�c�e��@�II�����<�`vP���ݰ��z�OT�Y8��f�E��ɠZ���v��zi߹u�H���(�I��_��ĺ�I�Pj��6�Rk�%���9�G�����%�)��2��5�K��LVg���f�4C��?�I�J��z�Bb�%Ί8����d�����ɋm6���!C�G���*�O���Z��[���k�@b�^|6���b�f�>�@B'�[�R�4�Y�>��H�&N�A���H�� d=��wU3�&a$��z�����iW�zcl�sԳ�aS�6��h������0����8;4��1�ױ�����e�!Y㼘�L¯ph	��P֋,����4�,"��ֹ��ߔ_�^���`U����@@(�X�KKN���e\/�~&��&+R�� �RO�zH^��,\��;|��P��OԆ�G�y+�BJ�shv�t�`q*�(�Vɮwt�:�0V�Wc|l�OME{/�Z�F˼^��el���E��i��B�Xs��Sj����������F���53W?���>r[ɣ&����s�� �E�SD�@�MRƮ��R>G�p�t��@�fl74�&�U�V'�����t)���k|���@3�m6Z]�S����<Q�z����S bf��P����^��9���ޙ��
�iޑ�s����y7�������U�H�3�|�x��)�\��}��ͩ�#�L[���@�~���n~&�Vl�Q�g�ʼ��y�֢vN	�|e|Jp=�qSj�����$�n��A	���v��-�B�_d��A����N��u�I$Y�`���5��w:��/؜&��Tn��|�<�f�(&�4u�
�o�F|$`[)хy�_�l,TC �p��Ur�
�mk���t�ŕ��
PYT�G̫�9F.�M�E`���l�'#]��mu��Ms�ab&w���b�U0ꋘ#����myT���E�Y�+����P��c��C*��s�c���A���p���F�Z!O�n�k��r^�#L�]#e�3sD;�;��ur�z�$7���e9������W�T6Œm?l�j�
I9�M�7A�m�U�W[�OP��1�T��h��S�jg�
��9����"�!5L���nf�̈_�M��6M�h�"�Fm8/��W�Πr0L�sX�jE޵��Ƃ�&fU��P�mu�ȶk�I��V���Q���D���e����#����ᆓ:=|���ʨE5����QR�{�w��M�`�q�����`�/�O�%��]Ox��A�'��[(���U42{̾3��εX��fV%gm94Jy��������r����C���Hb�^�O���4Uh,de\)����)V� I���'��a���BHb���U�M}3d{�I"'�l�q���ܨe��Gj_('��t;��VJ����1f&9�;�F&%Y���#�d���X��"��!������[��U���x̲�룻p�$�8��.�j���Np�"=�m�j����;��	��;�A�v"���9Vyh�o��(�9�16b�
d�$�/�'����0!�{���q$m�J��f������`w->��+F�Ã6n����c���l{�ZX�KWz{��~��A8_M��)E㮰=P�}lJ�&�6\8İ��:w6&����׈���>�	�nYAt�����E@1ŕ�Ll��D6�2\�|��(��r���8�W�	��EM7��o�xT�Qϱ0�~�l��9�17uɊ��Z[��V���.3�����(,�6�A�Tw��
�KC�b�"��Pl k-/0�7bLv�s$�^/a���Zq�r[g�u��7�R�'���Td�|����W��1e��cH��*T�-Մ�vj� �c)���<*^
��$�MU�Ln�J�m+�iPj���%VT
�g��H�u�N,cɟ�Օ���t��\���XI��.�dR�챃����oe�at�}�z=�hb�s���N%0ۖ��Ȇ��^Z>$��!��u\컖��J�� P��J���GN`t��%OW�f��Z���'����
������7n"|���4\�U���Y�{���P a���?��P�"b$�G
1�ѫﳲf�*�K`~mo�iW6c$!�R5CgdYnI,}I�$.�hG�~tC$U&.W�N�V���W����1�6=Ȑ�6\�F$2ы��D��ʷ�E��prT�
0Ҕ��x��d-9�9�U���&Ct�{`�+��[�Z�g�T���7�պ�n�凚��X�H[N!��b��tћ7ic���ƄB�Q��;	F�ǚx�ܣ�EC�9�$����ʊ��?���,�s45��F͛b"\���z����mҕ��>�������qXl3/oI]��w����^:� �׫b-��D-a�[p!.�a���fi�1š&=�2�z�5�)��vXX͂�yN��ڽ�Q�xt�7�׬���ᵓ��5x�'FS���@7f�ҙ��k5�����<�8�1��0���E���Ef31=�������:..�8�N���hu����[�Vrr1o����l�]�o_�����*Ih���i�p�մ��ܝ�&228�Ŏ��<� /�yBP���+��\��m��֯�v�����]��9_��̢�e��!��<�8
<��_=i3o�u����Ӛbޔ�]g䨖A�����B�1�LvȒk��x	󕖊%��Y=��W_x�Ù���$��*���3j�U��`BI��v 6$�<�w��w��%Ddʄ�6�+r�U5�����3f<��R�y�MI��S�OWR�<gp3��Ӷ�M�����)#�C*E����,Xvc�pl��5<��{�.=��V�R�zA{lM�����ܬv��xm��L��6�n��v�/�7ﲶd.���F��"!���p�S�g
�2�nh�K�`^��O�=�;*��FAב'7����U9�W���@�.�n�ϥK��	� 3Y�T�����b�Ŏ�#g����{5m+G
���V��m&��3�7u���lb���>7�t	�|���+��P"�Q�C�}�|���E<��i|��F���h5�b�Ȳ�g<�4����D6�6�nD�)Ԟ4MV�rv�_jop�;�;0���;�1��=�=���'����UQP����YVj_�}�������#^3��m���1(�XOG��Baf�)��dz s2��Qbz�.IZ� �D�)�E���N�K5L����\�������i���6g�Za_���;#�k���=�@rZ��f+�+fs�ϳh�b�\�&N�-�.�@�SkY!�]�7� Y;� �RfY�fL����9�P
�G�3Ǜ�ϓ`3�jÅ��<))�6��D����2烟��6�!�;�.�	�B�MU��'g:��a�V?�c+�o��t{50扷���c�H߿&ǈ��D���Q�ԆD��B`�N齼1��4L�m�K�4���7fI4�u0V�Yq��tX�Zd��8ت��?h��i�P$��/�~W����,$�b�~J	ܗ�/�S�An��u���)7܁��9���)��!f�_���[��$���&Ŋ��F�i��L���cr';��X(����7D��i��$.��5*֖�!O��� qJK���������c��&��G$�`�NV��>�9S�U�dz�D�C�<�*�9�s;���ض�AK ��>@�g�`�*�ȩ��(1�*�ǃǥ��=R6^�b��]�S�~~�@���8��d�S��u��cy����%�Yz�ƃ��UN]�'7ldZ�ffYn ���[̯Qv�X�C:e"��K%-db�^��k����:��v,����u�1ó l�#�c�I��?V�7�>"cx0�4(�/�<)���4����߫����� 
f�(
���KVr#���?~�V�r�X�2uE����'MAud��ҩ�zDS{/ F��i���D������r�N�)J8��]u�|�	o�	O��L|�p�wv�L����O��h�a����ѥ�7�]jb��/@J+}N��T2!�k�u���vR:�1�����IN�):�ya�z���G��ՏZd����˟�R��!Y�:YU��Q<E�FU(!��s���2���9I�s�߰]Ktx�Od��H����]�k���)�q-Сc3~:]%�7�ۗ�#L�G�:Z1F"��}.�7���묜��u0�%5��4�׫ރ毎l�f)Ly��]�G�규�mӝ��ɇv�hVh�I���G74G~Zc~J_�H��y�X!�W�rr�yf�3m	U�L�б�Ӈ��x�X�6e����e�E��!�H`eo;:rbq���ҿ��)p؇ Le�<�I��/>�4�3�L�S�3�[��ؠ'��A�!d7�"47��A�m�[���5���b(e_�'$(�T/F��XD�dw�so�KFnӒOvTxڼ�M\��(*��G^ŖJ$�$�D��0Y�SÃ���I�.��U�IZ��D8'A��Ų�D�;O��)��������7���֬�A�@��0ȝ}��v�����ț<�e�t�ӷ�a�vn��ȡ[J5>%ηiÁ�7M�~U6G����mmTJ���h�2Tg�v��tk"�,�ڼ��A	4��p��d�-��.�D6�0?�R���f�%�y�v�,_��\�<�0����{�q"~M'�H:p:������tU�6E�HN�V٪L�L�������T,�3��Y��рQ
�Ƣ	X�%`�&��C$��#��b���=��9o�վ)�O�ퟚ>��k�q�/�1k
�&��bٍ�i�7S�4���i��V�jX�k�p�P٬��q��Ԟt��A8E!��M�ߑ\���R�J�l�-�)r�>tCgP��[F�/�}wa@eb�ٝ.��x��%�ٮSx��,6M��r$/_�S���9�1���/��jim�ڴ��/<cn��lS���ȼ8S��7�^�l����H����CZ�s��@������>LlQ��D=G�����5����|��ot��ѫ�5�'���Z��r4�lr�!���=Ơ���+!f9J��0�>2�pT1��E��G���%�2�-�PC�z��y�p�0K�*�ոG	����w}���W����j���	�o��AD����!��MKx��UD��v���h �N�?^���K��Q,CqSSڛU�y��+?ɅTS�p��񼽬����~{8���f�x@��u���j�e�ׅX7〚���@���3~I�n�nh�x1�ՀT�3���!Y�+�TR��n��]7ߎ��u3�3y�fټ���!�kO�~���б���@�@_W�����S�"Ӯ����gfxU�^/^S�YkJ�'1�p9a��E��(t6�P��/Ľ}n?*�[�Iw`��'�������?�$��W���h�Ƅ�1����m��zJ:2�[ ��)վ}��[Vk�m�MB�T>�y&�����IŬ���3�:yJ;z��8�8�h>���
�������I��RQ���f�цlC:e&,��~�{*ϙd?![}?�n�Fm醾L�k��vٽz�,Wg8����%2}[s�`C�ڈdش�@z�Gy�a<� �bs�핝u��yI�c�[��s�ڋ?�$������6�_�8;Ӹ�'{�֯�A��V7r�g�;�«U��X$��{�P�+Ǒ*~�����f;��?Q�|�����J���'�D�7�i��������f��q�Z��+.�]��MXڙ,���G*w��zȈ��cKw7peP�\b�M�a�l%צ;>߻���G���J�l��P�]��S�$�[k4�l� ��}*;��y|o_�9��l��
����`�5���=k�M�V�d�Aצ�ǋ�b�ۄa��_ U�<���$[��AtD�2�{�1�]�tϤ���>�yh�W$��mx�6�6}�eT�G5�7�cW�	�g$:$i?Q��`���o��*�?�;"�yJ�I�bޡH��\7&�|4@���H�&z8�a&��$��E�x��>W ���:X��=ĳ��қ7B��n�O���_�S�ʧy����sV�D���K� ��(r4Et�^}�@A�n�k����i�;���0K��S�^����b6_�۸���M�)��	�����KNFu�ȟ��گ��2�\P�N�r.� %������н��{���G�2�qr�T�N��Gx�t� ԽmڳnY
�iTzh�2�&�I��i��{-�.;~ܔ��3�	��S������2��7T�HLhv��y៺l�>�W�t&5�A�;p�<��,�~;~�>�$��ɇm�	���Ax���@љ3;��83s��2Z�1�-?��U�e�_e�{+h�
�Rզ�ʅ��=_���Slg ?X�`c��L5v�1[1q�8"����Y�=`�z���k@�J$�*�J�h���c��p���aDՙ�(���+�(��D0�^�-���ٶ���g��T����ʴ�b
�[c5ƺ���*��Ǉ$e�6޶��������E�{D��7�z���௻ީbjC.X0uY����-HC�+ q�/�������XmA:��'y�8�1��	�}
!eq�!06+�*�<L5�6W"��4��*���^�U~����Y\z�Dn�l(�Z�=��ԃ���3��!e�]�^bR]- �����}�wW�b����,l�:�e�@��a�oiK0A�k����$��!d[��*�ַQ��x �|��7	a�|ӷ�
�&�l,�itH����4n�X�����GQ&�����[�R�^ij ����z�F0 p� P���#�Jg����ȋBA��	v���g��E&\B�V�?�x5gN �����@>UdvW&���7���,�A Q�����ɖ|`B.��$�2��$`�o8s㉏D��L�;��I�N���q?��-ډ�J�Rh����M"�Ř�X��À��O��#:�3�&џ�ܽ�ĩ,����>�5Uة�sq����|"����)jDѓ�o:-Jߖ��ʳ �l�~L��E�(Z���.�W�7u&c(��9nk��.�L����Ć�lW���&`
$�Rx?a�O���8��sϠ���b���������u0E��\E���8�k��:a�z��:"�c��yO��-�m�g�on��E	N%}����S4J;Tx�$�(�:c����ׅ�����5�Bӧ����;�/�l<~ʓA��_�;�C�Xuf�����:1Il����[����I����7s`��b@��,�or.�$/htI�9��o� ��[�������"^#���q��+�3l>��7KX)���	;[sy��9\ܠ�}��_���qA�����'���]'�x���:ե�Xy��!�a-,�u?�t �	C��Evl���.9�#����Q;������L�ߤyo�D|����&T�'�S�_{'2T�7q�i5�s.��6�ҧ��3
C�7Tۘ�B�#س�4>�D3P�*c��<�Pr���؀������R���c�,���I�8�3Nq�@��$��Q����3�<�]H̙���w�L��R�
��m]�Bv&�J������wQ�Z'��/��y:��J�'�>��Ӂ��m��� �՛�?Q��Y���D�U��kQ[��!�����X��ҮһШ�l�|�����zr�
�a�-��޼�
m�]+�WմڬkPOS�gԣ��E�4k���[۹6��Y��};@�w?mX�ط��`P�ۓ̻{AxL�s��r�[�MGQ.~�=װ&?,���1��@�:�Rg�Mpx�r����Q�
�@���S���PU7�n�I	N���m07k����09�6���x��GwRܙzAm��̛���/�,�"(����sn� K�Dӏ�{�����s��O�6o�р ���e-�<&~f�hz{�Z�{{�ڀfE��DQze*)����l� �*9�i0����F�S�E��@�p���>pW���w��i�pZ�4Q��aL�G	�g����+ʖN���rx�,A��� 	O^jǡ�q��5ջ��s�|����Hr�G1$LA?p�W�$[F��pd�r`9�����6�شOwI�칙��~�s������;�ҙ"B��f]�8��|HE|L����六���4o�T{���6�h<�Ju0��2�:>#���
��]\����J��:謍��g�!�ׯgGx[�:T`d&��A[,�*�v%-�X)]���a�k�;��J;�U5h�5��.+jo��׽i��QN�%?/|>��fy�{&U:ׁ|�Z*?f�d/CU"��9!)$L"�=E���� �<���k-S��/=N��1��1�b���6������;�ii��(����4&�5�|Ń��z��!>��I����E��&��Z؍�đG��Hi����%l	�r��Xcf�� �A��UhV���S�_Y9�S��?V�=Eql�VCbQ��Ph�d��>������EϨ�q�3CE�I��XM-5���O�`l�%�ۨXhs�5Mj����Ks����%!��D���CD���,�?����D�/A��R-�� ����f�K	���k�.��yn�u�_j�	t*m��2r���?瘷���`I�1Y�P�ņ�
���/�\���\���]�L��o�s6�wQ�*�;v���M�t�+��݃��J⥱֍�xce����5B�qI�R1X^XP�U¯a�;���W��I%u|����F���J�ƺӢ��2�+���IK�j��!�GH-���A�X�ꋇpAA��s�!=V,�d����������������������2���"RnΧ׮愗j盬�Ye-0�Ѵ쎺��V���y4L@'t□L~�ɭ�	��i	��<ː�b��0f��.��s���a�J�_L(�"�+�ۯ6�r���a9/_8��O0'S�@�vi+�Ϻ��c�`��G
���jʰ8��ъ_�=
�÷��}�<6�}䰍�=)% ����ipq{��u���bQg��1'�Ac�8V+	��So��%F�N_	j�� \1�sV2��l�򆘴j5�Όy��i��=�H��`r!~
�9҈�����򨪐�9����G���5����s�x#�6@v-���=*re�M��Y�3u���~9��p.�Ɣ�)�ц�5�� y /�_֎�2� }L�'�S��=uw�sʓ�|d. ;Բ�}�p]Ҵ�Ќ�!l�L��O'����E��d=���[Ꜯ�pH�Z�]��:��++'��<�'[ZS��B	�0�p �Psc�LQ�����JPv�c���� ����/<�T�\P̠��Y�%�>�'�u�.�8y�xs�1��c����X��u:�г1
�`�xW麢�z��|�]_�zT���th�ޛ��)r��׏@n��ݫnHbV:��Pb"X��|d�I)�m�����o�$b[��)��z� ����q�~ȇ�]�����8�f&�O�T��!����4g�F�伴��7Zy)��G2�ͥ\Y^.Cp��y҇�� !�b҅�<�8%ۜ����麐U�������X(��v��N_(X|��%��������R�˼�fNa�CN3���S�켞�h�� _�r�\��O�'��޴مP~$Qy���T.�(b��c?��v����b�
BJ��
?�����"@�"\^d���<+�I�KS������>ݙ6�9Ŝ���"�r����uYuBQ�R��(��{�d(�(��~yRV�m��kh�$)3�9��\yBN��YJ�ȝy�����P�N��+D�?�`~?��V<���Q:k/��p�pkUZewD�}���Y�w�~~�あ�%'���è���ط;/x�&7T��Ҏ�B	7�IТ�`���Ǡ���\+�(�Jj �^?����M�����J�c��%� I�����W{����u�h�a�Uf�0�\�@BZ�h9D�&Иk��Y�����|D�n���[�Ya��\0η<76w�/�ھ�F�K�^��՛�H�'/�ȱ�d��Yt1>���>rc�=�Z�he�A� ���zj����ŶA,�H�8#�
v|Z��2�m�Τ�`�Tyi�]�j�.�A8�ؒhQ�[w��C|/����Z�4r�8^/�����+�dzqZ�ܕ�^��R���kA4Y���_�,��CEʹmzgLv�G�39W�!g��sԣgBD~zj�PDw��2��蟅B�e/������1uIu�����o�G��+��EG��n��腵mI`�3�foo�����G��H蒵�3H胙@����=��p�FBW� 0���J�������[���m� �&2v��]ZY)�_M�>��m!ZJIu��P�iy'H����^����EU'������V�y5`D$�ּ�7�{ZuV���;�iϸK=R�ᗚ]§=��<���W�i?Yz�]�F,�)�n�w]�{!�Vk����{'a���]��P�w_h큧4'�_MEL�@�a��AJQc���,���l.$�w/��KM����if� �ͣX�#'G.�ʇi�~E�R��l>�N&��B(�j�q���'3z�K@d)�<������������x���1X8��FU��"9{Q��@$A�A����4sA���쮝ֿ�12�ܕ�Ť�'�,N��w��,D�2�c��+-�&�%`х�3VV��)D�6�^8=��r#|��1�H3=��F��&�x���q�J���2���������J��X~�P�LI��^��EH��%q<�}'�W��/-��	M�'���65ƙr>g���$���
�j?m���gf<8�Yq�&[�}9
���؁��ܖ�����!0���Wp�D)�D��ð�&�>�U�i���k�[���W%=�d�ͦE�]٤0I�a���#���\B]׿�t�=�9�U�aD��v���I#������"a&�}w��!�m;��1�/шR��Bo���^�����!q��Sb�]p��������y������3��A��NMf�n�aջ���� `Y���ʌx�W�ژ��U���T7��/UFͨ�^NR�@�1�ys�Ex(A;��9CW���m��ܿC����X\�%ZT�M���j[!��X���4���f@���� O���1y{d��� ;2�((�`���稁�F��GzQr7�Qe��R
���aD!��e"���!Ul����a9뇮7l����L��=gyPC�8�Wc�o���u�#�3�l�,��E
8?4*a�G}���`�7�3:�/m�_U�VM�^��y'����U@��|�3�u!5.��������MV�������z����DX	�c�W�8T�����[KR���8�͌!���e�fF8�4I֗
�>,���Dr,�\#��:M0�8�!����;�zGh1*�xg����5ق1P̿�$Dx�=יa�d��V��G�&�@1��z����g��?$��Ӵ�#){�=3_����%	օ�B�a�	��at�����%����8V��1���|�ch
���fYk3��F^¬+�d�^�s�m��귵���|lT_O�����=�Zy��H,��_�x���g.�k}�{I^ɔ';n���?�9�ܒ��S.��w���,�\�h�'��.ވW>|zr�Ι6��3�Y|���D�`k�s���o(�B������h�|��_SM��#��x�&�.�W��-,r��TD���4��Ƒ�ݰÇ�>!l�E׮���mr�dx�%��� 9\Tp�a�DpET0��F'eZc��[������Yb�*�k��'�n��X=F��7a2�����e�}gC	�8��(�8`^�ޱ��Ӝ�p��x�c3t�/Ģ�;��d	<�&w�� ���N�/�d=���&��m_�#
�"���.*_�{��\a'��M��´�dp���ͻ��Jl$�~Dj�@���j|S����/�����$��w�ZV2��aR�IQ���CC��5wb�td�5�\.%��7�_�uF�Qý�O��lc��DX�Ro'����^ǌ`*��uD�������ζ8NO�6 �v���Y��'���=�1̅���{ٿ>���+�C�	�Em�Z�u{���������7�[v3qYŝ���x	>�W9���폒�m��#;eG�A�9b��w]@X�9���
��#3�6���\�Z�˔)j��K$?lVP��F���=��� ��λ_T��̽�#&����v���;�t�b��;T��PH��;Χ|�A�2�2��@I^Y��ȑ�Z�jo0�i�x;�yO�[�?<>����	��X>�`p�,r�%��������.��B̄���Q����&/$�ɳqS�'�Yw�\d˳7�U�X�ȩ,{a��KJ�_gb(��Ť��[���+�%�o��9�ab��t���g��A�y���;�tݶ�:���:;$z����?�Y�c���tFւ ���ҳjϣ_��!*Y|C��
=O^�x�L{d�������b����	i�W�e 
���#�+E�i>g���!�p.k�#�KQ
;���9�ʮ5�|��k�������BHE�V�7��0�Bk;�Ψ͍$$��i�^������l#I@�T�s+��B�^�lB�?n�y�5V�������Me-P�ί#e��%�%�4{D�M~ú��"��Ml�W8^1�e�&.��Gg.R��8�g0�ԩ��,�;���z�����Ҷ��2�?�TynB��k�i��s`63hŒ���,r��iГ ��e�1Ql��Ɩ��G*5>�0�p˅�:�����-aLp�g,n5�Et�����X��?�bߛA��!d�r�V[��9�$�_M�J6CP�)�����2?���uvI^8!�
�)�d��V�� ֫����i4��&�O��V�k��["����C�e�O��ȶR��e�R~b"�����S&v1�8}�aR��c����<�_�h����Yރ�v��d� ��na�S^/gm�z�r1���b��&y�b����6-x��l~<{���);b�q�<AˊQg&k�t DU�1�.�����Y�Z�Ք�S;�?��,�Ty?��/��D���A���C�Z�0�Y�)��.�ڢyL�μ���l���A�g��A�	�62*�����~<�ߏ2ڴWp߿�~MGˬ�|�`yy����P�_v������O��;XyMU
uˁ���g�6bQC��b�k���_�u a�H�M�C��� W�;�-	A��1���ӱ��r?�B3��[��9a���6[����:8�����B������k��\��ͯ�d\��LP��,��!jq���A�B6���I��!�K�`ѫ7�����&ө��������Mxt��$m���g���Kt'��`K뤾!�C��*[Te�&�����6��΀=�x̰�g!݇ž�bR+�U�p�2�dL�X^-�>�̮�
D�_o�E!b�
������6�M��7�ŷi���o~Ǧ��S�Ĭ�y��S��1�A��x��3��̰@��i]�<��VKR9�	�U���\��c"(lm�Y耾%��B�?z[�ylb8e�Bx�{u@�ʝ�lۯ�fu^�$?�9�̯Kݢ�7]�[��02�t��G"{��
�A�r�.�'Щ��%�{����O��1o��BjX&S^��7�8%��%UM�'-{�{�����M��DH�3���H
����NɄb{{Ji�Ғ�'�Vq����J�\)����U=8H ����#=b=� �����W�R;S�G!iD�=΋2%o�r�b���	��PG��Xuk�%kG�b�]�|zk4�c�0����UKy�<�~9�knH}>����4~bx�p���_� &?�P�I�%�J�'W�FNN �O]GA`��
�����(;�y���ڪ�@d����Z�
�&!K�w��3
$�pP>��T��Ԉ�р�x���� ٬uv^�ΣEh6ӱF��pf]X��3k�8Gq�:�����?D�#w�
������p
�DD���{�5m���T���aʍ.xN�ifh$�(ܫUTTN�7���3��Zܶ��o�1u.�6^W�w�n-�
I��S�0��e����6PYs
��Z�ZU����U�������V���$����b���G�I���Q�X}�a�^n��JE�P��X7�/���Q��Bi��.���g���a՚FmGRI���?U�>��������8tO����Ġ�K���d�%��L��`����^�ى$NCx���y3ϰ)($l��ꥑUD _��u��~߳��C��+��z�@K�eC�YM��(��Z�1������ �)O�M��!)e|���T����x7!����`�T�Ͽ�rt-���0:
����E���l��l �,��'�,,�K"�������I[;2rxPY$?o�a^\JWMY;9�F+��b��	�(��{0�(�):&���T���P|k�/��'�Ϻ�0$xo@̠�o92/� �oJG�gO\�̋!�}[u�҅#��]�п�k>��[��"\E-s�>���Dm�	�B�_+$����L����� Z���x����lZi� F\S�6$���Vڵ`�6�.L&�5�PG��� �y�o�A:3M��\�Ƌ��}���1'`��:�:)��cte���3�ś��	�߁��l�.߿���#F�B
����$�T���|���S?n�o��>*��C~	s޽�b��\�[���/ҭ
��4���f&)�T$>^a=��qwSh�+�#��J��僥�2���$��.6}��V�>�4˭�����vq҉�`��e���ڰ�H�z��O�Mߝ�]8��[�D��ƻ���9q��_䎠���i�d~(�̡��V¿Ԛ�}��x�a+U[��8VV =��_6[Sc]b���)'�n�FMd�OA��Ӑ�
Al�$w��i�k�i1�P�E0P�N�Uoʨ��,��Kx'�ҥ��OF67����g�� ����G��}\�s��_�ҁ�!q'�)�y��Y��D�+��6M�[�6���2?%�s��ҧ��j�l���=>�ZU�����@BDN��sl>��Xb9d2��{i�������0�gR�-�ɿo3�Җ@K~����v������Y�:�X���rqڬ>c���V/�ۺ_4�E��v�d���'�k�tE7���>tz�k3�lA����u��
�ɩO�h�a�&
^l��d������O.�a�/��[��װ��ljC�H�j��0��*t�!��\T��5	��vp7�m������q`���b�p���`פ�y�D'�#�U��4��%��7x�;��bN5ޣH��K#�W�H�sI0� J7#�OF�QNf5ȟ{��Px{|���v��82��1�߷y �����'w��įba$y>�����#��f�)�Bi������2�מP���򯼀@��dX=��F�C�����W�g3q�$��� @�!��2g�"�8��3�2�ҝ\�����Q�Z�����+�:�Lbk ��*g������e�oңQ��+bc(�z�*0����� ?-�?�7����Q7*���=J�M�ľ�o�����1 �M����7�kE��{u���������C����&������iW��ܱY*nc��x��Y�>3'�-Y*�\q����wg�Z�5��`P A��\����xs\�W�F21"�<9wZ�K�����8��ŀ������x�a��+n��1�r?��Y�6�u8��W�,�V|�����Z�cg��˕U~�	.zk�ڊ���J�ѵ��u,�/�kZ=�.����l$ ��]�Я_C�0�}��v|E=p�
���"x��=���?�؂��
��K5*�������F��ҫ����W�@ �i��L�A(���
b����L����*iL��W]��^�$���WQF��[;�tL_�v��`VPS�<�L}`���4�HRf;T�������omV���?�8"����enu�ȏ�<�T:A�9��Ӊ=^�!��Vh�t�4�z;"� ���6��,�����D�z�;��Rc�P�. ����a�ĺ�[��9����\w=ڨ<��/U!Z|�.)��ؓ���$ð������>�H5�0^��i���foJj�O��6���Lr���������� G�՜,�\J��&��g9m���o�H�7(?
L��Ե�Yф����\T��́t�R���6�h��.oTtް�C��uƧ����8@!��<�nSo��h���l��J�6�:��~&j�z�w�9�${mODvݡu��q̥Lr^A������)[8;�9�}��׋��.��S�c��&�I)���n�k"��7?Z�h��u+���3�C�p%���|��I�Y��~=���2��&="ڨ�#��YP�\�j�h�kc����,��𻷄�V��:�>�>��n����r!��qB?�gf�h����<�9�����2��)gȷC|���ɼ���x�V�@=ŦI@!@�o����m�Ρ�1��%~*HV��Wq�SGk}~�.������<8�Y�~k�/�I����*Z��Vv���x�lL�;H6[���M��Ǘ,|r�|�������l�+$f��`Vt��F���I�1&eH����6s���{�F>r 5��  c�M��(.F���u2��6y�,�bK{�ca|��==��gL<��@���9�S��g3��N���D4��\��:�z�X烑� ��zY!1��K��V��a�U'<�Q� a+-��֢~�n,j�4V�d'Cl�=/wS�'�ܬЪ��8�Y~>�9��y�P�-I�M�'�QkX�Mm�QZ��+��50i��X�gUD�f�!�ً��E���j<w
���Ը%j{����fS����R�A+s����Q�r19���,?�z�)�-�eX�?�!CL�.� ������;�+	+�T���R��f��[TȎ�R������x�&}����&�wb������h�췵'z��/Ŕ,<�XA��^^�z��<Ah��&qG����vt�úf=�~����s�yM�1~]As���>�>�|�'ļ�Z��@���GlQ�^�o���Z���rG�
W���:���΂%��̞���V��j=slZ�.�z{R%���r����,?N��b%��@	�Tb'���a�`k���s��"�ÕJ�iB��$��Ҙs�z@%�^��7�s��c��.�E�CG�T�V3�O� ���	%7Æ'�H�qW�楲��~Ԑ'��.���Hy�	˯Ŏ���{5O��i�B�K�6���҃���l����2��sZ�x��;/\�eسz�O}=ӂ�r}�+��0뙿�u9��)
�*%m.aP���7Ȉ�B2F��r��t�|K������K�>��PQxp�;D�m�,բ<+e�$�����ƀ~�]��4�����'9��J�RK�5w6�I<�[�@B�����5NNlZ�y&�',��u	o�Zv`����R��{5��Ö������3п���lOh��<а-���	ә�x��nU��2��^[/Ѯ���w�/--�`��v��d/0;�.�c-K@f�A~Q�U�Pڊ|���F��kuF>T�	yp�V�D��Y���xL�{ض�	1�m|��>�Zt9
���l������`�'��������[=���~��CM0�w~�I0'q�M�v�:�&�py�b����>`�4l�%c5ݧ`p���@�;��/o�������v��p�UKP���h�t9Z���,}�@�����u9�_�x�g��L�r��G��Pv*3P
�����sz,Fɽ�ѢBkjF��Iɖ)K��+�Za�⩙J�s�j*���0�1��O�g����O4�m���d8F����,�q��%��m�ke;y0�q��k�1\Q��h�!S?_y7"N)�X&\�l�=�n��'9�}x3	��X�^y���)�����:�LmԨ7�b�uֺ[e>�87��S�[-������D<m8~R(={J��|�zG[e=��?�8&�B����6�۝UF����H;�R�T�T�ع����IS�Uޑ�N�&ٮ*�h$v��nr�v8B��]}ک�i�Sfi�� �G$�9j����x�Y�;�p��FSG�m'���bzM�i>>,{�fA�
𰑢�Jn�����m0*�c{o�2"���T�C�/>�L�f3=c�j����I��=0�嬭V�1<����(��A����݁f��h�����]H*]O�NY�#��,�=�� e4#�2����+��t�c-`�4�:fu�L�2Hv���Y�K�0�o����nh>4���/5X�q�K�I�:�і�G	�9(��T���_r��e5-��:��\�8E׬�n����Vb�CqB�ʢ��$���2qН��O;��O2��7<�!~�?t�K�E��X�-9y+=��:����ġ�J��G�V_�|��Ö.�U���5�NA5���c�C�ݘP��Q-�A��ţy"]4�xzi���Յ�篇��3mK�዆�o�`�^��e� �P<ڪ�~�^c��|�cUr��㯙h// ��O��Xc���0,���j�4ox>Zن�5Q��2�n�Z �ks4��t��"4i{l!��;�k������4�C�yj�EIe�F$�?d-�*�+)L�Pݍ��n.,�+H�l�H��6�ć /k9S��n�6�ĭPp]YR�p��.�L�[K� N��@9Cl���b~c�.�Jc�G���<+N���<����m��H�&P�J�L��8"�!k�݂��OdB�w�-Ap!��i���:�-�)�\�^��Y��d?=_ y4�J�	�c׷�����
�Ғ�5ҥ^&�{a����;;A,�������"�N����J1�&�N���Ӎ���xB�r
E����e�=0�5���*����L����}�?ǰo��`(c#<V�~S���>W�zv����Yi���a_���5Y�R�+�$�|�n�(��Ӆ$<�{8��V���S/f����=��;B$���f_��Jy�7�ς'��+ �*v㭲g5oѭ�ؒ�sL��dD����&6�α#՘):������EƋsuv��`��xH�e��B�I7[���7tO떉3)�M���-[m�7~����7��H��d�*���Gq�e]4dms�Hy؆cx��2o3^hΨ�U�G8;NP\�[�B�O@� �\���>s�[Kܶ��_#����qo��ǆ�ЌS�)�� .���=Y��g?P(���7����6~R���m�z�<��b(`�T���M����j
0�%0m�qov��`�����.
�^>uD�T�����v�9-��~�y�6aI�� ��?�ax�@�)Q׸d�ҋo�����Imf����|Impo�Eߢ�E��P�w�W�K5��1����qd�O���=�K�������e�6j�I��7u�S�?�4E|I��Q�f璦�T^	XrP	\�e,GH�ho:2�v�
�L�e��'+N15f�l�$ë*��?�Z�E��|D]�gzMH.�	��S<&��h[�1�ϱۭ$Ѻ�é"����;/�	+yZ
��:R2����n�{��Λ�fE47�7�kH�W����Q�?�����0��D���W��ʴ�Z
�.�"]����16�"�T��A)[w��η��BE�7%j���:&M��J.A�f�$\1��4ȭ"MХ������6��/����H;`�9�iO��p���qV�D�����=��d֠�JI(<;�8��)�WY�.��X\�%k��nyZ:7����wW��;�W}]~�w��}���<�'>}�3{��?������@np�̨����=�� ���%5����JtFy�ۥ&I�.@�Az/�+�Q:�Q@@>�,���Ej� �,�
��k �H���#niBe�'�i1s���|T��F�u�X!����<KqX��c��?�Ɔo�M0Nʗo�@n�<��'�8�S�>����~*�%盰�qY"����ɉ�n1�ƅ�6c���eb�P)�H��A@�6b5�S��qCK�L��;�/N'_�M�ٟ�T϶��'l�!�G�ىU	k���X��k{�Վ�ϴ�v�H�E��-L������cB\�A&X�_�tM�d��)��B�~�$Z�wS~��L��aҵ��Ίy����1��0/����+�0����/�J�\&�:-'��q1k���ͣ����C�3Qj(l����4���xb�?�A�H0=W�{�+�����2TQ�������HA]h4*{�G^�iP� Ͻ/���G��)���Ӭ�p%0�ںn�O])�䱳ֹ���ci�C`��]*�K
����]ԉ�e������י�kVq��]@S���d�q�:}=|t��e�=����Ma'&�0��'a,��Bv��hɠb�A������*�wΧ5*�%@3���˒�ag>֭��� 12g��qSП��x2f'R{A9̎�A��>��F�I0,UaBI�|��ǈ��4?Վdl6��n�����+ 0P�";�ܝ0x�9b���k���4��&�� ������k�ܼ������l�}�^Ɲ*<�=Mꃒ��v�/��G�fZ{Mo��
�~&?��m�udg��g��ʐN�ר�>�����br���T�o�e�8��q�8*���d9j@0���T�U�����A�Ϥ�Dy�h�n��V��uPǠ�z�.�h������$*O<q�A�v�c�}y+y��/���퍀�.O'��`�\�U�R	��T�+m�7SJ!��cյ�6)%�|��ά�Ty�f�ц� 3_�j�M��Q������2�D�L��DE/#��>��Z#t�U�TA�`W4�tκ���V��ip!h� +0�v�C�[U�)`|5})���,sU�Z������jUr]pQ"6��|��]�FZU�Aw	QNIb1d,�v�Z�}��)�I'[Վ^#��.}X�9���P!���dN������l@��{EP>��k�,��|e��q)�T���m
I��L݅���E���㈮96t�PQ�����P �$�Б���gak�a���>��b�x���w�J�^��Un�R5��_�txl��;����t��������I'���y
>@_7�Xu�>��D���~�V�
=�!��3��_v��1Or�h��c%��4��v��)$Z�܉z����L��4�t�)�(�dY���#��!����Đ��x`�̋�~�� :bL�0	�D:Ԝp>Tk�l�,	�7���bb^ȑo�Ƽ{��8%����e�x5�����Rp0ְ/�4&\I�`h�Cf~A��٪��{c�k,����}��:��y��^�[@O�����P�PL���H��ޝg�#��eAR�F�����4�D;�l�bId�vO�Ff�|�QEj���2S�8.��9�v�+C�߼T�{v��ɵ��������;��o�X ���N$cbc�zcRhs~|{���E5��$�j2������醠o�M�N ��Kམ��N-Rd�6��8kܽQ�Z�Z��>����$S�f� �P�}�!�����ֺDС\�fZ��zM���z�%!��\%�O���8��e�J��> ����ϥS ��Z�ǝ�t�[�fZ�[ x{�t�g���0k���[D�ý���,�`݇�%�$�*Kٰ��z�"x%]��+�?�S%��Ӈ�su��Ȗv{�*��?"��z����nk^E��*#5 %#��Z��<� �0,�{�ڃ��I���zo������иuw3��t�T�f��'���tȜ��a�O�kz{�=	��1:fG_4�YM��o_Ǻ�|�g�"�~�ܚ��ha-	�¨���Ru��R"�#21��i+�QA|s��J;��
������ΰy���m��ݏA��;���>i�ωY)u���U��ާC���@&�~:񹈻�Q����
\�z��#�7��b�w��4�b��\L2	�݀�]Q�8���8�E�&	X`\�"��?5�b�>�u�YG�c�9v���Ze��uɸ��pѣ�\��Ϝ����Vh��!ZG:�p^�y8�oc��N�j�(�;����x�G�#l���*5�{i��L��Mi���j��疈a���{w�e�0}�T�%X�$��7�ov0�+�ہg�(�'
��A;DTvytowxAbg�N�`�\J�n�P����ޯ�O�i�$��ɒt�"5�	�� �(S@S&C~���Φ�X���$V�Ib:���Յ����?��Q����<�l�������W�����/Z�{�� ��QPV�)�	]Z��s���02Ki���B�1�� ��툁��*���t��	~��������2�Z��:A�Ѧf�X�y�G,!�����WmM�ט���Eĥ�p��T��>ɩ�>�v�AG��	3{�o����`���y7UvDT�('�:;�#��#���v6`1,�k�g/�|-k��^4��B7��!K����@� �HPc*9/��ӓ%�Ɯ���]��t��L����e� ��n�-���������/i;���&'��/���2��!�ڕu�#��0��)����$�R°\F���V���D�P� ���8�-Bb�N���qA�I�L�5��Ҕ�|y�1/&�\���L���ke���г��XV�fK��ڽ�aVE|��d��G7�2E����׬��3�5�U%�vl�����oRY��s��f�Hf5����	��W�q��TU�'�{�w�������u�l�������ޓ#$[�U���YF+İ�~j��o�H�����+��|Vҙ��pv�X����c�� �C��9sZaHh��m�l����=��
�<⎪ϒڤ:BGɛG�O��ѽ�B%si��� >rϨZ^0����\���D�C�������O3l�$%�ǩ�eb�Xi3i��==�S���c^S��,��ì�l0����.2{�S�4]����v�I �����ݲ���\7N������ه�A�'��p����$|�s�[����7�eOl{��C(=D���
�Ud���g[:<�\��g�D���29�2=_��2Uh1����.4����W�KC}�m@S⍝o4Egϭ
��W^��k% ��x\6qX"Ķ�|W;s"Q�_VʤDkh��K�a��v��u����}ɮׂ�)�����Uf���f|t�@�3�C�tp�r�*ψ�du#}ޘ2�&�����Cc�*6���;M��Q�=9XwP �ep�ql���e�G�U����t�e�ϙ��J�C�]��
΂n֎sa���u� _U��/>��g��א+4.��S�Q�D��q�j#���e__��j���;�:�D-
Ƕu��!/��7+��6K��V�m�O�r�ހ5¾g{TYޥ�(�X�J_����dEp6���wH��Q���T,��j�f{I� �	�Ji0�&��0I_
��CK��^X���R}�G�pVM�����o�+p�F@��>�:�搁)V�zSمfu$� ���l�q(m}��	+G�;T��r<X���*Yt��54nd�O���R}�J�������
"�	���e06T���$Qx�O���gb��j��?ȋ��y��u����<��G �H=L�pB���N���)����!p�����)�s|t��N��r�-{qʆ9�ޤ�U�nv��Ƃ+�28�$5���
hY�[�oǊ�1k0#������&V�?��orlJ��s0������Q8ܯ���s}�λ�\�'X+ԅpK�7������{o��>w1E	����A����*ș * ��v�bmK���@ut}�7\H����&�j��۔HJ�
)�MĲ�uC�}�����d������ҳ���E�-Ap��k,
{���hs8����j�U��j�d�8�R��&X�c�!�,P�^#l ǹ|����܌sN��Lm�?�x5��8�^��wV�y��>� �wgreޞ���*�[9n�!G�<6�Դr�$  i#�u��pa�A}�%�B���^����ܫ�1��ԉ��ݮn��\M�% u,�2�<[`-:5�˨Ӝ��4�1��8V�p@ͯJ��M���ð��D�!"���\����2��`s#z�����&��4��$�e�4�3H�'x¥���v�#�;ԼުV�8׶�t�o�WM�����0~�Y�@��n���0��I�j��������g��h�m�L]�Z�˯<���[G���bC�K�҉&����C�{�^E|�*�4��5"�x�����u��֕B���*P�UX�Q]��Ï=^��6h3
w���D?hH��Y��� �9��a��˭@E^^��J���-���EJ��u��͝\��Q}�ð��%�~"K?G�4'���Y���(��?=�h�ņN���wI����
!ޒh���ZbX�XfF���",M΍PfR��h��0oNn�փ�s0������ߙ"��X4S) \�,��H�w
+��"ݤ 4cb� ��/o��Qx/� m	��G]��lN�ɥ���s���햒������P ]�4d��5G`� �L�3�V?�^��&q4/xuդݔU��W��s
gn����KO"8��1O��ھ!v��o����Sq�9;
�7�l��w����R�
�	`�i*��m���򌸯'�z��!d����.E�6<Ʃ5�
�������#\$q�	!/3Y����#�ڙپ7[���=8��Ul��O+?os1S��Ŵ�	��X<k+L�Q�����nb�rH��so��(� 5�W1�<�c��#�rA���A=�T��"��`��u��.����l.LT �"��maі�������8���ت�EZ7^��?L��n9����r��c['o^:wE!�כw��<�A=k�K�45%���A|��KP�ޑLc��X��HP�������<�k��ʾ�~�#S�C$�i2, ��]3ݓ�f8
�1P{9L���^��ͤthf����WZ���b�����/�{L�(�	��Z|�~ozV���hn�����fہ/`��'����2p{{~�5id���iW?��8�1�Ҽ@o�W��> ��tXJ�堎L�k/����v�.%�/��t�$�TEd��2��W�6R/����?/8�qd`
�򰈼΄���o"��'泖Y�-5��mو��G��o�ҿ����SOrR��T��{�>_���`݉�����/��@�UIՁ<�������8�Gtމ�7���_ �*���;��yS��H&ȡ�c,�.T�77@��m�$�"���}���4"Mը2���Q������T�����u��������Ɏk�B;6�̊�M3l���RI��}�9��w��T�Z�?j�I�-WD5<���T�s9�Cz�u�� �w�������9&-y�4�S�.���q���ȯp36-�Qq��{1�r6>��v�v ^��H��@k�����Oy��7���o�g��~o���|.x������hD�'w�z� �ͷ�K�j V�J�����1�ƞU0(��yM�?�͒�|�_s���/˔y�][ͼ���ZQ[���__>ݎ�=��Ճ�X�W�K����{jXnn��׭_+���MV�7hB�n�`�=��cK$۔���j��[]�iZʍH�+Ք,������՗�ͤ�s�A�2q<.o�����M���T ������kDɭ��|<�-<���V_C���H�5�Ţ�������a�<��@ 	WO����<�Z\3_�������A�l7~,�t��ň|�|�'�u��>3��Y�&�!�q�[6_OM�;�$�h5���I�W/?l��	G�e��C��e��� ��~�����q�=3��(q�t:�W�&��!#�K���q$�o1H�^G�ǋc�&�D*a%����=�`��P	|����"Ο{�.V�mg>K�4%�3;��W�7lB��U��Eb����W$�WTzp�b�|�8BGp���>W[T5aS���^��
ΰ͝��5�<�b��Vkwp�lJ���bbv�3_�51�"�w���G7"+.�e~���F��nr�F��k��`�e�� �!�'��}�����HXt��H*��u�sz���n�u��~L��>YC5�"���bR����R3���tতpP��L���>����9�pr�]$M%ۤ+�|� Iq��A��}n��rC\d�[Hl����ߚ��HEY�IfTQwf��u7��π�B������g#�`�E��i�qA7V�fC�\pRdq����
���b�u�S=ɂnA��M�+}�bIx���L\y�!�[J�N�{L�	�S�uy�1�sU��LZ���i�I���~Cx�aE��tm�l��,���xכj�wS����T�����ӣ���ێ6o��f�u��z�9���q��������x�Z��e�H�k�R�u�D��.�=j��|�ea\;{�g�έr�2�]����+;6JfĭNo�ؼ��� �~іE���E4�h�RĲ�����t��|��.lLۇ�=k�n��۞�k�!1:�:�����D��u�;`�'@�:��[�K�m�E`�f����N��2��Wj����p�3bkس��M�K�9PY��?�pb��#)��u��q�sJ�Dy��B$�����F�k#���&�Ӽ}��dx
�G*�ޘ�C��	CA4p��ӧ�I��Gy M��KQ��:2�
(���)L�E�L���G:#�6�mz`B ��E��G���7Ж<BrO�ӣ�� �
d�
���G�̝���e�E���($y�e�$�a⑤�{m9�j��f�WW6�i4�F�C�B���av��6�4��os	:��D���+5�r�}:��+>9���lFM�J�˜�7���P����p0��M�}�{ £���}�����wL�6�"%J)����?Rݑ6'���Fц�t�����;�<^��5
s&��Q��Y�3�V2�<�OU��ve��^Y���1^�D0 ��ҹ�''%��p�+���$_�5՝nW8@0�N䛎1g=�ϡ���9�}��56f�XƋ�6Q�����x��)��~"�W]�&J`؟X��&��0�Q����рf�x�Q;{0>�宍WH�pHHP��u��fD�U��O>*��^\�-01f���ibsG�v����DUr^l�hX��%C��!��VFo}xi���ب�,` (}֧�آ!���\���u}a����@�E����(o3������9:�N�1٩X�2�R *��?;m(M+��4d��-+������!P˞�۽Ƹ��b+���w��9K|���H�:5�mZ�L�q��O�y����b����	ᯪ�u$�'��J���®&�i�t�� ���ޜ�x��0�A��g���	�za[���P����*
$�6
���ˈ�.���'i��6�ē�O��4�t��s`�Zw�I\�b7��Eh0eE3�w$yiS�\���A�H�W��\hFt=dw��dȾ����O,��5m��\dX��
g�d��?�B���*��8��t@XOc����1��*y��r�!���R�7f�k��K9dہ.��B�yR�x�f��3��<��ȩ'�C�����՜\e�b����*^��2��lp�����S_o���A�m��[]c��j�-c?K"����ݵ���[��&�ڏ�r0��h���zI%��8�Ħ�L�h��;���u�fOMÔ������*�M�RS#!6�xy�a�����z��v�
iG�i�.��w�2�����pGU�F���AO���g�I��`�j����Wzʴ��a0�Pl^0�tK~l�u�Ψ�#����I��m�d�&~b���w��
R���w��:�BGČך�񠒸re8���~ �](T�s/D�����X,�%G�ᇗ���>��>/K�|$R���@��`��u�=��A��7��`��W* ��E���v��[p(z�Z��:���
,��ﺡq`�����7�����-o̻�zid�~}*���D�'�)�����M�����c/n-
:v���#F^Z�z�4�4� ��(�W�>Ę �?��P�U6�4 ����xA��K"���0��ICP�q�����4\T�_fS�@�d�>b8&>�8�������4g�ACVD
u!�ǰ�l��6�5>Um�&0r�t�q��=	�`�g�v�}!?�|p�Ꮋ�/T��� G�2U�(�R��Rβ�b�d��w���ǅwf�o_�Er���V�]Н��Y�fl��F�����7P�&��yf�+��5�H�*3��t��bA������y}Z+�Þ*E���v\fsÛ�ު��$y��J�V,2���zpKFC�i)(u	T�D�>��J�ln�|�����N{���q^�ϒ�`�\l�I:�aSy���6��'h��v��l����{�{ݶ�%��NO��>|[vw�G��J�x��з�F#,��G^,QΑ����V�Ym��.!��t?�JĹ���DAw*I��h�Ѡ����4� #�K�H�xpeU	<	�N�W�B����|m��w���\��A�����C���Wy҃�����J� ��#FBՈ_u�h�����TfmP�cjX-�4�w,�n�tm�37��b��uI�Rl����O8�azP�x��9I�.�ܭ��YN����{|O���s�-���g<�v�&��g��C���s�2gW�e���&�����ظP�x�]��Z4����펜�O%c��zi��М_ �1o��P䵌�7���X��/cl��.��+-_�o�/�z�G�¸��im��+֧��� �3Q5L"��M�<_mO種No�xR�� Y&S�����ġTD�Ce�1�:�:��qN���X6��q�/���w�v�������#���WM}�A�-2B�	NmS�S�8�}5\l/S���B�zۈI�-�le��I�|'��Pnp>����S�]��25-�i��?�~<�da��N�v5�Y�[��o��)	���u��8ًOcy��(Q��t^�8��	�9��@��Ӱv��^r��E�O�T���HP��>j���.����Aڳ�ރ`�NE/��,����|
ݳ�Ć;Й��k�O�na>�`�t6���!�g'���s~"�DR}�"�� -WMI��YD�WG[��פPEѦ�nu���Ya� JN
/�'4�z��)�'�<;y�� �����rUw���R���W���8)��G��Ǐ�#BU՞�&6:6sF��DCĚk8Z�$D�9�>�1�#��j�m+�YNl0�O�K�Y���A���~�b%L�P7�"��,����@/ۑ�WK�.��}p�y�\t�-+F��Pf�l ���<���:j&��y=3�z�8��~�<B)��H�MhDD_�ք�����ǁ?P�4��V�vXrC�u��a?��������ߋ�k.���ɂ,��f�󔌐����ѧ�s���3�?��aH��DgN�}PD��}���\�6~�H����\�?���� ��znr���涐��Ec� \8o�}a�%8��e������!�CYo�MǑVMo^
ȣ�}��M���i�3�.¸H�b�ԻxX���v��3X$��m�O��H:�8bgyt����`���ˁZ�gk�>J�<D]�s�r�lMIM!�p`�oQ.mQ�D��a���Zrz �Cv���ٿ��>�'�`����g�T��q�q�l�l
$��-eŚ�Ӊ��Q0qYEx�C`�����X��2�8�	����4��ۢ0��UpF�_)�z�8��X� �I#;���-Ɓ-���^^0U��8Ɲ�r�E�(�~�Ũ�h�P���g:�9,C�Ïr��05(�}��`�dbU�c	Z�K������a��q/B��i��������n����?�ݨ1����0�0��0�Vv���w⍼�2�䮌�W�2��grJ[����A�Ae�;�r�h���]d}UK���/x��������~���� ��-z�#[�1fq!�1�*���i�V�Eh���m�?��a��`����P�%k/�6[8@n���Ax���.�zq���'H]4Ү-c��`��dy��D�%\d؞
�3�Z�'��}jN��`Q��d#O�,�2g�l��'+� �cs���%��N�%�;�&�~�cƢ
%��O�7�z�U.B%�F�R=F��b��N�Eƥ��/��j�+�b\\<��
�g�h}t��}3�9$O�^��4@C�"X�u�q��Q������DG+�ʝC[i�B[��Eq���1��u�'��_ػ��k��2]U��8ٖE�L�9 �����ຆeD"�ޭ���Cv��K�=Gu��n��u�����KsV?���u/�R�m#|��.Ȝ���!�Η���R�(�c.`������Ñ[A9�[d�m���/M�P��@C.�F2��*V�y�8� �z�Y1�n��l� 0��|��c��k�R���0��nqM��J}�����[7��������r����$�+ؐ���l��}�je6K6̽h%�!� G��E2�0�;.�w��6<Ũ�]Y��l>]7�4V&(�N;�lN�1w��4@�yv���~Cbl��I9.��3{o��w�拊T8�3ow�?5w����:�Z�M| �ʈ���u��B1��@�\�cb�ns@���
Ʀ;Q&=dffDeLJ7�6���.��F�mE�ި�OG;J�qx���z�%����[).e.�‌¾��R`i����~s~HZ�&�X�˨ �ޫ���ʅ�u�AhA�^�O!'���Y������s,�:�	y�7�I1�����q��v"��Q8��ʦ��Tm���9dĺ�a���˙c�v��żh�֌O�-Λ������fv��9�C����68T�L�*��Ϝ���|�G�\è8��T ��Zl"$5�c�^��� m���^��$�~\(��]��z�j�i��hF�ՊB�7�θ�zC�\r|����t,��lx�ALě1�s�k3�6ۄ|����	
���o��p-H�#���K�W邨�"jЭj��[(6���hp�y�T8�)���^�!#��#��#2N�_����)Ѧ�wK���L/�� ��?)�{|��������h�%wd%�G��#��{Ё{$��a^?zCG��FHX��l��zf}�9缛<���٠��{K���d6�R��)YY�k����4���DW_�vF8W�/�.�C� ��)i|`J�)PKB���r�؀bi�P�f�8�U9�}-�@Z�o�bX�W � �S���G��ݐ:�1AR6�x��qgΰ�F4���%C׋=��Zͭ~D�%��PHAY���ip�^�q�a#���d�-Q*,�k��o�����WPnm�48�뮻�dT/%�U� �,����\a7w�=n����F���/�W�#cF��3��ҭ͸��SH��Q�e)�П�v�IE��B?����$cQ���&�,�3Ͼf�C�0-����W�c��	8�J^��[Z{���=2��D�Ϋ��Z�~|7~��=��V�R�hw���G;��ҞC�^�'6��bԐ_7�p`�H�c%g��2���Y�;:��^y�מh�F3�N�wD4Ba �Z��-�)�P3�b�Qf*`�c
��X �`�����
���JҒ\�4�#6';�e"��.�2�3Mqf!U���d)=P��Ȳ��wX�@j���������J��i���R)z�,��^�yF��+z�M4��9���*ON���}mF]�Μ�?S��}�x�t2�i�:�2���oȆ�8h���=I�<��m���M������M��1�>;�����H��g)~�i'C`:j"b�;�3PC�F$/f�a%��Oz�fH�ը{�u��C��Cv��&�C�"�-*�ȗȷ

{���@��&E�S��Ԣ#�"�����qvPZ����}d�|�zl�Є��*I����_�?�D ��m��|�/C��g�u���w��_	�е���ʀъ��w�HИN�l%툔@ӧ9�!���г��!�����sy�Z*���H_�F���H�_:�k���� cv��Ҫ�_ǸN\HC��rU�+h)�'~\��"����"����3Qh*���I�~�l�ʜ2w�5�,'�u��^?�oYW8�>i���^8�����Y�k����>��l���if
�65 �k�����{�·}p�VA��W��[G��Ck�*`��4؋(��wQa뒕�3�B��o0�i|�RT��u��b�G��Z[�d;��2��E�g�ٯ�w�RY�N1�w˨� �5	i
94ǥf�.ؐ�;L�t�~V7o��K��	�����u����[�z�h���2���ι�ɠ�����Ik����!{t5,��x�^���Wx��2y��ES��[�5�mb�m���+p�Ĩ������Ѩ����Qf�b��p���<OŨ7ÁŚ�\�C��̲��*-0�tשּׂ��'j'���Y�.�D�>}�2l#B���8��:��o|>�%MVЉ���C5��=�(r_��]Ϯ����jU��ėz\j7햪�Z�!dQL=��(Ā��2 �I�Z�C�\��8�F��r{�%�e��VA�b[����C�M4v��d?v�V:��ˉ��l|�ϳ1�RD3~��e=aɶ���i8��O��e\��.�{c����8h���f��XN��4�A��i�1<Ӄ/����rt�>h$^��j���{�q�D�#�݁�^�~�D1���{�ψ�'��T��D����@�QU+�w��A�+����.���z�� ��섛���:Z^�TD�鼳�u�	̬�"ec��+�T�j��[\�[^��X����`KƢ����߈EJˢ'l���cT ��|KS��"�8_��>ͼ�SK�b	�{)5M�d�\��	8�S�F�Z�/͇�6��.K��2���>����=�E:���� =Z� ~'�����z�QT�F��W�7Dd~0}$����J|�1�ϯ��,1�~f�~�g'~�q��N����y��<��TC�OzR���U���7�E`g��a$��f�j��is