��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$Rx�y�<��wA�*;�x���@�̦�W�X�fa�M-$u����n~�%���P�$��W��kYَ���P7�?UMfT��q�6�U��k�>����~�\N�(�����X�e���/6U|)�X2pF�]$h���d.���9E��WG��L�X"]�Ad����ľS���8od����e�GT?y	7�������ݵ�^��R�q^]�鍦�����s�ae���h��L��P_���ާ��YЭF���'\��68�b�[����w8�[X��V�F�0͘3����q諵�uW� �h�u\V�?@��_6G�_�*�G���B�絉�f������[�G��U&�����~�F��AׯK1�`c��[<��FY���4I� �#�G��x[X�=�Q1��`��R>(�w����R�O�?����7�,(�H\�#h(W�EH=�������yq��Ѿ��aF����:�U~m<|��.��0=�P/���4ǆ���T(���1�'��*�m��J��	�kUU	՚�J�
�*�;�n�U���#��+ŧ�~61zDiMq`�
�!H{�\Ӥ[�ޢLM��qW0�d��S�}��)��Ʒ��q�d��A������r�I�z]@F���?B�f�s�G�-x�D����zݥ��X$F{��}�_5�����7�7�׋�XI�6f�?�Ñc9ȥ7o���&��c�)^�do���%6�D6�Ҋ�]VG��`��.�ג�ᕍY&��	rd7Y���������ִW��)*��v�+��H�rEoeC��ڨ���m��0�8�c��ޱ���	H��G7a��Rx<�Y�}A��wO(&�����Iα���~�R�6����2΂���c=pѻĺ���[��N��� �QL����4�c	��
Bu�@�EU61��1��2N��ԅ��v,�JD\������,����T�#�PJ�)��۪�eh^�P5��L��q�R9Bo�O2�Aj��3 ���C�PJ� ғ�_�rA%���	�����ћFÙ���c�珤�?G�ǽ�$=߲?�)�:���꿏;���qx��I�(���AО��S��ġ���{�Z��a���mk�v�;�k�/��p��WB;oP�4K�}�6��Y	X���s�[d�"b������w���v��cH���6�`Ӕ�\a#ً�d0;�����7ݹ&R1Z�S��]o���K����� )����O0R�TG[^�zK$4�O\[�{��UҥT����r��c���
��)��p|:~��_���ᗡR@I.��"�qK�D=H��Rq��aZ���%h�� ��
�*�*:����i���p�S���`vN�3.e���0�1	���ʞ�F>��p�������u$�а-s�%�$jӍ�x	 Q$�v�ZBۏp��]�F�% B�.m�D �F��
���[)!/4��r�~�2P%��#T/�c���g�Ӌ,�7*�"�Cs�6��uq`�#���&}V��2��>~<��7}Q��(`������1��h��pS��1�5�*�ڸ�7M8��K�L���*8y9��.���O�T{�&��[�oR�o��2|�x(|�*�E���y��� ��juY�L,�����1Y��FrT�Iv9�-�t�U3��;�����n�I]D��V�2}6>�zK�m�A�l��"�gc#M&5�t>�;�XߏO޲�;bcqkV
x�4`��n���`n�b0%��A�9@�W�1iDRh��M)0k%� ��_/��.U��Q��[���B�lݒ����>e�+c����L��h+*�"�s�^��9Y�?����$@QA)�=b�K�e��/k��J|�B0d򉶉�+d�J���c�8��'Dy�s<�"�V=��s���&�\,}�و�Z}������Ϥ2R���Pj�����Yh!����R���xL��P&]��%�g�r�����V��Z�U����8R11��R��%�h� yL㰣}%�]�u���4$|�֝)ܦK|v�Dn�c��D��Qt�'C��{h�w�t2e��~��O.&���`�;������S�8�Sc�l1b���-i�A��L��.JoE��ȭ��
��%�m��4=,��הp�#�گ�g��V�e��u_�< yTcZ�3][k�`��L�IF��)�k��+L�t�������J�6Ns��u�R&i~g}�%��bu���[be���]K�g��m�1ؖ���H��ɺBv�+�O����j�_R|S�^T�s�� �����M�N�d�nx�N1���VY[����E� P��C�B��{�I牄+fED�"Obo�����{[n0h�B���+ӞY����z��(j.[i���_ Ev�1�?S�������(�����M-�"���:@�C7lD<�~G�^��I�ķA�HN��X�E�Գ��4�����K�|j:*a}��Qthv5��ji�>��c����0���
4]}xN�/Igo����R.AV���a�Q���@ljK5i^>�ѭ�}d&��Z���WM|kH������,r+%��1�8���C�A��w9���̈��ۡ�G�P�������T���6,��f�,s>N#��p(X������@W�I5��>#��(��=s����0���Y_Т�0?�  �ِ��"�����c�����&#�!�w�e΃]�$�'���D^-,�˫����0� ���l����5̍Lw�9/�\��/;+'@��v�("�������A��
�dBU����\�X��`V�a*^����m� HͶ��]�r�'�|$o
�����ٚҿ��i�QsR��V���� J!�p�i�^]�r1�I������O/��lK��]��)7߷S֭1�`�c+�ORb�P;Ճ;)�6��{Ւ�h'��]��5=	���e�\��9���ϧL&z�pk�L����@38�ڻ6x�9�Q3��vpc�Hr�E�._J[䧞�I	f��j��O}�.W��qUӈ�{F���`�b�8�`���3��Eށ�pB���OVռ��"W�U��H)��u�C#V)�p�~�Oѻ2�>�T�ǣ�����vϜ>�>�  {�K��(�7g�C��nR�l���u�'�)�\�ڌ�1��+��u�<Y�dt�ѥ�+m[�i��"����@�T�҆�z��tn>)������UL��O���|����A�X����B���VI�4Թ�w+�����X��;h�|�������;�\���u�� a6�(/X) )�Cl?a����lխm���E��mL����4�{��:�䖊	ͦqo�Wı�%��:��&��l�̄�u��o4Y�9�w#g1v���y"�X@�
�����z�+#��~�B��ދ���ֿ�h�O��LD1o^��dv�BQ�}ޓd����I���T^��>_bd��	���ê��mעU�{��:�c�(�;T����%�AN0;�۠b�<<wqzT7o�O���,��ti�G��;i��o��6��Ǎ}��.�Eբ�f��	l�SR�ck�J�ֱ�ZbU�U��k3b�F�2��rd�\����U�*����-�?�%PsA�&�!\N�<d�4᥅�5�NGg��A�i���O  �!)w�s���*�?/$���������{�7����AŦ�v��P�3_��jZ�s}g�׶w�{P�2�3�h~ i��RH�6�m����n������ '�O��2�?Ln��5�f����rnM�ٌzV'�)��\���wѢH�i��_S�sw�qV�7�e���Lo���1������lc��:�Y�� ˦��{��	�r��:���x�yi���^�7�o��ߥ����{_O����/j�Z�gCzpq3`y En�M/Q�l9���|�:a�^��V�#o=��w)XV���t�c?��1D!��kN�����rK�H�N��SH�!��
��0_�=�g�_�3��g�� �_��C�u��)����.��o\uAf���?<�~a���Bt@���]klX5�`,��ql-�'U@4o&�H4E�Rl�A��T<�� %~�&F�$�N�������d��9]xr�wi�d�bV
�H&o[^�?�e���(�K�\�V�u-8}Ř��*ǋ��4���%��G��>�z��[�4���&]�̉hQx-�7����^�M ͂��T#Ո(�{dhW�k�����B��Z��s����t����#w��%�)���S�K����K�uX�;�4tmoׯAn��M4�����!Eq� ���~�ڣ_��@�yv
<%z��B'(���F b�_�hp�
��^kl�B�c<�����o��a�?~��t�F�{�T�Ja�V���>W_a�V�C4O�:���"֎ߟ�J�!��Fj!�w��k���\̎o�`a.չD��O!ḅ`��:`�Ʊ�S��"cA'֘g=�ѥ]��3>p>D�R��S�X�C"ٶY|:�/8@�.b�ϵ=lB=�eaD��ɝ��rK{��ů������`��K;��,Wd8�T%��Ou�X׾$?ň�=���_t5��������+:�h�|�u�߽�~����3���W :�dlc�-�m�X�%u���~�, ��fҚSp.��c�	lJ��<�H7�4�z�%I�~��yO�4#u�dk�:H�����]�0ARk������b�-\Xc�>Z^�&�P�ٜ�u�{�<�Τ�H�k�������=�ntI�K?n��A�[�+n��=K ����+ج��D�+ȴj���7'ᄻ*��X��"�6��+�}��c��)�rh�A~�.}C����p�Q�<�'����>an�`���8�����B�H��}�R�t"��]���5�p~Xb�s:�o-�!rF���s��0��DF��K~���i�T怼u�Bu�\���*�*KL�=�j[���/;������6?U����G�ʎ��d�J���TۻQg�a����k�/���r	(_�ʊ�H{H��!B3�ؒ����c��ɏ&�N����/T��V��+8�$���i(Y�b��.@��p}�k�����=ϼtt§KБ+g-��
;>��/J��{��9�ҫɉ^x`t�Q�b��� �(1�lߥ�H6�z��y��q:i��Y�s
��)�܉����h!�L�v�p���̪k3��jwqƟ��3�)�&%�M������t���Ĕq�������!/x]���(�����s�hɓ!���Ģ';8qC����No~.�P9�&44&�ag�q��R���)ë%�~��H�
H񊪤��Q��ϒнRj����L�yB'EUYFt�TV[^Xz*EZ���=�:I܂!GxY�2u�:	���x�z �M~&p��R���7��@n1-�*����ؐm�%�oa*9�,����c7�| uwHMҖ���J�֊o]�|�;�	Y�JZ�Iw�=N`6�������z�k�m�p�s)����K%\,�d�މQ֯y�bL#�e�*�̟T�YȠp���~&��g�ͥch
%r�0>���D�b�r$�8�`��F�2G!R�~9����`�ɦY�c�����S�}�N
�*��Q5��9��:�ag��5�^h1.!y?p��XT�];�0�ug�&Fj8wdj	�j���Z�p��� %�5|S��ǺfȿBg����$��H��T`0��1�H^rC#a@�+�t�!!ٛ��c�-,=���f�2������%"�m����E�b����dIs�)��jCT��KT^bg��(լu:�f�]�$��i����25�:�m�s� Lߞ��.���0 1ǽ�z�������
��7�.������e �z3%eǰv+@BI۾~��c�fU���"s7�hSc��1ޗZ�Vi�L�EO9vAp�g��a�����	^���)_Y�w�����@��1�/f*��hv>�CV$�B̅3��dx�b�4����b����j]�PMb�M�e��R���hE."���D������'��B��0r�3�"�����(�0�1yą��D\�\_�Ͻ"��e��q��W���x��Ú؏��DuUwH����|R���'��yք@J!?A6/m��9l�T�d�4��C6�>,U�*�?��	���V����ٞԚ�����h�\1���{p>��skD��"��B^M�-��#/�/&�hd�K�|�L��Q��}�8J�㤱�}��7M�t��&Ѕf�s�t�ޑ�)����J�Xh9���K�j���X7=���๴�
�������x{_�u��al�P5'*1�7�N
#i�3�pW�m��A�oC�s�؇Ц�,P�g�P���%%zTp<���-wI�uN �G��&�y�e�o]Y}���6� .E����������AO��&�?�DM����J��'w�A])e��2���l�*deP�����_lV��"UO�qaʰ8�R�� ��	"߀B�*�@���+�+��Ij�������ː(.�B<�B�r�RʙJwE�a��5��:�S���@OfaH]k��	ȑ�i쒞�Py��ͧ����;�3������^���}��!A!�	�#1�F�| |g��q`�5q''�����!^yB��1g��+ź���n V��o���T�J��`d���OC)�@	������$o��V��R�K���;@��h^�\GjEh^�vNTO�Y$� ^'�ϒP*}�]S�]�b ��I&��,)�.�iM*�s��I]`�̰�)����x��W��t��m��q��e?���B$;\�����odKS���`�P�)�Q�7d�*j��-��G���h�Y�-��`���@��W�W����?�L��#�<#F�q���� ���T�,�¥�F>�j'��n�G��7T��u�ZlcD�k��Nh\�ct�*���.r������*F�XoQ*"�Ǔ��	U̱�٠�b5���~,!�]��,��_��J�J����]QM똴�D�5���y\�h������**9\З�g؇�K��e_����xF!3���y���e˰���2�ub���g���p�^�Q��	BJ����S�D0*Ya%�4�9|3�F����\my�a�+,�������r�n�K���Ozy3�ѿ|�-�__Ye9C�w>:�ɰ��yQvǴ�D���[(w��z�^��10R��k�������h���x�֗$f0�oR�c���!߳5k1����-7�)���%r��B^��H+ej>�iBQYɤ�EI�Q|�~_k@�T���Y&���X?\
)���<)�1�Դ��/߇�E�"�\���Nݸ\u��w�"��bѹ���?&���+��Mc���W)�٤����|�p��.�(͢1�@`��M�.��՛pkv3h��-�b���.��h��41��rM�`Xu���Ӭ9SNB�K ���>w6
�m��~G|�ld���X�X=����I��=��%��W��T���Ќ�&^�3 ?����D6����]��Qw�mt��*�TSْfU���# ���um=��Rh�W��;�'.|S�q�ٟ1.hx���Q"��+��Jo��/��_�d��y�����,����s �]$x���A5ʥ���ym�"�n� �i�RVL��Y�Ica;:9!�e/���3��%	ѷm��S��gL��a�	����6�V"�F�u4vx����bK��f��+�h��T�g��<����
E�p�.����d�P8���|�S�O!-O_i9��hxpD�9fr��p��=�D�OL�L�Y�S����Pf�!�/����\8X��噯��*�o��$��=��n}%.)+�a�\caT�9d��i|X�S%U�\��dG�,O
I��,����/I��5>�\(3��ΜЍ�-:D��b�����q��\X'<�8�u�C�CĤ�5�� ^��KȐ�V��D��z�0�r�W����Tt�!D�a�8{��2�GӖ�V�B"9��D�nk}��`�mL���^3��?~�)�%�Y��逆��^�oև�x���1m�D�걊*}�`�cCZ���.U��-3�ɦUt���!IbԌ�ީξ����Ȅ��^�cRR�[�]W��{őo\���0i&s_�C]�8�-ܤ���R?��R�Y��p�%�@��;©�����ŋQ����Y�#{���	����ƽ������o3���J�6���Zv��hz�#�QB�i�w��[b�K80'	L؋;���,��6�%��_-�d���,��[J5 �B��z��dI�c�I����G��XB�r����tufQ��a}�ˮ�r�z��ATc��9ٚn�tv��y-��s����W�m^�r������^���s�5�����#�X� S�K�[�0|�5(���{f�6b��%���HQ��J���{ܺ0]F�Q}�$���fR=��f�hXh~���{�	�����<�;�&f[D��3z���@��b�T�>}u�-O�XM�mK=�$������VP���!>��{/�'���cn���s��;~��r���`^]H���.{/�i����gkƳ�E������RhSX�I��汙�8�=��si�f;s<�	M��O.󶬻ax4�r�|Z�.\ڠ ���B@O'�?�Z&�g�<,d֑$4�=� fkm�yz̨�H��.��J��S&�����XۜF> �Nf�~e9��B��d Ο����D��?��
��8�'�$�0�Sp��<��q�:o'��.�v�*�u���Е�U��f�b�I̱���<!�7%}�~j�t	�L��2dk_��4ev�2�4vd�!�6�ID4���pV�Y0�1
g��U��)�M_7�Xe	�<��֨s%aR��%��K%O���TydK�E]���;���>�u���ʩ��x�~x�M�g:kf��,%ѽBRM.�ߪY�= pz痎�Bo��\`�5��"H$���/MF]�pɗ����:l�@��H��R�ZX�4�>��}%�\&cX�n�F�!E�ߞ�w�zp��M��V�lj{���Q��K-�^y��6IN]َ�N;��ʹ�eҕ2��wx88���J>���^{1Q�^�F��O뗿jw�*fq�����!*I��o���T.�Ξl�5�P+�N����DN)t׽1.Բ�XV+�Ȍ���&
�H�Ў3*x-�o<`x��B2P0�p;��B����#o#��5[}���ر�YEԹ���u�ϛ�ѣ�{�6ycj��#�l�pR,��"����Mk*5�ԑ��0s'w��/�gl����Ld�z>���E�y]�T#��v�+Wr�_�l���	$!>:W�@Z�t;X���P��<��U�u�w����nJ�D�3��$я}���C���^�(m�$D0<+ޑW�������������[2z��9�_6$�]��6E�9͋�Xm�f<����?
�,,���;4aKp����8�<|e��\�(�Z\����E燦�]���-
/�l� 5�᜘k�#�NG�u`��x�l������#�d��;G�B`�Z\��Fq�47[�Z�K+�974���b"=w����(K<pބ���F~ 
��ƃ��'	H����C�C6BC	(ZCaո��6�z>�i����2�
[�ՒS%�!&�*
T��F�Υ�V���N���k�kQ���F��7 <�;��r�<"Yy��HBGo��$�ˠ~U�I	8}\9r�"7�@:�ټ�Ђ�T�\A\?���% Z~�_ޕ@��q��j��s9�� �e��IJ;�`%��O3
cO�d�VcQ袤5�8O�lo>��î�+w,}��ʡF�ߎ��}Gj�A��{�U(�ed��<{�ܙAt���no�Sk��3>�^�>m��zp��j�sz'���'�n�X�V1Rn��	��w=O���M�fu�5s�B@�FZ��w����̗~�������Y�S�Ü#!p�к7y���]�-/z�<��=��=ic:�΍dF���ӌ�z�t	UB�{�w�kΩ��\��^*�'8&-�V��H|�_%������"xc\�����^�5y�x�w�G���#�Ya�[�-@�,2�<�}���Cا���ؐ��`n�s]!)p�'�QG�0�i&Dk�����C`�h"�!��Hl�J��NA�S�tܚ��ͨi�a�a����N��z���O'�Ɏ���`���m��@TQyD4��m�T$�_��c�0��^a�T�Ev$>C��wү7���xt��T	|��Y����k���h�[�m:uq1�vF=?C����VFx\��i�w�"8M5"���;��M~�a��'af�@:�Āϑ�t+��fxiYo8P��|{�;��w�-l�V�����I�EJ�����|<%�cQz.���;�<�&`ՋǱR P�>�S�������x���S��F�Z��e咳��H@�W������T��v��3�8B�?OH_�H^Ӝ�eAX�$�vؖ�I�](��q�a(V�+[+t��ׄEPS&��A�	�sH3�^�H�l`���_�X<槪�l�Lw; d�Y���(U����p����~Q]�c��2�ǋ���Y�Np�Н���E|5m)z{O1/{��k�U��G�|��'/��s�D�tA����]ӭ��W���>�H�#k3J�������	7v���G.���T�<���Y�@�?�����x��%��i3Eoכ��ma����w1c��=����)���٤խ��Z:�����kqʰ"t؄����ͪ�ٴ]m�k��ޜ���˨z�Od��Nh*���J{h��,P�j���~��:B=��-��5j�&������~3HB	mOQ��>�ǣQ�-.��
�@B��E_���7;������:�� �A#����Y�l8i�)+2YVʮ�Q\�h�R�
�'��ƵΖ<"�9�/n1����=i^�]F���KX7E�h�l,SWO�tbl��2��?eE��Z���t��V:_֕�T������%09��Y�3���5+U��տ�T����_��lQ�2�=�IG%_��5ok����)��qz�'=>�~�d�K܁�L���Oʲ�h�+��@�Qf$�L���]*��u�*L����u�n:[�"�WX�w�m��0�J�-e�
�K�.�A`�� [�=8PS{����m���͚��Ndz:�EV�]�!x�E���/g��
��iy
�G\h����#e�~������UML���)>�&p��N��K�1���v����������v����e��%���X�d^w�7���m�ա> ��&y]��$�t"|W,R���Q��=8�O!;1;8?�Tt<�fӇc���Q\�����6瘷������;�?������k�cmOr�fL�喔�RE
�v?�x����6�r)�Y���q%}HҢu' uq�Ɯ��@�i�h��&�� �$ �Xiq6���L���:n&JL[ʔ��C�*�ۯ|�N��Ȃ���Mȓ9�L��e�0	���P� =��|=^��. ��xF�޼�Q;�E���x����2�����7����}k���o���l��	�y7���(�Op��G Bn�IW���^E����Q]�X���J�VB�]G�]�����j ���p,�������ߌ����w X���bz�����A��OHK����a2�+���4h�p�V�3��TYdpno�q�r׷�-��1[+��G�&�8?��>♭�����S�n�vg�0�����A�� �s���� ��Lx�ϗ����絶Q�8©4=�-�}N����(���Df -��/�!�y�@����C��S��Ů�Y>Ԇ@�M����m��_���F.�8�� �
Z6�g�}����A�J71�@�r0�ث�	� 2�����z��_����_6qc4@9���_�i�L�54�4��x�]ץ&��n�qo.�I�Ѓ�z���
�~9��J�Lm�4	�H�ɰ��H0����c�)�������F�J