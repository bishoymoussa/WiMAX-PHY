��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$Rx�y�<��wA�*;�x���@�̦�W�X�fa�M-$u����n~�%���P�$��W��kYَ���P7�?UMfT��q�6�U��k�>����~�\N�(�����X�e���/6U|)�X2pF�]$h���d.���9E��WG��L�X"]�Ad����ľS���8od����e�GT?y	7�������ݵ�^��R�q^]�鍦�����s�ae���h��L��P_���ާ��YЭF���'\��68�b�[����w8�[X��V�F�0͘3����q諵�uW� �h�u\V�?@��_6G�_�*�G���B�絉�f������[�G��U&�����~�F��AׯK1�`c��[<��FY���4I� �#�G��x[X�=�Q1��`��R>(�w����R�O�?����7�,(�H\�#h(W�EH=�������yq��Ѿ��aF����:�U~m<|��.��0=�P/���4ǆ���T(��垝B�� ]O�������x���f����U%�twcI � 5�>K��%b��dd���|b0��N��e���J�b�j����i/�zثy���9Q#tR C�?�M���P�M���ҐK�Y;{�
0-���5j ���햹��Q�n5�N�^�WA>���1��&|S3L��C�W�;��8���b��Θ�\9��k��B`��kޖ~Z�k�Yqj�#'N�� 
��Zuܠ�����:�-���j�;��ܰ���^�sl�ݵע��uʲ��Ǻ|��7�i"�Z&����Э��γ�t\ݱH0�yܗn6�����5�,/@��e:��F~��D�z�A˚A|a9���Ӛ�+m�*i�#�2�z=�/M{���>�b�j����v���71i�t���(D#Q<)�f_�8���)x:�?%&�o�2�i,��~#������%��ƕ���C���mF�e�d��87�� �+���&����~��s���n�пF����	 KԏEb�]���u����9���_7�.��_XG��+˞�D�.P%hܩ]��#3�M��@{>�_ON�	���'g%Ae��{u^}x��(pG?�!-&�Ll)5�y��D_e����?�!�<� ��3@`��C]I�7";効Z�a�?��azo���d���4OD�7�f���a��J���Y��ƌ�[����fQ_Ր�Qag�c�~I�U0��\�Y�d�p���v��q�i*G��� Tk�6� [�CT��%��J����}B�)�� j��6���.�0�C-��L���t ��)ͳ��5�w�����c����;X�e0��v!)��Y����D��k��z�ϑ�����Ǡ{����jՃ-� ������
�S��#� ���Kٸ�n��N5���˴ǐ�'�x��U�����4��M^B�����4�����;��s�*1Z����ݍ����-�K�dMX\p�Nxntvَ�ɻ���[�W+�A:<�27�>�sӐ�ߠ�6�{��qn��56S���m%v�Ԟ׸�����.�7���boG�C���,��p���0�"s�hӭ5����༭�sQT�C"���)�SN��ؙ�e�zo�z�7}�o��VҞ�^�q�@�=~��{'ڬ��ol��?�q�H�
F��ŴiJ�x��w��ń����v�Ů��d�*�6�倰`�	:'G�md N�k$�k-��kp��]Ð�C�2^@Q���m��y��.L﷢��$�z���ʓX�'i��a���о��9	"�H���x�(:�qf��`��xJYU�GkE���ނ� �!����%E�F�F��x}Q�o��垂��qr��"��>E��@�V&p�6�`H�'�2v*4��[Ϻ4��ϸ�������;��M������i��֢�Q�IyE�91��TP��y��O�|��J���cU�h��_4Z�M(�~�v��'{r. �,/
��99���y1���_�Pn�e����K�_d&������5aj��I���^�rOxP�aC��_�h�����!?!=������'xoap"��7��i�|��M�����]s^H�y.�z�:�Y@"�o�v��]n{�9�䷸�5��=ކGuϺ���q>�hg���#���?@c�GI��}�ZZ�hn�3�S�m1/r)J�"<Ɓ�)0��E5F��Q�<����QGi�sGŠʆ�d�y�UY�}<pw�P�D??l��k���G��v=�k��+��X{�.s�o��0��)�湽��ӧT�}�:x�$�볅��xQ$�x~���oa4�pCG!L,�� (?9uܵ��ۄb���Mo�q����F�4�jRm0k(P>B�s���q�)Wmc����!��&��>�|�'k�*���<�b�������E���:�@H��|��ͨ�M�8���y<�J�Z�F���:̥�=ß�+��m&m5$�c�B����77kgq��9��?��˥"e,����	Ѷ��1��˰�T^gg-%!��:U +[��^�#�����+�e�5&� ��D:]��9�i�C��C��s��q�D�:쮝�s`}��͋�u���K?n�9���vn�#���A���_iW��9P���
��%��i2e����S�Ia���s����m��kղ��|�eJ�kl}h:	b�������<�:^��(�[�g��M� dE�w��u�.F?�r�&Yoa	�[H����:J���/Z)�o|����DC��ܮ�l&:?U+�f����kOh�=[�(�je�,<Ǩ�!15|�Uo�F�FSj{!y�����ё���⡲T����P��O_G�H
^"�~*�]�{��e�yM���h�͕�x�F8��K�N[��%�M�o*G�J~*���S��Ѧ��ˎ.{��c�������KT�^����f�%|�"�T~�M^;�,�k�ѭ�^�9O�&�� �� ��:ŶCN�Q��/Ӓ�+t[@L8��@H+���J��cT�c�Ķ�W�x�ڵ,s9'{Q�������LsZb�h^�$�m��J�8Ww����J2Ę��Ҏ���9�eR�N��=���8#��6Qp��8���+�w���P�B��:5hԃ�5W�T�p�G� �_|(�|�0ZЦ:!D������*��#n�!�<�񝬘���Ɩ�A��7I컶��l4�4�����I��f?�q�93��W�-�M�l�2n�����`�8W3}��@�z{�R2�D�嶛8�?�aVl�O.>k�(ҁ�F�G^_��7�BͼI`*2ׁ��o8Eq6�ۮ�~(-�=�F8��μ�`h1T6���/7���۹���o �� �j���
�xodF	ü�N�����$�Z4d���
g?S�,�3n�H�v��n~���������:|D[Xt ���~4�!��/]��;�5�ڬ\�R6�D.?K���Ph�8�/��J�C^�9{O�:>�=m7��C2�P�F�ހm��Sm��B�r0�-{I!�!��!Κ�-�S���|�H�R����Mg�v��ac����dbU��X��(�t�6��:ۍ L���R��M�?����Z�nʜ�O��:04sJ#��wm��`�|������f������i�p���C����H�?��pgW�����;<|t&�{J� �O�"ˇ-<�]�|Ѹ�B��I�G����LbK���RN鞲&�;#�[<o%Q,�
�5�hl��]��m�0$H]�����R�޵ζ"]R�aGH߽Ǽ����D7��	����X�������}�9?�gy�!I���p^EBWu�iߡ'Y/?��>_/p�Ut�c��yb2�O��h�2&�P2�R|j�m�U
�B��7U:��\�Q�,��g���OYL�����X�$����B���b�@�䉿5��0~��Q	�+��F&�Ԙfqz7�#���q7�d|�uG��CF�2t��|5��7^m{R{�R�ʷ
�<}զ�ٔ���hNюi�h����:j�q�M�l���+8��}����<�v�Y
;U��@"�Ҽ&s�+��2�@�����KF�Ї����p����'��І�o(��o �9�Ls<��NJ�"T8�='Kj1��&R�� ݠ�eC|�;V8S��s�������\�[t|(x�+�l�n�9S�����4�V�t���b�N���)T�\�C�����R�I̻ ?���;�G�0�
�L��f.`k�{c�E[R|e5�Aq�Y,�ͬ-�B\��;���Fr�ݒ�>���f[����	����������� �n|�P��0nڶ/�pO����M�'yznu�%��2�튧�].�ܦ�?�}xQhjӷj�i�N=��Hz�f�;˱���q����N<^����ز�@�F-`^xq41�[��;��tf v��[1^G�����(�"@1Ԕ���z�~����c���=�g&�PZ���{�����N��3N{��~	�~��p_�r@��IwU��vX0����!Z+�t����pI���5�	����5����^؟petN[$O��bg�n��|+�����r��D�Nq)b��`*=�)��H�si��4t�It����Z�B��P��{^���s>J/�{y�#��i�C-���Eq���"k���5G\�ܺ���╄�(,���c�"�GH��Q�/8�]uF�K�d(sFE��q���Α��M�����[�p�v�m����'�!�t��~m	kT��Y`�:��_
���`�oROkd�%m���>7"�Հ9/"�p�9m��!`��4 CNB=}�~���%�ꖨw�	�>6�,����ke�W�X����7)�+)��E�պzC��\Û����H}*�aR�4��I&��)�,3��
y[ 0H*���I\���$����L���-���^��s�>�K5�H�x���8��QN}���E�os]����X:�L9� A������ݚ.�tC���#�
/��z<Ֆ�"�j[,���5 �T/��X"�@t��(��F�W(p�{��b9�}~	�uiTV�Ԋ�=JM�]����?��}��h�+ )�g��S�j��+ �V�>��L�_S�������T/��-y�m�B����˲�[#~O�e�no�Q���I��������zϠK��BtQ�������/��.j�Sa6١�4�=bB�`�R����B�\��E2��P�$D�Lw�4���-�4��7b,�.�@j�n�&MMj]�y���=���A�zw�vw�%	�wE�P`R7�CQ[�"6���c����\����~SCѽ�j�^O��M:���bL��1�2�Q��82ۼ�_����ciJ�żݷA�U?��Ƣ�~e������R��"'��aG��q ��!���A���~h<�i��!�(���#A6ޮ������^Sqρ�(c�A"=8�l��#�$��n���,�M�}4*��^�)@"5'�`r�B��_=�:��F��]��D�?��n�kb�k3�ƎD}��ЧR��ȳ�Z#�:���O�ԕY��C
d�XD�cz��!�aL�	��99�o?�z@������n�D�3"2��!^B�Ԥ��s����-�䙃S
�-.�����h%�V��𠖯��U]�ӊ-� v�ہ}LQH�4k��Ճ�5�D��$/ A�����j����K��z��L >��cO�<Ȫ��9�660�5ME|!��!D�G��&�j	��Zp�a��0~��s��@�.Ͷ?7��p��p�z�m�G�W+
�o��s�,����Lڇ^d��9MB�Y$������1z[�'�twi�`
�D1KC����0��e�F��C0͜�ȋ���O;yp�&T���Ln��[�KeC�=�<ޝ�;����]�/�t�1��j���m�M=	%L��Y�p$����CV��3or���݅o�騥&�V:��b����l6�d4�>��n��7��,!o���n��z�Xg������&�HÊ��ps��&9��-��
�2� �>�Tp�!_��b7.����d{�gte�H3C��Z+3����x3;D|�E�4�~�<�PP�>��%Bt���T�8���¨N���
�<�a	ı��O�(ާ���B�g�:r���ҁo+��&��ĚȮ��s��Q�u��2� ��3]�|�|���Q��=�B]����G�3�`�\"�� ,�1V�^��%�iD�k�h����8j2"�@�A�L�j��^z=Թ���?=b��؟�1���Xy6���D��N�WfW3u[�+��k�K~I�+3\�	��_�Sgh�Q�H�g�MF��i�@>�&���.[����D�����&<V�Yg�ˎ��!B��梃�*�F�7K;+R��j̸5k� C���0L}��7�TI�	X�ܢZG~�����VΟ1����:6+��_ȼ��xDߢ��u����<��0���v�I��Q>�:J4�v{�O	���a�No�����5K�n��Gz~�r'p��J���-
��U��ϣ��7/q���L��5�����LZ�F���z�Ֆ�I�s�G���*mX�>q�ϻ�AS�'�쐇��{�����3������Xw��	v�O�#Q04�#�C�|π���U�3��/���t�hN���~��;O^�6�q/^�H��C�/h"Q�^i	��*Z�G�b�#� �@iI'<�2r�)��tÜ�>��SQ-�Y�$,h˖8��X@�秛F*phx�=���� z|n�O��S�����@ao�i�h��� ���$E[ioN�@�̷5��!�Y�a��$�ES�&#2���?�(�m�\���̫J]����&�_���z��K6��Ȯ ��P֌�wCj���]Y��k�N!�-=1m�B�s
�jSP�D͛��^�d_��Q,�&�{������#H�'�����m���+�)c���@�����r�84�`��~�-�0P�P⁂��O�X�PM�w�B�O�B��z��<��+��Ӈ,����!}��e�Qq煰�����),���P��R��LW��Y�Cl��T�0B��c:���_?L��p7��`�*�}z�_$V_���L�����򁇬��]*>�}:b�E�`Q.����v�0*�]�U��-��� X4��Z�\��UWAX���G�%9�� \��$���^�\s�����W����-�%t����K�_#���a�)F9��;�C�mOr�����<nXh\�U�qf�y�3�sځ4I���ń�-�6 �C�V�ih������]���9�xL���x]Mg�|g���^��v��U����N�8��xS�Se�.�e<�,��7%��Y�ջʸ����T7,�ɻ�al�̔�1Y��R#��G�H��-�S��uRo��&��I��,��N7�eǌ<%��ݔҚ�x�������n�܎���:1�T��"}TbY��V|���P�4^�>�l��e�����dڏ���H2E���R�v�1��D��5�)�2�
/��)�J��s(6)\����yƼ\ޏ�_Y3�u�N�6�3詯�~�#/���*w^�V�Ŏ8O�/bnE3J�3� {�h��g��ń^A賱YR\9�vj�r.�DqvfRv���F���V!�je?	_����w=�����	��ZJ?]A��]�V��\<fe8he-���I�}�L��mWӤ<����Ͻ�IܸHfΨ��&_VM��ȳ^�ݻX6�a�g9�/=�V�����=�n��_���_ȳ7`lwl��⻨25�?,gT�f+��B�:��e��J�=vLE��.Ȁ�o��ېHM��Wnm�d��(���9Z�>X��X�j���뭺�҈KU�P����h,���C�x��p�һ���#n�"�@�7�l��{x�
y��u<o�?����u '�;Q��(K�A�9�r�V|q�?;2ބ6ؤ�Fڲ�^軜����E�+Þ��5��3�� $����sW���0��h�-s%.��d�`U�3��ьo;Iy���Ɩ�}jd�9����b�F#*f��g��+b�)�����ӝ	5h�� ���?C0�����1C�3brXl��a���6
&�uq{�iB9�>p�N|�O��9�P��r_�3]�,�����UЏf1���KY��h�a���R��]�Ej���� �bR��D��Vg+�ʸ�H0��~��R��~�e�� �&sZ��6��{�UXa����):�������1�`��ooF�r�
��j�W��v��4FI�2���;�E��@G{�^#�
�Y>�E�/���nw�c�N�|y;�=V��L�m���a���=Ep:($& �ՙ��kR4�\�3q�/鮁S�Ve-�W���"����t��inEX��<��{p�}ŏj�6�<��R՗�����L(�KM�i5��PO��W��μ=�e����	�e���Wm-9TD��H���h{Zw�� Bo�����B
dnUٜ�Ttw�3��M��mn���	�P���L`e;�����E��V-��/V(�R�:l�s����.�H1&W�B<��*D5���C��*��v/r����m�~�.QN=]S�0�$���>),1H㋏����#�k;�)�H;e���P�S�$8�l�-;]w��� p>e��W��A�V����Y���Ӑ%�p��7TXQ*pE6��=���4������2�����L���IQj%�G��ո1��a͐������D�{`�z��$�M�|�*Cv���8�:��>U׻JyZW�E��O���w���2�p4�)^*�rM�5�n�(}��E��?;���{;�\Z�9�:�,��3_�ު<F��}�(y��j�̗��M���r�O���)�	��g�B��t�C���
�����p�pf0У�OWF��0��w�pH�0�R�~?<CQ��8��5�� b��8)>t'CF������٘�f����/!z�{�d�j�W�ո���@�.x�{$�)�r��0��s�!bH<-�-hP��Bh�:�5Ly���_
U�=Z���7'Ћ�f,�m���J�	p3�㿱fUjɋk�Vx2�ʴw�r4H�:�>M�7�MX�m�	�G@��g.G�~����@e���ۿ��xЌ ɟ�<z�g��'1�	�-C�X��E�A��0�:�����_i'<\}�瞄≱��5��d���j�C7v�Eg��ľ]+ ��EW~�y����=�wt��،���� d��)V�_%�R���l�����5Kg��Lj֢d:�ijS�6�͋��6>�������D�*�|h!b??�g�W�� ?r`&�m|ù5�5Ρr������*/���8���E�	*��z��{�7t��yƷ���S���*(�
m$C������)0��	���$��F�shb7���0$v(LP.AR	@��N�W�v�3�E���f�����*���t�iuhM�R�<�U�