-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
dkbfVp/K7QjrolNwhEYgEP9/PUVxiCKcAKw+BMY9E+i9mU2yw60DsSFQkuWX1TsYqPMwvkDjdO/f
6WCRQkbqunP021A480gcHhC3p4mN+BarKNqx6OEOnMix53w5F2sTUK+78/hmZdPZ1A01tt4kBeBL
i902PCIlPFiFIRSN6pq/PDxPl1rg9Rrzyl5RrRKLjg+VLWoZEVX1QS8/sTIkxR3HyCLsYjq9qAYe
p4PjlMSiYhymk7ksfozxDpeAsvIWYiAT0KS9d5ez+GHOLTfN8JvZovHpZjLtV0NDjP5LpHiyX+PV
CNBLO6MC3NQr2rRYWUSNvcUKps8Jg1/JKIJn8g==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 7520)
`protect data_block
l/YFOZQYMEUcAXuwGvh6pr9bjJLbr7FZpPKQgwYRXZEYg2sBD6wBk/zJZY5PyjNc2XE0t0om08Ng
XiPPqz+oD4yOpgFsUtyd2b45FwOU21JFWlaove8oop3WtM9sYTg5oNDzidaKAzlp3Jkk6taOtVbN
UIqFmACgPyxxsNABZbDbOn3SiDF9unj3IVQtkM75RKVjEK0gtUBcaL0RehuUzpi+6MlRMrrFDWG9
hvJ2hqQEonOIfmH+IbNFjmispRpcIMimEJfV2ICdWjBPgeMl+iIhhzXQCbphrsK5aOVWQfZs4FpQ
xe2kT1CjO8HNzsMYYfdOxaqGXAwZsaitSnuoI1dz2aKjgNcdn6Y4QyZj3PHh4z6cwJW7hG0qX6wa
ma/uU0Y6gkMLg2lri7jUympzpKV9ZH5sTB75FkTrfanZQ6aPoUxA9bnY1IpNmRdc6yf12HP+B/7N
nRB3FqxlbNbWHLY/vf0cpm4BVRM+ed/ZdFzCggPJw9/sUjUs0hGBBC07bOyV9tZ/0TGS/DjZhwbx
bamZsM86XlSH8xn+8MBqqVlztG8HukdkDz8oqGriH8ysP6HVGYU9wKzZvqTKorgAZ11zF0j5ggp0
eP2vEkidUuI51fy+v+yeJIILCZgKc/BTsB+1rFEtsmjP4onrRchTZNMHjhS5wUDEaUkIyGQhwx6S
rgADW8wOlYygLbi/BYjtSYAIVOPjCoMM4pOJtoRZpBoz92J1+CxJchTbbHqj+FV35IEdwxml9FpC
k7Nvm24LSkOokqidwAxkA6gxtGXTsMeu+qYKwdEThaVPfAc22P7pD9bvvYBI9jHKh62NypbqxaRi
SsnrMMJDHRxqbE7nkiKeVlkd6uzPp1gn2MCqqr+nGNDeKN7n1xyMrDBBFBWzT8uCctDfgfS/yzJ9
mkVkBY5ICFMci6MOtPTCtR+gtNUVsb4Ns4NCgctcW6fwi5W/R8nvoSkfdCPrFY2B3H5J1KJ8CVij
1opmIkXHT+sp5ROSvwT/Hhx9tXgWukmTi6AgNovX5ROfFggzfnpdxdlHTQcWW/CDVqRnkEmGT/mg
QTInjQTDT5YZ5gSpb8jsX3MVJhj1EFaoKDWGznv4zbIp+kYrYXV+UDaffJyZTPKj9w8dV7t9eAdv
mU30AjCArkcEfLiQmf55H8IYokR1hJQcbDx/qNrtkbIdfCW9iptrugZrxNM1xVZ3Y5+87Mfg3gZ5
DaDoCVSrLGJBFlCwZRjHxHEilFMkTtPTSgQxLPgWlVJ+rIvnPSUmEjkYTC5ejAphGw1RmeI57Nnu
Ig7ILKBtW2frUrb9lISP2pxxc6z/pszO4LT3k+kHS0BBBRuK4Lo0/7+y+nxo9h8jNkEmHXRJO9AD
cPukX5iJgbyyK6sWAK6SbE/ms6kRYfMkbWU7zeAracDbAOJnJLUiIE2nyrvhMb3sMFbixN920VOI
0Tx/vUu7msZBtgDhBbAnvYmZnyk4ajYW3lcggaOOszi3iobC64enVIGoIJ5++05o7fiw9otbASVz
XK6eCWoc4ADy9gPbzRfodIo0zG9AYuY+ZeDoyumJAeqNEEpoNaaX8qn+cV2VzHZU88wyQgrFXEL3
15yf8vC68EoaER6W8IQMlFelXmQtnMTM7ll3bRZGySRVc2joz64HQkeBOgIliJT2AvGtmvrSBxdP
GwDlbAH3GxyJChHyTCOF7qbJsT9pY7QE776AHc2G3wNbhlyeMk7x2y+1XNxtMq/xQm3tZtTJQ/jH
wHewh6q2x2/hrylyF4k13fuHDSpixGqATSUHjn+adx9gf6qQ8pi3b7/ptjmyXX1SBurpZw13GF+d
eRnooY8Gxg6ndK6Y7vcfn57RBroQis5WddG4eZTJ5CIMcAZI4x89FTzBhT+/3jJsjnan1OQ5oisE
PqBKJbgIKxg5hNlXKwpreLkyq7Wmhe+ZV2UDl+5sR1ZTmFQKCaq5rEQRVDQ4EzfeGOVQXHSxmq3K
TQXtm9qYq1DP6LebMG5TyedfPWpDg8s/fWWPx5ro3Xv0+4x4J4xz8DZxvjBOV20jGuQ3IgBqp+kb
1rcAR9s52pR18f1bgPS3tjM1rglmuZbWF9UfLXV/+8532ZQR0ICrXAcMMLGOKnDiwh6MCBoNIG1D
ZJ7/VzbgPB7WxVXNKWaA0HVnfCmcmDuVE82tNv5M786cvZDEhfzyNKbFKnFf3XT4Ywdh/r+KQCin
vBvhdJWJQb3qj+5sZ1LlPhLXJVGUfXBNza+LZ4ZACYZFm0GcidfePP+twk77I2DiI+wTOX2+g3Dr
ocQNf00BPagkusq9IKzWY+gNkZOPME7/bFJ3JeMj2575450YGsqAxMHP5lT/roBPyrSZFWkQtgVv
qxVWNMdsOtkbSd4nyKftisSXIDPYNF7EIsIf8xokXLH6HUlgCVhM6CCzCjZwyjmRrXAL/7zWTVqZ
RHOm2Ma2+l2j2fa6VJqjmNJ6xFPjHAvz/Di23xJOn2FMOZtgDaZmd1KRzKiPRFadOXh3teo+yOp0
BRzBmgIDk+OojTT1cBiXfW6Jsg4Wai/C/pM2rnIAOfcKZdSvsMlQwymGXpuRpRvAvaBkbjINWjpS
zlHCiILQRhOUqR0W/IFo8LzZng1MhVHPQwA3KD+rKfhmZ1d+kFrnG0JHvFmbOlBzWO6VL6TLp5WG
AEcfbvFf2+4KozZzXQdvN9Cl761g2EmcPXFoMyYiun0szbP8AQLN/Gqk6MSz0MbIqx0LrYp0rsOr
TJG2UGaau4L08cSkOcxndXdqlSIFwCQvsqVUAVzODvr5Le4bTbzHxdsz6jjvipupR6Z15zCgAZFX
8dpSLeMHCgeyPP0+VZ4ss7ad4Q9EvvFQDKvl8uxI+zPdK6vqUwBRDrI8E3Od+4CmcYoGKaAVg4Id
1K15/nvP/q2YIoVBhjETQZKy1mT8VE4jaY7lzOtjcwUB/itv+pa3/6RHvyR3u9HfMao5O+tA9KU+
9gWMZjYHvvdHsM2l0WI0gH/jUDsSE83qCN7DZnG9uff/2Qc6FH8xlL0Li2wwfXUi8ZLK3fKME1ja
+UNJzV6C/zOakRqEVjTO/vISbuAfzpo3oLwQmsN7swn7W8aixQR6Sn6splAI4M6zlafsxSJf/raa
p3KQJd1nE/PdiKuN+7QdN9Q+BhbBTpxZAV1gOkZeIQRmMCfNhilViLuiz5JxyXZ8mQ6UkNN8f0Sp
e7aI+BKO4PwcpkVY6tYbaUMmKtMxq/UJhdVU8EWvd7UXfEGyauLogXlFtgPYGDpmrVRW+crJegj9
QaNDKxIIT11ZJX5sII6F4BGQQvAuNVxq+t7HOVWb8QK5y1jytH5WOMgGY6TMOj9bb6DHHGhXDPok
daEAzduOoK/nXxwCZOnY/6X6KfjbPNPvN35iT10ebyFYpdnOjTNfL9fAbi8w66FTCsIhFVRyfOYA
lScUdGgCJvmp3eZLb5bwhyRNkV75SMbHvMcJsow72y3wFHGS79jnFb/yhkOs6ogtEsvevmsREbg+
JuLGMUmJxIcErALiZ8VmNTAFGjBxC04YthNEmjJSoOACOGik0cUh06Yd0pKVc4MGAqOgVWCD//rP
EfB7+P0LnHrCLmnUmWEQZv07KF3hzG9B4DI6YxFoI7q7G4TvtzbkqCJ3Gfj4459/OtU2Jl0MuX2K
naDiJj+F932YTTYfwkRA8HGTtOnE/bWQVQqWdI3DYIb67/7gI+yn/dcnTJsAFa9wIfkzOBff3Niw
e6Sy2FIzQWBVoAuQnUlN2WlQBhhWZWtfPfl159KQtuGwTawxc2iUpktRbZf+xq5+kuKPNA5SJvVK
xVCMFw+mUan4tdL70HMFTUVegj129zm7wCb5VKzE8OXb3dVlG8BM6275zjQyFlliTIYkI5dD9ofn
ByZu6Pq97SUuYFDnu0aZOvaw1nkGdAyQ4IZaL1/fP40oH/9nSJT5Sfht5VghQao+M59RvKUZi59c
SwI9E2KE1fJon+dS504w3+P8tvWaRoYY/llzqMGlKsdHJZtFDMdW6wJceQGMKrfL68Cp8elbk0ve
V5NleTolVY6GSCkzTque4tF6gXpSMs08LMVbuJiFQKoQk/Gm5vUrcWYKYmVAePk7YndUI/hIjVDx
4jtKVKu3yOlz1Dv2DBlFDXpeErlGxUb/BwHCa5+lHV6vPjeQC9zRaVCj0aN5pCBI3XZwYZawNygA
ZXkmEuUs0yt6R5kHr7YMdqGiL9Uk2FYdtb7RmYteekf0+WxLzbcxhIFrst0YAiruoK86CBP8xHsn
FslasfPrlP+z5d0QhmsK6PAxTk7v9aOpclGOWcx3BLaeCdj+T6zV1IO6SwprFJUYpNZq2dSANn/r
R/HQuham3NY3xxuions2pMmrAa9WWjQUwEE4hHt+0RDFpN9sVLv3601ul+AV+YAS2IoiTufU/19z
JA70YFyjo2h2hTXxTarHtAuz3hqCIaOYFVTcJVlrNeoQIU1Y4EdccZbKSbjKMOoyq1jt7CHglO9y
jdiuz3oa+TDx/5o/a3o+oIt2/vvC5PIuUvwKewKzICVwAyxyMYOirI4VzW+iIMMvuh8hAncFyUei
etJCFN4Vf9/7RDa8VmgVep/9y6OXaA8ncdrmHbzNPeFNIWyM91SB3PTrkUp1Wo3gtXN9YgqTo9p6
j9LkCaXx6VQrfIOmjeTiaGbojJVNNVvGbJ55peoWTPB1d4MuyOBzqa4qpvc4khcQiXqzAZunHFBA
nzDOTZXt9103EGu0nvPpmExLGOLQJGzx30qAJck3mUt/LrigpqOpGEDa8zUnqtPK4aMLx4tPkj5A
iUyu4O7/zjRSmibpXWUD/DVUVzT0iqY0DMPPxwZOwDx/+Q9bP2EYvhdldF4TUncLjkc7tJPsTCtt
LH/92+XcCE+juP4Oc4BPOgOAnwz1nHj+JwfxC85diXdNcM8tmb/JLCtdhKFsjq0+xH/IhIOCYh5F
NpMxc4o6lZgNcwHG+TyFDCCY0hRN1T08dRJmgtQ5C2NJGAHKkjR1JO0xXP8lyEmNderL+zVVzT81
LYjFXd6UBIz2GjFSd1vE1JsO0f6EgUjtA9mPf4Ekfm92soIbeP8lyvP1wuPZCoOj/vOFzCMpRRqc
M/pnc3bgfKnFseKoskxBdb3hBP/GAwWUheArqMIw1UcQR1rQEANqznaDowZ7V+kJ7loevfhweXsk
N5MKd4e4t4GYvdYan6in8UEsoqTVwnzVMFKk2kSwP4QPzNpKb8sBZXm70vA2N1KbYBERoDKFNwz+
PSY1PcvLyobpA+cXHNGNmfQ3EXaL9vNo9pZ6iSowbtbNAIcuQPAbk1P4QH9HucAcmDr2Kl9jbSm/
sbPcig1WENv2+nFFbAGMbN3GEmgT5kDeZtdPxjgh73Xk8MPBzJJJkkcSGKqnQe5SLXYUaymhujtq
EbiHG5nSsJvjaPq1KwE4O+e90TpZa8A1GAiQtt3A0EifObKggx0+1Qo+Ct5nYvuIhn96mlOJjtce
ATSJoiUSRjUcUg4BVupYtbQnYKrxc2EhA9v/DTBZrEKore5ZfCQ5HVvY60SBJ7HVjBrYBjqxuOtC
i8Og0I5m59nMLUgU0ztN5GEgkuI/C5UIJNkdECLdsB86bMuD1XdkTz2D/E3QTIWGjoiKOocL3SyN
nNA/nged5LJ2q0v2fIiroULM2GvT2kdR9hV8w/gEG7saX6SUVKbv4FzmzOPhAA2UmS5j5fiartoU
Rha0SVc6mMJ7Nj6WI2Km12Emr228KDnnd2D1U9VUlqWZZm75dGPzG43MS0Xl+UMZ3NoXzgW6QBBZ
nZFrIp+9VpsPgp9iMDEEAwCwixAdyzm7AMfN37jS3iBLjotUJp3J45RWkr10be2cYuBXb2fRhp/a
fYDr+ix1oTQ1ehD0bpusJpBrJSegRQ0maLqZ5OJZqlR4J+W8sQKYtHOYHcibYF7vHilbZVA3+0qA
5L+aAmdoiDDxTkmq+AITMgLBAe3nQ7JEcNC7PNZk7aQGavTo7qX5NvXVkxxLsXGVULCAGe7Ky2dg
wS4MY2/6p1xhMssKPU3FQrtpECafmEvdP5jPLHtwsGHTqDCyCJRUZ+JcABZuaLdEYfCLgi8m9NPE
wgGD3FdqKsAUKQONTwY159E53NPNjXW00DSgFAr92k0/PTPJf5rFg/LatYb01E1ojy35WWnFHLWw
ZGIG0OUSg64Z83EiSE6UyMmVFIg/6V7WKBNaTj2uqc+kQGJoUIIZ2zm2xTT/cPTYKYnwRU+ST4Jc
TbPwN5qnTOCBI2aE2lEZrtauAfF8XNvicU+SoHB3hyUs+Q5ofuzmCYYpLSw/En3Pe63e5ubKv901
GbUcKnSCzee3rg8m+Sn1Sszb24tEqpHHfVQedrSdaPmJ9fpRUm3cVfwLZtvgU0g2mk+Bq4fAxNHC
sgghoNexMMhH2hXJevlRpMQ8zSdRZs+fv3mUr1+caCfJDRDYBpAWjrUMVWlLkugz0YpED1ibNUtL
F2+/oZNCPDRoCb3uLDb4JDMTmbwOr2/TWvehTpVCOocOt/xmZ6QeC9oBoXIEfM+m0VP1TSCFjp07
J3WMpJHrRa/ES7by7M/uwhUP54Yuv6NNatu19vm7bfVS1Bj6Y3V4wYXlYeO4IbtqyP8Hj3JI53kZ
JouVPKUS5rWmbrWjU7I1SqXnQ8vmlMeZ35T5VNOeNu2TvbJd1zugCFACdKq0VnevRzitgRWWeuw2
DHyaj9ny/lXklBfuN76qzXtsUCxIgI/5HM2MH2uKFBLwj0KCMD9Jk6pyhTDR+vYh8ER01IsRhosU
vXtjcvz/IafuHOFemVW2Vmdg0Q+k261VD6kc3hd7qw29dA/Cn925fVYSI1OyIrk0GxF2NsAM5YqV
o0elWrPWEAaRLdLDJoou5eQtnm5y4N3V4HhPxKfqxeHztQeMjFaotl7ifnNmyaNFM+fp6s4jSw/D
xZjsuNbQhlX9m1VZAc3FrvSGgxe80YF8NOo0JJWzfk+p+0QpY3ppt0i2OSrYL/P92N7lYCVBBNvr
NwcbgXuy4lDl76Rz2PJKscIlVOlE+YFwNYYj7VsOPUR7UZ5fujqM0QIMtuAXI+KUn1X6PrRNjESG
2DSUynGNHvEq74Mdver/OB5WXSotUrocpJYdhCBPQSDTUyuhJUvdFNkRBXi5gQqNaSG5sZILpXTS
gFqoo/oN90gvaMQIz3qH5zSeBd1gw7F/2ToxCJDASYY5mpw8FJnCRlKE+RC7SIyoH5SWrkS8JTNR
kYCnxVmeBqvo5U0YggXyHe9k9XLtuO6Q4855CaFAzN7++Wz6bNd+3Et0vU9Z/tt7ktyW6mOk1PPl
E0AqxmhgP+68nJx1NaVSg1INDjglNvpbu4NWJ5ymXUS1CYjfJQRBkuGA4b2a+W9oGEq0+2ro0bFO
Onb/68NRjrxYR3taafh7YlqlBY4H9vqzMGkNf9VPLPqD9o1yRWJaGrz1+iFgqTFK3cTWcnDgVifY
0nhLFUTaMZisD/eQkAuTRliHHt9m4qscdOyxH2YbFSugYTf9/n89s4elmHBHiDSlWcHtdznFU7J7
Z9cMa1XPFOKKcbArHNG88N9zuaohSg2iN0OkJJsqX3xlS+YGl/g+tm8XSgLk+pC2MaeNu6VgrryH
cvXYzmdM6sPe5DOQZQDT7Ppm7tenMmCCymJkXF66G8j/3R0TvzjCML6Q5jMNh+0DW3QKgP5FWdw2
xYgHye7MML8QXGQfwDshd4ATOECABuLUwuLMNn3JLCoelHYu3xvjgSGH2dsdSr/6JN+unUYHyBpV
H1b0fBTQnv/uvXgOrRFyVcqjLEmsfQetULmBNjo/rdVUvdYCwFWEDV4LPISYg2Ff7XxM7BSjS0Bf
FXs0BgBgwzgC7/UIBPuI4visCqh6vBLL5mysIrmUvuK8D5tTDSxvrq6GrFbTkHto3qyd/syH8EzV
6l/GUNQOiDGtiHFv2g7SlVVyCQBbsLYxpZMflupgDOb0FJPDlDUXsXzrQ8hM5zmBbCW87A5FFBJg
6Jf68bgaCu+STDc9hElH/JvcL9C/ZfEIRelwvZDGFkp4LEh2E7S8t0PPC4OiNkbrlhbe/KEH0Xi/
LRpgrMZKco/1U3WHWlxqUKyP620lp6tCKwisklD7nTBtwVpBdc/WRcIdfWKNhaGgZ1zGUKMhQm6W
bUy2h/d0QB+iDsHzvlFdjh+cPxRHD8psNLqd6aOqX+Ly+zFG1+3DVB+bCoSLaG0o80e3L5gTcArR
e47BbN/d9je2lL7Ryv65CdUnxXyU756tTs9ZRYiy0ymqTkr29W/fpr0KjWUthOZ7LZ9pR0e5cPfX
VUzPKyn0597PYZLdwKeaFho0RFBuGduqAC8YXNVDbn1qXxYWhd/AQ9AvWJSO6ZEzdlA+FsZHdv5L
4hBXxxyl1y538UZM8dyCaVgENSzNtIfYsEyhdOtdDUifZMCwX7oLNmmb5MjrF9YmHL2TuuwnBcrE
dupNHpM37GMk1XBHfy/k4P/q+XjbHW1ds0ZQ2PvOovTv0pq4qKhRvaeLWd+IyTTDDGZXyqWMhyRI
fsQuuL+Os4WxLyknYNCNcwSJLZDam9FLDq9QBfvPsFT/GU3FrN63yi1EzGVkH2J39eSxeTwt30v3
vXPU664tOGEaBajR0O/VQkkPRN5McgGxmr8E8iSCnSctkq9maXCVpG8CDR0kzkk8iJgNQDNOBd09
+/lGzTfDmFkRtCmGFk32P1tdM78TFijCASLOYYyNRLdLmpc42qFk+iGyNu4Xrfhwz3WNwz3qxf1E
P4WQr6SLha0DTXTaqg0NCt6gw1mKLIke1qsis9gIS+erpK1CX3jo1ncfVBkJwHLidfl6EM2ZU0AL
j47RtNIqGGFNew22A8VIJXqndswQ9Rk6YCaP6tponKKwEsJdYEfhBtKSqjWdGeSp9uopgpdAqlBn
rO+H/ALCk0qc9xKidpPvIvqHtuyBqojPZK4FPSGLDfpeZ/wRw+H0qV9mZDG/MsoVl0kdVj+noE47
lGcc1Am8eDHR/Fb8Rwh8j99Kv+CUf2TbLGLEXoBZEnsa+ksiPX2d6kAX0kQdU4PIHiMPMqS6cMoG
22/XSHcPHPWJgYtNhzsqPewkxyIPjEDHA+nDyMWN1OVFThllYv5dP/13Nt8ng+xt7Jh11zOC6JaE
dWAPHBN9HlhDlnceukjWqknnLqznOadUduyMk+IkFlIhV5JfQb6SPx23Fqk52GiNF11LXltjwzVM
SYRx+0Nm/ZBhmAwu4eZ/46uWY4URHequmx4DKTljQpNn1Go0coxw+o226AjG6mY7XNS79mkCmXVk
TrG0mNIn5YJI0rmbVpqwioZdkn2Df4bjm/HFGwaXtWZHVy1byqtPL/WHrBdK8YWyF5grNt0OtsH3
M6/Ef3QDBeh2T2XpT0uT7J1ewwBUH5X/Zy4ShPEUHZchGkrp7nc3CXdBwcfpYFwBJOuANSN0kOfA
zhH82n8xNd7FKJvIc/uEM/JgD3asKw9LPZdW+rtk4O8ElUk15ibSNMhNoaCUlYlGW7EOD9DNuJKN
aVvpUAcQ27HKyDFh8yE2r6sk93fbL/1XVUcaf/0xbWasey1iug4almY2ypCU28PGPYe/wtw5A7LQ
SyYk0OD0mxcTaydNcqE+RwQaPXNWuFLZyRfolEdobnF7wFBEtI5zRo5lKbAP6NvoMa1JrUa5v64+
V/6v5O7dEI0KdmfjHSq431jR5TN7n+qsyObDf4K0cfeEPqRs2mxpklQivczjt9YsZXvNKxkssspo
UVa4OBlHpKpVwdcI3G+IC7GJLpnaZGWO8OPjFDXSyWT4on1inc5kat8UfHxBA1+TwvNGjseCJdR3
4V8bnjX1f/wvC+0chMhusQDV/ynbL3sbsyjtb3Ve2/3r4AQmSOcD0McpGtKtrQ+2mDhQmKbEZ6xV
id2xMRD2uV+cLm6+CP7a7M2ZF76NQS6RlYXhAKWayxULQR7P04Ub/5nN8tu/j/7qZ5SELEt2xDzk
Ww7wZv5nXSCqexZFbWjvZ/WXkl3v95g9/C+jg8GLbaVAciA/BxhfukdwedAQFLVwhWhxmq0=
`protect end_protected
