-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
PW9fkKcJeuTvPMTByVDpQrMddMKkgDkPUdfLNjEQQVBrvgy54Z3hny5wW1jC5nRbv72NincmbTjN
rj+or4W6KDn5zLtWcxtV9TMlWyuzmcgVJAdLbzp3LYjkwahvlTxeWEIK+Im+kF5kE94dg/xNl1LJ
RZEbwRDomaBzKTeyVs+OYqchNu4rivj2B/Ssy0bvgeqkvaWS1DikdWXsk5x22mf+D+jOmeJEp3P3
R5qnb9dreHXYG6DCz6nyq7RNviw8D4Vuuki8t8YJkbiTSr8FwcTpMBhrNOYbheqDDzv/WShfEI27
tRD3/ipohwlWKJwBFPEX0ef8BSkspNixrOpNnw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5312)
`protect data_block
gnVxaUw1QbgnYpOjoOwZZgRMt56+VbjdA34J8YXmvjLn5yplYwW86WsnclOIXIs3abqnClL372PI
akXizhtwjCKopJvO8cQxsl5NQGkLVisKf9MVQFmV/Z+OHX+8qc5RghPCrfKulcMWy/oXc3YZlxn+
gPNtUPQR05g/U+r7tnf1Sso2aDW0w3CyFzTon/Zgiv/APJiXWORnZgAmNsxbEiTvgnwV4O3iz7aq
4dJfCeUL7/c2PyPmlSpiSmObi1RvXPwiB1ohsmepopt2dyK4YsmrUyf21HE+7d9McSzrqUz3i1KQ
XlEZGVwztmgmrv9ZyPeRDxJZ2n4xigPUg82M4e6Oc/O3O9Fc9QPxXJUMHGZP5Fm1plWlR+z0JC0D
XUuoMUf+TWzujy5aEHgwRLqQJnf/o/M6Yirt+Vs4KozCyhlXpR6KPT7yXV80DQJcfzX5+9Xpsy6w
Qn8uazFbi+l0eBa1aISauIUyIjFmi301rVv7K3WlQpbFkrjBVouWso1RxPZOPvduCn9gSnuJHVn6
Ry/tmlqAnKwkTHi2A4rkTgEGe083WZ6HSTbK4wMo6XYCrtHA3JSh0L6DE8f3xRwukUPm/YYgRuRp
DiFyPYVajs7YNvYdSdSEuSMC7sqBiDBcPFNG8W+Wm9MFYWqbnRo7jbX32g3zQ0qhf1kBFF45gvFL
GUMHzzpwlm2uGsDSGSrNKpBzw0S2sY5E6jhV/E+FNLSDcHbZ+FzrxETv2iltPGI+NcxTsVrq7yST
WCDLpEKWwA0uczDnALezX586EI6AuO83UlRFWRfM59SxIWzMIHO2b65NXX51zZDwlKffFHPrEK0C
/tuJF7tdLELR9BEn5ao0L4doSxOHED6B73qsg0ZJi3C7nn7Jf1kOdUnrGQfiHcJovAceVjyn30Oz
YUvS45NZQzVUyWC//nZznEWFtS0MAkSjPKUOMMgBf5hmorHJhFFc614xOQWOVB3AhXx9e8XcuBsp
l/dzyPeVN8k+3CJ7yfM6mQZn4Vt5E9yDLhJwrL6S2NjutjVclCwpF1/W2/FDuZ4iyRDCW6eNWBVE
Llh3kn20rota8REUmQgmsaaLAYjqLwBiNzmSGvd66Tqull912TDzW9+eNCgrsH9Tw6o1cnQD+H8o
X9+IvFzAeqt8AXI3I/wauLW24T6da+Q8i356F/aEXL/eDBr/EhgcP7AEX0QHFDDIOqZgcUAJ0fgf
VFMIACJVLkiQixBBR5hWvurITdP9MoBUKZ34K1s8KKo0VPeeSqB4hw8OzOveXF+1AIhJAb+TwI6w
VmJ3JxrY88uMrRK4O0mYeXn/OoUpebXf29+xYFfQWhh5w9VWe1HiXeyu/TX6KhT/2LtKRhuQnup5
ofwLYSAsCouJ739TiOBiCiII6fKqaB2zKDWN8ZxOVJ2RVdvA6qDSq/vC/hXEfoPvQwQcOx1GzI8X
OVo6Bc7cJkVw8tV8MIhBfJzzY/ryP3mkd9rAHJha+C+rdyIS+58ojzuFjiGHJU+MRTo2ObnFw+aE
kS0rUAtTY8CFx41YwsmnsYwQfuA8f26aWui1UPAgThDsXPe0v3NS1OpjNjlI+yEKAylMy6hcs9h+
8lHBieaSJzhMhzy/zXQdajpTsGtLt7/FMuwbEi9nvhc3pxBvnUYQ7wgieNjK5zPakYrtfrYpQXl/
AjxDUqgNXQclw04jX2t4wrM8KtVca+md+GA/E4QuCm1180A/XD3bmenM0fjf6MF7eoSs4rfIc91T
VMks3jpkd03CsSdXwATTFyIP9xA8XT3zNgkwkbgjb87NV8u2U9RmiyKiFV9/AIEeJRI5UVaqc5XS
MeYnm2Iq/QiaLuEYjSMGYUtTn/U2Y95+DcolgYVFHLNhZZVCr4TOKnWnRDWYl9H5YlCDqjXGICcE
nNokUaLur3vHufegCNAXdLe3OU2VxxluVAP9MUd2RP/KwgCjWqIy4M8tfibs6R4FvimtgKNUWi57
QNAbpqoVpJAROf+FnwgQsVmLlpaBTngYzBzjxJMonCm7mFOTjnvDTHDnMMAP94JXnraLdGU2B4ON
LVnhYLTnrtCHPrGLPaJAZq+JmpphqOm9HEEMMnSeievm0qR63UNP8a3Ha0vWvx5R0k8qQXrmUUFf
mqHPTjRDCShnxaPFg2mt8qxNF/M6R5MHw2WfCCnIaomFCf0nY4wsM3nsFveKin06kBgCLWIxE79z
ELCQvWOWE1PEyfNBXJP5v+l4zNVwlOJrLRUO/oZKwngHU1pA5dbeklnkdxm/Y5X8uutmv1SHmut1
9G98PQGWNqyJeb/DDJzCeLnjaNRmjf2SSDZdgi/aDdOWy25ikSyhmZOY9vSCZTNL7lI2F3UUqW4A
veKK+cbOmsBFx3453ZKxaWw99lMWYZlHIVgXGRl/z8mH57N3LvO9pf/ZRRx96/VIqsmyosk44Laz
64sXx75N8ilhMSbaPjB5drMEdXO/FYwvW2Xfu3VCJ6EAJ6+6+HPTIrq8pLFyDmYWhEldtutbknN7
lMXeSsYucoOZz2H9Wrjp3OW7L7QgM7XYqgkyqA21DJTKmn9rE8hoEKpCZ0lR35dsRozA3f/2UZBP
oEn6kf6FVzY7UZk4p7smX4JXdc3v3W2l8tztESZnTrcAqMVtElhjwAr8E8DOVaJSPVjloTUvddR/
55N2mb2DM8QCAoOIGs7uMAXudPpHIGzqF3T/yWUYUtDD0R9Icsqcl7VjbJzmau2YAKshh4MwViA4
ZivauxaMd8BpO4JG0fA2hWGrNU1PxlwWqsP7tc5+wzGftHrmfq/0ZOQaC9ol2i20/dmuB7OUpogs
bcidR1Otv4m4To6aVnH+iVav+W8dZebpqhVukrmomE8qtQr7e8sS252LP6640C6sPpwGKiAVIWZm
gvdmZyYeI+xFT0LEh8HAXAYXKYcznX7nJXCD4/ywO35W5EltEt2RqMpv/Fqyyk/Csg9leqE371M/
G4RqmzJFX3kKz4/0Tens4c61SGb4MGIP0sV0XKgApp/qASdNJUFqxyJuDqOOBn3gFUfpGS7GZ0c0
SGqkqYJuyw1QTstPTsLYWPB0KL2UQGMua8CbZrc3ctJod6ZBhRGYD3rTtr472e4shSgnI31aSYwS
XuwBClfY2SVPCTuyxNxEQeA2I9/fT3q2NtGklcj2dMNUZxpeL4fXYyhynRNxue6ODoXKlgwEwoyS
yayXyjYuBy622dsyHCGuJN+0SffuXdkopHJaY8PAet2QNUvqlLbT9FKnB1iG62aX3dt1Lw5v6bV+
vGa0nrh9qJda0NohMImROuFdiOYyQ7MhMYgSE6+NefvKXhPKHQrMqIPidp6ABfltXcGmQrMJbZH7
B0ry0HVk6EDGLf0q7xni4n6CJaw/I1KuoLXhAcflUW131OnUqx7ACurS92oqhjwyt7Ya+WDZ67XF
SptxwmabW+TmcAUTclAkOgO89oDyTd1xTiTT4gwKKkc+XiKM+aUwZwVZv4eJIHOgQ+49hZ5nC20+
bmMIHQ690TVsJUiBjIqfl5Ippk5mQ5AKmLR8np8BpQhJ2+hTu1PY26VeL9dDYuPiHI4dnRoiW9fI
9FagsQuKopKdt3EgKW4Mhk0Fsb5Wvg2FS05gh13sZwGKC1yOP1tbMOe7ITd4/jzUzarsseyT4EDB
tKc2YJH6U4SOGyOvRc+rW4m/sku7Vib/QoQZL8vaC6dKu2du2QNATaAOFLEwLKwFQuy6svEmV6Ik
fGcblQnovx/HAjOkEKxzDvUWjDEBGUgCWZoZsbe67Zddoq5Gdm+EFsn7uFQ0Ka11NblN9zl/MT6Y
EHqgh4tKGLigQJaa4fi3MSqATr2WXxkMfoKAVUFo34nTTZUJxxAGUbDonXG0lM1nXSD/l7+fPZnw
hi9GX/4yuQ+JZW1xrJLO6hgzVIjbpGMW7FDd5wsh0LnM8wtB3M6vtx3ItVAiYfElU0Y+TYK0wpds
y8aPXphj1mERLsZ2bzwarsG2CIjKESUwgD1F3HR5Uvhsen9QfOQr+LmGYM3Hla87yoUhiy1TZWcQ
b+nwrXhqXugCdGVZTRAErRH5Ol0x/1Vy/YnNVTKAkAyB+WytN8KwZilXkOeH+KbvAqCN88ooNWtD
mcb1PW5ZaVE9g1HgCBo+xOwt/foJHjhaajKnTVp9gSG2O3u4iMxG2JCAexTTazyVwiFYV0eId3d4
2fsKZADyjPdxZ/kAutqdcUGrbiN07+BpJ+Z3EEmppi/b9uP79lKoBapkFIsxAWqEPrrcc68Nf5DW
/lVCcDGz2Zujp7mHu1zXU7sQvKsrk7+bLlw/putEDWUAX7hdIOK7IJALOnuNfBEx+gQ1QscxBnZ+
47pgv6Kz7P9/Yg4mHQKgqOLFSfCokJDF5TS1aIA6BewxjW6uYevkqL0dOdI2Oq0KEnRBLwODSCwV
V3JYzxgik0FS8m71fglVRlM4PFWLmYYJ++AFCsVoESlXbspnemBWygRTlksLGPAtp9232pHK4DnM
KphiCIdvTkLEQyfYt/zyFBbLXPj76t1Ev7l8S67twL0cuwDeH3qgRKqTBpp+g+ojJYJUzrRgu7L8
1INKx22Asb48jeH4K80JYeSVX5x76VXPffepOf0FP0BoX48KrTR06q96DET7F04KQcTHciYeMUTJ
cxy4jN7SkU2jeFHohBzHYBNXjNSSKxCxOSKiipy8wwdmlZAnIsFJWaXSIqG5mFJdFD1Qf5R4V2kG
ewrF2SbcnU/wh3wsLAGNPWfabuhd22lNWhvNfG9ar2jf6pc3np9NDoBpnfxpWdm8xcsPfn0+io7U
KfXm+WQWJ2v++2qyQFiIXNMylUpGUnftPkHue2F3DZRfm0cIOQwR1d7tSdxajRewkl7Qbnx16ZG9
okAP18iYVsTAmi5uRL/mbHHVjfNgF+4+LxjcjQIVjLbmrEp5yPAl/o1uVmIgOxVR8MoATSYEY3Gf
fRkvGh2xqJJOLftWHfz8SMtA+9A0Hz1mjZ3qxYqUtaQepDuk4bPQ4dhXiuwizYt/678mBQU6tQ6R
HgqFfytcabCq1o4rTZhHqlB5TuG3EclNgMTTadzsqlkNYg2YuSB0VREpe7VlogqKO+9YFTCxc5cw
YkNFD4pWwT0PZgR91bLMwe/KG0kivkhuOO8dOf2XozQ7rPSWM0plbIsBRnV2TXsNwtA1S8m9NYaB
LSOgDAIt+qPJofz1eD8gA+H7xK7Z/1HZLS9ikjc/x/WWutxLPTRz3PyGESnfkyE9ykVEaqt1tXdc
UfU4sh6etcZgW8BJZQ6eC0IDT3AUCJqvYEM7XV0Z6hsq5C16wIleTTQCRZ1EMLQ6M1Dr4+R9WuG5
mLm/hzEYIT9iD34DuHMLkYVMixhgutwJmVuILOnSzzZ8P3ATVCY+aR2MlbzNl+FgPbKxF6ox61E4
bPqGjRIVler+//nrEAIi7V9xHq75z4C98jpW1Rzmnf4Kc162aTP8hskGvkEJgbKVJoEv8rmQPD+3
LaEHRBW6jQn3LN4IFchrwKcHu2WIYx1lJBj7zj2cTiPX5+GDz2x68rRwYFzzp1V1u7rau5Acrfdl
EszROxnV2gj8f00IoqN1p/GWlBrnNqj3PBphzp4RW/yuQ2uYS7fuQXAWU2ag5jYXrcNV3Dn6e2CA
+wDSDNuwMmd3aFJR7KONm2qKW0NU6pnvM44HG75NjPMnLJ3HJd+9kkR9YCLsTjKw+lBZBkh3lvLF
ZIi3/PHSy8O/T6/QAXo5DGwmICE8g9iWMUXdJJQQ3jYjSjuQgY3sFDQhvED9inK7vRmJFAAR0n5n
jkpLXiX38dUWtvS+uCu1Rp6cc01xvp1O2h49I98fWgb1Wb064mDyHKwA0VprQg+t1LRLn6/uHc6q
fBpK4LCs5O4xwd3bdbOOdpZFqCEUg3ORO2wE44MQan5nl68irEoifggAHIQKLfnOwygz82ajG+oJ
IM9bd7IyTofe3yxGuDME/GsU+lODP5xv5Szpa22u6Y4M91/aS5abBYkTOfgSNQbJEMUdO4DW1PDV
4YDgqLErlzU579aRAiBUKRolYVq0yf4vbO7BWpcU/1BxaAS0PLM4SNpYaQvzJGGpDFSdlyo7eyHk
3Wp95zzSVpqXxltbZouqWmv2ceSNDBjhXVFKtusTqpWoN0tnqzpasmcdjCZVVz0fiG55OFjbcxsl
9ItySueyTRJ0RpxMiKZS9tOkrCusYwVKmzCMbyEXsnRuqh/u56QaRXJdvNQal9B8Sl3inhoLDenh
C5iFnzQx1lWOokwyYno8zeGdoMmk/YB97AaWyKrC5guEcHMb39ikjCpmPa+2m5D4BWHbSkXTdpmW
1lz2bfAVEJMQueDOQDX2Sh7PfN2SxRM8qoo3QuNry5qRl5GLmqc/b6JnE1ybzdEmGmLchJn2SLS/
B6WaqZbYuu5XwLFxNNfH5Nbdft73J/4c0j2pVwcTvZ7IYp8LRjxpgSKH5T4dDF48dARj4WG3HQs5
t1JIhD72AimyBSc+pNlRyr3rWpEurWPdhtL7hu/kOfOu+DSBOvbnZ3rw2YUiCMR1zujEUPrjaQGx
lTmzcPNP+oEuMif/0OCvk1R1X0BiY7vmSg0vhMO7OPLWpM5z1n70OlAa2yu4vtxjStBvrJNOgdsj
7+rt+oEqTdXS1Gh/YwkRwClBV+N5dNQuu7wmtjYF9YVZ7YDKX5sT7LVk/k0Ah9rHYjUOr9cio72G
aYx+XWolwDM5A0Uks8+mlOHcgduOJj0WPiZCoqPcowFuONBuITkU6Kbb/tm9U5Tr+dIXEzj7CK52
jMeXmpSItxWADHN0Rlwuo6qH0MajRgZW/niVl/cyFJVGjANdpcpmU5/KGragfgvwokoj2Jk/TWP0
w/TmBSEeR0v9mxg63ekHSPot0JmRfiFO0j+Y67DyBkMfa/Cu4/4J+zf6/OVr7NQxmW7pe8SyZAQs
jLKC9ixA0PtnTmt//zdmcvhzI+P9l1VdWwx7HAuKjmqGnN6iQqLR00X4Fq61EUhUdzYcnaXdJhqH
oY+Z85yuKeZm41htVllkqfkaEMhhT4Db6jG7NpqERun51je9HgyewCGPo7JhV4/+H9jd7gxVYAau
SOtY5gUNgV1ijPQ=
`protect end_protected
