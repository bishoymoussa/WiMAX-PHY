-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
YYL0Xgpf/AwDCs2/eRoGkyL+rPZAZw/holtIdtCmtuUcQvQBLtOZRJ0knxYpNlzV1k3h8NaMfK1m
dA3ak6xKjYsHsrEjg2hklj5SkJnlerqkZRN4Ezq0lVAIVIdT3F+rqIm2cQq7/fpP6NZdiN8CndZv
KxY8nFfQYHN6HGiIqPXMdYlh9JS5tM5F+EeM77tR4zkcXIpyvtkAMKp9MqgMAMn4PwfM/nnJ0Thj
8Fdoj8JVk2raZim4anPGrmrjwL05gD8DO9AeT0YAX2lnFVjDj3tS0iV4/iXCqqDr7P1wqPi4a5PM
4SFo1bPd5by7hQy6kpAg1WcC4n97goCvm5KO9w==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 8544)
`protect data_block
z3+qQgUBu4KyQGefBfdgvG2zpoW2MUSbhq/QMldIpfqfnU2+elWzwh1OZF7KxuTRfMIFZ1KuNzre
WUk1W8s9pGvu8yktUS5jIqrFAaocvO80VEVZ+qid6aI9dlgL87TzuACECLR7osKw2pwwQQyH9H8M
T44Wk5PZozayIlTiV4OnAalTU21GAquvr0iF+THXmfxVo2GAPP/eyFAR9CTcu8vX4Oe1S/0270p5
Tpok/87nKTRxouoyUivxJqWlz062CiP0voOzWw3cx7zH+sxJ5CSLkfKJP3d52JiOH/ShvYXWpVSS
o2rn9S+JJk7rxHtHct9WwjdknUiiXoCuwjK3oqq6EBxB+SnKBTPhDFju3ksV/sbG75EaAm8jCJ8k
eAvvvvsO+DPEB8cn7B2JOV25GS20mL5fs7JWdJ9mqqsDd6aj7JTMSbRSQZI69GtEKVmAq4RiplFm
5Tta59BI0hc1i80VtE2nv/L/fD5tKP7/zpDtV/w05fCaI4P6GHRjjWWw/KpFlm3FYwMfxeXhWr90
6QTyiA+6otGirnk15GtWpnunSo0irfuRh5N/FHIybLpwaqEQhhZ3sCsOxxmFIWDljh9a6moHjYvW
5JgKcWE7oXY771YEmTwwFt3rWiGje+HplYhZtMfz9ghIkL+5ylXXbTNDLFAw6E5Dw4o1m48hy3vj
Xul1SSFwxo0hz9Ce9lOXRBz6V6WZ+AAa9HAWKnW7kdOpct5j44oA9znweQOhPXgIqZqWrywi46AD
5NVhHWdYmpEG8QtEDtyOlbazdP0l86ssGt2mZRyAPq75E9mjApDQcF7RVigW9KRf4W0ai0HocP73
6Rl0Fxz3KCDs6tLWlRdm+IQedHOLGZbWPnMzSOAydRE0n9v/F/1q3QZa55S2dzVw3sOLjrzPFuon
emt54mIr2QrSz4Pkr8hseQ/YyCf9QXDVVOyFY80jowErPpzmG6+1up0FZzM4jqCOwL2jL8Sy9Ttm
ODGsfccfw1zr9g+y+kZj12mU1eBWv1qQnWlOlwkoopDzLKyKre5P+jeZ/tzQHnvzBXOxhepTZIJ+
prCl5rOEzSs/XpMetFaJXyEVu7HFIvhwMhW9Z7lzRYq63ItqDJXqT0ziUMUYa3zn+eQMmDQ4zNrm
V2iFAuEGMRFK98OQvYKvxEuSTCXavc2GVUblI18C2DdtRkGu8XZ1r/Y8eo5LKjBwe9cxBOUbalim
pKqMDhBlC/4ZJ+1URGZTvr+DHULL5Xeem/4Jnak1eq3DkCY3yapKin8ACsBBsz9a/OaFw7LTj9gw
HmQmx62ZwZkTOhNGrt0BJfvIavO5/VrgrQhl7HxZ5ilIhD4Wagy+u39qvP6ixpEXfgxU7BsqfnWa
VAb0KF6cfsVjdkiZ0d1V+50mAqSOtN6jAN8Qjg/BD+x0NSBB7Bkuwcp49gqXRVt/Kd6KMZBWDNg3
Oj4idwJq+7T4wu3t7KDUGCUz/icBdgX7ayjYxy1WlUmChJUsbsEErwRAMSj2VcMXL02oxikrWHiC
moK4uHImZYp9XF5FHqhkUheAhj0f5iEe/zXFxvv0t6f5VZ0gAg9+TK9OUWpyjx3tcW+9UEekB5GO
KVH1BcyOuvz+YAojshN+k2idID+mWldaW9+aH4f1qAMR+XxlfmfXDRv8Aeck4A+lZ3hY6UCMxGp6
kRA8qYmfQRAj3vUMDEsraoeNyoR6yJXlFZK0WbT96Z0lXawLaGIA0rj52R9CYOF6qfcoDkIheopa
z1JvbHUV8J6ONitPvvUDD46jq+2HDT5oBzSmTFm5HNBPXYZ+rZBIEPpOkmSgw96R0x3nVd07+qwL
BNPOPkqk2Qxzp0Ziq0sBs0p5WfifEPVhD7ZoA0jkmdxu79ANI4cwICaFO7GC6wQ1e+K4S/IXCzVd
62krRo+9Q+jPEysLIlntwMftV71KGRQ8dnsvd/56YRdfXCUS14JlU0Uw+HmdMK0ySstvZJImNYbX
RRXCvtluUush5JIaUj68vPyoRr1T85ogW5sknXpg6e1mWka69BX98KmhxBeOkXgrc32VYiVo2jO+
RY1qj4FK0udS7Q4Gs2rXQ7cD+A14BgzGf1T8+em70d1zqo7buO+yW6PDblyGS2BrNgixofLw50p3
P8rJo7pLQxr5skHPHcZqAbox+4cL6lqYdMXlx3qUcSwz67D4Iym4LgnGaopiwt9xtq+ezuo8w3qb
fpYW+ucLS6fWsrH/QwcNw9bOK/S//oSczLLqG47nEEUDoax5/o+ZOYGRU6qVXoaQYi/cOhaFS1Ak
579q6vDcTRVBfAODqL2XWeMm9tZk7XaFXJB/zbmHkj2h1wZPgDxha7PMXFMB6RfDMkyvqOXH2tez
I7VGoXttZ502ZHw+HI4/Uf0RHx8/BcCVDFQjCNK72ri+m1x/adGnRfzHA7a9cu43EMMFml3IJd1s
m+sKsHfuO8LjeTfejElfTxKNTXVQRfLQ/OGhYFL+TEWBYoa/6+Yhf3ubmDUVYlTXJJMEcT5YTipB
qWvcZtNtbFPzFELQfwnqXqPrbxm3AiKQiWR4B5AfvXWJ6hsVQBs53HeGXkxBzmBSGDA0e02if9X1
J2kqHine43XdYGoX6pO/yoEqFewnUYbb154Pz290aF9kqtBd/jRBBBr+f57VhA7CCScCEwgBBGFz
tuqJGMgk1codOdchy9IFnvOfeWqGXRLYRNR2u2zVfoSeN6jAnVJZogkN0NANeBViUiy0ZwFxZ/Sp
ygCPpwYUwDUgVa2N4XyxaPPt7gO5eQTTPAh9P0qGE8yQgngqYx3PD4zf4/OvRmWVCXkHVMuLF6ID
KXikXSsmZLebORIx/fYwW+C3mpEbqnVhX00DxnFhQwIcmnXv2OvIp/az1bV89eLuNGSRAC1oa7rS
VYM5NVcwxI55q34ROLEI5LZi7G1jbaQnHZyfkMyag6NXd6eO4AV+6Emwm0KZQ7M7OlLPcR3neqxQ
uoEb6EJ9820+l5spPrlT4ZoO1isozcbXMLzTIWoFMezh48ZlW8DMOgVwGGDbkVUcvSUEF5AHZPMg
LQF+4UpNa9VUVOnbhTJ93vX0DEB0pzkiHEr7Vj/qKR2kTGCTUu1WXD1kOyovmaM17UVTgd3IYT6Q
RITIf8V5QxwCXezJcmmFwsjsxmeEOZkYffHLmocqOdRoSLo8lIHRKUWfYPZ48uJnOz2BBNNPfXu0
kPS4QqaTg3IWbyG5gyOtbHRxnhSLkzZZBS7Um4EqFtS1k6zqltjSwJ85MPOTSfnxLnvUMvM7+L0s
Uc49kO/5Cva12APj0cifWg0XAg/SCbBGDYfmtfcbWsnCBmzyiOOQ+7rALit4Kes0krSN0fcg0XHd
VZCbt6Gd0s0IvzPTaMxn69lB7vau2rc4A0UUJPlR+xKcoU0oAohmPwYrnZ6LM4wTkOsyDRZXPaTi
22Jqmu69vIOsZ3I7ebGsYQee7B4fOfeHhnBE7W3u85aAxapbypAwRkV/9q1b7XGNP/wwX/jgpf9K
PbN3wGtBnoUMfcg0MtK+WSHG269Dye+SvZZWiJz/v0m4LlVp0JYK+138D3sNbvUlT7NWLFFnQsPQ
LyZCvSSMVN0kieTy2RwhwcRdEpQ2Cl53A6G9LpC6UHVxA81FaWXGYfSLLTHW9wOa9yPZ9AznK3Ts
L2HentNfPSjWYq80Z1sEVdtBa84I2ibErWmTSVDQXh8aWwm4wXaZTsVjCkjc2fM6KZtO32pAI/lP
HdhZ99jpV2SYaTfQRS6kM+QSafyxoJ/4+DgPsXUASYj1ix+YVGI/jPwd3N82yP+l759IExeEklNr
IZTzHfisODLvT5vRk+yDdD7cuW1gP7/VqhsVESm8L8F1UvuszlV0T5RAo5adfRVU0FDnQOsxMX4I
+UgksPXlsf4YO4WJJjcqocSZiIfRV7MyLPji4j1BQntb1ZtGRTILL+AMrPEbACU3G9MlCeIV8WYz
keK4ZRHF3Z4FsE4QBg/BnbDzREMhwI4IhXp3OSJYKmiQug8sWGIAoVHe9ICNkZpKjy7e8+aayLNN
6ggaXnG97K8MCNk7jTsfH3S8m+lgXYfkh0xps+EaCq9tchwTJuC8wHl+QZ9gEoQLO8OR3Y3XIV+3
pBhiC7cQNJ4qhYHjlbSqX2dvE9GJ0tVwldvRc4neYf2/Y/Xot0OWHOIisOAGqgxUl9lX/Irj8h9C
eQqim6elcU7P1R189uVrdx80AOAt2zmIvSAuIE63NM+EyW3Fwt0zvZVPmVRtz8ThG00U26YqghQV
dGDcgFfdrN1Epoy+LC+OAk1LHU5FtMwSAOlDvNvjGvv9/XSpk3/xJqqqa/gLCNojUl3wTETPwnck
iSliDX11na5c0k8plAjmg4PlKYN3NqHr4CeQmtdY7orPMkqzAlEYDPkUpBc7MTI1jnC4hcXrtcHN
JbKCLQPbNe6JcGtjQqDakqdrcNzv3RTuVto5yFEleRvSWLn2obM9a5anh2m4Tw+IB6rPUkTl3J1g
Af30ro2MMM3XTwPmI0yLeMOZ4hUTg80YTdWO+8fzSS0PA0iQ6rIRux1aptvtWPfT1rUWm8NertUB
TARCJEw1NKDDmVEl1ic1dQj6nPxL3XlVXiqAlpEXSKoTE7otOftXg7PO+aUqIG2GbtW7amETYXx5
ScqcYkPEwbs0vT1eQxIn6j2bsr7/LMP/c3Hvjc4o8ueRnTnIqB5MMnOO9qGorPlYWoOkkFyA+QCz
/xIXxNDlUZG5n1QZNZI57P5HB4er9TC3C+bQw4EzZMmGPS5Gc4OnOwYwPfkITmxoW0cxzNH16yrd
8btyc4UhjvBD0eEr0d3EIpl4nDJb8Z5mtbR1M4DoqNbSRuqyf1OYWiU4JW4dufuHeE6Ew6cwfxlw
zaVo5Y5H6NEDgOJRWpcMiMHVpY4ZwTim5RnaMgqBLfdUSg7YsqnCKWIi7NZ1p7YShy5KtzW16b0i
zfrUxXEVn4BNUGW4lIwORtHjWxSnKZTK2akOQCUO8FIbYG1gh7hVCQ+nawIxcvmTVbpQBm5XgSRb
596wuKcnn804lVx7gstnMMLxvFsPvBlKaTLi/heFMeOWB031bvE/y4qfW3xKtU+E0uZwnaA3uU3b
ByC8WbRRLTaK5Pj95JhHgRd7Zw8EpUeiuauuqitkmxNhJFcASD01M6CNn6lg/khUZzm1kmH3a5Bq
hnrGBhSCEg2Ns9aoWWMRPvNI+yjgWSfbp4YLj3u2CodRI4KJvDUgkCm7xOyevQuqROBqOWxOklW6
OuyYxWPLFnHOrE+0pMoZy4rEc3kuApYOV9uSX85+qdnRjY2eOoMy6+pmV1zAx029L7P3n60L/le0
tHgUf1ltkcy17FvZhsJzbTBwEjtt+DouJbXH4FYqpgDD/3+sPsfPXXVsmBaNm2zqAw0z/FVqyikj
vuCTuLhSPc6BF1L5UZdS5B94OrhQjMo7FJHE7L+wO2UozfonFWaolklWCccFm8lBpvpcDuUDqUfx
viln4dH6KA9Q6y7hgEYcymFqx3uEEnY4wPk24QUf7qN7DWmK2GH50erNJYds2GdBl48frDaLMTDj
WXN9MOoCay/6qJyul4sxSN8IfEdjCvsJnID0H0SS8rGHpc5xxf3+u3yQKIVlw3GmGYX6NAT3xvMP
zlCxRey+Q/qXso0Ws7eKL4y3fmng6pHvMPt3DnaymMV3IAN2E2tEva4LDemUAN/60s+DlGTNbMMN
TGhA12Mp6KpllTcy9QKjbo1YiRnWLg9j4v+SZ5Avc1UVnImT4zg2Am395RhakQzflKKl0zpoy9Ur
uov2pjbXUaF9Ggi261qBnKMxcJtWfH5dX27cBupdKBxaQm40PC/7e34qlg2AmzjuLU1f4diKBWmi
y7fN+i37WiHEdx7KsluMPU0isQG+uTm8+0e8SXdDJoeBPzcwjbGmpSgcxCu+mt1u2QQ2klqUUTz9
aAZ5HM8903UC8kmyb81gl/oBxbbpTGzHDxtSzNBBNKZQGEjrS4Hp5SS234rQ8vZpbaT9qFyWb7lM
x6PCxOh86Pk9Kq2ZIbV5i/7lY94fvVRapXdF8BWHTrl8EJQoypRsdevDJ07AXRZBtouFh96r29MD
hktnkXcwVbTvnCJlwl2XWlykS9Gi2s4sJVVCfaiJRxi53FJyBMe8Z0xsodp3mTzDBLE/jd+Hk1FR
gYxdhgPq1SGIz1lf7CRvABKoVyj93EoOZNLyLtasS5+6AzjkVx9AsMHuH64c0NM1DlrA4rxAF733
giuXCtQoxmAKeXyXjOxbBgeMy3bz7GtPYT2Bvl8SPr2h+cgF/rEWOhwfzPM6R9+nweIB+4cLE0Tg
i4ua5MvJDtf8YPI40AcIvJxV7noSQFfbsokhLjVRQrtww9mrNYqE9cRSrkDUC8fOyFkGuwmyFZ9p
08OkJhpCtuiyaJEONDFJOHMN6qKLwRMoPmgcXCxfHpxPFy3gDjroBbn0DGcXB7w8wmuwcuBymiBd
WA7hpt9nCzZHYxm1hVLJ3IZwwRiGxUXMOUkUF4GoGgf5km76B5cUJ1MhZnx9hqJqZcX1BBPe7TcY
Tcu5/geUVIHRWqciyVPRmJ6EqbYLKRQMJ2riyHxqpS39ADI7VXeIrBXB4o0ePVoX6oblDFzv2s65
FxzRs9Z3yR04QaMYDQrYXfGiP/UJuIFO1ikk7m3mK1dG3N2+AFCDNo6dEYiJhgtTsxLMgErewI0H
i12z8mXibR2SOAjYMdpsOrTpaxDDohfLCxXgD0YQsYKmS3nrFYPhJ9BHHHOalzq6ioQuAWQrvpkX
VbaCkBrd/WsXHDCODv2tSS3pS84VLrAD7Cx7Y14KQKZmIUWEnmLm1/NTfde9k1meIsyUmdgQjXvT
4dFBoXKN2SMbQ8bokLclau78+zqZan290fL5vEwjjaPUIMCJHao5ihFFFKCJEO3mfzT8+z02HKIl
8macAG8HJY0sSxmf1esAKEzIg0MdrqITAOJVcEiOoxFaekVaJIW8NjsHggOro24TMvhxijILIJmE
k5LJm+8DsYvwKuGWx//lE3up77a40afO1y6TZI0YeWsupeUsXoHMoDVxkB8dSnXz0xhjrWFJBoiF
fj6VojM5LZfLtOWquw3E8F0J9eSNpkamUz7iiqxlNSg/fUM8ZSqMoxoVnLboT7b2YiCqd/3vGhYn
Gg4tw4hK1ri9gycGFyxPzRySClnvJ0rRlbiCivU8U+XsaAGBDb1KFDDU20zv1ED4pvmTocIdlnKZ
SN4ddHeI7XqdfQOYomTUIrb6vdb+j9BrPwASbx26PBA1qz0UBYJG6Taut/kh7JTPc4tfITNK67U/
YmjAungB6Za4WDJpKRdU3A5h2fkOwznqj5U4gELxMTrS4WfGeQ1j6CPvIg9Q69bb4pVuYwjnvmAt
IXasg0MDZlKekGFPlFOhOlcuhQkT6aiXprd2Y369lsDL/TCrbWNU4GBrKxLkMTUsujBIHaKdts8z
s5bo0gkjV00SdQuZzp+x3ZiYJV2dHLNK8nfssnA/htGvD9ebZwpW87F0BPmTYBAwgtwOuxc+Rfni
6jv2dpMPAqyexDtzhMZ9nhVcSEhIfvhDAUTqtjlZPCbVW/yhh3MBXxPu+oLZaf6SPjY8poheyID8
PQc3IKqcu4KULOPIFkrnY7BnEvlBDqDAx7/+YAY4l9JgmWvQ0d1G+NIZs+lZgOBf2xem9DRkZe8O
eAsp3P15lmnYS+bcWqoNbESDDTno9vmEECrFLbUnoPA9rTbH2Exd1ca5H09OGT3GOdpYbsC8B23y
vk1OwJwQiFqKr8sG1rvQgcLnZ5w7ca7vIWmXpSCaukcsuAplMIZY9k87yYxV84ClIo4EKCIkRtjd
J9FzOksDkV74zkqSAzDa7EsZTm/1beTdUvcwt3WGnSCod77xcLRwI97flkXVmNdrMagL9lm/I6+2
y3BL5xsXeWv8YPJMIPi1NoxOeVhDGbLO9IIxmEe6Q9gvkXxD/0rd9gSqleIPNjOX5afBhXC0Mjxu
OlBWcT/uLM9qTqrI6ZLMQuSGC5n08glP4cbkIRw6TVIQU430oCC/ad5Dph5CfI1uvKkFBPaO3yqK
TNwZTaiHarFMZZ+QgA3qNT/SCyFPRCb2EsJAThszorhRCKFtVXuTfUBPBwn9Ba/TYn8e/ABt3/2b
uhFl+LBqgsRYJlS71tv+9ydL8uocpkPpvMmJKJv3tGRMTocfh470Gcoia+ToXTU1heQPrcLN5f3e
vrmkVlsCJOl9d8ZruKrhMzGBru8J3RyiFfoiQ47W8F9JAnZvKq3y9nAi2fqK3ehkmfoT4omJzBPc
qZwsoJoVhOwe49wxhvjZ7jcz6WD/jA6TuLdeaYQG+PkkjaBotH/c136M/hGyn0jiS6kZeEnKEtQD
f2i5bnNLnakIrPQcJZ0YtrxnPypN327ZiIgxojSQQ3QDSzhCQ9cUQn/FSdag7ktbg7/SYpLhDWPc
LlVObRqTMST4Q42RMrJkUBmWTindCYBAX67+dHlyQERssIkKLZhgU+tDeZ3txIjZq5zaDge8GYZN
GQbLFvW9Is1XzzvY7tDGPn53xW85Wp/IkC74KC0GE0uyIQzErcG/8InBZpXnfFcBvUycpZ0Hb0kk
5UY2VqxI1hgCesoqJEvncgQdNjF8V3PpdbU1u4pxmakyFxiDrM+JwPwkn3X/mCL/sNBQuW9gYUiI
dipySM52NRuTTrXLcW/jnfa13840icAfltUdiu79iAd/21ph8CqNR6LjmEyCF+ZAgmn4CLQIX05t
OOS3/OltDZ+dlzT7S5xlaX0df8agGkByzmY8UUiN6TW83Bnc56G/nbLMybi4F0nYOI2LHsrbnDRu
EnVXSMRflxXjh2v7bXucb8stGTFKyv94mXb79VPd536YwkWqnuPNIFGkSywjC7C6wfuWOLlvHRcf
fNU7vY13QJfbivqeuHJRj2tQZibQ7XqUbQPdSeQtcKNlAZSOnr15Tmwd/xa6sCWud/0aSZ/lr27z
TMiEbUTRRn8cRN4jYmYp66QswbRIL7RsqhWUVHUyeLp95vvGX/F1VTbX8hLdrA9+GLhx7yAgznfY
WSqHYl0EZVC27VCHsKBJQ7SY/ALcsF5CDXMwwLDv+z2TWRn+Za7hvEyvoiiyanvDacATpHTeFV9L
K//2MA3cDH6GixrdgwFMQnRlh+ux8N7zUiMDjbXwrOIMV11JybfdVkDAGezJ+nfBfidDmM4Qp+dp
q4m1KwtraOkvPYrSKiFu26YfHeG1DIa8PNjndJ5r03yK+ENpwiHm/b8VqfzPyEk4k1scRWTRTgQF
rDFqNF64OdxeNgi5DlpWNaWIcJ5h9GWciTz0lNmSxiI0iIBWFdF4TkcDxTslhngFejJBTN+QPHpY
A1r4VxGNKjxp7B/2E/Qkjq24/sBHNktzBE8tDvw7NB1vA5dgpEzfWpEKepX8RCXuRBFyP3UyktrO
S5T91xt60Jn/WbAPa1ZxVckESj6uMHVcgDIqPZWKP9eDCdMHU6deOKoHFQRcpSD95VfkFGiB/AQ/
igD2DhLLmiCSKLUnb67nGwg0W8CD8oGCUZYLknE0iA9VfT/B9V2VnPA5QYlq33GBCy0pyrIx7o7j
Fm2z5IUf7vi/FoMHwPcCMAzvjV1XM5gNnLa0koAHqNPYLnvv9gNV7VO53kbt2eM75O8Za1fcj65e
uhc5KLsSrNe8U9GT63+6EiGIFTx4DClyv/1XekBU5Us3lihBucOYKMh2ilMZOwBqzaD8V2ql3tJ9
mCkvPALpRjOJGzMqUSTtorsPS8dYldEfXE/sX+4ywCSh1bRkYq67HfxvHV1v38pP7A5Zhi4P6Wr6
2i5WbjSfS+4azoGk1Kpzdy4+r7A4j+YuaLWeOUlzo5XewSU+dE7HGbg6RRHXO8xD+UMbkIwu2/+q
EPoLUgyxUQu+6Hx/mgq11abqnzv6IU0BCmqfxb+gBT8yR+KRXmDYNTJCZSHMtfBtQr8g8j4+fX1l
3eaija1sPSfobaG7lHEPSPX4tUskrSkhyUNtxjlKcm4S25RxHbNhoydxjWETQgzs83lSIWAyXKBe
mmkQ13I1/51uWywnhcytT7hypJxzzEavj73X7VBrgGUPeSNOzj1kppchyAWRfubuENGZCmYsxKtx
r/Pg2o3UwBCLl2pp+aDHzPgtRH2EPs8soTwC6FHBemQcIGzeYpIi8rue34jQ9V1iVO0j4zO3jNNY
B/u60pmpX33sNgqZLK6WUNjl2aLVIP/Z3Eb5Xy5Rra8dTxxPv+zFc8YlPJM0i9rB6IBouW6SXK2O
SkvfcxNG6B4HGkC8oUvbKfkHLAcT2m4ZZq8p9JjOVsPKDwbgGRvPLATQr1+yrLYlcv9DXbA+iCaJ
1z/DxY0riX4imFx1ZayzmOuNzFG2O2r3tDRVEPMY3nZEWAq4I8fneOHRhv/mpv4Kpl+U3Qrtfm8E
wMAjmPQmt0ig53y0k7xyxbq+m7oh/rYOfwIUrVoJdgrxinaF3qDJo0KUN4xzK2Zja5I36/hJUY5d
SSoDTLLmk4W6Ej+HQ4W4uo7xje86RaQ0APzaxBguNeYOn9cYtWZ/mgrCHd4o1o6V+RhKfxRiSmCB
3mxtCof8sww8VvZH/Japxx8kyUZ75HZwcf813Do5+0qkAJ7viJMtl8cKpoWEzwfIOIdmoO2xBvPt
1i5RyCB9p/ORji4MHwUw3/h5QUwW+fgb8sknz85BSvJNaHJ37EejPqYzYbi218lhEwn6RkOpR8em
RgiovqhluMD4Yo43F3izZm9ZQQLTBvOGAcVs+HEMektE5cir9BWqryTDXrBPEYg17IytcYTXhdYV
pFDF6kaNOWQREwlhqin4JwS2HATd9ZzQr0ubpj8Q5zdWelYD8WTpyOLoE7oJbeXGEw+psBe73jp9
ptPFHLqDeVqVDpDCcI4Gh7di0mbar+KdQhS7ovWERfoertMT3z7EYuvl8UULMlFLJA4eO7vxTmjm
ZZ3gccFnIR/KPstmOeAKgyfaAa0TZNI8G3pDIpp94WDCrwe8YSLzthNh8yaP9mbl3HMCoOn6Esux
QfiSGZsNpfh+GfOIyvUQ1bvcEZpGHwkcxaDA3QSXBes6cba1t4KKrxwPxi1wPjYxoM8amuEXbN4+
qojQOFupBY4o9NtyZGvqQc6QVXAZaRo3mDuh4V4Wq1u9aQcyQu8Ci/pux5tCqrfR115yp+Zr70ua
DMcBfQY5ygZRLqKZPT6QDmjtc3smJgozR+AVEzF8SZ3IbFlMJ0AgNgmfkaYji+5ul53Ex5pHxTLI
6Al5gUvioqtxXYU6gPct360jVeBni3/N7zm0j1y5HcccktFxpTyKikJkdafRXAJvULD6N9eWjC3Q
33X3wEXzT5WsCAxrtKg47ANRX0EG583YGgSxxEQg48s7JRywF4aA+nPMBxrU5uicWZW6
`protect end_protected
