-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
YAb5+q4bHu97E36BuhrmUwALQAdA72hiUkHjUk5TCJtUJCKAaqVvNDBt2Cc36O15zumrZic2efUx
y5ASk38r2U1IaXudDUTOVnwDc36EgO7hcGixiRFkNU858RYByhZvzQImIyu2VrhxbRhNNxKScTep
vRI36URIrbCQL3k2uox/HCxi2aGg4chPCRHlsvf9SclQIXThoQ4EDC1Bg4+zv4Z8sZqucbEfi4MH
b2ZGravG4Nbcr/DtbA9uuqCqubvEbOnl5hIBtJNGI8IBL2hWr2SRio0pKOPWU7dfHdEpiu2bQ3B/
RIm1mheZ+mBXYDt90WVj+QaE+cU+h3tNHeknvQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 12960)
`protect data_block
icRdmrzqOBISNjVyw7kcy76LiPR7H3swmcw1nKmu3Tns0BJgTZhG1wUAkW+DrxrHm1Ho5BYgjmn1
nai99gw3biNsMIDBXvu6cVNa6ho/eEAgeeojlh3H+u8u/c3VZt9/eTq3zmxnvalK/Lkh1Smkb73l
eOcIB7jEknRy1q8IGAAQeiy9/pxZ6st8a0J75zDWhRtdF1zMRJxaMY5VC0HzvAVh7ieThJztotIk
bfiC0iGfPdH+geO2qLRH+TpGeqpOQGuZG+OsDPANwv6GTU4OhF1fuSNl8nRhY4BaJfsB8VNpmA9W
STPTMPRJ7BYA1IAh7HmxPnBji44Hb/htMbJ9v1ndxBQCVze+WYNBdMD624VQrGJnbePq5mev9LOq
ROA49K8GsSc/MX/74wIqIQqc3yZ2l4v/+A3Vo5KMJrb7TAVigEYPSkDbzk/jPnGtzMrLhO4JOuX1
3sj3BvsRC3bJBDErhJeVA2iK7/My1fzfPHSAvlnwj3oEOdpT0TaazyvtjouOD1zRKIig4rwy2apL
+vwmssYwzSqs2ryJBl5IcdmF4fbGtmVD+Z8hmPAJXwxp/wSLVLAHAsVXGBuzpnNoWQpDStIWfpht
wC+UqR5dwoaP4938uVkRN3Z3fEFjZhkPjB2h8Zr0g/tesys4ottgQGi/ij2Mr0bT4dXOBOAZztPP
xjYgVCMZcuAz+/hrqTGfigeqaf/5R0JnTJer91XMagYTmUGLN+1WuvRKHk+aZZLJDPUdxRf2XdqA
dMV8ZeRaFbwXFh2bja349emPdAHauBjQDvryYiCQBVyLndDFP/HdsAFCdbY1fsLbR6qK/bJmFodK
68qnPsPD8ktMnsMeCsdtZ6u+C4rJXnPr7FbtjV/uLoHyVwueeB8OtdcmEYPhytLj0Mf4x0JTlIGL
4Rvk7YI6KkkcmpXaaV2t0mHRiDwXi8l3rkk0GKT/vb9oWmvZ6YrIZqToOFTZWnJ6E+tAwQQ42VAo
OFYtLcrQrm9osaN8KtHQUx1wQyManGLeCCuGG9XRyNKlnlY/BvmaphYLrTUl8zroBddebCQCqm6v
68Z7cWbtrnSHoaawPSvqOXzPWEOIkO/n2YEJLZQgUsfzKHWFwBjD2tQSS0IwwUOIqnicWeLf9pyd
j7487NUEhAwk91/pPtNW0GoUzYXR0AGQM0ENQjlOWn730ONpPgtFnA7iJHuVqGH4YiOcFkKdTdLX
tJxAdMkeefl/aRnYDV51n7YoYAZLXcq2kXehdpMnnAewaiLi4qGyPdjErlvFHwr8kZp7QD7p/SFw
YlfVQlMP/L1XWVdoaV7bLiK5mAuKHw19a7s5L+9lmXUE6RhlrEFQ5Ye6g0J84PNLo3BFdxPLGZBF
RmNVBkOlOvM4l3d3iujNmmLEuCpeR0xrer7M0s6GxPtsU4/nBdEVVHyypGvBWeHGgaeQhQpCVuRa
6KpR1UeiUcVEf/HK6ykSdYRu+kwc7RKM9tEWFwvSY/iFoZqiAVF3Ej8bXnDdMYYrodu1+sQYMVoQ
YhSzApaXtsDFQ7+Z8masJOQ2QANyytTZU5MTPzIVN57zkoR1J6asmifwzVgPCSXMUCh6NSM/qhtt
BRZby3X1jdJ+0A2lEVpkzFv2n6b3QrxhvuSw+qhj9H4ngEyZyJQeTHYzFPVV2sE0dlxH9tuu1RKQ
8Pqn0avPBa5+9KeE/m7vcafYNGLZTc35nt0mg7Kt8+hLJaKdXqn1ntlND/B0dIyBXMNsGmOKzef3
Eab1vfce3/ldtJdeYK+oIOAFrwl5rVGg5syYKQ483Lrg/0hs456FhF+Pl4BYR8Eoi9atmgP7D5zD
eySAiKVxmTxhrLvGpJq3qLKCZrgjlJpdNAZnNtfgbTBUrTWFEBJBOwUtPmouwlSY3DFVqKia0rt8
W8vUJTpJ68onLCwuwgbSjf8OXC1PpkWtccS8TQ+MATpJPYUqy/tDu5ubCJEzRulv/xIDritze3q7
e+n5GCeL4POT35/eclwBrw/UB92dO0gXOsB5xkWNbkDE/rqJIG6Fgigqig34l0GTwnjFaiAy/u0j
aQiyEEATZ9aCfSZsiAVDyftpBXITitQ47OvZvJwRqGBxdFjfDPI32w/Ig7iW3R0JXCfAfiVqZgS9
8mLL3yLxONwJdBh+Wm6qNVOW9XtC7wuntLtwVrS8s6O+DGxBV2qEKYtwPf904gB448McUbbgiUYX
J6FDhHPOfinl4bMB8DBAe0nvJUmjfgW2xstMgarbhT4t4VQ9PczH53xwNHZufCNY5Sm6ZSyFlmue
WJ+WYLG28JvlYPiZ3bkTSjw4Ggna2YnFlqyLYrBWJLzhpC9yOmSZHaxgVxeXwrSNPmMiXx2+lEet
qqEs4n/q/MeRep7WVGqOIfUKbQ6AzIf96Wqru0Uym/DemUOBkAVZ6jP508IpBvxrOfG98N2y22Fa
Zq+bDelA7v1d9qTwQ/EdNSCsuRHaWZyVrJCb6R3GaPvG5rkCtcur5S1SpGBY0JynWxuQmUnWSFLm
M9P0OQ+pnI17r5Cvs4A0APtoFvrbu5qDhFS7kzVfARj6P2tfl+DiUFg6cUxJqrveJav0gUd3A1ii
54QEGoCZdi9j6LjrunzwG1PrLCI3C+Xgcpnz8wFFpnorVEoIE1RF40oywLfTU55eCo5UP9EyHKjn
cKB1D2S1HkCnTBw0Ol++cVbjoeMYPbxXpEDscXr9AtGw68srNE4P553C8LX6UkqAzNCox1zZTz0V
buY7+f3+0pnN1Y7iMsc8soQ7xMhoWcHOmrITXVA9YSoczsTP/h1aQXU/CZmYodp7LIoEmDOCuhIp
vIoiS3VO6sep6f/m+4SgLBtQ2E91lVFVvd1tc0zR/xWKtc/+NmdFjIzLfSU5+ZbOBqZsEeUTPzCJ
P16c5olkfr8c3KkzQhdMdHkUVy0XBUx6IzlOb1ZVO0ddiYnCvV/P/wJTBq6AEYXxJHwiDYDi6Fz/
qU5cF4NilPhD+eX5Gyt8F+3VFZBJfgsftmrQqi4GeS21ybXCg/a2Lohhd5vp11fF+YqUQ3VJnctd
xIuCQPVbM2RsLTmCiypl/2Zw2dbeoiU1cQ5fA65zZIbvNLX9QNMADqDrVfQe1TAi2ZrQ3QfpkjWC
NCt0A7s7/aDk550LKygg+8l6PXmNKHpei3mBgFhrUbzJjGLBFArPZoMdf0lXU81pHSINwNwa1f6d
+VsR9C1017VphTq7IXNTZBazQK5v6GF4csee8HeVFP+Gc8RNgyiAtpTunEZa89ytl9749qKnMZtK
7sABB5A2rtpMzYkS4bHSblWPGuv2dqB+KF5dhI62xFAk8IIUV7Jy9Y0qRPUp+y/EOWLtZnuDnYrD
TWuBpDKB5S7RoZggoQqJTx91UGwxyNXI6aolwfddm1O+RJXgL8auTBXH8p8VeGsfGaeISeToPklL
L9VizBjzDwueSGtLNrIwHGP8+CYQOHmkcdHt27EPztbQXkVBf1V9m/wrWDcFCHhp30YAFUWFdoA+
h1MgmrdvCvY40D94oI13xVMNTQtuFkfF+6HUH9YC1T0ThR0hXMsZksF+15P4BBOtcQMf64vcAWiW
CH4LWuM8luwAEh5nnZLwNrgrugl1GFNoq5pXbFl1PoHSSgu9XdmwIHWq9coPhQ5cNCL0MIXHPvoW
jIzYX+cu/1DkQ7+aGXpTwP5kkTB3o+Kg/DRlhjaDw53kD7a9waeVfEMAxilC9wLTSSNLPIakXQ8z
+ougzKLq6WPykDjAEya6rHBS3njTmVmGKq0hk+II6LPS3CjwDpHvoyV8wkVxCCXAAtmJZNJcQyVH
S9WX0T3U0pDXdj1qWtAHpJILEZWu3q4/1xI+lgkq6hLMfoUMCDsT4tgrUR85QdyoJx2eun4KNjXS
8IlUbIqQTJaq0e56PtKVUJU2GG4a3SyMT+zCcag0Yo9bF+A/E5Bq11b9Eqtth0K5ziRyyWZnfMf8
JG0xlyJ6Zwx3x4VSLwswIvl0zhVgO8+1OF0kI3WzxNuWrRQVEDB6R7E3wfz/14CH1RtJRJbzqq8B
2nb5kwSZuD3z1O/pXre5B6+0IdbKVKyzBy1CsVKTjrQDtBvc7ZRu1CIFvwgXYreFb5+W/nHMrF03
VJBxTPm4FQzNG7exvtsvdNQvJ322lUoRwLAsG8fBKe4qb380++U5qj05QJfAeC1QMUPSOzueJo4m
XlnJA9gt+1xr7Y8eqHGyU0HvqcCJZzjctuHEL4yTVpBv4POxuQcvhgpINg7EY3NVgJyUHdhLe3nD
rgLm6L74RM5TMaBje1deI1+SnynLQpltQeMzQ9coEpnocsW2tS9H7l3R7zrbn5AF0yNgGZUT2hiv
3rtu+yIHH6zZr/wey3fUyoMyTb2264AVuHJEc9z1wgUK0b4KFt2P/5M0K3ZjusdV+J0BCUwEwBTU
noy+hChxODP83eNQmmJshQm7UlbFoxIxl7FCmocLviAPAzrbKVl3plZgtMwege7C6c3KAsE+j16P
/f58URCsT9ExFk1EMOYJm9VKGWndSo+q1y7f/QpGluiIYj2Q6s+42cZv5WNneAFIq533/xjaldNI
1BslZ032zJ1662ZC9/c2yse37RDrC4MK/sz78luXhERxsPuHzWSnbSXttCvj/xHEjqOC3unUhTuo
GvE9LH8CY5smjs7rDujK+zoR7xnOfKjqME2iTWnu8V1wS8f5jTMZgyfBEOa/FWdUXgjQt5QUOwsf
1t4GkscARJZO9sf0eL0DsO2HQ7d3zoYPABETtpIubQj2k5gb7bOFIqjFIuU7G2L3WJKOrHT8eR9o
XlaxMkKgF7TxLP+P6mnGkn6U/+o5oVPIs5w+ZuOYd1tl01GilVK+Nso+XlPWw7v917QYCIyU40EQ
iZsK9bF6km07swvSZ+dU4pbySXTZK+lCo+P0Xtrfu8oOc4Ik7PcImc/3qVmsCqLlJrRwuCtZXxTJ
s3zJMDtdOxeGTuL62XiYXf+y+3urh7x796hER6oKrhGcchOsXs720BRdxz2jXSy22WDnbMF8UuWY
YoyBBjjgY46WBS34AT+Jl/5jrBP0Ey65YOvJX3kej6MRQwV9X2+E83zi1PUdHGdTzgLYFAPbvnea
DMjLoNBK3XPOCvXsQYFWEbWEkDm4IRSH+rE+e+L2HSuVrz+tm4ublvGr4aw/Mm3SSz0lF6qdKlnB
WR/MnoFHnXyc3v5QSvivQWC0dnpaaQY0Mc5vx3NYERVqO4SaLKssbxf2HAx/IlWRSe1lE/kD/BAd
COoH7OdTGUHNpYABNW7zvCnZFP4O2xanVEoJ+wQgmb5PUC8hbef/RoKDkhDeXJL8B1Ti9AyDErdv
0xBZWudA6OXydswA2CS2SMYX0zh0wm2QvWI8R24dob+2w0fQqGY7sOX/E251W7CxTFM1gjBaHUeT
YpEgxKdZ1NqOiowQ+5zFyPJ33NEbphu2CaCdfG0BJdvZwdzHUtxZnk/WC2rZ3mPiWMKVniY9Je5F
V0xK5XUaBFW8rR/m53afX9F0YQWvVkrSKLdbTbeHDFapDBdj16vH5uzODg8yfRjvvYfFo8VNdadX
BKd1shng8mTb8SERsmUjE9IVko11OxSJf3AZBHta9NCgtquve6IMKwNz6V/gOaojP/A0ODrmT7+j
yTunQczmj5pdL27ZLUNaq9JUguF4doHkOXYlQGJOvKyagKnj6N5reJ+N0/0yRX2WfNiGkBHadPRl
SrFhScLegyTU19JS0x0Lu6PJECql5DnYnAkoSMmYInGue9um/kaP0P5cYR4L8KbYPJYAusuRxB4O
NXYY04vylZF/fGZLJx5EAnGI/RzuQstY3czKtcdgh4yZ53mkyBdSWqcJnR+iB8kBlqWprh829vuF
riplXKR49Fvtp+SNzodpZC2lXixiV3k/kOyqY8fKJcXLTw14o5jzVv2ju0NqYtwVWcy5mMRTf9ss
4xY9PlEuUpr+WbhiPLW/nJaEz/yh5VtNNmB1/6ZS9HECHRI9syzAnRCSRVHTcSLGJXLmi9XRb/jg
FS9Ma2fZs5mXOfj7TRjr/WdvBzLGvD0+wsRidSiwCnHuG5XVDdM5ljD5B3jd8xIcP9pWD59cCIac
LyX1jnYGpy5mBdzwHx5hCW8il7dFEypBFUWCHdIcRVl27CKZ4KIvaocckubSFLNTHv/hRJk0mV6p
IjRlylYkP/czjVUdcmLnODXHNXrr1p53jIeqFi3GpqWix0ocZSdznsm1tLvkQcNbNGx+CFVAG6kE
w5HIrp8sForWibkY6zxdnBf04vv2y2RetNUFSciNdLvaXdPoRbPZFt7PNAjh+d9ROzDSyjrQKfXj
WzEKeUjTEdvC6dfM8m7qOlr7JcJzZVbUhVKSJD6KtAZk4mldrvScvRGeyTfjeE9nSKJ3bebVAWvB
fTM1+lGvjYh0sExBKXK4gBUObxb1ZOS8q19aOsfbJwTuttCxbijEYoesK5VOuuAj3WufZmKy4uvh
I70GzHWjidqwd/OcAz+oy5pQRepxzO5k29aciOn6TUxgM+NWC9P/f7xY/dij06ALuMU23E9VnnBY
B7Xuwl4t1hZcEMdKKIRgAa1CHbNOO+Y3fElpK4w8k6BBY4qDwmGGNS9i+pGab/17Fa0tAOS6obyb
IYmpRMaZ8UmfYi5RO/j8tz1+qwBsB/dWYqrh0YhqQgtlSsyvvMWNiCNbpmK8yUH/wkxMtbjKugwT
daAKkBTSBZULlFKRmYVQTomsNkCAoPzA5xg3dO6Z0jKibGJmxUtkB0S9Cp3x/h59Srw4RL+aYW9w
9V9oVO0435SI5fswYap2HAp9Aj/ZUa2yGek7fUZfQuTwi1VAt+iUbxQJRcyl2eLBQtexC4pHBRez
ImB4ggzq2QP2rPLgNmgE1wO6moWe44Yy2B36ofuYeQjgm/N1psM41zkhUq4jeLL2zmeqI9fI4gPf
cm+LTkZeWy4MS9eN9UwtWN20VKMDL51PafMLM3n0crzIrdqYrrUms+7HZBECd33mNeCaTs2n9/wI
NZVaLEsSgpQEMTGbiY3Zkh6ny5AvKNQDEraDTQQGuRIzbNwkk9M/6VJ0Sv0NQI/GfqVtmL4zU4+o
A49SxEzyWBEMXGFV4uJTyfWYcnPKSbEOZzEq1BZH4qe0YyNe7uuGfm8pgbWWKxY6woTI0hk9eZ2r
POrxpY21Z2WKCUEBnlV0H9P3bSIiIMiSvTOXBeLNbsUdFYX0uzLv4ECa0amtYw7iIhBSJRtP1qaM
VZQpJPt15PlnI0fzoGNW4Ux5sePSvUYo5rONc7oycDRc1FekLFdjffnhkqR4bDo9wjBhwRPNeZOi
P0TWm4poGQO3vSD7vuJ4HAkKMQ4IEzG+CywpzTGFZfJ286eJCX1ZqdJLTkuX0koa4p2dapIsGvDS
TNm9Qz3A2TOLAbm0IplZFVKavNVpSr/4D0VN2EtCyJeDXxGKP/djl4QQB+t8qvVIQoWCDBwZRcKs
LGsq/J8ZqR+XXcppDypYHFxqjtPjfE4ZB96el49ZD2mmcsdVt8/kCzUYsEbl9R7uR+mDNeI59uNf
L3U/+ncAttntq6A0LmTOEA8lOB/PidsZWCm+vDehdTMKtMvXRHORbkqIa49Ds56rpUNnKALWKpAc
wsnY/sONuT16xsNQmzDWyvD5K0RuvDma4YTy87zOk6vt0JN+nIV6vZC5PhzIKdLxqvgiVHBm9osv
SHFva9jbhjnbLkrtoMdqGe6EWmCsLzxcB0vshYhMmMDOxr2cqsWGxYjpmNRMQ3F4gbDs3It0EznU
cWnpn7ADZDOp+airounQ+0B/ijH2B7cr7rdeMyF+sxO2VtdZSus5vJ5sEgj70QM0lXZ6jIqerxMh
FtJb8Z23cv6ongiLEb9kqM1eNpODjHE6rH/62OlqDjQ2aw99tGzGeNrytWo4wGUlRxlWUjTOVj/f
8lDPUse222og84GwSWfzKRyM97K6E9OnCZf8QjhkZxjp0WO5Z5JNyA/cGkNBhQSBuyyk2oYFKOEc
P4inFmTBiD4I/mFzohzEyi10yl0Kt0DUCA+mF+WtQLUReCiXOWTG32uGYBJ2usGCAS0LM9MtJ8jl
iiGYcl6ooSWTQ46eivh7zpHh8xCVqSPjZ8e9LFp5vX0Ola12mFroDs88rVcuQRA/Dagob1JZ9s1o
i63nnsndvM9Hx8pvhO6say6GapKFCka+w+JrvcVhVBzEltOK+fmTetmDP5N7zf4tzmnflO17N3ol
iWZGNsw0PWWpvJJNoJgXw8L5WAIjomSlCe7sW1py2HQvJG44ATApLnFMG63XK9azcJxhNJLd5orm
D2v0ul0fwfofnLz1eToZyiAvfr0rW1WgUVIQ3vZV8ab16FiS1iZo9jrbVRLZql3WNM6d5c2gS6rO
gCtB6BckGn5dzuBsUAnHjdyXGsXhBLKJZtTfxAYgarQ3cguZYDcldJLLkAiA42SC2Cg/KieIaSXo
5ifi2iwQfNmcrSacOIuqJ8uaUkw9bfSEjYmn8fXvyTFB4Sv1GLmCW8NiAmsCbnnK/dvJztmLTBPt
KVwAZf3zeVfCfDUaJEv8xX3PfoEZhbVGjoecCyUeXqub1n+ROiirP4o5rjW1GPlts8sSCIVsETik
1/SII2F+fNeuzzaLbXjLedywfP1yh4ZwaYpV4sJgrnsz1C+R/TsG0/PyGdNonvikbagynutwBfi/
uO2umWnS2dQXDDFP0ouhCdXHqptK72ejP8g08AuzmRmgqyYOUSq5/Bs930e9ORk5c/UNboaS5USL
+2NNbtxY9SQbrKvMf8ZPU0xk4l0pbxRI1H13W5VCYTJdbwcU5dmCZ4AwWPUNpd9zHC3eCUt3jn4O
8Ol4VFtueahtbOvEH9hEUYXwjPbSCecq5LESAaYmDr32qV9uRuGaQ2AwsxeEUApAQOjRokQfK79q
ECVUkekw1wtVADoNrLGEYKzDn1o34QCReWokZ8e6ii49C5cEM8RMrb1rMQuaXbGsVHJ1GZZPDBwh
N2YnS05RN/sPhiheXiKyLB3ii3T82+epjE1NoLn3JJWC70CN9p6VJqIa9MG16kPxTPJoaDits77P
xZSDtLC1sxpg1fSQxIq45f6TIb35KHOpscpsomYxJiy8VGFj6dT9QaqBq4QBUUbl+xBnDDMEsaLX
R9GzlXWsYvbCJd4ybMqDVKo6RbWo7gCrEvB9SFqHd5vye/32LgUOcw0E3ROpNCRrY9gaKBJglcP0
pKSI24A+tYxNljacswUN0hzHzMmT4U8OFJmNxWEBZYilX1k7IpaT4IljXQ9vXPZn9g2Vd8PVVfAo
RLNFltZFW4bjpqKROjGMugN4a9qNsbPU7ivtekTqxpyg5nyhP6D3R43rCU8g6AC2+2JANbakbSwq
ZZQabnhgGfkRwxOW+11H3DBbNkFTN9f9BRCNLAiYrVa07c30Q7dpuOFCLNhrkBDQVQ1/OjMzbo4y
jBHOpGLlBezj/jA5j1thsaJcNFbHX+hIlOnbg4NyGlve5kk4/LI24Ah3oy42LC6V3y+EWAdH22Hs
jcZOnFtfKAYH11DK1f0LGbod9kpqJa2mEgZLBL1PZYictJIzBQASwifeIVaNb8cQsdhn26qDM47f
kkR4y7hVQ46VMhgYsPfVg7nKh27nlZWmcuVNEXXz/VM8fNpj7CoZ/NXy6KSmQAZlHSL84icLSg+Y
t8/Ti/7f25Dy1H6D1RPekzMEfHFbVdfsbm3rPvvyZ/t8eHhvr0R3KB8fbPPvSdJcKypVRfu3Ue1W
7VhxVYo+JklhVLKgAXvO97gzygfnTX6tPfSE3zB0dLcKfamSfTMeSFdX8bcHqNtmk08ezmMEktnX
zYDNUbQfYa514u4fyml71DGpjsb7KU7e+9VVAD1e0U/cxEva+MKAwT3XD5S+U8QRDhgvIQXt90I7
5R79Cp5bxGU7nf3tqHQEZOoWoLjUfDzWO8glmaabF0jcy2outaDg+GOn7B4TtA0ucpSWZyvrgErZ
4JB8Lm9Kb3NGpwoaAytS30ZDvwOz4vC68hgbhguohp6A835iAJU2fqqvR4Sx8RUlRSmRMCLFffnr
R6xJ5HtmlRG24+qIIbCd7RtmNcwR33NYByBlfiiMpF7o+ZvcprQ0/8DOjVbuS8chVZ8EQ1QH7ts2
4nHuC9XZGuCpbbWiMiFbVOmusi7wEM7ktZbs+bVtg9lrOkafEIEmaGfarW5jvla8Cn9Eq0wyKqoN
YzKEWCDWznb+YtRGAqv+qt8I1tU0qE+feYBc5K3kBGSfewVoAMLGLE98DyTF/tHlJR6ih/CwJzg/
EE9VuRL9NfE+Zq0s2rfBHT5tohTRYLrDgk75Hdwjc9/TDwfebXra9a3+4PmMu2/7hBGBvUN+IsCn
d1hUMqJiTTjQN8pLR8vKfRWKz8dVWgkiblyMtXKQ/0GIMlAk7MhH+N3DOHO05erQAE27Uq/9tmuf
tqwlYcP6LVT61QoMHs9HJssPXO3wol1RSQBrY82JqAN3auHyzndg80bppvIfviUzQRUhQ+tLTu1k
YoWj5vVYN2FLwx5nlPCOnvXVXeM104Wm+dtmiJShf4WizbFd8dNPDtwi6IQZZgBqZ/KwtsNv062c
K5eWE+xJKaIGCkLAahDzFsn8qzwasHZQ+6Lp45smHG/TQ/kXPB/1X/IzmLfp0DCHHQAXM6EGqPbZ
X2Ky7mA+F2Lzs0ZK9PUKmDsOUqBqLALTiaaLZVWk5HYAoBcgPGmJ0eTZsXkObH6+jHDhNU+YfghM
mYZ4kbHDWqkxJck1eRq3ww9JvqA0cpIytSHYtFDRgIjY5OpPMYni+dPATQiAZ8YjQdq2O6YCNjQo
+8iP05qeVZAljASFQf5JOzrML5QiVH9GALovFEzrS5u8eibGQZxer5tvjgOuq9bmqDY/a9YiCKYj
L3fseTvZ0tAmMPwjGIErYSOe65HrtOdxEQmDudI+EVh+cXomc/AJcDTLj1akZCjpEZ7mAJeoLGaz
NFutj3IVvjk2PM7CA5D8ZU/YlCMd46H+OyGGzLxyHVaaCC8tuNX9P7Fwp7E30vrkAi6RW/BemknS
3G7FduKsJ6cFf7J5zmVAIb8Yp6Kgdwet5pDHSBNN1ce3uAkZfV43x/uHpnPjifyKDZ32AaFqqMb4
imrvZw3tApew+HEIrOQjlujrASVg11NTooGQjaRkxZV1Gt46BHomT9aChzcb1el45HNA6wavCNf3
m32rqrySnJPdYFKqyi+gKtz8cCn1XaqrCYGLi7fxCv+oW7fuXtNLJsKNkYEftnZgZCZGWXotj/gj
5kyY3YcTUQptWsbb+tN2yOWhNN09vs6fV1/+/lUejtMLJGMFBiuUkq3Sus0j97N8D930JVvioYjZ
nSa0LPz4Xl6msDCfXLK0LJ+/rSUrt56LmQA3MKLNTBhHWBXKiPnAbiKbEPNImSTzEL/GRcEMHjYv
ALhm71LWzc8nKyQ5FSJY72hIDVcKW/a+kw5+kxV/DGrlpDqw7hIUufvP6PEZm9hsTSpxTmq9J/pk
7u/UvRXWSSqfspGNOTnEkl9x2tVNDNsUNs20l3aGk56f5mmyoZK2B+ZMaCN5FEF4evcnSUubDmu4
F0sZdu/Fq72UyZOIQ/sUX/zjVfDfJFyEMIc7wM32Dgia7O1qemFDWZ7DfjV24K5v51+Ov1M6U0OS
VU78RcI5uNgfyMPzpCK/Udb/vCFc1Ydne6inEqs0qQOOhwfDYjAp+bCU47i7cBiCeSdIEjThcQFn
tHl9Fxbv0I0IxoyTf+Tx3m/axz6tc2OYYoC+JdgVSe9q2uJCiO0naxk3iyBDxxm/Ix2AutNB8D40
PnfhunsPJXUQ6SHgNEzqaflf9uUUGTuT89+uLkAuGRAoTjtcDT5kCDuox53n2c9zWh38Znj4HyYt
MNFc1MVTgBdAbBVrvu8vePNa6UJe49o6R5kZhxAN+mNY9OacOfzO9lZfDh/++NPNr3CyTrtLJf3X
4YP2dqKRnBoAwJBy+Ur2kOzrI8uKG5vRRBcvCOa0O1bj1v7JWTLCFlx4Luy1jdLnXVqeQW/5lkjW
EgvbY22MTUvgtYwcRnWz9rwafYBvOvQVj+zA64/pARaHcGlTX1tyBIp0TEV6cH71ohD1DhmJ5r8Q
Uwv7L7hSKq64ZHz4+3Cn4cmXqtG5Ljm2pG2Pyszmx+nk5MY6JRzC1wrETc6pTNVcBgWHIYp0XGfY
2HnBRbJZmHjUAIwJy7Os0P/Dl3R9ya9hkxCfPV8y8oQsbQPMiSXrYt7+U1AwUIHSI4YpboIF3YQG
fl1k97on2sq5Z3FOvCz/+zYeYU+ZYmVJ2krxgi7bKaRtPZSjez0udt48HFQMIx5b1hAN4d1/mOmd
7QZcEunCkNnEhZtxGxbRnz1nvSi5gsLxFfdYI3rdAj2Zv5sUGzDTU/nyIQB2/i7Oo1+Q6RKW/TEG
iewVnehSfD+h10f/ubt9/XXQAvFT9pguLDmtEON/IYhtb8xFRN2uNWDVK4IXyLlzvrAfPnh3oWNO
gaF9bWjqGXGitIppOKCkzSNtwcuCD+dHKCh+dAr9J+qPeHpoR5d92Jl9kjNsknoLG41A4Jzqx+ay
LNdJbgeWnI9kc/vvQx9AkEbMa7sQkRrx3aMfiP2UokuftMZOjF//LlsEFfKsRiXKY3ByiGNjGAOo
mdl3bUGsRbiDpeouzq+gsCCQW+BIK/ctndxOB80RcLxtESxoskd+4BVtV5tW61R1kK7sf476Qzg1
EqNLVQIdDnpFxvMdp4rmOG3tJaGI86EjPInH2mdMbyR9xsA1NmoucNbvvzQnxIxEc1Yt+VtHHGK6
eGB4KhGurPsl8BRN4StDSevQ6zkQJDSc8hllOLa5O3wU7FiVcF8cvgfch/AlNqY9FCBp/2qssuDT
MX1heydnydOZdeEr5Jecis52ynNYRUUf+NGUlPz21sR66LZThWqx+xufhxWX6H3mRtgDKKI/EBye
GH8GBl+eZBnN1s9QlLkC1h0YcUTS/1Qjzg324yc3K72AtYltmFUZYnO52nFc/sG6zJeJvWsqmvRh
UKy4fkPTr3i9FzhiB8XJnqRy5F9ZLZQ7s35pKeGSXWwuNtj1rCIM5IZcWFN/3PiYnArlXmckUIr+
scBpUZAQZtK6fjlMJq3Jw/JDUzfpCgQJ56J/Os7rTYZ5xoQZ6ZJ4YV66vWQIiTUVgpZbwAo44ppV
ujD74XXEPfRy2Q5eisKnfx4kXU82bUV2+4wHjWvOd5wSZ1Dsy7/7JYgVwzEOzn4o+pjdV5eLIWex
NLldPyfIMIjpJdc19eQ6UtjLUBCNOnX7ATqV+kEdUnkvv0raR088q77Ssmt191rpmh1YQs3PFce6
24g3vHGtYOKiIpRs+1J1xrGFgSIa5j/pV/SaDmdto7ZdQvZsBdxEFK/jRr3SLHNOnuBcwiNoKaIs
vErk7wlxTueDg0sJqEUwIk8l7xTySBEI+eZYMJIxy3roCcfLSkDLcZbvqAQywDqe518OHu+jjjI1
UcUef3uuOgjwlQWsqDexijqjcmlmhkfrVQyAx5kNRV41MNbq5sA3A8HB2BGVHv7kaE9XrCftO8Do
X7bnTsvD+0iK6UtAENMz32cYuxFHVKnT9TmKKvi9JSjRUCjHJxizVsAPQmadJeT0Ju0xqFdRuKiJ
3HITEXN7SYoIeYW6rVOqZKnleAbuB/kQ327px386rZTTfcMwxaM6APeg0NrrP5sTlIjFEtmFZyqB
r4Kl6qPa7O3TTxvFo13SfnB6KcsmF505qAyyF9wkpkT5uvFMTNhWEsLWCxh2E1mVQ476HUU9DNK3
ZcRUtrGua20e42rkMwfQLsh+aWKM/yKT3Wpwid0DEN4G4xz3sBeT/lTNTzdMWDzyhkyNIhg/jr/t
2bIvfTd4GXil1QKyphliS8bNXjOfKqxKSRn0M8fg9ffVzz5Yt+IyEIawKdzc/CceAIGgo7DwOF1F
cnt+een5fSisVfeOHKpzeodrXFARp8o1D0B1fU3iYTX4LBe+rUVaYHTih4znZ4DQgBy5UYlwD8h0
1Yh+iVqCGN6YhAxCFgSN42sPPoltGvD4QZQv2PM7Ra1+mg2833oMSz2sbqmy2SJg0caBgorLcnl0
7PuCPn/k1YW4I33rI3q7RaSJVcbQb3tEWmWOj9+hfwTKrxBrD4W1meTdksoEXMs7WLvRfN8tnQ6I
Sf/WPTq+3tbnsn4EdiisWoGzXRJBf3OU6kHS3lYPaVixq6jzf8NsaVvuzyPBtHfipsrOPRBrHLUZ
Gxx4hY/jJzv8tB7ForvNoUHq2bRuzgQ55GFqdK94qp2Tu6j5x7FUmL9lsxbM0t/qiKVuD1Qg6HUD
8oJdV2J7k3t1yYQq/eMGNTnKITm9naxdNMOxFctSlvAibwIb30voPNfce/ZLe5FySHvx4iAH51nC
hqBVsCdgTz+sgeEIx5xrwZLvCc7QXXjzrbDMm0IoHn8rBtHOGRpteaVHc7K54rbJ6gCNfJaYsP9/
95dxL02MiUGsg0CAGBkChiJkT810Tsc82Q54ySF1U6f+REB2qlgxJc6ptPiuQhkZbhuceo+QyDe8
XaOxdy+oHYwVLy7lw5Xl0U0fGZzG0YAwNPcDRzPMVXyiT7bbR0c+w6ML1TET5YH3+NtpIJeSPJyV
UhfLpS0hU3Vb91sTHeKGBE/AUKiqg9hjwb2Hi03z93B4bW8hOZa0ZpdUcFMjeFZMGmp3XOrgiUJ3
mDkeh0A+nS4k5diWGjxzaZdLfaaTsDpjed9IUwjz8QQzwev8XbrLdmTMXfbclKWFzz52/lEpUvNh
C0XZ0Gua8VuoMugQCTRilTEHclOkus1CIDl8CTUa6XeIfhfsxzZs81isluVzD51qrYX1B/ggXSc9
O+uJst5oSYroxi7jdqdMLkn4AoySzOrvEchozMw4o5sdfAMB4TAormKShMa1hF2vf2Tx63Sp/ch1
EHJPdVAoxJ+XzDJcJpMsuBwmbfXT2i08TmCJH+YkxysmK+Mo31LR9qUFktOo5S9WOIdBKK3GHr5S
Df+LhjESaDIoNlLDg7dm0xQUghsdhgj2PElhP906o+esQDlY/VcFjI4WJykL/XYzVspqDNc3MT5p
Tq3zrJQ4FbrDSBLoF0eKVOlGU8p6lk8ImFj3ebKo78JQfddEql6zu64NVtgyco3DlKrORZ6N3h/E
WveYKHgw3LYuh/nY7WqmRwi5GQWYjfbN3dS8ZY0nyPfFoVttsXVsEzuylaXJJfbnRY9JSS9FuMq+
UKWPSXHtTyQHNeKqY/1IKdBDsOvikksKeCy7sN2F0qvUGVC6TyWBfakEO2uSHb41s5BqEDRWJ8tY
9mmgHYxXjrWvNWliWCQsvwmBWn505fE7WcFBjpQn0kJOMvlEZUf2VqI3TT4u3qqQ78NSEqPolJgA
3rmHj2vsTZz9AHrJn95CBM/dy9LIedtO3Hb2hcCo8Pu0lsyPeySeqfT5yNLstUf9IZhJgGvikncN
PfycwfuXTmlAJZ+eckiy1Z3gjB7viYBXlVkJn35z75Ov4SRJQaDklpUMeR5gmq3EAjiR1xgGW7k1
jKqhj3QPivkAMFzcfBYEaXK+l/sBAIIr1pSzD3IZc1MnaGrAdJ2tzRSAPncrqBZjDAsO6tfyTOBn
lt5Ex3qxfbPfgRSVkktxYfxCL8c2j+8I9M9kdpBBnmHZgxmejwEZFEnTuTPN7pqx+WmpTAwHh1SU
m1jvi3O0Lz9as01tJaNGOCe/HvCrru/kp8WVMAeMLge12u8A5+fn6Tlm/b607JSrDMTSExiY5P/I
2Odx8dy7fucLbVv48kaoIx0n/yXKUKU8l8YXerYCgmwZdBlKErVMkeIBs7I86yQMF6D42Y4V0Isy
mOvzeyE2+YlQBuqbpsQWQwRYR2ACrnvEXsoKZILiOTUR23ICQdwharCNqcrpKTL7FJ0YYyv62VMS
QuLMBoQYTo+XHRxwgqd45002ZYwoRHkOEvUYDzPmVme8avo1Z0qd05bsL4ItTt7XnkACVJPwu94N
DRiBpSTKVpXU9enG382QI+G8a+ZX7JydnCEe+G1PmVTyry9Otxa/Cs/sN+WNmm2jI+zIZaZ6UsUf
M13dug4DG2dmjL01bubeCGVcKPKoUhdouY4fNPva/v8i0QjxkwKxGN3kDGoALWb3JCWftTk07mAx
wwFQt4V90uae1C+HyhvyQQskQOHFTRUDb4SIEvRUXlbXJAwxWUx37p1xKSzBC+6lBO3ryXcjpnad
kwVih7yG0qr/tm8GgXbX56YIBoaLoyIHIj/pwXeP4zkSD0ALGDXAxhCjhJLJEO094Em7w7VGYhDt
M0dOYEe80YWHdca+3Kev087gbyWhKc3sMO0ObpGDnJE5T5QIYNxBA2+ncPtnOFEX3makg22gipiK
X4GI6Gph8Eih4kF4jf7ExD9yJgm2Gf1Pqh0HVwZvbyWTmPs3MeOMvcTkFBm6PRXoF3CkaTBurfYy
UUO94Nhhozt8htf3KNErP3x4WlC53XSNgZe7pIsgw/Vjm9gHzbCPN8NkbgpgS/0rbVu1kUQ77eme
TNuboAF/34AYQqX4zEn5GUnDWJKVC2RmBk+XAkYQvQJcAkf0FHddFbSDa6T1tB3uRt6jD9A562Av
ppmr8PpIsiF4YwhqYahwUhqUMVfon/Tla01W3zyKJaLbj56R2esYJHn0/IufvGV+xxhgGsLSeRB7
TVuHPnGyY9NtWz6aLFkrH/BYSNzN/CgGydp3lu/Z0rfFsYWuYTAj/FfGRwcshrL/ANzEe5Dkuw5O
2Oq7Z7iWcLTfxhyIIVfTesAiJKvCtQK3qPxAltPs3kga42SiYft3sX/I8WXtVGPBW6qvIxAVKjgW
1NMimOp3HVQvVu2MvDJbGJ4a7aIvuOkbGF+c1lcfo2q3sos5sSK4bqryAJamU0i13pCi8yOhrb7a
YxrIXAg63PIoWJ9JqusWDpwzVenBloopXFWfb2WLHHBziCNHX6Suk9jRDzUP1P1fsqvNGWOIgQbY
YZUZ4dGFpUlhR3XiYEmDpLppOUPIaYeoZVz5fSNWQ2IjvK2v1iBHzN7N7sYAI7NySWSD1mJ0Xbq4
9l26J7EXRiz18Onuq5l51t1ojLXbo8ZKoiTKxjS/Z0UoSOyYa/2NzrKoJZuVOz75XEZls+zspjLx
EL5496xglhaVkfHetB8dGrgnAltgnHbuKnelNlAppOgB+7zuis+3uuvnHLQHDHf28sGFHvXxuqFZ
aKrSeUfz/t94PncnZPKfPq2I8KDC4Zkho8D8+5zzZmBwsTbnYTNl0tktk2ReB/0DpbvGlJxIM+7m
MZlStazTazFdHFeRWNlSu/txFT4n
`protect end_protected
