��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$Rx�y�<��wA�*;�x���@�̦�W�X�fa�M-$u����n~�%���P�$��W��kYَ���P7�?UMfT��q�6�U��k�>����~�\N�(�����X�e���/6U|)�X2pF�]$h���d.���9E�	�IN�f"�\��e�z�y�b�����Oo2�?�qˁ'�͜k-�K�P|����y:����3�l�d���bl��ˢ_�d���kx�rq�mh�MذM�`aS�.�DW�mS�9���Y��+�>��!��!�T�uOB���,��\L�7m�O��W���6����'���j)n_�I����2:��$�K�2�Sʫ��l ��!���{�l����.�j4�	��很�̢=�����N��s���s5���_�R�>����ТP .W;������	�"�מԫ�����]�#7@O+?�⡾�Ԫ���e�O�\A�	�ͼ���ƹ�d�	@�nQ˰��E؁Bf���|D_�%au�-�'���w�*%��"AM$w�*�!��os���͞X�������mIOI��޸j�r;ZzO�=W��q\��D291��2UBs�Ij����A(�WüFb��� MXF�,n�h�Ƃ����-�@�D ,�f���('��z�������A�5K$�8�KGC��7�����E���=��{����mx�>, 8�[�Ԭ���\�I�⪞M\�á^�{���E������6	�?��N|��&h���*��%2��P���WP��U�f v���9�d�dK���,�M���6K��`��S�����j��6��8:��P�=ʺX"�C$9y�����l�x�v�x��x�ga��a�Do;�WTnV�w�kHn%f%^.Cc�d�Q�]�S{�ܨ�C�1H��L���p�V��k�/gE��9UO�IB5����-Y�̆�:�w��gBz9����5Щ�������#/.���@F�U�����M�9S�]O,��1#z���5<�
�i!�����S���>�T�?S�?�t�����a�f�L7U���E�N�S�(�*��70��վ��\���ş1��+H��iG��ո`Ɏ�(�_�7��f
�[��1�|���o9;A(�8�� �lh�qA��i�� %qz��xKyleea�w/,�>�-�6tisYQ��6§�(��ft�j�ш�p�'�Fk�o�o���M�i:Z_�`L����V+�m�u�lK�_˩�h����*�l@NpN�+�����ja���e��1v�:���7L�g��PO����j{�<�B�� <	�*l�h�Irx�����s�`�+Y,Z���zy�^�w9^�v�Xz���J��y����QI����l=�+jR�BI?�N��5��au�}�x��:%)vh�%)%�}5��q0����y�|A���0��b���矘��z��%��7!m�%���-N��AB��i����^dd��e�^�Q�DV!̪1AE�t�R��(v� 㓚�n�_���b�-4�����~u��u��nq\b9���cX���^ç%/Ns�^���U]���;gh�n�5�
�B�(�Zӊ�\(¾#'3��6S� ��(����p�r���)�� Oϖ�ٖ� !�z��s������ݔ��Ͻ�]A���Ǭd�L��?�L�m��XZG��U��+>��<5�PW�=��� ��Ʀ��A먥5/�����w�N��Zk����`��28�}K=B�:J}o7�`q�K�x-|{�]��Q�ّ/
r�[��苦��@����bY77�H�G9������>�x[#�|�83&Q�=��z(ɠ?B��ǆ;��bĕRD�w��1��[ ��0��Z�2�n���������+��7')�8��|l*:��G-�9&�aTx��\��,��C){�/�wwՅ<�nf�h���w��\�w�.�qL��a��;�
�F�ӊ��C0#:ő�D�a�Z2g����J�o}�\�����6���<��gbB���x/��|�֩'I���&G{N)������?�<B�����rs3CBI��܂����f,9
r�+�j��$F��-g�G/�Y�g�����%�>���o�Nᇮt�N&2zQ�F��I2I$�7
:җW�O� � 2���$_���ꗧ�yn�\�`�&= ����"��{����*��r�/ѽU�=��*Q�$�p��C'l�$e�y��=�]1�
�v��3A�m��NԷ��|}M��Ǒ�����t���TF�,U���c'�9y2C����X!�ͺ��TX[>�?p��7CK9*�N�ޏ�!�;�d�G�-����J��7���0�My���v�w�z��m�wR2�q�6DE�����P�w���-ϥ��1m͵���o��z�J��RJ�	�A�Т���v[x��< ̖'!ut��=zN�=IJ�$3�+fW�e�j���E���!�U��h [�S�?I����4�v���O�!B��|�miу;�4�C��/
� �-�vRC��ꢸ�"aI��i�r��CI��;J�A��$���?��vsZ�I۲���&�Dòg�"�9�iK�3���������z/r����)�)A�j���K��9s���Uo��P�puE���6tGV^�b6 ���<P9�a-O�Z��7)��:��a2����q���DC�474����L�7)�����^��\i�֬XF�?�$o0Ed^�\�m6ba�e�]	!��3��}0����5*biW~�}� K|9���w�2���ek5���s\��K͘*\��{��� u�r���ǰ9�r�I�N9>���0�0�f�����ϭXj'ѸML�8G��m|A�l�� ���5Ɍlh��@�+�=����zԼ�c���W� �=<P��)u����d䱡/�� �#�����S ~`f��%��� �&8xE}"W%�ś�{M��0��
d�3�i���&��3����z��mI�P"���t5����귽t��g���=V���R�W�d_����X]�*+hK���ԳPˆ�"����޼�w0��Ng�]*c֖��I@�F��.:��"�h��Y�����vw�-3�e��ۮJ���%]��.��"�c��#�bOV0�nR<�i�I��gة�2}l ؉V�f��X�U���1M�a�}ѝ$���Ɓ���G}�������Dx�cN�/ռ*�8��֎�>��a#�pX�u-t)A?Ui�)�SSv��.�^�/JOM�6��B�mM4�M�F�!�xך�0ش<�]mL��!܆�\���.?�m6.�/:Tw�U�h�U��;c�.�����;�$;���F/F��(׶~D��b��S�j~n�oϚgs��K�Ms���<�6Pz�>�O()@3~�"�(�wX%ү2w(�Dv �\4�T@ܡzG RΜ�>�;�oK�uv��M�?A�\T[bR�
���\�jܽ	Iܒ�O:��x����aG)�F�Y�:�)��Z�~V`
.c�YLȿ�YuʳI%�ȴ~��6W�\E;A���ת��^�i�a؟h�	����0�	pB���W6��2�"�A���J-�0�X�	���'s�Z�Jߢd#��8?�RS�ɭ���[�u�߻��wJVHǶV#���L�`��h8|IƎ��$[3D��[���4eY��/�`��ï\��Y�!r����}���棦kQ�����4��O�I��h\����h�$?��tZu0�u����G�� ������6�2A"�W>3�'�K�f5�����iP4����(�Vk�lۊP�X5�Ŷ��F��9�P�@nc�޺g�����.���t�Y�t1��cC��ļ�����Fjd
<Z�Q����`��:�p�+:1�?���|oXzA����E��$KX�Zd�7��*R�)���Ll0k}-��b��c�D�E��V�����6���*IQVs2��l7(���=x�B�}#Ά17�� ��0jO���Ӵ�����7b��S�dG� ��H b]V��x�]��
�m>e��"������+��RQʝ��>+ӕ/WBY|Ը��v�K�p��=2#�s"�ZXh�����dϽF�V��93In�:�oEF���A�s�@=��bC�*,U�?�C��b�����q�
��I@����/L�F��^��7�4˦��b��@ak�j�En6If�+j�6uO���wL�߂��}�E�A�Qee�j
��Cqߺ�T�Q���cUL;=���
�hW���4�Y/'���8����C��nӪ�77Q���w���Ќ�L�Ꚋ�w�6A8�P.9�k��٠Ӆ'W~�����* �}9����@+r���a�<W�3\>Z�
�R3���hH"��U|>8����hʬ�@����]qI�Vrq���飀=|u���Aޗ�"��G.ByD=s��n�a��X�&ȋ���s�k�D�-e���oxk}58���U��G�������oun�Ǐ?��o:H8"�K���~�)#rS�.�b�������e��<s]J�ኇWy���[ۨ�����rGب�X��s��6�K�u�T�I�="�8�С|\��/�s����fU����k2I԰!<գ�.&`f��1��v�9���=1+����p�嫰TM��|zC��!><@�#�Od�l��\4����ܣ�0�>�Ea���m��+���	��=(~>Q�����fiңCM���*>_��{����h���{����0�Cz~#(ܴ<�IO�j�BS��(��~<��,h=�w�������6T�xۉ�E�8`�-��d�+0������K�0��Z`���{V�d#>���ݝ��0ʑ;�A�Wk�� ��c�^c�& \1�)L ����^e
\��ʛ:x�����V>g�Yd]��3��]�]�/c.8�*��d��P�z��k�������9��ڜ<��t�yԬ��4 �@���Nb����ݦ��*gժ���� A�zPە��M6!�eyJ<Ѕ��Ғ�����%�S9Ԯ�v�WG�����f���\����,����q�J�����`_ȕ��2B�c9	
�w��%�2�K��wo�FO\ǣHW���|?�G)���������d뒁^�F��bJϪ���!����hM!,�����E�+���	�n�j<&?��^�zxO2�����	U���w���������z��Z��wl�MB���Y�}�Pm�V��S�=���Ž�F��6τiZ<��28���B��\���h{��ǓŘ��/�� �s���n�FV������I�:��*X=w�zs�l4�v9ǼO���̕���Z� �:�l�]1䋿��'*)��Ӆ�CHB^Q�
j�?j�����b�������7�0bc�4����Zͪ��ֈ�Q�P��2�+Y�%��{�TL�-)���w���}^�,�XsmS	��QQ�e���Lp�����`wM�t͕&�^���? ���8n�=�&�4���~6�p<�U"�|��!��Rj�IoBg�@̋Oͤ�ehl�h]������}O_G~R�R
����\��vJK?S�8�G�j��{�7�+:�Z��D���
����!�95���>�?~�"��Q�F�ZA����i���G!Շ}Yy��$��)����d�Rㅪ{��6N6���$
̛iǅ�}M(j����r�LݩE��x�׆�J�� �>��l#jq�7cs�5/`+�u�w��U�ki o$ҹ�T�]���cwX:)���%A|��侱�5��өNe��0}�e�5��<�7���b��mwRh?�_�y v˃1��qq�R$���6zV[�t�F�fh)�\�3݄���_������[�h�$��+��j���et���o�Y���[w����5�Oi�"Q|I,��Ʌv��㹂*��ٽFhwN�	Զ4�������x[a�k�ƃD2Hc�C^L4�� ׋./�L��Vȱf"]���=&ָ�.��a�}�D����G��)(e�&r
A�&JRaEL�/̰D�S>K�	����2jg�<�OE�\�s<Jp�q�۩\UZz@4B4�5����J�D���pJ��Zb�9�,�,IGy���X:�+�?)��y?*4����ξa=!XU�pJ�2>�L��/CV�v����jᒮ_:���W��ٻ��1nn:Vxg1�xe|%����ɷ���#^�0)z��

��6�oWb��R�٣K��7�v�[L������::}�V[�կ� �g�������뮡�v7��nЛo�@�>�z���1]S釼�Y۴�"��^-B����s�POq�j�s	7�C���q,��r\滽~hTn��o�1r�m�#���+ -~<K�\�k��q/n�����`@�����DD=�/�%VcRM�*�m�^�m�zv�vֱ%�S�����p�D�2b�����{�E�����@�a���yR��f*�RɼtSǫ�n�#���������1�q��QC]��T�\)�R�1~#��K�A.��MC����w��l� �<�/�����W	C�|�Š����!�h�$�r�L/��.�u�K@SU�C�f�:x�lį�4�k�����H���#�nsd��#�%Jr���B4�6k�g^�y�M�$&��/%��p�3s��N���%u�����ifV�a�A��qk��Q�$���v%g��N��������_>�(*
�Cܐ*����C�	NY�o���I�g]���!� =��=0(iW_��Ø�8c�{���K���?���*ƨ�C�9�
$x��Zق�Q��VP����vi��:�a2�?E2Ԝj�\z݄�@�-rOu�����'��ĺ��I����
�����j��Ey�zۼp��˹�97�rJ:� oi������.)�h�N���%��ʽ�?��%�� �lI����'�Ln�e�)��/s�Q 𨾋���P&��j}�iɉ�Y���`�/&2�D��C�:?P$Y"4QgU�����9�T�����	4�&�C\۸��o�������Z���ˉׅ!�b�u�!ѐ��3�WR���b���~Sh/T������K�_}��j����eP�� �}��)�!�(}��8���I�,��a���g���ڋ	����`�c�R@_��hI�� ��!�A�iW�/?b9M��,�)��~�t�4�SL��6�r��^�F��1J�Izά���11�ͳ�����D���ְ���OHļ��,\0'O�u90Կ�������'ӂ���֞�����-�E�&�����_���Jj����h�^��2%p8h5��po��4��@�w�$s��<"f/��)�F�N9|����C���go���OV�9�I�\ӕ��v��l��M��/���^��#5ASP�zk�L��/ms`v)-㙈��-������$P��PGy�%u���c�D���ITI��A�M�̷\����C�A���:m�*�'��i�FA��ѱ��hlr���I���\8���{MwS�%��x��^(�	���Am�Y���?dy{b�"^6 �裇.:�?1\��H$�g���`���zt�l�c��5D]���j���:�zR��Ǐ��h|�؅C�9����H��\��.%�b��T���8{���<�!��3g %���!j���qy1A�9�8V�Q2=+j�^���U�g#0��4�hE����07��#�d��*2���P�4�5�°�l�w}�=�FV���J������a�gy�s�X(ɿ�(���o��6Z����G�6�}b����>��H��X����j�~�W��0a�����Sd��TFG?�ҧ��0ku��Hb:d�3A���]��',�������+�S��*�9�9*����<��G���m�me�}3�IRW�[�K�}���*}:Unk���k��p����XP�T}�J�4�3d⺩^�(�����N��H��`Ԍ��h���]?�=b ���*�����B�~����o�x�Gc��Ff��D�~ƚ+(u��
����%�a]���z�Y�-#zS֗�do����t��Q,1�ͤ]U�,
?�� �bJ��7�kγ��zU:��cv�fO+��\g���oִ�6b�Y����qz���>�nl�D�sa��D]<����CO��Qa2_�_l�+M,��<�"c+�7*���A�4h]�&�6��r/��_����
VI)�g��.����Ÿ��O��,CѾ�����;<�mq�1\�m�6�;ה���k@�(/�⒅��p E�$��f��E��70��[|9}��p��N�������V���_�ş�W�.�T��?Uvq��oL�lg���d}at�zjs%�<�U�S�������og	���&籬Vw�bKg-!���?����dX9�o{d���߭	T7��PCb�x�r*��oZ�p	;�W�d�k�>\i�H
��V/*��Pge:v�kp�������[�v�]6-d�(���-@ƻ,����%<�U�f�a �S@�A��9+���[&��j��NR�Ilr��q/CݳG�TDG*[e��e<�Nw�K�ါ�ޛ��[�,i�/M�P�0�8�-y�W
�<�9g��Q	��ς@0p��T�FI w��7��HlS�Q�?&g�+y�.��h(P99�������������V�;��]��B��n��W����������+ F�V�NK�I��S;�o
�OP�k�lĲ�6�:�b�8�W҉�-d���d	�V��1�. �����+��3�w�t�E`P�R��	�\\�Sp���4�
�Z�c��xN�c� �eJF��BX�*��$�^�
o�T�Ѝ2/i2n��Ҫ�R��Ly��k����:L��|Ɣ��B\��y.�k|�nѻ��jԠNg���z�f�$���R��]���=�wz��njcw�m�D��@��R�������5.Yx��l�����D�z�E�P9�AT��y��8zO�E�a��b�Ky�zrI���LnO�G�P	�23C�,[N�s����{(��W��kiW_�B�1�I�.�r�\�����p�2�Z�z�]�>RE)t��X������*�C��l��[:Ni���O�=��v!}h6�Ģ�j�G�(�.�à}ɽ.��>	�,;,���oo���r��F��M��7�]�O��U�g�Մ�Px����8�'�xq�Lu��7�6M���z���U��&K-�+T���i�|u��p����?�W��MaW��x�\֣Ɔ�����Ho��fJZ�N �����:�>L��k�o�\"w7[f9}��4���LM���<�4����f��w�"�K�J������o�PE�8k���d�`��$/��KpW]��96���璲�(���=�дW[�s���..6fQV-���;44��
s, ��5� w�5��__B��w��T��ۨ8[�kY.�,���xY|e�d�@��������7�0�1�T���v:��p��H�}���D*,�dGz
��� �%�.|CQ@m��d �#9~`A� ��A�F�IQr�))4_��|���8x�=u���1+0� �Z��f��w��Z,,O�<M'{��0���g��������Ε 0P�����%/,��t�%U�Ev���e!�8�Yo���6C��s�n'?��p/ yw���)�O�$Qxi$|9�L�2�C	�LGB_] ��R�z�G���4�/C-��@�j芃�N`>w�*W=����j兾w^ԸDM$eSj&J�`���_��)��[b����J�V��z��n?6*z^����Q��}���j+��l��a뽤�D�Ð.%����EB�Y�s�=��5"ol�v������F�`�x=M5��n!�r`t�ѡV��X�iERe����m0Z*��@�J�
^�/L1W�ώ�z�/̀�B�H�-� ����b��Ͽ��M�v���ՙf)r~ q9Խ��]}q�j���� =�C�؜���l�뒁A�R��拏�@iݝ����b¢�Y�!���x���	voE�ѡA�YLk\��j���-0[�8;����>}]�u�+�K&��`+��-�&A�)���[�o0�ēՅ�HG	���S9~�Qal'�F\���
��B#JD껟���4��}�v��=��ʱ�T�H�D�1`��6���*��g븒J"���_��3��>\$	dW2%j?<@ �,���.4n+w�b����dض��W�1��j��vw��[�^�9�RS��<�N��2��Y��|���;�������D���i)qU��Nb�3�R|�۠��q��C>��]L)���0�)j�V;�:<R2�Γ��Y����� �k��k�b�gC�ik�ȼ�vIv�bʾ�uQ�85����!g��(�7>�i82Wg�ku+%{0�a�4�ɶ����H:ǘ%��D�,�B�<�\f#i��m��	�V� ���t-�/X��s2�ko�0m�L��HA���#2�C/Ǯ���D��+I�žE;�-��7Ϻ��c+�}'Q����T�O7e����K��]���X4	`7���hC�u;0_�Es8�a3�6����4_g�w�Q_��:��YQn_�5t����ሧ��"�J�c�����ӳe�9�u�e��*6�"ZK��$����}fO�*yH�ָ���*�C#Xah�_85�3>�l=�w+�yӭ����,z2�N��ڑ�a�%,����Ղ��h˽�,���L�&�MBM˹O�$3c�CC'Gq0�����2� *�J��y�ЙD�EF�� <\�w�V��0�GM�d��-�����-�]�ќm2G�d'ܹ�A���S�@�V�l,�>��u���9����y�������yt�p��`n,{E�}�c|�b0���R�M��9���hr^qϸ�S(/��*=�J�&�	�����CW�),]�T�6�2v#5Ioh\�9�Wh`
���䷧�0r�mWw��`��?�\A�C�|I
̙Ju/g�Lc����<%&K�9�ݮ�8�\�@_�XQ�?���b������n0�@v!���	c]��^��Mz��q�R#��D��||f���u�Ї{#��nV�~^�7���b��򞘞�����u�Q�����f+n�՜�$/@S�8i6rD椯1��*?�"��'�nK���
hf�5T���ʅIU�}|^Cjؐ H��d�̮Z|t�j�����iSC���3���6(��*^��)��v���N��؍ʷ��J�h~=b(��x�ٰ���cT�>�6t��[fJ�x���䌓���4R�t�ɕ�������_Q�P���`�)�ۆx�CL���Xl��*&�5��H��KӦ��4�`0����v}`Y�v+��`,%G}��V1(�!��|��^�F�DQWфe7 [��H��<��R�%��5Jc$L�a��3�r@L�?�l�N�2�tkyb����:_��{i7�{TM����+!��O�����2�����G�_�=3��K�3����)���d�V��6H��S���\<قkzW��;�j���+���n-2Kނ)�*��Cj��2�97�.�ֻ�����c���>깯��p�
�M��R�U�ΐ?��d��T�����E"����g�.=��.��;��o�'p��3x��K���0#g�?�g��<د�i->����^N���k��vV��i!0�x2����Dzr�����G�M����*�?�l������G�6�'��!F]�eO�M��<��wr�(���t�Ç�wH�K)���m���w4)�<��5�M���N�:Jمw��y<��b)�����T��.�I(�io��P�t$)���tl�I$o�k�tD�ܭ|�¤VB�3=�E�@�A�6�+7a]!B"�&�1o̕U���Yg�W���tE�Z&T��ط��aKw]�l� ���ۺz��'��I#���S��X������"�{�I���㞳��d7OB{78��*�1��x��)�� ���3�[-:�D��t����/�	�m���e�E�L7lF�qY����`{v����l�A�	��|�l��w�5|la0�H!����}u�oD:"��h���%��=׵��қ~9��j"�d�fr����/U���K=����i>gU8�[��R7o��� C� �~o5J9��ޅ��!�l�P(?�=����L�w�ZIz!.Q��K�Qu��dRr@}ϋPN��ߴ�4o�Qu/��%�?,"�_��25�y��	�W�j�R՞�+�'�T�Wx�r��8g�P_w�-i c#j��F���ܝ�3�J�<�����ƙ���B)S��q�����L���Oy�� ���r%����8�l^�7�q~�Wɴ�E9��g�ፖ�j��Հ�<�1��ԃ�9DK����{ܓ'#����O�X��0���6�z�tp4Y,G��P�P.O�"�;���2��N�
�AcJL_���C#Oo|� I�`#J�Y���#U9�RA�����p4�8^�a;��O�K���|Zz���U�TfB� �բJ��n��F�DðM�u���On&V ��r���es';?R���x��z�j��4�H��#�);ö	v՗2L�g�n���٤v��4�P�b�7/z.�t���t||��)�c��@�׊����(:X���R�az��+���t�4糞���SM)f�4�J�I:���R- �"�*x07y��ӉgX 5�"� GƟ�貋�-��'ū�Im:͢9��NU�
%D��}��`sg�ty��57�t����:z�ܝ�ʂ��A �r���M{�XN�]�jL=��Lx��UxE�_\@����N��I���'i�\,�D����)(��1����zi�>iᆩ�\��3�V�v�3a���(���Z��rm��!N�ѣ�
ώ�%qb�H�0�׉A��z�[�  w��Ӂ��W����A����qȧ�P���ס�I@,�'p����Ig����HrYK��?�7��7r�+ �.��$d
C��Y��+��o�7��8^!�1K�T��x�3��(����K�o�L�7*��3�=ǳ��s�1�l���X�5S�G�*�� �ܟޜl����+��{z:�G���R��������Q���eQhᤫC�Z����gFwu�6����6)B^g�4�;h�H\m`Mu���ĺI��_�Ҿ
���e���V)��,��ʌbhaTsNw�?j�?���q��D��[k.��>Aա;6��w��)�5� Q��+6��׺T@�Λxj_S0�:�{{��hX��1y0�d�jB.-~��2� dc�k17ͦF$ڗ��ܒ%(m[V��YxL ��BL0繠��N !�&)M5~�y� �3J�QE^�bص��+�%��`>�@��X�r�x��/��Q�Ɗ�d&G�<4���4�Z�}��?��з̙cX<d��?A��v�KI:��N޾'��EA���+��|#:I��K����{S�:F��c�k��C�:^b��b6�_;A5;�{n���[�G�S������2����\$��A%a��xZ���W�l�#s�������!���;��(�������N��#�iR0�I-O�10�)W�H-���s�y��#��z��)�7A�m�����5⾍����v�mO�&�$�Y��I����RY۩�>OQ}	|I�+��0���YNP`�r�Z��X�TT�����2: �W���X&�@�y)4����}S�_|˸{A���$�,�L�I���:�)n��(�fs������Db.����v(J�u����ԅ��(#0��2�R�Z��`xs$���$v������^Yr�����D����*����^Z�N����Sy|��~�Ù��꾴�I�FV�����8��0때"u�Sݭu-X 0��TuUd ��R0�Ɣ?�"c��OĂ����T��D�+���fG2>/���Jw��e���u�_������;{�V�ݶf6�遲�Dn%��9�g(�Н��|�캪^	I�VP	J�I^�r�b�Tt�:�GٕS�W3�m�2=�$���,
w��ǅ��Z���L�J8�޿O�e�����Pp�i�сvO�k����������8��x���a�֩Cf�(Ɖ�j�ٮ�BІ\� �(��BY���
�O��YE�4i3#r��+�u�b�yẌI��O�5/�QI��юIU�a�i�Y�b���� � ���9!nz�ø+�}a�f^���s��x@^�L���Ò��l���W�h�)8��QwL�Nٜ6T.�L�x�~ڊ�y�����Y�]�I�(N7t�;QQ*��pz���	w���z�F�`������目UUQ;��b�n�p(N[��9��O�Sz��,�LAS���:�OY�csi/��U B�c7�{<���b�lt`���zR�-���5�(�4)OIo�`}��mY��A��a�g�4�|��2��̾c�T�KF�Ҡ��"�4�8�����l����5��F�U�}�K>�*b3`j(��l�_�8�nNx���'�3���K7���FxC��a
�E��=�VS>O�`��hM���I��q��YF�&�A&V�:Qq
�'`Sʼ�K��IY����&��/51�<� G>���*�-�>����#�4�9�db���oy��/&��?�BjB��k��[�i�D�����<�Q
�<�[#ׂ@�"@cn't��Y^�2��zޟ4&�z��G:�A}�uX�����؁cm���?�[�Z���-3�Z��i��"��k�@��$S,!�dm���#��p��=��i+�aV�9��638��Q�a��jzM@S���*hNM[GOfuz��a��od?��r��jU;X��
\��!j��5��(%B�1�12r{+ؠ�W���3� ��	��ӓ-�'N>�P0��Ħ��Y�Ub�; ���� 9�/��4r�ޙ��J�]����w������|g�4דG$>��Ub<���]!1F5ߖO�Ū��'��}���&	�
��(��	��F`s����l��Ch�}. �63I�}��'�>�k�O�=�y�D�/{>Y2 z/��͛_�@�-15
�Z���;oM2�#���pם�
K�P"�d�ٽ<q=�l_�u�F�ҕa��ؼ�y�2w�,�8��TBv�[ĔH
 �/}`���?��i�Q�"������k9	�;�c���<N��?b��A�oz޴5���𛟏���̩E��Z�?���8�dF���DĸgE���g)��O.RO�ܷ�7Ǫ�f�H�z���˿�?��C���Ngz���3�x���}��t#�S�"��@�(��®�����/0��V��1qh�RM�^D`�Q�vش�쯻� �F}�(�Y#Y�Ն��XW_����wK���U��L � K���7��Ã����H���Hi�b!��V��p;a��s���q�!:�?����Ⱃ� ��+�U�#(�{�����z� yu�^�,}�7R�w¤<4�ؑ�%f>us�A^����r������ r�06C�x輁�n��9��Ia-Q?8S!�H�ǵh�`>� ��T2����ܒQ��zR�����H��2e:���mX���ӽc(������To>�6TR�8��������=^�ܐP˒�MQ��ݐ�hu�_�Rl�
9��e�d����}����^9y#���º��iL�}�U��M�gjI��2[����Zvjb���os11��ʆq4q'+���f(�f5�i��p��m��� S����e %�������ƃ��M��%Z�˗��cj�����݊�K΄E	VI+K�f��,?C���*/��/�rs��0s"��[b������_��������dc8͖r�+��ă,-�?��#q����	iIk����*v�rd�j�>�7n����``��rl�����`�@��	
#%@2~�`� � s�̣.��6�:�8ǀ,�Xʰ$2��0��}1C�_�/��Xa�e������,.���6��ۃ���Z����0�{�g8Թ4im1��9��}+^|�9�z7
�,M-������:�}�֦NM��B�t/&)!s �;%�A=�[�`�������`ZI# ��}��[p6��Ät������*�����^���&��,Hi.�vlfa���"���;Eo\C3w*|-�
�P��!���Z�TP�	�͕�.K]{n ����2��/G��͋j"m/[ipCƯ�&႒	ih�1��FI1"$����"��u�=�V$�9O��f�A��ԓ?b�`���b����Z!��ſK�ʷ+�Rҥ�dZ�V�'�Z�e�g|�9���I;05�-���B>�,Wk�C�z��x�ԭ��(��g�̡�(:���q�
�8����f(3�3(dZ��r�r�um|�=.�}�Xڿ�o�W[֨�)a ��L�a���z/2u�˚���;�'tJo{�L�iZ�6�{kꈞ���\v^�F؞A�5��R� �����eߕ�Q��Fۅ���IЭ2>헔�1cI��Z�u�^2�縈�6'6t�d��(��z��/�ͩm��+]��4t�w3�sl+e5�p��o��BI�h�M�ɱ��@d.'�hI�zԥQRi�	f����a\�q{��~�XdO~�:%�����{M� �M"K)K��]Q8�1!�1�T���I9L��=� )r��m�S~S��Uh�
��..���9�T�"u�	���I�C��|�����b�|~A0A��4��i9e_9p�mA0���r0c�]�O-(���U��|ee|j�l��K��Go\b�e�u-ﷇ4s�H�I0Y��koN������6�w�,���J����C�O�կ'��L�-!�����(��
�1�W�˾|[�w/��&qX�:�Ƽ�q++0|h4��ކ���I@�w�~���'}�ʆ���Xf�	�)��4]~ŕ�$$��j�6=tp���6�u��2@ꗡ<�}/�-[ݰ+�ݰ+�mZ-%W���߹���]�18�Q�����rd��գ�e��h��$��J��ͼ����T��m�.���-�I����@�ओ1�']�|2���}�#n7И�q�X9��ׂD�H=�	´\(@󜌩j��������5�f���xS=ji,i��*��<��O�o�p����	o������l>Ʈ��$�U�{
�pG͖����8�m��jb�\�dU��Yk�7�����Y5=�?���p���κT{�FC�ߟ�̬���!���rV�i�� ,���v�n�m������\���̴���qGի]���[���s��\�n�:��ҫ�Z��gܜj���y�Uk�$�=�3#U��P!��Q���-�F�Y�)������f�� F�2��J�!nfvLn\&Cպ�C���S�[ꆍ���B�F]��]�N��������(5}!,�<H����.2�I��5wX7�`�$�,6�Nߝ��}P���>�z��M��Ӛy_}�g��b�����W�ΐ��{j�[����k`w��3[�c�+�>���c(��0�#�>|���eu{Ф��Y��F��lAwo�UGO2e���U�lk��F$����R�>

Q�$(���@��B7�-�'�Ǌ�%�Շ���t1���B��aF?C(7X��K���u���VQ���Œpq�-TH1����I>�:�Rp Y�콻�!dЅz�iLmU81��k3�f�esp�������/m�/�]��Y��ܕ��;(�ԋK��Q4�,Vz���8��a�l[z�0Ϲl'�tXuz�7T��ev@��v�i2S��=��"0$䟟"�	�\h'�:|�=p<9���l��y�"�fC��^{�ܣ�˞!��v��ܺ�4FH�5ex|��t,��u{����D���D�Z��-濚Eʞ�|�#P��>(�D�A��0>�R�e0� �cw�#Ao�6v0)H�B+2�+Ɓ���4�(o���Ey��B�;��u�]�s����/ʋ}��|l��b���QDZO�|	�C�U@{e*�i�Y�6򘺑�n�U��� e���,z2+ӄ����e/Δ�l�N��l�od��PL�uo�\���AX��J���&�d^�h���ہ��(/1��~�&�y'��E�q:2�<��+I��b+��N��M�^�i�M��ncIEz���쏝zT`�w�n�OPq��zE
��*=�ܭ�6�!����a7S���k�<{6q=A+Y^|�#=�࿋�gchv�ቧ�e��\|辧:��
��JC� ;��?s��Q�=z7��\�莼��}�da,FA�@�X�����~��彘���[��L�R%	�©�а!�M,�ò	Ӳ�.��j����u��|Sc�Z�wSS����Ͱ:�a���_�4j^�5qV�zC�@��̊6S�Mh�A?"�C,̞"���<B]l7��$�h}�8�ׯ׋h���6�+��՝h$6�)��z
��BP��>�`K�
^{Qpl=bJ*ҥ9�5E�O;�S:O��$��z8c���Zْ�9]��ό�(e�I%S�A�˩=I-X(���\�ct
'�2����+*�}�'frb�Q;C��c��keg8{E$���bt�	���S�hF��5�zaCu�Ɩ����b��6PJ��c�HZmqh-����iPW�ШҶ(y����c�k2�ֻ{�lN*�~9aQ&w�؆��y9�[w�?��^O��H�lO&2�:U:X����٪�򵅟�8G�WuF"�Ƿã��y�Y_��QU��v����O>�l
Jn;��ʻ��lL�z�W��b)Z9��:�7���M�����UpE��׵Я��L��N���>�����A�)�����ʯ��3ۢ-{�cUM�e�QOb��Ԩ��i�ߏ���QJ��Ҝ���L����9y�>�*4���۟WD��@ek�Ϣ�:F��<Ԉq+�;���t�K&��N��{Т'c��=��|�v���x�!��S�]`_�0w��d���$��@��J
��`#�r�6p�
�� �2�hHT�޶=0��h�ͤkD��#�r9Z���L�+*��R�_47��><�$S��ϝ6,���5��,d?�.���^����v�O�4;�zq��єe.->���R���຺��j��G���[/P��uW���)�h7Ӽt�d�"Ӷ� V8�7��Q7�sdX�עW#rA1'��� �/�� D��Q���Pp3������!�k��h��hTB+�K�{�u�H��v��D�Sj�4��Q�Xu�%��粶��9`ry@��K������ ��sR���&�����L�#���NG�Swnwۯ3Jz*!<wDX�-��t���V��٣�}��7E�Q�J�8�le�}��)Dy���eP8�_���S� i�Y+��A06�16'rG6��,�*��V�/���������C%����z���^��+ce���s=��ޕ4�Uq�
ѐ�W�7D�tn\����$�T