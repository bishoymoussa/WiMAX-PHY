-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
1gI1LYT8ADimwzzSjmeD2TUKgpUKHjG0h5ksTswU++flMxvCCuqIs1fe+YhIoG2T5eYE3uvtWCQW
YHIE/IJKCbiu7n0YPKjSN1MzgcDw/GVaBjbkPkD5UbPEHy8jz1yJHBiRIaExWm34501fXo9MQ7cI
SQgIVUXTEnNFedb1RyXEplkpy5KYa9qJVp5at7Y3YUTprwJAGKerfvRZtag5yoBc0k4xRtvDz3xv
Jujn0PQvXZ4P1/KictP7OFRJKPMTgwAluBaxcwe6ezGxkR48Or59iVzM/H/fM9R1jl9u4E8DrQK5
p/q+DVrEAX+LbzU2v8qWbJ3fRVt2bgV70/QrpQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 82048)
`protect data_block
c8yR8uti5T28gUDsE4I/M4tZOwz8aS1qFOdsOLEiqDPJq+Abm4iUNuxebAHX1VLm/s5ZE1C8ZZD/
c9bqrFe5YjNdE2FZgvTEXVonDjtQLyK1VkWVLQrCrSnfAD0N/BvPnk7Il9eOdyhJOAdLDIW4TrDX
g+YTqgZNBeF5DBcU5RESxXFuF+W6EKzoUqcGQ0nNUj8xFhRPZX2p/Ora+7mb2qmw24L8t+psXBI/
nTuVAs4qYDsU7x/AWTTLbWM1xlc1Jsdd6Lw9lRb38JO27gxxMT1VuyCTfgacFWTknucxeUYqc5Vv
hGb3+h+6/cSQHumzDoPES7Zta3I9x5NwsFpktqs6CgNPy65iRh0QkB6rM1Uu5ilwzsWsUvVzHM6j
eU5zjRFj1WiPvR0TNcW+o+nksFFYzSBWJeBMXda9FdyHpx+EXpajeKxSyz64goKdL02Gb2L7Ne9G
rFx7YGgwXehbB2LOUPUyywdNBzvP4YQiaabxxRhPSltNDblC7SPw99flC4i2OO+iztqYYhX7QlMc
jDSf3sk7C53in0J2ZB/TeCYrq93MMX09Xpk4072XCUF8V1YAWH59h64r4err3qglVfoOTcbbHYGW
c25d2ErU1/zqXviXTCogrGw/slQUhWx9S8El4E9UZHbTQ4loBJ6iU5v0Lyztj2B1/tfydOXvIcnC
VN7F4+ingqLg9aVrtntWOIszN9ROg6YYxDASbMlNuZ5OrjTvr/71/O8xuP9RQ3O0DIPkgVtNpCfL
Wf9y0a/qyOI/UmXbY8fHTjvXfYlzLynGW+Dm+0HP1kzGqBk+8Gdochl2LMCxcIs0OaurvK7WxeXu
1aM1iUYAF0AYqVCPAoDyYCgRDEKLLwkn03NGM+rJ6t3pK0MqjS+Q1LfsUjN2r2JunmbHqMOo6DFl
uOcv3imqQZVF+PQGeGWXw3gnlGYnd1vtPzPMmRqZNpK+QPzmfRiWMJxaMnR+bMYHkqYWa4UJT6cM
G9JvCw7HYmXi4KhuAhKqt9mX/GrSU3s7aE/Tpe7EoHlhHt9GOMgCANShxOWGt/IfhZ3u+uVi/d/z
o1rxMB/ypSXbc8yG8bUqG/yJfv4B+IPNTMlgYYf/3mVNVNOxPPhabpkBcxOskSIxHJC1HEeTLLuX
deJHhNlgwiRoLh3goiZOONYGr6DILG4AEpVWodDoAO775VoimIEZ26T1sQ/oJKDKRJWW6AG6myOZ
0LjHKgpcadGVh7kjnJ3SOtkT8E7JemEnyM3oZn1nQoPQ7kIV3EpWNwPB27f81eOt9HSsG8GTk5CV
BpxGGxRcg6PUJJDuy0A5W2mNvyU4d9ptX6ZyK1S7KUdZrBX+4VUIzVsEAaUV94UIaq3fu+oA9Ykt
OAop0aqFhi2Lxw/miA2wer+DCFTD9LrB6O+HpkiD4Vzdj7ly7X5kORRjldiD6ri3Sg3DmnNUV13M
wikzT+pqvRO6NIAWX24EQfPgm4aRXe+JMveXU1Ww7fmcJb7Zc66d+YCjB3BYSMS7qCB3gw1l/g6t
041YUmPD/Co5ByUFbwg+S0qgd/LZhREvc6kjv+tuiCUy8wD2RIBrKYNTdgKiYSFIoRGwzvDNSnmd
AL+DpvUXpe9mTTXbDrszKgkDxC8N1UPPDIG147XIZ0Yu9GZmfCPqbnpRi/4CQdZAkp+Fk8Bwp9GD
+k/wzLB0bnylxJIhfOoB94eszpvyDuSy7Czc3L2mcGwUeHL7e3oddKN+Wq9lc5GJT5BdcFecfvrR
Q1O51VjxLNajJ6iFLIKv7tTbt0+pZuataKI2ho3cKcx1eYaBlvKl/JS8A3XHMhunzij1oc9oOOzI
ajtCgd0vn0uj7mhBTdpaFTY7be6REpKFkhGbBNuUbG17VoAkaWOEgECFhwSoyLqEUL3armbqZAnp
BXeIDSTST4ylKVEVsCHwtWpQOpeRBA4qCkVrbW/v1TvbVFpFBXcW28U8eHkPiWJ9tyvCl43VmQ4u
mHBkHe7ds0Ina0lxnf/Agaj/W/HxxDUu35aYtUipfooKf3qozUujywH6sTuhULfnYCW5aRkdgxav
yyTUMd3eTEz5u64lgmYCc/yB/rqciLn+zOEZu45SdawZeP9vRM3K/fQSjXndcsOsWtvbnbYVcOWn
emvxgSPI9oNRObo3ZHIEO/c3WPCHlfmexn+KNu9d7v06KJlMx/HA0oRmXc0ZcOx9Uats91GKRY2y
YsaGlTYok+wcOVPs+1mfWppok+CWfA0r26yPiAHkGOuejcts3GB2+1RLL8z49bLCgy9FXnhWBh8I
94cmFLZGr94q1+6cp24mYkkAIAsddoh4RYap4ttp2NCQO4gTJy0xgxYWa7cRREq1VedaMHBaV/kz
MPb16iZqwofBCCp0ffji5MWIWvW+2LgsRIbRW0x2/VCADMcWBNHeiFanpFpsmz/IMnl0WWqOZ3yB
/FmH6osRBvZScoWhon4NNwERmXUbr/sL4UPU0ppbfODZraLKhDH8rgDv1P8TVqizZW27xCQbnA+P
mi5Q7CEXX1uYlSFbWp6x8bFb1V9dw5IgpYEEbs2ZnRQw8seXfWDEI83yeZPpRAi9NL0heLdk9Voe
TuW2kuJVvFQJyK8C6aVYzTreLE4gM5DNHlq+l2ZeywLK0pcysPWnYDbGpIWC+ZmcsVdTWUM/RdmV
vMV55NOT3hmX4TN4ztYlYNYINCs7+yjb8eb/36ZfQieJY0AvFmWLmU9q+f5xHgXCbZ4uKpbSv/g+
CTKDCXrwDju7wTSte97CN44+QXybxaizmS4eBBKHq8EKh/od9pkDQrQF216JZvT9y4BsoL8v9GDJ
SEYhBBSAExOE/sgPxeyCHKb08S8O1QwMJY0FqrSrCBtZNfzOV4g2x5Jfr489bcCOfPVTDL2oaiUB
+HnGqu49q59q/Edvv798tSnfRXFTYBQZtAL1h7eSTwn691tmDxRRv7lrJ4O6XDZFt3RkIWjdj7ZQ
4W1ReBb4BZLGY+7A8JZcauOMfkpPSVkqCOrJToDM4A2zdm6QZa001laRlcJjQpnyfQCcYGgV82yp
hdGKu98hghx0ZC77yeZYNnOu6s/qNp4Sn8o8oRJjUdH2afWOPC90lP2DKoY3+Mhrc9fsFliWLSkx
/lIej7g3REYm/P/j9D8S5ovcphE9PiDPdsW4C8GFHDAgfT+diHxNy+TNB2viZm8AAO1zoaajyxdX
uRZM0lnmvhdvkkAI4svYJv32b93VgHPc7SDnMq6vki+WuThBw0spd23DkIHW/xWghV6Nn32VUc0W
4Vy6ZSWnHUnIHq+acGsbhgOLw7eGfWSkRZrGbqTqEsBCceVqJrCpBuGQcITcFyAkNK+1S4HO6kPh
BIM05HlOVEeD6Gq9pefo5aYiV2uAOuCXB7HgZJ5clWaJND9gaxWjWh/TdtkIX36tUJKWGrZhms0s
VvYr0q01oBby3BYra41PSSMj+BE/LgOp57LqU9Con+P9XBmmwf6upHwEF7FqvaXLNvzdAfo85WK8
n7en/kTXBKQU5HeaAbOzMK9JDXfHUvhm76IQVxVrUoOFYNYySFDyA3EKV4iEVgUyAnuRIm7ScgDW
vTU+sMDZ3+rIiLrUeTiiJK5xEZZZI7eniUkDRiONU7AzQ3GAjPL0Y1aSgAsLXYjBJ47Z0GMPy4jw
g6rOHKEv+BwGm1pqBaq94jJnlBrx4Fa8oDvPAR8yX3wcEIDPOUp0ULKhviSEs3sQ8YaEkHnIk6TA
mncJnmJ1sOi6xGR96IDt6p4pMToDNlbumNGid/aPHruMcWuRWubPXriR6+9WvD5ubYVOnibTZf3S
Wo7f7hTq6ndxOIpTCfptHXLIXhJwUlN95LL7t2Dz4kvdXJqhPOiAgR5I3Bh4eBZ0LLekcr5LQf4m
Dbn1vuaUdSBhI6utBMjP/FlLr/ZYdvAwYqoOQ5PHVzA2/oEz0DO19ttVjdJzYBFYAhpLIZNQHhN4
0pS/0qZS7zz/IG373RtMmZw/LY0S+k0P1ZtaXjLuqeM4536xIeMW542cn39cumFlpvXtPRDPXkzS
MjHhuh0rfP3z7I/PKGDQrCQUutWYGI7YPK4EflD6hWgFwsS0m7v00y3n7hpjCFwJ+GMYN1mRjJqd
zk/qlo6B+cmp9POEiWepnknnwxE0fHqs7mhlR/1Pj6ezrqUB3I/W8qbJ7WRtHQunWPnycX+5fzq1
KdGAV8SPTdkMfPZ/cwkmrb3LLrhHV5ymUx2xlwSogGGcinmZTxOJQb+murE1pWuckazg9KIknvz1
RI3ysxTiTbEa4kjsikmZpxzqXg7p4inlIyk0Ca9VRwwDCTm4mVRFJWOZH27I6kgjwJb1npZ2tAfG
S3AS9QQPeH5j56w/v3raP+bWgIqZWzXFKGLHhf9ovoJINilmc/zwIP9uhxkGvs9bA3k1WihGr3Lm
C9D6A+xFrJ8wHuSRr8IQHwSN+w93RsTpq4M5O+ooV2bua4pUAEl/L8I7cDueFsOr9Qe9NA70CtbS
jXMUY5T0J1dcHL280rJ+iDLhD0CNJG+My+fYkZmpTFGYL5XEPZH/l+whYhLRJChDyD4I6wdClPHj
TEFz5IJmC7ap5XgbwkIcOW981pk5wvUVvW8EWVe7pzf7/h7hXy+sJB0XNdyduB8IOnm7qrxiqFCG
HyIVUtcFb/e9l/+TH6wXWt7ZVSj63q98U8npxea4k5fuBOQuBsQ3CyLXs3KdPqoqc/BaQVnmO9WX
YHLUrFCe6NIDfJe0Bl3/D4hqDSiq3IHffF7yD3OWXbJnOD6Pzkm97LoLm0rA7kau1Ia8yfExRIJE
OtAbYXhBbZxvKcEVaIza6d+IWIWgPFzax9VaQ1aaHuP2SRB8euU+mq5FhSxDwIEfQ5fsO0DhSQBV
aXJS9ZyjGklAL8GI+Dp2KQ2ULXNRWlkZJsqrTRMtU9PgfDZ86NauoimZ2IY3PZMqjtBuRqWBS3I2
WRCv+jK7UfvJ08Nd/cvhlLRAsLU6uPnWsLBkO0Ytr5fZOS6NCWMwes0dY6yWrIvfvRMW7h5/mg3z
G/NnpYbqlFNqENi07uX2AJqamEeZsi81QNLX7ClmBn6+KRPA/nwOB39HeFLsGfDIxtQOphuSDdHe
1RjJsoWhWKT1dRAm9YuxjycaKzg5tjloavhbsovqAKf4GBzpSsWjtnNyneYhX2Tn2O5mnSE8hAkS
IqQ5nW0Sy/jUjOnMlUI5jIo3oxhmzNxYw9BUVlTjRUyaEvKsnn28xh6AKmbIldzr4zxNBxGw/bMF
bt4jPYFM/pH2Do6zClC29nXI9bbe4al+txTKwcsvvYyIHYN5oKQPVKuJ1wOXqpLJSdYc6VyeQ9uG
eMYrsUehpjf7Y8Fghzwp2odHwYpfO2Df3+iHFz7bqfZfi7K1rBqjQYwxBU1S3kyYsW1pnHalzDiX
tCzZS44zZ2Un+OV8+FaAbiXF9FCq2kN6cXKr8MWE1LqfvFJGsoh6ePAIxHfyNBU1ALHfZhAMrLoq
VyGHNpDfCvnWRfpksUsDyL6y9OGVfP6A+XjwnXRuLHU4LteVo5YAA9dchymoMOj/U6zFx1AQ59X1
U0JKeALV+NayZ8lncCnEMkNN8A/MQk2K3rZbX+sk2rzG0V1MNg8fFQVZyg5F12OZjel0NAqFOTcL
HOk+37ScBYzFyk1ewlExrecl5+ANTuzNox2r66xPemkcy7EDLvcxLA8tvebpRTgqajpJdHIRknbZ
qWnae9ZHV3zvt3WD4VbzbVWggevTVSkONIvHrpGl5Xd/L32pyrvM/Rgiaj6K1mC4TSkyPtyA+TvE
kz9KXDayE37zXcIm0EZmlVSiurt/mkt1n1zPx6YygbX9fiOmxBky8fj7qGhm0ZK7M9if2daRqjXm
5BTQEfU2GVyOwvvgP7p3ONDJiMsSqtqhx8QrL9M1UOmN1vf6Beklg4MXLuWPxLoNSi3d0bHFKme2
hqxvxtLW1pfLJGSvlfD+T0zdcumpQZ3Q+pTE1R8J3Q3o8k2JESfYhRSLS0KCfMKpTM5ZMiXOs1Zh
zRMcM9mpSYn12W+BI1GA8DlQ1B51aHNHd3W72vEt8QId1+x33sOzgViyUmhy3MtJJuyR96PuW5yW
FhKYSrmogC+v+yUNf5VEPIzgrS+sKOQ9biDRNPU2vxRctumcNY/AOLQt58cwLmqcQbKxIoxboy7i
aXweMZxnOLFesNvEEo5FS0+fiX9laxlePB7KzMzVSJxLm5MYYnF4uGEQSLpFDyvIKbc6/Q/X33A2
0lPjSUCCq77G/8RJ7cWyQxTPsjs4+gKzZ88wHNKfEBk8wE3LoQIaTpwx9M2ILSe5npfxO3axS7dp
N7Apaw5bCYYsfr8EEbkuhB9//dq6rYehxSvVEDhNfc5tBlTAcZrz1N93DpM+kdBOipZkUByswLiZ
2j6+p4hGLC/EZKgI6dJPI0Tm0OyfsSmVbRu8YgI8K1HyfYqXmGUgy8VwSXtJSbViRac+1z5LWrkY
WkqGDFKcBAwLM6bJTIEBzikWAEZg1xyFK6MqEuePDERg7IjKs9RQhjukdp14V+BeUj0HYqXmWMsC
3AqgCsRX+2O3aXY60Rf9NgIYXzrSe+AoraNyf7bzSmqgQMBa8dsPNgh2WkbPdbWtpm79sRAcdfiF
WoOIh5FcXe257aRtljXoYWUXmtlq7BC6H9W4yp6JcLT9O0JF7orWi0xZBOKsrQfp0RTfaOC706e9
fiMMt3r5NALKaG+OKq5P/6O58Rn1NyFJm9E5saH0p4xRJqc4TBO0a5nzoLsqc09mZEfaZT1fSIjg
J9X7vWkUbC762BB9bThySPp1dTrjevhYth6TcUGaE8C9ufmfkrvuVNhHD1rbApJiAbUSV73fy+EU
Xd+zVE5HqeLaHfJUg3DTgSi8U/Uh7eQrg48wPy/kVVV0Tz7oyixjQlWFHYeZHAHQ4ISyJHdb3olK
DzOlKVPlWlkW22SqjgLHzuKH30XFFAF6aFxiCtUZxNjA/h+uW8QLrT7Xx9/8ymxnR98sMJPBKDq1
GTK1zmtyDK3JghY9F4TJebKgRk+msS1MOzhKqG4TvPMq5Dt9GTbRduHQpkDDt0evzdHXYW+4cjXU
J5yOSx+MOjqu/xVanQJFxw1VlGFpC2RnqU0mjpiUIy79HK9c/8aM97Cy2iqXarS6bqGwx/voqGej
A87P5Oegm9H7BGAl9DBDw8+Ek3vUFh/hLO/rAKdtZ3cQghOWsdDIZMJClc6DcyygrExHnqyNcvnK
M3mcrc+ncBQsinQl2vId3iCXq6jpY7BCFvkPhfvhgptsQPnqiYo8Kur9uQ9uVRF0hlNGEYYeHfv7
Gva9uqH2mBVEKyjX57nw+/v2dVNZYhCsd5sDpShYbsmjg8S7xq8GP4/XKaNZKty9BrTkVbHHx1Ip
NQVLxslXsNNpOoxjRZi5rHXnyxAiMRMXl12zdG7BMYYvb5/blj0Xzl3eTL1ImcD9IjJ/nA/H1fmG
ECeWD0a1WfX8MQ2WXVuLe/05w5wVJQPCRHbteKDLRKDRtPm2X4+SZEUDnM/G+FkyrJ5BI2UeiwpB
+BzEHfMeA+Jr1qtwgxNqVtXWy843T9dPEdQUeThB2vZzT6U+twjMmEcEYo5JuAwVOdBWp9P3TT6w
ngGbpSxgexznAfn2VJBtZyv3rp+Z7QfGgDAGi08HXu8xTOPfq8eb+JJRHR9mLgWP+YaQPzLLLcIJ
Yf/IXwCZjfsPOdWA8/Lx04nIfh/5wdFqMIWdIzttb7YnJsQ7Gt4MVnf58T8xwd2j5n2/hUVlca85
Dd7fIlkG5dCwZZAc9wUZtCNXDJPkh3gmwPfTzX95iATlGblwR4GNNoG1nrKCNcZTkqUAHNVlQ1ae
Uvq6ZJxlcNN1HEOudI12OjbesL+BRCPn9BFCoxTh66vUNwfgAarYyOElpDRbp/0pBN0elnvWuWj6
++NjlhEWplz6NAVsw3LN90rOzB43nUTyxLK8L/cRJZwi/16/+3YYAChutX5htTODtEzoShM02byr
w3r23eCVSjv7es3EIZ4ofHl3IeOz/Lx6PpMBUFyeVt+jfbjNWKHpeRS3BrzWyAGHQD9h8aphbD86
pKNNHnGk8pQWwFlE9g/4mlpjRSdgyj7GqWtjgPRF5Culvh/5z0/0BzhkWsTkORPMzgqhw3+mJTO6
bANDe/OxGcBMN2AEIlSKStME5UoY3dRMcJA+mZSD4q+zub5ykdCvZVFXWwPg8z5VOG/fF0VDr0Qv
aOe2Hpp19GdrXvpkvcwPdwPz8Ramkvjs2lGMrGjLBw9/tjj+EEcrioxqli1Z4y9i8N7vyyPs1sLu
c1t7N8FitZixnfwUT8rdSPKHU+XjyPpJCIvIQJrRXtUCpwtk5HU5nf4N8C60EhWIPTG6UFoBwJDs
JJJ/g8/8ZTm2DOnO1qcYpqJSi9XWUFIT3SYS+g1R0quXuqeu26YETXQw7RIpQTAzdKH2Kt8JuoKL
ZHitSnsiW7kCm/Ya1SQoeCtItMIvAvlnNr+0czvPoAnEaFQyT9d0/eUVfge/qqkdZXP03v7lR+hI
kI7Kiy96bd6ZNHhMrrcDUxSB/FrwupaDdxfohB+pMlFZDINtiWQtHQnhKBOyHwCxsBVL3U1b0Wwi
cHg+6xB0r9t8FLo81F+l3x95sAd/Ccaw8BnGtJN+FDmtRHespWeuagnWHmeFw8OmF+Zoy2oxnKSB
ldZUvE0EeYorn5QMIMXknLUulu5lfkh/jHFixdiXG6m/EtiGBCLcyJvtBMKIpjT4bGCckGiyQkTj
sxIBFX3olt+t2rXIJI96UrV7Ixs6Dqczq1CBp2aBag7PW7p1jpjoOI4Cg3pJEBShqQ6gfum4S0SP
CQPt5/qectrjvlQ6J70Vk4nV0oH+hfsia/P7N0QxKdmmekuj37Z8H9Sn1FlNKk90/LQrrfD1LkFB
hDTw1xFBaCrzkQHEOYPvVelwx5egomhxI8gteXQGXkxU5x/OjS4PPL2Phhn8DBPjjiwAlHHznrZx
P1PYmx+v+Jtgs2GS8EluCwufQxnE5AW09vb/Xw4V1mKugjukGFv12PpGuXyOCwgpRp5afDaxx8Ls
Cc/fmy/O7bBfzOkmVfkqJ9ZVMRqj8ZzVsSkKiXzRKyceVFQ4M6ZBGEiTL+vjGIcNM6GWJ+3sAuAP
M40e4+hiArRYnLpuKBGj+Sr6XTOLeJ1WkHBk8MTRrGNdkZ5IrOJ1ROPUjqNpIL8den11QyTcYgTJ
HAS0D3TrYujJtd+UxKPuPsITiIK28SAqqCuRjXxPtNpgelBSugB32Gp6Jr86lbgcWwQes6gDfc9w
4Ou3y7A4o9o12zflVHXDAtFA/80WoZw62t9iQWB0nYNaKPengA8X77yr7LdLryVN3GyEc46QqWFY
uZqcRn6Zco1KTn2OjhSQjKQwIxDBIWBYjIgnGAKeMxbs4eHkosx78VKrR4A4KDYdtF1zA8U4uxdY
U7bDQvUJQAMk4dFvma81Q90rEg0N/YCT6kbArqBPK5ZXnOXScsr0E4fqoJvnzdQ2HbuPiQkRaj7Q
aXl7EjEkw7fjG3ixPCE1gJECs8SKImsi5nM0rDfvCBNuFSYZCU0aKuqEaMWvt6xBIUjJmwHkWPo2
A6rbCVT70vOKnKhNHSIt20W4pREGff8o4zPY7HEnBSonbbC1m4GojifewQGkjpOJYM63P1Y5oJaA
wK2pWAJtSZn7PXcr+7zBfwy8T3Ho/bGzxRVn9AjC+x964ZnB/hrtgcq5AywqNUnWMwz4Yz8iZe53
dEkuXbVP2OyNjLTq/CPXTwDAndvqIwvi1IdSs3acs2LBMFyZ2nbqAnL4LcphMfk4hkvx3DnpmwaE
OVVqYhFVPCHViOTAuwZtC/apJwGYgEH5PbbYjLSbgBXG9TxoolUSC8zExnghxhD+WJZ/HBVh3xzt
KWUbWc0lSAp6uydBmdnwQTnIRbT8L9b3iotBRSLiWKlR0A4o39iVFJK+meeXYyKj6pjlIPO0B8H+
/p0FGRlnILSS3EH6WgQcWwY5jJNPRP5d3W2pIkszT75KQvvwX6Pq/cS2RrAn0CRmnguh+p+PQyyF
w6tPvctBlmxzAVBfOJ2xJZ55akQGQNS4PAJOPlyXj6E7Mujn9OQHlPTELe62PWLC2sTXfvy5j4B0
+iSeU/Ky/I0/hKpnOXtetUgSQwakMA3wx+BXKK0UtJyM8uhzBSyaLxEQ9DLsxT8O92sRMw7/Wfx2
eTVRABd9UivOIpUdT3Ubc2pf8RNiy6eNDZxoFBMJToBTdz0lPS76W6A3DFRk4ARjjA89V6Ui6A0k
9/U+ZkYbUWfLZ1PSzAky4HynY9Ja/SWCdrIEErssnbNASAxdbJHgjCxHpNcT6m3g75KrixvBx9Ok
/qU5pD8UNy01eexeTIDjr1eoE9bxc7fZFMY7fY/YJ0EjTwDcAdrvKl2k7tetnFcUdbJhi06AP3Uj
Ip2OOyWH54i0RCMHIEJFqcy3cHknSJxfX1RjZiRH5MwBnV6IOGcKqZFmFSBEG8batwLr6Q2BV4NU
VqJnbPC8HNII1PDziGcUr085bf65ocrnw5qufXuuox+dzoYPWJNBN/QxqL6E+sKOf87lzhmIUQZX
sf1bj+kw+F+xEGoW5xgSSa5e7PZwiHHLhARRwjYrR2l5PFIlMUl4u5pkLlLJ0Dlty/EhQ7/n/DZG
RCP3bXBzbrz9uvBPiZ6fIfo2Aqcbe9JsMtt1TZJjrJ+qtsPNwpKy0DZtEaGvqXS0GyOzwfQCLGfP
GcyawPFUWxTwEaqUc57wzaDAyFtyI4TIcgAfq1GQxsx309ltaJU9e+hAQeGxd7KnDAWFnafylrHw
3U82e7txEs8Y1n2MJwwLF/RYlmpBG+cdh0xm34GQUxg/clZB70uxc8XxAtDwhWKNl88UE50L8zTq
dDkDRp75+qNfIF6eOOcVll+oXuEp63zSXPBEtxlV/Sfgcyer1fCbFu+wquQCgLVcqTK3Zx0p2nTZ
4UiMLRKVv6tzab1VysjTrOPI9zVgDKf4iI0FNL6z+gO8elRCOaFBeAZHqkxcwjCplg/VBgkDrqze
EAMyzyiDs67RX1kemJOryo0q7PGb04sSb7rcrO+bG2LRi7lbkpwYvVhzF3YpamlsGF6a3jdmUj/K
VtlO3tDCbz6hG3sD5hPeIcDYtPiipPmIQKOdOcZaXoFtmQfmcijK9e970REVJqb58d1YvYXekciC
HiAcGuOAMjQ/Oq3hz+fe6xX0f0EKkozqr2dmQCwxNQ3uyv36PXTQfBE1xtogU9yF/RHG9g2BB1bb
5XT83GVU0QMABViGP6+Z9CtRJ/Xr923UgkgwH+7aWDuHwnTuDQ1V41fvL0Ou2m73AbBdgJ1Km7KL
qiTFZ57vuwxsw5iyrjeG3PYbSNDCF0VT9xJgbpIBezTN+fHtywg9rTKjQj4rlJAZgpog8PZuf7BA
pZJRIT/UUYe7QIOwnPQxr/+GivrYd9pxoOMGG0139uX6+85bVdjauI99UsxjKLIyf7ydWSwvXVqL
VZlBJNcX9MR/djmSLUtYTmDtRqOkM7Ro9uwbNtVoxV44WK6uHlF3WOVRqvvfrzTdDo46BpIozWyt
GX+E6Kn0VIfjabhuyNttkXO8erMDKU1YyIf6IaTl8QpGkWGYi09xQNJ/4tuxXBUg4a+BsxMX14hI
7tqhxKu6CfLOUfHHjF8mC6hcmFsS39IeEtiMkC1IWci6hBkZkADywZwh/PjlQm5/XCLtROpVmPuS
SEj7XtM/4YAgm8pZd6twAJRAozbDjQ8e5GjEa3KxnSmhz6FShXJ17NL3jX4q0/GWpULTcXpWyrzf
l8/48obfmdJcladzKqNjcyp3dlnsOxXL6Q6gF0ix7Nc8qEPSOEzp/NGb13mxTLc1ZLmZHX7Qfinr
YB8e8DK/VrjyS/GDmZwzVonP6eAJIIiUIW5vRLoeXG+E5Bem99Br3gdaaqhCsMWHiCmLi14THsjE
NQeasCVz/irjmchus7/uszRK7B5GM1FfNjqz++HRuPd6gV6TATKL9Oonj6UPqqWykpXMtrIs/v0w
w7CpAXJlmJc+1yOAjmrzt3T4qFS2A59Lx272Ej7lm153zn1kAeihp+AZEhthoLdLs+KvW9RrpfMO
lEjiM/B5Jn+NSis0qFfHsdV6XyiRae/eMKIrn8jKs5q7SGwvAdcw2jl8NScsrfF83NU8n9kV/PZ4
WHM1cawLHQ9iVTsGDqPjxV0k4Tvt+g58NlOHi2Mx+Cov9MzZTqyBTPXevXMoldhXHJplicS9mxU7
KbBbeckGOReZFnknIQudL/zVHXjPTthuX8br9ZjKLnIGr/WpoFG++lZrp/7RobvuDJVlgL4V/CRB
IRuyXlvBSFqoC2uFhpTL1AtVmqw4NgCzDjK73capTbPyfMBzkJmcbTegtLIoBSTG3jvL34LDbRJR
yGTjtY9phPQn8+yDO8M+LmX4Lyx2u7TKnHFp4bPHtomk/3CsJ0S0ujak0y09eHHHMI9im44JsYps
PefujfWBU8ANn4xROaa8EFGJuqELk54KsRI2xqVaMcEaiV1BgjCDcGHhGzqtkymE1aXKi/eSR6HE
rRmlsVBR/dL7LzhXkAuab/w+TvneQnOUgnjz1HFN2flz/yJUVpxh6WgoY+f7NfOT56h1+etnjLcV
Mou/WVX8sOLhLfxD00sj8TTfLnt3D+DfArM/UXEZVGosBs4KEwnqhfMQiVMB819f+jJV/Q/jQkXF
oFCQ/r/zhln4bUuwUsVd9+V2/8DkH8ji8f8az+QMZF7e5XaKiZR7zBLocT+CyKx2nBs99zvPirfs
HiaWGPaTmMQ6FVybykRlKEt9ZQIqa7EbNFsvfA6qHi/ZzikOtNwpznvFUbzm7uiVQ1pqHWVerjxl
uMccs4BzWxsODb2iV+p28R+f9kSzLN/HCZQWsnGjjrfRKdZ/kzqgPKYhF2TKn/vcendN6tuh/NVL
JyiwTpwajLYnpDiVQZR9mdu3f05Vh0S35eVJaMh+zYO7A6iUqniWrQpmix+HSMcFF09NafEx/4zs
mDkRvh0DFvJNyjShnMWz8uLTggkeS8WwdJO575MxhfWitzKqbD6fElGwB+Ye184GbLuGI1SJxuUk
gVBAFyZlSbFwxwH4oOeOmsk72xqx0euDsPryzoJTG0SxFBHNp5PMN8fUwObeU+FqgJLVg8wz96PT
xlKCMfoU3CZYkpivlWO7wVnu8BesWKcRt1lrQ9NwIglPTQmZ7WdBxKFEub9yfcohPR/dcNaW7GWe
pIJLXq0EgeOyLs/1zPE9RpgSsx/99i7gSaGb9i7ttkjwgPHgyjEe3utq4ylhOuUgWFz+0FtFWb7W
tXqZmw8DesCAEx7JOPD5acM5X3T+N8W3I271qzP1t0RxIj+cbXZRw3L/tPNczKW6QgI2gvqxXcTJ
/8GFS+2Homc+f0I0pbbKXiFMZZgSJJLaNvCrs7msTVdnYlSf+aiI6VcwRntm1YtEUoXHaDYLEeON
UbE8MtRzj2pOPdrRvk9WWeV3PkXS4GBNPKMZy9ypI4fpNCPQyTMxzNEevLZYvy4kKwmAHoYDK2GR
6lCkDv0UzGFaXNrouZQ8hcbQBcNzD4n0qd6mnGeQAvqUyInaUJe2MCpQD1GBhi2nTyX1qryS2A2w
xFpKV2MN+kYIfyYV312Bvuy4DHdOw1pS5/GBMSZxRh/9jcmVY4dTfgXwB+Kf2UzyMY6bdgvL1cYP
FK+Epau/ZZMOwp208W9uAT7is3anopVQjwvfNNuZZ2mxegYZcagx/Qjq8jSidTxNRdGPAdKO/XXM
n6gef/9hbeyOsMUGVBLVlS8XhF5tXmTc9AEKL9+ugEWZqznnnsJVvQ9Dz0DKYeTdPW1IbxZgmEPT
jacKgopZBXHYM13byYvRbE6YGteyeXjJ6HsVKYAufxrdQ/fUl9p+3WxRFlKiscK7Avjnr/16i+Q9
Lkea46uD4Cw+ZE7m+D+/ZxITq/eoLnd22Btb0gOYlzlsU3rwmKgJlr5K7xnPocW8Sid3UprqKWSM
/ohAY8R92cgkUkdOtDfOoeotzVieY4aOCfk7ryTbwsn08GTIxkq291D9gqWZKcuCCzgDc8KmQMoH
1EyWuWltaVPHcCrdREmYpjoThC4vIUUA1uOZUh2VKczTB5hWGH/mb5sY4pbHwr6fF7h95Rb6mDkB
Xg3HckfaqmdrgJAJmY6vjDBhf35SVOSomz0+dFDyymNTBrkavO8cQg4MZSzGNERxRRaLEM9rPbOd
hNrDJApQBHQGr4IyXFlWStzp4rU3xgE/AXsV+G0VOasy/mqZonzK+5bXSDyaS9MySkY0qzCpFQep
uHIq8RSkzrlxgstSMspdw7yrr6JLxmyLfllAoWW4eds8HLSdIm4s19nANRlKSfr9KQ/4mr7VoMR8
hKU52nhEMtzXkso5SjwaJpqR3surZGJJ6crYVf9/H0tYmczXdmpqOO1uv18GsQVNOD55y6Eoj3U9
sJ8z94yQBm7LvyBSqdHvm43nkkG6EDep0bY9dCZBwFMVYnCSoI9UX1nxr5E7lSz29YOCYqqdvl2Z
82Rb6VWq6uvG3Zu+v0e32I6gC4iDu+8f17R6m95TMaor+7XezFo/rgx80hRM45ejm7ZcdqgAoFGA
SQ9MA8BrLfV5HsV0a/gQ+S7xyWCC7taM9Kf1sYuqBtJ/jmrQISBj7SPQtMEyppKCe3IzqMp83pxf
h093aLigOrnmY9cGPurKUABjqkf6nUsphPlW9HWuchUFcZI92yzlALJY9isPvfgYg4b7m3Zcdpyy
k0uI0BnnPzGXFE8p2aGQGc6pxaDWI2F9UjVTgQwSa8j01Hoe0At2tVf7oiMfY36aVPzviZnoj4zL
mCt3/73c9Awbyhc1QKMSMwhqMlQLStSXp5pyNfF0c7upXuVoDNEXxUQ4sHYv4IIPLgvrz+L5zuhy
XXw9txhVx3d/dj5Ibbm85AWfl//wo81cLJB9XtxmOl8Bca/ir13Wm0ca1JiGo7w5Epi9hikQ5uwp
8DVaoaX+AuBTCYsY10Fwsl32uLvIg0XC2r1uFnG8pHdSiUDTME3nNBDxZEH5hciInoLdjKmCH8g4
tHDr/ovXkVldh7qUFvPozIihrLc6WnzRLOBowXKfIiXFfbT1dtGk494OpHAIEXj1F71SfRyZP164
LpfuUmJGackvcn0UehAGAUYPDDram8ZrTHem+zf5gCxIhE+BUXKBmfNyxTphadChLF04YNcuViCO
PacD/iJITL+taRjB5o0FQHcPIN7hsrxo3xFfzMRqVzEwGYQzFRnm8lDuRI3NwpJRn92PBIFUFkFK
fiSt10rRHH+iysxQEv2547dQVxAdUzBMuFk9p56AQdDbIpi1DRfUc1oKV0bPjsiVBtTnUurnzfZ/
j/dh4zWGIXocvcPeQe3EHmIYirOPi0RikJUuRPmjGxmhVnH7eLUaOamLycZ9KdM7giQ2BvcmzFXO
WL9dyGIH2HmGh/V73K4o7v8IryUu7XanwwgjMoODrkE1fT2IkzWOlubQfEuIoow1MWxXfpMofhj3
HtUSIz4U0ZVYMCIvV6fdVPU4KGg7QVxRQ0vhl4A9hVcJOxQ8vAdlmw+QK/SUDTcXfPwbTIYXOrJI
1x2eES0Kmnuma0qLNX5sxFQMNGLVyFf/KX9cayJQviTyBHU6C62Lhx7Z1c9hzvyEwiNJnQoJH8Sd
eRn41YemVmzz760JMNRFBqlHxEvKrT0pHT9rKtko5ckTVGbHcEazEV2ty7IopfHUKXGb0UXpuFPc
EhbdXZkHV36bt0Ta9FlQp50zWM8xr6PKMdoiQyBtG2WZBWRl6+BzrrlIV41maH3fNgYdGCGRR/Jb
KVCgiXeOdatXccyQPNGwMkUQfsH6DF1DVbqCp8ANkVa41T5sq683qhasAGIp2M+4lEOPlIy43buK
aGA8JfIr/WNHDDKqlEvNxNjVF67JvRdXjos16EnrtyTGf5KgOv1xiij27BRweSODWKAfg2xmnjHq
w6F3ZyKCv5IIYAA5Wl1GRFX6c8YUWsGEFb6ax0Ae7AsyTzxqbv9JIn1hK46y988zBRCjRMC5HtrN
0/vETqxlSrBWZNCF1jIbj3d82FyfY1v1mW8jo0DiFlfnlqqAMN2ZIapsg3ok4tWG0XVc54OSK2w8
TcRiOwjfEEwUgrN7puzTHkxKYIp91EYfeKLXUOZjtRNB3wscgBRGg5T4Z4RzxuWzZZVzRXMWOnAe
B0rNG0nso0IwvuMknhzByBZB5Jkq/Ph/JVhTpTiQZUS94hdYz0mEtWA25BF6Zpq/RuWFggOibfSG
5X14AKT04oE/F0vH+h9AFdK/PQBE9u2bGV2v4IfN/m41juLizBixmQjB8uAgOHTntahO97J95rcW
xsp2pIBVKjcYw1S2mr9YxC/2XFhL93O8ptzj0WABvVN0CmYSQaq8S1t7vkjbseCWfHzUASP3Mfue
sOa0N713YKdtBho2w3lKRfP4KSIA+KDTylnZXM+n2nez8RavA0fP6CuhSRZ7OrtzxhlRylg/KyEU
XpAJ9hkKkaSYkGu2M7qQt9nStHFw4QpUk1BgaRKzSeCUpOJoUot59kDSJS+JNt0/kGS3+AY0QJe7
RlZk3Hps4JtaRhLdFogoQaPO0c5ZEYoBVuoEPde/PH8UNe2usEGz43R5pBtGbDO3Dpxn0XCN6iY4
erc/g0mJuIucCRrdw7UB3chaHk6viVoFOaDIHk9h/HvAvQ1Sq4S9KMZJkCXH60PwDbgx/l7kiisx
xWAVZDDClGPguZrwKuqdvIn96B4S2wvzKENG9xLp9b3qfHiZezNwaJO1kYuPRLaVIwkSKL8B3mEo
6EkEl8a6GrQDCiB3DROAxu9kcYkKZSq6WERAaTwXbwU0HLUMngjSJIvEmucZz5qJw4rL3n1IQz4M
22XILqYeF4Uf6zelV94CVCDdILmPlwUxG2GIuFVvV1taTTdsCbEEj2LTOQO+hxYlTqz6pjTBiUfA
uD/WLiMS06k7O0/p50JyV+dphZum4t3TQZbZsbwerXLCtP/0YrPTkVCv0L9cIkDwivB2HJpJZyGh
N9UVYfjFW82luIjUVTV8qt0wZTzCjNY6b/NRM/GB5OqJewUlqbAibupbuzzWbdYslc8RfKCESW1/
p1BP7jL1DG5p0/N/3pRo6jViYj7juazrTeByYqUYlaUXJsw6voQu6lNyDdbPETtf8DGwZ647J+y6
1989k6bUEWLdKXAMheCodX0atFHLJLZe3PQCziCHMTLftzIi6lQyXuKC50rdzevw6Vu8i2zSECpo
DsoRFE3EL+Dx2WixtNLXQHsNf5ry+oBQZQOoSttH/JaRa/zbGEVqWh5JnMMT0XyiFUS8OfnixBa3
LYmvgO9lCMxMpDS67P5nrZPGLuJKJwLFTdZ0inxbiy7U844rMFdCw6cRbU4eOlkv6lRjPrAl6/fH
o+b4dCxP+RqSSF6uW/Js9yL3Egezd64fEftmS0x4UhjYR1xcE0X+smb9QOUsaIQbgMrNHldi26gV
T9TTKLqYhU5fX63qMsC9FJrPsmCf4poHUVWQwgKK5869jkSUchd2/QwtFM+o6ju0nxFfZ0hoF3/q
bqLzkb8U6x/4Wkh1BYFYfSHvyWzJcYpiWboP5HMhc9bqltxzsD9MhELUI1vU0AWPl2gdbdheqaJN
vJG9CgMVYCrnQosvYkDuWcfFtuIJr4qc1PEFgCUraVfqe99n6aOc6lT/yY0vPFBE6j6sKQhQSJpE
oCrt61Tl/f0foUKHqn+tbbExtgt8ge35MQ1WMjQR5WiPvSQNgf6bAE5CjeesvmOsoYFc0W09aWTg
65v3YtInHy1w4+8IdsOAqqysq3FPnDq6EVUOdSa7yYUfvd5RtDi6G7n50hWWE/D8obRWdkxsMm5F
0f+vLEFom5cZoqv6ZxNoHSN1GC3/XacxwymgqZN2sJntHfVx2UYjbV7JsMbNgwQoSacs60jSMzf2
w+s3grMbh9NgPF4uOu13FtP+nS75bfkjO1zMns1n8urOozlvn0HAmSH8TuFf1CyzY7ibszTnqWdh
EWQAFKvLz2KSlWY8Kh634axBPbm4+x6V6LMx90OzJDCiV4soCmEst84cu43MTzklFrO/3qafD45+
BB/1/LUKK/URSJpUa231yhqFZW7ksGhHcV/E8SQOWr40mAiuPD9WRF4IK9mfD2ay4I5ZhcApxdPC
sXWZ4G9aR5Oah9KksIoBjVgsin59IuYjWBhqBvWFqJGugFmWW5g9mmY3vphBpjFnfKlMLZIOcVyA
hQZtukzL90OByA9Od3ICoUhY7jA2kpjr83Hkv5BYqhxX2zd2En9wr2BrYI7LF5XnrhjLqENtNDEY
O9mccwMrKWcORe6AHmHOcXdXz1h0HFKztAogD/WpgpOzuq98hvPZc4hGKZea9SeTmN0g0BBnGU+G
WHHeEL7ibt7EvvYaUSsCEca3WFl8yOfkSiaQQvC8D6N4njgzLNHamJUeDFehK9TlC7JJx0//HbL1
aQiuKfxUCe7mMufx5oSWN9AGrY0GKg5+wHdQLNDddv0NfLTHQ/p8455SYGvkAYh1LLC3inGLfsr7
MB9ZYvES8IgXJf7BDiH4spX8A+FdOFX77pChnnb9iXmw8NrDNjS8zzD28KNQJhz7etondAWh1rPw
ufuUV4HZo6PDLj3LUdIEU2NCmw7EpZNgYPj4i4Rgt71/UiFg2Ktbg8vh7anIEqAmu5gqnO86Uplo
JSZRouvYjrxud+ad8lNzp1rXpT0FSCwKJ7Cs9J8eM0mfqIemCFrif80yps0fahwmdsstF85sOdZh
pjNbZzyzfm/eapzvgMQfbzYubFNkw9n8lm+XnWSlALqWWpygRTS/cgV5rXiidsMDUc+FZL17UdSq
Ss9+aUG+JDOQSwDThOJY8hDlq/IHriaPiGHu3+uqTqcfJ2N2b1/kbaIK9Mbaji3VMVi55UwEXT2n
/H7z98/x9rziYkTm41ar2dSdgRAbk4opEawChYBeH9VABhxOC+mLbTpLTpnYPZ7h+uTRPvJRhX4S
xpV6sxSw7nBTVaP0fb6wxGE2kLKsAwFIfRxdv6Ql/b5pwnAKULZbmcKgYU8fO55nOPuemsIX3RXy
KzIg+1WBA1Jwqw1K1KuIN+N/MB/uD2RpGNWwVYl38KNAh/jaGTElMU8sZxNuLMfJw6QaxCcZ+xje
ENDdrslEXeJznEMotvDAJ5vYgtllauAf1VjAAoPH4vRZAT57bJBWlQCYOd0qLFnCM6U6Q78E6AOg
GqcO44qD03eRzmFGu0f4Gxmdb0PpEr18opbUb8LUAs7Y9k9azJJ5HpDikHkV2KX55CLx7c0u3Viz
U3KhQcOSDL7M6D0tySNrpPXy3nSQ/t8emjOnnaqRim2h8LsLq9mGOj+NzhYdTVx5r8vx9+hpA0rX
2XuM0qpYxTM38OT2HgXaIw/E4tZ7i5Fg63gZ0FlwEpYv9NwwsbOA+jMPmMv6yirKGPSlogZPGual
ZW6vgzGf28J03E4w/NiNRjGVeMla4jkr0bjyzv5w29GgUxmQbUVRZz+G5NA2zTwfIDHBFspApag5
gXyBWHogSWMP8+ojI5P1T59i+0mF8/J6autwgk2Oqkf1B7LD254zg0ZO8pySbAuscZGfh2MoN3Oh
iZshOM+A23bepbxCNPx4Q5+aq7TrvRGcK5dPSOQnI5ErMjX4P0p1YD7ya0S1YHGm8fVJRWYrxVGQ
TNRp8DP8YQJPTEWqoEbJIk/LZG7tXb2f89FcekKAVkxkgGpaYH/AMrUjLK8a5+sAPLeFi3DugoLx
xR0M/NF3zHWRGzn23eBw0CBuLmqD92pAl1HsPo9Ivs02WU6lgZxZ98M1WMKS3UR0ua771ztuTa5T
N8WlGq9m5foZBPl5C/B9RNtpopt436bbyPY6GUqKB74B5H9mB1r/L3SUNIRLqEL0t+NjjWt6aVFn
iA3Dvl9rNNysz+oRy6UXrRbk1fRvUF+iaqMNN0vB/Bhql1rYCKPibYyB4mTZZNrNPNukbryTG/G4
WfGn7DqUMcwkc7cMy2kvMzKXBhWWLrcYD96JjpHb0wBJAcF6880uTzj9UuLa8OAOFhYe9pkY7FeL
oH6kJ5FSoCFwEG2ZbChJTVNmOzdA51X7+go5L787eFfzZ64Vgpmm1LzNF/WjAWSFjUvW0t1n5FEC
dXZOKzsWIHY1l0M2PbrSOBgOOr+MNvlJ93GACaTU64VnREF66uNuAOB20Bqs6bjNcK1hGebOE4lt
ldUOSQiCtBaxTe+QbYoYwLvdIkzmpRwP3cep7LLrzdSlcibgXx42WQ43AquvZqDi3wPv66ZnQqR/
kc4JyxNIYxNEL8RcrwjuYHtJJ9uAZ2sKBkvjg+zqhloVeMPzrhXttBiwbIXgyA9hkMOS6NL54VGR
aEgnZ2dWzD/XjBrGybeCfl5L9Zi8rtJWIMJyXRqoaK2BF02X0bcO22Zx+kdGz2eDmw5U9TWr+DPC
6CWyssA3b8U0NOolRRhliJGScVSdU/tar3SO2SPYk2y9cLlc4xyTElCiZrXsAJBlfBFhUsbcf38g
OeT3iW0or6vdqbGc5aSwWqB+Epu8mloYRK8PfCHNM2xaed0JGPP2maJM+10qvV7lSvJ2YTxBHfVS
62GsGoAg6RVItMzP3SXx6i2mzNpJ6zz++ED6DR72Kv35XnFt2VMqnoh1V5eBlbY9+rBa/yLl+Smm
mgroF+eq4WrTzavRvjmjMgjHp896orZVf1zOTdaJ0ExkiwVFlVYivwsm5bfEOmGPINikUgGodn96
99yuKGvGnvuiMtgClzWdIy+wiu6tVWbE4FMEKsAD0MPSCz8zU855LrwZoSeMN9cGyMLchntPmd9t
uQrGXqee/1EpfIphknuzjGSOQ5vIWjgufAHziP3W7eK2LU9F3N33PGyk4B209KbmL8v4Ys3oInxB
uIoZ95j4AEfMmATvnc2aiPeXBUDEqMvgLOQmCRZdj0V6o4c5VqmACn2yKx6Sexo+/kFXWB3UvX3J
oJHoR/bJ7CAHSR+VEyVPDBRLbxv8V2FkoD1FhLUzdBZOaipTXlNuuQaRH0sWUMjtNB44RrBmgmN/
kY2Q8pETprAos4Y9klWmmnko4lxs+15nd4O2G4Hh8W+5DuSeB0f7AJR/rBwMfMoKpsanropxcDUE
N1Z4j7YxspcKMFRbzVgAppPkytrqh3HKLKin+p0mNP9LjItQ3D7QhFdQdTCMhINMNqyIadfr6TtW
nzDm+vBP+IDmmvBxoLAUd8zJ6tg5NHnuuUH2c0ceF3gM6tXIPEdKetcYeqYlw7JSDaQPWjYKUeB7
ROjqOLuI4/prtQy8/09eNnr/WTNPNzTQFcWumswbmgx6m/zLrIbXLzhHadi27Tj8JO7JrWf7zUDU
R4Hl9Tl02GlK3G+pJJFlRu2mtgscTXwwObITCnvBablwmsOoM7QZ74dEFMG6iHSeRZ3eUVsD6eYn
GKh17loCMF3KGyp5x3v1a5QF+G+e1EdC/wqH59IiSg7PgSqrCsDHApgj5aeef2f2AYX9FVFNf/qV
QeaHnsR8GpimNWJbblttbt7NlPbhgoRKLYXVNhbG1dnS/EOH+7rptYAStTpfe2dSW56PfkeHOnbv
PtIc+Y6QmoMJ+1cTC+NLXmPdxnNdCz56gxZhhlBIcSKfIwWGJm+2glYuN74FKhA9SaLaPM29lqib
Ws/WRIjOpqw3L35qGIu0ljZxYueZe5AqNb9FyGuL0+ib2U41YCBxZ1jjP/2pDzMk2oMUtmD7smnh
UuCXZgHF2C+k36CJLQGLRmaaYaSyrkVbQV8qAGOtbiywm1DyyR9rzCk96Dse3tcf0Bsv4ZyMdepI
+cdDjk5poURryblDnYMQKk1wEx1j3bPyChzxXa35gHMRMUDaQKdxjNmVWrYVDFcCEvV4ID3Tp/wf
Kr+D8OZiskPAf1U6ruXdkq/XgoHgfk26mg1D6CjTU4jESZEqYcbxneCIKgsr2dPGlqqib1bKF345
w+fC99ul34dSzqXetGpXAwx4b8sd9b+CrzYsKgQQ/DEYuI5Mtsc4ASxAnJelLv2zmunnMg8XDo71
bkQaJYhPkEV19nqrUSjOCoCnhdbLaJGRv5hlnrhgKu9lgXhqktURtCCKAW9vXyn8Rhe62ArzYdWE
CV3yvkUDoMVxg/WEiXzLmRfhAvEddePacXsTttY2+qAqFh/+U47yybqK4j6fM2SBTJdCpTI0LHIY
js6T2HYKSOMBnU+pDAiY2BH8EFBMlCi9ZMy4zDxuXaL98keKG+fTmiISYQ20U9z7jOZtBrcW3r9Z
3UHIpDanIWmsGcOFLW9tOOc94V2T8a4yEsI591HJpdMM++2N8ga3LjIEqBECyIgL3ChPdWjoXHse
sEeJT+qlgk+6X2eL0eU/i9/xtqYdt30npM8hCEJkv4AJGu+EWHQ9IMNKJHag22e2N3PQcMg2Phjg
/rnMgXpRTJOwpKfvnQxoLypbGpAQT2Ug1cNvrvhXa2EFJyjUXoGLVQGla5f8y+n7bqt3uIkpynFq
aHk1ljLmhzEFCdomIsVver865M2p9VcuCDtdiz6Yxz5uKYOZrDwGsa+uXuRuUnN7n42vqTEe+JKU
CTo057LVbV/sxGXiplou+blTG1lj4x47jSZxamxEYV2DQCj+k+XOKt8hWVB/ljpd4jPVKhiKbB3o
VzqZ+sE8l4uJ8QpBttpc12BLtO/4Ahja+xP7h+FsUB4Smmh7GULejMdcJYcU/NbVD29n6K5sj0kF
+eZJsmBtxQfUd6KiDxqZVe1OhHKRKYii598YKi6A46D4sPY9ANHmXyVZbrOE2oUl6pN+QkYnDJuN
xL+EPfkCO2nW5lJ6s/ai8nglHtchTNRx82epnFG6yogF+77hkxjKmxKqb6ycixYJykV/DZdcaqI5
RO3i1lTTgvwiB44MQnwVvUMdTBWCNKsOcQe3CWGw5mFP9k2jz9uauWE4FgDpzpHNtv7SMKKFj4RF
qiu1g/j00mkzhi0gvIY7mNW4U9p/7zpJy6nXSDnUQp5WM13TjRzfr9Qpd9O6PMcw4GYIm14ICTWs
FsGmcYQM5AX7LfWWbr3wxk6AHUKmgaW7BOuhGxGkRglcJkW93fjwm3uGK7HcUkujFLn1xEYsdiRT
jzO9G0ZsVOqrXfLch5tNumKkM1dmTTnXOSvkCAnqvUd3yEG750c+4fLs9lIn36HzIrCuYks8agAU
8j78IAYBrnlFZ6QG13wcrBl5J7HHV9T8KsHmLF3R2vvTx3YmMhx7fwuvk1erbGo+S7UoYYMKs5h3
M1kOfsWl1DoqFmkp8RpCsTeI/Bnph5YbFnOtatHZch+jikQHQBxULb3095T+WmAnsJNMvlsIePIp
PqYA2W5K4c4KX0zwG+gZT+pIlkA5xLUye2bZ330EozmYO9M/HEQarmnqWACZ6rSJlhkJ8zZOae58
ebCUDEakP0YvSKWjLASdEps0WPmF2gjtDmNPpNqwCaQXc9GNH8kUAgWwvb/m9qFKa/DOVI3CAN58
9ZMlklVGWuRH24m2sNZci7WKedJErzddBnfhVgyzBgDJJUjUJsZ73jf9KF0AZNIn8tO5DlgtRQYr
idOGoedRvj+duA+JqeCS+o9GwEmP6ts5Gs7r4UKsoOQjhT6/NF3tBtAIiSM3dGYpOWo83r9ibBTq
gcf4srPHZrZyNLajvwRS1w/L1PvXmFc0prHW8vkbbL0cItRX/cKe6akd1PHFIL3zqUGEvbxvNbuc
y5JtFXFJ/YIJ4REYKCStARRLzdANgz5aI7K3fBOqlfPV8u8WfI54ZEQHcsESsEGLns6dvO86ki6F
L70vOiT5MtYvgRfPxXcM9TUr39u8MXHjglzSKGK6PaX4LpPYc+suKFNmXHRf2imqupRs6Rh1AUNS
CWipfaCvyOwI2jHwXPfU5Z5wgMUUFHYaEs7lFnM46Ab8YuQzdT12JOArqb3nbq+D9Q0HgxO7FwFv
i885jr8lUQG4XqjdFfZbwIoI2/PNJut9I4K0w77K9h62L+wYVOew/AmHamhxe2dAKuSKEDR909Tl
ejYtd8/PwVdgRvLn4d6DrmFAOdpUWZ95jGA3aWq7pSUn3gNi/2gRLWOYnWplULCjh9xwK9vV1DX6
56hJCbt4Oa4CCn2Yy4XVdbyzyvPUINvfjiG5LTGI+gPulJV74W8nr8DlRrM7GiSuHWGpIOdoD/XS
hTwZzpLk4RVPea+J9BStwNoUNnkzCx0A7UMuegHIKPW28tXSCBmOXtJmiYSIBtgjuVy9YU8bCyRT
CLXYT9DSHT+1ZIihK6kWSryJfdCncmFdR6hoChlXrpad7JBQcZb5Esq4tjSeQhEGioqhbyGCsi9B
YZJsjNaSa4vVHRSPTW+GgdA3r9/2Mcz1T++CeLO9BHIOoyiWFkLGGZF7CKc1vj4Egix0QJAGathf
jinP59sxG6X668Oxzk9QHuTgwBEPMLnrfGO51Nbdmb7m4KryitGbDqJNPbsnUZvu4L3dClAez85x
GwU9VRRTBeOgoEHxLpAymmx/MWQ8VG2Tv6ZnYZqgV/aK/KrFaMypCAl9RvdACir/U8cIv6LyTeur
zDWk0ugE48vpDBqNWcAmsxzpbOR4xA5v6ZhKHG3gwoe8iPuu71o4APLpoDA5PfwJeoCXs0MuF92q
p9FaskW6fncb1YZBtL+fQW+if1v0uYNcNYHQ+7f25exjuvaLMMDh/lprhFXju26uP923fQRjkFYc
to98uoCCmhJyJhQo2Px1v5mDSvWo3xZKmisVAnwOS/vP37texwtbzajpGIMq4+vZ2DgAej3/QxS3
ejHMFVWoP8zsvBjiRGdmwVFmU8fS48ygjMBb7VulJ9aYs57aTryCAquc5ZoeE1pXryrQbre11YVK
t+sAb6YNUk968M2giLSMRTJ3qkwmYx86qQWzTKgPZS5E7A5fKf/+3UI53HaBsPRKtWZOOBAavOqr
zAcQbejHrjS+TlpfI6sYUE5ogxalNjEX1rtpa2HYCX77H48A9bBJ5dwMSoy/Jh04cg7nB+rbd10e
p3WeA0nmdOOYwYjoAxVp+H4mXTO6UnHt1D/k72YLvO2C785HDTd/OoGR5fitAKYgSbaUAgAzEa1L
1kNbxRLWmsoV5SiP5YqtEEyxbYCLTgRzX6HS9uMQAOYncH3nT8zFf+A0ZoP/AOoxccALJUE/JOI2
hyHfZ42cQKGMt6k1ENJ3oN18RNGZNGx/W8r98TAdF/EnbWgmQ7pDQvzuSqDNoYkdm5aqdFwSZH9p
GiyEFBcrM9wSuUjlXCPJDPZjdEBWZksmqG6154bVjFS8j+fMSV6AVPHbwuBN3+9c9fzhMm2J9/Ni
xZYnqT+ysXRsp7040yl3f2Cmf9AJWyN1h7VMozY2kaVUotyakBrfQiDnBkJq9IUeT2ihEj8I9Qqf
RTxh/jJyDlNLmB5RlXo9DtC+p2eJdr1vQnhDAXdHuA1qOhOZgE0ZL9Kok51MeZesUxx68U1wness
ZohtPTzlvgR0roVq4pS9YtWMnMl0ftZvqsO5uYwkoHrwjp2m1vW17W3R/aKnLS5BwJv1u+2RVuNV
PFWre7ZvrY0hBUsbDGtJqx+6hdoZJCo1eUB971QsbEbDlNolopRf73ng5xBKSe2s7cpiBOH7qJW5
Jk2DroCx4/sFd+AS3Zk4QjJIJZQSOIAAzxWH5uT0UQiKzBTXl3nDElkYY47JVyCdtRLzI5i1uOTI
gpBq+pyDIKF9PkMh9mB+6r0DKgFvaMhrLlUtbO9pu44glQFi3y/w7hWOHsbHB+cVUHsm20kmmqQN
8uxtQ7f+A25WV2qTXPKrhXn08jbXByAkX7DdK28FcPIlr9HhhUa6ASbxwImwrxMVl1XjOiicb/Lu
RA755PHjJgxVFVUreynNMtIoBmLJUp7mvjiwjp1UXRaVEGMVTo/p0kso12qS5lofkmCnj+aRfGwK
5+4ntEkuAUE/AXLlnLbdUh0ImT7tfC0KzDwh8Zeb/E4j84bAZKmtl/1oyd+qR8LrVwTllIyCimXK
G5Hla+/Lpa5Ubn1WsrloRd1qXO4bCx6EmVypzf5qNjTsclU8Ch2uZxCikoYA58LiOUBaZvoQ36DO
vFB9y+BP/Mu3GpNA3IHkmDx7Kb6QpN9ii3T0i6LvSI14rDHI8ZnIwJ9jPc7siwOWbSknbWeU2cVs
ZMkBAyjT7S2+Hej1wMDcxLG7qbvoMBO39oY1ugIaVvGdWCqKVJx5aIVQAix+P3jJ1WOm5Twxupfz
jeJsryhagNbxcFqEZYGwExDfhCVQ+kZAQRjpxpqH/QxACceIl2pSOVtYbSnQtluspPmPwjwWgPYA
VkrAxb5P6lBqzjJLtoFTkPMdtuMaJQeO6Q3DWDMyzU9KasBY8/lxyTbtiKxw5Xiijfu07KPYoN1/
OYAT4HO0D2tasIzsfNYwRnBSgDwwm+djXOBK471n3Taq4BLenDeG/+u/ESlBJPxvwHT7XpaTRNba
dQCp4RTxRG3vzE+I9OsOo65UJaT0WscrfrOWRdRJuSFpgnOhhtdwGAIwb9M8pGCmu4HVj6ZSNGhn
UOWJVWweDWieMgMhImnE+TyB/rjCLi+FSMCkFqU8ViNqJXrIgXi7G0Y5sF+FNwkRqVpmCIMDxk0Y
hmK8jjGebByq+Sc5i64+1p8gwO4knEvGbfEc0lQnQtF8RPFa+W6JHpgKlGzzv6+rG2d3rSrRaQRT
kqY87WTcj50b6fBUI5kux2DzX5PKxkYJ2OozH3WN4flhfKXJ3HzhZsTBW8fezMfLbNNSaETFhLPS
iYhDU4V6hyVcoLiHZZhMdLbI4kd+oi+5wSVNmL1+U+XfgsTfLGisA6YSjpLbM45zUq8C3GCWEMKe
XkO6dEmfag5zGbqxsOwcDgiI1IB2a6YuIs+tsVwz/ri6ciHRpWP71zMTB6JVWBPeybcXsxwu7Vla
ESfekvBO7nub8/HEujuZHfo4zwcu2hogEgQ1bdOfob+9bxsps5Hf/XVOJJmcP4Tv3sKbMZeigrfJ
ATUErqD1DEMsTZiIDLEuZnopK1soDRn4Y2Cb7zTKvrmR12tRZez60xbTwkyATDH3B39zfZ+piTl8
oTAE7xrsutcfftDaSi/I9UVomEebwHO2tZUHbwmEjhEbWv3KLvIOmCgWE7eJa8TV3GxmNQfQxmup
PVo/VptKD4/gonnzP5q1YUfoqhrXWRpNm+F9xbJFv7NHn4iyxDZQcC2yPQmNQCvNklrioHd4+3fr
xFXwBTV/BUgE0AsgjsywLL+fLRLtO3dRfkNrVosIqh3VEPyvg85oewEwJyrgm0cUoAdrP1MSfHGm
2bYuc7uTELSHKRoLLTO4nwMDAHfHt+k8uVVtPxLBhsQr7pNjS83BVz1duIJckSuhqtwz3hB0Vcm/
M7cGbO8xN6LPjXodZMqsw4eLiIz0VKz1I6J24n80GPbmuGymPlvKaCkgbhbp5vB5O3SZX2Id3NXh
gwt94UnX39EY6yYyc0RIj1aQBjhTJMw2YM3/0g9W2fBEffdD4atSX6EmYQXpK758AKQ+Cky3KCqx
aKfBHOqJBChCXDEjf6YfNq2Bk/y4nRm7WQ2xozTd/tEp5/vihVZWf7D6EmrQBIoh5Cd+lkxqP6HU
w91MQV2wkQfITdp6dOZ0X5Z5WpJ+qmnRYFCt+/szbwG/ZsILng8cyWzoRexFj2wIcHkBozW11Sht
aJgjAWJqhnbM0Ot99f7PGZIhdVVRZJ4dbqj6im5Rgo5sb78F/ddB4Clqsh+/G9suO7lGYaaF+lHW
h7IhDVddoVx7SbRcGXAXiDmhJT3tYZTl1qQMUvrLgvmeeZGcRt5/uA5eBZmWZ9sV2fSsH8cno2ny
7Zkj0jWMz8Sp4Z0vULyyyFeJEbCorrR8eYQdzwSkDND74L0tNr1OlgCkwEFWGHRz/FefimAbF/Kc
9yeLNvhg7xRyK2UtVtbEqhGDyl9yrq3wtYVVBrqVkaFEAZbSMkgrKLQjOExG4tL0ncW04skhRCwa
PHEuXeyPqzFLJLWkXTMJtOZbqd0Og/4q1avW0IDTTAhKVFJAjPmH58nBMn8HNJO7xCOLHG0UeEUz
R6ud4c8+VNOYVmtC7vWGiNczv7NHU16Ka5I8yImevyURJhmsj/8VVasqgeOxcBNhZDgwdoQTJWvM
j8fx4A+9gNrorjPg77ab7EYexS3HbacPHj2eSr95XBV/Qd9hGpPqJXBr0Ffv/RKYl6hGIxWO7aKf
dMZsBHonBOeUbfahrqj+FA4FCBhkCb6a7VIOQciMz0O+jSvNcLPMJWNBgppe1NIVR5NU7i95QtBz
o40Un55XDkbOjQ4h52h69Bgq2sEUrSKHR4ZxzGPqu9p/TcPooMGxFzfk5+FMDuY+AmQkHnjf+797
lsCrDq0bhaDlN2dcC06QZD0rHpDtXThugEvMhGJ8+/F9quoBjyUkjD/UYASNKL0PfnfsEY+BhE8X
AiTD//Eo6WRvX48BmMfO+vCp9RWZCAoYuh4SSavFEhROuTlp73/vWQUiUuM31hy8KYJsFY22Kqfj
ql1+ZX6fIEtc2cvG4Ek+5ifOGmDY+4AzOCWhvTlMVlWgAPnMhsqP06sK3DUgXtUeLUSC17kH2qUn
1VxbwzKUfWBFb/4dprxh/flLQQBo4aTthzFX9LkXJj3fK020U9Lsesx5vTWqmv6eAqJ4B8BeKtof
eXQYym2gyceHQlnAHGbV43LtSC895efWiga+RTesQbdH5GBOrlz8ZquS+vxGYkYjbioljJ99Nv7W
g/Shcgb1rnVX4dpgrsuxzJd/pWNVOHkt5NXXqioH4iChc7I2RrUQ5yqLF9YNQSCsqOR1Ix3NtV9Z
IJVC+KUPtLu60cebsLqCIGJEgJuuhGQAn6k6aIX7STY+rb4BJlt/Gh+uYsv/juYWj1x4/9bkUkTs
pBAkCsDKB5qBbVXSAgCno/agFx17DeZ/KGuPgaZ7sJfx8mteYEBYwqYlY6c8ASI/j84bSlrfApqm
mRSEaagQRpvMAaRdKTd5MucIAofkkjCVOsPJPj7ymnjZB2ENG1tXobboJegpTAX9X04F0prLcKe/
raVreFw2KNpphT2sjZpQmUo4QYxCAhozmMdpWo9lFPB0UVEp1hmds0kl4b66Y71FECBc8SFn91f2
FXE2KGaqq0wiww4JlvszD+XCm7Fsbo/pqyyRP9U3d6rHnUN/9OVwD8NTPisz95Pz3Kyo3j74v9eo
rWuNHiyr+hD0ghuUyMNK6ws3XSD8882m+PlbgnZn4CdLjRyw+6GltTfoRUiioeqXmiMCxx9VpwSh
Oc3rC5y+Qukdr/gpUaA8Nj5ZrW1eVc5FwMJHlA3sKvSkuG8YIL2AABQCZm3tpQsSbNO/egZmDRq0
MtIYArAwl6vEn8dCZoO7Z2zfhkMwB4fIKP5GfiK/toLNV4iOqFuBmKQFvA5croLGRmueqkKtJc6z
b/M0mK7LTrgtfAwtF63xdSolyAvKsxlZvxgD04hOKoeMDjRNrcME10qLerZNcYNObhFx5kUshNpm
foyc2im1Uy59ITcoz/Dycm4gBrrRSYhXOU3bH0kg1v13d04yuFco4CtbcVrPBfWXLBuT7TK/DuO1
EMPCG60H2/kkI4phxpSB0m8W5IWOWoTOoCWJZfPon0/pHiRHcc96A+QCy3gwmM2bsz3bdHoxTwaU
uHboL6KUjmq6Kv1VJitKyY5fr1aa19l4jgPgj+hftRzOC4uhUvrpyZVykaDpR+IVcaArbSjv6djV
gVWarLMaL+76Xay+MLnRxc3q14dKAwJz0HpE9n+ZBonK783b+2mjAN2OmRQeoH8jwesJgfR4TiCS
Wf4ynn9UU7t06/mMeyVCdUjjivzVY4aHXIT6SK+0bwv7iPsB/PG7tZ+j981dYQBaeDBuW6u5DwEd
Ac8f2YKe+6o17GtynUlPK+yrc8OmwmrNIn6xn9MU4DYzy4aHmJEBxyACXBj8yG+ZxOB2xqS53PlO
ZSxE9Gaa9bPOOBQ5nXtdtXx6qND8jyRhkHLzrt7jKakIH+/HDLjzCM1qRrJMbe3nVBcvbJDUr31A
nUgoBYhhYTshBNQ8rh2e9ks8fA7rBkNHbF0Qmnnyeq7Jq8kQm+2rcOAv/Rrg/jWidQwryC0Kd6B/
cH3GCNnbQNn4lNwrU2Dw4bQwq9qOI5aKlh/8l32C6ty2mD7MBNuudZ2BAMCROXpq07Zsm4ImaFBo
an+p82nwFQ3IouGb9j2DimchUM1DBcUTCuKHKafjd1if2IB8y4eSQ0ibJG52qCicf0fn3krlJkiu
FS9OnDRwqYEyhKrergyEzZAlCEaNzzxibkSxiiWcQT5hO+8qPZ8333jfV7tOWe8RnUQuLYmfTVuw
WW/YZpRErUWSF61gpY8wL+S5Ggvic0C7hFUwCd9uvmkv/Vgg1WzRWtV+SfawZunQX4qFd3he+iGx
yCkWaWwpmmmp45XN+shyXxlFQI7bQSu0OplmojpQjja4OFpmJiNA0318ItoKfmTcYKai7wn/Ff3b
FC+i9fPB23kX5ZPmeRl+CtmmunRIp45daXVxPiMiJij4g6JzgFE7YTjat1wmFKHHD817WkMXH13z
UcfuEr4sT0I22YA2aoOOCr9NDnKyXick+tmrKM02wC4FdIxSFcJB7d01MmBVatk7kKzupOB63Fb/
NHbIJGnDdYKGryNcsccmXauzP77u8CDlYqbscw7vBF1Ecy4R/Z5FbhEzx4ZrCokfi/Db9uI/cmF6
mWNdMm9ysK+cJBZU8MrIqEoGxIaI4a2KyIoh+dH8/uvCIjHcEK+AG4djimNmy8OjFCX/RK4pbNn0
0qs00GavhR319YZ5eLtAEYhNqO2Sp4/1hikBP/0g6tawzpoqKMKkbg18NhM2Z5ZUxhLFkck/ed39
xlwJTBBQiyneI0s5lKh1s7Ms8JtwMVpqZ/FPc1zREeYMjF7pIWMit1dvd60sqfL6pabtb6HNW3vE
m0MDsscqsit/nxeb7o91WxQWGzag8C+7cXw6MqRybkma8rRUgbG1Xmusc+VpNHQcSg1EOtvv2LCv
9ldUmsgn+4MP2znzqmqnyXufuPmDTWpbtCKjbQo74RlXwOec8dzGDs3ZBgkW60pa1e2NlOmOyRaD
acZ63IWcQC7v/SiOtkESnThKGL0Rs03W2ve3KpTmMvJdsBaiWuR0iVQw41dpcyjH1kMdImerP/4X
MgjVB1ZM7XtAYxHOyuN7IniidBW/IjnItpg2Mrrqu7xaNE5/KPDPzZVlVfd3bS+YQ6fPdNTvRaFa
bBSOdmzx5oZKnggsIRV/VVoXiCOJFM2ce/vgWcy8B5oU/nstaflmiX7Sfm7SFXYGct3G/sFvBGUd
8MGytErM2FH0kTEEoUGTGztkxgrAAm3GOqLpCtLlN/Ahp+ZjWd1vpK+h5kjClOqBuQfYcc0xGO9B
BkMOPJKQQcgGfgbEiaLLah57HOnNAPa7F9flHltPU3dk3vtLH5bsGxfZN6geIvPowkHpRa4Fmnks
xHfaNtavmrSJUOO3JqL2sN8Q7/7yYcTD75aoQYn1v7kBU/CAtdByziE3udiEpDkA8yMB1XXRwrCD
L6SQR7nVHzPT6Y0X/IIEU1cmWOeryo/jbSj/baF/gvONZak5qMatV4DgM/GjBJuU1ZZvjh6aivtv
nGl/GdXNiTmgDHLFwDHrh8GPymZa7Mu16VJFsS51+xw6PB8NL6STj1Sak8Me7OdrVKG5d9cvYukE
mEiMWRU4sksVEguz3fWqZgRjZizG2GTt9M0JqoeWGT7P9b1dQZ0ngsfweZuHwPdu7+X0/TurmQ0i
5g5KUgLKuqLtQkvv7rbnMyqEEKPA8KMhq4/ZvYUHFCpQmQY/00M+iEMkcgxU3B4SeP5BXOBKF46Q
8xQL9aCD0pv8dj+0+EgkHN2MBlmXggee8KROtmNCwdaNrDBMMqFNuWHxo8zL4bMluA//rGxmJg/l
fVaNq951Ya9fbA4j+tJo36WnGH/zTrijmQTd6HgMWRMdMhU5tWrIcdyfYZJGI2xnDn71jhvBd7sY
xmgdAPXAYijAU9Ke3NggXxbAzkzTGbvepqnAspMVB0Nh0iNuBcUnAcoScPa/giST3kro6/wuElVW
LKWX+5gdlTMW5ST9TTy8CivF45Uq/sN3vgc7Az4mE3eWz8o1KPCD4zdVISV9B0xq/rMtdxWJLlfA
fcIMClBPITcbdGmUQ2eap/Alo+UKbjgJO00YlpfMWU5tlLL8+qnYM8MdLLs/InFc0TesvPLQkLEB
yLN0c3K8+EMpQ8b2ihnvE89umCKLc/2Ux5bb7x0zvHKuWi60cDkaE8sa1h/eBaG2Wz6tcbQ6FVS0
xd6YcW8+Lx8xYkKRknXBVE0ngDekb5uhcviL955y+K3DDy5LRXWusZfDD9cvz3frMzgD343az1Fo
LU4J7CmCzoIzjoyuStfigEAE6uisLkK0oOgSqyrk6I19Bq7QnlYMqQx59lvulzcjjb2vqWpgAp0Z
zCEwQGrvtbhVjZ9Gg5AVvIuT74uwrX6bEPVt2YK5VqsoeNznuVjXX3LBlWnT8SgQiwGn75Zud0bP
cl1dPDmVJ6wX4pMHeS4Qrs9z5F6KEq86CiaobLCjPwFm665va+PSaTEfgmbPouXK5Nfe6YTLMVTJ
A1o69hCJ9E8AZWJpW2xLHYBi7bjLqVmn65r+Fi96hm/1hgGmYvTa1kvxYZw1Hc7CDnvawLMWKxA0
QdjZXqPY9LHw4qVQUVc2jqKz4U9gz8V3j2gIkEBmEza+U8jUJ9V2b0AUe4cFjx6JLOM9DvtGGOr1
JoDAaZdkHQEyLrkT0TVnPUNq/KSTcoz0XktGQzJoqNOt4yVzmT8OuPR/rAyD0Vo3qeEejsBJgvNL
Ohn1gpBS6f6dXgk+vhk9y3U8IzFJADlFEVC8lcFL87zijpkwJMZzHTONXS8g69GI+Pb/6fHivCMp
FoxT/7Gfq3te/oJwcdsL2dqD8rp/1aKiGZmRqfDdRG6NYOGe4FY6XNPI2CJQVJrhegIA3Fc1hrkP
488r5igxvoBDSMlsDiEVo8drvGtOdz3SZcJ3TcpTMtYXJRvQnpaDTe7zZvz8HKxuTlVbAb8+IO2W
K2nl2Tj4njDfhExXU3GURklqiOJNPBXuDhNk8QuSRBa+1clvMksjMMtDWwQ8hLSDeGjwUVDInj+U
CDMLMxVZwQ23YijTZaWuXjbAwgUtbyFcs4z70OoMt2rre5g20ybpSJbFVlh1dMSDpvK0IVOQKTeY
Jn2DktzMNwkfcj1ECX9TObznTPfM0Al3YkKWY3u5LfZDy+7Ycu3mMm9K3AZZ8+lXuEMsVZRUZt6T
86Qjlcd3VYyVlWLsYbtT7bgGbB/eLvQka+wkf97hj6SmbsThbYYEDe84/sc8tw29ZoW1nMj5gWGU
EG+DXRL0/f6sQILQ2Lz0qWCEPPlhxnKfoAtROQBxH0bIHtptXO3DQNIxfvLA3BdbPwifVr0DOXQM
c7FlG27RMgRuonOP+GZEmjxCPlrd1eh+ouWtvCblUr0I5ycq3krZSZQeWYeHzb1LoJmzBLZOMhH0
Xc011FPp+WNUytATtuxQEaxfJLuACrFwDICnt//rDd7FLKmZWX+Jt8I7pTlRK7FTa9WKN0MapBKi
wRYCBxFr6SuZuBRc1jEObKSjF2OrpMba4j6+c70Myapj2X7Ivya1cgZavvci1YvcXqw3bkw6TsbE
fBQTzGIazyRcsF0fsn4YAN6kf0CFHJJFa+FlnkazJ6lbc2i/KBkGn2SMxZc6HGFZQW6T2tjBfkbt
O2/Np2xClhljT1bE+naQSjvRXzRBy2mcNwUk08l7xnOn2QUcmM9R1tgjVV+NlILRoIMoD0yZxwcs
XU/CDg/9mjSYRUez8LsU+ajwjgsVsdl4S/6c0bEwKpQmIpG7P9vX+fu0/rozMh7KroCzEyN9jLwz
y/uN33HaphI6UaKAxyAQ+5265U5cnuFwRZw/9dqxN8Hae79Uo2XaI0VSNRZpbvDiKZc+xzQSPCWw
IB0ki3OondRV9aFsP5JDARN4EFn776Za+anMj3iBcoypVjaMZ61WPcA8LCb/GhlHYrJ6/aI5mwbB
vr+rviZPn2MYPaCc+LdvhCp+uwiKxab2Tqg3MeHI1NQkn0aU1Fp3LAXMAm2gvLMznk/pun11QC7V
CKnelQoG4+b0vv7VCofuvUJa84iUmytux5CSKQh/H9Pr9oBDyJJDMjC6zKZSB0YMZYIdr/bqQ7gq
sXkEx96nT2z9QiOONt4X55h7A/K53lhTc8Lr3S9ihvkYE3ERDDFLW6ZVUuxLSJXi9aNafQdkfz3b
fhORZX0Uya5e4IfsbNf1Gzor/evfrQIgDoAe/3SCZol3ppzNKjN8p+G9wVhas7q2Hu8L6eaEQxVP
+EewCyo6zkoCCLO0cBr4mI5e7zcsOS51WQ+f0wvtuRf0zENmOQYAIWQ5TjCypusd0qPtba0eGQX4
6NlLQS7M0tQCAMySfXnpmJ8pqYOZKAkYYnLCnCShLVa4YMZnikGTvY2bdlDcYO5TS3rr/C5c6eUg
6d/E6awLnFSGyGjC2pu63r0nzi4XDPYtaz6YbGA64vRluIJqTxXO1fgiqasKSIqPLPqOjG1oR3wP
3UQCUhX0pZXAULEX574JqQNeKKzD/CCrXgAcnplg0NIhEIc3BoA9okhCCM8FnVkc65M2JBOHZjo/
q/UyF28z9xd4c9hQ07VqGWAUYICISXAmwl4ldwp2iah93u9A0QVCb0aWY+cRGNMT4IWiIpvkaHMU
4c67YKSMICOchZD4hdEJ/DW0RuqYbbXZk8Q2MmiyKAPi+qh1rhQI958ES+3bk/fNwm6bzGVX6pVG
4MG6h+tDkwNXVA3jSkb4b7j3IblSm489Q8dRAFnyRfgwhjd/aQneidJPxQ8XEBTOwF3r7XyK6oh9
Kr5w9H1cdIFxcbWA/jOcfJd9ZFMuA5AO4FgzeuEtMoiBExTmJIc8iVuMu5Q/lHqKcdz3gfnjNlCa
+gwGJ1wvuAWnNx1ggzmpgbEgfdzQ+soMU9gf1j8dDBbFAOfXsmt06Khh59nyzT5kzqwKXMsCk404
cUGZESFkczBTpzrzI7erEYqY1boWbRXtbFsr3FbHA4Yn9rhLlLwRvbMo1NP3fWJkclTpVHOkg/B5
1sHHlWq0iF87mvbSD/TNL4ee5VzR0UxMR/h8LCCRQG3umhWiwKaHznNuveHL1H9RJYpW8aNRYO2l
b4zucigC8gs7oinrQcVsTSaAUdf0NuX2m2/6nIda6GFY8d6clN57cG6k+QqZ/uWgKL5mYq0nBmeO
pVuT7RfEO8TWq41uXZvZvXH08yIHKjpLke7H3RAk3o7EGCb+5iXhyEF89cvgwUUBdXH15rVbTRKA
cjiM3akQp6pxSsH5ULbMvvMdlQG/3joyBNvIQQbEk5MX7Dr2KpM5vHjWz9sK6MuHKzLLLEFrkYWu
bLt6/oiC5OYQVuuPcRgADcNN4wzvGvAvBd5Hwl8RYmOSG5ssjELjZyGB8DNP7ozvzYnUCBUekZRF
36iEcO38I2XmPJKTF9PTchiZDw3VabJbMWNVN01s3tBN9Q1LQt0a9KcGcUaaAl4OWSQkhblD/Yye
4HcjBdutBbRwBWw3wmUMXMYzfDS4T45oftuTvCtTKB65LhBsiNDfP9+0wb+8tBs/g9Y47hARlbJh
5a1Pf6ZfiIT2CF5EvCrxykxCIUqFAPxaYYMvDEufRHXnlaI0ipyWz2bp7rYSOvOdkV/Wz7w5SFQf
I3rtxmWsq+QglRuf8aBFRbMepJkdJ0+io6LBgaA95VrorT+cgRhsYCT/j2GGpXGcKkLncZTjxS+4
v0pzXZMTn+pZLfEU/g3+PTFXftxpjf343yRfTuXluMctaGejeCUuooYmzaH5DZql+gxKGsxhEMLY
HalbQLKfGmNoo18Jsr6zeWxtOciI5+BxrEp/01svmaAuNhEN9AwWeObOJxAj3uQFUyOOe4TgUGto
1iS3VoXMnnVTxIm5duJD2EqbSa9P780jyzsq9ZO3nSN5A7iZAM4argyo4Z7ozj6qYrnvM+zRET5y
LcZXVYXyGa4YcVZbpIPZJ+xHrrkeQAAQw3lOJ3eqgWPwHQYiTbSFWmL6yrAsVhWK0mi+lzi77/vF
Rd+Qu7zeXzHxpwgcWpUtc610oyhxFdoDdmn45ugutTs6akfZeegM0bhCeUJQOHALurVbsKFElJu+
/4DoB5huZI6UEH8or8WuRUvjhPWSompYIRp0znu7d1mHfTgTkkiAlBUMqB6EB8Cm0Cgnqa7cWaYk
miBXBM/WF5QVpm6xsOLEf1sOEuCNzetxD5H3YaoN5rPUYwvuzTi8l2aB4tKtwHdj3Nel6/LBU/3u
4+i3Rvc0lOtmmUMKG32ZUenhbv+zx1wSExdjrJ2lYSnG/tz6LJ6aiDtpQfk7LL6KzyNDpLup9y3E
eyNFL1WP679DUo/M6E9XyoBywfPuxJ6W6mOysd4PWLsRnkTgjx9p0rXGgAI0l+HhtuMirt4TJM6r
+iB57bgsX8rwGitY12/vW41S11oufKpvqgjgh17KwD/8Y0SRm7SM7mdHeSIoz+/cACIEflPwQPyI
RfxxzSEvbqd3QLnXSNMpwNyRTiqMqVk8RNnsJ4KtHeTrRvzPZHDZcGG953GAh2moHCRvxG7U4avr
krSnCAMDZyu5a2oEdtkBp88HPuTh/o5sejClGrxyZQuFk/lT4iZzHVb6gQenzYX/kyJZeR0fwJSs
zPLqdg3dI4CxEAyNODZv5E9l5nv9xErCVIg1ZmOhOV2KoC9kvDXjNMvAOXkkJA4WOFLMnNno+f6S
i2k2koqXWs4cZ+VFYuAqzkFEpXK7MeUepwBoFCW/JOB9o4/5TrJ8H774hV0SlC3P3DdweQIPD1nh
oZ5nnJYuVQkruP6GG5RJKytItrkHriP0AjekM1BDyOkWj5F9jCN65I4symL7uQY1u9mt3323nmkm
MNptlllJRf/7BRBF0U+a7OP0tPt2cVA000jZi0JLbN5LCIlk9NW7akFqiBRyA8k5zNu9VB7CHD8X
mkc3JmAdJIW6KJSuOefpsuvt8vRrVnZrz8CNEM5S13i0JzMQ29Vr3ueztMEnPwC6ODe2ewNpE2Mj
g9typuDyITe/iWC9vjsT9nmTnBoRgwZD8cvRtSzPB6sWznlyZFwJc1fTs8JBu/wKCXI87tSfw4WZ
ZUqD8OAabtk0upxRa3tmUp5HCg+kj2F7mrDB2i9CYqD/kxlDbvqtShqHiW66PhLd6n911X3jV7xW
WOsqhX6+BrcFAj0PhC8LD7Kj01U5Bmk6o5IJGtH2jvLDU+kX/mUdcWRC8q622pipWomBYh2N40yp
uqA4BW1+BLrOU1b1KtUNAU2KqvYCPdJyx+cHzP2Cy4Hkt6RRes94SZrtXRX2zojUPsoRoppH2EXq
OJc0u0czcij74Fqq79GCKExBYCNBNf58MdNzSnriggbyhnavyD8vxp4khSkEDXswqksegwoM8QfS
JHuEljRKhcAtW22ARqiNjuCRd8Q3NzbXAK94CWtJ9a51/MPPqLFjYDdOpdbVwEOluP42+B2EO/0Y
6AucnQqeDuqI0m2jrCdOjoqyfwRWeCc71mk+CnjuqFIN58XSWDDfuQNchrJyaFh1b/6hSSBx14e8
19/InehYIxw/GCABmR1TDmNCHwWhWjIcp2C2JUbBAOhT6q3zfjvkdnLfH0uBUuFRJpPMdJ3H6IMQ
W+jSHgM6F0BQmtNRQLrSvnKAP7M5C7xOt7UHZO95aJ2mG9UHOnFi0FOFlAq5z65D4Ku99gZdByp8
Gxaev4+3Bi2UvD3g7+R/BOQRYVc0GbgEX0f+TaTp08ozQEXrhfPXmBP4fyBhOp2Zp9KZw9cLovnV
sZYQOLW6yNl+tAx65PHkCCo1ST6yqW7grVEtJS3bpMAiB9dZpn9tBcz7cKcLUSNOqm1n1HfArjjH
8FU9g2x0Y4zrmCtlq61OqZotuWtl2TDAQVEKKi++yMut4n0ql37gkJ8Ud5vPhneBGt+QmYJrBj26
ErQTisIukNuNGbWHdwbCWdnBMYEeXIIbwm7gRmWIIv2NwXLoyKx8HSkPs003rrvgj57uK5GfasGH
9Z9uYTqiBJg3o74+sLN58ELripDOCFaIym8hyDjmCzXeY2Ur+ltKtAIDia4qVv5FMdJupyfpyzMO
0UEFgTUP2O1sIfiAjZAN/OKRMuYOdOietbTMbSRHMoIunxb3Rh/PgYt07bPq0VS8kxDg7+lqYrtx
f52BZ1uwXwsLNfie0kIrNoBk7YZ2a/T541syUcP+0FFzEJqvwhL7nS04nYdwYeUcd5Wj2ZXZQlZ8
YaAU3rD9fdFDPVDZqgaT86b92vPhwPYh1MBdePgTnPJKJDk8In5lTw61d1/1XL1ET6IiCA8osOtp
yRQRRya5HyGc6JlkuFu8CFL/5fk5y02xCsRKdbtLkumatmnyKx8XmB2QPpoWKMIGmMmwMux4XYfY
LvUaJwm2Hu8axNmYdVb3gqvqIC8AOzdoqSySvkkFoRwuWBWzGw/oxr8l+6piUcXSLiW1b5W2g1/W
T5S0n/yjG2lw5uRcFzMhXlxrFsBPiJr8QYnuIIBl2qGz3D6AyeIBOYcP5I24BV+/3UA7De9b4uwq
1h8OAQBulzsQvZxledJdHVxOpL4YHi3kb0ICKdW1Qza4RvDRoB/KRH5SKMgpvIXY/VWrL0zYpYAL
pXxf5pogWmRcaesLury9sVCRa9Tc89smoAzY17PgFo2YXk+PWSqoyxhherYuYhLjRweaLtkOfsgS
8eMoj+UxPNqiRHdemlCADGXEhv3+hoHY1V05guQTxySEnfqAp8v5vtMaKgsP1S4OhZGkGP9s8vw/
8LnKjoHMjbp/Snlc7We4JMph5rku+5XAv3It9yVTaeea55tZYWrf2Q9K74l/e36TLRMLxV22PO2A
Te/FWI892aNbrLlqzI4wDL9qYa9F+ttdoxv89xxuv9FR6ALoVm20ObagNZJKci68frmH6yaIj8TE
RoHKKycCT8IocaO1J5odVxNcC1pQrbBUufubXpzrd0VrelAJcATmvN0TxVzVl99tVzDWN+ywAb18
No5slSwufTmjW31KON8V1A8kYC/D3Cl5iPnQkGomv7NDeIX+9bRaUs30BvLX8KG+mF/dWISunkwB
UeA0CesFP+apj+r28/r3xSgXLJ57y1CLQqGoNO24+mJf0NjyuIZm1SogSELRnt9DuCPV/bMORwGB
rv9Y3A/L3PvRnXlgZLcYRcJxqq5dO5BEp1ukYNq6cw6F1tTfDqmKmLSCq+87E2yQL018lLQD7yU+
zDT1QiDy50ieoTZVFT4N9aecEOSvww7WQvsx26lQ+McmHeRDnTHWJXiBmptE/JzYACz2fyDGNtrz
dkcMWGoToy7gVQILFioHGmAc4P7WmmLD72s89/BTsf/3b+HMpykcd4fvv2e/heXXpltVYIlmum09
kw+rWoeo291pRIdBeXLFSWUb4SUGW0b2TdbWF0xfkjNClEnxqhj+thbXymxN2f6cxa6gqWB3hWhl
4xZzsntizg1YRLrl30sHTgvoVJTsCO2YwqHIUyrrvN2Kgt+wKnaw/smIeNoXKjsaZa7L53I6DENU
yxihReWjLqy7FrD/oCbu72kOki7by8kAut6VYBP4NqDCh8zFiU+nROQFBgC4ZlS6WFmHZsGxClCh
o7Cmk9y5i6UGpbDKM7LI4F1VYWYAbHaUhH+kmduvjc2PTI7CsYpZWEMZRLD4/aC6NKbZ+vZkuAUz
gjbmxnEipA2uSMXIyZaLyAILThqlLGYADn91vCnpkN4LUVFHgzghfg/OWVDSmrVBUAD/dqewvd/O
sx8QyPKMnUFwXyuIAq5xbLM/3gZ/H4+yuYFtHoj0lxcVjJoepsbPmcuQh65qgOeRy9ZnQrmDs4CE
iZlsN2gZEvNNvABp9d4EVP0YgDLeKgH+Bn/Ipb3Y7rtVLxOx9DrN0CA7lR1ZcO5sE062+uSSXdXk
FDJKdlAekXeRXnNJoWf0USvDpyIrr2GcrgY23FCqYRtT3Ft617qj0xxKjvCO34Eox6a46Wkn4Fne
1gDdZsUKn9UIYNGG7AXy9DyeyC2E3agG4k4B9zZZe9Qrd0LgZC24cS+tcvv/YEauTD+EQ8JdO15w
OshlmyYGqts1H2C+SDoeZCap7UzxOu1YUV+2PD3n5gVGPRbo5gosSlxYEjhvvKQoYMW4djUHnQBc
m7LuHAwCR3DAzKLx4yKxu77wCNI5+gWEO4hqXhVHiKl5is2uPjG9NvsB0o967YzLUMGmkREfrTh8
6ntwejeeIE772e693KCFy8nUC1RbXTfmmXKDwMleIYgBbDmhU88m42MYuu16EXrzuEeOysUtQILK
SkGrU1Ze98AFBOotR98JWXF31Hn2CX2mACweMpuerF7V18AjMmFP7wAv2BwEgbP5T8Ve9Ku2kzor
fBmkjaDf4AWSSF8VSGu5JEbbF0Z2LrHaJfplzDjIlJg1eQicNZvsiVTq4RYwCvde4rvcdO7IT+Qs
ChLPYhPqJNaXCf+4FZz/Gxl5FOk34qaiLZJQhjGidRXUcScfrpxo4IiMZ1TucgeHbsXJodLo/PFS
/m2Q8SP6liTXz0VPv79nGHurWY6eUUzGPbIsmCSV4gXbg1nYRy7cdA0fUJ0kR524Din9RAh9KEm8
CuW4gUlI/k/ALoSzOnPw7Tvqv+e1VZyCwHwVKQkT42K7WbGSqeOTVVFM1g2bNj0hpjgWvvgw/Rzm
Izw/vZd1TciFD5BGYR2uqwc9eweLUyQPfzfHh493F+y0hAp209kTLb5KuXthGYnuN3iHpwJa7zm1
hkqNVcuQJzRsnWWDEqLUUwOAoqHlfQSwGk/9h+WUrtZ0W0TVsFwuDOr5rIcRhOLlPTVMZLabhin4
QwJJrB3CLuLyxC6MO5PkoIHsXpNLKMcjxZ7lAvbiFritjJCn2rkeQMc2Wpwyu+WUYCfLMuIGY9vL
MyWitHx36z4Z+R9qRkUc1/2ucoI/sHjDv7AZqvJe2udhLLf7Y6ji0ejXsynlvs8yO11c22/P8CLH
JWpEYuT0gn7uvUjrMXEZgbmNoqrLJEqLB/cPgoQ13reMz6jURo1PVwjqgNlTzmJ7WovvRQI1an0j
UfZF6Haqe+ZLyyy8R3RjGnlB91DOgIcJ9rEzxkfHYWHVW2cfv9PEEFTOOY9WPAO7dk9jYeqgbpnD
R9Psu8eYrtl0GEOZZu4rUa1HcciSo+SOKBmPn1CyqJ73VK6EVTqu9wCWcl35y5svFEnte4nw5Tl5
H2aOa0N18H1pDQSkyH5ZabdjigDmuAcDFBqnYgFhET4E8XmlK1QuDwadIYuLBxYKB73MejvYQz11
xcfcLz+EUzU+69I27jOFw7O7GG2RSxV7CfCwJ9MnD7rAX7XXhxRFU8+wWvfU/XyxATGEljtKq7a2
aKDbv5GE0TBoGnoHB/dg/ZYhr+PJ70Lvva7daKcjfsNqP1UuwV1wtIMohK+gNYslUyWuQoRwMcAM
VMh7KyJELmYMfrcqiYYOmABmuaWakNEnHu3va+QeK7uLuPoSdgPo7dBPaoHi1MaNeBSDf1IGBtAr
+EyDo68TycLXVU8OeK6K8vzNlIcoTKBNWMdqUfpdGdTEG9jEWrbQHfY4f5hzb1iE2esu835NC5ih
/y8tIevEA1gYek0oXpr4dozpmnFZCIJeBr/raKagy/ogb4MMjQonfbE34wCUmzyq8mlD/jFZZAUV
Dbq5Wo43kpVuxYkb6XE4pmGggIDTUFD+tMWfQU/FEtyM9d4iQ73a726/9T1aoYSi2R8xapOmNvcN
pOAhRFfh9UepgzRXhDO37pODfGVVWiTrE4BP/ofKUP/K3jtwb7fX+Jl08TCurASycGwXjp8wj31/
KyNKJ3a6v7OMSIMJlI2tiPsKBcJLX018eZ5DpdLa1zGsqn8C23pZ236owdIsNpBkPbee2uczj50L
6dsBrP1ZSBPzxPRRRmMLTPyJ+UvL620crNwWuBtZoUCI69ipHyuXkH9RKx1NhiSKc5BDTtmMxaa6
nNuwZRj5pJIKnxAswqgJ3a6Sc+E1j6+OCB/7zrGTlv3hY0Cer36PONbg0ks2mfgUViS9rlSbg6xq
AgCrOEpkKTiXEVrA8Iy/wfJRaTGj1pBva5h+4epc9oPPgoz838/A6XgSIVltV80wWQsPpevYJNbR
vWa/lCOHbBU6OvhBDoWDniaCGBocZU5Jo35cX402lulyVeZwakbmGXYcVBtAvkOs7EW+nmkguizI
JGUJmz0NtnGwuAn05W2nXBhe8BAKHzhEOnROt1E3ScxTTtCxmOuwUUEDXqR+upbaHCjCysJp16bD
QA6rMu5qvHPpZOsuUwb+U5+/6m+RDJ1FPh+EXFPLpZj3LcQUtFGEsWFu1CxN2q6W3nR2Xhk+SQ1n
lqemY9fhiAxJHM2qSuiAVEKK+du5zUWdIBlPmnDFca+q0GiD7eTbRUh9gQd6rKZPB/Hl3xj0fV0j
MNVWRYNNtV+KjTkNMLM8O9kglnM4Q4OT+claInWWroWFy0BI4NZqAPO5WzVxvEFsB2lPcTzC0FkI
K1tXhTi3BqQqEeBuLsu5B9DrhGpc5frIjIfbOjYcDdJXXSNII1vECYe+Hf9uuDbBHmHzPNKZjHsU
Qf3lJ57I4C/qgPjjkyNP+9h1oRQfyjZhngHWnQ5QsTlj6/vU8+LcTkXfoUL2JjDUHJwFDikASoFN
hRnWfU3AxY16j2kZ/3aDFJy6a/vZ0DGSJLwvNLa8PunP/6QfLeRGLLhsQWeS3JMDCC5Fq3GEvKU7
K1OBADd65iyFwNhbE7RYf7QxM2hVF51yE4o1I0ApF/JmHIaP0mbW2hNnYmppyCrGW+d0v0c+qk5r
pw59JLsqdTGJVLJOzOFNkz8tZXpIltzvvfy6jMJ47A6LYWEcwBQTiKNjGJunAuX4kYeIYDvTQN/T
fIyqKcvRrmmHfEghvqoXItzkJvlPog4mcZQgSY3aUfgU/IoO7RYLOBpES6EYYJFAOFlXcDFeim9W
p7vuTtX/8VVnZ1Sul3n2QpnPPzJJxSbpKM2e8lh/+GRLY3GtE6Jdvw+3/t51sBvaakj1VI7QIKyM
dLsO7nuW7hwnxIPea0nVL7y8vparD+fY0qC1ne1HXiIRr0BQEwwcM7jGbYZ5laeMrbA2hlrSgjJ/
ieMd5j5n8VrTku+n7ZvEPpkE566JQsSiLzGY7j71eqWo+g93gpL1KffOtItHX+l1AMXtwT90Qcn/
Y1aPY0jdqySwZeXWbBxgbsOElkmY0PN9hxHEDtLa+NMzKyZ4P+C5TfsVIGKMkjlT+iGVh+Y7NRQX
DWWnV1xHNTWmvjyWFb42aBwoVnVbp5WsSbhwsxK1Rq0xHnWxUzkol9Q70FA/bHkpr9JvqLhInqyM
KH2Sb0WWH23nJyouSQU3Xh+sL1gqBVDsQrGk9f9aDb52VFwZnYObU9zOFpQfRcSorUKdRPVYlJdv
hsIc8G9Bgfjco5GEi03FmmEX/QjZ0wtFPd14dCbbGDDVlTKsrJEUa22N0h18zP2HYggLCvDfM6VM
JA1Oi6DDQ/4a9SVPrGxki9LdmcPNX+PT5ffRYb3TZKGAf8PXm6zq8BUuIF0yu6U6ETcEcBXvtGCB
UHd5UjmGlhQfh2UVj+zgKRCFoLD3zkdG32FOx+7Y+yoaFGOZWvo/QYo/o9t70GG/Ubl4/L9HZupT
VKb+ufsEu9i8dXWhMZOJ9aVAo4z2DAF7tZbqRs2ZsWicrPe6UTnrIa+VQLJ0sU+yCj0hI7v8+k/g
JP0NvBTgmhviQCBYLt4Rsz47Uzc19lMzwbIEjf+atG1LhFonTe8hUHs4wIxl9Cby6KwpGK+SSHcV
HVoP0qPWcWNeKaMJW8xdqSblMLQtZn2bBEa8Q8zxw8qc55vaoAzSAxUnSCI/btfn98lPAZISkJN9
O+lsrZy8GazbYIoGL8k9HNemJzWpJCqp2aX2TLYc75yP6QQGU23ItaTBPFeX/XgoAMmlQ37beeyL
tJWQZKJFO8hH2ujFvU8pRJQtSUVy9UTHq50g6oSdm32hX4PeXRd4oXyNG6xnp5+Yl78GvOlP2i3T
MAZt0pcaBpo6LiBvf14Dsf0NbNB4PlB2rJxESncvMdimhelf9T2KtJNQbnNUS9ss9YDeivv4d+Io
gCp+SrAejBqFSjSxoD8gf0X4QK3I+wNXL/dlW2vlvFG1ehzFGMTiw6w8jZ8dDwujqCJj5XF+J9dE
AhTdtVAsVEm9cmWxMiKNq+SA8CVSKvUUpwNT+Amtd6m4b684q6yxJmD1Os9+sjCtkXj4PbF4damw
0wf3EqLQn0hSVr2k3h3yVJYQRMcwb4RaqOAPw/4ZqcwMOKHx9rtfHUNRH5de0mwlIt+GPHP7pmQ8
pCmi5NrVlTUSAXSYOH819le5sCFtWOzVli7YV1+IU+ix2BFB+OKYioGJ7OXuyA+MNXGSjdyRCaxw
dnnaEJw0TVDTXptfu6/nH91HJeE4azjaKCV40b86EKSOrIldbA4nGoIeDvdNUGhpzld0Sibo864s
OScgUk/eOzOmhc/8bcI/34q+LsjEsCEAWupj1FrFlSBQVqBZc+O2VlSsCmGui1J2MMzrGxZ4Jm0f
K26T9TMaOPXU3QN29j/BP6aNuRFMjNLTFZdLdPT7WUpROreZzU6+94QOyameRd1Z2hlxRx4VIjC5
pI80xdU6cm7HcRHxyCZ2DzsWX1ebGRlMBGm4Atd60XQwAKe5tJMhDzuNF3uOSccBJZUCP/+DIFZ6
+lgbwqP1aOiR2pfC3QPKGHFsAdjzRO/39MGpKXtNg1Atrc+bFUu73hfX3V3drWIUmUmq5H5iC3YP
IUUh2Hl4DhVT+mvfP1VTIAliBleyMpCrs2iZPx4elJJcPMJPaHRDQNF/TA6M0EVJ7kEsdnve5HwG
UxZ8yIBe5g7oeBijCvJFt+qtoXW/Nirc33hdTOKRuNTqEOoTT2YdFGlmdk922IMj1zOkNQ01Ozhk
5DkkK64xSItudgASvgvamRtQerONyTYDkiFEdUyHkd7hGxT0qno26aHu/vXO/ICkBv/zfK+i7nWR
Op+pcCP+cwV5phxR38fCjPa4uHCRX9VSDIJF4z4pg7GA/IG7GJLSszDuCRfBrOm+hVk2djphgArl
NTFD9lD0WlnwZ3TI97ouFbM3vsDwAmiH/KMNcEizcypoIAlzMbpIhsGGB9l74n3WL5gQCf5iKkfe
fvIzY4IO5+l92nAeK5si9AvzMfFTHqCAWdv/+9fiko7v18206+mN4XT3bG2UeIliH+MLC1UnAWXg
unvOs2RLc32YgC+CsCtYM3cPL5KLOa8nSdJnSFr66LFrr3hvWvEnUF2ugLRVeQP1c3T7xR0aYRqf
rnF/TQHkhFwkC744ou4al0Dd8okd+VK2sV+e4cBngzQWIeuDoQ1b2CPA5f0z2VZv4pBAY4z5wiT8
JpSwYCE8k3b8ST9WGahB/GBuy4LfLsGjO76ZC62+luWNgZYvXzCnXuxKcTLZEKOFN/pN7x6OoZbr
a+SvSRYKUqTfBhhBxliGpvZ4uJ8YDwBiVK5vhJuy6JMIRxP+kWBlDiTHFE/GSrviM6K+P7ErbhvL
8N9686H/vPCO2K5E2UU13G93/YkFKWgwsgaA/Q+sgPiUpD95JP0Z6hFNjcIse03tT+3jhxwf1azI
ZiXWMbSNCD0bkVVGBs62fI8/Iv0Xdxt8tWj6pkZbe6ch840161kaT95Hv5eG4RNci9xlPIdM9iTH
SSKOLT8KL3Pw7K1sppvqS0f34kt/f+UM2zZUzOXY1xOBtoY3OSomloFBT1fZtLCxR/UsmnVc9pC/
eEY8pE/DaH6KX0l+ZNTb3jxgc/zh/RXO7fqjwu+8CpJ7Qg37QXTSZsw9H5ycLChEt2EpAJ25uvzm
nXpfCPZ2MAPLWCoQMmAO0F81aNb5imXE08m44FUrpuO6LlIhT4FYHqcQtnllPBhq8Cz69GRucItB
sxtLpI7IpCJCp+X43mPVuu3zDmN2Baljy8/1hLFtV22tUxZZ1KcaMWpgCv2SLaML4j3P+vzuYUHs
hy7SLpXlVuMojBVZuVnLlL5/6F56gUL2h0taSvtCBe9tRAijMs2y5aSjbmQ+6E1e8yAT/YoRNFyT
agB6h9qziQQBDvwMaTrFOEJKWTLOTsI5ClC9A1IXwrZyO+ucAVGXiPSHOKHLa9huihZACPL2v5q8
nrSJ5YgD8Kiw2sRoz280ZPEGjChTxOpVHeCZYfvy7ym5QFo7sG4IPKcJyUbOvnoqM4R6WpCeVpsl
4vKnlVZskMKq1/qrDneNEhunh5HBkyCZrGpDQTM+ywdHs/YcRIuMGlJr+u3ZaDqPAvtoQswIF0U0
hxqUMQ276Y8r4p89S0Txy/LJ27GMnosPItwkce5lorDRHNBA2I0AJYF1vUrynmCrZypcJ8YhC/57
DnhMJeLe+pEPtP8zJVAdb46Fg4X6eQO7MxIvrnExl4zBiyfUj5y/1riI8PXf3Y08H3bMj9esath0
eC79wwxzImpfdr6f7Jitl1t4giaEA07ck8rlmv1Yh9HyhzlkSRd/TRlosF54jNoWUnd6ljfvDHVZ
PHOmyi4fOgnsDabhJ5DNuMEQI5irdxQWmiO+XSq3ug0X9OvQxRsMSanOwUBCFVuNW/tNhUF+VHc4
WxjlM/FVZiWoNqZhw0oVzYWNXtTmhnA+xnTCoOaD/aON1Jmf571UUusXLIFxSAfoxPivkZdd1HBV
5eTggTlcHfmA9xBZdAR1/Qs7AwXTS+OKNIRvphmBlS5LHfu0yOr2c5JNGA4dRrc1Xvl4Md43o+yJ
rE89PSN5nIMFYCUS4+FWxN3WpVTzmFx9FAO6nFWCrrz5nuM9/DsYrtCV2of36jziD1AcupxhIT5l
60ZjpKzk6DJVMi+5ncTFADYAK/sozbrsZgJu6/Z+qcPpC3X5HwMVD4iPGK/DugtQHo6xDFJcq5Id
yEuMeUE8d6cGZIjM21r/+5qLr8OrI5RXlWh/h/NZwSY36cjjC1Snx8Q3m2Y2QS620073ODR+8hAw
rFUTX4ZD4wi14quyBVEBiwL7xlGicB84cXtxdJDZX27hLyTQhUoUFgkkqqv7pJA6A53jIllSSSel
bCyfqVONYFODmjEgBZgiVZqdc9AgKTqlY3HkfLkdOGs2jaLlW0T5VA7nvHZK4L12WLVLg1gmZkLe
LI2+SYzSysh9/gs/tApBWBiVLLJxnUmXT3bONMBh/dbrViYEzrGNdmWxwVgmS488Dgrkzsx6yVTc
00AJdpaSPwxDYssTlrtCCoJgH7eC7mT9IXLZoHAkOmTzLm1QCiORckmlolLNn4/Sb1ZDM1cYPyWV
7NQ/TE23/dTCFOZcosM8g8N0RE/1MSRxhz49RLKVwe4GZkas7EPB8qcKhXsU60vS7+hjpDFFHXIO
2ORvGvFylm5R8mKoWyDgmjnhf/r2enlIeKp9t8EhIp5AZrqna9bzUsDsDusVGgdeI7YjdWr2wzxz
mW45VP9PjrZw572KFnan9Kkv6bVPetTimp9DcOZ/jc91Z5vVtERaAoxH1+s7a1is0XFjaJNfaEIN
ZqDo0xtEpNJgpLMN55Ddmqhd4W9l0l/Bt/b2Iz1mg1CME/Wjum49pwj+z1otutTy2j6uWXnpby5W
LZMMCOzmg/BJwlSxxp37OZWpJokmoPaFkGryTUbFwj5USUP7qHrX6Xun7REzgAXYfeQ/a2d+6yAn
oMjxvU1N+Ae7yHPQRlVj12H5kWXaKAPt82sXCSnq8kpNTJuY9IuA0uUKb/sfgCf+Zjc2xyXyL88s
a6qEY2Bci1pxRSeMadnAm9P4eDAFbSN7U5YSS9dGPTwjcEHkl0vm0yCVn5JcDX0nUDU+UTzFvfvL
ub6bDFQxUOqixgad0xrD8GdSLs6+mfTF20NBey3XkfnMJWDH90lL0F1XCMZIP72+M8+AjO7uKFPs
gDtB1bqjZec9GBSsDMrJ61JjxTwzLswGvaNwGrDD7CsQ3YOCRvx8zxqxQb9pDZC7geEk7nXq9Gsa
CmY4+Kk3Fyr9LwNCtspFpzIXnG4hY5N//sO6gBWqqhMgprsHkkYL7rURIVp/3LjyLvdBjtmvp2Z6
2RjrmxOVzDIFcNmseJjP6WyA8GAuEHHhEIZThidmAOSmvxrxB27mUQMcwocIbX+5Tj+UbSSh3Lmv
rXKh7OazMEPbHF1zEyheuKzyF6JrzcZohMmbX3sq3yYdBFxpszBtJOPnK5FS9xu6U5gdnarTMZv5
PhEIBr1/pRRTyNuT3dr1ZfOajafFtQGiseb3wizTAE3hOZ9kTympSsdug2Ft6MQxUbVcDOYW6wHc
otgOwoz8EDH2rJ8KsjQH3tuNY5cH7dBK/MvJZPy9OVpJmngXBGP7PD5pLUQoH2Fb1iQWgLTopQ7O
khfpi4gnD+ApQZoFUEPz1lT7OMw8dwYfwtIF9SVrxg/4TmXs8c4aMDv6mo6UGa7LbTgKQulmT8pX
MRlG4ok4MoHTeDP57T3JqwUr1CToQzjC4mbh6MNr3Jd2xwPeURhDAmt5UoWD2pakaeNWexf5gjnQ
TaqpseK8pzZtFPYV9DpsqYHt69sk4K+XC8Uq2mVkBAIv42xxJ2iNSGfHN3zmzE4uTuXWcaI/2dRP
Wqx+tVl8JFfELLtD04XHVpf88rkpNtrXxBX+aJCX35xjgMQrxmC/pSgfCtBd9qFCxGRqPhhyZELm
tp9Xleov1tMdgoefk/fxf9LAOCREpj/Kp6eO232pOaUAN8AvlianlZxDr0Tr5qgWwFfa7qLXmFOJ
/sga/IwIusW5Y01uxySrx4aYUCPiSg3ArqQvrJT1YT90jeTqYS1ncxnExGdsmohQCCzjsR0dHl3Q
gaDl196WDsMkE0mOHxLtfXahpSMpYIYX9sssSGVdvNWz2+VaPrjWg5XdkuWfkJMsEVepD20sLRyK
+DHIGabNAnxnJKXN3Q3jTeL9HIwhiAoRcrHjUQvihS2Yo/FDQDY5oMsKbzYMC2M9OprSanriysPW
JVjI7ZuIImx3g5h0X3Bmq/WYY9wHFzTHzln0Tvrklcswb1+h+V1lcBudcdMuozD4xDfqrpuh05H7
yYljfqm/reWefB6Q6/DCb0dYfENV2CYA8Txy3yHzhOkZeJEi5opx8ZrtrXdyDe34dMPHfnxc93Z+
gaDBmMr+ec78Sku+WES/LAeVi2vw/VTlJFq140VvtcepWWDC/Hi0al2CRXFLMOtX3AI7DywnJ1S6
ZnG0rtExcKJA+o4BZ0DWFITQTbriC9cqEzaXG4mZaf4qpU41LKC/A1khlhfHWwXDj5YI3RCZe1ET
4i8alaDBT2JZ6s3REzxYyCG8dyd+3coeKjV+t4D/J28xuD20pPE/erlHd7MgCeC1t/o/SsGURh+g
93x0xhuAVI6NVywtai9IYWDrpXi85ea+9yQfhWvRMJKO2SQBX/d0UlLQfwMMVgJBFbRa7isGI3Gr
amiGAjlDyxHn4PeleFzPu3QumXLTf7NKFgZRjK4VfLAEW+SRwxeuDUBuvbx0/MCWinqRvCGaOI3C
z6JNYtSSzH+IYCiZRPOL18P/w5TOPu71uQ7ym+3zmzto85/qsuW6qdEWBm16WjfeAN/RFmtowD8e
z3SoZ74AmyPNHwxyjRFJ3e6VJSyA+Q8ZNOd0tz0kCW55eX42YZ9RuDVOCrwB3DhPqbqDp3yX0yXH
Vr3u0874IpcR84SkBR+K9/JAcra3/AYetKOWiPTQfhK3BPpgIiHYFaN53m15/DnsLOuwxGztbgec
ff8DKw6jzohMxW8PFp2WWc31q5zXLKnisZxr9YVLe0evjzo5bDznYdD35GOzobAyWdMGvsdbNGiw
7Ztdy8O77lMU8YcCuAL+HfOsSxk43U1jlfln5tPnxDkzWst89eNkzClI10BnToviA1ZLGBQWD8/w
8HLOEgGlnKzfdzzXFLf9KgRohqi7o37P6wUAzvGy8Td+ScFK40+BNZl5KM0wgrrXnW75c2ymBy5+
rK363WFVPyjVgv2Sq0+eprzhElwp4SCKBiCt2sq/x/zHUrnojJCfmDfyFR/PoQhLw8dsOfyA2Djm
39ZxxUkkHSGWFPsdcYNgTQg98fo3Q+0lwCONz6Nd+L5NZk6ABtfgaNGeHoQKCd70d1+O1feLxZtk
6kaoBN4kXIAS5rWfR8VRHSwVYyHXXgfIbVcXdHlDgCZMRnYdnMAl5mnh3mXejJGnSxtDVDJy8Xkx
bVtPggbomgcvnYRerA4yJw4+XTeP31Gm433tXLthVTNnuFvB5Gl2EuyKhk8j7pezEJEC2VMWzZqj
dQeY7qqiFbEte3o4lBWkSPxCfT/2VAdpKwXGjoi01NzQ6Se9TPtcaxP7uDRql3V9sHXoM6uReuR4
4+x2TzN9RqNG3I5iUgveIAK3UDYqIvgadk4DpCUQq4/2TJxiM9NRhIApi/7Z5BuY2S783EWuvJ7Z
SVop6vIeMesCd6x8uter1MMc9IRwdKGut9gMTCSXSg5c3JLSjq7lnWleNItsXhWsjKfnUAQ/cwD0
oct/4TihAbZDcTyv18kof8i7NBpwa7IAdlIndUo5x8bthn3YvXaYln3+Y2gn7ATjG2hEW+piYcLO
uNKjDdAmMA+qQzPaeQWxxlSefwN6p/o+fhhmpefSoLp7QccVLc681LKCZ5P+O82B0S1iWOI5IjDP
um69WU6xJmp6rp8QHyqoL/1o59+0V3cOMdXw/ElO/G9yG98ZR5VMiXKXnkl3YOHAjsA0CW6vENy8
bvQrQdlexpOjCeXY0bbgafYdJllPSasIqz7chGQTBm9ZjhR10xkn54XHUDgGJKpEJu2I6n+Fsjml
sGzMD0jjDkTgTeEgPXc0HhcLBunkGuYWxCkazrRzUCeLrc6RUXU3v38Uj2l0Wy9SXU5o2jg7+3Lh
CykNLGClg162pVseIxa7omVhnGNeW2jLmEdchz84VfZPxyPWYq1in9Cs64Q2oxXAu7h0PXgt+ibE
ooyqisa+0g8bt+iZ5es/rzT0GiPJbfmnU13k3cHgo2sz5XU3IFgxnjFYhQNDFAVjf1uDeU9KXJsX
MuPzHxyrpxaMw+pTBmuPKLtAN1OSM9ErxWoe7/zXXxdo4HK+FjQFt/cM5qK/IhAH5JINmCjRtzzc
xOoNvn7KxDB7JxjgrTi2KxRfvBk8YsKCIZ35cTA9nwqYGad2ZhxTrBHYctBrOFPB8IlrP+2CtnN+
3q7HI2bKnD//doBketuPPgZawO6Y6aaynkb1W6MTUsuoxJa3xepjUNexqwEbQ3CN2ya391a6W/8I
ClVkRcP0TJeV2KNKiA9Xqn4BwuMR0kEwIyzady83oCIdjEKrW4p1zIWeQoDVVnp1q1H387/Q8/al
d8w8AWp9+vldAGKa2iQyrqnl0tnluPJe9mYHcrSRhIraq9kLyFBABBcPuTVWwGhWsBfoV+G56SDI
A9HOdcXmxHpNuR2zgwQpv+0bnFE2TdJGxgWrjNZ0pbCfml7nJAKaUMVrXv+p5YxgjeoOGo7jB+4P
fd2VxEDJAWJLZa2P/GFsqydfdRV23OV4tx/6UJRLRmfgIuIVjwvEbLYxGv8ByFPpZ1dxAVGAXAZa
g5yKQXnT4YPuWpxwPCMhgcdmMUO9kWkpvoW20DtHVMz7iVzjA+UxJYCkoC+HwCgXHgafFes7S8V4
UkjTbCCJXqx3HoYTg8exc1c3+Jq5SkeMMSUD0EFgb882PhSC6pkwEdTY+y3LSqbXxzIeqa/MTEZx
HXAbVpY7mmX9haERfdr/KS1PfYL6ZDPMBo3F23fqwSNkW+fQZPMVU/uEblDvtUhezxg30XGx/O1w
IW8mIE046LEM0ueRsr25L4YbNUdhr0gF1D+O+r/KRNyIziC2BMsCNMKmZn+VtQtjYuhNOqk3oeTr
p3RWDzPbeAGg515wByA8q7ySpbOu+RDEUYhGFldse2+2FD+NSAe7xmOk45c5LLBkegSJDEUkLF+J
22VMynB7/kXYNsHuinbgulZownlXUr4+AlSoOt7iBn7j+l3ga/7vaIY1zHNT46E8NIeUximlAxDt
2cM1Fe0Ar6+k7HpG7ViRMZJNqRLS+qS+7S26Ad+L+xDjCJClq0anp6tJNp4mKW1W/4JoS6JAqiVe
/veUCE68evTyzlr2lFE3Rf5R2KkqLkr4SpWi8InxTEMtANfAfdA6EM0O4MTKb0vxiY56r8QGsFZU
679NHAuglhtRZxo+JLydKHL+zlzXzWl0fPwgBb119QUGDjCwzlaA447h5Otsh8Jh3xdeT5nbEg1t
EgToYnBUrfZSCo9Ts/9Lr2l8VcXiq1IvY5IlHr6WCmOMSZSgIcGwph5CJ1I0q6Vv3A2vJv8CN2JX
tHqOmqNY+mwsJF+sSDX/OV//Sy79ff/Si71e8D1Pr1wH7q7RtbYViGzyCdUmT6R/KfbzMEr0IrWU
YccfK44rq0fP0tXoOZcNM3pZdYOInkgfZ8lhhh1XD1N0LwYqbM2+Cblwq+y8lOEKJCAjvDsjdk3Y
d5+wjw+oq0XkcK7M46WaerNfUaf+mr+5faC1RkkKj/GTDKvbXgcBt23yAqfewygZV78fpCqHV/1p
dLWFUzIIW0snQ3VE5Bbri76lZsgJv8wR3PEXGQLpV5fujkZKHx1Tr0DRLUKqZiDoZAJpfIbJb5zf
NykQNnqKL0shtBvjA3nuSBrp88UPlkH85n7fV/OVb3LKPK4ktaUE6CBlAsW1tw8X8BdghaRaWrd1
WsTbONwzIb89cmPymWmuWMs8IeObTszv5C4K9+UBrVBfzLSgoPsWWsfhghlIxEZcXdCgP9wEwn3h
P8ckxwEgpuUg8wyEA0k86r5N4oSgs28ToLzlN9jEG8A2M2D3f9L57Nlupp2lbnO8Ryj2iNo7T/rW
SmjjC7iJbbH678sANlgF7P8tPm87b68hX8nuJp9hYRqdQ/wjHTBlB/Z9Cr7R1kMlFGI02p5x+iWX
K8bZ5LILNn4xQtLJCT1NfaAo0YkuwmawOA1tNL2CSz73pVtKTVnUD3wT5lqStngEQr1SSuKCN1jQ
KL9J1BjEd/pi8nz4WORKeFq0TcYNPVXouyA5LtRco6kPziMwTYRPANHBVLK7r0gtoKaSHund+zuH
2H+POWz1Rj4ulz/PNhZSZZiOzb9nwgruwq6ewZZihHj2W4MnAb3OzI3+t3tEDg30g0uAsgbtv0BJ
e7kpJO04rW94op0i9uWWisgQEF6Yip/A1ncwIxO5twzopABrt97XIADThZjGadNYET1o1DynU4rv
9yKmzsjuF8ZN1/OCDAjaDFMOyCRqt4wspNNQG8JuySLzf0w8h3+hdNNS0g1PM438n59bpn8KoFqc
IR/lIujPdTrhC86svQiIHy/W8JSCx7qPaavxJTU0yByEz8VX48IBuFwiIdJdxObdu4m809ZZsRth
HXruy0i4nSwBa5NKXZTfCIYoN+V2A1eg4TCXV5MJSQQd/VbPBE2tV9KtHNw02qAOOWETVocXkfXL
SywuTj7182pDpuG1j/r39Z+gkBS6bUUtilFyl68Qms7jNC99znUCkpMTzurJGkCQBHanH3cHlXgx
f+8w1Se9rR/OcJikbdTai6BXC5kVz5EHm98i17NU0WZEL5dbt3aIjVKca4VwAcQGeC+XvvX8NOmV
vs/0C//v7BN5UNQ7zO2jLiZzspdnETWB3CpA0uZhunmCsmu62fhH79bsYVsyclfMM/euSZsQ5848
zzRWsoTAbl11xJhWKYbOWB3yqSmPfSLYuJEPzlc4tkKpFjivwUatyA0BdvxWIKHTOndfS1C1Ih2M
80HIfqAQQFLlWG/hmCbTXw2zAGlD2JraI7WGxmd8n0zHzxU6PAYlCNvDV1A4txlHI6YkBQpjsPwP
oF2q9n8Ld2WLrWi0ZwZSjuDe13DCmggvLlWLJOHuRFbifgo8ZpTZQSOYaZaH2lfyD11BxWL8KM8S
rExKAL6e0dhOwzn2GoyoHVHHrfA/210CaqWjPRVf60Pfxe2D5DAiT0yuTaKtsCgllW9X5SvkYqXr
abNKMASiRTJnvKi9eMflgqMTRHFo9WcXpk1+Xb77jZokBEV6yURV7kKK34Lql6PvM0cl88ajozRt
pqtHcQGyFVJwSSB8RzLGVsCJthATthxAZpjpQ/4oXDtugJWT1AN8x1l2Y23tZyIDc5+wqtinOgDm
va6FYb2nAveqMMKmvk893lwsSfuG/UtIpoCnLojpXtuajVq2jbfLu25l/cGMJ0Ig58qXtkNrZ8Cy
Z88Ejd4p8gD7dZxwQQoYzAzehlBlPzr2WS3GjS6165sdB8ika/1Xj7cnL8CG2WL3e0U4BDKQtCah
33MVSj0GWrXqUWTSRhOyrG84nTo7g4x3u5z1IlVPxbUznUcRWB6SvraF0Xrb4H+ge1/ALc2wkBuv
cBwUWFo3gj6ev699M+S4MhHb34C0wrLusCj2wsv62XQU7cwYgEh9ArQ71fSfhd4nd7Jwn4DfII7N
dwoDBgrj/oMGfpFGs3M1sM7ZTpjprIyRhsfkKL5hFyLpA1qmLU8KTF72/g/o6STnPu+J+FtGBnRg
CS7u/lSMXGDjgMkJthBt8cuQoL8pzQKDXzYZHWQvoTM6QClSYYJ/Uz9bKcPzWjoWdHu7pVgvpsWy
NBb7JkucOgelRxlcQv2c0PC4eC6Ej5jG6MwUwCg+5/xd2tVuMjiIZ9KbLRX1ZDTYJDPlExbS00tY
uBK16rWMa2OrZuqqYkaDSH0nNfUqCYevwhMj3wD5jjmlKsIYqRWeJH3esnFYPIWAq8yIZNxZ7mKX
UDzFe2hh/4iog19ihMlBkqlPIZlxX06Dcjz5FWPhrSRtJXQO3yqfxpKOM2SPg3o6UR6s4Rrjfjrf
V6BiFjR/vNNeA8mwBHj32jOKXdRAY7A/qwQqOSNQUCOS46JVDTXINewHAoLh3X709ijbacjd+t5h
hNSW66U0VAJp04Qivadf/D3RneJLLrQVS7E6EDDm7iZX6qhyxWHWmsXEx9T+xZ4CC5PtUhospdKr
qpBBlyA3BfnGszMvIlHdH3+HnyfJ8V1aqk66K3TmrPb+IW1hCgaQMT6ZO3OEl3knRHS1+ad3yUgA
n8AE+wKZo88VB4aHTyTvtZFM3fYbzREs3xSq1uov/Rr+1gtQqc7YhNJD1BZKNHnMfGKBKJIzBK79
NMs8VRtCZIeAqCXC/pb3QuRvHkX9Igds77YuNEomiOcobB4PwM+jxsT5qpMIYn2gb3/enLWuCoGm
ujpZBZMam5C4W40e4dpQKKISgdSq+0P90IB4aYxAu0mOVuhOJPjhkpWZWkLPr9LTWpoS88L3m5Mf
891lcDCTEqsE9x7MwLXjdkwZMgiZGHeVMiF6kDZncvzN0pZWoIIzQLF/fT7Z/kls2DUP3BWgiKW7
/XADw7S0NhG8VVGbMsDTP4PHRweFLjFvZIVZ4pBUOMUEsSaj2D89t2+vDUPhLkazt+VPiGoMhE8I
aT0sZcHzSpizExPPjp/i6NMVowfeflYDwGg8Rz7Lf9KIZ9XK5xlA5bV9rwVE0/NwRUvaAmNfSgsq
4vv/V+b5bZ3Te+/4iD8cOskJAB8Xu/X0qOrCvVbYEmObcF3eY+Chn/kFywZ8FgbRo1fMkYkYG2Y9
vGp4T+cd7Rzai9J1CxPk9Y7myryBe3tC48YYvz+1XC/cZWMh5arovaG/T7q6x6wgDIJtF/t2xfAm
+DfJw13Hyd15kyt8Zhzc/pw9nh1Dce9/AzT6l7DG+MCwZsqoLXndkxImNDwNwMglx6AjtmKpld5y
3NE7wH666fTGWofECaKZxmFYOyzHhtWPa+Pj/3bdl2tPjoS9Q1WA6zOCycKoQDFNoXLzizvF48RH
DtCdoeSa77bLR0nzgRdv3zioCS4eclSznI/uypE1SDbJagsm5+ToGPhjgfqLdS63gGCDCgTpmfai
Kjk0sN+EvQmW2I1YTyjd40nDKXDhiI/YjysX8pLl9I4q2wx1sELNl5uaFjBUZVG8AaQUu+z8zGhT
kD0FuPRXcdTNMYlF7yR3XDC6OLNmwiDkG/CgiHQVTAoq7KFmjCREb2BsoLR3lGkL/2AEcZMQ8ixm
ek+1KrL3zvqJB1zkL32x7VBD3DCnblC6t8EDdUsUnlyAI14GvmBQFDzDMKch9VAsTOrYIBkjcn6O
pLC5+NJ5DXC2cPzypVyQZLF5jKlY9/wkbly4KOq/N1ghMV/xnhImA0Z8ouj1erlYhPaNZ3N3kMQG
lp4yUoPQRWpbsw9ViebLwkAfTAsgtufkkoOzXn5RwcAGb8MxFIR5e0dXmJbU9mv063MZeMh5e7RP
zCzdFIvsdRuoVNWN9KVbLd1y6kXNuA9dVRwYzUfW+JGUaje/4Hrhv48MAR8RNfbDdTHC+8JT2+YC
51BZVDCatApjg7W+ijtb0t9zYWYTEzM1LvtvVSwKZC4DdbHW3HgOcnBkt3ur8teijnZsZuAYJa61
trYeNaITRFDxMf8+gICYcG08l66hZR1t5k+jnGrGzFec16LGlNEwnotxA/JNh85NiJQSfVUWwRHI
Ms6ILXJLXhoh30NVLL8kab+euztMHVjvR+DVP2togbgLcmFt6sC3ymLFQCuTm78ruvl1Z/ITu3Mk
nW9HCo1dGvDWJVDzwCh8pxam3S0+UUSfqqOQr7USjQZxcaRu+dnlSqL/FhEej1HKaQLyhQEfRJER
wdnvHvDP/xKVgd5lB6dP5JXfD7GrhdyDvAu8JhrTGPQBsc1S0adAljtdwYIZQjg9LRkSxfoE/xNB
EuF47TxE9DEHvIvaSepb8gs5eiLa2KtK7IaHFh7nlFJqC7J7b/Arfl8LYgHh22BkvZCLY3CqZ+sI
xNL9Jz0nuRwO3y8en/g8DcHKoRw9IaiKfWH/OAXASMToLjh1Z5m0xn0CHVV/2yVbn8+yMe55srDZ
At3n6IHWNHlnPrmxQVU9H1FhpzrkQqZky/ZUG+BzgNTq/8D0a/2QFFoMbjM0K76cmlAuPtdKoHQx
n4DL/ACwyhk6Vfyyriy4uxqeY7qMDWcYUQOH+r0ayFx0DcWhttBMFRXbhO3t6H1FDtm92hdUA7fY
iZYmoqQiZAbhV9aSEvMy1VlFuO+eO7CSjT3UwjtSIogT9W2EWx6dENVvpBG70CEKBB8bHPOSJzHg
wmhmhcvJ3XtXXqmlSq1tyKOvhSd83WValtMV0cFc3u/GDj80qjgtkpn+Nh4i4qMXF+2HMKWRSEMw
05ZZ80M8Xmw5RsEjY3gjvx/wx1fWcsCmq73Y/kBEEnoOLlOnB3JgXilRTX8mi2I/t+eR+AyZkhX3
MywKVtk+aKN5obrZO1lRLN78E3MCF6uvQR7HPTwOwxsifTFY7oP0dIAZo+RIhvZFfPg9ZAfWBLoy
UTs/5LQnJu41YQgQl2wIqp2HvVR1iGxOiIw9huj4Lx8jLEgiO5PTg3icy9v/RMbk+QnJjE9LNbfI
V6KWgmivCl+AX43V5Pxok7MeummeMkGsqAjvNHx8fiudQb/ngoLg8pnVHdpANpKE7pSZF2E9dyYn
2Y5wOWaTJ4F63meiLEtjkrAhm7eC01QJk11tHoLIHyBdeHyERnlaNgG+CHyupb1AiUBxFf5ot1Yp
Lz/SLppIqxwrd/MS+WYzOYJiv1GK6cSlMEyi6dbKtqZEPS1b1F/b0pDiL3AtWidXK2Xjk4iwwZb7
SADpWrRQTU91skPkJyqy0T3lx3xgX2KCRNCwj+zL8+qOcq0F/Gqxc09Mhk54VdhbxbanM3v8sGcm
x5BaKDkcv602vZ91l5O/zloj4uDzn18CWQ8eALU9tqgKxIRcBlEedQWKHp2le1aGub++m0NAYLwR
wiu2/QZcfX7LXw52RYgnPR0bahO+uW1xQI/GbTDj5Ief0YgoErzbazfCBvA/PTvHYZjzYoxmXe6i
JzOnGpp1XO0sPDGjcFzYJircsMPqUbRfpAxeHNRQfYvYnFkCmiVzU1oucRgGVuZH9eU6U56kvwiA
eojbp/UJQWrNw2D8/KbjybVvgOtt9cBFw58FOaQRH+RXftGS8ud7vxWjtbyeeYa6oWzZq+zmj1LO
s1H/iDyIubLUDpzErAX8Ci70AhHY20SwRJuax9iFktkhAq42xOf5p7BorLr/JeNgmbIrWlkDgCh6
/sfXn3hVb6wYgdqn4g4xgY0V0UAZEkHIP2JEnGphldp0Md5dyd+cVLAuDyGTPo6NLpvsjQyY71iM
Ym9taP1svrAjB2TCnEdbnyxYw2/QahfK4NdNL/l261gVTVXPcvu2HVzOWHXhx9AbY1FwBoAqJDUo
oWMbUptobzXPdMSxnN95vku+Asbcdy8g3vzI6QKxHBc905diC8toFIF0gNNpHE+fZTH5+9fpvKe6
qyQ4whK5OT8jDIFIr0U0STSA/pgv8JDzkVMJzd/8zk6aw/IfI5KpelStL+9nfbP04CNAjVa+yF60
3GPdglkfFaaMep/yIBJQA+CAnwGAv6pu+QUehTuoo5uwSZux1HgGC1Uw5Fw43qEbPsaAF+yYTJsy
gjLqNdupwAUn4P5lECnyMx4fBwLYYUl89+SMWqVCMGIk9u/Kwob52/Tl3UU6gPOkvtVa1XvLk3dT
X7+Cve0vL3ZrLp7A48QJCMZqaQIaUHBvGk+WN5QaAWKZ0Hn5YQXlamPTdREV35KIQvVtG1Zufllo
p/09mwX0/cKR4c9kATLA6s0sn2cthRLXfI+abdI7bIQCTL8mU5BNUqMgL9NpgSNz5UWceMx0ojmy
eSIZ6InP+2Qde73hh6h16tPWbnH/8X2BjS4Bf266l0dk3M0IxOGE6tKpmT5rVB6IyZxDbpaGKuiG
t4J8RhsSJcvHkFtqcu28PQbwOLsb/X7uBq28Rzb5KuivraFR08pTOfFOpo14J5NwY7Xwhqy4n2QC
XdUr/bn3IDDMll0WZbkHoV6wjPsQUfSVoKUIFIq0j/XKxTecChKafpSmQLOZ+jYVYUmFTGkkLJeS
BLwqQZJQHQdqGz7Fhf89QsNYvOtrw8xNzubO987tpD+5elWjqyRjclRrdlzOK5lcTklFloOwu8uL
O8EY9ODPkaOwLVIoas3fKZSYDBaMex0tQK4tcNGrZ+WNuRcqttDinzMP9fdvLYT7NPgQxydjEzCw
Cj8AMxBvQ5I90+e6YuDmKHPsVgfaH159/9KlzyZ4XEda2R51953zjGFaINdmj4KWSivDmg5RnvR1
/gGZxwajUfMou7B+eMicNQd6KPdlUZ2uNOtC8HgkPRrS6/RX4eo9pEeSm/HqH1iK+UgwRQTWqXFG
uuVTRcywMDFbhC/wP5McOYHjoyqd/vcy3QEhqT8nKF4Qzl4SGUzt93J36SfepYcU9v56PnDl0zDU
sHMRyiM0ZMCDafxaw0FpdjPgkrbebK1mj3C3tuOGY4U9asg7geH8iqKUDxdptMl5rZDFVl2Ne/ax
ZgOYAFIPSEcLMTpASc63fg3tl5UcrQeIi3NR6txuUZIVT88WT0X0yfTwohTsdTgTCoxT8J7yfcKV
mw6zAgiXQxz05agYAaTxSuUZgmgtnhvNqiCw+5Cai2g/vXVps7XAGzdnai3UJ5h94EgnsaqiDdVG
c1OcVvCdR3cSSJf57LoLlZe4G73l6bDCfVmnngZgXwM612bnhVoV2TKxtl27m9d9c0SwooEVc6+L
MMQVvTPNI+HKWKl/7TI0fou/3DdxWAmA5lsDp3gHhLzxFotGknYHmKCfXzr3FL+B2KepkUVzOUcN
vGGx7M+fLveKdteiNhIYmseYp3xhQnD48cyAm8y6xiyEjUGTvonyxk5c+HGkkPAYdAmCKf4wozJv
wZpImE7HN+aPkc5Cc2AL7sPwTqtY9559BUCjKY8Od93oOGnVRkigStJFhApGuW0RxYnEmZgHvbCv
Fd9iYnP45zROVWv/V/VJywSuia5zDnhVDda/prSaCSuEjR0AHMBlE0AsbkoPMZgKeYZJIlvEdO6E
zScvUE/hooAi5ZAJsGz4sDMgEsQwQxnZ3lLupUWr9G/SL02KQHygOzXT9nD6o27X579Hl+g5MzZX
zOts8m9TmeeGGfwpWmnLcsbzdoghXxKY678LcBVu5HnXBNgBLxrnrMxErrEaf1U5KZyB4llZyNSm
unZtgfLtsZTUsrTJktzZgbUwZFry+MG6vPnLXRwSvHzTBZWiauGqRh0ZMKqUk2C6vz+TLeCVwhPj
3nPgQYKc/d6NL60sBgVoBqu8LL2NbECrVwn27dwxau4aL1OYsUYW6W7/PHo5lb9+UUvn4jj6Bpyy
S585xUqbetTrcbwFYWo+mqdWUpQ0AsUMd67Ps3rHFxtridMsv4ho/3IACE2zXtvOJbs9aFZL60md
lwtvsMi/itTw4eKA2kMcLp+DAdMU1JECJ5JUg83CQw2qbhklFnXNrIj7MrjYqvcMIdH2ihgVSK+I
VS92Q+h4O+wNW9yJ3ZEYKMcWvYksAUa6xlSOUSXRjzLCXgHnF9IXv2x8tabjCcF9FjSmCTVHSJcU
RQ3KbReka7OHW2l6XEYPYPm3cEcNKMGdRloKUrez4n90TFyJdbI8hxCb95gZX233+tquzbYp0+jT
KcIllxVV+oWbvo8RY19leM8fG2cv6pfMyTieRUeDNb/k/0zkJlXTzdUsFu1xdZM6C+UkRWeNbp2S
2nRHK8iuB9etC2SAn3zpSWhSj31dr0dGmnJiyWCRjgHdRC6GLfFkUefIs1RhRCOjY4fXfDgyXi3G
fvaeYbgJRwc2u5CDZyV9FohMlhQ7cFPef4lTtsNhtUbUYpqtTopCenO3+CxL9Fmez1WhjTzt4EW+
DO4VSuJyCVY7P1e8VUfHavX8yfRI+oSIctxuZiW/oLpDBWlTcH5L5GtaZoy7dEHdqpuxGr2xOZFM
0HqMr/sWpgkadh3dP1ZtbtH5YHcQ1Wf9KcAeasoVqLNpjELMq/+Z/vY3+5YfiaCkZvgQV8m1kPBS
w1g+MxHs3Ps845LKhXIXNHUQ8V5E/3PlfDiHJr2hkx2AFIwE2LbsEcP70IcdKhXZGE77U0IXA6pY
7m/ZDJuc2Kh1AW8mMfjQR9uIJUEEq/Ib7HvP4RoWAufZ3hcpRfx79vVySHVyt4g/zAbWvcuBzKGU
CUjHE03LoiA0mGO9r37wxZ+flNU6gBdExkPl6zqbWi1nn+N7wlYS8pS+dvyfzqgq3d+vSoCbFaBW
nXCppd4w6sXVd+YROFw0KvlX29pRLCzL3C3UcGJUpTmpquzjun6SYlmGTZZkhzfTCmml2PZTnveN
9DtDy6lXfD12cSJ72oCjY6wiC3u3DOR4YRacNwSY/PSxit+JHmB6lF8w3fIi2meBgtltIbIc9oW1
Eqbn4U97bvPohGxJ5DSnLKryDFxojELRlUfyFeTb2/rzHxJI1EAcshdtDX9nhd2nT2KetuxPecUw
/HEglEHfbf0W0SeRmZ/Fr18GApHl9j9/LHFYF2IY5gPCc1++8H5Iri+WP8eNlqUJ3HooFeflkyHI
ceChsvpbQMcCR3pmFlJzvUrw6NwUHBgae79jkDueMCJj2O7nBcneFpslL7JJirIAY0vKILXmr7GE
ewcL4d6UcmkNIqmOvWTSb/3kho3Vik7ZIT7PW6dzT7a6GhOyCX613KTblD6iPkZACaFrY+lALc3q
49XLBWh0J5GYyRmnX4degKk0MjXgHp9U9OwdO4B1L0iqWnjSsspN9bAcGLC9sfO0uXaLGfc2eslQ
yQELavK8GgfNirPNzIo3Z+92xXuEoS0vZ+KV5YWg3DJoH4AJMEWVjhotzc3f6ME91qTvtFnDJfti
0IjgLuQiupi1aThhyEXNWatldS7G0frWlw3rdEDweOs5vftb1mruFp1v5D3SfalTQkt/0ACO9beq
OQHGSc+ecFPJeZDWpFmrPDnVdqxFwvbkuXH/bNJGvw6KraufyVkZliXCkwzL71DMhn/t+clX2fNh
27NiAwnZ7Ay+2wLVPOB+Z8Lz8dRjoyuR2yqMwUrumrbYRxRFLjnWObqBRwwl+ZIo5XW8AN1whUDF
NgMlcNcSA/smQSTQqdXkSM95YUzQMe+qoIdhAtuvhkbHn39VuaQUEi/bZ1rnb8tdYYJuv8BCNtlB
8npFldox1KJWB7V/sV4rP1Lt9s7QxSj1VCqdx5c6jzw7KJ4/R42Jcz16qo5v7yyy2cJYaNgiLuJU
ahUcFJ9bjGxMe64dxuG71mq+0qGp7m0HPZFM0tO8e3NYBRH7e6jl4pmwBLyE6+tWj7doWKz8HQbG
7ncohWNLjkuKlZQ24uPrrQloWrcjBHO+m8K9Cr3hIxySBfXDOdYuHfa+FPE93NcneWvATP9YkADU
sTYy83NSDjpgj0CsyEFttxa/1EiYjfAP1ErdJNPW9NxnzZ7TFydezUqJzxJaWUAUTpuEbkWRNITM
jxC4Jb6aHT4rjSXaznMLGO087iMRWbmaSdvZNCGf4Rq7ezFZl2fhZijbzS3UNCPd3hd8r0YfAvnx
SmWhHsKaw6dN7mHAK5uClcZQ2gBbADjnA88PopC42Q/7aDZjTyLBBvIl0zeb0bkpqHPCqf+3qV15
EuIya0f4h4wrZ2PJ6HagvzzmU6wR6oQ02T9BdJXrpCGBpGyQk3AvmZmDZV7lCY/N/eBtwBcUwQwR
MsRJEsCQwgwHZn93u5iOjeHQmNoMzkzEzjlOAyEt0jMxClmoNdeSqLyXRgmHlBIkyQgMrdTNCDV4
GehKt+96irQPWfck4s/qrIrCcKN8GpKlOwI9vFk0Fto+cJSPfBYBBZtpi9/wFoM9jBDJyXtwT+CA
2vCX0XI+SnreXWClI6Hh9B0RnpC5NxT9H1cHq/oH1f2d/NOKhaJ1QP0tcMNAISINmiYmgofrhN55
WRn6wP/hRUiFYixvbN8I2pPCBJFYytG7AzT4tRk41g/cejcSV2i3B4fVN+FfzY26LJejB5gvogoO
yc+V3q0ICCyAmCeUzlh1YUtX5s1RrNU7J3i3DANJHP5H9KN5zH8fwDvXbeKMEifcZ4X7Xx/lC1rw
jX8yf4Zk51wJs0CVEtgSCj27K8v60EdJPVK1N6Ggoq3ZljuovrYYj/9Ym7H5/K02imleAKR8rXit
UfP2AVeuYm8r611C85EnI+mpZV6Y7Ue6cbL3u7Sc026oj4br0EK9TCcbmNq37Omk7fgtRkrKuW9s
RH51I8BSIdmrpf0/Yc3HS61e0KNi454oU1QEmi2k2LQ0XLo9HSbmae+w+2RP/l4/B4OMlEoZjQBB
H82fjx+jzatfkvseN+lPcPVad7Y0cI3FB4ghox493wlAXh6mwmUmAqkcAbtO1rvvd3CtQQMPwo38
nem3WdESLleOFOI3RMEMxt5AeYhqRencqs1TsCSbAvtEWEs+F83VZP7PPxTVUuiUFaWR2bbZRO5e
W2yYZTrwJtbavyxOKFkuoSGgY/hHpIvuCnbdXa0udmQyuTlymmqGvfEY1ZftyyAYDI7PNVqLdsKs
mdf5p4CsM507Ucw3FaCuFynkOjwCgP493+fphQ/kLQrfBzobOgoDM9EtlLiCnelsp4TxVAL5x3bB
INqAhJppW46R7mTPZ7SfyGXGQruNmvO+SUOlEVD7TxmBT5UY4+giwUZ136W5I+DOl6Lww/eeGKca
QHN5eukWG+RUoLwmS062UQa+9GC9nLLQbnmxw4q8tLorUctkrTi1mIAsZZdv5ASXDh1IE4+79Tg9
y9h/54FnaO58JJ1anekcEnfowvu3cCAucepNCmjC+p1fOKpeGwTxMMs4YHiXbTd+oYxI/1qB2kDC
xVeWOGqk9Gv9wioEejSp5XfR2ZE9RSrio3NtJPWbvN0cWQTfjov5eWOjjuKFYldTcdYfymvvB9Q3
UPT7e9kw5zSbIysSqeUR/62dbVmYnoDJs2kno4JijVngGy3wjyq06/gU2jQPyCZu6In7ao76zFvK
loXhmpSpNbGobgCCoo2WjYyY2zeqVXgzIN1zkXRaPAAYBPc8AGxhrX9e4bjrefitMgTaDlwaV18K
uJlO8TIODzeJ4eJO4ZClFRnbR17PLOXgj1t/Sx2WSo51bpLAi7nXcnQVMFH2D0qfR/AugWTFgH5o
OoAcbw/60ufNe3xFJKQ1NbaCtqQzqv2S30EiMoH+7qdkZAwMUiiyIR1szfJ6Cuer6wUkhHo1NSzG
ToE3CB1VUNfYQcWCKmK/iNz6VdsfbiqItx4YjAuSKohZmRnea0Z9X93RygNU9TRIbzkh+x/Wy1SX
tobFfel1n5neWLxKY8PPl231AWTUuMgxMXt6quYFASzJKOsY2tX9WQUndOG9pODIqPuYkYrwkZTI
DORS/O2J1BCHL3IHhCrOk/6+aP458v6lljQB4lza7+wdxWMMxx4tn3e9xnZlucYLmkBHuQiuq4bA
JS70p4uffrHQT4U2z7SaBp5VR4wZDQ6mCgSMpwtXQONCfDK3Aj2TKcH3Sus+CAmV6QSr1NjUazdT
eg7gXqQQ/RBAtbYDKlDLfP8Npvo0nFWxBDrx/TFMQ8fb/W139HPu3RAouZumyPL6bioQrrYfy9qv
QG4l7T3htaJwhb5uEcGFR/e6Ts6pm5aLW2BxnEySgY40B5QYRTi3mtqtrknkku5zHG/SK41Wbe1N
hXKXSL27E92i6PKdJXn4ad02+NfQtUpPYZiNfrDnKWVLQneiFwhxgA3jw1uwdEReMxqWvu0Ac9oa
/rF93Ubvo9YwlYTU5n57M/rj5yBC43G8sFOGnR5Iab6Q9pJ8+4ziH1e4IEaI6lktkYzD/3EGrcc0
CHh7hnmwT1ohwcBC2CD6bJm+k1jRFXE3LFT3yJNnqiPk0kZzbhAjrnJ2tX3zDz/IWyTcqjtE5s+n
kOTQNLVZjA1i2JS+eELXEInJG+khTxDU/7oCsZB7hUAawLZ2SewCbb8S9LaAi/EYZCx2pI5ZLXfk
pbGaNqxEgJevFBFrhNk0Rf66T2TB8d4ouI1zjmGNPhdw973xlSO9Wilh9LQXrGaYrsK668VRz/QM
8mlVyLu2r8+QfAoyh74/d+SvPbwAKUNxOPzr3gybziR28XIi0PrgPlugF5GjMc2ccTS1tSgpHmhk
jfhgFkaF+3iwDQFZ8cXkYdbUU+NzK2vzMCxSvMLKi2kHINXsM75MxpaJfYHkGez+IQj77dy3ybS8
9IKe1PDi5sjlLhPFnBHSawm13wOfLjaYStu7ZiQf/WEDv+D+lw3Wl2ZclH2cgC6J7eO2BFelhhRy
ahcEq28V8SH3Jz9y77n6ZjfZ00Ds3gGGVkmwmG+b2vt8Smr243+5CkMTCEs+g+be9hqC+y0rGwTO
kO6NbAvDSzEuM1eqxz+zX7y21q0VOa/ZAXhU68EFJh7suuRtiocNZ0gx9v8+T2J8iHVx/dlPGoO6
i1TM9OW/ofvAPP6YG6zf/FmVSPkC2nZaP3QBIpnywNZ0KiGNZUbxve+lyHlXNOVwppKXPu2RASQ9
H8/9rQqOebuxSwOJcQwtK2GV7xV8hXuBnQtBgy2W1mke+Gh0VJnh6AP0Z6IthXy1ks6qQnRbaVVB
d6eP3wq5iI/4Hv85xAL00P30Oe9eYVeKcma221YtYSg2CXd4RvoDabr66ZRK9pUywJmpww9TEJ3S
ohnTMzR+G8u16GJDlWbVAYks8URdl8GtfMGAgjVQhB/YZHJGls70IPctugCaMXAnMowMcULqVUoy
jTofjeUga1tn+7NJRmUJ7cFr4UqI/5fBwHGVBLp+ggyAY0AEmGPg+3JllzKv5pivz2p233C0fNm9
+nF0dFcK5jgOgJNGgDyQtyv/H6RMPHzobkd+smhsLqzX5m1mjDc5Atv9hrzZD8nDige8E5Jfwqbp
y304hvCOxGO63o808uqYtR7GdGVLcUh7DtJGUqYSAUG0U7R48cpLl+DGNOFdB9BMCl9drMohDNt+
H5cB0yBzF72nHcy+khcawb34IwwsNNAbmQQHUH/plwUC/LA3lYcLFBEkEBO9LTvkSNYuqefoNYaq
KbrBN/47vD1KCBiv8J2U6Jz11KUTx5HpwnBfvqTA8LkLwWc9f1FsbJt8Zpn5Y+okAC8VIzWNWSkz
nPY3QxY2DmOI608BKQSYAh22VxWMHksSM4NFNjPWwWkJtdIygSjIn4Hix4YFYNqm3ht5A+eLbUlu
Mfx/m18aErGQ4GztPr9CIew4CsmOR5g4Sd7VYiu/e3QIZHs5nlrAfjIa2+8XRW+8wFmitkkklen/
WV/0ait8mbUU3UQMpx16jemM6AqrPYUa9zJZjKWt9lnIaBj71/DEy4T1fwVsxDB+Aa3tiUGobMPH
FhTkP+zEcIrJzQzE7OiUE66CHMwe8XDVyZb+s3GTUHjisqnciK5PT5KdPKm/P8tNTZ66ZqzJlp2w
nYZJpMGn0OtXh0kAtNTWNWNRKijyyiOmREyDKl8Xed1LFTGFFlqXQXFbIsw4uvzuHbywfZiZvKRe
24tpbqwbeBT+9Xkpy+wrqAChoqm50Q/KSsD7oL0i8rnV8M3EnmZuEo9T5qjaZHycYtf8xBaYpJJO
+ZyscI9vzlnfcngc+qfgyXyAbMVYA5rj+bTPqtbVzMfX61Lrf//10RWSVImhqiJXOJ5xS73waRL6
6pPZ35G3dwMttN1rdhp7tfjSukwxL7QRHSlvOdqr8/iGK+d+YL3KsdtzOB0TCRYRLZw2AqmpFJYI
GUh/HeSWzb1jUnNh90zLCxtZ/XVVIuZMwkdLSMjvAwDyAfyB+VfhHwrR0va9U4kPH1rRzWycJE4L
jbW+ROMMaB+tdWggCS1ttiAE3lrdnj3Lr1V6qfEAq7qbjRM3tKQBnmuia5ecQjfMXLLexbY77VBr
FdrmMgxvqVcCzw57+uNI3rdvfONl4HOd/UkrcrCfT7iQb6OTJpqgu2esVY1gugzMPloGrL3J2jV1
LHquRVOB0EdW2ey0eWRc5SdV1MT//HGGLydSMFuRNPyA1a9zmJxMBoZrOCq5/e8i7w2KltSjd6R3
Ya5HUSNS39xxIqW3OwD9kzG7J6cj/eXifPq9mcdlLvYtomnbodpk7cPxgzYBkef69G9J8Npgch62
m0FofmwNng229O72zUvRqSvL1ZWvHp1031IdxJKzQI67bdtKtet8GYPvIAaNIztMIUstD+/NBXur
uHPbSu119RibqV5kf5IL/M+ccs0N2WMHp/jjN0LinBWjGM7Fq6WdYqTJ1M8u4NvzP/9a/EmSKFDg
1vw+z0i014KULag0G/AspycT4SePEyRIshbmmoh9/usNCvBAa4y6HjUK/bXhYVvs/P0FLtp29AmB
XM1KLyokWf0KeXiYp3WTo5FyNhjhkmW9ZquTFpWBUt1fKZoKCksnKADdQwHlu4SZhyXdB/mJbXSk
NylpgmajUBu7lECabccugNx1hoxuphLadb68RAAmyOQXfBxDJHgygbFm/7sHVO2AU9irzteF3+Eh
lWsvVyuBMhuHhZ1cCch+sV1rQRpvhzCI+Sn1IGldZWUcl2if+/O4sVs57Ne9FFC51n1rS/JhOw/A
oD6Siwkz5l88DU+JW8Ich7D1MWoylbwmlSxIG+wTZ8EqqeOPrUyBcP8/pAB3IcOAgRAH/Y5wuyXA
BSUqjXN4npfgnJqBdQN0ITBamQ0lkQ6QQxKQyQj3I0hPTY0ikCQvA5auaB0uesJRZt6y22/6/IHB
pP+AzOblt0BFrBpN0acWnbCW3ylQ7f17xWy3Ffyl7z/kcArvgZ07d3rYWJAZNjiA/JNPWEOI7uzs
AcmAd9ulLGxth7Ul2c8ethwRH+84XwLpCpnw/0nAeridiO3XdA38x++Se/paLx8g/UDkvjeqceEd
BlJlzincu47QqnWo0DnytK9lc608ojdgPZ16KMEv+qNhlp1+GMj1CTJqewXBOEDh0PYEUQpeTcbe
6J5anJiItSMmhywYZOiNC5aOWJyBMIF+oTfte8KH7lr4ZUXYUUpzxc1uYutsg8Io5GeYQuq/8DMI
U6kyYKlL2l4yLp6XH49C858b1cJAo/qmtG6By6RO2SY8tkWt7Uwv0qDs9BgYbkh3hn3AEXqQjsEq
SeclxOhPHx9v0S2/ULJKTVPhgvRU2Kqr7oS/2EZYDZA8frKsFz7GoJlEe3F4DAijlGr7HXzX5Aw9
zunVgGcvQFqyO2YujMDc30hNQzCG+hy4MgEr3H0TAOosJ+z7l8PuyF7vYXFYEIX2it5rcuQ+SI9q
gM1vD6yo6wyAaF907jMyqJ3JVd093d21w2ApCyVCql28img0BX4WsGNuS1PgOO+MCDp2P14yX7BR
Uo4XyPsKkvdggHtdDdk0o/9wsfs2tlNWYcXRRkd8wrhAr7HOYzbpVQmQbXkvfKLgr5MFJDiqLYTt
G213eyqpJqFqtkasHKGV3uQftn8spvzmxSpi4wpgq8uevK5gAWVt0ZHT9tbnxZbT1iZf80Knvu8P
+FMAfUmhu4ExV4EM1+0omNG6x03lCDPTOr8ihWqQu5GXGLR3cLsFmhlb3XZA+nNWwQwNgeR1pPJr
z3iOj0NKoOrNsWV1HAvCNFLz3ni+ROYWDFkeuCFuJ/QA0apBtI1JZUK8+cPMsI5hehnLe9TcWHX0
XCe72FY4bHsZeFXT5P+/YudA/koO+HK5GXmFEbpM7Z5SJo2xD1YexFaXSksQp9IfMuQWcjVn8Cwn
8yL3RWSszt9/wjKGCB+rHxYxaYqthkJkFt2l8B1XmSBvySW4qFqMlzaEr5avuWzofEttJPWHutwk
E1dGFKQiXJ1koct9rDQvUKnWdPxRWi8BsoPJ05BESFvUO3lOFNy40+uszDjev/7Xlb+36ArvsXBS
GkxNBbOmokqdcCJd7fnuKeQBP0gJMdxuJ7Lt+Jijr2E1CXEgn8SJ0gxnyMiJ9DEt/BHa2rjNVMlX
U0XhYpF6wlXNzztrt2YK8eRU/sBo3dpZz3UIq2wX0RUdA3eZEF4sVSuT3PvZfyX7LaNkk0V/ABTh
HICxqXtpCQ2iyYzRtPDaaXN0uWc4Qp2IZThTIwKYOWc7HbSUncxQCWhrD3gnGcIZLl4F4gTrDwvw
jDl/32QbpHbHzGSbRIuek0ROzHlHgyu5+6GfpJ1+ZkYTanRpoDM9mjPuP57FGzCBmI6B1JJnT9pE
Uij/MOi9iuQ+YyJ/kKk7j+DbsTxaTf/PcGTtB0CWE4dbhOaXHhxqO0OYXEX2OPDsAaITrEQx8g4h
oDlo4KSdF2bMwSbjypHBaC/4VsV2krNuMvBcjmbOldmd58PwrgybiE+rsu37t4qRXAmPSC6Ebqvl
w4l6Y7TArWV6LoI/P/ecgYlgOvpbpMdpoMWg0EvcVviHJPQ0TcUkkBQsLqc5xQanR2IBrimI/ViC
70zKvLUjyQhhvrHoMZDKd9Culoxn7ht4tdtgl/NHaDObdenFg1iWDgZe3EPamYBqJJQGQ7pPPs/9
bBKUW12wByajq5ViI0/bEFYNAacDqxAJ3w39W0BAwxNirDOazNbxFB2o0ZN3VLEV4uGA+U1mjN1e
DXXztp+TXqEKnw+v+iQSfvvIh9qSHMf0kTDQwzyhvwnLyFZ3rQZHoh2aUZyTvxqxpwTdH3kIsArk
HFpb7s0ddYGpAZKybWqpzljwE/TWIJdTotBo4fIYcqX/eM6ioG3tSrkOpfo7TyN4cu6mCSPCZqwx
PLe9YSq8AkYdH50Rzcxf9/T+3gAYP4z+H0wgzVyKYimIRnaH7HIUBsvMujLNnsLlXotaJPW9fdyZ
t35LF8XLj0OYRqTrIvwYzSIpFQ5DFFG+9jzwjvYR2EYUWAk6jEgWdA4vi/bS/JESdv8eyfHSkfvG
7PRlYXSq+3S0YqjHMreFZuPUDLgU5M3s00ewip9fyr6jLyp31VvtfsUz+gn64CczrISz+RHMde9K
+EW/OD4GULEKwiGhPwb+iN6TJcytkAxIuscjxgxi4UFN7uowQdU+wkSjMHiNr6gfuUZi8NZHGjch
iFssc4+hZPC2VTAvnVKN7Kihw0XEs0MxAOxGbAq2YDmKR+tgMYHeA2RnKee+WCHezfHngYLnEVqC
AndbfMGxc304rjAj046kpjmE2/MGg1Kh6Qh7WJ8yQVKwozTuth8TvAQ+PM+pmiNw9LgVdLuwWu3d
pJLN9iL4R7HNwwH1YxcGjNFjpUjqm7o5i0i8xj88iNjyBU6NCz1DMQlsKF4z6OI5ktLviCZbnYI2
lD4IDPJgZIgE+W6gmnUiK6gNEMFQ8pL22yPvDsJeUifA2zy74i7hSxXY4HhqFiSQpBGJv3JpZyEu
YGIQWrbqmBG7F9HFQxWw0FIsS3vpWdR4HrTnOmnzBHvPHCnK/DEndB6YdtuS7DwMHGse2z9dSQVP
4JV7bROsdQARUxbnpWMnB7lZTX4w8Vgc6h0biuOS98jXwxSqHPWspqXrODDFdcnP1bnVpaP1EOHt
OvK+fVg7cHFQFrYZnsOJTXcwCkkmepZ69MTlBgzs8KKSY+KcWW3QvCj6jc0qCgSojevoqsjcysIk
gHZloYgJ8VNiK23vdzfIQrlj8BAnpn2ESOz3INLQcCgQTdJFMXvWJHEAww0lf3ua48Pp+OWrwU2c
E4Hyrhiqu1lJU389w6ueS13X9uCy4lRYYFWzbD5FakfRVf3UCJhVHg+d4Vgcg3ZHbGosewesMwr1
HrdwYv9GD3lw5uoFpd8YNv2R2MdfvBpSmVVkzF3zMsZjrqoa0tl5CXSpsubRcYHBAeNyn0Uhjh4M
3vTtbsT6pSIj1nA779fTLebekk9IzCAnhcYDvEZrNbGS9gxHEgGGgyPaHwRnyOGH5y0EIkO1ZDz7
IMiuLcK2/kw3W3F1XSg/bB/YHXzx5U11RO3SdKSHMWxhm3aEZujwxmHScJmi2ZBeNbEtbGNdDk+M
SMWr45NxOUkW9ZuRtk6XwShKggE+PiN7fMBakkAFf7vmqvGUp2X4WJy+3nB0bBlNVi5vdLOb9AAP
kNAx53aqbq6/UqJncC3coK0UAXGsPC2PnklkuMuFOJ77zbxT/4APReEWgtSSXW/yWHT6Ca9H5P2w
gpnr8YOEGLRum612PxUlxYIfsrVL8EpLZf01qPJ36sofYAO+tIHsoFbFMW315UIrKXe041NfDWMb
maUjmWsCrEEvKjcl1XE0tV3+ssXCitmhkMXpTdyQk8AjCnA/hskeYPPtU4dsp0bNAg4hn4Sq0kHD
EthHH5WvQ+5gR4mBonu16rxs62qd5ePFZ/PWZhTUE5+JNRsc/+VZH4wVrKTKUD8P9490rqbgZnYW
CTYsR5lLaYaenuePj+fvmESvXK9L382W6KeZzcEBj0p5Y6OLAeZAz8zVePmcMz3SlIQiBPQ3gwI2
Rx3qjHhfsKHyykRTKI28uEMHKgd59Yy8++9Le1IpAnci+SIa9fgHAepc9BfsD2SPtIbsdwjDbXUI
c41TSTU8DX3zTgmhfSq24zfSeYbFjtUxyAB8l+09tntsOwv4SH/yBl9tJpXbJkxLIMjgOgVAMhpO
KYZHvZVKtfyIDxGRMN4pj4NqOWXrh6nAoidSDFNmIOpFV8tcF4x4xaVXyDU8giFMzkJZlLvK1TWM
jFir5PGtelkRLRv05QyhDK/kWY880O5n5k5uuAzIgbviOOyu7BrEClxzgziQoXYeDnBmvvCMmNjd
o1E5nhf3+w6ZghaezFdqi6Rd1lc9BsWKyG/t7RpFkik4COGWDIyklKALWBjOe9/mNfSs7mF09gSz
IWHFeWPaEhRIowr6ooiJ6PfW36vVdsBop3MKg7tzXiKn23CKYhkvU1gJ/osYl/7qc5bMZPP3nym6
0ZdzC2n3H2xJOSFFLvgD5Qfj4TC2Wc5LnGscXoOcF8FglBksJ+HAU5lbbiluuoXGbriydOmomB4p
EhHw1kyST4yCHlF4fBrgaSZt8/uHMJQnYhaob3+nBUaIjVe5mpKrjdkEQsRxGFVUdjBsh3pclULU
1UmvHKgJbvfe8X4bUfeXUJvgtd/VAkGfe0epmIRmjImeXCBP4EtjOXoZwVa4CKyPWE45x1TQ6qAH
iHl8dRBZw5iGHfSocrx6BvlLWmcCgclKaeurUlaELcXADTpcGuNP449zMgIu+gfcpndOsQAnYeNw
KZpu8woErM4i2QulDQ7/GOuHxg+20w3LCKG6J2IwyqG94q3lpHMIRMyZauqcIi2Wxu2tCnnB9i7F
ehgfeA0qFxa9hSGnPscnpoLmovd9nXZy3H9YTCDdIzFxAszZZWdIzP9NUkVEvapMwlmwq6vgWt1r
aYZdGScyVSaOYdq3yIakTgXCY/++FbiXu+A+g2GuwWzihY0CrtQ56Xbg9lg9JjRrhjR1cKqa2ZnU
XHuHdmrsOqC01ijw44abwgt9TFksydV7lUPCqSihnsy5m/5bwfHlziUT+bYJsQk7Ed4NWalUlVol
y0J0S2PGG4l/cvxXd6RaEkDEPX3bzuvV4ADbPgI82LIdK4kXLGpmk6Lea9j3fZgoWZdil27vYhve
WiAUhCBZc3HZp/ndq8WaFrtNpWP02mgjDkUC9ppIwrKOLn0eBijGTvosHp50Kv61XHrcIjkBqf9L
twLy6F3zGv9Ji6TobHzrktQcKkqFRSTfOJQn87TqxHuve3iyt76W4BgXRiHtvHifyI8R10PhwXIS
RqgaLrYvhtR13Wsd0ERhYXuoUU2nHl4ebdY6fxtJ5ln1WDzc01JqyYTnOtGSj4gTK/OtJKCdOjni
Ap5J+rbHcZnd1jGqybHoAaikaGKhqRrltLk7Y1xcchlvTJT7iXmeduhfq6UaEuF85UOmVLBHwsB1
/8dCiMYxToAvvAQ4+0Ef4lzc29qmIMwzUleIWOBvJRuyS+UNq+8TlRN2DGcNuNeL0SaFnSdSy2xR
vuP9BxNtjb+24vBfOqsLjhZefOd2jsHItlqjKa9QlbstQH/vHALi2+hQY99Nf+/zzfrYsMg1xpHU
60U2LnnJzrOvvTSKzIU+5CtCaqQABPkkCfxXMGbCAZWO12uzl8L70qhmTH4i+paQKS7cpPglbyy6
0WW3legke0tDQv1jauSjUvXS/fYs8IB2Valb2Z6vAIMevnEzNglcbzsKaB0rNLz0jMty9A7Ykwhl
sCsVsKDl8lMG4WK+qq1rodcPfqQLesZImPEUnp9TL0Kofp1N9U80vfoQX551ggdf1E/ey+Hb0Nmg
b65Mlv3kWrn9+7S0x/yUv9HeowrQIakhtiTfEVJ5FDUKfpqrmVmG2lwii6LZgAeiF7stufg0qlxX
rBcfmCi5wM1qv2R72ThQvoo8IQvoC5XzvrYe4vkN9K+QZCrNVASS5i1cwRSfHmxzciPjaLQeBB3g
zNwuYxKaLzvRcijsRCM3cFz1tNRFMeB53grcYKdzFEtXNsXdNYTpSBhrK/sznHpIxyEKP1892/Re
Iu4Ytgx6tyrE0eGuTEcQbwh7zGlnc3nhIgDBHuaAA7Xx4sv+Zd3CkJS+w5pSkWGBkhm2ON83mKkI
ln5GQUGvHPSwskN66vKVwIxq/KOauk2OsNKKcAqfMxzo+9F3/GjRsgWm7DzY+ae+KGQMoWG258Pl
UvvvdRabsJIPvnA6FWoqNx6CSEEPqni2uHe+QEPAkZjokPn/cSnaqS/bfgKf5acy+UIANkMDxnqq
ybFObDIkUkDGvIjuBcr3zctfW9fRlzN8xK6rHFGC+cFj4p0UwXtNX1eAKb7pL5NGRsQZE0TPhwHC
QP1xGM2bmCVaup2qS6ouAZzclGFsqLgoGlh2t+hvaWSFdX66+UPPpFYEvi7cXnuetXysU1OcDIY+
y7oDXa2fL0Vos7m42e4d6wkOUYv0X/ZyWFXEuBRp2bfp9B4+RuVUGcDGV/DYcYlqbFKMYkg9H2Ps
+o0JAg3n0ION63slHFppzDehCk/ri3xWr6OXvRxDno6HykqIY+14NfsfGZ14d4D22Nmaru+Mm7C0
fTNTmTvvMsf4uXLsU522zZIN/YaMXpIcXfq1/p/CgXZyaxMt8TFsIDXnrJw7ip1Btdb2YP9cgkaj
lREkZt9U9poJ5b8pfrWdWJkkQq3dvLZxZ1cl6kNVsBd5FG07zX2kBKjJlWGOYVxjsReC/IjvamDs
lCF7Kg2MurUdK5QVFiY7i3k/a7KcizL3vwn0T8jVmaEKvoHHgpUWyPfjjB/xWxWeznOuB6G9HXzb
1KDU0P7BSsXwNV6QJ9PofFkTCk8COsVcuhe+8st/IqlOIkeArsXOE4m/t/qcb+km7rGuwlKvY6wu
bZqXzI8qd93gV8kGVaABqaGGpkE+E+6Z5GtFfaizCQgr3SEbpMFUfoixgt+n46WHyDRuQ23GVGRy
d3OY1/b/UW6TIPPzsKoy/unPkeEpYe1V2wwU6zdllOHgedsVw61DaPsPEsRns9MJXtx779Ugzfsy
2uCoufOyHTtinuNepXebUAxQ8dy15HZuSWIbHHnppyjRkQl98NHopCc+/yaJ+SSprXfuK90gYF9x
zO3VbGaUmZAlKVfoq8QDPzLK9coGgo68SY0pw20QoiJ6xjYmMkSE2qKgmjAHS0NgX0LQPDvl5vyN
7UTBqsYaaHlknJNl47ckYhwLymOMCBzXaKHNPzwowQ90FBDqIXFta3xh8OlKMTLpyQDqsEgcuEu8
Ix+ba98RAd5FsEX2haUxSrz4/JvCgPV0KrSJp8Fh+Qt8WJUtYQX7VMONR2OgzdT7g8E3cgr6pM2H
MsZhSR61anzQ0pqZiDjaRbVt2NNLQHKxMuqB/fvEyee2YJm0m9ufQrCqKYl0ne+X5wuzoZBm07Du
RR7GXvaW+I9ebzCBBOSQc3syvlnHp8Y/UQkUzTM/TXo9zV1c0hEeCWzn2/Bef41ENGvdLZJEwPCA
WppiM/IekWSFjxXUQ8r3vI+HN4zwqP4savOvy7DidOeMQqSlaAbRSvC8eVSYxDv+Krndpv7iUQVA
uodMmLwwQN14u95jlEzrQZu7qNTHbDdtHPFrzKnehLhQwH8IMjK+SwJb8NmmN8YCt4g6dnWbZL76
cFpEIfyzqcr1kXgAUMKoCg8/D28hGUAsk9knuLSjA7Y4vfD/0NTrmUKOWP9xmy3af8DojaPMsm+r
mfqNUws41rueEfFXwnl62eepTUgPxXhPpU+bNK2Ocdl8XpfTtLOaQS0pxbRtAF5jJrxZxLwO/rEC
XXn1xDDNCUwXFX2lYuMEWrHZm4quoPQvWn0JmwlByGqYRgZHe16oMdHUWyXPTpcdv9+619DngoNd
hgCqRqajeg/2FFUCVhfh2izb0wBPzHNCi0Gz3Eq3X5KATV/AolZOhMh4p+T94xuAzYMrJPMmtSL5
1ak5pdth7+t7O2HVqKgX8l7snw+skUNz7ZKhKkRxWSakkj0uUkbiItEf8y2kAAdb/JiX4FzDufzb
ZQy5BJzzfXMfBA6Jv0eAClCysFkO64JaG/F9Z0KW3lmazCMt0V60TS1B7qaYip9pKgpPWvEWCHHr
e+heRf+fW0TxTLEG0WBmMYRK6QSs6W5G/N7MXdFm0JzsncYmnZKGyw61m/bWJaM1fTXdbnU3rBBk
4DJb7NCy5LT9mQSv4MPFlWykxlzR+GLbMllkgDQmSwuQNuXqASpVJrER3bAMU9YuA5lA6zJVRkvm
E3xeFHhxJdE/t8V89DtAJxvLkaMl2EuV2SfGwWryqlbdiix8ezt0oYx5oz0v74Z4YVt3qTSFmaXW
vfR1qQVAdXr+M2pqhQxlwbb4P0ALteq5LPHnq/S67nhTErTMbObSSMCjmEFaikOWN2PhndSCNuri
cedRA/JImlE29qDI5UWGE8yInZ4Ip99EpSJxS/0lKEaLchQbWfamhtMWqLFF1tITlvDAYeiyRwlO
sP5R6gUePbYTe+KzXl51LT62orsGK3HgFBnsLHC1ABLPAAfNyVsOUD0rWLzayrmbEs/LlhoRtne9
MR1HcRpNmO43wNFj1rysxDOocpWq7/g5jNY0QwmWa1cVOam2k3M+SpXizC2VSuY+H7Eu6wgj1pKe
EwPj5LTkCBZMrW2XQiFJThDSPKEw5jxDS/WjiPNpFOscq6G7ehzvdau1htq+/r/lZRIMyNa2ntJo
L4hjBicvjhLZFXyuebSK11U/4akwze2XGeJeBMIB1V+dPKyEkoXbACL+GeJbY/a850zPWj3h0PVS
onf0DioEFv0ZewotQnls8bMIp3+vlbhLmvF88NGB27qZ5YhYsGRwHTa21cDjQ/wgF/TfCfW2XMh6
fcyBM4jOeqxD6rJ7lDMPvXg8B59sAgID9FtB1ObRcEtZL2thvQBEkhYeFS3CGBa7S+MxtmamotuH
B6+tLSZNN0A95XfZGUoUPeip1meZT0Qclg9TNlFEHxcYpTGEjLVcK9gdt+FhOeMI/o7w9XmcH590
2xgbEaQanYvJUB1k4yajjrubNI10SjVrpkuT0KOf6wAIAEKjoS5dGt/y1w84bR7EibET68NnhF1F
BHlqjwlCd7+PTBB2jAWyFy54V6S7KZ2afZCgmUxcn1ax07QQZaMPHHxKSrs727VvnhXYmV08xllE
nL6YaCQQdXDw9bkLTIsd86F5XV+Inqk48o/sZT7KinsbjG4WrcwjmROU/h/u4Ktn45nLcY//g5wZ
uBkQrQtUZIL7VdjySztM/5OIvmzgACLuQ2OwcPtpZIppm30OBGMUEBGNO+/oRn3xxyssCnNfO6om
SLmT+e7OIav8Yt1H84jDbZl9z+/qB2kAIbkOoDg/JpdaeygWzERIKPjGsq8g5fueq74PLpdQj/Uh
v1K9CtjHDQQQxfv0wU40puAy6F70yvYW2TL9axIg8aThcj3K6uKJghh6UIEkssEVyAVkGZ5NtuN9
RSFnc9alxY+KsnQDeVfXgdhwunfzGMas9snUdlpkMX14LJNkguw/dlLtF7ie6jyc5hshJS3k2J6m
5TRWtnDsLpSykp3+U0mv4VqZ3xx7S8lrhAd8xIas8CahsksSx6xt50S+IKVpe/EogHFUDBVrJkQ/
pBtD3W6/5Rs/m1jsAjom6Jtn8rAufgiJwK8B0FQfzpNRfvN+aj2E6Op68dQbAVBJFHFAFk4bjz9L
ikY0AbzTgxNLMZpsn7ahYkE1CEX9F4+r3uGF3pbyDvRatPqXixmiEXDuvSO6HmO0U5JZTws3zVle
L2JSBlo67sySpicfR51GF4UcoUcP0G0aiVYNm1wD4nyoVWaXkvsQn2IWpUjpxqimG27dDDhZPlUb
gLHDK+LZIORnZa/wp33qAUfiY75DmdHSA9ZW0oXWb76WPYtSb1+5ARUfnFnii+s/zWXbSuCd4Hlc
i74sIvFPJMONuMeObtidvFI1LjpvztashWyNQGj1v4lNBJ00LaLPAGtnMzhGOUTRSIW75QaF/iQo
Ps5Ky8g6ZY+7yiPecEx9bvpvd9PCp7kb5puSwJ+gIm0ePLs3LkGyxK7LgrdRW92EmSxn5x8jNjhs
ylHqtpogt+iLM4a2zHczpCGAEp/+wv1zFeAuP2i8f6ua24kiYUTSQ2T5NKWINsGP6zBPoQe9A+sz
qhNedWsNhLMDCx0RUE6UUXfvNmNKsaCLhLfxONFj3eHKcdZavh0intKF4Pfes0m0jNqppB0YTqEx
adcbJxZITBXkvpF6uoyIoI7txs68ASNB1A01OHC4hFGwVpnZoK2vHTDJctUlBWuxPttiF9p29bs3
DgT1cNrXqVYm/FqvwI/1WDqKfYc/tJjZnkdc19tbHqstxqoU1BPjbFyXpS/BYLDkPehI4rU0OiVb
KUKk90dUaObWPy5eQuBBp3pe+32CjecvpmoS0JXKR8++fJMGI28lddKyGBlzA7R5T4WgUe08PMeT
QGv/RHrFyChFl1HxreOFVTL6RF0UoGRTzCNe3v8qMBS9E8viddhtwxyE4p608jLFtjDk5FlEhRDU
28ORW9tUhg9XdQSzbslA/OQhbyFOPgkpsh2Eir9mZHke78KzbtZrePGEGrQOTekHAs0ilPQmgmWR
xK2v8sOryD9VVphIGg04SIMXCqtJd5WYFbPIluKCfK05S/t3pwL2GmcFona0cjUvB37Nv2MxzAkN
6IlMWp2Y2u+qlatmixLk/a3dex1G3nKLBM139sER6vtakQZdaVgV6dsydP+p0QzSdg/qDl3TvNl0
W8UIT9qJB46c0mLWAf4BqTWdTvcIJd5bgX4f63XtnZ1s50nTA6CN+HsLYmgk1F/CmVOuLWlM4f1P
LWvZ7ZvjvKZiamrf+eNEKDTFy8mWC41V3o3Dm/c7djXRkEJEFSQkso+vWNn8/M4D216Y4594dF2H
VTl0UUIUi/v02K21vDkGE0SuxQqrH0Q8uG44Sftf034mBmiJ90enLEqNwGXaS7OOVvDFW2j4dp4i
I7AhYG4mN/4ODl+9KbINKe5v2SpUmd2WeN1IjkTjd3J7L6XUyqHs3Td8xw39WSQbQIjZaLh0G+dN
q0DaddpCHypcnwFbAb7uTj9uJb4gUwfLLKVfKOHn/xYSQFocSREW3Q+BWdTLDeIoFUda69NPDKSc
+IoVYVAd5B0W6qwCQGit5Zxjq/dgNZq3z2cQurIwHpk/EugGEz9ou518fclxleNLpFd8ZHlvoRuj
XfIoIjiw3hBsT26K/gcx4wlKYSGI/JASgH4h4f6kwzDOOjMU9fehDSsTB7BhNtWMK8y6UbNP493T
FWButZgHGBL/Xs38wYJsx2cCTR8ns7sLjzIl44m1Re0Dr0U8jbJhlkhxav1aJKvZRtXkLIaZin9J
KmJ7gb9MTjbIilH4KJznZc6yWF5hNPwuYUYUtEQbP6fLnridXoNbMQw5cYAIs754IkuJmcssI/eG
+2igh8nwFPCWT9sirztjAOpAk0CTpgZ0/GR2WqFT+Eu3Amk6qJEpCZeAHdAFNcixBJwS5ADeoCn4
H4/avttu/g0fXHkg1u85+JATdQdzRRQWKRxv4ZY2Vc5D5CR8NNk87vit2cLS9YV/E74uu81CbSi3
r3c6CJ3xqeNc39M7g7aXK559dVLIiGOSNpCzasB8GmgNWwG7MbJL2ru+TyD5/+GYtv48gGbUDM+G
TcH3YHGCzpTqft7Gg88JkoqMTHYzYcxguHQKue4RiHIkTvGCCfsTMcVGVHqzG9sjSTYqfYNBU5hO
BhXdLnjWGRGj0gbkKdMJecrq3GKF5zhQ3VspoyH5ik8Fciyk/gXPe7bVy/eIUa20eLuRofZIe6Bm
6usTizAftQlEsS0JkCmEon+tCQ8mvt6w0UUD9iImDe86Uwwvugl6sTuegoXVBolP+qfGGE2KPL5f
/+5iAohXAM4lc6afp20F3n0+IL+CmfOPWRKyJhJl4pZlC2X/wUV2DZggpJ2khm0BkHiLQR8Ce7Cd
5AyRPw+YVufKUvUVSFlmF+6Ur+DbpDNi+G1KSMGEIxhlo5aGrVdI9xHJQKsONAjYKfeM8pYWe351
l0p7QrDZLlqttTXJQ3x0acDpNA12ZFQI/ya6n+t4GPafs2N5YL58tEyDeR1pnku1Dx/v84lPqM8B
b4htMubilWEMrx4OubW0qJfqLpGI3OJKXjqLa6qM6uIm7wf4+IBzRiF8rII1vLqPYL4km3mt7v50
ps9zwSfwW95yWrPCrWsil09xQJn3PHN0MUTocINCLmhxYtCX4G7KMoM4JlpLAvLnlSxK8KYX6x7R
Xk/XL98NPKWlstpeYHlM1V9x6+Rg439abD3//chSU+jYZeLPpTkjI4IFtFl8ef3nCjN395WSi1Cg
QKxY4Peg5nTl+kogycX8MieA9jkUSqihXJrFoZlOL6a8MmbBQjC5vICVmcOPIQ0Dlk3rM7TsU/8Q
R/nLSQunp3NRqcbB74IfbzpmVdnA0Ws5mudZY41gMnZESjXPYHibHvkBA0ycgdHPWwvFFjgGtB/F
oyQMV4EFaTgXFYtTFLVTA6mLGtN6J40i6WQhSzd4mfmi1SfYbjhslAuuD4ryyyxtLrDvzk1N5+K7
XX3MMRGHM+0FmEh+NphrzAiCM7Ql9nmuKjGiJWEO46BIe37C2dQk/yM0lIZ59yRlv/lnTAN7K2Jt
tiIOMOdHd6UI19ySPpWC4GfSavfdOgsUM/7FER2s/5G0XKLled/e1BuZBwLZ64qOgf+eQp3gv5SR
EUGN63lOX+celpyceePKPDqTK6EmbS7SkC24Cma5E4E3w1yO35c6WFoSQYtF6H0nfOvktWOmE5yh
RrwGY/61sr4G8xOAgZUnacu6ECdT1FRwtsP+sjf+lZPTrFQNBpFY+AoAxnefxnj7xZJiSTQMnB5D
J8zif+ERqyb+pEY5WObFppcWbN4gIX1Y46ZXgNHRHKbuLhtHzJg0cewU6fBOCjtq30OoaDhh+nbw
jcRrhVQebLWMch+wnJppRBgTquv0S5bks+HGuX3vkdMlSrrGn+vzOxRcT6Z1/qIE10RUKfuCzFLB
VxCkSG/6rSjWXb4Nnaz4mnylRV1zOYsBNjlwu1P6dIwtRaAVytTHrBb3dbjG04W5d6NEmfcx0/e+
8nikMmyIFPdZ3l5HAqEU2CPG2hpnpWHaZe+DONmiDD9LPVni/m4iB+RSHkGU3/vTD9G6/lpsV1ik
UnEyVQ9GtH4sdKO+lENL29AGANmzV2jvh7LypVYlG3ng/0DT0FNRX9aqDdsuglRCV2nDdZP2DHkQ
tiVODBYTSnytRfQrNubCK/D9WKwOSaIA/+6zGfzZG6Dng65yPxxav1kJG83fRTdf9ytls77W218g
wJ1DTD3OMACmb4dGpqVS2x0jaab5LYMHkdH6cAhUF1slqT2q6UcF/ZYhna1J9YwPDjbhHB6NvoyJ
O1ZS0BX6dmemM0feX0CIq3DKfFY3QS0g8h/04n5ZPJMALROk6x7/5RCEgLYCEwk4lusvenmVmK6+
hR2h7OAhot1pJbhP+yDnq9wkMx4nIjOQAn764t6MWKT802+SF4KIBe0VbowmpJYeR2RqrHHFu1KT
/F0fqgWQo2p23RuYt7v1qdeMdTjZ+qzLHS5DrPExh3iJ/gEw64i72R9SlMw1xCSRP+yj+k7GNgCz
SAUnjUSsTcuuLrVYBG0gmA2jBlOv365Xx0t3lSPXrOs3PBcacfn/gYEXgrXwgFq3X0OqhPMeBowU
7h+Fny0Ir4K7yLLsnmPYZouRYVZVEm7BGAue/zjhv0r9xeLVOnw2nzx5TQ41rxN1bwLRBvnq4xIC
LRAjLxk8IylEW7bKhWMFy8tNOWe3VTWDM/QMx/F/nmdqxt3GmSiN8CjREsYVq/Fs6AYbBApgKbsa
+JF2L5rPkNZmCO3TiyZbb6l8ooJbP5hlCtr6FNZtnzg0CM0QIi2g/qiVbAcuWRCkL9ypbH/sArRl
NiNRnKFnmt5VTWeKUdsMx3aG0vVg/NOrstwuWitmXe3XYgCG5zTplwymG3sOSmtoHJUqG3zjLWnk
K0WceQberG44QfNmEgLjA+rlZvn0i7cbPAdOGX+TbTV3EWrP2DdORFe4B+Et2O9JNaBGvefKLASc
+YkoCMhHaXKuYNvcl/S1ZvgkCFwsBLDBCzmQvvIhL0p+4YiRAtVvTFSIRwp/HU58D9T8aXMFENWz
qHtF8j2elx3R9m6NaX6KuvxOkKZfYPw92hJssKBEYw7uS7+KdlZSBmQTW3oMv5b7YZW7tC1xIEB2
jkHFU9HGuHbtsBbY0xzeCfPmqsjWp78uzI/9YRhq3W3bLJ8+sALtw8bKlo3uSqCi1jWPXwtMmuER
sc3b9YRn2QL5oE2QtCJn+TH3V7dmsOTm3THv+XCVkZKkZfVF8oigJkPqARNptWlJJNMG09O1Y/HE
e999Ys5WF9NUkftwK0bjyKmGHuhr5P/i0uz5j7Miqk9qF88rFh4mF5+CIUgfgHhYlZxWM5+eh9EM
KK+uU/Bh/gYpL7p9duMbd5oeJ/hEvytALL9e9RJ56Yc4oi5m2j6ylRLGpxXOdKsFC4VtLvCfR57b
1rJz9Bhch2bUZuxLJe2K+WC73QgQDSVznwP+szHfzPf914S7Ou0W9gqEKDKtDE842Zj5XLkTU8SC
Q3QdHcPU24mEnBve487vHCqNuyIvgnc+3nFU7NYVTxxL9SB+HE2cj5D5UM42ht8ddMiliq/1uy9Q
RmpSVpgXdXShlSv1bPyDU/E1yq8cDQUYhutXYM13ZvWokpNddjU+mpIy3aM33W53ogDJ4LMkyGFJ
J8H5ScVNTYrfHvhc+Kbl81SVikSFKwEE6ATwuabw7wl0UeOKm0BiibOZlBGebG1fJyBd6wDkb0SY
t+Ia1YHkubwpnYwj91YLyC3LAk2cfCZb48oRgCyEVF3j48BgWUMRfqZ5xyKTIeGGkCvi/CiwfQ/W
uh8Q02LlHAq1xVptIJZcBiDwGl/QclaWca8O2QBuBHiw1cWjlyD6FZukUMQk7UNV6NsFjxRC7JUz
VEeDSTNfO3agrPkpfielC0nU8PeUZS+pqlhWySwfzzY8q2pIcOw2uYgLl9SHgicjKhOu1NE/JK2y
gZju+PTHg4hwG8VDbXUOczjVsH9gmhkgDLHNhwfMc6MZid84D5Ar01F9z0VXXifAOWmX3ZVD3Tni
GutnuFPMWgNDxsjg0Gz4WaU4p0pPZ1qXx86lhj2DjSkLJzyiUUlj8n+cNpdsTcNFQhCrZpNo5zxb
+tCfgV8WMnl4PP8cg1FR0Sjt6kxf3WNVPwaijZeEMEnRSB5gJQz2IaVMoK5lP4ax68w9fjQuR2EK
DqgCecHTI4faVThVBHARp5Idom5lFzZ6Oe+e2tDXaQ+wBWm9FgAvagHnBr/eZ7pQGb7CcJA2PWQh
tKkMdhLs0AFlnm45fAhW1QgFMSgXKEGQ4SHZfZN9q4oI9JHKE0ywoNojd+FO2zBzI1XkxVcbXKSD
1djkaYKHgbS7svs5xeuWzgZA5veylqf2x1KfLGb2MkzDbRr2Vt/E8NE7KDzfwdm+g0+ECGaO5Wws
JzxoZDrsS536jfHoego0xP7XGkno+jcCTeQ4cnCWsz/tG02YjAgfof3Q2qkF3/D8BL0NgzXsl6pf
wXbBX3uJA8nFQedh7fgpE7J4qP8rF5EZGY+f1qiMPgOwQTQ4F7q4Izig2VmTLCSAwybgpgkUnhIU
ZWYSyOKb1ataKxIn0CyhV8rvw5H+nrLvwnoOmNUitpn/y8X+vk63R0L3iEf5hZbN1KaR6mld+hXW
pgXzNDn8Hh6BRwkr32vjxiyUm16iTh6HO3sG2vViEY7zjT/KWDrX11C5AS1D7QsJAqormX/55mtm
OG4AYyz0uUBZ+eIV3/ADZDcWnHqq2KqtvI3I33cgR4SAq8QOtMqMMBHQrFvsbu9n96nK8nZfg+P+
i5GrOU4LuE/1bbpsA+lcRtwbPKs4H/lxOc4MOBIaF0yITyhZMhNRPfgMqI39+/gduxeept+GOMkp
JEL9JDvxMlpLfuufF504hvBLzspa6yE+p9xyPhhKQFmWp6Bhl1LT0hPM9UX77qu03b9VOR3uamZP
iLD01/v5i2xhbNL3FON0PygYjDpcmT62BLrxHwnJMp3l3CSEAWt/wC+7ywTE/EJRKPqw7fgfN6WJ
/PpAMwcTv3GZdK5vZfV2o86L/h7dWyoQ8WBwiunCrLkXPZ3U625taXky5er/V9z+s+m7NAqJPX/U
9mLmCrnBIiVLUmqPmCSh7WkkrlrkMGv3dLKSoiAiEBM0Ii45b8IVB1hA0hstYRNnIC/ZY1a0WT1/
xxrenqJJYEnHHk54bJa16EAnBeUSdTcMXRh5eh3is/LdnHnbrctxUWGCW2/cePgd0y6r2HTrSnoF
toewhi6pa1Cy8OWUsMt0UqgMlUh0YkxGxBvFhTOErl5AyneP9Y0SyegFRxQlEncq0J4NVF79Gtg1
tHDTlcJIiZ1gGUWN91lAIZaifvP8sayaSMEyJDiQmIoolEUk+CRpy/rVjeD+YsJnrYBB0zokQ+S3
nTbPkmCPOvS3iQUhR6KHG69uo6SviQ/oS7d4JpbKfkMmuGdLL68t42AOv1garTjJqjAZgLGpHLoH
3axSPcJy0N3eDj0mtruWyLUeFAON7OZW2gQGprZF0C/wC2cHU+36yngvbsH6uSwsWDRhBckS+KDR
xJALS+BMqAIzDfUY2ARYGw9kjihUBzhDRKFpgSgU1KS53xx8m779yFcGIYMY8oRXCYyFAZuAgEkg
OY1J9ZrvbwimAZLkOYO3JIST2BWXGNDkAXVNB1rzFXAeDJF2n6JwYaYi5em+G+VLDg9N+aw+JvXT
D5rimoiLbxlILbMoQbRt+bZAYz754zaRhgMgoFFsn0ueSw1fRe6daBSUK0J3mwQAqeya6g/zelxy
WmZYuixAMwR/uxDuWgrlr5Vqn2NsdXMfbNoiYOSyrywXI63SdehXw9rax+3F/imMDNjrO6Q5FzDQ
zopshn+DFSELEVcZYg9km2PXr5yPTv60Cdb9aqH6t/ddO6lLDRYdTp/y4iLn1dmFYihZw92gyBiF
FKNc9UK5XSeXUkXG85zTFKPsNB0i8vLQTKNUTtlI9STXeLHBdc3Y0lVuopJfIGwStQps+RZlXOC1
XMwhcsijEubPQbE1ilykSSioryLK0rVciaNBHzbBkb2q3wAtwi9e2LFnCWddjm5Lg+r51l+mhj02
VWOerGLIwhIYCEibzxhupnLjk2FZxnz+qjOc8xKFcgQ6LZBt+9bLg39pVFn3R9YypDSDh5mViRu7
lQJOsVdvy6jTWys24YknKwIhwPLtGcnzmPcve3rpXdtK2fhFNMpu1yqxca5bY8pQ6yy4iE/lq1EM
N9kqp8dtJ7kXLYBgv3Adwkxnn164n0OBUcD6+taF5m2bmrxEe3hc5weuc1/18ec+JaHbAIjXU3f8
wHwNU6u8UYAEqvMooFHZxq/NfsPEXSN/Dfc9om8SxLQxfyQpMTmV+mPQ+EswS3gUEqV13O+gjlpy
dk1GxsCEkMLucIiBmXMTX63d2jGIxjiQnWgJbQSN45wM3kR0qEJlJ4HRdpjyvtBaAVUJ8HZFHXJ6
tDoYCSfvDy3jW+UB72RRGncSnvm+7zbh6zJu5hzjg2Y8Z1WEAmNC5/Z7VtTgtRMmtHlKEGz2vod1
i/s+VtCsqSM45aO7J43PMCadYjrnllhW1WgDwwTwyuLPlbhf7Ql8jzn4payMV8B0La1hg1KigDMi
xIjrpTKN5Y/Fu7Te9n0T07OOcFh0gFLbJ2N6VWvk3Ov10mX+VTdO0M7Z58B45g933+kuYBEQdY0g
2F8R8BFabwzPMAzB3IyaH1ArhOE6TFc6uZnXBHS6uwCvj+AUKwDKk/b+RPu2B3mFsKrR0tD9+lKn
JZXMh+YWrQCHDj2u//R0xAXXqUzYUxBXDn2s2hxnLuiIUj3CAiKEFnTVeR1NQ+CeJjUb3nyh0MMt
bqaF01lqRStXwq/1/kTbEm+dJPS4jWUxOkmXoZF38iC6BBWeEb/eLoAlTHZLKL+4iJoYMCxGkrc/
P3hQ8QavsfrZLkSPEWQBRiY1NncsNRl/iRpYmJedAm54MjiSMG48wZtd2RtmkctNzmZ6BaUFzuRE
6uxxeIUVgHTJtagBh5YrFgoRABQWUXlEPCl6a54Tt7mPJXkuXcceuyzNlddj/kV7b67Q9oDHXcYF
Uz/PU9xwX4jClcxPe082ljiAXwTG2nSKJx5JuewLtRpKC/I/GNBs9xT0sSTuXIcgOImVg3ZP9GRK
5u90IuL3UpUjo/mKyeZItacWfblTRwZoK2FmOXnxCZEMxX4KiSyYSMGQ1jEsLl7JxYLdy55NdXXh
Y4cZTnPMRA/gfZEsD37Ih4y8XgkggDm4UTlV9GAEk79vwzJZWX7HbTrR9wK//4Q+EL+8sSwWVIOC
viJpHscxyShHh6KlHK7ZCm/XoUdK5Ruo/LTj9ers1i5tvFMr8i1U1KxJBrJ6sqdq7JvCIFR5JlQv
fbuj7WTyjKIENaHtMzWoleZ2wn8VVj0jUWAwnjkg7XRt89RYKvpF2wpvGyGW8c4GqhH7yya29HH1
EQmCv0T1pnlFALFUy0GoDXToUDngLXvsGcUIrjqCDSlVFuv5IefAVD+EypeNkpfPqHc5HGXYZYY9
s8DzxerJf7Zhkvp+W0rAaKB1aK0LL/PIZC5TmurYBs5O0m7LedM492EEB526XNPRufblaZSvqRHX
kY8kdvq9x6dtnzeCagAOrn7GLckHH3dm3z6tYMnHyvGldWUmmJTXrcf8EY/BLK7lHhAF2+o+PFzH
HM/umen340U74HraDj5XfrPbClY8t+J4I5PKG/53ZJrKaAZkv0XQ3svruvdsmZANGotnVnEQ3OXf
Ivt8/BgT1Ut65YXCfRcvWeATwcM8tpjJPYDImsQdouGOfuRFxe4ILhIlZ42ymfIQYt1BGfBaugbx
bS5NAsp5A4PTtk5Pw7q9IN5CauD5z5ehMVJ5fHVkRkHFTf/0vKtcOcvmWgYfH6XQdV7HCTSWXmhp
2/2yuftfYQG6TWJobHH0RzOMRXUhIDGSN0WM/BBTuNJRM9ENNXbU+0Ljv7lvYsio+aNVrkg9aGJ3
WcpbyX+ZocygZ8aSLwM9is0NOcPPJuhnBjfAR+fcdiDqPP7IVPN60xez3aN358Wf8hS49vCcswVt
ajgILI68ZbYB11zxbmuCLKUUoeza7lKa8Fzfdyv2DpH3++t0QYFXrINTamblesNxuHy6Hf1Z0zC3
7pAAXDUL8VQj8yl/4XM70+/ja0J93yyrN4/DUaLHJF3TfibjX8Wee6coReAVMRcCD0hb6hEsfabk
ADy2yimn/BLksZEqMTH6+Z8W38gGNm+EQiJNFObQPQAtLWUFmROGdkS/1ZoJ5/RGTlS028VewukT
HD7jzxsxkuggTBr0hyXC+rm42QW6YyezNX5tCY5t19lVT3/iqYXb0Yl4vSf18SFPKND/X0RoC6IH
8nUE26cuYIGZ4OmBVd70ls6BA6RrEr2WlevpVZr3jQNf6oywI+5oEqkRAT+Cq3mB6Ih1NZtC+Uf5
Wyw4RC/g378jDhkeJUaBZ/mdahnYSiZRbuDvAV7PctbzShrwDEaIfxgxTi6du+AD3FNQsDHI2QSm
YD+L6QzmTtlaJVh6ZrwQ/i8qW/efFu2x2D6nAMmcjEFH0mICQgU7wNG0gOrBu2DRnutUWLxtDEBb
y7JkFCUK3zedvS5vu46uIZArry5S7WQdxlXxrEStT1IFSw0MLxXBYJSeILhiwAgFWhU8AuxBfHoI
mJaxy4TSZOYxIgBUDFJnAODfz9whM1SJZUrUe+EAp2vVbYTQKAMIU4b2xVWQwIi/rORR1g07ppHO
ZF/T4KDiOwvhUKQl0uU7zMTfSnnqc3dPkKkGUoz6dcU9S7wnWQ6hpvJehBuer1neirtGuRcYGp3+
nJh3s3KnZgQUU6ArXklPMcTuuy7guYDTLIu2nA7r6RPOZMpQinuJYU0xZdP4KxelL1YggrlxNqJH
kC6oLwkiw/PuQ1yH8Z7Gro0rW8fGbBB6cgfw4ZAB9vjy7qoJlYC9ngewHKA+F2xNynzr78O70AEE
aHfS0dHt4g1CM2CKFIIqr97t0VcK4f/NjrQwIUuiERcQYyzTFbqNNLVcQHMQRRvf5o3WnqXpPEEH
UZWwjLSS1NIg7gRq7XridvjnORUCeV9TKOYMpJ1u6+UqpYlhdUv48UBKcsHcp+ILKMG0gEriN+E/
iJZPTBtR4rVl990z6I/rIIj7E0xk/+azz9G+/22QaXN7sDGd4nDqr9vljOUylypElcQ9mU0TE39B
cAMpVX0AgAS157pq+XmIH566EQ4tfB8Po0FWFx/ln62BcxYF3HOHnGTF66U9nZiP2wvWUMhFpbzk
XBeacfJ/cv4i0lt+gvewmW9cBE1j902jBxJE5hPnH+PfyEGx5LquKatdsvgs/1GPXI7G6fi/KbEI
jG5KJsEGnAHKmRU0S1Yu0t+I9YZwsBi419qmeu13yj3Nltcu+hZJJSwEJdewFGbA2VQk9yXlKCud
R5N44qByWFyKP4WxzA1pC5dLBFESa02J3lFqYMXsIl4Ko/q7GBUyjxCl2qD/WSEWEUrxPa6s2GH0
9sgHQBuAUAsa5e47Ew3cK8o1dqcGKKmAH4UHUL0EmO4yReJCGQjlA4sgpJlHovtYItY9uLiV8YVO
kJRsClavP88EVffzvRGrO72HGo6u6mp6TT7NRALNel6uHR9OtfcJAa2tmEVB/Wb8q7FKmN7VQQ6q
U/pr3w7nheMGjg1lQ+bDq6eVVosLDYjruW+nCjHptJQw+5wjDiYg6+NTqRJKMuXd22hTolLv7qnT
4FOTLU75zUGytuHNFkeGTcKAGUzemXMTzSERwTkdkUb/yU24ozH9dhv6d+DQH7xXhqkLKaL221h2
8aLnN/QN15IF+fXQ1OXP0VNbb3DN2NEatfmE+5QrJLdVheZ5fTyDcqgoenoE1WZevvlM2mPvaOqf
QCvhG8Kj8Gk/E/mZdWcSdc7H5zD2zRZCS+z9kycXCFW1W2UPV56muKZdZlCe3lhQ+TN78ubgYyIH
/ZgQ2BwM7LgVnEhW5vr93NGUe3n6hhCt7muIBsTBT4V/CqSBa13QY3vsk7AES7iqDi/doAQXi/Ie
rFUVSnpAVMMTmkPhAxnjmsKFi95/ACHrR7gwSC4BXP0fhXGrzkeSiWh0YdpRc6rXtBecyBwVz43E
e14nWkINxM8f0S89HoD24v3Ap7Y/8wBCG5hAoYnCGZE3BQ5loTWZkPY03WyphoH1cKHFgzNSAjf+
d4iwQ1kPsbt/2JhjTv/CWWMMlRBRigZy6NEDnKghvLX0WUDshGyIaY/eWPJ7cxOfW4URjYZItAPu
kcm8+O5taUukASoNscX6WUhdo4xusUYAVNXZ1Le0KXTV/ARLrVbt6aXmjRXVyNZQoLNewc0exii8
2cJ6wFmilj4DNSXenoJQQp3+Jvb8aJnkZPvAxsSa99e1hcgBgk4rT2mqZOm7kWSc8k9M2r+JeKyY
p4m8bV7PXL5eTKHET0Kbgqe4veu0r6Jb6VKW1x1oY8t9dqtkMOHfBZqsCVCQ+gl1B+u9ewaXR/xQ
3xARj/qURqMI8mFzT5tprttLDYpfxQwY1i/tqfMLd5zWPrR8+2KiDFwjkphKJa7cBcob8v3+CbVo
QtlAu8qY4sPGXzT5EhojL0Iqzk6+0E8i8eBMAZSDd9zdWC+kyr1sZ9hqjKwo9b9eHXnzTVIwfQ7n
ZRoy9jgyYD3hoLyySRREOoEUBrfACkNj0PqRfEXef92zKs5MOFadNp8Z3vjHA0oJzEFxe1j4IC9v
zB9HOwn1kEcrBgtgtJkk9Mbn1+gIjcYCSxq+XGhUiBJiDNGe45reQhoXRSpypHsMuMhuf1wqPfpG
kTqUcA69FxP2QkaMT2Io+qeY1FIBQe+JGwDTx3PRhlbv0aaZ/8KH8mXgSN1cUDUGC6EuEQflzgVV
0Ey27G30KI/FztGJLcC/qreu0TkCm/oeZ35hZnEhKdn98j3tYXRbmzZLP7CjFCEeiGjYALlIVgbn
bl0h8uGyi0IxWNA9LIH3DI5lYtOUIe2jorX1iKrMX6uKMBwzkI7T51Njb95Onw1GtzAHLE2xvZGV
Hwv5U92ZnnMxPLjSr49NDliOHm0fZ9t2bvMFyzazxCBBhU7wkTe+m8lm4YAJDAV1AckdDi2YvCOP
Ggt5/W5sadlBYbZcfINcvRgX5dGU+NJKRhbgRZMEIeFIkKNmL3dPV9iG1JeWTlfXoHsH9a1GU2ZF
Q75KBYbp4xIRNYETBc+741/0ErBKARxs/ffr7unolzSfr/66QhGaqiwgjlu8zogxrOANuSV4Wzk6
CLmlG0YMbaeAYt5jcXH/KWufgVzb+JC33RrEFuxdeOYU2gteBKYtUL1aO6+IYjiSClnSV2tj6SfJ
/D2sC9Zkul7rDTtfKacamgKB5GbZ34TWanb2GaWW7hLfQ2FACv6Jfm5GeYDbhWSZ3Y1K7ZcLLjJ5
+vfcCbAN0/h9KJ8quMbgci/YmsgxLm0EkW8RpcnWA/Dfr2+TP6xs9R5a0H5s3xb3IRTQF6lFNrac
MrUMKQ/3F77iACHUsjvQ51sZk2OGRLbxiZyoG1mCmiV7EiMBkx76LdO81kCFyKoyLIZESNS1bY2U
KYms548QAAoRCeGAlFl4eJwiYHvpY/r80cu2KnL3AjgeTnBWF6W9zYx11RxN7aOgMNV/mBB6rJup
0PmVwp+tZVK1wwBdNp070mGpDewBY7IWEr12y1YwLc9eBvV41ey/ObfNYtfjKaOvcTxC7mFvciz5
7F46MDGzuBKHf+vIcBHtInxn4hJ1ib/9KdVjJVwsbcwcICOzlxFbmkrrrf/cPA6lQoaROVzEH6Tn
4Nj2d90JUXxB1Dm80P6NZvzhQzO2UUuUBBhTyKXZKG3Xp0LOQ6jNr7+K7c8z/LwV/l9WOJs2SnAl
aa173UqQIfJpWm/AzcH0fJtPk1LoeJDbTsdBFaIGmeP7KD1WE2JwLB7hZtnpAwifmgTUdSA3EB2x
YCGbKB4mzonlpq7kE/KtwU2JYA97B8L4esFM4z/MSNvM8wsYV4aml11K3e79MqjHbv8407izcqSy
MV/cpJBh0Xzo3d2ttdgsc0TPAmpWPO6Od35vkXCDwzem/HBVEVYpT2OZlXk9JDcgq2cvmXwWmGmn
ZZYB1fI/JcUFTeO83O5UKZlq1UpWiagzbDciu0vVSG2f/jDGYQOkDqodtUBnW07XLuoV25i+EKeN
bon07r3WPtXsCrvfq/h1B5iTHfwUtK6vY9GVeCFf9OPtjxAKKj1ynhCtT2xlmYZ0TL9V26knnxH/
kUJ0774pQmHTfC3Wv/+0Ra83cpAX9TApDppn0bZe2t3Qr3tMDFQAnmN992rZ8scYqAmh4BBBJOVZ
ahM8SYLJPes+wZO/zmt98vsv7PgNoPghOGnBeG/CbxTRiSCEzVF0kcGcYi/obTQj+G5dFqXVncTw
FDpB86T43GoHsjBOxjBk1ooGCA3eh12nOl89BtdAjoep+b+NSS8kf/sGa5hjb9e0w1I/NWridi0e
AGFrp666g8X8CNPpIIbIwvLRKnZB7SV3jd9gznxMbrAjZLlOtp1ZN0kW5LZ+z5B/NMFXvZHhGwCC
0YwKrGsC18HXOceJBQ0Ir+IJ9wNNMBamNeCY1CcYZlbi7g42U4+gLlo0w5F2IszTJPg/kOwKEzwb
bm6bGXoolqZzbo2ZQVd1fmnD21Kf7JhBh41S9t39KXg7pMKneix4OzI5zSG4UFw3AG2jpb2SU9xe
tQ3/+Kh4H7/apjL/2MU2SWZaJpfCu8NhIcCSuX6FNOfEGWj1/YKTb0YzsqTmVIVxf8sNYSIZEFVc
Mo2fiu/49Jo1s7SkYyd7qY0F8nWQZOOKEMTDcwXSsDvdCzCjwoyS0mXvfMej9jJ5Ir+YNFhCG6Cd
iaFSIX/tWKlSv7f5vzBoTTz6WJZKUi3GmD/3hyGuWGR0EvOxtdM7F6ZJI3dTaVPEX2zJ8DYo4DVL
OaJ67ILFAeSADQF3QTLM8KcP4AUEH2yrnrvWVO2+jlCQrjDimWicEevAZPZf1eZYF0TuzvX/df0I
qZf8QVjWknQZ6HxLDNnx0mVKBsDz/iUwYVH2v+nZnaYrloYvsgkbFyswCrpMYeXFO5CCBfRGHJ0l
/JzwPzhFoCZ6bAopTbdwyLcFVDJAuQV/YF0fhbREe2taSU4GbBvyPC9RsoOnMLZw9o6NZg8n+9gs
dIorlWcUNkK6zs0gTkKVnQJPiackxt7vFfIFazwL3xk9kv1q15X6oGTGaI182/KEI6LadBTyf5/x
hc8X+FqQUG0BzvB8pdscogqB3KMIZcyQ4P4RGxV/ltG5Umjbn1QodC8rS1Qf1cftNibADoXUJ0BI
X1Oi4csJdUt1iM76WUw47yyboX0y7fdSJ9EIWPWrXBWvmcv8BpmtKoFr7eRRoKImX8upREZHKOz0
AKkdEboVhBPLiYO1ePusE40UJcF9vVvkg8Oanq0S94bBtZRfJ8zG6wmAxVoa3lVeuR7GlTWC5atT
MtcIL33/w+ZrAmKyqS9GGipIzQP6X+bVnBB7F5U83R6yknZWIyiS0R0WOn0V27w4WiDxr/Ch+I2P
1RsIEhwGDE9W1w20pm45biI9hFnE20EuKOZXD2Cqv5XXbJY6UpviREQL4M9JYf9XQuU2Pqm3r4wk
EyHXFQtN/cb7Y/QCbxdsGRi+iUTfDAL48uYfhlRJiTPbJHKkK/kujII+zQaycg/dNjDgfOJpd3OC
07rtjDNH0QC9gOVryUXn8Bp9cTV0O02jri+wU1OIcfhVtkgEXhZI+FVKdx4cRYQMb6wi7bKFpZkF
j9AZhs2x3+mXoG3JS+7LvAbnXyTIn9ELHqbg9ToFcE46DHeU74Q4j3thS4ONUAK2d5pJ9k8UzUyW
dLAFmF2qXaOhsL4q30EE2irEHH7M5qS/h6mynlSGLpu7RnczQ60EwyqFsHezgoxJETZ/3/uUFnik
82/Y4qBDTYfsEDowfLFVNE3kkQubjdR+cSISwvdC/W+hcJWfI2KX6kBtw60DPBtBCkSJlz7L3nE/
0RKHctKC5/4A8cszkscnvttF0J5tOwG1D7PzO2iDXcTleXU8HePIZrxhIx3XvW3HRrxsxALkvqCf
01mK8Jyn7Jh6V7y+AGH7IIPT9gdp4O1VwRmpjBpzNTVJJ+CVF4z6fvFM5bk/iLh50Avpw/C06ffN
9zECXPCZMjdHGVGE2SIGoVxvN2ZCEHxy9eESIdB8egTC+77dp/pSqmDogDe3VXHqXbPoMiLD5BUd
aAgrgkzb9d5Tt3gkFDhVMfX8j6EZktSYfc3yS/LBKNSjuIY+aKDoLoq+Ajpkxw7N7eVOVpv9OAfc
Z3NxCLx8ogEyFdZqO6lobIIfwy6uQn9Y+bf5M+33P981AGpG6VfW8uGQ7cjNlHVdtd/B/qhdp3bj
M/iPo0Y2a1kjz7ThdXrm8x8R3kKm769inXW11EhZ05PbDzuCj1SKcZ6yaxemBUEPsN5pQEo3iN+U
vnPH7PhSZ3CvHC+iB1Q/AgRYKVn8ng42n5miphOAkumnbQgC/HxvUiNmnV3Eb1cP9YDAn8sO6cO5
Fj85PgrMmqI+W4JxntF6MWbXXC+eMWW/W/KVNMmvGKMLog7ZBNNoFCpV7SGmFiMvH0wodeSnaBaJ
GmJESLw88JMInVq98XIEQE92yiHFZ1CQ4dEVFNGuguhysWCDlom47W13G20K5yjbuWsDzVGrvZ96
qf5G0n8ft/YRJ5it3jI1er8pMDiFytls+K+U5uimGo9o+svxTikm3qY6/5M7HhaubuKZNDBWDwRK
zIISuKEPX/WT9k8vpyCTT4apvbjsuiZBgk5ePy7AMUYxO7LdD/gqcszIVDTZEeA5S7PshGSh8cZ3
LGvj0zv10bvHw2OIERAUcXB35NteULCOWx+EQnYLu3bhIG7GjYTkE4/v+UKxd8D32KocELcOz/Yw
Oqoz2YVrlKb3Trwu60hYKjulnxV09qQPgwm44VxyYJ2AqhqLguByPdC1YiYBZxxFK9JMHzBGvWOG
R7174gmMfIVR/cgFHxzO5VcJC3ciOUtQ2eDfTLik9EQNiyhfjx4HHhSkRvwzhBMlEj3SdwI2r2QF
NyT5igJlErvAQWArDV9N+t6gleXukmB2T4jvpR1Dc61GmYNgTcQywlDslP+JDptI2IKbTa1Ovy5X
yVH8Sagje7ecvNP48eFSW0usCGrMJbyUYCQ+Teo4v5Nu3UdH4a7LBLPywcrklrZeK1AZM06KdB7c
QrQW7s9oIEmtVUFJbLEfpqefakVNEddi+TPU0szeI/2SIPJ2p/3da6blbOdnT2b+jFuE5orZUkVK
jaoYUTC/K9XrwlLDkL/DNhwjx4gdQGjzRfXMFoau9ohqSgbM+qPrWRutMHhejEIf7ayUftxm44o4
gKrOZMIKl/y2pBVYvQKHvf1Q0pR+gcx41Jykmkp4do8MglzGxlV+tHI8gjg4CtCOoNY+Dce+xVTt
hW/eXRFJojOL/rw7UGU9lFhL93ScLjui7j7LUYNhVBJJAndFC3aTsGy180hOWV7gCIPWqhC4UyFj
/ZvuXnjkoLDr/ScpmBpcNWYGW3NW3Eil7kSta1xFaWmS7aSS9xH9A4zbqC20W+qPbBAjpiF7n29H
+dkL1TGOHPZWWow6YjDDgcv0/4VxOuyXyfowuIDhQ33e969u13YZJgb/HpZlpaWpMLjqjCIoGm14
70Lm2VkHBo8J+nP9DAb+H6pjlJT9hcu2GKXkkAWnMnOJDLOG2IPeEBrQ6lm2YlDktJxT3Jq0Whgp
fRxb4rh0SRliRLqGFlLYmTduyiZNIzzTeIpYGQU25UUtCTGW4fgKtXguZBTsKcgbWNw9EBv1yLws
y1Vv2OhqenrvX0OatFvh89yyvmQSo5tFt9GKT8pigIUT7kdfVqXOtQtZRpya+0IegCk3Iccm+Jju
tHLPC5oR9Lt+KlDczgnMC6QK89NKFCjxdXkfQSajYPZ1eYma9cu3dso7hCpp66pIUfIrP9ogeWCZ
fJ58V/0Yj+3fEuksbp6w2IbwFEqf91qp9omRYE1vCTWYlVVCNvCMcZNhlZArH7BK3KAc6+qg/OP/
JN+37oVoq4SOoy0c2M/wkFd4BbfQBRnbmFq9dc7tToJagfk83KUtakNebrvFBqfOrKW+/k51caZz
Jxndbl7sYTuBXty1JaMTZ5yJon9GnhsqyGDbb4gZXDoVnEEYFodWaaVbv4vr7FDl4jc2BMuaw5sX
ROv+xYW6Ns+4w802R1ubMiXp0hAk3e+aaO7YZ1gCiDri1AOVv83bPzqO+IwbdVvn96UwJctbzJMo
djQm/yA16MpOpyQOMcg3B96nLPz0mB2h1tiIw0eAiPlFCUx8KN+2pAFNbUXGBWm2HngMj7ntbBmI
WuR+v9DPd5wcvs/pXLKdzrGEsePSs5mmGt2VEOk2rdGh75qwcUZw61lDhtSlYz8bDTf+Bp+L/Vpk
YjQCLIw+N97xoIzNbIcpJ6Q3S4Geb6kv/0w2GOR26DmklumpDRfzuLPV1YhfRcpiV6aLktC437Fy
1qM+EQl5Mm8jbkLFEpw5D4AdrLNQUWmgBevPhnYVNciWTqOZZZhb4KgeZedrKK/fuYRjf2KPIaKD
A63VtpUW9FRqv1prwEtXJDzox8AETRmievhkaJIG4fw69E4y0peC/tAbjWato9Npfl6/3WsvG5Au
dkAxaaCzFMN/4tUIYtOYgl3xzHpG6HJraqFDUAIBdnPT0lo446szu8s1a6fi20k3GIIhBcvW9YzS
tmWvDpruynhSUwReqYKduHcF8XCzd2WGlg9MAHZvVwqyu6pPV4Q2nMNtxe6tRRg5p1r8l6rfuqjH
YlTAdq1s3muTKyXjv5C40f8eos+RC/1S/xFvLv7VnhMnsCD1pNVM90ShfW4Mnxz4reEvoRAwZU1U
ibdBpp7LD7az8+b6S74PVnxEBeBzvUb3rR87hIMF9Z9xHtSqTqA6dgz+t7Kt7PiajqvI8GI1AaLa
fN3GIBB2RKplg7hIbKFSdh8Fjc3k7wODdGa8GW74tU/+zjcffpKJbLMa5VqE4yTpIdx0UK5L7KH/
3vmrb6T5h4Zjkyy5tezT9Smc7KHQfz3Up6aCNmKyVTmbjhQ5hP8C+tGTBmcnEzwqP+JwHajfg388
IYyR9JvsI1Rc07Y1kAnFaoqRJCexvMGYdHRzDHlG3gxwHI40bdrVtXll2saSr4qYKYveu6K8/y+l
UWUb4HX/p6v7wSAV7ArXpdszBP/4Bs3LqRn7TXX+CxhmutCu6KUJRcPeivFL8t/+FZXY888v9o6+
t+W1oAt1I+3cQVX7ucrAYD2EVtntZdn5QLFW0ZWLaI+/PHGfNbrMVIG64xVA3MLWhW6UzTy3WJON
MklH+U+3bO4FsEwA+oOxS7itM9mSgNWUbAl1oxdgWZJ1jgr2vt4mr2iKCOpBZzVA1HaMLoX5cAKk
uoR48rNIsMoNQUfsobs7HwegHnAt+2uAfWaOhse4i01Mz7vXezfip6vqE+UUBGIhHFcl/9YTT2eS
cE0Kwq3YUiZ5bC/FiLXpuPC566msSXzGix2efLkCyGRgGpZBwVVKNvAb78NdI7PrQyzoA1REHUca
W8hc981CH1U3nayhvi+HPGB+AJyaE1qcpOLJe+Rplt8QFGOOIz0xWPJg8rAk8swDJ60Tbi8o9jXD
DjqnU5FcQxflgfV2ZhSCOXR/QnSNenccPfuYOogm+jPTUiM1w11tig09umYe1SOJBhPqQ194wDuE
kaUnm3XeW2sp6QNS7nrrzuucR/z2dpvyQHYoY/0EKkdYv9626pKTC86iDWPJ27GVH1E6t9wXSJn+
8w5eq23zjH7QMBbrDpOUNjlMDwsiBWv/1ZE3ZURyee3pIPQEzCyDu5w3GD153Q8jQWTNdxH2zJyz
gaGN+TOafvwjTb3eAlbAjTSjGKkExPZrCGyt4VOFX9isCZdmJsQFavDl8SvbilKhpYvCht1LccnJ
4sPRegSR2mDoZy/6uUaX35+tzqOUMlTYqqeze61WRCpVmPSqQf81cN11PrRY9h3/cHtVPYyTbzD9
zk9lvRsE1yu15LRBlth0oln58omQNK63wZFXy0cPD/7KZQBKf8naTfnMOplsXKqseC3bick2zzMR
mf9nZXZCz3k4AQhDhIc9oXqYxzDtBt6NNI5EKp+XxaJA4FJoLWNFLYSnIxaL5G3VrfLE8WVcopXq
vkcIFt8Cm0duO3asXo8hIC3A3DxgY05CbisDR8wCUU/p5VJoZFgSQdlximmS96+d0e00JYBv3ThR
7sAT2ji0dSfPES4WNuBsG9LphHkIIsOu80TyEhRP7kRHwNe6qdHrGyTQ69VofaOjqAmNMJbkY5Ol
EQW4puh92ochzu4IwE7VcDtLIrPowiPsH3JR3V6aj8joznAKdzwz27dMrz+UbahlAhPKXuymdt3d
F5AEHAWv6kdQkLFVt3eDtrZ7PoSXfUEM7hGvdrS3mU16ct8L3cp2ymZpcj5LKQW2JhMSv0ch8EVb
EHyRnJMMRWuufCFKNLf6MKy1XEw5PueRtMehbZl655BwZyQiqGV12gm4Lv6Dj9cz3spIM9FjBd+I
laQdH0rNyu22br5TMJYEe4tF/nxq8tvrek3TusFp5Zfxh08b6of9NxowEcykpPYOMx1lpReS0a8j
8EPuxtCCssHI8fz+a+BkV5mIoiMxJQ7CTxxlxRP70ojzztD8l28Yjy1Djoabm1WGbz66bzD0llOw
+o9Dt08xP+YBIAvrfjfIUi81XKn4D/taA76FnMi2FVrA/Qi3fXdE5/GdebsuQj+r+OlWRyiEtJCi
ShlE+5PwPV4h6QiaL0k4YrzB0Uu75AhyuoxbP205mDbKRgzeZUF0CyZL2vWMzbrfz0RRGDitNY/L
nkN2ZD/+BVQt9Cpi5wNNNE0N1dK/Z0L9MUSAwH9NZ8bSg5gIMLDTJInuAxxX6PqwyYZOTrPf5Rbt
0HdjocqYllGBi151BZALLLPkkzpDNcN5sv58LcHmGv+3PX/wiL325hbwtTV2g1d9znTNmqP4Rqlo
zfFK/G69t8l77YFrG1djAwu7VNAd+RiFSsCBNi0Dw+g2Gw3SSMe2XoBR1BtmaG0R/Z+ra2uimyN9
SCXxX4qo8Qyv078ioMJf45XKzRL95/aRtArUZqbSlersO6HjdAQeeiZRAxHLSIJTn1jMnpseMg7e
22+uB7HHh9W/Fff8/b3aC1ULqsQvLYZUdI/Jw28wR37WqJAJy7y/tZ95HQ60anCoH9+PSKRoi1AH
tKohcRmT1xNNMpJu0rj/32QBBoGPzYq+Sfc9uCN7b6CnR5oTZSQTyOUKv/X2zkdZQa7BaqTh7O3L
m7CgkwzwzgXRxmllfcFmOrujYGoX+f51BE/umi8VrZx/uZ33XkX8CzYahYQb9BGDX1yiDVqLy03Y
ojnYgraNvXPIdkUkJgI95RVOgbah3kx3IyRyK7EJuVMdBZZ/HfC1a65ctMa6yL1Q6pD1s2REYDPi
QaYEXffq3brTdGKoz/EcWS+L6HUVsDin7ExFJe5B/9TJMGj8p/c+fL957kvmzPvZ2GdxPltn5k9K
kOuUUUKAU8EAsE+5Sum2KYJSkSspWlrUYPm3WhaZkZwN0geENtXiUd94qu64J8fLO6ibnhzRJdNM
gO2ks8fD8bvE3OLRJxktUd4LEJy2Y1MrkZV+tmQgIUXsy49x07/2NVITacjE7aurTDeSMhLe+uQI
yTJrY3qr6+1cERsJGzPiVUkagc8AgS2MfAlRm1dLqTJbgLYzdpQ9TBKMt7LlOB3J6Q0mBPSYaXIl
H4WkdoAr0D6rEYBKpulmOVnqPUcavUrmth+MD6DOxX5QC1UUgbwCjLysiJXoK9nRQZXPgRMAytLp
QooI5CXrB3jGrR4p6PYhkHQF1UasyCyMQWzl78KHphKgrK6YwVCGXZunmwJsZCiH9Xzd4rn1cTk7
FNDYz8rKtFucymNOJcZVeN2lyVWnrIhlI/GtGHUV8K4z5Ixuzu6SkwZsHCKnZXK43yFCV+DGJoj9
W74Zr7OqS3SNkEV1arW9tofVoDzFxW8Huc5LbGEGof1Up+VzwZXRldRGzWkDsCsAYChef7xutVaS
RXM9I/Dm1cZCygac8ICwV7jSbzWwGHboMmzGyfg8Gq+zdbAmUTdBbWM6V0+RaHVWy+lNo/iiGUdn
Z2UlreJ1GaxyzckKR7gVNCH26LmEoSwC8wDh6M5+Ff1SKOd+hNTu1fSyrSWS8ru9lCj94Mybe1+U
37eGuEUjGqv7t3rLaY9w9z43nY51FAw6pB049TVGkBdU6XANojs+Km67ACKU/1T+QknwqLiJpghW
MewZ0DPAkBIlfiUQLPDboKwVu9myUVQNCuxi+0Oul5NuGfCVOVP6gTLJmkqoNOx3OOiQ3eqtXi5h
bYH1KC+WG1axahCklqTqJvIiYZdkLjZ5d9RSkl27egTGvWtlWgjGhhfudHDCkNATAZAT6Cc9f3yk
kJwMubrU2OQj8ug4/S5qUiQWYEK0u5iWZv9ZAc8PmVyWACz03kICCdYrDqJZDGOHIs9EYYfzNRst
gJIOJhg4YXxLeCZlMUgosmHyD8Pbz/84Go8tNPr7N1wRGS4jhVLTD1OkKPB8iRPlOy7wgyOvNbUD
RGDYGpnTsb9pWh1/JHF2HnOrOGskk6gChCyFOKdb6Vaa4DVuwRg4YMlgXkatNDd3gBi+5B2oy/Fb
amos7B5nKp17BEG0QfNSk6YhUfzbTeg+WXtdr0/+Z9z0clvIGNdn1Atyi+SWb7Rr61shQYcLWOsv
lhUvjBlwlklop9jTrWvhgVxdxFb7BCCsX+JteT3p1BbRXPa12gpc290kOW9XDPsiWs2BBtgakeLL
RlDcHO8napBsTswt+aQlZphOH2hUrJzbFnfRebbw9VfvBye3HXezYAMaqA6bMgYNSvJpL2yGQAB6
lZNpNvdlVlvE37oSd7gf4urud9/wL6+ZeHe8YSwMxlP0s0pjGFPmyjET9opiICm11PcQl5ZNN5sS
dG7L32B7/0Uj9RDY/u5PS4h1MzfUUxUXCegdtz2He2ERvdGEae21AN8zNbSN6AWiYU+JMNg152uC
4/3u2K2OD4qFxYlCK3o8zCsc4K+xUOv8pECIjC29ZxI5vqp1WTXtTvk0N2mKWqTdVK8bm6GdIv8u
ysfkQYFEI1CVTDzrAzmWb2jl6wCEKCQgWxPJfX24/rHoXgjoD5I44GxcHv8n8AWNkmEcxe9aHlv7
+z5lLw0uVn2JwyUloYCZTixh5ARU1WpLwNV6L3YB4E/zFH397ZtFTS3VCk2xDuyT5aXFe99g+Pvg
J7v/j54Os47S3VLlcMMkmuVLGJcmOrrmzONaaYpOem037ht/mX2I5piSEewiNUxiouFBSY7g4yGD
0+K8uK63tThrrs0V58LAlRZmYzfvYEDvMItIg6YNx+3UTmnyX1ygfcqhJD+SHuIVpTNA/H9cM94g
BCNlwomo3CbNftUOXO4IPgo1I2ksx/QHTE6bcdFPEweeG4TZCTuS5Q4FAUZbRnBGcM+LaGAFXXaM
3juiW+nflrJVYtFeU3Lngh3umptK8RgyKrqWdDKZn89LkFR0eJd4hrQRFmKcFYJa5V+DCc5HdIZg
BBkpe6mGiVxjvc8rTvlX5RjN4Hr+7kR0PW0oK6Uk27FmxEwq1YpgpjnSTqAm4hW/27WXLXqxajBg
4k4Ozmx7HnyRDJBGs+6ZLFnYNXZQGBpCMn87KfQLGjzqwxqGz2TGdc/9dsD/4PnWylfM6EfrxYZx
sQNvIZ8LQp9je0LGgH9zcgFi6xrz17Io//Xta0ZLV9dipyj7uPBP7VCffJDB8kzm/s9jhL4EXA2r
oUBlVkJZw549Qyue8enZkPDnsNMSocc2Kg2TkXrz0ODKU7xWTuAHvO07daCe2CcIOMJ4oA0zfMhJ
EdE+Z2mcDs3WrVkpA0SgnkZkxcV7FjeCPnG2nt5H2EuZXhP59qd0xe8iZczTKM5ol9mp+XxWGHh7
UQtTMDg1bjMe6QFvP5fMcvRyX1uSO7zsmujk32a4BEfFRsvZY4j+49QMz+lNAOdMVwb3kgbXnULd
GMVJVTuU7ctbDwKQFLDF2EL9A0v1a50wMpIQycINkpuhKm3Uk8/oDEsZ3x6xqOyFBuIZ0WgvEEVC
HV6bAqWL8TSkjPH2KWMaDQlFOR10t1Pwf2fCUThBtJq+11n/BQYpjw4Ju78Q+B6sURVBAQV77obP
Mx8vP2egK5/xmUKvQu088p1G6BPznowXR09z8ILQh5LQmZXlO9GwGDhzNm4u/+E86nUC1707o19L
xz957cjUnUx0JnhTdl6Og1UKCkIS4OX0z8X05FkdZMgxoU+81h19taLVt0kj8tJSlo//iBk+kTKM
2aly/xPbYt9v5eYKyLaDMRu1/fQnF3O5gRKmTbc+AFUknywydjV0XYNWVuE9poNhknmfmky4kIlu
jC4I+5wrV3sQI9vG+ma/mkEaQewAZoFMCE+IgxZUnDNWh2QHCNK8Oi9dM0BgEGPUS0tV7p1n+BfL
RI+rGKVyg4p4dXBRv+4ErnQy6n6UIK8AvK6JdBR1egfuSA4l9UPga5NQuwxQyjcQUPzT5HIS2A/5
XB6ZPdh4QKFRl2EtQzjy3NW+cBmcw0EF9oF2awnPZ9ldAkO5PKPTdoE9szkOUTNoYQZEPquz5WSp
mCLEZ2P8BPtFrvrCIDnBJs7KQBhzFNgZFfRIcxHQdBhxDjMc3M+p2jgZcOzyxMGT//ARCIQ7htA5
8xRcxq6GGABoHbLqB2rK+nQAh3VVNbc8hG1r1iUeU8DGv6Oo1saVaoO9f9yx9qxVMz7wUTsmEPro
zwEM04OI/DBreX+xTls5ArQVN8ld5Dy3pT120hP9JJeyDlp92MuIfa12vM1P7GIiWTodlAIhIa2Y
iN+uSHg4nleZDJXfywI7xtYUTZOltL1hDjWGVTRDJsxrnUACtIbfm6YGBqNLaTN1S+/3G655MyUH
INwx6a7mvrGlV+fXYt3c+FanCXiXtgjJPyabzS38mfd+ZntJbkyW7BRmzDMbd6jSeCsgxmpF10so
Fu7wXxlQ+jnz6CxPvtYCBw3x40Zbgtac58vjVhHWYjuq6XSdzFfPhc0RAcNnN/dDE4+wX8bFn28v
Bvg2lIfur9KGc1Cd222sqcL6Tb3YaK7xvhooBWPKSF1ViB1INAco5PQPuFCOw2es1WTZPChrXDy5
hAp+JJTYd6KkOp+LJrBBq4Xv/bT+SoOqwTpb/r5cPRQkYVhgo7PbDLMmGDvwXQLj1wSsDThcqrbE
nUv+epAhmzOti6xwaJCW65GNydjkMNGG4mXo+4pMfqbFm5Nak5IsLj0YWdCo/33lbtvdCSf1sf9+
9twKPDUkKBtJaJTQqdYV943UmCZF43QI108iOpKIUjsdkkIaF68CxeSl4jYn8U6aubJuoXZIZA6B
3sQawuNfszzyOols5MPqVznG/9Eud2RWPfKf8H3dqCNtawdWJ5uotBg22NxkguezUqLxWJ6i1oRX
dxxktJQGi1zipV4SFtLNluiYQkWJ7pKp5KY9TYGi2prr4e7cL3OSXhweCUlf1iA4b6ZoYgyve1b4
T023bKQfrdL7m9xOGcnxMDoWdBVibmNMK1G4Lahth8471O+FpqWM/KkKV8+ZnPu117gQIwnxfu27
RbcYtgC4H1fh5Pcp1cFaL/xIFEKWxe5MMT9D8QPGFiwxWGmlryJ3LGqa7CsVypm6Rrk2XErefAwl
zjK++zpniLA8QN5scdj8qlXwxhJS3cBPg6cH9suJLSHvmZZCj2Ax0ztVqFLRP+Qt2OMAPcnhEzkb
s/UCC24TrU/qlLmD2+oFr+Lkjm63/rRseZggnQbUY/AyiPa8OivpVEdhbDwVay9w1QftjB8Rxo/w
JxwXQK/Agwl0VId3DILi58qgjflGL0+6ZJd6lZ7WJVrlduFUpeVcEf+jtKuxOK9XZYtrORNzF0eg
D/NNPXSyxyP5Ea0oBFmoijawEITxuC++lf80aphX5Nn+qZwQ+/Bc19dkA8MIJ9jOLC1vNpfTRC3b
0KFehR6D3On+3ntsORRcZztHZahh3fMOYeboYqaKnyuvhdzQ+crp3RsJUeIWra4hMa9J8423DNR9
FX+pRIQsCGhMzMtF15Yrz0V1yt6dzlYLRzr/XPOsBPFIkymnx+fwfy8cm+mEpJ2f20qHvpImpz61
aFEqx3EAkDyleJtEmXYS8Wbc6NLYzXAHoWgaNANWLyQkLIdWA0411PxFGlZ3TbIQHzgFsqd5A+li
RMcjFmYCEBaz1Hn0soKWYjcWisjjCnb9XrBWZbYczRSqWeYuP09UIsmSdzuyvntTu0lOvH+9S+P/
FpLbx91uEjuw3fvGje4ErymooaqNhZp43No3UlUUkf4s7ECphu9B/pFoBomet3bQKecuxivbcnI6
KeKXb0BxeH4JqkktliMQxDPxT1b88MliG8P6+Av2urnjEDK0t8hE0BcpX+u54ODK5gAkNLJJncUu
xfqDq2+NkeEOVUyERs5AzO9XCMKoJEUrEEh8o7Ng1mC5iRhbTJ1ZhjEpq+AC/RWcMLsYbRsuRUOU
7hgBt638jSZLVeMZhT/SV84bBDYIhxc9V6BLIZh4V8fvUBYp/nd03ZSVG39gasOK6V+ZJeKdc3En
Ggwfn/WGvlZ68Ol55ZBHR+NYeIt/m6cuMniegnqKI4Oc4I9YaYSPf93WLcS4ihVmJ9HkYFgYfenM
/+HaZuDLB8J65mLlDLPHDMMszDHlRiz2Dyx1kxX8w7sC+/6R+WOPWJZ4LmDk03ibtklCo7AZngM8
uYW/9p1W7n9/F7qCU8Rq3tplo8Xc+zQssdd1HS3D7rlOiSzkFKi8nghB4ABem3toZtUEeQmNImR4
pkLE2oC6zTTs2mdkbPKhyZt05q+IPazU59d1VJQurpwqOt4KUEEPSP5DQHLRAjEg3wcI47+udrKL
bFAFDr9sPM5hUQOi+YaduXOk7hBstbQfCaKrHGVzvZ25pLAvS5/hFecEKlo1OrNcIqTMIK4/SVZx
xsW8AVH6rQUGqu3U90S9dLDXiBKoCXr5JViiQfqtr1+HVKnM0AurD2zLyR2qvPhxzq/RTobhQwYq
tD2r5AD7If6sHV0jB6Cw7D0D4N55bUg0rglE4s6zZsIdlfU8kk56rHgBU9N2tJPhKe8pIW/8toyJ
8ULxdTDn8h7xbHtMPX+2yqAKO87ZR5P/2t51WOAT4Me/aKO7P9k04iYahfl9bT52VMny3FFyg4hJ
YDLHEoXh8WDgaqCtXQY/ALptOGsC3Pcaw2RjQepV/y2E4pjFqLOtGik0ZwLtOvZNDiL3yL2L0frL
h1qRMKJC5hhSpNR4dyiXZ7wFPwmNmg+n4XVCsVU6JOpZHGuashBsV+NEQSzkioontCdPLUeEX1p5
BH7RP6zRyEeFQh24QQg8nP7rA1cqZUdW4kv3WvsWUobkMeAcAc2/7ntOML2SKEY2BnPHW9iGXS02
bzMPvkOJZ1egON3UEq8RfHuYEdJqq2d2QiRbX++eZ1cAl3mi2tCmByv0GT7yzhEf2QNKvG3KhWb/
pAUgx/e/TP3FWsTSry0voUztv9/hFZ8dXC75CMR+T6U1LJ3lcYE98LETfXSRTlKnB8U6h2HrgVmp
bMh42JfXnxZLuuZxow7c7Qn40byOxGkKudl8wHTqPw/k12vUhbRz5aUtrqc42J0LO66Pn5JlPy6q
QU4PVywRd/zlcdWmJwScPbOfH/igEKKXzpidAjWkK/vlYEO0BmiAV3SRQaB5jrlsd5jEySP93NE2
cCPDczz7EwKu/rbkAozNOFB7Ap+b19xYFiSeu1zD0IIcgQSWWRsdnDSWR8f7f4Gt6S1jIzDcV5WF
ZyzFu0doUX3v3M/Vwp5OUkBgcId+1bPVn80E5DIQ5lvwZsAIedNXZ/+zPK/pkikxFlMW1PfUDCrU
G4uKpIrNaZ0SE5m3qglp9BCYFZpv4mSUEehF9blVR1x9sfm3tZ4lxOPa/WtZvPFVLWBf0kWpYrxX
AW+fEF0/x9iG4z/VDaByNPUzdgfjpWCLLuYFWMD8S6wExo9hT7BED/kZPH0KQa9gD1H3xfySUWBP
nc669bUXK/u+fBt4VzHmOFUYK25qXlScvOEI3yv7JDmtR95YEDi054PVTIKZqxgQ3ae4+B35bDem
6QKw1MqIbWNzceaUtSTswv7gaFhh1tkfLLn0jcHsEqy/AKL4Ai0jKUYViIaVxpsMal6oE0hNfaPT
8aTgpLc8Bs24aZfDv6eD5FLN7yMhZU3cHw4lCL/KfRRtYFtSLF2TrT0uMTcp1Pgcae4AZW1Z2DJf
c+FMi/roEwH3EUKPTHUikXCxd7lPlK4wwqIdgVMUnPU1NJXH20zTPN01/Nc7vZz+StvBufJZ8DWJ
sq622kjp6IdONhQgFrul7RocwlqRGih6d+vx5WqIO8IW61MsEmc0HxOfun8xLUrg24pEWQR9cK/m
54KaiPuufL5hxbzyA79ra2Ujxl3xSEdvZt5i0Xod3cz90VYE8kg9mHwjYscvv4xIkwgkCApb7W3J
32h4TZX03J5rJNT7yIVt8a2hRWUgt6Diihc+pAZjkxF+bxRljHFCfCzuYDWmxhGW/92/bgkxbYYK
kpTDKyhqQYxFHJdj/gi+drMCn9C+3uWejpX2ssq9AvSVHxyzLukCWiewxSu+PJVk9003iI5kQxNO
36/8xHdv1CtSNk00ol0M+aifnKrcljTXzzLb5cao4sx9GUaxvOyXjjneryNlUn8GM8HK0gEPZHKg
otkkmMuUhcSeRfJhE1Qsir65HK5q2A8xV8gk3gorBPgkE890k3mIwNAwKfw8X4ze6EPIQzwgdyx3
lBEsdWU0v/rH/P4B/59WlBh7jZCTTDTR9zqdjLj/0F54HUjAH1IQsjQleyVhvQVxJa8kqMEFAE0O
0PuxijDt3M84HURerKbkSa44Aq789h8qQ11AIHxbSqQKemQVWHYH4dwPw2Bt73zkSs50K+fFVkDG
a/d/p2zuclJUo5iISZtgC8tK3MyOudQpsURzLE99J0dRUOtZ7K1zZMla1TE7pc5Hq28Hlb1aZ5uo
ztLvHqZK+DHKyKoxEmxv84HM9ewS5n4FrGANn4IGlmP+x4lBLHVeCGGWLztb0wOpgp7t/Y0XCSjN
2ZECRLqEwOB36/jhHy7I1PbMFzF8Tz48RCtUOw6l1Mx6XnPzSO3sWwUc4VP7bFhUoGSFuviCR4Uz
rFOzFFU7/XViC3B+LyoFNcBxbyNd9MgLlW0opmQLdTT7bkGq+UYOI56XW7otPbSWTmTLkC8DCr54
+UaxrjcYnJaI1nHwh/zy0ma4EHk+Q1U6em7vU532IhTnfbeXHKsjepJsC6zCfLp0Y29Xh90WU7Ra
JD5ABboL5omP5314QYqq1uL32sic8KxQBx52my4rvlWqInJXxLvsjVD+K3sz+4lZz7BwhCh75Bmr
rNqWh6PrjwE9VO8nK0kp1LKLROdqMi6Pv7avfML2i3L+Vn7+f90BFYwQqnYsIh2LRfqoA/dgh+ZO
1+iJCD6OdRf3I/ivrBdtcOMFFJzhX8r4jCzICkPuOxpE0U8L9ygwBlm6dNcXcp2HCm+LP4/WBFzN
zypfAhJelTTdii3eWTbXe2W/E24ge2aiWjDnLPo5Sx9KveJDoW8qPJOe79DHzHPNM2lvboSS0t3a
81n485/IO6FzcsAo99aysvYn10el9trxj+ZBZUsx4D/rgZY4XeKkbBO8/RoZxCxKBWZc0DUZYf54
07qkLinsBoMRYmTIpFye8wCemdYSYqDQBd4D9PSzMhp/nSejqQT1WP4w7l77jHIgDvZ2dplUHULd
ZML4woBYw3TLRot9p0tQxrtpcUy9sVPztmC10KRDNLjR/dVE7jFB9SyGKF4wnQIzh4au2KEUWWka
M60cOa0Y5Nug0oH/yXEpJKG0Ae4FHt9gyhp2D3riAs29+FxFC85JogY6s8c1VqrB+54egVb4qMPa
QYareKk9GaCM+3/vfeUH7vyQRcWM49AZdUPUPO7z59K9UI2SQBXE6oYc8M39N9BrELXkBH/noER3
nfZd+vorHlBlQPwq2HucXVzzsqn7XcCsXxb5weupBdZCubJTviffpObYf9cT1w9kX+DJAlvW0uZL
/hEVnAXuvIUkySXtqL9PvQ9CKKiImhEJ55Uo/CMLDehTrnnP6CY1givKn8JYFSMl0RPT5wgOHYhv
Jb8OwJTdPXtms5snV/O+1FSqDZExRVx2+qPQXrd2HttkEFJcAHXVhOJfrJWRgfdnfz2f3+04XQQ6
axgEw72DcBq1RRC8URDW7824GkkDhUCScr3N/qUXAsRZQY/OnnKqvqTNkOOnGhkZ5Wo/HVuDSG9o
l4GYnEyeVAiImvFLMlA0FL9BQsbUU+RXigMmgEMSovMNK092dSNHcZTu5ZLJph5D1QPjburEXooe
ao62yFedAcRgaADHIQ/MOjNPJl1sVzu8zVt2zMdFPH9T8d6Hx8dEsgjX53SMIsoMpRVhLlRRgVNs
/YKTyo7CfJuGZuFaw8P+cMEoDEWS9mMyiqu8XHKmViiLdTiSlf6kNZrgjOgFaqyNn5JEP021mSOf
r3Ue8Lcy5nG1ClbecSr+K8uPzzBmu4aawLTb3Y0c6waL5xr+cp9G+2MQ45JX5JTUMEzHgicnmch7
h9ETfQtPO3rAZ8eIYBMzronJyBAwp+csaYFcHwyDhi77gYMnWbaQJ5HIgaU3u6oVqYvDqsHQylRt
WgFwJ2moWLL815MIzA89yg+9IhWzC4oDOWKQ/TveI9KDMpk8i0V0qW/DUf5Tcrj2b40Yi4ErVwWF
me7BQqBKp0hlDVIDMMqsJRBoCVROcBB/ruG6fhEnarpsZs4Yu1ipYfxWRXK307I67euvMoUCOnG7
MfSFY4ehLO1SX06yfT19V95JdE8nfHeLUIfpwLIRi2OyH3ya5vtOTNioukymMFLushXiObXuMTdp
jWpJhJtlCjXsIjNfEBvlcOqUtP98UvkAIQeb6WLfaiVvwES9/imELx2drsY6L4AVrLy75AnqpSpc
pseVr33I5lK/iJUUnhTprUxnt0RDZvGOnmGbXe2QEuo3LrX9NEl1fKdttSaUg+5QfZOV/D7p7ke9
7DlnsE+zbYAJeQXzQwcw9uW/EsZ+CV2lY6bYg0ABwY3LoQ+qUWZ9xZt2UuHIKGK+yg+fy+yN75D7
83x+zbuoI8E5rQm4h/092NS+tojaXYDXQdzzGxVZenvsDskVgyspEkhY51JTn5AWP520cz5FFvIC
5xWqqsr76YykNjgmN69PXCyfpRydT49bM1gikWZCZ6S0ccZ1o35fwfnfJjcG+qgq+DdcuiFzoBQs
ic2kuxs6MXQY6BycTQ1zuk1SanOo3O6RFnNO1lS1u+1YEzcGWMEgrxW1Nd8rxMK0FnvZ+zpOrD71
3W8ZUROiqQwQ8ynzaiBNJU0LQyK0wjjFgSUGLA6zxqHYjc97wKAsfq5LK6w+VwLi9y3SIarIV6ba
jI6oWyS43Zvt7orwArX0QaxXiSSZcoKZe3ZnWnCsWC6jM8jl+eh2ouub6bK1bbLr0osdZNraNn3N
ph68m/jOXFw736Y/3XjoN+re8f96iGo23vRemQ+I+59sQnmEqBU/YCoV5YwKAsxFgvC18IbX1WKt
cRFDJx+zZdZ8UzyhTsyHvVE1/z8yTLiS+j8Q7MyxgYJi8hqALgvaRtP+2G7Tv3loHFgq8vpyNv8i
amzJKySIVTa7MAmKWksR2ocVgNa64zeCrwimKqDxAusiHQ2F4gGl5KQvBs1GACoXWbKnrJa82S08
7gVL/VOUMlQHKEdooXfZuPKWoCqNINpXMhDhkBUcjaIEuEQQ/yODqF+0EIfUS+BtNQl/9JDGdDyX
p0AkSjUJEM/Hbbpc173pbFzI+ElcY8GESL6VSz/QrTEHShNH/94lQjrDBupw2A4wezgDjbTrg9GW
1xHnEePGvrUcYjpyrJNmhV8tBfaz1jfUGyzcaldilbe1VSnfg6RXP4NCSxCJaMDl/mpcPH0h9ot2
DoBm5Aw97JJfVCbwviMnjauoDJIPnQF7OyF9Hooiogr89Eci7lKN3+Dog4YNIhwwKr4SPGJxPjEl
5qLS1x0kyF28nh6OZY02KSlTt+5SAbYeBRUvbE+UA0xBfuCbKDdsPfnzTnohsNva6IYk7yyzDleM
dlwlBg5frCwspcnOnkr5LB463MGyxa9ALbGr8bGSSv4EpLMOWYCpwZxIIZAqMf5a2uOC/YtOOnST
aBNNayRqcQg+1BD0CoCilKdxzoszoxVGW+GDgOT6Piln6V4ZXVYJ3OEXDmx1eSG8jDZ1s1baDyJj
RgINj/S00Df4kyVGQXWQGvyVeAS19z5gG3VOgiobnYTuL3aF/4gbqhyYNbHBm9TGb/Mu6QYDWGB6
qdETNUpVuaYyzzdribq+su4WfNpqoJgylaSphEDfG8qUDeWM6Hr7MyfohiGDS/JJ2jemu0zyMdZl
1zxII6tP4q3BvUlngjg3DCALwOoQHgsai6G+UQAemRYcHoHwjn5MCCDPxmu9OTdJEoDojsDFf+Uh
yx8WY6lEmMBUnK/USs3ns3fbawlXwMCg0R+WGOWQrp6BKklEioOKX+qCephuKsb+PpOHrpSEEseO
ucGk9hirT6s5IV2G47hIW7B4veOxponLMBLh8URkaU3jt+rxtMz/qfhetanOen8KsG1PDfkVzyZL
Gx1fR7Td4TRdmh+JuQYmp4/2+jEFncVHJgXJv/sGNAvru1eOXxpKmXLCqNhSZhrIvJkNWw9NXAZg
zYNk9J9QLlzsV9P3/A7lsrim2HwKyoXd+Y3lkvmo30FNCzqCd587Bbf4G78ihKN9G1QwuIVga6cB
EPU4n2NGpQ/D5qyxexEn9wlrvkfKctSltFCxZCnJjos6BT1R+VgcR3PerK+GOkVceVk50o+2fwQI
TgijIUBCyUsYGLKL0IgFEev07x/xTSvoCg==
`protect end_protected
