��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$Rx�y�<��wA�*;�x���@�̦�W�X�fa�M-$u����n~�%���P�$��W��kYَ���P7�?UMfT��q�6�U��k�>����~�\N�(�����X�e���/6U|)�X2pF�]$h���d.���9E��WG��L�X"]�Ad����ľS���8od����e�GT?y	7�������ݵ�^��R�q^]�鍦�����s�ae���h��L��P_���ާ��YЭF���'\��68�b�[����w8�[X��V�F�0͘3����q諵�uW� �h�u\V�?@��_6G�_�*�G���B�絉�f������[�G��U&�����~�F��AׯK1�`c��[<��FY���4I� �#�G��x[X�=�Q1��`��R>(�w����R�O�?����7�,(�H\�#h(W�EH=�������yq��Ѿ��aF����:�U~m<|��.��0=�P/���4ǆ���T(���IjS~���G�f>ܙ2�Ҩ��D"a��}t#���uc�ع����qHV(|��#�pH6����>��>������z����dn1�f�|�=��H@c�z�un�5.��s{��Ɉ��Zq��C�)��	�+"=	������!`b�8�
/%Ӱ�;F��C�����H�d��qxE�*n7e$��0���V�.��'eކiq���x���~�������
��ڰ�.m����9�v}qR�|�3��!����>��Xy*#5���n�skw�(�����̡���bfx�
�pMTL��؟X�[��]�H�qҴ�u	U'_�NۛyQ!���!��������ڸ�2xͣ݌�k����a{O|&a�3D�ʨ�@<���Drs��?Ō�r!4J˞���!��jA��{Vkԟo���oγ��%��lߥj�x�[~�aE�3�#���{��N[��4:�`��Ќgʈ!h�iW* ���*n0�ө�|�iT�ڍ��Ā�y5K��&M�/��W�?�4%��z$�&��d1mky���Z�X.u�aN�["��dO���x��RXBTC�����.���j��C�'d}���f�_u����R{e�"b�w-SHP����"�T��tD�qs<�մI���E\�~�]�P� �?۵��V���zZ0:|�gk'��@���w��|4ס���������P��C�om�bH��5��6d�r4�⒱�hd5e��s(�֡�d�������ab5�銦/l�K�%.�_�#R�f��]��0�U�4�-1��ĝų�V|������Qs�́� =���B�Y��A�O�I%�m�i�0�O3j�?s�q*�=�ԁ?�����m���X�� y.���T����|[㢃�v���B�'� �D{�i�)�����35$��0��r�5��R�f�R-�ON���'8��0��W�ۂ��Sh�_؟eTlČ�}�Nca�V��8��6P�y�ݷ1p܁a^�u7E��̖���d��5hm��yT��wF����l;�#o6��zB�5�G)\�1��WR=!+�"�\Q1�o}R�A��M��W�
�`f>�_|w�T��h����}�f�gR��8�ė���jg��,����,~|Y�R3�/Xv�KBŕ�?:薊/��M�?>�լt7mY��{�a?PH�?�*���&����y��$P갦B8yE����P��}w��Ap9̹��R\�] ���Y7�)���%��/�S-6s�/l���njni��	�^tG��M���½2�{=:�:EcY��!����E1�w��L4f.�C�ȴ�o8���n	�?K�|�co��.t�d;4�":c"����p%Ct�>�V��8\���t�zrz�=8�h�n`$�%Q�7nAx�zN�	³�aA���A�D�ӏpҨ��Y2U�khO��*�ݤ+ЄFҋk;��Ph�	k������Vk�)��XЋ����B�p�'eyW����d3>;
	����Q�=�x�%	�p�d��d6!�)TT�L��U��#��NǎX��!m(y@�v�]�Vyf8-~9]��%nP���˖5	Ŷr��mY��C�r^Qd5wA�J���̓O�����u'e-��[9�mz��qF�=ò� !�nCr�4��6�Јr([��X�
Q@r�QWv���h�>�O����a��>qm<���)��.��T+@��cZ0�C3�� �����f�f	}j��,�C���tu9����(��M�5<Z�	mTV+Ed��Ӫ��1O��	���0b��'n�'5Ԍ��]`(p5٤u-�X�e�؈t�JS�AM�
�&��j8l��oy�>$*�D���6���xJ�VՍ �er�C0��
Q0�gxOE��ǾB��y�}
PjS��<�`�J|����\ђ��ˢ�4%OU���$+�N�]qT����ñ1�0�hu0$���5��zr(�s�A}���U�!=�q��@�`���SM:jW!�e�g����E"��4g����S�N��IBe����>X-m�EY�Uþ����H�(�7�˫h���D����T�w����>�ur2y��K�c`�4��j���t�R��7�M��ԫɎ�8�hE���F�g�z{"�/��b�L�zj��
�ꗎ��ר�v>J�Bv���z��֠��e����Mnt�k�b�{�ڵD(?�@'͎��4��r/C}ݥP����3�U��[3�e/2��:6�0nTRX�R2T���-���~ujҝ=���u�(��u��3)�pR~܅�Zs(�iV�fۋ�w8����X�qt3;����|綧_�vi��3�n�C����*���"�Ӝ�>��eT�@� �kb!ɱ���0��!�8w7��u�<��Z}K��M$�����0z��ie�$q_b���)M�u'�H�r,eș#!®�(�d���!�ɛt�/�^k�����i)�s�AHNOH.��6��{Fa��dHݧ)cbZZЧ����n�Zϫ+��	��<�`�h�ID��9��4���-j��	�,'nD��t��S&��n�*Ea�+�rl>lsň\��d72*Ibʗ`�S�=�m�#��&y�!B�!�\e8G/��G�j5�V��ij���]+�8�}D��Q�<3�����݋�bŸ�i,|PI��i,�Z���]uY�a�3�����&0��WNZ|"�i��653
�Z��[�Q�Kx��D롌S7����~4����ᢙ�_�0��L���6�d��or$��f9un�	<ܴ�K}��[4�5Q��������u^�]\�]�j5�K�Q�6��Qߐ��nk��OO��l�.0s}�LɐX��h�h;�O��0�m���C��ך�P����|L�TBV�̾
E����1���4�l�����'U�9dw������qiԽ	n����;��IMTro�~6�)NK�������!3��+�@��y�!�
쩶��h�A����p�x�>)�>>�B���dO���q?t�9�7t,��Qmac��"�B�v��c]:/63;��7���^�a��L�]�N��u1r���I��9��]��h5d4SU�Ϯ��&��-Fϋ��#��i�Z�j���o���>t:����i�������O:��P�,4�U�E�F�cJ��#�,+�����mP'����.D�8�2�3��/bb���,�ѽT�$�����y`y�?ΐ*P �Н�<m�J����zO�Dq1�P�[��~<k���jp!��V\t�x>����hG��p�'��gD�d�6΋� ��b�~l�<#	1~�&���Vp����jx��+[��:�(t���+���W.�8f� ���B%UO�8��{!�(
�c`�|�*%�\����4��HLB(*N_l.��������PzP�%c���\d�(G���y
A� .�5�Ϩ
�����M��~�F�a0�Q^(���?Uqi>�ݍl�A���+��wp.��e�#T2!QP�L^GUW^����[	ǒ�
&�)K���??�Y����	�z;P�U|��#R�K�� �GZ�N��]���.rb��b�g��*#؊�z�"� �<NB���}��n��w�y�J��@뉺Nd[��/(F\B���r��O�J2��*��9(��8L5<s����q�Tq~ŮM4�,
"ou��m!\����1/װ`��S~r��4�I����������ҁE��_k&Ї2p�*ǄcȆ�we@$�?�ܙ�8����!K[c�u�$���%�,� �s,Օ%�.�ՆH��)h�Q�C��ȱv�+H@�$q�&���o���G�[�j#�Y k*�cXQ��Ķ�"���x��zsH��F�@��ĥt���.��,󐄷��� �0܇W��i���)�'��7׫;]�k>I��M;Qln�3�՗���nD�^,�B�s}�c���c�ܨ��y	��_��6UF�)��;=����EQ���h�{�!#��$Z*�:�Z�@�/0�/qpKa_o�c�
�����<����m���������}Ԣs^����T���/�QrZ^hp�?@��Z�P�Q(S�<�e�/^Y��+�sx�e#���Xc�Zv8Ű���$.0bn��W���	�O8�7�Z�f��<�'��١Iv=��ڒp��{m�`�Y|āz�B���"><p,~@�[���`�
q��o��[����M=Ϸ�Z�����T��us�"=�V�=�k�G�s̘�~�
�>���1�lt��]�R 7{���q��SHm]�p�_����zi�t����r��A��K>)�Ǽ	ˊ
9���>��[�z�o x�>o�
=q��.����J7��C�P:�>�:z�[��z���!%���G칢.��c���@��r�tvI� ��8��:Pt2|������aV��[�&aG��?<XP^ј�n3��C��Q
{N_訶k_r����R���6��8<7�83��*�i�i�L��.>ہ�F~�����S��?q�������ȍ�O:�DT	 i-ZV�$�}�hѤu�Y����Ŵ��Q;��(_c���M��l���1�%��F�k�
 ������k��^Gؽ�L3��:<t�6��0�9�*q���	����錆��V6q(M
	M�ZD^���dZ��@J���2�[?ii�����ؐK ��dZ|s̱Ps�s�$�8&@��q3srx�<hR�)o��7�_��nh�L��h�v! ���'�+xy��m��5$=�snC)�#^EL� j/���mI���!��Ї��������p�//lp��,Ƚ�X��[[��T�#��k����}�Ip�q����K�%�{3���-d�4��H��@�}8�H���c��"rH��4�����Ʊ��p�;�h��AfFb�0�=��r��ɮ�d�j�D-U���t�17���ʕ�=�������$�y��y�����W��]��$�[��!�u�N�����cR�A$�%�(\�y%�IUÐw
�8~���`O��8A��
��W��}�*9�f5�t�[��X���O�D$m_ҡ��ɧy�F�3���1�F1��`�*��i�l.ɔ7B��%D�U��a�+�h�/��v���2{�k�>,-�&���ҤT���<�� �b#�F��{�ۤ�qB��:�yZ)��˸�ړ �r��d���f�^mH��~���"s.rIc����r��mZ��Z��C�&��}���<�ƸT�M�:��g��G�����h�j8����U��9� ~B�"P����[�lv���^R<ŒE���s��|'���xkUw^Z����������{�v6=���h�ƑL $�E��o���ݕ�wBr<h�o�%YX\�"ǭ�Y\����1��{���H� &i�Aj5��#��,�O�8���D�Ȃ��n����o�t�V�r,�%.! `A���z����I8��َ���E���c���a�$�RZTEtO�k����i�t	���缀�{���Ǿ�)g�y������d��5&$�������QB]M�ED{e���um�5#ըa>F��`RQܪ��S�T��V*�B��]ɸ�^�( C����w�ۦ���ς-olV0� �*9f>W�˜\�B���B԰�|9��F@*)�8�`�6���6�#(Q��؃k�A�q�hv�����
��:f˕�t�����f�ĳ��@�#���3)ee�>;uXSFp=����;�yq�( �s`��.-=�����DRJ��Q�-jW��"V��Zc��rF��Y'�K�Wqmm����x6�qw�8B	3b��e��E��
Kv(�8qE5�j����+���(q�@��| t,&1��D���:� #����5�8���|��R3��u(��V��0V2�v� gXmoz��U�h���������8�$&�z�{��y�����
i
L9g�A\�����
���w7V?4����{{�u-j�K��'�+ugv��\�6�zG��߈!m麉%g���W�}�DW��D0�  ��uHRA_������#'o7cq�E������X��M}ذ���P��{*�A�/�^#O֕|�ީY�r�ul����X�<G>ā���(5D�+��j�Ctj���H��;�m7�vJ��|O�W�������Z#�)�HMM��,�5�H�{�Sk2���������l�{(���!�|��3���$v�!Q�,��f��7R���1�L�=�CӢ�`/��Ⱥ�������J�2s���̼dA�*�k���C�����"hK���v�F^��ݤW�M	��1a��]o�_�}<m������ʶ~��	y_[����M�� =�c(^�V�&���9<�О�I_Dr������'��g���M}ӽy1����GId\���r�ڐE̿��%��c��}N]�� N��6w/^�y�T�;w0d(-�N�
߁�u��X�i��>��ת�P|�实��]4���T��D��<b��lT�	_�r\9;���K˘Ό�.��� +��1�� �=Af�\W�T�h�T4t&	�g[�A@-*�G23��y[-�_��ߙ��+=���~K���� �ea��1_Aqz� �	�/�!��ʺ�2(c���v�MN�J��F}����Yו�&^�͇>�$Y���V���tD��t�:pz-4��*m���W����Q?����\}��V~���Eo+�I���53�J����yn�Pjp������S4�S_�M�Xj!�丯�*kYI��6f6��f��!"�C�d�r�������l�Htj�0:J��U���vߺ9h�ٞ���Ώy�ƍ39���-�o�G��˫������=��'sy3�%���`��-TPC��ç�G¥��T��EښX|� �����´�ix��y��:дK9��� 7�l�2�!���87H��J��Rk���yO�
�M�n�P2��(�h�q��� ���\g��S�9����~�Э����� �Ӆ���c�U E�Smtk��SVc��ل�U��fbc�����^�������F�	A��f^�?�a�����7R����Jz��\���\ǵW�:�Ut�{Æq���i�u�}[���R�c�iաW�#L"�<�.�`�"d�F���C������8�(BEŏō���dt� f�V��3/d���WB�?�T���p���������츖�/�G���ʌaa�����W�:�z��rO�}����A4�����Z�6�P���B���3�.Մ@E%I�Ppޥ�����bͫ��Z�E��[J��0Q>����;8� ���
T)f|���g,]��]а0��p[:�\T���hz�D���\	�s�8}��𼪙��ݝ�mj	
i���׃����kJ~�o$X9w"�7T �c�dEr3�h�J�ɮ���߈]ކ-(��O��Z��0��Pu
�!{�⠼�
C R�'�4QT.�r^�\�0�u��<7�~*�p�Jo/!�͚�o�|���7� �og��X��|�S�ٗ�z�f��0�L���=�(
o���<E�ٳ sZd	+�I�����T�P������yJ�@|f��JBD=V�oއ�����j/��[��$��U�����ZXVٝ�Aa��v���� �&��>��h��^�BAat�u	wC!�ITT#h��B�,�a�����gQ�@y���(������9v$��Cď�B��x���IN���Qkl�a�kL�?XK���<<��M.�����ۤب�7�ٲ���y�<���Tm�s2��H�OL��&�+��$��olRd��=s�e4�W��3gm��.|y��mB����� r�r�#]g��J'���7�(Ȁ�f�N��!�/�2���C+�/k�y�z�c�S<�VN��i�Y�݁�6�����S�,y�/*{�0����U��wR�o���`rI2��F�{֗B���l�&Z���5Q.���q��G4[�H�#L�rr+y�R���c��
�sNO5F�yGc]Ǡ���  �ozty;[1G�2x����X�ځ����s2-|�Q���Dz�R��F��g�U�s��FuM��%.An���N`ϡ=;�,[�׽�^�ȥ��:wQ����N��e�~���_bK6��5�1��/ 7�o����j(b�{c�ʧ��
^�z�Е!�dī�a���vf� ���/�*U�b_�>�b>�Qb�1�(/J�u��'�M�l!�!�SO��?1M+�['�$M���N�G��a��4�D��j��4N�C���?w�=����4�e,���eY��Y4�?�OF�����*��[ް����+�<�����/>G�����y�>J�!�;��`W��Z ��a�����hq��Na���8��'�^bJF2g*3z�]Ik��y	�gX�κg_mQV�����[%j(���'1��)�ᾙ������C�{H��W����M�n��.�G��V\7���C��f8Nw��J�yL֟����������������~`M>sU�@?��ʹ\r�//��3�r���\S�_�q�I�LU����^i4X�ы�J�Y�iU�����uДtr�ٙ�M01Ifm!�R��-&9���H]7���]�1V�6�q�";�J��)�c�R�/���鶴&�-��&�AM���Q���x��	�r���-u/66��(K�h�;�[�7^��m����e�T���#���e(�:Q4-n�9k�<�
�$ֻM]�ZO��ȣ\�	���&"{�)ҧ���r��n��T�7��������\~�~֘3�{���g����2��r�Gc?'(�y�s�z��+��K�L�n��ӪKa(]7��x���r?��#k����BMq��u����Lÿ~-0����NW<�V+'���'��N{˩�ah�,��`��O.�S	S ��Ա����4.{��TW���Fh�1O�`���0�)���v�����w>q�-»�+�}oL�2f�O8n4�Oxk�ñ�Pq��@�T���+���qd��5�:�ްz�%�+-y^!0����,P�:���Wڰ&������f���vY�M�o=D~+1����0A���k~Oʭq�r|��(��x�l�������f�T�iK���GWN����%���FN��l�s��QY��F��lTX�M#o|j{�8T]��*�����H�M�C&��C.�w�Hn"5:i��7U��<o�]�+�tZ�W�'_�4K�m�'_����bG���CfOHZ׹��t������*������d��鉆�eVzl{_��'l)��
I� ߁o���v�#1_�5va�`?uѮ�\(�&��	�E��ځf�ͼ��:Ow$��i[�Z���޳�@M�b�oi��+��fzO�)��RMG��K��V~�Kqۿn�����b��z�[����Ҍb%6� P�:�s�0���$�-1��IF�T��bj'�2>tJ��RrF��1����G���IF+>�m��Ih��:N<D���6�7� �k��f��9@��/���{X��� ��F�f��x�F�#�@s�/j�+S��n�7��)�Y>l�D�R���z��� �'���&ǭЇ�K��[��?5�U��G+�9�	����^~�T�#[�*�7��!�l�Q͛Nj�ZV����Y���!WOQ��b]��XɌӷՏ_ޓ�4�(I��\�G.��>V�O�:��i�B�k�h�SJc���R�V�ʗ�K��:� S��N$����!	C�(p�*�*�D���x�U���R|�����\.�1�f�)�Hk4"�Pjm�ϕ�e�MG�	�ٲ��7�&k�G��`�����	ެpe.>è��9��`�Jbؕ��U�l��=�;J��o������	�o��p�8R~��/�L		2�-�^o��i��D���1�l��󶭘�R����cL"e3�ۃ�L��*����mb�-vL�֓�Z�� ��dou����O�E�Wb�p��5��@��ض#�
���y��eU�����۔���-��Jv��/�9}xd�PuU`
ʶ_�mϻ�F�c�1=u�?�Eo���ۧ~;�7ȡ���ś����SHH)!ЋˑUևP�d�Go�.pG��ޮQ���󈠃e�tv�qvq��E}z��3aet@���h�R�ۇ�1�M%1+N*��� O�H\��K��n�aU?$�
u˶�v���pG���N��d�Z+Q!��Mr�?Dg[���u4}��N����3��?Eȋ�0,���V��_N� �G!���=�cq�P�s�V(����'~��>���K�j�M��S�#��;�>C96�{&C*(Nr����1l",2�P�������NV�*��t��`]*�zꇵUg��$%d�[�W �c`�1Ϡ�+���T9BsYZ{��R�~��Z���>��~�v+�)���%�~	
9���6��*��U�K�N���_���ҵ�j�sѾW���8�N�&�E�־�5(�$�w��R��F¾��}�nɿc@*�o/|�ڈ����� d­�-���Z�_E���-� �MD���2���W�I�I��.?��'�pJ>�;? ������1`�3Q񙴆��|M��Nf�� _sM�X�Z�m��S�/��@������#�M����^'/��� q�E6���~Ѭ�� Y��$1�	Ȅ�d*����{:^Ǒ�+��W-N?��4"��b�V!�gg
V3�2��o�V��k^I�t9��kSW�<�4� Ѿ����Yܰ0�<�����f��o�`cS�� �
e�
�
��)o�6��K�����gfp����Z��V\��<�\th
P�x���~6����D���-��/�U�[U:�{<�c��.Sv��1ns�'�4πj����]���^�Y�5/X+Q���Ѡ�p�q��ا�7��|+A���:q���E�mA�=-�S}��xi��'��� 6�^9L�g�y� �tG\���`���74�`���-W��1̧�J�Xc{f�b]�G:�l,��s�z��_��x��g+8� ��<,ۣ�j�	�^H��3�R�ޫ�Uo6�����`����ii�f9�v�C	�_e�}�������קs�w��%b��_S�/k���@?B������L��p �B����W} �HeZ� �#�!�ܚ�ێ�r��Ǐh���JM��D��j�ITS��Z7HZ�K����`�Ax�b�/�f�k���y6�������'����RSA�ZBE���"��BKcy�(���/4&�?Y��e��ty�B��5�v9��q-��� �)�at,����;�q��� ���^yf���������?.���|�*�G��1��a��~վo�8�� ����y;���r���O��)=4 s�0�^��l��h������2��H�+~(�Dj�6��pNA/g;��^�&�o�k֢�#zkw��;�A��%�a>��n>����'�̫(�r�%V��{�~��D�[��ȣ�uE�����������ߗ>��G���y6:CSw����%����F�rZ�S����g{oo��m���M���4��O��|�y�t���ŨJ��ՙ!���4Qb^�"��1	�v,qds��K�aᒫp|Z�Ǐ���+�c����8xk˵�N�&^��`�!�x���ؗ�0�%|!�!�Bѭt�A8P2�|B�2�����)\��[�=�<����HJ�Sw;O�]Q�KZ�)[l�)߮(��v$��D��"g�?:Ò�(ڣ�Y�,�=Y"��C���~��w�y��W-u���|i����1�`�-�g�����M1)g&IL�E�s#�<#$Cy��^)pJ�~�
�ی��7]E���<;c������67Θ-}��/�u� �HM#8wMs�|�HU)@���������.�:�q��P�"��?����o�XX�|h����.h�<ʧ`�0N��V�m�)�I��ˊ���!�wC�����~��y�1];x���-��
�E>��ڰ:G���/f��7�I�1��l��6#���!7��n�)(�I�N`�(��b6�q�ȳe��W#�9e:���A��q�e����xJ�b��a���O>�h�\�BkK���Ta�L�7"$�wǞ&$��_��=��O���bdw�au�i�I���q�$����
��!�����/s����ʢN��E����
~>�ڙv	b���d�H���%�5��$ϕv2=pڻ�椰ůQ6V[���S��=D����4���97�L�4�Ɯ�2��;y�.P��$
Tv�r���+-�^H�ߍn������u���)�Va۷F��Xlqh�ZRyGl�Ɋ��$�O&t`]�L" ,��u������o3p�Woz��XXP�^��H�����0m]`�}'o��{O�6C�P {��7��o���1������� �#K@;����Mw���}�w�d�g;T���F�eĆzft���G,E��3�Z���<�d�>&���iě�.|���ˏm����������5���p�Q��	�󆏏3��0��$�!�P���o0�	��j\�_�t�v�T�eg��/�����;l̜u��e�uD?yZl;�`���4����B��gb�����`���2�T��v�f����h].K������.�B�垸�N��&��U����>Y������� ��� R�t$�a�@�$������uVn��g�*���}U[dM�K��(�}
�!��A1�u�D+�m��7�t�08�;82T��Pe��9�[�4ɢ���I�Y]����tK���Q�l�!�M3�=���"�+�sa���f9�(��·O�Pֳ�,���r1}V��:Sƫ�7�J�'�
	�(��ݗ;W7i�ǪzY�.�%�_�4^�f�ΐ�O�&�i��(�����u�w���$)��^�m��P��?���(��@��;��ĎE�]�
(w[,���j��%v%i&�%%��@����Z⋺�����5��U.B�&^uXr 9���Q&FO����1DnL�m�=��y�{��q@��`eQ��[������4�u�(�	%d��\��~��-Ѧw:�j"^�=����C?�&��#��Ƒ%�x}3q2b~���9Qm��m�X7����� 2��`�lY�-~�i���<h%h�bL�h^34"۹�]t�!�.�D��wA-���ٕ���|�l���Z&<Jt��z�r%�Q����w�g8%|P�.N	lf3{��:��bc޹��v���>@��4�V��L��W戜���L0;�����-��C�TH�|hnMO:YN5�OC	dLU�f3�-S��w��/W@N[�ฒ�Q0/����<���z·H���2T�QGM8%b�0���>iS�9O]h�q�_y�+Q�j7S�#�㊑�\�
e3'��s.E�;�m��[��*%ŞF�b؂��Qٔ�T���>.��$[�<��?�������Gl폜JO����[>�o�5�:����A@$�;��ӭqo�
= u�}��Ա@��P4��I�������]4�1��`����֖�p�#�%R,g��͈5�ު�ğ��2�<�3���ϓ��01a����r+�.�ҕ���6"�1�1<Jx0�/kʙ���-66�M�X]F=<9<�����N���Ʊ>�=��݄�8���3�&�t�i��X���_Q�Jح	7�۱!�ue�u��W�g-��TF��eHv�r���<EB��Ξ��]!�Y�mVd� ��)�j<�FY�J�����+,��o�h-��Gy��= �>"�m֋��,��\�*����6��L��n4Du�p@FA�U��:��ި���i11*7z��GT2��NI8�,%I��f�+��aep b��2�c�G.�Z���$�B;(��}L���zNs?�_�o��=� �%�S�#�z����9��	K|���gen��a����%PkK�Pm���Pd�Ř��tT���Z1o�w�0Aj�a�-�Q>����05�� ���Z摣H"�WEL�̈�s���g��M#��h��z�u��*1u!L(\�Ќ�n���Ք�E�5��H����E���\ӭ��.��"�^
�Q���on�y�0���$�o��L�)��'/iJ֋�D��L�\�:�_�1�͕��Ά@�(.��u��.�c8+|Ͷ�P�P3v������t��B:Ո�SS�f:`F;�D�?��[4
|�Z�5Ae�c3i-$��@;}k
�=�]�DX��������z���多�c�A����K�/S��+�J9���V��CرKf����T ��u�§̰���s�k�_���SS<0)���WJ� 08\�j%����:���O@-f��h�5Gt�8�&!�?�nx����<X��b��2�����:��E��z�D+Ui�ꭶ��JJ�~RH,f]J���o�_�i��^mEg�3e��_�`�@hhkJ;o�+%7�������R�u*T���Q�t�%G�\�|��"�*겺�9j��a)�Z�����U��N[҆�l�]�����;KE�Ț'Tq(sF7����w�=�x&U`�R79�@�+��ճ�K���F�4���;^�q'������G�"���2��!zH��!���(�Hע"M��ߤ �tB!*Ѫ61�b�kPn�C��p���7�<M/���{P��q�?�z[�nJNa�d�׈�2u�Ihzj�J5bl�y}�R���^�� 7�U39n��5�&�G��w�R�q�(�E_v�Y����?br}�LX�ɇ�9H�x.�▥<��N�i��l���ʳ(��23-�����{r-t��Y�Z�Z@�f*k.:O4�M����u�q�D.�}��s���%x�aU�0^Ս��!���7 ;"���n���j�.5�� A�T�z�;�5@zY"���v����"�μ�{�t�q��߸aȔ����K�g���w�vJ"��aD�s���u=����� l�d��YA�+�B��R� ڃ��qK�(7�m5��!��͢S�$�m��d��jV�I.�JO�Bε�X*0�Kk���G�@@�����y^|�k��ٖ�SC�q�M�����2��t{�йȟ��z}�^iN:q\��"	���v�9hwiJ#�ϙƓ��8^;D���ү�A�%<�� �cG`{|�z�Tt|P�ŉ��`�SA¶� خ�9K+F�֟��h�`��b��|X����;��[@O�����&�����_��ϣxG�G�a�l��?���
�'����>d�=/�[���H�+��'f�tеl����/O���fBW�g]`�T?��;��b�Kx����fS� mLQ�U��|<^=�Iс�3�K��v�n��"Jܺ�F��6una�S�J���Έ�6%�k�[_��y� {bO�τ!�=�"}A.q������@����GS��-B:�>�|�G\���60͗�Mi}��g��������5-E���^aTĽ?�B���ür7��kC/�[���ed��Oi5ٰd`�gbC��*����:E'����)�2&2@��E����hE�R�F@��+��iB 狪��d�P�Պ� ���_�x�8�aO#D"xԵ9��OJ�uU�����$�6�o�g$)׸4�G���E��	q���	���:��d��n�8�U���4��	(R���-�z���BI�5�PQN�;����I����<-&�oQ�����'���T?-Y��N����.ɮj��O`�Q(kd8U����'�=i�6�B}�N 2���MUT"���.=(8��0�[�� ��N5}�<�"�gg��}�Kvr�����Ha4���f���p7�=��f�0v��cm(&��h���:m��N�͞3}���wL'R�iv��RHo��{�K!1ֺ\dY�W�M�;�0T��3U�-��7��KN��T�d���Az��n<��M����#�N�Fw/���N�BX�~|�[�=��l��A�So`J�fx��|�����2��:�<$�Eyǝ���4�$K�Ʉ���y� �"p(��p�:*��h�ͪ�{�-_eF��-��Y�r�U`+�{���<޾��_���Ou�}ޫ@��$�MF,�nr7��U~�X�+B%c��?)f�?e��e/��{��#�����Ox��;'Q߿u���ϱ	XK�XgS��!�-�l{��/�'�U���JB7M= ���|�T ��h��W�B:���{�(����5�L(�����1̸�_��x�IZ
P�uY���J)�g9w0p�wcּ^�㾡�����p��[���	g.�����v��RK(��Dp�C�8����"���V�[�:o���u�zyng��0̘��5��m�jG���y��4��-�m�c��Va�1�C�#��q򃸰��(��SNЫX���/m�a�\u5�[�X�:A6�l�+����s���<h�`\h{��0�B׸Њa`��	�����fr١ST�� $ �t!3�T@u��]�0�����(�B:�J���m��ꀈмs�3+xL�#�g���kx|1ߩ~��c�Բ3K��'5��!`�����=�]S�i	��i���^�ҜO.v�}���\Z��{F@҂q0�:Ob cٖ�?�k�,�[�2��\4�J�,]*jeF2�^(mai`S�l$��Ύ�d�y��1�@wA�g�&��,�/m��~��''��,w�v
���rS�K��é4�@J�K�fn Sda�h`��%�
0r��Z�A��I[�Z��
|H�7>�GO�u.Dz^�d�A�P�]ɳ�d��T����l* W��pj��G�*�F�K�tR�?1cl~XT���/�\x�@��Yp�g�+�Y�
�]:ɹ*�g�EhA��8��p�S�x�֭A,�.S�~\2���X_��_�E\Ҋ�h�b~�d䐐@�J�5���p/CQ�,i{+4*
���n�ug��mk�^;k�M��گy�l���ᮦ�x��Xj�8_�4�N2�R��,c��G������<� ����}�z�0���5���E]����ٗ�� x J9G
v��Ru#w����4�fnt!��p���N���n��Qdf����6�9������2j�~�z�]�����Qpa���"F�v}:�+Ji;$�6sˢ����%/�e`������H��>][�3��u����M�3��G~<:���a���KS�ƨ��<���S�/��J>H���Sɑ�Z3S0,����DNtv^�|��e��|�P�21b�%_��C��r-1���B o�s��sm��7�e /{/H��_a���V/)��ٶ�%#cJ��2(�?7��m>j�&��?/5���MA=x�m���I�U�+���G�|?7��#)O/����|���~�¯F=���Db�P�B d�˜�UU(1�}pI5��.~I�1�PB�&A+k��s����x����� ��އ+�A�]@*�׻��m�j1E�^�q2�v��]�w�ϕ����0s�x���j�y�3 �;۲Mssң��r����I{N$錱����5�G\"g�Q^Zd���\��i%����#c������g8���QeN�˨7��Ak��?�h��Xi�!�^��K�vme8T��-�[ցt�r(����vM�����Q����5O�fV:[�Z�ˀN3D�<�R-��A$� ��� N�Mي�������V�ǹEڼ���.��S{��G��ip��?��R2����$�Z����Ą�*P��
+d��ٰKq5�Js7�:��vt^���"�\"Зl܏��{KJ�q�hEN��b���Xv�I>(��j���f�,��Z�4x����u��ګ[}߈�l�!=����]�7w�R�z�۴;�a��������;�4(Ž2DG�G��i&���r=$�SnVz�1�Q�����+W���o��qB.���
 �����������<௠�O�'��5X��	{.��#�ӮF���?�����̻*(#�cX3����Ы�(}��譶��1�|.	���J�3��wX��ʉ�ahߑ���P0��R�l�up�����E�p9S�_�LGgϲZ=9�@<���C��ڵ?ee?��~�I�c�::jS�j3�{9�H57