-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
LlGPwgUvD6MhB7YNYjlX6qi74TWfzf1iw+mI0zHOVxRRuecTxHE4kndhHvJ3Xiq8Pq85kPij2AgO
ePsrYVjAMjdlYVEdPGOjiImUWVtvJcYOmEHvJfNPB+1tmcixKBLhDPG8A1LJ2XSP+3BgOV8h3698
sytxOwzp6QQ8pJoyZg+ciuFL0o4HBgW/MRAYwpwos2zl3qhDbnANCAAaFX5QR9R2mQj/Bk4LznoC
cUeP56LwHrB36CL2J10B8zd1RwBY1gAT8e3wHmOl+kXW1vzYCpTbnlgRnal7rnMPWQ8zYkxzX14x
r+eN0AHsrsASOnjy34QgiV3bMr1Ats3Tl22zcQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 9424)
`protect data_block
Sk0SkUho+JwM0h2rhubl4+y9nT1Bt3dop6F3toNQZQgQJIUn1KttVMBRoC53zi+5tvLuMDxJxz2P
Yj4ei+qD1nHHa3l59Zvp+QFTDzvnkIkoc4Y46lv93ZO8g1V+K4gszfp1B4Bq73rpg9dGVvfCw2a1
tb8A4XXfRmMIcTIVWRCf47vTet4d26liVfEYGQLwYFgc8vfKfPLvOBjkrTDA2E6JqGkQgu5QG7O/
bB7Htr0nnXN9I1zwpOr+W9AvNa7wlG/Duu6TGM4A5uGYAe6v0vfl0Ad52zfOWcN4k9nricwx4GOq
31JUl11S8OaV/ARPuiCHGnEHSOWCgqlUDVfRwRMH0Om/U8fPMS7wcLR5ucOP8Cj6x97/thtyfRlr
UxuiPAwZTdsZ4glUZIuS4IVdQvMGKig+KrP8WKGQnybxIJezVNa9+9rdTZUDW66q0GDfnxDGQeDg
+Nzap19Q7TP+2IhLJ3byDzYsbJF+CWvcVBmejnI+/wbsNG/EUtkl2y+AvlTrXRl9poN8WiaEngnt
D2wByl/6yUtGuEi7j0UzQ9Ln3X6ns7S/gyKW6fGH+dJTMfAYZkApAjOvRgM7fEx9t3KD543c0SDx
MyE+/TI/Myv/4ysr3mMCHENJYFaGKrJZaHtlQ3feEiNypeEPg6tju3KbCCnxRCNgQ07xvMuJ/80X
N4Da2+XPZnEiM6IZXc7dRM9S3VKERn1+zMmIwYNZQNYGrvZ5MUQfO5M3S+KUg22Nr7Dc31eQWE/L
6eRRx+JpWzofetR/v52bQoZKYmzP5rgYP+/uejQogemCeUrIMKScg8HOcTw786CWPOwkJKOF3Cc0
Cn8jB4dAqLSjO2GjCva8vqG6APzP6jXLn4rL+7vvD/NM1c2vQc6FRPOU746LRAzdrjuZNKQpmFFj
iha4zbiOcgSlfd8bCBT+csB24mah0YQtSqbDmtRcRVEkEbIntcV4qxLCw66z13lJlAVFZrolB8Bs
+gm1wF9zWIiEQI8vkQyZtY7Ua0dozHZwQy0ASjpE9XN+qC8psT7PciECRGsJlM8rZUy6d4eiEmS+
bwu7tIanrTChvMC2YOGGFRwDjTo0Vlwn2hbM/BRtZY4yuVGcsa9KrEQQ+/f+/YrodEw0pF6KlFaw
cF4EMb0SOFP0loVeMbXz0hCGmFbwji0oi4N5hmFttwvVYkV34ZsgCbRLKGJ6MVDjoV3R4Hl2ZP5r
9c0szD7oO7KFQIZ9veh+yMbRswnBZoRMEdVOoHYwOMnSsg4hX5Ri8K79tAaMBl2LwjkhmmO8Nuax
DxHCDV2sonoyYXGalourlbyn5f/RHh6Zy2uhTFS9PQh3Ke5l9W+UXTsrBDRss5P6O5eHdriZFgOD
GeniH94lwZQxKmpFRgsP77CNXxVXVg//1bFMbfVKq2aazCcrC826p9cV57seQY95edEjyWpCAhei
6adP7/8XPbVgQmLrUjPzEkGvBIpuncc4Enrj08oWruBrTMRTgYFsU2NacAO59aTj0HGaR80hj+l3
x9W4EKxlUUbSXv6H0lxh5vFGerEo8mqRHUF3cjZngReJNSD45l7MjHBCQDNPrBkIWo36EVSVbd/l
nF2cDuRFxu7wmbDf0GXDbphyhP/VcygBycJHE1Pxam0Z6MmfTg9h71aRCQowphF+iQpYUoeVAEPN
sAV4D5YQGmXoQOvOziTsFBLUQ458FdgEU1CskiIuH66EqNFmptbJNS9pAu3M5dwPf0Ftda5nP7/a
Q3Luu96srC7R/5XKpKE2GZn5AwdR/zJMqht1gDe1o0LrkKCBw3k/FVy97Q1Y+dMw2nxV7tES+ULh
fJlsnhhlJJVCIpNt3exDtabzJERREA8/xcTREItqT7vIAO+NZRSTm0KlQIfU4v5CiFFIbtf8WDfe
RlsCpGIjrH3SQnzSk9M/Cv0Xq+BSv0C8qr9d0++6BuKnBTFpRmA0NcY71qrsOd0zwBAMFI3GHo5M
XETcsQ/hOoUVYuBC1XNggH0BP9BAFD7SEgPnhrHe0wjTPf4QX2U0h/fNfxln/R0iJ63PZH7ACw5+
wFiXFLOtx7HNbn+/JfsM6Z/AiC3pUmhqC2PsTiznCDnCrRc5RI0whbguSyQ9rv3M3z9QwRaaQB/1
xU9aSSMbHbgutVE8sQYQQ89ShBdmGLljXSqZbt8d6NS67SKfV/BO0BLCE0qC4UJ0YdgfWRbgUVAK
P1ZpH5QXkS8pTorCWx6T315lbJDm0F79A+D0HftIe4FeOgJUBoPBRyxgTNqGpFhYnDFHJOSS22Mz
w7bTj3HY260SSOpQOVrs/yw8lbfyWWlW4wByrwoBIaK4KhvHp6OAP5bTHtC+T+Tnm27YwNvJ88Ll
KSsaj9JHN1Gj1X0HOmAzVBPAoOEwxnEMtQPxUDcJHJvTFCd2NS63L2Zomno5Mf2Og1LPXlUlugtf
haGfRLygqkOKYVwS4FBUMp1BKH8odgcezXJvffl6QKntmxl9eFQ+O1Wht+WDIU5JKD2CotqrAeB4
oCAde7qwry9R5LsR2Y1cLJCBC5vqcc7PlOCtZR4E8ecynQnLRb9sZLJMo+iRfsBhw63uzzxnXptx
LWalhv+ksgwP5oqR+TLJMfCWvThrPIs0ujN4hDcynXul9uZPj0CCndBtqW3VRj1KLqpJIZGVmXeb
NDo4Ws7UtJLzgLomRdaY4m3/0vOyh59aNahV8lgaoGJBtBssIPC9HsgO+yXzuRg81QXBwo0seOST
GJDvCKWi6JzKF2Q7hW7KaFVCN+3hhRNfwUPGEPPmpnwAHx4VkDQtRf8Z4JOSDhPeOtamYmgHc3sY
/lkk9pCuG2fLzuKiB2IA9YBLMrk4tNbR3LCb4hI0VUpnxovJVGJZWv30//1NTxLW0i0wbbeOkHJx
hx+k9dsxsGIMGRFpgjtRkGLbvX1wU6UkTqFYw791L8soV8AYGW3LWP9kyGIOKYAvodUnY/INr3TJ
kHOBDD4wmLtnpJ0/enb7o9QgCIrDpXZtlx/GH7tVU/bCCNEobmGj8UVwubZl4oLSgubf1wDT2dOv
E6AkJ9DIiYAT76EcwdPhyhaQEJtAicThCCFoITORMAIdk43IE0cQa+TN4Ydjz43NmJb1UHDhNm8W
AD/c2qKvYARZokewWiwbRO3OJnd7FdqbhaP5Q1jogWGTMl0+WHyEYNA3ZItrVtjYCBJypdfQ/frh
w3PdnyiBWEiqpAbbUCDe0oyko8P+1P2VCA/fqcano9AHnrg4WOKondhyzJVKn+TYA0g9cb+FZRdJ
PgA14JBFi9f4wyi6aswibOVRrbyxccNSXjElpQ5Nhy3vR/SUZw8GhkvHnB23CdbB39OAQz37B76k
Ugz80Fgc494NFAAaQGIE6xOdcpItIM3aOaz5ADI6Dducm40gexn6H3fEjeLDHsoEi12icMJFjfop
1F0Gfg/Nl1pZYA+iXkpVEFIoSEEabIrmdv0S7L7t4aAiP8R/bNaOL5upISRf/RiqQRnr7eqBn22Q
l0m9ppsWVSIR8Dwg9pQ2Zivx9i699Y4k3NRa9C9C88tUJtf9DMkT416Wi7ZRy6FIO9gXc0V0xiKD
fa2accWLiL23ihU+jRaoHtCFlIEz98S8AKAhSbJes8TCSz/fVRj/ScDDr42nti3F7B4PxWjLVXqU
eHM/CgDzlqUKNTsaYvAvrmw+mDDAaD3AMNof8B/6oD1igiNSilSx0bTyqA+ZP1Bv0Z86q5qwB1pV
LKxVulHmz0YkvPvgslY/ATJ6g1HykcIDZX9gncp4ySn2DGUzm3EL7rC16AxXqGUUdaMbsgEprGUA
xubPcVYnAv2F2eU2ut8u9066GZVmOSd7H4SoC0JYboedJk9ckhMCus1aUhAID9Dz5XvP+lwyqgi2
KAZOodZoV1CsPowi/gpnu2SJ0KCK/SqsbFWzCtzEKJBfzazJh8N3HZnY7UjT4K+8JRlLhActRpHV
1/T+VXw/onB1uc5NqNEP87lZF7/5R1MHDSujqaXWni7q1nxmJ8FkEObpiPceWLkTGTdNzLTUPghd
DnXKVFidhVlWBuin4B3xx3CvZYszn05c6XiWvwzAxIn1YBV1wJOP/xLIaKoh9eP4pzvG6ZOSASCN
2XXXJNQm8WI4/9qqkfaulBYw4vCHkUCUQyqlNuxXx6W2IXKM2my6sxVAxpChmjU4pPXZMztP9P3V
tmeVbSD7x2VCt2OqSfXuC/LiOp6/R1Gu2ylC49+nveFDt/KUCAZvJKtepnukjM5XZJLhVttgyo/a
Qh2bvgT7eFTjbVcIFifJBgdH7WOcUM2HP2wSYTWT+sIFx0ewAXIx5DqLhWyYSDIIFu6dxaNLtkj0
bBi/fmBv+9+iqAi58CaiempT825HaLzFZiIbClQ658btG19eyBacG0moWpwn67HTl1HrCPwTOuoT
sc0P1NBGPht0HZyAZMJ7h1WFXIRyVRGCwaRelERSuIZTm51gULeierfksbzxvSECJe67Yi/gqBl9
OdDKsKCC6Pz0cm/Mx0AuHKjxIR/YsuzbU6MMlGocn2LKWUfYNjhQSoyaFZnu0GpHoY1XXyEwr5Sa
pO7cOfzTcrU6ez6ZvZMswKPG2vMCVPpa/ybfbmRVK0avDPmiwX0CctAddskhAhlA9zHnkYn4wSF9
kTip5WOeJTodYkzAS2IQfDtyitnMTrxXAKJ40d2CRjyCutcWJJxzq6OUMG6VXwxlMK9/FkmNwwD6
t5HxW7tHr3yNQuafThLxR52Y+//PVw4QhFUIq8BTEEfunTRgglDQXJ+LQbhJmFEW3fWHQYOREWWm
MDgkRFOEAXkCc9zMh231KpDAy8xw3xSRlAAgJf3WhIZZ6+zgFb2u8w+imP7nCg/jtVfOFULu9+uq
7frklE+jwoc+fAHcFF6srzxg7myAwfkN6e+1uhqdYuzvXqmaGHh0DJ7MHaVnzpyCHIXRH05CkfXo
5KvMdzZB3ZWJ2P88sLmruWW/2zb9BavkKwqlYpjy1SlCGQEWH7UDj1HxbbuwQHCyCaNRSTE2mQkD
bUqChSv+VZbppv453dcZnlwJECmDOswCb+bA2UVa0XjiJLjZLOMKguWvluYp6Mdhnt54leFli/Be
7nZAuxvEWBcFOZXO1JBsIfxwmXmEK3+5BrkhivZUnaSGzIcI9bwZx/qTPMajapLGZmt2KEmlf7V7
hclek/3V7huJ5n0jJU1fmw0dimYJM3IguD3E1XPfIy6GLTonRWBnOeyy2x4UkY5iv0CxUO2BQGy2
VR0FOuRAdZBQnyQb7KLt+CUVOm5MQxUIFiqXJGga+WUndlYhaud31A3RmlqzAhoumuDrKugutKhR
0xLrdZp48v3kvqCVlA0MUNMAliL1m/UsemU4hJAw8n0mArljet9/WxvBd+ibfHMlQ3tqX+TEIDtK
AGIFamITeLh0hL+J1giwdWeiI76l5qH9TFSINIjQ3D/Xo8PFv2sxwmX6YxR/+7Pn4mOlU11VYbcg
hAz6ah22Av86b7vhHxHnuZR6/g7Uv60ztDfVUrhGBFytRoSUonQm22+ZGlnqpzlkdTdozqeQ9sFi
UQxDqAWDmxJLU2DUKmuDbgeyTm87sizy1wxfTWxg4ABh8k/3ukOIqJ1HUdM+Y66bX3ggKldnk2Rt
tSfhoJSMUsBo47V5a6PemLySfPhGWGEkkoNuHxbtNG/+nbp7nOZjexlnChIvcrkiOcofrCgRSDv3
NbsORxZaxn47o9xXb7mlJ+xB0/aqxlEEHgD/9JcfjhmBlfAq48YU6eNtlTZhbNsZr/WAj/LmKdwU
XVVN7SpquEyOfUzfyZIJfb/2zbe3A8kI/UCoMMz8/+Ar+kFRDaKtKexWmPmo9qOZRo0R0cOVktsb
5L8WwjDrpaq0EPxNLHpBbV+QPVedzM7uORWt7BRprse20BhYCQa6OL3AcWPROhbZAjnJmds5KTNU
4e3BBYbILIKdUHJ/G7y2Ve6FESwHLTE3EsN8jwF2NTbEadzSWWfn+hN3QyfT6/uDN2L4vbAv9aLM
gV/4iNO/NBbOAZrknR41LQp6900v0ltC0xzUeKz5yVfTA9efKiP9+pkZLyF7D1mMt7r/yTHRlN/0
vDp7k+V9djZZa47eY9xpMYBWXzeISms+jvMIq3ZmiqUekVxN9bAj+p9LZ+cISzmZ+FlSNlBrKj2S
Ain8n9yI9JN1126oDh6DqHhDl5KnBE1kVaGBP8ZYGwbrSE9TwiU3hvIYK6Ivh/9frag07T9eTFXv
IvrodnR7LJTMk9Y5eBbfnYVRXxVf20t39xwB/swvWOuYB/jwpYXLi/H66oguNegFcAFywG5/nDEF
xYwbiS99TqOP6PLWTk2Xt1Yf3aUeZpNhuJDhKdqhLzjF7UaoXoke4/FCP8IzhZ3Y2qQheHbNKdHL
jPvhWkq8oNnrFx9kcegq70qh22zhSAK0IFD5i4NOe03c10jthMhqW6bWHT3476rQ1N9Ea+HKsMPX
6szmQ3HT2IlAJ1d+TJN8w3uC7c9JCRawK7+n+38T4NNEdW6jJ3uXFG14qOeCREEu1LmGaeIOpGLw
EfRcvGEzbuFkP2Bhx+9Fvr+IMuWrctt6ghHYI28ZnDEdyxmpHxy8QutBpWWd38sWPpvYhuzr2G8f
e1UK6ir3hpBIicxvxEnTdZJGZU4vmXw4Zc8QFsyidYlVT0CSoITznssr5vZIzglGTd6wEOwbxOdO
Ood+olZ5SbeKMIzIUMBRwNtSY7qmseQSsYyQWffoXkVNf08spaqQCTYDrB2GWO8RpygmgEWIpHqk
EJdPQdqFtcaHHxCq9fNfm3lSpO5VoPzX9pmyHn5dfxJDGBuGnFu/0lapg9fmOZX7o/ADLN7fksXv
GUEgQg9ylDunwJeXom8YwP+gCt7uXBRY99TQJiItT2kUFUiUCJ1MRs9bDk1SvFI5+9+mg+6Vt1uk
MpGkystk8ZhKEO+dRaXdw8E37h6iXiVza8N+rcxM6DZb7/lWlTR8yHIawiZbuGu8VlD/p4Cvcjd2
pRW6Ry53GE2dkeeWBvndd5TLLvVsr73parPDIK42GSNXCg3BhHcwApFudKslY9n6BjJh4/p6SQtl
rmzfaT7pIv3734Nar0VoxNcvsUv9XXz6uIbYFpXmYA+0NnX8aJA3begeoLMUlYGzj1D16wZRHQY8
hhfKSuX4Xoob9Z/1B8UhGWtImQE1Gvh0D8EYxr8TnLUZB/YtuAIp6E64Vm9V6yIISsCxQzQQktaM
pDuVNfw6PuAxdjx/Vp+kGNIbBonLpYGrIbAu0RCn8I1qr7HI3zb/GoocO6y2ntGEwIhzANmTx7nw
zT87PZKe/E/gW6x9/KL8HqDGkNZqBdB12hSYxvuZMQmvFH6jdkxqWRkqrAmcPzXOazgnCIZDhz0q
Ti0Dhdo4o1jC90XsxCTa6nwUIVIEU5WG59fjgypjKHrfbRECEJYjv61Nfa16SFvB5oicb6oNKidy
LXpukBtOhgWy/VbetRzgxlUVA2F9OY6bIxdcXmE1vS1cPmsq1tEQ44r/9OAThP497gKVC3ZR6ojO
ucccjbtMHHUwpATF4AlxqXmxjS7lXC0rHDLwq1Ou27CxKc9uoXp3P/3C08NlzT5BDMO1vXIxRphb
x/avaBmvc5t9jPQfQHQzqqLeHJrPIDRWyTWs43N5/gjzblSB5kTLr9yflYzoYMIAC5VIZToO2wmO
FTATtdm6Nma58Mo/BPslNnUyGGdSHuqVhIm/fCJAqmzSKaLfta9m55NaRvYx5KNlaL8CYEUWtjcd
tK7sNr3PuZeKoCvHz1ZU+oMK3724tVflVa9sOb24PUzKwgqgClN/6ZX6t4GLR53U5Dslf29YAwgS
nGQjm7uyCsf77g+mbH77CefxzD8dqpS7K3oP/h03DJv60+aqtCIwgyJQmasWPjGHTI7k9r3D7Jpu
qlywV3ZYR2BAEUH1v7hhVmNQlOklebyN+P4C6ZmHXM28902RbaKlx7GKI6JZvoC1dUUOyIGhzMaY
DdMOfmxH2VzjWy8T+HNHkd1VOiwJrHxL7HbqAozyEmmXCJUhUhl9fv2BZXHt2RO+XzrJTc/L4eSc
5KVjCOw2jEfH3Q2xsazdTHB509NkcQzrEHAJGRQh0in9BBYRoymrcYTi6P+IyRHmUyl9ugnIDTID
0Po+vA08T6uwAZIX3RP+GnSHKHvsqtPdOoxHzVvObdZCJLcU5Y80mkDmGhfVa4eTHI1AewBPI7jH
k61DOYg4KtSuC/goI+31i4K8n/Uo3/mQ+NY75iF2ZOoJz5RYkj+clDmUMO3X7dxHwxc6JzAzb8A7
/1tX2SZJbMeUIqm5wTKXT5GKt1HG5e386DQ4zLAThchuooEUVjG2viXQdtyNkkmfu+7ZzUMn0rmu
bvF8Eu/jvZLZJu8+NoNXAiTdr24ZpV4856Pk0U4XwBIw/e0nGpDbl2FPYOCrIoLGZZ3BIUucyaIf
n1GilxB8RISGMMumq9Fs02CPAnYmrCKxi6kpkcRGu9TZHUnTAvjSkQdFD6Ik3F5SyCDRPz2Ytypz
AB4yCYL26L5HZW9Lc5oeufReFikPlfHIesjEH+rq4qXvImUnOZEL710g2JfDwNBTNWJYBfrWs8Ov
Yw9h4m2j/qrzF3BjwdrkhPnC+dNxFfJdukysvyEp2I3ysg3cAvsnhjVVWL9WnPe2W/rw3W3B+gur
yvn3vPZjj42YXmQ20Sy6cpm564K06jRvr+/edboE1QCOo7Vm0zUBQwfV/IhcKHzWeYj+JM4FlBU6
hqyoxMhtuLTUZpL/5XsTbIgzFtGCzp6lW3I6pf7soNaDSvUEc6qh1SFkneQANsKct5jzcwLG3D86
XOteUT/mLBi0FM0Dll0EillKI1CMjRkEzVgQVX9CHWITL6thnCd2aBmpeWC1bUkaG0HMy/esnMeO
gxShUGiDpOoJasmBR0zgxzE42Q5xXLMhjXvIAx35r/CxOtrg0TzWFwMVm9LqETOYfqLbyYWowwnK
seS8FSKU4grPpLz0t0ChRQ8stmBOv0S7clFwFx1g9vuR0oug38aGkHgjTpKqBLcRRZSK/uqK74V8
wsKX13W0pt8seThuPIMNq8Qgr8HVc0PndBYas10tpfZO2plZuEEmq7TeiTEZeMI6uwK4InYzbIk3
1c+48OLkK0wwX76l4wKyuMilv1TmzY0rZ7s8Wag+tn6H7T8fkxqOh5IECMSkj9fnqAR0rWRFZ97g
GAAYoql1mXlYgaD56Nvv1auQKHL703ZbYAh+pT5JPQP+BvrW77zDTiTsP28b2BggD5/iqgcvV5z0
BfWoqUkE0kqj+oRdGh+N1fOAzqHsoGJ1hHVUOPhdnSDMdIUQEiF4oXKVSL28EteoqLBDi2f52sqe
KTSdAFLmdSu/JxRkXxzoIBFBiHlKTl6tO0m9uKLmiQKioBDGsTDRQs57yppqA9x8gjmXVLKeM4sR
hwRTWumkKvgfdzJmy/bWJvOqb2rfZxOvZGSiw/e5DmkiwKnnpdZELf9EYjBD05NHB+cbRSADUq+m
kwwgwiZQY7og7pkl6hl4U1yFrE72JyY4+bW9QEu+jEJJTF89k1stx6EvgVKlM6ftQO842Wnx/kpJ
1puaDLJseUycwzXCznCbdLOOIV6HhfjqkqTcmmvmI4pDzFr0TbbtS4xuNBPY5MQqYcCQOP8e9+ET
ve7Idv+3LHb64SOjdSSzSmfSYis22forQA7sRkZ+ZsT4TYz7BDcHaDBYOlTx/65kXkNLlmHqmFGb
mv9/plq14XKoFA/UAfFog9ylZkW5Cn4ooLnAI8Ke1V5PplGS+CozgON2STcA764snVP2JrJdcqQ1
u7+j/wWRQ9v/GK/KKzss5DhHIOXOLKZyZTvzFMxrCXSm+vBpGM/oGgimdOdf4cICxlJqCnATlxq5
NZ/Ne7CioI6DX8HPoJhjazq2rg0rHUF9+TAXKka4EJwHyXg0xJ9fvCtrOwTY6VrlXBgNWs2ZicvD
yWOvO3keMjqODsOr1MZTZDxtFG+HF5Q5MnOfKpJS6lH9D1SPGTCJGrMxm+8/T9j/F3J6uES3WWTl
qbb17oSImz2PX2a1RdytdfF/14iLW14Qi/W10AaT4A4RbQDoayb6PH7BilDQk8muL/wbwef4Nybn
yjYYQA7lkkKUF9TC0jhLzUMr5iwKZa+QJYrasZg2ZomdJLoApMzJn6c3Np0QSgS1idnoQyPNyCf9
FFXag8ZpJYuWVibHRfYGzfJQM9Dh7nltOdk9RjTTTbyoW8EBozmQpoJTZYUZp5ew8ANZUStir0Ev
d9RAsmx6IgZF5WBeUe2850dri+1pgkYT8DqlLjhTnO486I8Ni9uepw8+YsnckSafNXsqBTH6aXtp
Z6S84qXHaXOAqqSIi0lbQcT4z9mDlBo5rdXAYSgh86wuV7d9ZQm/qI3u6xdEytigcWh4iwrFu9il
ewZn/rWnQHEtAHp4kJtd/zAuah1d/vZK3ZyFzsgyH7DVX6jVdL0l3zciduXhLq7kliNrxMJILMCT
lbLh1krynh7HvMwhgK8QgnixpQIz6/QEN0XGmv3lwgOZHMPkFhOw81JLbjdPGuRcLn3ah5z4aOuc
ejJgGiVS20DVz4CJezlaYe0XviaQBzWn2SWsvS+zELBqiVviB4/lIYwonceOj/ZKVr1bmlmpzWYN
7u9Q1JHVWM63OUmPZzzR7VqxSlcqsUvN5oa5ib/GqeVt3/C782r2cNcTNjvlNUe1vK3MFUrUakYq
6GTUXhgF1HF5vISvmhRqHynRZpLN0l98xguaPazhYcSKKcPa8CPe3l464o2/A0Pax832EC9dgI0j
YreZQ7jRF4eQBeAxvgbB8pagiTHKTpVnIwg7eGw6EJUtqvn29bCxchxGl7EYtVIRy8VPkGAenmwZ
jlR8fIzEFb81xKjFXU6r3wcFX+Hc6gi+n6W7OyDmohV/47XhEMw4IO8cLnxS9ROjUZdFrhEZbQ8Z
rMUi1hifUSRW1gL1QYlX8sbeKWKFvDUTdhukKqXuSwru1sRW4SVrR7cOU3xPHxTTGCIua+vs23vK
v3LAur6HW5aLTL6LFP/7TgLu0m2nZUiprB5BWBWNpdBfQk49892Giqi06Ins5fg9CnK0Lc9nfqgy
8uFJzShTUIsdTbG++/MpBOmd3tClIshbSiObn7FLu+BaOO5NjYTIMj388vFmW7LiSG46RjJmKU5t
75ye3Ffsz/sRKNHeFbpMpHzFPuTQ+eBgKXN4kW+YzRGVNaMBuuQr7XhZNMXSXScyrbnhXAHxl7GZ
PlLj4Vh7x8bSWScQ/5LHotrb69w8vzvxv5RSTltiorHKGV/pylhFng0QvfH7qdFIt8Yt3u2j8/u8
uDTjdDSkYkFmcnvaX64lqthK1KsdM5NBqdaYpFyY4pZi+1r2+Ngd3PYZOmRZ494x5uxCJABB/c1F
JneD2zTm83f9eKfODqm8/INDtSZvHbJItPmLIwt2R94PfCumhP5/y76you7s7GP8RSZMpbun54jp
jQb1SOIPZ78+Pnl5/EvmmM78s/lhSbKNUm9IDbh+9mU0qdVFjlbmaqOQrRXQLqgmOzo6RarmQ1fS
pc4ANuiVKhDkcIn8QpHQ/8KYBM/q3kpRaOLU38UceDyzsyeaejp/INZ6wcCcNdisePx0m4gawwTr
G5ZTUC4MTPOQCiS4mWz0+pOGwy5FoPqTPgIeAlxZFHuqEQxH/xIXJwMergH21HfGUdWSN4rQI6Lj
/t5GKFd3TcX5Pxb0w8YiQdM4WtJ/hEfPTEjzOS8XBwSLQOwiajjeMvBrgSm5M2JYpaNoifbK/UA+
61e3AwAog+KBAUE0X8shPAptOKfX+KOiksEaxuUaoSAdl70ZDLhzwlP3f5vEKfT3hamA1yP16jYn
6xqYitmMY5n5rN/wsDxH68PPQWH9b58vudvoIQjawRNSeevY/7Xl4MjRFMQFULvkF2SvMxe6LyIk
oZ4K3lzviPmRLtW8B/J5vdZff3ZhwqahNstQUhQSW+o2dG+ii1ZTHAYpqp062lCf8rPFo2KIdDWm
sLacROKyJmkHz9/n2AttOmxyWcegXtwJJEmGj5qUyDyR6eQK9f8QwnTLjvfmiPw3cVjmxldcS1b5
MCV4D0e/WWg+jyDHlYRLnwFs1uAfyzl22bH8toDw8hqSg1Im1nCUZ2fotR/cDF+oOOOTvpFtTM77
TxXIoPgSmke98fHYZpoRItfjfiaku19iX/zuEYR3483THOd9sUFKZJScf5rwEp755HbZ4+ytqT/m
tT1/T9LVvwiTBHRsYrWPDtTkU3jUcnSYTEoN5hUEJYs2Vq+FIs4DeZ6VkYECtX2L2MDjYCWACIay
ZeSndh4/lgdg8bowzE+Xb9XpQmCDvbrqOyjoDvlfMs2DD50h8JMHWSgI5HCl2666i+HSwYo3Q7mj
uaGQYK3r6uYw/M7niZe3DfhfkW/anmNYYVAA7eFxzt9O4Lx3YJr9vl/LIeTHlirJKWHZ0Nu8x7Yr
aiyxYAAzE3Gvc9YeW6DNnUcPt54ZcUhZF5SOGWYbJ36g71FbbdqHw4ajHFtelt16fJ7uUSuY6snr
w72VDpIAIgGF17ySZMzQDJ6LOA==
`protect end_protected
