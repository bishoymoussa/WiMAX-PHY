-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
XePqQlYKcckBlcH0sVk9VG/L/fW5zF8FszkcTYCpx7ZbozkZPEhTlilE10wGrkE3OhnlsnfwiQ4w
kX3lpf7umrK1bFu9iq1vRY8vA06OwW+Yu2rT82lfBNBNBK9rjBvLD+iZtNKc5L1EvUpMoBVRyhGl
BhM6ZkwvrSBKk57DW4LCcbNaQNgz66VCPDHliD5B1gUdVRRFTldQOVu/7HIrdcB+T7cY1WllaUFh
tAnn7hC+J5pHiXb6t/rok/O3i4zsPyP94YQUNk3YlnEpW9HgkG07qMugA9NZ5rCSVPLMdmp5buuL
d9YQa2fTf2giyeIPBZHLY4bT/ZFdj+hA87aHbA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 10608)
`protect data_block
+qtJpInrSqwJCT0mPpd49TovyIVG0fP4TvHRBGdJQdyWBoJSW3tfHsQBbKPgtmOsHJfxmCMt5k0D
vD9wpNlmLGe+jpBVzRufG8eNmYMo7jjJGQu9xuj3Sd+QvQaAaTqjIhsPYc9WFiGttj5W4aTU6uzu
9deTNyNghpV6a28q7//YroHIoZ/Szpv2QUoJ0O4DFfV191m/5qDzAWYtD3sEMSp0lnAppkoE9Hvc
FGfakZlNf9sE56Abq63qKXX54IZSV8ptMamas6FyrJU41HBRk6XwBd2EJHc3gTaKfEZZ5I1fxFWg
CcVkq2Em9mfzPbNacaETLW5T3A7rIHaeEyvdEODSkQ/iCelBWKReFKHiLqf9i9EDUcIdksXbHUCz
KgypSNG4xOa/YhuMMlJBcmeIzRdcJYPYjmZtBmb3iYf2LNujd75SDskSoSkObmgBTvtFQWUtzvsC
1fskNlIkVq1C+O8QPVGeQqZChk68m0zD7ELnIovHGr1lZGOx8mxTK0STqc9FPbJtVZvLjVoALrKF
KF4pBGDOuPrlEolQGagV8uX7RS4+PDNqoIBQ8cW+jqJ0RHFP7QPuw+QD+/6//vEHNQ6FWf07HEJn
Drdb96p/fXg4/Cqx2WXwPJ8s/xc/E7rNlFj8rOSfsZHLDchknp1CwB0spTzZ5qmHegKl2ln895ok
mPakP7+ZopUvuOmZPoF+CqowSqTtuYrQdIH5sbPuqmTJrnR0N3cT5iWDYYDCeNmxTYxmJ4/IwoCJ
i9z5EWpE9FX0jLGUAwb3AvI+m6JduzySUl4U9rDL6x0Xak1EUOrlFyt0SnsEQOdYK5f8R8fALQG+
sXwS2KvRcjLOOVpml3b2znI92IY7F1qLEml2QKCDtWd8wCsA+lAIvrJA2NcgxyzzGzci/Giowg38
iB3VET4h8DwWAxw70PQd1bU+rY+zazXbsVKqjNZdIJmSdM9efjQosWj8obDmZfE1vtCeLpUHVvdl
lOiO4Qjem70VOHG75dRv/O/DGclqliwhXJo1jj7fQWGpaMU/KNtMTmsPwj6xaHApl2h0Q3cnjuTA
dQRoncMH+MrIZxye/8/NFNZLCOVNWabgvFOdZDPAHgXtnUwuzBHAWZvppMuRo3RPCv+nAKcuEYJ5
posxHIO4zLUKjWObB76/JTjfhBVArDM7BPhzjt/6UWjBUWwTo7Fkmx0UN/vMH6IQGz3+PboXO731
nXRYhgeTqQi9xnSatAJI3kBLhXXtBgDs13w7ZOIElbvZ+Th8MBn3KQcbrtoD2re0Y2npBu0xsfdY
KEPqJv0FkEnnO2cI8JrtNr+pN1uXTU+BcxPsOCOQAeX1zOHddXH5xR9BZuD1asO3oAccclr0f729
B82bIJTuz39OhPZ1f/9P3bkZCofpz5ShgNdrVDUDWBLNMQXPW6LwmxIYcjUlieMsTUJcvlB0yskq
SteB+MjuqVJ3K935fpJxLXRmxF62Jqe80hRvT615Rm2WFzoxxSutFOo7da4/UzzVjt/ePp4b29ok
iFkYtfsiGjBK6eqgeCoqI8A/uP3EwZl3IH3qUxmMPHghfUKv86zbWgwXL8iGGpRnAjDazzNDGtXM
f/12AJRMsLlUqvSkwJ+aoZvOMRj8U2D371sl0C37BQcSZEiObVdMyyOwskLvDCkyW8NpwrzPMtiF
rLZDyG5SthLMdfPyjULacelzkpQL2knWFpE2q6E2qGF5oog39W0jeWqy/gO9jgr0bpVcOKk8Age9
qb72SGifFnm6RoYDMIToDIXSbMhrnWsIZaRLQg4/7/EgK1z5R/GSYfCYdSrOzffuq1ETTie4RwFk
1AXXFS04xLCDqBRdcj4MXWEBmNc7sCIirzKhndYqEwmPGI2i5qfl0Mn2e8onSRaCy6M+DpDCJzHP
pkYPSI3pt2fU3EeV45CRwfGXs1BvyJEOQsn2JLhxVoG0IKuNK84UCMHgiXO4SmeItlYBFGqXMnfx
/egNVwzfK0BvbpvUX2scCko2l5WuxZ5bzntKmJ6Hksh9ft3evkUp6x71Q85Hozxk7zmqwpiNMdop
FvVGeN6e6PHdr+Tjy5GydZsT4ZZbva8amH3AtyezIXRcMIIyR03dt1zSzbEdWagNCmhDJUwgPoAy
HkKBNd6VS0vvZNPrv2QGK5+JUDcDiMlvmWRCADcHaYCN2dg7kpXnUhsWMd9mlmV6hjXsKeIsrBa9
jTDdLva5LHRW1k/2x/Nif2HrB/dIt14SghaP889OMEKrkbW6d/R4kNssNs5L1+ZI8R+pyabwzC8+
rVPoIOQ0KU/I4ryojLrCbVk4sZpYFPMRIDuepcwUi+e8DwvXsmlITqY7KmThDxOlXS0utDcHUj+h
Kov75ZT46UW6U1s+OAmYdzLZpnUzYw2imCHVLo+f3qKPuZDiWsq1+k7NZ2lsZroJpaq9R3+S9Dob
SkT2Z3sb6JdYN6vmZaPlXiOGO5KCh/++yiPOphfDEDQw6SeanpfYBQmohbBCrW4VDPBMB0cCv9zz
gt36SOBrj3Ho7MAS99ijdEFrg/7roy87f8Jzn7+CgZJWl5WLzckFHk4pFAIcPd/7PoeYY85FjPuO
AxWcuNOkzdpvkVKuPdWyI1PkioX2csgdeb0+8g9UX5oX47ZkiDtOPXHiO/0MHOIp+r7KcXVncyxw
D6Ehr50Gyb6XWYk+sfR9FgwMVDMH01m0xNy/rNTLk0ffKuMPT832D57TZAevDaGgwbx+mQ3I+VqN
ABlSLl+gLE22XS21VAT05Ch5uwWjqRssq3Ki18N5n3yOej7RdeB8n5Bp2OKUEYM2aZSwmFI07PnX
QWpjQpBZNeTIxOlqE8p4UQynmeFJiibkSq7k2O3fvQPSVF1R3OKuTZMtF8hubKFbtz0d3xNc/1hU
mAZsFTFV4FEDYXPANOhZMTJ7elxvir6oqmUvR/opwCv5eNhRhCwYlwhQF/2djz/7VX+qMzpMIUfj
xS0LaBCDgHyA/RUW40QM2JNywkeb4NU+CQMLEhTYtQaeLME6qhzKuKotKrlBnsoQ2wh2dRiAlhuY
BqV5Jc4N2Rx/hYurc3PN5Ca5uA6WCPhzHFintXKwmCW2tFim9RkoZ+R+WYiNkm6M0grXprzI+Txs
esVGRcKFU0oH+IClur4ZNUPG9HDqlhzccA9y89NZZh5bnEKU1tbYytqUGJxy3usoGxtp3M8GE+VV
OTF6s9EKVXty/ePEsCztdQ+LDknKVefVKi6oPTDB8b3oLbe8ZKaCncAvHpWFMRQYcnBzDz436xTE
zzcYw3X5iZRVd22wbY9yEHwNHd0iyqxjD/7Xgr2ppA1qmTiSxHuTKlq3+LrCu2qIhKXNGrNOP9CF
8Po1qD/2viEjuvuR/8rrIbsahZJPQrpAG6OWR2vlKNY7uy5AlXAAOHxUOaCX8AZGYvDmC5KdBYXV
Vd1RHNo7s1WbLU3r315ZOL+OMTLNO/ToRZMoVwZfvaQ0whc5Wupd0+aGdTWv5YPNfoOIH22yz91B
RUrxC2dFHSl+TPNJV1m5dR+PggP1fR4lZGWfzB2MdNzlQEXIcV90v7qyH0Nsz8exjQhRwFER34L0
nFVF34+Tw6Xi3M1wicuzoYxA5yrD+SYVsCRVeyINr1chLr77AaMp6dXi7tKqsM+aGumPRKH1CTm5
mXabznMTHZaYlqi5cwnHI7kv6WLA1EXXhv1yuk/SLbEfEYTsjN54TUk8UJJF6r1qrZuqXCl/2st8
AF337pXoweGkt7BSRmY7L3tJ6ue6TmQJn+XRRPY4WU7nL5hkjY73o4A6Uj3QkT+Mc8ctqIbGyEyn
tUtdJMj96qPVRinuaxjD3rg6bNXGYGtj2i2m0H4mbQa2pmhPjJXo4o2a2x6dpSewcI2Divhhnyyh
lcEmRU7PQlz5t+J2ppBvkmLHFHX3izXBZUKpA2nxmq9PCcxQ70B5yhOqZWmysXq2zliBhuP3LvxB
zul/MBSTHzHlyYbDGCOMFUHrH9nrw1XAe53xFsLjVmXTseYXjalVTASBhN//gC6kiP33du+eAXWF
mvvnua0Xja88mwLHpLXeuD4TrbCpi6sH+yvj8oPu0dyGQ9eT0Oil7nx9r2jKQQVByEVkK79Cwuh3
56c2fa7PdJlZiJNxijEpMLUm5KdPNRuBZ894m2+nu2RggB+k8CamMoR9R+VZSbnuNAIUihN7yyLg
8xHjgEKOai3xnojDch7oNZAf8gbDI6GcDQJgi427DSa7G2YpWH2TJKdBqJbjL5Ga4Bl/hC1S/Nuo
yhmrjj6ZOfGo2AR/KC+M9hJXUj+bJPEPHealGfshEr35TzTEV+AkhYmbOiUljMaRgiyW89UlnyqC
Io7TAMvMz9ayN07k+3Zfq+PbRNPuAkUFfffvbQQT4O7jEaVMuSg4/suiMLYRUGg0SY+HdVl7NPzB
wyDVp7VpaavaAQq68B6EXSaJR9Cfdtjx3+fPzNhzhr9Yyn713+PB9N5acQi0140L5gSR6o0ZbmHx
io3eHhU0QYlfIUO6LiRjRU3FYrcRsvs3WmeYI9++ASZGEXFk7k7KxyveP3Z+zW+oWLmjqwGaUD8i
XUX7bGxC/KZprrQKuIRG45ey5/+PJoxbO/LbR70c+u5nxbtjYbxEyFpW/qmL8wZiDhS99jaf9nrL
IXqVHBVIRniEqhPdgeMz/DF0NZkhMaGgCVhQDHscyss50Ta6BdV2h1u4hSFBXC9+YpgbrXPzUq9n
RJ7H14Ca2JIUIyOrY+24rwRUOoSY2H+Y2Ay09SUu7vGfodreJ5HqEPDA4yA6yxvadDiCp4+DsBhj
VLmLirSP1P4FlweYzsIgEivIoSv4gXl9PafzfOCoOdPOPaboG4Nar5woSfW7zLviGrMz0QHbEJ+b
Y9Zud4YeQq+5rIRAI8bDBn4U2hkYTvplcXZxxogCQwlyLqLNmfciesVpxZ3aDdkDOMkQKay0NmOm
WINJgP3UwxNQsQfHrWz6V4TQ/t/5T8ZDb+jBhvYVxaOLqag2fJq9w84ltINkgAkfbEyV9SVsafGQ
uuKHiVSsl2JCD6Xzf5O5IHn8D1wT8LHKK3GKFrLeKrTKIikX50x6Asv3DaPwIlTC0cF/wnSjG5zn
dxDS4EdVMiK6b5mkLHK3WFHGf/v5a8fPEhWEf9LKd2dkylTdoXkuvi79/YUOYQ7iNPuN4Uu+73+a
yhuPV2FjVxLplo0FuzZZCumAozUSjnN4bm6Kjgv+ocReNwB1KC0htYUkMSPV06QcEBgBckUCtTO8
8lrLoAyV98bdtFVdKHCF1rHuUrXSA70TtuqKD7/XjVWxZ6bhaYa2KPq8Pv9EGJzB9IsqfMyA1sMk
c4EJTGHjLgqb8tl38hCiIzymUWbKavXfn6OPYdgZcnM9FoOQgRhd2zFdW5Okgo3gC9FVCTXdr/8E
d4iwNliT5svKudg7dTFlTIz0m4j2E/GakC8BPO13qQ6xX8tS4TgutfF3o/OZOkMikbwsH93uJi2r
GM82COHToiqI4oP0on7X5MIXvGSYlI9fiE/BBp/c2HzOwDc433zMZFKW3QDbeyEn+TYQ0tTaSM7I
ttN4y9t89LXligd6aYB3vh4I1Mg5wm/tUu3SvMIEg1bCZ2rSobOQbxlA5efH+3yNB9tuw+vJn+b/
xEQua6ABPYanZv1zjjEz/2XK4DtzPJaq5RiRMwYiq4/kOzPYUGMEdztwwQgQ9S3stP16ujNv/eDK
oJOhZMEhMzY1JCuEaVRbVLwFjj7FSobt28O1A3JvJt8CiRqNjlUQpNn64PTu594lUnVJ8bLm+Rx7
qKCQ+QWWv/hKae9vVEouWhwm26fFDXcs7QWqgrib0Ni4LREzyoswDy9IClpQ2Yffon8pnR/51/H3
h7Xhe4fS02AmcAf8JmHvXIban9DpxK5fw4X92J7kDXxjjGXnkk1cPlyAwaTzWRdDcQV0gzfqzhEf
xGA7vOFX5LM7TeYuKWISUSCEEooXRDoi0kSS6Byo76K3aEhWXv7v3cAJOLiyMpwz1Zyn7m0gbAOl
otm7Tp+AF1WGTUkJYIhFWPyJ8FG41/+Ouf5KY4QJMRb6TBwzIcxRJh3AuH7OnbFDg5EkGYkaUHMU
nG5Y1D7GHM3i/4ehh7MmfxlEw0Vz2aDgrRr/XGbSWaMOMkZ5/m30vES643a4yaaAcTeeWGhHWMAA
C3i/C2GgpId7PXMbMebMvUq8JY3Q+GgWVSeL1GPtMLC+yzfY4BpYt0nCgaWxsoB6iSlkNTQCuQ8R
9dhH2bvt+LG82m4GNYa3rHrzcUfrZ4GzUuudBqurMrPKv4QS4FvjjiYEJc2t4LHsmF094YSnEodU
6roEmPCCkWwsivIhwtwIlV2BzA9PXxVKEXqH0+kjh6chrOJojuWinZydlK6y0X2SszUZCMUmQVWv
jAg7/wcJYVGrK09XErNcqNrjFDJ4pHsnc36aQZgqsEV5o0gipLKXws29wUW4iZVtdStdNSaslNwZ
+w1ERypzvML6YNVSGxyOI7fSaiOHj/pj1ZlY+Ea2Dxfq1gZESSKWfQeOdV8VXY3i9747Po+WtNZJ
7DDh6G7l2wJWIXlfuvYpq58CVxjBhE5JoyMjDqo2OTaVXYxOlRoJ2JGpWEt2A3FK1m2gcGBUWTpk
H68kE9x1M66DGW96eHRb1YEc4aFgigq5cY8gDBY9d2G1z7w3xINFMcrCnvWtU804kNfRUjo1DzB9
nx9fzw6goEELC2aA2VLodqrC7fo6GIyE4aqzuqf3GYIwY/2h+TAQCUgOM48pvqwlqQx/qifOwUAN
FO4EheYDBVUyfK67NzOrDWLNhqhXofg6CQO+pph5DV81QvYMgK/pY8dTuZCvYTOY4N6ZWlAeANB2
+qdzbBRjnt+7vOYATU8+pPGuwWfCFh5dYWgRSqmdbHD5woJsxBRi7rmBBuW0mdaTvTCnLqvKby3P
JhnpDO/0X9btzQpJvtJKIRSmeEO81osuWLGw2MOZSJKkpa47pU0mA5Yfdb1pHiofNm28JKXnMvxn
8Od2b8liRfzNw2KWJmsvCLZeueEAju4N1zAlcMKsGXFb79wTwF7dA/pL6NAcGnJLgZDBOa+hI4g8
KNj6mzMiEQEA4R9h6lfca/2hfYSHy9b8A2EaRnEOk5JTFhufE9EZFrWGHYz9b/21D0XE6jc89R+Z
6ryHF6OlvF2IL/7EJZmaQmxYTe/Sm5LQsQ0rFDnIBKjE3IFDhq6iISDynkShk8vgPFG/jvCehplJ
CO10xMAxMKBYpxZjdAAPRMET/H2Vtg7B5vsAPph5Y54wfvNKIt+RNLWi6m6mS1o8nFK6IkmLaFmd
jjB8XFJ1bVAAIK3XSRHtjMfvemN6C3Oj1vogHf7MArdrF9pLYhyYta0v9XKYQCc3fNHb5qDIIZuG
gOID5jnuW/tOQPDPoQP6VM1JlDcunFBQ7wCwzokfv61f2vyK6MOi2MauWEXBuPWHHdBQSIRQYdca
uhvQm6ib77s8/fNrcBl1W2AlxNx0/CE/5uVwNmxCjV0oKp1Ps9uKBSkZmvThAtETSWF1H5UU2kW2
rgKsqTja3Xer2qwQvIgYikMyLceNL7ZMQ6HR9p1LmJtsH1lVd9+H/Jnvix7g1fnhpp+L5GLQw29q
67qKmghqQ83bRms+rDfzXBmC43G73hq4gZ3V2/4FCNvAHvLOzqXjuTW3NpK5w0SULcOkvO1gMf3e
Q42or3lQXpZpw3cAxMYfIiLdsjsmx5tKiY5AfpxHP4ruSXqcdZszzYSYwoqg4YZG3BRS4CrujU+g
gIdDzxy37QTyOaK9C4Q1AXWdhQvHtH17KIZFkJ93GYlu2ZOCdsuO+C0tVg6tswhpiY1DwmXnevXK
K7385EM0/cuDY2tlp76ULcGhf/NkoXOVAgK3ZH9bfxEBQdJvgO9+Yyg0FAqntDJjcnb2eBFT8o8Q
e6EpI+boCf/uS99w0kVex2kxUVtp9BSFyRa2OOmPx3e01TRR5F3ytwmRL3j4NhM5qxMMVap8nVsI
WCs/rctBK2RmGPJSYqU9YfAoiNV9RM/W+uYARIrV1bxomFeq67fVUR3lEm9ZlhlCH8rBqo7YVtaP
PtphUW4+EthRSVpSdvEM5urqiOYJlj8JlXO0CkscvAUni272cULl5WaFu0oppdVufrYjB15yEEnd
Ufu8eE4bb9bG/r4acBwM6QfZUKLRWuEmWijq0F9LsngEqIvd7stZ1btwh8Gc87R6ZxsDBItgNfhW
yQLvEAn2Fyp5SIowQqAwDgPSoKfroUY4H5FY22d99R73woFWUCyAmbpr/JRH9OB3zx15WmUyoi2+
dAMJoOECQZd/DlUTmlgS3ia71m6xH+cUHTk96hrii4ffO1z817j7gbYtpbP9obNHOiRqTJ5G0+Jp
pp5AavgXpsGpOyRIlYd+SoSm6GsTY+X+EFORqFheiOSCATDbqbWAgKy0kqMOF45OJEVRYWZ5g5bm
Mrl27P8ShgGXMXwPDTBydLTuuLUt1lp17s7SKIXyZqqgyfUKfTFMPtN29DLD85xnTbgfju2a6dbv
ZNwLt/tD7k4674fOqNq5onWGCntGsonex7kIss0F5QZVnHgkBvIKc2lhrOsV8jBrJnm8xKdDFdDq
DoEMTKYc+2RPk5WB5fT0SNaxNJlm0v962cI3CtPZ1X/Tf5mAQAV4hawhFRcdOaUOdJUjrltxWgmy
ovnJlxj04wHlmW527/xUCvA4cHDHBd0Lk/3DFXoHcqa4HrPJsQXgZDWKk0Z3h82RcAm8x7xAGQcr
Clqd+Z5UM5BqSCGlOQvAeH+Oqqw1CrfwSWuA8kxNJTYkOKYkUgXoe7fMIx9dHW/ap8lv/E2miMz/
vaQRlzR/7/RhZPGpyLBjsAQIAkPQ9ZaXYysXwG8BFR+cWCxKkl7GasMTcM7+IMNUXWEVCUxlF2YB
4gkg+mT5Vm7BFin4tE7UQOao9XKg4lb0jVBVun5J5ZMa2rtezfD/KQX3e/2wGOD2RLQGStkZoQhU
0Td1PHsDHQzs/0cRh6rbif7SoY9tXVLlUrA0TebDU6NF9SKzssFs8CPYOWpuGZgv1Gi40Cv6QTfM
KexG+nsFhi5Egavw+Zx6bndFtP7z227ssNt3/6QMxXMS3yeqaFJbRPcfbUqVueUx8McQtnJFO/Pu
2QJMmvK3R/ra/YU1lLM+Q/nw7ZlC9eY3qrc7XpnqT58FCIkT2EWmfiJmJbCfWmEF8+G0jTEg6R2V
4Re46KsYHjFBd2wX4w44tH5p5lEXiqfoYw8cHepsNJ0aL8jAhbQ7ZrMdXwiOWwTHmyZQnbNljk1a
7xcZDPQH3g9bCBS1KoWzg9QKysLZq9LkRliSCJxXh+QcwEGcW+eFKM3MfiKM6ekxVZVPKEUfzZSn
V3RIEDwbsCjaxJU1YTNpaMd5N+Ux+9Js0hIpnbs9PVfuPq6o2brnkRrrnM6pZjSSYIK5cUgqGZMO
IBrxgkDxCf0zrgyL2lQkpQISLbW/XeiWdFADDwOMWM/uOw30lLmIAz3auJzCww6MaeCxWw3OGY82
0nSuYLl25YwrZKj9DmkB2OQ+9x/yjamRBMKHQKz+yq+jdgE0jmoqp03ClXr0XB2JkYqqg2IxFPFS
yVOGENbgByFI6KOfAXZBV4WvobZ2shu5X6iHPIg09E5NMPxwDW1FZPBDNwmyHAdcrjTC1wIWPhS+
uUvFjVqk//vgPtsZbmJ9XdRT8mldbFiYdswCoxi+k4aFzbfk64KGIGwPcwHP2roI8TzgiUQ6w4A2
KLdg2+LBSM3KQCkcsnQPjsZWlJ39JojtXH/RrFBaW4Bb6eEGvyTOlGt2r0fM80odYGbW7bOOODJ/
1B+FE7EDCAacay8XATXWpc/5oA+m3Lq35Gz0VJiXUIVCBKR/eqC4Z2rr7hY0KL1y5pbzfFEt/BN0
UWeQl6iWPVq1EAG2KZWcqiEZyJTvf3s2iWyelpAsVwhGMxaN5lr2u5TLsK8P8pd2BSN99PoONlqW
Ezn1mqfjEydUYaW1EpjyXRqmNcWukAyYUjeCylZhXlXHMCeGjGaxpdyMpBeHeqZjdnZKKnLTu5fl
jma8yABPaowFojil+Z92zFKnOrlYGsErVatzbRAGMvX0SbGZakUABvEBNXCAj3ypStfGPjEOx9wY
RWb/lIU0pI0Z6KTYzNgBR7oFb+GhGjQHUL2H9t826rnMdZimQYwDy0cYFyRzug7XUPXo2zR0DQN3
MJ52murZ/SVfjSvRjEqUlRPrpTO08roMm/W4/R/XzqNSu1Hsv8V7hAKGduMUbhnDNXiasOfdLRew
dbIphzQ18WXNzPyBgliaygw/TwsAeyqCCboJmSf1klTfs1oCCbfXHYfoJhJWIQ3Cc9RKFu7QN67d
Gch3FL9T96Dm2fPQLlzhQ6Wwuw3+mj+ozkSeWggTJl+7V9zGLz0byPV1+PDqzIa/p//pfpYHfNCG
u/NpzO7G0RLkqYDotTu63jN5+i9zNO8aqh+9gFImnf15DIYKbHwogHIMwGNmpwyyhKeEVSIr0JfN
/CAJQZx9gmb/0YtPd6ruNZNrT5Pcrg9zUj0UEozazOiqfoLLSSaEfLZpqxGXxQzf2xXOqaK2kRXb
RDJ3txgncD99wnx3BlFPtvjmbh2x4WMtlwK3la8YCH+hcDCjSGhGz7NrOHpBCxXCzyXyVHkT6/LL
aauyVmlN3NQpAlV4PZGAMc+hdujWGQOv3dJCiLCn8X3z09HYFWPRdLTAXxNGRXAl95txLKRmAOEO
N5i7GhuMQqyySSO6xE1mN1MT1pI/HNUieFaM2X0shP9shxYvwlz6OeNCznj3LTXAjebvY3Za0BAi
jPDG3xEMM3bupBwjst1z0FoAzF9VhWQt0GEPokkuYFacUg3xLVSoksHx8x2HdRxEEp+mWxk/DoZr
du943Nva/jKr2sV0lfjCRk5wxg9YjbWJDLKARTKWxfjAGtE8OUssHliJIDImbelwqcyjumNtXML0
URPDoWeTw5rMo3zj0VCCdQHmx3IRt2XaVCmM4XaAFe5cstZfa7Wn9UZaT/3k+NJLePDeyCEQYUi/
t0nlFPiDfhlDtbo+S1xlhLGdqNSVH4Oqq9pwmyLEkpoIgwA+QKQoP/UzNHK20iKCnKYZi+q44Ai9
qzMysq4GC+GfMjnMdy9aBk4rguO3VSAE8ID0MaijvqczaBKVFgpnV/eyADln/k5KxXGmYNDMgbhw
JaGB4d6o2HirtGlNONQ/t6FZ0Kx/FviqwXaiNlqLMxnZonF2ETJu9QiMsHoDpM/5upjZSZTX2EZX
Uco/rPSWIccYiilNrqZ09eBIyP4ELWcXxk6Aoi6kYO4MjAz5vUYTTgjeR0iNh7L3Lz3EMgy5V013
KK5AW7qGOWkeJOPoX+sdL/3M7BoLze6BfQPgOICQC7wwZ78z2OZ0ReMUk1aB4gJXxmutiAX4xA5b
ZUBSfOR10PnhZEyo/cjvsQ1D18U52e1pzBOYXa4sQOX3ET0uAI5JS01pZ8zUslvD69PtRggFvVQh
wAdJmvmZYgZ8CjQ5rnv/2jnIuwC/7c3f6aWEMHD0f5WChYktx2oB/whyHNX4n+IlMGpYHRHdF5sf
o6fa+aXaR2Gt8Bs8T41zqhNZ0x2iD/cDNCoW9JKvDpmWdnxKq171kWArhQ5RURmZo8CIaznmUeBF
UwFC77yOXnXXS1so3KmilUpGxyaw9hCNE3UYQBa/TFSAAlVtWu8Y4HrE+E1lovD1gOnfdeiDTX0G
ZkUI6dOBWlCm5N5lVkBlAIGBC6NMWV9HmBZv6CMaPBKAhGsayZKXk5EE8VtRq0JnLIr65nJcFJIV
vSxwIvWklxlCB9A2YwsGE6VfVSkoMVtlYwqQNwm9kqkpGigHS+UCWUbcIq08tTRC1sjxT2XzA137
YPIy/hVco7/NBWttGeTi7k6TUDduYvsUsW/HfCJB+dn0W1pQe5cHt/6n5A1wkcIieo2x1NBoW9ry
0GqlPf5gYB6dYRWKmU5hRysWa2WL/xN7ndH8dy1HCnTiN0wb/8tNO69sV5fiJPYYeFKW9Z+M6mT2
AaLcoPT/GKXKM9CFPrTnT0E5p6M/f9AYxXaSM/GVNsXF8YFZN2TuXADpHXdJqhhQel29y4Xkd6ks
3wff66+OpbYS4ctAafksBzUJJR0HM5HeYO2EgMAAz90aBzt0CokuqEpWw99QL0O+y0Ez+4E3I9E+
rZAm9ly5ZfPHYMgEGZqQbZa1KHkEET+jzU3Bta/+YRk0rkiThzrFw1zzt/j4dbpW4f6aTl+1NZRF
M94TQSwpST7G5zz5cOIt/wMyVmdzEL0DbB5XXwQbI5c6+0wceBK+8RfbJx1HDOX37S3+hhbXFhYC
uetc5eH7LC8IRCpNaa8raTTdpefI14L27qqDWYOD0szZjJwYEKU3NchXzS2tyaSBljGoqS8ZN6uc
v/yeV8e+S+8QQ1aHAwG2j9NjhN+qnk0LNq4/VyYNJbGQCQ0Hv5j0how1jnveFLyiOOy5BUVuGl72
v1QUfNcMAyyV+tuLF8EeXEw9mlbpKMWEetyaxx00a3oVGZLYJUguExEnDNIwmenIV/K2OFWA2TE6
krapxLJIhTPtHEDCHemFtEeQ84JSQY98NQB1Rix2vExaJFO/tAW19p8bZNY5yWBDPY7R3qhNY2RM
tKCTOGW8gSgHtA5D7vNo2me8dOsLQPl0vhtHxaSb/kTiltM8AKy7NxJ7LbBStYeA5Xiym9LqJrp3
GQecld2+4r7NeIWVMePHQ2NgEy8BlbABocA09ti16vfH4tZ3xT2mCbk/oSPPadVH79lXhb6uScOA
uKH/5P9nI6eLLAUp5r3+lDyIFXX4XGAwvHe4pbElY/xYdKUHaDTQ6VYDbFdEgFLOwzM42gLIosCc
wh2r2J3ptTpaFw7RJGZk0e99datjwp1g8o3O3j0dgOuhDh07/C3Io3tO8GIuz/SXGUtMrosJDsGH
e3doaMhCrwi63Jq6aFhEBzJKJQACy2unv4TBSsvuPrsKqC6T7UGIYBpy4vwiTm7tra2U9NuxH159
vVL3cZxmbrS1HQTRC/LxYV3JlVCOczW8Cq6o7rl1a+0BmdwxMw/29M8qhAb30ugYS/T/dw6tkG4j
FHCKYG4rnEYLjPSpXDO2Vz7iDHns0Q8kXcSdVCVMrKqsUgdV/UsJ56lKQc6ot1v8n+iLDGjJckEe
e2Aqx1EVmj9/T6Q9wXOveDCzPQc6HIjXWYRiy1vHSBG4QNMAk0NkwaifWmW8ebqG7+x3fXzS2nCT
nGB2sB4PACFELlQmDm+Ul3FduweeQ46auYsFDVDh0hlQPCFiXp91QiARPc8p8yWAbTG2KJsCo4P4
D+hmoKqvdQZvRspmVBDCp9fgBKVBn348MdcV9N0JlizMjDmFULn2iU/EIyzDKLtOWjI+w7gRhKQ6
qkrmcBTJnFWAJld0muK4YzUcNKJYUUXifSszeNyKaAgBCMfTZS/ngbdmiPklugJtvT/p9PhCUjc1
O3I7JNL6rU9WbuPDsLyE/ylIRoHgj0x/719JykXHtbQbyk0VrY1I3lRHhW5PMGphbhDrxUkbkElt
phhYDifbO6Zv0ofYKUrzQ1E2zKkX1PAtJ8WtQPqekzPZHPm94g2wg+cvahAIotQLnsOAPZIDAoK4
IJStamijiBKg7ZmEp/pLDogro6TQzsM0edGcB+rjHb60+Sy7WEKvyR8i1UFtBglpNxSwsrWZuByA
Me/XVS31CFHg56/u70zuSgan2nKQ7D4BZpU7XMqZwGEjfIwb4AQS6nTOYT9EO3a3kAcVlg5Q+1f1
zY2bOn9JShRUirdukXXxi4SYNZPTwnCt46aSnWEpbD+xujR0MYHbEqSjYQYzaod5mriE9Gx8j57Q
bu3cDJPU1mCg998VcFVCSch9QjmnxunZb1P+oTg1hxIV74MnkL4dqO0ZLBVsHhuQefa370wFq3HF
Ai45jAQtMBcHOmedt5KcBKYgwDCDJtL+D5ElSMb/l9zDn1l1MoKFCX89wHjZRALVgnckb5NCu722
wII2Zny+OxdreTTf18TqwhCdmuWVXu2Aighk5HOAc+hhv19pbeNwryzgg3XWTEEG1WvEsWmbCzR9
zj2wlSuMCz5J25b5v8gCq+STvLOL8iy3t4h8PqSn+EcOKYuU5DaWmQnOAHi6tOZUoXeBzH7tsxn1
GxS45XQt
`protect end_protected
