-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
tBCFgZK41jJGnVaqxFTXvaWiJ6q4ToUEIz8dtGJbiKYi1fzIOYxm9IJA8VK438agCTP9kcZsrnUM
yW/E36EbBJo5N8Pw0u0WwbD6aNbyPHR4DS9LRCHWUQHMtgtfy1LyJEK4IqA+VxQUMRvpdj9VJ7TH
9/417UmLfqgzC3WSEkG+3tIGDSPYfEAJkH5sAmG2GZeyprAeUj32CxERg5SqOn/WX6UoNW+EMc3G
VDtGWiCnH4d7sJmB8cBcbF8Xr5TvFXNfiADrY3RcKe3mf8qXMwllTYD4dm80d3333gRu7uu+2hKy
1ZOS2AbTb6OshvUm2861UIJ45sH1tN0VjSWm4A==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 35184)
`protect data_block
8yT+MU5f0zTAc8Gwt9LY91JtSR1ogaE75LeO6hmzvvCoJR4pofXPYAoOd9Vv9Ig6XGZq+NeOocYb
HBNo4HfSJus3XmhmdiAQPpODw4yWlqi/gqN0QqsF63sTTx8SQU44aVytEj3Jm3I0hH2Es+2qE/tc
1/zgw6Cp62j8ofDXaN8Z1oivdFnYxUTqCKGAsUbWzg4uqSopW+PzurA45XFUm9C3UnA3NK0J9RRB
/ZxwO3MGRI17Sp8GZDppDmj0/rg8s4D3LXJSIIqRvFuA1ecHoKykf1sZDzzhtMrzh2rAUW1u/jyx
cht+SwLPrcfKbMA0prUmTOzH6dSbWDXUmqv4JasjQMFuC0oc/qRSG0G5UPA1LchTmg2aaPFplRrI
tmxcr3ZJ4v7WyeZz27Dljt8PrPeeNxKj/hPATxBT6owXF6TgDIuIV+2GdfxDABDHvPtfE/Pv4uLm
PLOZWLNRghEykeo5Pwrjkg/AMA6uIzp1sNDsljZknaWQJMCH/D7vYcMp6xKKQhbAJqEeRemgk1no
yP6W5o2ZYXAJhF/T4FqCC9HOHoSZTkBbGZo0DdLcql8INMbuk8una0Q/B0H0LqNhC1L4/uzcC/Kk
FZ5ik6EPn8x204gnViBLFM3eRUGJU8Wm8aGwJvo4AN9u1W/LyEqV4Zk7yylrV+nX8TW9+/8IH74G
MnqWnIOO7NuvcRDdLkeJxdbVLxBJhw3QBw4ze8G2gyHuHwDxMnl9Xm+HlYgZMEypFiNN+dLtSny+
+D5tPlxYn0RYK37nLfL2Y2MNlySjG48qQCGc7Lz2TxQPppg/7JEoAuUdN7qtVS1LsxHlzkPj5rLj
n+0VxX4/LV/vuDPENkltWQXriojvwx+Rj+JNP8d0TvbtFSmyN+rSth6IjUFDBKemgBPoWL+DKbdX
ZcwwCkun3d1keED+D2PYf+iliE1NZodV52CZ02vvw9TAkAkhj94bDivQjYYsSOtQH6CVv5lzlcye
cNVckFMEmPtCw1YMSRFEMV9/SIJgL2lfJnqsS5Tf92zyhFq48mvBWQmokXQNn+ecp5+vHfyLp1m6
PZJ6Guxzwq7y4ne2AmceC/ILiL+jZm87Mwgiwj5Kye5YN0FHwE1k2lWCcxo7YHs8n4R0fJ7UvvMT
eda+rpLkK9DMSB1oh4ldslNNyHlqE5v7ajCAox63zbz9ydzvideIPD/qJf92GiSLskWUmha7EsTJ
oaBI/zaplMSFbclQwPblGY1A25AeBSJQztdcH9gyzPhvrZ6iG9GbVcOberoun1qLZXOunGPTXNG7
egtqtRz96xeZbRNdSNlWoWU9jPqD6fYHlxB7rSdnCYwy51wCLsFnL0WMNjbfRgbNpjJJSf0MMBpU
/u24oLIMZlkVOVeTlpjPjORzI3RuhqzQXq6bJXtNIKsYpvH7ciZhCsjIWOhk46JFk1gi8bT/J6US
MkgwIv3oRe0+kfbDrx3NCbjx+ingco+B3dqIbs3WUdJB3tkxXqLb7z0VaAMbm12oOawdah+MYTP+
C98F1UkWGo/jbP10+BbKFjal4zIf06GPq0A+DIfGIVC3dF29akGvbOE+KX4Ecz86fHXdSVEXsL6m
UoeM/up+6HEevIeMta3+kncqhmvW8mHuLyIsXFCJPAaCdm7YnDCh6PlorxZqIz3nMe51JSeknXvJ
Yu+Ie5dkQSlZo6SGEJCnI2LzgU68qQblDQtt/VCmBiwaiLu6+6D7vZg+ou9TahqESiLM4Tubqe3F
e9K4xraUdIpJdKKXV29mnONgQUTaOA3aIQLP4PnTSXRPYXFVkZE4mj0l5bJlReLiTvPb1hId9Vi3
mflB3RQ7zabVhJfLpG+qd7bO7UP1bSjjuRN5puXIlTv/xaeLST5mEkvoHyhCm2nbD/RgxeD+lPht
ePpo3PdL5GlwAxrl64VoQdSHwiEC0FvDQGRmmXA4HhpXZ+xPogEBMJw6RvfREu2Nvcx0785PObFx
NP8AV0tppz5jXhQFNLj09fcjfqiUR44753DsEuJc0X55QurfznziEm9zO6ATi+HNAnEyYGUnU5iq
+Hgqlda5FmIGfu6dx7y8gq6W1IYhmBk2dpxHYgAfWJgN1a5Ecb+FmHcj4uvcZ03Bx9s9ExDp8+ND
uVxiInNFn0eNctP7m6+ZCZAoh5kyTSn0cILYfNwnxSpu5wBijVJNatXjyuBxEEnQCb3H2q7zEp7P
OOdMQ+Gh9SV3HeqRRMIpukKm5i6SN726sN3hzZ6L/+MeSZqngKfov0Me0ZzS+wPN9Aff4wxaPao4
LYVgM952gBL9oSpNAE95ILqJ0WLk1xCmVDWDbKPJeHSk6cmH3rAGQXBoJ8JpVMDosltLN1dBcrfu
Oy4HS7L6tHEsvF8sWRkLeBh9/zC452i5xCwBBtW5OppdTRTFtaNZTpP5PHuuCE6P9DqMmS1Fq1bm
w3WeI2PahFyV44uFKUvjzCertORhuPQUfmRW57tV9VikRdEoEBTUdtmEen6RoUlRpjgAGVYw3ehc
C37n+aJCqj4mgbIwCFSLLmJNU7UuBHy7l74XBrBmCJNk0rC03YD5snRWPavzXdQ1J91M3FOM6loI
VotXnIykt14LcuIRn1UNJyw61/3yW6Rr64ECueV527CNBG3xGjwXcisHXUyOjedXMTrHZlnSFkgB
R5XEE99n07HRl1py1vF2w4+nHgBwSC4BPmNuDUFN/8+GwM315+ISyqBT1rnaD5FvdafBEqPSzWnX
Rkp5kupOo6rWh7jUjUvInipTYDI2ZbmMzdEPHpTwt8VbdZF9nDDSup2oWdW2y2IdLl7DgvoXpDH9
jkCreA/nKdMEGdqlX3LO4yGHgCYv07nZRSWKBVxY+g7S/75Q0aoXM0OH8TkvrZtlXeS0rM8rshKb
lJK7hnpjxenOO2iscdwKoW+jyaaKSGqNTNWUxYEUgy9aKOWFcLhmab4Crxcq5aLjnb35yrz5qnAF
v+0awutKnHIAlBqOLwln59oprVL5mqhxJryXv0Xtj1ey8rag7on3ixgKhzInOGBMoMEk+ceV2nhA
wjqU8/dcf6hxtbyOR8UiV+AoCXsGivij1kihq/i9nOhEjGfM7NIhgvqp2Zp6WRIlbdkPJkJ3gik6
nph+zmxXUCx/KlPHC8dY7b9VIydWZgke9Doy6RAHzUcWECM2didCq2aninHQikJ/O4/LlXSNYlJf
hb5iJs+xBZtSjQJWR47U0PKE3x4YWzQjI2OLf9zQ8XpbhgtD8rOZ8FnB+/jy972uSrKVtuZV+tyx
5Zx86CmhKlJPDs7cbOw58ggQr3CUHOYPRir2qj1ImoQcDY9yIECOaw6BHwd86dc+thQoI92q6/3E
YW4KrjA9pcUVFENwwqXXMXWR8I2ynIOGQKhEihHAJBd0tyVA7hT/xIN/kmd2XGqceFaUyUVSrUk5
yYNZEdceh33Ovcmjn08gIbKcvBcMc1Px2EQXpzG9yjJF2o5MMpcndTfITnmTtoRiBd2l8rZY/h1h
MgPGKpfNP5p9i8RaAorNmCoXTtbxiw3uCrqktSA9jabi28f3EK5CQIpC+BBtktxzvmDgVoHdsN+5
+ycQ/7p06uIyxf010QeOgSg/tyMqfYdheh+8IEEgxpzMh43t13y1dUurorzrJq9/14LCGHnlW/3R
eC47hhy0h1KKttZU3hOrtbLe0qoDDBQWti9tUV03v/e2d8KPBOZxz9dSUM8D1wuDfo2cVMrvtALo
Y+eWxKAlcCVZOjkCqmjFn3l9rBFVs9zqhyJdrqyMv9DFt9zIqyRjfA1+CIZXXtcZBipV+EUMy1d8
VPpRG7B5IBAIjMZL8o1tUXQB5C5OZjXx+5ajE8fwgib8xbBp2ZaLecWchjTtW2UxSvCT7sKyC1co
IW8fXaoCoW7J1iVP2e1FPmPfQPkOOj5yzii6WuVpb7SrFTTHkI9e520yXTJSMnXjBWp4IswJA9JG
S7o0h8H/DhMyapopBkPG49Tvbh3KfMhhXinT3P7okEzdZIJyVye6ZbtA/wcTgZ2OwKs6TRwKResM
laMj8Q180rnH2ITE6kH6C4tM2t4IfyMgUVl2kP6nQN/jgUikfxRfURrnb0DPhgrCIswHeXeNVHI2
3ghwkGIW1jDZoL+ZG4kv/kh4Fq8mL2ma+rR3d2cuKkyGFk72h/wrDdsKvCzPs6J0oLJ7Pmh5v7Jt
g4eUdTP4Nn5VOT1Fqmvo65aaDOCIcr+o1KeA9pTkTuoZLju6hNtco8mjlqjDkhYfqL4Wu+SGjcfZ
e9pkEeZPqtNTll6cy1fwNKImlkc1job9F9Aphtedhye9H0K0vSfN1lxM+Nq6IvghpcOIDGKuStkp
eHuCKBCC5dDLmvjO6YmWLH+AvJdy3xRJZV0ZxhN/L24oqnKGxapOFA+XvzJrKkdzx2wqbgabP9vI
Pq7D91gu6Gv4paVcwOhumM8mMKgaxpg+NtT/Aux4gRClqbkSEJVWi6PVyEiaWgLH3HyKYDHkxkJc
AN5H65g1+kVeAj0OT3CKztDffPKsg1FnHX74bgymQBo8KL+XfZNzzasGJ3doFFRgIO9H7PqrG8iZ
1nuqyKW43noD2tFQEM4KUtLuT8xntNTOYrM1HyZIzfMUbDESN4cGgqHYKME4DbQDTnMJid1OR8IO
qdme7Wn5Hc5AE+XWrclXEBg42d+DQhuqWNyIMUR9tK3wGR7nqzYEG5y0WeWr+eiHdSDeBBfoXMj/
AZMBFAhH2/3p5EZ35hKFeMUNTR5kMQnMGOm5buDNf2E02aRSs3COutp0qGJ4D7Y6Tq458h7i+J3g
EKcWC5mNxoEc7jevSh8oxdNeIKw8vUCJDJqm/AM8g2I5eQ8skxURJb6JrNWdj27tCtutlBHexNtH
7cffOieWTwixX3MqHe9utSChnqBloLsvTp6ouPwjmklW4/EiU+R+6P9osSvBeJ+P0C9sMzIVs1T/
hyeO0O2nO/3iEITCYXQKvlPSpW3u1e0C3jnz3FTArRHHbrkBAGpaH5D+L1cT5bRIjuzl8Vo6IaCl
IpKXEVB9zGcMojUfkY6tpjyG1qU3D8ScPErPNcp3Via5wMrY8xcdxH3E0US9qqObg7O7ufZSGrw5
3nJHtUnVvWeguhxdz78/QPkgQ2bcu8tpXA2d2KVLv2UOHX4n7DwT06sS4EUMpAcE0T5xkuatZWMR
aNSxSmcVh5/ojIoolTvwpDEsbcUDDMxM3pb6ueZYzvOVYX/IoQU0G1wEVGN7Cw1IguewudwoePAL
J7U6cMVCFeiVhhw8Si+rvCDHjtbeTDJzE/cP8wsBIRACa1HINi+TuVnHBjsLyJ7pRjiey3VrlBNq
eJQbHNxsXRL6IUcyIX8EL91Q7cfCGNrGYRxg8NamiZ2uFmVotQFiV9VceqYDqcPcHjTpYJVgBRff
dGJQ8qsZ7b6FgiIVJ1oQTbOQ7FwIQao4dW7ldxoEtXioTicjr21rWSE6kKPAJvYTZewZwikK+0OI
fK6itG9aHpVkUlTLNNTiqSNBt/HFutTzNlYWnsr6YQi0wo42FqEsPurjujE/NTh4tRDfmU3fpSVN
pkU8jaLrcjHPb0i4qWoKAPZEJtUraRtEQenzq2fgcehvIXSF2gx5AGnjqyyGnmC+i1auhuFk12u0
fJy3HEyaGD6uNhsmDhxqpgOi95H9e5UjWbNDfXd18bxp5TLXNQW6leyCA+swMFmmOCJA9GEBNbE2
xL6zEMSd1/QQqz4ql3bCsrq2yYd6o75pCPbnptNyl+MZEzwi8hhR0EP5Ti9BFeO9dRmh5I6TcF84
GT+Mcu17QhiyyhmpLCssebzP7w5Wq4GdUIbZ6DKueuNsesKvf93lWIeigiN4FyD1fLnHIpuaJZ5F
2DFUqlhff5wiHswN1W1bDzIAo7Mna2vlAPMzRxCa9afWogj8so/MDhxQAvblfh9+bywEYw63dybC
6U1dYSr58AIwJbUBYoKRmP5cGlVDrOI4OOKVHctb3oajfdCTiV5wvlcdh9eytUNQzhzaMWGrq6wD
li5I/VJw5JrZZhZVw8UBd/cnFxiuOkt5h68/8hp4oYsAt1hRazPL4+IxBk9YfsnaVwL9++onoWc/
2A+AFwZNhXiZ9FYx7wNnoa8R2w5A0Ah2P8+mUa82KsWt/ZIbBidqy5OoP1G+Vt3kE5ECwqEvHP+M
yhpDUpyrF0WnS4bkxa7P967lc51uydqjNRTsf0vvzqqrWvq8dA5T60B4ZOEnz9rPNIJN2CX0K5Dz
6hDhIrG7vYQu2NOpqRCpvWvVzoMvUncPdptin0XDIj3fhGcHEgORYAZcBzmuruOUO3ybcm8p0pTH
LOl/n+dH/41sgmZnfqHc8CJSntgRduLPURFMfi3og4MRJMrvxEj3/dbai7NO49YyhozR7isYmN1f
eM8KZE9KP4eza79OfBtxbEi4/UsnuafTjUxH3bjf5lJFPGWAqo2YvSDqKdY48xWAXXMmN228TUlm
zxtBMqvfh9StNy1QSqJBdu3ZgBFfW9wt65IXAn9vIMXlpGWAuKK1cXSGrbGJrPi2o43n+OdKJw6O
4/2jMqGdk1lfcvlv++hzarr+5E8pUXMQMQUvl9MFhuMvEMmHaOJlKRnOJrx1HitT7+8c0ynv0bYP
aFMT0gl8A3fbs8yzBvBSzf4jfrPYOcdn6JQGQWy/3wP+KQjnb0MN7jyUBXREGnVUyU15z7msKLaa
Q+ynA9ezIeoReqBnkPo1R+j9Cqv0urTSshLuYq3qZ9TE/nLj067kzXtE1AmaGVndoFfn0Ln/IXJ1
0hN1DfEU+Qp3P+CLHU9jekLQUnPsN3Sig02NUcxKm9jBF128rjp1PMAUsKfUS9+rIv4Kt2dkzKpf
GiyqoIevoI2ff4VDtPsnGsK3WF8ZRLAfEcWj6G/D3pW4vZp5reatBBCps4iw+kh62rYZnEn/etdQ
feSETsnBs7mA0NaKNHsb/wUBQ8DMuHoB2tWF3A3iONX0wMho99YK+SZhBNw02GbtGqREMKVcYMoG
H84GY+E1C3VFNwCD4kJhvYDifHEHFiCvgpkU6HaBQGtxrAo2w+oC4f4JsXDXNn+PgA0MEKYtRbIl
N4X1onEtqD67oAxk0mmdFKAmUkLrGB1mEV+xVpJcv6vz5/qX1BhHU2a8kT3yxDKnkvT5cE/1XRoh
Ed/LAOQ59nlbRJpDfM7WfUoNA9ttIbAVrPCnhWu57gSNYpbHQquWwe5vukBxYGyMMKsFhrBPxvww
xG0Ai6JUBC2URhziFEDaIfwmq2Z2qkOGfVHuc5ZYvkgTEZJQbp7Wj8BCsCHCXQaltUiuy5ReSpax
+SveDVELuCN9fZdZ8r+/3kPlWN+5x/RmOhOkNTbhElN98ibzGDfje5zuwBKhdasGkLoDfXnrWMqR
3AM2JnYdvubHqrzCzBGkbNx8crrjxtWaIlf2B5XWGp9VFqiescXgfWUCtxwNVx+4Q+ZYBT+Oop4x
Am6D9x8hRQ/Rm+oy5WtBaB0xROnEb8tCTDCzLdzYs/hHmP3lHtwi2yNE7n9nFXHloj/NMfEHCE2P
N16SoE75XwsF59B3d+3KMXQ1OlD7x0AZ5IaXly+x370WDs6fTMxKhTG/2z8nL3YuNdRRUxvPIAH9
8h2ojrK0lBdKg84oPYwpXm8i3aeIj0NSSBg1hC8mmcrayvl12TcSqfpxcARxDErtBTS8ApBDeN1z
Y5ydwKUDk+/qdr2EYwmFZ/oh+C6j0IQV+6vdEUKvKi/fssF4Wy2MSLg/ZlEk7Vxolgrm5eRVlK/m
0nBaK3RymCVH/9etwB5nLHgFzCVq8AHp0P5n/MuO8H/ZdEygzFAokIqqQglO100kiLIla8GYicVx
pPrfa4+mraryCdlVdp1EHqdFy6z159oAYg2UPET5r6PG+N/E29HmVWai104LYj129q5ktaQqAuaB
qDIY1D4lhJn81ZUSeHidWsUoH3qNLRuOc5ynCJk0OzGwdaNp7UkwKn0JZiGifzIEslTeDF2sp0wm
RZP1Je9f2W0k+MYx/ZwARa80x4Kz2A0tRcE9fyUG81APwuKhsUeQmuKLsNelZRlJafuin0PM3zX8
Zkytz/7co3Rc0859sPX6MZvDMiJ9P5X6xAhrF+XTsAxUOkdOax2W9ljuzuGo5VcrZPv4C1ZxVsWa
T2Nqte9iSFeDLPod4P9ODxhwegVFda5oJVoC6kZajH1DCmYtXPTrGoLm4zhqgl686GjSxdVbHfkQ
aixbYkAEBec1d8sXXtiaenZpIJbCXfcKdq4qOfmqzOIbISFWSBBFjwQiwXT1nXsS4hL7c9fAKO3z
EBbxUISOUseZzeXMH29sdnwDYvfIF+XZEWVWasundRPfGhGKwlHkNFrEUoV657wuPib2c1h9HXBk
jkxN3RM4KUQAsz6ern37qZNE61ML6NrTR9EBta7M931en7+v32JvmNUJ8f9yIMV/seSKPk6VrxL/
W4zxLOTkimWWKm7k0DNgOPMxbrLD5pKXJs3XcHaW63Z/s/Vqpr1IVzSJAedHbpC3IhqszX53QsVB
9ICgCNb850EHdOZVAehMLQjCX73u5bNeofAcNY7mflImEWGfuXoeyh/nXfW83m7tYU51DUntqdl1
yBON5HvtmHp9x8p8F/aJjLBKjk6oXvDhKOM7fJHE+XnwDOvMu93pmtZ9unC7zq7O0IIm79IPU6Ye
I75jXdmyHVmVruYKoCjDZQ9+d8rWibwinXwJUSIdu/+2SsyL71Mlm0vjPg4qU42aDTnLKnDz2BRv
s2R2Mv6ylauemMfY3ii56wpz0jj7GGTJVAKuabfYdQQzvd2t29OWd/FDd+4FXff8DfnkMPvnFP1j
q46kf77QK8F/1x5JWvGl7t0oBStdNpRzCmqE4JzkIc3Zoggw8TPCFk+qcB6rUxPZJGflfqvXyDHh
KMPqVUCcgDJ4r/xDRMIIDX1xcjFTIBItXiYyhZn70FIlW2JZRAtDjecn0MTVIBp1SgiOfxKqA9iJ
BVDy5FF6K3mQu7QKqAV6tuMbahoJb0+kUVjzj9s2fdfVhA5oYSSVBpfsrKvPJeuCdPffd8vTW6dW
iTiC9DrsRvmUGAn3aGzhk1WoSwK8xNwb7uplifSk8HIuu0KiiZyhsZbthAsyoqkVhtUxL1cgTgO1
mwYmTGC8AvP4FVyNIX/0+kRoYvPTOkxQf8Qj/RtxKMw+iKNHWsqUAdNH8p5DSKrbro57QznakjXY
j3EG9g4TCyZVP9LYoAiJPLcK25TCs1NnYjD5m5K4YJeZJ2dsh34nJwlTxxPjnBEr/hLzV7BbtBCi
HX6K5CYctBobgd0tbsEpp3/vffWURcKiCd6H+SX7sZ+SAvKfUTi+985jcfQFJiQHHMMU8+K9D2KM
nuaHpKbDPGiZ2dM3YwcOcBoCvyaypRNfVhN/btRRUYjW3jrsXoAkazsapIotMpw5kgC+JoveSkpG
B/Y5y2T1mrfEo7ul8pbSVdArH9v/1KVO4MUWYxXHDzVLjJff4tbMUoDnN14C6K2duLToTFsqDGeh
eC+CJhATTBBpIPqVkM0zimHrSZn85NrjQfdZkyRriSnncQmFJGYuDegyYccDs6r257D26JerrhBd
959wKI3TCW6GvU3fz7skJIZR2A87lVbrvBnHyB+SjUqvkKsKN8H7l9JOjGBzl2pDQuxXrhv+0iL+
k8xenHVgD2ydzxd+WaDSGkhlOjgfZ4F+y3Io6grIZSb9gbnHBCTFVwSJ9M8mifigFtY79ELQaPud
LjDoQiZZ7pvLj2zAoRqbN5UA18rHmTrC3P0dLqJsMV/E2IMDV3oc3o5/LuaI/lDyR8i9SCHpfW0d
u+S2ESRbtC96UJnQGrmGqoajtx2OgvlgiLDswgCeAbVoSEN8830yqtZNGLMeC7jVG+a5aLwClDyy
eoWyK8laR3Aj0OcerMUS+XPOzilMYQSxkhojyBBWcziHlsqlVl7fjPr2quUg0f9dEZhQK0IIWPRA
TI8jpDYMrE6SMWRh5vHxJV+nH3FZDqBKbyf2mQI9KSdYCFnT/Q/ap/V/TPGQN1LFKEA5Azezc54F
LLWcP80GLqF0OJ2AufMHiPCwr6DKwPyUVzCghpwHte4UMMrg0Z7hDmQlInABnho1b1Wlgh6dWltq
C5eLYEYuhiGeS2+8l5Tdt88AlEiPMFCPRN6mt60+sboNbSBrlwQfHQCJGrc4x0PR3TGYE0uwmJyR
RWw6IHifz7kn68ACwmjMN0lFndtKTMpUNd5aKqvUys3F6jHn66EG1NjXsSpxoY354uWymE3rhnnH
pBn4wWw2qXXXhpP7ig3v3AJRju8b0ydmlMpLylHs5xl3N4Yu3hb9cTm1H0+GD3O8mBD3GyGV0Um7
LsxK2Wamm+SG17AlS57nTMgBJk8K4Wl8Weq0tAG1Nf4glgaf/i/2EjdvHeJq8pMi3DW4glIHeVFd
U/0E0JvfSkuyu12bHeFWbl1HJvDqlMXzZuNGuroABSZOM6gTALxLPrnfvLBMmK5p/kbIRtxQEs9t
gcIh0LV4yck0/kKvaon1iZAjeAnZ6N75Tpq8cxR715ycKDxsK1Rplqx1iGesnj6mXJxPAL0tb/DF
zSRQ27C5+Bsgn9FsCI+jhhn9glJj7YYWMCYVuA/Fc53B643lROEn64Ap3vWO4FPIiJj2Jd0sxPyY
dCdWxvT/HbI+HZuZXB6Eh/ZBYocAACCqEU8qsoiDS9qncjvzrfLaAeHVSgZoX+5mUidCKZKmH+2d
LQs/f0w+IksvlBzn+cuPbBEunwHYw3cqLJG0f6fIJMBpWkdsXTmPwM9OsDqHdxXuRMD9paSpPb0+
4D8qUa3vKrQr17j/4XT/lzXAXEXE0XvNaBq216pOyGxkiTHPQngUdsUlfwG4XWTAwB974hGkJ5HT
qjpKGPg+xw3X8rDzrXRPQbhNxa9BlXOHkrRvnZK0itbOokorOoXidaT52Dme0sXBfeE7R6yKXEF1
8BmjRHmSt9kNH8/liginf/0iyvYuJI5g3RI6SqMWllYiAD6Hr9rfP87Myd7LdibS1Q/H7kyQoYbL
uRMV7auc0AG/u7tne2/FkldP6/4sLr8uOqdH2MgSzqJAzJLt7/ALufvAMNsJETYXUaMygUzg2HnM
hHWtGUZcGmd5NVoXl7VTHVOtqp87n6tB4DWlQWRQ9xn+RPetcnl9/jhaY/4UmL8kyjnOtcgsPGGe
hbrY34rZ3a9D06et77YNIiojn0EjgO/yQTDa2w38Xz/AuAgjENgepufoSGgvujmhj10PzfsozHlb
opjS5Pmr5mcYVTIs3qcUi8ESnikwlewPjsi2ctx9si1Fa6sQcVsdK+cTP2nO47gWRHxLl7VTVYH0
aXv8PqnPKW+GtpcKBjTBi/jFGQ20Ca4O1JlFZYnNGvP23vuhgl3USTB/xOlFz8a39BqErC/za66l
ne3JM+gx8xo30JBY6gc/8uHu2Wj6819jQOLnoayaWAmtPHOYLrPiptln1R1s3uO5dwyg15Dtq1X1
TCg7/4ZQ2qJr5pYLcR6V6wXAad81hj82Mu01R1cH72IJfLqtqf0hNZpyHvwoFA17GIdV9vpfaQ8r
O80uO5InvI4RFNY1rM3quvLd/Ml4Ek4xk2hc+ZNEBinyaS2XYNDlBKSWJwD6j0QHCAIpYfp5GTLX
/+1rqnnUltHri/sxqcAJpUGs82glo1Rn/+SP47A9hfQbNquQYGvobn4hcWfU3M93B+w5wfTIxqCl
lJRfWT5c3JB5hGLVWWT9sSVkljdiNUZ07x+YVgvzvbb8b4dEBWX3EQ+Uz+GC6LwlJxG4koHYxARp
cJ0VfvRmbXl2hnLNpiBrWFy7R1wUpNRo47EQVt8gyNCBcg8M6Vxanf5O+EONzId/dXbYZ5Bibqxg
vtklQqy5uONNE4qDJjqanvZJgFkPlX0RNHoeSImpJCzk5xzv0vP2BBgatey0iz2x+tGXphJEufLL
NKyQtAo17am4wZOjVSh0l1kaXgz8g+foNRLNbt/5wd7zISczWWkVs910B2Lx1gkjP/nHPgU+rRBQ
ResAipwWw7W3AKvFO2kFlczuzFXTxFd8EE5buPLefRLXxzwRBt/Pb+H6rntse72tTr6yO4zFqzJP
b+eSDrUX4hIyZJaNytekdaDp5Jo9SkqhXwLqiUkEIyelhFytXZnMPDkm4NgrWTKVnCXRkpVnDEMI
Gpr+RzSJJtJ/f3mRDNEfHHsrA0zmh1XvN9gVJsxWxSQE1ZrdhjQAy/PF1xbJxze5gx8YEiE5g0ki
e74l1N3OeAKMEzk7RbeUodpxzZJIOguVwEjvQ77lFtmQbD1+rJCqb/caqGglhuJlA/BeKJElRx2o
aGmoN3usgDc6EQx03v7ssUqU5Gt9+gcxQEfg2ulhg5mUJRQg+BkGuWWqft85uFlvQxdA9XgY1noj
a6YGJffGmvpwEDqBiwfQgxeDx8TI1r27ExKW2EfOrFsSoQH6Z6Cc3zKeh7pX+SWSsQu218M85vIY
MRjokQg7T7Ud97WXRqTQBCUcNyoebTnPwwHMkJyGapVtFrL1eVQvXIgT0F8Lx0rnojAUDtWqtAwp
+xJdhrEXOTVtKaV96yiyrIO/kSxUNCiQjgs8VKQZkcXY03cZ+/Pdf3rnbCCjm+AvJwakpbJidIZ2
rZ+G95mfxTCMhmqPKvY4uJLKKSdNpCjDw8VNdD5XhUtaZlFLoa5tDSI+VPYNjN5XISWMPVItoV/6
9aPHI/CQyYw6t6/C+++v0qEPkCCfnUb8hFR4LMQheCecNIQhl6gxhUzDP+/2WUj8XnH0FlwIWu9T
0rGyJHrAmE6oo15kgadfBBN4CkNGgIL1TfFIl45TdzAk12hF3ZJh/hhk9tU6XvskoQeWLBwcxfiE
feza2JMigz2xbqTeIvJ9mgt7bTTK29AVHfdiwAqInH51entaHx0PF5NlrAL1niI6nQ6s0E6LWD6n
qyXZVN77OdkdirXiUuW1lPJJ4GWAML1z0TBtogbBm1yJlHlP1YMf2kdpfOPG9YbfGbGrUaE/gq00
5/L7RKypf9AxHgOofiTK+3vdwpqFlHUwzG+BUG3dT7KlpBBRxAld44NbbTLViX2Lqbz+zz66EMgK
FuqzWc6ZweRUKM5mnozOOi7+PYgQvXpws2vTiRzd5SCLmerHCHtWtJeJHaKbcVGZzcZ5wtbmMkPd
z4DlqNtUbnM5odoHeqcIUBCEQ6eqyQhK6QRD7E+8H8cK1wPcwH+ro0CZcQjOGdum5N3DYlPKeX69
MVYFskcZBlpVGsQcS1d8IhFEVkZSsZqW0NXSIOTnkqSzVGZYTrNVl2ohtkKkuDs/G2fduncUoz0a
/6qhMh6nX7xAiDfw73JHtZRbnwkfTeJpGFmOn28jDgPhVVEUAWeVkh+W28SBx8yqnP58oF4BeM/g
TVE6Brli7l3cAea60lqOpg0NlEdMnQfswQu/JfrJsHczjt7YJLqwXENf5ZQz5lOWQP72rsDU9LdU
ERJQSO4IN+DAbScB7hhjDgHdEt70X6/oUvV9+UDXzu2pX/5PLAhRNcWPzZqAJNs3F1rcEGspqDEJ
O4R+nYDs6CoQh/icLLNwVFmYYHDvtmW01JHNONmC3vTD39TJhMXVFpkVRZdYyp6I+sq8Ko7yugb3
m7/JehoRb3QWzXpVLnHwdOApbBe/nfZ3f0KGh0RxJLOFzfxG72aGL1neIHETGSYYAJw1v03rd+5e
dBbg46b21j40glI7+WS++zG+RotCVW1nzMMaFggwKMUz3+jh8Pk9TBfeFasNmenoHuMqIrHSnYCz
RJdgCvvaplxC/LBK3f1X8DA+5EKyhNtXsrjOmzsJ9L+FFfYqj/jI6hpZI06IVqPXDhIwxo4dlZbJ
ULu59YVK5S3pISKgcj5RCbSbfb8wXw9CbblLtDU7NfQM5R+ngJybxFkvYyiQHo4C6NkcXxNdsfo9
/2pMp9KeBdY29QPqrRd2fYcaU/nMXSSTbam//0DsebqjtLlswoxxrk6g6t9y6XFba0Ash2NbOUzM
Z2EHKUp4Ke9Xf2E7k++4bXd0bLS208cia+Lr+eidp5MoNmTQjlvlr0k5+OSNcqq8Y6A7tAxvtf2w
ywjBXsfDGUw8VSzFV1hb9VReXFfczTMwybPKbkyiIeoE/KvTy4JzfXMMr0cwIByGzw7EurWdOAav
Guvz6i5LjFfwuW4+C4CBDZ/w1qNSuCNaPfN+VSo2UIise95ZskPWzOB9rmKMB0oc/he5B9GtIkhd
DMOEfiw34t5jO72azy4WpUJxRtgYCvRAMi53yFNUTggKDAoimKxOUx2RVop/LWxFw6sQu8rWIY92
okLPKmOUARb2cmh4rbwe35YjbG7MsCwd13bgr6hjcJxzT4aESrnd0RLYJ92p5ow/kMMQkPafJY5j
zJIvlQcGsgXZLsNtzofxerF4XY54Z+m3oYGcjEbZncZYs7gM1pQnfFPEXbFVzSebdzFW+wZfO58w
+6LekKnnLPUpzQjb/QBKNE17dk6wGxhqV0ICu3djjG+bWTj77oHNF2gTF/scnXIIjLz9xNdAWbCt
SD/jYcLeu5zKgd2BJXuh5a2vvCP0NeghTnEqTEM7Xfg5obzmC94sr+OU4kNTJeTQr3P7Sjz9JmJt
3xNKPal+w5qYLFliu/7N1v5X7GGM0ssFpM89tVpKsI0HDdRIIH/riF0YKUCLZHwkPOMKXT7KxiQ0
j+aqJifFKmo9xDAYGY3abo99S3AZbkLCoekCOhvqEjMyj7v2ZXMjfG5KmkMbSUUep9hCtAy111QX
SIxQRQSdDOw1Smwk4eMSFevW9p3Qa2dhlinp6M78S/T56t9YHezURtPgriaAAMvjAVyiJCkNSdGv
268tKi9GPn41a/dsZMLMorGxbrRjfUqC8nqrczgs8aa7WUjIv520WYtX+A6ZxOlGAeyqR9ZbWRM2
x+K1I/zVIBVi3NvjhJCK0OWZYyJIHtVr4AHnijSswcylaLPegfomgPGNDSndpHBYXkp/MXh1D1FE
R+cBBSS+NFXg7IdhMaLsrCjlVDG8NV9nGKznkTSlm4Hvw3WcrQCY1movxA22ZInR8vYtMVLZUB9c
Htnnnf1GH7a91hhIgeCKcZIt4JNm9FFQK3G2MMHXZo76ofmGplSBpaSc/wSAwgxDGRwiGXQljvmu
BbB38+0vUYSTK9YL5/Dfq06qUxyLUUdf34s+lko6aJMYFM5021KeuW3r/fL+p9Y+IZE5++u6aOKA
5CDxkpmd3grN3IYFcWKVa/LSaTsqyF0HN5HHn7KOde0T2Z1YRQszQAdoHUVk2gThZsoBxZuPZV37
yiD/uSnnpVG7DlmhTX0qgicqBg2l0guTdcNZAeFBxU2tTnrtEs8YdcGyvY3D429uE0NMJlZP3Kvo
JdA+vub5gQYw/0eDEISnc5EH+tBDqka7BzGCPrcByYfNBokkmGtv4S58Y5ipV8YdYv+ju7QIl+Me
PfLKBXn+bMZO07r+aL+bNy+6xzymOLnUx6t1i8Z1uoTvGaFsDx1XkHtaVGb+PDmaplPksZh0ZDlB
O6c7/Rfm8c36xiZbqZXnGhmcRvFx8I343K4AbZaTLwSzEAQSpDu2utbeohJU4lnwHszLyTIXT0pT
5L74uCj7GA5hM2duiqgtLPBoA7f9Tn/drXJHD3QTQOWours6wG72oBElU3rNOt3TcLtq3MbLn122
rHEe57YbbAeoO15o5tWUas9Ze5djDhzq6GVpilViluPcngQ9ahdfecdw0CTk8vgoMxyz1ltjYET3
Ac+wFwcHUd1U+WzdH97sVpKmR1CYSipbzUtCFGspb410sZFo9BbCkZ8YA0ey3MZwDqvrKhfVZ0r5
lt9LcPpfAu38s8nv/ZxNK2DvnpI62piMqM8x3PSi5O8GqTqG7gSjYhAD7ybLdQxjBIeafWXrzFtF
x04wgusZ3zrQ/yTVihApRZ27xauX1OZqLyQGqNXXqjoy5DDtfDHH4aDi7sXK3Bv+vXuXV8XLupjF
4xgFjurbiiOOXYAzJQIYgb4Ns2cpei/K8Vw4fMJ3EH4x5DtS18fkBPwGwgt87b+Zok7lcjWaEosT
eks9Q3mTVNSas6wTuagHELrFOBSmI+28nEX6JgxqCz/ECA3tMIqdqS77J13bWBbNzu72cchFRQnd
B3Z0c8+b+tAuOXSNsDOUTtWWRc3LIERXJdgKRcUBgM89azOvfRYhiqTlcdbAuDsFkGF3yTfT7oJU
B/in5u4h4NCUfUiUXARWcEcQ6OwEQwkczfY6Vqmep7XUtquxvNP9onpWd8yVx1idkjYqVIewS0lF
LU8k5/Z1+rsu/r7USdwbW2XCSghrQfA1LyHqg8DrOkh7KweeChTBL3iKp+R2QNoJyHPQNlw4T3zs
UgKu+uqrME3dZBTnjuYQdZEt7NVc6sEChNHBKnI1BN+gAwF/0/f9MLT1f6dliXg4LFp7eDdrZPkH
lM14fpK7G85ogYtvTEQFi1HmFrRXH7MSGsz7cEyY931ePw+PdC/xnRZis3xqDPJ+lUhq+58fiWpC
2/DDV5xku3dhIT9I0S+kUa5T51Ade0a0sAZqnZvXvP1dhXcgzO0hZCYOBwpEWVeczQffAWvzCH8B
/EIHOuBvyY1oH0DAlYqpG83YZYsMG7OwaaLLyharEKjvRFrKQgb+wMDxXwTQHoNx12QZzuyH9hvM
0CYdqa26L4IRdmtdhtkbSqfAY3w6m4/c7paLm6Oe/W0+5o2EtHixEL7lFrjaxq89F6YJMh3jZClR
rJkD/0hnrj8BqwgMGsdopq3H2ipZHYLh2B0fjPT9za2HD9tGE4vFE3FWZ51gnS5OSQitQKJvB/EH
gUEOJrb2Y0gwyPmf/XgN5ciharIpCgknUjbcKScoRYVMK08Squdemdfvj+Qxj1yHd1dCGeXRw6kT
HZawsL4cwuEpVlMcSFhCIuWckd+Ohdug8KH9V/WzQNGCq01WQXroWziEefwic/iwPmPZ0Q/MtUIe
8/Mu+0TNYiLUiWpLAqGsCuxp/TKFoZFtdiwj6rLuLX4s9rhSjpWCERujDhOQX+vFg4rVvaGhrn4f
2xpHzvdIiu6jQkz2YYVVaxRiW4dkCdqno0O/p0HzKOxqPI/UJR9v/wF7UXzcDSzhKz/tUdpIi1XX
CpD5tgTDnYt6ONSw7ueG9qsV0fLXRTn1swHrymvgDUAo+3di8NGhYqc5IfWnUcPn1MiDdpLNN/TA
y49iB+40SeZ8lJcsUEwUcJbwZfH9pCye+RKlsOEcKOc1vLULYplswTSiyQ9uehTNPmaYU0fpQzDd
qny/7+LhtCoR3be8pi1SQebqII5VvgkRydjoYbcPSKQ9HSxrejVyqgsc1YdzaXaI9IM6ebpLYDTy
UDwO+RfPb1+qZQ/V6NWjr9sVqxYM9bJ6j+G6ccns/dizlQkq+q7vdPU68hnKlRPYHO2W0ZlntbWA
uUO7MvTO6hwhKKt0bQbaJdPA6tRqTepYHlRffEG/oSq7DHjLsOlSiBR3zJLC9pPT/kpQY5gx51Ij
LIBVYdOYcMtXdBjV5qwwD+nwbY7Q1744aEsFO2UFc4Tk4VYfngHFlakLNJlBRSmh5b5/Ux8ivedT
Vn3dZ4bhnhH4jt75lG2OXTKf/5gnJfN9wXtJjc4WsDS4YosBv6pZDrKk+AEIdKS24hH/Phjzpavn
fTb2kmNLJjZCkbNkf7Cj1gMFVvcyKG+l642X059CsL1udFpTjkLpXL14krYeKeQBXwl0C9QnZWVD
//TIB39jfHeJM/uZD6A2fvFkg6BKJXqeTe3O1fJtg4pJRHKf+o0c/7ea/jCgyVAUk2KLiraJLTZw
WR81lDImtQzY8PjdAsxnMRy/Sa2o094yraZD9O4bHr/ZprR32M0yxNArzuY9d5Wjxig2XOmYa2O2
f8Kfidz7tksqmjK4oaT+PKHY4+Htv6RZ1gPQY+Nwa/s15OQioOiDilZqlUsqVrQaK5P0R/IT8M8i
tdhGaIMjHpG9DbY8RHres4IMF9itDeRjjMfuDE0rULmPWNNdJ7thAvdo3i+swX+99VtpMVjrA9V2
ThzHg1JQIVKQnNnS97ZDkAneTJVamy8Vg5gpANSJGECRxJO5zbpwvA5hAo1RA3sgooa7uXV4n8SZ
llUn7wR2b93S/duYB8YJKRl9iU/qwbsKz7rF6S2Fmpr2Au+Z4+dJ3Q1T4X1Ky/PFlHIYy4lHQW58
BNKMjAVX78s8wuAqrc+NeShdsS8LQqKE+3aKXNNmGy5gNO5zcEsjRWgI8axoQ5XhLrDG3D/wOaxx
VCbakyu4FQBSA5k7IOJHAGbnFEPDKu1/ZcDdpxX2IPS9CuEQ/U9owZJc+nkiiGyzndKCdbGh9biH
0Gyk9lq5UM8pu3g2IxOwP7GC95mYY7d3tfEnef1WCYLLO0BwkSBB60U7tmN0wrLlFQ/fyA/Xn3U1
eoUsjHnN5lyenuYmhcWmktUzUiscvfR3lXXQtcrLZevSjyK0JDksuVEkZtxEmLSredlNdwH576DZ
3klfJUycoOa+VpzkKRaeZFRkTYC0lWxENNF45wzvkvIYDK3739hnkY2gouQ+7jWEkWxkg6HnZVYQ
s8WbXkO7EaXJ3Br+BD3fUW4fG0Ah82dCxcgylgvTD4/G70FGHbSfZ8XhgIaM8/pcCY16iCdr7tHT
I3slmhbhSrfe2zUSgWnScPxHRPnN1W7KFHc9vhLCUWtzfjFhxEG7FZ6Su6Md/gU99dl6jqs4+yIX
oWiAbfaTLlCC7MmLTJEmt3mBJrqPdCbZtk0++N2F3LqWdLQh7aDT1q49WnDTrIbu8z1TXPFPfiSA
TCBo3rUUAJOVXEJGvkyj13mJ2xjek+Ct47gZ9E7EyItpBh/CFHas/f9MbOp6ojztT1rQEcozaWCw
Oufg4uGvCvgwQoVWPx8QyILEw5AkVrIhjTPwA8oZ1cQ5zupufNu8JTj1sKVsYe7QbBMlO9uh8QFn
xegzB3NAuMo8y2xlEEH9z+HbmsruxYHvsvylmjQP1EUULBsR0gs5PlPwtFCbuVnRCE1QfyfoStsy
DPyZtAKweMFbSQPu4OnbXqPH+O/O3fHhObhmV0cbQ3lAx7rxiJayFnHt+d9b3EM7hRCscZ4IPMFo
l7tMtZumic6LPKaH0GYlCinLz4u8J9JLfFY1AfBa/EJ7d9VAk3WEjIGYx31Bu0F98BS/bTuFO+D4
tlwwKqHAtq6xoOKBM5+AmFKbx/5yioDPP2+jlTkV5TErJBF6nPRaqRzTOI0ZMazAlckTz1BHxJ6O
BafoSmDEViQWKvolCRzjLHxBM2kkQajonD6Y6GGGpbaEyt07BlWKFRVlL1MXuR4Uxba1+KV8siYY
YUyWRn/66qIqu589zApUxwuFs4juQH9DZbV7duyj8XsirW97O4SxF4nJRbNRrwud/1Bn0a/ny6aV
ZNK/9eLjaXifCKEUWvL4tQqh3AjWZTX64JgKphlWaGkb1aXbGRKs/BfKcJbojMakj4NEBLFLGwk1
xm2EziZqr9pnmuvKwRdb1tIjI7hqQz5FnPCs8dp7tCc4x5yEI7NUCLkQuXjEldwY61IPu2N1t2fl
RrHrGBEKr8r5+2lbbgvv3DQK9rE2chDy/aol8jzauHOSjzZku4hbQpvaBfB/3LJBh+32zo9RcHyq
4Tp88om2xksx355SJWbBGpCa7ofaeqk5AekXx0OxUAGdyIwAVT5YchJP3rs79aiqejl2ncRBfBVw
3lxG+R4XTtTR8TRMmCcs+3oyl3WI6blmLZbyGwpRLfFLes4iEeMA0ITBFkzoBs27wijOhe8i1zXY
tGR21/kIgQpvwTqZ6AeYbm8FYJkY/kapaNGIt4392A2WeoGlO97bkLxG5c+MGeuZ9t+eXQ3ph01v
h/YBUjHl+tHacFKjTxwbfe2YivXuV+pSv4H+JJYYi1hAevja/dA0MRP+xsmdh1RM6rQPE8rbYmz0
pz7pCbFJekilAnS5kSdoNNGC84e/WRnXKCFeYmf0CzT0hdo4NW8manJAGYaOL/r8tx1cg0TV/uQN
UdYlEf2e/pjyOOvtFjubIEJYa99LHvgm75UyN5pHpkuXzlyhDyr/XRybLk8Gh9r4ZPTujOBkW3J2
MfhM05TyPdbeZe+0hECi5HDVMfeKZy74EHd98EyRB1ppAjduwDz2CQEkX/SUVxp3GHeLhG1vUDct
eJq344rhTM5ex1Dz9OuThzZUZ2851hdU3dp1/SLM695/FAYPD7WLhS/TyNZgLq0dIowxsKGXGb81
ugDudvLt6BCqFfL9UVCwq+7rHRDIASYwRI9T4gh0JOkXBqZMBZ8VLYPJnyoGKm6gpTlO184YAyRC
nTOqUYbVy9dJ1qa23BEHgB8rfl16+rhCt4t4Lvsgp8gUbIn6GxWcuGBDirV4SvZuL806Sc4C9IEM
HC3DdT6pq75/AejH/Q1QdgcaBPj/ESTPerILLJa3u7oVU7v8u0J1ZXzCfc+PtkkkNp3VXRDq8Jip
8/CFQ2SiZW8CFC4pEkvJQNtWptDsXJa1R9PmJSz4aLgNjzGG9etqceBLC49CF+T3jhABNAAeLZRx
Uy07iglZqhexNEip/PSDSb1G1H+f0HPV8JVU1e0p8Fy4m6W+xTFa5dMwZj7iZCQrEptdHDMOz2Fy
b4pLFvf9dw7UDQEjMCgm1uVHFK1lMEK1zeeKOMSk6FC/PQ8QsJQrnI2yWuxaPpUiG7E/xTVje67t
orR/l10xWFhw8JD9DZZk4FtcHFX34epcCY2TLhwszUtCP9hWhs18kB0060BvMuZTw1YY3wHylAr9
n6D82CFzXtn7dPKSCo6CG/87ap8dX/uz5ZBT/4GZj5MuLHlGRzxIYgl3vqNycZj/SB8tB3T4eaVV
Q0tpuOWlNy0nl8ej39nJRFAA4q/l2q+N50pxTy8UxIE/F2vedrAAbmA9nb/xJl7p26gE7lNbyri+
D4A8g/OBYOafsTGzKH9jUSt/sz3DBvhRCuns3M3IwcNxEkz6UFtYegOuwrOnmlsJhBOgFmYLn81I
v4UEE4Ho+OU/U3QO20G6IfbFyYa5f7z/gdBGA3QiLAE1jjx2gKvdoFP0pYfOT3DFBP0q+PGo0zRt
bUEt5823w4Ag5oyU9yNmwbskcRaGF9APC/MEmfh6vxABcI9GlvA4SSMNsyI522M1q5CEfYF9vKNz
6+GgqNR/+gP/PspAneo5H9HSqhgN+w25hME8tBvyhb5vkgfbGDiTm2DQBLuM8O36sIGiTRjLD3IL
sw3YJhSdjpmKtcXykkiInhYEtPg10lkAvCSNlyXxru6qzKVB7zSM5MEJS/98CMvaa3Z8QnaUqufv
O9PEsI2kh1UeYFTKHDJD47Gcmi/aMtDv8sRFfdjQfu64QhGOsjWHpoqfwWw9Rf0bmdyfUOOFABH+
l6pvJPPj21jngZqBpn1n2hD8vDDsmdRcbKW+3pYG1tamnd6+SWN2M8GR/jJeR4FVry6sKrqBZHb3
bhoAu5eKbam6nyT4IInoGLTjHqwBnFmMYFd6L0i5fkMnWPJPPpcnFF+fxv6v3YuPT9Kw/I15iIUi
BDc7tWKYu/485QaexMM19bIMSb2vIPevUjxDY/GEj8gKwKfNboSi6EKzxnVCtXfXG3PkMBhQ0c8c
IIBQoIKNH6UTNb+ENTCRBsVYgKTlG5wlpWszB7X2pHeAXdqw7/QzftIRuvvK24a/Uk3wqYmH5ZGN
s2sLYDUq97bjJpKx3zyyJKjUYM3fgwSQtUqZN30WzkGzqquCeltQkeKg+6igHPpXouGjvcGX+hUz
poEq7D4q5hXJ2Z9ce7N7FweePw9d0U9m0XD3p07fTwkjSwucX0yjncHFPYb6fR2P+NUpXVxxTe+N
uuot2W+oyr3Yk0QQB9GJfZc+Ne7zErKwfSIMevUX1Y8fU7FCr5QIkDXptxEyM+ZCFZR/8asy1gnk
3x51g9Vv0jtge3XmBWleh/s75g0gu31tKPtYrL9viL92pwQritVvDe1x81GKqVq1wMjDkS6Z6d7Q
fj0zfUauM4wt03vFwMRwCHrcpbulN8a0bm/+QTMTSxgMiT5+18JL3mszCM2lEEtMbKbKkJRw2LPK
/tUgp52DiK+dVhPojX1kadxHVlO+eaCcDQXlllUkb+k0oJPORKfDyqERoPxpSYZxHMpHQCK/sSBO
msdyhtaqsslBGB+L3KTpth2ynRfZu0XxeHcNchkHzG1whZxdFr8G1MkBmALSJRCFRKQJ/ACWgEA9
7L8gGlZ3QCn/Hf04J9POsyETrImOOUuXVNUYE/XcQd+bmbVmaXPtWqXOnAYJ1VdWmfBQW2ybxzjw
SG5+6kN9rCFGdV+fPIi/J5SKvX+GGAzZSvQQ1nUSHlQrmcA0w/2D8vsizv+xRXX17ShBadkbHwgU
ESw7C9DZsCt5IBW8eiERDmRA4qDJDanG/i85ru91GEtHE1nPVL2tBOiqyZTO/8B9JIsTmL7ofXx5
AEYzPZMxi1pH6+g0pTT+N+RqOWk4u8lbDpDiFzhni2M4eBK2O6EEITQDLpd/IzPsyQ1OFquEdpBW
IvTAf8V0btRp2IvcmYihecG7ta0w3783fSb9cGWkbUbWgThQsdp0G/0rmp4tE1PgJHGEQYyJMwDp
PDKMx+emhgJf7FZFGMGuQ9Em9QXdvD2i4xn8DvayNvXfud4IXKNy1F9mCjXMmJDVfR78lUB9QIq6
Q3vGq2VTRI74QdghuqioNFqviG2zrlfnkF623o+jd+/ZOtHI1f6wVnJF5K3AY0hVraEJpNCM+a3J
mChgANJdSKjD+1d2eDjmGsT28sEKbN/pLku45kKMdcgG0ru8Pt9OtaSCgjF1ZYLund32M/RNqFD6
MFk1ZBFV88PWWnO/lriT+xADYsUhW4UHbCj3YYykPhOgz05Y5+E1tUclMtYVhCMY8tQVBoYNfzEC
Ste1EwQeMMespOso4XLFh7BvLjjBVln1buDcw9eRmb0lbA8raus54P75LVUCoW0prxq70Z8fTk+X
JX796xsMRqRQRHNrSg/BUx3r4/EFNs0Gwn1IBkiFginHX2Dc+sKGYi5itV2ivTNqKo7FalTqKQxx
+bwfGFrdempyzdjI73WhQ7sAX1UyWau1euXFtJGJ6G0qafd7yxIGV3ow1JH/xlrBv2LvuZgy7gdA
Mf+N8BNJVZR2HA7+dxI6HpnQKg2bXKiYDDIXOO9eKn+a25+20hfJRJN3jXJydKzkMDGvH6yOuAcV
VIseu9HVIY0zfrvnE4CCqvvq2GwVG24koGfm9LLr50OiUPKreFqOfJ8yEKrZ2QkBfaY+XDq0nu4C
K+dSiST5PkHiVNL8zd9D/DPB2QSmZE6wGovj6Y9QmOdI2X6RlgqcD6ewbmuFghqM08J7wHxLj1c6
nMTWAjta6MIRXEMQgbiGIWIMP27XLNxmPgUTDBOG2AOH/1cLZ+SMTVs8wI3PVS+kXq+PeOqkRpb/
dAX4d9vp/xqHjUgzjRzm/YoIeMriJGDDR6RdNQipxGs0v41pdC0mfjoIckgrGFC91vB0EVGPSN0G
HG7CpLP+KLVHkVEoynpzLwjbFWxyol5eBna4sYL/1kQoefjDRS5biHI24cEl5GHrLBVN02AmK3ed
MY6BlqnQSITQRsKQ1N/v9CLXTxrn0hIfrupmH3VSnIQg97A00nQt4w2g0xFkj+WQESbOcq9Anutf
OuHnlOy8j07HHx7TzKCfO5AJL6KEVAJYg4ickA/KR1Wbi26/BRiBmJFY+tJFvlGLhdGXl8NrZQ5X
gLzGPEsPIDIK6LjAK4uOOyTneh0tYVTscQ+W31jADWut31E4Gy0FLeTccRTIoT2RYgJrasIQwFxz
J9FzPtX9DSnoqktzwylgI2qcm/VmChl50LAeIRivrVU4oFPFOpWFjmrr/P/NLdbBIzWubodSeH2Y
DKgDioQYUriwFaG3QnE98l67bbCzu5qjXze2Llo2XEvtZtlvydrwlQKR395rvsEcyJ8fqZozrtu8
HNTIVasvQf9uZlpdno6gspbacPZzODOfs1j+5qLSbSHvuZTNPidNLoY80xEhJIDKYfdd6KQ95wU9
/7fjSFtLLyDDaQMCZbe6PjEM29ZFJkwxi4Uec/RsJNgkRKAkOVyZvOv33JMcCP3fS1Wepem7s4YZ
RlvgRrxYpszAFrwrxbMxU8yqiVF4r3rY1ET0P4/kLCjE9Mz4WgsL9xqnf3jSTR3dFvw94B1vlayu
AUnw63/WoSts0Sewp5cthnYEKOuypz42VT/bLjn904sficaIt6NoEmw6NT3qPsPYzHWAQU8zje5k
C4QqXK4nBOxxZvZGfdUU083qd3mYcDAtNN64s2B+8H50opwih+rlbN4nsTpXKJiip9DRHjgY2+SG
F7b9PPfb6L0An01bIqW1n8njFtEz48YFtM89lWdxShVbyJBzPMHU0FNCLNNGUZaYUP9Hm0Re5SUr
dJ8X+uHSvF1Ng+ecABSgK04OqM+7e9U3Qb7KnfF1kRVLBSWroYwrH5O7tQPbpKHY2X3tzX0kNPVf
T5zh3oCBChgA2fmteQ13D4Ar7E4WEumlVTxCZdD9nvG1VhNl788NH1tPsgCxniD/6XgpHr1KbaE7
G7rJLf3MWXkFhuqoAKiZHtQZB2cGE0qK/muc5ZxhePg7K2xoV4utIeoo7f7hXPGbtGqW+Z+r8jXy
3SO5i75651dL9Q7w6Nbys15OMARpotFpC2z0mnKKJvA08qelGKB7lfhnD+TS9YCgMyOxKPuer/CN
JKwfuK0K5j4wDiY3ui1Pw//cmzsRCBz66PYa6+8SBqnDGJ3wcvCWGTW3Pp0dlbHxYfA/mJvkDhNr
Ux2rnF4EEtCqn6X5Yvc9VATfykwABZDJpgMIs/bfyO4+3p/qDsR0lKmGVSTJR0fwf5AY8viQ6jzf
LlkbzPfq3HraAXOUhxjFJSPe3BT1y1FXBhEc3vOi2AEw87wFeMpgeVBqHxceCeXE6s8nWjvRBF+k
aXAa0s1EFLXZ+Xgxfn3c3H6I0NThu5iLzJtoJ3RdXw8fvPaXDxw6pwWJ4uA1z4MVW4pSQAN5Q5Gf
IWcxFM0IOR7f4A2xByQNSmgcOP3AVlfH8lOoEuuoLLNCUrT5RahD4Yy8jKOrPOOTj9eFqOxo8NqG
ZlpBA+H0vInrHs+0GkQqbxoye0eTycAm2bb6rU9cVql32b3p8oMvhLcww4RuRihuZqU3M6kDkeRY
6v/vAMDaVGr/gDzLsJMq0RQB/60vzEaU0Tx0M0HXDZX3I1VU710w5B/9IjDD9N43ar5pY536zGS/
DH9Vuw8a2FS4yu1CdeW5ukMnQhkHLMlxWGPlMdVImOVjuXaXgE4TWlN3WN7QwA1XBwcXQqjLyuTe
IXz1FSMmB2U4J/RorlZ7HD0Ym2Se5AIOQXBLLlaX81OO32AnYtj4twXC7TDNYgIdwUTCGewqRKx9
WI+h6vMULh1d+qM2/b+Db/SNGNOJkUsm9Pde2GmTwN41QdKkRg5Hfg5TkNMBvnN4BMa7llsvkfDQ
y9cRhmBIjbq0QPWb9XhW0TjDo+wSsyZtLskZfxqdbOKa9/i3yhw570B4kWLefrTWa8fZCA340MAn
h+nHmh5Tb85WAtXo5VWHNJO8bzIN0xSoTyMYmQn8gC7RH7Cm1DoTDNK6w8V6sJZM6TdIUmFyDtv1
VMSd+E0j50jnTyoN9sgTOnOwLoFMTKIPc3EVjdL/LncOXwHtL8hIm/c8LkTMH0cB+H19HH7D4Esu
hmC5VDOpcjAQIQOYPJZhVG+KK/ti8/nOt6wig+ZyogMG+yvebp2Lv0gaGGNgi+LLoHLZOctktduL
1IRsvLsGI/xD2xRxRCK9opyCCNyGt3C1hcxyC1nCQB/jn58mrTfuMRG/1bFMsDJoFqtrWmQgpzG9
+1SQx3n9gEXvlNKOdCb6h/miSrH/9kypFzwfCWNABWVUYs8TadSayovLsuUGWnGQVpRBpxttL+I/
+ITxrG6puJ3HbW1cjtWZLnmuWXCkHCH2R5SGcLIXlkxKM3Nq4QW2bjaNnTTtZ2pLbK3yr6QSk8H/
8WLnGhzvC5AKlRUdwrsyp1Mt3XAyIU7qdaijfKyY+r2ifDy0d6xHhC1ojwWDEidaejVmdv6o70L6
04A22WcxLI285M0ak9yk3waWjw7rk1F/sCOrIBeTeEKm/pQa2AfKZ2O6IBF5g3NfAwxQXVnJOokp
DLiWU8RomLoYiqJu12VfiK96dvX7AD/jM2UP3Ne2DAnMq1F0ACL+BjDmMwvL3bU/XLjodwO03b4Z
cnv8vj+RgI7mz89nluX/j29PYMmxra7qY9ngpFq8kKdKh37w/m0xufKq2AS/ZwtE02syq9QuVVix
lAq0PY5d0wwWulGWcmdEwDgWNVJRL/iFvtLj2NdKGcTAtIithjCVmoEcAkRHCSJjqNjyLNKwBrJJ
5GkBRVNaE12fbVGinq9BV8rS++2UPfmzPfgwX7joeEPKyH/gRZQpUhKBRSKjAb+5VBizaZNHe1uc
tKin5VZmFnu18yK6GZEN1PlfFrG7l9GtmeMlkKUKvynCt7xGoSfzgKnvroRPTfexG8JvYflUU9Zr
JVPFaLkKe3mpcK1I8YYae7FLEw10Gz0ssonTc+j9rHkjg8P+uAwwo/LL8o+8bKqBaAIFqlwxUHXC
Q2ZdmLDrA7O7NqVddSiMNYzCOF12JbMRYDYhBey6Q7ilUq9UG8f8RhQd/1wy6GhCge1jatfDvAH+
Yi9JHyQgr3PfbTyOasNN0TRZJYc0bGWO/da82mXlMYqDLESZSflNEGQjKwYy1gQVG2j9rlQ5TEl9
0rszHUkHUoo/qGAN124CQ/89d4b3EVW+XGWlDj3tohLDXa9rCu3+nRqTUG2pfJXG5J5XoF0z+XLR
sMaGecfBq3QkWb2xzWeNcIcOGVuAGOpeTxwKtd0QkYQgsfqae0eKUGFE09V3WpZOYw2IwzlFQ5vE
DVDHsvfgJnoPuLsFY/GzxVOXprUgfcaVHUh1149j8F0fS+PTI6o/UI0+qypQa0j2VDdjv0Ju1kqM
AzSDWpLLZHTXxMws3pIj/YDCaPgtrEwLNfLIIYCbrJJ1lohzJVbIhmopr+pqKkU/VY7aJGwuS5H+
3nDnvQGvxM8El6Lmsf+mH3yKvORElDGMRtt1xhISf6nNkAQJI9w0iaGeLBnS8QgzgWbN60tyJj/I
oL2u4QnWqXl9Z8MAgaZfyLFVHkw1wbeyctBphIiEVaK50bsV3MhBT7qdjxmireApinGRwGelD5H7
fi0H9rbUju7qEBm6yosqyjJaf6phYfX9HJnmjVMswmx7xJ7t+tcnle5zCB9lSlG9yjNnfz8r0sLH
5CNwWoeKC1WOpu+MbvjuU+YYS6irCC1KVDSSlsbuDlYnUOV1CgynU7BFJamlUrm2NBTUbtm52juG
eFLXiY8/tLXe/uAwgsQmtOTXUh+MTt7X/5PkBgs6j5hAKTeEAoB3UWsoXyji0Y2sNMuWxhnwXGgV
NQf+CBK1hvQwoQBnj/EzkGZVC08kNhbCK63OTRnPFetHsypoamxZzhBHFQwevtQUI7RlAbcZv1EX
53q1u8pWyxM2pKq+o8GR6k8/wfrV+5wsm8vyI4ACFzKfss3zgECYU2ow8SYddMYgnw9DZml+3dMR
TCLahRwurECxFJuHfpW673sFUnQtc71GVlXOu1az30yKQYSxCUBbprfmc8GjBGiCKo2tzoIB+aF4
WIpF56WXrqJSxe0J5iDpUEvzEu/z0/myWmyxj2LkVbM3G3qb/24UuFGHL/8z2gB7P5c+t5sIiaET
m+kK7HvNDNvXnvm0co+aMPH4VKBivyrriPfc3qxl4Y9cbzlrSBK81zOokLrm7yEctuQG9yMow9DX
XlKX8BFEeZVg5eJ4+pdG6f0B/axy/oUk4jdDiuLFxyRQCXTUXzuusU3NCODjnCTdlI0Iytf4KSDn
S3jGtXRukj1kGdiYXaPKiWo8N0MbCIGJWsrNLR7Th+aLN90uuYX6qx1mU08ep4oFkQalOHWgq3Y6
hzM+by+aL3Q76nrJ7zwaD6AHl+8DpZtkVzJlGuE1s08DFps8TVdXcetFxoHw2hf15xUOdVccPqVq
ihZUJBMMEHAi0QrxeYiUeBwp3adsWe8OyEXe1t6xd3fhalttOhrkVTMyuWttO8Nl4yCPhuAG2hjs
bS14MF5dwIxAvalMcjnRwhc5ZtIPP/H23MBNw47ckgmyGnYPtN3qSoc/JpKcZCxaKzr5uvW03V0/
D7WP1eU4YbvT4M1ml1T5lIr/uwu5sUtFRDlCuPSVM3UK/0ypQo6brR5bxiIiubFmN7YLWZ/h3lnu
DUJgW1T9zaYdU6+kvuwE5XlfBfz6ml/qPwelB6CfGlZAcyxa88kF40MweeOaX25yiyWS5DJrVa9E
AGmexLYVZw1nh8OQELbjnVBEuMcl89nuGQYKGMncCuBCMT3qIk9HTivdKS58fsJhE/gvIb61uLVI
2u9U8NztzDTkGJaIWvjA0mWVZlV2AqZM/UMXr8mbr3GnqYCC1bHRlcJuyl3+3AGnkTXCckpZx2bG
U2TwleDk/2VSQJG1BkYASlCIBA7lbqC9gDLfvvxXyxFC7RWgOV3TlZUN668dh90jqFpwfENS6ash
jO0aqpa3aBPyi2I6+ON88W3Znw2aGgkNQAuNK1JGwMIoT7RqMi+YwZ0AgdjI0ROCcwHhZpri3Ge5
HubocAjUqhjvvKePXQqlSQkrm7wPvy/bSaZTHdBt2txsACagRlU9+nVmuAetn1DqX7Mr3cE5mpCZ
uH4X9dqlLHc11B5X0j47kq5Y7Jk/FPZRqh8B8spUgrMNMvRjvInrlTlSEGTuSp+wsnx3yLMWqD5h
66AJScUV0ijJw5PDjYa0j1pcPCrpJFAxEDkiInDBucUJbwK+qtoy3seoymTUsknfJ6JsBA+kaV0r
7U43kEhgcb8NPux0kJAJfvZwdKpo1E5S95RUIXdhOjHwIx91A4PejWjOqha7P+3rnD4xHQ8XFKFD
IJUNB9bsHhzgJ8JiEem3rPOZqUMsp+Pc+NQ4UVgIbw57NPu3kzRdvALkXKGueUkOETkXM/ib+2TT
C5ml7P3ZFJd/bQnCLlW/g8GUljv4yXLqUDdLtjMQnG+rs03o4fXzQi4susOLIzYn6kCVoxB9L9Pp
mBJS6XsRUg5cLFh8Y9H87bNKWRa/hBxEAHO6IpGRxgO7yHVBq8Wtvh60DvkRm/Mj8v1SdxBWyh4k
E7NnqWZT2Zb+SGnscxCkKVmKrVMZ3VoCZH+QgmvMUuMOcRqSkwMkwNDnyUTu/NDG5p2J+P5hKZVz
BY97MpVOPArrBAwJAh2scx3QquHn7T1Hx7D8LxhuJsakmDdUuWeI4DUeEKwU81hljKrj9B4nBEic
dWoRjFh2Hqs9r9HHjBEqYTRx07LkES2ju5WRQH8vh5S8lpXubk//KrFkXF5yDacNGj9coTnC3M1n
QqFmCD0JO0i1QeGw1FXG/Q1u7DbXwEcCWihgcQOEfMTUwCI3jwpEusvPe2Z1BIjqJB0cZyhoitIE
+5vpLXTNXvSSB5HWogVa803OpbC33VZf5+9WU5Vr0XsyoxjkT/EUC0BL+4Va6ki9rKLMqvceWuj6
XZSQp9lU8ksw0m2TBKeMr0iH7T0sruxbh32gwMT5TCbnIHICWHtPbZGJ/lyHqZ7mkFgEr5eBOC/a
046ot/lFNVB+ZZElG3qH0uwdPoHq7q19cWtvHJTaamILOZCxL9gvR2tTTtwRP9kfGjIVMWPSrhZb
G6Kk29gpK5DCCRRG+4sZz5mG7bLtubP9WkhuhLRwzK8BsSvD7MDt8n5rWmGpULIDm0bp0Xo68uT7
Cij64KbpJokCvRIUES97FVMlrgf5N0eBgkFovV7sjG7q5H+FqplhWmyjCItSIepltgF8JtcssRB0
GfadwU2ncMJqteLuJ7c180iCBr3wr0fBBfu4hOIsI4zGgJEtosVSk7PgXZXkkiuhxi+jABrjsLN4
230nrvyoKYF9JI0lrQfW6dT4HXpDgFz7WSqQGqtIl+GsfyyBB+4o5C1hTJmgqH2XLCi1xyFaBGXH
9wsCc0wHYQx9XI2N+MekA0TL5RSeJeMy/lAY1nU70vLkEOebUBjt9Zr4r+SnCj4winouPd/w6qrs
aTzMd0npgOaSPBWQf2qmbzRNt05q0pUo4PcYGwp/CPGMBSUTb4lGAkPB23wrTPfNfmWx/u8BKU8x
9oL91h9Rx/c9TtQQiCQTJQWyIpZ6i99ptopCXrJZZjnxQDZdHZ6/CMbuia0pXPRoGk95+9esryUb
MkZ3Rw7w8Y6OvPfTvuo6HxsF50ntx9sISHQQGRlWriKyYLeVC4ZjdAjT/SGs0wlPIziEoYulqTiQ
7EUdqiPCufbL37QyC1lWeN6lPpYppqXbVuUWz4e8Xq9A3ZE1CYNQtU5BV0vrBVBKHVrmZUWR+Td/
iQHBVKIey4iPWHZ6dl5+1d2pakVYTbZuy5bhSrPZBN42T1Epspe/UcPYMIMLHITObrTTQ3RI4ZzV
JgGp0EMZZ5vvAHGyokI1M/4vx+PudFGXDp6eDx3A2r9B4u1+HwCFN3rN/IorQ2m07ihQ3GWiTUyM
mPKP2Uge8bLEua4nQKlAngh3ORF6/kS/wwF0eUnlxm9sKxCkp0LPk6YO+z1jQmW9RWkagfPCIbLo
ro1HvQ9VL1ObEUtzqm/7BtfYuOsMOeoCIrUD/J2IJdkyFkuHjzkHpYBiTMuzCeoWcNPuvkBSKGsT
92wTKXo8RxyWu1yCCGgY9KwTlti43avJS1FUNBbmXtt5UfIJoy/OyQ61kS7zSFojwAdMtBn5htxe
32g0Bwr5ZMvxFWtMOhS7LeUh9FlaSc2irRVPfO/9iqis4vaZwo6d09TScfJM4NgRMbK5WSfsyHTk
AkTdZcpQRAwTQo777yglaRQZ9FefyBBLNdufmVVkRQ8xrt27DFo3TxqcGoYN400YMQeLAvWq7umx
1jd+21eqMO3h1zkfLL1SSodKAwDFLrt0OZRgIH2aQH9zMLphH4XWmH4jBj20OWwPIlFa+CFRKBlo
/m9rNSM5yR49oVDhvEzT+38w4Srd2vIjrqsZgBFGkhlFv2KEySn2QHvWXP/AJp+f4SXJAPLefaPj
nzZIJrRhEAZ+NKu+9LXdiGCERHmCyHSq+nt80xCKn5yY96toRl8pFmLR48NratcKEZy9JG7Il/sG
nHUF/i/mt7mxmkJ0ujOjQqfxLlucXQ8dezg2XXhm0dc7D4oZbNHsiF//TsFRrnix05hInpT6vUh9
FM+7jC5rysLztcC8/1xqjxTPhe4kg9Io2MvXEP5OnKBT4lp6KKPKChUEN1FBt9U+4zNeEIjmZT3A
ZzTq8fDJ0VGv/No0MPz3BAb3C2QuOgtDhq9Ckb3JiQ7vAjalGTCv0YkWzpT7gsJowjaZDHl3yG/+
sa4KxLhXiUkSBrs5TXo0mZc+FHbRP9vwjqB6wAC6daq4LtVc5MKkrblL28l0EZSdsKg4w0QhrgPZ
aRD8iUho+kcQWR2T9HIZmnunOTUIGAUuaQsuoq4KHqBVM4TVeEWtGZOrdLuo+z/O9QFPlxNnm696
KPaoOENE9TciGc5LhTm2EXqaIBg6g47CMuv0cb3Kw5Z81NRxkRqPYgJbsjdnjYU+s9of5OzsHVR9
h/b+F4SJgeYOJvw65/Kpir1YPFz3SWRSxwPw+feZ6Amhiz8BlJJ6OJ0OzszTYZ59gMfEhiXaQh79
tqpO5ptWefY3mnXebZyfmYNiz0IlvWGp2A57oNoYBzV8bqMtXt9PwqoEKBA6y+T+jdXRKJ9M2JFJ
cSgCFhc+TSnsrJ4z0QEpqF9BTWcW7ZSJOD5+PuPS/1F+lXxRuNy6sN4iXN0Kc7r3dGQDuS2aE/71
W5cEEHO65ZxvedY3G0HSy7jaao7097VGsYcm1GefwrsT04fetZbzspjTswfTchOiJsrBxo/bmEGl
l8kqb3TXc0orY0IhBphyEBIjgpzVbcAQ9lFEODJOpKKWBO8S6/IyqWPZO1GhI2qzpHOIzEe3t6/Q
Qoqg+BUd9Zbuam6Pw1/ZVAljQY3lQzAEeuPIUuVnRzH4b7AQOc1d3wR2Si4IqYrlLuDJOLyMZVkt
cjizWE78tp729wXnRrqpGXNFHyu6E/hrIF4uwmHyYJfzDS1Z8iAmRniGEIeKylbmKtJ+QqFjIjm9
wn/4G2LzayBZDaglY+hhzpWdiDlAZYO6aAnBsFzvcQ2J8qMrRgjJTIyXnYGm5xKwgRUPB5Eq0pk2
iI4usdnQfckayDVmyCyeSFnFwzPJfkNz32XWTNTY92JyjnW+7QDDKMr5vHK2MFQS34U2aKYynuy3
zTIUmzcZwFTccdsqp2n5H9MV5EqBCNknz9gjSW8NlO3fuqemXicHNKZj8HyO8LrC7YWGAoRnk4D2
4J9fIWOpEMkxk+fdoim9P2mrlFTcjg5SYx2njZt5XmfT0KNuNY6jX3v7eb+9SXj8w1d4qa/pggDi
pZnwF0MUVpYKuPo1EWwpr2ljb7zFsc/ZudvUFldJiEYU5f1PVlayKQ/YfvpS0TU0ViBLKRrpygcl
povMx6rCWrtb7np/Zqa6RN7OiWRZP0fxuDFrvSTplWmLxLigVzXo91/Gg+ro/hS1pwB1cq6JO3oF
FNbGZDW8Zabgg/qiagflhlzfatSP6wW1p74wU/s4rYi3tof8GUhFlprqvt5KYHN4Bj3cWZoRs1Va
tCxVoItLL1+0q33IXt2Ax6YVotnVWR1M0X8mV0SSnSPp7EuQ4u2vj88G2nYczerjJXosL9Z3DAMU
BW3e8J/bA4heL8yckpnIKGefcdJ14viRPq7MMOPYGPW1HBkw4uP4ShD7GWLQLcZ3+1KbnOmx/tDz
PwsX4spD4NILJkD7TkNUPoVJN+amyTqKuf1bYGbiyz/AM/4e4oBQBL9lCqMl0PKov7zG+DX+UGK/
ULs3V//eIh2HDPl1pYRS/F3D+K9Fz4Ys38JTBX2kDvvVaPzP5/DScu7LA7j5ylhPHKALu/Aob2Vk
jZH1bHiIQNtyIBh6NQvLUAeV9a9lDwNkU9fUVXRk1iS23CeeEXtDY1Z6z7wxuXNlVFsbjslfovpu
/cOs8amVbh6OH25/SMW8RktY4kXRFQpEMQlk0ZN3vuyFePnLsW1mPK2SeYOdnLVmTszbD3Se+38d
wI2IAOp3aUltCqlV1awyYiM32i+bCIA8+G/8t1irPbjd9rbYhFUaOjcW0huFxGW0OwjHMuEqMvHp
1/ecOn3tpeDVMhIvA4G4Va317x0vsA81c7cguC6pPC911o7kdhtmxY+3II+SvgOIf9wAuv2bFD0G
QIuvEOm+MVnkxrcJ11q/akjJBWjhVTSI30u4Oo3wVB1xBB1uQcRo/WH2EnPChBKPlVH9MAmvJT80
cUgahkOYc9EqBnNBSFjqLJgSdqZy4vteEmxhyUOSKhKD7Rqv0rSzLtQ6ZVqDg88Yp2Fo8FLi0Hcn
VPIrAGXgl0ymuHbUx0XhH9pDuNbSRws9ruf4WNvJbo0OT2Aj8gKd3oQ+m/+gNlhQGueWXuyGVbYX
l7ChhBLqtnPciDV2Z2XvCKfe81UrVvtcHa8loxI7tf1NXjyTf4ie6ULS04lbo04uDrrnuI/s7vXj
EBx7oWyOdmiqBKbefeSlx8jZtYajAiRnm0yxH3kb90Q0P4mmjKUJb46Me0XGYTdWqbSKaf9sfw+I
aSLmI1Xt6b+Z7ATNv1kKrGPKRFeMtmN2vViTP3tg8fjXuCp29sKHhKAIs0SP+ad/Z3p9MdQF/oEO
Jt3hZebah+0ZIKk7eCRE7NUD2qGAi6W+gDD6po1VLs6cDpk/c01VnJZU2H/p6IdFHNRh+VhC+n+I
3Num3nWf8bkbQflItGP/NkAuN7Iq5MxfFXg0yr/pH9sNwW25iqM7H4hRaBgWNiCA3JuertLPtlCE
7T2SEgKL1LdVNpwHSmwimqpHfyl6qR9CBXUM9tTvd03bPcpcc7jqcwQ2vQiFfwi7s7FH5gjgGN4S
m4eKkXkfebhhnJaEZOa6GAdOzCzUwDENGYUsNS0N5pvl9rUPlwR6TCY6hHaLpUv5mHr72gdyzqX+
SeR6S7LGhh4Wn3Oo1TZ9fz0oS9WEjDvnbKhhaabEf6Nyd4ef/nW3gL8Ci8KjayNoZ6ewKkNZxokl
kj8QJ3kF58P5ECkH318sKx33jhXGOYw3T4v7aUw016tN6sjsP5OmSF1w8J7eihb0gvBTGLrCxY4U
c1sIs8EHZOTsK9t/x+KvqHWD5rogyPmEUtyFtuO7FMMuEkqEvyg10Tb5G7Xfo/M7YOdrlI9APrbz
lDpK0UTQNM1cvyrFMVGEJkxWwh+a6GMxOgIw1HrWnY/qlJM9CkvZmDTH4Hr7TjIIEsAt45lbbjwA
lnpwryaL6Z/isEHnay8kPFGi9LJsy5p/+j4VpEt06YZdZJA3Z8nSLWw+nkSvgdbm0M2FMMOCQ022
AA2EqYaZ4BG22COYf27wjrpCrk/sMC0qF/om9iHVTePwe/zgxlPW5k90Kwo/158OhJYLOV8GNjo8
fAo7i/QKIQ7iNnNvxeNUVKHhhZ0JOPBFjEKR/ojsJ/wtEFbCMmclu0lH9uIH3X3iNq7Yg/Kvj5RS
Dls7gq6AcrXyq8Kya+KLCb/Aa/+ayg7oHJ8P2GcKbcVmQeDM/TpUTga5SWYiZlIsZpEYzVzMxzl9
jlkcgdcKUEgy6GAh573OFL1i0wldgS2i4V3ztXPkbOt9CRifq6NrOG3EB1Mm7v2bQv2W1SL2qXlw
TUhmW/KihiefkkZmHTs7xU21p0jnVTdEaz6mDHEdhJZd2/wM6yvNGheOWwihHvUyV53n0j6FTi/g
IPeGMUYk5u4vXKYD6s+V9SwUi/kqrENzDGEEhY1ViDe64tqQIOBmeUky7FOChUQsunqbqC+DFL79
cADB2BAQ1oWa/A83wFP/6ijizmw+TGA4WlcBCkcl60QyjXAHHfGdAXUsTODNDE/aIKP6mDFWmrDG
A7IMUAHIa8CIQSyqbJhcjCBr34LbBh3HQSGb8LKMeMd6JDvdgFg4RYkkrguRZKz8oDOxLo8UYDWb
MqqsKscNuzuUpPRO73zFa3xeH9SkUnSkahhX1dt2Q48CV0hMP0ROTbUBDWcZ+M0kiRD3eGT9Iboz
OqOalYcjKVvmQND4acCqu9Ocvx7HznaImEXtJamVYCQZb3qiSqEvHBr2gxIRZjvQki14D1fehZJv
uTOz3pUWltUAjzcPztN4GyFsR86Vnxlas8lkiJkSiv6Mzu5u+9NteRNDmibVS9bjbn/ksMrAQCz6
eostwsK6N921q9j3kh3xMhAs5KIJVUudirkg0gPiM5Y/Qjnr3VLQbr8ME2BVujyM0ABSmW50gfuX
q33b57RhkhI9mFrOI0rViB+sej4E+4nIJdV9W44LuOogRDsmsfSN8BMrvMfrZy23VYS/IJUD+fGT
w79mCLEf+B0UG/cMxWpqTF6T8XBz14Fiajw3awyhibT7uof8YIKkG7gmb+pXE8HC7xyCXZb4IFbw
geiVKYhjHxusEakQD2I4lgiSQlleYYjGpWz4rlB/mqnunAAcHNGN63V+4qgoqGZtf5/gtglAehml
+N6DzYXVApOWTVxIbqGbDXIXR/fz9t6oX6vh9vPKV0oD4DuJst0vaN+w1+I1Nr7kvglDcAm4ISXc
NTLeVIAzg61qGAptWGp9Fe4y7Mbae/CuhaHiBoGOgcb6dmRh/BXuvwODe+k0gMX2Pwp/fTEgus3c
PhS4MlI7wOsxaGafSemxlhyt5YVh+eS2WFb3iLTMXVLREX7/silMtmazUa2+yvvKRMPUkaS382bt
X2sENESuoTay5lFWDbjW1RcEDKonMU2q9UQv4kN1sbK3GBp4yywYe2S6tJkMs9YDnFacCjQGyI8z
Y36O79GnBpqTk4nvu+g87AqY01MTi/DBjtum7YEx0EKSkSWgU3BJ3HTVgJFKQvlVyvd80OVrppH/
75ntQi6MmvwfUvOToN3xmP+qlzy/mRTEdf2uUyE0wr+CwYmKUwXL7PqnQuhFp/8kcZU1k+7bEhgK
YJj9zffyXF3wN4MekhPh2aF4CCr8anzF59i6uMlYHrdIKu6hBhYDOBYW4dTbhFfqKkbsqtauqGpA
AaStOr5x6KY6GU8u5ZvGcK90gsJOxa24zXAakEUi4lAl38h8fnlQjg//OI3xLkF92/BBayGVB2Q/
c9TZmfQXarG4kyZm7uoQnz/cP3tOE8NjDHXjknIXMzl41+bVApzr5hRnw7lW0Esbiydiefp4KgIQ
TuBaAYB9gU2JQ+JJse7VVCT2DM3gtz9uN8rRCFf/UEhKG7AOvBdpJ6H3YVVpZyMeHGbTF/VcVw1z
AplajI8XbvHVLksWIfV40B6nJl2+r0x/1rp42h3PAvb2hMFkUSSCgq4o2/omocn4zoiVVLsjPfTP
EhUL0m3CNIuhrwO/ukNMhS2AwdukeybscDh1hNB/i26Z5DGgFY9pwxa5F/wkQ46C73ahtUptfXm8
p0l6Ct70/nUNOOrDupmPU8b1kipyduJ52kWMwyw8bIkTgXPz9MaVNj2OZ89CjFoHpoSY0sFmRE1s
bFdyp3dUf9TbqBVBS+aMSD3hkhYCPDaPd2pBQK022LGlaD2HPjcScd91vHBHP1QpRvuRgr+atrhs
lAfmlZEBizvBB/LGCAsJpSgCuOCoGzcs1OvXIY/Pwp5LDJS62eN1vXzu0M5Fg0YQBVj315P1dqb3
3IpvZhHzpuQkrZBgIyDoOxAwcMWfGmyBC+Lu4MNZa/XKmlbF+lpm8vH1xr5esamdTp7APrch6jk6
Ml5v/QdOMjCFNJYo6p5aYa7imeMBemFST7RgsgFO2aurbemfOZUl/6UkdKCeJiIkSmva7Mtw6dxC
JoKfT/BmYugqP0mwaMH3decizWnOtQR9vdZnojZcr/JgNTDEC9MuACzipTRCAKinxGrMAaj73Yfp
vp6FixBon+AhtjWCxsDkD2EcnG/NOV8+q1fvEQ3/TjHlXXRD4TjF09QvppGQFoDgzVRNIM3LydKy
oCI4mwhj0M0eTqS6CksCvgnq2wkWdDm/KjEYIQaGUNPeLNfnFIgLrJv2xz/b+1imSv09AYRPGSSl
y1971H+xd3S+N2Khi50a4aZrs7m73RwbU4srYmYw3k8ry9LAgpKJ8rv05jLl13pDh7S6lWdb6tzz
tAvBdgPKwPvjUnre52S6//iZ3GH1FN+0C0kpf9ZcMA79Bu2WpWWrPtyAjPOSlkoDARFLXJEJRyyJ
jGBdRoSyFqrrXRWM2ZWPBDwX3NwGgOguxeSpAd68mEfqx5Zx+u0TTInCcYq+Di/SozwZilWiMdx6
f0QY0ShIEwrcDVm9FCaabAaDKCWJD54s9H7xFE7jVjQaXN4JNyfduRdNRwKHuRTxhd9kAUT11A+W
kVHoCk7YHQXUDLF5HiD5k0AL6sQ5dCLWVsw1FdaDdu9wDfnRj92TIMnSElg10ZNqdEhpkEHhP6p8
ohLoFrBKPkV62icYYOHZdxY6K8/M72nDaF+AT3FKzHydDkjuID3v7/rtZ+MMZd9TYkxoKYtROiEm
8PXEJBvgb4K+jZQQlcpTVpcKDF5UKlU7MBT8I305C9j3LG2FQjEn6YWyWrS/EKsHM5p1oJmk2LTV
tbBFfGuttfYwESQ6i9XUTTO0Ljk7yN1NKqF+gNxu11W/SonRG4U0AtBpwyZLbdDTYBBMgG5Bjvll
kkNqhHmIGn9kOkhDwMn1LfmkcuUP8vbuQs/h5tBXle5kM91enEcRxiz6T4NQrjvDZ6Gue1DxDDk5
Z0yWtoULzDRghJZvuNz0zuuJM+F7glA+1K6Z5FYkFEUDxw/SoCr478YciVho72sQ6LvA7QDfP+Wx
kczIpP9Nsy1ThSYHM594vBXKpg8vaKliRIKR+xlhXGqcxAOYymmlJSfqf83qLaA8DeRysTbc/RnJ
9fzhDqt3VNyM2xo1l8t7N6qItCerKOThW1wgLbNSac8oJPM0HM3St1BV9SgmfQkjteaIWGYQhNBe
kkxUNPH8viERIIZTPgEtBmlzOFdS/gLa2kgZ0Fjf3LLtt8YeYqDgBkjPj39zwCAX04tp4BQ1UcDs
OKz1NkDaPoKSpyJcp28Mk0xNe1gYHlyA94AaLOs+9Vsfu0BFnXBuuS2x+DOyvx3GpACBijD2jApc
tyhjub2ymEpmeJRC7U3zgxQZWdkWvgX3iwPDAFtRsuFvWQeSaWOW846Rhx0+jyw7PfB82OHZRMtT
k31jWhOj8OINVf/mib6YbvV3hfwZHaGr2zrtewFZYPJJa3r/Ji81tRtVCEFK/iX/hLTdWLQ0Prgn
+GgdecUHQVlhiaif9772TNWe0ZjKC0+uj5tQktCJJuvbCPG2B+d1Sdba4ZXcTTJt1i1IysGAW+Yg
X8S4uNADXskzgP0vh2AHaFoQ2zs0rIpJK+pVp2lhtAhp1zpv0r49TUsyN/znlEeoATl/zENblQHT
RlOx4CeugOc3LN88W2EevrgkYbZo7C4AqcqlPnApVGXAI7jFrAYlMNC0W2FziWln6iE7Zflhluy1
bOsNxdDEiA850IGM9dCX+yJ941dV2e7PrBPR3UXv9/JV27sEsqnMdOZIj3tsy6bJahAs7WBsN+wF
UHywnN1d7ghlk5nx1fkMklobAMmBucwrKQ6DaB9BS6mdw53ZasDAmic6Jmg5Ee1TmE9YNmF4OEMP
Tfxr3Veeg+cqGd8NEztdo8oxuKP2bDcMqyTgzsQvyNh1zdX33EVoTBCEqbM0zjSRs05K1xJU8bDv
454ctM+AHCO0c8eZGDY+a1Cwdy2YMaWtNmpn/uGXq8KDe8qeMXD2BNbKUORnBJXyKp9Vg/seNKlB
K6gbWMSC1uVG7Fp7/f/W53ucfSlOcvwiKSzJ95gXCaHUTCv4C1pIowGaitZjiIA5e4yndMDX1VVT
AfMWvEUadoplwXxz2aCV+baU7nKuizgkwPuNjVbs12jeCEaP3Cw9EAspYAsQZxAIt0WgMb8BmnBs
RF4CbJUKrjBlqI7LZDmkRzbHcg+llMwWzTPpeyOtxlgWsMPCtC+vwop9RHAvUdbRQ3Nnxnum4/+W
zCPD8OcgyLh0IxuTGxpB+VxTfwX52eE5ywNzLKLzGFE3piTajcMa2K3oa6WUt5XKk7PsXOkcnYAj
2FKXB307BsYMyFWMDATDteFjfayr65j79k//BrW6AsEO5F52LVbedjTe7S/IcuBQvmW/Emve131h
HCa9QBnpWW0Tfr7HoTf9oj2IuR7bkUPWZpbQA5lSPh1KxnxkhEOoT9kh6vRPnR5SGJL/PZSUUDY/
TtZrxndsr6tad2WdptbFOVy3QfEP8sPd+vsR1NniLlUQlbgeuMkABwkN7zIGIGJj5LnKsB8YH0xA
yfdQ+qyA/CGH1GgSz2UuXMJFgC1pd3ByIWq7/84ptMJgqtfo4/uhtIecnTeaOoeSV3VefrJCKpdA
izjyN+1wgLdwkAeAooNv+DbfM3l0sdVIxTxtJyTVuM9n0s0763e4TigoDMXpL4PQDLiXcGT84iDk
ieqvJDDaAZ3uzRuMUNgxLfAr1teidGXXuZGNsnGQgcGvhxJskWpq8gvsJRC+8hxg+fbqt6uBYhhk
JsCfc0816FOVa6LNU+NE1HYdAn2sTLYLyYBixAi01uJ4+RUupp9jlTpUGMQI1JXOSBU43lGv0haf
qAvrqiUQsDCHbTQFweY9L72HEtQ0jo33EoCTKcdB6jZENl9y5789swIwPhVtsZI0+0q0OgqLvF/b
xJZm37zpGiH9bLSU5U0oVbN9C2qQwT9o0M1xoNfYlZ2rC4NSSe8gkIc3yNybJPg6TRQOfqWLzQBW
GqgBy4htIX91X8gsxNROJNmHjq1VrB/8Rz5UE5TL6uoqwfu5UQK7L3kUOw33sL6MuU2MBDCnT51O
LqHiNidsbvLpFiD5fKeGWb6i5LnpaLfYxJA4KEy9WR23kwkWD4siGdVJ8VxZrrkqB3SjhpLiml1D
Cle9jxmTOMZ7QskUEct7tFN1VKS5JFGWodvMy1EH3VcO06bUX4gt077pOFdQmiWUrdRdAlUDOfJW
A5ASEzH4blsg3d63ryrMKj4Tb1EBC1AhDE1nDMWosd1dPJEgdaVtRh3Wn/ug2mBDkWJRNBykTNDG
u3iyH6w9rb4jxoZRSgUcYC/6p7LVENGKdS0uHBtQ+sCyw+OMvqJBLYj3bPd0B9Z3Xhlo2wC/Oavr
JvMDVzlmMbSQOlHFaycnT5WU6SsEgulrqevw2WRbmqCZORK+bongsyodE8z1unu+zAirBYtwtzrT
wQbkRKEXjuzKBCajqARfIJc/xNaFUQ1X2X569fx1YYsxO5tx5hmVFqCd3HGIuCyaIDeAEgPqhv6y
cBe6Nr627VPca2CSWFY9ryybiKS2fruLMC9UV5whTyO9asVmtA4lJrVzrm99CLxacZm9k2bC2atZ
q6iqw0t3+MQ+C3qu7gO+5bU2WEYqv1yjaCFshOCBgD2+tuahU1Obj5lBSpAhNlQvZEnUJpL//ViF
Qz6hmfX+aOQethY08O7tlkYvDp+ku6jnqRgwxTmitdbeC2jox2jsomQ+DniHAEDHN+l7c+he4TgD
cpqeYVKEyFcRYrx7/mXaieAyyqO+nTmV0FpwS42Q23X6K2HizcS8OgZA7Kjuss6BSNwmi5ftL8vO
rRp+RVmbMcSE5oKaO7p7zNp4fvFVgevaQlsFo9xMEtVT3qDoCgaOHgv+mDTIg2Oi0NnktAGkFiTq
hhBAlWtlYXZjznu+c2aoAaklPQOTGF4W7Lps/JvVfghRtJXKObYrp2hCNBaAgQzlkBH+n6oSrf+U
FXVDhjYoXEnKm+9mQ06Wu+CEI5sF3YeFnLGtGwpSSwF+oqxhf9IyB/Pm7EvXjsjKPmZTl2qK5u7B
OOa54Qo8jkzvQEkk6IH39ERPtvIaYdcx7ftrYKNnYgsubKMVr90X/2FcwQCthshpCihf7iYIbyXr
/zTvhH4bmdyQa6eGsPsPPLNUlSkr1FKjFovDWL35BfvDK+6hg8yeLlkP1YjoH7bz+dsycTCetxJU
0WXHy4II/LXJweg8rV0/u79cV8hhl6xPwep8U+shC3mCvbgPoGSDMexTICv+77+CmyKldh6LHT/T
a+vSjdHi5fJlBgzCG7VoVkkGky0PvhYbud3b+ZWDe8IQGirVrXiTwWuXeYiBmDYW6b4KaqmPCQ4P
07L0IEFeBrvqsK0z2Xy5l+dO4QA47pIZFpVtAsY1Jng68ksyQcEAW04cRD5YvKFwsnideUINTHrS
wB1HSfB/6kShfIbKIlx3IyCyvMBFyIgoaqNG5IkP5hxT/ljJcxUCIW7j7Ew2sgOMoBLdWrOnIvGt
cwDTiekSXd/CIaXk5VVEfJ/iU/TNA2uS/Q4h/u4sMjYz4bkbwt300eYpaLIIX2IBZa47xFtLlzE6
bYvuTOGDqNtOcaEYnYh1AwEppSZ4Uu7jCMR8phV5ieActm/MrWmDjMjaOdSOHOOqNdChC1nLarqe
XLHbOIWO1eG+vNfeBdQ8JGTupr7vXrR557aGJGRmzCOomSBYfRrYlVZ8rldERr31skBoKKqseJYE
V9BFo1Cb1qKnCQnrDQ981eKLHJCWvdB+dzdlo45ZI2QPAQmaQq+qYgY5NCR66G/gZI10Xn62836/
h9KrZH+AqOi6TiAPu0oZmYxwBML3h67wDN0eot9y6C/RONS+KBZkLHife+QpsqGOJbM1/Ib4qOu1
yqXP3HsRwpVf2UU7oMqWB7xlYLs+LOsFt5SX2vmtWpdRacF8bQlIyLY00TDmLAMp9z+bKpNRAjKy
5OGZe8KAtyh3T9FhkHycmTvT8+M5zEbMjfPA8wgy2CssYHglTCn35C+2f9u64uRwaLcALGTa1yT3
dMUHMsFLFSN5sWyUarmiSfYtVLsOSWK1JlzfTrShhOskgBNR6de/kKIRjEG6EW8p6ErW+pwYE6UX
5wbRdg0eP60V2WjS7HsvvtCxQ41E+b7EXegeLmhE/DXvJot5SMRn+I1qgpJODhCW+8IXxi2kX84f
ByI+G4BUrkI0FbyOxHm08SRMvzYUz28eHoNWu9iukEgq/tsAjQcuP/bVglOokhNJv3MHzWCkRkdj
M2c9FCJPGhmGH+I+bhHa4+IUEoQaawSmZm1FlZ11B7kT6IgeSkcMxhE435iiv08tuSBzbtoJQe8L
mlm2lI7OC7eNPiFMDFceyvU+rjUtbVItxgNY2/PJ//6b5ttoYoFwOwNugf897fm0wu5m+xG9SN5C
Lm0Fy/ghh/AtkExcewlPjlbZ2/y9ByRbX2uQFHjKAl3XsMKxjIE8lQ31+u9TwJQf98ul5CpCda3s
YdyEvFxjTmW4ebKe5vYpNfagftVEaUpDxX/hqqBV85sgNbo2J+3CZ53xYuvjqAsH7J622fqelJNk
c9Fm2cSbAB4AIvcRrzBDytgrGVwW7DiERIV5JD+oWEPGs4g4d/v6u0F+CI6p447Nfc5GgPjsPWiw
cTm+2bCuyi7W0fb65lXv0LN2CDf1dzBi5bgJZM0Wh7c4UyRLnJ+Jya0EOZinNZEFmgQS8ts+mxVw
bXTfFsWGIff07WmMsFOV784qpbXrtRiVBg+wQ6lADHYujkGHc5a1p/hxAkjFculHttlb1RqtWTL1
R2J7KU6PnJyi5lrWxmRbNIOqtLWE6D/Es8aa2/8vnp+40y2oJnu8YEpeMIR2AICwTOYm9WPz6FsX
roXN+IMl3B2dHQa//uMbVyQK5PgUR8c0Nj+sceo6gllBGVh0Usq1nxmC7BHM2SnOl0bqAulUHdBz
92IV230wFO0s49lO9QAUGoePt/fv9zuohg9M7rnW6Edcu4Q3CJkCUFLPZdzbDHqMIkdUz5AQ0wRm
wnmTYSDpZE0Bx9+ajxr5p5jFMi5NnshOsPPYlmEVcnPnPooITP4MUDc+ithtxNwsrlTV9l5R3cwp
+M3pdV8mKPX44zx+gNeQavp/MHNW+Z1QixQsDQFALwFdk92dkRVCcqZNmzG2uKliAGWUewkTSIcc
1g9eS48u4idpSFvBlEkN0an1mCC0ro2Y5tkyDH9J7A/zt99tMTescH0BkQt7x3WakUhLTT+QuM/v
9dG/pCwgx5N8aZtdPks44lK8Wr+aq3WanImi5iVZy3Te4rI4W7Uw5KdC4VcYBBvFKAoZObBMDu8T
67i5L/kWEbzy56IX7ovc9LsZR1HGHawm1BHy0sJmw5UpI6YGUzgHXB1Rx/uJigvWyraCXxhI74Td
JonK9WcG6UuWTgVsrXDvFESRJAOR68wYj27jQfHUCbFe1yCHinXXYCvM8O5/UFM0sWMS8HwvRS5a
DQhAgd8M76ulqooyur8ElcITzAE4txlpTTxQyGsgV7XilJI8H7WAt7n7cqOYAKMaSp/GiwHw24r2
DMjQi1tT0y5rmrupS5RPxlB0ft4Np3NK9aKoAKdIjFR64pMaEq1PAzxJEtaj7NmJxtCe1jejOD3f
W0thhxMpFti5NPXlWyeAZpEBXHXiWMPkwalfBveaaHbIoQeUB96SDqWfKT9ov4FP2N2cfPGcTdTg
Hyb744gIw67IOgTz6EXdMMdddcdLJUyKSPFp81bQwUAOPGS7SsEOdcXK+eIZtqA2yuGpKMIB5hYv
02JR4tqaQ1MEBQrTLkvCvFKskKw177eafrlxFXpsOnznSiPdZDoWQ1mG/84LSW+j3B2TF2/6ZNV9
vSYoUgNalf6ui3uMnk7F166AloDidSDzNAOy1QNUSfjtNZcV7etxrUVOESKYBQ3pmfvOvEWkBIvy
jcv4B5hCbFN/eAG4uInH8UkvgLvk8EtsP0lglDejuCO8Siy/fdapJw+6CN/P1/IJ5zqQQWGAUG6g
IYkl3iMxhvBIxo3Jb1HdYpu34dCrnLgWA0rACks5C4cRYQUxSv6EQRac0IhL3wP+QjV/KDwzGFxF
11OXlsp1mir17aKLD2HcyLWoaB/oEEGcsWF1dJdEtKKM6p8lG8PgDZWykWS9Ty0NDUkUmxaADWI3
zt8/Egsn/b23wP6vmim5IViO+5Ubf5tq+i53ZblDfnnBG/rwc5oLTjLXa6DufYv+TOBrPQsumuSr
j2yTYyYBDxd1seWnirpRfRxKG6ZuOty4N0ksdmZFooIXrbrQmniz4O8EQuVysVNlg565RHX3nOlc
VvO1zjqzvf1oUW0k472kL2172MXUgpQNAC7c0qwju53VAwp8PBE15YgA3Tgz+jLkYkVkBLl02svm
OKPvH0dFQ9A4cXm09FYrx4cgeLHN/ylhU1/4WLUyIuDNXXE73qVyreA2BNS0DywWwP1NKv+rozOL
h6qWlBC3H20Ac3x23h23JF/NERLyi/uYEpPEsIIT6wTX2H/0HCJS+8l7SaveIaU02LhG/Ebx6u9e
IwbuBYArT5Ax2l9WSaKjmLoS6W+UYlTr3I5U7VqFNTVDzwfxDf2qGp2OcOw1sq5HMpU+KUVw1pU7
hztq7x8SOUIxMPoTDAk13HbpfPcgE6w/gqoeMaIzvJCVOmGl9Lw1hZ/mEjolFz/Z0/cnxV+BIHNG
L7BzaHflZ11UsH1YfigUFScr0Nqs7VwZlaf8CQ7GtZX5jFPULg7x6kALxcQO+lvsYQYZEpuyNuPb
AUKNYGa+YGemVhZQi33QXpcChgITtHvFvfSNIGhP+arl1UA2GgnJ7PZ1rw7MK5oz8k6fl5TDOjLJ
VLGwz9syrdPh6q3LA3I2vzAIfkSQFIMNF1Lw/Ml5Nz4Sghtbbf5GapFcbwIp8CMC49Yq1iR4sH8t
g0UAud3mw3FJ8C3KMN9vbgeE9J469gyhsc+jcCGaJbm2VFr2J0lYR4houFqAW0ZCvp8et8MUGKhS
FxxCg9V6LKB2MT6JFgzYwcvaVDbOonrPAvs/D8ZtRV02hTsYYlEeoU6f7V+dwhmY6Zlpn9g0TMAF
TMUacxdttf97Mk+nVF4+NlP6FzZ1c33NGGsJoX6MoXU8wonZV57eDu3vfivUjWDPkAPQoiRZnO+z
xhD6hW1uiklg+HZTpdcf1YWz9L1DvacFWGJBGag2eeB/9RJXQQj+Q1n98U3v9EncAI9lRy0mmFac
9qFNAh9jGtz/Tp/93VwNtHtYwCt98ivn7pZUhE4PyPNwFMY5ivbFv+sl6pys5E01hLt3HKzq6GVE
vIVEvpJElxfZmjPBXQxbJ/kXS/0cv2cWUPuX5KSor3FnGd3y3WAytALdvD6UsxHzfW6HhI0Jqk/2
9XB2qlQblxw9NgJfda8Yz3/5HsZ0SaWcrWNygEcGorpCQk+2GUpC+ceU4Kxx7UbqE2gX2tDXblCp
uE6gtquYL/Vq59OjHC4IPAze3hP8wdHsCy4BORecQpeqt5U3n8KQbu36ZSjoSwH66iJmJturv8MB
p9FxiNek/Q66vzrJXxE+E8hQT4HR/8BRoJWhxVHmsSoq2s2vkbu9c1ghdwlruVTsM19HzrwVf5m4
P6fnQZetVjy58V+pJXYX8LLVxkQ3O3ZiWQZ63dsE3D1hwHHE5IAHisvFVbDfZPE2T6CjwJBN+SDG
3icRb39NYAhvv/Zqfpo+tKsT6kxwJSDMPmP1rt4nvt+be++qO7v5ZTkQkXd43ci+Fqop8CwLU/Up
hVSW7b8pGL9mGLPrEznuvl71k8mx6FlLDq2vmMDIJBO82k0b4zS6AN+6rWDwHk2MR21f2jjRJOUW
PUKxgTw1TAIem/x2wVI7vl7pbzAYnd4pMeX03/lnPxzwc1Fxh0my2DKMsib2eWHZDmuqTNmipcAi
fA27nnroHHWeYL1A1zOy3ocrtA1QOGG04//tiX95OMeHp3gwmCjeYs3PTawLZym0gwCJGkNrtXPX
GnfSAyouyPRuOvLBY3M6D8ewPFssQBhUkSEQGS/ZszOEnYi/hDcbA3rYL2Vgns7biPZmZ0RuCexe
1J9S3kzKmkXva1q7EsVw0GJgmL/wP/O/G1m0Olb20ifegGkXeikdof1aa6uMJ7CzCtHpMPPfcuuQ
8JqLeCc5BFXFZEmJhKYBadwaXTW+8De9x5hqXqEBYZrWILQARFIwo34aC4I+N7VNI2/UB4S93a38
+0ABdcqt5ABcs7WpZ6yGEsGqJd5VoppRqxnyuODjs1N0lQrrr+OHixTSXvOnNq4bkYQ3qAdyvftH
Nf6xgBEW+Olc940yAmcO2iPW+43M4JSN8DhO6bsMDHWG1iP78BnxV0TsQNwcdosM3INIsDhNXx3I
cBtVsyXiys/Nr7sz8FN4hT6SrcV0rv509Gib87x98fMYTFUv+2BIMASL8HZOhbaWWmff5ZjW8UMU
Lk7oWa976tNkU6a947iTfK9ppFd9/E6IVScv00CzJQBucetRSPmlj0NUtcIm2tR2DdLIZVwtGJPU
JCSWdshmjpijs3Rwd+ErzGIgMrcsXssm7CsXBsIQHVvwVanHPesE1/ZrZAdON56a/udiQs3L1p/E
0Ci0s4Wwlq6g1eO4+7j/Jz6zJuMd0VVvQ+w4M+dhQNn7Zqi/cIlE1EMBAjgNsPEMmCRbGU4hl4Fw
yidJRKI96DXcN4I7XawP92iBNFsOpDkHQVt0GrxMq197UVMPwau4qy3aCkt6+z78IbEuO/gpWqF2
q9GcBNWtTZcs+ie2/9OVRZIWepQ/BZtH7pWp8MoCSQ76yNBCQZQNQAGFM+WxxiXNs/w3Hd5EUO5p
+68aLnMTiOeAclolQYZakpFj4NJsVi8N5h9mFM73HPjJwUZ64Mb/qUU0bIdhnBLQ4ytL9d65sYW3
vjZ1vJiVoJWyzKIr2oIwOM8DHtcwilW2tOJ7wvzUWFgqH15JVjlVPFHuqCKAW5iKFap9pfoJnPR7
ofEc8fi4j5sK0eVD5xfbttqZNdYb/q7Z/Wb46fuMh0E4XVabciVem6V2mSbPkNmK7hB2D9NEwf9n
ofJYAMPtG9/pWYzpzkjE
`protect end_protected
