-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
ZHaxQH0ug5nEkb+sPLfJ5YU1YAcfPMN5T2awHfjdCaaKmwA2l/jvYlYaJPbl8b25zNE/jkW+5axz
7bHl1tjSZLOmC6C2FVCZBEX4zbRh3y4g+CLdw8wnBEdbNHXSxRQxfQEpYZfcFrFijVDNCwuLRKWx
lzFTzFCBcvalaUNXpqTpb67pgJlbBQMwpDKTpbhDtJfndLcNa3jqCgtxOegsYUk+uYaneXanHhm+
gOliUDeF9lRhpgaXnz6pxv2ieVB8CWRUTtIeL9rxYd4yobqTxtwqxxiI/pkR+mriHJCUYSwQOu9s
utMp0FEtJKJDobOQmukn8HHFSAAQJ+TRXYtPvA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 30528)
`protect data_block
xCSKlUVK3e2y72GjSryzurRYtmmZhr4E5AHSKprqyCR6d2ljKxg9VoIX4oySR1ef2spzBOsECOjq
jGi3vmPf3fFDLxs+I1GHS3VhGSV0MFotGdcZrPZurBnzq90p5H/nHZxfJI17jj94YQtpbuu+axI6
uG3WWRk3zpRlknF+2RRzKRhndKgLaYooN/BKpq96LRTnSeWUnbJ4vEyravVLfOjW26Eet3YORb3w
Vzw2VFMxFTJNXMUvKaWAbFaf8rZd8XTgvQEFMAdmEX35iL1EDv4IL70QuieE2Q95Y1na02M6p9W4
8N6Nc6f+cdiLiJZBpPa+KJejAG9/deh/3b66HmxQwr3MBMiG8tUULng7Pe0tto8Qz1MPXtiaNd3u
U3uMJgDPa9YXH/g2ho3C/KI1q+06MCBV23QSxoLeQzolKSOgS7PSiNgebSXQgVdEA2j/hmg1hRcB
1mf38lBGbldfFRetBPP6x4schz9cgteQSPeF+bg26pM/aZdIxY7Z4BODQsbI/slR9h0pBRVh3ywi
X34OkSXixl7CBUuV6b5IP9aia7C1/TFiIccpPKYtK/mX43DjDARNkj5LkhqrjFiu41MZlpKNx8D2
k7wyJ4fnqaQhVgsVQ2NI5iY3aZLao4jkfI083KqzUO759g1O8IYk1aYYvYhyacl0xVYeVgBd1UMK
pbyKrgNGcjj6DQcYX0eG3fjuawN7eKkn4HONE2sltyAYeUG2vrj9bSgog9YtClEnQTGXGvWly7r4
XvCJsACfmchokxwI9NbSjFQuVZ7CRjnsxB/kRoHvST6IEiC1zdc7rHKmAk1LZrCBIua1I5aPeF+T
9cZlUlZGRxWDoYL0cxCz+KesySTdD9Zck+VhqURqZrNCdsV0uHv+b2OAbnJNcgjQ73n+MZNCkhEI
31PiEo1LoFbnFoUsdN3y0VZ88Q3K+cK8HoihivcpXtCuulMxTMsxjp++hRUHCch+b/csBHb7HAf+
12wZC9cPzFj7s91/pll1HLDR4u+FUyyaFRPoL/uyFGvNxraAunJa3aukQN7CvYgmebO3bLZxZrw/
dOV921jINQqpzfTjzTHTkQ5B3ls7ZzGKONvt4MUMO9w7x0kXkig/1ignGQSJ9URVOO0BiUFO1zLt
mOyTQ39fSQpLzzQZdvoQBZwxJ802g8wSxJSLY4WGirPqEPqgcQQZ+tnzvqIijDxZUbvQAT8AUJ5y
dC5wKLvDkIc0rA7aN7QjB+sUo+sKigGw5dhY8nXvXvKU3wenBNSY5RApGt3VmKvK9lfWrlR56E+o
cdUfB1ZVpJTOjU3ymZgTawm18ILArRSGIdSJa6W0pkb7NftAgjfA7DCgAv+JvK0pwFjkS2ByNGxS
ql28LYOEOXUjmmxu83tTfHVkKTs11LwLiKPWvqQim4Nvu1eDpke+kw9fuYejap+Q3X4qiQPZbFfe
TFDq8gHTVkrQI2vspRpaclN343a9E/DQ9KgB8BJPXuEJwniedQDX7dqoeiEQk/79lqM/8pY9/DNS
Lz5CdmuZ4iK8nNE027sHSy51Oh2RIL/mwfk+xXtQGHV7YQOfS6REvn2wktCs8MxRZ1a5mjaxLz4b
/c3cPY6Vm/fNIU+H8ocZ30tH4l3QfyMgGAewVoPYYh5t5gccZLWwd9jdVnhS8kLudO1Un3eb08nA
WLe4LvJz6+tNgEJCwokRGWg/ucFrLgmUcwPf1wLIwbkoHwZLpEFdZhrN2CzghdjKshVRTV52ugOB
PajKWsqDOSk1ZSBYj2TXOML+xpwWOhHhk2u7ZJI72OvweR9E+vOs7YRDXv6tNbdxlnwH9sTSwVzB
3UogrphrxmWLDwBjyz7LXG6BxtqMhGVtalk10zeCPGm6l750Wepfb+/NqgeEWTQBrM/rtBiPaJPz
Y/Bur62acpJhDja/HBua5pS/DnCMJ+V8ITdioiQTo2CtRQUm5HyOgbHJlm4pHeiEZerU3Gxovp68
OymDV+NMwx6D7m5yFy8tEJkUvUkox3s55wuGvk50ahQvSPdEEBAdWLLVx7//CmcuWnxLO+9JSyRr
ldtmmd4XKZZp28ZmXMy16uohJEfC16TlpJoWCwYQkc+IEP3x5ZH70WVEQZvFDEFSVZLjQ9II17Km
QFmO+vca0gW/xadJc1PA/qGVxMoY5pFk3InsB1jSTAhlMOml5RHlVuqiZ8a2hVUs+0BfSX4k0QGw
QWw9On4znNCZvYdv1Y5pIYAyUR3UnWnEr714cVIcqWU7wlnuUcfuUQAIB9RJ7+QwffiVPdiz/mc5
zFGVTXZ35XlQoe5TsmnXNmXpvkkuzBM6qbx2jGGhIcxbBp5+76mekyYqB+RS7PJRSTBQ+mnYgcy6
6MV8JE4KWDkPC24ccYYIrNpzw7CusCd+scMZurovTVF65Gz0hYysBrludLLpQFUE7b/FmFMZZlaP
UAZYwUEt/wh4fKPcqTis1GENpDOnmTolfgTEjAk+FEJVU/CmLL2SarTzjf0a+m6MTQEI20uhktqx
vQQzS8hElmccDbmpT6bBYH1E3XbWxK4WlDkoGaMbTOGSbFWXBUHVtfiRwCbZhf96Gg9mrsF0S3EC
2259qc0Iyagsgn7cDe3L1Kr7W3QSOgPU2+731qnxlhUEM67e5fu390OZhZct6DDLyARKlPkwzkLg
1V3Ec2vgdt+fzJBpHJyFUrQNUh8k7l4KLgYjMCmJjblyZogZ8KXmtIEE4TzcotZDO9KEi8eYEwbl
MQvvT662vlFXVKDnzPhGxwa95Ih5sTBrmMDsmnqjh9eyIX6vI1nXTX485/jyk4jQ6yNcmUg2iLJQ
oBoxCaEyHkW2xwDsNEk+Z9moMZvaf59Iag4tnd/NGPE4vMSv6kBz+05y7hJvZzbe4wvG1j5CB6mp
qC2lvslsyhDfHiCjFxACg9dgG2CaPCw63cg0acjs3+WAUyNCGqiElqnRwSZchnNecXKNViFOx/OP
EXNy1Q7KO+azf4V42U4cfLytTOYepne42LznEPfSAiIE3Bhbv5yMSB5DjC6KouDrMPabqRuRRHHQ
ddvSgyiq/FNBHGNbh6psiXhfcJ28EYkPXG61cURg7ELZTirMXekAdcs2OVQbc4jz5FKYNkfUfg4E
gryF0+cq3C2DXnBk9v1GpsmKu3lzv0nriVu/qj0BnW/n1DcGfzkIcDMUvR4K2KbPGdzAVjJ1RQwc
o1o2FEDrnqMWmp2NGJsvmSvsm9dKGmE9DNwWrcw3CGuocfQxD/91SRI7WUrKI0zZjTs4UczNqYqa
JZQx5ocn8QXsaFTjbQo6nWKlfTqy24gEUeEddA8yhnl80uXmCpVFB26NCCzpfCnAnVE7WTwmp2U0
dXJDs7eAgwOLQdKxYwSw98pcYiPf8txZMIyBYUelduXNZ+KkpgTogStSW8p/tYq64FpBrojYwQIx
Am+fFcnd1ejJYwiW48jyyJPEsg6o6gp9clX+GTfTSKmbmhOI57Po1M9kUmvOJi7r6C6ZUWJYfddG
opy2gMcYuNuFuLwYESRn1wr51Pzpr8x5GVnTp4VPnORbFcsLSGHyDWr+MduihR2a6uxRyNbiu6l2
eaKyQQIZVDLf5IBhtTRcwWIpYu7ki4G2TN43vvIBkEjISwPDP6WPuvaxcgZOvy84BsgSd5C3ei6U
938T0xpTgqYdt+5QsV3Z4xSosfmQMg4GkTolV3e7x4maWn290swrYNQI3NPoACTbeRV29yTv9KQ5
YhNld7YZG88GkP9xsnug1xmmQAF4GA5S9t400wzE9c02Ch+6WOSDe/itXBF38388UjvKM07LikX7
yHeXFE8MGCYoa7EuPifXqCtTdGn99AB/oZIz5jqNCm7/YrMPAjPCteOXraIc4G3//jMiHpAvkse6
mi0IAVhRqc3u2WqvSXh6VeVei1qpSApy1wFfB5qQnq8MqLyvXunmQGdf6obtSW3LxkTqO7YfoC/L
0kxqkoRXLbRW1xQKafAWdWwyv7aEARXEt+H7PYy+Vpid+L9yXxdFfQISCVq39JfyjAI2dyehKZL3
HdXV5EhpK4ote9Hajov7vtBzwEc1WtYUUoN6buw3Qs71evtQRrCpeDuHrAYUx+nAo87quk4alBDX
OfBAHfCCaOwC2oJV2bR8B7/pZzO3cqW0Fdg+/54wufOLSbqdDKINcSu3otVvv1w5FFIToYDcGyE2
EJAb2AAmzNQgBQkpPRvEaW+GuBuYOp9Ci8T8E2anqlRIY5y4CYcyoDYZ8Ixg+HjV36raqsAXrSD/
8GVX04DN/vPqXPu4RUVN7XaMC/WXNa14zzxySsykvDdU3ELWCdnTQEBYf3Y1GMFkhfbTLIjNJ4EE
clfgZs9AOlosfJXhkbDgPLXroVsPzwfKLV2kDEt4FUdduDx5LnrHBMfYzN3pwEPcSSauClXhVeCx
Hw3SvaHrbRl9YlX4fbJIx7CiiV7+goAHO9UrjTnjnXHqEOS9XVb8CuULB9s5w606VpUVYs2wsls/
PFTHhPlc3W7Yq8ZVJSNPdfjA7QPnZheVj2EuiJTuOYDomIAfaWMOXQko1TZ11pqwW2I9I5afKgQH
8QQiFFdj58KD1v6IHRDJhm94XXxdGsz62hknKg9i5SgQXuM9Eb4jZ7WVbparAJbRR0aRgcvgOiDi
yKPqn50lo5Nad+E01m7b0pfXOfAQWX3unCD1iAxtStGsFezUU+o6G35K6GEyucJJvNEKUw+HkAIK
phFAXUmMcOnJWJPXy1AZJDxdvsvVm+ds3tMhDj3bl1jmH3gugo7Faa3VIceTpqU56gYn5Hc+u4S+
b6XBFgT/F4Ks/1vMGyDUipWVCxbItAOUVvRmQM89gFDv6iGBHNgHx0Qi8HfhusasHzXFrZj4QUo2
yAWj5hEAyEYjUzpYjWP9ZO1bhOZHehFrLiIGUw6X50Hq3PXz8bMHmiiLwn8hpv7d6mfAYD+DAQNw
0ehFex29R5stCaEbeHrg6y8gtnvy7VNR/69+NyzzDk9v4XhbnSBL3j3bAAYwuWSXg0YrqHPnfaJr
BIIZ6f8LEeWFS3q6s+RKYQ3HtQ+hyfZUfJPU+/lK1KEuiEtJBsFRJj0PVmDpCBnMA9/RrfWYprQk
yBMOGZjzxjfUoOjdh/SgtcrpRLfhs7VXgo5Hkdro9ZIP2GweXi+xtQ01u8bL/U/YQw7CzzVQowDT
5zCHxENiMB79+DqLEq5oQAHAILGof0bJIZmY0XByw/+RNo37GbNNfZlyMXXfHKLYQ0UYMbuMdQ1r
+sTdsuHqYpTC1yUCzz4qSjUb8Nn3I9YtkUIYti73lyCKd1VQgPufYCuKAwMc3e5kSWxfTMJyLVqz
WxR8wwx8JAti6ONzhoSmsl1owz9qlDZ8cPH2PqM5izlWy4Leltqpjk5WUkU2U7KzZorJq4hyKGFk
6UYW0kJLhh3dmqAntZoyh4W6nJ3ZSLQy95HpMQiRjQZHzdQbFS+lL2gscPLVlMzMISbaMFFSylS3
dOg9ADgT2xzedpFvF8FcFtcCzZ9fUFHsJJ2cjpeiCexiwc8kwIo7ibe+7iQorhk4d+cevBViWDPQ
9uNc4E57UOgZHUEOD5XQ81y+a7LYVn2j0a8rGqaYjQYf5h8riXKato32NjGsELBLn30Ya9V2eB6J
hVZhfSy0hyZQxvO00/fG9Ixms0Sq7NAwcpujWvgVbhILyoL51KqVjyV0Dl2KV/ZWe2EfJ+Lw+fuw
HNQVR3hkt2WTcKf2jmjrgLpULwNEI9VB3r+zhJM+e31S51unlKN2WD1j+mVL+JsNFdz7/lkT9Gh7
wKgeQiPG6D9AbPAgvDScwE/hDa6g5mJ76URfTHcn0TKgWL1kI6UpM/8tlT9UrU/OlHp468Oxl6Rd
wxpOxdDaZ8nu1W2xC6fGJFZqs0GnBCS7raxsjrCp18mUq6bnP7KgNcNNxcfpkcKr9RPmBjOB6Vz5
lJFWGyYAp9SnjI/MP2WALNqDqlzZ8N1rya9zLtDX2nNSMysKtDJkldWOm0rd6U9siXOJSsGCtp6/
MwimpZ3YTAuFNOSl7J71+scH3SWxH4RJ9VwPTf4wkG94SXNmEktHkE06ZwbTJh2ICbv6lUGyQzXG
vOVAFpq9/L8nXoMvIc7lo0ikz7dOdx7DIV0n0dczEd2waBERCGAB9ljOk7ZsmG0otfYiFLo+k4J1
21r1PRatiioKImVmrsQ3PPRF7uRoBVzuZ0LvzTibDUyYZGmh0xaIF6/z4qQFqZ3cd3w85gOl7UQ7
6A9amc+DXU4xQ6lCsXXH53Zl4+SX14kQ/C7nvZNEXdBdsrRC2X0FxHYqNOtELdEoTaEMkhNXF3lO
uiUAlp3ts8spCavevFJ4IVJqpiL9rHM+2GODXhPE8psCS+LXFHitZswF7R3cELWKk4B9pw9VV48F
VjCMBjJZwcaJRGPombbBKOrZpVBzp11xxnjKiLvKLFVTGzVH7pCT+0TO+vBMesZnjqEDqogxGpjE
U4l1jQSaIfnRpH5gi5lj1YWtC0aVi2CesIr8fNdsAfGWq2sHdrOKNhtqmzf9GuytL5WtfXK/b5JO
Z6L2Pb0vxj6ZXjDJ3CPN/TvJcYQyi2XIisHoj+lxbMt4qR6fCgDmPQcr5xH3xJImC9xAFSiWH2tL
kzfwCWCrTcXx4IqVTpzm7epomEQs8febCfFiFWy8SV8EfHvAk7p0bDeRY+7unlU2PcAUryypnr0+
9La+b/lJ+pSd/HkiWUJosyWS8Gc/ODSREDNQ07k2PnIOxpXE9YLL+gn71VNlxQfuDqgtIIms9IL0
TJ41LRrxr6uDtEU4xlbdtg3vNZu8wdcUEi4jBHzA8N9zaHGjbPjmZnCPUuiViO5GpaontppesCoD
Mng+qVHf6TnvpiD6WX8SuhTMEWqQay4sxsTMqRR/wFFR+MxtevLMmKJvwFyHX64uSMan5IAfQ5Br
3sS6O1clUL+d92w6XbEnkxocqKRiSsDj0abhNmXs5EHd5CVYujVg5eIK+E7u08TOEnGYx9CHH+Oa
ploAFrfZFVgA7WHalmv5wpk4atxBfwez81bIPRIFkLjP8ku0mgezv/plpMRiDg1DB2zfMCVIPKtV
FjI2rX11oubYfp/pu04TEhXg7uHa0oDgbGyZRo0NUhfGI3UFVMaP0yyGDg2DKzNuZGK0Lx4QqpLI
LWWsNAOb59YsXW8bXS36lRofBShzvuBU1RT5lA0aRgqv00bsUtCT4w6Zl2gh/tELLCMJdJpu4tbP
y2aJCtahvAqnUB9ag4ZXI4NcenVf5xv7hSKoYOzMtJMpVV+U93h1F4oX/Py9X0u4yx4aHPkjNZBi
GmC22jv63e3I1oLRlJIG2vBxTS0QUZy4LDKMCmfX5t9wLz/x7YT5HrDh0sG3BkDiNL5vdUrZ+xs2
P8AvQ6+BHKggjFOYRinxR5gNKK2dGUlsNBEIQNJmWIVFZnQeTT+Talx8SLGD+caIBIogsI8vSy7R
Q/IwHms6P2WJUtGg1SL4WkFveNDYkMfJWdpsOHoSKlwMOryfdXCfKHERpJbbKGc4IvS4asUdX/8L
vAD0I53z/H+p2lbcKzO3YVAuZP+XAVr0dQ8yEEPVz6XcmT+LyROkVVmvmaajBh84ygFWM3hcl/qU
dk69DkY3XKaQQb1K4PDdAVJBCZX1Dx84Yy7uMiOfM1OWbnsQrhJ6UP2vbzyCulyM5tt5PGHea23J
UgY1VVBZgR1jLrQ5mw6oLj8vmTWcJnlemrbRj3Yn35W56qeWIzya+piuIKF5nZMN8AZJdKZvSFOl
o3qUojNDMTZnwYjKCa3M5V8LDlowpPcWMYobBE8pkdPix7aF8DdGKAYajY9AbdKGXo0AzpAVvnPc
s+6qZEI5N3M/vbbkV0CBbXpp7MiREMNMvD2xCP1rQWZjddiCQB9Hisz8z1rNk8EmXPOHZmo1rpis
b/8tk53BLfBVjApUK940ZQYo50GYxJMx/eMGlpstHlC9T1HRs+cTYbCH5HJ7GVubXNXy167gAryM
t1vrWXor7+QGyFpouwQbSjDV5aFmSmHQZUJAMEvFaDmFKFKnARYeBF91k9Fyu2o28uFF8Md/38i5
oirhCuS4uQU4yNECVKDqc992+WzdzVajVdT4xWb14HGGKQBgs3TJzxkREZnJB+1DTdPBSeylKgu7
5HL8EKmUh3FdLJkRKsDP/IQMGGrNGp/Wl+vNs0Pf3t8iN0VOHQN8oyLzP60k23mAF9a6sOojsGzm
UAfgrpXBR6qHiiD3uGCp3TYMz52K1TBLfxPR1CB9eoHJvWY6a+TLNYz8K+GFNByfwxqHZUHH7jdW
bKm+tUQj9n5HGnxxEcfhMqkBLgYg+HhQPIkc/MEi37JDENSsLDVfkjL3WcOhZRHV6YNuKSDjOvk3
l5x5cXetKUm8rJSR3thM0R4diI9CJsdDoQsiQ9EWPx0/trpO8dYcHT99XG7bcRsk350FTNZd6L8u
sQDOmRxVnAj1isztZsWH8rgUCQ+sD0jZDolQ1rZaVisacf0bdcKL4TMdRvyrMzB+TFmehz6BYiYc
OMWQruoLMXOss+LDRViPmT6IquiPiTQPapXbf6rYlEnPAiHYzIaO7GtofvhLmXxAC4d2XIxxbw1f
mCICRg6wddvhk9zVLw3SfEfOlmC5CK3uV/sJ6+aNh0AFzQbXs7tmkEiMNz4ezSAmzE9EZraoNZaA
s8hWNfX3YPmVZC6L80hAn5ZqSUhEh6Lh0dkGl5p2gvNIqBmEsCVagDnXVIgEaLquiY7gjKMEbflp
4emgiLsnSE6cK4ZvGh/IcdWT4jMDZhgIf9jb22UJxhDdNeIYMW+dgXQ7FbVYaCxxxR49ZvhaB4a5
m2XLjfL/sVq8qT0vQ1h6vlmXH2DEK3bNpPRuyePGH9a+hgFa1KKp8C0PAcgOPJxatU7JaZ37FVoB
DsqvI0LmteKNgx3Btj6viYDAveLT39bO3phrA8b62ZwHHEoRRn93EffXL9D9MeGL3AUDs/dju5YZ
0U1li3BkfBW5KPhIp1BEp0krpyo5ctbWIoMVwM9TvanFC9T9pCLT58s5BCcIsYkPQRV2JwQRgbaw
ylvOO6/MGIcQ6+i3dKhGEdCLHCwI2Dqy7RUxJ47rX+VDl/NMSkhTOsYGNUmp6NNOA1u1Kpg5RIRM
FSASMwjmhsigmsozu5rnsXEcIuS/vOA+wJtJuQm1X897jLfeFErfpM0ZL4XZNE++RAjDUeG+XaOz
wsb4mgKLdqOjhFh9mlE/758FWwxiWW1Ppx1DMGvFrktuq2pTbpKOnjRciQxHK99jqotZz+arFilz
iDdYalAYBCK+QBUFL/cZC6TwGdSwoKvFQLyjGSakmPv2JRB1hwcBQ+IZQVyCzW4JWE4vsNZMrC2o
UDYIm3xumAYIahst92bAyi8DPZDx5FjVjA2zieN1//Gd68W6+MDgvZ/mF1Nn+qG9wUg5duGAmpGC
QCO53z5D5XZnhlU5IQHt1FWT3I4KYx/LUbOW+AdqJGRDMD6tKMWnfY7nVfsKkM2ARm28lNVaaMLn
hpynf8I977lrXzcDRdZfR9C71FKkch+f3xxqnJ9QRmuoNpjl+R4tZgLZlyfY1WDuf3gpuvZeZQuH
0Vq2MyuavpnerZasZTg/upt5EOhwgoGh2xoVip8uvOEbZb8h+0iPjZKQC9CkaBvOM2PseCx1IQRk
2t2uQz0Vh4keCdP30+RHKKUMMNv05mf59MWNU1vWipM4CLm2KPkVR2Pa19DOzT+dAV3m/F52xBY4
wZoHlsQuptuPKfjExNw1jhTc2JyJ39g2GgWTWm/JurKSyka/arE/9nxie3jpx6JQJTYzsuhVHGzD
Ge5ZodBLraTVgS1aBGMl2LmS1zUasEZE9NEutPoOc3VVHVBgMpU/e6x29d7qilRki4BeCN64Srb+
bAQO6IsQ4w47z+UHh80GIZLHg2oGGcGU6jtAkxrMtOY/dYUM3HhoGqOsW8ti6lYyLz+Lbxz8w+SB
vLVhpbkfkwY7UYakIoZdca8JvxRIYOw76Axeov5g+KI5BqxXe0WXnAfccKacdI1Mg+XGiE8BpvnY
fbQFranu3jzImAuLSgp46gvLe0p7ZtJwxuEFmJzcPIO/w0F1lqaszMIkzMPyU3X9rAUzAdIXm+Zc
4ZL3HbS/zYezka2qjiWEXn+tf9sjlcVicfXDz/YzodtKQRaNqDXX7YCC5yKt7F5e6eACMtftobG2
sf4Cb4QGcVK0YdaE2dV30/75HI4iQcRx1dHavESVBPFPZbb/10yuuUlsNoQHCTYC3xlwR2miK/5f
DFivQmSllEed0sJy8LXf64FJu1Ra0OkkGRkjwFzh4px1O/3USAvPePM+aQVCbo+k5mNUgynRpGr0
5n71k52o++U52T4vb50C0id+FpMCq5NoLQ5/5v1HGLwcRR05/ev+ZP6oWSIJpFamLsgKlRrO8czj
fqfiVuq2EHYuFbwkfb0ci8gOh35XbXtUhcPoI8rNauELrjTTyFewu9JmLqB9hkxk5Pby+w0pJtq4
3ava7WTfFu3yf3kYk8XGhpS1xnZPjrUy0Vlga2Yb9X0/m9T4mBDwDeyymXukIBTA+m+95aUO11WZ
zO2qX0ps6uxdIkukWiJj6OaYN3LLc120dYJG3lSAuEbROWq6dcuN9gQYnbQiM3AV8n2P/lgoDFx8
7/y1Y48SmGDYJbQM9zdY/BzMj/awJJaITqJUQy+dMqWL3UYfU3u55tBaacfbgcV5xqNWE/SZpIqf
em2C6HIIPqyepOzGnRNHfcTR99kiRbsWYoyx/LITVtWDsJ8poziwwlOdKn52BkPuCNZszHcGCuBl
bBsWc8wo6HE8wIaxKGue1OFsZwxuxcvuz+zAJX4ZJNBoWcOc6Bbzbxrthr+QsvAGkOuSwJS1GZCL
P90iOuozKWq1azgCnUY/XEUSe6alocLQzr4H/bAI0iZv0FwPLT2ZzODftumKSc1s7y6EY2JtZE7T
HlaxhI6YOqRj7zjphErl82ypDedSrobdkBlHT1fz9yq64g3LUrPQroyYJGx5Ts2x7YXnOzFn0wKk
SFvW01rr70Urcy39pFuP9mu33xafLnhPUc4ogQsrIVnSfUJPn+29+WGA7c92HniOuoe0KyKxpsXA
YZu2zn3lvUiLizWURkUZmnNsAmXYBeXgCu+tV+TTMbd4TMjhkcgWUB/AFda5sbiBSJKt3Z8LXLjl
TONjXb6vplLqeZ7BQrRnql3RaefDVD2YWvDDkgmy88pu9Y1mPHdPV+wIIg+L/OSNfa+C/bD0T6XV
f4SQV0HlVvirJWWmt8WdAXjI0a9DB6j7VAgDx5VrsFe2c+A5MqEaJ1x0/Nzuj5nDPtS7bz9vuk44
hyApG0Y+VuVffnCUsz8fayYfGjkfsxkuiengvq6QEd++ZRhNHhITIVAKc6qTPU1nRk1fNMsza9CZ
wf+SXlGaDCYVkCXF2PtZeWXCJlsQVkl1mRnWhZWrHOITpxjDi581K8/z3hk58GEXft3ElDqZJouM
QPHs+fvLmr37W/tTFzaMw0G1KifjjVyB+9yAMYFgAQhLY7RQ2B1XVROCnvFgIC+GE88pxT8z0mgd
m1HT77EWhfA3cXqSc1Ll0ZxYMVsNuLv+RTXfj4q0e2dTzqDsRZ8C2uva5iNVUBOKPWTe+uzcD3K7
FikGzR0L/ZS824ntsHKAB9u1dEGKbJtbyLgE1+UZJfeOA7ODlP2t28bVoq8bsFao5IDq5mVFfYif
gEan+2OMbIDL9XzLJV1lVUHdL7V1IbCxeZ45075nvcOs97qlpHzUX2h3PcnxXQE4SEK1b9TG8A8M
tp67yejhughrnUgPpWwYrFRLKHzHHpmp1AKrGw89qjRqdVOxTqS1n9pBraeMnLTzGMETMEZn67rV
DCG5T8VaPYYHG5aHPi7GsSFr6tUP8J3XaZLukgjqn4yOgdBdy3ZAzJXBQ2Sb0vKZpvY0M9/mTXlP
HNn9m/ZAQXtcNIvGJlPBSsXreASHXX9S2ln0QebQmfKkFrbC7P99ihzweKaHQHabcG7FcRdAk3Uv
mUEJtSXORO9GzEFQFeXftQZ3NbCMRbiDPjYM1aGcP7cL0ghKg8a/BG6IpHolZprOJ5JTKmH5wBFo
sIs2+ZhH/RiW+rEU8vbSOQELOyFAz/cMrVFIdqBHCTeqr40M66menkye1R4jX7vDMfGBWZb1P+Zh
AwCrx78YtN1WUoadP5yeQ7LBDMWhVey1KJBfODzQTExjhZFwU0Qq88vLxESsauwQWIfd9vAw5bxq
neRAqNZomxlvrbt8SKw2SIdOJQIM35u21T3/igbRWP7ClJje17d7/V1A3uNOoLf6ByZh2AEzH9O6
+w2iA2jC4cTquyG5awV3kFOzNsZ6Bmzsw49HWiKLLqoGEEqza6wSml8KxcvmyhSloocg216vTDr6
OEADo31pM8doLbjvXOaPZkdyYqHLbh04a7lpjLBfV9SLxpLhvqZkaRCkIJCVIDlt+2J7b4qnpJ8X
O1kCLpTRAXVWB60j9lLQiwJZVeJ+tGwplmV5ptiFBuOKmYxnFWede0Mfzchc+YBJhHdPYqAUyjol
VajEEj/VCZA96SsQ+q3EOfvM/ErGXwtW+nIVNw0TYTsWUJ3N8kzHreMEmWuQwuEsk16e3L5MPVQ+
IJ1N/WclU/ZmlLecAjDDg855z4+l2HHV/W3TMJHAgiOmhgBgON6J9K8G0Ygr9FyKyhRCnUUWH9/F
CL6zSkn9MxNsNZQH78N3eu59ZBGnZkzoYal/6k3CRvT//PEE4fE/Kd1V+XATXpbxc652EIDzXy8h
N8wsJJ6RCudGJO6SYc1jQ38Y0/AnbINgFIFCfJLnatZ9T/rlPK2QYndzderS7xwJNyMvzsfm8Xzv
009PYx0tOnrgu3EaaHecRgpxhABUdCGENP0UKK5orCK2cbs1esROnvfno4QnJLGcqRiIVMEHEIKA
OgSna4KfGHRg+GWpyZPsc8GyoNAAhC8lAZ4Kbec7TqMyjBGeo4MShqeI0siHJQ76XKveCLcGb82D
sziRw/SHjIcZ5bjrNpcP6+ICHvOMYqWPnQ2WIA6KELXpFbcQHo3QcBToUxMz0peasMLf3L8gEmxz
VatNR9+V7yZQ68eTrLgEmzp/N/II/nEpdPBUk37l1HyRVqm3IaxuSkdTyK43c/oQWbWz06rc5yaL
QNXLZNvKP4jSpbGitersK2F5zNvupc6FiGFfwqqqlYe0LwZeH0rjiXAh4kx9A1GJvkTL6bkQl2aj
mYZR/oh1FNAERKYHpxMxY8jLwUtxiaaulnOUV3zDZAoptxyZEo5unK4idTRhnl8HGKOxHzJh1tXc
71GEUyb8OdtghAUYBZkHjQb0tBkJ9uRXq2eDfHtRXLJhWE9XoXK3u/20oxtfhPIyHgPE8VPGtIeQ
/yjVsBFR8BJ657jGNjallzMcsYJk9XS8ztemHe+B+WeCPwVXHuSNi0W3v+Pm5zGVyel1roD6iWIm
2kssdFkd2e9j2iUWEbyz7wTCQBZlR/g2fP7+WP/9eFjP2HvjToSfjyyg1I8uAlmawgHtu0R77hhA
Oo1DD09s7P76my9LXay5dK+L7dtinhWbYcsKpuQAWrZ7jq//zq7nf7ChrsG5DsiKIrm2xXr5Uh9s
QcvzmK4z5u4rPlHtjfpAjnZOymJq2ytzXK3Sr0x+8+urvZzHcbHGQ7g92p6tJaCmBoZS5UPPX0+v
4BjiAwsC9PJ/riHhj4kZQP9V/k2ih6BMVI00Yic2bkkBCwKLKH9/2l8ts9rPHW8L2r+yGb+2vO06
FGt+Yx0WPficqTaIckFAX6PtLhWyfJ5VpbXMZo1jc705vnRz4jN63Xoetvg7NEtE5f5Tun/GGFqn
888FAm3AhMKFyJ8Xa2GtkRN2xrgkWQfEK+bQA9A+Y5GzKyWwU/faC1gDjEWbG+IZYFRL14lHBANW
ISOjHymjcdcrt5kDJZaAssFHR6Ys1qTdxIEJLWHarM2szYDFiJDVIl8l7a1RIbhktqE2wVl4X57w
4FkjkRzBwnuDSsn3TC/PAFEzAydQvPobKRra016DRa+jr0iF/0H4f9cBKA8BmYJG0l900cHKaExe
lfAdd4NNZZEQivg3hfuIOswVftzzyEW+MLw6B0I6r4AtZqPJFOIS5S60V1/dPOr6ucYNvGS/T6mn
7CvaeGmIlf+r/PRVXqhOw7Y1FO46B8AnErRKlXGfHflb1eco6qnSX5fIpvMSJkQb+Uo9SX5G/V7n
Kg1XnDKCCbUX2BfL0Z/av32OyIxnUOly5uLHOy1oXClWQ2O7nZbEGairuHF5siOL1i8HP4tqO9VM
pJJnxyO3sfNNAwWXyTgaZmWer+flUmIqI6Ft7MSv3EAfgDtyXOVTxnsYj8aEC7dadBL5kf1aq6Gq
ul7CUbCuvoUf+Dy6NyxRzXsQK5mYDgH5Y1Z+DJqmCZN6CE4Iyx9eA8pbKLKW9Jh6lA7fhwlfAEHp
77J8M31zJf/kkd6bIt//Gqle+htPDhZLAHGHD3BGCe8Kk8tFzUpZHI30sJUuVHJmeVcneylVEaq4
DiAvG9QY8mo/RgRfew3JpfJ0rHEWoArf6XcBlYqApoKFlO7RlviZyY6GEt6M2N0xwXXiGcI4/vI/
0Tnutdm8pa/dDJUM5Y55ih0PpPWHzWgjr8cpbRITmg8fZfzYwAtv6dD13c+XohQqCrDQcWJ1hKAd
CFj2/gVuBYdCAqURCJGlOyIsb7nI8j+nxWVEHuZ4NKPYL3dsyZ1Q4jse6wm382yos/mRDXsrSNwF
kTq3Ch2fi3GNI6q4fwAnGQ6LMi51SENIxDGBpEbulk5EY3kgenq821BHuHLrvcaOJSCKRtNZS8Qn
p36JD/lx5hOw6TAEdeaCIPX4IaMooPsaZg3eXxZZudAQv7UNWRKf+dD9gXXszgshyHs48MBIjepB
m2acLmua8XYsWfEJTrxk2Plo2ToTzX56VTfKFKt3DM2nS0dpClCnoScNX/F1vZSGaDzJKTJa5Aj0
hAuAgPF8wb+DsO5R34XNjpJA5B1LE1fgL3V2jvrvhE0rOYM9gG0UiRJiymOGNzVfcMFOyD1eM8nU
e66UqMxkM2q99EPrmp5hs7vuggANxZOyw+kTn8rpIj7FOpyNbkKgtuM2m6Fnk1jqGeVlg1BFiimE
pL03+QOUc2aH4TKkBp13RpphPN8eDxjE3yMnYQikAgzURubpNo0WdnPpJ8n+jbV9AKAKT64iz/ox
7tJw1WpY6sOVqQoWRZRtAPbLr5rWAoNmGAmIr0aESvXL7RpCVk3Qb0ixnR285MCAb2V7N3EnhnDc
6qbGLqnz+wpkJYQ+LJVRQtVGi+/n+Im0ylGZCHp1ntoD521PGXE+U14xg47vMXobx9/8C98lhv7V
k1z56QJcpR1bl1hJZ0S285EXQcDkj1za6VZ1ykOTY7wPLfi//GOEqUA8G9Ckk+vkjGBZbpe/hTVS
Np34fQgw8/UfHqzYsEZrx+VnIi5kSWzAdGS55zMw0FtwyKS1KAi0LKNUjlrq2iEds9tIM/pp+7Lg
u7oOpY502xiukzmW+hUz+T5tNjyDzAD0NWIqcTqAKaY+VlLN2TblMhbq/glImDWYkZveXVPC7IQD
uuFtK4CP0i5X78hT4DDitiytcH/XToK/DIy2FFmtiWUL2KlBVPzZbt5Srryp+ZdBEfLLiSaG7ooF
f90Ct6k+AS9/5KuOZwhtaNjeXQijoC/RdEbWBunn6mpeNMyYJwBqNYgzGLXT3SntbX/EtlsbIkrq
ySjS5cOuz7h624elRhq5yJYkqqLhxJvzgnE0OqI7qoB4Mx9ToGcfRkBvT73M8zIFmRh8bNDrMmKL
XMpgsUdnRUgU3ogv4YpKvh3vdTC9nM/NnbF5dZNSLXbVKCyoE4p7kbMtrt6WgDBhDtBU69hgEGzV
Az/ev/ixsnylYmBvTNWghL/BTA9DJQ+9xKaOkgMRFT14vJh0IHPdwdZ2nrdZKWePMPt4W6pQnuj/
UhxYtjph6pF7F224lYESnu2EzeMnUF8sQl1a1aJUqHBfivxVNkupIfsQoU4jdUaDbUUCl9gENFA4
zGFhZlQSdSqG3b8u96R+HI+3MajZgZv/ZSUkTDvG+uoJZqkMYFVy5k2d+k+yAW4WtrsFHjwNlEMp
NLv2c0YwCmPgsxPvqjETGvtFUe2j57ka/PVSEMMm2kVKuFoUMJLMe0xfBiFDSSmuMjd+DT8qv+kL
7HknHwsuAoUQFpHtJbQ2OAVjpOWgaVBvUFadHORaBTjI75dom/8RWirojCTVyEbFDb+I+YC52p04
gB/ES5TSyAkzdB/y/nH0ZFrKJrVn5SMc1NTqzbViIne7gqAuIFPyiszwfxNhDhiQfC829Ood4YJS
lvmbqE+SBTqZlsS3N/YQ88OM+TAm9yi0xpaa1McxMvqN4ve5r6OupXMMG1WE2aJDlgpLLUtrRHAm
a6Pulf0HSxeVbmJeGt9tAHiitLww3i02LLnLsRY4kBeHIEutCDXsr/ynbLgxGG58EnyK2rndIdoc
m9EJfxa2fn6An44zog41z9BpLXGQ/t6OQyrN7uZSw5mF8M79kKKb2uYxcVgTs6N4zZbuzaW5XIDR
/COJHA0Uva/61rEwHaS9iyJZ1BvOdS1mUiQ2Myo2/6LTqq3pQLHLrzGuiyUdMDhNVOZCrtARnPz7
svyYwDFUfbM6cAz7pmEgmsOhJ6RLa3j65IZg4dX/faNL8VP/gBBJ6rMXdqQzT8V/TKL9Nfn/XV1O
/xdF2K91n01kPlChwX31kkqar5JxzWu5bXeEYBQLnTlqIZEFECqDy1dIBIpGWJ+jVWt/1hne597p
xdIqszsA49xDM5aMmmlMUeFMjKW4XQWCV1j6toSrvqjA+1d+LBycCw6VQX2tD++GwqiSqeCE3ota
DhhlD9I1MrI4gNS6GgNe6f6a5snIRPshIuyM5YrFsUJINOXQbnTGrAl6IFMHTaeE9pJWbkzAQuG2
2/3DdMnlMlSleWaN6frroQbSP+5JrNoLtbSXZiAEBLG1hFJzv+C4clnsP0wuU+4bF41WDYP37PRc
2ZIUwCYNT7ZMyYfrCQBkJUD3j3RGlrk0QDcuxLnXyjhq7Z2CuSFGovt6ccqh9f5erqhGs2SWmIgC
/WMQ5dctOnZ0Bv8NxPNVIPHEExtKfmCbB9ayg2Sb/HQgD39LLHYqiGCh/TJNJ5oiBWws5QqxnYIq
vKrK/PSqL3bLJ9YZO+/HiwBtDBOiVRIstFS6/2X6HlJsLCCJFOUB1R7TvG/oS+Mkh1ei8A0dgPRb
BOPqi4dnzbzIdjhC9fzNrhCyulPNZcRAOmPl9FKxt3vseTxCFq+rRmbfPBBixRRXnM2w/OM37iHJ
nHEJcr0+FYYL0lKXKcPNr7oHMYhaQ18j1lB+CNLOek6FzMY0b5ZxLo+wF7StTyKHGG4h9jjZrpBa
CR9fSd30YAVny8IM5pCwQJMIJCP0MXsoXToHVpxyThKPy4I4Rs4HB7n4J8f1LeUbIB5gPnzgm7Hv
2YsSdwASjLuR/aZDCKMvCeirFO4FeXEA8wfbtdpvB2Xj2mDmWqYImUALlU+yUzsxYolmDmhkydrD
GMqMsMUKX2Fq/QsV1sJx57Lhb7eTp7dncgmfUh4xHuWL0wtgfNvtybJhEVA23dSjxTIaNPIuKN/r
7fGFA+/8K+qpx5KWg+stQzrpERrdKk20Xgwy+0Nc1SKgUz2lU0Bnk6chTydOzrslSdfqqwlRj1yy
Pq5edX+8yIPBO/0hPaMJBFUvhXyjWASza5HrTL+armWtBfkJapL0AbHyECVX5S4hvivhh2/1hr9J
xK3lNr/al2+5l9qE08wyG5n3wil9A7p1CQmSZwC5iTChXI/Q0+EPE7obi2aHFjDsbX5Judn2344D
m6uUFWQfqi+qWL9+dcnUUivDACJ60arv5p+dw/RiRIDjpuYpXob6sQzm1OreVWQ9KYknQKsEfpb4
suwM7rCQjd5C5YfFMWwVMHavnl7/WjmVYV3B1c78s9znfckKt5GKSAhY4BfipKYaJAidMx0qgpJn
OV/OtLOF/bRcY5J7HgzlXX3z6wAlp2KBeTN4wyP0qIIflyv+lugun4NdeblY2tAcs+6Dj0bXH2y7
Qltt343G9Od712dOQQUa9EWkS3ebortAdMuBXo1i6cmDy1cHbkcAwyeugYoJc+1SI2lkFvQ0PyPk
2DXGsNorVW0uLmceqH7xzhBASb2AsZRNrS0wa+I7ZW2bN0On5glsL/aVwTwEn8MWHQvRPlzryV6O
m4y0Y1FLPNvyI+GbGKJ/kbNICl2URKyagobUtB2GqtELmte230Iav0Ay+0GSfYgC84GT7keXr4/1
rlyvPprooBTrz0yyj+1Bn88n2+U2tmj67ivsEdY4bRUxwHk0KwNOKDzftI/hHIu2hA8NrI3UbhY0
vnpe1jCkZwz2m833EBcppY8QjHepMhITlDdW4pRG9M3KkVNm4zaWu0xHqSl6ngdx0ZJk3YFAvvAo
CZ9BhK6TU+Ktmg3s2W9abTGLt74YMlwu/rsd1z2jMGWN4I9Ln0kQWjolMjFFum1OsF6X1/I1HiEF
1Q5M4qjFeteR2s2ktQR5j8mJ6lC1sgADNE2IXXIG3GueQUuKdAup9QyJJZ/AHk1NH7W8xnHNhTaj
FQeawshQrDD1igmbLGCZ3VyEWiivcuoH5Ds2Az6t392YRLolwm1disGl+XNYREHOACCguyy4qKsw
+kyYhOMxogYWIFMtETbz08vs0abvwHXWBCVfi8Z1RN5Y0dH7RodlOMv/ZrrotGsqvM7n+VUkdO6Q
XKF/u/SaEd12EdktJrdxu4egQmahjsxjOET0/9pBYh8kunAC9u4CcYcwOIhlEAh3QWq8aJ5/uEuF
FZ1jnpUUqbKf1owpVJM9kpmIDZNvqiRUqJEOYw27fzR4uehTcEdLJ8V5C0MsWOzT1JRIvrbfgSc2
b6carI0H1qMFRbEfmsFpOWqrLA2I6iGdBXv4JsRnW3Z4S37mcTG+vlM9BFkObBSpFto76mceopmv
iRnfllufgo62bSY1bLcNxOZ/+1CxV0/1Fwj4QXiPLwiQMT34URMqLtvkBE/9oxaauHCNKYKcO8Fa
69Ly8qX04n6kB3IKTLokdI3XRPpf6LeO9gApN7fhM2zjBXgYffThXRRi5ncnXJ6faBafVkivqN0l
1FimFu2uGKXbpFiP/CixTHawJ9oCzw33LUyymgj0114NK0IpuBety0/7uWrheBR3o8lJFYKtYqDg
Jl7UWGDZC9S0gYo05af2zTyeoz8ZociKn/Pt2rcNxfCCMiiv98dTTjmCszNuYzT0HbpUhMxlTdbv
A2KHs7jGMrhiu+NPD96q4dB7TXWK0tC7SP28Rqz7ZwivePmxOYElocT5TRk+IneGSTMAtIkI3Zaw
6v6b/UyrZjnsfbLkPRMiPc0SXynTnF/88g4BZCc6CndI6lu8lQDZvg6qJnzIC12FSF1Or3eCtI45
eIFhEI2CIZY8tUv0v3GtWtDTsT2TjXRNjI1qYkxjKmpT44pLe9eMCOedXgKlW0WQfxIcRitpX2sQ
/BxzVFKM0AcYrjYKwauwezGgYT3csTw7Lbw2OD8So8izT+2jNUho6y3q6hevJNKKNaVDE71Gh8gJ
UHXGjTO5eqY/twV4/ACJAOH3XC2UPMfbO1Z2nAMgh2b1ZPmCBYoHh0WX4RsQRjc1cxyf+PHg1Try
ia0lfuEP9id3gUdZMHePyF9//V8ouFLjVhf1EbZflCs9kXqxQw8O27hmFAdTRHttUpPhpklXjOo/
wuvuMgH+Hql4r2wZ3D0V4ZPFSkpvrWn4P7nMkesG3smsx3WbTeeyw/sLKMmadPpm2C72616yjL7g
31ZZXatU3LY884Y0JndItTa0by+Il+te3bwWHgHqzKtMjltJRWvfqNlTDKJyxatL//PCMD73EIy/
5SraBfy34SnR3xcXHAh2bTZRLM34IOcmQAAWGI8Mkip/RwrkiVn/Uj72qSjEot8dHV981zH6c0Jq
PfZLMzthJ4w6PC2r1+UP8nTii6zM47vtLJxdtVRvXGTMctDkScK2AEu/x6x1y9RbrDUQHPK+7IHH
Rzz4yng4Y2IQakRGONguFPtFPQHos+unyS/7Emi4DB0MfeSKcpeolJo+0SmzANuFRERfKdWWvImI
mSUxsGQgsWMCqoctY4Ph2gMbnGRr2DCIFXgWFj/fQtLHztAPRnktde3KWWP+7baApA7nrpk180cf
8tf6FeiO5TMFaSpmKyeL8O+HyyvAQrf5U8T14ziHkfBDag65NjFor4rI3KVMUjPkDKtDlLSbRRYH
hngt9HPuXxaLk0CEACEO6hILRkwpOei1FnkOSBwpE3yimPRnsNBLx+em/mOUYF7jUEiyOgxhDzxl
u3bQM7v2XMbqWvZhSL/IYP8lIbwOCuAjhUDozgvHeErnbhaY+XkwU9Sxi4XO9H5rDisvTbPUDO+0
/EOWnuvQBIOhCMnVMXTl10S04MAu1i5NL1Rchtp7tpVkEj+8+/4tA1nRPHgAXkq/PXbEQHLETuNP
m+rnrW7Uq/pYJvZUhuWvnwWBP422U9KeT9O1IiitIzniExAPENiS5xHx6gdwI2B83XqEmqu5oi3E
8+yPJDesfpmXvBHahiIjxE6D4kH37gYyspMEj0kFzKOl4y/YGAaQ9uwlcTDWzA31ieEzEH8DnrAS
HtzQOrVPL3OZOUZFQQO+Duea1eksKySV/uBGYtJZbEnzNfI4LKMk0xzI7ANOOU3guUA6HoK5d0ER
FrTAr2pFZyD7FdIpHBAjqtuCbyrjYIlpBdv0vD7XrEwfQtBi+aOiJCNdw1HWM2CBKTBhq52dlUop
BzkELTu2MwNFvXZD+TuO/1a5Q9RUc94usePvLtLyhL/WbKTeG21pxVhye1ojZOF8KGcY8Caj5bBz
0T2qKEQ5rmXy+YvZTNwDD2hb8K6bVRJ7VTd2/VuzKVPLkajMxgou6Ntj4k8KmpfOV8GD1n0UbKP9
aoP+6oIMwf3LU7QcCx5qkLPWHY2GGBEQQYtOf0mS8FoSkfgsZLbeQ+P4aVW3KWA2eZDOnR5ToJsQ
uswD1VxUFCvZ5fhnx2a0zfcp1Ye3LmPCJp5ppEqz9lcJVhVGsnWBqmJPiF8S+JTXm9K4p4l5fvBw
W5gr3p+kZYGOgbBsdOx0NOZY1+ot2cOzTWLc58YLTpq3yK5L04Z+uc2pCaoBEvPsgsOzWaMJAqRG
x6IQiiWrhTidRweq92nH9AZTDaGCHUMy3wg7aR17Cf5dYNBLT9GzF+Z8QRdVNefKAHcBi4VkmOMQ
FsgWctYX4uWgV2JINMW7+CyvOftjMFR5fktyPQ70KZ5CPBx3ABmGI0qRjxCvI6lBfDqwJrrameCY
wy94tydaPSHi4ScaDcQVzkls6ycsJbttQASG4XA8OSVgzhpFamh2DYjDolVEdQx9nI/i7rgelXPc
kduuJgpw5w2Oe7x/4qW4h1eps/SCF5rkA/8MmAkuX8Xsw8ekTHYD5I4xd9XVk4SBSl5fNWi4Vtp9
DYI4f6OCA3fyevVXUVmIhQbOcZcUUk46FKWNzJ+43ZKCJSQx/QlGWnqMPVJ1TLVA37TTDAfVEYfP
hCPYCB1IpvibN0vYPxv5ufIMSJwkV7QO61biFZFUkMnXWfvvxbcnuN1d6A8/AZjhC/+HDydDcS+j
dOFQWdyuk1+y3UlUEZSKCcraYYSbAOYpe5wGDd4M0dpEJg/iw+8o9mquonLdq8HMhzIceg8OYdC9
D8vorCmqeJuhFuoukSNSDOfRaAxuUFcWv4J06tUwLVZ8eFSD+rQmwoTjDT4Xfxt9EiCHFHc2Hbek
LUZDtMA61LC41u30s9ClMcycUYyIVQDQGQY2L+2TWILKnfiHsRAmuDSFYkHENudBkI+ujoiqCbUE
E4JUEOu1ev5jZr7lma65tFEcr8ExnwbFrPQDhLFyLdiHiPEhQeah80K9yk8q20Gk1Yy0SH2lNegf
+eYttp/ywoky+gEgxIffC10Km6E3du5nxo7v1t0Jn3X8QY0qTxFDpKJrZTkTQYq9gziKqyhbA3kJ
mKcwVVgv25fH6mwmNwNXlHp+N2+fboGIpgi4q9A3hL3I+cfXrJvvDx2yLDzOYhC9wiKBOr1oTm1y
XTQsSi4hGlRakh5zzKyJc+SKNuKY0rwZTsZPIe+dwj+riAicHZ3vucHF5byBjJJHKGFzw53AWXy9
ItIIYKTxDQam8YJVLcZGA998S0rI7yNmxIWkXOP3PgUgLlZbjRWEg4zjRpXRcetaSNb9h0OA/+4e
I1aIPxy9igbhcxzQ4ZYW+gNpClzucsKFS1QOWSkkrxIeNzPLCqTZcJ+Sfx9OpptZ7qK9UIuSOjMQ
oh5AbUgXs9WJEAOfGmDRYjAjIDixgVUocUjZ6U9lssLifNTBXKB5F5oXXoU67NdcwdFVgPCo2Pdz
ZlGph0/LEQyGHCEZZ+x9HQIITXuJGOiI7WfujqGzdFOnUnXfS4BDyP1/BEa77368e9JBmTN6MxVS
GFKpwBXbI4TveKzuKWV3bOX5qnqfnU4d0U9/k9Lg0eFoWuXO57z272w3UvZN2J9WAJBhoZ0WvEMT
K5nuwpHVwr+0bPd0T9hqmErRNWTqnGpw6Cb9T/JLYy4OE0OR74+V/O/H8tEfyAkt7HcUS9DWvcGN
2UFulIiwIreBBhTYNTIw4OLBDMjbYn++IGTQd4esiMI3ukwMhSKFUZr3MohtMUQyeuWcgP7aTUdg
JC+KypAWl6/GYqqLGcBfPmu0NNVQmMXnYdr8KA+7ZBkfFUbNIVAjqkVQtl6sZfLhOo4fMXF5s/GO
28uat2f9QDeKzP6E08VcZfxTjNK8yPljMkQOMdvOub6FBxYLeJaN6GYS1tO/GAwyP1SnwHi7Y150
bS42g3IjozOZkCFVtyWiy1GcFSuYWjYOWlz9vOIsCZdf8UI4p90iW13wAVXTqRoWW5idxs+EcRui
nxO8r59rwXwqU/LKc/78gHzEIKiHU0rzdL0nPjOEz9EIxLLWhd3vLhWwHywIJIeMQVsUZvyJEjbV
P0aWHwGFqiZo3oZpzHp0alP5yYqkjrQDHqpF4EyMGTmfOteo3NRbcMNLpPGnZDa6+2Gdw93gYvVu
p03Djsjtji9e8cV9kPW19gquqM+3DKhUHUHrZg0I15fJlLWiRRKm0NxI1iNyzT75VPjucKMCRgSO
GfVLMGWyc9l/F0K5BH9OPimAzJC/hZ5t/hPEGiPEcZ/yY/GfZJT0WY3DyUdvKZ00iVEi9cDBqJKO
IrdgQs7aCqzdMfll+g5LUdAz/G5p1l/iCTetJ1yBy9RB9U3nFL3XjsqFefUjoM2f0nHXATSfetMY
IlrFzNU7vpIeg8JpxnOTjq6yb2JxnKSivFh6EuFDBPZ8vlDA6zpvyoTtJVo2+11zFEFueWSqy3bk
FJJWjZnDLVki4z53HeEA7YEhGlnkOithtMNZuDpvzkd/8imzEoEDaoNDsHburVQ8FnVxSeGYIk2I
48We+avtEyGthj9GiELhN6DLqMsDO8yRRtahUvItnDQIXWrQJ22TOFBjCShJr07HQFk2b0zb26mo
PPDQi0mYEfQiKO8oND0o2pTU/+eEK9RIxAKv4xAOpqQXVGFtmBmlaOPmS2tUbnJdod1GCxdPX/kL
vaQ5AQZEnac9SR+7NnwPfY1Dk+t3aB+QQeQxGfBPJeC28vpyu+jQjKqaex3QxLpJNv62/RdG3GnP
hMxrGqCO5vK8QG+G3J86/1hmE51Jub7Bc7SXlmAzQkkiu1CFP6UdEZw4cOfeZUb68XCMqtudWyI2
5kLkO7p044T/br4c34IY5NyQ78ZG1RdlVs6kmjRu4npbXPojSQ0wGP7bCClQPlbNlB1XfU6v/jhh
9CB0yZLCWnw4Ams9xgrfNf0PqxcNATeoi9mTlLz+zc9BlLwjtOETTIW/2KtcT0cZTnJlv39xHeqP
F0QcmZ1Fu+0UUq08TsOvlFIYhrTLXXAkRT27gOm7z2JaJOPMfp1z/kxaziaAOjPRSJI+codEeVGJ
6N6iWuwtNCrkgNi9yKpRngSM1U6BMmUu3RI/uzvKYUyiD6j98Ij+styEB3DL9akyPL81GUUGiePO
guRAE0Igg2mTkFDlMU42k45BqgMFKfbk5YgMq/YmlafESMnelVoXQNNCYq/xp25TWAcGYiI9e14x
azbHkiwfvNfA3HFHtuCGBnjGjMCqQvCCYfJDe/K+V5V8ShXY83LKIPvCQwj49ftRsc0VgYAb3s8t
0y4QjLLgeobllEckHk6HWP2BHXmjyw4I/rvU2mVcx4tynwn/OnlkbtlhhnBqWX0JrYyEckoPH9C7
pnB8IEa3KevRtzrbSoLGHsQD/QK77vHAL50hm5MsDjHN+RChxyH2J/Rj7HaUOsR/rzTYLTY0ZCdv
lT8F6lBcUv1Po4yCRFsxKYUdeYmhZCCb0W9dHZcxe06eWJ+c0Vsml5S8a0gXSqsolJ/HyTsdEL3y
wPwjlyhqOrjY5oEBN7fmVcfr5dVSBdk6zE9zGpgTJFzcsX/GorYtGI9+usE3VoDE7hJEsrcXbukM
ITvlRWRkb3bZ5UvzObSeiG6UuGhmQnSEp/v1ndUpQXPEK1rL/vlmlnkptFbH2/FFpiWGzjvHlX+T
gcQH+3WQczQz0tGRXsUse9gKU1H6+54Iu/V5Q7CoAU/eysmtwsnkzsK0jaY73Wry8kqkN+0a2Jdp
H/3R5XgKz8T4/YVPEw+iLcA3XNK3IwSzOvjwqD3jOx6dFoAizfCCkGCwRloSIIvEkn1eKls3+Bzn
Z0iJIJob8TsnblLE5kzzJ3qgiYqAOXTMau8UypI6peTzw//6rEC4IgQji0DMLhh5sWoBFi02wHDZ
nd01piK4CZ/8LtWB/oIrBdS/Cdm9RI+uQx11GVWBpXYBs7ZSPw5f23sJPmX+bMJvlszysUX3UmSn
Uo/SoIpS0/u5HXBdC9hm2LObortKdIboKIEHyK87OG/7ViSeCWdUcQuVOF0ffZzDJu7UvTF6vW8q
N0BYgweVR31VtXZ5a+MSof3lcNzW78EhsPB0k3NtBsvOyynrtZOZDz5KC1zdKLhOg/B5KHKSVnzS
1njbdZ7TlkRS7WohYU+bLDlfaiG5mbvigT6QhGCltwJKRvC+/FWjI7v0+EgAlrnQfUZ0UxqXX6pi
b1fa+zD7fSGaEjkGCgSW22cVUS5tWi7gNE4Pvsjq5iBAHn14I19vxfM5v3u1H66tKzhujL5BKOY3
vZzvqzjREE/HSfuBFKFqu0namsSGeVkiWQPM7detOb8O6hDDCxT4Di4rKNJX2dRg2We1UHFKjd9g
hjim5Wy8zfpeQNEdYhqxeKYeBGFbH5MgnvECKgHBT9ydQRzsIVttJrZPr8oPnV9g3bKvl8dg5l0T
vo4nS3aBNuejhHTeMNUof/Yh58JiQJfyS5vaQiF/nXWO4O8U6dM4aVjXi8p9cJ12VmsLESei9uJS
emjoJQSl8T2F0xwUc+b0X2QDkxX5fH2wZsLvb9fm0mCJX0E5ca4MIappTBwbb93mykdhSUAtOmGX
Luoc6Xa3dOoVI8buNkYhUc/dJ0bI/2iWYGNK+aa79Rv0L9gctaRotojNas4xU5PQJnw0iw1d3uFW
5YUtaqPZKHZbZL/qNN52DAGHIf0rDUtTBAhsJ8Umupd/IiCtgr0Rr+URz4AU+EFh1TimkzDxzesH
F8VIZVrNTmoBlo8ZBSY3R3RnF7DH9sDViR2MyrD9oHSHpY/6LrX4ocXTwiRSlU+D7c6k0EsA4zak
UT/0kC87xhDXxXq787Y9fZy8o4NMDTYjSbfvNyjoMLm4xsqu4hTqpjOkfG/79CRZiCTDK4Apww68
A/vf2+/F+Hl8z3jiHiCM/GSbbK80bpl18WozOf17Tp0oXOnTye2tSKovgkfGeXv0E4MxT2NYbRWj
cjZrCKSVpuYV16C2KZJBcnqq6XtoFq6szb4f9aQCw9jp3v9XmMOPGRqzSvGLAUTPRDl0pzFLDA0a
5WcOuCW+uzBtz6vGgM6Re+XTTXNI5vUhFfeVKwwTNkDCjF+kredauu3eZN1z/c+WUemPjJfUD+rR
oK/JFrFT5oE7zyE5uFaxaZ7cofb9F9bRlPdrGHPUD1kRKsozyKhMjovzp1jAIv8z9P5rIvk/aese
d+3HHdyHM2FghWx7eJxxNkenX2L47OAnjaoN1LO+Z5AS0ISFIqeSCwruuvvpc4JYbSRh4BrIc/5j
p6GFZc62vQELJZwrvPx7phbP8S2Nj65cKOwrvQVhz7OEcnrdoyhUt3/ByfIF0vlQJXbd1vNpilPK
0TGYPcd/Owrx2moMirUtctsEpqvNOFvq/CvOBzwIJWYk8rd5d65v2ogWuWn+5MdlkOw3YaUDcCRL
S6+pTmSK00KzrYQPKnvaC/rc0G5LIzOyTdaXIJpq9VZMzg709/oiRIC5GMrRvG7bSqFSLv0QPJ7M
6nCrUoVuiIAVoABJvzIXbVcZqfQ2co3cSK+Ds2/J9ZXkHryssJCB8iME9jE2h+c7L0kmmR9Wz6wg
iCjLArMc4wdZRc87BagmVr4yanirF/s8fw8GdZ1Jd8ewihTN523alO1lJ+ULBiOMUFDCd/XEi6kw
Q2csaCDbXY77tbtijDdaKUvPpIR3eLuR4NjXIh5jb3YfwjmO9BXSvQSCjsly4dv/bUnDbecG/6lW
N5c9pgmE1EOsZKC5x0OzNNvDMAjXMVS4gUd+28fYg0kH5K9B2aa4itfK6/5gsO49SHBmLYkgeDVI
ywufZnG/HoWvmrQDNWExYlEFy4Np/rqnfESsPbKC1Z8Xtl2H17sF5nGw9k3B134AGWFELz1oWinJ
hvW19frqojKmKMX3Y9YRXCNwIH6pg5uOc0Ejar91/mJzRYXZPySFCyRYQ+GUITc5/Qhek5GDAEsm
d/yFPMVYXS0NS0mojI7VvBW8VnlIr1Wcf2h8Qq1ZaZP8XryEO+phc8MCOxn9nhibA1mM67pmSn96
Vv2tO/HG9o7iDLewySrwwij9g+B7G6+N+GyTIMHej0ICZE1nGmgwUyGJAkzE+38b7VDC37tBCyYt
l/VQrNet8qzbSKPmf1rb3uYUoOA8jBwmJj5xb1wBkRQoXmp7pNceTx/1L6criZaruGINx3+XPUyU
18YC2tn0OdDyuKIY0m1yYgkV31P1Oe7ma25uGv4q6sVb4yXHKS9I4VjkktG5i1Jn6vnXIGX2hHqE
MQBg1AvrPYc98LK2JAMeMuhzrybEnNTaLU4dV2ARvYMoMSYmJaR6o9bDl/cKTML2HBXs6y0a1kgy
v21OLErgi/FUIbQeeZ8N1imgB1ajCOajKYeQ0/Aktp2DXnXk82FPF+Pn7b1kPybb48cdOh52WdS3
pH3IcXHIHxzWMgWysP3JoYnDNk8vx9ERPvu2wfmKaKjxZiL4HECLTjHDzaUoMBNomBv8JrjahxML
4R6qrh7/Ql1QXfpukkMfbkWntIbE8bRi2EamppNYqXOFXHvjfPI2QOyxpdUENtYoFvad9F4J+Vxb
a9f9JQPj11jmfWDuhoIhquey2kMXihCIjB8nG+3rxdp3zaKh4xWF6xsoXqCCqwwoifJXMf7H+32L
c/CPz/K4zG6RlDvPlElS25upUe2GVs4FftE9ogvT8D8+errHEAkhR+JTp8wBtAvL6ssxWF/hUJSR
aW2MmIx55otN8x79G0emPCjPE8O++i4H1cDD+OQ+x9lYYfRuvbD9qQIW27SzQg7SHRhDSK8/hpe4
r3C98C7ePc+jUcb0i4fq8IbnRHJu3UlxF26WtuBVi/xj2yiJFBaymnhv057qAGm+4F/5d6C07Ub6
uPphmUTdaH8nWhMsW/natDoEKfN3XDdfuUVqfPTmZKWVALr9fY/eKs0lh/psXzGdKLysRTdnpikn
ApP0ATIL9I9J0l0bMyvFN639h0c01PLi6FFePvRfBTZ9KsmcuB7MPG+R3zIy6X3JrAwTDKQlu1Th
b40Inec8E9hmVgCzCP14ttReWmT7XoB2Szsnvzy9JmLmDabvzruGNHJW57+eDY1TohHCUG3aWyw0
blc/B80jn7NP5rfVyJQfFy19T84K8PPIq1uErFd5q0oQJgZEcWcuRkUGxtuTe0vCkaw1Tro5UXeT
z49zQGZ3OonuYnqTW+fb1wtPj7hDMioQdEKMVuds3Gyn8zSevYKeAR22w3U4rErjIHZngYcBV7YS
oaMRkJUyDd8o4wCJ6ACQo1OJVnYZ2Gt+bV8xBI1TF/8Vze5krwxzd90dj68oOu3PX59jE9Jnium8
1O+XPr0e7uBMwV4o9hlGbPXjUfHLe5ONC5eKk75OSExmy2haDunwW3tRRUvy4Zp+j9WccJGKbbNC
4HW5C4W1+rWwlIFz4cWFkShOf7Gm0pTfrnsNJY8uPKmd5gk9pynfGBclq7kdB5hadiCdRTmgqgsA
F8T54e2Tgl+tStu80WM89pFAWQ0LYvhIHKYSwjO1+qY5jwJ7DmJOqBCf7gPO9ebah6nT6ajlzYYi
C/4wXssEgAcChQBtDakT8wJeHzgbNhaPo5/cg3jLFux3jhiGNgS5dxT8OYfqgE6ti1BfJ6h+se4B
QQZs1Clb73SJUHv+QBXb6JO22JOO1210zwxvep/7AaVZfiupg+PQbk4eeYvkz2PsJNUvIh8LWLRe
YsZNzC0QYMB7hzD8AW0kRVutf2P14TCU3dlfc4IpZnr1o8xASUQwiL2Q5NddHKD1CeWH8VJfOjMg
9LVE/8JNxFfhDt0cbHW0Ru/s2bp51UI7BdGw6JIhmQPCrt+v0+iKwE1xd1Xhdfhrk+NXoz6/+Srp
cCpvQ0reUn39DgSS4oOcIa3kttw137P7OiMq60TQbMDso30sLBpCf/vPqMfc7ngu1KuHUaO3TwFo
qr4/9LULqV2ooHCb8FpUajyTm3BAy8lFzBhr6J6Dza8W+eJKtKNwDQgOuHRAXu3BzvdHlno7xbwL
kmhgFcmpd2WEOkhgm5qj9ls5TKKnN3N4beQJbXdTxyEUXpXz2EzQgCZXOlW5Mp39PNQTMyFPphgL
b46d6AUB94Lz44awzy7k2wu4z7XU6IXX7yPbLQIFFmm7vwwMfbtkf74XxsPi072cxGgegS4I3djZ
a4rV0F6q8rD0PQnVk1aeZHrzLmpuuLcPZXmlsCbFko36jy9C108P4YjivLKVKMdPdzxqqdPKXeg0
iOslEKnGMJbahig+GhyNxDByCdAT0JOCJQu5Jg0Viedqk/O9z+XKUyMepiRbpUMDiSOUitHWHv69
QtL+OGh2Bl68wbfoNmEfVLTdWmqZYK8YL+UEt4uxgfJvnmO2tEO8yCqWU2Qi5nDKhaGJy5PvfyAE
XO8fsWFz5UzxlUPrm9XkN+xThHdJan8JDIWQZ0qu9GTjAPwqzk6UJsKdNTUo5RPayPN0BTTIi8Jm
M874AyUHhEr+IDYib9BAD554RgW5xLf0xrdCtFm4hdYcqgHRLGAnXYbc6Nh66x6zv9nuk4bYooHa
VZDJQiRK4tlaqiAzBmxRCXpTb04AhxwIeTibtMNxDH9mcx4vSY61EPlEZ+srTzzzDv3uwmBZbet8
biL/j00/V3GFSSYPoCEP0/AT49MNHoqTlc9PiZ0wW9E34z92h+p3N62NZKyBs9GN5iSE+2bSBfor
Rwntdky+7h6KRRpqK4U7vhMthRcbZCnxhtQ0tud/zib905rp0xUAbXxa6WbuZN6f/9YZjIDqNvcC
332Q8JhsVlDb/5dZKad3KW/ILl6hLHa+iPABMy65TF7kCDRVx/X6cvLi0XsLy7tSF0Sc7JdNkaSf
vR24nruwhDCUc8zQ9eCTYjUERvRjc6+YpLLmQHuzO0S5TgA3NThFyg2cTSx67IKpCWcBr+YuJAmy
VWNJeN3LUhtibhAOk62HWQ7BtuMZfpsLrQa5Pu9dkPBtRhyi3hzxhrO4QpG4j8seMP+JH5kJKNqj
uIsuxzdxJAFuDymA2eObZDaojiHxQb45GXSzC0lMtqr9cIWag5f9+ZqJyGjDQuTvgNeq46Xwvh8G
WQ7CQEti8GVeO5XRTI84B+3ezRuZfiBzkQQR3Cnb5vR+2WOQ+akCPfTiS0Zi8Z0OGi6oRKgh1q7v
O5RaNPrh62Hj4GL+xkH/xzKIulFJCOoR8NPEulXgYgeFgKDkgH4ZURmqZgmliqRYqOC+0owpAoKq
ok3FaMssyBiYsSDpQrElgjIDKqH19xxjMhjMYcUlNVTz3IF31RJLaZGJYNOnAiQUXADFGuJM07ND
N2OJeM5y4LdwyW82KWXjf8qoOQVg11kqtI3a5PIx3xPov6HT+G6obTLMxZ/TlmmuHn5WkaaDA3g4
tdG0j7peuJgjPdniQVe8gYljEqarH99g/7oeSbYyQJSmul0JAtDVfgrHfI5zfQjgSH27Fan/XqGW
jmEFj/bEgh6PJ2QqTEITjRxwOPg59KvaOwIHhPmV6NA9hAg+ZAdW68uxcPDZJjNLkZ0eNQwKErKp
qAAWhm7YwXi6esgH4XUDjLj2oTKvvhkdTicVBwNhEr1qjYNCKkF7nvKUrduEW+oUbwIBUV3ToSl0
iZYxzzdUc4BIrM2AOSWnefjjjmrCE29ZONxDKtdkuVDQjEhgqRd8j2zZBAjk6S/srgrzh1xRcIjj
4DrPPeZ03iQIQr86qG9FiOZZzLERYoxKr3T5j8elsXZjEbxkoWD75qMA/r0cUUTllGRB5cDXLP53
7AU1HnWkOPe62ovd9/FdbDsVsCGtSB1KJpeU/+vK8dviHP5kwN6xIFY/Gc1GdTf5TNNJSZvNSwU+
xXluCJWLhvnjBtPDCMSqmYJMx6mTjb3fTGHSWTI2RE4Yt4Bni0HrsQhZ4W8fJZylzslFcYG8+ubk
P2V61xPgtUem9CIwrRrzgykOFEZUEx16e7kzhx6h4JcrbklVkv8qnm/wqoReKg3dlWaSLPdqkK22
goCHFCKKPtd6bYho0/lvAZBRQlQqIQPD3xkzpCtkJSlhtOwy2xbXtCZRyJOe/L4Ge85R7WoQ6R5t
ycFDx/Xfw6xOq6/WF+6ZFzAJrs9Y2wxsiWic2x6jspmgQGm7budWfuP2KIUVQhlwGhm3K4GXMcx3
JOElScOk6BffCfYSvuLj2z5ju1/KjwAcLLYe9HygJNcXm1ODQYSc00NRkjxuTuCiCQLmPpgUexlV
Q6DLpndtbP7d/8a/khR41jOOpP6k0kB8JJQrldepiLxzGyA3OppLESNFceFASU+8Kj8pSj6TTKFl
EFBCMDXjna3fLN5Hctuj/ak+8a4/zPviyQZn4nI0KnMTNYYVWH69BMHziApndhh9yxVdmj1URJ5M
TByK5hpbna1TZAUh7daeBqDKSHBuFxzdBMtknvsMMZkarBC+QGdoX31I79BKMKf3knOVcKCUeRvJ
7W4K0+y+SnuiiV+tr3o0K81eW5HtKsw9XXWuy+2xw8K2sQLvrAorLC6MKFEkZWmYO/+V9MVaXfl9
a6MvOp4X158/pX/mOXS2x5HkQq2M8sk1TwZuJAFqLeEtWbSAe/spqlFTz40VpZ5OPJxMOsSfYWf8
WKUeWdhm3+C7XRt4d9Bh9jH75GujIMDT8aEw2UnM+EIXCNR4zvO3y+Y1FSPwEFcMfsnx2fXzurxS
+Ref4Jj0iERrLnuUqC/qM3j2Z/m2Qean4/pKv9FtzYusiLsSdOY8ebOzPHtdu8dOdETa0iAVVxfd
9xGApXTiCpUl+F5by9TOnLy3dlyfZbsWkzC8J+BJ5LahpAp/AKfNEd4bIVI+FT502Vh+QXtv/cl9
phYap+TjyCIPEtDG+fA6YzokC3pkc9a8c3c2zBfWzdbvE4QspY1E+hGRM3FLGNa696IthVLQ7nmm
hIt17kneRRbZzWRsVNnoDybx7wQxWlPqrh0RjhXwPWr0PnH2m5f/YwQOO1Kv4r5RzM+0QtkkI62M
UwvUSGRO+cqXxFkpTShVxLlPA467DTPW/80mCKzeeF/QBxxihn6G9moAERyPQpKtuluRycyQd1fo
AIfyL3mqvmQ/AkxQaXFw46LAKBAIxqHF+jM/imG9djtEqEaZW+jzI+Ht8bELs9ELYcv2BgVK8wrV
uuWNItp5AGzL5yPuHycnSVfZOBVj/FD5NVdBMEqMSIvcv+Pm9Axrn8oaeEydt5u8MOQojjRCS/kt
5serB3xD0cIf3QgxWkhkNBCwUEK8yl1jdMSU1RhU/tvGErOeF95oAF9mdY8cbBdc5rq63h8rtmKk
9iiZgeO9UPbHiUcJtvxs41EuLNBhdEZu4edcof/7Fz/w981KDpcEtuTMap0J90V/VyF2iTflNBzp
HY9qEJdhMRmfURGpccJ+VOrYJG+qCjF9ncqIweHe4ZnCGzTDNMaBW9sFCb1lip6Vtqy4lNT4PkTY
CMc/uoZoMF1QA9Tw0V2GTTbDAXlVSPzSDHOIX8CySfANXw+UvRAOcO+DvooHH6qCsNTT1tpVaZ8X
7aU9y5mJCtfx/jn+rLpvr7tXPUJ6lRcxbwTERZHnKPaBN/9pVVNX0kdIPKtEV2QkxPbFiCTmuFed
htQW8ScFRADYnVK1Xb4lBV78FYE5pSGeDOdC/8lQYW4wlqQJbnHt4dnaT7lnZdSXILiRQYJTnkBF
SywHbfh4kkigsrNis4U20xCInSXCz1vuIlRwTVY1JBjEENhxhTaGEC2R6014Jol6D3jrwMANdEOB
RRITZC4VL54CC+Y5+AkZVhLG6+2uy/5C+/TVh906B4HN81NJtPMcgojQBgLxk693OmvYpHoBXgP6
grqJ2KamLf+VJ4JX2QMxu0We4RXmc4PHPZ4pSGoQrtKswOJbF4/tvTUigJVIQFTHLftGoMZivpE9
PSpWm3Urj/TsaRWVOLGEJidJHLGQ2TcE7LkEl5PHJk9u1VvuGfhfLBfoookptLYSDxryUTK4Qz1F
ABeS4gCwwms6ousOpVj+UaCdtv0PINeE1YtNYyWKNZDtDTz9CuVKcBEKKp4TCCsutrcS+wCt2syP
DzmFiri20s+iV4mN4CHS5azW8ZtTCCY4jiWehGLuAQOTLVlaw3Jojfo4gOdAgTNFs3SqYNWP65Fm
6suIe+/rbslRcefUjKA3izc12GA7/Df7aumuaaCGHf4TPbD7ATAsXe212+0AROPxANk66WPAPD7i
+ZYHMxN4INf0enHS70WvG0/EXoS5/7IStpFEViNCi188oza9NTmu8/zo+CcRaSIdlIDKPCca9SBQ
BnVLk0Wg4Ig9jmPTVMMdYRmE7O9kcZTA8MWIzfy+Th35w4thvWMUqdjfyxsM2QCj8V0spkz+eCcX
L5KNNoVB4AuhTH1HvchX99hXbYTDKshLql7lNS3QaHvFoc9Cd29IYctKwxGnXElRm92/brZtG5aV
hamxUEg/ZRKAkSeU8bdYFRpxrNE+hvDoYZ12JBwWSj2uN2xVbVY75URAglv9wtFZyHkeCq5u3nB6
aZVdAZiBtcX6vn359mUWzMXUpsddJ3XxQzHsPv/O/jKCRR9Yef6XO9QH9GV5s9Ni1NgnElzcXHDv
SNwaFPTZ68RaF4JVdEalrBj5ASfscSZqWHYPOsrlauiSUAchHSvKOMmG6N1wyTgdE+wOdmBB5P1j
nHX2ePa7XMH8eC9vLp03pbed9dl7XImZ/A6mROdfmgtv1B0X3Sa7Ews4F6V/6Khm/qYKuB3TdH+f
o2fR3HIbrpJIY5jU7HS+cHUWdErKvvvAig8fTM+csYrIDW5g//yhurxyLsxsYq339GTT0yDfGZGI
BkwdKDMJAcVcXFcbT07kPXr7MmrWr4i3+RguPDaHfQ+UkrVEudLXOmoIjtmkc1rYgb0hzRa/I0SW
vouQUJpJ6bc4CosDj7fde4Uz0ZuZd88k37cDfDRLYK7L9sUZajo6369mmmtfaPOzlTttzzA5lBX8
bYWQWRv4+2xZ1ZTq7FeCqDwvktpeJx5rDNTbzMjumOaGbZYaEySnS8PNxaVh2kl1ZGd8EOe3unOR
M72z6p5R5zKXeKp+O95rYgk4an+j9o0AZ5Mi99pRtYCHthQQuCJSEgmLi7H03k77oSwJ2XsPUOn4
Do/GANq0PQBmLTNsmRtaMkZk3KrvUYPNfM7cAGi/afDTeDjP6MP8eahor9Fh8OGagOZ0kXY2gIw2
G8uhfhxFsBS9XfkHDWbhmkbiTUjAndZkBHyjpq6gcR84+yBbtZR0Pt1gNMJFYHXSbznK9J69iFUp
/Nq5bgUifHmlY/SzKAzcOa6/RjCEJnJ3TmD80QsHDCgTUAYclTwa0zTuZuMdbJOmJhQV8IRkDUJl
AgkOZkGR/1z7mQ6UZ0UM2w3l/0OM9m4VsejIFAC2uYBnzZPwW6YxSYYlDeP5Zj3Bq5GazO+GQp1w
bvckW3bsO6lIB0g9WMmODPdMgwJ4FnoX232ytafXf7KNviEzM7hWIZxj6nYtlGJfxMEauDd/cSC0
YxKzN6xkYV6QnwL3zamD8XBpFVuIRJhaRIuFE0GT8p5W0L+I8+NGXAkuEqc5IZJG5U4TYv3JpFHZ
URLyMY3RqYRiEQPluXkeKl856CYNCSz+1QkmMish4tkZeB4A94A1SOWuj6AX9esZPeqjQ56h3iKB
lKSWvQ76yEN9wQ+oNh6VCHdM1fhIpAvaH4uV4Qc0evqKvPznWQEnE2DZlpaqBJA90WVZX6yFqVdZ
vCXiGjG88W52Q+iQ+wflvNubDSllulrsdQBhDOjEZQllDdcOKc67qoveJH2PYdyz9jixZD8OPuHf
Ewd4RlXtOEYWMw2ycL5sz7Zuh/9w39FqYVDyhDLZOD6zAOfKWLCGN1zqlGZFEbce/pg8ghwtt1Ne
LH+T2YVlCU2zPqt2FNQM+POb157r/fliDNAxzcS8wmi4NG5ff4My9l4fyWC3oTsuKK7nvppNQg0s
LVWmJDVtZlADrDwTkqsn40MFoUwxWDZ3kSY+eENknKpeeqGOBAvyZRljLIT5Xgxzw+62XaXDalnd
YFdnHf2RneEtqjMaNlA6ufSduqHcuK7ZvzZdVpTL5CZcEosBO99idW6TBDgonRWuqCIPXvnmhxhx
wm9+NwNRjBTI9xDNcRGFUCjRX8nrUClVra9KxPNH0o5T3JALjwYQM+G1d7hFBL4XPB+u17MemSBa
gRCI17PeNlak7r3omfr6yTyAwMAoKWyUPwSUYD3U0vxnCZHGw7jIteHvSSqVkFx/gt96Y0Xs3BaZ
r+QjAB+PbzH8tV9qZg5ePORdVworv1674woULAzAtPlTzzVF+JKVJ0efTqrHDDnF7mC2CKY9EBzl
qVHPjQJfziNE+6J3whsphG2QQM58zKgsh37mR+wCTDcoDVZ0Bysw0NuVnVRjbi47T9NrPPf2bx6H
LgiCGh2buhcSliFLrT/hp8Z5m0YZ3pDWF+qIByzHGXs7yg1kPfK57ZoY4tULr2qia6ycFIECkGVp
mX6IO23KZeWAJBH8DnoyYbSbVtBBqBRw3eA4MjwcJOHjPdQ4B6YebHE1IJdQEoi7vsFVdw/2hfV2
9g0BYAPIwikYOZA1VXzq1tD6BGAu+R3TPIJRKAb6fIH2eLA4RWHXLGFXKjgmIgAJfGSFX9M+27FH
+1S7Gi+57H7siGJBVsHGW6UTHu5Bk9tktc9YI34yW638bcfMTG2DesMapNxZkXdpq6mj9p1/vcfW
OmJshGPrYxGaCyADRsPda5AD+hUolAS58yMw6hEUnozZeAnlVJnxRTtJpnKPoB7k3M16B5utHLyH
y1/6FoNsHkfaFOstOaykXxjWNhOFsxi2vIsVt2iYn5eBaN7uFS3gQeQLs1+dhsn1JpvCEsmDusFj
Uw/3DeX2mJPkYJzijCYWiNFiYKKO6dsqQMw0nDTK5RRjQE5uH/fa5sAIorwzUxIuKi0h+p/Fh9Q0
7j8FIqZCnyu10DCBiwIiyuodIKhSZPqPU0cRNk4XpBl4FnydemrgdjWVWm6qyD7zwpR2VL57xp/+
9Pxf3d96mWm7awNhidTvQ6z60a+EjnaxZPOeiuMRsydTo49SzGfdXRBieAx0PKmJm3+YeVW6azqO
0qeYE9Kj7PKYkXasYA/Zfos6xL/JKsgNflGu/iAjE5JY5OBi0zzb+i/bVFsmF9dyDvgFf4ssl6gF
eNnv4DwW7heoOcmul122cuk6dqnGHiS7nKFeCSJKpZ0/Ck3ppNURPmtyCTp6uTh5yHaIqq9wyBAK
YSLrJkW1diG3O2LcG5I6vVKWL0U3uCdZUJN44WD5p7ipQd/lA/I/aehwm1geQ9j4d6yhRlsNwjQW
dXs0dmlyMuUvNL+z9xMax273Rz3zCnTjxcRBPIlKi1S4w4hlpAF7RzOuhnapMPxSP2bRlQ0RSLBY
1R0JUPjyVjURfpm/iA0ENF/AVhaLrUSCEZ9Nxnmj1yTq2X1e7fHYVm3HRp65OZw362MqV6tCYrmx
Fo0f19VOe7+xG1gmIqhqedimgwnvKJ5I56GRKuq6fCW8yZJ/amSQddWzZB0w/A60j7Dq/Y7mPc01
VkcanjeDf1ZsbNdbZPlDoAlM1QvnlhOyZENLCWpW7QZ8vqrYaUWH+/kGrzmESOdkFyb+Pzd/Q2Vr
/+v2AEpsjJ6EC9wOqPU9un4j+sXgLci0H41zFhSrhx+kFlVe8leU3aE02kX0G49260h+/nzZxHTm
OSgE1cpXBAeXBrPCSLmJYQBzuGVlo8xdirlbP3qOZjosClGhkJb2RaCQdHl7m+7t708YB5wOyDDZ
nLZ5A5V2yQKZk2jK3zdHhMtDGObXWwM42f6PRlIf5ziVmTk5kgIUJ22Fumk7jD8foOE65xg9qPeQ
4FVtT+zQruCII4FvibOggAQBaAMY99HlQ8oZOTV4dzc/RgGn3D/NQROt1hLnHpyRvwmZT2hbehSb
P4GrhcSgZ2QutEc4bZLCGoveyevSfEVOmd7OTgGPZROHFVYddzpv242+fQMPokwZJ0HAR4AGQt07
/tsgFcz/b4icKphmkhUPX5NpOOsVAzqjF0UkMfv/w1OK0xlNOb/RWusAKsgL/6uU1qCOVmo3iDL+
Mo4Ni2O5rqTelYvf9dluQ+jx7hN96U1Q6xhm3FSxt1x+VVuTAkw8fB6zDPGwhBcuZDRmk7ugKKlI
qadw5wT/J8V8ml+bzMHHI4IIGtRLoVfXS8AHl5gBfXkhWmkWhT5Xj8g0CfOi9Lj5+U1mN5E52ek1
QQ/dRpFXkNtCNm8o/jENnELZ/+2VrWZCWNhd8Ey7cQwUBZyP3N8mSginOwnFd7OiyKt0c8Gr9kyt
CJfzZp7Sz4YjCIsAyBAC0hR8h8ZqXU4j3AHIhI/ERFKVf/hq66eBnTFN/hFiO6f29pCTQB+lnWRR
wteG/7G2UDY0hdWuom68h3fdifujNRgwnED9aWuLT29XffuIMcYXzOEeQL607zP4y1o4kzSEwgh6
NdqWeAFg1lgZGF1qyJv5dPSBuGPmC5l2lnvjApAwtWhckcfPjV3MiUYBz8Aoo+IBdUujxwyXUCjq
k0FI59nczje+/YvXVA0ZkMjCL7iyaikj3EuyJ2FVvW/rPl5LG8/ykDDGceyeyU5r0rMwus/q7VB+
btQKYJWvlxrvm0wv9bJoWOlCHeZ7/PhTRmvp+QERBeL87M/4bvd7QVJEGxWb505MpOynuzGRKbpB
G9slrC6uf0Js35IZyBKiDjSbUInRSRsLZY7+xJic+s0sSIXwsPX9W/zeYeifN74GpElp4TTatiWo
iZvnpONYTv+Y9oWRI1YyOFzNbdSwi4wkWOZKTUVHkVbrRG8vevHnBLEcj3DgdiwuRAjkUxF5PacH
3NiTStn+pUuMA/Vtt/CmwTZBP68k5K6OmNE0qUYyTWg1IzTKeFkF1U/IAbKQp8p+hXW39iEPQan3
qthEdDrNgu/oN4Fm06u1FB6dAq/bxmPTPoGdqLvPgQTaoJxWtGYKpttxdD0OxD9L+nBIIf1L0Adr
Pb5Yk1HzZqgApQXGZ64OiHKUbV+Kzojglv0sjVtqpDkpMo4MpKivJaso/TC62w6pEfmPycByc/ds
NRtmVi62OkEwoYZh+9kxnhdxV34CdCEU0Xul/cwDlToCwggKjQnGox11Pezcen3x0yW/k1WqQCRf
a0OEfYx0r+14mFevWW+yCt7F65BxZKpl5apiBLghpkc+VqW9/BvOz4sq6cZg8dO1vLPYBkApUJ1u
C7eueFpgbRJaLqsmKSeKKAEOFa/LEdlCodoHrfpKmUNctikJevTle+QmcYd3dmPJhXCvzNg8dI3f
CIe9ytU5fgEDhUdSrx1e+OZxEFnwqjf89lSjuISGf1nYa3e6yeb8djIGcRVUTivWL3jUJWeBw8vh
ZKSMjmv5gzSTrnMN+bpJVH3WwVBw2SzrBAvZ+5IskO9CQ+aVl7GlSvagVcOC3+VBzxBo2GO1rqgI
PLC5FbYg2DevWmQIL0AS7rvHgZFWqZgmYII3moCztPANUdw+X/RCws25DPBaC+1JPooKnGF41a6q
v0XA9zTQ+HJxYD94JM0mNHVVlhiZEJdzqKAoloIVPfT/Fy8Bzub8W6CxSGrMDkksMuk+idb0Ai2H
ybkMzGa1i736xH9ITNDKT8XVvxwewntL45r/ipZ3TMDsXZuXQtQ1LR/kBp3nDiafd5RbN0Q4t04Z
gTq/5uR7KrcQ+j6XOD+bq0Wf8EkobgliUomfIUqarXrzd2zHTIVn/mYdLVfk1UUz+96SE194lWXp
D4OT/EwQKXFr75tkAx+n2qkozPfpSQYzDOdExLUg9fqEH9h94fUixaoYtuErXoA4uwHADmKDaIbg
ZrqWdBxc/nG8VdOFMmwGiLMa/u0iJXGY5/MX3+hzzDOYM9GsXy24Ru3tfqLH3xYXNEHITbb9pb31
r+UC9T3Fc9P7JBgxPyp/1Va2c9JLvfTTN8c9rlPjMtRB+R2kT7LrD5USBDYOmXLGdOt/8qepLqqw
c/bImjQ3iKYQrHoSc4pw2MRKX+W/sceGpGh72ox+gn7ij1mLYtjglcBkIO2OsggdAeBqDMF4rSQ8
6pKrgNUS290OVrqZl0K0amc6/mX4/3Qv1eDGwU6KZYUa56ieyY+AUJ5oEwSLTY+HTLhB2l/7KrM4
8LFIXqEKUeC/iy1GhWDfghoQW2V9+pXd+CMypApCeNK6ecd5RduVMl28Kpw8V2vIgGopM3jYPSJ8
eq4hPJaqi85vuYmEOQ6uTKGavXqC9ABLFvgpaNf4Ep+zqfRXXeLZRafSdPcDKi3E1Ll+HQEPaHyk
+K9zwAq9jpLYWamtGnCQJduQI8dlLqyjWk4zRXXD4oQVz4qdf+CauWiC7gyh+UzRYgTNaeZXl5Pi
Z0LOKV58iSJaVn7iqHCTxvZHwwlPIesMDBSNddDFLb+CF+Op8J6TQIqmWcC4l6X/AfQRgupcLqeW
/OJFhd8q33wwTlY4pdf9qnTIuKjL9hTNVzsuWbDVppsTEvt9sJQXf7CV0exYws5q1U6+mTOga+Xk
7HSjknV8goL6eC683+5I800t7CKGhQ5V45JvjFq6WhNCPK9JG05zVr64hneCc0BY3QYOQQ4lVMex
X7PJjtuSV9nMFTPfr9LMF8myp1PaxkbCBfV975vIsHgV2iURfK7FBRRu45X7BxZAA5lwd1w/a26Z
0qbTTOixmb/cIrGdI1czEKQQofppEnpdIJbXXuhDvcWtcl+1KPQQhMqUuljlcrm0VQnCcd3hUHLu
QPKo8aZx+FOuJU1wM7i1U7NklGicVaR/Bp2pYVwxldbk4CNl2ruIuRMvFnuieoIivGy2mlDW0oh0
vds857sJY7+0BgVV4yVm+zEjfjjNd/oSqbzEgWIBrhHSvHqJsHtaA1LUIW/Gi+c0hOR4CQxVYgCs
f/YxLzafM84HJErh6kziODAGt4Z+YBE0A3GL5p6DjidIWuCmBKNAjT6GR+/Pa5iNZgduAmGwQ1FD
Ds9v2UFG41z+MbNqua/0ndcY591UsUHPnH6ifTaU4dJ6XnJJDMgsyeBiytr5HfmUittxEZBfP8HE
6P9uoM0dxs4rOz7uoXBszV9I9Xhepta+kBSAtU9NbXq09qJFQGker7Y1WDk/dovEZ/AAj+09m8YF
eA9E34SloSovMoCWCA5q/chM8O5U6dzCuXIeBbpW/GWmptjGTYY00YxxPBmAGKAGeV98mBkmhezc
wEL4osoUVPbisDa41ryC0iCicpKYdTUATLyzYQ0tRGkVBE6AgcahL9y96F0bPtkLCkL/8grNgEJX
YayLC1n8yr3ziWaf7McnZJ1odD8FSmlv1HfJqVOYK0DJasuRRhres1C2zIG66kTqZ8XnHPoAr3Vi
PDReZ6h1wCMk07DLU0uvSgazvtiCwU69PpZVlzCqVinfhsVouy+LOedeBAENBVI8eDzCtTfgXutT
h3cEVBiEyhNzxGNlIFdLgLOlvhOV6r+tcKTu0LY/oUhg0C44ll4m/n7euMFITCH3M2MWZZLBiDvn
bAxRX9GULcYDaWOEXZ7l/vIZriuYmuUYsU5Z29nn/PNrFmeNLP3dOw99xuJi7TZYBkD7N2BWmQUl
OBuGqwftawrOmccxtNPg5psmMu8dlsyhz/jR3WdsAn2KkO9r4QHnsFn5Y6IVi1MfLYqS9rLJXF8U
pki3ngMF6hyKFLWlkqXSWhPUdgndmxWTNnN+Icaln4UWnJhowDqmQFggkuNuucOII+uOnEBcViUs
bTUzuhkYwNVtTQuaLe44krbC1v23nH2tGaHk6AdgFnT2
`protect end_protected
