-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
sq1aBEXCdXGfEih01pJvBZXWONCfjZjqCHMQ4gOyFrJ9ITeaQ8Y3pXaZw7n50GCEUr1csk/Qqnjd
qVLP4YM/rfwKMpPKk8OByWGFU63S+N/2waHuUUYQD+8bLKWfaRt2MbOiT2JOVvyHdNEqoJpmsanb
evLFh8Z9zInLoypTYunHcgnKmyaBLZAklT0azOPUBbx3jTuytQ/3UmYZXseE/naJWAkDM0nxIf7s
KdB23OXs/gnyJWZFuR7HvUMX0e4PGG3gnOTkphsDvL6GZHNvYxdQCKBw4LnxDnKUHaMFX06OHgjC
1v1SeReFKtX6odezRDyH23IilvIE1xi4Q722vA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 90624)
`protect data_block
14FtYk3Ud73pttY1SoUFFpx74k8jfMtStK6COJsJ4TZTml6c5Kw8HNoPYJc0XQv/bLp0RA9/uGPn
IbiJqiWbMLQVXE33u6iWLXDvP9SVUpc/3dXPI1tieRjKs/lCMyeAGquCLGWlu1m+NSM1iYNDehBg
9T55OXHzMMjH/0HvWAmMDM0SJGKeGFF1OHVzO30lbNyDKqRSHFjzgjaRc155+xiP2Bid3ErknLkw
NqpT+jkYwfKGsejirk/bKcxEIVYyXWFteLc5HccvQTUgAdWUsFHerdTlrQS+m4K3ISIu2s5WzzB7
eq+qqLnc8mcGDX2bqB1Brb3sQOnGoD+w+awklg5Q2HcQMAoXigpsXlc5tTR/eRigZ2ToY6mj5oyX
A9zqQIBmKOUpGcLI1UoGtN8HKRDS3CbRNuikW1HFwIZy0btifdY1e+XDPD/gmlNML8ektzwokUQv
D3kGuN652PrlBRe3EQDYDTfU9rUNI4LG+ZB7J0q6D4i00t+nHbzmoWoKZ/rMGi9v7m3qGMgDkhGS
QePyJLDGZ9+kZiTA70NmZHzhlbabfnd/0moJvQiCvckZ0dx6dDl7DIyIecawoOh1mxn5zV7tpQjg
V9kNab4Z9hBsLZjwa83gG0JJOgCKn9LZ2R2bF+X2YxupQGAyBdEokSi1nWNcmV0STybcoLAmYi3/
d78GnHHWm8kippsO12o+1+95gOwY3w2akQdc5yszUHsA1QLXL4v1PmRB7nxd4KqLeas2dCMlZWSc
ed4cAfHTdi/WqDZUiOyM0K8iiswCoJABVG8xcqZzGqdf4c09Dx9AlTnloNd9e0wcMjpowtGCPklc
u3J0xJ+JukGJ+9IHSI56raK+0fmvMxaL+lKNPhBA+Ns5M6oMtbFJUbTUeQtHlniqY45vUS62Cov0
+F0jtqs+NTkuWPgYd8IL5Oc7PXmNrFck0gEaznPm/sUFNwrgyCGXXzAiPumc8tWvm9m8jO4OBN1P
NABf93xLHRcGj8lrL4j2nwmGI8SQJvoBOWjI4Np373/qDmjVvxgiDixHZT6Yn1pkfXSX/rPl6ZXk
Q9NSNSxjlhYJzVKs8Q1+b+H1l2G7sdJtF4TBm5bgxb4s3IShUdsDFF4wAfOYb2BQXMDxqA8j1UN8
aa2lio8H6X7p9cUoM4rNuD4xeysWp44jtPkYOJU68VbnelueaFtFMF3562NYhBYTZVZSTWJHWUjj
PjTMFmrSdAXeDAOcj4NuVy4oASDsHZEDamHIraOrczTP+2tj/fTuZKRNRsYrSYllCuV1zukTOqJx
2By4IsRT+/DqueUfDXU1Rp7B2ZAqFBET9zSATRexXkNlYf5xEAzF3Kuf+ftsq4EQRgKlXTM351Lp
6LYeKrlkkKGeDrbN5Vj7u1GKAC/NrvV7xrJvtCFnPUFpOrpBNEf8l66Szz56so08EAoiXG3htl2J
oZUDyI8BIUSW53QD8ZrZ8nku2FXdypyZBVoG7TippLDrdIRVykyvnEWirw7ai3TpZ2S+f5LPy87m
/0O34XjhGqYDf5vQii7fWsDv7SoVoTENCT5QVxzDqy3GZrC/1dtsYNbfFcP5CIOgjQT2bAOjR2BA
CNaIqnTGVzsDT+d7rfkFiUGjnxyx845Btrthuh0agmM2lIAoNvZD8mgaDNpJsa9xubkkvjC4CKwP
7s9G9t/BxOmULyr8t8KTO/vAuhrMkdfFY4m+Rmsg7ZTvhzIjXlPm6O7QiPwlGPMPHpfVSYliyli3
Ma+WxQdGPkHuoIXuZRPC/P0JCKJiUcxj8fUf170CdnSP03WYDdyotmFP0MT18mAVHOIfivgVpn3A
5doueRHFNBqZJ/xPgcGmz/nzJ1zpi+OFbXGoFbxcnzdo6WPXs/EqbEDNY5xpMfQ8Q2pUHfHjBiOg
CjHeCDmI5uLO2Fp2mjZwOLDIGRAkzNTE3SQb5M0NhmcLqTk2RrhwCRPgXIGaMOIbwFWeuv1XwDas
x/A0K/tOL9+cwTWwyjaw2QPPAFE1wPHvydqUAZK3jxzO9eYyvMK4wqGRUo+lQCjyPWcoLeAVkcla
IOXZoHTfqMCO343Y11T4QT6T7Dh6U4ObSSgNWZwPJ0bfUdYgEU+0o4hJ0wK+l/u8woWdBvHGLhoR
Qu+F/Qfl3OFNS/3lNhilG/GKRo5fe0lXtpGrG6Mchq2FEes+wSxNZQGY78XflUNBz9kCAXFv7vFa
ErDEQCJ2vS5l+1NpW7embKeu/LsnBD1Pr/3BGdhIovygbUECtisSwLzjBDxG+z+80RXV1oH6Cvvq
sS8LkVT/B3QGKAfXTisBHWFL9rhTdEyU9bJ2FS5+7Iyh1sqpyAkI5Vs4+DqV0bUtklZlRqAbdxxG
JFELlj9kvbzExDDFSM6ytWbJNjgicnUrixh49kMamdYL6esHkJZ0PbvNCglW5DVKbKVFZrPIkJli
ZbiaAQ2wpf2Yoq3MkgI/bQsBvVfemqjUx0IS2dvLSzwxvBo8x+87xtrXISfJRPDhRLW4zMbRUnr0
QFPAeWtSQW2O0mlqo4yJPhZA3ml8PZo3GerB5lv5jpeZ4zlfDAWFcZaqX61qBcfYUlYQOeBsOWHI
BKudagQHB6gBm3NqmzvXmQViJCAlwsqGJkN9jo8/lEwmQsF78J75wQNXVNqiVqoWI3/eFFpUEwBf
vNQg/xpesfeIys3h5oOZhSA4sjFoCS9X+63UZkQM26FZ78nep96Oh53tfszbRoOALZsgoXGAkgCb
+AFaeEI7+jTPhupXcJzfwWUNhiz2cphpq7+n2dOceB6r6x/lKUFrpvrUn+Ao8X7qFWkt87G+UaWT
QHVZYrmG2VZuOpd9pmh8ljTG4CddKk0t0kaEJQWQEBSZeONh5hE0LNp6rKH56uCCJSDsRko+qJnj
iqJF8P1BiK99QFsmaxFZ2pNVinCfACoM/fshknoQf2lMsQPinXui8XqM7HKJzRPjiiI1lg93wdAy
JMzMk1c1uhTw7wH+5+Qz0bnIfcJrfq+8kOs0s2+DbhI8QOLBmu1hcJ5eirbQu6FSAaWTCx/KvV8g
tk6BI1KOi/5NlVj0UwA7Q1XyB+7LHjvyCvFBqGdk1dw9bAzS8xFEmvTSbvNmlgZW91g5ItVaJak2
IFheIXRIN03qGwCk08m6o00W1a+pTqInUwzkr8Bgi6vhwPAwqS/73lbVllXCD6SneoX5sbfLjriG
ddNcFE6Mi/Ej3cwos4Tr4ERSb4uM+MDzj5/uAVjamebgOSEF8fVYBph6ENY84kA6sIv5/fCKZj8A
rknVh/MRZ99Fu4FeQSx2d/BiFYjj+8HljUqJbKUWl7kImrY1Cl9HCCJesyI3/k6ItufT2CbThfPz
7R9eGtEzLcnvxhwdye36zD8tcHdBdA9rEvNL0n/1zGVH3wEf2OK/lPH52K7mGH8cdxBLAhDMKpCq
t01u6IxwSzEUMXkkSnPkNt8S3qx62MX42jIvZKNBPcSU1O+EXjEhs8sIgF/TeVznce23jKv7eCv6
ffWjNKSkQXFyQMDGYFkqY6RgtTbPw/kY4WUI1lp7/B5Dseep4M+yigSwoqSElMEO19LU0dB5VFrY
lcMl9Rri22YNGjeZ8PHTZeruSG6dO9D3NHj+DKmUXyM8x9tvhHa26DWLMDXnse/ofqeaBCFxRibs
+sw4f9X6onnFV1de8smTPlD9HT1GB5XukBcZvhHsBN07Df4GvwfyPL+p8nhrvWs2z4ocIRYEOutP
gDiyL5YSaLpk4I7vGpr/HMLGweARJFog/OlngCi6HVDzgNZ+S2QWX7Z/XeJDH0NM8uy9i1A3/sD9
BZ2y6eibmf+HcUeEm+X/Szn0s0miFvI/ZwSmxcc6NQyMsGRslQgcBxbKcgqNNMAuRXCnz4cprDZT
W510CqQ7wIkAD30c2Ce/NZBN4dyPUa547WfwCtt54ys/F2LUXsUGZg8NN7dU6HslAxY71H+N48JB
D63J4Ixkn5dx6dRJVBmByFG0cT1HQBBU8jXyqePf+pSeGqtAIWMwH3AE3Jg3zGH2ufh95+NkPwUi
j45GgnW17JbYe95YsaSez4j0C3ARLSc0TVjaZQTE4Ova7RMWJcAfMWvLpkMETomWw1w6IyZtgkou
YFefxXczNYiXO52Cgv0TnFrHQ2dlASCPP4vOb02Fi8dCkyLVryLPrtfgDJUrcFp8u9kfRFuuHk/l
A1iM7U59UDeq+lwAi88YSBTFOFdgCdSXiipzgQwsk2YNXShDEjaAeuX5PXJX8UVxN/j8TcLceFlw
Mb4GkdrZ/yvLCPmO1ULBHxOxfkR27NNlh7Q0fOhAxPlN+GsYSE5YsamL3x8hamXOeuymgrLROunF
oqfYNbAHfYjAbl8ulKiRqLjCvW5H85Z02erEdIhDlcKezX76/fu0r+5MdPjDi+3Tav0qeCeYv4QN
+kRIz7UJp1EqiPwOgFhckaWJb97HKHWirmU7aBBh2pei7Vew5bTIO5NCAQ2m92wktdYDV93TLTzX
/iPxnJM1mQGrctncIH83cic2ExkSIM5uzNbk0RHIfgGAOBVv6IhQXlfLCyom1EloJHK2OAOLZl2y
6XdNJ5Wb8hf4vYN6I5C9Co3Bmfyy1yVqCbuz6R7tcOReEdZCCerqhZExxC4MWRsA7ZL8A9Dq11dt
nzAldZwVz+ioAq0heh2McJ+GNeJFFweD0CvTdZ0QpxVSFhZ0RNNy0bGexsnqL3VUECqLHhfWHs0L
fhKazk/oZVi7FX5E+yu+g4ZSGBAWgxTdTqdTAuxFVU8tffPwrBaN9zG33k397I8aU1h997g+vjgp
/+3OSno/92KTFTqt+U4gscQI7rlnUXwcTO2V/Lk38E+TScaxQMztC+boE6nAEcvI2o+ak2c/xkPR
CN+m7lX+2RfTtk4DPU/BoWuHJFeqfaL/AlXo7dJVxdjyXk2LyNR23O0Tufeff4Lj3siVACMERwZk
v5U8TgZQm2E2O0dXvWqF5bp8l9wqU/1s58P2vrTOdXwzULuvqm00csdhHJCceRGArDtbIG65PU2G
ebUxa9XRYr4VujMcEf8M2fg5Pto1wycv8cjf4lDw7Lot4I0wUsfcdtuktNg0aBOHt/on5dyiCxZp
UMMq2ZJV64EVw/Ib9VZGH+RUey1su/2nLLzW+NumExmOOIsdtL/NAvzuQsC/WCh0eI2BVFKqFC0p
8GJ0dd97Yx5wDu7rNlvBfwnppUpjTURSjoKB4c4RtZ/P60IEMwMGt2z1zfVfU/o6moU6kZ5/7sGM
A6otUXfGF0PPEX21yS75PzcPigTMtd+ksXC9L4NRgmtV4YCubjVV/vEZwF1VYJb3jucNx1cNHXOF
NBSFr/ClWPUXY219Qe1JxgL8YygTEgwlFdwWWjbKMoy1sTYHxKlXtbid7v/7oKU24pA+R/dwe1VG
b8iMh+EiY2yXz/GdEY0XdGKwHy8vGxZOMvkZ4pVh1SdmgY2vR2fRNYR5sA+s5WrF+thm72p6fgiy
x997Z/9XjCkQOYAVPqkGRISFFxv6uw57LIbUjcanwKADiOh0O3wWjn3y/PVKfpYau2hxQYtWQX4E
L4f05xBwEWLJcsK4oL1ub2a2pKC4twd+HUh6lPNPTvEQgB9/OWRGTRx0AHmgZUWyNgqAdhRWLFAt
Sm/P1Bfvvxm/3y/dZ0YuJCdY/wtr5fbeOls9FoAIi3JjXnrTHtqPWpgco7+erBXIkIU9RDLJiXl+
t3J7Lc/yu3fTO19Qs0JUC+LTS4WTyByn9ovQxZ+dMYLRXLeLOOGN+xP0SxPiE/KW0KmZQGbW1/Nz
tjA0EoXTD62UpFLECClexNdeuWtSs12azmlmf+C2JLescW88AET69fQqYpsaVIWifBLLQarrCtqO
jMdFqLbZaV8KWXCX0XjLKYRrzs2Oxo4dJL0RupxJu6mDOwqv1ddI/dV2oGZPQkieK8QpGWZcAJfA
+Z0stC76UxVtP282vD+yXcfBaOM56osE/8g28Vgxzehd73GHVDlfuKoGE7FNUXvB81sWvpRfzuEG
/BViI/uXmB29rYm7rYD5y0yOUE2Vz+On6PjuTPdhyWBPhikFYPwO+wGhdmlmIMq6OXKEfKpfHyeP
31zUCyQM48MaYjovefDb4oee6v36tKSU9EknTW7971WyG9fhdV9j3hUD5vxidRrJwjLgY8CrPOuJ
XFhpyBP7yEXD1uMyn6TNvUEohap45QC1/5+tKkZPCEC87Yviu0e1gm3shWcKAyR8ucoCAxG8XgRB
0Xqp7mpeOERtitZZggnN0dXOy1UAsWpip8dU2mBVTCfqPzoJK4g3V5Q7tzBXIKKlgy56T0l1VvIj
waOESTcQFqiTOiR5chEbXhcfdx4p9I2IA4CzJ6RwTIDXx6BWDn+kWBQ7sRUCR6+A6V05RYKeU/aJ
bWIXU4o8N0317+CGKNzUI+sSpUGQc62gWgWoibRIiPlaXKrsGms8t0xNrn4o7NV/Ee9SyZVIaMzE
SJlLTJAriskroNMPi9ukvJ/k3VnMH2Qt3LsCoHP4NihGSUe8ORSj5Y1WXnxVE51RbyuldvJiCzvs
l9Xi3LtNdAmLlmPS/TQszM0IKS5dc+tKeZ+9dGGPVJjs821sLRB2zoJgWuA5x29dUxlTYuil6pvk
hL2nBKidqcr1lPQJ6mrQjHOdzwOWsbTsT/WfF+/2gE0ns/vNiYL48fOV8oJ0kee7XI7c3t3NhnPH
4vLUYGBlStoOfFRZJvhj9N7X7qvY7fQcZjn5WwoMxOIonIKFOpyyvCTXt/6pTd8srHXKtYz+oN5v
LfO+x9uVS8K7gQoA+8wiI5n75V7ZJkw5D/6htBmQz3V2XCawdksLdGl9g8F8ZUG2wZIahdf23BGK
fXbrmPO91vtcrf/EiexsTLiAKlDW8fScchEh+qBV8oU2MdQywq7TpsVsKIf5zCfCvqyFIG5KbC0C
Bktkq9RmMNLzcp8x1yRXwEaPTodMifxMEm/WIeGwmzrcvJ62Bk+ANIEc7UCWbJcm2gdFnPhKJphl
Nuu+hMeJ3uFrA9El3Oz/oAFD30yShInM8iqrNspGN2zPU5wsosu1Usq9pLqjLkdUr4TsnD0J1Iim
2M4gktdHNPFK4vmKbI7Q6UBVwP2LFUpMSq8ODWSp1qq3EwCHuWFFaJ3blDfwRM+3jY9e4VWZQAbr
k6FGQUn1lEBZqpb2ryZaTAoDqUcvB+G+KXBcdYJeBnLLDdiKe+r77WZToI4b/LKS03VFUZSxTQR+
mQw8Z+Ou+nN0/PimPXPYze9Q8kvUGVgIHQRC+8QhuB8eQYgZnrhrCHMKbi/R/WjciqEIat6jomxr
SFgJn6eI0D8tGCN+j1pq8XnXqyXsY+Txxgpkjf0OwpUT0QShd/X6Zyy0GQKHnkcCNKZdTA+T75r0
zqTvZFrqJgPM7mLiM1B+NZWOjoXFGI9zN2SednaTNLRpiCSVSPEQjDXu4nOmrhazBSQCsVNp4xGx
e4ZQWIIb5Mmx+A98YSH3s9ZWHZ2P9EM6lDtyF4zjBXl23lVMXPDKKm+x1Nj3o0fV7Qb82IJVPRdq
5YAu3YpQ07bd9SLuGMqBEPIVwPRDtTehaGxrKHnXjGrtnZEbgDTp2ldBg7DFe1y3gr76rrSsNkmN
SbTPAsGGSvM0dAEU76nFDeW2Q8XNYdLtNxO+mrSbWmQChvimpORaP80MWFxYRNYOnXcGBAZZv9JZ
/KCQ6TyD0E0gkfdXtSxyxdA92RV4vZNvAR3RFKVJOYDNXKhgQzqAVxkrRSX/M2rb/eO55+IwkfeM
Pc52/Jhx/7KVQpPtuOU00oitvRD0eHkt9bI819Np6IwHg6388KaG9Qc7sedc9E0ySFp/PKt/jS0p
zmqzkHdaoaZ7GCNQzI2b9cpajGoibq+LzprYamsXAteuNd5iKjirfr8FinmrTiYyCyPjHEvjtX/+
UasYIqy87UQ5bnWYK38HmEnCDARpmqTsv0XhXGHwNOUj1xW9YQ9m1NrzKBPiUrm8YmgprmAP0PKD
bowlYFQjmn9cCLWPidHnJ0LRlLYA5igemn4+HaKEmpUqnWIgbsBEvH2ekzUCrgndKXlR6vweAd0T
XqH40V4Qj5Q+9vQPrPg8fVq7vDad+5TXCnnjhetl1CPWo0bFQHfnm3IyehHsjL8/7DRRCSkYC3Z8
9nQgXDack9WqdnfSANJulw+ld5TXZLwASoLvSKGOYssz+4XO3piEGJt3A81VjF4GAPNNI2ggm4pS
xl3fEssPtE1JKV1L5Sc52K7hstP6qrPX9buZ3z3u/Lmb6OB04nJbaW9dDBIFZBV2nINLOXkNR58M
AWu7QmYsYPR/XRgLZ3bKhNLLGxdMcIshmzVi/xwTb7z0KhwhJB4IsU5gquyyvG2UnK0Sv5OLZagz
asHR4nwnT4+/mAJoNWzk1jLoSMIiZ8r3Abui4+cGj4BHo+656icNS/UO5RF6pNuWxnDWS3kShgZ6
UV3aXxrenSVljE09tRhn1eoEfKgayJyB/kor/b6cEGr1yH2u/zOSlIjY7DIKfITKsyz+rOIMNP7G
TTpbWzDB8+6U8TvhuZiHcaGrOwRYuIohBbKmLRbxflD0DOf/xHwBh60OSMavTIT9iEEvEIlCIY3o
2GuLbPklqVCZ8G9mWR9Y4Uz/nk+UzUk/t9EmxgddAjSPFwC0BVMDykz82webb6nM3k6HEUr8hB7C
T+Pakvf8VgL03W7ymLVpOzABShlwzRPMzo4E6w9AV0TXr/tYV+4BrrQxAZRcwVIs3nFSGhLItQVB
9Icy90hwhreHxnIe6n1tUp33pYl6xplQtxdc6e/ql20Puu4t1rb4VgPXXF+k+6M8DJuk5zEJ+rOS
W1QlsQZpMrutfk7KT6ANXvPciG87IGWYEsicok32zAPCgkna4rIK4hCznA4bia+4Yr6Q4E9ABuPp
1wBjvHn20KtkBu4lQCya17AegcnWqz6j0BeEsoWrs4Iz65uQU/ydXvcbkKIR8JCbqsxHXRemE7Jb
KlhFQ7FJipiglRZVsyEM4tS6+DL144lhd+Sa+I4T802wKymT8jb17upW5YnvQVoemP8Jr+ksZo/J
VFL7VuSWSRbmQv1P0ScQ4qimRN/H/fUmBE7pmb46HbPKT7Me4SeinA6mCnK+rmLcY5HNX1OpILNS
fNyInXVbstk+q1v8E3Fwg2keMHo8p2Z/s6Q/I8bGoJ1qxNeE4rv/gMZVxrC8KEWxKupJq2HMj4Zt
jEcFZjq3Ny59Nj7oRqhUjBnX0UbWh/2PkrQ2u+ACNK8oC5PGDhgZ1Zf7uqvRqF6fym9Kk4hBgapz
eK9aUD8Oq3TatTPmBwbidik3PS3QJ3piGPg1QOp44kLypDJJPzggpxr3TRzKnQOlZg3G/TvIwfxG
iPABcLgpyfuHE62UJBSyilQASH6/NRJOjT3zJ64emcfmzYuPCMtY3uHS5glxO42nOx8mMzb6Bc6H
XF5rZWhhZBrhgiKHUNuuCpolppfebWragINjYQ8IZQab+Q4pInlXGDOZJ64KlSIwtR/9dr8HuoNJ
0b40Chv89V7okURNY5rsDbILvepf5NtRNTtR6/yw4a2gtJ51PzvDDO2bxR2lbnntGw+Q8nM/EMiO
dbCsGAEuEwklkz5rm1HVTzGvsAtJKVoI5v7i98xq03LPRNniV2Odmgq1+/Nan+8c9dDryDKa4b0J
WCjDZl2I/kVF/4PkdCfhe6OqIiRfcQb0hb0wH3ggjyXZ7DVzwYPvygK/39IBNU6rs3sCGwtnxHZX
ISbcLGq67UDw59NQCpIZwUtmb0nBmSkvFeDrNKnSzzFjhDh3GtPNqjNbobMHwrCiEov07tuxjZ0T
7Vq/aEV9VZ5JqigHSeLhpjjA/j+cLCbVjiYWrhkgqkqOSAoNv37ijxh5szG5/ClBmLw7OQU8wb8E
DRWucZxh6QdQBcFW9OUK4/rhrqjPM7sT85YvJFTD8FU2ZSAUVNmkhV6fxcle7FXCBn5mT1Y0HApk
1Mi06M058/vHIh4b6U34+Wmnenjts1xqYdjRqoHIs/f5OtuOJ43QyELUCeyOk6wYlNF0mzFdTC3A
0nru8ZeMs0Xv/r4kITCab7AtXbQpom1xBfjJ2s3H0D0sUe54Z2I103g3DWJPcm+AEbj/6ZIAtts8
KX7vyCvR0FlDt/uEHyN1Cac5SO0VhECQWvLI9NR39dmCej3dK8tdV7xtNyS4hBbQENrWOjfantHz
ZcvMJnzR5SlpO3xjF9Su4SCB687w5VaNkpWXysyZzpXE1YNDCNibM6KeBMAbsWabLz+THSJOPLsw
BczJ5O3DOjPN5Y4L9vq9UySaOFLBvYuRpbE3HQV9IpvPr5JGLOSMwvHunuUnrSpjREv3SUEz2Nvy
O0bVHOxBY4ngHiQkJGbnb1U/FIme71n0DP/Sjg+FqJvSzLLqBLRZmyd0vu2k4jfNUAqvs3pY1d++
dMbb0c1nx+8W9w8zpreWr1AdPbNSpbTnIXKUM5Uqst0a4YDIz8PP1h4d87UA5Q8qCcjo9sHquWbU
4NJBIFE7BJAbW13gcJZkNzieCJrCBzYHlZC+ccEAiraJQ+NYl/AHU/4pUr1BA5XTpwpBQn+PfVjF
TiS+8rRQasoCXU54QMJtp/NUhhoUDryQf2FGgsWbsc3rQ0azHeiHujPnHTN8Ujs7IPzU1Lr288qO
LYcDFurf9QiRsFm2I/LH28IrhZn8a2DUgie7fWOJaeYbUIHHCrEXNbeDdkfAOM8KN2IDwtyNhzvt
E7VCE/JMFpKTJk5AGCROH9h0VdjETJRq7QYgbGPFmuKI8Pi5VdRRWFuaAnaM4+DViWrlMyulzulW
5IwJqiDIe2ulVauz1vbjlAe9a1aczHDnUzoUXYd5kh88NxdtdsGRBKulzbCAKUYHczKteVaaxszX
xFBTDXfQY6W719/YquR0OUSb3sPeeJDlkhezLZL+le08abDJn2Qkz+B+0N6U9lLlUEDp+iNtjpZb
R1y83+sE3mi3uYLP8d1jr/ytDjYI/GvEkSWTz25W3jmZZU8dTgsVB9+wttDxenPIgkGEo+u23Rb7
HTcvWjBzDlIHWdEzfvAV4+htkvTHW7T9Ce3YLXLRxn2irCMZ8x5jl7S7OSobFTWqNdSNyC4CsGQ7
fkkohXhkzS4og8ARMdkhv1GFBkZGUC1b9Xi68nfLuQzcr3P5fR/ypgtAjUHg92gJxPLUX7XqGg2d
p0a/7ZUUuEpe6rpwylBSTPIOaStnQamrGddFAN9hz7Np6z22Uep4eJyYaUKeZa9U/zlW1RUNu1TJ
2k7Lu+CsOYiXHwICHFP7j5O8Ol9ING12snJdkPg7+2Wdh4F6m39hOmRRF7HqlWNGKiqsVSuDO5uO
uVu0/1Ptf1g4vy0k0ITm/xGPX1WOAEsP7ibvUl1LP1vnhJSSKD8MIRDoldAM2AZ1w7IQ68SNe+Ez
3Iug/4gbGXgVg/R0kLQFi0eTai8263AJP2GjlHgS8SsD3l1r3k9gMz4QoAjWRAOiiS6v34+C5sI8
G6hDTzK8DEYpaezl1IS2YU95Zs+zGwNlDvSjW8U86ZZa3HH5Nx3kGT2hPd8U47+4/12NGHVa9f3t
aQE8oDHf0FqOhbAavJGyGS4dLNJaS9yHlbjtvM0snthvE2uf3u8kgZ+Bfxo6Gfek6umL9A5BytF2
Bs1344Lh3TRGpOh7GJgeWykBmEYitNVX6DfiN+OgtOgGr1tdmQe6Dw3JeBCjjTZGo1kC/tm1JEIl
nfcnCCY7E0zfRU6cuYNerhkclXhmLJUecpbHTQ21QI7i4T5/P0shak6DtYJ0Jqe1IhLqutGEM0xG
dbLTM+P0bdzN4FVXILrHwlKMn7DCEFvuIJyDo68byxQIif1WEEYz9gxmdJHL6gueEe5CLIgAo1X+
90j7jaR3n/AVmvIt2reBiDmTPWmWMaO16F6HjkNug1KizBPbAryDlvfuoaGKlEEMsFGyrvoawIVH
u866Hz4EzVb4mMi0pe3FlAcN3+s7T6yQe98tz0XqzaF42Ey3w/iaCXP+iK9rcCe42EbeCJu+S9um
Yho3ECEIMpyLx8vVe3H3q4mOzlofmxycqio1HmGF6a2lwxVJ8jE2Yad2Ulx7WeM1VhLvNsSMAca9
esoDzEwqcPAgDg9K/Mu3Vv4GE9qsJOG4/RjQ+Z5JKJBYp8WCTSX9HGmq90FVJhKFzwaJRA0OVZY/
4aJd5J+6UEPqWXpkRyhWePood6FNJoas1cKJmOTEdP5W/KkprA5WXeRY4BJUHEPvt1WEdmjiQD66
3l1h7Vj+OgeB/CzsVF5z1tiNpSizPe5yflVG/fVP/zkfOJhLgCjUQtsa4fU9rV1WwctyXxEQFZMR
cXbtRQf0GFq0jfX67jLzCvVuDs3nTmFRQwmfhkxDqGrbkjyeJ+vpuDnwcbDnZvTpK/2Jo7wIsG4z
e3ESLUuRiKIfUtkvPL9b877N8rrEiWTbaMzbAu2/INTxpz2sWSGoUwJudk6OmIdVuQ2iQIe/zMSm
1uqAH+w4UXeBSdlptU/B2WdpJ8cJQBqL7+PNfeCMvm3AKfHKQXSNcWNlV4jSS5uaB8eOJxDNjpt4
y9jgBGDRtlpiaSMAy4bcmfCBrjVNNW5tznw/Mk8lzfZVs8EaYndCyqkPHdBiey5D8m2VKppUARCa
7ULO+S7AJ/m2aYuuEDi7REBtV2vUOXgv46+lFfjjuZC/eHCiEtdaBpL/46p2SRyfceaPX76OeH9C
7d44QXiVLw9MZm4zqj/JOTZhw58nJ0eTyH6iE9XU+kuxbBxqczaanFmoKI/8Jk0NxoEFrKUWPrst
TFi39LWNMtyL5KZkUryWWOKbAAwuZr5NVas0Bk5vBI2fu6F+NF9zAB3dMzXB9oWYXjb+8Sky6lXk
xDgiy5pm+/f9ThIkfmwA9Ci7ETwR83TgO7lkUP+BcdUC+D4sRIqr/RBgmeuboMC1IjcPhini4XSz
kbC2pPoOrIdl15wv00a/ZxQEMoV7XpqopRGtyTBb+RCvv+09YzEaV0vbZHtoglpe3yewzxtvza2I
b1xiSYcNpTbVL3X71T5moTgQC8BuKO+BG4+iDgbObUJJa94+mbxkTzz8x53enDIO2bFsLKHkV1Ky
fhiAmGspEzf3KoxEVCpCtp+DkJIyqwM4zwUn8TvoAfW1ggm5u7sy/oAF3LnAKFGFZf97BRgjEiJy
jb1T5vTPaAgCq7dnqxdXojvqhAhey4pHtrVc1wb76tyqakzpS9+Z8FLxTmEfrgdZiPGx9beyQXIu
flmqD7KqCtBynnZjzWhNBK5K7wwqXjGzQT6XAFXPVOC09/3mWqVWLK5lCDz9McbvzwRnE57sWPwC
saY1DTtdWccqd+YLExJ8GSNlAKhEk+ka1ijONvEif9WEMWgYTmIQABMaUnndJYBB0/yE4jqGMZw7
Sa5dbNBm+sg7rAnAVlvIZ3oF3YP6fB1PthM5XqC4GKKLxZwCEDutpORx1r8w8Cg5hMFo4WA5jNe8
MmjjY4WK2bIOEOFRh2kfFaR7+4bYKDFd260BqdxyvPEduT+fqFEiru0TQ4qCmXQF/XCvuT0bAI6x
nj+KqldEkpLEHYFrRRwrXzAP4Q1JPQ7NnNcROeZgpxNHS4OECiB/0MAtuHupIyXkTlkoVId5OQYO
dLVu+mVGdQRSz2qWF7HqyygEMELl1AGnp7f71SqppXfUpsLq36L8AQ6DUjDPvMOlgxg+XD7ZEtC6
lKN0w73D+syELvVWtbmwjz5crkdHClX2bW4gk2mPoFLx13QtSt2hMEvRMc5FrGHmLa6UUXfjKi4F
eoKWT6uOyg0qltxLKVbzUR6pakUw9vfsf2IG7Af7uEsGJ7+zfNT6XlSqe3GS61LE82q2FUBjt9yB
YUvIrIxoNeKt89CXid0zxcW0bTMZwz9OQSajCGlh8KTfTAGdgUfOsQi+VLpJb7JWIOLdtVWZwtnf
jPZza6dcKmTa1QxaHSL1I4n3GNqvbgZT1vyu/Ajgs/zgVEt+GqKfpVltaB9eydnR+oHBV0VhZZyj
21ZWqdnMIvjf0k0FjKpIbMKswOu/sxddeMBdyzIOxhiWu9U/OBUujnuJMju3el217+rBSHJhma+D
6g5DghWEhJnQR/WXM/KpxNf+04ZgMV8ORRtgDm5yyFVgKIy33/4j3Th3aEuPcOsFjhpy8TtlZTMy
nWF/sdOExMqjbuB1re52eyCq7NocNZQD4mzUcHmwsXus13aDLOxrmTNc9c5S05RtfFbgF64/p0hn
O8R54h6K9CIEgau9o5mhDS8U2XAlrlTLJGTmuj9AZ6iqpppAx7oSZD5pi1XrJjnN/sre+BOHMWaY
2H9H0A8yT1Dl0MZDJm45FcMnKhRd+ylaQjwgkfDLqvbd+R0vFQl2Hyb4yq6NhhTdr5eg6zVhYGEq
I9mSb0fNxeV+SKskPMnUuRxxnWlqRAI6LwiL38HRLpR4y4X7CT7s3tGJf/4HCcwxDYz+1wDJudEX
CQUKf+FA6pn4Mm1cbrwczSCjRg7nDTkhpea/XLobni0YHU4A0j5TqbPQbdKfccOb4NvO6uwNhHJR
x/oYFgcVjJL9tD4FYjWl6pDQPDxpJ2kbCngLYZhjK4qiDDnFFBM+T6JpHh91M2MGlCNDvQopoUIc
TCdNzUC/4+jJ8+3fWDZJqFa6CWNLaxvAWBrOV2kEmjs0nokCsm6NNl8Jdw3i05IHmovWUvStWu7B
fOFnHXj4X5IP510Q50HA0CBeO7beruw40Agj8ccYAJy9MmYtK3xQbjTpEsiMUQvL/lxTgIeuAIgb
f/v1aau9h+T7wje6FKpeATiwFTwBG5sSjfuy7PwipSGKkVgr9U+/wIAyNH1vZNXL+SgBIikSlLFq
7cgLZQhtaPTZAJjEw3XicFKUSA3egZfQosAtgRW/Kecm81pFaSJuppCOuAv6vr22YMaqan6tZO2R
QKUqLIl49EjaT1HdUPfBTSaLw9Hu6bfUDV3/Zg9pBxac8nkRk0A5k4GHa0qBRwJHxg73Jr35bU6/
r0ABFxTR3LVvmNqeAcR8mx5IBvLm1ZldG5zlE/2sWufEhN2vg7tUlxRPQdpiSUXEZjx5ZBMn1QPO
Fneeh7J5MFU4ZMsuvM+rwSYGFz2ekhcSAVf6bjqgilsHatm5Drtst8FTCawmqsGdNN2doUxC8l6l
c/+E6t6iclEAihFJ1208vHhL7wkrMMQBpqXcqEvs75rDJnisJQRbJ8Kp0aVXe442PHVoq3mekpPQ
N+XUgUdezmtT37vScKnl9WYJwQHaQi+ea8o1+yJlSVeQxLGl42cm7/lkHkARzXHwzykzVvJhV8KX
W7USV4BzwgoqtLNYfirTD3xSzNqgzH78smovgQuuFVYHsqtyxiY3f/6ERxaVxN6n6lJyNh4sH+tq
h2ljNvrWwT/JuZQ7lwbDXmednxpnmopRsTVG412S8MLe3LJ0G+AeF60boe5Gyw2N32uPmzNvdS2o
WTWG7mvNwrVToxeHkOO45LdNSXaIIl4wTSR560jwE+f8hD52QTC6/5uUlfPCUwRdDXnHBPsflBgF
KEC+5zpvowl9gozoF4i/qpiTzI+z5nbofl+F+HkzEkewq5Ssl1ATEUY+8ZgFxBKeXCg9Sjcqa9+6
4CMbuxrQFoFIubq/Ht7PeuiDtIuyOatdaW1MZL0Xcxn759ul0XAJYuEm446fsRP1sdalgVMccMMG
wXCzqIFntNCm+yv8uuZ3mHdbqXzdua9yjUlBZPi+WIXab87ueAl49jUIeJMBsYAmu+jLrpMQE9Zr
9i+vMDjQzdd/r0kGQPlZkabrAA0yElXSg6JXRIU/z2CFpEmUwRl76Ft7zbKMDd14v5wFqjY6Kg05
9XVZapKiOF8FkkifmsHlyEt9Qg5cDxuKMAcZBAl1Lc6nZcTZ1ppvPBhjmGnGZiK9zcPc9ujROX76
vfLN0XwFkEvBDernphTJsoNq3pb+87Bx3TPN3xHeQCQrC/iem7dswrvBc3k5xJRWtkBmqdfQTF1l
6z1Xpgq6Otvfd3K1AF9boSe9xybDNZ+AvhSzKyqwu4h/Yk/UJuUlDgfQwkNwc74HAMO6CejVkDOL
PhieTWjofR5fjqAEt9TjE3X/QupdYfvGwwl4FsT0A0aFywf3rUGleC7Xh0THnbBLYAw78PAs3GsV
zeTxYpSufHGN6cQL6IbjFnNq/Ufef4v9u06P6t+ZFyGN9P5LaZZgxMEGbAOKYOg7uTfeUZ5Y+rap
6SiDwj3iYdzfkDyZowT1ei7TPDLuprtZc9K0AnYolMhlOzbnJnJ4Igu66HbSeJcZcGSpEZCE2lj7
gA3uciPGhHYB+jFn0VSAPcwELc6A4lEPnun4btnJnlxrnqZgFzZMugMy6H8xOHBv2WjC94VaepGn
dO/+aNniEKFfSeHV/hJRLnw/cKaAAKst67wksnxY8SjYb8bB4tjNch7kfmyYRFW78tSrruNUQ+xK
fJ3ZmP2kmI+ykMdMvjAA//ASylzhnX9qdrlBTDLg/Zebevg+/8p5Gt+IKssiuUZOvUlK1iVfJ85z
sDv+A1QfqZ+C/5plkgXmdj2jhMEIl/zFs6BjDrTy6kfRdJoEgHxLS0ayDLiVatl4cSBrDYPs4B3K
RZVh8pI/iPyrOcDqio76cbpcrBwcH6Y867BxFCnPguwr0pzzbEMlhcYuU2wNQ+AbBX5BYt6TeUJP
6ISUeHqStg25spDTNqZJv355mohVVhy0gEJ9GKJ/0p4AbbcracmPm2n6CwWZblIow/w0k4KAvl2z
V+nnrBCRQ4E3qzxUKF5GPwsT8kj72huVtPEU3uk81w4MwZDyWKG/l692/c+b73SM4t/QWisGa5js
mt9Np3fEUdq6i8mvGhcGrqoBQU5GgVsISKlVUm6nImG6WHgxcxaqjBLpgPj/ihc10S/UJffnmFUT
Tswmz1QN0l99GyvkQKuNBtDyPnLcq9Jif2ODQa0N7npJt8/Mh1v/k9P8/eWPqUDomBtFZn6hfuKg
NLTf+dSY4lz/rkKr2Pzb6o/LOh2d6BAQJvnDRe0Spg7k5WbBRV68aEYhHEx4xT56aItc2s3NRY4f
pb7ZQgMOI/1AFjAbRTLUR5SXuwpoTkD6OyeIziqBcB0ot1uMPBJgIgClxmRfBff4pw1/MpqAAwHE
fibQmnFDRNk4l1Slk7soFhri5bHkYmcY/egcbNoLlDgQ0v7Opz1h1O1TFqD6rUIJQdydrtzqOGm6
ebz6iAATRrWl8q/2czqkXj7Xw3t3JMEd6ZDM4BJy+DxHGzlhUL4Bc4Vdses0HX9D2nFrDIYb2Y3G
ErKRZjEf1Tby7Zw7VaNM6t7Jh9cytCE08s8yN5dvwIN2R0K1Ah0xn895cQZE8NaJTKLi2vtMXFiu
M4hfZ6/F0RNmCj4ixPraKNmgd8GHJfHb+rsoqgz4FCy/pCbqapq8cBXRaR03FV3FOzxWQoHMJ+Qj
CsdOQDztLhrYPxK6mIt9TFDjlcfQeGNALS7aOT2jFBBAGwHdnzmrvdpx5eO5B46Ufq+QwkDhcdxy
9CyRn2/QfjkVpTg+82J4A1Dhq2sHTonTzDGjoJXiTuEHhWnUOSN91jSOUzO0Mwl6gB9WsRT9Q63N
5a3Wk43NpNWd/aCZVxKHrx8hOAh9iZRUQBbb4DTBSCTXZCuV0WfhjRy0Itx4lfEOtFR1toGbpy7U
kbpZl7Tg0fKLFxGizEoGEqacxAkODBKgmgNqc/gyE2RpbPBk/yeOhXGbhX4GwUWh4u7n3e3muoJL
ModN1zmNWbJYR0+br6QxLWntpPx+mGlr8XDtWg58qDz3F2vQhizv80oyvIbHkf25yiktmGHDsmig
mvS2VmGc5B1x4UlEuQdRNhUaYFQKrV4D4MN/wqliMm4biS8lgGqp9TdYAKzcPVzHeRInR//3GH8n
V1paYpaZksp+lElJ8Z805Fp61im4jzRiyffjCxa8of6kAfOUcFJdwxpV95kVM3KSlGU2yDmWeySX
aYfTvXA5El1rhaOVEkh+BKXsiydBle9F8CNCYrwNcIn62QSbhk8a4dw9Su3qG1GZYuVCB8HDq0Oq
/g1dUKwDblL1HiUulkvi30nFMeUW+tiZsEPj5Z3kEgWT1R9G1vxWOcqfyM61jIpdgDXhAGpa3BmE
HlCLuD0e8rbg7tuCxYrrosetrE/8rXWntwbzNpAiYX5oh6xR0Noqjk3KhdkXF/aCH2GHNToFCZRo
Fp1sqM0suZSVPiTe9BHVqnvkyjF+5ScLo0mVqTBj7hTTCO4p1pV1yYL27Go7dxXCcBjANhOxlPhL
UGvAYlOUVUi3GlBDKFLiD+mwgREByKIIJnWKcLsGrDg0YIZ2X3IBy2aE/Za/h4YA99a5sejIYbQr
WoDWDy1ISr29vQT+GiSvWU0UKRfM1V2/um0delTYvesnvLUQlKXqLJlLgvsRkSwyllrCME2r1Ed0
IRITuBgJTpfjyxX9KvN7ybso29m8xZUFiMojwD9z7X9gSPw1zUUQHXtj0Qdn2PDt8XfUzIq6IVhO
c/5Zwdfvg5zpBtcFoqSWI0dTeHrnzrZHDEiobExUIgrLAIHai4s9tE3vQBjdKksOz9BVnDtpdueG
zeJTOajmILrXza/rnShucrP7rVd2sdu5dQ6GeQ1eojpMWS4rkE6tLzfvzwfoyzlllFCXt/Eev8k7
JrNFCCquZXKlDuRmqVE0uv4A0QTyWaN6j6soJoJTD2/0MW1Cwsph9URJgxp8U8ORArjy2VXWzy+F
ovN3mL712Cidf6uwxtNfOce28YBMyomwVm9NX08D1K8PlQmOyrihFJM044PklRpoHygaOdcb0sK5
wq+6hjTn5y0hSBMC1K0PhFxCyhcn80MeW5gkCNdAqL5Cqo3AuUbHaO9QH4Hkz8GoXxB/Vsu6ulXK
4S/m6eZOCRNASk3N2bLYJtewPG/BMog0RRHuyCcUP8e59ZZ+MCCUK82QwZR4zRaH9zT9unSxaMnK
kphqNnOgRUGK1YGmjqAqdw/MraOnOXc/o9HfWsf9chJIF3hFoj31PPj0CfUj6wgtlerEuJ5YsPj1
ludq6pckiemFyUMr2aJmxn/otPY1TrJizhjV1idGigfMPSneMapSbtbajKRp4vQO1hD5EyMIGFLQ
oMPRDIdg3BLXhdqVNRvXaYwxE40E72k88QzEZ1ofHD/+bxoidMFZVUhWCvISKTo38pDosP8QOUOT
kvdyFvpNvipRjv8H7H/lPZDn1vUF/wGPZYptUxz6dVIe7haMgxqugDTfNC96F6UdsDdVX0amsTp+
h1mFoSLi5vgnEi1GXBAKx/bJKQ/YyNG8l2aUKKi1B4baaDE/FtLRdEExIxtpTX9dNiZhMjrnqoLg
//l79XvWMoEEdOCFv0oYxqtJDyNXclCoxjSrwpTosQbx6oZvTtsEF82fwj+5lpBDXQuW0LoykjmD
bjC8o8WGuJpTkopWUBxnNo7Kyn/T/TbB43IAn0JB1L/KRsCow0aR7F6LCwln8j3I2jeKchuDALKY
3Q10Sb160Cc6iivnP1z22FC0arMy2fw/i9HPjbGCKOobm+r2Vqna3dLq0egBrfpBMm8+RRdE/L+l
OVuQ7sLnQNzqwj5xai7OYr1QFBpuOfo9Syjxi17utMSLKgu94IOAvbncV+wBf4sQ+VWMP8pO+CI3
E/S+FNZler60T3ICBgikJuw34EyBITD9MjwWT4CkTCIzXr0xejxxetujnYmmf/AEVpGA3XgpD/5u
cIiSYWuUhuvGW6mc9e+Bj1ekkMj8y+wcvB0lTndslIQxzRXIq+GBo+t3NfgfQFafTwas43iDrqDv
KfdRe5AXPX54C+wJ0mAfH204IeRRJy9gDdSe9nGmsTKJ3pCiyFZ4b1Fm0dq+8uP9FLE0v5tDgr5q
s8EgBMKMDKwMRgts8qeOxvlMib7KRuSftPSE8mjd6WeRvEEnBHOIB/1ko1NjZykcLd1oKlA9sA1o
UFH0DdHZnhw+KeFuyVlfB4DKHSERHBZQ3ZoTjA6iKy3wYh/1L81YTUGm/pHuBQgKdgcQmeUIw/9/
VNy4RiM748R2NcAQM72YaHTpMulz3w/Pjodd3Mit4M0g5OPRmp5B2vvaTp2qdYn8x7avnxznpoYQ
g2BUXQjdTt6X5cpPrSe7IRhAGsrAhg9gkO9AH6JMvSUPIXppcCpxMx8HLPDZwOorL3mPlXmG8cJs
K4DftdG5QeYcUjS1jmmdF3l8ChJFgnLXQ21a7+Xfxl1PauwpcHDkNp40yAh05FPStn+AxiAq/3+e
fnn6FHR+PxuUGRFgYK0hO6GAVu3o/meATPYyuDEhTQGob3Wajk0Q1YvF9eE3Gg1S9s5k7Ejo4+qs
SKitMRM01Qp22GLbOHmeQUIwETy4D+3XjmZJT8VvECxOmKGhJiofpPo90VucUOjIJr3cS4gveJGV
35dCCIpdm6Wo8GZPvTlRmF4hZil+LqhIYveoj5GFu34Igobve0YmwxVnpowyoNmk42AzMsxZHs+A
If3OXakmZeOPzU8KWPY1/hLHx1sgPxOb/5MYIGlXK7rapYc//mXcfqqBNODkiVqFwrVRYKSUm4vQ
NZKLXUg6s97aYHobfKmdACCNSu7KqqOflXpR1drWno1GH8AIdqk7d7ngCLNTpcQj4n1NlIal5iTt
amskb0LCDtOlwwp4i7c5QN3g+GK/ggvBZwelGlT33qhUUiFVenoXWrr8Vm8/1GDJc9rewEjYpTVL
K+vVMKV1lBC9BpApwH3g9/FdmZueNAtxBp3sO4asT8gg4RVPco9836G1GRbe6Jc4RjFqFQ0w0O2U
RiQy3AGq6+INf+1UzlKHyWjjS0sn4rIT7p+kE6QoQhOl+spZMpC+w2qFmyIv+Ql/zklQZboWyyl9
qcUapKDnc8ZyOOXcEMuK/hiGeyfhHOexAdDXpYpKWAZ2vr6jKf8VuOScnmykp00iPy7rAgxY7Yi3
9lIbJ+K6avmg+ck1uGQNnmys8AWKKsXeArn4VnbgYE5Gzmn2asdChPKWp7qzygR+xQj1TD4RfNYV
40dVi7Q1NAb31BHiq/SkeqPQ7RoiNAkX8hd7yLBf73C1H/UDdfqWErFd1xHNAVt8ix7z+AH+qt0T
NwkiTRbO08uuD5T++DlrL/z9i6Ht+hWH2gWVkRMXOKsvO+VTJhzRb6EtchR0XZOEHTUSiDao7na/
1zt+5DUrS6nR0+pa+kHCerSuPIihWSCCZi4C24dGvAl1FZPgo1Ve5UkPZFvlKgQv1iU9k0ptkP+L
mTZk3Hj+R7Ggx0qkFZdxoFBpjWITz2n5xWAYGG0P47v7g0WmTTGs/3mqK1tt4fiC6b0m6dtJJVmt
aKr1/Fb2X3rO8PFeFEGQaZX7b8RU1Q8o8qeztLyefqIPBtA8ry+jR/QPZoBad8ek9MtVkqeEVNuH
H7m+eSrqOKChpREpFkO6Q89FR41BLrDMWAx3k+28jSLe2DfjOm0ib+f8tv+S0RGD4og3ziN0/Igy
aU1SPG+Jqjy6SZT0WcQdiZ5u8fXLwsYsgC2AI4iTvh7sPJ70CaZ6KbTYg6vj6ZdAqIElQKIGQvbv
ZBZoiHXymPRIVBadQfFeEL/Vo7Rw3d1zWDJiGXPqTO9rgG+xhOieqOSBgmcW4s5KVNcA4FJi4zC7
TJVEsTWf8/XnywdFvwgcTftjuhGxqTq3oXxbyaAeyAFRUn0trowIEN+BSCKahM1JTJ4OnVcxsQzs
U96e0EmwKl0k5U7C9/Tyji4zRLgoftHreot6LrjzYOgaqzqVc+C4gHesR0XNc+Y9f5X5VDcfZUkv
rTbeqvK9MCy/FKXG25kdkDrw56WuQS9zCed+7AfPsKJI0cRFrdSZXxXFMgc59lfrUNs6Bg/RliB+
2bdR2/fR9yPfdO+ZnmZdKsSMxaPexaLqezX+QgjFs+dgdyftzq3x1t35yDkfdOlbbcao+mx52tZt
++31aZvrrz9gua/sbTWeQVUUOSz/AqrxTHlYLCqGYxeuhpNmNklJKrwdqVPUuyizlgOC8IWNjnI7
pt8DZO5PDpAEy8u2GS8MtAQUCfQqsON+gQ66hpj8L69nXqxtd8yUnC/E+bHDH9G6J9bMnZ1D/eQH
m7fqLqayBalSXuv/woKwmuDZlu2hL4NyxS7b+etRLage/9rfxf8Y/2RxVWThJZ7TlT4XdKq1O2AS
3VbTUSrVDeS2eZ0NKVTbTTMDj/YiRfRNoKs4KrKbowL9wa14viNjol6l3+PymLoI9f3GBOaV0bUp
8EAyGsyz3v1BwC0Z/e8BkqoDQQNt/tjwTiqM+kgsQ1WSTsLJC8eRuczaaaCiEUZj+46+jrILiQhm
cFkdBHYeouWd3bQEvDaNoKIjcOt3ajinvmTxonSQ0DOf0FG1IZyWRzNz1LPh5tE0M4X+BpmrxHHn
FOOKlMfQEifedCdqnE2YDG3O/7t4FS/NYJd39Q9SffmA070htJWjtvjWtdMw1jX2BC49gZKlZ65H
p9f25Y0xT1K1T4rRU/UIUgdtA2vhjZMmOy/+7naYK3O4YPm6ZovFS+bKddVP1p/BQL9OVJkiGlrW
4TZHwHehrnrD+atXTQ8AuVhWOg2deR0ARujRBStwTr154ZF5u10KM3ilaBOBQOTo4LwEJ8NlRoE8
5dLt5OVW9hVIsaaa2C9UYtGvYGRYkDx3S1w4CkjxaZryTCspruxr0oVDLR9p9/RjYlwMgXem78bZ
XqkOk6dV/AW1R9MWWFhkNhdupsRr7WZwWMQtm0LM6ak+tlYuFcoQBxk4WcXIO7grmh+gXkFSKRyX
bhuVTfF3pw9z8VBxBexqtwV/nsFm7++FNlZqaSIpp7klIY7Kf6K02DnNV5SV9IGPVFUgqoeEb/9N
2r6dBCgeD+WtJDYuZyRe/cE9lw8u4tqCamOcNtRbdj7nG0ypaHfwZeHw4excTZTEwaqyk7Zz2T/M
wyvQsUKGtGD9wOqCq1jP4iM4GbdNiKpwWPXFf6V1luzlPKiC4V/3bB6Ye0EGq88TJaFn7rn7FaK0
lE7b/EHoSUdCvdpt+a0pp0vvLrGpXudRggvCJW/ujSQsnlj24E/iR6bkO8HjERiS1lv9mMEbMSNT
lh0XSCFH5ATZLMEfWPzrdAO7qUWq2NwT7iJ+mdjLLw2f1qL0bMOqNUfSC6bJPCNCYGNNK1jV6rPh
tlTE4PgRsQQb3RiNf8NNWVJPKhJit4L3u8DTbiCDocj/NUN+K+pl/cF9bi3Aglmg+WUTz3RFGGdm
sEIQTUUFSx/u40Fn3HKOKRcHbNOLLWLj+G8UAw7vcWnDqnuMPO3QKWioGb02U536SYqFW02Zxo4E
GSzkuwRsKPodUMq+kPyHrbvjciAI6Vs/gOS0yZj1fFiE+sQtg75GLrpIqTIkvrxesEsPZxxjmHoF
ueV1ZBjQJrgR+mm0NAMTFjZTRRp+P+Fg5tlxwglxuIstXDCePI1MuThi4qvdJVMAy73aVngz8HDX
bLO0rEkwu9kaAjibLXwwSnThkgO6MuUFSAXPKJXKP97MwzoZGYGn4FE4Skfaq0x5RmFCotlmc4FR
nSS9QBWTWVWqbm2A/UoBFTZynth9mL/saUXt5XRDBasM8ACgdt9RLE3sj4H5OEE3ePHcrbnSBDrf
upt9fTvcsa1bUgQfCFI8pBkUBR1O0kd1MAok3xKwlQm4BAnhWOyKnu+ueZ+Edo4cyxNJhsn2hScF
IR8NbjUBrunkPmPYhLLjqkaT/GRO+39cZHayIjTQMtnaYwZGUYSc4VDHe3PtVm/UP4DzbM+T33Tn
S/yeLnuEbh98wtDCdqz+ELr6T4fz17Am8S/yyB2C3gNOjvX/X73XoBiXe6fuWmeVUBcGqp5tPRSi
5AKnsPO9SdO73rmBfNTglKaVxoMZeTGa72SOn59ZSRZ2V/pPW0HEUvmkGN0W6ej6aOgdP2rzztZv
bDsqFLCkIKD0yhNvx/+TVwWF2JLHItYOI1RWHHf1yaOCzsyowmrDQTkIS4YZPrRC7Rr3a3fa5ndF
HXjheNhR5XPWnj4D8qOju31rSLr5v4ef1venkOyNU3y/F9Yl/l6mvxPcFnO/s6a8HPio7q4E7XMV
tiUmkOWzm5oERd3LZuwnvX5bxOw6QAA4zlB6qktFnFw2LujVxdKYLrCgR5+MPNVo8h+Cs8q/jeqc
bZQyrEC+rXpgOLkwADxYcsbOHYlRjR7Yv1vvrjtd/lMOLml2XF9AkGgryhQ10XO3gxpIyp3P+qHm
AFO1jwu84uNuqZpBlJc6ZsjXLCGG0qsDqaua+E3s26Q/FeBioqO9pBkfYomb/PROxkQT5nDgWgYI
B9SYBI0rV/BGyTh7fw8rFdo0EC4Wai/fv/URkq+7xgDtKv0k9v2oJhyXuGJkIqvLL68rdP2UyO4B
egaIIpgBZQAXa+cjt90dGZxT7vO7YWUlSgwH5WVeIMmD2/Xr7JjBL+i0gkmxikfl30MXgPOzwW2d
KeaMe/cvzmsqhMf4FJ+xu0+kfqJILaY7JfPLZ9a3FQkSrNAIvuySDHWO8dXlDD83adTApNfAJrtN
KVPbEjKxfiFFYzLCoZ4P9hOi7XTEdj6Jg2qrVHWJJizGejDVyBXOCJrornD+W0iCWUbQYV/CRgMm
ZwjgaockW+pRW92IlwUZVEaeVZGpBtx3mSIuRrOptrhvsTynRX0sMZf4qfI/3FZM+m8QaBiiFHwO
Tznp0wB2xB/yDaKd52HPp7cs/fLM2XzhEUAWIMy28DP3bBvfycHx0YmQsTOZOmV9NgpDOH+KXd5A
B/lsHn9Tt2YV4rVd3Wavfob2x+BUJn9NkT6DcLXWGywhEpvCMKqKZTC/QX2B/1OV5hlIXYrRUhJj
C4S/M2IoyGdo74U3ksegkAv6M96pxv+WlL24jkqND4ZLkzq1NB/CXIch+sSp8uC8aq5/HSpyODxW
M1nOWJdDbJiA94UPpRxdyznidJ+5dGJQ8899Vg6d0NgbsPxQgDhrxvvl2maSwTG1O4VE6erLEhmU
4p4Y0Neg9qfFwz/mgEIe7DQWUKeeyIJDjHWCvl2uyFCXPD5O+U4wGzaowS3gKas2uNVH+uhhrcIw
3iD7S6Y3sP+CF5JoNI6lBMFL+RN7sZcJZmLUYCJeCluc4J++izNTHQRENGj9jR7XL7fGUGIU7sRj
IpHO+ZV5nn1citGxuuc7SGUsRWJr6EV1QvE/YC890W8dcmV2Ub4ErBD+GhnHufTGGirpu6P2D4Zd
qyQ7PaK54i8BGKR74nnwxOPsbDDljQz+yfWjHziNlBVR2ptUepjggZ7FaFo36CuR0ZKVjUqqtwQj
9eY6FmjntILkUxojKVHrT41N41JaGvy2kx6PMUHQSHUhGAaSv493JXINRIoqrO7xUOq8ZYO1bBnG
SjBV309bQsM0E6V/CW/hWxasxg77uv9cvBBMTix/966mAlr1qmczmw+JZrqOjbqoJdIgB4qrVzB2
RwCK6Y5T0cLnZ/WuCC4E6T+R0lonwU9ds452CONYLq1hgzGGty3a9PhM+cHYAfC10EdQg7FlyuLR
CBcd6wHRBA/quAtZdbkzGnL65fpCZpbNUfuDuoauoAoAwNHrOgnK/6DLje43T6zpccPJPJ17QN4U
VVMQmkowcK42HZ8kPzGUdqGKA1QouctY3H0wuS1szn7Z+WghssjGvV9ELIrP7evLElMdkBLxL1BY
xkhOzCGtz0aFBhRuSSsyoQyV+sACyyWQYmkop/KMCskntsyDfWR09u351Jj0ikVcBNOESW6e9HMp
AKsxp5zo1TnimiIKPDd1FN6gXSg8DthDTrPJe7L4nYf+Yas5GIRr4xf2CtEMWggsLcl2fzsPZM/A
iBAwiLmR5XP+l4aGnPmNTsow1urhYV8h4CPOFs+kk3zLC6fboYKIGSMdyCm3Ya7I5W+zDG+CfY1W
ogBxILD+TMcl5gq+UexRpciP2nNCyrGHyRxUCdCw+JGfetTQRVsoLuJIMhl7zqUyiVIPDLoUtACV
JJzXMrS74qbyVnwYHiF5sXBKelASfSe7htZ06WLN+SSmXi8snXcHsXXYPsgsnItlgLVkLjv4lCjW
tv1V3jzksILaL7WeOey9NTr5Wjr3mZydo2igu9hywtk8kUzMHnwvD/9MAqyHZQgyxTy9oimDrXwY
gKOqy9yUt2MpLp/WavyVbpJ3YboEjxH7V6xDPbH8hdIWsm1i/ItH57s1/cTYc98UkzuC5009QTOU
xYaFtf1xtOVVdoH5ECU/lLFgS+m0nNR/3RCMA1nQ2oCA2MQYOD9RTKIt/0f7s0Csxns5IWOkHjcO
sO5ywL6nk5H2pogUrk1h6RBqWsW8C/h2SWQx5sH1xpEDtTnGRc85VM5TfEP9gWG/ziolEskXIkQY
wKIxVVnZ7pzPvxIs0y/wVonMfVptnn2r17/JAeF1wkFYHpBeCdwOAyI/Z3gy2pqINAgMWtfN6c1v
YFKeLxYrppunMdPOC0S1J6mRCMVMkirX6ekXUMSG+KG06P/h1hfDnBs9AW+hzuhqz8++5uoUlqyQ
n+kPbYxINpgfsDIe4mHXU/kefjEvQhUa4lH/pZIDyHBR0/E/33z1E/33WXLqSN+3pfQuliadXbe+
Y5jFaCRB8Lz+iUU1imICbcGtJSLZXRlD1/OZj55owMt2fzeo5vhgK8T9b+Wq3CwBA+BGop4qk4bI
efCI0xDJ6uIM+4a6UnSficZi9qR6xbsnzM9HHwuEYRP0drHjWwrBjs06C53wrv4NNmsa8hyHlC4D
gNDakf1lJSsKfzorAjQHEqr+GoFPrf02LSQPZPj8+zlMZlenoCn91fz1VK8UAMX8SCHPXPQ5YWgW
F9FuLUKBRFnBXy7RHq0KoLfs8TSq8ymVG5LpEtrUX64IW0gNrJYpSbja3CE+OjLVpFObw3th09qS
h3Nx5eFNSDsZTRffKRYHXaKuC5WUWT5tsilTVegIoruEqO3jVJR9H2Mj/XGeO9ViPmPd33GfAvd7
WIN2H1P7UbCw4xHsN84L0Gi5ySypl55FyMCWktqdjPmD5JF8Th6CKNE6hAkkliSoc3XZ2g/exu1H
GAAc4iXwKChJIMo0bbVNd+hVLhV2WHzFn5rtcBgEWLsXHGFTkYS3yPD6JAMFX9P+erMA6aYS21RE
98e/8tDn9WRRwhB2Bxy2WeCQDmMvMKv0yGQKr8i31Mq34S+Y1n39UhT0mG8+I/p5wzK4o+zJ/hwE
+5x1NuiMDkPxgfRPQy5Kw3UiQwZrAbh1z+k4U4hx2XRV7mrSCZMHGzCavl+Er3aVJq5iqNeAnHFk
iQNtr7v/qNfZ/E2QyVyh7jEQ6YEN1uNVUCC7mukezmzgC9UAwBumPnM1TAG3crWwop0LMjdbjPnI
v7eOLwRHxWFwhMDvR3dEiskfM9KpVdG9DwDYN+DEj5wUYcBJvKgQZGdl8xJ+e1U9at2WL3ohgakB
e7LVNam5bgyubt1KVyA9lBr0r/tMIcc7/AgLkhbS6R55yu2n+nQILtD/QVGodONbAFewILQz3PQY
P4FaEH5OJ31xsxFurIKtUoDjFjrKcl3xHjTBHEax0aqSSHnSAUp8CLT9BwscfqHuaqyaH1Z9GJD2
b4+pN7MmyeFMp0EqtoXQQnIhjL/XIaUlE0M9KvtVbwLUO5pgGEpju7TiylyG4SFUYJNAdW8RRQ1v
jSHN7yyOjbYVzDh9sK2tiQosLYjM/go5tr7NEYnXFGxsA4NFrdpLONkFj3wa49s2lcVb/ASryPEm
1nGaUXhKNmt5YxkFfE+qwxSjMcEq6HBaVOO0xOwhO9ywu713+vKUnvadx58Pf5KoIykyoRczMjNa
tDYN0o3ONs8QptVNUMKhhF+dMTozZMmP5dt2bfGGjnyy/QS4dJjf4Ur1y5OwVxKiZs6p2wjPb6ZI
AGLDjjt2cjTIb09TZt4uy5fBGwPucqPbDynrgKE0Z5PN7lO4l7cGdlyZmHKUwr+02F4ahUcYYbPL
yS6ZGVekJfumS1y5WIkZeaIaDcPoTuBNPSFQBax7nkZc9SGlY8AXraWq9Wqiz5hK76wdPu3Okb8k
FsiKlQqAdHUYbLO0izmyKrNPJsQa1J27/bITZYG/N5nEXfM7SR3gkhrtMklhIGV3VOqQzsc3CRd+
Ygxsi/e5bCUZWMhJiQ5elIIrborCn5I7K0ii1aB4/A3/S9zGvvrP+TGZg9AgBa+WedkbHJfVMcF+
TEGojssmoyNJYDedrh8FIv6O7NwKSVMaGBkR0MssuVOV7MWu8/0g6rXVhxJgaftLw8Q5KKCblMCj
+HyRVWs9fd/MjQxjtp6IZEbwmACjLia+Pz/HZz0TSbzLYi7Zf6esPHmEsdXwUQsbQqXdyeSfhGrY
AO70shqoBTcZZkLNr98rXv7btBQPRZZIk07hOgm88VjmjM5iRMCyHS3JM7lOPkNpToyghiOMPKyf
wa/VCBeUj+qp6iNiXotogSGPFZ5ELt0o/7yjBMxVuM3Nu19TE5Ac15VL8ior9CITSylSlRFnwpgt
H9VFIai083zRbiy9YRo/i4ESTjJPjfv9ggzzTdYYpw4fjJiV9JiLAYA448G26ggJKse8HDS+Fj14
wnmnKWngyAeObD7NlvTKL/jYhUFqU9blI9lI1Xm95M0c4tEhRXuB0n7g5MKDIeEtw0r40N2ZGPPr
lg7oCxugSb6GNyAwe1Um3SGsgkSzd1Zf+im3g0/8zxpih6wqkdnR8pw5zNoJ0Xw3ck+0xFTobd8D
HxAUcc2q4QN52+cWgOS6FqjMoEkNFI013adSrP6CAtUxeBs1mCvK+Yb2TDIJ7oFM4j3VS++DG1sA
zgn+ozoYYUxwVLM/irf7A6dcAT5zO9LQYGDzlQTioOBLnL2DVIQMPy4traYNgvutpCSe/jLK6TYM
CEbpwnj8df9prybCPxFdlu/JzOsBRgkVy+CZTFDK0XdsVhrm2JFRXasOzbnJZPczF/8+xS/9Fp8b
qS8P6oN8nP15WK/H6SblkHb6nXg4MuXLMY0rgxvTgUHgBXt61TD05FbdNbwTDRt83wEuzK+mvDxU
wwqPcRaIUNLfxoF0SXMwtiQNQGzZEu7rJUAFJoG3C6jFv6PxLMK9J0YJ1LDn0lL3kyfZXMPf55o3
eGlUiUTP339tgLFCwBGgUrz+jaNYJXgQTr60mvt7fpGynMaK9R3kAlWXbYjpqkcncT+re4+KkOrc
LtqVLD7Vj2RW5u1rkIsSeW6AsQm7x5HHPvEZ3pRPgeuQ5NshHcG5BM+DMXP5jd4F8cIF5jL4aGtw
wkzmG1RFDAjfyBMpKIaB8Vd8qs4A7VdQNwpc4Q2dUiwV33f1IZstdJBr34P4iiCgq6RSl2VZYo1A
+r7sXhP+yCTWfl1Hw1P/huHKUlvsR1g22lHAcEgdSLYQyMla6BH/Dt0pd8iAcAwGH0s07TeYKDEr
vkxrt3mmTa8lP/IAmRZccWjeYyllQF0z6J6Ck7uMwV2hAZYPXbY4MZazLRQU1+tUUwE3ltFDQ6W2
geiU8pudLBuSwEI6+EzhXSU1o0T/8MN/aqFXe5J1I4Wiq1D83/0RHZ4oLeUQU+cu57TugipJDVxi
bcxmnoMe7iYiDGCqoD5NgBfKA5Ko8NNaCFgU+KPFx87saEi678xw3rnHClma9xJfFN44KTWy1NF1
wG29binmpjcjdlcyaPd46D3C6CDFfJjSLPlywsBO3QaoANgJGrG300jFAqRnk1P13gfJLXgxR4N/
GquX1UR+OM86kiHrv9ablm47niclZbp8DA7HIygpH0jbzmKt2o5oEe28/HcHo4VX47KhTWE7kaJf
QLVBjpCbajsF372n+8Xez5WoLBKbkmNmM9M4dZFxGP4INLq17jHIQVyITGrI99lPMkJrJrjDKta2
VFbCmvZ/We3nPPgtiPL5S2iPVvUnXCWKKgfdfDuYzVjj1brFupWZE6GmeULdXGVWye6YT54E4D1M
3793Ogij0Ymm9A6/XL/VP+v0UgKVcqw0padE/s1iJE9pSRfhOfYx/pvsaeQJ+1qGtnVDdsW9jetA
jmIYBjHJwJyjcrQFj4TBMpSMkBW1iX4LWB7kwKkcO/KFCadb0761RtHvbvg1OCfmmqIVLH9a7qyJ
YZ3R7nHFIvmlrUJbf9kMRjt6PCJrUCPPknYyY3gvA8xEnPx9Jk14k9mCZi6g0Rz3HZnKf7Cceg85
mWcctw0noqZjn0x4yddDNzDkTx4Fz83OXvxadoNAY2nIwbvoYk0gfgdl7Cg2oRFshE/e3j23C3n9
4cH0+QvpXp9WE3QS4JS7rXWlWdmAEuiEqDtPpdeKb3xI925EpKawV/ESTqm6dMld6KC+BlAx49KD
ladhqr4emUoQasRcwMKZ6cAy/c9Rm4Ddz9Z2jclxkM/G1GJPYjUo0fjD7PbGQMyK0c++Nlertk6U
BM2OynsmkpbslBUPD1pgCvcpUJTUUX/lDmsL838tDBBzluQ4b4tHwIAuLqpZAB/RCzHvsaiTA58H
EJMQh2sJLCuMQ32+ThrWXH0A1Pxtsc4nw3gxuqa2XbcaOspRLLjeIjqx5k4bJ6vDerXHZiJvEqi4
oeThMDTyH0t2S/Kwue1emwpUBuPj4C+EvSgQKorhtk3De4BetJ5FCaqX0uytNt+6xu8eXDS9DuyX
Us1goQz5mdslbPMtF4ny+L/eu1C/AOM3c9l0Xfd1Amv8vyBiBK35kX6aP9hYBUmtKmurv5Nd4Vk7
ZUfniZE7ApUWAe6JaHZX7G5iBhBYQDqfSAe+dO6SfovM0p6DgA37AGbK1qgyMkxggInRgXDkOksP
sPeGuZHh2q25W87pAV0wVJkaqJBxvuB9s80lSTtp9t167D5JuvJYPsYfsUvH+7zKWfycj/c90o+e
JT7j5cXZ9NACiDAhncjZRlfrr3tUSl1sI/ccEcHtpTDwvAyUg4Z/YjGOVl02FotSA9IyAXrys0jw
ELVLmCcwxvbppCgCm4njFrx7VRi49nO8kR1nDTmZJosvL6Xju/wjx+fE05WD2ca0m1KebQUfNTv0
RX8QwuhuyiqdXZ+UhlYF2rgDnbZZ59F2xh4UfCJ1DIguKayDAA7PDORIoRH43cPUCWQGcUi3qA5V
DGjcRcrewoQYz9ENe4Xa13nkMp7a+X5h5o1V/4LLbYpwTHCaNrFRl3go5ebtNvgmf7spUvSXRFDX
ncRBClC9dbdA/cqOV76sI/K/db4qjQ0V+tNajwCS3rxFL5RQcRwj7R9Z2/yz21uPDDh9OJkzJzs2
IIu0UVKSgw8AtoFE5iCbPxlbW44f+8cAxUM18lXLrnq1zPw5QfLj8DRhtcmurdsxkMIKGWrHe/bi
5gkaWJ9Z37oqvPuPi0qCFsD8mK6vm3qOmCqBwBN8Rkf2iPO7kzxWkeFSHShnmqgQadpGD4GGQssZ
q6SgTsqeWwDXtpvjGsHqYYGfaoJCBeNFG1TkrmITLGXUdVqRETM7ieVl6HzXvNhRzXtiVV6XVFDz
nfPpePOJaKK9+4S8jHWB3tZdw207TI6dRho9HxHdXLLZ1KRE5jRZWTbHcw/TAYxPA5VkQ0QzF/j+
XVd/fPDZ4IIT3hOnNCeTnaPdoLgb90bOYjCWK8JLb3oM2cFriE+lZ/ADn1qUctUiiXCkcbFDNOwh
u/gsPMnMdKOLKiek5lRV1faz+2wS3AgRR3aTOc60gIOagO1N+W3yH5KM1ZmZcjOFOx/BGpIzLzvV
Egc2aU2ByUUlNyM8+ZAKYiDwQ4D76kyHU9zQpQlX+9UJO58VmgK033OI3tM7Ap5n4UBWVVojox2+
79KRIO/0fzC9/R0sOOYO8xBfoEVpYJ5Wux1EEzVvBh1JRVRVc+I1voOFMYbWS+KXgI3un8i8TtJ5
XsD43UJBmlHAusp+jgS6Rn//Hmmx9WPsGZO/fwEx8rY4r0i3LHlxPrVMLVEW7A+Knr/KyMRXMHjM
MINtZ57fY6t1yi1QOIk8CD3IymD8KooavGy+jCb7vtV0YzKMaBmEOFYiYiA/NbUb03w8JcxdYvK4
uu0JsQ56wMUHD9Zjq1Bip8nmvAOpX2nWnmhOdCDhImQiVT0+cYMwo6XWSCVZxzxfa2kBy0glf5Bx
l+Qt84WwYkmGW91TcbNqAo3cnCTpYGR0ho40mjzbG9DDBHYdDbLeP1pGD7GoE04qXETXY0E24ChN
mvnw32hu+nZCaR2vdaMiPqrazHoIY9PTAYwIUZqb/st4y3qgaArs/iTRsV3FF3gcc1cLb7Hx0Ng5
K8L8pIR9hxBqYoOfqN8g1mCmkVoXJCAE9Zu7hVlDAYQMi+2xzEtnPSX4mPICf6kiex0HrgwqhVoJ
+03uBNBlezXs8D+9f6fnABSkDXz/+LOgO/j3TQ1QOwo5YNWl5SkRHf3muzmIGhpcN5H8u/Kn37P6
6HErLnlEGt47M7PuXXeXbyEf4Tity5kRz0DQIs9J7fQNuFs1j9z70N40aVaW4V7/uyEcD4F2d9oI
3ocfEL7boiu8IEbwKTOglCiz2U/bubcMCfx3b9Re1GWHYJwh3+VOnOwMRLj3fE7um39JSJAvmdCV
wHwkNdic8E8Eaj76Uj2oTHcIM8uOy6o+Gk3E5BxooeHU/mmSe4yzz8BIIq8928jjTHg3Ek0LunSj
3XjHFSm2/exNP1kFAMNjwjBgZ1pnqbKeE/MLuAqQysRDkcMuXyt9BcM4SwkIx91owNuQaWKwNo5D
jJ4v90hMGVsjwqwWOcJ19FYqWJJgqduvFkiu6lgMbkaPSfmvH3IadkdVaMb520S5h7I6Ew86yP3Q
Kbyc5bXX7R1eMssk2/m/mFu3vV9+uaPaXcxnQJ9TkrnLRiwMK/WnecN+IP9ZHTjRAsX/Rf00y4dI
S8tHn6vVAH3BeTQFY9YGXZt7gJw10qUjiitZI/I3KKwBfozI9Rn6wOU8ul6lXEkunKxKoeRVNBNO
erEv50KcAFWiGjmLPzZInrGBD2kXlOPLiJegS9rjxQwvNWiEp/sXd4MaeYrEaplppqgzFrVWdoDa
ejGa5vxJ0cg/brbLW1U3TWnz2Sy7X/T+ZSrzL/pXLsvFh7raWPhK8lMyv53x3RLCW4rmF2sdT2bG
XxUUXdn+kIgfO+K1cFWq9MkjoxgHTcEFiXw9VLoALqYRDLwuTY1NEGURX20Xm1p6tAWjG9319hvp
DpunhSErtaTzz0PcgHWFy+qqCQv8ghssbAxcXMZLElwi0+ufj9u0ofyqJU54LQXSEtXS+CiZf0Lx
oS7CUbcDFq6rhOO2RjMO2DW6VmHRPDv12XbYNT4sRVsIAYi3b2mxGh3/bAVPBJvMG35t1DAitvHR
BITb3MnmvzRQ55eNRO7sUJO8qL3JYUMHR9N5opEvTpvdwiyXGOliaQFMb23eactipcGsVMbYvoTF
kOI/gvcMVJt4Eld+un/1+ZD2oXm1V3QQRuV4VGvdIxR/QN7/l1qJx+p+sZI24mLvvNk8H7HFoz53
8kpGnqbKtB3i/1Ms2FNm0Jimuhi9y0ZkV+ciFqWLSl/x/CnYiajreR7GyaOrtN+VoqCYkneFy4m+
Z+BwehNjiPRiSeEcJF2yz9oYvMaSPNMiLh41U6OyoZLWdG13IUTVJ8VZ9Zdozcgn0xHYAqwYYrCs
t+ES/adrVjx2iI/kFpu9SinjVtHx+o32iyQyoAHxKGdZuEsImtysR/5x7m5ZHwDu/B9pZpEBmNXd
R06/QACSa1OZbWgUgxjKa7afyV7kQ49SyGLX9mQB1LB1pDvzbzlpjGEuzC24IbwUCzqqhvqKey0I
nMwA7CqvZe9xt2N/3nYckR7IlZYnDNT9hzJfBfJibTJJ8p3Fl7sPzGEd+zhkZLXc1ckVBIQFblXl
nXrRLsFtMU3QhK22YMDBGqgx+tLLohSn6D+q+6SXIN1kSMErwlBycHC01FWLP1g9FidC5SxoQkIG
u5Q04ZaJ8F84P5DkkRYHLLTevriD0O08/H9dkV/5zIbIpascgXyC4qTQJdI+YYLchuogY2oChiJS
jEidJvo2Ww0ZXwRECJ4iLJV3Y0xdotqyg8zQWb8ztTqozy3tC4F+5OMb9bPidzFv+Qi5AdNdthqz
nm2AVigWuHvGTko41hUOuBmsW1UNDa8e/68OuBgCIGmNE5kWK4tF99pshjM+4fvADKcFNkGxh54L
qMjkriXDWXuwKjDkczaGk8ogzngVjGLGIZJJ0UzaQyZcykFF+xc2PEbIUVYGu2bWQ2wJlF4lVJ88
Bn+6uFVh7TPbeihbZi3c9KiDbP1lENb16irpJIh5mV1JDiygbAOsUEqFo29asut067wJxpPvUKdr
lPguzEzDeBAvGq6nzvnWRuHdPikvFu7RCPtBmtlM96r3nTXLBa+jtt1qEPFqYJYVc8Z+4QBLyCE7
gQavmPxu/Pvajam9dFHPo762haoxrb/jSX4dCLhHJQKp0mkdhB2hBcnNFCAeCPpNEiH22/M9kKur
H7xQUbJJXz06qt5xn5zkFFMHPVqXTr2nipGqaGWa253dlcb1AAlOYcpzUA7x/80SfbbRlrA0jinE
edSI5D0+BdGeTEZghnN1kGUW+0vNRZl6w0Rdw59b3EVTKhs+cx99W0sKr3B173wE7apGrS+tu9z+
jTS233TpPDEa5psiVavUQ9wGqHuKUOsylAu7cqH7lHEtiOq717mH5BsaezHXqCHyOQs5uJ5C/Q0c
oe8iTWsAJEbfXZ7crM73CG+4kHYO5HbjOCU22WzDjrqTMhOKuwLymzGRhpktigqBvNkvVPMDeWr9
T3bK0GEa2W5QaKgFsfQcApsJ34oAh5I/0HV6c6HmBJAAx92MJ0+XccsiUnADoRC8za0mrMIKNXla
Pr9euQ4luCCg7igKSDzQED49Qy4SsaxYmrMUIR3o6sQNAstKv7R21X4OMcI4MT+Djm+I5Cek2qeK
sozv//DItFJX+qpRwSNXF+GKAoQItP8jwjOPYfIwGJSMWjPQNXppiRC1HdLP9BblEi0ww/T3IxSr
bPkHYF69UZZeCHDVI3ImmrXffPGonNAoJjANcGBe8CUSAqn8pzopFskKmp2/7Kbax8oUf1ZuAzuZ
ZJT9Cnfd4Zw3n7JLcR6WjQwttEjSgNh+GNN2d2W1Sn7V+GMohuZqgjnwygJNrP3JEjaaca2uoLQ5
b2zvdjllc6sx2aXvQ2oVh8eN74l/GFjJmQv55/hTsM52bIbffJrzfuPnIb40wMsgqkmscOQeEgZN
xAm2qzI561845kkmg4YpN39A8guxFHSI30y+ZVoFIsmcliuKM/hIQg/cTBlqiShKheCBXBcoMDia
RpCl0YnZACMsKjg+5gaE1y5YCiAz4xXjO+wrzK2gX5y0Gep/isarcAgW19LNBZMXnd1mb9h6Y9wN
8l3UQ0XYl6LKo591qI3mgKT13HXLWKE8cvgWBL6rD17XXXmY6bE4ztymR/6HbLIGjPGZkT6HffEs
f0LuPz+NcM/LRKmSS2vB6ypYwqoh7ks4XbGuAnFajF9lFuhGoJyfcgF73NE5W0S7QUIEEN2ZALMb
DbjC8DIe9dlf7W0wkKntoow5RPWHQeYQmNYponO6FYXLITvt4HzBTk2h1DsYWBFvTAsyv2zdtN7b
/6KGJTmzPBw/WunpgjBTky3SYZVp+dzF7E5Ux3SZC5Av+je3CtZ/xY6lfo3CNN7L3lH4aBR7FjKI
7BvuPtQg1WSnXYH5y8scYkOzqXCGWeysT+Y22O9ePOXR0YaCOoa5VAvaSV6GdP5F6h4i6Eu0FUSZ
D8VTmWt7zYazrMR5m4FzffNgQjKNGm2pgAlbsTqVDBXzDKBZ1W9nt/NplKdyoEseoxfX9+ytZkpv
OeZOBhbjOoqTO76tV7pZccEkWZ3hcDBf2IIIkmlpAv4t2NPcma+BBXIOwrtj0Pi8Chb8pVAQ5Bgp
4M2r8nCgoL8gMlW1Ne+BL8hj9LqWI/8Sl5Hw0h7zd1zmJ72kj5MjO/SZatW5+I8NFn/jdi5AnKcv
Bxd56f1HFIr2oSAwd2kRiUQgQKTZDJ8H305pc8dH/y1ZlkFJiFWiq5XIrEFuRVX5f42yOOzS6Ffl
8E9QzKphFPAcOyCajDpjekrnYISndYf81UxriyC60sPCj3GNXxZV55mwVQAhPW+9Q+hwW0+apfms
BsKNUhFM4OkK91gT9o4PMf88i9eXByXyA14nAGQeJ5Fn3CJYu8FOxU34ue6wuVkW8gKSt8C08R56
23Z0mwnmfE5RrRyAmllVCy8MHewaH8GbMBKZJJDuaJSvivFbO/6A+U35VMMDCofPlaTTdemsC1ON
GNz778NbxOhy+R5CPGBoxxSO4JtzgHHLK9JlLb/UoBJLt+YjYRYijBjaaF2Wvy5WIXGMEW7/nCsb
TJjU3IF+mjmo1CVcDLE6HvXeTsBePi6yDArKS4lqMq7gxpm0WyMvkwAqF7Cv3461IhS7KmnERpGa
lotR9YSvRJ3cwwNXaHUBdSSKg9XGI73vUIDZCk1gj2leEFRePzEzYFv6Di/Hw9hgJJZtmXSyxDkq
qBEBxJglnExuirNdaCLgUY0BMtTTWUqnoZj9BWZEwG/pR+CtYiC1Ab/t8k54EdtB2qGRaSiyva5d
2pSMK8vM5PEt0pMkk84xhDM+gKmkjmgr5wGwTR8Od2i6etUXTbC9nq7BGpMOIYrWmoA4UNchIMR8
QJf6G1Qn6wfs/480N0OxHeP1vIiops30xZGoA20QW1+u+UpjkHupPVG1z6NHiZuSgF1CVVRp3Nsu
1dAWYUB8XKYF/ZYY3410+4gO7GNNdpfQv0J2eoIvkuN+JqgmnTCaEozM9CKmsxkoeRbG8z/UyX8D
/1Uo11hIDtWTueVR/Q0091z6FSCYGE5QGm8u4qV+BTky8I8oK8XMHygiedm9wh+HuNz5eTDYRu6y
u3RvMpbJ2WRi8lyFGUAcnJVAcOyqxK0KzmKCkl6o6lxL/D+F5Xo27xiKsl7VPZSa0h8b5k5ImLPC
BLluFSaoQhrTAU/KhHCOb/vyaHYJmAZmEk3gaggkoxjNLJ5kYdxo0jW5++2InUlFc5x3BTY+zf21
euFS0RLuCxOraUMX9M/XbFye2JuBYI4rxFL56HFXa73nC0yqXJHmsuIhsrlWE85JduXNe8g5/Y9c
2EOz7dT2yOoonMMdSxJcuBYtRH6KpZ+N4sQsN++xipYQv8YiFmS6IsyW3HKbLS2bWPiYemp6HExq
+rsg8wFbAMZORhqYjmAYOznOCFvh1LvROeTPp+Vshp9R1M4bP8fA2vF9e/EHnzzQod484SPVbDpK
ZQGncv81Zn9L+2y37Z0j7eTKRQODvoaZwml93XVnp+Fkm8mCSkUz/zphkkhlm8PeIsoKMvW3GRY/
BojcKBXXwtk9+vvWwyUQcaNJq+cX3In4PJzQG2+BwZ8pKUmLkjEuihuWqSxuzsVdNRvNmyU7Ox6f
nDMTZDLyAI/4djMTgva2vd4n1dRib/ay3z2NgVy2HFzkvcvpHZkBpTZ7afW9rMysR7XjXFrMhG0X
NsFf9X6Vx+153MEIEN2AQfn3C1pWRe/z+84KaDuNw9Mt4EQ3Cti+0OmKXWABPezn0j3msMD8jfCp
60ftrtRcbeF+rnxHeryAX6V8egINoOguT4qi+OW6e9dDNTWupl0P50kjkrrz8jQkj0/DtDPo/xu2
oMtfgiMske3n9tmS8CqmoUCQGBoYcjdeMnVChiV4Zx1rZQBrHoB67HWqBLIUVzen7wIyu7j9zDao
BtDTf6cyv/T8qXX/aLh11TDqU2j3Q5iIvTCyegDVoj8EBJ+yw6rggV1ITnPiRE8M+6bWBSGH3Rd3
nIwMhubVDKAd+8p3pfJMds0yGaevArRvVv0eQgP+pZnruyhJa7TjpKpsbucknD9vE/1nHxnN0Jrh
rdfKUftT0FMf65qnwUl4kFVMABeEzzHHM4bdeHTkYfn7R9RzbwAJ46LD9VXaWGBXO6pvayxVlBRZ
Yf3OXQ52P9AleamRzfnHrjyLxSXOUXfXaoPHh22yVvURE4ENx3W+bl7Sie8Xh8Hyurmd9MqIeHS4
3qg5x+1zP9ZFHPyJQP1dCrt+Tdp9bpsUqV2QR2dZoVuljyzIRlBVXmrP8Z9//UlcFc7cKU4KYziP
MskiK7UhLRFRXWBONofbRwU97W0Z+e8ymw5v7bxkMwzEguE/9VXd2pCGu5AfKXsvvhmYcbWRbiej
Z7OwqN3UXoed3hSiI5MZ31sFHKhEG9//QVPQnpqRvhUM2d0CbyDSMKQfINga4pFak1mZUkCJt3bJ
JZ9hU62xCKvN0C17OeoXJV9xuXDfOpBPsv3WgC9fwJlqswVOeOwQb7mb43MunUNmP7Wecsmj2XGG
TRTWaB5JvCw0xXqGvsQhEF2ss4++CdnmynawiFGSUqT21Q4aFqyHSb46WC5qj91hq6VuHFk3vENg
3bp1WZAosuErytZKaeUgeIxdN4dIzkSoM0qMhaxsEx0lPY2g40UWWDxpWnT9H4gUftwxlMlmdmDA
bV80pDlR9UBVl6tDKHdGGfI5aWTifhhh31rWGR4m1xHRXiLsM6vqLajm/sJFFoDm/uvTlG1Y8lLw
4heSKWXJtxluI8KLW15oOV7TiZ1lyrBRj0PN4laa3+R2//tmsO1cUMeClWctytt6A/eFdfp5r1+0
5XBjrjSHDs8iToOjBbIDMg8zfNrJU+j56+A3xivBpFBkiwqpiJuDb6HTRIaP8qo0w0DiZU0MPGD5
qywmFbWZ+G/+gDvRxTAZma6aijLnd4TFssDcdS5xCudMCZdUG+qCKSfPOGRq6tiMy7Z5z8d4josM
YSut1cQGSz/HF8hdpMyt54csJNvnEiKvNw3reELIhv0qwmatUnFH0H75RZBmbYs0UM6SShNRsT1k
58UTmj8bVkOfWeXqU0Z03pU1Ezt+lclspNfaBJYAjmXcC1j924uOnAHlnML2aHqjrhT7XDEFE35k
SIFsl5J188OfejITtZezxNyIkU0zo86P8y01Ff2uC7FsCQHWZOxpcaGExxoFwnpJT6ghHFyRqXYv
z+RNvjme8w7kc1KX5qvuENIecKhal94aEh8D6W3wBdYlte2ousbH7+IDDbZPaKuHCU8PFryrViip
sockFzvqHLBLP0QH58a/I0Qjj2zxy+ow+iFVSip8ePq3UnL8irGvG5pBIBLNxVCGGImxRWPOnCCh
DAy0WdZ7WAwUDkBwqguMltT42EF0DFyfiTmyzTlFrBfGnuflog+2aIv/pXfGsmMXV9WoNdyRL9t2
ZNL/j7gnjI/JSKVkJzdVGzIS0OSO6BN4e9LWc/RpPtUhBo4ZIZsO6dkU2z04QAEFEdTi6Q9J8wv1
bZfBB/U5CjgOr1dn3NGXVHqtzOO1TJUln2pQ7sTHyP5qTwtEDd0gHnliz6UJiIu38XKlmdUQ8A0G
Z10BARRTc3JxbSjhXuRyXnw4/QGo8Dd/f4gguQ3V0AeiY/ZLC7Al2f0qkxkGL9X6jdQkDNuyTSsb
EWFA7UqlPIWknBzcaO/O1bU74N3pMhI23mA8VWQM7Tjyihpzuvlg0Xm+d/UnIbTL/magnW2LuwUb
0TAgnvoIrPlvMLR6Ae3FPNMcqwX5Ej/biuR4tFhgXDY/Z4yex5vS/R5bd0qlXZrfy12+s9WC+OuS
xZgtzvGn4GO0hnw1ESieZhtFR0sWPnksHmEpQ1vOLoL5cvPNQNEb+jP5nLSD/1RyPwtrdafvYf8Z
2JPjHjBnEXp1KAj1ATPYi3RWUa/VHbh6zAodh5n5JLyO+as0/vOM613/2oLKzgjEFehqvR5DSoxr
V0mt2UrNjF6hjt8vak0ocbzkYMIfqCH5atCyboYXvnlkkZ5TtZcMYThl3XYrzqh3HOQl18szxq97
GVeZI+99DDKHViw8bgYeP6BfyMLusU6a/LlcldZHfS08v2bK9VOLX+PzQALDM7EJyXlszXqn3voO
DZgjT6pk87RnetOnlnXT4nYUVbVvDbKAefFttemQCRtOw9NPMIcsBEqsDYUgAh/6JrKJqFdZPXWg
yNengruUtQaWmbdnJotsr7w5I4MVM5hYgM5pp04RXw/oU41KBNou+qcCE8yWbRdooJXLHxhK/5+t
XVVlW7qwPVM8BawtzUOMUzSkdTnU8CuNes4Dwsb2RehmW2THxrGjXRgl7uFYPynUlr4ISwBBY1vx
y1cEgYCb8weuMAFf5Vu8efNGhYG7QQD+gJxIF5ZGSnbQYlBH2jSwvI1UzwsEJ78CHu6qSl6nGaNr
vSUQkSMEDe6Jp4p4Hl1smHWrxhNgvnzonWSZS0UEyYrtTBgTzB1D7mPr94Ev7LrdI+qzQe8klEVu
vxhT9BgagCBvTsATEHOzwhWnF13ve7Pi+F4DKCT0FSySsNwI2Fn6YBy5tJNyHgON6OARWDRYEB4G
o9tsZxetW/Rk+zorIyS8tc+LPZ6kRz3CU9jr8bD+LkjBh8bLniVQYmcpABhdbGG7drUbLF0wEWbT
BJacRwoM3Fz127y0d1XnBGZLrhc1ROxGqCRyCMfYDXlDD8NWnqqv0qZnIhbZE2EFCenquFx/VIqE
t/rW2Aa/LMSWD0ud3BqgdqhbH+/ChNMPlWDUCSRz+gUeJ/Y4Byfq0Xf+HGcxCFNjSIO3Ecd/nhke
3JCtoYawQpAvXxUf1AGd2AAcNier+OiO66/pnzmLiMu4NF3jiWJBDV8HilI2dgqRSFh/E7UujXXH
JX3ghcW9cgaJ0+Knpp77dBRBoQrXHWwnGzwYc7w/C89+Mv8ZQXHGgE5Is9GS4jn+ZKkXb5W++rDZ
Iu046zUUuHy+sOG9zNYRBlOzafFyVybpSlqpcerz1rvMkbM8UBIsCIF3UHVQRjfS13s3riBwHORk
YU6FigPCeYADaILCprYwp5v6ZfcdJbf7t+Qo6X81QOZFflAow062vBVB7/iOtEmAhQpX2dsjeV1c
SWvcTNHzXdnRvZ6o5FP3Rmg9dtPo95QHNkDElA3EQhhHCloTqHCV211zjbXlvih3Yep22tzdUkKG
QRw6qy9sV9XWpWObOs7z40TvVGVl0XxkRjyZrzcXkNbzLRCeFJHz6sASLUnZP4rlmXoQIEIJFimv
3b+Sr5bLHC/CCBt3619DJm2SH+M/Dg3SCaqFRfK9SUEXxgrz0YS9xy9VCJvT65USb0/Mt06/E7Ka
cc3HSLP+uCCcztZxaVZ7zz5aDrRms2ujnhrJHdk6l0t92ABWyr47oWRytMMiWk+7UtEXjUWI/4vg
sULBLppTZKSY1D2PSHh5xiHslsf6bFuq4GLmhrU2O1MVzaIOuvh9za3Sw1cdQBVZytGjAkweqSVd
5lkBOE+EhEFtBsaNnQO9zQ0ktkoOn1mRB3NNHmNwbpKUF3TL2l6sRQzFRS6sxZ91wfBn6Epeuj07
InapLlzuOgtFT9gFgVYx7bmzwnmqUhV4YSBmsmQzayWl6jLStyUq0M/Ma3+gIh13eFQj/JPw0w1u
QuLZsz/2oCZ8r+PPA77W1ZPDxJ4XwnIqujzKCur0TOKh2KJZCAqcb6twINyAlUktkeryKzPBDkFz
b20os+R6uLqZeBJ6/PtQvrtJIrT4PvHyey/lEd5G+7/PHoGmyfdXPvE6zZLLX0g/jP2CePKb61LC
IRJE6tEV6UEDrHi+lN82sxA8ixdbcJVt/tHwYBtYA0xv5vLiznE76JtnJFhUTFLbJvaQeesnGnEs
ZK/jWNjNTrcibpy63o0WGlCFkrqR/rMPLtvdvkuCpJJlWuAUWGSNGNsDEuYpAfrQmjd4MDJJk/hT
VowfQCknUH1cBlmiFjx5ZDpHVc0RNCOc+HJDfuvmQRiXdULoy+jNUmLhPV/Yix8wr5FzYoq5dJU6
4HLYLeGH3VaSbkpqpBc+sgUdHTFNouxfjKeo6MNvYukjFOIoC/TXfnE9W0A2Yn/QT+NFZR4YfHwb
n6f6kvE0ruiH9/vw+TfywoFBNELqnCLemK4E4IsbHJ9WHLQN3JepG4skyqzIKW9Yc8VG5C7Ejjju
Wx5x8OEt3qHEh0vYLLaLyZG+ZPIQUdN262Q4OS/BdXJt8l+hTzPG0knLJKjG4vAEZnSUahKOeyIp
gh3syfDo5iKQWi27g3ogUBIeMJu7Bhj/atQ5umnBIwWewyaiQeWNuHVlAQplywvC4OIuVP8mpP3K
zwcy8tebcTTEFKZ1owNR2y/KH49umbhZc2grN3z91qSbj+I9QG+thwJ2KA+nW6mlfY0olAWGzIu0
/FRph++X6gGpXbtCslNtae7wDGz+uLFjwo8r2tODfzwm/pJNlZ7U9NodhdYZqFf8F0UUMJ1XSn1+
b1jVNW7jy8USTs/Yw9f2/T3oxWla+VoYFcrasSgZ5mYV8Vej5uqoC6iw3vaYi4iW/a+PiwP15UTg
U1esWix/atgX63Mu6qyf9PklKx+JanmLzW7OsQsvka6kPSD9qxWonSTVks1MEj8H9z0skwBk55qf
be7e8VBTie3ZrT1ektfkS2efibZxOkg07Z7mLI1Jsm4/gfqDkS17bCA2fDTcM8JmfkSIi58mJKsv
Rr8J6xVPayyKbg/fJVHkYonMUeR5SYzgRs3wxeu7oOti+HXcvl6ZlWZ2vxnQuLRHomYOcgcVP7Bc
Rql5qLNduhvqKpFRtzZgg2bxzo8ma3DyfHVK4+QhD/1kWJIhoPCEpdL0u//p2SrwnNyhq8A7AJef
/I56IKuvKE1Nvh4NNFqxzdDkfMwPjLvBPJf14JAUh7UiZ0Et997iFh77Gzpn8farhdapiyn60ii6
njobCdX/sdx7gOIgsjNLoevF6SfkP4h4pQzlXszg2jDwF0LUpKk//CroCqWZRm87RNOEgJhbWiEs
Yr57sndUbBvcyWuVnFm7lxRIs8ArdWF+jbHr2lX+qKVcGkwjyQi7+yUXfDnE4cQFk0yOvNlQdWqv
TdjkIt/l7T7Ufb5sr2xW+7kGY47KBUjwc10/lHKo1htEoIUYZXRWXQOGL4xSkvf5nESscinFvGO4
YBrv7X9L/RLi5BQPHvobQ91t9YoNiM3qOce6IPdjb16ixpzKEvQY9OFCIrFscDkVCO3tAwT75mDt
CZMHqkz+HK6TS4Q9jZTcJlrar4fNBfJpeIDALOiWG8GGhQOHE+eRgxM2QAiVbRI0kIe1LG2cZmYp
tF/pFlN/7TGyw64KWssHf9B2tT1bcGev5cqkxpslboaLdisaB6lQpp6Jgu/4HwtWBGMXmDyB5tuO
y7mnWFCMc+2Af5c0vDxrQkgUQEnyEUgihqi71lWiJ1Pou4BXOiDFf0kg1v5BU6FGCg0nV2aIS3Nu
QKVfo11zn5E9FgYVdXIJ9W3xYirhX9kQNs7fs7dF8K5L1f5BufzbkMzOwjuPypBAKFXb9K3pGy89
JomSRgj+4TrOO5mWLzVI05zFai6I89QRDw7TOWrn58DDD8u6AM+msH1MXDV0q4bgsp+KNzja+iwq
ZwnqIM/ItrfN/0mix5nD1Qq1A7l4atikU1Fo0hEIoJQDTvpKr1oFMMsIbbRMDGo1R4U6jqyoA+e4
bqOMWYNiwoHDywmOLPlUrE+LNKWYHAFGQgz7Qf9BJUGbcXmVLvtqglgEl+XN4Gh1F+ZHoZiog/W3
+cfBmOXn0xtLpfVgXF0POlD7tPCNvVFDrDxOjvxlJMQgAg+bS0WLGfWPKPFWoY7fybEQuy1xhaek
XLj6mxQwEoYt7ASbX3T1aEh4q3vgGhmpASMy9tRlwNb9V7cc7EjpuqiTITCbQOTcZPN82gM3l5vJ
I5Tf7YIlcEf0RuECOJ7dfK9bGAuZgVEgcXHaxNEKEot1GIAhwmtyP4d7AVXcJJh0hMyqC3aEAVWy
vqSaUkq6TYbME6mKuLBcADJjOrl22V/mM2/CXaCvBbseVRFxphTyV1uDZIyN18hOL4Mde41pVtUJ
MEBWOM5ZGEGTDRdSMa20a+ua6JsVIg9fM7HscsW1aWbaGfcuYYfS2EQ0Z2SVCyYLhXWXh4sluLX1
cXOxBtr8ln+fhLB0Lzl3GijHwu/bi7sKhVE2wEQgiUXOp8FNnuRUitjfhWgkvDTxwwLIYheFXqwC
VHYD6j2sdVIqLtbRq53HO8w+BYnQZLiToOyiWSWoZRHhbozc42ytt1ays5DkbqWry3B5D0gCIqjd
GBflBX2w262Ftpe7zSq9TmZ/j/sEIzTUB//6evOLrjy1G8chrMNytymCHRWqmXLp+E5ipuzerJTM
NilMVfO171YAvrwLbUIoNC5AZ2feNmP6aE2ytH4pIF/02OPFTt8WIoWnDFgjMN6PopIwlIDmfc7U
rCOMbjhuYxahg4K4chsBySWIz728Ziz1WL8veZnAxU9Ft8vg8JHPIIytrYxP8OYJ/zs6DA0tET14
f604swfwVfkdV8Yq8v/DM/6W+VoW16qI/qS47EkV0WBU+FIOXJmtJcf04+fjeGfjl90n2jfWqMpA
egUoTFx0HkanRW5hRII5o6Jnkj1Jps7p9VK9yBVr45vaDNB2JyS1qsBlt7a8684Be3jECqfadrKf
WDmO6fXFswRKLoZnSKF+mMjArFutmECaHvbcEphO3iljPKAi36dxl9OyfzCwUEXN6QKAy7p2vkvr
tCbMtVAVfUIuMg6n8MdD5su+UCFyNnAZRZ+k3p26J7W60J5rYv3d9MQ/ALG+1v0RSe6eof8zYhz0
qyFjcIoyrv93Rykg868SurQKhzgXNmFnBviifIDulYAqxjJMbfX7Ipoc0j7AT35U2gjnHVoF4/n0
jitub3AhPxl5g/1ePE++YEsQy0XJFPgVjXwc0QqmQWy6uQ2Rrbi+Sb/ItwJDGB6Q/3DgltPecuV3
MvByF7BYIPUJCE2i/UmqJqmT0Rej3tUV/UPRjWWBhZEQ1rQQ/zZmANwchuALDBOsBhZcyG4cLNQ9
87kIJ/Swui3xxiDn5j2wVup3iwdkZCvADmMnaEBUZ2JcEsnPsiaj+U73KhYXPcCgMWzLimiReIoA
Esag0j++s+cNREn3YawOWIrXKCx/LwuDUh2YilKM4XTU4d6VrAbnQQUlkAK2YrvjYEURgm/sT8HB
dTnNAaNTJF9zhjI4kIWy4t7kiH98tsl62+Vhl5nN1LeehrZjlOeU/MENHSaLRV0YdoPy5GhMRuvZ
qgRlfnX6HUqlX2avLYF60ChY3AHRzMemieBcnfpsTLW/GHWLPIeIpqmGXOLqQSR7cjELbsAQsj5L
9hr2jQP0wJc1G3HzBk+qHdVGlkRS+rk47ZMcPD/i8eec7DsnRIlzeyAhdC9c3E0xYgX4cQUc3+wR
Yq4UDuX9W0HE3j53GST6tIJ9TyE0LxjBDn3Vfy45k3Tz6eXlfZGOtwr0jKsKwakluAs6vHRvYVFh
HJ1RW7nB7qRt4kXNzrQVwhw2ppaYfbnRLglxvv15H5/siFjyHNP2szkqJ/0mGXXHhGjg/eG7L/Ab
wRx9jn1z3aHeLB/wNQuiP9envcgGWoyw0966g8sbP7puPLM8v2qE3uB2HbGR8dc2mwzdLpz4VTG1
PSfaqJ6a0PMgq6BgOx0gHyr3jT1OP6aqIw3xX0y7cb/mPe+9FqdeWIheq+lvoazbiDFFFgI+LekK
vPbpIDNfDstcISUt3ZAUIIFGu7ZAUlJI/bsq2agZySICW+TZYc02L/CT03BGLEuAc+diRtiWWt5q
Y4ONOzlWnBhL5dBl6OBdSHC4MH4REiY59ap/jiccxuHKKdR4ginxy8mpCmUZ1+BeIXwuiZI/S/5E
ARgF4W5J6wKyU3AdNC7wfgTZDKRS8cdBZeatyPkD0QDUOGfFmTSUENY5b6KrArYspm1jVHTJipbT
9Wf6+VZw71f8YFJwenPUhYjkeRFLbBBjizKu/7rZDuTubYCKb7FfqOvTMUnTWHFcdCXypnoz41oa
n4W39x711fhT7+HPAUCe5SS6D8kbcbZ8aKEe0fIGPFS3IJDXSw3iiPmOJMLn7bIngR7ic6oMHCj+
VO++QWjDUcA8y6qb2Z2OLCn1z5olPONv9G766KFpAciajNM3g/NHZKS9QA+qbyS4wFYIMX1l65/d
AVQwgfwiuruWYcSlWUrQI4lK/wOzrdOIpJf9arc9zjn0nYwps2EIMpVQkfTx/gCB7Jt8jnajyMGE
D18X18qesgoKSiVMXZiBwl0hXm0zqSvvzNGE0UQEoxRZD0ZUQ3elNnOdvGi9kE/kVItC+jX5bv6Y
4INfHSWo1A1Ix1Q8hKESv4f8cOR6jM94X0pLTES0forq3TqQQX/jskjHwMA/xvYeQzsLEXL7YFvW
8sm9sAo9a/JBYrxaB0mbE8c2qKef6tsLemUn57AppOp28yggWrUtGtm6V9eAeFfTDwxc7ltzgcAW
D6eL7BQSBWm++QsJvuHXytUDfIkP/BxmXJN1yjebNpuLLv+iU+KDevOvExxQ3wLA9ZzmzlfE7cxd
DdOdY3G++P7TALZQCRevJnNzRtL/8kLq6SvA764wU70787SjoET90cXAijZA3GCIWqAG4RfGR9se
CweJtwbFw+DDTDVvLGiZGZgnNZbE5bH/kJgjdEW0Wf6ON+5SyTED/nWTrX8MacoYjYtGDiJ8+OGx
m1fUEn4oX1WBgnb9dpqcOFHCD6ZxjoX6BuEXOFbIKrIub6RKkpF6F6K0wIaFAkXZgojPf/0kjqBq
j0Evz7W8BFTBe+Acir/02Q49W26n3QrlSPOd322FFns4egj05lZx1jAFhSlMKDKLnFGPyZrbelE0
3yFiivFOcF782m2wGayPErIugwL49FsUAB+tQZFpjWSKw1WUjKvzao0aERUMDoMGJSzTYn9tsBV6
gDmX5NLVYuu2Oakjb3wpYGchfxC22OBk50DG63BXk4PWu1r11EkcU0WlpiXAAsjdpfRjjo+R0qPF
nvYnkmY1sOSjoSg/yaYuH/rvwl/2dkmdtOIBrTPKJ4ArHletnGBu7k0Pr+lZ/bVpnszYzaCAexxx
Aw30AXtHHcl/ms2lVb9PEamaSpF0OMQO+JBEjwkhDlRao2ZgaBNRSGKYAnimtMDEvTDFadvpW78E
cjYDyMNY4jXRIGaQbl4zeD6byxvPTWXm223juk3sF9BuT5CwdL4IU+ps2+Tegvocn+5kRSE/wheY
BeOOqmbj2paT1INtyrr2o2UqGC8jMhUDa6A2Hrl5S4kDJ1E4GD6vlF2KngR7s5Hz16nKzd41lCYt
Sr+RDHZV5GsxbGHu0vLEdS+UxrP0vfPY9LPCj78YUshmjcdJusi1ZZmCFGawSwEDlVHRdCUrTgRJ
X2sdH3Icr65GVsie/0hjfH74i+DEjKjTdWCGILDcr4LotYaxhtxwq78Nfusb2PWRgkuYUEpmTQlr
ShjXaBut3iRmlI8CqkvsOirPSgb8MXgGRM3OhZ1IDIAfK0nwe3TekHmE+Ah68g00ids6+5eRe95k
IdsPCposbnEeNEI+uH83OZ09Ta3VM2BL6rJCmUB9zzobRq2Bu+nraYES4F9SHSB+h4GpRDUmY0P0
3P5vkzc96RvHYXZtmmrqEIZ58M9B4z7VCyNF/mzNUiuv71uq1ljB/4C5h+6AnJLizmDsMOxHPIAF
Ax7nROxH01F7cG9DxN7dlYDO2kYcPlMIZw70M7nFyVndFA8UY7bL9WTqFkBpSPTvwZdeflTxub9v
N5eGqF747GkqjNgocYVB0LmNVAzLF8Oml+9TERpk7K7hzgp4iwV/XExy2cxCldf0VBe/YiD6L6Ca
3VId18sC+dJ6zkZVDrCYOMN8oXsOtS3P4Kd9YY/Po4oh6oVYm34P8Pn8whLSlyZTiJ2UJujwzC0W
3g806TbmXAwN9z6sN+ZSlWC5MqgeY+vGDB11+QPeVnSegDRT6uJtk6tdRxEeaCg+0sRb4F+bz+ug
PvGyWQWzzIg7vHgj16y2VAJAWRPskgicKj7f0L2e8TjnJGPtlpw0s+JMkESrfBk+CSYVgRlYOwai
9DcKBvK0WibzlAPHH+wHPVQp1z2OlaycXoIdfzrLJH3aOwFGwciLdeEdO5ULJ0Wiy50SopBwYRjT
ATgbPM5DcTvohxp3h809QuCaxRGqbC1mYcWfTK5qyOBGTV4CaZES4plOhd17da8gzjEdMaUzC08n
Hp5ZRb9QBbJL70m3v0Wl5om/n+5PTIoTVVftvfQISUBux4223GYnVSlAgYnGkS2/5CfPYzYBq97s
gc8keuindtcNEFFQMlsRQWfWSVKvCL7xYUw9qdR4rrLGZPzi/T4AlxqZvgenV2qE1hoRdoNgGhj8
A2gDStvUYizsmDy6YkI3WtG5EknccLC7sU86wlrM6cgnLEAHyfxsAVO2rLRPcHW9FlJQmsmc+KuW
Zcmp0XoqxFwvE8WB9bcjsGzjRf73WG+WX5D0E4nyEJZFRdkLZzjSsOabBq7qAwtSrSCz+lSXpqNh
mNbxqdOug7a7k4ez+Di9bzgIIz/1lK9LBd/xzKQTeMxryxkxEGenPptg1a5hi1j35n5Sa9vbr2Zp
w4cYg10JTk3Vu72XpU0Y3cbqSeJpWEXq6ZbKQHFwpJdaIuK4t+1Rb524/ypyh9z0ZeEs7KpBUpY2
JHW70Vbb3kYyzIObQsXGqyrRY4lOWlOakvbiemL1G8s5bBNzysztZHdn6+h573zEPlwg67B8+5sj
ZPgqFe7+uFpfHLSFDMHbe12wWaLMkKOxO+HSID5feqmxy7wqlPHmz1qkn9WGBnY1utVr0MHN+bsR
15ruvXUn4dvo67y2WVC00yCxI079NwQY6A78tdT+FSGrvAcgPVDQ8q3YjS0w1rC4p5cK80U6XCUT
VYJIk0wOv88in02yuK/Jay5au94VU3CrTVZhyIsyd7TwpV+S/2n279YGOv+TI+B3+PlK0fUpHhH1
sIQbXiW0oQFL4+e8nCAUv+uQU61WDqDwVqVm0dAqTFs2fwcqtTx4DTlwL2l3VUaR81x9/UmEHYKU
tVP2pEP8zptKb44U1cp7ewAXZGxf8+bJzu7NSJRuly+qR66M/vYbMkFSw+liqCu9FlXt9RmzanlQ
/RujFJUfhUzTDQaU6833GF2D+gRDAziWQzUNobo+gTX31yG3JbNW0yhNGbIANUkF+O4nET02Pb6c
e5+Jtl9iBnfkjFNR8CgMq/dRS4trh64mBVL8yXwsSQZr3tJYsI6B0OUXXsNgIUd1mPnGTGUvDRNb
R6Gz76lNsV5ESpuUjEqBzML8cc7hcnntNaxLGid9Lrgkcciuzznx+OQhw+g5mIozBVrWREosPwZA
R7s8vpV4TdHEhC4dlh/3ypU35l69KrCak29MwM/OXrBlZCgWDkwy3n3WBi0r6YzG+wN4naKuulY+
EWX+UC/WtH3Fenidd2bwuX0iWVBRxh8PnZlJMDyfTuPUopMCcfcV1p0J0kEqly5QSiogDcgUQh/S
sj8m4OR3tHeWHvSxknJHu9BuFW71Guf1tEiNti5j81BY/eLQmx5G7cL9JVJPFhJ1lUOZVYmJi6Q3
NNi8O405nendrTJ0MSQlLiy4VLNCAD5TbnQ3TIsr+4Ub22lClLLvKWc06iliLRW6RyIH1PgA2a36
5WQRJHMgA+a85kOPYK4UsuH+y94Ij3kvzj3mGKH6U6pKp1Pkg4WSVdVkkIRTFAG74n0vOcmCh80D
GSBMhldc2lEDSE+TTaO2TY2vhDY83E3oRkOhGyp8vc37lkSRwJEb1p2g8dwZH4imAaylMrjVn8/k
SpinHgGQ0hHVR26zbFT6y7D+jgDV8ndWayTqd9/LzXPa+8KGcHxThlnmmyzgeSS5Gih+4nUgYTy5
3JJko7gIymG+Q91AfRtE45gCjOu6GIvM6t5O4O1aEtTuiJ3OVXxqczZ2oIB6IICHXNeFTJautEPT
YlhURgHZCqHElVk60PIQogVRYfLL8LCAQmfbwN1McycAcOpxblsVjKxa7GhGQboHM0uO+w7OzLJv
u1mow5r9s53xk7cFs1F54OzsOq2fFJbn7HFmxtOcZqvUbmVJbHt0ja3u0FThkYUVnsxW/gEsYE7m
CRFOgRoU9bwNtOWPGyqt7y4WJaXoaK7f0JSfFjmbrrGbFDRwmMw/SWCrOp1Lf3spU2oUF0IcuidA
984pkgYQ2Tr9MkxG4umJ6Szs4Eg+1FrVD2ReaCFBK16jaDAMRaCW3s1yxo2t3jHVPLt4VhHWORf2
o50mfu2KyRayXKkhBwDAAPMYkD3/XtFWah2hWqiH4LNjUuX0zXrnDBZtt2pSVBE+bx+RPeirpNPZ
vIU/T0llFnu9NjBP3SU5/2BTOSqJI4570HrVt0HZqmY+bV0WTsMBZNsNS/gUgaC4+KjPHQuSrHmN
2Ts2hwk3wsayNB6PfM/OMOTYkjPsljBEcV2CVMQF5zEpjw6ljbwQWfA8yD0x/QNikwf5HMMpjEmZ
V1PSQM3Dawq2PKfcJ+lmRTw1dC9aMvg4V/+qwrzC5Rfgzf1nBemsb8iMV6pMgDLuI93P3MskrR02
/0rs8FrsORSUByZ20hRYQQUQUP24BtFZsFYQ90VSmZjU2FmznrTUIJNySxNwKbm1YjdIMiUgIeNL
jdcNBm56MIoBX6vvSTV4kjEPAa2NVhN/wJC6nkYhla9q/5auNKWvaTbTJg8E50ORLbPfUmRb6NCK
lfQCs+AFK6GGb9On/ilPr0WLiKK1yMBZaVPkKqWuUyl6c/8cYBo4Jcjf1Qikhd2K16bGhy8lwXGF
ynZvHAEbG6njfuUh2wBXVrbZlANB1vgYO7FShVi+HVtMEqoZgNgtmQQzchR+eCgDkygC0ieClkix
P0aw/0DM4Dpm3B+at9xZiLvs3/EAvVG2PKgT4HVh/SViwOFh4W8j6MpMPhvqXVwrsZF83vs6qtL5
elofAIdcXj+nt7Bq0eNXC15u56uK5uUx0VWfeWMD3l/hF2kI7DuxowObf31w1fb1h2p3LmmvUoTT
gDpnK+uB6LL+QA8dqsSa+UhsVco88MVDya9Gv22wk8QAM+//x3HC97vOn3veXt8s1cN7WX8ckjqA
Q7+K33Ey1GF0B0DcjbJRlk8kqQtGLhKKRhGaPPfLi960AsBHWNdqNJ6uFcbhbihGNbPVysaVzliy
vHbnf4e/x4lcPCu3I8S6N8b15cSl8KfNo6FKAayOLpItUJOV4zIbGcqbQv+RAsoE/bfFYNqbUCsx
gqyeKa+mgLtpIJKDVGFnGQcaBbOCV7FspQeGv0068Xmjdjj2YqIKiRMoz+6I0Dq3MEfwUGTxVdLJ
Ha1+/CkVdGNPu9PDcTmXrb2TgT+6FBdIKIBa5MbsQzc9wRNuIN0OQ41Td0bKBREhhS95Kw+rPnYO
skP5wpNV20mjfab23m7WkYOm2Oa6UV43pthA8cPdyMGBnf9AurDwua93u4yZM6np2rfpE8xWw9Oh
s23b5KzQAQudXImo2pYZsVKACTbqWWjCtveHYrtDTP441NN0zlRzeDe/JNhvpKheZsLtQZ0ubMyp
w6nuX4FaKrLUVcaxbs4twLrIdIkp0luAoUKYEJNbotnl0cLBi60F82hiilj5cbV1+FURO5ApMDQc
ihvDo9Gt2Wh8VlDLG6tA+ot86wfzXH+q3IsGnmWftTJUuRSdPxAiXX19gW4oQNnuN4hiCiJxjTEF
DBW2njCW2MF8CL+WYVBXjlH+FaLYacVZ1RrsjP4LZIzUyD0ISxxMtC7otsZw4tr3blndmuauaO0w
Eo1bWAwJRk10c+xnokttBZE3g/4alUeDcA5sVHK2fbOm9ElgJGy/d/7/q3dnrhSsEL9pqH/KDMVn
H4fcG1Z/8Aw6QIYSwz2gHpK4kep5GojrXnMSOO8kvCYqLkeMmKVxBc1dLqGjvFF/GKThkPZaofKX
5FCqqxbRwnBLI9P3a+bOAoVmveDl6EB8YoL/F8wq1GgO7jyI/ugmL9H3R14Ny8IA+yjAOEskorq1
osCRllYrRywbQC263qALkXJZSmy8KeoQil35sGk8HTUV+mhWMlwJwM7KuEF6BKgBWBG5run05Y7e
gWyKKRXz8mL9k2sUD+qG6xUxO3OhkTmZrCpsrgjy0sBb3Jrk7/by/rqvtj5yPi+v15+KqcrR69K6
zpq5AkP3IlNu9LG1t9ly0UFIyf1a3voju0G4KurYuxa1OjRwt11IaL/hM9PhbtC+fXkMv+GlO0A4
MjInrrxO4TELZaOMU/Lh3/AsGjIJ9u/nR5gtgIYwMBqbgTXlxybpIp4QY+7PZojWmrN0RcrdkI2a
lzz3e1iOzihTmySTdBvY8ydT26faNVLKWLA2TjTouLfcqJt1wavNbAUQWADAEbJF5dq+b+9bwWnS
5XZmz3dL66NCkPfbfGdGGQtbuHP4tlDiQ9ODOAJh8kvcYfILO1VjzEFNUwGm1emLFFOT1AbymgMd
PvRNC6e/XF2XIYCICBnpyzt9h+EZm69YK0D+3hCButz+jAdoB3KUYELkFRp5RsRH0c2VWPX8D8Qa
wOjlnQ4OPlD40DlnItuECjGnpnFe58tW6oRRSy4nsLDbYfNXD17iBKQ2sQcfp3+O1t5YgNC5NFyk
I5vpUvaDd9w7pTucpzI6XZAs/FfNb9A5rKBT0gO1E+OH0dIWOJwSdHdugsEawJWqV7HpG9r1/kId
Fz8J4m8US4ZiaVHfmvUEBxQrj5yxiQOAe3SC1kQmJJ9u8G+2A/OkW3dHBWBU9WqpZYmFyz/OEF/t
5hOoTjnyxXQ/xbNVj/AgzPo582jG4q24LU/SkJ/EThOIKYcfWsKLN7fKpHlJEbxp1s0IL7i1VVq/
j8r4q3k/O8uuO9PJGTAnmxP5kTdgeAnwsh+gCZwi/fZckZ/GHo/GPGVW6g2X+q8AcuOWusEWE21p
ubddc/WUsgFHz8oi3GYRGCchR7xIlGQIT/62Chb0CAUKSXAzalvF+3ylWrTrVk8kVKHt2FT4MjIC
JHJg1kX8Erf4dHdA/D7e2TWvZOF4jUixZUynjztDdppD4585b5hwYS/9+aGiHfg5bsAcaUxgj7Yg
cc2XcD53qfyIuZDar08HlbTWOyvlFBXFtE5rdpH7cMJRzLgPcgxm4220IUwlzcenTA3oHVocl8qP
D/PNEOGswyCqW2LFeAOcqHstfLRASADdn5rN5KdMG994gJsI6HA+vJH0Kt+I2cBg6feHsWuzwKfQ
3TLh5QkP88yDS7EJuvg7dHCeV9G1IM8Qij1Dv+O7oxK7B9Z0etuI7GkaSeVpLlq742/OXxX0IRvK
4+KYehLxyO2ls2KJ7Ak7vnydQh/5B9txl8Cc1D6NpEym0dU9Xpxs401G8Srg39lQdjhSw+hi4xr9
edrnktoc5DTMJSxfpfaf/3zNs83lAggaViIklPq5QPD223BTv+doEsRXXCghdnQLb8yHL1iNvp1J
QfOCZlj0NBVLFFFxDNnb+lRiekSIIoie4vD4+W4MqGlJx/my9I9O1lLUXDrz7+xz+f7w1RGKFFkj
vQAhUUh5zSdgDzeDQOH127oMGGU9ifTDIVyJpQ7VxK/foPwaEuhdMpoMTx4gSgB+tpqiUA1DSsUf
NztmOT67jUCIkDj8TCcRGiTglBCozuWbNiLfZVsEGkknyt2zQ/Ga/819lRDKnh0kZPB4fTnG1jqn
wtt2HM8LFns81tpQJ3zycP47u6bvI6BwBTmZCgaXLojC1k7y1ff+hORNDogep6/cMmF0ZN9LbFFp
SFfQz7BbHUNJUxW52VeWMoZ3jqgJC6CGB4yLgO44nKbd/j4ppdYYTqaPvIkNllz8Pj6Du8c/YWUh
VFIcO0lpAc3aTA8C9it5JStbmQTJsvm7O2uoCtfCA2TKJsSrOgLVPys/ra4IiHTpfNNQyg1b8vKi
w6dJehPx9CekJDcDQYr37j3jQ5FcjA6O7WAyvNl3pgunaDo3QJ71gXjfxEPctPXDtfl9yX5KG2OV
Q1WYDYsfrnZOFD8NO3UsbY1qsPdHaNRu40vk1djHtCeu5EhCd5DKJcW49ijkEuGsc96Ky0KyCNYt
TSq68gKwf0Ik1jjuvweLeqYiGd7++N+iFp3JX0b9pFp7wf7nUgyCe5d1fnX5HUQPnQK7EehPYmmG
5N8nn0Dsg5aF2orsNpP9NbvyK/jtNAmKVRxTldgOpaEIOgiog9wLn0JJWQIw39Un49wwj1eS9De+
yn/JzFzutRee3+6mpBJCfc7DZcMWkCFb5dffqPwidzTeZyxidr1aWKGQTZrQd6rw0HM6j21aDJEv
/ZUO6cNKCkW7hW4bqhz2n/XBxsHNW5lwwJ9EvH/SOBizo/27bDapRJKCp4+mIva8I550AwZBbIj/
yyGKG1A00rxLP5vQXgBpLXBI4Y8KN+l/xZXbakQi61RYvGQzXtQwlPfqFgaTSXKd3/OikYsNyNXY
EUzFly8nzdZP85AnSFZwMYphlHs+A67p3EgA+h/Bxz0DVNTAb8EfbvbW1t5kzr/DHJw/14NoD1bJ
3ycz3JCS9DlbIcbZR4iS/ViQGpLe+GyISYrtfvMZr354LRAmsd+dpvj8r8WKgdgDIqCo+SHyZNvn
UWN3eBzcTvUUgX7m23r3qmWXinLs8VwPvzyM1Pm4Cn4W6WHYmuA3hsghaR4S6vPLP7Zqp49Jl2C8
8o/hYEfeF3wxXHscitqf9ttzCeAi3yQ1WnRdq+cKvPRToJyYJ2q9WQ9wvCH8L6iLvW0eWKAQ4O4m
Tv2oMXjCBEOHPlBzSJoua/kSUSVJMPPEUX6HzHN7AttrP6XptUtFK6aI53mHR9T3nSSke9PkI1k/
Qd+nEFfVbC2SAzMgpycPpLbBKct1e9kOoaNXloiVfw4WhiQ2k763dqkTvIQ62TfOhQScbQCdTIzX
9yHSdK7LJaLjMbROZXtrbGY+V0geN+b0yx7AmpYJt78bMChWsTnE9SnQi7EJDvwzYExtmaw/Z0Rj
t10WRyvOJ/sJbmCUUy3DWHx1Qe0EEXnivubxLGTSs8Ox310oK9U25LVdrgT9fbexTcSCOQ8RIzUI
nKuZ4ny4r1ZE87IUgYi1Yr+fPPlLSZz+JxY5DOtGVjPLyRDt0kJgA1iW/L56N5nR/rXod/zmoTpS
2fooeqQGIjKG4vJT2toThdjarnRVOwsPhuBSfeH+cEAp9tqCRQFEumy/O/dRMHTyRR75/HYfkU/5
9GHkf5PgUHPseig5Hkoo5GlWpXteTrYJgbiRiRMeAVDl8ynWmt2iI24N9giEcTA8BfpagN+jFfvO
UDS12CyVMAcOWgpHFlCba4DzsFSPyVLNjNRcNe/hDw912fE4iK+xsvl1lASn5cQgH78sc7MHCxps
kKeWdC8t5zswPCKOgWcZATt9Qcf3VFgcmRWfoInfYYXO5HUAxrgCyzA1LneLdosu1Wcc15DqPv+6
wnOejzYqCVwhYmUq/hpIaejuCrgyjx8spXT4s44tSx3uA5An/TMaX1M3xWssDMOmLVjfF9U1Bdck
3lpWA3k4CWhCRTXgu5N3wOlHncw6LzOXCLT21gT08omiAOFC2TEJyjvRemtfjcXxYIdPsfUE7h3O
s8BLukvAX8xDux2B/30AXlY4p6djG8TBO+ZVov9w/Gxy7TnqU5+0vVJr/tsRKMlseECNIxzQHC0/
J9lW30shfoN4dhT+8GMi2ZRaVvKIZfpoQv/WkTWNCG9KmuLVcH/zIRNSjS9PCfls8D3HBQt4GmM4
4unb/UfxQZd6DojlbogtVOKkEiNe6Ix39iGIW6nHUR1zQibzgwUrSuiCqJ3Y/qzrD3Ln6OqJBSZO
DzNHTBdjOTHyzPab0hmUD93uy/vPrj7BPD+W9pBCMtMFJynWftj/VM8LXvCvePZiGzJTWOsjWdm2
ADh/sJIKwWTmhv6vpdD3zkF35mQ3ysqBCDCq08WF0ElJaoiASCzR+HUdZKxq496k6o+rufmKeSEZ
3y1MZkwpSvb5/Xb0XM+Z7und7ZcvaOs0zyWmmKewFdZd6e20XAdIX+GNC/vjSMCm0bLLqZYG2cAS
+qvoeMcVPk82oPp7ay6uobTHM1E6M64nMepTz5ENjknbk/RaMd5NivBEMblxxQexGV43TJWJAFgV
H7sZPZoZoRx8wnwqgu/inxaEwDh5iAYpS2Q2e9nLcBvkcqev47rnW4sXCKanMWLWATJeSoL1r5cb
l+cg9gDLPVQKS6JirAP35EoEVjlSeTnMHk03xiXmnI+p84s3c7RhcH+MUBj4wDkyXqyLu8xUof+H
PH6FexCmfxWtceAsDLuHA9k2KSr7a0lc3+Ke9CNJHgWTw4T5N/EdP6e4bXbnR9pwfHVXppIE2tFt
ZvxJpbo3bR/MwygQUbnJm5QYGe0tgnmez1AecvJ6UN6jDXVbOZPBghGqXcD+43xDZBtDjXye8jDa
0lIGF/l8JQwudv8r/1B/ddV1H6ASYrGC1lCsmnVpX4YyQohb4a1T7/O7OydW7+Jope6v8ZqiK4+5
BrxsLFyjI69AclnBBYtpwdHqJRvNasCoGpOymjidjpeQLTRNtXYW3ojjrIf0D1Jg1SzDkFcWnoCT
mYjd2zviy0prg8kVs2Lwy+kLnQ/Dcr2E4W6VwykKxFSAC8CFBdde4tfTWcjEFmOSQITTUUXkgml8
cwQ5OAtlwq981Xw6Fprk7nHdl8zlR98fcMMHRheEc3sdUHokr/CpU5+wBtHyDUq7bz96IWQqCCMn
u/FeC7LjgIVEahk/ll74GBnM+P8ZV3zHFbriQFbnA9Okx8l7MNLCtmgPYqLj59l5iR7MdpcCvmJP
NU/uVx/2w5l9J6G2c7PeosGPtm4dlVnSGxcXDI6RADMcipm1BlejQMf+LQWN7VQuw6+t6UDJYxDR
uGU9dq2NirVhX7o2h+sg+1osYStdsdKTLw1467LIWRTZTvjpVuuCzW7McoihbfYFVVZraMBp29rm
7S/NMmAaQIbo9DbepPhSOiOWdOHd3hGbIuqZgAPo63y/bxWYlEvI14iLffuUnr9+kPO42JK0U185
Mbxu6LCsRQ2dxVLBeNvSDgDWIUHiwlPbIbsSNjyCbUuGnfPO/jSAE4+erviG3STvpDLFWYZJxonU
CI94s1N2nloTy4qEBZGxoS+0wFJ3DSxcj23vUvAR2R3X4yO2EiFhgvWwp3dcaKo+2DaVF8ylJBup
X5QqR322qIyYycw5ehZcWelmzRJM1duQlKhIpjmutBnyK7HK0cXMf1Vm7y5CVqEz6/34haAF/F7u
BOFeuh+Ru58PQgGODRdWd4KQb5rP2RJj/XQNGwg6hWiBkRMH6Cur7FJDxK3+PSqCJN34eERCCMwK
wJc3KZqu5W9jDSIpUpKtyWVUWU6oPvXtwf9VduC9xmByzBm5NQ969mPvuIi/YtuaS+YJPSX1rkII
LzYQV2G6TIqyklGOyE6z8WNr/+q8qaNr7E+yWSq7xe06r38QYsfuwrPodlruYm4GJB9wcUymOfZU
VKznE/kHdj6zHZ7sf/EicRHB0UTwKDVrCo6p6pkX1suGff31XUBSM1EWEpXGUUj1K0MYUbQXpiAl
22bthRdwTY9r0engHVhPgsBS+MEWJTT0BKeZcD+OXxc/GZjwACNOOUg5fShrv+FoyFddUc+vN3iy
PGu6t+IaJLLO9N7ErkUSo68k6ekHA0PFaNGp8fU5Cp1IHV99zUu8yMC7KO5GrJk6ZEN2Rb8pTC1s
ZZO+s/f5zHTxv1yhNZSuj/AmpicPQ1pkohos7djM0iIV0C8j5GpdUXoHMjMOkFh8q3nkC4KODRCG
uBNZRm2ay3ex4gUn8KwrmP0pCFdL/Rsbh7rR48s8ErY6TGYhPsux72tB542nl5z0lAo1Dyd/CrQD
bmU8IHdZTdRbO1J1ihbL4MyFgbNSWo7DW8fUcKgNWPmj0XAvJqYBeir7VvVb3Jypogc+FQMAHwTt
jqXbRh/UtveHj8OfVlYhc24Tagxc2b8NdnBTbVFeuNHH9/suOdbDHA6+Mdb+8wYXr2/7e7bY3Orf
sHJBCh9g/itO58Xkoo+IS5gaJgosnQZD7bdc7nxGcKzczACuI3VUUvhPycvnQkdgxReIl7F0eudF
0LRKq3J15drHd8eAq7Ifw+kxwNbb3U/EQ0LqVKL1UXFWQeOPge6KhHq1cD0dTSeM+MWH+rmYvw5z
MdgRQkwEf5gHJEWEOiTaongcDcH8y4B1pbpFALyTkbL0sxrceqMdAqbVWIWsZOaZt2jeb5dPOfN8
jueNLdVL8WE+WKmdSrGNE+oOssdRHcUQscfIoNAIOxr7ik4nMZaqE0NE8O/KyqICpZPZT5X7z12P
y+LSeNvCau0tTgXT232rD2k2DSFcTfzcoI0JXMj68DUVNt6AhqNk3igoZpr6PI4X0b5eQ67mpYTj
g4W7VkjFoow1Hmb+WVO9gko4ScNnWtz2VOFXkcROWS+1F4hXAGjRqdO72aeZP4Dm/qaaDvdC46z5
E9v/5O3zHoDsxXNyl03QLfFTcGDVEef5jcahH66gIrDwMtUZEzHXneMJcSkxD8t13oWHy9yYzEOV
4vVdGCVbc/0ipapKc4si1kWD68cSkH01FNVL847+1I/1MXEk36bRHuvcQhGwE3DmXLGRxMZeW62N
id5hIrYHjClcYY6KGvykJBg6w3OkD2JWn8wtSWjQq4E1GApsSrYLITtOLDThOlQR6afZ8tBy6TpD
iJ46YjHrLvE5rm67Nx7wIGyX6/rbB7ArUJsvyvwQn7ybBHB97vVEHpNcZdgWHxOIbvo0TRF5cJub
wBfPgBCXaQwNfM7N1Z97Fotc1avDgkHjbibvwTO7uSFrL4RGBpan8OOVKq9RQAND2f/t9WDBfzZD
nLQSdZEii4BTHhXbKvUC6NBbEE4rxuuayRx9uJv5XHxoksKq2Qdhh05NFGa4VuKtMuI/6rwKMnLY
LFVzEhinaIjh0m/84gNljRVoZRJ5nyzme6XSMLmIQTu2Pfl2DuxKikA0HAwAofgnOBatrBkjTtwP
/qu7O8FeCIQkicZCXmTlUemnA65X9AZT9Vw5YUfb65sPEeQCxNXnmgI8JoHJzjIYFsiwj25k0ezU
CDRogR7jA8oQx8kkpiq7GdHGt82d1ROnTCxVOUiykW5685XsBHdZV6nSM0IH/Wt5FYiGB0Kws1Jr
rWODVV0ju+6CxA/8JQp6W/j99ng9ADlQRG6jsyZWheYPuthPfw4HNP8SdIyMooM9ntOZKJ+EsN1i
FkHXpPV4YnU9rLm8LFC2eeYKQoNNkIqalSDAWavk1VrwuipVAlMzCymfOuGZHVam7gDwoSKDEdtB
vkX+ZOZOd/xNvjTb7dEuCuG79PUM+Ebr65IRry495CieGZqZMJOmVsWlK481JZaY5kvnnAeEJM4h
ZqbE+2RaOZAc31VtF2c60T6h6kBAGS29AouSiffy0ug2v5bH4vOStl/2DHdIaf5L8qS6RrJwkhlP
piujunNVQg8bYFw5tCcLWr4PC2V40Q6wWAZ22bUIW6EA6K6yV0fXapwZXXxDGnHBtuCeaufmPc6G
AmcKdAoRFk2tEtUgfZvwwYt2qVNBbow9LhkzcDgCQ+J2x1bHsUkb/v6KlzDexqAuonmnv2zVO4Bx
XN8oU8N/25EORbRZut2XlaoQOoae/bLu7vrHaR9pxmWZnHpd7FPbzjgBnMPMlfgHZEI7EEvKiG8N
V5xcm5DcNBrYOAdySGOVWEIz+59p8n5DD/9O20XIzHUR+wD42z+RDmQRtpODBSCjQPnqAu7+Bj1A
y8MC9LogkQtN6Xv0iLXphDF8Pu5lrLDKYsKGmguBDw0vu7sZ8TKlzF18NPINwK4wXiH5KkL33aVa
y8JgGcS0rqzAdd1QqCUhPrDLxkLP/ACz9hTAuTCXrp/tR1NForUkH6bTo1GSFliwxfTLRP6c7J9y
u3f9QYwFmPari0YIF98742n4QAo+HXJtTf0Ps8D0srCS07o2DLH32jf3dHQ13rJ16o4m3fsbR2iS
zs0JVVrQ8xpC4lFOEUGcS6quLTFbGjtAiHBrnUlZRgyLqhPdRuXdw2YYcZXXBnAQnj2Ar0SBBen3
BgqMnra8QN5Xulow4Xd8q6S7k9IE3SiBMZueMuYm5UuHG/ZZuxDxQDfdmu00NxE+Ar1Ic+PRyo+8
aarDJLomw8696VMfRCTI45E/BGEg1xEW49r9H2awjV/BoOtK/BC/LEnnPAOj2tZp+go3EnXIssMo
wCITl3fT1XdAD6kQesGqQzSFsJNUB+JDQ23zRSotNRShGkPf15H50fu5aqGiajclTYhE0ZhsBvSJ
E4eqRR3wrLhU1oJ9c76jIFHsnatKaoHciT539CewEfqlGxOF8+hHVQXNmfV+YtN328FNzW0qEq63
EyHYIjuv3u+PbitbuEHq1PFdumVg1hE9qexqhC5bSWvULwk6B9lVLlIrMEoHECzLECl66GT2SAgF
JyEfhRJbMXrHFlaBedgp+wr3e1scsmEv68072dAKz1L/nCMyC2oatnSVH44UqgGVJPimsLSRnj+Q
1C1APqUfUBjIZ7XCTleNWYGXoWifdAFAi02zuPBIEVVv+2BmeOaxsizSkdKzvWKWaJsfj7uDQ2yY
UpMvm9H2bIO+nDwyXj32LDF7DMz7Q9N0UxuNvkM6JHfH0rpDuqHEgBoDXKyZre5Wgk63sUWqFOMI
q17fzKjXVDwdm8gOkKEOWvGR+pY7pJ1BnL7uFhMrgEkDqwUNVrZ5O9494H504P4OyU4Y53ONS6UV
GYtovi770+ktybdAElB33+vdqUpw4n6AVIqbp6HT3wjwjj4DvYmdGEtmjoiIS1ckzxaoYT2EWZYZ
rvMDnjf+IQDxwmgRRa0jfPYRWXzH7s1X29LaUAghqEaaFHrjKrypBWfT1U1mfhOcjS4RE3cJjHgp
YBolB5yVDBAjjDJKKm5GIM479quwP282CvhRbQnl6mnrqnxJ0PoZNnYomSAp+1WGrsinzVfSc2x4
3aK6ioj1mzcrR/vbAvBgIEIbCAixy7jldJvLw3QHTOfmkAScpA8qX7WZnqI0rxCpqnaTzDAhZQBU
uLFZgEtzDLYq1KzfzgRnqaw1sZ2Hd2y6Xwq13uz0BDZnQZ4LUd3+LRq1Q5FIPmR+JBqRIktqDcsP
HzRvvalRc2O4Zzh0vVkZjoWBi2+C+Zy8CG2Ds5ibnqUNZt+cS6107dX7+KYbquN9ZMWhRgyjvM7X
DdF6ebXQgJgSwZJnOF7/MG9nihT5wEiDMH+OWtravZdV1sEDDq3JCUAzP5ruvmweufLWbNPDmNgQ
F/+kaZs8iFT3SkuqdO1MJt2oU3lIhVmDBTSGb7upmSLMEb/xa0mWcsO6tohVBJUv7QXSIwPbeM+d
IWAaBELsSnh3h8p4mv2BevXFhRxpqO/jJ/mLk4S9Q53h14UMTlFw+VneFDVXIpo1XPe/5vox2Cei
Oq0josfAwJQen+tC7D9smxIP7ujs2PIFvHRY0/OvHhlExMjc5qQd6O5/M8aG9TacY/4/AS6EZ7ab
imIB8Zez09gQuDhE85LmYTcc72bbNk4sUHRmvVNwW/s3po/liEKEOJQY+oKO79Z5beZV4i2+u0Po
Fscz6E1vCRrZ6FPstetCka2XP/WF3nir1m6z9xYGh5cSFuG2xspjsk9nAyY+RzHLouMcXJz7DigJ
a4pxhEnaZiwlXDiGXhyu/QkxrZy328C83FJhoXhLATGJgVEHwO+zhz9qF9i99hF3DbAWnLWJETtC
l0PNr5Dab4WTL8CPLIO4vboTeQjc5l1dATs4maY1SQapuCot2mHBCrjrJyP0eeiH7ZwR+F/DvT6C
aU8gx/EuLN1CvxjW7CdIAZaPC/IQAPs1u/O9hs/ChK3led6gZ8nUtNoQ3shtAVQmqUpzE90l3Dcu
EwY1hEZChDoBWPlIqZrbJ7SZMyt1tues+qUUQ1sz/2Vesz2vnaKJsFJO6ZGDIZN2SMiuySEDOzU6
tpRY50OCoN+HDqGleCPdGmkO2ofvsVUuhCe8XYAnoW4ocwXigqoSnYXV0jNgt/Ak83B+L/JuA54N
5MC2haV9TLh5VicWD5eMJCnM6z0iFaTXxRowmTfTev8bhOzfcyxNC98L54suwwvNxDuf3u4AXb3q
FHXMCtbtInWMhiHu32pYO3d8wzv3yqER6l1o7wUTi3cLvmIDJ6T2MJxaDZNB1TEAm7HNk21BQugF
2C5Zwa3ehJdNEV7GdEJln/moseKOs61ZOsq3WLbNYjvJxkXF4hKzNrOtPO1MwYDFyUfbnJE45CtE
jTsu+gmrNa+y171N9Rmqm3PyTJYjzalXlJRYEA6a+tEPejvwCrKw6aYQLz3Ie6QihOTDlHQyUl78
eXJ/cP2K7up+vgn43+DEU+XFss8Z1QjZ/cevi70vZOUQ8H8LQdO6opE+6ncIZW/goK7UfmzFfmc2
ULWhkfMu9GgeW6cfC+ewUBRvi44wxU+xYoKk/a5gnHibjbzHMK/qqTqMc8/ip0W6u7M7QpyMTPTz
y6ezRaRyl0Zb3LdVTTpII27y0z/qy9hn3YjihF4O8VfXLEdHxYRQ+mEeo4d6tC67k1IiipctWrg+
c83bNhhd1mFePtx3DHHVwXyMWyKkBHEyrvJfiezoDbaFFYvQ4HnLb9RFQrolLgD5Kk3o7hMnbUgx
Hc48PfGe24u6mm1EQXNreqqDjHjhfppIQkcIxmDaApRA0QnE8HVo62+gNIVaun5u6L3LW/1IT8Ck
hzq4pmK/bnPNjQgolKL1NxHEkFB0p5Ym0dpvzkZCoK9/J/ffQ7n8UhGAXbr0F96mTDHyslR5JeR7
sv/IF8C/8vW3r/Jrzhe8T+ypreiZIRvYPLacYmXxolqJrh7C1HNLxHi6HxjOCMnfgYd6ov2m0I9m
E7G9m7x8Z5Ch9gh9X3chNFd/oqrcTOO70C7QfjMQqbQnTba+/FT+fGBQXEFIrpELh0fH++9y8GA7
AmxOawCHkV4ftgPyP3MZ+VK2ANt2kQzIaTJ76Ast+Lum/OnevP8SlZcZv7r/Tq441aWW5+Heo17p
SvlFR/TIPhU1kNccSj3DlY4wHwaX9u8C90nzfrk999p2bAEIVIOJdLvZqMCMgS3vgr5bJvs+BF/H
/xbLhiT7w9NSTx+tCzfTzaRCGWt0oiqz5LUrdTI8UcFmOFkCHdFJnjda2VP7GNmpCCdkUS5dGmPG
qjTyOlKGs28IfcKIKN+GxbRjd2GqfdXM93J79BKfDkheM/nkD45mBRvadBr+eD43m4Zu1J4Erz+F
7zS5fDaTYlEUH7QZ2VAaGQLhMoOIqHbhKk3ZVq8WGNQwHMHymxlDylDeBVo1YndFs6aRFze2npDN
0VGR7TXEtxvmnU08REAzGEBIB0DD+uhpUNaXmT4WncGMPvM5vm12z7PFo0DLQ191WERVP9600KqM
gPIyYVZeFQxDVjAnai07ymkeVmnWDiTfQRPb4P5YnusnPYOWzR397jt30hYL34Od32dINfNWD3fo
7dP9tuKcwFOf9Xx92LGafKiw/ag69tjirD23yNLXruwYozJoesK5jqVsxgMRpz61oR9xBstX8q+2
p0s2Mfi7D/QeRUymZq5gMVncWY/85vdZ50XQV5MoE1fs5a8c/U8eVBUgqgqWN5C1wRMQyw2ChrZP
X8Y+U8DWAU/JnZwkJ/nzkRwLF1sJcawp5puNdRppdOeDJy56q1LpvG4t02Ug4k4fQl7vEY/Of0cj
8gdQcNB9/PdL+MVvIhRtqZfwq6wVvOStLAtZScUr9hNzevH1J57KSH8TGaLMiYT+V7+gXi5y1xLx
+GuiIueMcKYqOoTdxvG32zVzvSD8ZUwDcbYSw9IRaQr949vQTNnA6jMc98twozt5sA2EEFc2EC/9
doMwhgD/uGTWaJ/lYhzTU5gjMunqjxBK+Z7GO+VGlkGWEmhETyYOOInaA2B1+Z3rm+D38W8x1Zya
mKzPq+iyyfycH+UmAxsUZnaujh+07f2xgqplZv09elzdUWawL3OqOaAR6M+Vu5/tUs0aDRVIBDYl
P9iS+y6eeqaf3z4fWlWk8REM4ErYKe15UozkJHXpxocG2Zsk7aOBDOpJTipfa5wAqMBNefrpJrjv
xvogQrcnPHqXCL78HO13A6je0ZMiJA8/VTlXYlha3Wf1KDzLUila9GaWM0LuyHRHNdmGwkliWoIx
kMTHgG4a9FtaE+JPvaSX8139H5uCDk+6NLh+xaBQQ706zC2V0jJrxsgw2/elJAOZk+ydTSJq5WFg
Pc/20Ll0b5Xr4FwBczRzjVJpPesG0eVs6Wx5sOXSJ6SbAl3lFvnQFYNnINziuxRbQ2rXonYActd9
R/cygxh8EJ0duzvgNstIR0WqX1X0ui12uJdAVnHNJNqSsUAKgysxIm55kFTBOS2exEwDYLttzikW
H4Ouv2hWOaC8OfAvPCmIZf7rLb9H7zh8PAccsEYYSX+zG3hiQVxtlaHpHbp/IA4zb40/+zu7B9KP
ORLBYB8FZu/Bx4w+yyHkb1xb2mw7Qi+jK/2GgVw2LVWqtw64MIfCS8Zk4VHvE17SUt4jcWkp940N
9yv351+HrqolqTgmqDLax0MWDrxQku7hV/kHbzIUtG/HMcHIza7iXEbLq1OG1HJ/PROQMTxSHdCT
dM4N0asF78Ln6WaZpbAG3n6xdI0z1CgHIjVKa63q14t/XFuj/bDkdMKc2rMEZsj6mONeRRg36XTi
ouP26IzI07VTybhjxSiWluw6wdN0HNJywYrhdu/xR1HNZXe8/oEDKg0v8qmWc4T54BlXbczR4i0U
b9XCzRHBeuMWatX+TL42858qlZH572+1Z8jLZSmco29t84jyNfg0CsjQeuJS0uRHv6gSY/xIPKv/
c66aqooHGcAtnpRum3e9Nz9cmunZMr4MNgShU6mDETdqyhzRWTGPSB6bGWVbpZaGiD0YNkSRDUZT
OoYhdyLz52cU3Xn21DMDqrbuW/NZrXYO4ifHQVt/5AcSGPdQ6+FANQ9wggOgNjFpFp0EV/TcHm6R
cZivexYqoSUa0ebU/0GgSvxnugpoRoZsGyYyAii58w9JigIq2klKy5fLq4UteBm88Zr8yiphF5Dc
a5MHhMdvmE0MbCxfkB4YAkVWE2BzUMucxJ/ACk/scKlPFpIcZSGtc+yCsUCI8T3OhVuuyHjpbNpj
dr2sJPgKguJRbFV9C9ZzW9hs1h7HKwZE86I3+ilAPqKNXJFDiZ7ADiro/dcdjrbg6gDWUcO+kXO8
38lzRfj/3T4ETNKrewFeSHLdS8Uhbyn0ymcSgndLcIHUCfRzX/NIfpiozKcMJnKuOF18zNvwzGKj
rTCruan0qrEsjhmSAWc9JTtxsgX+VOEeq6Z+U0m/AFokdg+dkjuB6jT+e2pvKLrQ3YQWFknu1k2f
ZXtRqQJxljkqqRtZ3OE2DTlGDnGvNh+6xFHggAwnI3okjtU4GfQbwM3+wIV8uViRlan4k3jAy1S+
/1rSeAi3sxqehdivXmL0g0zhlI2xl7wsKpu1m8dBpSsN58X+sBUSzncbM3mBvfjBWw5ycivPtRzU
JJIKE0oA6NmIa0GLruZkXwBojcHLOXavMmVg8qOv1ckJzuDFgmapeVZQlbAEhLZd5iySy214Ub7U
AQrgpkeC69fsOCYgnxGrav+NGBHOL5wKRkuzXNNqrQXcYJcgSeAB473trr55U3hI8z1bjG2RUbZT
4eD2sngVpbchs5MUo5Jgubcq3P2cHXKXBhAzZh6/ZDHgYCS69QZsBfJbdA9HS9ZIuAwfBglSbV7x
syGxqS+jZuHcTIQm8YWM+UHaw256dPwKJGAgSy3yVgZ0GPdiblQQxqnUmOsukf6c6+w1iEM2es+L
xrESWVs+69A6Dp1yJXVSkbLrQAiNEluiEJkMUBAnTn/G3U1VvHwh7dI3G6coI+nXJ/6JS1qcP5ee
oOOsnd9rnoQv3Ju0DMiP4caINMyC1xAskfeuJCKRuKzLvJadakBSit5wcvCcE3h+G/ChHzPuup0q
WaF41YmI3bZBxrm0q0OAVybK5LhjpxR9p3juRmZ57iRj7flkt7jRrzCp8Bgh26RiHdmftvfBSQLL
pEQW+uxG3iDTC5U0hUlrWXQi9zI/ALsrpV1QVu53FHJR2j90oxsgrUbSJ15P156wXXk8GAj/k10R
8I1pYPknT0I/j35QyCNrcu+q7H5qJ8IdZyJfl4JP7vN14iOdHZreFOkBn9zIEvD7t2UqCBdP/lC7
vwHXq+cpJhdzSMGjvgLZnpGnWMN+QcPlmpNhSCPr0qT12CZFyYKcKwkvkaCAbshs/btWR41BL0Te
fYo14v2N06NwdcFsGHxicvBaJxiqCfB7oyobzikpsKKPChyL835LROaURDvYa2LPnxzUI+C2SUIg
P+BpJ0BRZ2hM/Y+Td+Qx1cw8iCDHBrZG2sXQfWDf0c+d6PvuiuvxIxPciG0YQK6vznuWrmT0Qymw
BpUW+lypKaXwqqWFdiELYCNAYDzRzDh3jMn6dCnsTC7FWXhrSyzx8fJlLPguqtWha+OnMxCOklOk
3soJ0uShn19U0+egL7jkA9GWEOX9dm1bRuaZ3H0M9RQu2CRWL9F0OD3PRVE1NNkR55ERiYk7j41M
ng3DGoFx/rFu8bd7P9tR38+K5TWhkIi7dz1chtt8T64V4PONbKj9MMIC30Ry5XBHeXPqzcq5b2jF
WASVEis3M9mQ3FWtC1tGjJHKmDn42CHbjW5kDHMTDOfHjpAFVCVefJ0nLQN0GtTLPR+j9hZu3iFG
+5JKnZDVAE15RkU9yJsoTV9+16tbZKXvd5dUpaTYjowl0ZYUzks23LPCPsfRfbQWrH0L74zvAE4Z
hdrCdwllQdW8yNc7KO0lgZsuDUL1EN/8I6pyNeG7ZULi73K+rdUPPd4koibRn8acDyPzuRHIvPxP
QlUkehDnn0MLqeXKPxl7da1ZTEl4VQcZr/XOJ1X+/s1DBXw2QWTcqj+K30meNAMn9NfCOH56Lbzb
YeX/KEwY8L5XBg6iVGwfzULiT6IFE5bK+G2jyhyqRbXm8+GYCLWx7kIebiVh6qPqZGQeMBhFLRVw
ZgcXrg6LwPvM+i6bLbyl/jDn7FGLydyXmU5CQ7Gx3ltLZnleEfuaQ7aaWDaFhVLGapZTygifgHW9
NpBOrHPHvTlpZ+2lB5MxQ/AsfyHkE5H+2LE07juPhdYII0sNkCjelwTa5U1yZ1D89Nk8GLCpCMv7
p9+1BOse/4Kq2Rv54MFjNHJFcXZ30qZ9RquIjOzEKfOt729qb2TLGvMvLmTnHtTFcYIRtcO+Oz0c
FeWqkhF4vVxoxBPaXKCwZM2wqq+oKnz3DLivchI/WvzvpKNO7lcZC7Px8ZN6nxYxyk6GX49miDSp
kEJwUIRWK9woLLU3R/82uht0CaNXFXcyYXEmUtN88+crEqhJ/hd9ulr3iRok3U0+968UoP6ZuDbD
jNpzU4OMecOSodtDatBRTgBm2JvOtjHUgTXJATu3+jQQyfzvDTsAduUYQnUCgnQ+8fB+0edaO57N
hpONxZM7l9+kguR9uqNXZXmpqzT3p5F9VoM5Eb34zgLyegZ/PwQnytD0QtrwaomlCpdjPisM+jFR
zgmqhHq+bMxIiExw3W/3CmhRleeLDW8LdH+aumGf9zXKb+jyJmEm2iO7glR4n28IhkFF2EFCezWW
Is6gc3wpjVttqIsB4LTdwXnHs9YSE8ZjC2CHIKNeAKJC3cyi7oTFMBLQHFnQbrGPKpflmT+hZ2KO
039jhAQiq1lZul6j930yf4je6mWVYVkeS5GmKbh57Bj0G4QPwfm4ClIJeu4kupvv07NyeGyYAgXS
zyzALujLyVE2pte5QJP3f7czh4JkAxKDOCpPxbqAhmuBZmdnbdtIahUo+iL8fqOTj2vfpFcwenUr
1QcUYyJg4/gNs8EAl+XsD0hGP53ldx6TtGC2dUDYC2AmJTXxyQ4Yn+hpgC/RPz7eznV7dvpZ3At8
tBUK7u0CfAc4+96H/bvmjAVHzj0Al64D9gO5718DxIcHLyw0tQj/QX1qi7/AHmWYIfiZKfOhYz/f
yRlU3rzkuh3bZU8F4wRpdIAqgDDMvVKqeM6c/xYyULIOnVxiiNu8vV7yxIQI753rZ3LeXr3V18Ut
HhUM07uevApjUD1JqB7CBlmVxhwUvjBHJRx3iiw+669MxUMCE4M155BZu5Aw5NcvUdLSUN+GAYYW
nNtaXRaYVULbkIvok9ywyTbQzm6HbQzj9fKACqw4EoDSOsQBa/NpvadMvKULDtAkvQx5NaFCHf01
ZcX6dYC2UPGHFezLDsPNqH66hlI07qhRt20PNeql9lVJ84bCFKEP4OLT/MkcsJx1s+4TD9jL10zF
5zEn0VLs6hJF8XR+tR5hRukGCL/WSshhZHI6FhvxvnjUHSRgh4BNnkYIznFX5MRs+6/yFIi/I8JJ
PVtRa3/Y+KX3j4mXfCrX2PHrF/Yf8nKvGtMASl6Y93i8gi89LJ5E7OPAuNft1ak/CvhGFhWvn7VI
GcCV1p6jlXzhNsZpeNQ9eEwGJaoBKU66r87hkhGD+2rDGYUDdMhlLqIVy40dirYrhZembk6WgX/f
BiVj5AlSKQHoDtiVQ4XZdeTVbI12KhzusTqhMQFeEu5jLG9NeNAg74AZoTbNSToA4VtRHLCkduyA
k5koSkCYKEQov0LWRuQAozhYDoqOuh4DfAFOKFHoRam0/BUtsbW/m53EZy1ApYf2hbxT6TCBWErO
if/audRph2XdxeatWYdIrlQKMIk56WfBVOCz4ShD4Xv1JC6SKHywK8uEzrbnHfaBf9Agh21O1GxN
1IQkb5cfX46WpO2uoRohErCSNwlrE/ktiyY8mmHWB4FO5/4LHtN+bANYjuFd2MMvhOmExUoMJZ/r
Xe4heunYk4XSlh7nJpMrs3YD8FtaPdnOYplPn2D6JMts/SZKFJjcrSi3Li7yRa1uFM+kIScqTIfu
ilOIJD3amOsN4Gf3mpBJHAdVItWCqQWFYnm5V2CFrIDqrXZrA46Nq2OrfmCsr7RACMJPv+rZ5iJJ
meR/s1urr5J8EHz7iZCvjbxxA6xNOhJKWGWBDHoGStQK/jVcr80oF8Ekh1G6HUSUqsfArV87kifw
tkS7XYxOx7DdBWyAs63QABp4qKmTUEazuYYLTkYWqRb0XjrFRFLe0tXCSybQ+2GWwj4yQi9MOnXJ
ca9MWK6vsJY1fBfxefoLj9uHgnf5hHj7uBRGRIPfcT9QiEH+9bH/2hFnGg7HuTnins6IsdwuNPZJ
Vzt8R0dXlaOVQlLcRKDmtyTn6wC5lh4M6AoLbNOqa7agvcOimOXjWfXna6JTZRU6qbALx5V+krof
EDOJjPTovtDcFBnfhIkCpGF0SjX/JZ6u3CP6pZIFJR5eqRqLY7mddfBl5FNixBL/s/+JlsAUXMq+
RTyuPwcLirFSXrbVmr5fssw4D/GaiCViWrlqN29QrSLtTzXMKjXbSQfmgyAnU2Wq/5v8DhT/8sI2
1610209QybdVvK8RbBTO8z5w140DRF+NLw6rjxVNzErUwH2to0MDrU+DdhFmf8oOK1uKSZor7HMW
s6WJikqJMYkscIEE4Ipw23SiD+SZEbuA8T8kdSEO0InxaxF0CSrKoBY0CKU8+3DPYAIT/KyV7DTr
jtmg2J0DAvBh4vxqiR0oXKDr+MY50BSmlKxbQ/s7cZVce25raDK+9Sc/XY1uI0+Hj4qXOXFJn8vu
xjxSuUZSt1Xl7Zg4fahnMEvPOW/aGyQAfVZGtujrJaZg3Qy+Gt1jeVvhORxqKevxsJKQwDS+6AKz
jhG7oNW0N+mqr6nYfI8eUjmHdNsaErPROBSF5B1QI5+L4+5zgz5qtbL9ZpOdFX+VbEMcC6p/KKLU
ZrboIudQLSYmBZa9JGmOjb3rFBah6AYKsavc3fLW2sv+n3xymLd5/+fwEDP99kXD2mGuRP9o+Pck
csrmJCuqW1HCbvqYkbFBw6P6WeK/8/Im1a18I/lHyKSRO/JH2TCY7LXCcMF5Js7DvHIKOA/9psLv
svfcmybk4Hob1s11wa/3R9vol7/uiJw+pC6C7UYMI1uh4bIjw53PulNJZdcOwPH3UNl0rX+amtq3
0kbRwZwUq1CLHB09shbGTd/jcYycBlkpTay2jgbyjc4ntefGOnY695GdmsSZLQECOR7B52dS361d
PCcgFGwgr1+BnqrGYUfzUSkuUr7wc3k0+eWK+XU638dikPSYJqc69qrf0kIDq2UjI1yJ+9r2SLL3
gm8LT/8osB/Dp6z/EYZueY0ZCc1CvSwEBcV/Ymaw0pIDxpc2s+vReiLJKLgFTwtvHsMVMKM+l2PH
76tOxiC+s8yS509PR/A95jhSYkr+/jUqmkqcOglnY+k8celBUWE6KA0TiN2mD5w3ESV6Nz32kZxA
/zbdr7UWJjOkL0yFiEV/C2LaYve+0dBdntNdOO/+OnY/fhfmK7Zt0eIxIYciscHsAIW5vTSKJmd0
znqlJ2SdJiscKDKYFSv39H28PvVWHoXD3rmlWxT3BhCgK7TfJcdI+kTgy3ZJGYU1LhRRh6q6QPz/
/KjfYi+Srn7VY1QKrngm5fQpm2CwWrZuSvt1PEi0fiVoUWTHMVaaAEC3YZ9rw3oNF1wSYOz8nNA7
ETkSPRnw9s83UAeLNHZ93IVfmY70duJXA2bspPGkpvy4MiyeUp9bf9VcacAdMQReGjVM+MfmpiHR
9n9b5/r/WAbZmVX+k4QgmCVGwqaZmbA+XUGukPJVjKHb0BrYG7Y2MNAr07xk6viyZnmYaPAO1xnK
uTmsPDYc8j2lVK11V4zDjWlCJTKDxv07uy6kG18iur2mI7nTK/5QT85XjkK+oma7W43ztyOWny1I
fxgHYU/zIv1eJMtsWV7sDmrVAlQSJoZVQfpMRXLeuiOLt8pJ51o+57HBHCPYhzds965NM9tM7sGF
dOuBoAaK102NnEhE4VqInChxv4rP55sOIXw03AUOeFwYSBbVpBv0TtuTAPk0OU3wLaXkDSqP5YJM
l+YpxkiKAFLbjms5uND8lwZP1ClCicSDPcUUvtWUnlGJZ022mH3Pil9S3Mnh9V/qsQ8CrrgonwNY
gLcRqW+nb64ccxuYUZkmKKLaX6/bL06v3jmArZBezQdmdb6bNKe7HPWa/HW6xyJCYdJadEnt6aC8
juggE4+AqXSCQHo8guVSW7psCvHim98JQ0DCaXCgB7L85z34I4Vm86dmeFHGO49ggdi8duTKhPcw
QCs+P/37Ix+uNEBoSWdzBs2Ng5cILxlA+VrekxlWgsxKN5FpOIGkaFc+i6DtRSuOGZfMoU9Bv5zy
LnE3upN7BsN3g1C+vwekaigwW1II6VzHcjBV5dv9LzHBvjydhNvWZyGCWFVuj8GIt9FrJmvrh/93
O3u164PmZQXUFUysRi/BUqhxCQex2j9ORc4/VyIvqPu/Yoza9mhxdDoRiT0zse5VjWoNxgyLf8ez
e1D2IuVqRkigtpH7hHJrSaFhcXB2sWjO7SHYvdw6tT3wKoEaRx72AJSE+UtGbDkR0GgjkSRBf0Tr
8I3xRSrGMlHSZm3xBe0SEIMHnLaKd/xmZ8ABIqhZ8srj5zF2NY9zgiWu9Rfo+pNqWFTwqQr+XxyM
GNlfYSDeo453w9hWcLfifTpZrRZDD0qJr7kA5VvpDWTzMl1CX7zhsDhzYI5D1iDOL4F40Sa05OWV
w8p89QXHC3NSd8Ht4ZZI/lo5W4uyqMDXoW0fqefcOBK+EG4LtrYiVhDH1Bs8R88TpDiHhYPi8uxC
aDbbSvY09Dr2GY6Q4FxNE1G0JyZXxpC5BeLsVsM1x5SSFlYKUtTA0Mnex981lTh87v4apXIPENfm
ZUy76qe3RqcLJNeuVakBmB6Hvhfcq6h/r8CM7l8TAdTzOekuzMVw2E3Vgq9AU3M4MFuFl2vW/WjR
dzYOzjk5DM/UfusKaL3I50xvUnC4uvhhayUq++k61/PUUtmFO0Bzda32qHYR4AVZn9KtK0vdWTNm
nva3WBmNqKzfAEM1n8SSSakhg8KhCOlryn1QgunvHlEfCKYwPLrts98jjnnKOIbn4G4N+yOZdz3Q
OCsYHe/mykyeCMe+npOYTEevrr6886ean5FifxhaPZ5AAv+iuK/ij5spe7eTnYHWZ32d80EHIh8L
0ecUaAHxGo81IBdXRDLcv+aRuFTvdLiT3Y5f0oodbpBCmj5M/F7Mggy7U2eDvU/tjYAvV2KaATz+
2XTqtcixpzLUHS8IIIURFQnm3swnWTOWD+XrD6uCBNObonSYCuAJE6RdnYyy61vJVoAoc+yLpqRK
xOxLeKBXJLddfsQrG3h0MT6UMQj0JvTsX+nvrad9j5VzTDPpAOEkrXtepKYhw5dATfT5KpueE/Xy
7mIxR14sZ+WuYoGQci6DtHTYAanp/X/5Z8Bi69xXTx7nq6QDcR4fOaTdqq5iY1HVUFIb6xu91kDZ
WiZvmU25Assmh+IWFnghMcW4j8y7Fj9RZ244j+OR1L9fySMUIDfKttZOX1A0q7U7a3Vy9zdyDaJ7
dCdTi6suy+b1lUy2k3Uc3CGBj+jyE0iSE1xZPlBZQ85CelpjN4vbTMqnn2cGUGxzGPO1OTIP8p9N
b1pAmi70BIShXAiFwvsny1xlRKNIHgsaelHgVf31NKrmUdQTBe4QghhhprWL2dv2bCe5onaGcZLU
d5pJhqStII27ZhzRojYf4d6fVs4GHt+5E0PFQkdXptm5amL8ZPAS70CL7nVZY47dbPqJ3XUoNfNr
JQdjaBa93uSO003HtrU5WhV9glmJRtVLKt60MaA0KJXV3Q3KZpMR+haq+jizwc9Gg3mFkDLbMjqe
jNQRjiYRArETg9RxdC3v3dz/kU/yZsflNtgKV7miCEdE2+Scu7ZS6tf1ImoLa10twRF9HPKqgTxx
oPzHyxMSfRdwzu/PCH6uDGSZN9bPhnECoI0u+qNoOeeWJGD3f8So71Q6ULji49o8FYUJZkC7fq0j
rHbQY3NaCd3ZkeRuaX+TZCUpQwZlas3fQbh9r1HK0A90JVGJZEExd90RUO2qtL69TSlRsE0VpLEe
lphe8NJsFZbKGfaUKu+8WD76Ra7Lmb3k3mBPQNZ7BCXc64NCL9Z+CdI+iHIOrp3Y3a5lYVsd5Jdy
wfd6tr81R9dCbGGqkszTyUpK6E48qo5BRuUVgfHg807pV1F2anYH28M3yTViCZVKIU6TUnQNggI9
wc117ldtZfaQf2xi/VbYH2HrBh7nbPmQLN4qAzskvYZkqT7R9jHnzcjtYyODlalT8WkcOvgDXDqg
hqT7batuTfVcNMGKA314uKLI4s5vUuYmqHWMPRAz0rwU0MtP8YNwTfQdFOyH5IdS12gcuJswx7Hq
baW0sN4AyF1rimoLo6mGtaF1gV5uf1HMiTenSFSLzGf45RQHWbi3ilVZJqpkgUMl1Cb8zZXuhw/g
TNHuvpzkWkkPYVqNyPjIEXylQNQWaIgwJhCO8vNXEzaiXD1iu5ym34ZKcM1TqqIILQ7AN2gd5ljA
EDXxXy+3+UPCQV00Jr1EN1qgRQnUtOJOQIjbX6mCd/zTEQntQG/P8nYCVFtBldZooArhpmYXYlv9
RipRByfj5BZRaBoeYAoTWDGSPIonUNWFsebnSCyJuMjy3UWVvd548HwIKghGTdpduUpOGRG5ofF/
XNSaxJlxuSjPS3iR8Tz5I+C6No+Ndx/iR+/5gvw3OeH3SNXJHH7lhZTccriz1isM1iP0UacE97PE
5i9rNpOTNcF8ZsuPWr/Zv880I8lPSc8s3pyfNZQsqc7jFCFHEdsqQVOtLkN/kcc5ZihotZZEt4Ip
A/NtSzOa1r1RT+gA4VlTWhfYPn7YWhsV7SdZ7ApFg8JHfyfW41Zw2zEWtgjzl7Q9D9yOjThVqDeq
VuTSUsTahHVTDvJedtoRTKEstIqvKdc+XQ/Pa9HZrRGbeNvtvFp+EbEXDFH46e8juICs8c5hOS7j
HAsuQTZszYUNFbDUczwTfeuBsgnFqmyGRo0qfA0JYGUDVep/00pDPg3rk5UWSHUfwtmy4Djew4WM
O02bCZpg7teyKDW78oCZH7edGXQl7WIwsQGAX51OmDGTK4OGdtq1ZRDS9MPicFL2m0vQ+Y2qXSvt
5JguyDlMVC35SJoGXhFpsfX77YfpAi32tSqbX7G41d0QTX64h/WwRJwqdJvz2aofxNMmnG7C6PCw
2pJH3sQ3dRZRIIU4kJXUB+hEUhZSJ/ksds1W9GO1+62kmRoe7Lm1Wr5RCMmRe4Uk4UJFAApInJcC
2WagwRT/AgcD8B+179LC4e4hlPT+BHsKPCAHQOaIp6M549ptR3rnj1JUvlZBZOHUaI1Z1a/3jjUm
wK+WtqAQ4BXfB/zq0GR2c10zAmriBKFnMi5GNtoKjT6W7H3ezCmrOlRHPRIyEt0KS0OYcCrJHGOC
RtI5Lo+Ldfh2aqJbQLQcQ4HjnKfowFlicv1gS83hMhYbzCOk/r5kmNLI8dnDdw7O720f0hHZYa+9
XaDjM5Om/d9tALZUlY/05Tfz69tf/ic4bqMVP0UWybh9V8kB2VzT59nOnoXSJPeufqFyZafn/aVc
vTv9WYCGqf/C4+Ourf+qVgqjHyh/2XcSwxn87totwB6jW/w6zsTGgvhLRTnVPOaZjuiAp356QpN/
4HifSvyoCQeiM9P/VcnZZ+ha0VjHwU7mLjUNy0ne7+JzzKb0qs2uUP0Gi79v6W/vYdvuPJwQ1J5n
wkxCQuVzEDG9GL9LLa1xnTj3F03weS27p2ljvpNvoSopwButLkcWwHf+oAYE+PR+KTHV5n+Ru8C5
uOJMsVN5HinMebY9aTq4FsyLc7jCzfcdFNVBQp71Ox7xJ8u+hEdh7dQiJMXHerLRPGtqJBx6ZwaE
WzbKQNMvsib3hHHRy5j3lvfR8FP0BcT7R3HbS7237V6ts+F/23EBtv/2ilPmW7a2YigJU3Q+0kOa
EdBxKLxMzxoMVVwPBWVBmQgNMEApVRz2njcbxyT6D03IIAio/4I8/P66Xt1uJwuzHGdLYIFdqo11
Jer5P48utu1yYItSIrzIl+s/3VJWjoxZUvyQAGACWMqArDWACEt/Er45SWY9b3m1DRsvbN/eSC+m
dzBSi30BIEYOE9GAC7x6m95eZeguffGrijjwtbfmyJJCr6VTLkEPNKBBCF/vvPSDlyNqdk8M37dt
peNvZ19DTWCr81sUfgwsXePIuNyzGq6AzXDbo9I8wVUszFIzoZ1JDsnnr9oauZ1LeqEIU056xhMY
kC/3l2QJ/e+eXt2kpH0GfI1/jjZJbV7qkx2ndlYc1dSckVu1kFx9BFq0ZMiPY5/do7OA06y9VlWy
RoKueiaV8tepDtZBtlNq6VBDW893IIG5rNN71G667fLw0ZQ8sBGs+yES55zxrIFwkYYUNFL787nh
7Pm5Ab35v7AFg35TBSSxP8MRKYZAd5r+e96BUIU0YsI744SMdzkH95pWU0i3jdmlA1gXg38omr9H
A+kNWItUhBOc4i+viuPG1MGSupq73mZ3wp50xCkdUzBc9/IWGdc0GYFfxhjIx1qFD5gyuf0WuJme
1h9Sl0O386BcVlN7rCkqWisj/MmdvfDsw5fnqSgms+ujEcYn2RscwIKJLNgtF9CkUik7iCUvOAyN
uRWXWRF/7NYVDBj/cxIU7vEBxIH449eFIPhWuF948Fhm3eB3tF1CuWECKc1BWAQSXWE2Cd3TpXFX
0tcMdwB/X3NMzccoRSkwQWLKLs0h3ptiV0f52CVRq+SjteQsZXx4hSWNIPtHZcZ2MY9RQ/JMSO7n
9+1HMI0Q1Mboro3/kp1xfhYCMlCfQLA+VZzJkZlZCsVnivWpM+Aj8yvqA7q2wRJs5YQWfH2/mnZ6
NlhYQK6lt1mvUEZ+opgurrkzDTQ4fX46jRAst9MyuyxLJDiY9OWhs20vgsV5I2PgjHMLyR6sVRGY
6GBN+lQZANhSd9vpnn0XFTBlerYzuevDwbsHPIT3xLMLAEE/UYeGjRpLY47IN5HnrJi/R7On4JEC
6s0eRUtDDKcyT6pOgM5IoSL2fbNWbZEGzoZBidDsTuEUbk3S6Q0nt8uW/JmYhdQDQ8tXwbQg44HG
d2+ws/O33DSzWDAo3FPIQ4wcRs97ktliIic1P6w0Wj3eZ3qb8Wy09dOnvZcQx/OU+t6v2pkfv+TQ
Rx/jjMANbRIMYHxlmjqQp8W8Xxz90RCNKL84TVvKP38AsQ8bjc2b/k8vxW6bTvENF0JXNcIcrMn0
Z1A/AG643j9ofU7fUUv2Ip7fYVHEIIAanN3qbEhghgnylxm2fzrzZ551K8TNilcAiBBqfih5Ykc9
h8BNtOldTnCJRtHN6/rWI6mug6evRIg9aydTUnRDNoMgQMx4Yt/r2UjDVP3q32nBcTYVi7kxaHDO
TwI1+qzH6dPW4136Se+3sNxzWEuHWhABMueUulzCdDYxofWCiqA8MMsUSwSlbc4j/r+IyVzaN5Hu
CmrwVdwbSfzFw50P1FaNc/dY87nQAD2GNollQgAXdVcJsGstFjjjFt6WD3h4OyLD9ETWP+ESfYnB
KGv3RDPC62xBgUa9sU7c2uxavYkN46VDFhWnW9DlHBz7ZonltT4yfSA2Bv8a0dKqNQlvhEEC7CbP
+2lfViGyZj5Ds/fuX1IvCjeLNTkvpxbpReiVNmPHnZNlXhbgvD3vY8jVOlmOhxpWB1wDka35yTj8
/s0JcUHFsfIa7DsDbujhE2Sa69HPrOfDFlSVqbVygvGx4T7xIB1Ars2dOCvX3V9AgtyvB7LSlfFj
SxlyWRajqoSLEY4CyWl/7Bn6InfSUV4jWnkjHuQ9jjYM/GueZGZ9sGBrHy2fVdD/snhBjHfDkEe3
RrKth0axS/2OB0cFWZVdmDxLc1afwZWuJe4KCXZ0kHZHcug1zpt1os2xyXqk6ttuP0RuCLx8bJUQ
zFsO9/wfjP9fXh3mfWVNLO3tj2lfE5qIkRd6bx19aeDrWjVRGQXWZSowT3OSwgn4q/pKbaLLCpPy
2J58M9ayuHdFm8JMr5nIrosA1nKaD7iEg+tLTWjg4WzJJB+48d3v3QHRclSq043G3okipD5T2EYu
giZY28hNSghxJhbEmfrFY3gGRUc0QKnqq3MtCKn3IS6HmwUB9XY/dRaKh1oCOXWG0sAhSqhrcfq1
VRlrFapKhfnrbX2g54i6us1onrDXolMPP8xH17oBJJx/94pZzMd5ggZgHsHBE6z4onyVK6QtRkut
zF3Ye39CKmW5o2ItNpjmr41cgloTU+x/XYLutUeScPWnVH5WEhZCXKa8BB0Mr4YrHJyj4TnCo1Ol
L6tpfrK009I78pKcY/KuOQnSe4zescP1hsRhjsFaHkxNfkLmF+qoXuvBLhxg4Uq5LH4K6tFppfjg
FvpMls1Zb4keQAJ2Bf7J15xr440o6obHcuEoxesR9vQ1iRM5xvdOpzduBkC3mBzZpRUhSZi6DTe+
YvZenN6oxPH3oxvvOPCpQkb5WKG1xNvwMWfO2HoGTn8109CCDoyM03wIyidx4tRLmkzuLyc1ljU2
lulJ3Zw/cOM8+y6x0Wbzq1wZRO1vvOIT/uKLpwdSNfhfeupSTDBLHYlPb91tHAlIqPs+vLEwd2a2
k+Ar9OUOaOME2qy/Rd12pE2SW5OrDa/ST9wGxK74n9LcxkHeIHPBrjYA9sTN68TRpR+NM6znR3bm
M5jKtgPs+W0VLvFBGBpPww3yEiJ5dEe86/xbnxuRyhKzTYzh5DGG7htnXMe2XqDOLLU/vbEnePoL
HkDzext95E+LDXlVY28Y+zmqsRsseRA7Ni7HkUO0nGYWZDwRZO+UZM6jMeD8Q1ZJXlVM9WGbYfDz
5i9m3Wp/8dxeiO7rxrdN66Y9jpnqCFKmcN5ypwWipuLDM/YT4Zo20wd460b9fD8rHFstmUjJYUQ/
GWSBQ8okSJKqhpv6ZjHBb9axyn/aFYG1H4gHT2PbTVrlv/8kxpRBL1igPOVOzYJmstIYFpnSlSRo
VfLlW7u4SV8kUzhUhF6feA9i6KfwEx15sq36Hx0bLdZ76FX0B0mkXRtLDZ+D7riRZ0MTYL9+JwJA
75AYRIzFiz23p6Tp8DbvYrA34MuGWOvVm6sCgTmMoHOtCdwypP8qDGFvw//ncT9KMJZirwjYqjuK
Bc0Ycgw3ttWfrJu5Hq7rAuD9NNUc6J0s+M0hyaqmR0ifG5zrkQd4befZfzw6s7mDxA/VLBIJdrhv
hLGtd1J+we6m2z51py6wv+Yi7W6vto3jwYhFbqbMxtW+FDqX3Uav4ztj7+QobjsuaMulm25qlhEa
gR/McXblWTymwK6d4x/K0QJKWWDZfkA5p6NbaszY6Bv/S8lr3Cnl+UgbqDPm8iQOfvva3vO99tW2
6qWxUzkOI4egk1F1SUCPlHmtBAaPuP+1qK7f4ewhJHCZRP1FnlAhbj2dfPyWMh2ebIf51WIcxXQZ
6xcQrMp/wSEpv8/qmD0R0Wha3qUy24oQiZJT00C9P1wPzboVIZ7yUuZLaok6IzHubkzG92PaCLpq
tXkgOOlYdn774NjdWE50+FV0usgbnDkYXu7FojSfMRSPnGBiMQGVoivQg2rV6V9KnK4+vV+efEsb
lVnYTfPotNPBXj88ZlwJ0VdnUd4mGJGUody01GbwA3L+HTDjzEtt4gxkDn/vGcVGRfYKm7ZBozKT
CDbh1svImHPPXv7+geia0a2uUR2M8t03SsGSvczjHz1XvtoYWPwU19J6MLTwdiLysYAx6fMV6Otz
X0ei0hbywP0aOOd1EGx6JwWuxl08z8Cnyklb9wNLBihjI4nsLJKrDDQTW4QhyPN5MTRvN8JfKpHt
n8Fc6gpJvBv14Zrq8wZvwvzvDH110c9BcGEUXcabuDkaeAAsxfuuxAztKM3bb/KuU0HQZ+FI3xea
jkrU82Aq9yvRtZ2E0mKEooG8igfVGNMvgKi0kCNuufo6bbzdOzm3z8gaw0vnFFoTQffCUqHzRJIp
y9lcnMTL5HlifSPKs08dQPyCB2n+36n1HBR9skPKHB6RBu0eqXpQGlafGLyYRoAJMUJi7WYqolQg
TFMsYYr/S2bg47fk97Qc28rdx7mW36aY7y0QVMdm0pAbxjw6HoRuxkXaMsS5HuF/99v7H/5VBWRA
v5r/JgWm2t7uLosvvYED3rov/NqFwVZA/lfGrdBVuo2dweyokLWRU+wW/e1gM2oUJR1Ol9OZ7zOR
mTq32caC/S8L3nNTbAT3Uwygh/Ab5WDmInkmB+cRtYfWQTwFZUWwqsoiPBbo6wFBJr8U4/NH/Q6+
S4cuhhfl9cyB9lNHMSgFJOs4NihHLuP54skWKEmEl5btIjpwPmHzpMo2NxypPw2B5SUQr8ZgnSF4
oJPfQmvlvbmZRgDMUnV5yxnggv3FkHf0zf4KlxUdCIxjWyTUPeEvNedECKxlOV6I9RI66Qvo/x+X
xu1YTKIQB68vDml7vBcJMYCL+h54pQDHtZP9lyLyS456qeoMCsal1JcWhCIVtUPUe4Jq4jB5Bcxo
SONQpQRY1PA2fQCU6Bv7b1uA+ZRWrRfDbe1ZyJT58aXApeKrgiAVYI/SzK5lcgdsxa1H8gStK726
kB6s/a5QSzOWKuhcf/+/XImWo46B7Wk6OqtoWrdfvge4hK2SvDBvdTR2l16Wu7yv3emAv2mGHNKJ
vStANo+w7xG1mwveqouVA8ivzwmBDCgw7zvlme5ZHL961nX/K3vGreCJMnKv/R9BaOuRbjlRjZPi
Ww7+Rk0CgSxEKDx+1cCq7u2il/S3KPKR+Rs8fEKe9CITYLAkDMXzU/20+4mos1Thy4Z4oUl8995d
kvdYg8HFuSqnXhbBmL0uVeHyr+C2llO7FLLI7Q+NinXWsz7fu8z33Xg22RsR3SrgWNRd9xldXhgV
3g2J5BFdMRx34Huw46YH8SljXm6iPGWWKktBRbLjAKoiDEUrsKgikTD8C5cS9Xj16BDsZEg9/lkF
Irf3UzrO62jWHyUrpMnX1zNeyyWF+rK2o9Mqe0+qTI55y6MVvJSznM2VosHaoEMk9X6FJRuy9nKT
o+HnPlTRfHvjxtKD1k1BTEVcnQr6bfuyn2+Y38OkMdv7IfO7UyLnjKY4nRsA19H44z96voWzalI9
crS9tCfvAv6YxZOEnJu0AWJlGPUfFBvuFr9L95AbGBMiPDRJyMTshHZdbcAcbUkevTo136NCkuw3
qiynxWPyw3js46ocd6pdcsnICfmp8zbox2qbn87HXmPvueiYnuQwPZtvfkF5WYf2E52LimcdBjM0
Ih3Lmm0HxG0n0oOO0mcIx5ZPV+ZdkWoE1Kyq9uAxoVLIzq1ID00kP57TYkwW6LCULIawfT7hwTf4
4n3JQ/weKn0/OSrerz28GLov/YJ2m0pr7j65qMBucstCfKQBQ+9G+d4IZUe7aj/DZn3dJHFxKm9p
OlTupEbkk4YNnubWAQB/+bOni9U3Uc38Bp1zJ72vSFXz19VS1g9GU4MHZhFB9g/Jk620wWYmLiVu
KdInaWa/jG9Qwgl54uijFRZ87Wl9Xds/o3qa84DFMi5LfX+X1uv/PVfsE4oeuj7RKn9gA+FhfBfk
y0P3m+tW1xmbsdVVrijoCyRSi0yJzeaJxM56PCR9Z4jY+uhGSGOMw5RQNu47NgVAkU+KCNyQPeQU
iPpKogLu8mkucTXGY5rSOwBPMems+eDUg4qtskmCQq1OGZXffgjBL/shfOoLzHf0kvfhe7HdeclH
E9idWIM4PFXji7HzM/FSwmmqLjzyI0GGR7uMXHdna8cea9op/SvYSD5V368n74mo86pzaDXYsXMO
7E/H0zRELq77D4S1mprrRrqYwWwZu7FOqfmqtdQLmE7T6X8UK2xBDxSQrZwEfZI/iOBBmK4S/Gpg
ZQNmHAxEhEc31Cb9VzUIsewsIJY2vTbDT9L3Ir/CJP2AcmOlWPzggla2Nwz5vA1sZgASzfJPyLOI
JfP4+KvbTs6zx0QS0t+S7b4JkYF1WH9Kh2E0FS9Yt2ve2k04og44sD82DfLayvVBdNBawUWYpV6M
Z+vxeMtQJBkeGp9/Y9WPHz1q36ZcnBDGbjWHTem8jzNIU2O9aqj2h5phl/xc/jx/ElSXxXiNn6xF
j9m6tuSgVj5H5LUaMui2CYxDeK8BVlYQKxX8H+peYyWE3zR5VPTGrcwGRY8GD6L+oPoiSaClcTei
Oi/nZWwmdyhx+czzeZA+9x4BqN9xhPHPD5ta+aINJ6KLqC6r2Lem+sR4D4woY2nfyfTw0LKEsOdz
fe5By5w+HLJWY5M+FvK/CTRZ42uaIvOoAQLn+YpSwNb7dUGMBz7dPj67HeZa+K/uG+crdRiIWjh6
JczkJlLCzzlagKb5/YqbGW5nQHwFI33VwMm27u9CLg7/CxaF2cIJ7Et2rIk9fXMDmWgo9SmW6eZ8
b0TLizwY4wX3bCfxqD00rRYwF50PoJZ7IsdPm1bsNEaG4zGi/pDe03vA/iNiIfBCdLj5/lCf6Kgg
Ka1gMKqf+yD/opO9EFitZXXAuTTz/aXz5TZospwF4pQpRCmkJJqScb247g/I/3XwMH5IxouBvmUL
N/cWk7lR+smpbNXQeerBtjVK6qu2wKrXwBSg1UOthwk5NQvQKeEe81y6VwzVvlm4BmOvHNCKCXep
jBODrAdRyFKZR6hBHqTbn7f7/WJkraXjN02ZEJFnNbPIqb0hPn/wq6O5tP4kXp38j/LUZDROPsgw
1hgVagwIRLGO0KdIemr+V58iFqxLdw4jgPh8xPR4Y6BjgbW1x2Smy8jM/GvHN2qynU6XfMKWA/pf
+ghtgPquW6c/ir3mgcKLyEkFx3r1SvJPPJjTtzo5gFFQIpB8a9mIOIamTvOw6X8mpBT0nzP0m6jv
5xq7fKbkPbOThLiI6TIx8I8zPtwOsarbVzweeKPQx5cJYADn/TzLaktKlD7LuIOBJExTp40DIq+e
V+XV6CO1yu/80jjZTq4ZKez26N4bPANWbz5BLSLYYa9yG8PDChbAnWHTy6TA7STd69MGXK/dre+q
aauHTv0ADQrPa5JjbcbWPijmNGl6Ik8CaGn/SN0FMJd6O6r2w398ElIuPSw07gZ4JHNbYAb0pHm+
GlrnojVZoc9agFENhG+f57+eig0dQHfa6y6BM3VkGPZSFpqQOtSExv3tck6r3g1v0bJkG4sPDg7o
B52kPw5SYrXi9rPU0nTHdJAeFsPpZ5r36V6ly5xmRXsG2TFVcNFO3nJ9WQslRaG63ZfFlIgllL8R
Wu6geK/9Tbmtn1BtngJM41hehGob3DXD+kjNSlgjyNrZU1uc+TLwyDU068nVlYNQY9Mxx1if2Ndz
FCHjRuL3t2PLDkL9r3M3UPsvNyQN1rX3yeWsUtkBqDr5TxWebM9FHUkyfzw3o71GlZStbLIYYJhx
U94BARchGEA2MmBd9miA7WWCj84jvTIfmDOH3IlcqJOL/BlsMEvhhdb1xfhu4km2tIdutrXhHtMv
MbWlX0kfJD9JGHe0SCzwKdCrvbZ27zY1RzXlEqa2RfhRXWcwPMYyQZ3VuRuT4THE+ZjunGmhIkyN
OGf3gpxBBrzlAUvzGuEqr469/Jvmb7zE086HDNmMSe1KK9d9AgGXOUR0T7sqMwfOOKQr+JGDsv2H
lmU8IBvmWtCFyTA0anfWwgYLhRF66xi+MSGdeMKtNOJ3gp+tASZbrhvuF7Yhg4JrFhF8c4cFX4mM
WxKbFDGXM6TlXRJ1pisJI4LOKqP+4oyjr9QPllnRsthrOk1CpPj0FN4wvyr3C9FF/rc2nq5vs9km
1DLX2CQj4WPcUiYyPnKRqG+VghaV1wLaVGNI3pJt+slYdQ1VqjDoNDmAczQLNVmrnwA8h3VL0s8y
dJeNiqY98DVmA3zp5/pyZ+cnFF4omTw6Mrj8Hm2/rI/vwN/vHUdbwitB/zaeztfKHQQ8AYM5obCc
dqmPQRAeIMkjKkVgaftSJZFcrhvshYDBK9X3aIbtRAsZOYv69UuEoXyZ0cn0MDS7TRmEIebu7m7a
QoisibuRgtqWREAc30ZrCAZFdTB91XwZNor+iMCaIDb6BrR/+OiOzEeh0Tt2tBNK3p3A60DpigSj
XYkCBiFmdZRq2l4DYdsZj7TumVOMOhJ1ai8KAyRlTbpq0l7X1CQNKO5q1UCIB61YIRdj8ZLlwyXe
BSj66rGfx91KKVh+rExYDkdJ+6hIieNZDo5oeLnKEBtijl3VcfubaMKSGSUWnH1AebaNv5lRB+uQ
qd/MvabbI++S94wBvKX7btyKQI7Qwat8nKiqL7yrZxg/lSMn/+n6eTWn0mBq3u5j/Sh13G0wcsZT
XoIPV8bNcAJkde11l0OA+X2Zo9UllkYilMOW7gRh/ZVCg/Qy5CpILDPpRuWIL63+bDKSBT7C/n7V
KfG71Vmv5ghizwi0Sez93dsblenp4yxgaI7UGK71GhPSPMd4c5rixAu1GFlfH6r0dL00wbdMg73h
HtKJ/TCzuWd1zgo1KWZmCPR+OZ3gBqw0vjoaOUkORX963L/UiJMZ4/Y/woIw4Pb8DBazX6lgliDN
EfQHD6gKjd13e6aUP4A7pcBDhTTx5bmz8hXtnjxx5NBYUNZJqN0h5ZSegYwsvFXRG2DC5vxc3Lvz
KhmSiTQsqwtUz50mjDx6NP//pN0IMAYQjFrywA3C/od9Dj52XQ4JNathBVve9JXeF+qt9f7lbZv4
efC1in9w9nlM9dxhFpRzGx2Bi5H80jifzOb2GwaRekNXl468LX528MubSAas3J/DGGlVUfIVzx6Z
UfODfkgHLG/rS+uQ9hatyGNsr55M6acPihajJNlTb3lqBJmb1VYRIV1JXmX8zyyf5IjQSb/CYR/+
aOfmra+SdgkQ3OzH1+u/1CTNyFlfvDmhzpT0HAUy99Fdk2m5BGYdjHaOzKnaLyUTW6wgIB4UCAOc
WBBNncv/ZbWb/p8BzEa19RpyU56OzW5U/hJnqawjwlvxdx8dx90g5L5U7XBM6lb/Lpoi6r1SQVDR
TqR9xHsQGUBi6sv74lro1zTRE8kRgD+MCl5z1eH4b2aZXn1Psf9PgpqE98QQImzUYNOTOTb7ylWI
G8upT9EyPqNCiJzCz6h08oNuzbtQqXp/UnIOc+N1DKou3TyP4aDcHuexuW8CbXKe8wFPucARq7nN
TKASsY92UE7Iew8UV+JHB+JeKOQ4YYor2lvEa2ZWXZkjyhgTsckOXdIhc/LW4cQL6e3fpzIXWW+/
tN3grP45nE8IarXCwy0j1BEqmdmwENOVBtx/7EEsvvrp4Hd1zuBOuneFbCvyb4/6AnwLAA1Tdyzv
6hVYeClEDDIXPmayt6aQPFUZ5c3q1NtrsaprxUBuBnp70BmqWJTsYXvSDpoXLRRK7ODZlTii6bHp
BN0lzAkX926DHp3PwlTXkPvl4kQDNvvp7lnvzn4xNMaviwL/y+RrYhzucGwUhVWtTw9Yzgoh3jPT
LCChoiztWzSkABtErZKDjQtcmvZsCVZQhfYEhkQq+1cN1N3O6Zl8fALt6pl9yz8VU2Y46bf+GIMV
3qRCzU32ryX73vyka1j+Ft0j/xSg/w0Ys92Jo2WF9SvMd0LQ20nBRVrImpd7Q17uWH/dULnaMr3t
AzXvujUz52qVx0K5KRg2Qaettv6kjyZA1oGIR6WRbNCeltSVeKCUkh7TfgRXfxOCLClMXRSA9jEO
oN+JojDYfLwupEom4h1tYybcFgtmKwPCfvamlbebNiOkVC0qvvfXpQgP70Cz1MyrzDGcBelTkCAY
GH+RtXWSJEPAxdwihvd2yHdQ20+prPK+l7/jmbovTlFCasNuhuNn8fGBjIB/loqs7fvhSID/U6BY
o3c+1t92gTRnnsyVOs9y+sge2TwlR/MbbL4pK6JIgfHigNYgVifz9tb+PztXStWESHjQ8NwqOIOs
VHAPHH0vkZY06cqI1KfbcPYglBnSIC3xN5c+95SBl9b8RZEsuy1eAjdGyQwCuPKUJjyI9aDS72r6
ucmm5FOK13fHTrSMYxNBL+0TTbWWoaC0NvsCaflK4cwdAKcQ752eGKaO6wtxhnS+GEjWCOBqePz9
RP6p/XC55CvMeTnyuwI40gT3Z8QKkI/C5Lcp5i5RUe/Wo39PVn+t7d1f08CGj1EiFEh6Y7I5hsTb
Bivym3pfVbhSkwXDwSMj5wdd88t7oynlK/KgBRCrtQ0O/4qcAC5KWkk28XLLYdViiUmOocJknNSY
87RQUHq1qcWN+knlRNgWIy/tGN2A9/bBmLtTDD5EPswC9OvB2GGygvxzxmRmqhewwyfdy2XUkVEn
ersTgxEhXEjaCxG7Fj6gDS9qp8ynl+Is9Qe6Ka1NXTk78SrhVIsIELOdxRmz7OGwo9QMd+4zekK/
x2ZQHeeCQE1wgn0g3TX2HMv6lh9AgdLA9VhVKVqaCbzPymMRdVaUgqc3Qmdz/XnQo31oLvTpUotn
SLVX215FUAf704Zxopb9SAlKGI2WoTKCMXs3W11aJ4fB9C/CFeOr7/sv/ogYHwlXWb1AFHZP5vJY
rTOPh6/5aFIsK48EutueERy8y/oH5OYp/a8phY3kUwolMbhB27ViJxD4nwUXeTDZ9MdyMEgSMWc7
vBFcic0sDU1876NkNaVIfwzbVUC7goUhzg4S+D4bVBObSiqXTcN2rcaI2XHhNnbN2S708818otWY
wTTf6a8lskVZcd/tXzG+tLzbKs/1dZWhTwVzM9ArUw5s5cAHZHXxYpf0EBHhraVPOy05gRQKNLdM
iLBiRZjz+sYS/eeZV8qdl4y8/UG0ueLMEHFyIgXGChsEjdWQgztSF8SJyN+IRDk5CSJM2Em/uRgn
pmp/6CiY0xoX1V1iajh0S0qJlmNQmO7yjmtauS5G4J9KzWwlt/PJuEL0SEcm21I3pgQGHUEi1Cng
AX8EImCftmkILjnbmfd4xzDB+G9CaSgIR1y/OLXF9AGFY6KQxgBhzq3/g/auOnUMhde8WwxnOiVN
HiaxHgzhPuTitg7434hXrJ1faa2Uut9NnJA4WXB0qFrdJ1xz2NOjQGcxirDHwD6/jDq8RUk1umTp
rsSSf77+5eKbY+WTZhCsi3ylU3/4yUDZBPbUplApYjbcosvIN1fNiaYaqegnkZi2J7sGP8aiwTDo
8tGQFVoJrkRxuJmnZFJNJNd0/VkZfpnqR96GxxQm4s6nItAX9GH5cnmjfe+VzZaE7wzvYClh//7e
9u3Yu1ugA/t/lGA0+mR3a8mje5NR1PTlVXvox0WoUNojbApE5eoD1FY8/QqydiRy3mdufQJ5aWCR
MxA+1r4benqaM1SrNUOxM5IDKdZu46koiEIWl+y+HjMzBXoBhdpRwHYUeMGON8bqD9hyNqqtLJq4
/dZTCbMa3BDt0pV3gk1H7oaKx3s0IidFqrk+GGM79U4yq5ZJ/njqYTPMcYiaXM9xfBT4CF5ZPHtu
JmHO6se7jJusntvJunUZS72DPshnqiR7Mit+x/jOlpQhh3dFEdTLI9rjmdD6AvwtIq1wAlQHVt/g
MZ3QRIvCwFsfCx7P/+87K4sj2YNNk4QKGAMj0SVgF1O7/qFaO1CCNqXT/OpLWsV/vZEVYGke2LEe
+OsId3cFjnuA9fhmhmHSABeyuICjdjAeqJ0nq4twNn+KjeOFspfohDvmoQ/Fsz993Ta0dwgcLaJ8
1oLwT+a60xPLmWv0p9g5J43w8fzoQ7ghulWpefceUazqvPe+yNVF8z5YsKASRJVAOhbSOYaZmhXI
n6DyY493Qgv15OVTZJGZ7lgy5eZ/n0IFa6atbCJQ/MQuD3/caaBZTiZT+nyonr/kE/VOe55D45+r
t7mpPkjy4ghsWXeR9DuazK5PAmfVta9lF1LcjV7MIc7GMdP/92a2FxwkBQNLf1Nd192dMYbweKyl
B1UjvxeYNvNOYE3sw+Wipw9e5phRNhd+CEIXSzeVsR2aXqo0VDi7iIbpsjirhrdn/0eVjLUJuIpD
wWgjDBKgqOJzZKE3s20QU3CkE11lALfHhJH3A3Mnw4FX2npNwMKUeyzoQUYKjz82U/JbTss9Sk6U
QFSpchx8epvNpbSaHYUA4ZMDUJtufyBDXvwX1wpEjsO/wP2mA04ea6Z1Plsad3AE03mzw6/gcF9c
T86ptqj1SQbhIohq1rp++WsJCUkkffsC0amt8ZsBYALe6SMf6F73COK2wWB3s6HcJRtMXw2Jab48
qK30bL2fGxd3AJ7az+N4vWaZoWBcb2+HEEbo4/Fpr5rO7eTDAmdwSvkHbAJsiozVXvj0FS7AW5Qc
wgcKbkqT+GZYRmXSYcaZ6eveQ7wp5ocqsNyJ188hqjAB+kiPNqzUqrKz3prnbzgbhGZiV0ycZDzV
r7tO6KsGEkJClKSsOmRf9a7YOxAKezX4IJ6r12omsLPwNXsLcKUR3tmfHmSe44CAg2ZHTjrsVr6U
BnbiN2Z9NNOF1UjRmastrUw2EuWr1sJJX85OV1Q6cn6uUDSuz5yxFUeK/oWSdwh4h+ZjC91QG6MX
s8kqrYeZgyW/47H3VsiQXlXPSkdevI3a6jsUt/cq+x8BcxpQvs8y4JdFZpTeeP5mghLBqeZytRdc
k0FGWoWApUs0uvoRpZvdr8lUMZ5nXQOsFkEuc2L+RG8DOmIkfzWplDowRtGRhZovVkzIBy4+83dv
HaeiBTOI3HCr4epEaTEll7YphiERkOBO//XhQ0ETCHU+bNSkJ2tJHpPqON01SPG8Zhk4PafEI0mK
VS+AHcMrG4Koubojbt/epKnXemSHYPyx0+vymA4xj4DPldGYcZr8gIdSmgXAVmiWcwhvRNNTyAg5
siZPpJiMDiDAe8gD6FRDALP9rzpY00Qzycsfkm1GEgk5K4F2cwdn3g0hW766pe39ddD9pv+Wwz0x
ow7XMV4eesHFZbFriinWjg9MLrKYQZwae/+0WDLfOWf4H/X6ooa0AlZ3/lt3LY5MvuBGJ0819sLT
BRmtnvNBo+shaz+7dQ6455TtFbW0QN2DloWFD6grg4nUSqv2ss3G+Yv0+DBPJ2+iKuEwOeAUySOz
CilvhC3e6IeYJJMehr5SK5qAHNWZjXEEmW4CuqBZUcBGP0J7gBC9V53hGyRPGP9ksAlFOLE8T3wz
ksbT8AbOQW3nOrs5TUMAvIu/YEalK7jvsSFVETc7yMmD549SDYs98Gc9f2CpZFhFHYDvzGXg56lb
1o5t7ct/K5aEvcZW7okRycvcRPXIR08yCx7YBIGDUggd0RNM4NVpkur7LybGS5uCqnNJqRm57yvB
ScIwVBNRPGgCzVA1oC5Le0A55fFySVDAqlBhvXSVwrfRnr0hkAJc9MRZbordu0cCfglBdStGg7GR
vNzt/G6PxfxY7UB0N9nPiJHCHu/4zxH09bXbEvTvY24Hh80UjMgcWnD9jhwrIfXfkCIpRzUQbHRO
/X/hUtk9dyJTjbZ+eDUKBEj9eWgSx5A0P5rVYmCCNZpTPgog7eFtpm6bKSOayJdJKox73dEYP6Xe
vPmewZs/Nk6BKd34eLkXrX+fzXL9phBBrzUXdrHb69dr+TRxhmpFSHeLgUm2RS+D3Qhl4Ox2KD91
FNl6V99mQIctJWYXBUTygMxwrpE8wqqb+S83SVbrsO0YJXug1A78h9KgK5ngZ8PFZJnt6BUAjULz
V1Shv7Mt1bOgB9Cf7GCMysSf+NTREhhKaVsiLSfopu0LmM6Aqiddz06+m1qfXaFiXFc09wfxZXlR
MLeLkP0q1+fOBZw2tXSlbdCeHdV4CWz8FoWteLFSB4gwYto5FSwqTkRx9ljIKy1uwhuS30UBRdgl
TsMBZNJvUNvyilnIJky/p+wKcz2Ut5nuISNxQ/EzMt5Y7fCqkYBNd5mtkMkgtUgxrlEVOmWtGNwi
2lJ04PIKCIbPCujPKJYWKTnpBKuaoCCbY10tHx41DVgl2nTdYRTccGxWU6QhTYjopLjMS46LZfAT
Dj0JXTxQ0cIl3dO6lK1teXoZC+INXoAQNKjdFxKHS5OTz2GieMYzmI0DYnzjiOF9HievRqaChlv6
f1DHxF0Xhw23OmfKpObocM6fJxWp+g0cMbfxBgrzyENqQTNz9B2k/YUzZ6S00jqDkVLYEt2Oz+Fi
V76g+I0ccwE5xcp0ynr6waGEezpI/+sXMRraqg8Rv8P1ajLRbpwlpapM5X5VvpaP/I/SeU9VD2kd
//N5odbUFxazQUmPhlNczT3iQ1ung6Dqw6imnicfBhgL6H+jCB+xXQUxrDiv+BJ5iKcjrx94mINk
lCWq9WwJwh63FOFt/WWiYry8Eme0dhqItn9wvkAmpwElmziQKhUDiHCT7q+ku+Ixi903U8I2SN4B
u2A0sdWK3PFSPLjgomMBbu/jGgw4JX0FLB2qIR3FZtEBAQeYc1QiHGH2scmt0URmDZhuDhWMeyJc
PKAtkqsSZUbPes4J7Iaj1XzXIz0eV1ZbZPTIHBVeRkrLVbqPJtEW2G3hBCXFcEjmO/Qkkenb75xQ
QarLg2mkGh3cbLq4/n+uDd4X/hTnWeu1jq0+26luhUDFLx24QRRergILxbdG1PJC6fTI1OmFQFUR
yTk4xlcQ+wxO5qcd9adLdK8sswUsVICUC7vNMS+Fmw+JzxximykqQfCQ+Fccji9nRVBnk3qCf//P
yj5cytNHnSUXWCkFvlLxfYmKS/azJgppL2Ak3bmLng15GOCq9uUnUAlhabGZ0iyI4tQYy4XrnfRB
BdpSk6Skro2B1DiFKb3CRx0BUrwIpk9z+CY85ft80Exo2hA3JI4PyVv1Z1Ut8ZmyX5TnMmfX4tfx
VyuWbEEcNTIPsTQRMNJdYsUA8aJyYmjna5vSXJ2SStgoMW8RWUsWhiLnjUohDsQqhTHD43kY57+Z
rU13sZBvDn2RGhHlCJk65ktZkGqUOmYlhBSso7E3Auepni/cvsd4M04GFuQNq7yKA63oZrTr+4Pn
JbWffX/2HrvIiLw8gKjOzo8oMUzVFcQxNrb5DvoMfhhW9c7kDYYYDtG0C3/JSPuTVPVXVJrCBzxE
Ys1vJKITXEiI4MAZ1h9dficjoi4Gqustnf2SWCYtEJVVpY1az96IAy1pGpgMvvhYLDfv+Y6kR/LG
jsep+d9B03+eUK7gtVfIqttyktXSX2BZ0FcgBTFNLyg5s8L/IUU+F+B7fBWUZWnEJM2InSQr5k2g
97m3KJF3cCl/y8kYA5ksVtKSt+coFYi6BKOfDWCuK5E431JY4Wj00apyZE7bYCOk8o0DKrqMDMOK
XjsYV/gbFcQ8TiW50//0aMviU+lZkrX8w4m4V29KEURa6+J2opYuyJnFI+F9m7cntH3/6ADiUUa0
KWSizi0iQHg9f3MQEcY7SITnNTCkXDzeP0P0M593sKk+OSYz/3l9gHOdTGSMuPkktsX/Uoegvln4
hFRrPSytOd55Zzq5eDGWe0YN43y3YFX3hke+mKG/JJV92IIvZBY++eMV3zvJEsV/T8Y5O9kIiBof
HHDLVu6wJHE14w/W6wU8T738ZJO9wG/97CpsF8SspJJZ60Ouz82CsTrgsci1Zc1jmxcHqAvU0qDI
XPIWBoukU/jaKb6unWo0H8SgUlTc+1E12wVG0VF6jFhZ1BP5TW+1E84TlhmntxGppF8lTrv5gHzU
USfwss8Ii6xcX8m/GsX4CjXWb+StQhDGS/KsWBw6rSyqKo+SxjK4wNqPMmnEFFF9aAUWGydpuinm
uql0p3o0+B4R/wIeBX+U8ySWX/yxFJ/Pl54ptl8rf/8cqDHA/MgTVgPAKJUyoUt00DiAgiFi/nBC
+3s4rNMNm10noWjQ2eTyLwLZAKxy27106TViSRMhX7I/2IC8SDKia8AP2cAA3tU0VLvbMJXpAQ3H
zjKhdni/vlIBTB3s9oXm6lN9MyWft9vgB1kXPrX0ELYTiVQZTxjsPk+FjhliUCxg9ZIC2cFdXK+b
N55e4IeLG4o9LoNYkQn5prDsUtNp1jnBKCuAmcjQRDBpZChbZAvaXkBo9l+ZXVC1twQTfKNEcvVt
uqDkoVXoAOAkqcmOVyk0Xizt0KzVFR4wQuQOcpRgZjqacGDCgsfgajnIZD6+Tc59gr7apicyMr2F
bro1u6QgXJSHYUO6g0h3Giq28pBeiHznm77XRjda+VC4adWEtIfpNcZ8i9H+4+n2JQQ2npg0Q5wb
Wc0wAqr3RojKDbMJ5SBwxxgc8zWiolJHANomXW5mAD1JjUZp7q0NKJFgeOYFoAvbNRnN1Ba2Nge/
+4nMZa/n0IR72fkXpUitzve8tnxyh3WaJfz3+xsnArzqLqb/hbvRL5SfaFu80+Yy00sAbmR8vsDH
6UZWDDeXxDAWvpqvDqlQ5z50bK86sBWTxDRc5bVP3CV6REZ4TVQZulbJZ9Un9hOonRa8JuJ8+jvB
ZD9TUL8yPJHyydEJylY1ynjC/Bk5z30xbxqYPSrp1ZCiINFK6DJe64N6ErV05JdzbjSBve79OvgG
WHp6xBwdt9XTxnLbZwBWuL8E2YDkxp46zk33k3YIJy6HsgCCbMF6k1bRL0RdWKzAlqeIrwDeCpv5
GpvdA01Sg7mKO3vr492GrJku4BhlJGLv4ORH0MgO1kTTQPFMxqZbUREini9wVTxFI1zpjqRjpo3Q
qKJ63O1MbCAFIms37eacD98ztUCDA5d2ykq2SToZfOvDbPDQqgjg86BHcdnF9x+q0HRyaHznlh/Z
Pndc2J3S4FPGiRQNDvjD7a79Bju1eZffeD8fj6n9Xh1KBr2YaXIQVh9FpalRGAb59POnBdlAVqDi
cAt2GhXklj95em942SJ/sYeHx92w+K0f06Rj4LusKpQ8p7ePxv6BZvQQvLOHRoeUzZI/FHRJ0ZHR
GGYviEHkuwKsGOEPNSP5tifloMpQiCoixBKH7GAFxvUn+i5C2fgUtRHHcyyodw1PtwGUeVe3qZTm
x6R70SomJj9XNB2jtnGnvjiunJypzuli4Ssxg4/jms/iXLPZ5X3PQI3caQxZbulw68O2V78dG9yp
FnbINpWDOBX/IpRg7aKNObXgwudoj39iNZVyLzFBydiTw00MovrAL2Ea+HTWMak4yi2Ee48Za+6E
xNbqD39RBrwTVJZRwah7z3AqX04gk1hdO69L+qmUtJtJc9zUNST/rrM5MTrrlA8a3lPNw001LV5T
MkGfApxexF/VwHZzZpuWoJDPajQfmMXEJ8fBPHhbi7kCGbTEcHbGtVvvmmItDzT6u4cQAe4kHeJ0
eo8WzhoTMUNMsk843i+8oevjnvpJm7dptXdu6vRjzgpOFB4MpkGvE1cNTtHWdNAm/QDQfSschs5h
+ds2DbWUN+rPmGdT9pLF6h3qopHCmk7uEzonGe08g3AeqJP6A/CTA2MjzZyp3OxPzv4rBLnQnMhZ
dOcQox++itjCtgJJ3g7S3ouelGZv79wqA/dAgI2cD2bGD1XzPVw8Mqi/lKZynrYQF1/IeLAJu7vm
dRH/g5iBlUATAbMbLYUWxPjVSgdzbZK3FvjDD6VQ5TWMXoE3GBnCDIirm8/WDpRY9oMzFsRlsSym
8L6QqbYv5fG3zGOjYEziYmaL4/d8oC8EXTPieYwS1JGklitzIpDrqWjJ3Uc0MOAGYl0yTHPFiEcd
egS9deHUWpU+6JJfoO95GS+szJ2NETOT/zD2ZAnGXKSEjzRk80unSGltOASPi44fgTKufl8C+472
/1Ei2kJvbU1Ho1s10REb9nIosrHkCIqq+XepzugbPMA5F4NNqO9wBIxg8iDi+eikwnVZjeDgNpQb
qedbTg3wZWBfT+PngUcjUTc8brcogRfkugiCii38SlceplgRy8patxb4ag/7Swf2XBWaX7aN5+MI
gMrPYGjk5v5dBi8JhOdDa34wmY+HkOoZo8IGIZ9q52u1bID4MEZLUUWQS7auAjCMZiLTVd1sfJC1
EtCmpnT8SPiM+T71yM04VKRMUxpnmTmQFrh73DvLIjpmQBN9k+nyQcazRru2pqcaDHofYhx+4ikv
lTIXqikJcUYHdD3ZiMq80xFg1Ar+llaWU/gr00Y0q/OeBncLcffFfOegvyNpuPvGw0hl87Zo8WAM
3CqSCce/b5iKOywo/7EdtqEDl8nXwsHQhXTnd8zZpw3n4AZO+ihLNiSqE4iFsvJGnq4j5iiOGPfn
k5INGp8ZePeDpmlp6Hp7KUFGg3JZTZPXz+1lJdNGzZyYcVdXcYGa8Z/1U2rPmXq/slCDF+gEwrvJ
+5d+b60QVCuOnrx0lyEG7u6v5uXwsKuNscMQ+yaKP7qM5DIwY1pglF8Q5wtiJE3wd1V9T0GKmc3p
Gw6EiN9nRhe9RmhRS6t/aP3Jg3TGJ5CFRbfUT3467raWXGkdJ/kdYL/UJRBeZE48d08UKklgGH8E
sxaskYxF6tvc3Vbe09qPTsDy0nlomAH1hRxU0N7X+X422jn/V8MJ6V92JJrL67MaF8haPzM/bH5W
GG3i1ZPMHn52pUPpc0npULn0H66ScaadVlx94MKLqSCI5XLtMpkGcKIu+MelivKsgTcYxxH9m+Y3
LZAluLszddx+R07eWCujvnSy7jLIPhxFCFe4NvdM+BHw0fpfB5DvkA/QtJnexG3T1Bo44UdyFi27
vIR6o/4q4IVdzrQSKl7mfUK3Scvwwj52Hb40/8G1NqRxx2dBs6U3fYWIIUnKCC9IT1tZipeprRpA
OM75rCWJFdCTIB4VJbcp4M5Nw8zwiWknbSrUVuIk3M4bZuJ3djMalfJwqX3Qa2SjUrlRTGfw/ah+
65LMC30kwY02yoq1zPc9imnYMHvG0oIe05yTFmz35EVMQ6Oiy70jsRJeVOFj5pQhXXW+sk43Npoi
BowseYpLFOAkQEgIDaBXwTxzJ2A8tzkephMRfQbUG8A0pax1qQHuUxklVmzLC9LtSNRZV1NM1aaP
4GM2mYilkGQyhwcQxLUx7SIHzdenyFnVn4U7K4wvQV/qwWM/Oj5jRjbBDjOwYY/oMTkZJ7xOgo1V
FuzryW0o1i6hPixjgiaHXnugFrveCjkq4PiS3lUFGLbfNHncLPCVeWBmyOYPYUYYwf8rgrhe2ZxU
PnQAaDIfZKPSudiPgcRbB/8dokno8Pa0IDAc1xh2eiICkDClOhHDE9k6eKt6k+HzhdWOBFBFInH0
PusqefqQ7KNgFewTIaK3WaIyBkGdTqTHcPQlLPvzoTmucO+DReaqDXkTcNwBsd302YJkqws/cc3q
zZ6qoDiL5FzvkwyME2vQdJ4hs7EgVr6b20xNDzGhXoeGmWUScS4un/PnMDkA09jOdNK9BCJQv4wO
LP2mH/9VbuDi3Y5knqjDCnDgxLaPC1fJhjolxdYaSAC70RzTi0Hjp4itQjiYYx3WwthgfJPqjrSY
yBhJDnNJ5J9QVjjRg8QksIQwJVC0flNSogfJ0lTacoSO78kzbxIjm4CLNn8tmIudpvHLsN0M5k7i
TY03UjmiNiWIXkxlyo6GKphw1sAvves7dGiDYJFVNwRjNzr5XUVzv8TkQJLTRSXTjY4cCXlH8as2
G+ERB4myvZpuk5JmZkgWaDCKKY2zo+p8JO5KyohzIygIg0sYzGG8Xl6oOoQmLCz/tXqsIzAEgPEy
NArPLgo7VRKXo1winRG0hbaJQcjHDmv5dno5gBX/10feD5oGfYAog3SZo35heZ/7uwIU8WJ/fDhT
C6gAAVmia0vr4R4BppskRo+inUo0ChaYOpkN+lL8xLgdieTlHA4WBNKJbe5shAr/C5eQXpzagxNP
31IfYAWE25L3q7mU4iyTpXaDJnZTWPpmEtXFEnx4OKyDYwZi5/q1WPazt4ARrTaISZ01yRK69+h5
PN2CXvhIIXmXsldQZidzpvlxdvucrpbSCyCu3gdBPx30tKftUGUEcb+AvDHxBF2zAEcWwXu6708c
AxG1Kh5FTdY7qeH6/NvlmY9TJBCO1WO00sEPcwi6j+RPk2mrqP831JvFY8dfB1lhoCa7H3ShFZc+
urnB4r7lUKNyciT+rZLzW7sy8bk5HGy+z/o1ANQMWoIFEanTEj7C0PijsQ72J3BXx3c683vFA3Wr
vxkENh5cY9m1lMEcuFQVbRr9dA055t8FaG3QHPYwAdHrTuYIs8Ri2PH0WBWaM8sb4q3Iez7xQlbC
WCbIY/tnlMtrSv2P+TAdu15muRj4x+fAWFzERjk63XPYJ1uuytEYZ36MaBHvnGAQtCqfa9lY0nn4
gedaLukkRNmVb1QwI+xhhBnHiVBARpGdyXTRkaODDTF9IanMGOtk00MIq1LiTJ6nj6fJOWkiHg0x
P80BJoiuPenMktpOQ26A6Yj3KQGFgOr2BpuWI/xXzqq57cG67/pn7cF3Ml5KIz8C2bKDDT1NniaO
MIEvuXrMvuCqTFGMeRqNW6nfibgg6s8S0Jkv5KiD4sgnTpMCRVEZpXNiYNsYWGROjmif3wxVuHR/
pJR5uSqiY1KIqw4GORvLDuggaZ68hdLpAKfpxAx++NYX9eSKbmmnd4MGM2Z+xk09a7poUTD3MTlT
sn2TPMynn+M8e964RN1gAzYDrOnpYFm/v53mIKX3+y4iIMNyWFgxls0KZlSXqmYty6gnmpO5Qw4L
m3KbT4SnD5fonN6ta3ZvcWmBP/r1qNyzDCx3JKQ9ZprN8031Ox905Tu2XT9H7vHMhIZAVOOuOC1e
PKYCJhOquHVsjD1tUi9vlHAryNU7LksxEdL9gz/VTtPL0f/CwprIP6pn5T/HjqXxLDxc8b9Yf4Yb
vo4Xx1n83lntsZE9IlBlLFOvbERZOGp77mMWm8RMJFga1IDp4dF71BFJUlYyfVHc1AIR96rHZGb/
tAIgqesrCL5evq0NCf9X9wZcJr17omkojTXAf0uNrrb3z30rBz8wKHX/oRC54leDTQSwOCywxcDp
C7DXnxfgjWUhB8pMg+sca/Di1g/sEdNfE1Xx/GwkS1jUKh5+I+OnfuZxnNuLCI0OpOIsR1xoiR6q
WTe+rdvp7Pd+lOtGKkkFKGDLPt6zyWjf+9DEzWVvD7kHIRQPFH5xN9q0k+T5sKeKOqleCqysYOvf
/3O5t/2eOGY532cCeqf9AKGUVGS07tHJyDRvxWXB0vru/vaPgZD1ZrExQadz+b1Z/HDwCcIDH+Jg
uQqgp5Wa+MxrazwNaDFgWwWJ4LRtUaWxWW9/sdcQGiTy/sEU3Npr3qyDY5f3AHShzpZoZw4GenYr
Y0gDBmBsCrDlEzQfrY1AGvl0H0Y22VvvJYreZx7gdyNHpe1LSM+Dp6/RBrKcOOtUTs28U15GAMlj
T/u5BWgMs9F3mn6gUxvmJbxe0sPHxw4xdzIUF3ubdd39deSfS2mBT1W4HLwrhbHjxG2zf0nIpg9y
RaQ4BMKKFfnvccrlElQJUlpUOEEmPuTn8UyFaR/ZmbMZisIzXxYLR+3DN8uV1h4XcZOVB2xd1LFN
IjGdWNEnkMafw1NqchebjySHMghzBMzrn6VwooRoY/FBj5Ocj+4cPeC2LfyGpTORUpHgcsB88Hcl
7hur7ktAUwZnHej1dSSkQ9JOMu/KjHfl6L0NksRMTZvCNmBBCAuJf9ltKHW3XnyBDgIGiLD9nPyT
K0RQiGD7DUDmICixWdWCVrzHy7xtaKVb2lhMZet7T8AjTClrrf3CvrYbMEGgIRkPSjnVDT4E4s+j
48ga1qkpGYZyVXP4Eg7QG1IGEWTWnb9P9MyPSV8+TrxOpnmah/snf5m44oVuxb/3IgfN/Zb2yJX0
35t4ERL73Enb3C10haZOeTjvk8X8w4LyX32/xO0DY6DykgLFedkGzMgnFV+Nxo0leSKjOSkdrumN
iLBhAPeSSi2gTfGenY8NMm8WbgWABaNpZVehg4GQIQD+DUVMjhbF5t+TTAUVepXD72VdQ11QACdG
6vUobxZXqzzxheKcFwdUF9a8OHdcOKE3MqChnXjli//tox59wZ/6xRdTmKI1a8is5l8XEsqRdeM5
V99WMlFePsNnfxuUzncRKW2uiUMmuMzmqviU3ay8MbT4qs6iQNgxzem5kZqdF0QiitBWUMFCuNOu
K4wlIo861t9xi1lRvFyZn5HJuWFxk2VXqsWUxmlJgG5JPx08vZLjgfKm8BG++jVw+S/DgUiG03CC
MKsJyMWw9jGYtAKQNdEOeRSQ2WWB/SqbZaswWQh6lMwvXSFUe7kwWyfJLZxX3Dx5RcB2+VcMqqj/
GQIdxa2yPA72/NrNr7KuNrtOyjnJWiHBCxf+CddQbFPxhdiB8CzvjkinqpOOE0io1crO4AiOlVkJ
mPKgx3uExDrQ9o8noAoaZboT1QjNGNfH91VXUw2N7CiwLyaDF+zUNkI1ZKfKdk6sAezBr/skcqdj
Xh3iWT+aFjZ0b8mdEdHP8PRZDgvE8PWG1pRa/utiTPxMFjpp9teGaJX2kI0IL4lr7wVf6ADDy6DL
ZJX6UUF+4/XyeJf6Dah8JD26Oos8D7VRMWpqCbume4y/XZHIwt6Oifro2P0rqny9yuwwxcmAI1JD
8ivj7JLZaPnVu2atr1B3MKa1NleU62ErXEgT1fj4pM/3AM6w7RhTeh8M9y4COi/5GUfdeMAZqAzF
pvSuBAAbUyE7uGs4GdY/Gwj03ioGheaLywKKdK1bFo9oCUYszjge2b1qdotHhBev04zxMnpVx1hR
ebhxw1J9DhyREp9q5Wco2U1BZItYEqA+yYYL7bDUoI3XbNwGegok4aafD7mQfVT2Fhk6jcZxQPH5
JPxwh/yxAWvXJUpUaOQhZTqW5iLITPA/7P/1E/hbmFDND+ok/WAE/hOIq0VozWAgItoMAWr3+Zwq
1mp6/28lWgctdO+EfyrJtPwwiDRqzyTTHTM1c4gbGkKHGh15AIVHkuIKf2QYZWIwv6eVWRwunigp
kvXKvM7n4ZmUdrI3B+0LoxDMDBXUT/2DXOZA+8adZAXjXZH9ubqnvH2W5LoVKhDZzb7aLNL6FGoB
lvJuLjRsEQQlxVEdS9eI3blasmOXnkuQhUOV+d/HNF+sjiOSIp5Fn7cY9d2sRwrHG1QBcbKKJweC
+fQwNZMedI/v2sHZGql+wphyXw3OLLqswu4U5cn8s4rR1GvjNHCkeb3hkl1+NfxSbg5qf3Stsq9f
5mjvpavqXaTsHSXpZomv9o1z39KYcdSOa0X6x1mzwMwRRFdRKZu/Ahx0eZhXUa7LJICbkGOXHjfq
EsXayLY5wY98P1Swgc1bk0u+yqBha1JheSgVJK9simUmAXzYjxANwb4SGRR44ZBRuI6riX9UyWxe
ePLzNiJZLJoSY8JEJdTkAa5JiS8k3FRyIEyVaDgflmel5oxwbOz9nQwAv2tpbzmLsijzGcsOvIDJ
4+2w/3oz6/3QthTGvJzzgDQwgvM5flIULWA/fHn+dQlN7zSOUOWXJ0ARnj6vMbQMtidflzqYOJIB
yWm/QfmhpkKC0AT53Za/lZ37QJ2d6QVidvLinfGY5KH25rxpuvGxLjwRujzEviuNnTcjb0uP18GE
7uwN8sZKhGaBmQsG8CFubZf8yeSSLe0YO8kTsvlI5aki0iqqwFLam5uIRD6XeQiPsjlTzU2bFzWk
D9adrA1sdgCA2VOWahLW9dpvMWTfFXEdQAM91XiB5u0B76teN+917ynWTnhKKtL4rZP4GduJ+1BE
j82582mM+tqaGiLUtovUUfB/WZ4Onc7VXQ3970IZ3rR1AZaIbAm64rmUfoQcJy2mmMmS3mFG/Fhi
7W75R6ac7wp/F/mZ8KgOKrxCx4O/pPVrI34MBwqoyyJcFvX+t5809zoRFwWvba1hKJQx96T4HpEp
59FkxisxNrPnS5hgSDJWiIsdiqNqheny8VwCZIaaj7JPSWL/LPMhuemyRw4DIf+q9mNYuW+DAggi
FYltEo9pZDTF+njcDeRdcxb6uy8skzsj4Xm7m5GXoJu6R6cSdfu7Acv6Z/3LBu/i5d5JlqC5KIHs
qz4oeLZEzwX0kZGf+2Fp0qbjRt62jVODoTO9bx6EUKdbNYSSf10FDyDteMLcJx5pHqIfoV2jWVgF
fjBm8LBnYpsztuhT07at2M+0qMCs8KxBHG6ZLe2notsprj/g4stTAmua7In2YbCrqOC7Mb1/ROrf
SQHqvRGKl6+hUORexgyjEElC98bj812Vo1lZZhu1rj2w3YFpVp8fmc6H7irnC9JgQ1im+pFhM8Dv
unDDx7EUGARjpPLBKc65J+yjbmz8i3S6PL6lp3F9l8wXB/Tj4g2NupU6SyVSBgFQGTfgHDOG3NlN
FVMHc9VgM0m9526qLLF85E+Lrah7wMUU098hgk09MSkJBdtgGJugzqRT/4hdw97LYf2Q+05X5sll
7EpQUvQAFwZEdH5OZpObeutRP1uJyzJjQIpUP+eLFxWNnYkc29Mcm67GsHVvqO+ThcovSNSIF3zS
wu7CibKpWrXDOzCa2Lasu211+q0iocAiOqAP228XJUU0lV2oSnKGvYbijgE9/hBRtE4XHwcYpBc4
qDClW8s1N8bCp3gbOMOusCDBXj8blSgDPk964tjM8cKkho36HhytTdylFGIlUKWRhhOECKg4aVSH
anjxiGOOYmyXRp1Z0FpO8xW5RvDf8SkA8WHyzHyH55zwuZjrx0/zXcIJoHBlqvl4hQ4Fi1lXGRzv
/L//Q/dDvsyzeZkWOabvjbno1hMXsYbhgrAeQzAIutm+lihkOlDbS7rQ+oTP9F5Dm/1vnf5UD8HL
aK9KN7nlB8Ex1ITPv+xsb0Y6SwAzXXu071y4tKQ9KcOHR8EE6PhaTymYbm5uTUmPhgIwNk8GtfrI
Q6BNE7ANmY6QkUAQbn1GK6CLheKfVp6ejIi2AgvNsDTDEUh08s/MFZWLy0SQT48U9bL/ZBLi++DD
vS90jzoclbCW4P7jK1YMUnvhZFjxOSoVEfdXxawjHBRXwtN4t7201OGZprTdaHx7HV2DAdWAUZRQ
r3ZJ9UK65xA3A0vW+sfHZF7o5SPQu8Mqw1TbTlok5vpImbjU0t3IiCq0wd/ncAyC8LEavQv2N+zq
0KCzxmn4CK+KNE2CELwwWSrqaS5re2NgQOTpvddULhul4XbRuvvqtstxzT+kGjNlW+YAKs1opNxG
hvcD4jEx+4R0/gvZDn+0ySzxBqIIMQ7kwiXgi0uLppV6vDD2VvyAO+0BvzEmqEGhsdUaMAY1vIfB
EQOLmscjxHLMaPRJf7d25Ytu0NHc7jfTlZ/okD9zHKmRX/E60uycGUAbD8nmruiDUA/BIHXGnPzk
0L3UV+i5eaw+k3y6bFLR2QkwJs0RwfhTsDhXDUJbAwGbV4+pkPPLBJu7i1VdH8WNrklTkRZzwBsJ
XLvjiARUCZIX1RPaqQ5JXbUcc2IHXp2TdQTwe/r8Dg491eCi0DBYXQwvYFOVfehRpgoqvdtYTkiE
Da52UV/iVBBPlm9xUPLBYnp5h9qwmfiXoJAgbPGRb4MfhQAedxMPpIB47FhWO9EIEQ9fMN2cr2du
mape3AnG82fdNsvgRdVQehmg8oZjFmkbr+J6qQCHnr8HAeJndpa2+d6PHkA0KCvZnEo9bxtgViFw
tAEOHvBSPBfzmKhCH/2nALglfuqje5N42SNba1+Yn8eSmQb2U/E5iMVqAp3MgnwGpZ62JqxC4hkj
eQe4WljDt+bXizaLmfKqA48HEdd4+MIXezFb/YaTxy4prmYnjK7UmVUPeEesrd/Oa6VzR0B13Cu+
7edmkrilefRmg6fiO2RaiTCx4ATnMFfZ3jSW0e8Of+lJvGUVfceTvPgE/hAxtkW/EouEfIt3d5Dn
XsO/+7voEuxcl+ssVJT1hGQ79n2w7eM3mfTr3Ab9AD+pJECTLmvMa4yCv7n4fRzZqPWhcFjTYXVu
xe/sSYFXIhdvAB31V2KN1vXBrFpaNzCGf7ysFZ3Xdeta5aIAqrS97l8lIgxV/J6DYOlJD7VPeRb8
WpOe/CQqAu0velHll08fo4Su11XoMqF1ACouDfY5m+nACUSQC2smQ5eKbOYR0pjtVupZcL/oqnAP
G1R8FNE7JdKXe0VkZaUBfHdvR/fYDu5wANwj1bUibqah03mTWYY2dEXDOPDHVbfRkC1HOPGXirRB
IqZfjbBIAvBYp8+NeO6wmfsgwjuEjLQH6cRJDdTC0+ElxYIFalu7GtGvqWJEu7lvQnxTvWHIkpoC
ekzJbP/gklq4NRuyOjJ+sPAhCHsrf5FMPQgz7sFPjJZ7DsKsUNFwPxTw5EWZL47YDE2dYd85w6Tt
eEAFEYznxTpSz0LPeJBKgTKFBwabKF/3ytaIYez7dU10ooYogm29qfqiXkSQ3TbcOPZ67SrWWRkx
X+4OJUbtHayVo2pjtKLgG5vd4esMnTS7SodVaQDJEk1V5SLimPiaTG/n3ua0uAuDwHWLwhjnVWkv
NnZevThcPKVy6x9L4wrfGKuEH3kAr2SZruHFsgHpi/PRAoRMLXCGpLXd4HPrWAshUShe6ZVFBtNj
+IaYlWV0NCZnfSr8BkoR4cz3fgH2BDSW+nDF0GmqF1TZJ3yEn0wgrHFmCbDLhV5MFGzHsIQZ+FDe
2KPuJLXUJ1cxLBBbz4J7OSNXrv4s7NnruxGJL8a/c24m/c9c8aRJdax8K75OIolYKgZnUqvMcz/a
dxKc5TM3ASVu07RkSzfEZBiZrlBx1cU8ruwXScr0Pk7YvTCvrMyLeSJ8x83kra99cMyn0Hwtm5Bj
+K7Nsy5KltUnhDRoBT+X8934fokEHo4npD8Uud9tusNpj6N16EI8u8FRexunR2A3a7AQWNIVZoHk
pYDQN8KJHhve2zcLqU7cNYe10ZVPYhF69W9FRkc1HcYQxMPZN/HK5+GG9WA12AK3fm03AWI12yr8
sEhLimOS+Ta7fub60pSUmamuYhY6m4gBOB6JtikHNbvdo8rlI4efgdxRwlG88+wFzZo4vft36vwN
kg65b1u6ln6tar4Oa3oVYdtDNFZWRNt/S+6+ZkjPtYOHP/OyoIXNwah3GX070zs0DY0S4Yt7EgS8
eRV4mc3pGKRhBSTdCn1NDuidD6/+j6AshHrws52ZBvZ4s0XvOSYmK7tJ5pd8z/pAR0beoYa0SH5a
zOe3yG6gH+BA9CKJgTOg2n5AJCmztFgIHAI2akRHDn+OTf7OcnfA+0TOcfRUwoPUEChNkF3Ak1qM
2gC7q94E8aVtJ9W1oCX3U2xe/liaGhp1gWpZf/m720xFo7ORfXyVMxVQTdJ51ptz6vXMx5d2mfNO
FxRXODDTKStMaLeWjFhWGOGWknmeCJd6KLErahYhaHf6MniFMVM1sQZvRG17I7LGfkPQfm3gkEVI
yhLhm/tRbtqZRE6IKWQzRO6FEWZQ8bsAoZz2F6Sl3qeTG+/X+ONny7rOarZ6qw5mvs0P3h7lwmS9
vS96S7VkuknBGF16w+oKl9xPPt9awSX/7/IF63KD0rlHFMo1d8XLY3IxRfx+y+gp8xVvM4nZiEtq
ECq9F90fz7skdBlHQ9zLIIjZfenVchZmP1IbGbqGPm8phrUiySIy7sBTfDRm3ZZN72AKvzHBfcIO
kqvBVgXjoUPhOWhWWMbjspRZCdwGngiMDqjtsTL/aq3c41Q/TN+O9VUyQJXlBgfzG23JUNum5rt4
q1iKsIvXK0AGLQP2R9g3OvGcTnHeqG+IU0Do88JKcSY6mVWFLpbHsg6AILz0vaWciSQoFa5tfse7
anpnYr8ha6bTojI8ykedVkbN2viYOzVI4TfgSSl9G74b5tKG0wfEjKSUQhZT3WqNix6/o1M+btug
edBvl3RwxXqWuBk3PCwqLzO0n17ZnJf4ozrlD83Czgxe3qgOj2D57HBq3Y69fzCT1BaP1Qd/D2aC
d+4G8/0A5p1Ez+4rjGuM5GrATtSH4BSFcN6ZFxkFNWNdrMhhC5ad09FYhM2IWOaQIrWNKTcEGzyf
o4UrgeBixAr7rfaFNcuDX7mw97JMzgUhj2SyNlXeJ3lee+hTc/9e9QXFrC5Me9KwcQcoCu71s7Pv
V20Cn3CJkcKKZnSF6LSln/hfbM3my3jm5uA8pw2bV22ioWV4P82E93EXK0iLyjZ4tcfk7k7qJ02m
17Yi8LuvV005LrHL0PF5djx77lSiF9mnWg19JL9obvJd3sucB2SZF0Ga1dt/j7lYAWRBe6AKk0p0
AnpketzNl8PYPVp3LIcDIrY+zU5Rv/wKqglIBV6eB/MMesnFR+0zSfrlDDhjSLnWKSWnItuFy+Y6
C6bP+X3HCRFfUrir4/0bG+Ap+840ujj6YKZSdlCukoLuwSwIrML0rCHtA7xBwkBv+T2+6yGLUR9/
hVs24OETczIAlkQz08RF5UbckrFgi7MH962VBwd26boUaLLFe7PWl9Qf4s5xOywW1OEYDwgmRJXL
+SLMa8NGPqygjCpLqSLPxk5IWuhKnhZ4oH9AuyEzLvtESJtHL/vcW+ehFB/tzkRC5mvSmvai8Ilt
Ag//K35SgAD1JwmHrUZ7fIDZvPsQKTRh2PScJVqT1WoDbi7PIZGgAyXVMgBl5I9LsUe8Y2fdf5/F
l/YVPTPq6Ax+gDwUafrtvrOqzu4KHUy9paW31Um6rNqZZ/6yJu0n16KJmEt8Inye0L7mYqNSoY2V
MUfMbt71pdYzF/MgmiiHo/VHDVosi7OJD53OHdTRykQb8U2agTvydeNhYolFu1DuYzwHuOxLoGma
ijOs6qAt8oMTzPSiVTONb+CsB3LNFl+8dC+uyWcXb2EzYe6BnRhuxVE0U+6M8hBDmFvKDnpFGHUI
fcrAxqn70gtPu7xsAG/KUiboSM5pKM3fS5eOGqQYDiExB4fv0LsQwVx7kOV5NMmQHqCGv+UxVrU4
c8nkXvcQDrf3CCxGXr2KUnGefvcHXRww0i3TKayPEUlt8f6JHofWlqYo4Fi0h/axTlQPfX1HRfkT
lDEH7fp0rLAOWgqm7AeVtkdrU3Qlg6nbRL1zo0rdGZxQ7t0DUeQcUPXIiznf5XJ0POTZh9KN46oG
Qa8wpWQFmwOyUA4xUvMpDftj9PajWhE7+f79ewd3eeFuXiflN8Py0rqgBmxoAgW896NLxS3Iy/hA
bOIVFRGdZb+Bmokx3feLtsuQ2xfCUsIiHFTIW5MH+IGjEJAroFY/K8sgCTg59pF97PymDejcKYlR
4OPqp88/I6nU+4sZDZ+6/76QyrCoeRsLWbW7ma+YdW9Z6qXlRH7gRFCUQBltv0vjMaU/LNi2rTiv
mH4ACLcJ/Yn/Wtit4+zeajO6vzm1Jp9wZRZ9AcZ1lowxhLE8vQSbi1om7ZuTWAt5X6FGnZtn9mGM
OLLtf7vkEBXJAppsbqc5k75dtirPmvTz0kjw+N08ODqRceWliEcYLSXJVA98NhLpCpBSiViFt0IK
PV9Q8qpFpa1oLKfchjaWs7T0O9xomYkrnzA2kBqEZTl7EJnyCLZoMkXKtGtZZJ+Q9NvpPgUEpwGe
tZG6zbseutcIPeGf7XO9eX0vvxKWED93nJBF77qlCOm5OWuepBZMkgN4Zqmbo8rLkWnW17pnzFXh
xU0GIRoqi0sdWdFy9g+4QdtfKEjW7XcaNSSuljNeLCqCMiE348NDOdTd2SsZSCJ4IoNp5bfq9J4E
6a5vt9uvnHE8DNBC7sRXQUKz8SUQKnNlzHxt6yllBdnfEwCM8SHHHXlypj3u5/qw9HjLw3axM2hK
9qc897168KmPAaw3bVJCBC+OmW65MJzSeIXdSNFZPpYa1jDaqI3yvEDmfKa5oUYxYgCC1uUzvI3a
GplXXPnL+mzPnEvRmH0+fyDtqZQCg/gAErHwNkAZbJAwq/P5flbP1R4ylL2+KThNjz9oxOw1/bYO
k0ehfqWMGaGjZF/aBnRJqNmzAcJl4bfw+9ZEfi8k0YdGQ/CQx9h5Ak5s6/npyBLwjn0XOAOxKWBH
7+cBc9YMHg4ZYEQTnttX2sh7ydHdNVadwubyFqzVdbUPMjmYcDHX7SaYn2ES+h593/16Wl8n4hGV
HO0edwHiqTSdTWpDNStUZhy04Ye37uvp01kZ9K0+buz3RZJY8lLW/goI0gC1CQpbrmlDn1SjX2W+
Le7btI43nJHhQw8YgWlqMMR+8Y1qQTXbyZS6kYiGug7Jaq5vfpgRQUAjz80BlW5WJVNAP4wKxa7P
M6WxNGwSVIfWonZ/lHKjfSudi2XAjGlUNixS6KcmKbcdQIVrGmqYPAN3DPyRipNHbEXCv79X17ru
LOum0MAzlmc5eHnnnndhxNA167bdvmS24MTMpReC0zL506KnGYn8jv4Y5pp22VC6yFHaP7y5+jQz
8c1Gmk4vCjeQWiyt9DiNELeQ0Kd//Wyw6DE4rZURN94FJ0pCdPms+CTJFmyNwkW4FsdaT8mTPTGZ
3cFoG61ly2SIEQXsxkmOUxrQRpn/+I6VRsy4/hzFqjQzIua7sAGogf20gi69/NkGmQtOPQEk0Kmx
oeDN0RyKntO4aLK2M86wOUdpAN6JT1kWLphoETpP91rXJqJPbtZ84Nyl2KgQG8j7xQk5trbickq0
7Z/yNLykemxc6626DrC1NaeeMHX7ILvyNmHPeG93cOFwl3xGyheHRkzFcmUziXxTsn5ngL4+CQ5H
xauYEvW1wgMqOfypNVD76rrC43diuxRQALLmXHfpZux79DmNhOnaUbeX2VsS6yBrNVI05flCOBDP
YxMV5wxAekXobzukf7JNqGWLkH0VYMqatxXe79T8f6XgTlcdT66yawEpBgg9g4o99iAGmx3k+ghD
4kHDh+sSo6Gvb21+zb5m0nbYseAcjwbZkTk5+VVOArnjKs6MrokAxGO+g13A2Fn8MxVmyjAaawuh
SrSBgAC3Co3oxCR0155BJsorBqMyQ5+rL1xBTkxry5oilITXfSF3KqIlFIJ4u1f1UD9vyF9qOEc1
faoLl4iYZGEn3iM7EjyYP5sXc/0LaH38RjZoEDJSpd7R6vfZfWukf2GsgcQPf6x9z4EYUvBROmfb
mHXhAO2W0NWv8Uj5Wb8/8JdlObASjPLFi3g58x23KnJY5Q1UmAYyh0QE6LgFvUCyYJGbfzWa7k8i
8776IBof35uL7UxR+9vtIkWaMTrl14XaVG06Btz5ag57j/uV5j8zCX9IvYyc/omLxl/iKkGLBAbt
CZXMRq8B1soi2BpvwKXGTlS+4HCGn7C1h3L4NKGpAwDIs4MyOzNMiYcidyogk96s+8zV6Jtar7Sv
j1dvvjmBsezUOYHCuWsofLJMbIrh/heGu7PdkzOUeFXNYFYAXlRVLIBTz2pwljJ6iPJBEihAnwTB
PoiftLaRzmyxOse12Q//N5FYF67ruXRZlJh6K/Mn3nM6pEOsNnwgu+AXajKJV121XPiwzmkbzPxn
+AXsdlbttylIA+88eDTXUOmxedjJhYDhWPbfZ9+6PHro+BlvDHZhhv+3WusaGaUMBHVEejqmnw6y
rx6Q7Yg2T+EuzRDAxJS7P6fPq25n1Mz4QMZ2srd/NbAO5gzc7b84LZ5uMh7iM8Rid4e6U9wkef2h
q9B56rAMHFElT0hC4+9vtJFmOXae9SNIwrl4aC8Vm25UAAxj1UAZGHZ5mJ6o5l3xFE5pGtpM5NuQ
NTP6SnorVAua5xRMhlj0nXxfqonQjnGFpozmmTzdzve35YkoMYkX1SrwueNeEKfRtopO7b3pjPp5
tGdCX6WLUp9Z0UKC9rVtEX+GGKuOUYIkshlVK8t8Djwj7ZfnPjdcyAmeoMwKqMzOEmY827oNoqO0
XznnGrzTnm1gOaJP4f09h5vPffW47fYR6nyEzFnYjIMXu8HpOzqSLKC3xN2NEUQgqOgyefTw6Zqk
H3GDOGdp2W+KudEnLDb1fl9wR7WOaFgE7LsAkKp6gSoBfTtx0eJnNcqUwGwA8ZPZalwiUPWnVlgk
lfGjPG/Cuwzz2U7dA1AghsvXPRdR1hUX4Cc+I2rLME/YA0txHEJ6PL5ZotYLZBvdW2N77qg31AnN
+K8eQ0yldQou1gakA89q9AAMI1xmbfv7+pKfNkXcfXlzqTm4ciHInqiDCN24lTBgBpCgNSKurzHg
D0beSHed39JSWcj2TtxddP+fkEdX7bqx2WrwZXrOEQz9wenfVkP8qE0LjVbFwDSTRm9wOWcC8rde
Y9IxiCnLIeP4GlVGqenZplnKUTWNQvvlaxfAJmKJ2opVKdYkjZ2JTGw+y89AnWueVoKK1/p6nT4N
rfa9LEmxKOwtqai3UeM+/kGTGWOtoc+zYesPel3igZgPviM2gcNADRGtJcnCU8xr4LtztqLvHk9H
qkN0suL7ak3KTDe7Tnc7M2Qmq5oKbL2O/Z5TWh0eYdReScnk3iXZ8/EUXYcufiuRdjd+SywQPVPy
NjkOHC8klk6j8VWoOI7chUdmC2dC7eAHfFY3S7sXpviA8Ze06srtErCJs/JD89NO67QoFsuUyZqI
ubXzfvAXsCps84KQ3gnkysRyj+r0SlbLFcfawaEvqLubWgpONYkVrUTZVEHt2D2gB62uSffBZUWj
H2c8g609do/9JtEEi8vYO6uxEHSh1L0MsIloTsH/wrrFbJKXJTfSm4nyCUA3EBzhrQ5LFzcGGDG7
zYs5h44I0tkp4xF+Aqr2rRpf25xEnjpu7NMl42kEGAjqUNrSZXh2z4bnUxNYENtwgmMfeMkMJNWY
YaoVsExBZ45OiCE5tPsollDsUpPY1DKWywuLOZEgm7Cl/nfDxnz1PD3Ca3kaUzFJkz7B720Ywhbh
geVNesIqnFb6LUu6HU+ASDnS5xwSYBJ2CUZVlZn76IuCEWf0ouFMKCCqgJONpGuKYL/MOX+vNXBi
kwO/7Kqzor0GUkjy78cHyM1IX5JpiZSYIqGl4pH0DMqUuco1PU9Ex/6DyDsATH1JC5C495CV0IFa
hCFy9OllUAF8GGmzlDQ7OSlP4r5PGward2JkvUPwopSfQKvwm4Rb8bOsEalejihVQr/pLuwlhr1I
xqU7fszfCDnDGyAztqCN6LEocjm4FHhlhlZ1XT1/Of+LvGCrVWJBobbbNDd79J9ZViptkTJNUAcB
K1Y0Ju5HwfAPFDv5WPMKphJsW0yC26CoPh7jF1Cr7HjSK3qO7VuOHBiKV2onwpMdcvboZOvgM6hN
tkRTC28QlJ8pu09XdmUeXLVsbfee2CZ52/HI64yI0RuvU4asT/auVhlkDxLt3bnM+rh1twcbh/+3
Mbj3kAmAqMnkb//ZsX6KrBtY2vQmm/NEtZ2649rdUnzUDgy+dLvztTwgZHaqIoILXkEWuSc4UyzF
rjjNdfo93YHSB+/TwHE1w44YBP6U9WKfsE8LFFWAh3g1J23vDQtCPgkM2bpgqgzDEND6dXSU2YR2
47CsVtHdVGLjJDCHW3ca1Z19gtMiDcyVvFV9Udo/xg6vouTeHoLoQt/N0xeaMc3kjm+ZGQ7pXb+5
lsLzO4YwWLNomGBPYOlfCiWMKdUg6IYflsgeIxIrr1Mz7s4i7vJnGsLGklr67ni7wba5dTFb9RQg
2R5ghG5S5Kof2j7tX1reSAmZZitGeQmkwPzY/JRNKOM3sxQCJM3IMEQki8u2yJKM8We4X+NipuFu
RePR6UxOKPr4j1t9A6tubftDHPTdeUNFezO8ij8QPAMA/9fpoZBNbipws5Qf7OPhIJ/l7oDwKznT
hBKVqtUAnbwc3VThrc+5Yar8R7VP9LWjMEJaZJ2/pAhuNrkGbcvte8AU+/5UGiNzHxZqq9fpdqu1
ZENXgzvrEZ5m8zCJwkO1D1xj2t3PCNOEGeQHxMVWmc7WuspmPdaMz3oWDq4joa0fSTthLiSdrtpU
64Krqqp5bTG3U091vAsTTd04lJ27hxZvOzgjWZ7yQt4KE1luzZrUkle6JwqILp4hfVVoApYDOCtm
lhXMp/u6cgwnDl9gTyDWptyTHRs9O0Nms1cddwSnydaoRQ5o4VzwTUwv5tGNePDhZ/JgelDwSX+v
FF8lormpxO53Xj432wu9WMeLd37GPDs4N6Y8JnYzMpd8wqXavQHaJvckVEzzm52ls0RnqiW7HA8y
PRm7B0fAP6pjwFq9tYE2Dcw23NaadzEdndg8Vi0hSE+lXuoBee1f3UX4j3Vkse2zQcnKtZeAsB3J
TrcXZl+6LcVUsRq+ckNpPVrCQ1aI3yf4sfJv5F+qqcpWS0apifRGqsiTsUH6NXCTIU7MCpGftjwG
InrlsNsT7zPItrCXdc6zviZ8QvWjjVyTfNO0+pC2Z4TMkAa9q06UFW6ep6tkDKzom1KwFmmn/FoA
dlX3Ipc9ky5GWDjxqagyEJm3N0pkdfJRQfLEDbeI3df/OQewgGgkCciyNt0cypadVAgx0LjfuZx9
ijOlSF8Nz7liZ48raGnzfm28F5fPT4bSqpYQxa00USL9Rx/pr9IGTUI6Q7PvoqHciDiPjRhMdaA5
cVMMIQfMp/ub0cNsopwhnIzdAg6AO7GtaoatynhFqghtQw8plqZanDQi4k9f4CR+LyuMhSMDE3/4
qzuuWAVYRcQKxloFhNNULm+iFYx0VFsZGeCjI1zysfdvDRIEYRvUXZOja6ggFbYFznA/qEZX/b2b
xJgLRj646JUpJ0s+12x4+lilaF/oNN+hll0Os+XvKQ0XTvC+XJc3UBxI2y/RqiqT7qr5A6tzmWvc
61Q+xPIlMzWSzZ6RmEMA8xEMU2KWmT+WaDOG5eToqyil2o9sISZaw0TJBNGm5FFFblATcTu/DyGV
8+uWC8bokS06ntUiNMZSJqCmw6lrjUXJcrLrn7J/hsIRxyGJIcAZFIpjTU2vaUN9gHVjCfvQfcun
wmLcPOevD7jV/1zbeGL0oiYYuxezdMUUrUeXxPdydHxROGDCTdZciVh/yQbZtVX5cZaJZypyqoa1
CsL+yT3fkx/Leh2CFsPA5TCNjUMOPS8iMPMKYH0XnUWn+eRBc0lnyO/cyZqGnAhykfLTg+5jaoxc
Nqe5CsY2Bxhrvme/0QIefRO98OIAK7VNiypgVDZYRzFVtgCYccAZjW3fAR6Q/Rq/1T4MgBtBWy56
caPqy7cbMQLd5UGYUTBHF81He8P6vj4pKYjau5Ri0dgECsB35bnp4Q9L6xjRYJgqZJBKEbLyoG+e
SBPFvTaV9UXkbvE6mRjJW40mxBNFalX+mmTwv2G989TrS47zCmkMEKxRWIkKcMriEFEAbSoCelVt
4xfY1RniGb5YQxrl5UnTLn18fUTLe6kRRGBnZkNriDI4O7dP6A/gJRYsKVh8KuRmoM6tggbAg6D9
l3kRQduV8ytDjM2y2xHWTvR7oYLsyZzOJ3GxV4wk280SKEdXxVaJ0H5VvLFZ8TXFVt6vBFX+v3LN
squ/SU8rmdA7keXhig2sk/C9M0Qov7MvvTUAQJNsKC38d9gDD2ldhjM9p+AP3FDYXlp/FaLwhVOW
pVrUfVgUlB8CLC78ciZxXHZPXGUeTjjYABkihps1eWiVey/uOqsKqLeUzyPnfECwAC5QidyovXzr
pAJQXI+SIYNuCi7k81kLiTXOJr7isRyYxpOVmRdLydQUvltXNF9050NI9cZ0sKEU55cK6FUpKstl
80OHOmdtFYi4kQYR5tmbIjDwGQW0nDfVVgdH4k/YM4pty+wT+q2z05zGEeIST5SMbbFL+heRi9+u
bMxqKbAApxgrGDs4YOmFmFsIYvE8u9bilcNW2d4v5zd92JnK9OLMTTm0Fp4xhFt4pBK1hV8FQpw+
Bh6Zc+Ro4zeeuuecGyMXJpgLxuvzNdTrTZRM0AskOPjNOsks9FUAX4D8IrFJPY4u3HdvT4Q6GswI
younAJj4Y557HhlRcDbv3+Jh1JMoBLfKBxihtUQGEbdY4FBEiQZSjSdjPj3+vdq08QnSroClGciW
RXi3LOWZBYivuDgpmHr+LcsM0+m3ljdl4HiO+7ZXuN/9eQL1JEewvAmGjIwNXUYrrf64cwZOSwcv
FwjzRgAKYhBAf5GqnTdqm9BDO6LASiyr0OCnIb9GwuroV7sOAEbwQn4QHs0TItGCzi88f1OPgv8P
ktUVarK+cZs1CqmqvDXK4pqQT3k8xkhqfNFFSsw0FHgBgmitbSHIw/Vukq0TOiRVjvdJbFpO6aeL
Veg32s5I1CKIpjzo7rbJpceFhz31+Na09aEDpPT3rv/FyL7dhSUnR56dxPvJ31dkbA/K2oHa8kr6
WN8HJL4SY9J/96NkkV52Rv3fhguIKS2Am14AiVI9y9q/MyUSNaigKFrA+f3u2ajXscRfkPbnuQ1k
JGfkmu8opRJrCuySdlM30xT7+wTJ390qTRuAZL5bGKsWxkOJfBgodnCejiLA3xyoZLqBgWV2pzpD
jk3NlBHM1u1pBlZCJUX9haD0qEAP+bVkya9LZqW0KTEY8aKJHzZF+ATli23uj0vvt4ZlUBk9ObzI
LLIDE6ihWz/h786Yr4IJR1j453w1iO/25LVsLvgKqaIrS+pYoNqHaGt5Ta/OxaDQqO9Apl1kOkap
rVtmu6HAhxp/tPkaai0YH14MXBODvsTig3MuPP0oKTb+/vmqLPufhSb32XzmkwEpsXT95ILHhuB4
BIiBuvgIaq4QcChk18LExVht7Jco72UQYtOi4UyLVm3JCF5NiOpUnodqBEIwynPIblG8rwJjJu1L
kvLayfqoXuXSLr/svT1AHgJKzirRGQ08gLY1apw+aN5uvNmpT1C+GfIfrXWCfXuCpAlVssLRQ97p
rcW4KWJtME8SL69QOzQnRxfAxJqWREW2w51+Ll163zLSBZuoTQaFtzi9nFRTESmPxCLwM6bTjATG
QNggQlj/e4qw4kDqKV8xOFyGtB0ZJUX4Jvm/izhbyC6SdIdTP0uZz2kjEaxaRXXZFLinFGLKVHAw
vrLaWecZM7Whvl4gjc9VZusKxnNqzNSFz1R/QO8JTbZByGlNg8T49jR22cFe+rGzVilGTmNmMxLc
GxnKSLwBZMGBybNKamzTcKPHeHnIskRMqP13wL5TIKYecvllkIEQWMce/jO4bqLcFBEVEoSaFCwp
gnn9OYSgaPlO/ZPsxgHR1ddpxi72lP2RmlLDlqzihEcNX6HbHCS68kvwPPFd+6z9MFcYvKJdTXqL
eR2vo1lpug0vLO22/7k+YqxqhnuzO93R72Rdpcmhyb9wGX7AprpMWdWU4L6gZFMXNH2PEF2dmH1e
o659I/gLmV9Q9T85F4mgBaqfZyUjWp7IvsBNhCVABLbBIMDkk4e2311+Nudnh4Cb0So8d3bH+qgM
r5KsO9ky3P/8l3sgj2rWH/DTblj/jm04FIDov1NUIZoEmJgmmTsnU3CGDlepnt7470iUOqe38m9a
vuD1kzyo6wblmKXW1TPTf7ZVR5N7XuzrgGO40m+mMX6EXn/QBzxaHeEQAwdMj7Ktu/KtlD2N2Pnu
VxY23kEckSyRSXA96qvr+5PMnAwWbgsQpvwPmmn0tyKdsOSgTvaxEeL66m1t09Zbmi3BdWvuCE/3
sC/G2ZhGfeWBH0mU2yFPx21kYEyDO5za3ChdiSvC2bL9UWWdQygaV4tnfgkYIps/INF6c5KyJQMU
mul58zOeUOwctkVZmy3Ogs7zpQiJty4cW7fMF4ldWg8hTKXzrA2dyfj0+AZfkoQBYj353W0jgdW+
DJmnXPo9ODq3MLv6cRIOh8aUxTq9nT5wWdth0J20E/SbLPRsgtC6Hd09egGTg0e5Zm9eoG9nAa0V
1aHDaYRBEvbR0qRy7wDm9sy3h3xVNbjKWjqQps/XhZkF26PsrPGDVY3z9NwPl6jVB+BTUxWH06g+
sq/MDJkWyAxAz6qSemCNI4pPRmK4OjD4ztw9kbFNPbDkounF9d88V/g40H7Q3Db4ispxgvo0KIpb
qToHI4iIKkEfLEI2IARyd0UNcT4UY3QYdbbZZAE11qBBqHBtsl74NCvC6cGmUQ/dr5SWEAB5Gb3q
sxlpfCg3HhPux5GbbQEqJdhagzRJQ/LQgA71X4zY7SqXHqTe5rLT9Of4XXnZb5OLgWksoOwd8L02
rPEbV8hAs9kiBHj1oJpD9ZIQJcYFnUN5WXUlGkk4G93XrEaM8u+aS6VuH7RdG9z4zuZQ7nvZ06l2
m8mwr8Rsp1zFU3LDQCRJBdQNgjutGLdx53lWanQJrHjxrEFa1rVR9CkO3c09wfCE8sVS0RIK7ns7
p+QPqGkbzci0omumepP+xQPn/mCXEsjFgtDPCFsggLPotjlEq2tKJzadGVDpunwpaK1LZWRJ1/UZ
NHKUxcCfW8lN3lYtCQ/SLqEczJPBEt3np2eB2W0XQqyt7HLFy1Er9T+Ue5lCUdULWKJwdwOcQTIL
HWKqtDsMQKVgUwl96fIMGutAbTTdPs12uqR/4uUUPjeZ1yPC9NXoLiOkwYbQzE2I40Zb6XrhPc50
kEuS2T7zBVzvpP97MTrW8DhxUTinXXx2YbqK/lpzPSBVanfPOemD6tDCXXif9K7FArw2f8BJppqR
FQJDGDDN4/JcqPcllFwf1TaYL2VTN675PLeBf+P9KQ3Dop6qdhsDrbTbCxNNEtu88TRPdLrg2UGF
IftEmzXSu1soQirtfXjOfPoV3m+gzNJQqcMK8Ppml4uWj/fKH777FnaaEG1OqMVW7V3a7y3Non1C
yJbbEdLYavWciccU/qCOl8KAAtbI7PdpkNbjqOSqMJ4oDB9Ko9cg3PKyN/OY0k3ZgzOykGeC/Iup
OlQS9IzquruFva3Ptc25fG2Iulg5wjBnQAqMfii7woEUg1wSWHJrtEne+oezPMPislM7BIY3w+eT
1+oPx3zRyHwuDw2scxDdQsgcy+o6fQnxX26vJkDzxFc3GMCNJmuf5PeI3TArADcw+XrLwE5mdMTP
oUk1EWX8mrIoEpQZ220m7saPE/CUTEbGmKeB1rcFNnMwUfmHzAr586OAB5Sxu0OKQ5p7RRGCBqoL
Tkw0cZAVJEf4MPBjYzhzd8SiKDSHSyIYBSgXC4NU6hwyw2+R/XLJSId/NSaFJnzQNyuWfLzHebAw
dSjn2seaOFDxuZNeCoCaT87KFWIwp76bfqXGchTTYvEPKglDFx4rO/0vxEg/1TUtWjKpCP3x3rGm
SMPbIKKvS2m25o99xSMShTqoxeBN9/hxKJx6uPNq/qQc3V+2WzuOwapYG2vbx2epJgOGjuArlNeT
lKM/iTyLYOqlRj7kKwCIdWel2PSwEspQmeQ+kU99TRpuYGy9ES6sTLi8yMCAbwyc6Lr+Qo0xTCX/
5SpAy14tzruZyss3ft9VLBWEtsiOh9oQQjp6T9NvY9MCXnUB607LILEWlwc30iubumTRMXjius3A
NycXCZAL7exKOCHblPqfdNZ6VUDlOMaJowD/h5GfFn0n4yy2fb1YOgcXNuVN5stk8lSEqlsIelf/
crPgN1uruT+N/tg8shieFFzthHC3x3/wHKS8/11ImVD77LuGkCAjywwoIvd5vF/1tn0S7kVsbF39
/TNmgcu1YSceRHfzOYH+/+8soZwhT6Wyz1HG9RF1648IuPXwEKji+V4/RyAmn/yPKY89OOS+MoJh
L4i5SlrqfTZ3z5d/J962U8mbz0TgKgvR9jUyLbATC8IC/gtM8t4lo2eHM6ri07q7fVoC4+dcxMNQ
GHrCu8STSLEOfmfqLTAbA9QnvaR4R1/xFYs+wR3D0MwIUua0W1yOxY5vGNIvUhRpIZq3dW0gh9tc
xGG8YfnYAhzEBLRN9W4NMEMj60cTGb5Dz8nXrJIjaLMSmsKIJYGLMQU82cnC+O3iA0mjtg6Wgs7c
5zAv7gg0soIjRNr2To9Q1Cqvcu8k/IBGwdPVdUpj/u14+pEl3s3WA335DvZ66NcXKRHITYoFb8LE
s5ilbCIyMHMJLTWRxKVP1jsjF8abPEBFhFwTuiLyC8fXo8aiy71cYLyl7/H7jpgZuI6hTG++0qj6
4jpAs6HaDsId1V7LN+c9F2vgfvlQ7kqTIFsHXHb7023OtzHUaWk+kbicqbztKQiG6QwvxVPfL7Ug
ev30Ri72T4BmxxUgeMiOf3H+OdqU1nVlRBGmGz3WfDw0whlnv0KEYEqjKAOhoMenMzBhACuKEJdf
w3PbIyomuOIdFaiNOR0qzZSIUwUT5PlAPcjfUduHTnaJComHFZO5VddOoymFVqe2Aa6PDz6ZeAWX
Bw9wDY0ktiMklbMBelGQWGCSer7pAaI1Sv9QJoLioTe0gCgGXeREinhWWp9SQ2QS6p0arVVC0VN7
U1FrtS0/Il5IrSyFOkFo+PyF4yxMD3EkRBzs13QbMo76f87rfrIt/8AiCqNShvve1kNYbzV45jFp
32pG/TMZqjL8H3lzB9wsMtT9uYTh56sntZ6zgMyFufnQkG4tT8vhXjZJimG0KgDMd/IijFoLbWPn
co4FMz0GK2mFeRELpGTTsXoQ5CU4VEY587+yoR0Jx4rBe4p7RAOMfC3wsTFWXaZFS8KsG+3P2oM7
Mo4ECXIXx/SIKJ33DKWQiheQ5ZAR7hhzLJDTX7ctsdxsCl4ziMVYDbwFcCOVioUh4n5J33HaWBXd
+Htm6O1OBLwtogopxXtpui68CedpLbAoezzHWeeFL3FGxIDrTIVmARpMP98QJ1YRaq6Qg05UXbef
qZeuq/SZDQgrR0YqVqXiF1s3aQ4Ale1bm/yWNh2yn6fBkeeynf/7skbOye0oZ4vQ16HzwZLMGioK
rgSwrU7h/Ctbo1WDyOy+Me0P5HzNea8v2IPR7MgbGw/mUDMRyHfqt2W9racLi0A1jn7EgM3H3udU
w1u+cUjKw05mQN+U91o81bwiVhnWKy+dUerVd1n8FaM32meMl4n0PcdW+cl/g1q/QJJQw475r6eu
ZK9MnoKNeU4fJdESqfCOkwlzii/6G3vpARX4L2M7CjzvzB61hBpgPGlDcYN1TPixjjHc4U3szk/g
1SygRCkPHhix3LjCwbndRdNHXI1KvdHNdwkFP6NYulTQ2OzNCUBxGFTvjDznAU8dDUXLjdM8gkKY
WoLkMIVVMizIdovLRmtS3aR0YlDSZFwAx+EL9DRt0gMWK0MbpL+JpVyT0EI3aIYTs1VzCwyCHpRl
Pz5LOszJIEm1aJhIRqe0R81lTsHc9Umdu8U2CwEMKNWntm3/qPZekaZvvxCtqYi8jV9IupFQJ0jb
YGSIXgbHEyG69bfxuZs79nGRQqWXs7zD2N39kbh35ZiZ9uQZIX+KcewRwY/jB5nJBOXJ/xnlk3j/
JQHZf65F4xiLhKyd2jpRQAMNNXJTkON5xSeOpCfHdiRksYrmIiunDwTye2euGuUt55eKoyDHU+Lz
dcgIr7PiPaCoUFCsKj/f/b5XVIGR5zVXG6KZDvPiW97W9Ld89E4MyuAmaGClaCzn97raddwtEbvm
0Enmb1NFnu4ssQ+ak30LHaVdSpPk5v2HEwVPMXtixJNyUABuM7/EGS3kp8kMFkPmWolcjJAP2dHx
h3TRfPi0MCVYxmFL04/3/jNiOUjj0esfF5EWewPcBlgiQPQSzMrjSWKfamLaB1GDdEleewkhch94
cbXn7kWCADkiuFW9O+l6OTE3ViRsR/glVbla0rbkUoAbGhDU34qn1WpOWUdrvsUcfYKV5XVm0SDu
lQzlEooa9hsTa/PDnd+1WouA8GPnl4rLwPivFatvP9y7K/EYqTm3y+2QsQK+HUF3DX5jd1oHmOWo
HPu+4vjvwsvlPC6iMcoi+mCpBcuRl1yh2aVMjZ8pYcxhyk+HdQIDNOaS4ikws/GfwbSGaT3YD+4P
LC/BjtsEKglTTDzpnUR1ul+H3tEbbbR2LPWVtj2P6Q8PvQcYw8M0qwFmqxUDPi8hnN5N9Srq7cxZ
LWy56Co4leNnLzyHs0so0KtACpuuNC0w/KQVOmq/l9Mz2j3IdJ0PkwITGJF+ygNO2DO7B1ODse3t
lslpMbZkKmy1DJcwmxY2nO1acateV6FThOkhEBajGMJeL4hdWOD0puW3HtEIcS97LzRPxnPYSD1p
lWwC6LVsOBz/dgEaBDfhF3y+lOnWofZqjwDDCBNIgACju5IjD0hHJeHOgc1PYSkd2Gij5HNgiC2c
+5wfbrE6cEZ+MN+FDD4/BLMpB471f7GvSGRlEL9+xD/DuWX+BwKl+5o7g45pFEOsC7e9UCRJx5Zx
Erbr8z0ToXkE/UlBDZ5I7blo3HqknQev13h5qVNgyW3eQ/chs7JizFZzwSoxaNaby/aZzLRMvC0s
5j/Gws9KYFd8TTksM80CMuv0gDbQSdC/JtgEs1qVGYxyJsCRBut5cLqK9DlqcaJfSVPIOCoD/Pic
kocNAzIj6IUrt1puh5ioZHZUr5f+j/wEnvuzW8ECpBiriVOBQrxU9lKxPpRhvuRivoyyDulRMajr
1H+TuRoQk1xccR/y3qJ/vfCEQCZ0znVsfC4lfIxB9OzmFT52/KmMenCcuYpSMqdLZTZVbH+OypDI
AASAvmkxM2OXPS+XLmZ6kze+CJ05TgO73uJi1kQojMkDtpTLRycITWSUmstWymkfRdlHpiXMqK6h
6AnI4jgmp7fJQn0hkWHY4kqsCPq/Ej/hDDyQ3W9p7We8ydbBmmweWHaLtbAIgnFcS/ZMhGt5fjlZ
N9aDfG6j8EA8qy4nEXotCVKZLdr120lAiy82nfyqX9pTfREMdtWU5vDXxOk6qwQuyPuvmmSn3JIq
F45EMDc6rC5oUwlG1w+nCp+gS/1mxqC4n9K1VVRua94v7zhIN/Rif7ix0zqD519QAtTiEAjr5tTl
s2lNXWWr4uDxNE5zbU/mB24gtUTCI/q7FiYQ7VCDoIHg3xaNU0FRQzrzc8PVzcRECZWLPM0uv1nu
m4Y9hPdKHzJV5HcYKK9jhHJx2ADd9Gy3YJM827OTRAu1sqKV06fpv6lJboDqvdLYOL3AVa2dNNhQ
AsucYP+hzzQ17JwM2SVJe61K/I6l/u2I/JouL27ChERXwHo0osZ3oRtmSLa3wsXKgrshF27nhKb7
yUHTkRMU5G5Fn5/chtG54ZmfET9bJz3i60z4H1WokIYRbCIYQzi6l/yUpemlCjn6iNgGGseRwc8R
P7scfXIkR0dOLubLDxz0L1wiUZOEa4RWHki0JvxN5/Is6UlMysL1tMvAg4yRaHubTUsT36Ka9kiC
+FUZ5xEFgb7edrtiod2vyau9PQbwg3SqMSFfEH0eM806WfpX9yEQ5St24Wh5KebgImXgmdZd301T
hYOsvs95CvsZhGkOJgmwgy/yg72iyk1rnrVF2+3Ih3rvhi085dOKrpsJLYmRVaEQGE8JKcc4ME99
1ByAHZzahkZ3tsk29IHTwh6Ku/gt11bktGasMhbc27qoD7qMQX9oBKDUMYzuPQNz61KNW0+toly4
MWWSq8rPR04ATeR6KadTRtjezA9PcRExeK3HCDVvhRjvwzG1injzHXZwJbF8Z7lAeXqhh/IIv2DY
9UJIgLX5L9DTKPEkI9ck4VtOjZaEO/ZaRKXn65altH17NrkP/bZXF5NPy6vjon6qKnP3IkhDEUtf
hF4/gq4jWHrq809jIcbaib60EOqU4XmEXbVBYe1C1TxsfpYgPWnLdFodrb0wTlPB5NPM5pj+XFEX
pB35Q/pspZd6DcS71kWXjEGIDnmkqjLjuC9U494rL7vy9bOstRiGOvkCowdAXWU2ZD8sro2H/r3y
6iMlvbYNSwKLa7eaEqXBy0H0Ju4gMB+ftO2vp9yFCVx7KitbS9NOyFBKzvf/vorvvN03kZPL55Yw
LFOtI6TWua4ArqSKLYWWZgahyz19mXfI1OcD4I6vwrKxfqIsSC2V4XzcUfW7ijZpLgiwGU2WoceP
qUMOOzb+c1sl8B1hzX9fVLXK/IGAOAd/gubPfQKoCXoz+icp4FnhRO2xkcE4XC5sE3WtA6lJvu5C
50ZiII8GcB44OIcy0TQTT5Rvja1YQNY4sXtdIgGSEr+nIB03JGl47JsaGHP5zRvDORO36G9q+FSw
JBCQ0V5SOED+O7NwdmW4+NW6GSck0zZi76ALW+LT+fuLUjdf5HS7SnH199zutLq5KsVSM+vzLPFS
qwjHrbuKmSm2Y2vxCxBLohlS07ZMHbpw9zfl0jnx+ZhNluFc2tYlbN2pSqg/KaFG+L70AVU5GfYb
YI4xPfdxBNqY/YpKqMEQ5VWJKTmDH6w8hP0EgJia1tN6z80quLsUFgCN/SlbxOySl40KCQtVbbS9
6re+o14nGR/K731i5T8Qli014jnJ0BmeIIZ+USFaeCXn7LeHiBxJ22Z1RWMl/nR5AeoGXJsh5hA2
FEkAOc29MmKxYTmbBuIyRsYmMaGXlVBNI6L5FLnFQaTOqfL3qOk2GWYn7obs7atZQnzqbCe5CEXZ
QHmFog8vgpj8OqusWd52IyA9F1gIzIcaESCFVH5TvLk9aWIII0GekWGRNwlgXOMvyBb6oOLYCFcs
iAOmUJ7f9wx++DtpNALDQ6wKCe/etqklmdNGfzhDhVDLY2LYbJ47CRaY3lEEi9yyBtXoG8d4QBuj
jHfjkKm09PmbIQj/hmLe1G2G/s6vDEhy97IzGB9myOxK2rC5GOWNPXq78JEltYc0ggiVKEPOTGmk
Fn0WU+8FHLCj8ibGxkVOqYwII4Zfru7ITtdPnlVjbLOal752TMSY6WPlNg7mMxauLJuC0pU2F3C2
q2S1tctyTFOZtSGONdcghAr6iPMS68+W1VX+rALhmJ1iOTCWbAiDxG5P41r9DasHSbuqoSnlcqhy
KFSAClzh0m69lZPYl8dZMAuZHNNYFV5+JaEU1qGEXXU1Rj5A8++xZ/MGNcgBz7VRJBZ85p8Umkjf
SchhCsv3/J3CbtJD8KoEPq/A4kI61CX7WmLYODQmBFgqMTZow+oaNLGBmItgVbP+Lo+1/76ZL573
lNBKZFzS4gKU4oCqUQa+0NDt03KI780PvcKirjKmaKd8xU1VVKFQ1O+2btw2DDPsKRtPNL3RsvTp
jja+ZkKrQ9pw/MQs/lmXfhBHRIUJf4g2AJMaYhO21hGouUvlXRJrrjFQdTrlO9fcI1GljlZSTb8p
jwqQQXpJ2+L7tqCtRP1Rytcdz01sdhFoPkoAAdKVI04jxnDVXaShztxIq+sn0upY9G7NhUtSP92D
yASxkYeCeq+ue9dpuBZtasAjl455dQPNzbxuUzyXxwTDZztZmxcCvTtAoWJ1thYez3qQrkI2ECoF
FbtEq1PWmBiVkC8OkJZdC5rnoPi5g4HUvxGapt6aHrlHEG8Q7jr8ezahuovDcrjAXPNw8ztaUc3n
AibsN97SmoTyjNGy4GJXQyNLh8c/7aU9MPmH5PLVKMp11ylbJSxo5AW/Pn7yAPCWOE/a/CbiBfsO
yNE8h90l5qyQoGBMu64r9TpdXi5tjXxDm6mDbnzTa5EtkYGIEPFZtXj+WPLIqv5Fpchkfeu9yAZE
HoXMgaBYCAHvyYixkWssMYV7n+WKR5GkN3wouBMIT5Xmq1ZZuoOxi6FZVxab14z36PhyfH8yF9l6
wJcDZpdQcM6IhCASifqOjAfb3digCBEDiqs3UajujyvG1LiaSPgY94a2FjkvG1qnTE6w+K/i08LH
WsXd37hnTmwTSJ+CJ44jHjYyGYSA4CORAzYEpzbGE4SsLY49UKq5m7dXu1tIXifd67YH9cMVjAWZ
9u8aMAhEoTF4qP+osX1g/xqIz22x6bsJbB7EHrBaGd/cms/N+qqy3O7aNy3ZlzlCLm8mIdS+YfW2
Sw2K+gFd8fwTuur4xVsDi9z/klzD5e6inpEnIJMZ3ApKlx/I5EHccP6Yj6MmBKxfp8ptDghwizzb
7Zj6o/T9WTCCdpacHr+4hCXLZWjTfs1auW+y4rjnwAFgq2dtEknCeN3BmTO2/e2Hseg/6J4AGcpX
Oy3RKAZVKFEKAenOgoux7JsXz7I6zSq+ncHQ3kLPjuCdsl9x/o7bwkNv4L3OGoOehlVtuSEnDp0A
Uf98oW8HrrzSz8PPq7xrxpeIb+8v3S1UxDsR8skwTzu4Lfequ19R0HrMlpMNYVPG9gsKe5t3kXHp
+S68T0P9PLlSzVo4Y7ANkbX/C1T1Rl7gUpVz0gu6xvcdxHowt+g9E5I1wMPY9VMqblU1neEMNC7o
TLnR0fnr9AO1+6Myy9s7gNnFo6zPIrctZCFF7R6rarcrwP2CVh6O+xvflPi7JZWWmlwb95890xYo
+f90mnZxIEBMSQSAglIWVB8Df9+ktRG8rHqkUtdFrZmHOsO8eWPNn6WAPmyr1eEzy2em
`protect end_protected
