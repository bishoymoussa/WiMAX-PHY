-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
VxLEyIiF4D/PJWZu+BKffOdRDmumgEWO8QFQZYSsBAfWfTyBX0JpM2vXrHpowB3JReG/6pLWPLiW
Z/uYVOdbAZRfiikDwQsgP7CEwJEYLELBqHWD2NZ+QwTmBbI7Wb90ngyN7q/vBrDsyhZfGIpPuccP
Yxn4MUNLT4W67FOHWFHuNEgmfoGT+mqyT/wcLLriRt0PPUhLKm1ZYHWNqzajOy/MA0N49EbJ5+PR
jhKKuSnpA2xDbIBm7DBnUhRDle9jbadtoi8DlQxsP0Jkzvis5bPOFxJzlfhEYJ1COuuaeOmq1X8O
aoDVK+GDXW4dPX8c4qOreB5PGtAu8JEDoWrHVg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 25136)
`protect data_block
xEAfsSJRSYiwUbxI420bHyx1urTr4LxsuPMuYBxX3ae7uUB6B15nAAfEkj9V8HEFZ13uMY0yPwne
YZvsSOsUg4tekvUGl4/tCCGh7z7daIBLaVZpDDCxzcW5aB8u18PQMDPw2PQiI9gWtYcp1AoZAPt0
W/BUR1e+psHrh1hfGj582GwBJBa6PgmAmxxHj+Pe+90eDsaM+oRzWXzQunjMRXNU7AnMbhhDNOuw
poQrwFsBqYxiqGEhPpSvfP2AoIMjpaIsB2yuwptN6zT0xe/fb/+IXGv4CeXDOu72nrR0W3vOVk1X
3sKCGtkKfPMnu4yhFkM+Sv7BxnDTPYmt8rRSJSFgmRlCYdLtGhwyjyc6pEu7WYpQ7/39w2mdlj00
OhvIlB2wq9ipgPhy6TMBXum2Wjg5/D498C3CcxPWKZNzGd0KgikKQUnlOAkT46Vo7qe2mkLUegF8
AoUzBpnKCRUqa91s61MpQysE770ut7izI7CG1rE7n4tF7jOb8e64hqHoqDpOwlmS388e7BUhrVdb
0CX0CscLba3objHUIo36rF3sj0RLNV0xeH1jvAjTVoW+MXcAQpDQHnFjkI11MBb8n7a2Oswx61qw
mSTJCitIHbdqrdElrz6NONOdYSPIVDQkUIhENjzdd9aCv8EAMchkBFFo8KbfAf6OoaiJtGAwpZi5
u2VUVqO2mHeCFmVlI7tpQv2duZZOnRyQ+3pXBPsyH2P30DMFBqDpvxIH8vLjiAYs5c5dyzADjmZH
IE/b+wwDDKAX7HBUXkMwu7Brb7crY8GCAA2mNY2um34Pd+rXQ365gW+X7jedODpAGRMit/iBXY8D
7EN4Ce5mW+N6pBZbI62E25lrbLpSqO5BYkdLFruCktX+fgtRf3Kn3TF4+/9Gw32xl/n27tSZxwIH
iNNDM1+uob+IxijEPWLYX/Wenl4D2MLY3seHUm409z128Q35ta6+5z3e8/F4qjU0OpuR+lK7zZjv
WIwJxaRB6ch5DQ5cS8FCJltsp62CMS3p2qQoxOW7Jxnf+auiYrQIrtV/1anP2iLUbWUwwShnD802
dr1OCZk/BkASUeSzpBo8B/i3kSc3cwcWGOhtY1cMFsdGM9T77ZE9BXIvIgHA0opPl/LwjXVeVSyK
RQpiewYzG5GnszZVoyQsSCidMWrE4B4Nuc+BN3/mt+etVcnBh6qGtYL1GBlDvGEOrVZbete76LHb
Tjygq36UrFWB43AlpBqj6wzHzg6UUEI2DIi2WrrDenEH85AQWvGCcvXlJteUcIlVsIBakhw1/JH4
zc9ydt+fGw6GcFrqb8NNyn7S+BkVuD4XfAyD1pdE5jdkg644om4Mqnr8X+T3egBbNOWp46nHXmsv
xi9acgxJK533CnfCzWFCm4D58qHMYSfVKGEx2kfVq1L5cQqnMTI6TvkKPayQ4JcfQaBNE5710JV4
SAA3DmR5IjhXTkQziFFZNPiBtc5DKQO02VsGlqI+h18DElMcWbARfjkN+gjvzZj7C8W2yxeYmzte
ywpf0XOpyEsAQPL6Vbn7Bez0SHAnipLdJHp2cFObpS+BIHDHyWzSF3tL5BWyuX8IE3+C4jWsiWb+
DICf+pKalKBMQ7nrVicHYAscO2uAYK1V5iH/hfsyPA2nHPOmrmUXT70+JF36bKsSF5VVXr4+EoIS
ObS4wv4167Kpf0okgHV6fkMIfXzX0QhJ+n6x3DMPiSelXCx5ODOWALaRr+/ptr21aPS4njY1cSwm
CAK4A+fxTIsvwlflybTaY6AS4TDMhgfMJa4IeQLEOyqOVMVvSTVsC84xD1mnhljpGEOr6D8VJ+5V
aZvTz9gmLF7JO07M2Bm2ybOoDH/hFVczu6omGM//wb7gAzmLs5xgGwRvUqelyiuV/nnNuzxAiCdo
Kc6s9yln6CGEQqufyPlGdCacYS7Za516TvQ8vyLJIsMmMei48zSlzpJd9OU8OSTcquTPAFKI4S2J
ol2CA4I1oty8Qazsf6qCC730GwbSKYCHxCNyzK3DDtpRNNjgGDT77YvQYQmjcTwv7CRe4/pJ6z/4
DbQ6aDF6ROS5KLkjN/36a8w7ERSx9QCsHMML7t19RjsZFyY/eNHwk5Y3x+PoNBGiU3ItsBHua/2a
w5GvlLIG5Tn6uCypfeIqu1ufRt+g8zratRQhng1fY2ewYfhoU4ygNza+S1EvfDfXnfiSxCVzeDjm
qKdi+xTDRVJSLMpUmTy4eHocV6IkaOzSNqtu1sHAVUwK5e5g/ccgvE+0Fo/21f1AvkKdWUzk6nDY
TGBxryO+IrKIynyOWjdkUrsIe7ZdF+JD00VKwNR2JVj4I0KQJC5jLUiOnk7k5Uv5Ln7+rpvFnyjm
pTqckei3WPzl5/Iv21JX9YnSNSjn0RTYMFU/ZUQ92A4CoDHnBrPvPAbUOjDC2trtxyE+7IFqc1VL
avJZfn+9VzvHDa0BPh+cfEOxKUBht7HtZyd4tBfpzayVF7M9BUfeNgoyMtXiUuIU4/CHN8CLcEcV
eHerd2fDEpBAgmVoBtQ91kJ3UUtyCKZEQGgZYyfFKkbv6xsEMdEnuLOzyvXTY3GjNzfHq+JbDmp3
X2u/PDI+pEv8n1OxxlTapK6ioLienixHSuoylWWDQHBs7cxbksn84K+lbyJLc3pb9pGwmxwuRy3a
UxWqZ/fu/K8vF4o6OgP6oRSPJhxmL/r/eNmYh9eCuy58+dTc/15NtvvZ79e4mK14rxQdIXU6i7Y+
p1mDRlc9/5AEx/6PR22PQchhatZkn8y6Wxj8VX9bjGPY5K9Mo0JaRasCvoWv5Kiglpx8eJYWrufz
BFYi2wNWz1disdkdsGI/0vS/9MqUq1BL/OFI/Ya8LJ4N8BnscDSXNqyRASLMGwooJ7PiKgxhKBIn
ZAjp/+hwJhIcSo+M2+KJirQVgo0aFhz6oHjaiNnxRYyGbdrVM/o5nrmoe5wejj5yWdMxFlXzcoNo
jDk3Thuhwp3dTKlIO/WHNIJ4AY6XmWUlyzhuv00h774i8imv0D060UZ7weVYnzdHXgSooz0Z44kX
4dCpvTtI+vSKAL8YRZ4cwqmemBs1tEgkqqRt3amoDfcAZ8sJPHL+hfaDLyeXpXJ3sjwWBfbSVrFq
kkdEt+WCjkf3flPiyRf50mP1cUMA+5ncUIVCq+iLJDg5FE9C9Wd3sC29bxX51yTrNRthgC6SdzZW
wNaeaKVzVQTMRHj0IcX+kEJ460+Mo7g2yc8c5uLbRNHSMFV3gZ9TANix3zmWc5cZj35+++1ZGqiU
YQ0+c2ktqzI3nKjsMZD3cLt9nx1OIOogmUKhnejbO0RBBNiu8rFU3GMQ/eVxr7jeVDRJWVadx8p3
oH+gVytUCGDzvrlAhfDkQbt9Xoqq+7jHYf7S2CeSIhbnaNeIK7K9yGc5MmPtzUw8knfwHqwIDID3
vm0/ZoeFl9SlNtBynpFO3Ki6xyaDEDG59YGHPXChDK/5/1lkTP6mQYlVVnakYp9lkuYXmx/9+Z3w
n005AM04avsw6YyeGMWlzkB24hUCNKv8dodnb56hy5VPdTyZFeqo9ubOojkbbyisMxpzdoFMm8Fu
HMgXuKp83O6B4KN7ugnnZegn/Zrkq87O6u5wtLBhKcA6PX86TSErSxi6PyFJZc2L5aYKRtZbvbLd
P6uTtJjI89k56S6MCyG2DtsnGSNcr5Wgh94o/pG2/Nb/P7HhpTDsaC6VGsu5EvX9TsRfIRwZzBTH
DBQWvfqSRRgG/JIL7vISpGzECHMhak5rcNN+6/sQ1fMWY/F4r2YeoxILE7XfE7mQ47fBBmtw1Jnn
SFaZQkSaRotFXKE3AHiNn59ZFWt6vI15XwW2T+ynAvyU1cvBb17xvw3Af1N/P2/idNK0JfwtmtMF
UcPiVtw7vY2ajowENhb/WBsGT80uFEawoGsEcUcI86xT7TnMBYQ2sraqzWObf+q+f8B8yWNWbrr5
JBbfHl1cC+21jc6JB3Il2pdKc5z7k7I2eb6+9tCbR5+C1emLXm2HCO5EgjSPxtHTtHULf0KJH7QB
ck12sRFJH6EZIkWc4T9pFcIg5yy02Ph6iFX7AfoQKL+ge7QbKBOPjUmFUo2aQs7Qph+GRQcPRoGy
HZgYCYprqGZsvo7TLVMEtQ3+Sb8S8ukK70xMs/M6kVszoIfroYwmCAMDIZJ/zEsXea61Ww/7Dihc
99TItezOD2yivtzQLgFCMyv7tUAp+VBgIkWV+VPYB210+xRuzOF122TWPplrtVwOiiQ+6oX2rOzv
dwiyh4BAOsQNE4WnQ8Yzbr5BSM+Z1SYx40/KYIP3JgwQYLGxgpZK6sB3GQMc+oNFNr23hZZPGT4x
+TzT4iXbxjtBkkwxAPWMNEc0EyKTHW8HBjI2sOmIUzyvWK1I9cE9kQ/+BTOw2oKhBFXEu/sOecA2
7JzeSWKvb2uxqY2NEHHXTQ1WCLPI7mVD0Ad2HwkVCzO22JwyYNUec4cE8I0efeJU6NSSGTjWY7Ob
fru62DvQgXbxn6HOEEKOpkVpj1Izp8tUFgNoaKDhDpcbjXInHiC7NbYScn26D2i2CU7VPxFbof0T
O2Hfl+4KTsrSpvkF9qYSatvNezFwIjY3XGV6E2ixnVJuzXhOZbI6VrMjU2cCzJeS19HOnbif2y9/
9SF6RRNDEHYXtZfBhCVF6KmgTsPfOh4rJcQkXUwoBIjNvvKV1p1PCZ2U1KiLebwBRKu98L9M/uG/
ae8nId8+XmfgBU5dMbxUGVUjV4ja9MlA/whgHFsN7N3ugBr/yH08QMt3+aO2am0tSDNL8u3KFIwx
/SMFearO961fL7xSYkAL/4VE/+50GVUX9O6UIdendGGNaJl4G72XltRREqkyQEZ8HYLsKhtvV8Mz
IiXfl7yZPMdP/v0JpBiY2SiSFVGbh1OIEIKFrk/zdaUyn87q32BGtMCMGuGerZl0p6JYjXBA0Y26
ozNj1C0qPFX4XGS8vJoPBUJ7aej+XJhObdMeJECG3wN76vr1rAQaYmACLYcLZBG5e4ygQJd4x7dB
d0hra+9xx+9YANNOr7O6wrTqqWLHuEc/zfHDyn36NCXMHouiK6POaqtWMNXL6cdM4tayM5ZNzu2n
TXueInOwu1rddwrhlKSTymsEwITJHE+zNKC7vxUIkE+SCgNZfKHGF/jfbTWK1IpdWHmYKNu6O7hL
cN/ULToIA03ZXPC5TGshSSUfv9yG4w5C3y5EzBpZ92DfRnfPWdP7LZfgYZCRMdmTm/kHshXOaOx4
M9wmDJSStt+8FnMJdPPWCNPNYDDkUr3tAlixECekhhNCW3vlL9wAnD6rizI8pDxZuk/Hk4iFwbwZ
yxquw+/4VrbV4mgSRnLfqeZXYGv+AyI9fiLhlgxoQ28pNqo1KKaPrearbojbh5cZCLf/arKcVVuu
FstRKnz3+pfA4Pk+Rh1ZPh/8p8NbYUxFnMvJZbuEry3rntTkMzgcRmhLxc70eQLracMguR+SO0pf
tondhcPar1G1V+aqXoVH4LBtNIK/+Y1mYaYudhIsDFXS0EApKs+9bBL8mrnf9sPo0vOv1L2v0M3u
9CM/jd/Nc4ywIr1Rb55j1eHRALIYxK0VoiwcpuHdIcaX8EZmDzGdYyVFyNZxG1anu7WC5ptmTQRR
db9EqxT4AaGw9eOQBU5j1ws19wbRNYWXd+yq6RAAQtmwD4fk7e/dv5XjlHVlRkrkyuygf9ZUKoOy
lveQqP/6VzFgI0feRoV9D+q9XZGlBRtKEUSbKrsXK3Oz/yf4bzlQp4ji6BZSQXNWIA0D1nkDe1oL
idglmHZSFgO9npyrcsDSeXEmTwIx7QY9/O/HOJUNRgW/fozeSFa8hKjkiceJpm8AC0NK8dTEt1H1
4fqjjsF1IllYrNMSk5jQXJYXAxI1F8F1GhSYA6MCiYc0Y9Qw6mRyJ+jkTBLS6+A+dteM6M6UaY1b
4CZqaLrNAasUzwI9wH2fg9YjL7GazpsIhhOpIQDQGNQpQSjafPXXpDhcuNgff9yuZ3fUsZpwAnb2
YARCsiHEaDkpt0cXbD/Ct3twRPHd5b6YuVYKUFJ19xLghr1NshHQX5lpBSiGJdNX7Ecs/N2ZrESo
VR9awirB8syI09BjVMYbX0NOI80VL7Mw+zxfsCT3Zf/N94o1cN8unGgYLResO+Hs+iAIEdL9nmp+
xXvLV91C06xa36sWl0S4EGSamPIncVeX6OsATaH/32DX+GRE0U/mNV4BE+MqUc+x7jGYIejDiMHJ
SPhe5j4WCiYFSrRPuMlvEFHQqyqnj/iBIRDcD+BQfadBKu3zYxYkDqmrU7jZN+Pzo8PhJLmyLvls
XsBMp6VVh+bvMFZefMuCTkfTJ4JQ3KU3as5LaiVags/EkIy6ke99um1oUc+4GkGiBfa7Id+FzY+h
MCwWAD/VYrz4MsGNNFrXdHlEjwgSxkDAvASToG7jx+jrrxAGW5I67D8Q26eYOeRx1PeyyZFXxcNE
Gl45LE4IKDfZD2VYi7K1hJlxbtVTa2hyHX8Ksi23G8sp/+wPAXiKtBgufz25E+l1Zkxr0MaHe4c5
Bpe9SE3gI4M+aPAj1ePvXD65jfTtVd0X0wEH8bfElATDzXTkyxoCu2pIskdS1uKY33Of8qUF0RYb
c7vaZL8tGP/EMcQ+XB+H4jMgCIzSHGhiMHTBy4nwr8qLKeyP8mJN3W/u4bZjBBL0ndZcvGxdk7Hg
R34RZ2GQldK6D8z0VKSEP3Iu6Jg2p1ANLPkYwD6BC116BLqDuqoklRBuBW0LvFOJlR+uyZySwwSD
nCbhAPGcn9OlMSarLTGHJ+DoS+U/AOl6AtNNH0Dc7PFjgkYogG1WKpvYHtQbxqeEHl5IZj31ORfI
Q/X9wDUOMYcUczjwCLKQLNbV4sRO6Nk1KRbPAJR3/+NljWed4Qo8pME6S3a9OW/iBxD3dhVWdg0v
FZhh0UAk6356Ol+RlsvH3oULCes3IUTWYpJajllT6FF5yq0jJit9fe2tu2bZnvKb+dRQr2NANN7r
4xkXCn6ckxBMmkkNeF38+SRd8oB3rmlVz+1ln6d3WP1+9UEb+QjhPH4MU6gj9jS49erWlj9c/7fn
6HM+0V2xo9kEea3k7fkewHRh5tAOZsUT7zap7rK0L/zI6ynsmlh30CWtuGaAddFzz+2NF9uwIud7
T+vfeuRcXD2C+lIlsm+8yDpG02j1e0UYH5VN65O76vqfnFUoZhHgeNX4jL2p1FrlaGiUCUKr2OXC
Pa8vsUtY+AViRDDQ+WRyjNGRIR1DWg0zGEwnz2/j7WRUO7bpqAcOPyq+8o0mQcckfaFEca8iWKzo
1gD1JAqYwU5BSS+1vEpqRsflsijFCoCw3VU90tFnKOvxDOOFxYKoTWqeJRgYkb6SyTgfYc1sV3Kz
4gUqhy3f4q5/l8P4W0odYuZ5+Uq7AQfpe3sU9Ebgkmyhp7b+zB8Etld3GKTd9wurnthNkR40V9X2
40BQ05S18S2zvp9045LXTXwuYvlg6ckztL6ChEJMXCx1gS9wdr4LVs7vixBNyeojsIiVl8pl49KY
G/lc2JJzS1JyLCaVIZljWq3ntxLhaJYPn6D4ceil00ZQEensTpSuQE2O/Vv0o3NYckJLB0dKplzG
0t4iMYz+QZow4DUkcop+95B9ZY6iKKYq2XVfbn5KuVRSvljeRZhr1zB5w9FlN7F3o9GtPjzz0V8A
uBqp5X14JoX1VFk/cW34Ws1/D3qZjh3ixfnqcwWvk0RF3GA1wqunpuU7psvUHjmKNjJI++RXIxzb
RYX+DVGTcjMQ+VPWJOEHlclKTxw/eY1hLhpfddTDf1kLw+/WgTAjQZ5pn6ZAQgTJwosbwrkJkohI
2WdrdWn5+yoqKw8TctEf9kXTdKyBar7S06VMb0Yfof8mV4L8LRsWkHNlQW2Vgo1ScfyHEN2+35m+
drumk//F40yym3mqZXKNzGxDdhkEZECMMo0MFtVbWReVsAFRbAb493PSYlnRMlJXiL5mawj/67Pf
MUT1lAnj2x8sowRNzTiOYtE9pT/R5Fj6YyUCR9cAeF2URIzEKrBNGfTR8adoI/Ch3ArRv0+ksDnh
KoCiD7ivAqM9TKLpXV8bQvnlBokZzXLQYmzwtZvKREcwdxUC5xgt/Ikfo6rX4Pw7AGkFMif1g4jC
g/nNIWjlmqsfC9fv4SW991xPRSd84AVUfNsfupBSn9pWh/8UjTAak+CwJ4L5PRCPsKwGzelHj3kz
Uy4uqmSmj2rp63DGOzHrt2BX0TTV9SwXfznl7AmyJ2BrUv6HHScxWVtZIMCw6gXju3N2OUs24Dn2
OtfIg2LS0gYCyPAMRBO/xgJWx+PW008T+1ZsA/BX6YtiuHjI2l25zapcuYScOn5N5E0GdRFN50Ru
DRTVSxADrSyo6+s9gnADqM561KJmvdBMIsUIWsmgaqccLf5xARqeLkd9cLhp2m7sdsZP+mfTgaNP
R8azQ9WHwRKi1nzOshSrFYPLn/H3srRrrAlu7XfRRfnLlz+Qh1tR4J4g1EsMwInuwVo7Mq2xt2Xk
CKdiF25OqyMwfF6kCZ7VyjjSJdforwDHp/iAItBspC/zeQlZI2YwyeTsBafVxXw12/tzP1H3ZziC
i2/U5Zv7hPIi4NaPuOiXvvBiI67vjpOE9vBiN+RTf45zA2bY+YzyuafGcGeq8LFUYTKlSN7hM7Eg
IMOcacT83IN/lXe+Z+qqLhI+vDLzRAO3jUgPf3Wbqk0bszw6X345dqIhzmgzUZlc+dlMm4INfJLu
+owgAFj2uBuQd37vmSkGT25k5kxrAbVG+GvUA24AVGcKue97ehW+O3tv8vUVyQ624g14LOyj/A5x
csPhDFupqZqBS4/8k29swHjKSoMuyQ6g2ng0NVgNXE+7jtThjeTGwem8T21wyGuGAzkb47OozwVE
BEzeEl5hBmsXoAZ20yYWaSrj5J9LetRMD/N5VAigrgjMK4Iyy5rqu5dVfgZGvQtaz0xq5gCC43tE
PPwTwQ8km60Yxz99mVv03xuySpEWWR2fg89gH6Q2RaNZlBgZnXc2QExwizWn7Hn70GtLJrLrbMfD
vW90kM6Y8eTyTP4TLd2mOXC0V1zysjmaaKJxR0/yMEm9jMHClo6+ZQmmeGywQWhn5YvsMDnFDfA0
f0aWR7tLZAEej/GLAtudHXHl0KtpJwmgmufmEUay6tSZ5MR1JDesYTeXWxJy7lpwReICZj2987M7
rM1ZWOqO8zhXOhv6M/kHBWcGmJ5ycWxRS0jJiSi9HYYhrHEPNAN9BBpOS4S3HP0fPnE0WsJklvN+
6+KBi07F7JP9HPMkAJO5jB8ZXPD2U6LC4PA03cZr7UhWQ1PRIMBPo6VuuSMDsWr8BReCv5c+o0OU
/gobtfqUlYzpqLLu79MGr3k0d4hReTfgoap3+vkvz5N+OZfz57yeTbLqf6GzKuS2umLbJJkWsxD4
aDlvGm8otDWG2BJ1gLz7AbCxmY/LNjqZlD6ycQYcUNfF03CCOB2BZHMtrIFnpHvxN4gsM+fkmHW+
1If6XpSN3R5D0HhP4Ovys0BwJ2/8Q55lJ5oMlG/ey9N8EJl6BGlzwGzkhSA82+fVK9afOEmrEuJL
XVK58dOvmc/AO5Kc9oejGH4LvwiamZyJIdEghl35RYdI9D/UqlKFonbf9zGm0hlGjDh/TZ3ZQdPO
U/3Go5pD0vCikLGwtznXMEwwznyeQGm+HdXxiqSeInZAy1JmBecCQK1sOKsPNBmFqcxl8VAcJdZu
lZnUgfhd/49vK5iWQ64ZgzGGqnogufFLgOzZhV0ya+DiubAwRDCDHkaPzrdLIXO7G3I6fSyeZ+mv
dl+Is8GwPvaXbY4yGFmB6p/Qll8T/nD3SrP8rJSzNGRpWE9cww8b1fGUnX1ZDZSV04qoRLXMt8Tp
mU1DoR8xhS/Q0mEyTycGYhejnJmTbAEhTHYOBdsuPdBjsoGm+8NRX9nLrUUozD4D9u7El8GqMroK
rhw9KFlhCquUbHXVsansNo09DgIzSzp95mrJ27KG434s8tuSwZFHRKYKrwsCa7/BfzIot62eyFEb
FvR730Fpp0a+0YAVBCCwq/a+cNCyvHdHIl98rVMAGmkeNpw9lgIJMsjlTVGqvyyMP5xo2u0FnSQP
GZPVubmztzFSQqeB8yW0fAuNjkeb13qBkVmBweYn+J9j9MX2iwk+qdUGnK9itt84kPrGrICtzlWE
aFa9R/Hq/9qBMKh8sHVsC/4nBRsqQoZBvjKgkmiLihVWcR7ZZ7YOuzUFls0VgwedIndIv3+IGNbS
4VU9Lyeu0KFLeSSXq7jIpAyFOcsOUWK4pHyapftXWkfCtQ2IO212iBOuvUPD+DpHWhSBmH1r1frN
PafAxh1sRCGbCTLy/RFnh1TQstVlayGKvtHUHDbL+ffrYgx7LXocO4yYhCUpQSByxcc6HQxDQ+cA
EMlNk8E84JIUmWxTKCd01ZFJrZFW/rWxMaPVXMpvHzyOZdsLVu19/isYi8TYtHdg5EFdEuTvy82F
fMj6RQy64Qu5smrYIeVAjCLaPvIO4d4tGibRM/0hJa810300AilM2pw6dnoIPM6Yxj22SxAWhe1r
IeiEbCJZdwR8zEZmhBQOs7J7aVZbxHgHn2FxgdPSRaAxwwgYALNkzjRGhHeyNUHhiigQD2bPvJ77
+4DrXwLEk1XK8RWMjFR9QS1oQrVqW2Co6L3jH/X3zJiVavbWSRbR4aFavmzcdNSAgVBztz59p1Sp
kwAWNmRg5IBvskQcAJs9kxOIJk/cyI+Tx9x/ghdaxRx0SBGz5nsMC0cV2xGcMoML5HLoMS5pbB+3
0/Yy/1ud/QQgLI7rGVPghMRVcwi3CJODyrpIJSHPPAvc3QQ0YaA7B+uAQMWEPY9c38yaA3lC71Gy
BvLoqtnUlXGtTTy2Ep93JR7d1cnhuu+vTSCnCNVR56maI2hhTI5xD/NUIt/7JV6kneHytqbXy84w
/E9BT1afskdGMSqo+e/ipHLOufCzuiAJbBTKmXfcdrIhn6ZHpdVhJWsrNg0f4dHdmExS0y3kRLtf
rbFYgu+fSBLBMBfxEX1T+bFwvg0VTZeXNjuUX794ITB8DSCAE0+rkitFcvmbsfafkzdsyUcGgHLG
v8JCV9ZF6N5FVM0u4CWano14k7+GoIlaRB72lFLvNquUU/xOvOVEeXxCxCxOdtO3RorPakMHl416
OU1VDrAVGw68oRRWtfedu9GRnL9pq8UlmFxeCqp0ujTt7Ch33HNlt2AY59vshFYvs+UjyL0nGa+B
J/4xpJhb6W4BY5f+qL9tlAHv6l6i+2f0OqS/7DbxOxsAJfQlX+kRUPtcfCMhVT91WqXdi70tGmkN
kN+Z8qHVEsUNcZpkC8W7SKIjwS/2HKoaa5ObielkKAYCASjwmFJqhe9hfgHBELIeFfgcyGRj4Mx1
JZIzruymt6G62EtZfwGFtEfGVmVtGwOd2fhXXiFyNTJxO2C5zJUi2x+70dRXozPD+M8G6/SpuwPz
N7lUJinWPCkCGkeB+4g/BrXFb1TzD1hyhIkwiyY3drfWDJtx/zZB5jjRFHhIRFGp49dE4k/iUEnp
rAOZt4/7BnZOGML9T4AtBHmDuKYNTfbFzLSoMHcXKi+Bthn6x7xulxrBglBX9pQeS1etkP3U+Q8d
h4vq5ohf+P2pfYawR9m8Qz4XG4/+rmElaAI5CPMbuHszUWEJClSWqj27RLv8UjNQQv6nRxtW8QYi
hgC2wO5BQsi9nCDTT/X5y+GLh81DZfvt4ZqLpVxEoGJCM87XZE9RSGev832TgBGei8Cq49RyL9Hd
qXroJMXdLfgbYUAlh9dULYHtdwVOwiEhVz3TNeYJy+00WGqrwIlKNnxW69Us8ZxOlaFJ4Ccq9wFE
8Hi6iBCr2DEacJKL6VaNsTekRm8sQ76AX43NRBTetSrKNPrq4XIbT1jriyKK4zpygCKF8Q/o4kuX
xZXVvBVi9iTn5OpvQuNWVId2ys7oR24+GJgx+oDHuRHtRAI3Rfl/pycXi0qluoo0e+iKm7c5yopC
8NvF1E5zHVXSE+WZFz/9JmWmHtMi5YQOaFNx/O2BmyJtf///zSGxOOtP/X0rkL7qpebyMBjlz0mk
mZfLQKKTVPfk6CxqktxZ5BIJh60rvdIh0rSU3HZAXKweSFoFmuFw5sp17q8z77d5YNDO0foiuHup
FqJpYKNXs2mKK3T8zQpRmlZsXiMGUJXUSPp12zAsiH7fjiCox9WosN3lBP2KqSVq7WkoVDqodvXV
rQRaovrTaoCsxUBuzknEFlj4CnAC6PafADEGoqah36Un3WXBUfqKSwgwm1MEKoqty+x0ZTKZXimm
9LwCzpjpwk2yvWWyS7LmKqyULdITfGLSXqwbyfRQ/1bW0JRJW+U8udE04JmkO+Fxsi23aCCc4N5Z
AabDXUaZoPcwLoowYG6UhRtvUStiYWaOlkwimPKcp2/3v2Ge/JFjXq5u8SKEmW9reqWwVg73t1IJ
oyUWjELaroaSTYe5fz85BCn1KeMSdkofsY/t3vB8C3Srp69IB9mU4cppnxudVEvylHGZPkOvR/hl
p6zEow3o4Jg2Du0kEy0oaYmJL3ZGYgRBqf5tyk7nAbR9RczI88PWBUDHuGkwWBUoR9rQmqkXBckf
Jtx6GM1RWaCQiFFP7canYoF3XqzRDeVPQemG/0t0KWq+pBY7kKgDoeVYge4VsTQQ4BRLUeOCd0as
IDXUUcGoUrhpVDEpLYoULrwk3gBLlUxeayvAJogs0IJPp66GP0K5iPzzkYlTS2E1lLApizfvwwH4
mMfge2ZojwqdE9eUGJK3LdMcGbReMC4CXnOvKXET4hOpdXQpylhPaX96cZ111HS0/qG6HQu3ZTR4
5QEH2vClwLjWSqel48iB3EaMpr8k09cKLVmJbRJG19pgEUlp26cTdMRt9rimsKF2PVO4TvvTIliM
bb8gF1fC/Wzdgu+EzVTFJLY5KiDAGQ9udNxAcuCgOdkL//9ps45tXgSu5q852upVo5gBgCWZTCGH
bSGqoKe4DeTvcDiDYbX17KpneLgdjYIhxrWIvmNSt0XNg9VB5FonVp/IVAX8gWHCnW/BIb+xXmrB
SffGAeFE35ziEw17IJ2EW9E8Xq+EMYtxUbygrFFQNVqrKuXoLLZc80HtoYF1UGZ4HoKLI5kGzHxc
qO0Te/87ZnmAyL8y5RDJJRpM9fujJs7/EWJEZMB5jkrk95Y7ulrrLEjn/1uU0K0q6Zsgg2A4El4e
HvktRbFzWy0ukBzftFp/nmvYRSSyB6YOrXsL4lq79C2r4Hmq92h6epyQsZ0wIEufna19v0RTsJ3q
WdGlnxQOg5Dx9kpvFpZvUuHSdxbH/8hEc1VW8NNE6GB3NXtniUFs4sVc9gxvNyygNuvIkgCgr5Z+
aAz6zMpkZni/+USsJDPTy3vT1ULz7bfz6jaIQllKOARTzJbWPykz4AKvv5h2YOv2x6GiPsxXdlO8
TcyU371bohBjuWJm+hu7owVGvTWfdjL1xo/kAdM6ptaavOx1ssgDEYIyppCDe+a8X0TNm/zmyYbA
ACwg76yaCNdDccdO+mnkusAEuPUW8GR2pnO06WOEqIEsZHeK4g70u++M0kQPwH1FPfToAHPM3pMJ
nBZCnx0VgdZqQVGI3e/ZfPqOkFyL+Y5e7CUSTbHSepbTyFaYcNI41K9F5A7p4Cr7hbtnHvjUO4n8
U++XCd4s91eDRW9JrcsC3/abPZgA+H2Pd9mrBo6IDgQKRGpAOxRAznOp8KLaYxDkYsgcvhE8Jp4Y
gef5OpoyimJ/SYmw8sD16shiUzCkAw4ps+EWYKWA0npEgodcN40QhMO3o3NHK+Yzy7anMQSfvMa1
WBKSU3T+OJXycBrhOXv0F0LPFNVS09vCdlp/yQMog1Yu1lpcTf/1pAcW2M/0XrfofgeOA7uTxPCP
7/RFr2FN02PHRyBHyI/5Jv6005tXBSsIeCTNo83T3zLnNrBiTsWVbPlPPkOPtcDdmNfO1FBaDBNQ
EWgcdYUU5HemQrVShd6ZVDhuy3aN6n5KeOQHz7OLG05V0+obYWNyWyvS+ypfjpEWBGhVp+Tzo3y3
BrfBMx1dsDO9GaSLu4vS76j+kbhNL7UNbWbHjPHmboqTCq+ACaG+4oXEdRLvysqxZObw0dG7Mu69
gQgs4FdKh6Hg0Tg7OJjPdEJptXuaRbfXkqJoBKQeXtbfVwYxJGFGuWlrze1f7Or8ubqOM/kwpl/z
M2iGxUodwAGMivdm3uQ9WYoK9a9nAHTAVTc/88uSivGTvTwC3A0+8tP0U6FzycncsQIMs7otCPni
+YY0HREljytmoitzEGQp1oHQQOpB7MHm0otOrWH5YhDlwSrNLcsL6PYQf0sI6Rigyznk5DxW1XP0
8uijjgAA8uMib7VYRU9qdOG1UxQ4ukfo0Iza3q7mzSGY8gMNDODk4bvZOkojQuUhjZek/3C909Yy
jPET8FKsOBQ/eLK+MVKQjyXW6WSHAynnqrNjQhfZu/c89sG//cQjK2aKAv1X5lsycrLIp8Qk9n5r
3Vz9nH454AlqtZ9DBkmC8pI/uyOa+uR1kCniOz0FBDEjfJx+ReInNOkra/PfalYWfQVAsjK4jThq
XwsoTiiqJ9IHYdNcAnyp8NfY9KBpoh02st7ysmxq4NaevXUJ/LJW957YXuPXOC8AhHU7ZhSrIwhL
12wqif/lqAGh4O0HtURQ+V6+pJC65bL9xxQv/9IbtgLexBqW7itVaZ+EqFG5/9hTO24fn8Ay8vdE
QbUagy/854Rmy6ZZ6HxfeG20OX8T1Lpztg+KynCCH5lvjozjgjnYUOHutohvVvtpYJUN819e8pbh
Ng8dp+NOwjVhTdiklWyPWHRbddvV8tbyL9x36h2M8bF6szJMDWdCND+n4gvfs3cPzOX47YNG/U55
mRHC24gC1G0eGVEORn9m1ZLqmgLLwCWSueoIk24lbN6s/TkTxLWlnB3k2kV/1C3ptIfVXAtgG7WJ
Dxj8qVyOPrvrl8Ew8g+lA/2Zo4R6fZs84+kUgkFXc37feeHop52zCE7ASZwWmqweq7HeTbyk37SA
I+ceJhw+qzlpbfiwFcQlMpgYenwqUBaLoZ+qKP5ErZ4Ufzur9ZxqRmC9XDiTmAt+SUPL3IWUJ5r1
e+vL11Zq+BHy6nFvk5poBpO8fdamJo6r5W/7IIKVF+Nqg9EexynIpNtjEUyM/WUkoCZ7qz/6sbFz
3U/eSGXi14IOQaNS/iLSSJB1WATV7zjhDCRY4Dc54Hn+T6CJQzm9dUZeFNlqJRDtSSzy81QnW7eM
N688bX4dnSz1HuEV+E+1gixbbs9f95WrCPwhN9BXMvCCySfkg//qgd+2huCIEnxWdKtpY/cWApHo
QuQgJ6BIL09p0KQAcsmeqfTpRW187cWSSQxI/+h5pLovVOxF3B/Gih2EPoIhCoywwpshttEufKZX
K55lPj4uwhsKhdlxrAuZXzpt63aBxIn6wHDwDu5UWU3ny1J/Gx81hHrdLbws9ht4b3P3kM0fHZsl
1dHQANEmJA9LYkQHsB/KP3joxKLVTdZqnnFTErS9DSzhlPJmpodiyr6G1/ViA2/vmQ1cPpNj9kU9
/nl0cSQa3QzCwjqqH/UggQ46zLZf+QWwUR0Q7DeQB9uomLOZDFM87oMWus0/mthvVv7UpC6Bxwvc
/ckF5+ILjcTg09TJP/tKg8aIDXkAlI+HVJCbqmW1MdJwUYMIKOoHZBF04BqxRu74h8EdxcU7RseA
Ec80Lgp8Uzpxe81pXQWsafqHAeYIV4sJMnDRR6pRdpfZIU9GhGUwfcSeGGHuL7AnFe1N8O0enWD3
cbMFlNx6ePds6u7GQrAPUinEZlGb6UWO19gl4QDzlrfRpcFRHDjIqN4gz/TzEa2z9n6hNRO3fUmM
I30JQSNaKwRsc6aHa9+4dfeeBP7CSEe0//+H4kiqScuja2y2eC0wi38NXe/B1nbbfJLMLAZAFYMz
rpZoW0ak7WSfRyd4Qud4+AEcscxl/eCyoy9Wa3K+hfKRhh88uYTH5tWvVlhUvPo+C+K6HgcZsC22
s6sUELNeyv8wfoUw+pgablzI8KS1kamYGiLrRK8fP0VQmi7jfKFF95t8zCdk92AqoCo9Y2TOZ66k
IexuvqwSLyDZpjfNL7ev55/O+tY7oGA0StjlCYuwYhs8z1geDrDVYF69otxeVChpoWuQc75798kw
vFPfgtn10HGCMOM/5YFJmxHUcbFB05tuur/etGGeOgSL8kG68ayUm1wwITKqFsLPbZTcv1COMAZQ
tYybKwX5bvvvjvqBOAEpvFJe0OnDGWlib9SrvzDUWYIilFBX8N8U1d+y6sF79EVfKoBmOG96iu7Q
6wbMpHgQDiF5V7zipXf5kADcU9m0K2lVa0H+LCQubNYpjxtUKNNJM7LcDPlJudwjDzy+6r5NUbcW
N/peia1MHv+7YeZPAT/7Q0HsvrPU5R0odMsk3GcgGrrz28GTN3TqjWQXcEqaMUsfDf5lgzcIZZQe
wbYfVp8AfYu9opLehx8QSqHo7feTtrginpRwesSWXTTDA7VHBWD72euDsAtfPgLZMtA/orQ6UxUu
brP/Qg9/jmWKf1bld1N0Igd9W+VDAHsChKVVi/XTbGos495Bm4hosmOqxN51kE1IxBe4cRvydkFL
GT+oIDjClHsJOPu1kqsszDMmeaWiQ+oX0aiu4VnqIJGjlmAnHGMf6SSX1UYLX9wdyO8hhnBBnXM1
z2QOiw0AcixJ0pl3LT3MEoGSab7TSQS6AahglP0JQPvuZBip0AoXpvrXZxk7xXk7Y9b1vbqcc8dr
JPgkDvwp24ewA2u6+Bkb7U4NU2LMqx4/cYl9nwQna2C/OihnNUpsjflKCxkSvNokN6FQQlIhTHjC
z2ZU7gQrJc8JkW9mnmSIAfYJr9z/493eztbOw8XTDUGrIPNpW8k2SFVfUdU1OwnxsxTZW4TVnV4Q
0CX9kzXkOdrensGaabc8uJrrp2iLO4Wym7TNvZtnieRuR7Otke/DW1UkNo7OO6wUx+/YPBdP8h8Z
t2WqM42EeDWUG0eTSEtmlD7PBU33/bVCOGU8TrWYJtL2f/1Oq6ln862ZmC2G/X0Mgr3khA537c07
PJw+5bMw00Fe6VgltTOh4TdysN36F+dNVK+ESmkdyFUKE4KIa2R5hzlYr8t3ylOtMYNFdpbcB8b+
RCCT5QLSkxYXyOKBynbCDlnk3l4f+Z7hWHeopNY7DHntslgDPxzDSF500TwXARmf20WZtYInQsbk
VGfh/sviOl7F/r8OJxOwaQTE4OWUL92WYFSRic67r7rKcwCdWdff2fEn/V/0r9yimpYqHbThd2qy
r9NlidbRwoZCqWI9HhGo2OKmQjaLIqAbWlDhsMaxodEujVIHnTRXWU3kj9OmrlUj3FhLvUGiJt8n
3pESsoazYrq+GazYsA35IMfmcDPJ/cjEodVf9YqTgPv2k/TU647BCnofdvGvOG1yNWlAgSq9uoZZ
8j8yY2xa2W5QCux1K03sJ5bLSww+EXpAKYcAhK3hyI36vzUX7usrzCT394goVQHtWzpokl41Mqki
DJAcPF8qkOPOij/IAIZ1CAOosTyWbIenAMVI8JH3MKeP8WJ5jzJ+kUIhYmJveTUqzvFaD8GXOuwA
kOPPIgGFdh2oqO1hOFYSap+Gc81abSVyzQgszsF/ID6q3cFwQeXoP7qs5IWvBxA7HzY0YZjsfkh8
vRY6CFLCL2Y/rtREt7/5kEGEo7vIEy/lw3imQds90/hbzMcpRoXBZlgymZE4ZFp8/sqR0YhQaUzV
8iTmXdwuesWArUH0OIW36znrF/wmQ/296xAb8lFad3GCbCxE/DJ4/7CEag6OzRueAf7B/CSGkxFW
lOUJ+souvvWMsNazQF+7MrybIlunQZYzTlwqQU/iDyJC+oQe1NwTOWzJdEJlxnDY7qyrWtN8DLrS
r0jrFwMS3rc8ssE6AZHLZnawO5subpNbeNetqAlOiGo94HbDza/L0RjDQPNDOqR0fvC3V1TzgUiZ
pKH8TWDrBLASgVQ7jJfx+PjUTMosivuBe9dctWrw0SvmCqmYW+2XYqf3gUVw0umV4ckuYAGQeuq4
60gopHfiX1+z05DsWke67xzWN23MGTBY2p9IJBHsMaJyJ4LfO/dlvU6P5+wr8ytVea01uVHIntWA
lIB8xn0Pi3ITEIQdKCsM7Dn01PTUEUEwVYGxq4c2vk2oIV/UzLv+CbkwPRHRECDIxMgrAhf4W7cy
w+p0QTdWnwGbT4leOea9pC8pAON18uzI47S5Acc3MfA0xzxcye7byBuj+jMZqR3XXp0EPPddJ9BJ
msRE0P0f6bpFViXHKoSl72DgqUgdo7CCQkv1c3YXBmOPGBn92f6tCWGRTnCAe+Q+FOhcKpthMgUE
scBE7+1Mdyv/ZojoTGKwO1Ee7LDaJQueh72p88JVl7S4wsKL4WbL0Cf8sE0ukDeYRmZu3/uw68mq
BYaNqwx8KVGt4IKQq54jhyVslvaIIthvXNJINmixxGB1w1tR7/ZSsTICXqlYUHh8Euio94opLhno
iSbkp63cmgELAKde1IcvwzjKg1KAX/Ww1htnG8pWYru6INUID8YMJEcacK1jzoizgWlGJwLthq2H
w33V3P6giMEmjXvWqVIp9JJ5bgpRHdE3VjN93R2Z1N8V8esCGRvSObBQTPkL+p8TuAlqiaFbJM8A
Eu75U2/WpYxd4YFLhO6qh5F5qBgoHKhqbSz/xCFDeeEqeZ58WnVTxzCweZ0bKo5QQ9ZqSK9sK4p1
2Oh5U1hYLu0h0DO9csiu3yWNS3njuVdFE7BrjJX0yY4u9Uo3S7RtB/SqTS4NT8s1XkcbAha0UUzw
9vX6SZ2qlh75wM2tqsxkF8teQla1eiIOmnnRSLFCv8x8kBBRYBZewrCGqy3+w/Vam+pPC6tq26of
8hRs0SzNXA4BYss/QXD8mba1fIupByw37WOSw24xAXfSr3PRgaUon1/i0VeLXlFV7tJyg1kt69/+
Vviq8u+2ybBo06KnjtCSwcdwTMesBu91BHyVll4h8Xbh8mmlvurq+LPrzeqEI/F9IoJeciEVqmCm
1eCR0jGCRm2aAL1b95qtgrTTe5EnGuThc3YAFj+YEA7FPdxrqzEqmNSCdbX9AMfg/wnFSLCBU2mn
TjDCHUkiPB3TZQ2imytLcOquXA57CnJbI9aC4PxABHUzZwYn1iwWOf4jT7G4utm7kJWWSnQ0Qp6d
JIt1r+MqtqMjp2b3fQfgz50KCzhT3OeKOf4/uJODvotXmGVcwPhhzw/GONsBcdD3L9uIQj0qU1EP
8fPZkmfweMG3GuQu2lnu+R5TP3yExoXJyc159AGeZixnP9IRNa05VlfRrlDqD+PDeJPqdQAZChDG
/0cPPxewRzvfzYe6I41qOxICtUGC20xdtqJW3MnuFtx6Tgtc5k7AuerVCZk4gWMdwM6sJ2K+K0Iw
TC8E47sm9c0gOZAEWrPMq+63r/80Q60x8SjCYHl1LykUCyf7sUTsWsSZ/iib6Jpca7g7Hy4Bm1MQ
mUz+UVnSTcoSwwhoI5PpBOtxl2inRA3nT39DsJ/UVEh9BHbJ/EafoKLdjLjjvl8VSj7FO2I78L9W
2OIlTYEoVlMBD5mFVFTUcoZ9t6b+MR6I+KxvmGnUibl0t4eNQQHNlzhMKb66+ZrpMX2th6PghNOk
lC5YxvjZMceQyM/iF36ByVe+PTqbgWtWFySuikEh1ovvP/k+A390c1te8BWeTYdMC+UFZ+z+FGoV
aB2MFmezGhZhXT1MTfSmD/yAa24YbUsP+PfNn9PYbdJhF4GQaJkcXbmIV0J3RlaJANFE+7EmNeHK
sGnS0s4WMGP7r3npBeNd1axiCuBqItHJ/Vj0ZN3yc6dRMTnZpmPiIrAvSgBdN81+EDc/aXL79qfN
JuJ8UH40WwfG8aVHsI9gupwz6YyqTCT1XYJaB75hEZ5/XVA2raItM8jl6vRuN5y4ErVoza7B++o8
zs+mV4QNvbjM/cPksLTQgmuIo1c1UYmOdELXNHFne3JplibP1JYIpanwNojav1kSS6GizurG2Rfc
2sF5i5ZBf9+ChXA9orYL4DMOTZTNGlg1h9fFIouzpkrDnkbvTp7KwfQQk2q4fpAVwlW8PyS5IBsZ
FMFbTUvPNawdnPXl6syLRcTnUIdhgcl8bKaUzTEBVwiEjYdF5U2OLXMeRCuS8dOsIMkL7e2lcpGG
XTSm4LymXz7HxPr7T5o4tUplShGoits6pKObcew/eql7RgKDjLe+flXf+E67+471jWA3u8P9rCy6
5k1yqR0/i8Eu4xI9DTJG+O3gl7XFCd6PojJSZazgY0HK9gE7FDbEKYVAXJyl0rvoN2dRC567oc4P
Wg+bZE5Y8phnNj4/KUZD2ZEpnqRGvbEMniVSo0miC8aPJj6844FpLwnFc3EScL1ESk95DuLDMnqF
en0hQs+LssiEDxKsFXpxEEyGxKJJJspwA44NYVmDmzpVSMbHgxI+jzTWqjPrZY7nY4mm1fO+AQMd
fBMPcXM+UpeMSnML2g9/IOS1BW7lyTFpHy36hdZrZ49Izb5vDlMRnjkLtME1qcwXMol15jH5P05F
E6biaXy+LoMMvO9trZ9J561wC8GUUCSz81fvL39CeEpNNllE+/hT8j92bYOuL7XlR0y7cqRt19L2
f9zWWNXWrPQhvWOmEo9Q9GvI530qEaIBplVDPkIeI+7me+3VJfZCqwldVlmXjDGKTBktDzEt+I/V
WjyIn0HvrdrIW0IxbTyJpTAEo+8bl7ozkLAKtKwqEUGM5UNVJkfKGNSJ4uinzeiOK5WB8oGCO+Gg
Zs6fTr1E4Q4TUAThiZtBT0M8eLs3Q6vaxl7pZFWnejwr7PeGZfxEa73G82DBKbvKQx9Ya67u1z6P
3kZAUhKSK0E1ToSNQfRENOgsw/agw+r8cYui35/vH/r9TLnVLBgKLhQmtptfdYMxU5yCVzLw9kOy
NJqUdUR7g+4jpuXxw49psfaj3AUfYMKlW9cS+rkUs0KLSKlIdm2qyGihPBrvUAVgmmoFA270uPlf
BH4qE4Of2WVx8ZnCWR+IdBvo8C88yAePvMNeaVxP1O2OuCdPEgsgEamyvWIPO8TMxQcPCCfb6Ips
zYXc9ezI+jiS1MzOMhEifXGOLLO72PPfCzM30upXqDg+XZeFC1tZfA4SjSkbnyxJcACzAJ11xXRG
5/CfS9b6gGatXqxcFkX8mjmnZk05p5iG9gyPKop8a/Hp/65WTEmgfBRjYWEvD9Y1T3iJf/VnaEGV
yh4vamHeumHmmTH4Xd18XOmxlgpX7MvFGNRl40Y4PwC7LdwW2kiv+42moHq3wwfCyL1WEwV+xcQO
h4kgm209qjhZqVONEtGgEDV7glEiWh4XzRLQGCGfWTyOveI32zZf08qkA2pGG2bJMVsEASodn/xX
1RdHsnuAUmKCu00C3hLNIjsZ/Yx0fxnL9j80Q3IzoVQrn+07cyvH7TSLfl6ehe/N55FJm8rC7XsJ
LiaEtJXyuo7Uc1egRP1HsHnIXnJ21dGL8JPCZU1toSf7SOkedMJQUB5YUDJXD6pNz6eiprm2JgtJ
vSt6OBZkGhkolrws9kYyvncH46dkQ4pRtrq6HG74crgegvVb9guMb916haW6Sh4v895qJ2Aa+18Q
CKHi7W5K6wg69iJEGirLj6BPRHf2ckRSWqbJbgx+6m3CTQD7zrCFwIcc2SrZduOdqDkHEDPaOqQE
mzUYZteNHt6zjN+O0pZHOdigGLdcNfSuih91ltZ4uTxH8on7sm9TF9jHk7sRXuHXo8lNsyVQDg0k
kq8kCraBt9vLXjt62a3CFksLRWHLs00gyBTds+ijS4tgT6jaQpYlid3ss8TUe1lg6KrRlTb/a1VF
ox7gnyzZj6OHNfX+MEnOzURdu3sslbmoL+OuhUy2HNp7EYUmk0oXfQFvLWELgALth02ohkxzleJb
sap7hyUC3xfHLw/Zoi3Ex4VozS8V2GNgWizDnnIjn1ldb7sf//l3/kTqPn6BrcwXMMEXvnJ/AVRs
vwtMMnJ2kAA32is+/A8llrYz887M9apxEJN9mnuWi4tCbK77MpwUEbmCT/2q4KCGuEvZb4gU0bma
OfEAVWheqE7kAZzVr0tErc5bP0uB3THXqBkJ/z2EzCblOy6ifLKpfRaoeu6H6HJXT2xDjxeEN39A
afgskWS7sfRcffberkH1xrn1wpjcaPdejQILW3D+OaC1DE5f7SYKAUL57m17l8KwVPCBGVyH9/k5
A8DFX7ibYRcs752bFWTfSzqVtZc36fiTen75fnElFsIU0VU01OSl/YnpFhPHt4cu2fns3iC+zbKK
7h7wLUPHtuNiU5hkkQu2az+VPFW3tTi/UOxXFA0YrbX/9Sy177stK4fJB5rSI9nv1VDNEBufRvfs
4j6L29NdAHvISEqM+6d5F+2wL3t/nJFKY0vKNv3IMaeMY5yjNrN3TRn3yHH6g+igk17qNlpsQgit
KoKHs8zSzzV5mancW/6QzRw93SQ7G7y+D3CzDmbv4H2Q/KONfqx7FHjWvGRGi8MuC+FaVTGIOLTv
qZrHFXAppB6TBW+vVHR/R/2YcR6ufsuojD9SgfPSUh50gY6RY1t8ajSyFSBejjiABaXTXsowMQQz
6eZ5NcB6tJzbpBX7OPZGPRhwEZ98e6SZwae/66n508qt0f6gZJzZyX1o5M+ZFui6zVX4L3nv2lur
XlLqWXl/DvDI8XzoxkeIcFjHQzP8NyYtpQXaCzkkqKXE38fMPXeMFeiTuyUn2dgsTt7d+eQI1k4n
mQ4p/WT8ev2T4YpGBHz4ERT71EdTpKrFuJ/MU2pjUjWXRQIu3500Xkp7uhtC9oAyRG0v9FSAiDLQ
rAR1FXcHOvkGbpBjD5BeKM8r84YzLTS1VqB3/a/X1mydhDLgRluflug4XFicU6i514ykNYMHn5oP
E82FgZOBFZbPWPQJFTceu3LNx3FggWx7SrEVCeDpv43iU/PyYNTk6QWIAdW1l3XvbG61R76p8Haq
2nY4WEs6ioQ6PvCK7ZC+rxYpaMDbw6Xxr5vHT3JiaQp44fJCK3BQcoBv7jVSw3Xr98gu6sAlDaaM
8XU3zStsKmSOew42gd3Cb0ExLvS3aELWkwo3TN4hif19F28e4h7N58MP/WwJpYS3nKhz9BGsgOAG
ZQo6KNeTljPHoG1QUt9YYl2j9FWjdQbPPM9vapRmL6wOD1Mp9kSmVZzkLVIidNFH5Dm760rxRPcy
wKTIAycscP9ToKw7S5UAeCWAYl07xZ5yFcl1l2aRxEPwNMMw3ovpdu6bQyvroyoQsRMY1VAuSeuz
OFwW0AV1+A/+b9WJOrPhR3kUX2uS+cYg30xhWYNqWpBb1JcuO7blosZR0RCeLmDafy3l1r8Frw5l
ThElpWaExP4YpulpfPryR5xksOYDqz2/UZOw0yGs827NfcghbRpkDn0BC/1ybzLt7Y9f7pjzeNBX
UlMdl1NszmwU7ovfcejlQfLWEjSC0SYnW7czgcjuUiPj8CocDSlNQclcqbCPXnD7euuCtSk63GvV
csHW3wCHMchJeMeh/h4NGm21WKy0xSVCEBbIRz4pkNANIOq514wqScVh8CFjN3YPWSgfIwR6c7Pb
ZvdQ46L+1rqR0BbjcIPF4X/HJjdZgE/DMMy14UpV8Xebg5EYt5pDdazwMFXOWPVRYSldFCOXJAQR
lpo86C8ZoKGiQp2rEdbc7DqGleCOfz3IZTygXgJsVYATxc4oU3XOapiQ6swr2bMkDU0vEk7ijX5V
WqMATwLayn6ZLdX1UP+dDxo/KJ5xKcSKbN7NTylMqsQB1BxiOpuWw7cnlykaZwU4jWNk6B8IrfjQ
T3EwlqWp1VcdiMWy2ULOSvUJjf50yia/3ER1dw5kJEJ+cWEettBtAaDYPmHs4kkY9V3gl5eWxZ1Q
4FkvnYMF0dn4l6gYwb9jqasHb9e86YX1hKKSMzsqeIBCsor9qOYV9U+9MT9/YNCjN+ud3CuynZ49
wk/FlHAZRh34tyLm9f7dF3Z8Or7vTsaA41mUK11c3Tdlrf8CW5uO5xbid4M4R/ZeXN4WZohnrCdv
CYlYq27ssWKx6KSQc0Ud7DR4w5aZujWicPwS1Zm3ioc4Dh8HrNsiGMjFZ8K87GKw5hmd/w6VkPxm
HPeJ/F74V4FIvvPjPSC23xv2blp7RKJxkquTzCIdPvXqTLwq9zFnrIFrVf8QTvfEUswipQgnMjrM
AR8YqJ4AXVgHQVJKYysFsIBTa4VHdaxqVPmdaosqfuHDScmHEbFo4ZmYPbc7UbYs4bWgdUwjnmlS
vqYDokWfKp07Kzmm3t3CIFbqcpdbn+ti27v1G4NOQMkzbcfleTZ4gwqr0dU2pI+B+j1n/f7MdUTT
I9KMQeAc0reNxOp8zP+xOO9LQ/Z4YquOqsGBxc21QBuocZ+0aHeT5UG9S/dwdUnuuC1CEav9EIH8
03t3pyiKiVyVKE3HT2fhwz0lpwBWreTI9+GtxJjImbG6zbx665IIbqjAuaoO59qbaa86z4Q6Dr0R
iQkzwW/aT1W+aC1T4wj2PokMizlNO3dCJNeWN/mFsnbsFeHgCEi6XUDeE/YTrdFcLzlQUzONvUq1
sGCHYqOHWJiliGvNH/YquhFOfzlqflGqP6HnSb+wHLrGRu1gYNTn67ze+Plu+i96HOxrqX7TBo2D
RCYsggVAoqDJT+PYwtZW4GLvjfa6Izfvxy45o19Nbh2kZdCoUTKvU3aF6GJxV5VAAhfeQN9KbKjZ
F+PWqoX5JkyQvc5ez77NfzuWW9DLzeU+siHCrii2ABaaVQ+E0nwsA1gB+09Bo5Wt9WoCtEDvAxF1
21kfMLvhv8XTDXdHZd97M+2tiydLqT/nOQROlJEIv0hlQHVvmLyaNvJEwiuwNUQGZbCGa7pcU3cB
G0Y5ioaNWUox4mxP5EqZZ2cS07iZEx9/0F0PbRN4cvxtyT72IQAsWUouwPb2YGrhS03QUSKkfDeC
FYdwGGT3ofFgVRxaMHOF2f+ooui3M1A5Rc9UCJxlmR+LA8SMukNTxclP0ofuzsv+gsHWO51Izt1p
In8fNZolnX4sV59uYl4AFvPPq5rX7ryWCF69/q7vfzKBgrBaDGFQliTTxlLOS0ItH5QIQvFS0hAy
T6pKrg05zlTXWI/5LmNqaYnoKbdfOw90Lps3BHXGb1TWwcPPbKCkDQIMQgAZb1iwyBGxH8fjwMMM
a3doqc56Ez+VpQ4t9kLxsnKqMUbrSxz0k/DNHar41cKq0xRmhwYkSfTqHbWiE7MF8SGBwfDVhCui
FHdOYErzYJLlQR6aNcwAyXH5XLSmqg916ioo+0jCoOHLFqXEqAaaXH3gbwyTqkc/FBhYAat5USqw
1HBsPq3u2EXgWIzLrvHmjdAcx+HrOdnXF9gqxJm0GkOAOLTfikafUhy017jLQGmHk2RH1OYChQIh
+aYAS/Lrt8wLX1T8f8UKm3fzXdA8O6o2ahf571hb9D58XtDAqpAkMhrLRnC0+QLI6RVFKdTzDC1X
t0IjVUsf2Dv5uLvOsGp2LAbfbLcMQN2NVv4U+roPSg4nb5bz6DqXnjcue6E2C7P899hRgE0vjryO
PGoqB5aPIWSzxl6M2S6oJ93Nlh0+UBDUpaRY2z82UG88xNBtqVOB8AsSn7cJtjifprsOco2ejvHm
ySsTCQ95vzwQUZaih/OkGa4raYURpc8OZNBdtWkdFkXpWyjZViOEXqE2v2r8A0QTgivm0wapEJ1+
0bQBvspYGK4t2iKF4btTuouIvZvRuQvGgZZ0sT6vpN98iFsFlTLpflrkWP7mk18sVnktnymw2gD9
NbFB46tJBVgfL0avoZD16WbWw3KtFxNXYeY5YsQEM8d9nHK3P9nTmYqrft9vxKo1oGQezyGcHfuY
m9bDLLd5gJvtfJsIICjioH7eXntgQWJmDEver58zLBdVIWcCjX63VXxDkoZITex7VdsQ66jvmqW2
0LIubvvXGuoufykQ8GbBgeR2MxoIXeE+nVqB6UYp5dLg/+WIYjaAvGHE/zP4rijX0iRgI7DVVqXD
4EYWGYUlmQ1hk+1yERxKQpAJpLm06Jnzq3EHNcdhsjp4hvS4CP2C+bU6GatWlk4/vqtTefbyXevx
s/BMvkytt0Yc8LrglHiziyDpfGCKAyhmMFQWYYAO9YZkUtK+F7gVJyxG3++xZCYxCmb0tJOPSoi7
HFjG8rNQAQIO5uXoKlscXGk2w87foo0O86b8wU8N95CaofMTwTMIfFHg2Us9jDCV5Y7GERZPbTw8
43kUpNJdEgf3R4pWODhLPfxM7tJGF6wbTha1m31J/DA/HDhUl1C8FNZXeuwrVzjxm6kHe6991oUf
jF9OkA5+1EaEfonftItAcWwc5jngKYRuGJbtI1VB3ZoooIAwAC9D/MVxaKY2NqQDNI7m8gXASZNq
koy1q0ApUqPeowQ9jUAH21FNQT2QmDJW8zK0I4gb0kDXCqFARf09pGESsl0BW9Gl72JpFGXaYwSV
Gnoigc8/HuyL2jbx3aQtdYP5I8euiLESp3fqAOkpaTcicPX8XNVt/+MkkNNAIhNKg2Dy6me2T865
tLh6+vAzz7ScMF9Idv7v6YKMfFQnRz5iUeyEeFBlZntXMTUhjFe3DU4cp2h0lIq4KO7179wuxpLy
U0aSlWZn84DTd1YUO1/BB3h3nGQEGLMNI9CNTvCd9eqzWUO7eXPp+aoNS7kMinHRtOCmGhyneWTC
rm/Vk/3mZYc8maYLz4hiTBK4uodEfQxQIN8H0tGwD7W//bM/Og7WutmJn4ReRQzGjuFJS3rJtfVL
cUY1pCKFEzAIu5HXSi3+7tGuUIUiKxUvkKe16EF2hdjvSS1515ueql4Tc5KMZ5jpuMYsd1JhdcO9
GF0mDe4WUkEFK5THsRP+SoCYM8sTDYy3o3eGUubsq1CsyHCoNxrmJr77cpoPcSg9jdk8UEXfId6T
EeLDsQoinLn96uDTi4wcF2feusARsDLgCzExFzzgKlK5QRlnL02O1zMFnaMmxdf2GP/mYBDU53S2
5mtTHjUBDnOnJ3SL0RRYbz9gPNBb86gImBlU61cMSYd9nd/gB+nr4+OJJMzPYBjd+EhvHsVaJWX1
Njn9lvkwDooVbKH88oojbpTd5XxCPdUhQxZSTnZ2/VHkebZ21tHqsER01dAKfWnrEaYGDHgPdZBZ
Te80HQQkR1qLqhKsSCP5iHTXGl+PbGbr2EDx7LycORmZbq4HNbiuceOP41/HNvTWV5vIIwhafoas
IimZECWJ6A/ATs0kkING1Bd+0x6CFzchNREiy8KpkCw8NuVhBvIwgQp3jFjp0lnQNNbwFsFgs26S
uNkYOf0x1BN7K2sCm01C+FME4rC7I5AL/2CkwdlxunGftyU2E1duVMn2wDMW/DPNbPvVm1z5/L3h
6Qw1BaxQ+VnnAIKOmVLxqE7h8Kno4FkbHcm8JovcReTJB122UA8daggcuj9FxmzpkGLHz8qZX2sM
/A0EJP62j67wKPZ2eokvCP4QyKI4XIpv+NflZy05dhMn/RU1dOpgoaSI4lblQevScwvQxxJlXDnz
I7U1v+IooavAwYnbzrw2cP4k+B6/6XYnACuUE/FRg3wfs5MYjwnVNiZ4+62qRz1y+qjbtajXmTMg
3OUtGU+G8428ZWZv6kJdS9mpVHXLfMV65rJNfSsQWiQ9LjYYHmEHuk9WCvTXwHZ9ec9Fa8lfsPjs
lexpS8Wyfp8gcnpkBqplwiLBn+v4amg/7Z00Z0ctA6d3p/B80I56kTzxn1wanlWFOLq60LZGbDBa
XcTbfm2wN35qoSPtM9ctTLR87wVeZkf9MOmxFBm6dsBeXei4HYt3SlkhYJpJLWzN0BRs0e7Ps7u0
NXpeKlKturb+yg64b4CX42XBwkOu8VAPI0eSo4f4GXZYaJLzCQakyfe1m/9L+bv1YMvfWF0Yeq+U
w/bF6njKJSNu+LvNc45CQlZR5msSTBUe9f7tGmMr7Joxndph1VOpzLU7MGa8jqD5k239EIOWhfjo
TIEccSMXN0E0orN2TXzxFhNNyH+99edmSKyrKDAYbt1KEsz4qlJnH8KAgBvna9zy7mo1Qe1NUrq2
4pW56uIVbGiaHmY5c4eCc9LNBnO9SdU+TSQ3xV02F0ctnvTTB14OIaiVvY0DQP4Ad8Z4NW3stLRK
eN4I6RwlRMzJMk6Z4EDT3XbuM6WCbRExL0WSznEIA4vR9bp3zCk9zzzcoVAzyyct79OnQveF5MrU
sSr0hLzi5dihAKPLxfwZCZuoqlxR6UVzx9hAL7hE/VUBw2MzZFOJSz3Lr95zWSIRs4qI1t80k03R
e849+SkXpoMAKP/xCtPARSzk1U4lwcA4Tw5LmEXmDyTdV+sbotRVrK1bUcfmaG9eVTo7ANjkOhGr
SiodpmSqtwSyDduJIS40+9vsOUao2oTsquFqcGAhhsvyJtq1uDoT151v4Xe/edebwCazK6XXjO0h
0+m3+JpvbHHlnvIneRR57l7rtn6aOtP70IkcTgJ9zWd8VBxFmfLbBOc7TzatskwV+IedoAtGUUK5
XRTHc1sRQadunayYpAD37CHuxO+0TQd6fTgIhYkjmNEyhExEDU14nuRuEMf3UeTGXvL18mQenUPG
YLc0eV5FCvUFJlpfk6UEe35pziITni2i9gTUzMbgdjeZEDEdk1Cf1D169evzWgCalRTuJEEpEK+z
bw1MrTkGP4NuY2YhcFg2zdlYvD2Wkf3+bRQgyczS5rXP0SCsKYYAG80B+2lV5ChqMatDsuzcNRnM
ZZYDxoAcLmHcoYGdisdqMBzyakuZatUlgByvvWFRLRKemopzH2dpDR7iiOAMYYf9D/4PhJZZ+Xzy
gfBWHRjf5Y9kz1K0YaquBRSXOuKslH/wifDKRaaTK0mi2faPW726jIC+QLvRlQ1yOFvl4Obq5gAr
xWd8qw3d3TZN+odoexfa/yoojDVlJ4sdC5uUKbVH3Poh2sQd4hH7szFRaBr4n2dljLLY0FXa4cyX
dN/KwN3U6F/e0cbVZwA2kdIXElIZxWaS0jwXQISRln3sevo92aA2XYknIXzV2loafvXlQDXdgwlh
fLJV0t0OURq0rnvACfA3xFw+OMMhgEaquRPJq+vciUD6UYBNLupdoImOKYMkccJKuWxa9aBHtBFP
52YYCOct34KRp5ak1wQaqYkDn9PRRh7qzZhBGy21rvsUcylb0jghsNArDeymchp678wDN9F8WRxO
7yahH2oqdssJMg6nWJe/ZrKs159ciMW3Xd0E2dl8M2MR29GgneGzbJ0/zfs7D59gzoTycQTnUPi6
mfP9kuPsjPnlLwXv2tKBsbMfoOw8XkQF0EU5n41KdGplebHoJ1i+i0yfoi3HoIjjYLcFZ+bX1Q75
7TTJGflZWwTTJ2Lyyffb4/zQqImbGo4Xcnb3g3f79mf1vO9zkD6NqMM+4b1wGbFn/xAWDF6mYOMh
npuc24tas8H8qJRhgOKFJgVclLgTJpuBufGWTQYEORI2A7Va4OqwkZwhZS1MtqJkvNeyPOFTHZtl
9HT4xOgsvBXYqiWDUiS+qWjdHy3kO2tRKlFTgM30Ar9NpmL/X4plderUvXHRVbJoSreKKgLCtVZa
bfzGaePtsBGlSt3fa8LxuFSnE3aVjwFHWwvvbHzZpfhgfLfQEHzA6TmC8VGAdfD4M+n2kUlSZL1i
tlDAXnapn9sFaQ4+b6zx4IYzh4RiFoEeZzjTKq6x/50s2m1jz9QmkR8wSHgrVjXGH9AOz+PeHkHG
Nr5JT7Kv2jDHy36YJajoPuY4CtSIGda5LmyrqPZBqMNOo0yW8TQ3O3PoX3WwHShs7E/m7tab/Ngg
EiQ7ZkbAnGcGh5IAQbJ4kLjV9+6/aWPSfaDR7HcOFQekz8HhRxa3vw7EmS2WUswrg0nksqxP5EZP
+tzpwdfxLJtN9wlwkrmmXSO76/fXJyVWf4HA6UGRFfPbZ2cm6fWiTBDkPnB4VR85ADe/OH80AxBO
nhehy7CyWxeHuzRtO44Y7K42ycv6Rji8LC3D0O5+Y9JADDp+/32Rng9XEjsXNNvxaY2cfA65ZQy3
pXhCo4dxVy8hlCSH6PSB4IJWdh62LxsruyYcwIqIwIkeGSCikR9IwaUpn1CXjbVsgVb1oE4q0dMT
Dt183DikaJTJqNWtUHxYFMDGEUJhtryWHjBMf+q3FTKV3PWr58pRj7/wwhovFsUw0glbEhb7B7gc
AM0rVjnh16x6M0f0OwXI4V0a+VFHQAhERX5fg65enif/yKMvEwcueBL0Og3gllYYz8oTJsa+/J38
d/HIPxvbmO5Gg8UGg35Qf2B6607vaJ7Y4hd7fYHnA2EzTf+wraSK4YAqUJNhh3vXyKZkcCQi9XJg
Eh+kbgxCGhNce1L1JjWWyihk7Hxt6snYSalWQ2Bxji4Ky4WOMu3cSLZ/fjwKbZIkM3hDRyRZfgz7
9Jjo4QY2dl30c1C8+CUIbTedX7vOUkteRmzd1IbHG5kViJu9cJocl1CUkc0JqxXd0zlOxr6AEYth
E6YYdQIEoUJXYd275Eoi26ypo3NTUUm1RgK2aI4BaY4iuf8vWr32z5bt5ijNFbuFFjSL8SiWgvKq
VMbjJCVsuyzz2jmlTo+RMYX+gFmblXr3HB5fkHu503XReobmCXLJY+M1gCRZhx01HXpBS7707gib
KVFOuh2tmVR01jM5/W6hihHnnAzdozCvb6T+enbw881qDIpQ64qYf35v1bV0/bagDrFc0gW0ZF+Q
URLp80rw/LMWg31XEliD9QpDDxu7DbK0C9Kls3cM/4tYk7t1hivGLl3OxTIE4Cl2PKQ+V0rXaKDc
EMdJZCYQinq92stCFACMpVKCWOdpKxhD8KcBrEDRDSZQBnGLzIyO3Gausj6w0ZtTtai6q8mq+SPA
j5/ngfLrgVPioQI1Zy9PpBjEnZLgWOXEUJrBUthIetqgJzXaTDHEXZnR/ZRYcifpQNKXGPAgBHcw
GjUIs55H4hltADRiJIhi5uxnzrTVPFD8+Gkj+fpKLcAq1kUYhJ+wPpUxGWlhWOh1Y+5q14N0FRQj
zs8cH4ztSHUIn8eevjeXns/WXghZMAAKB3vl2VpS+MUKblqBaUcGqI5waBxxkv7IfiKkjqdjdTsi
p8N5k4pw226Nso8LhU+GaEAVcMJf7cqUGMGgIanzz96oV86kfQxvxELQTjGpMxVEWPPrWSKTDXcR
zRzJaMoIKD01edPoF+HU8aaBSNEHUcOhXKIEhNbi7ZnHe0Qf5ZBUzbLgy6fG8G0r1BidHjAYyKnJ
QVEO+lGHoxuC1MN7HQVByt21MWPwdkTW220RhKHYEae5Am1OBAEohRqYXRl9wjrT0qDPKbYMq2Kj
ku5fd0+rRzJde6QOeTAms7wfFSSAO83XOk/wVrarCgqrxCAxsS9321lejrWvjfo31haXzBtTDkOH
xX0CEVep9ZTNyTsu/3m3/Z11B3wBwY/baCTSOOMkq3h7wxsW5rDiefFWaUHTJBemi99pg/qnb5t/
EuU7jgD03hlBA05QpVi5CkG5odpEzVkbNhYmpJ/+PH2aMdfnGZffY85/vxsSXu8EfSZzY3rwUNbr
Hpbzpn0cncdpJJSqm/m9iRpElE/PA8TcPsG+/1o4e85ugVHERG4/BRQLxA+SuXNF8UtZEMOqGo1I
A8eNrMsve31qd71VLPmmCzSoTU8RoOVyyo5JFQGNJaCdrUE5EAV++CNCSIGtlxFjlljxZuR0rJFC
tL9JMdh2cBMxmKpqe37ccnZd/Bxf7USzu0UrG/usuoWIMAO4kUgPe21UeZBEO4T8yeFLbu8s6MKW
jA6nZ+ejFCrSinx0JEC6qull3KYwWtyiLEy1bR1YBtzbSNNdtZD3CjtpbvvoW2QLo5yJmCyihQAF
JMo6Zyezy6BNm317gRt1zBT/i2lyUXB6Jnm44tX1pHeE7BUam1vQlLH2byloe/s7XiEo8Ucyco/t
XGyXQGaDONHQiqZf6PlKyo4cvBksq4jzjjFMNufkaPrjjAlhjyosOJvosn4L2TWdAMalA0e/R7Sk
DqYLdrLJAzTOKn+uxNqOuYEACvuRFeG/ZlgIkXUATA8mQH13h6NKpO9GLRKnyFyHQ+CIxZlNQp0o
JFX7sq3UExld3jJki2tmLytoQihG/G6olc2+ektkJ1+pPnI1Zk3VO39VkB28UaRdnH+6oPTG7ilg
hAiiliEs7DYvR5Txgit/pZX+9MaIQhMDpyWn71tcksqPd6hYxawMmigye/wN6/SpVF6dzqPT3O83
BkxMdnLQjmCPbxG96djYSfyO1Bnu8tYXkXQmtBTn2oit7j0KuRSxUQa8MLKTLkenyZZ+D4MCqHhX
/5nr++Hdy6skRq2mDu6pXq8ofh4Q7Zh+j4pcRp8fWScw8PAydeVBzH+lUJnmRYvrzzLuUUMB9xXH
uEObqUwslqZ/Xd8WUhgDZX7n9Dzv9EsU0Mruw1IWOEK1Jay2FxoxxY0OFnAM+37C3njT1A1J7Sdx
ahLFG/6y9w1bgEBVcLSPRsmz5dcyCjsDSx0s8Ej13XKRM+z00Gt/3eb5oem7mqSEWjF0n2P7QG/D
qgMYKCkUGpJnPqxgDEJI1+/bWw1OPMzay4EuwAJ2LgGqnhz/mNPlrD6O6u3km9n329o27wWZE1MO
9BkXLMBfkIeXrwD5HIiq9o8qN3zGnmJsrnxG8y33xVvkEeKgfO1JE9aJqFBK9bLE3gVbM6PDcG06
I2QqNg6JJk1iYrkUN1U/hcST163kEJsUFFqkA5OjR9FbFWb7MzzfcWs1aev/EZzTtVxQ+7rfvew2
eGCx91xOjLqxciyHDe5B9hpqvMJD/b4K9u1/1twIKRMRm7QSrcNwaGmGdmmSfnnQX1UEgmgX/YTz
G12/VTMdwGOfaRpTgJxuS8M9DRZmoEusyIAjepTnoTDoeZIgqa+5S2bkKr2iTVRXZB8dbhmAv00l
3UN7PB4O/A9KWHrf5xxCmM2f1gcQkANm6zVfxurb06zkvRlg+WuYxLk/c25ptlBgsFmx7YL8/zoy
kQkj220L+MbZ+Vxckp5voMzDL9dyIn0IwrARBuUhIKwAzSq8P/e5HIRVj7fyl9wiF/yxbiInC3yD
1cgwnWMwNIdkqrksyj8i59Tmo+VEE2L+yJCl2jazshRJWVv8uQxlmDeGQmPsQsxTWUfg7yMsFzyd
PREGYH0UwlRJrT0+898R/5Q+TVLNFm5OUjsrGLcLrmKBVFdE2f/Bu0Xj5KfHvJ512LMeVHgi9uWR
PHBokR2JH6SB7D7TV/LwUUGeQpyWJxFnLG6yevOz9mBapJLKAmAK2WnawvwUvJDycMdW9UxjPloR
WMG5HcVnAyWx/3X7eIiFjzw1ePAP8BauHUZpKN3G6Gjx23RpK3T2fwUb9qhUM/FvZwGFQNtSUfyX
WCWQTmgLbwCTlAJaOl0WRaQUyUJ2OZYmd5f1xPL7uM+hezK+6H/L6YDnIoISaDHJ22PLVQyaMbU=
`protect end_protected
