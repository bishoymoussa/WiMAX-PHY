-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
xUT+9cYdblAJemMf9ik18lZB+m1eKgqJiCbTQNwyFe7NYbS7l/LSUnlsBlA7DANDEgZI0+wZK+QI
HmHoqXXEGXhsnIb30RPwAHXQwTPTc7NGLPJ5gDIGjOFTz32pmIpSJZG56B2ss6uzRdkJrUyuhtrO
Fyegqr47xv9ZUgnqEljwlC6RhmPvN5sB83SrRYMkHjMGoaJFq0nfmLyIQOw2RFwgN8z7ts5Vsp4j
OyfP9cHi7cJI/B7P/rLNcAyyEMIheZttlr0KbtN9gQT7lhqFsrS+IeXMfNw7WE+lfU9t80UqpSso
8ip98UYm8EScBS6W1PBDLElBjas4UT8yhnJWbg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 35184)
`protect data_block
SANyR9QOhqLHj8rHCpwCUKo/pVZgVc91jW7wFsZ6HPqC8P05i4Ka5uo/uaSqk3LaQt976JHJ2K6d
eOCkyW72Jp3wwpGKt3og7Q89tkJbDfDH61nc1MfxM6By9eWkF9r1xENnXCPInCKyORvWSTqMbxxN
htKVSMkdh1NhZ8anvmqauorZMIj4cd1WofqXDla3Xf93shIFINSCdgRzKfLObHxhym05WveT2Z5U
/OQTIw1NpHYW78a31VO97JvLAT6R7tzLbVbqcKQZzCoCk7/fI5uiqDNdHaMw8u9UhlnoV23jOBrM
E+EqpDiZ6mu8x+8qHKwZCo7UEv/pN6jKCLA3ddoydRajzAZ0q9A4J+zlfGsRBmGafn18ppoX1CO8
yGDi4V2XLaSXqJOsiRXoDePjXbY/dzPbX2DQZxqwPHcMG5lSWCS01I+SqeSJPDgNguoRsANI2Avt
uvZNKlqzG6fAa2ldlrZKUNIbauCdG2g1jnzTR8awiVSDuG+QY1RK22lOtjqF24Q1i45StKcD6cwt
siqUT6ojILYgYJ9DnwHUCgyT/ou55Q+SzSlejEv6i7AyCrbmW3E6rqNcdXEzzSn28mHtN++du22V
SFRJjnOV+z+W9vKKLcVXiDAjhJ/ExJQq1g9YlVk3iR+x7oTsCEUxtM681pzcmV1Z+howLGlfyo3F
1+qJmLZ2ZoBiL6lKK88NXVYMrXF+F6ZgBM1sCt7zetdjEaP0nApYo/+ukYLGCbosh31821cykQEf
m47r+IxVAowUWPaeUBpgi0qadypvL1GrJDStHT5YvkoeQSfSLfPYUIZWnjZckIZnhV/IMOvFbQy9
UqwWHjJWntmROcSF4HrCq6OkUO7T0gOAu1p1iqLKNWNesMXza3tKKitCg9DqtYhNGsYPO5ATL9LR
5Y+yoJCcgXbvAOeG6MKjKlOfqKZ5Dc2hXYWDnNlo/bp2pXzMmBQiBCDrcJ955n/g8oyCPN0VicMT
OnHXXg4mYG4NEQdh79ywUvLqiXtUf7oGgGwHIe4Hrm2lRPyA+Kz7EACIYo0ZyhqxTnR2uNkTWe2b
gZnm8NuTNYtPohWHQcTfy3tP3fYQ0QJrZ1kvDf3vmWgivzWhllKfuwiB5iH3XzjzfBAY6QZu9lyC
h4Coann77hj+XDcHnZpPU7X/Nyls9FIQkjYX3Ta46eplE4IHJZJUNa3R4685zBGGqMAluVE/tJvn
N/Bss/OEv5BAlKLcj/Iq65gxiyM891ROTi2l3AgE9ST0/FGf5YAF53R/GtwEQVjisYFl4XpTaWgx
jnnMXJDF11l5ZUqiaHlyc7LvgCbcIJAdIulG9Yhfd+WV33ofteCmyCuy5mLXRkfqTvi0fw3pEWik
QOPp5mHYOkVgRqBruQvP1YxGgO71bJcCB+eI/0d5wfcOQZM2EQQUvMmpNu+3WWEHBBWGxcETfyHl
K56MZIXi8B6p0GSG/4I4Kunwl9jeMX0NC1CSUy5lCtXGSc2+ulvgJQZmolBLPbGXy3EXhEn104ZS
D8mMrX4JwIe5oMZRHKcbOG+EI0O7O/2KNkI9aL1mvp+w5QsEVZnl/s79SUeAW+3QDgUcYAijIPkh
VjfUBBCXUeM7udos6fkATEIdU8HAOkDr/+APcyo+2DOr/WL1UuUMRd0JIQ1KMM5sxcHAFUWU7PLN
5LZ3YTDRVTobPo3G/XXksgdKpZjusNwuHwJxFgj/1/MyULPUkW1mHeQworaETRUN3wK0grAo9dVU
CrPH0h2UZJNMeO7IqY2QPPQ+/RoPj3iz6H2bGSFVXrnvISZCpHux+dFSLR07NetBekryY8Ah1xU7
4y0Z3+4JW3wuXfEOIpFk3n2ft5pGlatDQQFsXdrtmIC2pTHf6FAU5nPDXHo3dllSpwhydfjFwBaF
LWmQvnI9iudb4uI8Wok024xO5EOP51i5n6W10NY9TpclxCTHgHRoSYPDhorWsPDdIDLWBS7QiUcN
FOwef0Tj7N3tEhKFKOMKIiTIQt5C+GWjBp8cqL719tRjSFaqyXz/I2vTv7ZSv7SY1evlA89QX1I4
P3EFYlXzSRyHDJ3RuGJx9iqcZTZrkyl4G3FPnAqtJXbvx/QiFk+ILFSXeDx1LEAYYKUe9kKhbjv2
f4LcFPg6Vqx9sfPvXtunPXQDWDElKZmjUqTcdrV0jjRQycDMHC3nfdLyR9KIbv5f8Vx3R43GxO78
tTv8Ei5s6NtuuJz0qsTG+Nw2b0zRu6sG9W9Bo2lt9Y7b0jUaJRDnAiZvCTAyjPKAMoIBEqFmOL+D
zu/SzACuHzhuuRZbz4Oe4YDscMED65TiB9cc98NBTyiGzdGjhOBYPztk6wdxn0ETCYvbcxog372V
kpvy8zpBK5jJAqOjuEQ1prEcCgZyUy0cIxJ8hY9j+ql+/fiPzcKHi9yCsHjAhTRHX4xXue5aarKM
we+wrZ9uc7f4CvhuD+89igprzsS96xNo3zGYRP7Vm8NgVBCiOJwkLfJP/2Xxoh42YhZsRePonZtJ
Fupovj7bz/wpFFGYhQiqXAAFxoe0M28RcHT8UL1zG8/as2pYNK+qbG7fey4O7dPx547eOXSJYCYR
kwG56F0xTuPDNydOM2OAKZJV16qL/KMeTPO/vF+sgEPohAtgQVnLSIjejFclVkAebTPwwai701yk
QVw4XVCq21bQb+9cFKgku7NUzV1S+OJZ3GByYeTTdEdoCVjZAk0qZ4iYRUte+SN25SHJMdaKm0UJ
qiJCd63VEUZ9WWnc+5nPeUfIh0z4BzU88XDMP4B78UZ5C/cTvAVvK0K8P6s1BZDmGRHyup2Um+Fw
lXq8RIS6ZcRwg2YE9BrmQ4up6TUAixjIUNYrG0E+RA1vt96Kh6qo0TI4Jtj1+BVraEbRa19nhteY
Cy60W5FuW/LXNSuKQR5V8biIK9P9umAXqcoC4gM0prFOw7irCrdOiZVCpoBboW8xI/Espik4A9LI
Qf/F1XFebEz32a8KJ/ns+0vFhs49e28nxiuLu2OoxzWTrYBmgCTcj3e73c/ovIIlwhczLMRUTWQl
KgF72MOiRWViuvn/7XLLHX3oD0Z532CcYOQyacxoVGGDTMR8VcpkXMxxrTfo6vIpAvXsFxpjXZIU
+R8lWudQeCWY8SmMuFe82sA/B2gNwb7PgbxXHf5xLVWgcyz9un3UjPDeWfSpEwwos0ybnRuIQ/nQ
dd479BXCmgQvkMqKpSuZzdNH/ZzNb/ppTpB6FEzgxmBLcWobGUBWgcQMzfdL/T4Rq2U/iIrvqMOu
x6SOBEM6vfLlttUtFwW57mTugI89nEWuDHTG8Uj3tUPuODlN/KfeliNdH7bOH0ScEY1wqr3NlVpN
0JGj+fspjSdiAQZuUjUIJ1Yf2IeVJN6+vnYzGtEKaHIGvBzoxa/2EKf61fYb0tUV7vsM4JnVxD5v
rF+LL8Gym4R977Ff0QpkE5J96sqGumYT1/xKb2jJ5JZMk/C1AEPsyopQyhCwQIW+Gx6iE+f763D6
dEL7mWvRy6wwbc2E70gd9O+Cg9oizqBD3S014DVPzYv3OmNNU7Bye9mKnaNRozKLmN5VjogRAtmW
tU+fkyb7UqSzbB2M4tmX7RZ3ZPIzoThslKfANh7gvW8YVMGPE0SDDGP6ha4oopXGEfthcqVFeiw2
ojBUKv818PPLBJaA2kPpkC5UjRbxkGEQH8klX6vxDL1wgnQQNW4F3WWr3dfif5lPfhgDkKjK7oE8
rVZxmNXW5vg7OfiKvSsz2IyXshNBIEZ5UT9uJNHbKsjSouMuAITLEgDblllSY1HIbglZ9Czgeb1j
kOF8jSK4gXsvUKIRRKpUte81Ur9fF4195w/pJyHRyMm78Jav32MYa5mMclt2Iw/2NlCVijHtAo4w
+ieCY6ITpO3CrcDB0TuUlIu/5oby+IR7Po+ue8/zzfU+TlY8O6PbJL43ZPpmCeaHY6tX84ocQxDr
2ztOE4LIye7kBVKKLaqQ2Qh4sbpdq4BAlRsONEH9wrjmLxhFS38X+OUnxaYTJRkL4a7R2ftU8GLh
L8hrS3pBmodse30197DTqbqAm6yqJiW1Rtp9yBW4B+XDQZpTmIVdy4hBFIFm57Te/tEa/EJCCw85
2YwyLk3xrjYbbZX7wvC6yO6DCHjQmoA+xLTSBasQ8Zg6dywaqEfAU23MoR/9pJ1k6MtQlpRvWjro
HRkR5SNTuHb1AEvPIm/v6bsjZoQqmEfTZ229SFc/OMf6CJI0IbkY/rMP/l5luiTN3LqKJima0ljl
LUiVluM9cpxbhS7QEJqa5fDfzpe+W+zd4YiHKaGS33A3Zjuao/NIUYiqSafAaqhZRkqnZj3f1abO
iK+V10S24ZMwg1D4kEsNwBHfKyuBytyNmlV7RdG0MvcW+VX1znpKAHNYzsKKnCBUqFFBneUZiH7z
2QnGi24Ku7M+bpIVcwxa6JtAmpIlIfSqbllxZl/Xya1A/SVsEAEZGneyevbNMtIAtVZv79pYM5C1
6MZTT8sYzRml/Vm9VZgQI7CKy2WZX1zXal2druuLQBG3ASRhvtHMzlzM4BMvi+vzEQDCerutomL+
TOZby53/N4o/BxJMVs54RRmxm40MAV/wGvaoeCbS5JUk4wSDIqtiWdiyaqrSfBldhm54m1BU0ytr
JP1RIl19BECmlII91lxdg3z59lI3O4LEjVvkLK5znNvzsoERxiv7JKMoYiEJoT4ZKhcm5nx3OmUA
JS0G/gv/lEiI5rP/qczMSXHGo0GWCaQgi2o7UefydChfmvos/uX1b9rahVnlb5j+ruXlfIfBu+ax
Rw2eWBvS6ONDfT9pAT2fyAlpSVHspnEkePq70AyJuSQd+q9i/39dpJZ3lzeshmSUaVvuCiOoTi6/
UBNpYJVvxXBgPoxFt1GMFffByumYj6KOJAQBQu195hSZR8tfny1AEIDK/c0RbAs/s1Pcqf6xKefJ
fGrDg9hTMIypZOKlB5tvwSpavc9q1L61BsDtfZ7wX9FKvkgqnMQBNf1Lh7TS05rsp3bXBANNtNFe
uSbT45/CtrtawEWsxHx01Dvwmm57EiVF9/6bVglOLlMaoKLtecYD+CHfnz0+EnLFklW6BJj8TzMN
Ad9bTOT2Mk/EPTh5IHMjdlsvFDZRo/cfuLUQPZg0V7dAOeJHS5jBVxRXz5PS+lKaADbvBhjQpqPI
LWtw87Yy+YbxNYjH61C+sHVw3VaDiMOudiuIRyHyza7yrD6V3jZ2XQzGNgG1oUmjPzzcOnE5IBbe
fVdUopx+JFTXdQMNqevpCQS8CDVAoa9P2EUDbhU33jOw/j5QqvgXXzZclAfSTbtPoGZdjbA9pS2L
4vYBC3ak4sJICOVGRQE7ta7mAU4xhD2mXnFps1IFjgv8q6QhkLQbgeeSd99Ldi4UqkiaJuBC7Qgi
VLm49ejwbJSiAwfa/7HnvEZXpmaHsL63my3gsKzYLCICOQEm9uxDB356YYfB4Wq27fjMc7WeFTgk
R4Y15kYG9jfmfUQaeKS16M05+ItNJe+O060Gm7jh3ml0pqdVqGFjhScbTgdYSuv/6NzL9BYj1ch6
/p4x2F1r2L/bA/3D2jC79zo/Q47JyETkwIKDtYenPzWFIFECucfyM8+nc44v1kQj6wmcceAJV3H3
uw0eimZJNm4w2I9bp5c8gyhV41RrI9Gs1A2ao/wyuc9gOlHfvvlu8ulWKnhc8f9cNHxh8q4V4rnp
JVFmP8zc3GMjnVoqBVQYVBLKcHTqBrvjzNr3aZPS6nfhBF++duLA6thofMWnyvBIq2xa2TDI7jz9
O1B8swkRyyeq34UBCtPpdLdjfEjZhDhHbYo4KrDausQUz+KAMq2Se+2OjaNfCWZcT4xykzA5rVAb
WNT+78+vgZHnaUS1Ql88ro05ag8bnMNs23gUbKjQEPThuoB/4z/w9sVL2OSvzwJ+aynRf744/cyr
60N6ChYVPd56x/5IhdPxTaPnLc/sY1frg+bSws4M9I7tRjZOCRH6wQMQl8MdzwJuhz1QICtesNNE
LC1+e9wtizD1WFcxA8RRkfYK6IA/wInwuEdk/Kjt39h5Fg3sVqDsD5tV7mpy1zcIEoRWHetsmhRg
bMSzlFyxtiNJA2KmQtKSrnfY/REaUxlexjBqNxNw5IC4Wq3hfpmEIQGt419hOPqft34nl71qvj3h
CM8Zw0u4Cll3KYX4FTkelMmsBvphHEwHaHtZiZgOUgQAq8kZ3M1ZxFuLrvsR/ODkD5HqQTpZAPPc
Yt2fiUU0csfS7pf9woU8fnDmizveSqwjXXhLDXjI5PWTCtyWEU0XL/F36VAdwS3oLZBEv03f+ej6
ig9qjxWHs+JGC+NCnGdKb4DhW7NwrejCWxVsQ1ZVmc71eVzDJGIrHC/jmiC3VSNqlieP/Q9nBF57
N1xzSU6mu1VqYrcdgYziIT+RMjocR2m8I3qKWfcnL01PmTSuaWG1U+qpqRF0frzTIKxz4AcAkzHv
6PCWGmlsawROX0VYhUkzfPsrMioI/DzjTFGy8lRbpf5zo1b37IjRuyIF+gVeZCmq1Np4xkLK4s94
RcMZpZqX6WlwUkNk2ssQLG9axl0M0xr4jvx8bybMRXCsRV27aoy4vTKxuILcW8hKyO4Qev89/IAE
8WhjOK4ixjDsqoMfhZLj7QF9Dj829cp0ENCd7Ry1ykHP78m7chclhoXtNISFMgy0VGy+nfzneegj
COZXuHbFO2joIZRzgRb/eW9DhRovvNGXpF972YHRFlLywpvNXhH5CR9QOHGz3EhlzrcO/xMG9NMT
ASBXGXHQhAGLNJsMy5civEfMdwP/bNyPQxxNj/OHJxxljG5xoOklE6Bi30vEf9x6TJne3gYqAUcf
iqyiK7UzF4LAf7iam4c77ZVMaDJ38w6Gli3YrFF9WpEO8/7YACcMvJtsNIN5sclZzYNyZgHPeXVH
oxSri4TErPhnya2K5OtYNaz/0kpWCGHUQmdiwRNpVnQVZDe9d5ADte+LHVcCSKXiYnA8Qhgjelln
7JxgfGplx7qTq4RLCElqzs2hdBv2DXlMORYvrejjPuKspEUcfz5b3iglRb+TmgSaJkqa0oqY9GzI
bZHRSiyvVZwcTJnUs7tliIExZ59uMZklx95cdjCv+uQSxTiok8DihZ5YWA2T9hKzHFIN23SiTm9O
AYrZM2KCmu9ZoYWZav1KS+SlW6JiPEV7hOFOx4h6guRGEssT24WkVAhA1xxT/5A6jBqI/3KrcIwM
ydTkd0Os1SxnubBxnjfcBLRTEzpU3Q8uJyetl5FEqVUyOVXcssvyLbPzlDXVq9/oyqELaLA70BuM
qkPzI0oBCj8dlA0C+Op8ZMFToH/rhfPzynAc2kpPJpLU2DEr5pEYGnjmp+JnYgRb+3T54CRH9zcL
ozvAQpZRRlMv5ga74CfXSPNuio7YwhST430O/ZHFOeoUUcL5zUqz/NT2Jl06pTkE8XU0NQ1dQZKm
SI4U/Uqv9AQKn80T/GsHl1FVJpRj7u90RFv4uCl9egljzxKlfcxp4f4djGB/nC1/fvxKMORqR5w4
jNwTJ887eKKUQgxV3ctBxQ8X2txpUI8f0ADGZugWZdwNOhuXWoZhRVq503MjaKkUiNQrw79lr501
YWeFbt8NwzjdCFFDYCkJqoSEaCHjCNSFHqKJKkfDs7bVQSwmRS5zfqghdQKb7osofAqphOcRBjJH
NKJN6ZScZjqA0h4BscDvTeUUJLaGcJL95WtAZt9aqMF9KOWFyyIc7Ng+1VTzGKYUuQ6ELg1c119j
loUTAfR9y23nyo41OoEbbmot6WAXX/QDEzz/EmDn9lR34bNl2GD7Ns6IHpo5W8Fm9xy96AGna6fb
ksJRvF76OdcW/41WPfT2o4JckTs5tEVpE+zVUIi73iTVBbweCZic047qV9i1Gedolx8YrbVReUB9
zaeLNIjunJSD4Avao5XHNj5zfP8qQmPKeGP9UdDseKGmo6laShdo7Mm5jItHwJDG7TKQOX0zys2W
RBmdovozzqyhUl0/RbCY8EJagDRchG6g437iVVs1LlZjiaiZrZcJld66Xb9g0wzjHkpEmIVBuzqV
BCtEWdWk7wK015bYA+jZ77Y8WJeFtYTKBaCl3mX4hOKbFurTM00/wdWHTcU5zEiw4MKh9vElBbrc
risf0jC3duNUEp4Qp6pEt9mfeCGgueKEZpcYedkNOzEqP1TY+e5ZirLeYBEibDf81/rPeg/87IZJ
QGYkxvIrh/R08lyRWgH7MQDGiTW5SP4qgrSqI2f3XbKw5t5xfNYrjEQw4IHHlLpq81PiZF8Rakzy
J/qR/IjUnxIWxYSDjrPLsy/XgGle21n2BozO/DNzw/VjcQz6r+SXsLI5FlyjQLHnZkJbp3xKeXMz
PEHjmVkoJF8itXXJfzdHlUQW6qkapCakanLPUKBQB6iNsM7/2eJqDhsOwxWDgFEGRJHIE2wSoE2Y
e9TCza4gbSezxX6IBH1/ifOk1qy9yKT7opOMi+ymT15KHSqJkIq4kv2WLhdj9bh4zYkLqP6EY23b
5NhL+HhgzwHiq762BBlYJbHZkYORJeiutQA2sVwWMiA4vfUMdo1E1eJciycKIfrioGn18mphGsi4
e/j1tAHxruQ2P6Lv2ad1jd5U/C3R5HjDmvja+Mdjj/OHykRzPhg2PtSaKPPpoI1+F1/tRf7YEruj
mK8g+XyMBGlBcs24scejkjMUuEosxzem+PBQRwjRDe+fu+OVKwL143sxF/0mgSr4Oib0XO9Lbisk
j9OSfdmoPUkjZ9G4Dx1pgxedc7s2b41m+Fcekcks39N9hCHh5xboPOJ1VdU3ZEpHaYr3ItjKycz9
aVSmC/nhGVoJEgAkBCyuZz0VaeX9PZqU8t+yXv+vhfGkG8msLDI/yBHjGcP7ZB92Apc1TW5pGXUv
lc9LZRXZ7jsL/LCKzty6pToEojYmnUe1RS9pb8tK2YqM1ebw0BKhl/MLykULVDQyf3aQ3pP7FpkO
Wgj30C0KPJM1JKfA9l9ru0GxpX/TEJoZr3de2GtwTsgkLlg1/8P3fzOTB0W2Uuzz6+jXdppREx4r
tziaWGUAdYQRyoo5mMqm+4Q2KYcGyD/i0IueBe8UFrwcnQmwd192sgNkEY4oMDvFlK7rZKSUvVef
YJ+2FLAJLdj4ZDWeeFxTSSs8xZPVmZAQxiP9QSImzi+VyCV3W7yoL7IGMWvGtwvJvgo6jKXRQGaI
HJzePVBNwNKpdPak9mxVbENSr0Urb8VmMO4iZoFRJM5HFuFBtqA4DlnFfIjOdGkQ+FomICB7AZtv
PhdCZfun7r1ilXWvqghTcoGz3x4acYpLghXh8s+A96sXH8mlWBP6v/MWLE4bdzVa8T15rizUkWcU
vmKze27cwXf8NafNmUnmTxjxXZkLd/BvqZp5EXrtfgTYMr26uk18aehDBENwBBopqChu8vlGtXaD
9/A4SbCo2W/D42t49L1fIOkhCjiSay7wLJunJ35kZvoiUSRr3ynm/aqjkVgFm6Zd8P0CC4QFVpZ0
cqHgRe/22qJYtGybk/ogkx7KgymAk08inLCxT3AQr2Kgdj+4S+vtyO2E6llbbym0TIco1STuG75M
DVCoYhqxT9uVPmShrbchxmtZXOgUQm/4TcpPLtBg0RbaqIQm5O7+PgWjlkHhiQD7Cba6Ru+CouKE
2krJa37X9tkQ7C1yBzUc/erU7bdywTWWbi8rkiq49a83exQAJshZdPwNzV8Efhoz0d64eze8KT7n
/nSHVRLCAjFsEOCzsBVtoLFI7mxlDW2FFRp9YndQUAbIWZLIn5BLGBvTXKR2HW0/YxrbS/b5F6fI
23ZfLcRK9jH948B+A/RDHPfROX5lEEr8X1SMGwziYr4Q+LV7eAWw7muiqf/NDA0MIskvrvbyXJe/
0D1qhZ+xiN90a4ORV/XFdu0riy4PCEqe5zmD0lIEiZ+ptqB/UAcHaLkGZzz4Vc0P3JHeRHhvm9l1
FEzwTEfcQuC6jebadYfSkpyUkV+uC03xuE8izsqJVPHqUR5r1hquqotUXz3U7yqbEpjrjnYtYAVa
wzEcW8hQM2RsHqus9qUJTMBE+q6jT2u+tp9fKVS+62FVFPkzPPO999rVR4Vs0bzA8pr8YLhBRa/a
5uG2hE6b8QT1yH7hGGdkXcE7G2kduhdmJaxi17geTmts8u2kLzJ72IHY0VhWSbfqlydbgyR6f2FW
1Lb9+bKqVHokAO0Dx/yK5HLaQKAN51COPzedkBscNKCCKNDa2h0MCs2Of6OOtK0JEpvvltaL5sgx
LFfaJFuFQ1bwIbW6EtPYrpiFUVAjeyxzdVgde8yOx+5VHcWsviuSUXuUZvMF6823JirXbvjzwotK
lCoCcNlF0NSbZ9I+Jj+BkPXCmQYMTYoBrq0aTl6QfsAiLyxCMsYMb2uLNCYmo7J1ax0CPNunpvrZ
oU/qU/WvRRf+qg6+Gs072xyZ+5lIjAxi4+hylzKwAEPCFOWcaaxCZySwP76uJ7BAkaMmiUNhMBpb
ORfPd6AiCEKZH7hX8hbW6pxd33nmqKBYmykQjcHQojf/xMXMDsV+pYPAVYicPhWjej7O+YKfZfPO
FuT+ty0nmzGhmP27b/IOOqatDzSsIKtk4QsBLIg/0VX8N6tBA+2T0yEOmSJWf+BOid1+TLYAnqbB
WDYVmhmEmABzvpp7udK+IboUdhr2rX5aJwAFGFTeATH0VgMFo8aSo1daCSVv+82v91OC2LQIzDmV
MRVqaOqROs3nlrmgUOGqx0QRNTRcuY4EkF5D8LYVI7nFawqfTYD4z/Zx4q7xqL8XTXvyzKvDIJBZ
N6AL9Ks08+T+B8GDFe9EfT1Va0pmrt0Bl/i3NOgm/6nkSQ11SdaBRXGYAtN81dso3B5KkrhRa7Sk
tf8cmWfwZ+tTRSrUXEFu/vZCb0JHKWcmEVeLmFHXs1HaM3NHNnWIltxJ8bZ309Io/PNElRbkBXX8
vmHJLP7KHykJWkpTDfa9ATZtVFOY6czZw1Iz30S4192O537HRQJgxA/g6CG6BXp+VEYoCbaHBx6d
5Svv9i93vHV8sGHICf6zm38mTed7PBsDMg1lEfjUOkY37GCKAvFVTKJZCZ7EQWyObi2Er8RIsHup
QUpmEOeXParkF1vJyi46WI53foogL1ZKRKYJSupuEjrqhh14U5WQunVblLJvcYsjVZN0ipfWY/qM
WcDZCACCJFZmHsqU+9pk7sSxPE0syeQ0ysj0TlDNDujZc3sip9sTQGPFHAdYtUeoUpiop1YPg7ii
TKjdOvU/XmCk8V5OFlFEMXdCQtjAj07U5bJioQI+MKZfZQkcoJrU0edqzVb0Ulrd3GsPz6exBTXK
q7eP+tGBMf9OinEyZx8t8c12a9sy8ZUX6uOtELxYbM+078wg39hflWuA/vm3OBXJ0mM922Lj2UX8
WSUtY+0cYBXcfuKRaDMlzEofFD9fXQwmhNvhgPevFwGVuiS1EIudUP6m+4on7gIG3ukCMVsoW3Ir
Q+muc8emk77QVLEqPio5+6E+mcBBNbBBA8mQQht6+8tI1L+Sc2I0Ez0pVEAx46KplEe7AcF9+grK
Uc7BSccHJXvVVfPvciySDH0sqqlrttw4WS5S3W04F8PdVBSh/3xvFNIJJV6jvcjDvwRZ6H0001Rt
Vm2VwUF8eTyhvbfbuvtgST6Y4tS7MRxYhLTPMOyRg5eDTM3HLqsMLULUx8O1KOmqvRecJvlxHjei
sjAamAnHMuAej11o4bOpjv0+Q19LolmxxrbCpdYTpJKgOEv/kFgPnikGD8afwfYBB+UPZFaQJzye
EdN4lRUFvj1JLRz9iN88jSjHLe8JZz6nesqA2CDyOSkJtZlGW3ZcM5AJb7d8glcoPHvJyu0TOKAy
5vsCG4u5N3QoQ/4X3EIobn0eRCQhuqVism6+Nm2QgW24KUJ2IHCEBHij1Q+xFySNhgEntN+ubuuL
jDaFFip6N+FKOacJAjFv05KnrolHI4LiSaafVJuWAf5nj7fze7wk03w1nlSJ4T+vOWS4W+d/T3oW
BL+6yuxhCiYr6svQH6lZFyu1akPlIhkPQmoNkVDmfGvENPU6YOfMH+147bJl5sY8yTNPECs1wZVJ
1qsynm+3Mw/w6iLSASpNK31/yxz+zufvHKtZO4hLgZcctd0Ei2OsGICgiMua4LmvpvcHb9dnUR1D
VmiGyA5Hsm0bD1i5YyyPUBkEukrSZXdl0QrmZR2nyd7pipeQ0s7mKb1wHmJOgML5DiFgnkVebS1O
qSpnA4gO8FQouzjoso64+Wcy9XtFZ/ba6iZz+bPRhLmfndUcpg/5kGw6lhjIHpr2dIUC575QdVFZ
EjSnMJjy4Cw2r0FxE++OxN13feoI86RdrG8IfeKLOahVJr3dXogOkQ1XQO90xtDRb6m265uCScsh
y6xlK44loq2Jx031zkhqJRtpRpZKu1v9Fm/HGJ/KIYhEPOwsHCLPB9fDEOlsn+gRTQtjee3+XnY6
ha165FNO+S2Gw7DaAuVLI3T1q3XUT+t57gmLGhTzRUo5YW8mssnWUb6JHsJOfU2QBtUGyclKKyx2
VgqOr2aMNPZ0U+qGBfm7JqX99TNHQ8hXx8BjTszZb4w9szwGJShtx2RYdu11JTvFfUdjf9LeX9pP
GLGlsOAaFpuwAeRox1JUAoDKUZMfy5Wmn4YNPVqyRNPIQLYiQrBnvZIuQ+6Xmthilm7C9BORIsiw
SEtJwdK4dwGj3U3xf7h1vPfY5EgeVMSfdlYsVkfCzm1W22vE8Ufxhwzr028wkOqnIexzmgfes7Gz
n+tCp0AiZhJ3BN4gHprxKglTgpt5x0FIoB83oV8OCc4YuVM1ZCmFdJF7XvNxQwkJtC6F7D8jVsvF
iodTdp2ZcImVrY+0AmqrGd1pd4ONLvRaSBOcsg37dQf3YQIWJRRH0XwiJXZDczp5aH6cVbyvDVeE
zLmj0BVG3s/r46j5dIQXxblos1IsuawPWhJMEkE0GBVE1mRSU7HTuXiR5n1Ue/YXza/VmqcCKCMK
xY4HEWBresMBwvK9OaMrHRvvZYztczFAQIjKEMukFSL9BBUwxINIID4ssv99Cg6qmiGxLUnM1eF4
qmLyVAdyUTvnZ5PqWekWPrArM7mspRk2LdZzCS+Y8XLxC5e9GkMAual3LP96tvm6979Jb3rq2l4i
cjvRWzOgjcDHVxlctzhGJAh8zqHTaAntKUGgGjV1S1Q8Mfz+zSzPr8vLytmKWb3FWOQeHe7aeDJF
YLJXc3sKTxgzHh35hwCRz5pVXBdMitdwTsiL3K04CzJBBpNYeFJXt76hW1z2s35p1IvcnXOuVX98
Z0pfwbdpnP/211wyvEupbWs3D2/c7J2y5mriO8Qw/bJRJobHFOpuzHfDys+oaqJ2DtmI7TeaPDan
8JYb6LZuykeRDTyRER3okL1Uvh+uJkTyIhFyD2+7Z31a5LfJ+z8XgSMHeWNNgihNC9723UTulRb6
17zYLS5Nm/ZZvqb/LeYTmTLszHP4U3L/Do0Jxd7rCzISgO0IsNFmTc5OO353GLT6+Rgop1Y251O6
Lz1xhkkA1OTGRPs0QHie9vyTufuK7MT9/kLoFRTjrZWFQ7LlmriG7mMywvfSyhe2NR7UkH3ITOI9
Ibm6m1p2FVxSqZ4+qELnCrlZ/L+aIvvri38Ib4ATqYn2aPy1AyYp+v0aJx7x1NtzUrNpYusSEB/Y
SfAQ9dknqFbe32rI/CiPh8lR3Vku+u/9RpYvCic71k0GrrV/he0BwHpDkfGJSz27PfX3g1s03nc7
zH2Obstmlq+CBblchPwlAdI4VMf0LL9N2JEm9T1SZcg8SCDatJRALHbTHjyH/CnYZohsjZxUcqKa
6oheggyQVo7Nt/Qr8Frtl5/M4hm+n479sL8v4dlpTyE37Z3cKQnxqHmBpIXLGcVSruin1EVmiVmJ
vB5iNlHBqkpthQiQ6AOr3gALQQNihyHwdFh+d4OJo1HYHN2TOrFxGcf8ewSZjrb5DiqBtWa0nfUP
DBYAzoiM92b+CLFVgNt1lR0ai4vG8NhUQa7PGmyWdn25uKYp+6Eyy/OViMly6l8RD4efYaQh4c2P
4T1ufb4C3Wb6s+Cm3Rt2oPZi+nDFURZqYvYthgt+/xgtllnwf5Po4mEMPfDtQAm0MlDLgjvn1jqU
gRYF7QNqJKWVHp1H/INNjVo6DT5qrzhI56UUQgqZns3nrSvQPyxdDROi0STaLdeOdzEPDcCq+sfa
H/+Bas0TZzb0rak797B1PjSfMuW78BmBCkdp7DjTx9VVszaWd4gk4++EgAQ9J286QvjP9Og9gr/f
RqzztFCKJUfmjb30c/0Hg4ACfhe0L/4TUeeWmLUch2a4aP1iyzDJD64NCcvLj5Oyww4ZrPpev9iZ
zaJtAjdYGLewnGM6vvHqX8zWFwlWLUajsJnpa4TVfWUnuUNt+tunGc6caHOXefdcPbYgGRu4IAiy
XPAubSM6810bPKipz3eM8SqTO5CLXtPbj/T3Ov+3i+7AjL0pCk8NVjnqFcbwJ37D6kEDjeiyzzqz
vhP4J2jutvFSjaPFCmpwtnaCabHucArqtI/zMOfyuGQborJ87MSsv6LKrV4rLBej7k28iGe444nK
2JR1R+ZLqb8NoLfkwpRr6E8OOBgrruQN0Xp4IfoBrSBZZ/y8DtNkNxd0NQGUNexQ8MEMQC/qazER
lpq+GzVVqGAUereW1wjvIXDQjIIhrGi+e4DQYxIInU1z4XCakTDrUyMfx5OhKAFW5XuygCIXZe/m
MnztcSm1WT422vuTUWoOPmyzX78QTGa2CpF43aYRUvINxw31wTSlhlz6WWecXsuMZaOkhiZP0dZZ
qJV3cCu60rNX41ZmuqEQBku1F1NLPTldi835AG5ORpxCwK19RyzpyYFBfBU6FuDHybUdxqEuq1DS
dGHD1SP9KQ02dtYPho5HBtl6LdSSSNDPJhOPrqXyq7YXwwOQOJQY/EPwvQlZXMI8GZRbVbvWbyL+
gb7PMow3nFur7vY2khIcPxlp3S4mmDEB6oq4847N2UkLvMtn8ZlMIa1gjIr2A3QcZZNcabFTNnMt
lhdnObacHKvT/HoS8a+pEAzjltLj00LrjXapFL+7wXBZYITaIWeSyqnTnYjw4VML90/xz1KHQl39
AmwpGGi8fysiwri4jfCpkiaXvpxoAbLA1ON3n9h8RkFCOyxZxpYqGKq0s3vaBCEQtWld0dUZeVeR
vQWzfCdjKGWvmlx8qvHeKYLvV8kA5S3VPyPOhFJoJ/BYvQg/IGOf4ZHQuoCPZdauD+5kU7CGyzHd
FLxIcGpW4YUo83r/zmwmQWuo1FeWGkvsCk3cxn1fpYs2a2diWHYPK01CMqHUrwj+/+XEa3/h5Kmq
Zx9TPkIN7GIkc6TF2RO552dX69S2ePq0fM445qyAKoWVkaXxMfpWnWwS/jtcC3hdeYy2nkNdeTER
q76v49+RwvvgQdwiJD/wnvNxYqKxtS9FwkX2e/x+WXyXbYhWLmGH/jCo2pPRiACu+4YZ6a/jIc61
E/gTND8TlP9ar/MSugpHdgzh0bOswoMHa63ZpPBotj0/CQU6ExceiBnnL5YheUEyQhWHgJg7rvtg
pVjTO0wzjDQA67i9lOzLFRAqg8UdZIxOqiKK1FYVf+NuWOxMPnX1Kbm4vAyY7KsiXs7d+/DQBjUy
D4mlBU1z+L4FBsPezsk49yr587Ql4fggpLyXbeeDVOei7gYkr6IGE+bhAvGRM3bbMsSCmBAeUko4
S4MjIqz/+62dIqzNsH+DfN2ZhyQmekQN1wF9TxJsm9MmMJtHYNXoTNqzuSKybL6EPIMb5VyGRTG+
oeSrtPxl5hFjFlnfVFa6uMEvBdJ1W8CGAFfr61ZUDQ2eukjOaZPSyheXGriEJSuJ+9qr/fgi4kED
4ZOqnSWJwgOZ3BuJLX2v5yYrdxqGhwbOZbFMeN1BPifIicN6qco5ZLY8CUW/IBQpB4yZMd7Bt6hK
iA4RJF96N6g0m3wNyhTZgcwmn2le5xexlzOXVLehxwjmYaoCuSt0+VtUBgB95rbMuR2ESLW9NUhT
0oImeIVoj5KU7F+0HP349VemuMauOs/IiH4FzQJu1r4V0U0C8B0CKk+vhyX3BDQv7L2jYOf1dF2u
iu8garoRrrvI1Fn6T1LV05aIZAyEIo4/DmYgWGo3QSXB+As6I7M1P9SFe3kYr7k7fdTKo3+228FV
giRwcnHAKpEl+tBiVB3UepPF9d//wvZ1bMAPJPEO2nx7GGcry3QjaxKJCo31sLbPY1pan+H8UQn2
zeCufi4++HBIsMKbVKbRAN2/6pSqUtRNky59fOH+DzQKfv9nGoSVg7AnWH45PfHEjctW0bgFu1pU
vBGpHMbVvxkc+025NKGlN+lemr/2aQ7elWKJf1rgYsx4vWVilNakUs/IM1I6Nm4tctTFDCKW5AuC
RuH2N3Hdhg2SlJ6J23s1COoT4gNVjLaYP3PDwrZuyUiDo6O2EzPSsP7mlT7uHsixtKCUyoHQZWHh
9b67OwhaPKGwyiiIi7sZtyZTkBRkyIEQ4D58fZjxdcmHTcOE1sMaS0eQdaaC4o4vNPLS8OFvx9zK
bU9WPDlKN9gIefKJsAt3yiTh6+j5yyDBtRkpSkuGKlZQgTe2XAwXpfvJblsA1RC9HRNCFc29Fiz4
kjurWsXz6gYQv6UJem8hR0lC60mSvTd1VQ/SlaeJWowU0OBsbJGqzrwZQG2s9qLW6JOwtWCh+Lz1
e08gs3GoTMASzTOZGE0MQkdF0G7mdRcLd9x3g4n51meQOZO42wdhhrJrzVmKA3qLKL1MTzkrG1tn
2LiqlbyRAaWngIRSkEqluq2basgkGpJCMwncKBg0l8gMDCReASZAYtRaS9okvbXirZIGV00BHQ5q
ccY3fgOWw1UnSJlrGb2bRl1wEByuK5mD7ILMwjaVJjmHJHyTe4308L5WdHDXbMcAB5hsRT+iSy/v
8dRNsCPx0ON8tL7A/J8e30oyV78yyaTZEz1F0cvIazXZwTGB7p6j9PQ4Vy0sQkScSjB2NxZpdIGO
i8KKpEMYxLI/q+tKiEK1HrCUI9zG//fLsa7xaphQQiApU1/fbwhgkmy/zcorluWNUKLuI1t2dyXg
rZyt0uL7SCWiuDteA6uiI619Fsxf5tDy77PKkRwFMfAxU+2G1rMV7NSuyvbxMSyBNIjU30jvugED
o9O2+u+yB+DdfNigB2kh1WvLJvG0jNZtENZLYnAqXEFBRA0dlMJ99jg91i1rLdfhV8GzBP6P99GN
IZpdcVK4gzdnpJGOsfXJvc92VyFtXuZg3MwkK/PRMEtir5+Co6zRCp2V4HOyPVZXr3thLOr9svRc
WmVrzSbE1MvaJ8ngCuBDnquaWpMcnKiAd8Z/2hZd8+4GP+gZq8NYmMplL9M4sPXft3G600k+xElX
TT7KWdvcyzoCcnLBB8RmuA9FNel/Fo1b8kXfia8nQGVfN3TcZrxaZF62Dd5eyGtMNzqmpcJzYT0M
rwwKKDpRMBZTklD0PkFLdyJfZZ1RfKj/9COHqZKKjjdpOrYB4LuFeA9L6CyNGFb7Qoe/quzm7MIY
jgCBOSKeBs/oCQNuQxuHyEKjmLweOyw/gEXGwOh/QitJq/rlqyk4+QXfu2UgAoqP0fx609I44R+q
qp2sUrF2TWQIxhbS+4HdF5Wd5dsu25OkFjMBoVJWM/622rPGbfkv3HF7cg6XxoDMFrrNUfNAs9N7
3QSg+flned6tocWXnoXxSYFWDczc0cbvf7HnQguVh001kQ9FyJtSOHf1R/sfbGrTpThF+rNxkkSV
XcGzDugQulFJUZw1KDnaN63BH0gNJaEdqjTViW/0e3aYkZvvpZ15X2n28H5T3xuqqdyimPikX6Iz
iNFVaomz/NviqJZ5NwVjePB3bLaj2ngDOWXZxDg1dYS+JqnkhVOManFUURbR6bbTAvCC4PXhBesB
2fGdeHABtc4M/EurRk6Gx8Uv0JWN6NqWTEnvWaD2E96XxRG+BuqmIaYSLTq098fkVM4CNYtlrTT0
g7SE56/SEdXoagZqDf2wxIQP8Hw8LYAERL4hc3sWhBug9aQ9dHWEIt96azDA5yeyXc6PJdhIwSE6
TmyGOBH8HhPHrLlnKgFA+M5VHFeIJHMWDhh7jfyqhBbmqauqZF7SP4rf0Bw+2wivP0vSrnG3etw9
hWUNv4JRKUtTOrLH/H3im5eK0UmO2TKjg3oax+WohvSbNc7MARvchh8BGfAIPiR7NEfJoLV3cGbU
fOhMKVOwrYZc7GSHAX1FNKEzG1e6kj7tOmv8eklzC+riiS6s4IFa0G0UkH0hBLg6ShnGvxLozjqd
Mv+nq34Txz7t7RXAJO9DUAnkNMPcNNqtLPE3w9WqwHKeJaaUHBiRQ5D1QUSFy7D/k30fpeIqgK68
4rTtF9azRpeSbLvNhjU8FY5IvzMr5sQskGl9CzHBiVbZimvdKFEtA2giwnaqUu8twQxgSEyl/2eh
pfTY9NF1nZqfaPzT1/T0LDBrnK+wJA89MpGoxoUwzMPdbBMp2WxxuGOJrOtCR4nhRxiqybzIWvkB
CeNzvn3AAdKdYrEKnUlazIU+NKhe2xtCb9V4an4VDycN1oGQc9AH0aUFMyMOu3QStoWG0ZOx7VHc
iRAQc87DT1/MMjPnFQ3IGUaafhKQk46mPBHgU1D0t1x2OFN1urGJVyR+W3ef0VnCqDr++95VDhU1
9qWL35aFf5BWNeKLtcfUornciJA+0GBed8Zw8FSHi+3ZT09CScq57qEiT6rCabYOmLiLa4jindCM
3Ped0ytRSNV/+hFLifvfSwuBOZsSWw8C66xoK/piwBH3nZHIVs6xds7/5hixOU7xtmb+MLBILIVd
JXMMGEFqehP5TSvA2RvwgXRvoZkHBzIQsdDA6CaTnZjkBc4g2wnezWRtFZ2o6aqLf81xqSWDKUVt
+8tOzCf92k6+Q+n0Ioye6Jc1vsjpssEppFke1dZZzpopx5TWLe/hEL+P8cEOX3n1CZpFblGJ1t45
cvu+z/HFK9wK7lSnhJJMQDzG54k3S8Zwfzn6+k12DTE68zNOqAldAVZNTauslnrZ2R3v6pKixjWO
PAKqy2p/RHBqKpR2iK37JU+538PpJ9iwNPrUoUEIwrNd1z3vrRPtXSBtzeULZbrUcSYN4M+RNNev
FG5gMG3LoX/EBlZ3P7GdCFy/jwyagKDqu30pOOnj5LOjhZKlPShdZYpOPytVxUmlyrC2SqpyFcrm
vJyaG1eS1AnEY+IxYqidmcSSZEUzCx/L5ncjCKzyfugdLweWNFvs28iHQh4x1WUAfEGWLblWXocB
unJhKltQZg9aEYalB5LBt8uTdbACdyt7sIrE+Bhkgg2sveXcK0zaIMinUOYC6CIV7fzX3+yRexK/
XOcI5fFe7fikT4ZbczUx4TCz2jAuzlNOMaCyrDdp+4RmbhhNKcUvObkkiKG/2WB6MvHyhk6VgLnf
DN66yVlW/XeGTMkzF5NfJE1gafr8816b4l2sQSih6QXqeiKsTwKMyf96/972v4pFY+4E5A4jdztZ
7c9Owm7vX8sKkuoE/YQyPfpuHOCnzSmJIt1kUYiaJPxFIXcqtshVOxW18dWecmeZ1XicAeN4YpEg
Z9WJXj09mqvswtB5dcsjYmmhWUTLqegZuUQUllg78SzKNBiC9XrDjzWZz0PYKaByC2ZP+I985j59
ycSKLWORClqwv5lFj2fnUD18Q7UHYHTFIewxyFQxcd7nrNAqltCtWvFJOqW1x4mH9k6bhV9zao18
n1Qg5SD+DFauNu8tbhYAm+YgSAUgxz1jj/n1wH5/SVvP2oVcN2B43mF7cS2NWdE8K9+VBL8F07fO
+XfDyJENXa9c1DarhZBK/HokUSOnsd5ZPjxeSZGhuxOpR6zjhETKvBGD63jJoGNAnEZtbs++7ITT
W7Pu9ptWy3TS7UHBkxks8djJlSBCA0hNXCIxBwmJuzolW26yCsRRvAjghwqGgLQPBbBwrg1QXU/E
BlrZ9+Su7VZIkClpTkOIxrb/mGW3SWGu0O9qz7QurAcpR5uTWWt2oTaHkLY41S72Y/O199NuqwQa
5CrCqVWEFsiI0brZ9D1D7xS7gL7xmfPygJHV/g4G7k7yPvBRY1OXPb1nRIX5c7l2Xcl2mnstI1O1
8gPuB9S5kI1Vr3dvNiYnrfiBYk0nItw6IE3mpGHjHUA/4caqdJoP7RsuDru3OKTWan36n/USm4R5
kzKT1nZ8AWmmMZ99StpJDWb+KNyn2m3zb3itIKP5aAJAbaaXvbG7dE4R+NRhJBtQfj23aUTKDwed
BytTjbTRGjBBS1/GLTK2m7TzoKMQi2/602J3KRB6YW3PeI+Qi557rbpKMi4kbdXrTYcVnoNGK3Fq
FnGy7bJSNaHd710XqlLWXnvGLZB0am7eqNBX95bd47WT6dbKfUgZle/GlSWjrXWKr0mT9E+70ori
uM2zN9FHjEW6OSxj8SbXo/jFwQGH057TuWwC4TZ5bv0Ezqfy+9l4Be03tgQvZKMdyW34D7z6et9d
aRI+B6FDGDkBji0x8vy9vTi4S/K+cVQhbK2g0K8W6jSA8QWgXpqEooIBQj6d8CMt/8lrDNAw2oXT
B/kKnmrnK0kQ0c1nP1NJdi1ia6eK2CysbJflbXMr9jEaNSc/obqGO1SnCj6rURtr7wfIwEkQ/ldv
Z6qprlJ3P+iRCncj85sTFic0rCeiYPohgfvEMGTmcgtEM7HyhdOHOzI77ikIeg/2M1W1EKjxgxjX
1NniJkA9Vf2zvm+iZpBCX6AyuFF4CSUGofOzgCyLNUE3H/pvGCYP4bCoV9CAc3nAUCjF9ti5NM0y
bPPjAF7sTBFDBTRlkn4Eg1vWJ/s8Rr682Nr1in1q4fjc5vKU9WxH/1FJRyzJGyZy71awYPQcwuui
vkNZ6IVQjOXVP6hGIVjffn4FC7udd7MxRJArQp6DEnpUNU8CPYdX3kjHXWXfu3HXEW27di2Vx4CY
Jm/sg4DOJ3afnVrgGGbw5oqZ9+CQfLqxmRn1pnsBaKbHmLMAq3xaJwcHnWzFwJo1sRGih7C7Js+t
TjLnAjxkdIRBzR6pGzvYut1+J1VFWZeq2c+f8JNnaumuqcS963IIkItYj6/Zce+XS8AFP2m7uCPq
GEb17r/IiqUX/fldk8bkD0G3FmHwNCWB+c080DYjG0dHEaf+1/0f1tzXQpZjj92vRvGWkb+L+6T0
+HHndIEtWu9asGUld+W8E4t38C2M/oRAbi8kJOHZJlWeYREBHCAJBKFvwrIUcs/AauaF+wzNfUPN
+eTPhbVZnT0v7Ms9vrPuvVpAoo4zEsfl9QK/cGjCP2gnwqZbQ9lqQRwPtW0m1N9vy9bYGQT0MDSi
vaB/9KA6+mYTvjFrtz5noZZOsBjNA+SUIAm7QW3sDT47au2mA3dRAONLO3uqUcL12lM/dFNTbNke
FvPtNsGqTv5PuzDEa+wl5wDgAVEE6GTtreu9DBAJIVByRQoXpnlS5jacF3vE1VbrzVYn5rrZ/+dZ
UpSPEaH6CqcNKljNT0pbq717e+bmWuL0ayAhTaUm9+0ecEqgBrMGTnhOzqtpwZKJoO+0UqviPEtB
pguI5+fv4EWE/m7Uuna0b2DqFxApV6o7X3DrkcXPIb+S/N+NTzR7X4mq+ZOL6cSiirhw6jbnW2Mz
7a2GSlD0Ah34VQ0urPCkw12J/B5x/xd5Rqyt8giIMUATn2L6MMAKXqI56vXEKJKFCYCNqM7IpNVj
ULLkgsyIaqB83Fwi7SMaIk7xy5y4r3BYbaqHIh0s2eouZTED2uEai9gDcfOxbwX8aIhtYcxts/2V
9o0mXwsbSq3DOXMYAQNNNABmv5dX2gkkUhvxIZcugsKRqcC2tCDOEX1QzQS3jCDkqbZIQK5nNHt3
uDsc5ugstcdhl1gYzzKU8nHlGfVt7/DnCJoG8H9RBOKCkDsPYf/3p938ft0YLiiYnLrrUvD0Uam2
RcE4CW+MUTEG6puDELA0XYLXazSwm35E3U/vevcmgXaNtzB9yeiPjoG2VNjM53Bt0Bjp9Xtt5Xkz
O/qumGb2AYm74fXRCEiyCuOf1WmM0DXzIDQgQLQUBwHEf+k7Q3qtr0ibjb0QewB2Ubc/TPHte0xJ
GtbLGNXtdNl/PiPrd5dhF7MZDVe0GRQG6kQH5woMs/4Usp+yIuLvlA88CglI1AYTNTEQl2qzgOMg
EVHmUk0CGdeUUHBIijY4UWYVBXB+gT16XqllXVndyrZpghBvyp2I4VEyn2mzn9p56W0JPTkZw9xf
gMg1tZiVbgYfgeTZCLBNGcIte8aHHxoCGgck5vOVo3hdabHGkCDI+k3voafcV/tBHERyTC6/jAGw
GkrN7vR01JLzZ0RRik0UcdrvAhs8inMqMrhVeGKJo0+Hw3H94zeVOw3f6ve1+ejJfs82HaQgPb1S
xyAgbUhnCSAMKVo9ix2byRWMmdrEuvZ+vHL9O7gsEUg8WjdwhgjAYGWbrKuK6zc+a0szT2MA63iO
KiI/fC64MBoY/epyQ5CJlHfPMsoMg8ylIxdhZdra6c+LxXYYkrwFEo6VpZEH/Kb10fQIPasHkHYV
ryUqc96KJRn4ifwXWs/iIafdGQh3C5riZx9AOQ/XW7S8nV5K9WkEnaUIKn90E4YrKzq3maUPAAy4
OmqrB2a8nGIOsjp15HDDCSDp7kts7JRRlXzrWf7FtXrm2mnYMRRiMmMnDhCpLxrmu0LgZHdbnf4O
UB0bhm6PD30EMxxhl19soWxFo+FaC5YMO33pGEaEjE6sZf7+94BhunB8h1FlEOFdiKtdHNwhO8MS
QWxMLmIT79+nxBvPZrZfLQl1ql6yhpC7Cu3joZFABsbYAopQ7oheiHuOc6qKWrNT/xyS+8DC6y5k
QPoeQCNf7TJuUCi0t3rCU2PggvEamwi6UoXaIeu9Wttmlau8YyO2Y/J97i5IvNLtNmYjcIbDOcQR
vJn5Kf6Q3K7WQWhBFMopttY939WCBmTkhGJhOfBhl3M0RD9iDmrqpa/AJNu/dL9cTA4o3/KAApaL
IjvgOW06RNffeymEXmHULB/Ps9NAagH/KRP394u6nTAZJcxyK8yIUhCEbeQigoPN/Xkwjaodj7Rn
RhUtsk3Gg17bQihqwdZYD4VnUo+7HdORYI8TK7c+yNWrJ+33QMX9dCHYEd1bjfw1OPEvx2xnvr1g
Zp38sxOukfTBw0pnwVg0DoNV3xpX2umAjApMw93X/loVd3tBXVz7ECRBMWFKtu86OkQCYONz/bcQ
kxkIGJ196CxKhBJv8B0G7iN85lQs53yoT7+i2PhShq0QreTxyxnSx/sdFgKQkwa5PIZ/es/eMVJG
96uC1XPC25M0IJptAU/y0rofPsI5BLILO1hPH3Nx7maaLBmVdz09bG7HIk1qJAuPPo9QSZ9ImZ7Y
pXCZkGEZXbjNcTsXzvbZ4os80Nh+gKYKBgepeUJYD5tXDyQjfAc1T4z6k4shrSDw5wPoRTvd36zO
aJk2F6ww+L0fFgnsSrtsst4ePML8x2jlQS+RrzlXclDdNMv2s7FeIv7xCAEe2P6/qPp7dQ8xX6gy
tTGYpbVAIjzXg1AI5D8X5xbbhvNhSTOyNdHWU3BwGigrzwITcUnTuvPa0lbuXiFeNVUsnaVoJiFJ
xumV0OOvr24Xj5w0DPrF3x/vt12NqCJjcj6Gwip3rWPgxc2Zp2wXaPiGL4cX0rj4fcdHtmp8oA97
mkSheRQkvXcZj3TxUNs0iu7SIdvPVU1Ip6MAgyiWTYBiqJTS9PMxgU0UPjD/leEbHXYAFfFQYxsJ
aGr/jhjT11N7f0kUalSS/z+n4nRrrC39AYVjirWLkJUIfLqUgAKirywq39vosVNNGsAZeM4qY37u
w57pLFiRr8Oji2TfupCmnlt1FHUAKak+PGMFrMHm4UzlJdC30YbGEP9+NFGb5TFipmMTwYx0syXF
6twBZMvi7idv6PQ/3gwCVJco5K05UwHxAj9X0sDBtXbEX2Su44ulZ9jpAa/9g3LIId8TbLs+6s8c
r5uvm9lZq0dE6tczMwqtTCAMfORsIiO4gWEBzipbxM2KrtmX/wR9Iov+YDaw7KBcOMqVAAfeR1LL
f2Oy8L1N2SxzeN3f/sXDbH5tb0+LfHqaA/xtjvq57zH5s1DAk5KcOFKcTIOwjM+GeaGKUClVKMNk
cOygRM2rQeVHwXayPvTYARBQEPMfP75mmAM7H9s1lqgrVAsUIxfPgoi9lAirKN+0ktwxfznNzAe+
EDCg7vxgsl1q/xYTgT3I+lkNO+eaWFUubWrN8zJEupTAgA3HCmGx85jmbrjUULVcfa77LbN902Ij
hEIwgysVC5PcVszo0CsNiKOSMwytpbfmARJvVcOhwpV9D0uoGneG+ttNI9wg2+r+HVI5hDpAjqyT
+1Dn3l99LVlVbXy039ajbdDjifs96e9qkugpkJBoynkWr6oApwl2ZhkMDSmCfCFj2uxshd/Eyq6u
dBbsKaBa/84fjCnRlLVv84ZBk9YtFVSNOrM0EFU70z1hwi/73uI4JMFD/8S6PFpqrPTI4vcydWpr
UH9+HTI9uJlWjvr/U2CFPqpeifyNYp/4+divXLJWEG/+IYhJI1fa8tEKY1ibo696liISCvV3Gyjj
2RL14M8CV4W9ixefC55Fa7gwyu+BaghSydLMu/xJHzOHIOLyK55cNP8X11CGfSlwowTDvV+YxmBU
FWWy9n7AXoji5t1Kju6IRc3sviqcusNkPGOB1MtlbzZG2FOG8TEVinId+KY+/E9MIJR97EniUUcL
6uN+fa1XkW06SKNYQ1YSoh9xP1jQYgOzkNgu4HuMpQft/fnW3Y6Ce6rbBHu3KLk2VjoIJbvuCWRK
V0cnk9C4iM8TvR6H0Wv7s2K59rVrdG3w2IKt5BAIP+4L7NmjlkpNrnI3J2hEMVX582S5KcwJETj4
LPdPArjr0hhKHNnyYYK7KLtzWAWSuv6TI44k8LZzxxjxc+36lNUMepGmog9l1SJ+sciertwIcLm+
MZ2Yz+d0Ow+yAz5ooNXAM5ElPr1J6CHTGo6H6DUaHEqgyuOBed1htihNI1yVzrZwx5vg5FEj2iSV
e0ST7svTbjIdmmqEKZ92LRHlF+EjKTRIy/l4eR05+maMhfwcBS918vSbJ/4+GAxtO3RG7KMMHNYh
DeBGXw6E5LFe+nRIbF8Euf76hRWA4iWEyB8ynJn8+zfM0njQpzASpmvOPc7/Z1Xrh6LrW+Z7d2Qt
DZnTsPhbrPBK+Kk1u1DrgzbJs+jPM0y+dfQpCbSM78JzvC9UDKwL/WaS4Gm6eXGGySIz2FH/RfJV
KHKVs8DZF5P1AdD4QGCmVlC70JmsOgeyYSB/ALJRfiIxASfHfH89hcMx6vmKOt4MjvpTK0oVe6Zl
hulk0GMvG4rQLfLdsE+CeSOBYxC/FZGQnqUktfUcxqjBq6xYsDajljWsIb09+eFPmv1b0RKVT8Lz
7todOYS/fUoP3+h+r0OYAdsBm1URSYovdB3itc5Z/5xWHv3rnCrSd2Y+iR2YcfLCvUrP5lvAEpt7
HvF3mvUqZLSO3LzBU7+yutVGgWEozhnrDq/3CXxZsHHsLalEZVTUt4wkCVi4/xaSrM0irCzORQ09
ifhMcfi4SnOwDfI3swfgMVrhT+MojrDv9spCrM8fWKCA6A2KLw44miADd1KdGspp1VQpuq4Ifszw
s76gRO2kH8v+VPHGc974GH0HcpwKXTcNXGCW1aKsDtVa+3PWxU7lexY8k6PlHEH4RxD1AaFfoQPE
dsRUasdVS3LssTKPYq/SturEwzxjbhTuDf2FocWfR0EVgVpL0Iv/Qx/fxPRwDgxqbMtwqdUhgywC
uvtYqV3GDhq8iutxqpV4L2QqnAuiUBHuXETlXEHnykI2/oQryfOmcRN87ZJeOFFLXsxFM22dNS+Y
iRcTSKyEVMGYtJbbJhNlZ0KddOZyG1GPCKZvc86d4zFxQaUWoGMoPqXdpE8gYIBBqWQ8yT91b1/i
1YHilidd/1E/ggN9TOubDKNnVvG4w5tWOXb7Fww0FOAYTDb4T1o5Jh86HpgaBLXX6lzbt71iE89T
0vSziblJrNqLOQHrk/KM1XKdXx6XDCYRXVmlXZnO7Uvhmn2QMVqFss7b3pnKzyyMlVpAyEXKT9t1
W5roTONc9PaSRnMkrdE7+QgO0c0KSMyPBUiDwZbI5Eqz3NpKG9zVKDLFW22x1D810nwwKCihNJ5G
KIf6rWTJ4ZzOmZJ6gzl+TqW3HY7QtFZ60Jlen4+g2oGKcM1yKWKBZwEo/uT6DElpWaYbJ1AG5a1c
mvhIkhlkptIoDZ8wxVwczJxPNrZT8iGPXXymWyUUQ5X+q2qgrb2v4tvJ/FRbC+VN33p7rulML3IS
0rdtlZMW3eS7SOSUprrKUM0AhzUeQIhSOIj/mzPmb3Vdd8mS263D3dpPNFjffx1EiHnvXfThjJUT
Pxth+qXNYPjc6eni0ROG2m4FKHUW2WD5pEG9eydpRo6MJbQIQ+u4X7VapFkmQgLIrsvrCbEuAgAX
fDDnOQ16ZtQdbDFjDHtTjWghXnCp96QJxk13RSAA2t/M1CBIu128ogf9Un9Kt5pTQtWlbv0Rz3NF
lVXPQhbNByJ1GtV1mANIKiX7pBdFBekS1p228WUQi1XlAmhEB3WlPYsDBHFY5BUI6pCKDRqpoV5z
jPJjukV5AYiwj1Kj9PduZfNxON/VLyS0nCZvkv0t/7cyCUWKjZVelkUFuPHzKb8hojtL8vdOWgAs
PJ2ZY0WTSomRy6PYXLFST1XPmw47DamedoI0afOm7TwLyd7lnAo8Oaqpks6Y0xejPoz2PrAfXrma
V9fnIhCpB3bIun2EuSdqy3DPZs1C0dN3Ee+YrOVWyIny7csZNHN1S1VoxYIiTIqNzRYSp0x1Flf9
XzbPJd61/ah/9ohxhDecUsajQERgefejmt8CbE6QLw69rwbcI0qH+3IblwlSX0TqIjB0lc9OLxQ2
IDZPvAgK3dmSkxDLnVGi3iwe+Sn2k3F+bxeTP+pLz/7cy3YUDCneeikg115KrIFrpxla7KoJRPDw
+XqXEa6zO+A27c0lrWRMwTL10J/LASKq4/AuXvq5aTlgf2uWbOpOfdRooU4HJPm3OGAKRdx6QTz+
KgkFLxq49/zS7utb2BMkauWbh92f/E92zMyx90vEQFPVa7gEEUiFlcPuS3cznGJp/QjHTE7oDrUS
nXk3O/r3h8jdk5tV043tXyta5uFU3VYZzKibQrZJNWoG+hzZD032MI6jKuRDkuONXIkztHxG6vWP
Lw9zN557zqGcLLpmLFpkGQ37GFwbzKsQ0lf/+oFxFaWFnUmxSpaEtKdnyPw9v2ywPPl1zjk6Lfxz
tCAJwLYH0oIdTAVb4jfFvOc0uwDTE3mBPoAhpXWzifHrds2YbQt6zyv18NXeLyf5L6hz9BvClNM6
6Zzz4xbRAAP9KY/3sdwOVdWVVJBfj3XC6l58AoPV8+hgSjwkVd9Q+cpHqe8lYX9zj6SrNGl+QAMx
hRY5Zs5fAhCjs3dOfnLQcSr/LU1wquKXe9xp9i8g7Kkoamok0KeS3Y914Kwy3RpT8XRNiIhJOrD7
tx1v23yFoidhu00vXQIkm6HKT8WTFtVD1ZrZxwKq9mp34tJor+z0acmykH+MheRemd6kMb2xGILG
jRza9YjrDJAjSXXmiaaJCSchqXN75wHWfAqGuFH+lNHGZbtEJS/0efvhzNYS2JoBewnKeVFbwqB0
V/KTBTbpaJUjSRk4uCz+zsiwcCUHxLXu68ruaNqF1k6X0PCP8Ran7DflBnHiCZrR0tNa4VDdHt6v
k+8W0xLImSc3Yxkz1Aym9sV1Cf6KoB561fQvkdeA/pLV0xF0S3uF2I4GYMWr6IWGGEM3zO7soUGd
hWX5Cam1wknDVJRogqCdKWip5OdYhW7oi5LZ9OfB8Y1rdWCTm7rsfCDzIXN1EJUjb2eGdx8zQKGD
1FC1E6Ja4zpqFMsg6JNq40/2J8+FG4hOQmdb/bT66g3zmUR1H0DqZelmAZYPSjkDI733v0bk57Wm
IP4/tYpAIn7qzfNfsANFi89Mu/SRS3hnGYvFpFnLE9cQMYZH714WS9cCcU0ELeWGb/xAgyA9S7IH
menj/UD/m/0l2GorUaFxRUyMoqy82tT5BSFzqU889OAcwmebqC1oIUwIUmO+e/8OYap2RMG2Vs+i
HZDW4sFE5NBeNRb9hy1H244K2feRxzjTxn/3ApYsP3+sHUNtAQhXt8ldmd5bhuhr280WEMQXZ0G5
tfb3hKkGWHPIkmquri+elYtgbFrFiiDTL8kWfaf0htN/5AQzt7/CqtDmRotw0xNE53ayCJLqMeoW
QFHotJYbZjNYkp7QcORliFej0eI3/otQfuwakB4l8D24YWJnA4XvdPo3aRpceBsVgcjZCxYsqP4X
PHXeVR1Oim4YtCD5LSjsfebjdazTTRA2goQwMKjN1lakP4ZKOaE6TnJTDZ8Hr7MWUBcWcQ99i2Dh
QIEOdvdVlar4ODK5Tm5d8Y6osyQfcQt/ZRue8AJ8Fm0Q2Gx+0AZBij7XiZTMkmaDSBHJll2mLksM
gy6Cx4sYYrC7yQbujhyV/Jc7Y8rtNT8bfKNYrfN1n5ib5sx1X+dZX9Q9NaBhgj9fDWg34dER3gro
8ntP9rba/pzCvTOO59w0Wu2LutuZ6KIuWr/yDCwmFaf6TXn7LWkVRR5tzbl2ifpm0ejn76EifnBx
60UhLPmm/vcPj15+bdh/V0sNApsvxICpo1IelLTxFKOpVPw6VpHn+Y1vFy+YzKtFL5YmCxxQPqaN
bGMvbdt4jGWwmhHP3QeCOdILVjQwH0h1uMLj+JjHNLW/SYK8z3cX7UoKBDqQbXRICs6cAKy0342C
BulVaaRUVoNFNDymGtbCEpROsmaFLv4w6oXi3HHdjFq9MVcFIaVWa+b0+EOge3k1swPeUDqeM8X4
aJKIaEw6FM0A5mmb4v3+RVMVSgq6JOES2l5+WcdE9g3guqeWNeS+uxd//94//Ad1RtcNhCqj45u5
xD/oWnFXfqvNxZniJnnytCn+0Xy75gWYTRAr6b1bZzPEF/+8kiTvaFmW1uOvL+ctTI+anwaMs/C1
OlwFkarg5soqX6XlRRxflcjVijLya3Sbhs7XCmF4D2lXtw/3vpZwijrDtUR3zm9rcw/HSwZD6j/E
S0qD/0aGuHxxcXUQOjvG6i2Ncb3MRB4v7J5kRkdHYEtzprh1AVF2HUdRKJVQtRxez1IAl9+lpIb2
pRZUtY+n30tklgCjbDHEsQa4LKxCWzr3boG7sZrnudUAAnffgmaYqClr9MupRWg0G13+8yVpjc6a
fxr6Y9mTS+StWEB1rTM3utU34q/WceIz2GEAbY3NJv/7rp/IOGIgx8L9lU9zK6H95gm+pe3ZyZGA
3/r8FlLa4HT/38AF7x7k8wPtdPX0qQjgHj/VRj7gxj1gtNDtmplrOQ+wHRYxc1i6cmGxXV49EdYv
7at3FgXXG7WhjIgIYuR1MBrGENRJG2mA7X2H2HznU6FppSNMOdHkswVAJ2kWpQV4WOT9Ebb2qRMe
tKnPjkLZYP8eKI7Yg1DzUvPJhJ8fSGReG0r/ClQiVlPOI/6itG3sfW2F8BcvnKTOgUHrWrnbBY9y
l//wLNuwBgKxTwwJmE2DNmEERLMPN8a//OJlJqpHUG2wdJ/J4P7MTnHNSgHnXi2F3qlZd2Bd+gtG
6FcyNRIF59Grk2cIKOyA0qBpo9bq3zRSk1LxsX+GObV26DE7c93yFAVRmPhUzGDfvy5uCnmD3a+h
qR/nEg4cPamuCDhJHw+XBpiEYK0f9TAz+rDSzkczVjXqOzXHqoan+6AQkGHzDmk5MOzZ0VBFuCLc
GG1kzUQQrzTOj71ul0ccP6cSNbXxMnBqYiCh6HQca2W4ftjVLhHAD3elKdXki0KprpT2ncKIICkx
WOHibJIL/OMqpTbb4ynXfOE5cLD9244FqRPEzV4d9j3K/gAZACcn+5AY1+sZXqac2D1UVCDagzHd
uiDspBoNQvsTAztiDAL74FwsjvnNKXmr2+bt9MN6fj4mLcf4f2FoZEzYs1fxVOe5xN5YTvpnWs5s
hiJE7FNQ4UZemObItyqFZfx8oprmu2IRFMvQAcexnGakwsRO/wzWu2L31vsmMOMA7CEKZHhail4X
P1sTWW0nM85fIz/JkvpyFRby6xsvBZ0CN99H8iDBaJc34BUDVmGnlUsB43ZCOcY+Crcb4j0lVVJc
x3CqX10lKV1qJNc+g+8sJ84F20d0/KS69IzKFsViIPoCakZ4UDjHh3zqH83xTS8I9Rf5Esws/TlK
pAd/5bWMv82QnzCPgSJAguqmMwS5GF5yvBNViUe/n+j6P0f7q+h1bvY4Yf0oN1b5G9y0YZ4Jjz4Y
Hu3vbniQe1G7oa0+rrtUaaUE5YZVVCekQP9bfTZGjyGK0T3msIpRfBzEkZ/mOfQ33EzBx+QixNmo
COKaRbPuZiMzqu2SzxB/HURN+Qnkrz3UfSPAjcQ6mj/Tvd+sIdGDizhXKxDcNh3T4MHzDQCEMjAD
7rLsgoqi/lMLsumB+ntHIteImItfBAMfchOwThotYlPqx8ut4kcETCFkbd3xQF4XtdhBjMn3bmOk
J3QR1Kyh1P+1C3STOrGDQV56kQ9mHtozUzOOY6i57yQuCsGX2s37joR6S7sAVlMusFgK2cszN1DR
5HeBYtJCSCpsz9yuOmj/hQOw7liu/Nc/2PavC3NnmmcLg41l3hyomS0PrDazElRH2ufV2Z5x17Ec
xtKmqPhcv5oBmOkGFe8sTmRyf17dEd6y5zYQRxHNJK4n6f0XGdANv7pzNF0C9SRo0ejYVAcUzWKu
q8fR2FMJ48EK8WNXU+nyXlusRvc6rCQ2+mypZZzKGT/roTBTtzKbOC3Mnt599Ld33iiQI5imy2Wp
yr3KsrLK+LXCy3+0yFx+pnnv78HtKpj9hGiJF6DIMgIi5qXCmm7t2gUWM1UAMW1xFhRzlZvt8SOy
GpckuDYBlqWe4uQKfgA9Pm1TOjMF7vYomJk02FCMDTpCbsfI+I+b8Q09WhLgeE0UB6ZGVuDSDRwy
PXPeFO7RePZTK70jDkhvyb8MzmmFNZ6PtHFYbznUt/25gV7SLKWJxEDFupLVJCjlux+185CJvbPx
J1OUNNtbUGfkrtGSF8sJGHN2YcA0tqNIHcqCQaBGEJDC4M2hU9JnXe4+Vbq5rxqR3Nia0/axxbZ0
UKb3m4eA06yX/GzwTVnK19DjfbJmBwBrtYmXtT4CBoawqfgINtkNbpVbkE9J2tqgc0umzBVpHOTh
ptKMCaK6LEb/HoV2ysIBZOnOOZTtui4wf4UEM/qcuVG16FnfhJ4dHHyACeesJcnAmK/U0biWDg6A
+FJ0dWp5bq85nncX1cvCbyVpp1S3IG6wiQRUsIt1IMb//kVUq6BJdOVngDJO4cH+sUZB7AzcTU6B
Rf1nxU42c4KSbLpKtu3aSZiDrhwc/ZOBFsnlWrhlvMXb7uVyYQTUMSOAJ9rUKEpt2HXTabTSwq0e
FPHyLDo2MeDC3HmTHkqbw/ShQMGRK9Td3zr58n2LdEPiGoOD0zrSmBgFrc4hwalMzn/dZiSO7Vzv
tVyf0sgDn7prr6E6DRo9GzKRSAiIAWw108E9Tf8s2Znz55Z9oN8esiqClKH2HsbI5xl0yiSqMFlS
SXkbzcSQJpU2ExOM6iT8/HXLBsb1vf+Q4FhUBJ3qwhFl8bTfq+PwuwCO803tN+CV/QwN2JEqw/wa
FQ3wS8/LlKu/lqvJoKflqMNfBzpHyEYotB2fBjUrRvLqgwe9o+57rnNXAzYFq5XBjNgnXfbqXPes
mPe2f/MXXH8A1yWnRDt8hTsPdjAAj6cNPW3ZK0y8kJveX0dE/1cJ/gTubza2Z4uQB1MOeE4pDArd
SDkc0gC1wQ429gv7H52Eq+2Yp0RBWP3kCLa3tm3V1gU1Lb0e0pn6Vx8Re+tX/y0d6TppN7MZ1FRT
vrcNHl/R5TkJcCjWBbgbf3mOv7RSCniOgvlxXIgPH9dkpWQg6UM+hOMrdIL4VdNXXuCcwCs/e8S2
33ICsTjQ2rqEPwvBD1/QOJQCLpHKoKUZGn2S+YLUScXmJ6ZGf5g7CmnuegAYEETle8q1zQKBETf4
wFM3ZHSFujsY6XOs5PFMH2xotimy1oJM8rE6qlhHS0E4A+uniT52qGNULlY3Gl2dwZ7GZlA7kib8
R/PiW3/mfEdbYUHai6GG5CwmNAxtN5BmO2kE9lrj5KQji5vCshUPZVlfk1pQZH4cwPXS1w+wPx8p
CXswsYJar09x9CjGczr3mowAXHbtHDGwFunhoA/he8KUgmvAJD0QcBa+qCnoL7FnGN7kozEyo8dF
OG44MdgwM7F7KNr15pEg/NQWAbUscrwsNZ29g4NG/zxTSriZeYW/rHq2Sek/e3wUXf48YfhPSJyT
nQnUwh0UIEOCklhCQGnnN2HTaecqIPNcm7EGRqe7xDbu6HK5avzty66yIB6bw1ic21GsxWQQIrAc
wq9NXtqVdnhjiS7pB4TmDfnBudanIBkL0ByjEqjPVwgwu8hZJ7QeiXYIS8OOIylZMb+HkN77ODG3
pCXWqrdrgT6bLZE2c1n7QXZ/PGWCJGtnjE5VBlx3Q5etqO5AkRU5bMVXHb5dTCL4I57rvZNZUtCv
3sI7epSL+2aVwP2YE9d1t5VJGLHaJuc6w+2uo9TCTII2H4QObHhxLkpi4Ny/J/IWeFfMQQ7g1E3n
x5WMg1S5fKRn7KJ5BLU02MnQQ49vre0zbZxwKiQkxdqOsILPFn7x+sFslIr+gusfTVjiXHd6UP/J
dKJhbz+wCzwv1KefrZbtofemC4gmrVu7Nbl2CevmNYen6pLRaYna6aQdOr1GexiOQn1/ThxJZJMc
STXAwqA7ygj+w+s2HSwOY7YLHuQJXxzDdcnJSz1nLGEumMmFpu0y8O/tCdaIVTGBisz7MV6S1uWE
yAXuklYMq+7sww4wznw51gspay1Z8XtKOTV8om7oaYSsV+MmaSs/aJBLblpG8+YiSsCxNVI/bN5Y
1LxuWF8danIn1I/eyNKjgerlZhjdouiZzQNHHr53rsb/dnCmmR68idnbUfvrxhhRMXpnx/jR1hOy
UuwnYEoyenK2B2kVvGhUYt7N03HNJj85KG+ErLgt6XbjKPsNpDSXS9ZOzTzzDA/n0TaedBC7INS5
Zz7F47+mEqR6fstbBrn9kEw2mMyI+qCTOTT9IxctPLBLZFFjZ34nM+6TnNPuy0zDiIqwuOD1Qqop
JYRaGW3aHFeVLDVdZ2nCzc/1V6pjDsv7km5y1sOxEEp0h+TWyPdNaZ/aXxAQJTAjtYKA3j9FvsL4
/aKp6Uk5MxM/Hf35K50UdidXIodHMAtDlPBZVfAM3bTHFdB4x3OXjdnhz3NnQ61ixL86hAurNA/4
a6cMO13OCxrbQSzvsnyr7tRv4GcvKHC5I99xLfBDthynAxHT+vqOj0ZjI0N7ekSKPvDU2B9Tqi9O
SrXPTzY1I/Oic43SrTDUzbTs4iD3jmDeWKvPnveW8z65P6mAsi58riCYklz1JG1TQ1MDeMoSqqHQ
a+7+s77qXrUtgvvLU1V6eGzUMS8RAPofSaLFaF8o4ByiWLahFNQAMrq80I9tjEOcj0FBUKUMIoNi
AE76uoz01fzO38jbzPVESdqG8qLyibsjjBhCFCAGZkMqYEZDr1zhHTyy2fpyh7h7QC2gHUhwcHMC
49Ng0sqPPDZzHklWQoT0nVM/ut38823MGJQis+e+FYQ9QqcofEZvkRWTNu6cdzkSVUAWMiLBysbv
CSErTWhY4r1i02Eg+XNZfbTiqf5UJVU8Q8XX3IKZO57J2hpWODwI0wTz6ywc7wnIqXCZKfAjLNR8
DmnSSkFG+GxG3SGlWDHn96USBsqhUg7pKGi6VGsp1afU2RJVyXeGKw4K0I7AOEH1XUdwCg8GnftE
3SMWChehyrinztK5PAy6+Dlp/NyYk3jnfRERSo6dyKIgM/Q4pN7g0DoPbH087H9Zzf2SI9D/mfHK
RNN7jU7cjyQyJoRusqr9i8fAD/uFlZFo6d7leNwBDFACa+tevs2s6azMuMDZPXzy2su9b1mVJZXB
EJiz9WOJibyZNPZmLBkIt1QZLbNspUdYvS4DRLEGR1BTdw+mMNiubmMYQp7qT6utmigskpdB4ZER
1zB94I9MuyWE/+ys2mzQewKMrgWDKjMRNwDnQhM49ep8elbcAUD7WpnpwR5HYviIr+pzh3+/R1Lp
bsucHAE1+HLzhjgPR5pWvX3SMKmBsKL37fx547zJ5q0ImXqFO+yizG3b315Mq6vvg1EzKYkh5uJx
yagEuLWPISNlwbYGPZWspWtC9hC3tbR4b17gEMncEFLZPhqQD0mrfx8w3lWoZSW67QBJffunB2Yt
pgmV0t0MTjr7rcRyhV4x3eX6EQRIcGAxGf02aEZ8EQ7avHp3trDzzHWAWshxT0jBTbXM2SYQmv55
fa43fIRAc9Q/QaA1mhVIikLdajrihJRGdn0OghY4TYM5JqyjJB0cRXCGcYrPShC/i0Vgt37hvVrj
p+SQhrIvggGB3TP//IRnJ44vT4YZHQLIYWPWSdFIDTlVqg2Ox8hrkS3fLKXK6p2Rds/XcWoMwFW7
B/xPfvpFAvEEkhfDQ9c++XrvbPAeMrLlM3qJLol8tEbcnWD8iFa2MUexXv3pR5ENPakcB60CgkzG
NuyWwkE8ft+GmnuCegMrPPHWEj5nvqa85Osfml/7y5/MrsL+BeS+v0oJYj5xp2ItXuCxzQdvjB7q
N1n6yNPi9X3kA0yyLLtTsiCG0QOfwmwpUK36Cv1uI+TmGrx95fPVFFM65hjOPe5tkuF7Vfz7e9ih
iTjCe2xjhhobNBHV0cOqPQypMr1heC4aN+mI2uFl9iYHvzYe0RWQAJtcLNVYSqYYDDyOL3qZxW0m
oIhbX+svi3n2kOAHd+3Y5eFr1CG4+hsx0KMG6E98dR1AwuwwpqgbkYHrmzZiZSjNfGJv1E6Q7GUQ
sSuax5eB2Vmq4VAOTMxNxHkJMGILqZCjqCphXLBZxlvWXj8C0oAWgn8LbbK5rWNh8GRYW15M69By
IdIWuzB6X/QdstDovDn46Gl0qBmrklYYr6SdL1Xde4PHgMSDijnWwDQQOWbJTqXlDlLm2cOInfcK
0TAZNEjJG0xbEMF4Z+w0+IxwMuffpvt8SNFSU+yY6caG8ZMt4vIxrzoLVxBKrzSLN7VFhAW8g1cM
o14irXk9xXNGJLTQk+XdaJcndbyVDGraIc0uneOy68X2ixylYGC2ZQXP4YMK2gsYd8dAgSEMKVQp
CcIDOJADI00ECDYmcgfhWJ7JjAKpXLDrYUwFuBdsQjQzdvaRvGRvJzhKtjuDBlJ4Y05O9evgf2On
E/JUI7zO0a7KHts5ngi45LZLig6fGwvLwqmmaWWl5yOyCCFs5KYOcmBN7qTrT34J/PkUbKSftcWW
4xd9vbdlwqTl85EWBgpyH9CYFG1Z4Zj1LA3S48qMf9lax+J5eKEknYReRlmiIfFRCcaB/qJiM0Kk
Mrs9KeB0Y/QWMYReCGgXYwKbWJyLvEMOVHvyeSqe+LTmVFp7ifzWHVQRcDAvtSdNkKa9dbtQX5/H
je2+leRvkxy7RCeHb6s5nOOu8ggsv154xXhtZnDWOzEv7UXI24jlYOkbFoh5in6yt1RJX9aJiAwc
32uiTefsnloG4HTNht7IoNnWZQqw4T6by5QwUdcl+yBoTNutg+i/CsSgG6JcexKsKC4kw9JVC+LA
SiHwi3K/Fv1ZmqzcZa37nfwGrCOaYoAgBaz1pdcQn1KDeEXrIPsQ7mX/yLh320NoUKJ1l2IdtwTI
T4IuL0Nii2YtupD6MTHrlHEm4ROQJ47wkcwsJQUZt8TDzNdJmCQr2npcQPUBFU9i+SkS2vVofDfR
djA9a8X3EPPBwljxl1ea86Ig/KjtnMCKClMY7XqaVhimdjdMMXCdwWa2yP11cP0+2SVHf0eAZpa9
EUgWfnjJIFh/YqRUIWA8mlcsq/LVaE+OvmKfN4lzGt1Ml6f7SIKeUfPljvRkYhGBHfLtWjZPW3Xk
FookHaratrJ2rGqygaCW/yHFv5K2Bk5wSMNSws31AClgqcFFh2T0M0wpBjq3Q/kuMrxfXZkxh7IK
z05YhhQnr1hY3eYppEzGbMnNjPF7gVTz74d54DafwR9XO+Y6DCTn2GQwKm24UZKVRryaiyeD96zp
FEW/8wTeA7YC4VePghsPD7ukh/zgBmjagDNWdAWUn7FjBq4h5O8Q5FFntt5pTM2feaIJ9sfKXCAN
9MfAvrY/l4z0S0qMrMI6fPjVnY5gdUAgdAS9FFQmbFqxKx9YtqIRTftWsnr7MKdMunVF+rUMwrx1
N/tx2zmPX1bMbl+MHP/v6+jup0mRvUZ6Z9U3Ap6s+pBy34iNlKy48XvfycpdvZEh3JKt/nRCu2kb
h/2ztScsy9cdx5F6Q9BXEYtu2XdWPlCVveM2ohc79C/5JTkd/Pm4kjkofYT6W4obK9mlVnlDYg7F
zNVGQZd4dyt+WsMRSWWfuBLcQzALOk4VBX0M8aIv/5uO+WyWJHwfAOzXFR2nPqExDg+O6lBR29sK
fdKE5NrGYsz8/Le0NA3dEad7xxfPlsa/M17XW4leeXSE7i/VWcDgNvz20k5QdBIyotELdOy96s5E
QrYaj//wvKwV6oWLec67mfJxTPsO5M/lGeCv+tk/RTRSeaz0trxzhmV68mzxSqoWC9UXcBXMRVnp
lw5DPGxZyQXZIBzJzeZkf66E6+Q1H92/J8t905RYcBhdW7uavz3VTCQ/5Cdshv0jwklZ/ueZYTjE
J6Oj4BhIe6VxPnS77rHU9VKxmfOy5hxV+CuVf7Y8SzR/xhat5jbTwHqVWFFrRb3r9MwV0LyWkOkN
HqigtMHUU8p9XmpWBhbgv5YlQnqgVCFTiW8enW7N6xq5NDrnN7KliyP36OUIqKASbDErbKMoZ+8W
/QMrYJlzbhs99dmZDPG2yeCPz/u4i0DjwlIsL7ABKbVPirVWFu03S0pd+/hYb0qvsOASvKVroD44
qmBHWcLAxqi3e+1n/KS8R+tIDPNgrOUjj9sZr75ZHyt7g9OFT7U7h16ct8F20n55CtTQEllCJ2wL
PIxSJKd21aJ4oWpv9pEJnRHDM57IM4RS44INbwmp+2EvFur9wJL9eCFtW+NVVGLi2uFm0e8bbRTx
t6mblHiIKLVXgUlrlz/90n1rJIXpqEBWuB3Z4XtPt14kC6tgrZ5Aq6BWAG2AePTz7blaTuJx5jTL
avyy6D913q4njyDGX965qbz/JH77/b52Qi+q5ZDFgRAyim00k0QfeAR+CKUd2KnRFgrhbqzohxeX
ifdMVtlu7YDi98+thQA57s2NN8i+eOxuEiEZB0/woqc0NIFf2hIb6Au1cLLa75ptGvtc26/P7sT5
DeSXpPdluPiW7Rajj5X+SEnaM8owjpntbZ0HOlbehvqSjbBVQOWU9bAGcCbelLuMjQBNirULHgSo
e+UId7RgCdii4cbdrTyPQlIi1mrw8IZpcKQabCXOBXAV8u1QWtuueO+WtE95ngcUEOwCrjCuVdj4
vQ9Da/Wcdw341pJiuoUnUBIuaZ9E72a7RoqtI2PeXGncTUcTGtJoEi0GEFTKDwU4BGXb2USkA6+H
Tzo3O2zO6OMv0mb0WGJlZ4YRtfSk1Ok4zGBVqXacGWdY91xAPP5l1sl2tLKdGtWGxgysLB5K8Bfb
N82XpvzJ5jzRe5KSQ0xwmbQG6tCmIR2aC7emEetJiNnpPGLb1hgz2m2HJ152qwHR9dLlQUwSlPYB
erx+zhg8kwd9gvpOi792kk7iRD6QeYIMVs3qRnuTLx3ltRruKAkgEnvzwnJ9MD1TgXRAVtzv6Wuy
uDkTZ76lNy8ks6kMQF7YTU/Mwc9OlojbYUaS0DF5Bpw5WCtOabd21cXiDKjDUklv00YN91lOOA06
GGZRK5svyoZ3ze0V2GZ1VD0HPZaVb33/eh2yfodP6cdkfXHP3TUlIiuOu0iq3UFULEdC4g/Rd5oK
h199TFABS1bOWiJ8RrFu7y2LXlvfW/uzW1NpNRkg5epJehI7fbLbS0mgj5UCot/NKP+HygdMo+3u
BDWqtulR2c5n3mzHeyVqomygMjBnI/gkf/SpTo/mQsHmZjAu9gfYImLi34d5DGfettakzx/JA2DG
I2ohQrxnfRb/OdnWNT+kiZnoDj3HnTEbcCKy0ej9fYL0wnMD0SDW1BFNW5C+cFiS9kZpqVakk1tM
ZogAGb+2770UprQxb8olx4muFEXR/ZdSWirjNDgkVr7bQTueScU8/45ZDWaZrMQIKt2dfYfPotOr
yUQT3tlCD/PKx5/DP4/JkASQbKbYVltRxaQL9ibbZdH7TCArCYveXPYVJVWf49Bz/qGnyclHuQqa
bsoWuZ9XXUz1f+YArCHzB0nPqbsSOz8BsWagjIIWG4O476lKikpt7s7UIIIrGeHbI1OY1Fy3AqOH
64UkYicO/IhPxTj7zdw89XaTkd93Zj4DW3lSAXdmLlZSMu4bXKxuGBary37WjvWwirPaWJblCYJP
WH65byRAdC8OeSSt/drZAecqUCVlvOHhmTiOquBDdi5xkZLscmvjXCoYV5UG8ihYsrDt/EFPnE+/
Bg713rfzkkJCeTF42wWYgrSydTxIWcRyCDcyYqqUJK7AONfCCrKXZoIILvudygEI82AWQVnTszs/
cRkkz6Go8SMepaZBDQyOTK9pH24QbVjtEvSd9rg/zeaG72rQUcHjznFHrYTobjBT/6ecSUYdm8BM
pYMuU/2zYHx0VNa6zFDTNxdoL7knAy7gOTmiykScwjiddeWO3DUE1OlhczxRf6rc7bNI90+XRBa1
wwMFSv6jK0hP9u5IB6mvrbZOYfxMB16K+Qj1FJTqAiuNQncYkMpotqVGxooPn0XJB/32V6iCgj4V
ooKwFoUTm/5XrlJEVG26VPr157Nsa9B8ItkXgH1j1dpNitmWJLdnnbTxsjbuu8RT6sPuSqxVe8Gb
pfYC0orgJr0la1s1lOnNb2j/pfhEU4W/+9rnenynHcMUwfoCQOR6Kcuhkuq6z9TzDXUoRW+/QMBU
RJp9TByWk3n7SOzBxslYWrSL7ScEmcggDyO49pGbt0w9RI+ONaXXyg9kwD2GSSvvaFd33Y949uzV
RxccYVJDRlKI+jO29klXMXaKvXjZ0x+ArfMzMP9JClO28ez4d7wqwZPcr4AFbP8aXkcAX/kDZOcM
agJx3OVWNAkqcMF/qlwLpUViE1ppjmGlXFPuIDw8HMt3TUWWKOYN/Di4ofCvKx8+uQDLl8mfmQGC
7VR8UV8SioEl9QLiV0batLskirtYXkm4UOwiaQxkrJ2CtoTwiS9ZsUYxHkBgvUDWFlE2YnMnLvlT
ZeuxePLKvbKIkHVG+YHNjzFnfNCrxPNbGXx5VJ3MjWxZj/GrDsVgpOcPdD/jGDV84ehWxA7kI7Z+
X+9pXvlB3seRxxcoArcP+uDltm4I6GP/ksMQwNZrflkXt/duStKc5W6w9rlu4imQQRbgEwolC7vu
iTq2N282Ut7loUcwweufpGW5SY0cV2LiBb1RglrVpdYj/HrJQvRkQLJMMOHblYYQlwfPKQMF1NR0
b3/IwTPnzELAoOA8epQJhlIIC/5ytxd7A/zqgCvIzcOgL4+LTGh8I4OaRQtJKGRFTo7x0TkQAQ1V
Q3uB4CuOsrWC3J+ZMOHIbWQXaRV5FyMVmVkeXaL47EDsMeijBv/+2O94B+BnR+/t0MxziKTsoVeb
DYKlP6bx7TZMg8lGZqZHdTfiDS+BXZmgO1lLBnkSMuvUWKPE12cfF5wCwErKInOrKXjlGX10LZcW
qq/CNaRL42rPE0Z3vaqRAmT1/AD0czkCRp5RnrZ20kaaek9x0Z6EiXyCo3hh92Tz0bnxfz88MIyN
uqHXHiW1d1QXiseZTURM91FLjOSJWuJSaxIcR0jH6XcwCDizePCY1hMFvWAVv+0NDVCnnQ1kg7oM
kLA07B5Ust6NDEfSQ8Jtv8ksFEd8w89odGS0HRUIP0IR5HNAK3SL/kCM+cXU/T7RAwYej0Mx7J5c
La9+z69lEAOnZ9mngoGzgzRF7sjCmzNwcK0qOJUPCU6/N0MWprYb+SpszpY41FefiYxd/IQ7rdRw
euWEwMQTl0fMVHsZevGZlpCfLOWhS0FgrufkS1SGh/r83+Z9ZgFXf7bOB4ATu4BIh7K3s3ys8b6Z
yWMOR+tRnFPD8TmSFwFBygZegesKqQcQnofS1xDTQpTnxjaumk6dG/KMajn51tlhvhjJMrH7kYZ+
Ddd82GzQvbyKlm9Excy2/Wv0DyeqWARTFiiqRbxQ4DBOhxazsywNi2ZV91/MTovC5BQ7ci4ll9il
KqWKakaS7xJehiDk50PFwt2Ee+YfTtt9a9a6yKOPNmh/8frazehrtdqJnxJvnqFiTnAFbNw0jOCz
I7c5RTHLd3vmr6AsiUFYjL7fHhMHQ7SePrB24RqrcWMKXoS8/FGmkdBugImYKZTZ3bdW8B4af7yQ
ORB+emFHbXMrpAfnUGwJ8/sifSd5ZtothAd+gRySYX2EVE85MVAHzJJk0c26djA/KDJ7854Sgb5t
WjmZJMSy+TSJGOLjeKsUu9sBp9a/ZRY/GofbzZTMwjNAXhB8F/X4mlssztdHl9X37xboOH2LPZ/t
xnC5b3O1CjhKo34MoMagW+LEndx1vrcvupjGXGW2LYOs2p+lxnV3dB+GIlCMLFjJ4MDdOyD6Kzfz
nKiamNJzP1E2UJKM7j2DxL6e9/5xY+2UyipqV9Da3lArfgV6s/sqsoVOY58AU3iA77+gDrCQfJN8
gaphT/CKjQu9x7xSSbOR6TtnnCiHTHWiiQh+pax+lb0gOiOAJh9G+4p9CmNyB9zyje42oejIDdrl
UYbFvSemeswdY31VicXd4AtSHed7SKuHiwExjdLazQ55vWsHohVbTI3BoO/eJgNBUKanVs9Prreh
zbvoc6vLQ1CCoHT+G8UJyC375uj8+s/aGrxlnxi0pkO6tza1USZfUgBSrTr/edJtwJJFgGkpkgbQ
HouFW/OBjUICVAxwHbEAuWipn79tMQpsXDXcKYqcsa6H6i9DewZ70Ivwb1Cta6x0TGjSiUkyMVZG
gUp1HU/bGU45yQiiUHYMOmT66qDxNJfZTlYmBu+uYs2n31mu6yA0ej9R3P4qz8rYueEGu+H7BE6j
Q8uRkJ/5SgUJpOYIKhj/JYYvjI4x+rtS1manFsT92xHRnYo+jxmD4dxnJCePXIdwigDpkFQljjGV
OlPVPBstS6xIPyD3ChiX6kgd1vEvRfa3GYekTlN5Xsq+lOlOzKT1k4HbHr4gCxe6B+QbrPQ+HZLP
gEz+b+Yc408Nq+7IGlj/XyjMeW0DMpma3itjK7TQfh3xP2jGaRHCMOavpw5zbFvcZ6GZIA42ceAr
sslb+gzt2DQ+3szigursu+afNJ5m18nNF5kw0oGlU6lWoW/bf7jiynarQppbLW2GlU3kQlzzMR/2
SqwHoPQ9wIKYk1qT/6qWnBTk+ms9T1Pt20T6nrzhrPpkPfTfRRa1nde3VKyzt+9Qxwt0sCO3MVoQ
XO96l7GPDIbnif3oDl0zG/tyUq9t0A/6uf+7m2VEmCwfI+F+WbBl4ZhfjCtl/SOBYV5DTpHUsn3m
NBxXfgKVVAYErIQ1Nt4VTw0G4FldKKPRR7CLU4WrKEH+6iZuDMLII1ZcKBUzU93xqpqB2yabbbfc
ZFBkOFlN5E4TwCyG7r6JSuT8NdrHK08A2Q3khudYIMr8yRHzve4uHPOiCPnupN2mYig5pp2SAb5B
Xa3z5vFyeMwveWE2kbknJLIQCPoUXGEMmYI7MvkNvyq6tX6B9PHOZj1t2Q7Zqf6skfDbuJ2TNQMF
8QjZnM2lxHTaup/I8tetAQT2r2geOT6R6PZg8j4GJeS5viqD/FZvfSd/uMVhRgq4pWXpR8cJ07ia
Vz/N5e/abGbNtox3Wmz1ytw5DDaWDlU2EKeGUjhbF/5+y/3aUuecjQZcs2oM79r1T0GWVS1TKwP9
2SbooyISDMj+BB7Q+F2L9yFfKM/Uo29gN+JsunyKxmceYy4a+vKn1s1I3aGf+H31jvKqthgGmE/U
R2qUyT4kU8ZKAnHuFqhtzseB4QCgJMOsdtaaQ5qvVoW7vpxt955JZ7ouk8M4J7N+7zv+d9c8bgRW
g6NCEKzO/auyHbmaWiN/SOwETJ7ZogFWQ6BCAvxbytXJuxmTLMWaZ1HJ63U7IRb6kqVFkv/7k0CT
yIc8xlYKybAZiLCiQMq8d1Mqj7/NEvUQ48qnIV1lpZfZ/7ZMyx7zTYhI7+QG3IWsP6oJtxyfW+ps
vmTnWdIzWND1IbwJ1QVXz328qbOXmajYTjzRz6jG7JzSdrlgjMke7OrwLcV0OuMpIpvFYcQMSuSy
/KlVRq/xUTZd7OzbAO7VlB0HlWvjZzjqvN9RVSu6DueSSOKJpk884JvlPefYNab77RfvAmgdaIBj
Q5Sb4GcuW3yG4HvCLnH4K34FSktmHrkSODN+amBTHEDZgHV7SgOJ04Q4VvkR+0aRtk79Ghzxh4Md
5gXtFrGnXLoX971oMr4FSq/u3uEaodBkvFrRlTocvNDrSukPHwy6Lm8DjcV/8qLOuxSKyFj/yr8Z
X6NtyAa10KQgdcFIEAhqqkYeK1P53+1Sz0okeJcIiVsaHTwhW7JingNw/7TSfGHIbodsgzethe6l
dXez/J21oXw9NlFPP3ntOyLP8GVMYZd8TlrhadyhcYFjtH8ROjGdikR4QlcMqEs3qgFNJ61Lpb/h
+PYaQv+JtLnCAybXpyr5XsFLAxxydLCN8lznqC7IeUcUlipmUevuaFv3muxubNUqqJAHHDGI65iK
Furzyi/35qV8sAum6HWH/INLIBNkhKLmLpjK2rgUvpzSQWq+1DbAjmT+CCT4OFN0jHP7IUTm/T16
TefUP1YAzU9A1hFAWU/Q3mzvSLXr+1GdO+go1jYcM8HqP/N2tDU2ogohMCrKOOOJ7HRfsF9SCt8u
b5c5xTs6slGmMkL7v9RgxFwHCf6fGqS33WZgPMzic1NOIQbwVNQU0xaGG9I2xCHUJX9jQENtFCMA
Kkgowm7ArQ1DQtpx+0zYyF5PkrcPIQHLG+IzstzctAGjCBohIjaZcqIN4AhE3pjUTiev80eU9qQk
8CAJv6AW+1yYtVuj2u4MrLNtBfZcI9L9MdhwoTA2ZtTrM2JZEKTBSds2lVq1MAj4jTZ/rr8iFUSW
VCE3W6FhcRRwAVdEnvHtub1SYayEwEB55BYm6QNdOXx2pQrwUMFZHUvHuROBruz1oVLNVqKwlBzi
ywORXp7k/xMnIZQBni74fnn2QVC66/zL7+/NzZl1DpgelRF5IxrpLNmuimNaEn7Eon7l685lo+wy
YH1PEY0MypGaShQXrgbYZ9x4Sedmr3hRTXrIU6PX6cUaGlAwTuGtofOx8dkcZuaD+sJusIpUulyM
QYlPyaKHedZEKfbbTmMiJ8BT13OIFfaC0DxhaELu2SBuWacg5m8joJIhvqAlQh60V1ebS2IJpUna
h77XArthpurv00pyAaTDiAgbIpXo43m12JYn99DQQE/gehh/kgmHIPC2Ywot9h7S9MrQfcJgdmNF
SQ4HLEXIu9f1Jfw90fK7tO2ykUAhq7n6JnBTx5sdAaOXOnxhDfgI4sKsY1FZx/KxJQqh611is5I0
71WG6TCfvPU9yncTYGUyueYJr6bmU2oy5+pp3X7mztztoAtaq7Zg4R2lLmTS6awuCUBMpLRhRTlJ
/jrnvMQRBrhKwrMlVSgFUAfP6u2DhC319WPe+B6fYy76GcDK8A0WLEjOn7CxCrP8/4ZDQUl3bQRV
yNHswhVhwI6w2B01Qxw9xEZ7VuFy08Z9gAyYbtqB7GJTqZQssfOflOgUCmKaVV+f5P8//gfEY1yW
JnN2mzjw2Ryqvo6+v6hi25rUm5F2JPGipO2XxWhQoueoN/6kcZTorZCnbL36xMyhOOHWLjNv4WvW
Z/eVDQlWFzBKV0yS2h2jzbz7X+t+iYP/ejhxwjo04VANKPXDS+d1VMS1T9FraZp8edlwGXF4Z/W2
JltCXm9s5cvWtamcJ4szDo/tP6n/XgVwUXfQji0xcWnWuN19j3vpdrZS+t+6fDmc31RPvXaUOdeS
SHubQXz+qyZLoilxdPOPert+BEjvfP3nhMkdZ7JQ/VKAVZ28y8htrulxin4yMWyCJ47LWdXun7DD
YeQso7d7G9sARLWR5lEkdAy9AFXXOxJqTW/PF5/JZ9t3MLanYjtUgW2G/lIvuHYlG4MlZwuYXDgu
PLOoVeGo11dH51rk61pguRwTDY9C/jSdpJHAGNOkQknxmCvI2pOa3mK312BM43Ze/dAGozXC72pt
FZ4Z4L/zjbTXwdK88q+EyyLkW0Qoa0P/WjJLk36loQSvKk+YSRtpf0tcm3G5Zf8Tz2WvGOKtd8sm
gp+255AV3dVPQte+eop00iE5quaIywDBpQ3QXamvIjX2fWsCCXbbuKEa8s5LABzqh1Rdax1sa4Bz
AncwYwWdXLysgx/yfejFKSTaPqdUX+heZ8Guxzct2W4KNpsiuyo6OfvuURzmtNv/LWmwbXUjqsp+
fnm5zw3657hJJ2tn/dSTTLgChGmiedNIUHP2soaG40OhUt7Cnby1UTb5vulEvE3ZBPGFF/6ITb66
fIchAvY0vMkj3mCmTfsILNC+r6IZNr74g7BnjM8Wxx+T1+ZMbJ2wehVNMXA4iQhHwxTyy5IITL2a
AkV0HljwW4A7lbqAaLKJml0UuDwOa08c5d24LxVwGP7gAGP1j6IGMRS+fNXxEX+WxkqNJP4PSUj5
cTcsDB6I4hYeWyI501Kd3uJgMFsOxNplhcsOQmWJQOB4C6/Rc3BeWBjCGieqqvbU/JL8nxEc3+JU
39ZhgCtaDc9sS4C/Buw+ZGFwW681af/lme4ztTRhEF73M1EOsQWB9OuHqbT85bCcyCIXtNX/Vvem
szg6bZME4CkJ/UarsbU315DIaBpoVQnGTMj3okMEQkrnY3ypyBlqaTWSJBZqFGT7eAMxkvgDGvFk
NA568Sl5MX9aCya5dJLji2CgcVrvHvYL5GhKrmpyLCfp+QFiBcl6N43ixtK1SbBhCO7E/4KVA826
l3n70JWQh+o9B68FjOWIIBfSRskAqijF2FP0f2mzeqHCPeOYEg2dUea/+Zkh9PDV3GKJldsbB6o9
4oNw3jSVy0FCgDzO6VobvQCZ2NfSOJj9axzwT/sbOj9RRSuosuGtk4k/DCqSU4Lm0x4uE3Q5k7XX
c3WeqZFbSJFeFPuasrKgy+V1HUssV5NUkEbKq5r1E6m5EKxsnuIVuNTHEcnZmVYedloke7GMXNvT
EnnetaSipHvoDD9ybjnT8haWuoG3YWUF1W40QbHlo9S5X3LHByxnVa0My4z1bFrjL8fpkz3Ez5fF
Bnll9BLVeiBM/0ld60gXCfMHWTP4X59g023SelN1zGHQ4n4+aIygXir2eYGAVzOkmFDrlbUtZAMF
zwRwnHDNkAkQu01zzU9AA2ODK3WW0j4llrDTFy7YmJh6M9QCHmFmXKtiYzrmSsuuTOmzqSURmHOk
6O+YR8rDTKlckm1rndmlB8rdAYYJULFtwdDKyzaY7jQWqTKKkHA1ZAqcIalo9+Q/FgKWdFhlMWx+
B3zFxlVLukFdQnnGE2ein3VRyDeMZu878Q1dNj97dELeY1x5f6dFCsja9WjhZ8UoiWDEvYudhSaL
EU8Gx51l373C+bY9IZ4+lbg92iy1idmK5Jrj76jQiR4W7tXN9TEBDaOFmeqg2KEjb7sn12MdvDRi
5RvorPNXVjt1UfgJM70rBz+s38X7yswwP2RhRQ4H/ez0+GpKgloEzxbeJ0efgCB4zxLgQQD3SfLk
2RmwWYlHsyoHxC1OvcfF7qx2pLdKelAEASPPWJ1aNyO9/+R8TVaDGdxXQi+I1IfRXXPB40/83tFt
DhOYtGwOd9JkDJJeD3/hN2gUBBdP2nQv88BEs7waO87qIJts8YEPt3yAz3H3SUiEbKKNK5jd2xlz
jDnSA9WC/gQ7vvg3/OgCSg139sV1jMiL1Py0i2NXC5OKPYB1TDn8HmgYJF8Uo6k0WgV6MCpSHHNe
AexFOpk/0yWkPCr6dEAQ4xI5DG6F+H2ienUcaQ7WlhWxSA+bhLE8h6nGoQKDpYjtTjT2dIusvlCP
nBgwJaLjfbAWf9YIMnuRMbU/ISbL8D6PvdjMbwiiqaVnkOzOWY9xINYX6NK8Eg2r6XSSwm/L/lKa
i2gT4siFNZnZklzF70SwfOmsiPHQSgyyoCfwNpCI6lc4rZbP3EN7MWg1cRJl3kmqisHmgSGRgKDO
PnPHpHZmBlmEYylF8jjO65QdGctpT22UuxNhdKZI3NOe8YC6jfh69THZlf7HwR3w71rHkOxGxwky
PYhlxfnZDrEHe7HjL9bUfqiOduH2ADliWdRUZZ4LmXXK+irI9f2XtdjhRcmL+tDkDZq3MqZA0hQB
QdMwSgViEwcxdCBBvs5U4HIraZ2GD4E7910ptC+ZUoOPIc/Ys8ehsk0dBKUdfqGGLhfGBBZ4pH7R
XGy4NUOfX3Yi+WGbqa+R6Izj3Ewb0VGCDc6QKc4Qy4Pbwv/ZQVK2PGjw4OvxxaYyYupvMCd/Hgiq
GxThTtVPHA0KRkaq72m2eAeVHRRznxQ4O9nlOyvtrjjjEV8q+Nhd/pgZknclh/Q3qtbIX6P9dL7r
v8UdCFlgAhPndmh5yYYbZxS9UPfZMWwV9qHVZ+XWT7G6JHWoHp4BwlHzt/7lqu0k6UKoHOlb8EJ+
bWl0V2sy+rJbWeU8HQHy
`protect end_protected
