-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
BGKYNuIoda4/Mm8cI2ub2jxESo4+uofgwISzCj7cK3RDQslOQ40tNmUQaLa54CMNx0i4k2fP/f/G
T9jXH2MNV+aRJ9cJmYsTH0jfnhFDGFJG2QFGMZsKPlHnbjKSlh+ivSO0kESwb6A1ZXQgvGfotRgv
pJvq/VB0fqBwx0M20OYSBkAoFNzu2E0ggi8q7CWQflN0TO22En4aXH2OMs5XAWu8O1+m2dsWyyjE
2Z3zIIeBVfBn1VJQmiTlyPSHSgUHTqA9zu5+XyTyGCruNIRgZVA1pE5MUoxWuigo0XMqJ/rC+mkt
RV1bv3KusF32DvqGV1pLkcmysNkkz3Ros6KNcA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 9472)
`protect data_block
Jv/G6bbIWBUcvkfd3yh26d3RR4a5kAJ2N9yR0NlznBbSmYAo3G8hrv0itJi1T4kYoHqt0o2NB4cP
QLDYhLn64qu9DZ/ow0OuLl+UDOGuuWM9++zIXjpO0pY979K+Pwc63m5+2PbimS5JjDrUxp33M9ZI
znYNuFQIQAk2wjYvwMgXM5UIIoQdhMTTqOeia+4eSP2WzI97I81SAYAsHFtx6kntLosSx5YNHukk
VSMjPkR5V7sTRbTWXS3rYmrOFv61U3MINLQpP6sVrefKw1dL2podQLjEqxFg4Do7GhFPeAzN6Kvo
tzXIK4dqXBn2G0MI1yk2uioLZbaTPjXYy5YEF0/EuCLn5YXhm4/zcJzf04iE0WbJ4i7JEDuOR/Me
V4FxI/ymYwuZJn47Fp//qs2iNd7ZO3W5ilBtUKgvmRBi68vCdxPAIFuklwVxLw6mnoaVUH0QHjAY
WhmbTCBDujRujwvqQhOSUPR9UH7vvDsQllG/Tj6PBElCMzq+fdjaQ5Hg8uqofWMUcpTV/4IxbNwk
U0/aSLmYRAzYOZSZ+R1S7JWoSgaWN4wtO5wpKc4dB5xQefFXUBvvbtZqfFEvO6qblm/wDJSjIkik
gzFf+sNfu1Q56a0tUQ+O9EH1JBA3mqHNGfrSEYGYD8VB6fkMRCWS8qlRyHbd/cyVuvhRq/+GvlK3
0wRw1sjZUe3kYZm8QzqaMET2yvqf4qbxDlq6sKJdk3o5kYQ+GQ9Oo7SQTcFsPlLYI40yESB2UuhI
LxNZh/fNJ0yFjotp+2y8NxRbEOtgSv6WpbkW6WNlI6XeQI8sp5qfQ4Qr9mSLe93WPqU5PMILqPkJ
yh3UAWq8bXAO5ZGmNd8rIPUoWbhcRAB8PIlZ8ZyiMfaA3/KzByD2KUHNRliJ9Lj/9IGG8etDwSkj
63NkB6TlwNQgV482l28xtHciNlREW93p50j9icHlWFuiofrBv1PNXb2AaBhV3gP7Lz+vqCPVbIbf
zTuXyhol0PiYN4IhgTUGZU1U+prCstk4/8Pl5jRWCITYhcW30+FrNKVaWWGBdsvcDOJfExAeJqKD
E+PhxNDxO+c5GurTRPYsWjwJ7hTJvBQHYQpIeBVagkQWsbdV4IKxHAfdJw4vkR+Wv8g1AObQ2JH0
nVvGF85Uahov7Hu9KzXYqNe3zGkBpDAyjJ4ThonyYTi4u6usKUPVEbGeNmnbrPIELMCsf9v0lcjz
AsPKtp0Bl8Z6gc19uIkZRsL2+tuINOfmSDVs0N0uSOHx7z7q+Oub33a0TykrX4f3OK/XkdvKlhU/
4YlkmvPFyE8iJ/UR+497Ac4RxqYMg1/8azlgN88emjU0MP9Kae92pSTwLh2RV0fq8cSALmkghnV5
zddo8hdhJrGyWIBGzvwXAV/1MIFM60P+2zNxgKn38A1DzE8+AOwSDV67L0DDKo6GnzYPHxYb7q8J
ch9juznSc1YCtXE5Rk9aHD/2OBmHQofFR5pYwRCkvz9TyIwlF1UhnSlSAjp4valJs/Uis1XbmHx7
0poQNFigrjo5lr3WdybvFz9qoJSZBQ0zhO4tWxsISOo9duyGKDgpZEBPWEZYWJBm82xOdh47aimP
6yXhA+kpAZuSshpQZm6ALvKcoZsoYxUgu2L5Ur57qbGekF+cI3y1N79wzhRPE3pIVlDyL66gOOqD
x4xq8r+FPzSn+k+2lFe3q7ZHmeWLwQh1ZXtbYZgplfO/AnKxirPKW1KaITcmKy/PaWPamOykSIzB
WtVDXSyoB3PUvh+fePio/AZCfBsqcG/22mmGvRIHZDdfw58njrKuFYU9MeHWWpsApy1WCxpuVrXc
5uRbS6ptuw8Sm7j8/rDnaaePmKlY5B+lXV9bYT9kB7vhNlR3HBJpgMLmr+RVflscIxJIP0SWq+BO
UmeKpoinlNtHKGDUCuvByzJN+3n6mi5K9FN+GCwXVaszzWfcPdrqR8d+8od780uDndgkHUYXk5hh
ffZeAVTbdyGhzo6PtcYe6csaRWpE1OM9x1e+p7wvpDlegyh/MyhNSbDs26dvud9lpVT4zsOBc2Qy
/4hGrwW7uSYYremONT7L1pUkeUmWkL08JLXAA+Fiay//JY9Ze7F6N31zTmiIu47xuAJUBOEuX5Gb
fiPbe8cSp+cAYPYwisvxrElrCKlUahoBV2LdODb6XcP3g38oCPpqVl0HD2cNafugp427cFkXkISf
ogJzCvMfB45/38WQ2AwGmNxZOIDxnmMq62xZpia3m+unTvYRgpER9KZFhjYOzHoLjSVwWWhLbW64
HjQgu4K2TUNsCVC6tErYfJ0pSPmLnekJuB7w7tsShnnb649Zc42BfSuoMc+7VYO0pT1BdoGOI4Q0
1Y2vsfGJw3C0kA8SKsazrIelgGzntVedwiBc0flF4ShJ5TNNSefOwsXKK9J4nnSIh5BMersJDxtC
n/qx7GX8+Ie8eebBlwqLNq5hhpkg5qPFn55colF/S7H2sEd7+D29nlwoW5EwyKXbdrsxqoHMjZXY
GatT7qvuK1DXMjCoCPYkIYrV965/A+yFztCYv/w8c0pOWZrR22wp52SBEEFcYHfMAmGn2Ljsms0u
Q2XQMEDDMYHf2kMFJYhdbrTdZgBz3KLtF/ZFDizvf0+0rh7RJL5fBWQJWdg2/dDbCy0dnnxg9TIR
fmBxnnYWB8a+gKqSHNsU/cpmQSdC63YeSUcAv/5TaZ9tHffghHTDq6eZrep4BMbodTkUHKh3x6wo
gqdf0CH3rWxjlsxN6mXEJqzmJCbUoi4RQ0HEtzcw6MwFSVSs/EBcnEW9P+XjcdT9nW2KGduJT3Uw
lcVmk2Ay+kt9RhtTWLdlanJIFzYAtTRpArY6Bli+LT87i2LhdcLnX2jVG6qkW/zh0dzBsBR+k7Wz
q+2VmGKsJvDNGf2AKYe2ngZySw500OzdLIE6nYacXT5v1/xe1zxD2BEiuqTq9QufeKY8GphalV1g
3SqTEm+zYTIIPC9JUv/gT35dSC09/2t3iPppbGBSFptxx7yYO0ESauXdTci59bQH1V59iGC0/Qw2
mOnBAPlyOMehB7ZCWvpVcE9xQNd9Bkb6cv7eY8RxV4BfCc78kFnFQm6inb50moxXMk8JIaGyAmkZ
27tm0HomDj9wsU6EhSRY/5KbF76XeiV+ykE0MIT8y13qqyUTgzzMcEkN+WPA8sln3WPGdn8xnuKW
1mcq19qGbcG6bzTvzGQdyd9ZMcSPRfxfzbK5w7qXTWsaKdiTQ0hUqpRZetmZ9YHpXwbrU1DIygBP
NmVKg1lnaACxzb8VDZx1hD88mv0feDjIeIr9bRmp46AlYH1bfbWH2pjGbPfF94beGwL7htc+KqhQ
5/rDuGPejX9uaQpeW/dVG7bplMc5FuJSeE70mY5mMJX5ZrQwRAUmHVpLSRvCerlJC5LFJMecLhTA
JIzyMebvMyDWZ/TgJSoBH9x7+Xq5E/lJhvJ60sHsiYwmYE75r/4+FzCrMVEVYwcrmSlFhNkmc1uP
6tXLS+B/pRCAGubIH3qZXN8qVhpj/dyAKRgL7FfgEq7ZTw9TFAeIRupLr26RECMp8wTWhSoIO9gq
AtF4Dy7+iGqgIZy994dKyH+XBwUEwzQqpyEs6qNtbEh5J93RPa4svGy0+Ec0f+BUghcezTW/2OcS
C+KqfXx2RovVNuHMXaoNAIAVv9EBddfl6I5vvvP3hIR69eW5tB1duP76HRBBNvxFFSq7LJUE4G+j
3oFEX+tIG/zAFMNDKIbkqXwobTjD135fVgdTPOuIr1djtOJejos7TtIIvHWVHd2zKW7r3IrppcWD
mmqIerQ2X9KvOCl2CRI3Q09b6pnY++Jent48wxHhBtgm7atCBYqKwjF0MqPhFV2CqEHKKT5cyJws
NPId/UDl8B7txEmgkfPZrAwHruBdyOeDfEectKnOetQZRxPq2eKvjj4P09pMBmUu70gD9Xe6OQ5c
2OkXB7yhScIADRhqRysJqFXCu3sEmq8NKzb159XE08S6lhPbx9hCramUQgd1z8PKRoymEpVM4glq
w5TkhiGHQjnyjVtpA1Dv+uKy4phrCAtS9p2HWzTPEYcNrAER3ORnn8QAIhZtnUAIg6xewW33Jh2H
MnnJouyqJi1ySe4/p0goMR2ZRPMrImjCXW3V+fzXbrCXUz9liUfIJk+pD/AI06iH0S5iaLPT6C9a
nxyKa5T+2ZFjvC75xHmYtysOCo5pN+PV2o+yHZ0MXiZF4r6A2ymB2AwMxgwb3x6+DhLzbYqqcnNU
jlTd2Nw7gpesdfpsT8Zcdo29zqszFSeQ1T78+z7nf2hwV8MI1TgWoHNXAYHYH4pxSrWxsIdpXS3/
KZe59F0ORq5PvDSi30tJlcfAhJp7Bhm4DBSQDXiLIuh70KiiE0I0ng5p7W2JW8y28jycDiRLZC4x
Sk50fM3iJMef3mShZHLp05tswQDg9cfxvTw50hh7DAPNCTwSagoR2sNgqFxvYqWwFyIQCXVM79OT
my0ODEcTrLtoPQYA5boS+aJbphYreZE8izbYwa05KihnoWzXYkCg3f6/CPkJNzHn3dxbV+/SA97z
dZpoUI/Hsoha1U3dH5XTKE+lDm7I4lR4nFMXOnLJPJztaGXnhpGU3gNqXrB3yJAFINePjQw7P1e7
bbnNdNMMVQbPEXpmXIecbfuVSAAV4BT+mHSKcYUjOf+V9oo91i+DI+4Q+S03Kxsi7cxsMa/603UT
KDXdBHajisaGN2arjq8EBzr6FGtbofLNW9Ku9sq4c/iu4Gbs1uR6LicIUab/lCW03ZpZmtdaeWbx
6kKXCVeNWSGKSsByQcPbdn5QxGgQOP7ggHHD6JyvH4sxnkNTXyZVMgDV9jrNZdBBVinHoqEbXWN7
bb23IasP/TuCPa+h9oLdDubq4brZDVUDxFnsbD1an2sqqiWX/2eb0M5sgLzsYJVzUf8H3odweWHr
kyGLp/Scp129i2qujrv2xZEuScAQTKhqzIDYO93AcbsAM9kXXtchOR18Kv5Okl9prqbnlZ012ez/
lNWkGayHKLyvcN1WUi4qJT7lE6tFFD8S77tUi5TP0ezNxdco5RpE1nz6TgRvF+qiBvLzC/tKsG4v
UwzopSZNVE0Hm+P05QBaNnoboYtOQBVMDe0h8kxBsZX300VdTmAT+5vxp3SnaS6k5QRlpNVXBSPR
G3PTFDrU0VPz0/0tLdrAmUo4+wido1E1CszwHRTzLLMdxWlsoC3vpugBcBialx5Z4HAKYsvHZ6cZ
QRSzdYhCsGwSeMOGBmBDEmvrmPwKmHNjU42Ar+Qo2btmZtGPOLM1p9HZHHQ9qSJpitWiT8KV0lMH
baZAv+ljjGgWJpzEXbbb96vWe9wtOfg27E8vta4qg4PDhPuENaAlIzoCCLnh3Z9OheLAGk3qRzic
Y4tGVIC4QpMOyo1QIou47VUv85QgueE8oH4TbGZYKOmrUiXh7JjxBcyJtdQlj7Z30cpZ3J8mNPe0
dEAK3i8diFPTPMct7v1OKMY5s7vXBHXR4JQwozNHgMu8VJzaT6p2VeemA/LRPyonw5LFDfrxk0Xr
LabWsslNxZSHTdHT0CyYdBAe+J87ZCTSpr0OoVoMz/9rpBsxGOE/srU+sFus8f6xx2MFw5sAA9DW
C/7Dh/QSYXq25RzXtrI8FpmYkRdxYSOFa1JIw+sNZaPCM68N9GD5KvIIi2j1iXYEvnvz+fqW5a6A
Noi3dtlZBzEFrRs+uyuAlkeKCAbB21eWmRUa/zudMX7lHmgYaE2cgybuGszTyGemDhhbobMEn5hd
JX/GRLaW037hX8RVw+3SZA9ZQsCJNPqi68PBovc6R9deLCsbhcHPd/5ERiIJurinqFOQPOZyC6/n
JW2NPMlscXPEZbxY7haa8UYbjHdMNanLeBO8zSm/4QP0h02pGj0mbFOiDAoUFJb1tki1mvGVc6eK
MJMCIAZ3RGFdFFTuGCqDvvXpNpglowpPtA6SQVQ3sgPK93cCPvA0RjotUS9emSfILv2M+Ry3tGPs
bbatgiWpzhaUQab5NaKH/PYb2XkAoqsgLl2e1JJjal7Rr/YnYPlUfQnzGKz23cGt++kPnoLP0/E8
SyFs0+QUxNScTvBf22gpjNKiFEr2WlwP8TMYsxTHFFNovD4FKol8QZUCOGscI0VCuw0J/Hsq5T/G
iFn77qPTC7wtTQwBXHhyOx6beHBsGojFA42WyR35ncDcmb84DbGRQ3Xdl0m0Tz9xqJbmVyRbxEBa
X5eOAw1wwQQ3bYfIMf+mx50LcmGC8ApQvknCS4kIr5ur9oLryJ0tH3vYNYnstUq5xBloCstiPKZS
XIPfzxPOwDGl7qJiq6O9Fwcbwxg7VBNp5qHpKdE2ZQS4wO7C6YuyyHU/7AOtkqNQc8wDFZGfSg5v
HibK0mkMoKjKM4yYk1eMZd4Rfr15yTcC8EaS59JFb9kE4kRYVFlLVnIbXA33gmozqG/8KToG7flX
gsRIFm/qRdaKvOWhYcccwjEU0dPgNW+I1AQ4zKfAOd4BkEN0t36155arvm660xlPrJ35r5fTPdxy
8qKJ4ZwRXa5chnYoI0oDbLdSqcYu7XyXo36GHjPECGtv8+bwa/xoEMtVVXX5ICrP4nSwQnQ9GuW/
Far/7sAbBFRYQfBY64wpA8x9X4YZJm3DKht3FogDrL/LNTSZzfk0APNqj5xMHmostWtPjrLDVbjM
0TC2/PF2xUiBeiwNv6EPzZ0gRhEOCJse+O71uxiOofpAXhnkacLloch/b+GNz2WmoKIPFsUxYx/s
M38kiGnZbXugfqmMKdch/wkWPRqXBTB4UfObyghrxHPzsahJke+hUDukExKJ9H/hCqfkuFjkl5VC
PW6sr9hrUAOkQE2x8IyPHLXdHUo26ePwV7eU+bLJRI+L9DCtvBbifucM8JV8A8C2f8oRfjTYtt3E
KJL3LoKfXbCB5DfR2KBP9lHP8kVOmt+fER/H4kDZDRgUqZqRLk+/SEbirHYNwYf97GbCvp+DpwQI
yUKH26U0LXwvd+8fJptlQBm2iXky3mEOHQxQccX8TlnvU1Vr/sqVX2UwRaJJ3KVK6X1TitfF8DIj
y8HYO96lyydOVWP3yAW0Md73tOHmcGmaKMDo70+fIDly68+6FVUicMR8Y7X8VvqSr+8Y9At/tcCo
TdR/TnjHHt3nfaY9Yjon3Rcl/Pco7Y2hVIOrhyJ1y7VgTWEkuiRDIrhIN0aVuBsQWxq32AauvBf3
s92x/0uBc04MVDEmxJIn0yE+7Rc38R0AZ9vfPheZL/5ixORAX5KOfOP/c+CkmIEHvha3v6/YZgEk
NAzp1cEJZj66IS8cFpSKeyIGCU4Bp0se77qIPnw+awDqA26cfJCZgOtU3s5ijU5FbTOmt80P9G1X
0MGTdPKpeDTPtU4j7xEQxAkky4ESW/Sn8Q6IicPsMoFkPa6GzB37JZDDOCaPVpag9wWHgGeP109R
qzJS040B2X9zr1JCcFBAwhBwE0Oosfq7vxx854DOF0j17PmQlCLu7E2PUCgrDA2QgHt4RHom8T0x
Bq0rFJ0DL9KneU3HhVJ0oA1lHj5QrhHjR4C1aALeHPDG8Ry5R5Kz25/PA8CNelDauK0jVzjR3Ffw
ICRkv921+QqCM8ISjS2FD5NWMqwkJRt/gUk4+H8pYFDRRzglRl/nVQWOoHjdtfm4ADIl3q3pzFxM
3AwYnTbG+TZofkczdnQQc05YHU2tqd3ZfWi3EdQtbcJU1GHanU9Ag/3m6loai/Conh4VnNHGBnxB
IpoCZzvzp5gBVUSeiL5VZEAo5wDqdCapDqWP9ThazMfJBSL5HEGPVync4rq37H81pZIRdIlgSo3X
nyMeC4ME76KbT+pBeaqAGHMNE2WoASGk3OuDYXjhymMJEXjDBy4qDvkA3s/dgthPtV1gSZWinEYO
WT313+y/HCC8fVhTSqHjKDMglNYBjG7W4DA7WRqLVNhzRl3zTq5rcjqPTyDaXvsvT8lQdO94QmZ7
q/ziq755jJ/hX3gFxR1yua3b6eSZOPYXkdFB+e4pEmNWZ40o26PjNohrQ4aOsR26NkWxe98rwEpp
gM85c4jCnqtQs4cLNpDXO6LEFbuTlq9E7/UVbJiG1e+XjaveQpRWhTHniWMwdVzwyLn3eHGq7IIn
qEgF1IWZS/XpGC4eJAhOnX9vjpZCApwTcGctapTeS0arw1vplvUO4P+j2PACE4S23lv1IxneF7+T
0QLWha+YXOypstBkRojruSNgiPPv7kVwhRdqwwxg8D8lfdJeZLsGanjHRGIcx5U+zGy6GFEkmlYV
DiMrziByf55UMgVtJz60mWXN6oaKaUdianax2LhREMPAe9QX9qgI4KmLsEObFmjX8Zz+rRIGWo57
DYmLlNt/HIHU7i28qQp0fbR6JM2sGOkuDlFl4nd4+r8TX+ILOE4iNN9JQwwBQgGK1QJ8tmp5nMfx
r+4zZnS0P69ktJ8IS/6+KqFFhVNZaE08mKnzrDsBWyKG/uRkbC88ZkLnXARFppPiKUtA3shCWN5h
01hVwiLvhK/9ZaPIZ5DuoA9fRvXdEUM+NdBYaqD2oXWH2k7arUkDjPCwQDJJ6t6krAKMyHDraGDw
2bocV2wz8HbnXd5NXW/KuiDy5fgqnMO/5u9MeEiQ1JUyMcljYgv8JnOMoQj/nfLS+oTpWmqeK2E6
CouQ5aZMel2VHSAbqRMkFIaQihXxKsYWb3nvDIoYNOMovBxRe+q9fLRaR5ZlZ2aurrR/vafjt02K
6aC6t3bf6/AdtlJFSIWLFuFOKRkdUWF1X0FVyXcPtd6L2tCsWpW8i3sZXFCHNLMcJLdT6QiLFaUt
dHo7sMNz17h7FOt4DsFmApcsAe6+YYEMzck+jAbsCzkdh7MRbGJiP1SkZWfay77W8k3L69ua5dPO
uEAR6n0k0kYtzzu4KVOPJeTF1J7DQwg27Vz7lL9QHOYC2sBANUNlGgsQmpy0XvXQH9czakrQ8doR
bovDOI92rWgkCHjoBKbWsxKfHyqc5zAjO5wFkV39iWMQVPIUZKXvGA6YesF4qXk28U76VXHWeC9o
vjBVlvwBeWKB0eXpOFhmwwwBfpLWJNBcJgmFTYoQ8GdDZ8vNxNw3XQJPvyCuEahniF36RSH6P8AL
+FmFYZVI7a2kFF6h2y/+k/MpYIkGPSbOWLHCzx3I+QD6hMw2g6xdxVWD9O0uz1EuoQ1zf2J6h74H
GeiBpbsNWEpTOihHN6zsb1qlfj9Wuvb4QdE94QNGJcGwaaYbGAORO+3aPMrznxY7BhWJCeJutz/A
h+IHYKGMhoQ9VF/+N2rqlCrZhOP7w5yP7YYPllB83VnRhNJr+BL5o5aZKbJPPfu7aHMjDjsDyFwc
FgCv/Y486u2Ahw8Ooj9gioT1tkJz7iAITqzJVi918ajBcnKmLL8kGByPx1YRVnYgx1QnIpJibIaS
mCOzEEL6Cb1ng+kwXCdubN8FEzV1cBZMLSXqzsskLzScwCt8VFTRDPFKxohxUECZOKgI3rPxq6YR
ljneZ2NiJjIHusLgCsLtIt60IxMJlITq+v/QcXdgHp4M8wOl/BborCY8KZgUzUFJovhUKkPFVZbM
zUiLijVYAipkG4F9gL228xpG+lzm5tfJxNg+2kUlV+wKV7+ox8owtWvRwouWdGMcIdWOYrTjFODz
tNRwx1cOpOlKANgVdxFBf97AijJ4PHdi6H3lsnAGz/u2xXDqYg2kRRhUysWeHcRoTarZcruC2pXo
wsd5m3yKBdBrjkMNIbsnWkMY1jhK1fHwgA82YRD2kamo4q6IwVyE8YDY2+/6lpolI6KAOt3RkuFC
2y9SDzuEB+1Wr2mGvlw3Myy+eeddhp6dN7N1qO/eOppJmeozY5dFcBnSgmNPWMpA4QCENH0OjSRd
AFNObOVoNsMtlpueBSXgU5OjYOw26++GM9EI0LpfkLc4Pt1xQFmvE1Ta+AyRvxv6I8BrAC0fb1d4
eHXElPys1VUA88pzpPzVTS4+Jjx84HIO9gNlgp0CTAqFCRdZ8mEkjm/Wa6rEHfumQkLPXy6SwWQi
VnkFiezApWh1FOt/MUz3RGRIUr1RRd2i1OOyjL8yOz1nEhozApmffYPU0GIIqGCDQvbPk8/xvnhw
jqR2XvnoEmzrmkup3Z1WxL+6JRrN+0aKIzrvXaCHzpI7l1qDvniCg5ysNiNc1Y/OOHePBgEsI1yy
xgYIpp9bnXwFyacXJC/zVUrMc4rIcn7GDqRee8G30spT7+MhNEtA5NMP5OehEqBLgEeNOAOt0EWN
sexjaFq3xAN3Bma3f6HU1HwqzIHiGvR2+Z4BnJYsBsh26AO8RK6J/PizXFcZXoqwBxzqcj2GVpLZ
8A1tCqsUnDEi7X9M5Rj8rZSwueIFxFL74PbfSPTeKqxSWgXSHf5wBhfhOxEOFVQ7Nt+A/4kogFIm
cjhriQuKKWcNKJOeE70Q+XcLr9MRwc71EYZhu3ogSgljudpYxnDQxFHB6MJ85qsf8xUlw4bn8Uqy
FhmUccgqD+UDKc9S5ywtQcctjyTrvxJckpbPPBvmBF82pG2W86BdSW5cyxklLhnipBZkyOhQ4aR5
HuyN4AGMGvh+3KvlyuI7o3duspDuyUniCvU+VCZ/C0xx3U7R2XC38iKpihBkbE4+TjkOPLESwFIY
dErjl5vuYTR7Ffly1JBw4E+v91l7cH9Z6QyVLFigBbdqOd1v8FxmPjTZJYokw457ZcqVWqwENnVT
fGqEFUPytjAqWraluAB0aiD8atMZTrQvfHvuwFgXuVTIggEL03baTYJ7FpdQ+UmvuHMokSmsmNmP
LSjWOuCJBP5Un7PhmFLG/2KEO2BMpEugWCViUVKziFX8UYdORAIYyW3gsDfeMAe0U/ilRueBrwKj
coWGvyOIeEJGunlTLTjWudSMJ2ZeXppWEP6hNcCAxljOyh5WjFarHW5WXPSmA/j47rfdLLE4QwFs
p5lwm0QcmquYb9luOGGKKMabAVEklyjtRBUTKrRzNIcqbI8Tpznf01URUZPFwqwJuzG52d8R3Bf0
Amba+mN23GLJR9z9Rqop1A6wsLqTkggRA/+vNT0nUYMX7cqqCbtKV4z/a94HgfWYiJC0AQSUxo0j
trFWFFGA4YoVuDOLlslN/EFZXRpIIaVrITatkwIbPy6ZC/28WuLWco6LUCimLKgAV5RRVOQbSS6i
7EbFfIqxgz8b5/3Yunwoi9b5wl28l7m0JleqxWBiBtjSVU4LnYbikZsD+DySmxrHyb3LNJ8vEud3
7T5f7ajMK8SG9eiHAMXA5pKySMgJ8F8/YBiIw6hj7ezblxogXBOKEB29hq05D9rePQuk9tUc2vmH
yYfFvcnUN8iP3MTvxq5TcHYn1NIfMA7CRXUHg9nzePfs8okF4T2u7ZUsuFUG6E5SO1jg5dcS5NUm
Gmq/F4FuGGW0IjbKncafgdMvmmrbj525Khr4C3QwJk2NaIEuu2sjCE0RT0TlAVNFRNKYMaI6mV9U
Wh5C8gD8XrKShYfGw+zZhSUxdJZIVWThRAXplcYV1uGZioUEQYME6602232vmbCgPJAtDGyY2BVv
O+F9o7UkeF4c1Yv4NT3eE3ZUx7MRy8UpNuBMMR8ITDPafgA9fb3ynMZT2yP98qITfPEwD+BAmDLt
R7dKz5rjspuAa3Q1ku+6am0yr84LPHxMuEYQxodCwv1FAPxMBA/AGHFbaCgaCUBWc0Jy2/PUpZ+V
yzmX0kLOE9q56uPd7g7wM6w3EgxXw4ss8kj6QWbGOIf/nMH1U//tekdB7Sg5MVTYqmCwxyPKJefN
EzXpmPoVv+ewveCt5Drj7nEM+OyDxjEWlxRJpDgj15Md+pNYNoLDOm0Xg58RcyMCnouLP6IYOOL2
hUoFRgKTYm6V/gYOPikZ8ysyKFhyCQX901cwF0buo+6Cfhn4MLJER8LsZz56xQurl9TxkKXCCON0
qjZBuGIphhgnH3zZ6R02tEk73cL3ReOBE6QxtXNM2CtXOs1glkhKkzJWlpKpTXIWiTiUYesPOZrr
rIsZPDi0dGJqb1TRT1UWy0XGbYzvlrZonKG+f7M/rTvt2VdIbiSSwU2iMjT5HT5KbIEEGYLQGS+o
rh1wop5NNEDv13roQmU/CMAwfKlrUPzcE2ARuUcmo69+yqoZ7+Ksl2LZKLRvLnJShliNlaehDEZd
TDS372ljn+VqtrpZBbLtPi3ZVmy+c8Yj9ChC3hR1V1fsTS0mGnoBLObqS8hq9rc2k06Ikp9y5pDQ
xuyt7BPtXwQ0sda4Be0zG2GjzhNSbdbPYjeTlDX3lLx53gR5i340G2unth54XZACBQGym5OFO4Oc
yPVMydxigkzf5TbFg4Fc/Q0axevBv4hETs+iuq9E5MMxZT7thWi6oyjDtApMuDiCnufvw81z83ed
V7HrWuNd1nf9digtm91ySXbUDP4XwQamdeHpm2KUAqLXlFw2I10hJjQKk+Oo4c7EHkakXRGX2uud
8FjjhEfIevLC+YtJnn8y5n9zrJb6C1lzDBnx6Rhi0YHantsU3asWwjHdfBwKy45VbpjkzdwFmUf0
XD0/uMMI2omFdRy4NYinagd7jAvfdQwcjn+aEP/jjgVld4ph9+SE01kxlnf0md7IW9fJX3qVpiBI
pgrGBmfzWb04pw==
`protect end_protected
