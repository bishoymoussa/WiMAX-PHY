-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
k6KcjPvvsVAxO0oHNtBXCspPrWEfD4juufZyA1JA1m8ZnLI/D3ekrW+7dAPQgKwYVBvMh7zbjgpj
KDFpC+veWuDZd7lvWtB0hc+NUNhqv2ISx4sTHflTDDrRv0oJvDL+npd637Wda0IHVan0YllnDajn
4Rh40h6iDxd+jd4gOzUyg3+FIFS9d9mSWMjPNz+gLOJvUi835+zLiRDkLB6AdtvCljFgjqySadOq
Gsqsh7RDi0DEWOJxMxy+9XSjg005CCAizNFCazRqtnpy2/earTDIsl0vWXvOLzqkx9409VPpIFB0
GH+BFYMoxGP2UrVT+b7rE/Zx/CScgK2iy7Kp6Q==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 53376)
`protect data_block
Z3X6gz7LE0BCqfGCS3dyTJ5yjUdQpCW6lUv0CvorDVpsofwZQL7kJ8AWss+odBCIQyPa5fLXYR3Z
gRLhcLgoMNqnqMfYjIa1PoauCGbt54aCqAGRR5VQODkIE8CCpObmcl61SJ71Fy6zFCWzBxUfxO8u
MwwKWIlVhu57JJs6x062mJvGBM4yFAMHmeQHtYYijhHAo7Cg7nXADWrOqhsXkDacJlN69jSN64Cl
uVU7DZ2Klle/ADW/j9Gf/RZsl0vPZV03CAh0eetps8PJOZJ00r/lz/zFi+XsfIGbN7ZIIEWtwhTO
beVOYlyzdX+ZaQImCWAlyJaYgisJHp6U3He6elv1F9yome06R3oBtLQRgCW+fbKii1Tbq9yocXns
y0yj/FpSVR/Ou5oK/aY/TFWv9zvJQRiR81l91lpx5YZVGf0P6leG8jjca9+fI1Q3XVt7+JNlRPk3
N5dYbVbvtbOxGlrjKVhXV6CeFVmxjoYnFID/tJ3BU7mmmEYsCPguAFs58S/cb5pQKz9h5MxaBNoq
eE4lSuDJpjcp2wDxvv6bPet+DfBBnL7Eh7Ptg0nrBsxhfCWmHQeSjcwYON42mAkkDp7eERN0+VOf
pdWCDRY6tCZAfr6pbS6Oac4ILZNETcGeQ8cg3DVfxNzawK6P9ySVpb2HU3vjV2yWwp7jwDhEj8JU
KF4t5lYnxxXwyDudkh1E0vKzT/lxwWsqQ1OwySewFwVZrjUhXq+vD9dkO55EQB0Ywnz7mjIuQp6k
LhSQzaKLb1TVa4HXXA+I18rj4XPUovD1chF1WxMUKRQzDuLr/CxQ6Rbq7rDorlScem8nWcrXlEL3
4PPH7VIOSlIl93LLMfSB1U7JAnS7PiwwerdDCZwzS6Q30PFl/Rid+36SNHOn2wTmudY2JPr9drvC
g8vOrRj5zhPnGgAJN0/4yBiG8hJw/sbrtRDwjXGjJuJWL92dOQ7imsYQFIT88KeqFolPw04NB1Fv
lg9YkFNKvX5dWdQ7VkwEg8FmXUDKunoAbHQtI7zwvBVGUktEQMsMxN38eY3ZVVz2hQqBSXjY2Odv
Q92Gdvm+WyJl9rnZgvSawCwsxXffyvyTbOKiG0t+v3/Xz5q5Wbj9mIFf0wt43z8czqoy5b6jAvS1
dR4E1Xy19FvJVNvdYgf5rB72WWBV1sSWgWqV4r0WS620LKR3hCUhWzb9hSlrbOtfd9tmfmpML6mI
THd7v1VJvs8l2hl92MojN7OrX/VAwliHP6ykLPQHCrxWrv0tS0cio+Wd5Bpfz3ixb8gQTu/TvAD1
kv7OQIq8SWX7Wy2w07yLXjgoscykGzuXGbEJxGfZLGdbbpqdAVZYO96p96uHBBtzY1ZuBxKZCNLp
GY5nGxeDEgAxXQpJdoYKHc+dzpWu/EifUXQ9lWVHsv5gul2MWysiegEg+sE7OskHc98vRoMHOaIv
y6qizvBhZ4ass3w4esXqBbg8asUHnzSJy/obtlRR+dDfBW95ifqnnBgxAzqjXMj2dV+9jO3M2tjM
o1+3PpQzp8stq/jra0gU6FjKelTi7yU7wsUcnqVkWF0FFYqOgXmiiwK4UtBPndxd3KVGmTSX0co7
NnCf31TyaTmZLzS9LQgz+tZF8lRY48AyhLCCU1wgg3ymx+CpmPcm0DZFH7CKrpUQ0vkufRPH35yP
3STnMqlHsSYHx946YHbm8rlhNgupkbTyAwAkF5Y3MuJyFTbZ9bEVBLiAga8GT/O23V3qpuVvEqgD
Pp/cN2dONRr4vUcQxQChM45OevLtQsaA387TjypDxDDk0yAGVlJqnCm1nKrIJyhpPolCX/rJY32v
LfuyL/tiJAY20zA1+3ssz5ny+Bqkb5vraSOevZ/E3HpXJL0Qn3WXWhmGdVkJgGHlh66P+pnMDOb9
E3CS21wi4LAcfwT2wHjhg8Nqx4yV13zTIjkoLvH/jTOeVkmqgPAg0cZ9Xvoz/DmN1HAFauh/yneP
LUWj9YFVefWuRtRzhGXH1ROMrvT565pE4cC5V8cgw2CsnjobOwT/3Gu1CXifx/2c1ieAAWAu172T
TPVRwey9v2PRKOa5TMqEe1+R2NcMJMWkc+lwpVhHrZ2Sdj079eVYKxOp2DcrF/JOsJQXlvMBRr46
uhc4noOx3GddB+GKciS36SzoIOtF+2JSv31OheN8dk/ESjcYb+N7Iz0K3mcwWLftTo4BlED+orHw
kUNi79X5kernus6lc/a1RpZRZfoqhOTpsjo5Rns17UoL1NMgwKVAu/vQCR722xOOqPVV2MbClnMs
P2bFxFx6LRHlq39eoF1D2aRPxdZbVFjHJ4PJNYUN7qhybRxDlMf9F/SuIAUcUwwEXqCp1MGkFydb
c0lNtC8R56MyDqJaGmHI0DeC8n90xkyyV7PzPrqGY1L7HWa+VDazox2HbeKsCB+MtHav6+BQxnQv
tKwPwH/NqqUZedRXZbtxct+NatNthct7S2mkVJrTGA7z7PNiv1k3muXD76JNs3LoTbl0srXySV2O
rR+2S8alU9KWRrlLdoQ0ztAcPS93R1qgUKJl7mpJa5XSDhQiS2F9nJraISVpFWURS/KBqhD6hTfG
aIijM80FlTbt+oRnoML9R+iHwj6kFMDWb6b5EOxOFVgqYWRasXWUizWteOYXmZ7OmLNpTnAS+CLq
zYhGHO5OXcFCVgYPR296Vta6HOcjtlkIJZk6MUEbFzT7gDGPoYyHXplUrOr6s6Fr+w0+1r7kUFOS
gP3UxBfOoJlIHIVMwuIwGBBveigk8IO1WgH8XeQv3+IxF2DpBtZVHppAKS1tfOHaaXq4ulOKYwMc
fFgABp/HGk3hMqRz1omHXWnqZ5U283XQWIbZCc8/VB+3K3sS9Evmh6WuZ0fewrqoMzs1wbco0hvk
DAdtRH7EYEwPAKhU52MkQNDOVIoPxeDY0tRxUbG5tL7LeC27ceuRE/W8GOnFgzV5mGCK6cJdDmwK
2A50HLIuu/Ac8odyvJUgFKlhrCJLyCaHR5f7leTMJuEqZKgcNZRJ2CS1rL/2AxU+wPUP8Wguob1X
0dWzG1m3L3nF74kzulS995/DuSBNIIoSrtqMnHcOzFTBfBkzKVIQ2bpJ7sR2KMDHuoJGMkw3GJZw
EbjAmgaVWTGV7+51zAHEIIHThzaNqe/CcQw4Bmbm9CC9Z5xx/hm8UvR6ZhGg/NvfgZ1xWkqLpp1K
aMuY3dYGqusxq61irN4tGZa+0ySV4BAfG0RKp0xNczGiMayi2TGXtwkNOvSb/2AP6hkWIuSrl5+I
SWVeqlmbot0e7UvQFxQHn7UES4td3tFQZpzL1qNNXcke5+hnCP53GOQOIQdITTIhw9IXCMBhM+BO
YIi6R73ct9ugytpDZF2ihs3Bi8vVJ6k0pEVCPNfoQ2C4uBahBzNDl255VT7wSoDaXeaMx/HUYhYK
fYARP0aeyc7hHBmjdrjAIYBjJvf7mABMiGOcL7VDkohxPo6szsJxTAIBe8zxqXS2aWVyUJSm8o5p
whnFMJ88y3EhgVOP7u4+oOxgJuzj6ZrJ0J8hr/GIvojjbGeIC9lHd5v//vMt/nedC6ehH8fu95bz
IyVj6CRNFUivjm9VONnHxhGVrrr4lVTcSaPDdoP4WAtocTnMMJDTMgS23ZkLWfMDDmyOxVFBiT8m
9Dwscg6dSy3GFsLUlPTlJkQw6eCXFw6E8FCeX/Zhf6fn4Dn5r3Dzy4nOIGwa2RExmDDg9UyAh+XJ
BrhvWLIad4JqmAka23TWw6+Et2iiWAHO2dNvWMSzaPRu8uqxZpDIVIYyTRpitEUQQmEadJPEv0eZ
M3KA0aSyIXgmjp+jw/pkcHCmNbcAJAObTopFZKa5XTC7WJRA0CTO2vVCB8wZfDTMpUw9/SPJdvCY
xcRkjl/oFe+nXBBxrA1ZNABDhRohTuUKJk1gI7ybhqMRjc5EyWjhozCd3i0mLQ5FU5TRWI3ZsKMc
qCZAMVFdBJgc1uEqMQep2rK4uhduirsEAkgBy6yJ9acOj7Gk+efho5CvyLkG6CqeDoYEiXRuXzCt
JmzVNPbksH6j7rElcTw6xIzeWy1IgYCSeWwJ0nDBxriyivhLmgO5ZTfv1Su7vgDErQRYkgWE4OP5
OWKv5aj4bVwSSaZj9MFRCCEbRUSCO6txGcQ3y3DwdgaEoGwtBrKqamp463dLweJmxRIyEWYdgQs0
oU7yaFZQsO5v67dCnHzE1u2a1f0rzBaA8CI+AaeDnkiAUqBTglQyClkJ7h8y+JoJ+/lottbGQ3bj
gW/k0C6PPFix76fpGlGKnK+sq94Ty65b3TToPRT04ymFS2ogfjklPstJqU+r+dTEP8Z2u5Obkmz8
DnxxKsoZ8uFzAzStKRm185/3brMJh9dAf9QJIHNXf/g2XL0myagQy+MzbU8l5i3TnvatZlF/SyLO
ZxCw/u3AiB7NADUIYbhEyvu08HcabSAYg7pEHDKXmAbm+tP+QKtdPHE1qKn1Il6tn5nSSMJkUGti
vGFZuAunUbdwLM5nXCUGpWlNytLDqbmxZ7QV/mH8AsfpB7GAQ2IgZdNdklpI4SKg8csSF+ZL6QcI
7pTMtY94OLafTuhXgW532fbL/thcUPjouh+S2Kmq7z9NLfjaZvMHWeGDQ64rebzdmq+xDFuNtJSD
vCPWC5gWUNqnIXADVKZppZGOgvT8ecueML8fAQqnSeJ5JUUzkMQdAqfbQ0rnCeJ75WSFkp2cOBO3
IdU5zKcgS70qBIw99P5WVEcD45tWt4sIFlcY5mqujD4SkIJxh3d/hmwTk4OGLrlyMmCmkhtPnMsG
21L1sIXQKHEtoRqDUGQ8HYHovuYpuTZWmYdaA/14NFFzjknxkiWkmQPR3og0KCVHKA33Rg60aNEF
VOOLYfpR10Y9Gmh/QQsKQkSNwTnIeCUux7t2L+wkDhnDnYNyGlS7Unqx5RqZPloD5We61wQbB0fw
CNq7IsG5mVeVy1bwhjjMnUylk07Tk9WbMalJ1oY3RujE6+7KJiCndaVfkDYXBkr/5yoMz/SzUa0X
V8gImI6MXsnsrXTTRMBNeFy6lI32v+uSWCQLccZgbF2Akfy++R/7pHhmebxhuiD0vty0QWsK1oPD
TRAm5NFka8BknWmRnFOLqEzU80UQBVrMkx6swgZSMTXryg70C3uR75DNDUJVML5Kk/+qGVSwB9mp
CKbmhsY64p2Gf3xqbhpw5wIgVs9DOTVnvPaPwuYggvP4P6zrTcC/G5vff7O8b4oPg8o6RxRhoZwd
2WNpxOFRJs3BEKzFL3aYII1CbD9jMMVsaSTrwAG9x/C0iWIcBV1mpAvbHiIvYr1Gogxmi5U/ladU
TxZyOO8YTqi+HPl1xrUgx2qsT5wFbvk2WBhc98/qFw22IUGxzjuB8myGUdDP/quPtoxCz30RAljL
TURSku5pYJ+mpUfyVDtxKPdizTjU4p36QvEeHAAagtvE89HMp2wr+zontaZCZExJALRoe6XWmOT3
SUD8k2I4DieC/Vuc3lHUCatfxeSaNVY3ezrG41ds4VH+gIzDa4FuaTzYftLBIAyOwfSJmf3lHnMz
kwbVn4IkoyzRo/LYfciRddXtzLXv+womqMGTgVDV5B8W6ZU6Za/3vAF6yTwqO5A1ptO0icpm0spW
23JYYhUru2JUMg0b02XjZiv3kvtfgoC+6MCcjfdgEAhZLeqe2WWRSo5R3myjqZ21v4p60kDLMQMC
EaTWP7Aw6pII/PS54fbed2v7xQ7vHMWKByVuD1N6A6RQCxToT6pJmWLfkcSW7RY8297oe/3W4JWt
CYqAIKEMNr+ETDdWG+nDX6t476lOs60rOjaJmqOmBxc3iSYBD+zCLStME7vBJxAzoogMMmmhjCck
+hfWI9YsJB4OVHJzrpLdqv/UoULX9CgPx4dI8/qPZvj3KUfzCnLCE5OwaDigj3ltZUGCbW2C7cY9
f1AzRJdEukiMr5nLCOl5tl1AqKmgSThm3QTYqCKPQ7sFMujm9BtJXdlnITYkVYCvhWd56R4cnRvt
2eoYO0BghoWr1B/UBbr6p46xHj+qiWODlEYwVHuWCWCxQ6Dx5VJcgFaSo9/dL6o4R5FHMn5MMil5
YeBTmE90Ml+zKkqVQH4CvNNDwjZoPVk0PRQ9FafI6lfIPWsSjxiwXUwxXPaCmQ7xUt5qXX4JQevK
JdyOWTNdwYny9zUHAYNQNR0ZIbSJe5WJ4eylTAEEGKY1kI0mX0mflLROMH7TtiEsUaLkzzSMnm4b
cqQRgYu8I/abBeFb/3ZoTht9zTpEwknDVv4uvmIIWOWD24SxDlsQw2tvDZeJDPvZtTr2mOKkvjLv
hhJ/Mq+qCEzeYOdQSA9V/lXPrzMeIMJ+Dv4kNd1y9wDaxiPGnIAtcPqXrTlq/4EIu1J0sS7dfZtV
EwOtkXzCI0vVHiA0OGdTR+tsAeqTR3t0NfbWUakQiIL/LSrlijzZ/7pUSjN5iRRrReksp4b6kgqU
XyMKh7y35y2QiXURJN+e2JEyjuLXLYpwJouXG6xX2hdlgc5Z0KiNuDVvAMr8pWj6en4P/laCazMW
pZiMt0+YPEM/1QCbJVqtNqXo26VRcZvp8kg+nKxzmCwcVjqEmK/L4v8IoLtjHX7Zet9jUpcTaiRo
wsuzqbYT8XSTsOw5HADQ4jDhpCTseuKVy+HApdYPgxazTghcjHDGpKnVzAIJ1dYNvvwvhSpg14Nf
jgkT0YKRqcA/XV+goWvGfWhCpsFwGzFKW+/lgAtpB0AaXIj9Sv+VlZ7iY9Ma9BG9B6AvpZPhIUyM
GFb6wLG56z9Ey47hlWcNbmHCibQW2NY+aY73Av+jQ7f7zymkAWdgKexIQLGFOX4eGKj8ZkvpE0/O
xfSJnzGHyRY4s2El5pEkN6OPtoZuXthWdy9ZlTjeC3DI1Kp831C2L1vukYgIZBEelVQTR6keriuQ
rMoJyPSYUt72Lp1Fg/k9RlNIFwx0OB+0ajdXWNEJYCCjvT4Yye0EFWoLqd7I5XeNq5p2P+FDuMXI
XXZwLy39TZ1USRhoMwd08bWfDd/giUf6pwOCs1gUWRRkpiixAvsB7B6rhNDVONF2OVvrEKA4aoFc
TqAp4gSEp+u4km9XFhZK17RKLdWvQSfAJr2P1QDuZoybEB9Cgz6zX2Ei3EwHvb3TAwFUqChJPnmJ
RNoHKgo90QZNLz8ytFLYdOz7VsuMrilz5/E+HjzicsddHtH0SfRz4jo855dB+64zvDkiIkeeb49r
TMf7R+Txy/2C7p1B/4WpyDyI1pol5yVowOph5ysAdawuIYY7BfGT+ccfG5KwzxXEG86N7JlHPt5b
NxznJVo7e3MEwJbTG8wfoG/41UwKyAKO5YJ8chjsDdylGlqVetDTI1az/N8V7JPaw41c5jy1xn8Y
ZJfkD7sMkbpcfwioytUDcXutToAW9DY39Z33k7/IqilT7nX2as+IxKQt/wpYctjQO66iy1YHzjKw
UKGEXwTpVz28q9LPrqznHe75xbCv1eLthgaQR4aaX87eCzdVOiIDgmOLpFoQy6GcYiMiuYAG4rZ4
hgSTlI6iuc4KpuXDVlRuMmw9mrARXZYUPhGr60SjDbIA8BK36WTqh84DZcMgfbxb9lW7ibBdKXaW
haA0jHHuJcqe7xEGCaZlqqBvavColWCnliu1TXRBl0mVeinrU5x/cvVEYreARowM2NRkw+DjlRBl
eIbb09VsvH/BZGtBjTdH37ati462h8Jy4fykMMZrzjiPG7lIsjLsT3W+XUDsE02rGr52iALBvicp
dghslmEUp3bXy9XQRp7FqExhm4uLsP5GkwBK8+aySiaGp+LPkWSRmZSRMF8nI8mOcpP9Bg6/xFuS
y6INynPIvJRBSWmiTvHf+qhyEoe5Jkx5ftKTzVZzXL4mW5AZVyTaY9EkXXQyiPr9FAMJQk8JHiFA
UqIlPva1Zdsy4ZnDA6Hwy5D8GpW3e3FBt//MaF/SqWPPYMVnSQpgEMQKQP8arf4HRFSp0jOpD4E7
cyIXCKofoy8u0i5LfbdTh4pXDQAz+kR47obSmk6xvvHMu6k4vg2ZXX/li0qy7RhB47YvlrZ2i8JY
3F4dyd3hSp4Pmey0ZpfySr/OXI+m/7yLZzycNxHd00aOuysHUZXRWBMEGVKt7ucy73pNktZtqABj
c35zvW0hgFnj6Mkj8PHhsFWpj6TswfhdeQiRMsdOYyd7aRb4yFm+y7894pqR0Ac1P6UAtQXRy4lz
FXMKlw1YYP3jFTXcQk8lhzHyew9+yZwlNiLJ3Xxw7OUQePI1qYUNXCV5bPoTBJONE5eIOSxWpXRP
kmKLWN2563LjFawlKSFPzgBybDy2gfsah4PseV4Q3px5M9ChMxfwTTKTGEVQkQN62bPBncr4sFHz
plz6RJkzn2P0sBRDY7AxXDgWT3hkpyNm8iTg/Wdpot1nrJp4gWP+o0n5GigUK7apAziqkdD9us4o
6enmgRs2WRi60BnNZyFkocX7tnlUrDtphrUo5laRmJApnWlF5pwx6O2I/EypLQvoGdzdF9tFM/J5
/XWtr3EsVj8jnGAe4u9E7Fy+ziQIxCK4ijh6ztxoBtnVzJ/vs++7na2lOBBPHvZ/ab49vOFG+UXl
vPf6MO3ibXnIekPoB8O5LXrgHSbO2vI1vZ173UQlyTy/UsWo9auHlf5GKOS+Hl9CmTs1jg1ZOLBy
6scKCePEAU66RGnsY31Rw7sc2sGtjQoKWx5uaZ4+c1vCmteE4n6ZYKoqPdEH+mN4LVp6A3FlSGlU
ufS3mfEDEUD459s9LDKo69UxhbZOHVxLVKiWHcUOqUboh1AhxRIy9Uqa880nvJcyT9z/y03pKgZd
WpjiJ/G0Zo9GDS4d1/Qk+46yRFMsXGlR6cMed+gugLI7rV/a5UvmotX5F4bWWosVUaVIknua+Hs0
awXLWPW6M85WZupAPHcGoRhQUjTrmCl2+5OZXKrbizorI/Y703FDGqRKrrE5AiR7kLbyzaGqX6d1
hJJf479d30Lwf332Lt38iGoME82mg/EIT9xvzQakJQ8nVjnazJJoRyxaiNGDjqV4iiXXXCh0yLwG
7OLqyTImnjzejo9qgDj/YbaQTQEx28k/LvEnMa8q8IBLZTB1miJM0mDB9birolL6RZsoMNUuY7sX
T28buZSPAjfAJwW07M9p6f8Rl+ZICmw98Mmtc3x8AL/nBm5BtU4WwhSlLmQd3iQm9N4mdpyROdlH
JG/bvDJFIlh6vZ9DHIzyicm2rVerXytlF5D4BtzFWXrk5+BJhomXCk8MzyZQZI0u1WVVYLyWtsZF
Du99XfbHYfMv6hDqLpE+ufrEle17K51SK6xv16jB1ezpVVVJspcgEob1LccbGaPFFlsa2slydQ+W
aaO94D6Is7UCIditkKRi9VNA+1OyKisO8xFjB6UrqwsHBvqSbQtbmwN+Ebu61G9WNUsLoVs2NWwP
PyEcGXP3GIeaqkMjn0S+f6LcTGuMJiwKqNfwwv6TDBO9qGgttEONciD1ECvAepHvgwbfiXO+UfVS
MCgs03hhZolQCjoUtzJVIkctX94AB03iktLdGedlkAm1DJgZZ/41Ywo21GHROlShc1WUGE0fXCKt
T3QtiwrMYa3EwNRS2vjlxIAGsV+psHUO35MgX/I10PBIohXunPqjypATOvl1EDe+h6vo0g7PU7Fk
CJfUKJdX15eOTSk54HHK76jl05Vp/fIH0SACdso0bIcnHAs5j7Tl1Ume107gdD6t314UVUUCvjJ0
48FCtRWxrXsmWQtLQRdoeWlEbjx0lgvsHP8+JvQInOsVbLdgZ6isP5Xhm5UOOtizf0i0ACienNTr
KRTVBSKhF+1iOdcfCyYCvTViZKZP8Yex4Y2MBderrJnEG5vzhqEWkrRKU9aI3ZMeHuRkJBvT+M5A
/FFC3dt3AlJ7UTzDa652SOOw1o8PsiXupVCSnZbu2NSMAR3nFH/Q5PRjw0xXLHXrtp2sZJQ2sFNZ
iIOtb9LpoZPtNlzopwipCfUzkhvlT9JBq1ktgdE6kjf0PqxyS0+SHDjgJJwl7xfeAFy5ITbxRYev
w5vEPMKjUXvuTsr4gILnLAmf70qBoqaOarXoNdMSYtm7010E2iNU/1a2RjdWCbQMP2+4QAbF44lu
OtcdxwZnZIcGqPZ9X1Tpmid3hboKayw4Rw1nX8Tu8CDrKaFpIIFTb+svCIntUfmoyw/0t0qfzsFb
6UbmnHIGwIDvZUj4tNmStGtY8nn1Js3cwTGmyoeRCUGj3Z9b8izABTTY81Gjwpf6ry+SARbGJl4S
J77YrxmV1XERR9+v57FJAWZJ/NNKhnAbKhwr0FWu2XAEf9f5x6DqDkm97WzmvjLGQXENqlC6zXp6
FYhRqbZvy00cwMUpti9GZLtNkJixUrJ6tym2vP9GTdWjkUp2zrCUXNe9FxgTOL1pB8bpdqKZTc3F
luutd3YZdMpfeHlTqRWEbwEbxJcGcdiWA89MgoO0aesybh0RU7sETb6/46SX0cn6pt2cx0fkUAsL
4bi8zGnY7uRMBfDVTiNeUWt1PIKylzE26ECzd83plGIYU4kSd0RMnIaZFFuHkxWXgaUmyriettSA
UV3PbKQSBESrnDxPvRz7E+IFwslkqGEsg1fbMhA3QRjDKyXCvNkLuJDz1FSn7AOz4JA7Dao5hcgj
oAAK1LpLDWGHcD9ZmvtunF+gQxZ21XHMU3KTxl3gBGyDzE10ocF+GGxcWD6lH7VE0ukb75eNI9NZ
hzxLiLre3T74eBZQVZxB1AVEy2XtEpSEKxTJvQ41opJEa87mSv5xppyJPgAvEg5X5sUhAnBp4SQH
9TG6Ffca4FXqgLbaDMugu6Bac7TYjloJG6klZjnl3a/L9xQUQm8fSRyxA0Z4y2jyKD8t9cXEzNzd
V1f9iL4D8TlnTkqr7Q+l5Ufx8dkTAK/0uD5fXi1aM6vrMfTVRclU3Dc/m87SgpZeEAF21dx3wWTg
gRRDBE7K6m1Lj/fMzeN4QTwtwq4tbHPv7bB8ZI73HKYWA3z0NMlG7kUVT6DODMdYo8aPhjwsYlI9
uf4e6f5GEHC0dEQukaK18Y2Q9/9tIzcljXe0ICPfgrvw3+GdZYEGTbQC9kC+/DrmLUNqE9SOZXGP
kt68R8c9yCl5YyB2/g6ZwzgsmDm+E/8ZOc3mn9UOotIDyQwFKoHxE+6o8uZCNmG07wfD4QdLzobb
JmZ1dsJr5yBS9SwvRZTqzYFMnMbcQ68Dq0/CCIVYv8JM7TNIvzv7njLFBqLCm+jEE2bTt2ozD7V9
1CQhK2NPIzXA6ZN1sjNv459+RsJ6Us8WMMHAaWHE7b+mhdxFK4LeDI0Jor9XNzwUxe3O71HWr+ex
vIlTd0y50Jazx4KDwDbQKvubEcEzsUogiY35AG1gRkUqWMuGIofJxnRI4PXlz/qyQYAcsNaxCLGn
yi1GpUXY/wDbHF/ym5cXpYilbsRYz4BAMZsV9/ubNnCvCK9zk4CtomN9pdr1S3Fz8U7FHVgucLXs
C5TpJyojEKVC54apZFzx74nbAdNfMa2iyhu4BWgAKywSytpu9ACMe4IFoZAiCnDTZW91XKbr1r+i
irgZHY5K4dttCa9SvV7olLbamJFxmaP2ht2HB8CxJ9V7nryhOZ8DbR5BAyBut/CQRpTrB2lIoTz2
hREb6QPJhMhl+9lcaiEnV67922s+T4ov4gaEMJltPJ2bxVbNPw5TJdL1e4zDhGZWJ1Zstf/VRczL
j5Hat0wY1oQ9/1h6rtD5eqdh4Az1So6KkWs1yFQpfNFW7UsLAapbP7Vn9ioiTu+lvnbyn1i6Q8Uf
P6mEMOm2mT7zDp3HKzkp5jJ529bCivXmOs4xyWzGClHSwV8Pc1IQBBw9yU1KO8OWBYpZTIXniJ/5
W8avGrVWGIcrFVp6c8m9gIHdmHRPG09cTqB+O4lQUgjd/Z8pWgH4M9BrG8x7iN0fRyVWvEhEoe/3
fvuf8R094bFP1bIhkRxXhP5NWKpyI8oDH3UIpw8wVXGBczJzClHOOboJtc7F3F6g+aXP85qofAXf
EC1ZBpjclZNs94SS/eoR7ouDqXSw+yT0MkMywTZBZVw0FZsrVuCjtps8IKl32WJBnP1++F2Dhr5k
4blEDrSqhDfbdSS1ySVOmyqenXqipZbOjNSnj264DG0gtQogKgqmWqJ4q5BSfNyy8eSDfg7ArYr6
9ZcWQF5Ko5hA7onlGeuTlnhW0lLRUW88Mw0Mj+oai0Ycxu4EaatUX1FL26XJ6oem+EQUF7MpYynr
2DJL6XhmDYd53Zr15aQbh6EPgghMbmWe1CpTZCd/2ZwNExaAu7rRdppxo63AMezdhsVfTw5KM5mp
aggYJLwrUhS1uTQ8QMCrWEtWZz8hvOR4YVqzGec0rsA9lZk3s5tET7TKwTu8Vlp+D2UBYBpgZ3FN
O/ddbLS7sTsLyBEqyXbkKvrjaLSQ8IZYo3SLCdGvdCLhnPgRiPBRc0RHObNH2FwEDbzKh830ACSn
pq42JgDoKyryKbk0/c7L1E3d0LL0UZAyDRDwGQGrzkE1fHUlM/v1bp0dYgyRumQ7trZdotMKrEgZ
tevlWgFrfxFzyeGL6NKwMW20NBsttbV580wa46MmudtifQPB0redj+i7Bgov8ZtQ51ceM3IrPHfQ
5H+iHI1k5sAHnwBMTqnnvGTAeGNM4jPFgOilp6F73eSln7ev77jTeYMf/5hgoTjuNe8AZBr772ZM
7lHhVLx+nAALpYd3P2ZZUBHrMDjuFb9tR1S3cjNSbPiSDQsyjWgQ9eyPDNLuTP4aCBwhMF2fdRev
OxdYAH79gsN8/7KEwwxaN0q2aZY64P8lLbxv55V0pRTFb4XuOzLWiTui9yfVoYyqeQqviHQFo6Ex
rwkL3BkMb2sMX+IXOOUzg732L9TYw9IeJQ8QDyxavAjuOaqIMjwfevkLgxqXYdVcQKRjRpRzr43D
vWCGLlfttgedxUOi7HKdOjIJXu5RLm/Ceg4TNqXWaGvq3GNE/DXp5mYQlLDshglKiOi5w1h9exjX
eesadbZz/6NoY1LqtoBFgtbfH/QVFdjGGHgGaMTn3pAP3/2MdeACSl2HUoOjgQOgQvMelQrXG4QN
j+mC5jbuNDKivELByqIHtpxrI8/3x1gXSG14oI3ZuZB/HJNOsCBQ6ZPx/kE/H6uWVKirDj7sJzt3
crriDEpQok+oPYncaheWB4AZHYDMPckLiu0ai20L3ULXjHJiQUWHqzEY9IiwMfJfSGPMMnUl/z22
tzxWMDEMtBH7Hm7hFPrSgFAB5v4PwNZjg2SSRenLNP14bHDYacRc3KDq7FvolbqaNUmeRRcSn6Ik
mtIPiNQJLFwQA8x0Cl+OP18tpDteZUsd6Rf14JIGtL/6F8xNj6XsXtnP8MFU49wk/yopRy2C6dI7
JqW5HSj0EEFzimKjPJIakJhyGleh98b3206nBP6L3QKiaepBi2/6TCDdsjhtSxCI8nn7+EyGnv3x
CCGabDwgyft8KfNeRaNeKplxgVK5CUQ6//ci4iYpbMUquhN1/UMx5tUjCLT/MBX3HOTxB++dJ2PS
Iy7QpPiZeNByehdmoJxlsc9Fg4v+TVHT4jKR5iO6ITJRlIayxRH8007cEGAkCEJbpD1K+JEE3nQe
o9UE8GguMpBRJzL2RFs7FrPAS9Oa7cCRxVwuJvW3Jn0XyDOid7LLDutZ1TeHvP0fleorRGCbZTjF
5yOrxsBDQAvtZX6Dtzp5wIFqZf7ZJU7fT+HjfIf0xGU8Pm9064nZIjXN3pPQRczvq09JDgbeG8dF
Hy7R37k4uLDQX1airi9SVFjdLZ7jUgmacvsNCEgwAnqQwdut/2zxdI6NnY1OZC50PZtcHNZyVc6U
XiiQxfqehsyPPBYY/yBnL3ya963OaRu0WksyxxsnievkXN+qZptnP5qPxUII0NlNB82DYbY6fivR
Vrnx7+oZM5a1QHeEC7xk7hz9bw4083NlPnEl41sEv+aKFRVCyfbylWOiCnLjjhGQ2LKgxWE1hRpm
AdN+T/yg21SgzK9R72h14AOtZh0ku1lc1i/tTmJ70qte2k08Edl2WB8quNuIfxxl7JLme71k+F8p
iQkxXQp9TyR3KjQsOR/4+D1xvoRV8dkiCgAptT+dgdHIIu0RuQWgDgB3nm+VkPx6HNIw99kG3OFb
pVzrKaBhiSvYUHIv+PHBIYODqSoCZQMsq2hHPxIbCzouzVPQwDPct8DcJ6mMrNqLDCCv5SBdTddx
mvTXzilwBdFiMYKatPesK75qMExkIXVUHXLC99meAPv0SjR0wHX/6Q1UOJ4mkWypeykjVmZ9MD6s
CdwxTV4zS6/WT3N/iEMBOMOzlPvjtTUkYu8zTXi84ea3p2geRiMul5vuJL7/jMA5kLVGyx+DbPvY
2FfR0rjQjF8mDak5Zwxdmk2+9xNxepZRIt1eW4W91FeQ7mvvjikmkZR7HnC+bNaiaR8VTZFWEOYt
CMwhEh9jHLAe7iLxaMFca70RdWBOIXRZuCp0zumBHhyMKrr9JfbIR9gHcK01CWfoTblvMm6vmq98
sZqDrtajflNt4+5/7FTzR6P0Qd1euCK31Dy3c4ozfxuWfrfuVFjX3nl4iSnxxG8Mam2Max7K5FAS
K5TalwM6LwPIhn75ATjT1CoGLrgjy7wY1SuenZnlRUVOIHZBzZuD4DkD6EXvtIHnrI7b7sjJMviG
48SlIHk4yBfl7MbiKbOiXd62VEX6rkFoF9kPjB4pjRccLT4yzCTCLgfQi6blUtlJDjMQyPUmqzSA
rh79bW+NcQ/py81ASHZKaqcGL1eutId9Kpjd3DDVO+UGMwQU7B2FMU7tYfu/SHwut7eb1XEcMDyG
e9PGI3FDfgUKYTRJeU6TC8uJly4UDsnmAz2bwWjGriQwcQYXz6I31uppH1nbx1iigfls3uJ/bkh1
lXlfQE7iAjl4jW9OACegpLw9pek6LeySj305YPFwdqw5gBqU38X6lgaV5+05q293S4dSZ7vOt/2Y
cfqU4UFQfse7aQ8KCYjF0b7e0KHyQKzpLju+RvRTxCUQfOP1AwS1VR6PcTTepU+nuEd5HJdkHY6k
mabC2EKazUUtGLMQ4kDTkI4n5zogFCdnATGc/V8jtsTFT+Jnpo28stQqlUzh78VVqMBYG6LNNOCW
3rzBU7q+XOAyVFeOKA6W/AeuCfurxsaYS7MyKtx4abbi9SDy6ouWwlQWW9s2MRXrZYsMbU4h3VUa
7Yep4OHJxdVXWBY74D1p4lvLAubYcGl3Uo2lf/QMp1fzAew1XZNRBrsOjsHIDgT1+lwOrcSyv1WW
4KgrS76DzYbxKPSFpbo+R0vi13eOTaXdUoFE1D67YdiKhRs9gKH4GSfITiJiRcYjwaWElg2fLVN/
SCeFzS5xFqb14CckYPy5Ynz5Jml4F5ZT2a+T8Qx/equs3dFL2qsKijM+HGDk4pcJkGlMUxzpsnuF
vXsvVvqByW92nlt1DprpC5/RfLEfdxG95d1rUcpZYhuTejvLw5I0wXf4le4ebZc7MCjd+qOJtmqz
5bikykKIwsWa3Pfd1tSSN0mWucfeo1t6aM0YEws2q7ucXL79EgeIlnBKVDTFVOSxfBn0gEatlwrq
kqDCfYP7VN86/C+0q9gmOITbgo0/AnPpx+VqU+pxFcZwiH07WeWEkzpYNwdmC4sJv8EL4CevStBI
a4KA1+XBXqvBN/YCPzaa3X7DvCD7xqscqi2B67zC4qWgwwWegADB1dZNK0cFzKD/3hCpugdOt4YK
vpkrVnITQYb2OotDPOUWhY+eA9X8tGCKRgBH/xcuxDHwSLAwtw5SooZQU8JFahQt2P3mIDlJN0Sd
RjQaVaRDdWU44zXDHACIXkbSWuz5cXFuwaYJPZMGkICAHusskRH85BBcThALvlaGJKsRRT1CeaAq
wPoIpdM7RsMHwpNdIM0EjpAL9OFc8NT1gvXK3Ziugr9tNrKnPb8IXEG/76R+yOooawxtR5lsCVWj
qklc0J0LoeMgn+nB8PZIJLLHD8ho9ayLQcmQdxzMVev0BLNKYXT5YtOSmLXvdlsFo692c5HzBkfr
Wf0+cGe9S8poaugg15Xwj+uYOVrvKUfH6fEbQiCYvdYmWze+XI5ODO+k7HhNl2AhAGQ1i1di2SM8
iEqgc6mFjNXDf7uw1teywyWqT59dRxpCF20FLfV4iNqJiwxynBLlNypKIvLHYg2TZNDqLZTFXr3t
APE6HAPcK4V7oe95BRBK+Xhx0mTDZIEukO+czs0M70SzUG/bw7NlhxIVreT9y1Cu1faRYQvVuFgN
4spc2rQ7UBZFHXCooirSs5dcM5EYS/sf+G4yLKoJUil9skRxnyH/oexugx4ZvHIeVEL2AuRhzJt+
krcB78aVf9/kryt5FVOfwYxtfu771bNkHg2GcoWWMvL5cPSNnO3DcH/kTqtTqyMMLp6QnNof3JUB
v6cVV+gNU3XPYcBqLG2PS1PF4GzUTvPEsG6lQH+G8yJc+MiBOFcbh6XktxVTDxJ5yifp8cYl3/Kd
tvg5C2hJSKPhJY3ONCZ03SoQ69FBWnkK/PmgyXryDid/L/uV3Md0+64eZE39VcIn420AIT/m8+eT
xPDkvp4VGRr0JxctefH9TzKD31uFgTEOGG7Xt+r5EnfXYwewJL3pOH0LoZZH0rJiZKULpanVnTR+
fJc3Z5VrImKIDMebpFsu2y7Wv436EusLw+31KjFnz2B2SQfUjm85IUNM6jysNpCgJ7aTwy4bEbJp
EEg5JOc03oiBi4TvH3CdjBu7Ukt1qLrrF6iFL5S4eQw7wBYhA/zWKm5s36HffxtG8SGnzxxALWmb
/INTi85kmloSeFE2V+vRa1g4jh0GYLyH2/efHhZlQLBOD0fsxFCVFmnKwV0g1OamqMaV/XbD0OJK
g5bd3ZEhVr9kY69A/p+tABoCT5L5lqH7zprz/vw+HnJOZiiVYfSv+jmJpU+YsxZ6F38fzUJ+q58K
eSg5Tvx1agOXyOln0I+aBXnCK3RkSKRSzSzvezLJstS2TCmf6QRJbpzvrIo2bjIh5zxnsd+5zLpN
sQba3uELDXG2wBJQrtGq+wHD18oljF7eVXvOLGEvtYGp6a6RG2sx6R5P4vwgIunQvMNH9tTfhLa8
4lz3mZPeb9Ns4Tpp4uUC8dAQRx1aGzCr2hI7uuLXSmKEDpzW2quV+UIpOKFPFvNRYtRj1Pvt4P2I
IGBBjnRb94ZXuMC7U/pDmOAobVP69k0l1f352pf/Wzr+sHfBZ7ZcogIlQk3jw76dhOjqJKZg6EwY
Gk0iLr81ZxOp/zUa2mCT7a4LTF+Mzth2ZNmMqkrvbroWq42/LM97hYQYQKoUTMhlRLGVEIoMVRLm
O58KaZki4y5GiCw0XMDfcqJp13bIaFFawA6V2hbDc2f65PMZYcwIO9HKbv0BOTygl8cJ1yxrLF7i
fqzq1W1cWNp11MaNupwzuUcUXFV1jE2vo6GmoCbVjHqSZZActBHv35rRpa0lVKhhBcfk6VbbOeQE
5ax5RZ4w6Uy40mojBCSYoTfp41+uPK9mya6unGmTxTWnl0nZFosjcncDorDhCiVbZY/a+xG63m73
OQQrz6QUhw0korU/KN9tv86XQxm9PdH5HrTEahgSZctpHporrSQFnKMR1FlaOoSmna5q4QtL9JO5
Xh4ufsdClNwq1mjqCh+uvtEenA8ejJVh+aa7fgC2KdXNTcqLp4fttJVD57I4L8nbhFgC3kDFY8Yh
VKI7RM1w6CFvu2nTdiy/JRSvZ9B0LO9jCO0+7198YKQ+2inezumqagvIv5Y4klbHU8WdsHkYmiKL
itUMOAfVXCoRN3uVbQ20+4pzSNo22GKUbkVFNbZCJv6NukIfxC/fqwRW924jGtMSSY/2+PK2UIw5
kjSy8YkW5mjfeXkq79110KN/2PZbveIPMhMmiHYdaJIQtim+ztX32nXkCL4Z0G9q9GNNgj1gR/Xw
sPYxsEvacW9IxFLBn75YW/ADZvhRPLbxX1bbwaR434KYi1yt/hilKhnLp9Kz63qQxFyh/ig/z/7J
OI82xuAecEXdZD9v4gO3wlIqmmC02O5la3c/8LfZ08i/3mR4mw0bnXRINGouyJkCitipYtugksoo
1of+D/qK9v2XMo9PqvCG5mEsfCsXhDRxcxkZ6SEdsdRCWLLpUFbe00PTTZteWph5LJNn4iO7/BcC
lYVS/to4P12pC4aP8wo0BDqwFu7kDIobyIEgrwftbj2uqeb/xawdjni7H/do4T7YAkI3XFDQCeZ/
yrQNfoyL0Uhnrutl676tvMLQH6MT6j75kQ8IqWi3pK7l5JompeYvsOzzZ4hTvEY3WbJ55LqDLRro
4zPctX54FWF9WjifgJagNXgTRcTMq9/DTqGmDMOALiHLFGdkJtG7FBGcrBk2llsmIRrA8huqTrxV
E9h9xDL19DKhGcTnRkVDQj3Swvc4Nlwja86fQ/s4YPoChkSoTG+ElWCxWAuwF/USE/xZ4oIgUTVq
PfiJygaIuq1TmHr1H3BHBUCmheWTsaJUQs7GjwwmGUrsiBcYE2qe+wTvZgzxCqn7QPBJu95KWcIZ
xaiQAkdkaNAZbSVamGgMDDyMLr6nNujBR8IiXnu99iAYTpt9P+KjHXtuqTOpjaYcglqzNC0NpGUx
/9U5k7+HkueOPIAvr8clmK63Xb3i4z685y3frAhpCs5hQygKc7GqDVslRZLCa6bfNgEWV7BSy2lC
NdAqSozr/l/HS0KgyiuSw0cWcKTAWP9xjjPH7wYaxPpIJoM2mgRhg8eSFX5u0KqlLgcpbBIN/Dkc
cCuQt6GbLl/QH1O74+UPtohZCYQCMxv9uXBHhBjPv/xSuiOfCz8YEf6YzbokpkUkI2pWMZRThnhA
06FGw+bovNalW5ISr/hkFFhyEdEq4/YtgnWT0kx9cD4n4wzfNG2x+LmwOUbVxl5ZE7bd2st2oUAm
IVwW8UoPMCkPMeac0mXVaT5PQxN9cPXMVAgdqjLMumt2C8xGxow3PLJhTgxiTkaodU+8cDTAw+jf
ObE0lVi4wgMkQq8/RBk5QlWiFxnTCWdwfqenXYOjVjMXUNVAea/GUwVOa9X4GbwJNK0SGjHEiKJz
FA+tCycLgBgzBjc9LyEZyrS+xHe6r8ad/OSifEqiQpJpfd4D4gXazAD1YevwF4XSNUoZjCSGHVOh
Pa5ifJMsWnKzAmro/JVZP3j9WvPXm0Sgo9da5x63xhNNcWcNZOMnuy/4buu5udThdAtLiPkULiJg
mrArCaKRGHyM8gMR35qZbYcr5CCpF6KQ9PUmSl79h7LJOb0Xk6xGTQDprSHd6cVTycn/PYhIILY9
6RKprQGnfw/aGdvF2CGKLegn0jqWR/68sdbanRB4jXOHFIfZRbnDpmolt5DmUM6AVEDcf29k8NOg
RnGE4k5RZaipPY5BO2mDiRW358t7g5rDvjpfiTR1cP4iHV9hwkKdBytkdlMpZsmwnwcKO4CT9hSY
7qwTPmcMPrTTmKa0X4uLVmOGqwlIzQEoIntvLXyf1DVm/Uk20pXrvJLNp3fmuI+RK/xD2yOqgjXk
uz000S89djFu+PBXy7MudaCAg0QR5zO9c+B7N7DafXoA3OLR53s51aFSnWZXLbRAQXHcik145l2w
x2hBXSsY3ZpzIGvZtpb6qPMYLr4cOhHeqfbC2hr5bbS9xxO1caguSkWyUdU4c7ow4QmLN8GbDZT1
KFTn0CLqZ1JJbtB8oPyrNeOIkfNBr4cmwUCty1CvqFCCIlaULLVc54tR7e50oYN70nzHL26aTmcn
OJ6wsuAfCLgAwCFfhn75wDKD5bNSTCB4G1ROLJwkeWK1LdwCEf9ICDD6amS+nr2KCvFo2vBEJXe5
R23iXzwt/sIY2s5m/TGJQ9u6GRlNreTEcQzlBzUJVjpb7MF73H28M+3sYAipKa6Op4krfw2L+m2d
1agzdpGfiAdlV/0hTWMqmOlxJIgmapjnI74u9gJjIFNfqVHQNsW8JQ7X0pJjyiuXuXHU81glQgOE
vAme3MUHtQqZ2sy6p+C238dtjvxAGzhPg18Gdxllr+lL9LxYWUP+dQcmHXAIkXHBovisxrDgNxqT
EzlWNLSAXJ81MepJYFL8y4VDC3x4cZLVfMqSw1g0Yl5Hdv8Tg5hvNR19Em1Nxdf5AiWJDZptXKDM
aG7/Fc9SHDySQiM53yYQDRdtvZrfHsHXJcQbBUBxyDdnATSb6IVnlEWcb9L9QeeNp7ZfI24FG4OR
6hCO/7wPZN5BYi4mjpuIihudZPoezKFcMGuQHfb7gdhsevh44opyRbfiH5klQ/mOjPEOHLxEEnef
B/l5t+ygNirO1h9I7Z5xIW8Odj8HqwBLFPRFXtsy1tV4hGERl4SMZ8dMPCZ6ADTXP8iFcTa+tUAL
f1tWm68nGBPm/3nMadZv/EAEynyz5Znw3qHdreO5upjRMs5/R46pr0juQGYR+2veGXlAZDHaLJJ5
AqmI2aAEG+ZFXNn7ZryxM4IjGjWFV+W7m8g/vM/fJRXkCxyh3+sp3k1zW04loAJwpa4QGbk+yWD4
1d/OWV2wPheDeiAuFHNwg4HpE6qR0V4t2Lw51j9KsFuJIE2KyD5w+EV6XccLGmZmsre94hUZhGpJ
FQUm2sYaKDe2TEfMgqcX9WNVPRkHE0zoYAsPXTCBOHU0Io6kWJ5KrY4rvfF2Fvp7j3OedV5Clidg
tsjRL5gLAwoQcyw4z3PcDVKSHhWYWxoTWTuXlsG3rljltuB7NkKPSwg2Reu1WMQ7igQhplEGBCmn
dS4C6JgLsGmFzG+C9LnmQ1Q/7ZwrmR9vPnYDfXaMWrMYFFqofhIrw1P6MdiXP2TwYkuUNTX1BkPr
ixEgqnEVFZnNcWpJrCY4L2Qc2DSa0MEnfkUoVm0h/LOw4xAEKe0QWe/sKLlo90QwXmRdyr1L87PF
B+OyHt2OE7wjeAOdS6Ph9u7QJFenvcy5ZN8QjIOfOWErcQ7XFCL5jNm1wAS88QpsfkUD496FXMMw
qYbJymlRsPqBLFQ1vL3zS78EaOXbCdPG8B56BX8ggxXLSRXjS1AgEqt9yMVyqPIkW869fYZB8Koy
+BgvW/nEJ4SYjBQTxv1WFQw7wt6KUiz6cYcIKwXbjDafwyRturwbTPYdQpMJXZNWQUWiQ6R4K2al
LL2wkEcuXokHHwMjOXfSQlAfEScMMpq1FsHGEQr73NNWt1Q/VSVGIuOcqA2hAiJQPjSp/kvv6XcV
yFXDjKT2vG/0RBRtwHZolXQpDZNLYrzrFsE6AfoEd6XADHt+Ypq16Ru+MgUVSM3EDlNxAtaiGqMT
U4PBuw7fqNajqGFE517r3t5iUQzjp0/8Gv6n4aU6EDM3UMWGji7ow7adlF3Ika89WxA5RHIWzJUB
7qn+gRA9ArzOXJVbbBOQEEmuyypWO3+zHzhtxRBNZh3ZrKh15M0wHXu5p+C5gAAFo/Hm9wAOpLma
d2wCL4631G0TL1FYpP7vn9N1o0bby7PlS+vwV2Y7VOdz10LrFQkf1cNuEGE5gyy69U8SqK7Ekdlq
hJc4rI3IZcZaP/puGoK3n9IM5x+R557P38t9fAe+zChZfAwsmaOV4RJ6CHNOIhWjnbuX4BLjVE7d
aqpa39lwQZEPUgBBWb2RdBmU+O/t8APku4jSnTlZS0dI0ucInZTI55vcXPvVsyEt1XSjBCV+YqAJ
nBu6Nnxuiz0zrbidFE8fFWjfOwTpXLDFpGcD1ZgllSCzcRUJ7QKYyHyypuz8pdHyiPr6G4gQo0JK
1owGBHg/fUk7W5VPoRRRNebHEZ78O9K6O4UlTuqSJeepWZhBcz+mWoNiB6VGmnTxuzMThfB8yrOl
YxJLK5FXt4hElkqnpDiW4U5BCQMHZXnABxwgkMNxK0fXFCHKTXiQC+sMGBsR4uN5WILniW4aocMv
duDakiltd6EjE3rPP7q/ZscdZV4DmbZ3tbwlEE/1nVhOnidaQoU+XJN7RqbgDpKp15vjByB+I4JR
9qpeMW7jXoBf8WNzXchptCwCxhEzMcfQ4lr/Y3xs0uqUJehxkU5tcqlRtHNlda9AyZOaqyuA+mUs
aqud+owpY27ITBGOft+MmgZJ+oM15VhJTPdcwriJtLVO6eqJQ80Mzk5RmDJB/zhIW6YnndPFIBiz
U/gv2OkArweCkRuFjyBfonYCw27uH6PDLnW5bNXRVvjJRHaWN2qQTbZnqlwOA2BEQnw5Y4TgFUF9
ez7iOaUXol0e3zM2j812qtat8lowQMJmElGOczgReAwZjJrRZstmLIna6DtCwNA6tjL2OYEmk5wB
h22bVOO0uPDQ512sm4aXTEy2aNUIKVLjp2NrB3jMdJydT4VXXAY8p368Jua4WTtdG6Y4o7d6sU+s
k9zoF8dEWoFzLDxtznc/KYpt/7K57T5mDe/FDAENuWq99aH43LPI5rLy9mJnJGknM5XHX9546HCV
umxIj2oE+lvc0ZaYoSvk2HgsFNg78lgLtASgqki3l1NDOvqhqKS0AeYJuDKIBH0viP2qGsz59fLK
mA+ldKbkpLDfu9Ca2VKSw1o8pQtrKFhbbU76mNOpC0h+MC3V8sIWX0Vym1TJ3eC/4qnZ3T23b0Gc
8w9V8DvGCS7ej/Z66p5AsfHkXI5ttGsIHT9nKDX/qob+gR6jv5yWx9JfOYXMLovjY9MN/2MRWO1w
CqRzI1raUN6bIg+a5tN7sHnnx1J6mfT1vXiwk7HI1bbtuoYvdOHm9IoxLGvzMaBEy/NAYfkBWItJ
rZQXXTK9SxPA0v6HLJR9xAuwZpxkfIUBvSm+CrFwlUt6s6b4TAqQFnFC8eBwLGAJLbf9/bSr81L6
+5QOa494ZbzCp7s0bw+nsUk0LfCZzsiiiCslCp359mXGkilmqhyPV91MCAvzJqORFb7c0+FsqqTK
uwTGmgKFMThD82plmmI24tTKRDCIvqoFy5Cs2bHcVYNRtrtM+7SUFUJwe2HzGssdQD4HeMe+lP1e
+Z4372HDwfwb3MqGktXnxt9gkzTYfcJ2R7edDDNQuPOarbWaaYaOWxSP9a5wk3YOi1Gg8euT8FMK
99R7O3K7mubXqfBSH2LScaEd6zEhK1ir5c9conOWauuiLqPuqt/WKyY38dNzD6sjw5MY+3z5FhRw
pV3TyH5s1Td+07wBw1L2lAGZolGETEvuCtSoJkvbLu4nxLApq47WPh1WGtvTGcft42nbAraaTpz0
wQmYQ5sabwJJ4k6vJGhrNjYAji8Vt47dDa18+ZQPJUiS92/V2beeV8BlhAJgTzchBZZkgS4kzfXV
ExXfcZMV9PSDXMn4zOI8tbHCknIBLAPRg9R+0xjgPOziQsmgkxa3c5g8CEAVBgbEjHjr6GEet5Fe
OJ/XHz5pDd/R8wYd8H3jvMklSrX38AdyoqgZXLjcPXoydiAp/Wg+aRt6LmoGZZgQqnFHbfV/RMPN
JrO9o4UBBSijFTr1IxcZbJWsalkdLbNgpUuD/kp1OgqgoCFlnyftaoXth/Y44lP7tMynI/IYRVIj
C56y23qJZ3rl16KJeC1r//6lYk+m+edpHjWqQL2GaasjzXSyyBHgn04k8BfB4tn5Ve0v6Dd6stZ8
vRz5o/RAebUyPXGCkTtmaHSDi729aCyHQcejAvX3cQrTLUmrF7z58II4w0z04aTWSZrrjovA2WyS
fLKicOVu90PQMXyaPz1Lz0gx8uKFQ465axsMgIbnuoxUn4qrMEYiRibqwnOS/7U7hChB6fXhE6QX
v146lGHr8LPL4G9jTXv5vawBpECdqC/IYMPFpPmi9poOk6CwqHkvjWZ1PcbfB0yM0k2D/Mvk4CCF
C0qo7xH0XOKXse57fVG4WbamVGpUzcM/m6UxDlrsMqPf4/v3ufahU352g2c4kczU9zCt8LOrrnNs
Xr1gFX81dK7l0IvUJPlH7svpUtbycDcUmqWOSx8AZihqA0e8zp77L5aH8XLhCUwfpALmeE1VRS5u
BFHEzrDqbiAEPA3Ovh9Nnbu8eYttLO4wpMFKAw720w7aIcNM35Ar7jBUTnwT177a8Xv7p51bguPY
b7ofWDd63Op3Vr+F1o9wrX3fT31JBVA6yMKiZ6ju3GXm5dVRT1JouhCQw+qDHDStdzyrrVlGA7+m
v0lBng1xrD3Jvd7QDOZqURTp0bWEk7pmkNxk+fHkqSQg3EaW93YK9ylAAhXprKQX9SsfrAXtMAUi
+eWntcPjpEjIN5ObwII62MgjpYy15/dkEHYnIzKZmPQUlNsB/cu5HXwwkb3z/zVUUDYcYFZnO7Yc
S5y/rYUEm6Ic8wy9grPgaVzbKadRMT6fDSifEh1sCA3NOC2WfStP4P1BL9g/WY7WsZQ3NFe0OjD8
P8qzk/XDkaK944dyYzKmAJeHf40Xcci+2r0Dz5X9dHJc0FPsARDIvlqxzrKmXTZpMk7nqyrp35U4
4AENG1iKMr7Xb/+ZX6bat1JOuPP2E7vAUjrJiFm/qjRf9fWYXu5hE9JabhTRu/9F11CV7e77Zbqn
oCEU7AzlfwJmsXbIp/E2y46n7kP+fqzLPi8d9iD1MangVpjE/qGEgwY57A+KRPOh5aejeTa5dWMo
5QyvhtgQAx+k9M8nzaxdOdnn0R30JbVMYnH6lsaNb1bEFa+l1aLbx5dd6TinzBJw6EsID20mUwBq
KPWR0uWnxmXEXIOUen8K6KdBkjzzhgcsEabKs/3AIraO17L56S3EY+3vUoyNSeJPbNXkeRmkg6r+
wM0EE2T/nxUQt2BJMELDjVMhiCzN4kgtPoh0n7DGhLjbQNsT07R3qOIXol5ZWuvMv7RpKpnxf31v
4Aofh8b44loiQpQIJtzRbcIpbC9UHFL12053Kpt2PgR2dPsNZA0cLfkYP5wB2Ch5PTku2i2eZoNQ
Qfiw8q5rfVMRSb2xGxJUh/Ry++bdbbhJPOVVbBIEvGYFKBBLh9bVDMXaneQYcVehYkjaJEZxcfrU
3epCUMBvA/ABpXQBOiNfmQ702gur6oNejYmKp7R/Uav1EoJP5fMlxu51qBt4ybQoYrJAymczJrmK
qXPAZI0Y9nAS5jKLLiZoQVtMYX0OhIaTccLqfRLUkE+fPlEh9h3a/CQUWmymYp+xpunJ1HBLBfre
aDYPepz1NAEJcJGIcKok6l3HuOLpmaWnsp92eIE1ZBNORbY7sus1E14sgLj4Gr4sYPIBP9CgMfhE
0zoR/zhrh8GBv9vdtN11IgsE3uD/tfAs3igNxLdh3Jptg/Su3JiEGN+kvzLla9HuaS0HVnzA/qCx
WZmDe1MNGLuJiIXCl2tbFfy5S+DEPvfh9bGhhV37xFQVrNQP7KD1V3BUdKIWur5Vfl69EA4djj2O
JnawY6ydlEBOuBPnu7HLJG5VZNbbqAGu2UnF6IM9ulcTtrUD9MnLsCENIGIHKhWyOJ3N6r/5D8iu
6pwJMXdpeTVufhtWn7IoPYLxRyKOWoEZ3cvIAqoCiGQc/Hwp4cBlceQnqx9fkjvFJfh0UdS62RG5
QYYi7LGVVHbEcnaGOYDjF4fTREuRevbEUmHmEVRfSPIYE87UOZ+lJQQ5v3BYFU2RFroboI4qKngj
HHBzHP2VDRfscHUL6PBHVTlKKsVBxhkuYcwJmBDiiew9klNLAC1/D5ge/QeQ2nZ6y898uBxncCzn
BSOXfmm/OFGc/5FptPlyUqB2KBUXlaT+fMe0IPn5s9eDc9Muaf8kzQS4P8WUY/pEohOwYWKEacgZ
430TlPI7758FGumokg7fW8kRVs3a41uVLf8hFQyoB7IqZW4a2pLCSC6FAcG/+i7BzQ4KngEKz/hH
4EEiDqaacijXWrQUIVeGKk/Jw2TqmCVHtG/0TFl/1aHRo6IDITIKGXDg+Rk80qzMvyz876ehYaZU
8Xo4mapTd755Id4CRJX1pb7/PWFJvbIk0EBAo0sFocuU0pK3NlxXQ4UvgYRQckC7ppcFupM99sYl
STiZjGaMxys2Gy1AlO74BS8FXRgIPdgpg34p3aPCjdqLL6UUnU9hkCybHrRHaTLNglYPrewg0g2w
mTgwqW1leXQFj93I4SXct+iKylpimx1qC7vAfk9t5fnBeYbYgj2ma0hzW51eJghH5CCyCHsNzQEe
tLRWHHcgu9uBT+Pg2RnoKdfrPC29l0b85kAHfG+ToCpKP8kTx/4ntqQUOm7u49WHc/RnsyVssQfI
8ziryKCV3QPGzUvx+moTzSI6mfXJbcIhXAg+6S2i7B0akwbvBQlsYpWihFlke2vO2jtZn9L2RVOM
YazR3Yr8XJWEp1DvKOmolf/CywwfJoH8ooY3xAPrh7MsNuuQHBtWfTJryADELHxkHQaLNRtjy8cE
V4NMQV4Og57i/+bu6rpEYUTPgHwa+sfLZ+wmT1kVRYh/dC/cLIj+/g/pceQleT/C0as5/fV2kLgI
Bs+wdTcRU+YLbmPMDkXDRMs77tZF//LHrAnylxzhRcKpzkbPTlvhMkUHlDROzMs715oj207MKY0e
nckKxNv+edoEwvYUt6UaagkNk1CSJTA7g3pyNfZcQDAR4gyyEbDDP9xdy6Yu3JK+DLtxyXZpbLyz
L9Jw4w6vscVfCDIeDd96jSdeVt4wqdOXircDuXX/ZUTanDhp2KVh5ecx0FMjkiKLGvEfaPXKAHc5
oaC1JuXWPIj08FhrU7NRgqyYywJTVRfXKn/GuI2tSYSU1RrF4iwy1yq6xuhb0hmizC94dogtY4H7
vEEXCKr8yeL2KK6YoLZ5ASp/BSjyG1tlymx5pATM0WAeT+R5HW7eJswDwiiFo8SUHcBe8bh0ljF7
nWxE2TttfO71q7gEFEHxiAezEb8eOmX1ihDEoKT0ItCGW/NnA23Bx72DN25/6daf00d8DoDTZlX1
WC2A4ANRwxs2Y1t6boAhggLCjlmMSq5GpICHiUuPDvlNd0CaGjLQHdQVxhB5n7fXG3OURNobAyOs
RyfU3d/+LaKkfNxA55IAQ+amENA3uLJp0vgG1pTf9GxcqZCk1tkW4x4Ypd0aC2PvohhRf/oa47GO
X9vU7+QKWpealR/Dz8MouF4hcRR1TmJbjj0TwKGzelPqXjRIwHZawquXfG8QNArx8MeEJeIXe9lA
1WRzWq2yk6XYs9RJjFOspR1ZDmsUj7vUnRmn/l0C2A/uXflx+XSPG1M+963Z4C7hddnylDpEShJp
3nD6jg+uMPpVC9aSPExeofUHKi2U5VJuhTdp84qnESJPZ/5hQSb/2toUp/rXX5XO6GNnVIhO+h66
bxQ6gxLZRmIHkdemFWpUbz66DEyd8CSTZyGO+Kd5cXveGalaEXXGqA2deYxXQVbdK88mfU5Oyecp
FO27ghr+vmUMvSWuqmEfScddOhdaOcMZqAMlj6Uwqgeno891US22XgI/lEZZMJ2y+wIRZbwvUKFl
/p0KwqPLuvIsx9j7UVd2guO5MTE4/xOr0fS0tex4ZjJ2rJ2rWzXk52S73CtgEjL+pgdf2Cb6ZAs1
3T04QmmPVKQgnUC5fDBsYmkOnDiIvgPrcEmX04dvfAApAWWEFJujv5qQ2l0vq4AeEOvBK0E3nyNE
SfVDczezN7AnG3apz5swqFW6Gi0f7kZfYQMr4UrxjLyZNJutfY93ofcFZlBavudVFYvpf89CIrYe
KdHnp9r9JAY+j8EqfZDcYTKZj9HXfq7adAEaTnqw3pQiyDcPtcYq1WlJwpy6IOps+ATgghKSwMB3
Af1Bh1V7jy0jqjd2d+RESADfO2ZmZci62FZjeRTWFOR6OH38WMgb/ama/kghfes7QqPy1KeY9vQv
K/oGAPRl4psQKdD/N3P27MMEFAkZHAQcrbKi2PdK0mC3RfDxma0iusznkBmFx4Eb+fSRxPNuspGL
aFNAJiIpaM4o802WOI7z3av2TU2a6tueulw4PmIlzylUTm772f8pbAoa3+t+VeFiv9R8nAHBQsz1
G78td5W/dwtJf1/OewbHXGITr3h4/U6TiXL6NHKxDCWc/5CKiZx7X48upA4BN0LTQOdKthCG7Tb/
FrvaJVu8mk6exUVofx2SB/mKaVNuREYtSAPDQycVbEtOr8D52r+2pgV6VzAo3tVjdfP7tAFbFshH
+/FVd+wn6hcT7H6nL2yUehRcqzg9kSDd4Rk20TEF+1BrfMH3/f3sB3EQkb9vE2CD6QorjCse5/e2
sTirpFKNJIFY6moDm2GOBqD+4L/rCgIjYOMd9i67NcASq8igpxNHn6fv69oSWksC5PuzK3ctYOfY
E4PmT09WCqTOQK6ayaeQJdHcVDC2WWn7+FzdAwB7rUbEgWoUR4MjDBNM7phO7/5Laqg4z3CehaH2
HN77fscwpC+HzVmcYvoaTZ2AEfDS4h/ObUsREOqYxZ026VOq0JTp3HcD6QiaNEA1in57CeC6xDe/
uWMotVTfV+kKZDe5Tc//wGMxV3nplLunUOroJo9+qlGRgF5HmFFZXN59zMS1ps8gkPMYSNCuwyP+
TcAl/AJcj+guOWb/pwXBt9WRfkBmj0gSYyIqZHruvk+Sb45wqD/wUacolKJcF8FOtmXD2g+u3K+b
m9LtAyBvDk6+1kYGl3XqF5zSHvp1cuugTnxFb8sSbYmUU92bt0Tb7Qunvua7WVI3XvY1eiiSWmS4
LJtaMjzjE1aaROCyVysR0bCuhmSpkJQbRAzEvtAjwv2Hva9VZCNVt7Oz4TVOrMTJ1gwjUOg6/7iz
20TCZ5cqbpG1Z4+nKwpWDnqlejd4uEqEYnauIVBojxJH9Y0h0R8o64actw4kWTWyGLnuOEKpP7ji
MfZR5+hHvpdkK2EX68WFpFr6cB9pJcxjJAW+R5F/NtbN8at4L5YaeyS8r2XjpLCl3S4Oaw9QMlh4
gKG/vqo4Rd+uYy5IwhZqIK3pcxRovP11FxdUfky9ROudvzLxBNhGpgxzWXNQ5epu7mdTMitOGydC
lQSw3WYT7FeXsREhnUfQ2IkWiNOug7gLzDuTz7ezUgo3/5xr//Vhu3IJDMM+t8wW0o4DTxX4MJzV
78mNz4E4wc1lWuv6yXJdEmqM60jDUFeZIbnxsPzcTY7JBKE3RFdK/+zKTi+63ImSmFggc4y029MB
JjnFLPTF2eYeBEUBK6Vt7CQ/lrC17mVSVW5DT7G03R972Dpdt7am9VctjtB8oDHtBVkYaZTHGnKv
rfxRY9vBS1FKu1scYL7tiaXD6u0wYedzVcxbKyybYxuKiDn3n2aV2/aL1Yv6J2ZX9OdErUC5A8RH
4KIWz5LXYF8jkUlgkEvDLCrWGudJSryO/tP8TQtKLka+C0njR5KqcLg7KYcHDZG18WngqJVyQZQ2
57J7Sm5cj+5V5uRmcq45EXbYtCrk4folAG4E7gF9/g9Y8/c35fjEuZS71G4DEKTFBPw1FdPzmDa0
6MKwwnAkTHCy8yNHTgjNMAPI0qov1zxhOy+Hnpa9Hx6KAjsynmJorIPHbmg8AvjE34wWZgjXn9v3
3r6IPdC34wpRG5qrL37pnmsDsV5YZ45iYvODAT9s4e6f/t0opjEgOot5t41Qzhkzg6OuO2wvAt4A
/G+1VlKXVfsmbKnz4k36BH/0++RXNJBLgYDh7S5ZOdhlTiH/Sqb+T43MxqWaBBB3S8k51kYsd90d
St8RqrFjl2X/dTtZ8Oib74r1XOqnTMwKDckSK2c0N1UVrAZt9bBrCk66RwIZzbzBsqiXJRXc1xdr
k1wefbu683WJyL3MlNa7hFlpno3s1TQdSMw0ZURqv6fzpCnFBf2TwoAIJznBqPJ95b0chDfknUcJ
U0oXDbn7mdMEz7qKWea96BTiBRAFL9Tq5xgkVuAGJ/bKiYytraoUDJXmBZHpqsz0Bpq/vT5k+Oxk
y3DGBcYaaSC2C3kxQaR6kpj1fhCBkkSo0jxh77azZ9XMGTtUm8wu4tvvF3LauQKOy2FsKOG09QRG
M1z4zJ7+b1LADhkrJvM/rta7VA9DmBJT0k/dFiQD5fTQLNafonf1uDvVPauUs2E2nwNNQym+O/ps
hmNSuRYJ4E550OEdzFSLxJOSTHLsYKWwAOBdk64jGNEJ3qN0SW+Q/QTrz7XtXT7ziW2E7AbDftZl
7L1bCk7YCdHmt+DewEdDzDay47buE1gu0YZR/9Hlztyok41962OOQwZgfwye7ESpBKFdgZjQwLRu
DZrkM720brfExN8d1cv8xEza4mIuhiuim6S0eDlPVuCSmZll3/MHzXpTmweS1sr4RiQcUvKQI4nX
yTn33XYELAHktkbFyyGaSLgGddXBR6w08o12/wP96iIVwfSsRQgNADXtMz7+ukyTn8RCvItzRCWn
kB+Yb8HPNAH7WmQ3EbcBz1yxqAtmg//8KKGXe7vjyPafHFmM815VNM6jfK6+0hYuB+pUCh/c78nz
WiyJD57fPVCFXir+5hNn+sXYJmbhiPgrlL6QlRpFioRMEemYwP8oQ3zB/MQC3NG7Sf806uJasvFx
FHC9fXLg0hlHKiI4uvxgCNKlYmVT1DSQ70F7+b/Uf2OieeR3fumOu4RESVYeVCrFg2oJLPQUbUKE
CokEmFGqt6GUDIp0Z6hN+CoBONPoxg+E6KNDV9t4JQB7c2gxAwqJ1sMaik9edlkE8PE0o1yvajj2
2q2SToFL+CjlI/QtHkLpKKbW8/Xh88TDHKXFWFX7gdkqhBapkJYQ6SPiOJqEvV8OcKf8e4B+m8+E
SYKUaQIa83FOa9RuXGiQ/TPkF6SQD6R68WS0tKbXSBpK2pQJjW1/ZDetfGG1csXWRNUTIpildKJb
dQ2huoILLLnWGpKbFBCHpkx+Gp1zrcxUTf/GI7iQ6FtbuG7YFq4rqq3STadXWFy7Uq1yyUrSjTFR
DckQQ2YIWKkxxJ1leERPZGu4J1+BVeKVVIPOl9H73o7nstnNN9z2YYV6aBuqKWtABfC075GiESkq
eGnGIArPRquwzTFL5SPkQ/srKgji+FCU0YmssZmRnyRpcWnicgHL8IxmWzcjWendYz+W150ifmvy
FN1V9D5p0YtVmGoasc735SCzRkGWfHeQ24m8eYcKQzEAnKYxvj09IB9qdV60ETH9di2AaIu63pQZ
FN2LTddoOD2kmFEv1iyE2iRf/o/UvJVEDrnc8ve/0HWG7S1Q7Pv/WQ/5IpzBFhouNsmb3elZgr+G
9JWlkDO8UBhPMI8NqKKPIREu1xgnCP+FeDuIzKifLZ4csbPkhRRuP0aw+Qyz9SF07kubdAy+6Fli
F1mf+5BEoQ7z/paR96P9kbuNKA4LYUZ1TMcgzYf2EFVr4QsmbEIjyGyx6s7jgnnymO4qNYakiA51
O/CyTr5UhUBfp5Rlt/vrqKXSSLpcktRXwrnuzNpNu0DlSsXxHFq/pvD5wBEbDwOlDP+Cjfz3sZ+I
lDcRSOlLREKNkZLibIGE25Qv60sU+6aYrbTJ6lgazEFBa//dPcOR1DrfLs1jMARfEnfE27XJbMws
U2+6zmAkjHEx2GGJ3+G3DnBWqUN9CqUYjCT+gAhjwNm3PXc1ZG2DeZBainclR5gXlWDL++oLsaNt
J/scr0wPsEoNnkUikZ4/DJ8qGz9KHvks3imI0DW1ulgUGZA6gG2upEZ2YxuhJPcOIGuiJYuytg2D
CbRWaU4V+FixrLMsVdeY4fagsPQXc5DYwvJqSK91MKAw8ld9TPyuZ/ZsyUMpUy+AX7JN3oamUV3V
Xkfq334T7HxKVPybe1V7xi+4oHnLAJWxwkrVAJXIamW2XWmjM4/pP+ia1wpuuifwpn1wovrFKrxj
mon9I9yb4MiuE+hwO9wY3NcpSfGM2L7JMx5zW9IyTigMeW8Uj9usAic3yRiYwgc9VJ8LsMA/xdnN
R0L+JoMyAHLkufM0xCcT1jyrVPpi1Zi+rx+F6Ra7z3BrW7uGlObO6Dri/asJz3XnSpg4aXZhHrto
ZXKGNYRDP4/sElbcaeHBUPy55o0xdOkHqjCdUrMIGPOTc6fnzeOTKPTyETVzie1W34wzkhdvdF0m
hclgK7305Gci388T0bqnLSECTRjH+9UvhAT/vXcbrqcZIK0IxgeJadpRlfiS9IzSdMVXztmYdMg3
9iDRNVVXjmcPPewA5d/kuRdGXVWkwdIDJuET+xkZUl2rM1Gr8up0cXsBdth7fvmwP4vASDfirMVH
FkBCE/iZFtB7ii501T807Rrb+tST5d1Sonvx3BXTneJ4gBNOkyLFL3d/10XS3hRBWqTw3+NoULqp
Fp1iEozj4d9CjINdmq+6ZtIH6Ye+8PwlJzxMpz5se+/4dJkQJpkjg54CWaTTJPY7tJ4p9DtHEyjJ
2j2sjJ5VQxfNaInZ8vLRdyKJ2IcDtNcqLwfX2hPjS6rJORmOou5q+ISNvCQmtkD2Vj1wkJHKVCf/
k6Zo7eu2eyfBDwwE+0/b+0Ri+Zxgda8+o85LJ/tKcxQgTzB63dGb04Ov3KZ1JTJlmXfR/fxPqVpU
YhDeT+CgD6fUXoxovP7scm7VRdGyGDXL46yFPg64EH2TTf62zJa3w5Qt1tx+TaIJ4dFOctZ3PSvB
ihgfWo0jEnsZpLiI5fDKdT3Xv60u6yQgNlJaeN8jC3QB1Ygu+dPOk9cLD3+NsFa69LD7V0YDti3F
uiJBXIpDjdo/0tc2Vzv+iNiniluArdM2Q9Qasozf0DOm34oYe/guPXFKrB0Lzg8MBzsrTxEW29lP
3LWbDZPikV/qtA8zXaoGwUyDUqfM+EQp3c1XKP6GGHnbNRKkNidbjFLGreee8FqrMhzWFZ2NAhKp
XN9WbOoXPeTO4rw4MdWqvY2L+QwLxhzgUtsseFxc9ui1sw4KRQAgC6fxJWfCtOJ+7yO9jbQ9eb7Q
B4MEdMBkfhc392KhccfcflBn2qVg1Anbt4W4hlX8fIULoYxXJeX0McOXkUT+tdJt2VQzfpeo5KxT
xPgQRc7+zxmIOvniyUqtyEO3D7k43BBcLbj0iOk7GxKdDR/m9cBBUmxCCExtb+3j/fxC3TmBKcrj
a3YEKC9Pp+u/XTxHueEyhEsDQ7wHhMmfAdJaEPSePcFDkhy+VyIfNTaLbJ2aT9L8rA77rtj7bu+A
IcVDfRYnM8uMvy8e+OtI+3WE2wZw8h+2RL4PKEAz3cWgxNyJtqBu2VyP1nC6VJnIYsB8iVutJ+mF
Bizp5q1PnSMbNGufHf1xvszyIMEPU39tQDuaQ3ZCT3mjI1QM4loaFd7F28m6AfcaiCld6fuWSPoP
4MQtboSOvJX4hRxBxRa7jEMEfdLjY3yvR15slBTnDcseUZ2VpCoPaC+M210lOd+Jkk2PxHTzuqAw
uEo6NYDxHhoNfe1lIfluvu6qUH+VOGh6Lm6Yc8cvMh1PB2YhzdMXD47SCPNDAa4Q01/o820akxRX
bs4e99UnLe+NJ3SV/V4n3TANDQ+JmMW1QqCJ9fy1Qx7ixExb5w8QDMTxPgEsQ9b7qGBGK80XOCEc
IZzm8ZVA/QC1PTnXMs4Ka5tVxReV2HbIHy0/6hsFwmktpAoDpNwopZ5Oc/sDb602xlxWVQ8uwgTm
YLFFSWKuJtjamLyhea5AXpLQ9rP/OspevWGg5/0W6Twtk+mqHoiC+mzRcgOn/Rdoz9lRHk2MVhq+
u/lin4rfigmpQIWONSeDoxwZbMAA6Tcvj3jcEW3XiOKj4RWFF8PhsYXwntAg6eHea9U6nmlkSQRK
TDtFRtVjDcvQamnmxvbt4H4osfQE67uXaHS506PBni95K4CeKlsj7xL5jhymzVmuXpxXr9MgTYy6
iuOuVFePZk01f9jyT2AiukfKHJs4ERTUDbBnFU9Ep+3krAXKPnlIbfFGPRx3En334jikVFJB7Lh0
wlby2b7M+1tIj7j8IwncT9I9G081f1HyujbSIqleTaemQo1dSf34Sgmmm7S5k4qjgD6OkJOcYr5S
M40apHFIjJ2LqtNsCkS05TJaiE+4PNdJWBcGhUjOVL72KCXI5PdKdeeAlkr8sopHxEvH6z7swot4
riQI1MVlW1o7sNLWTXnJIzpxBD7oEDlBAe583d+JiF6yqtAQBQ6WICMwaPSGyWCqv3X95dnSG8dw
udtSCgAL5SUJsOzT2u4tAziNK3odF2yZPj8IyH42Uj3H75E15Urgwxeh2O8HHx5uQp49gKRj5Td/
KjzNG8TEbnLjLsb9IMkwwkHG6jqLrsBEx8rPkzBDIDV7fFxIL28DIsRbenj+fw8L0duIlGt2wl9V
lP2tiWLAcQKGrJ433EE1yDyrnvfLNPKIycENKu2oN/Ife8vAl+iuzYlHqhypxVnV/fZZWIFeph0a
10Gbq6AUz4l1lYzSpdSPNQInGOYotQZW7+inpJbYLPGShlg/7+Z/w+s6hOPfEWuRfEY+35jjre7/
HdfSyPQtCackszayrKAOajelmTto/GTACWGz5HkAk61sjP14JLBTrBS8L1CWeNOKLldZS8FlB09d
PpwJl5bZPGbSFu8LeTkAkPuVCw9VZX1Dp33fZnypXaa/M6cObSlA4Af49PJq4XxNiTseHckfgRtG
im7oFfIPBpfMW7ySrXt3x4N193H4Oa1EYLenLBoZQMwf1DW7gl+Om567sTLQ0fH6MUEnXWFLpGJW
j+HW7xZoxAEYI1RZ2Sw2a8SE2ozoE63E+2Wgq7EnyYHTzF8+YiFQCeTm3jhv4HvyFA3GaIXRilF/
MIVL170Cnh2DWnnqjIIzvl6LQEqYAuDXwzzAr5QWiKT84bzIn20Zd58LRQMwPSJjgH59xKagv5Z7
qbXFFafDwM7Rry7K7rLFEDHY/Bcsl8GR4dndu2KK0hj1NR6j7pIdbnGiwVHo9He3hBhsf9mtHoMj
j+pDVWDwHFM0bOXK/e/WoaNk6/CJNyEFvktBsuU02pyOmlKFAczTdzhHK9tL/v63NAgnCYmSp6rw
LcG+owobMXV0YH+tSdgmUezAyPf7JocrvXGobwiwkgFCffjs1lYmw3hBMVwejjaQ/YQQihHP4pzG
WmhcY0emBqN408SugFUi4tsxpPmwL0Ud46QEwWtkCpkmpAnSgzQR7KHxq1jgKm1i81DWUWVZ5MKr
1Fyy3f48Mvl9O3mhchacuQKRAAx7wYUXiXC43ruWI8sixDC+nwCjSIbBImr1KnMJLBCmy9hlP0ZJ
J8OAiRiN8nNdPStKmlUXJ00Rz1Cgr75ebC40N3EuWK5izC+NEtnaleZtIwTjQaJZ0UTl+EHVMhl1
7c+u8qfWDPkt6JnNSiil4ihQrA44OH1n6jqHyEM9QLsuTJK5gJZrBcokuKO3t8inMonGe9S+1ln0
9U7odRlLebGNEjjfyQSOdLq6axgd2zmIZ4sDPXX/xImi6fsCzS6GYLnlB1oqVZj+oq86kEOlScWA
W92NnZgCtk5EuD15xsN6OSIskdntyoOdyGOL2BzBDKy4N14Ghb6KDHp+1vW17M4VNbm5Uie65CS/
zuMmMce5RJJo29YC2aODAsP3fj5fCsTDCdXVcVMaFypIjT42XMi1/jRiSDJ07WcPfu0pVP5EcY+H
Y6GJrlDXZBAINqmxZip4e6n4t6VSGvDWp7v4f49oW6u7De6XDPk0HXJu3FutklP9moKmXp4oGolD
Ub3qMSE473aoSOsnzmt753Ajc61BKHK41xhrsv1w9CIzqROzcwp4qLqu8RMHv61o2L5gSgng9sSV
rMC7F5RdVQDZkUN1bLesNT0+Myu8AAfpXfhcAvfnGXiKSZ3rNxAfcYtp9fOI6vd9Ekwic8T/Gz9E
IzZizrqziZ7VwYhQtphNsPpKdgDm1PUtrrST0v6qdpJqlwGaAO9FTt+nmkItwVFCjn2qrTtB3tRI
Aqe1r1upU6pFLfrLpdkv7FInCBd5igNLE8wFNO27jqD70MlRm8RV26bw0DN2dE8RZjiNtXbTEYCR
Fc+eVWRctyPvzq4UIuNvdUE36Wq91MBONkE+SyR0sli3oper67MlSW/7t3QfO9YHBtJedaFBaZUz
lwsokmQ/a8ZIZpjyVZncF/+V9UbWq0U5Gj9fYddGTkStl11tjH+IZ1CKksYbRasZBPJUQam2xXds
67EawI+g6wthSnL7rRU872WXHYf2TIAQ1R8VwgSo77tyYcFD/M4whklEyRIBsZ6aFg+L9v2OJ9dR
+vX1vTBEVm6P4HSb8qmdJnRCWojLEhxIox95T9k2Z1bOMYqtftUf8mWWfUmsIlRxTC7xXbfe+O02
bPr7749Igeqhc0kMlc6qJ6tkI1mm7k4Ilm1tkakX1LbLv4DF3yesSbyCN9BZH6aKzKkNNERFM96W
7r1DQsjSrdVvw3whUKEi9xaEr89IabA/+DSqRlywFlkwhTOWaXyseYpRhgK32b6RVh5pTcaU1lnW
42Qu+RqJehMvijjhdZva41BT7BokYvQtyb/uu93830ns2C5nHqTDrpqY7AKdUEbqxg/PzkPs1UNJ
sn6Jy3yOAvn7+x/wSEMEEpBRsECWXdtGXEt5hlrMrB073jhiRGNCkZoVTjCZBqVqtWbkTZmu+8Jv
6RetcbRfVLPTHVoV2VK9F9j7yvAbzYJbfYIEH8gbUuoj0m1g4cp+QpOHuaCH/9f01Twteke5+9f1
ih8nIGZQOmkXLx9lKoOqfI/9BGohC0VHzqy8QseOfzIhrqKbl2fQQLmkHm41auufg79U4vMQsg2O
+AoGamf+GdeWexw3LAjZOjCra6Dh1iZ/Q8TzcK5VWYA/rHY/pguiSDXy6n5X/iqFwUQGIKUftKM3
2yrVz3xAXUxnLHQpXdS++Uhkv0ouwbeJUxMsqbGur64DQ6yPNpLqTl050hjjIwU+hoXZkluc2zQR
AZv//+WXSSsmGGH/XAa27YcjqUAzXYVx+ssYf9N1Rczg7/saHpomf/PC295H+cxkwWYU/ahqZ7sx
cNP6DTrBLB43WHDV5KlwMpHU+inLDkIXCFiT79Ig7jmY3c3L38gNaVNQxYSIkE9Udfj6Pd79HCO8
7uhgEPKdVZAa4F/KiHEq335RU+8PMHC+nM5s7xos2EnhVE4MN958Pm4d2yvujUzvQ5w5ZfDTTPWw
lX3GtyASDigAqFKRv5jswQIrRNFsSfVbBBE6jTRglSGBF7/cc0XAoGqC5v6nMy3HW1avCDC532md
OTI9oB2SmSwtg+S518XcRp4vahE8WhP7kWwHx4FmXpStnpofavQ/h0iwKmmC2emkbZBSSKTDZoHY
oHga+7im3hnPME9wwl/i+ovUb4geFTwhLa48fXAUYfft4gVMooHhFkK2TfaniSKeZZ68oNTSb5po
v7Q7by+5k0D2pRAG+DTnFeDY4D6ZxpqA/6/FTjBHV0TjGXgQvtDr1kdiZqXrqTRP0dtxIOTZWtTe
b0CvF4UpNjDKVGR0tCcI3Z8TQekMbNY4H4MrhQumM85+MX98YDeYVnpzv5QMkTm0lMzKvuqBVUPU
Pp5SfAkcY8ADpUIVHFxJ1y707JGPqeDxcYlDTJgfiwC53SMLTZZjqTPyDkq2UnqhUc1hnNNzFRbo
eSv1j2ANiv+IfL99WecI4lXP5efu5gPiAe9PJ1HT7nHPum8UNg6R8K6U/4j0aIKXYwJwKOcw9sb2
DZRn1q0xo8ZLmxcarae35cVobllUlGnZB68E5EnSNY8PJJc94tUFkYjSR/CVtyRk/1RbtqhcSfQW
mBXIO7hX62xVEGj5oowaRU4kBcwyYBTiM0DJchx8Cri622GGYG5uD78ZPIRDxiQK3iS2DZldNNXD
XCTzyg+0ow9wGOAQV8XyOYWBgSbrL0n3plr/t6l1gVqj+UymDgxuNo0t7duzvuWfyX+U1XRcovM0
rc6ymkwJu6RmfnaNOIBy3t9kZx/XuNe4LoqCfCZOS8zepB/Axv4G7sqdbWHS7Pq2P3FRbTr8607o
i2zjlfz4kuX2h/HXPKte68evKOLdHbn/MKsF4eRF6yQh7U0H0Hd0nDvLc97we3runv4nOv/zszyH
UoQ6KlqEaQsy7LrfDzu6v1Wid736jJHadlbw+WvjFgB7LQRXOVitbNa7mcXm6LyiUjxCai87z/Uo
cVYfcUTQEHGWD7gl+gMqhjaEE+jqT5goHRPuvOOhxv91X/Ljum8LmMim2XGwD1sXAViV9INzfaEw
WsNThA3pgsApJYfymyCQ+meB8lGlqPQ15hx4E788L+Qe/Uk3xkLRE9TY1eWaIdYzui086AQCFd/X
7UDs4V42gS3txv8ABF9HHJl75cb09zVEwAoyTmY1hko96TA0/PtTdoDBK3U9ZxYrjHnQhwb/612Q
RinDtulCoddMKlq7VTBvJbNZkbcVIUM3BkHqe8e1zeSL0JmAnKMVodxlxwR2dmxScF7/dgN9UoEv
vP4j+r4AWg/PsldDezTxBX5cirIpYtXz2Got1pZjmjS9URYHWcUk7O+HmGsUULSCzhFIHYkmCHAf
PSm1WtltiJIi3DX3nK6MnwG2xzfY+YuOR0V33aaBqKBUwUa31/X8l3LW+Lim3fUmdEjaDsR4HGcJ
laiMNG+ThnQ6SREuPrX6AoeOT/69mQorKMV/CK+pwRYZQEXioeOAHMxor+GErcf+lRWoPSQ7KRtn
sL728+tQ9N9oT478IDe6ltdiITiiDaI7bABKIXTF/Af0rNrYaUsf5ZaSAl2EGdGU/eugDtrHo4bi
okDyc/4lPC90bILQyg1RImI7zQHt71Q61V3ePX5v1AYh/Xlzej3gZsfEWXs1Ona5mLqgd8HRQ2k5
SUKxDqQ1WwN1UuRKWDA1R1PtKOMySbIB4lT1qp3DXnj/X9oHnq3z9p5k/7JkmI7hCXcrcTE/EIzj
4SXzwOd7uJzOVw7x4fRO+1p9e4XZRbLoYET2XCexHpzcOZxRu+gtrMXpvEvjpdCF6dkFUmFvQIDP
paMsFCmufOBQ/6Fn3Y6odcv0YmAUZBQTFVDrO1oiU626jU1gNqT4eVUdhaq8Roa6hViK1fBjUDYY
FenK3gZJpA6sQBB7BqptcDpaxjp6ujKX1/cLwFNsuE3B7hhIzLLjIu5hedd/F0smQHzdmPX97acc
bdsAlRTX0WRQM0F0CsRfpNb6kUz9/Itx2IM7ETQHyTa0H5Qce0QlOSK17QiFRyz6pqJoKJcwJXYc
sVjIKoYXha3hXHA81oG47sHm9wlD7a6BDcm+KGpXDEAdC7DjTLL/8v40utL4XchP/mVT0oI0thEG
chB9ObwINuAjuWfnkXE5UMycnOmaX9/drQX9Td0G/hhGCsin8lHCiMrUXUZF0qwnyKCEZNnN3CiR
u39QDJoZvP/Ld7yTKBC3jAorW5tueWeuL6r9qE98N7OdZzc64XzCebGsruATNXhFe9H1tl8mEUtn
2JqzxYEdt/o0gwrT6IqtS9d23+gIje5p4gXhJ1tekqNFMfmmMK/GF8W7d4s1l624Byd2GlyIF+1E
m5ORcAUSP95Vv8/0S9+L39Gak9hKzUKCAwgHvL0nTDVQDm+tI7iVZ+7jtXrk5G/FDo9N2cYB1uaW
USwXhKihEqUZv4Y+xRB5GGaTX1H53XNfJsIIpbPdxX76x8Hcf7ZIL2z7eQBE8bfIROzgQ4zKxqV8
nc4LlKvlvOFhm93MVTfbIgjWjWb/9HBAFf0LBEfvUd2nX4IB1zPpNtIiOzWigV4/JqyJa5iUFwwK
v71ZIEg0AzZ3EvSGXrejGetEPjeJdsufBoVXSLYMl4SXf9RvHRs4HAhG7N+ii5c1FkY2cpSYe2mN
1o9uHWuN3uwAAknMWpW1MWtrvrj9cP7fikoFY6YoUDlg0Dx+ON/G1akzcJJ8MFY9LgUPrfmN2ggo
ArIP1US8gMXcxycKseYuAJatq90hA5TuVwazeCOooQm25GPxldpcqgm/YhpczQkSGHCbrdKlSsf8
0kfxOUtt/PEIbGRGSumQ4gniiJgF3rDJIGl/ECP1Y0arBT+3nWKdVq3+/hfyjDZ6BOLPG2/CzHU0
5ZlfR/Z2ZaWQCrp8lOLXE6qJzK9t18kKcDsJeVMgPNp7EyGY01QqaLm8NECzLK/FvC8Y+B4AgOLa
ZDaD7AvKtt5M4UXaaNYY+wHUwO4x7mC2Bl7e+HZQku2Kig4cdHJo66AdrMkUZmDSyFdP2MVx02rs
QMBruse1u+d9AC5Z18RjKjDzrob6ZP2tJttbzHUoC50nw1+kORtDpFgglDmycCSoBmkNfNta8WVk
pitc9ikjxjVfybI7RIDLlNZY8C2e/bWShsS8TMIQyDltI6DjgqeR+v2X+GwZ582Nwe1OgApR22+E
x2LD/CvFJnivKEW7YA/ojuf1MiGiKH/zjKKrFJd0yuSyX78Zw2WjSldOdi9rs859XCNPap1FZv5W
JPwi37hy04SYzyU03Lh8btfjTBaO6hby2mj7ZNHCOlt4vBg7gdjWYL2PJ5qgwunMJmkVJac5qmfF
sBv4w+H6/n/6dbeBq+SzM1cdZ6AcmnF8GVMfXPVj9KXVKvrWknIFioYFAZi6hoRkaNs3tYOhM8Ro
R8ffFeiA5NNnMFwOD63Z2qv1QqxLeXwEMxkEmNONYbjEyIV2r88wpDCHv9gXvSl18/S7F+IdG4np
sW/1cnpkyH+jYgNbLJkVEXl0gH9iI+78iB5SQ9Ia7lfq0fEfeLf/EwopyGIPJkNJIOdXK8WH8iXD
wXmODvl14Qwfy31WHFt9bRB8RfWlVjysqm1MhXX1iuES6bzpqiXpQeJn4zeXkh4LYQ/dMPxORACw
ohGzKY9tqCP9i3kHhq5hvMpz4L4grpNGHxiXEaI739Zb6LnI/uN9f1hVkLPoD+0tJDfpuar3xV/4
T6XfB4B3qbtF1Tsu+BGS5pBdXB81g9pXBh3KkXEFnhD+4gxwmKBhAqjr3fX0jfpYQ0pLp3x58jJt
8t4FSc8GNQ7ZdvNweIlfzfIActN3WYjnv4/BAzG8OjYhlG38Lj+pMaKJ66uVMrkQ/ItY0bt+I8tr
QTakoaqG+AvEJyNXdHNrIaHCcedwVBzhLu4ow0KbTGUK1EFBPO4zmejhi44sWsjxZ3SUlznqZGum
L7KGgjsUc/o9Eh0Z2QMkpdGKAZNArbIKXkR8Cqc3Do+4kHh2DGyCz855abS4cB4EIPkXLE3GTmBo
9jq4B2843SDmEHB7z4fNXZ7P4M8ZktBovTD9e0VQv76XZ+4Igqpn75vJKC3V6k4xyAm/4abcdqrh
4tdURiBMOE8wKUspGCswjbSBhIJidvwn+dowsiwhOMeHKwqpYzaeRaQvXh5FTupkFPBQEDVf/U7i
yriOYisoRIoh7SW6kpET2kHF8jq7dFXw6gwde7AgMxyQHjPRYxHs3xjUFz2VqPRpO5BRkTKYpAJc
o36pI3oXI01sdLMBk4rw5DCmwLoq8Z2d0dp7rrM3QVkhfUG487QmQld/HapR/ytUeQ3Y+fRjroJW
JezCq0hXCbuOn34i0zhcIBWVQMf2YSXgIBxXAwC4/YZTHGSshoK4Ae5nec5wKQskBD5XY7Vm4kms
apU9JIzzkaRE79D5Gxb+OpUz8qWHrUcCa7a0WoSzKa/jGfqDVRyKNdzAUlJiUQuklxEWtHychXxM
cGJLViO1XFGCC3MmP1fr+46uKCpxg6AkyrfwFwSAt8ZGXrUiLOGssq/gfvegsWnvvtcC8ggawkZu
4OYbCO6gFQyRBzNnuH65pzqz/DDhaWy8MKOzlz4avywZEeDjYFZbRFcEfnG1xr8MoX9/8YGq3n9y
Vl3k60baAItSoc4NB/+dHldDcXaHLSVjTIgtvDYWFG+9mAusKkUmry3osJ0/LumHU2G9oIwuibUv
KfGyJY0BxAAd2ObNA0zC2R+YThDLNMiYjKjhhhrXhBWhce1lfEzejWiZtESVejclrzHsfw1yFtP2
IRb1w/XxYARZNbCdqtIrbLJszHuFohM0Q9KtfYx8Tz+6Rg5GrleSGbhLSE3FzLVOgZzsJY92SbwF
5+/BDWl3oCGV2ZeiAn+k+prK/4//6cO/YYpyvgA/W6ZdItfHBcV3tV3hEvxP51CrHGAKBPGBfBoV
hXRv4H7+YMkmEDS+sfHTqLxTkcpejUXq7Hx8BelOvzaMC/zMw5OIc0Wcq4ggPuC8yunKWMHFaoaO
tjKkqczcucH2WmgrhTYZgMFi+0UaFFnWdNi56DM9RxulLNduAORvIxXdEMU6ZvYlV0VBvsVQjN02
WU+t5HzXD0uYv7BP8H4kVXzFGc6NrnNuJG6pIzLxqjk3EixjBK8xO2bx7T1zvGy57V5B6cFSO5Wg
jRD7x57raU9lHOrAIX/lDwgVxVdJb5atJ6mh9XAFW0h6JLQOY9qx41WBdRfVEneno26kXbWDJtzP
UY6sHy7b2sHCYrbLo53X8tJomRRp9xZFJJzxbVXKwasDwvXWaqhrWadpIubYL16OPg3kyXTOhggX
Lhhqa/iX2bFaURzqK5Dtfsnhm/tVxgdWIQmMi+Rde1Z2I7boHFVAs1Z2pTe+wUa+ZItJdvmO3mtW
3oYdO2pDfhO8hhxZrIJoMVLS5CRMVPlVHz7okYdDCx4aitGG9YQRAGdUow/TThQvqoVKd5VBmVn1
FDwgXTYYqOa5Xf4cw6NI3m3GXrQMSeuStoU5ufLFIi4rb0B+wfeCNIM7R62nQVPqboC8xzuknCME
9n+o0DLK2PYdEerE3n5KAy+dRhL4Kn8a7RAMx6nlAG+zGGEmvGXuRt0hYLtHGwf985httBoLLn/i
2nJTtZarc7AR0T83neaPeyOF8frkLNaTWum3cZLMSOmzjc7m4uQYTNU+LDWBCEJQocRQqc3msA3h
gD3A+yhjgopzI7cFae+wzUeM/bEGkM8YoNmDfkJSrlkpskB97GYk+YqlZw0sFSl3cgO5CcrCroQQ
miG26E7Q3zYx4hMebyN/i7xWJHALsXLk7lajo9ehOpGfy+9EZNxxR0L+l2HsS7JCUxlUFUK72hjB
eIKsSX+7KZiR1He+kafmn5euQbsIdyCWUdlw2fJtDEw1eUtyq3geDyJnepFsO0fnMnB8sl9NThEw
bpB99EACHHBYnQFQCMZildUGILngaHKwaapDN1Ug3Z1ZKZXyOZ8Kv7cbD3fzpoWSkyAXVOJhBXQg
3oMUKy+ucLF0uNuF9YcFWDL1F4jCl9PDKi+px3uSFWfN1O7Q0+Ma0zGTCxGZn9zggJ1xxi83rp5h
mUmuLclHph1VYEvr/UDpmt8ERi5kiL5UFqJYEAYdsdxSVJKncMw1dt5nabGWOXF6vRb8a2gn+nng
s3N1f3Ein5P0/CTQ2Tn0TBwIc6/mC0z/97Kqbwyx/ta0goWHDr1DHZbYILjyfvP6GYEnZ/nTx/Tw
PW4UAn3HXY4rfZeAVSeobfGQEtL2Id8NW8vzr+PRLb+WdIcJZjbJEUYqdOmWo+JuZUx/UBAkGZWs
sLRT5DP8jgUbTXFGj2UMilh9WDc4uj5gKKyEH76iKZ1xDjiF/2VC8wrWjcjNcf++SAKFAnNJs/fr
S/jYPesHqxhDMhLmlx4XFD7I9AhTKP9ec/AmbWzKiL2jTO1plqzWJK34Yj9K9qQwfXH4uu9FHO2T
RfRhEFhiQNjLglDDdpqY6flt1IkwlLr8Gm2xA4rOcLccAOkdZPo1h/mjAIMzbpehLzb4CmZWoqHu
B9kgpcnMiO10RZeppfNjNiENTuKXUpyqve3bQxPeCVxzmfYNPkkmgxejgaSDI6xoZuPTmHRHnSud
DT+C0AUDwExEOcfo+pckeJyaVju7UvLz91/wBic4V9o7BOun94gOzapCDWK+ucvwOfqfB+Lq2EnN
YB7p0hkcGsvS2/uBtr0iwy/EET8dIfUimqJ+aKkyt6K8veAS9LkxLm/Tb8RDbBU+kZjCsOVlqOl4
k6L/GGxrNfiB9I8SQyijA9SaRpdDvCV2CCsX95hAZTZk2KvmJ87wvxa0IvoZfJitpmsDjC5OyBY9
mmfr48fk3vjcWTsalB8CdYbtJkYI02h0AEJAbaxH8+0CvVXtEfrweyOlCQv9BR/hJKKbngGVIMAn
Kx2MMhWUJltIkZ0wZcaJHErBBG41GCB6HXLmMbbYaX+HIqqxmLcTd8XREQ+tGiRRXxCVKbC2z8nG
FxWcnPtx0UeoMMqxVlptL1GwYh5Ghjs/4uryY9E1n0gIU+k7218L7A/G3Iz3Eilw9pln/i+MuLT2
NGI1dr5p/S+Q58xqpHl082ybASduJMwBQgmWT5gFw3Y9g1kdRQOtcAvFn/JKnWhBOz264XWaqHEn
zQdSKXuAE6rAxZTHiJt19BIYyn3VbmxfsHBjLUaAF7Ln6oOZFw2Ryr2hGSKQF1nDWaPthlo0qSjR
jnwqLlIIMUkkpROpZH3qC9WsHhlDslXztNvWJlqw2fF/vQckd8e0wN04UI7+fN/c0wlyXPLiZ3rS
lkyxEKIxh9JiHpRsTMiWJTYGySk11xkipvNR+rqLcXeNR0lGA1SoJHCa0xfHHZc4M92QLQW1Qlnc
UBCc9tzWGW1gLY0vMOdWGqhFPbRIJUw5yEbWB+l5+785j+Ge0TARBcxoJPc9MtXKQC3MyKnzZw5d
bvQJrFSZxRe5mBLJdZCSKFWVpXfw+dVuLFMgDEehiMrnSpucYNAei2CDsQNcKkiWw3+4tjPQCbAM
2hT0ZHd8brqLhXcS40oprqEv6NHzL3AEZvP5rcM0zkIabpp618cWnANCJDcgVMJld14aAcriTBPb
JAFTv/VUQ3YLrT+ycQGnhIb2TDrURSzFrijZcSmM4mHy6DdkJkkyhgHH//G57gLlgTM0wc2OC9Us
NguqD5+hZ/o0d1ChOyiBbwcHjC3c8eW0m6ZRbuHrRJ6qu5+r6M3pAqyy81dnwwuoPWa5KGULu0qt
9JdevCkzO1kwbHA5Igf8apOwKBnCsJcGF+UnwQKHJ5sAu8117I0PwJQTgHrzbQiBx9OBySepF9iX
4mpRwHUvPZTARTQsMYzcfqv1W+w2K3QJqcPeEVneV2e9W/ZnhJ7CPGTaPhwRhrQpXPgjst/mIwqa
JjCPz5t+lIq0ItaHBvPh/0o11LbLBBKiF7ciud9UnX/dTbD97ckxRbpqne4udhIN1F7mZYgIwY3z
kyZeqf+RhnkGmG9JhnUDnHisYz5nk9MZIRQ7uYfxw8Qe4deYzvK873MFOi/b7mNCUSyh+8IZA8x1
XVQU9a6/RNlwuOiLlVvQ341KiKhBidED7F8o7Cy6KU3flOAXQCpUaSrd0qpU2teoxrvxplWl6rIr
/gVhQBK9mc7FWflsb1gUoy487+RFIG1uCFxCbZaUoCYedMN6oyD7QOv1bzUOECZ6Tr/Skl3XmpC3
h1Akbg0xwTjwtvVsnwRdrUFCq/2eQ+pgG1ImX4U3mlGo5T5mEzgq5svYqgVzWA+jeCNcQfeeeI/H
HdWgG26ZLQrBry9+vkpsALPgsNV336lyDlbkGVPKtYyAXU76WweYYpggGw1+fyPxQD3LJDdsag7E
6mmV9yOyi+twL0g5Liru27tGsWZdeJe5AN3+g4/6paDDd4laO7VpdBT//XhqhsU+0/TTknydSZ15
OCMw//FL96mVl5XXjcoK5ZyPG8zkNK9cS+2pJCwls9zm9KhRtCLl4y7WrTciW3+xdhcUs+zu+uGI
5gliCixnZulCX+65121mnnzR0eGNMnm6krH1bw4irIyrHSaMTraCOvswrj0xgj+B2RsDkMOd9xZe
4PAmziBZxCOAt1Pc4C4pve+q7kqiujDtzPnIIpEUXszQNoXXvpR+kIRS3udKpDtFYUGMldS9RnMc
ICM3mR51gP3cQTnKuOhUQd52fAMWXmbf8R8jf0WXDB5I8ID3tDdl+EJQsdT7r4w72bUryht50PEm
AeurNH+bPXlUZjVWEGO9Nbb9jrJUl2Ta8b3Pr4//M8rdkpKxL6+aoTfdYukh8rp5n1qvvzTIaPzf
/oMaA8tgUlp9MDur1lkuVThk0avLqWM0UNLo0ZUZ6eC45xVDdgsmIZMELxfj+75HqRenknQdmFSF
dWzhzRa3PoLKvRSZ71aPZ8kcJ0PFA97sm6HNA4yPPoubv1h+BWOrwPh2W0VeFL+Ky3PY3iKEKPHQ
cvu45YcUEgdB808AaGyoP1EF287ua7dJJwVK+ouPhklXdN2keWFS4Q71QssUIXkmN5a8iDgIvEry
o9+PUr4Mr8h5RIICpWWoPn1yWk0gf7IXvISBEX0HAi96cn/dOVqcBf6G+jlOCs8CXyZKUY7/gc0v
CoNT+au34FhIyAKlSexTxViPLXlwTSJmEXdfcYYToYegXS3ILNzIaG6Jceu+Ed7glbaEDnm0mq3G
Ta5a97e8DUj0EyM837w9ZcFROCGaqaapMKMS2qstOPBa8pFnwlCY43837cSXEX+b3jevCONgLBdv
y64exoGTsmlgef5Zqd6RyltyGsELoK20BxU8sMHdoJ+5U/GyvOT1k30M3ammmG00qJVI4FOwKuRQ
mTEc7sZvHqWQKCo9i9Dc7nrkY6+e6JndmRxMn60qz58Vz8AWQyNPkJ3Tc7bA071RPIGLrGEJ7AMD
3fNVFXe0KwWgKBiRs1Rg5fewFbJARFfUPm0jHwJNG2IDPLUdEzNuRu/mXz/y8t20MyWpH0N2jDF5
lz1445tQyUP60YBZaoSgvEqpgYYOa+CtFh5GCnv7FcupvQ/R0sjI4wXyGwCcKntP6ZtWvuThSyjB
Tuaq/HaFgHvo7wBpADuGOSw+bj/OOm2T9rH+6dIVz052vbixpIeuHd+a3LkvF+YFYsM2rUa24Cmg
ooIjQ4SFtzYJJ8MXoGheqGuyH+NJY9M3cHdcbhWRKYTuXfVTggRqgfIZcrio2IfbTsJvbtTN4oBt
Rxm/mMYkED/qx3GfeelJf5mowEhk1mlGzVkLAVxgN8P1+rrNxXNMqzJjlrvrRggIxMkXT9PSBlfO
f1DyTHjqC4OhWmKqS796NB0i/vwgH2VlyLZ/ZELSG3EHAFOtN9nfR7PGoJ51Dq2lXaviwSGBQ7FH
R0jcPDwQ8nY6vBL5pcpLVjWlBT6eVgu9h/WCZn0BYBbgtSOKAdYRlj133Tl3VDiYh6kY9vcPoz6p
81qmLwiGJ5cLso7Ma1/HACvo1axgMn7k4e1+fP4TL7+mTufjKOFgGYpwpf5PUxZyBURpedZelHL4
2MjWMkeoya6OUr/PSeX6sbnKlvmH6RuyyGEaPcG9UovYWskOpMVfX8kSSAKyjUM20quStFj+u5kw
udNt5vAiZLsFyIaz4aYZZoHC1whIWtCTY7nA4rXqPsi6bDvNpXALEKuP8YLT2n8jDeJMgsVN3eOs
L3jZS/qh1GSWJ2N8J2Xk0jiTGSuF26bwSJwkidklr+LY7OznKQUbD/c6YljckcEWOTKXrAA1L7rX
Z+Ea2bMmjzWfKQtswLL4l9xBAkNAnAzfQ4zmGJTp0S485Y3WkivYDg1UJnLqF+m8PsO9mDmKJYZ4
DqdMO6b5inzD3iMUo+2uRGQpoAn/QQibBZnuz+6oYroSy4lezB/G2PSIOVEKe0K2yOmM0fE3pQ5n
V/UngCHgPiS1OVVB61eFXjmrfWKPKHKLKBW9CXNigsJWR3HHN6KaWaMXBzaw2WI0fExkPTnmmwa6
9vwopfmfgZYhZFiLLoGgd7x3854rfAY7MorD5Jb7fUaPPciY43t4QUC1e15cvbtQwfkleV82cNiX
USJET+4qpb3dwq1IJuJUQwe85r5hKz5NzL9A/khIsQTS4hPdRA69lePucDS45ynXMjvcfXuZBjM8
i56mWy9VcI07KtxjoChThm7CfZChUwLa7GOUxXzg9GxaZ57/VHVnNFrZcKOg9pbLeq/sE7kfpB4A
CnUJOnO7ueYQ8Esufs8U7p5p5E+7hwBFTfDuklOC+6WkKhOqW3DyFA/0Qxuw9YLPcsJyEx1NuIXr
e9+XlF7J3h2pK8Wg9GSWIGT30pav7cgKgONF9f2YDdewbYkyEfGYzvdnwoySyrWqteNEOCnR9+Vs
q1DeWSiGufxE540FmyPJN+0+0iHEo5H30M4kfW3Zn+VJJ0iZxO3q/ibCHWA1M45BLVzCLqfb9c6m
M8EaXA995IhTl/YEsWi7imiKvZf2Kb7jL6ld0ddtAplZ874CpqmpgdwTDe2qKjV6bFVzOEEqzikC
7JCmc9qiiw9c6i2GH82LJgKQ9J+E6PVJCRbes2cqKxCJMnFWOqBnfYyGZ6aErsJAguDCkdU/JBHS
1xL0F8ghOHFVvwywRtbHGbmTj+t9skljVpyYehItsDoK5EWP6Ga5Sn++x/TI4OP3Fk5pEm7xp8Jo
2mDbRjTBTpVAqVfISv1I2uDvGV32dSvA5pMTldpnYfuiFveoRcS1dlRC0wr34OQsHy167dqH5AlS
tDoaCAjqZ0DI/sWYid+he+w8skJwJpI8IYBRzZ6CYEg7uPr4h3vA3zIJLgL8n8STrkEW5N7kw7xC
qoXbdu5F6QssCzbcR+lFXZcS1/qoy/9i3Ahe4T4xWgHk70ZbWICJB2nt6CVL7VY/jK4fad9m3YX/
O2djMEXIn1Vvg31167NejmH3FaLfkMP4yG9c1Cw3LRr4kIov1co27QESIu+aPKaqfe18l4xRzE86
M6dggsuKvN9vH/8wSJyJsRWu5M64vU9EKeVbc5u33nxZNShAfYoPgzC2GmrcPMQ4UQISQ/Meg/wN
dEvP/JAM8rQIAAiQ76HWEoh/WdLtz4aTiehOqlS05GgNSv6RVAEBN8cVa688rVSQAKVYB8qw8tCF
4iAhDtVZxNaEkjUOQISbfRnjHlkFoG30RHdgd5ykvC0b+3ylbHcPCxZDXux+BJRm3ceY5LBlbO/T
ui7p8cOE3+dGJjSJeTZ29mxWQkdnwDoIDXMH9r5bsPxe2qc9+6WCvJrIwaxmPqR4wwqQF9om9BdQ
zdQgux8N9yFVDzh7a8XP7zVlHSh/nnjU6h8xMpip7LPEK2rHs6SoyvaXk6ff3VYBVUt0gfx8m1tc
ZGvabfaC5pnvHhgKyd2YvVJHrSNG7SMzoV7/OnOONjv6ymtL11Nt1nE6ZZTRE7iQ22cMHyIwhbY2
Lngs69aUFch5Z2tLvBchGoytY5438k70yJMR/Oa4iZ0JkDDcAEQju23sK0N3+iixqTk//O8HneQU
vo1pjACMmcgLcSSvcprAsBlhV3PUBPYviWYK1kSvzzEoEDUp/lbp1gWv0EmmYYN0Xs+6XfE8XAaS
sSzJahM2W0KksP60PV48HAQhekCgN+ZQk10mEa6sm4vhh/8c9s6i+uzO1aIPgJuCJJAI6Yn4Auce
+TOrkpzsofpbTpZN6BZq/QzvFnLgJ3jpJb1+RzZavi9VBeHUz+P01gGZcAbPH4uGpE696Il+wGq7
ceEgTVYQWxqCSYTFvS6brKv4Obs+MZqtWQGT5+g7LnInmuUoSSDrGokCFAjZPK3LYCvtK/7DHyTH
hPC/xQm7uo3tZiMDKqZHji4gRpquMYiLppm2tKKRUVGS+1mu41YQ45jhG4KuFc9D8Qj9qOUJVjiu
kgBUd39iy16KUVwsgBPJ0O3B9KHabcew2gBlUs8mMUCy/k+3/OJ4wWH92Cs6Y5zq/TuoHOyYV9O7
aw0Yx1rpaHJbnRkbnRnqHzWPffF9pDy8ROKf581rpYmtL4Q3VPswBMEnD8jU6DHhMHLtJos6OM6i
yDBJcGZy7qtDUR2O3ckCom89oQXS4p6s8HmoFEPKP+YFbH+4ufUtkrH0dmf57dADhUvcxozM4bni
e1RuaW4QLWcLNd6GZGU+NFX3isVdx9fhWBzgm5RCKhUoK96H1X1QReoMjEiFdhvS6q0xCDSdin+z
AUh9Uzs7CLrp/zk7Ve7/TZY8WVmtQguDGe+5180souuQgsOEqs0aK8l2rXrcswkFh6FaTakazwfV
Nu+bjybVYuAfoIpPn8TV8lVFbduDGdkfCgrqh/zG72iDDuf8r9G8aV0Mea8BkAsEwO5FW7J2PEvI
AXE/6XG8mvQ8X0x25IXCXagYmr88GWD0fsxwGBE6/fiS7M+24zEUpuIgLcKnyXXCz0Fsk0WtwI6P
Q7e5kLuLL3ZIqdm1ZfUxdO/qQGwGbWAp8BHycIPoyO3V7tpaE13TL+gsXNtNdepKnvpMNbISz6TN
ZiuXdqWaLDO4AxHcBE8paC4TO2YtyAbPNEjjLmnqjK/irz5Cc6FI2t0wSOYu3ioN/mGl+LvdS+CR
gYaErAJVgNtELsfj6lZW3yTlHesx7ukGEBAibGpveZGii0vHUL9B8WRpU2unv6EZbPmNxsV/6muQ
aVhlfKC6bvjsx0AYmrcNF7n4xgE+9S7c/nY8KuouNTVL8WdA4JNXbDFlpaFeeNYLBVPnIWLLXE1L
GXISWFAPcc0PHs4FSVgApCA1LW432sisR31+G0LeVhf/M4DYpLL7weVwR+dTZFLFLwKTP9RJNV3a
CP4DSIMquGEPf6bB5Owedp9f2Cl3ifXKwfVtz+AbR7lB8I0J1Xhy5ynNATvCcAKJqBlLFhpTiq2V
eotJGtS1C116k9ilmZcPqM/vZ1eiRxwZK12I1k6WHJAB5CptEv+tT1MoquHImiV2rT5DjgOIv9Qq
5bQ21/lOBtthS0tKJFHSPC3P0OQPUa1E0AEH4/SZqEbZjq9ZX5yjlFZ8lpWIhh5mVGW68zXOp50q
Zz4NkCWlj7/bLlupVBNne1n+x/rmjSvUT8/NvGoU68snsa8WJEAeY8CQM1jUICjiv3dh5VBngJxU
yipO0ezXhERjyepqJU/lIYpiAyfMQRmBT48kvVZQzGvAJG1HkJtOTTfwXhi+Jzhy+qeuhpxM0oa5
NHrndfF9rIs3603dujeJb6V9UU2kdguQo2ikg6JqkT4q7/SfqmFw081asPg+tvrinOcuciXzH+Ic
5rNru3humbRt/r39LIJmrpxkW3NfaOn8hH1IcigXo7VGnS4w3w2ILkhRBB/s5bPZSbUJ/S4j91AK
uNKd53PYz7MQ2ep5zxQ9JQP1eq3SM0mtPAIV0fCE1ZmqQA3kULNGEdW0S2H7wWmyVUEqeiL2rHVJ
NupQYovzrQKoxA7h7Q+F3b7MNy9w41dfaHwClJZD06m9J5YBGJ3m8AKd6i9J7nRnx2a26fr+usCh
Wzv1ElLVTDc+M7OXZ5YNKqgT+l7kHf90R+qosiJua+VZVkm+LHaktezLjxZCtG3oiOryH4sYiA1T
G9GBbkWxAPBZWT7AYyuQF09pVIYiIeDVyx4f7JC08zSRP0qEk/qToXKjyr9I9HJs4+VyeG4ly5th
DC6CZXssCQmK2MwS1tat9/xmSF+CoNa4HqV5yH0SJJ6LfPP9HVzk7jDOHAxtIfUEo0yazCgshTyM
BlnLaHljtERQ535N+EPYAyTvWyS6Mw8fJ0QIdv/FqcOX5z7iWrKntcxV6twnhgPsKPvskwWLmU+h
GT2F4m8uXLFJv4DbkiYb7TuKCOxHKaMkqz9hyIsNsOP4KNensKXsLACfaFq4ZJB+hMiBC45XqM3N
cYmozbS/6xRz1p10VZg2NF1/fZHoQd6jkzTf9pwz/1/gK0nwslpE1eQfns9f2QqCzNi+mu7O14xn
OH/DKaMm8qR+pIMS6uuOy3dYrN9XkTXVcSrR5vifoH2glMs18YYdlDMutX7B6vvmormrzME6ENo7
lpOUshFob+INHzcRCeHYtydbzE71KKyXZOPfgQ5V9H8D3/xuCvg+HEOzmxoMT4u39tdgFv9/yY3Y
aF/LJehSA2pxJ055nM75YsMToHL2rf1ta7YnbyNLmMutAuSM2sdCvodrDY/8b7ktI50+LLgL0kT/
5ARWf38atoSd1Jkx3ynYPtyB/rS6MdJbH74bk6O1A0bAsH5R0gSiPlP5X9NvF3sdoBiARZjXOAQp
643EXIFrWzsqNpX0ZObasu6RhJvEKNiqHsML+4jd7sCO08G8mkwynRpxBi6dH4S+ptIsUwY2hmG/
UAQfxptSEmnha7RoVpvyVtGu1ukW2R2oXrG9Ab7gn9TP6HVdiAcgsx47A8mCjFVCid+6HEbINFFW
lt6PSvjatd5k7H1pQ4+ffTlQKWCUjn4izIHDFH+IiSkHNsRE70cCe5ebu+hSg+MTB9yUnImliysO
lEEyl+YEj9jLPRoya49Ez/NI840Vhx66KVn35NZHU5lEdjtIlKzTzdi6y91G5zZhqPN7F4iE9wH/
ZKAegi4JNFOQd7KsPMuhhFtuuuk1z6IXk1PtXGyuafy2GuwmR8PYV0Ygl/+8MvYNyvODKwS8yp3i
2AreN6T5umlUV0nd8FxVbadLgTSGew+Ic4LbQ8Hubap9qmCy3inf9OwLahzZdNiGQR7gc9aBaH73
Ps7dA1Kl/+Aa54Ei192lvlKtevO1OIht6zUSw7HtR1iKwB1kpvLN0mHEjKiLaTG1UjYJFHx9uizZ
EdWoTAHLTpJDtqTvHdfvpibh7h9H3zv4WLHW501uQltzw33ROPeS9A42xbY/mjtxaWBKyYOB6bSb
AV5VnF5qn5QNM9px45CdbXYLpgwniQ/cgMD8Df6clmxBouRsojCUrWV8RTO8ozBBxjPdDn9GjRGK
q3VtOlLkf+8pLVPfq2OHpgxUFB1NRWAlN5hqzlZDoirD/46LyXvYw4HC2bPp2U5QBHSB1pRxT/Rh
n5j1khy6xDUQDo7Ech//gHj4J7UK3jF5nVkxRTxV01VHrz+A5fuT5FXD64akkIohe5hk0i96K7jg
y9SEN14uDp/9gZTe74c/k9YvlMArHC3qunzRWVbJ4SJ3vSLrkeVeWkBZtHITe6V4wn9MyfZ3Uc3K
fQcGVYpjbbcHLqkBlhcyHlCP8sd6U/IMNMSEEi+eKPCSYRQbwsmXGkFygcaV5ki6zIoJl6xBGz5j
80Jy7xiNSesdBpS/qnqm5nv6f/brLhtoG1JsHM8TeYr8X4dAp80KUO79d5GIV25xy3vTvrJONTMS
ZWS43XuWyfizHEQbq0iDXM2tLnCZpg6qYsiANhOasE/cb52ID20I3FhtDo5+FB44TDyDJ/l2j3Yn
1cuR90lukHZ8qhvcFJWowXSqcBiK6QPFSm9pO72f6Ltc2hxapXW9D3Jt38ou0uD+OtrtkkmM3ilp
7tyrGYr858v2tek6KH4TGUuN1QJkMnCSxj4Pz4+lXAXDXjcXuHhfvkvQt7MLHoe8FX5M2T4ZCuWk
rY3kuf9yhGA8q+Q+vnkz2h987hxpVzuQCxLU2csUpFiHkLpHI2RRhx0qokH/4BvaVM6NvxnmiAE5
nqf6AxDRbIFRMI3d4CthgbD1CNRsDVxTLOI7A3Nll++CtFVy87AEl7yJzOQXcBD6oJcPbzkELjCv
u+w2nGXM1pwH2F4HPiPNRusgMUd/lzVhDlbhiIMXR3kJWEfIw1azojv7h4qXKM9jmO6YKHOI4yRQ
rXcq1XGwfByo+rnvc5wWZ3iCEK+lxjXdrGJgec349BNwVD/SuZr9mi2IyFL1Lp03hzYBc4c7djv6
6mv2zVgfpcU0U7PaafM5rIJRTonDWR0PS2zauTrcSjKTQZacOiing3s3KozyColVr5eYdNB4UNcZ
8i0TPgOHa0dHyrGFx6WnJNiJM/46xRgwUoQZPJ6ZVUJCPxpmk5QhkApqpEwPIqxpwYePwSLZ222N
or4i0jdPj/RgxoixiLEmgNd8XyquNfymlA+dV+EEXT6pYxWRvPBwHiiFHJMSlU9wpf8dPpXIYfIY
/6+WykMy5wZe1V5HGbY5GflUlcUjgbD9ViaBE7wtUnqLtH1tbgaGND7KShhqzQBfRz0gIt8PXLvk
RTPnCyOk82Lch3Gs3zlh99APHdu8OY6HAGL8iORgMFbvalAUPRPSYvppEIg73AwJx4qhVri9tWM6
FUqfnn7o0VsKFK2c4cN3xa6Znwz/GyEGq8Hsr8kOBVPKCcJA2XruCqcn7xkmgfk7o3hShzRbx/qP
pqOA6IAZgIy1Qxb2/ODAV+OhFoLkQ4u1a8VgN/AFRLzjI5CkcgxOeY1JF33106q93ePPQVhrMa3K
XEInRRaCbUeEn3KmuOrYgHtwTjnvcVd2ClVbRDWq/RJqOjfwfxzMa29CfbwEHD2l8xQ/d7QGBPJH
WpmPIc4Ow6UhQRrz07K7l5ZRrBoqnioRdZvPbaqekrJnGvzZatngM0R2QmKM9fuECchcs1cUWUch
QeuvMG8uMkBACTkC0wNwfCBkw7sVj6PKyFU+VEwDGhDYotQ2ncj9I0P0mVIQkJrFZ5rloDceSbj0
pH7OZ7EIupY6SgnjYNHvgJRVreLfFa2O+R1+CRqBPav13Rm6LNu1ZIRvimEvJHvTcI3HKWIAHndl
/0A4CG4F0QQlamSYRGgsS5SHTeoujc74VOCJAJ2bNTGFT50vj3/fbvyxnOfotzlPg7vHNHxkyO1Q
KKufE9DCiF54C7SvxAuS/odEdTTYienkx71Wsw+jAc5sEtbRjxnAem8QekuKj41wrumcpzC5CbM7
kjrRxxN6iVlde/UiGPxGKa87cZ9uHOjsupPoTYb9kZCrNYcEQP77YQ1a3Mv3j5O5OXr7G953Hzz3
xkhTQKo5U+oFUZU+oyJlpmUKDZSMaGA5lZKI6vz/3g+SJgxxcZ0oIxUm3GdwLuLdre35cTgXOSYq
WiSUYlC+lNrZrA+DypfwmdWXgxQrEv5b5iVTMd7Lz3nhf2DcUd9eok514zf9OlmGv6cYsNkfkoHU
IsfbYjns38yghEvmeHhnlWOw5eATuK6Qp/KzQm1fvBeIZgoYmqYegmnQAv3tQUemEcp2cWW9z+8z
nx6qd1PVcUHyV43UcMDWtE6Lj7AEWLYjDmsL85eFHMZKM1Rve/Y3rOo/Nr67D2q58WI0OCkCON0r
dvQnvOhmJS+ZM7IOVfWauBBwEUupZdnNIJJVe8nf9tS76iB1zzfO1Rdr9NW/WZj0UdlkHJLVmy3i
h8qSFf1sM3SDqyHv+tgkEnfMtNygpWLq+L7QmfSEtA7Q5DChTjno5dl44LlsyOJByz1oHfOWiUeq
HO5LNwe0ggAqUCuTCyoVqZRHTICq71wIfOcufjAL/LjNBudnwmMIoLpy1Q0Uj2WsJIldWQYb1C9A
V4MQ0XgG9WriRedfSWapo3jb/HHfKgKVH/CTSiqRbnEK81cv7z4EB1decT9404g/DjT4ziEpsOVE
E5UXIB9psnLc5zG3d0d/rMkYEhdi7QvWlH0MuhvmSPN3FX3Q/m0zzW/LlLnIRzqU+hZ9Od4f6mWH
70wMgNFCxUFSex/E9UAZmOcwbjPoVPCEiHdP5Kuy/7HgEMz57RCOqgMuzr5ga7cbyPOnJsKfZhQ4
pLVolZkfQSj7oue0XnW83lgeCKd68SaslnRzErKEcJGyxkLJ+k2gjvZb4OuWsos942c05AmCABxF
CDe3NPXNJIBoS7BsZ6rMmEDx4QvaFcyYALLAzZAJH6O/tyqLhd7tKqtW3/aLqE1HxpM+bWat0eyp
+f4d0vzkBjOp2oqhOScFBbjonsXVkwc6yburQACRpigoL8tJdHSKg6ah54ZxJAvP+DBSTzMFRMSF
fu3dGPqH18hft5nlvrHXkBjj9D5ZaibWUUphvnv0wlwqNIlVb5Yirrxp1QBexe8i7FbPskw2Wtyb
kgS4jN05+StLGA6Wx8Q8Uh4MWKlmULjiLrM4ynwJzMHthOMt5PffX1AguvmJB428yU7qvGHfPIdr
ZDYj1Jrp3xX3ZOZpM/UvMD8cx6NaqlGDbd02A4kR72jLIWA9/YbqqL95kAcJ5w61s34RJ2JlklCi
wi6MyjpwkwXw7jsVwkHCenTxfqkR44Z8vWNDmBH6DPW9Mph9L5B16rvqC94kwmclJWja6+Iby6XQ
m4vpnqyBVQ8ZVxrtJgVfESNzpTwdj+IZnzV/0r4zG4PKfVU/uLS3ME4m2DYT5mJXg8MlEMAx+S9U
gRX1OZlWGnDNZlo1dlnuHOIIMM3pwZHoyKgVbfgEWQwY4GnmDSn4SlRaw+M32JypDVWsmD8kgFFk
BVKF5uWHhXy2bKczWpY90j8ppKFqTztEy+ORvGqpc/+O1GDv/gsZLMvta6gUED5uUJSpZbOkBtUS
wiquVBGxtCgRBHJVTUI2wdT25SfofyspeCpcMS+tg+bj4gJ9vpY3iYNdTel4NePgxLst0Npr9ryJ
OJqh0B86vE63eBQr0RIKMuJUMdpK8+fgDhtfFQMFi/IUX/YK7S5DeXcu48aXdwRzuvFQgTC4zU+3
zOK/olWOmVzENoAqjwJT4WyJ7Kw53DykseSy+eY250oEuuMYSbl4EKlq2WlpTO+/gRKlENuv6VNi
F0eWMBdWlatq51SNhZ2qhCvbd3dnDTf5uFMNWOnAatBQ7tbRhjM0d1YJLxWCJPLjRsrUUP6FPhYP
DTbP5unpLpaAGSDsCfqn153HpSthb3TwpEoAdyRyqD+EQDvbUCLOIc63cYo6hM8y8tODd7exbGV1
pPTqAvpyARFUNpruv52RC0US5nZ/hg4zk7Hjn4FIadHz+rQ39BE+ip2jCpVNB8Gv/oxDmbjNgmH+
eROSAIK9DeiDKm89HfKUsPgQEYubJWVq9f+BBZdiCLzOuCM02FcO5YEa6UlLJce+YoxJFlOyBaGP
S+QJeGocD1AzZQ9nvBG99xhNdBd63/mUEdVXfxNf2GfhoVxE2s//8ZLEkkxGzTQIZw63g3wZWJH5
gnKlpmA4HczY4dYJLbai88bAybIT441YmzoORd4EOYe07L1b406tRje4xGImuKbJ4gDwRMEEmp1s
czdIBGN+Q7M2L8OLyNDazmMRUNqntjh47HJL4s0Jy3xReNc/TcbdQt2rhenXSK1YK4PmOG2tuBVn
kFMXwfHbrfP6T3F3fPcq7FtpBxnglHkzNZ6z7xAtCvoljL6s29BDUrTciKA2SPPbVuvdkLwzL0GT
OJkvByzTE6VrN+ndA+vASDvmY67X0AKQrKM2znHgwEdsK5tl2fTBl3x8XEO5qWg2GAHpIe65Qlj3
n9SuYNPtWgS1JJnL7YS7K5xyIUTnnmwq4l5NfV0bQrDr3XUZREsGK0nr9nGsK4css6PTsMY+QKa6
B9Il6IAzobEnSm67ib/GYAjiA/KcDo5MHFzxjd0DCeEW8buTmlQZYpwY+5Xjkh4GAZ9dJTf8zFdQ
jhddKqhBxHOrJMG3WfuzDVjHqv55nuCPYC6kdYx7Wxreab/arB+rzxh130ZzqV52fcrcKE53e6ct
AxT+L0OkMXcuxruXAIouvW+Nk/TiBt51WqEKzipychFdmU0HP8bDccbq7pK/Dysl2PZcNKjiMChM
S8yCAYsnjnjAGWc0J0ODMDXbeYIOMifJm0InFeZtFMvsv9yfBAEBpKl01/y65Boh1hnN2C1MAhGp
NJTYzw2KpNIXyp725A0JQgxtwHtHfLV3rUef/r+pj8YzUzste0gFeKsMbFqGMPw6cf2Z8so30RzJ
//Db856eLHMwLqIXVWV7yaM2YPcJUTy1UbaT35ECWr9TjO/XoCBYO/qIxLilG5ihQmlQ9EBv3AZz
jxKHL4SkcX/bvHe5enzl/neH91zLhIp19F92PsMvQruR2f+c8UwToENjUZgpFrLzVhee5IcK44bW
0VKP3veaNRcrKZxx7k5PlE49gMS80dpiynXcqAbovh2OHIuunr9DzJFOfHkxJrcWc5fwB7I3uAqI
Ic4D2yoeyLnOVb3B+apgmg+FZ8CCMUFa/ppHVORgjoOcnXBhJ1jc1DmH1GXyd1oeU+z3lyQ2/rdg
cEbDWNqWPB5xhxsU1GovGsCw7wSkA932RK3Pk027FxGCwiUenZ5NTLMM6MYOZHoEnNGD5VeoTnej
G3qiTUQEO2/6W2E4exS/jrvjwUQiUQnPmWn+zkuHoRZvuNelKwzb7KuDcAaGUG/I+mUEp6CZj2qs
6PjuELSHVO/cqVMb/TazGFpi9OX+xHgoluFAR44lk7eQzV5Sfp98p5Vtun8OV09TD0kwUeINh5D+
SNj4s5P+op/nLlwE1SXBZ8efQwL92tbdpTS5vzZtL0zMqLBot/s2V8Z9Hq45kdvxzqbdDln0CU3y
iV3s4JixH6CjGs/1v7NWI4VTdySKCX+/y+KDDhQmFfKo1zWVxFyRWN2HTE+UWfeIZcm1CB6ZqWgY
GAx7pyD1XmSfpyQVhLEwViMtcXs28d/s+9fF3VWgLCGiEKdOt/U7JJne6OESrHBw4ga6gcuoU51t
RXZBGCQTkP49AMcKW6Ltdi/IdI/zHVG3VPSkhvaqcllHnJA5CLYOumxystpNNGKzcIBC3UvwVluS
BvG/RPPcguXGs1AyAxwSy2itR8PrjUXHPuFEculovD/esSwSlUgSUz65QIa9S1xLBthV8+6zfrfO
JcpkVaZYOaIdqcuu064XqQKvRTW+ZWOD3QL1hQVMyRDTwxTRmalQ9tkOY88tSfMkH5SJ/14R7KNs
VV23RY3dQJUDZeVudrtGPCQfWOAnBHnGizuUFFuVi+sj8XC0J/LjUZbfFdgj/YFesdFKwEEAC21D
FjFemllYaJpSZp1RerDPdEHPcLa2jynaPKWywJA82GKA3dW7hof/wHq97QN3nd9nU3Em9Ivnopzc
hHSPSTnbf9MjXe8I+z6FBQCKEa2C91sNPJCLzemowalQY1Jwo2CEthAm2e0XAD4tCB7zqhTQ+xdc
Xt/+rt1LNCYegZtMQfshPHecdlxTiHO+bAbTawfQXySL821Y8TnnM8UHVZ4LUiGaM0BDafk8suLk
ar3eWWECzj89ccTbo8pp4qygj7VekSnAJioxGuEaasoIO/WtM/Gl3GtmPPWHPsYGSIUIjwqe8ViQ
Manup9DXJx9zOB5se7AD6hv9Z3BATbUbJZBEmIkm6nwPoZ09sG7ovzZbAS2Bb7H1fG+kvhX7Z4NW
CSPBxAoNuqCIKvUUc2xadmnLaMdMOJBJXjpePoF3d9XNZyXwyCj2OpGqnEBTCdyzq6SxXQedo9Xu
29Wwv25Y78H7TXSzcPp9Y1bvdkBgkwIjHMAevTwSxQE9J4kIcazr6/3vbRLE9H0QTdZsce57uFJy
/5RSrFu9xZZU+j2U3we6R7UiSlc+TJcWu7iSTOxpfFkbezYu9X0CX70+nsgCGzPMC5QETU5fTY0E
Mf4ZdHceGx81oDaFcd4oQC5DkO+4YvS3ctI7GpagALoTSB5vEV2bWonerllLYpJY4oQR3S6WcQj/
V0CeLIifGmOOqbT0F7iItqlerGnIH6gbbH1L+Mm9tJL5hhTMxw6SAryIL5+QWEDFajniWq84J+VV
5Pxi+aDFI1o1S/lycPz+6UgpKomdGQnX/+rxPBMiAMICwkdjNIhd6CPvFWE2Q2QsmiCNaOm56sIL
hzATOlwRmlhrU2fZL+HdFXjQTz7MdwA1K66I9Rby4a5AcE+kyKRL6Yg7UervQpolowXQbRxZU9MM
g6fWTrnrXF75FuWiqdk7f6CUluiX0V+IOlQ2vSYlDmr3H2bjG2n+n7/48hlJ5RPjikEXL+qlV2hu
QmX6pzC5A1+9X6ocDCgY0VP/Whz5P0uM7/Ao0Yh6PqNUB/9GPrUgvENE94lNbCRpSK9cJl7x3+Ym
1IKO36ErFy91/dmICZgfbRU1+iyQDrn9j/MVw+X+choWzGi3fbDarYRcxcKf93ibH4EZPBhkzYoo
3txCENXnGhZTsJrauzTroKW5za0zBqL7bLbHOsbMNUKWw5jnW4GN83gKHbGV0OGElUBB5xKwAgEz
SEmjXOzEBwhnDxzNh74Z+cfd1QdZcKZnIOkwRSlLBTSWNeNaD1cYMppFMrtgPSuDKvg63sQNMbNQ
yXKZpJ5js/HWu0q7OScJLHq4dul0NilYzbeXjFQQJwsF/Wwi/gThyKvIe2iVJHzt0v6T+wQR+I40
yY3kTFGzAMgxK2c1xW1KgDHynoT9ZAEa4OxMsXDvzucHN3aPm276cdW66gpImQj94CyJn9Ae9V3H
Jgr8swLYBoI/KPeufGQhTA5nsfEXEwP8SFGyrrgOVRu0fkaSg9g79ytagL8yP1akSz8zOaKkbfxF
fo9JhUoBNBTNkdej9qg0LVWtblsFqmRuXSV4WmuXSSjwHtc1E0BXyVfWXAEHFVewSuIEkCxfTMf3
BK/iAgmX9tC/GZKR6wGYPsAlwr2hIwaDeMA5AQT3v+x5uu0dfZ8yhNWUennSRN4EWyUVl+dlpAHJ
qkgm49QHvVp34CGuQpgAfoMWMs7ikaIwOwLoDzUpzjj9MAwtu5yWdW682ZX6ciPOVwUMoVRFlg/h
0wQf1MdX+HHC9bDPk+XXV0V7p15d7s/dPxcf/XOoOyncfSoxqfhnLhwZRQLnUx7IXMGarJIqE0tw
WAqfERKAXP45W+FNpzneW7KZaJwkcr1T3q9PijLYQBWWEPH1JyP1FoH52BTHMJptB2eUAPYcI5YD
MCD01uRz2hK0VAm889Gb5HQllHZ/lsmrwBnDD0TIxI5XG1rrQk+3iiU58JJ43pgpzpEKKLHqzHLg
yLFf9d/KxrCPiMhYZIKYC7MJQO06Rn5YR9imRmSCGHZQGaxCB1JCd1EtMkgWuFF6XwkGmX/mopM8
snn5bOdrwK7r0N0Bg48YI7/i/AUQFrblgzokIP4eI0CrBXI7GDVJcCEXxexILP+9nIF6vTnRqvBo
c7ak4BG2ELoksk3oOWHOhCytZr8kzETihBPehDFf2pldQnVbJ7FR9VcdKk8hs94Np+//lcqrLVeb
64bBk10oPBruI2/TQscaOK82mIJnmh/x7NVqIxksPJVgVjGiAJg//3rfzGI3Uhkv3iyM+Lo8paiF
RLwU0IiTbGr/Kd52Z/hktmfs7qH13pskI4Zjv9vBIL+R/ArAkGtawoTkuy/C4Eue+FWrrLwE4cVd
THOl+asYRDOaY5gQEPa1+/00aKJuufOLFhCe+gQmE1hNchb4w7XD65WEJef+tliZdOpei8EXkzoy
JyEIXsje0mKO1n4GToEL/V393QI0bvCSbvBfheVbSSnlx0gkpH25SaXC52P7kgo44OO1Len9q0OI
M4RKDB1yjwv+OKO89YQ5vjhLxeCBDyRW37qZ68pBN/qAAnxPuWf5ehN1JeFf6v0KqUUDgQW5rfq1
yBWeEUndMbB+OGGlLYpm4MxLbo+0nvoGyfItmvZyHKmWW+8C06zffiSudiNIuFZfBGDWMJcuHs3o
qUdKki4hg9i9k3hgrD8mfX8gcXqOnLH/J4K8kBCzqEvWAdSJH9kZ1UFfEy69aRhFyNXNa5Zqsa6+
PMFLAj/RydIVdSMxsQ1bkpEbXYA/xmKMJrr6Hpol0FFK0m9hTQtEFyRpwaQfIN3M0VKpxmciYPRa
6oTfLKxD2m2vSYonN43oJuwuodPABJfvieuwYc8BEegPKz32YsaezvhNcx8UOPhy2LkrV1Kt22qI
EZSdyvTRRq6ruwiuo84N4Tzp2CoWZqayWYlLY3yv/jmHrcKt23AiW/tLnBoKiIfYjCJXqRxFJhz9
pnj2t7ce0M0wd5nNNUhT+dWlVAIuOs7ssscIIehmZ2Wx48X5CnD2KzKYi+KgdtsX4OVptx6aNiHW
VXqjdTtwvEoV3+UsTGCBdcnda7aWrLqZzA0Sl3dqq0VzfrpwXN74o25LqaUHILruqnKHmuLoaUXW
JnhKiQqIYS4F1wkf9ZrLI6r8R6/AihkVVDDJm8puYEDLqd7RB8fqXnBAZvG/aSiy0D4nyTwRmPkQ
EjQ6qyaEaEvn4L2+w+fnSUX7OVdkaLsOQQSn+UDainBPpilxX/NHWp7TebxYf/Y6UL5WihfQUHki
ocRgPrIYRsV3kHnr2ZUdYu5P1M2O6Hucq5L6zY73Tf2LU9KIzURos6hdXEiXrErG60VE5P4o/Vvn
Sagm6q2Nb/THiqi8Wy6YpnOIcospO6IeAsE6qCIhvZ5+C9UpRAWTT918qHmM1v2uEKKloLhuEj0m
KlArexLgtZ8iZEspKSvviNnG/k9k6iecKiBvZygattc6e/nMx8BcJQxaHj4hpLIbFr0eYdo9+Ksw
MbVlEX7CJK0X5j6ZYHVyoTZHGZHpZ95j4Xasl6MuQN1lbc6CGyBy+bjvhcMfFLSnlaN0CX6uEflT
jIzNhJFYfiq5yx3keuTYcVPu7FGUofjeKW/i56CbERfZ9ztFTgjud4MIIyRt8iiFXj7n50yt70T1
XlVs0DvJIv/8AA6pbTVuEABADX74ftftb/kXbdApgoSJHeG/AwXEfcHj1aywW4KqfMmZhxlsEgjc
05N5WuBV6MSfI482s3yYkbnNms38CHpWsDRUIpCQb6PGcWRrXXhHxJI62uTvLnnGt80g3qqwHgBC
tPjCXUDIKoEmhEsLNEmd7aPBIHKhLYHhJjek3uRDJFCF2K9XFQrPuJ8T9NcVXF0R/jiY5RjormPq
rY7FpjwqP0NxsgHoEm7mXXlTg4mCdRtWwb8KV0XQIBS7dYGNlC+1KOZgymuBp4JKlEvRxN2FLA9P
SM/Z3KwKb9s2EjxlY9dSgKro14xH6zccu+eGyTwqhQVA7O/jOxMGRqvHHMRJSkjoh4AKpG8MsAfo
F85B0PX7ou8AyRrQhUTQkJtPfTmjuW6JTGiYoDI/g8g+BLjHqqm29PxQw+uIo+HAD74DQ5G4wdck
cbh2y6iwF8S4my7vQcAQJtilK/RcRuCROZ6NvfK/4cB02r3KsOcBDv2gTzkyfmPejcvsiurYpYb/
zb9aBouH6tpKVddl4IiUD79NlxH+uJBotjrIByU4fm7eFIGxJhPBgoU7esN5+rxIZduQio8TxWJZ
BEhTGWD/Kk4l6iDtT/JWvde1i4DyH6XHY5F3/kjsqn5akcffU8lqpdeFUljuHhr5cIXUVTQz/j69
EzHYTUn75IqojkBy6yyvq6mepWO1C+RdMtxLryCR837il1kXlrbC4lsZ2GZuIyOeIHLhRdekLkCV
KgGEigrdHoi2d8fuXdw+LuwmNT9jLOeZYW86HgFJhLMQMmEmR8CBWthjT9LMVCDrpKVJbEvoxQNk
nvfuItRXrRhoboMnA/dMb9EJjPgouooLPHmU0XIVt0velHQ35dVP0OBS3z+O9oLQ+X6XECX5diWK
t2dYx+TIdsKsPaS2kBAVX6G1nwOSU2MjA/TdU1iFMe61xg53ivmc54iqAdomdbi9yKD0ToMTQvxv
VkkKmV+HnkW0DfBf871nel0c382+nT8YJqp9lykMIayuffTK6Z5EDGQbLyNx/WjlOF5Zy4fh7lsV
INd5tuRmHcrL+q7B4ZqFXlf0+WiKft6ghWtpeMJMZd6p6hZdThrao8XguAIc3TAZgA/+R8XWElyi
/qDcDpI4S1TC5i4/O/rMldak+Ki5znDZVrEeyu9RnrODZie8sICKJ4pVGPgWCM7jtDeegy6YvCCu
DohFfYZvT4hA/N9U1RKfXOBfKS/Kyv1JdcNu6HTX+RHFNNadqiQHLpIEUc0H/DXFmG+J3XoD8nk/
rxCUIOarCT2rxzRqhjuwdiB1blSgiIVaLpJEUVzYhrp1LvKIpQGpqyysvoXjONbYIL4PXYaje4M9
iVLCgdTgrdnDSlZ00rLGVJsS/fISOo1CgFJ9pLaaE0kBF9QgKLc6Wd43hJeEERikOUM/5RSc5fHq
UeZyWbUqvasSNHHEpcKeAwdEqRlxzr6jWRASjispmJ/wQa/isXKKMNtVT/nwi7klKFc4fjl2HeVH
6ozXY7bDK+q0HMS5AERdbt0ww2oWF4/nCfc0Vf3pDJ85okSWpwnzOkvtvvaeFqg9/KkSP9Kwqpa4
wRCjcEacrNbj0A0TpE1f+2oxkeiMLMLWGovTlzw0MABEd37hkSbZj8NXxa34IonQ0DSA31lxZ/g0
Y05KdlwuAgIT5Zjsti18QK0BR7suUfmekZwFamlk+35rzoLkGQhdMakWJyENmJ2ak1SYCcO1O1CX
5o5+YuUb/oqWmC7MeiPhNKZFKajSpC7FnP8cJXrvuPBPQ4uMTVY0cyCxL1RG6tslUXlUdPEEFdzq
+FQeFFfQm33ql996m9eo7AwvZfI/ZeJ95Eh7ugVtG/+LOMMulXOCblz0QiCU4gzqvIGcCO3941+X
y7kHGIJLoRtk/l8txM+zB5I89Iy83v4SfOOaaH+Rfy40Xf/gED0ESlJj4QttGcJXeqzsow8GOXQE
6ek++wz2js762X9ShUTL7NCDP7kwkDZAwuOpI5imeNx1rVEmWjiANOJ8SZ/sFWLjGX+05ddi+4TD
HqokZEfqfVPeDPSL7Ifmexj6Cj0bUGnFul4/EDd8RwiotVMQ/GxX0/bHK4ZMfDqW7AXd2Mv0sJAY
7Wg1cph+YFo2VyvtTniZl0pZEN+x7o4Poy1DvFX/C2dAyjTGVrywlUKonhPmJPdEl3ljakGdeTDb
e2CYITgQ848YfcPOh6QGZ43LJ3yJKU+H6+ELlRrtPcH5Whjpp60Ayh2b5AqzTTZYtSvxvk7GAXYR
gWw5YlW8XSZSHTRy7Z8kAT8tiMLuTB9Zo03O2MopYOGWV0oAHrTrxnCixlbYCBXd1D5BxQ6RZoOh
8Ot0Eup/Yghv9kSJB+4id1pKQpMo1/wvM3J5JDrHuBAN6/ka2wDbS8va5UWO6MxvS+h/P/x3RN6o
6k6aGowLj62Ay5E65KAfkvfgJFHgwwrqMuu4qi5TUHd9zKVbeXDRjamyN2OjN9iP4HwDzGb7Qd9t
A1yY60WmHDciI3Gs9mGmqp5Vqi82gabFo11OUmNcMmgEE5vuOVyvKSJWqOuwjsOymzRfyMrFpomO
PSqIbPYDKh621gwaHzG0xOPB5YN29gt/pVHrCPZYROUu3xLyZctBzw9ptbxUtndkHwUOKbyqm2up
fKti49wmMUcRNNZeQlaIxmvVpZElDYyacsgz9ULscqS/fa5aJSDb5GLyXTPbRupvHZUv5aedKU1M
+qe3deBhSlWd7TQ8Rd3+D7zITvTUqp91w0hKq14JV5uwRxyYsp7BtzdECHGxT+Vmd8eeqyOOwMim
XcgN67Ndkwlqwt+bqLTq269fOHum/46g7lwK659fPscebTCe+gYMhNeIz9idpCkgKiffSNawQNtT
olLMSTPjXlXs4vxRdSOWHkbReVuP/ETHvg27+NFhtDcxzZv5vXXC59gHq7S+QIZ8qSjHjLpAgEpz
0iyGz6SDCzfPi5iYpUkNIH0PaF9HBIVxlH0KcI90LJXRMjVgZrAX+trCoMKg3O55IA+SXePsCtYS
AO6mWfKKoR0ZuJUajK5DAWmN9Cuo0bIGFYl53GR3F22+Y363v5tYjL4KMSqMvUzvmSapv02imim8
668FYnZbAvz6043ZDUrM05H1OL5xOMsLTR9kt9t1mzaNSkHAkDp2B9rY9l3MeJg1wacOdgUG1QsL
YQIEstFHaA/MRitSBfIAfgeqNM9GxD5InCHNqGwJ2bsFzzaWLfs9sZpIx8xaCiYvmkr8Qoq3sNCy
iOIe55uL1AlAaYK0HfJRSk2Rpqp+Cknm0A0FUZ0v86gT5vMwLIos42Yeu0MaVeOmiqkWLj5gJJuq
oAl0fh8j19FV6KkICK0oxAPPE995zQ/7TJMjjFZB7YBk942vO8WfMt1RckINvYHWSERePAInzeLE
/cl8DJrTBMR7CMZrMe5DhbX9yFKDAs6Ic7e2nmy1785+W4dV2i6H87qlDFE/oLGB8C0Pyjc159QJ
ZSyfDDw4WuZ1sMMCarkO0zQJ+v1nK998DORIc5L9MXf28w0882zeuoGI6NrNxKvO3dtXALqLGdqB
XNPzSUA3PMf8Zg2tpYcwc+SIJp7i19QkF7i0OiPQx3hS/vmw5oR5rOAB+o7fsbJYiilbekeH+D2f
sRK6ZQjKNUndl2TmMRTqoG/0iG1XYTp9t1XHBEVQK8kKByYFtXOSr18VPVPkvtw1FkvqL339AibK
A1r5X//aO1qFD9IF8WWe9t3nY2RP8SCN0aEyR+QpWt+Y1mKtPkmRu2inBXcCaGtVIDXXrRoGYDIn
+kLyyBltK34+ZFJkKewKxw7uo2kR1tEO0QU5fPPgfG38duVQB2QVmqIbsAjxcYM3REr94vZo5wiv
6j4veyc9dBYCD+fs033B3yUwHsaVhvhPJSF1+7XThhHt0cxQlkd6O/FHlRfpj/DF/BnE/mHyPIcy
DFhNuEZPH/pjuPJHZIJQ7Q5enCt3U5Fv89HwBoK4VuLqOSfxsJ2e2JOp4J1YZiQ5MnopF/W14Vzy
JTi+65fq38aN0xjEsqIJXETGpVbgN0CIU5+JSQNy87SmVskNe4kbWmzkVlf/2QrNjIDN3W+ROD1u
wnmh37eXcw2my2lLdRC98q3KOTmxRmqTOAl84vbOAKGKixR8Pxukbh79ymc0S6TLhy458Pslw/O9
mDoarXeSpPte9iwfJSpVFolkEcq+NlW/K08ZXD4R2Gb+mGkXbGF85VlGpZs/TgWqdzcI98cICQcY
OXkWDYGqa9A2U74VOgizbpw5BO89RpYx6bfQWDEUuF3AvB3kliLDGxL06lNYPtfoz6Pl58kapSAo
ISNlVMXIoz6LXCoKrnP93DIqh0vkMIJUubkYWRIOXZIUt8BS/OS8FLSm7IRpJGbx82I1ihWLvy4t
/IWjmZXtDVCFdlfEMDW8elKwumIH1X/JKskpG8Q1r2ySlXmb0E8baFbsYpdrG5CfBKFQMXv+fCWm
UuPNL/4tk8ywNEqlH+xNfm8SozjOf6lE7PXQmr343Zft2XW7XIDKIaqXGix+qeQ8/yDSc0N1iH8G
S8wkwWN0OFcvAALbjWah+L3UnMWaC9pds8VPnmKkUWNnJSUgNvOq8DHBlBJCm/J4XEXv+5aiJ9qY
Ds2nhSs/NK8pJkn1rNx7ZPfu4nKI10P5vbKjzwS1aiFNluvrQw87NdLKwsMW0tFsgPhFF7laODag
GsMwC56nFjFwf9AUUzv3tRShHo+0COceTXUCmZ3qMpkcF8+0uButrjxufYXiRbIbjdefyYnUN3B6
IUoAgilSpBgoXbvsHb+j9mXw0ZCjQUxiFF//uH4f3IZmU4JrR6B5ELYCF47VXRrZJ2nBNEP6edT7
YaOy+gDXW8KZPXNQQA+tSzPGrIZySVBxosn6MBIlOhljff/vGIMAs9NipWbXVmeTN11lfHITFKLa
OsPEU+9wkG+H+T/XHUKpYQXg0KGPakIf/ELmp70Gqm94zkKw9G+IW0o4opFX23Aq6mwdsCaidd7E
Z7TJKRV5i3FsvvJtztxyqeZk/148eh9IQiyBj2gPBhhX1srBAYjvrab/4AieVWUvMvpxIOw4ALL3
gYu34kr5OnZfh7hfUeyBaUk0kJ/6f4L7ouQHxs6ALJ15MxyH01e6FnJF/A3JteyqisRMoXH4aZ4v
GXdZ6v+DSmmcLJEynMT22ND0CfvblW5TN1XibMjfoVNg4/LTwTd10Mcy9A3DRC9/B+Kq2lkP/+Ez
9VJrrwphlzXY3K5DPYYZesFljTOfi3rUf4g5dNXMAWDXXOr9ncOokA9MR61f3ZK/hg6zKfOPU7Co
c0Hw0ev3/dEJdu+JEu/2cDQf+UcdRRTJDqGg2ahSafzHu6u2QRVuFXDXMqL9QMkgZbQ8WrZgnWt5
H3Fp2Y512WpFY/nZIBc8Zz9pEHjW24yaWQwtFp6kOIYaBPxMLgQ10J7xLA2SJD57yMsvNxxWQm2P
nkko5VxuIc0bhWx5GuxX6b2r5nSULDh55xDZhb/Njjhx0is/RnIiL0aE61fqg3tdUSpYVCeil8tc
x5gErSb3SG7QmphU3TFMjciRvPyqbARTtuDNLT88rC8Wky5DgwI5DsrqHXaC07xR9ehoTLtdMdzs
wqkqrzen0TZRvlmNIaZIZKbMQ1wUspfBzbF0gf3yUrFgmXhVN5GyQlYe8D9aerG1Fe85Ej/C9vaa
a0oSOMtoUpvBUlXWtgJOUe0wB0t6dBoe61pUwW4GJZyTZDLwJb4+Q6dn6TrqTiCSA0xrbO5dxYbC
ff8BtSyqpGiKDtz1zIMDEwccd+n++/NuefFfPVXEOETe3c2bL+6pBVF+zNohV3XOjZUOHe1Q/sci
d6wezQ8IXcGcbMxD9rodDOKH0mPKMq1oXD7awyYpS3jlMjkdreMqdizs+BGTnruWNqdoik9CIJGA
3Ykxhyv2a3n56HuhlDrUla/eIAypldz0YnilqD4g+vAAvN3NDpYG/SlzRDedTvOTGM8TufK0prJD
2v7A6+3SAwkGByC5n6TRkBjSZhO9gCWN9O9Fd6ywUIjnOLZtZkIkfPytAbhquGuQoeezdgTn/rz3
R6S1Nfb1dPGWl1mX8ZDAQhFFt6ZJkKBdj6O7+fIbqO6UYmK/SbSIP5YaH0UUJvVtLEfgao1dsc+g
a54HykksruAckI0G76b2D6r/qldo6JOqWWanI428UojQSZwFBD0uAtj/IAEkCHSWuRFfgMHCjKQ+
p2aP2NAVncoUXiXOh1c7ZTo6SdzPQ4Kh2+qU0BAtXJxN7mlLpHt/HXiwoUsFGzOSIBdaZDkV2ZDx
fgOmSW+8pZ/iC0uDCCaGUEF3Q36bB8OavUvsrYkRqgNzmiuBjO8aNnbCHgb5xNAu7zJlJ71r/Ks/
9kwmYUiHzibaECNdoBLmRKdeazbbAqgFbDzgAO/ECS2BfVAxDrwEHUI+WISIUTSntPf0DWqqe8TK
AMfyDFvYNxGCXdLkLeK2k9r53Y6vJ6e+8gEl5IMw1wjYM06jyPGAf+j2gE1KunJ37wvseo0J75wx
QW8ZoRhww8J0FfCv2ma20hKIR0d1l42+TELYvTZlcw+HMm6o47tnP5alw5C63u6P/WCQ96N6P1Jr
sx4qb/5GsqB60qmh96hjCrz5yUi0KROyh4xOfdwxvUwMT0xf1bAGAnUbR4X7hVcUNlmyVSSZci6K
H6QnBLcIA6i3TIOm74TXCHGP6nB6iFFExD8eGQroa0nrTpxTEHU4t5VHu1xuTMRNo+Mdd6a3ydcb
ZxzbNVcDXxSfIFgoX0VtPhL9q0GQeY4uQykC0J6S7iTtoC12UU+Du2mtjOOCFEuS2hLSIEg1Zcfc
1rjwfJyg7Cpu7dtJGx3DnaJ2gNe9P/4VJ9rTPIyh/N6qXq11c6EUzKGpKs0UKEVJByzez+8eUpUU
kB8AZ9tVjpPJUbBXSf4LJK2W362rYsqPRE86N4foFQlySHZDEh6xiccnV259wtZXXyYEGD2H89hK
/0UoUt4nr0kuAIJqpNVkeL38LCUIWBusG6TBfszzATBeU6s2syBS1Q39vpDJ1+boDrduwIW0CBK0
YYE5jVupSQd1IHF3WWznov/+Pv0OU2CpBNh3KDQ7YtAPlQMShuntFbw48R8hlENICJle0QUb4O3s
AGHiL0TmRdIzCyWN0KS7zngxb9mal3Vp8K3yZPfQ6FzPUDg6ir6S4W5EmY1JmVHwKX3S41XOb2Eq
g8OpXXik0IJXRblJ5hEN02wCZTahot8cu1k9v/uM4gZK1hMX0dzjw8Fl5jDlGB5RcIDBgA3eIk4W
frCpr6lTsRjQ1+PXSEl8OtGVZjTHcB5unwcLpcgUCRmFVMP7L/3Jo6uxY4UaxzyTfBH/0uiQrtNm
AZBOtxCZRkSv4L5A8MEyn3RhAxb2bGcplXjOOqRaAAdPep8XgKE2MwLqxlF7Z8mM2T8EvqI2lAS6
jWxHhB4Te+CpXzcv7QpioEeD5AxbPRYnGOdCNONS/gZwD9Xz4+Xjh1HBu880TRDENZgXqo+meGJb
CqoAs48G0TiW7dGsGkmUFhLG6+Zs3Y9/IivYTLL9jyIh4ewjUGCZsecEZm8ZfqhRGAemQkGtPy9N
/o5DUFew2MVD/FU84CBBHCzpCcoagzmtEu4a0rGJxLVaknrF/dvPEqAjmHT4zJbh0aKSarHCCsH9
GRnuzVZz2Ilcdt46IS5RJrqv8RlYcyV23PtWRenEyF3l87xcVgXKxIxYBe6DA7DuY/7lvmyZ1KZf
G4eb7n/WXw5ucsniU4iJVTqn82bVkpPIy1AngkbpHMr8wYaS0egI7JrQOMut0Z7lxwM8sOqdE+BK
C4oQ/CmTrJK/TYXAwA8iJgLyw4LiQFhv+K6TU+d1HxrhjS4O2F4McxLPyDabMd0WvrLp3TR3arcf
RumLtsL7kmHv0aeejplxIf0VduaNDPAkwevbAzjPax69//9rGyetOPtTJCs5vhxBU+fdvMyAcXFr
GhAwyyqHYwx2AklVx8PqzR1oZSJvd7gfVL9AyOEvLxCHnZwaw0OgIFjUMDP84iEBoutzFTkhNmK6
bq9XKmQdBm3hIu4EBWJ6ICUrnAEqjVd8XOAp8JtZV8WSD1XWl/hSgNqVV+y76It79o3hUuyQoWNe
hsApts+510vY+KC78e18GbOSTNJLZy7pvLQSf94lD7Dt8GKcipp2JXLvOVdJCgepn9+dWYwnGCy2
lEdjEQNQpw2fnSr1zQTNQ76uuZ+WeMvBSdXcRD5y3njJFqbFZF9Edl1YFzYe3dbZAAC7lxo0VOc5
ZbvhQYtyltaOQ0pZt4B6hizRci6B5C3uQMkPhqqzL2TtwNvoae6NlPWFDVsK8/HYcbQVvY8cD6Da
HRRpvB1TFMcOtW56LCSCZB6pOGn6Txfx1IFE4eBDZQSQWILDxTZBszYQwnNHsDR5XUmorRubYdBw
8ssGpalmX5VpwjZ09tFOU4qsVemN91BwmptI+OFm8PPun59h00iH/bZUXBA7AgafSWZqZ6Hde92X
wnFtD32OcfPHqAix8q51y+300qfQHOWOStt3wa3KSCYYIzqjhScCeVOzMie1iU7qApxks/xHoWPi
dsD6ySv6JXtubGWM/MkLJ4Y5X0CsBuSH6/ddSW7hbXAweRcSNcoJLICp0ko1y4PCqc9tlsUzzfJm
keF6GZfByE+t08yoCX4f5kc+78dt5XL/44jVnHnICsKqu5NilWny3uPnHOwQ2ebytoIWLCE+Uz25
y2KStvnmGlRxIzaY6PfvOBzGan6fnidGGOREDVZMlDoUgWtrVFWLDTPHgjDyi7qW/p1HYTRWdprE
YTBasSahAK8a52HLBKprbl8PL+uBL9fPpQqkssHHsmyl7l0s8Tk4ulXxR3QDZ5xht6U1DmnmF/aP
fbl5+Poef+2v9wvqOSZOACOuqy6rhlzMreX6SgZW2g//aICf9o1RwTADBOY52Dip++sS1yldqKNA
ID6ltWq8LrpGuhorSyzCMLDuy6+iTP5oj2Bq5jZoIsCkLlC5yYjJN33vX7QuR8yWavTvUJBHI4pf
j4636pv1lMmjuHqHOWSMmgetJxgqLS0FVQCVf5SfOTDqpo/zS2qlUF/rAj3cNhBjqtk8InthMsGN
wAUWqN2nOd5UsZv8WXC+kxuFMNmokO3yHVOLPn6s1Q/IZ+QiHUR+7yR3Pu+6br1A3UVB5gqmrXId
CruTEPl0cL6sFn8kbVbgGiPghuLVZQ6M
`protect end_protected
