-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
BG2G1YLJsl/ZnKYQsFgygtw8Pr4vMvMUi1+hS418nYDDIYfYZyZlFZgJj6MM7YJj4raAvyfKvoP5
Y2QTA1x/mZiNe5ECeDOAjVd99/MC68eYo8SuCJ+j2xCBmVylZHgA7joQMzs7qCm4qmBjDEDT4xhf
76ST3IZCk2GGKUyJ8x2C82NxTLu9TWeQn0P+G55vfQEnS9hbC1/WXuamAjsqcL6e0DDXKoDLB9V8
pAHa3FY0t0UyjJXjWt76Pc8FdCDieso6hKLP3bwzdAmwb6LFjN7qHWalOdL+tjQlUSSIQI9/MiOe
dIejUeSx9Q+orZJE/2mV1ma+Ge3SepKHhKNOFQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 8848)
`protect data_block
A+1XWHGCnLuIJFNnSidyYM/pjpgdmth+hOJINeCowwP/Czcg1zlqJcb7x/Jnvp8y0bAU8UlWadBc
BzPOEOREiLpz9jCQBsHM4DVMVgq1EpGyN6OY43DxttcCAlIhjbCaBBHERw/oh1f4Fo+MibUoCBrV
9bOMGhOL/iaa+ti6sa593YSCi3nH8hnBF9a+sc46KZaO4X0KPJhVg2Oo2iGEjsRbb+pzi2GrznF7
fUwovSZFVYYhGWR55VEwRhf1UGNTa4G0SC0QFSuZtF2o/GkiJD4TiXFyBx8K6218/CoKAa+MUiFk
9yNe8BTGJ/qdJmxtbhOY2XmZ5UT0Hpdh1UQ7SW/zJsEVIjCViKYN5y/gsQmpg62GEspZwGPE1+Zw
mOSM2oDWwdFenA/UF732DfNhWC2qF3JdyFPe5+zls5KZjmUkYpCgAi5u9Hj79zYF1HbiXCKsyx8t
cJWyg/VDeQupPeqG4gitewgRui7pQsUlQLmB5m85BGowGZ3RXVi9m+37hV20O8iL3GHsTRdLNzLP
lH7VWBzygB0ZxdgQ6lC4FVLc6y8zs0Y2BAP3jjcLOPWuK+9TYd4L77JOFbb4TvnKbyAwkt39M2uv
pg+Mdg4aWEaO6P/ssQTNbDTnvg5eHCh7aDZzKoiBdwiM8yOctx1tmhIdnsWaBLctyWPlpCnIbElv
h6WNErgBloFhYTwCSvIgIJZNpo8KyHO5RU1LyiYutN2wBUnduhLA8QUqd10kBWSEVdmhMzN5LL8m
jXHzF8jRcN2ii/6+Kc26x9/OEFn5Nt5euhUiJVM91Eat6wppqseLu2E4zvVafZx6sO13UcR8pSUV
yJdm/zI8qdAm21XK2Dzmv7uF3zKb6Iq0kWQdFqoK1reCjZi3ztwMFmbwRnHnGA2LZKTw1bUaFEts
39XuRDwnYAxJE2oIDldjfGyqZlwAOOHaA17rmrSwgG9K1j1t0oQp1ud7cgH8b7Cv7zu4JQBR2Lh+
CdFOV2IrUBnQcvaNOHTXYYR2lIDc6V8+qktNftg9HKiIn7/a0JGAt3mKfROzosyso+uwQaLiA/qT
pGesXRDAbUy4+EOlCy+MsDf+TG4sGV1V9aRRAN193yBB12ZHoywwxGQe+UpSuNeodr2yaSFd0KOI
rQwGis96RCJDFN5Ez96OLOQZafdQRX3G4e08QqfscU4sCPOmfFDmSn7DaiVWxzcvlq61vrIkB3ms
itIF6dbjj1CL8fQutQifzLkCUgMmSvTrdxi5IohA2ZNMM6DUI4O2/KJxnZpqdW/W9EE88b12rpwh
QDU9XAOtdkadfXrqQIjLZCkb3BMf16nCvxdUBq7v19iYkOYJB03ht2XuHpWbfr5DmcPhdn1LM9LW
hRjoST/GzGHLAtLpR2OX4TmiebpMQTb2g7BnSRd/cBU89kpOuqj33fVtGXlZtgSA2Ws4N1VQ3amA
lg3/K11iHn2tY1052BdbHVh5xTTzmUtqhA33PtdqIVXQljOZM6wDli6s7PYv9qGzt/uqlAEgfV/Z
/PhrgfschoNYwDZiRlI5dawSQ+9HbvgfbnBffTsBkIrH46R9I9XatJl2pxUtVtr1m3v6Np48MGck
hFaZlSET4qj0wAA44N0m7JR6WsiMvMwULU96eGonDt8PV6JU7DkRge1Cftnrt1j/5KRkY49KqlSy
iG7QLA++Eirckxd2jPE3ErGz4b/et8LoxiiH5ot3/r7pE0JdIMwIKVJtKjoaf9GaGdxVU7fqTOra
Duti/S4jvKqP1EzrQdaKgFFU6kMffLhl3XY3L20R3fI0ak/dSduyk72daUTkC6VoVETo4a8UbhB6
t59Ci47z/8AndBux5lGgI92oE7NpiWa56M/3+rbvBEg2H+r7VeKXMvyferPhBSp2deqvuU4RlU+t
10nwiwHSpTXRblYcaXBPEMEtbCuZLcOyxOueLpVJhKTcm5DQTyT94sQ3jgZcfUl5znnZxPfAuGTb
9hvne/HdglAHKVW+ZPo3CTM0NUW2BWUkFk5pbsHGgbHHOPLQNjns5cA4nU0Nj5UVePSPhzS8SMJZ
tVr+Lnnmp0ia990MT2q5Th1s1475hW4ftYl2M6cYiYB41md5eYLI3HV8yLdGrG862sxCmHwDtniA
UPKAxBlguwUKYMtkWMYUC7x8s8GfTr+YNmGUb3cZfZPQ+J6ds3fQPHEk0N5U0yqx5YuusH19Nm77
7vsfntroQzdFG5vqL+oWcRcpWiIZObtKeWgEWZ8E7niktGo92Amv8CFsiUXI2RdwoGdwnpVHkiVk
fm9iQm1hdQxD4pdd9drj2shNvfRg369/Zja3dJjkU5J79+rHJ+4D8z8YlBz4B5MkdIiFwjazp3Mx
qWscgxakP5Iqe/6aQ0AgnsTYcc5f8MvjuBYlAj5Pv6loeSod7T/jI573Tt4Lpr0b8+XIJqjnIO7Y
XdoEWAK44PWTpPz8qFXZO9DNgWFt0a6QF3+sFkCfu7zWvbpMtaRn7ibmcRvYI5YUmMxy3n4QbZq0
tk3MQd5XYj0H/OpPD2ZZNgfjpgb/9I2gtW2IOh1NOaYu8bajB/GBSQOt8vEJb34vrrK5PEElaN2z
Pd8w/tcdA0ftVb/+bdaxzpT0yGvVdY+KFeCpqn3TbYi40oU+IrT+Qrbt94gRR4+7QKogxtzL1fyE
3QPZQkUc2ktCLrJ4BCE65XGrPxdOmgeZ+BNTz+V6lFatb6PmNb7A204uO/1Z2FaUcir4+zvTF47F
viKlysP2ZHDf+nKhFpBxpnh/N13iTwpoR4O9hKAEjRfGcY37mGDHM0AZXqoUzvX18b7pFGvv59uO
umSE+3yMnLkltozCUqPwftbgUPwN/zdm7lLd+EymY7NoNUEWy4bouzOitVnzdhOauaL10JP+sDoy
J1L5zQ3a8rmG1ic9fDpLNaznV/kxo+GLLgXFA+iC1EVJGxYyUqQIcZ2hK/Ydpmxy4Swny0GL5cYN
Muto67wxCbLM8Z4QOu1D1YxroiWhiwhA2oCfm+Hsm212zWCvVFtVF91GZ2G1QEn+hF6BzJbNiuVs
pKuwPN3OIjQZ2wFE6mCTrTH1e39idICcEfo/BTbzThZfciI5a3mJg1tgfQpb2LH/rcdEF7Jiul6d
FNC4Zkjn3U5DxpXd47G5s0wQvDdXKNlhLIaO+XzMT96t4jjE8EqlYzwNtz/oQwV9TGaqGNgr2aU5
/r/w54onk523T0pQsPmYXUESBiruuW696cqP7svhL1yfTI9FBOyKks1TpLMc6wnzNVrJ3M1jZU/z
a72PnPKwQdmkjp3wen8nwiwLfPUlI2S3WRej5JAAo3r2cVLmhfB21H6OFOVj2CQ5yP5tE/JDgygg
L/A65oyUsIW3k6tTXPL1ZG9zsGjK0EhIv0OIXrV1P6Cg6xGYcirc92Rp+/3b6z2/gfAXab7ToYe8
fKBL3rTQokXsFUKYIdJuEMiTK32WSM7ADPGgtxuiyylLk4znOIKd5QtKMV5GSuRGjtPzaKOwjwU9
A72HvcyLacNP0oIrlfaveSHxv7/xwFQQHBnWx1oC6cvDOTaB3ulgzA4vn7G+YRewH9b15wCgPff8
XrJJS1W8jJuzoGZvCeJ3+3UCye9xDnYxcUxOIgvaCreHstQMYx0LRyf2oOsSOfmmZkX3K5MAIuCs
G1oUGnyB5E+VZ7wCCIK4NvETWng+OENjqGurC1gMROYr0+Tr7Vl8iS2M7JnpVPd1JMMThE5XcJ13
7w1XCTPZuqIR+t7vWqVzIprE7HEhVq3aIFFssCewpfvSFSo7XRDU9gTUcb820MIhzsyAED+8yRcO
WI0+rWo07i4uJ/hqn3gVRyuuPpuza428VK0QdO1fkQAICDKBxUSC8fjoGsrbqEuTpJvfonFlWBgy
uG1hr5zMX5OLX7EZbbvKXN2bC5V1jy323q9WcHbervxWXt33Q+IIeUNCcUWpjcfrMgva1FRyQaUO
9e0Sh16AL87Q+WAA/6HqhxaRdR7vABmdbAUHpIRf0MLJ3NcglgGnJk6hZWsyGhrwQT/O8mwkFedB
INVgX0eo9ktuocUhD7NTxKeFBXqZA5X8vdOcFzrcXzRXbAyfKOQQ9nSgY5JIpRnzX4eEPQtkrKKo
KZnGDv7dwmLT9nxErt6F94b0F10MA7vvUIJLwGxxp643rMwc+CFeDT4EyTONj8L7SQvVlsiBzdp6
MRUv0GxQPQBlgj/lLpOPkO+rkL/vQP8dDnDrNfBxk5WYj1zpUQxlY8W7BgAX8ow9IMWa0Hp8092s
30iAcAtBCwuFIdp4ygPwvJvC1Vk/jJLNMmnsPIao1Q2Q4ckwtl0BGDe36o0/XvoSxcwapAgxA9+k
HkrDOfRN2h+Fgj7CE+ivd6uN5sadtoPZ+YKAaBZJGnMo6z6b3MlAn5uWsv/L85BPYXqTc9lZHKdg
nQtgVWLNimzly0gsK3WMNiYtE6GczNR27JQMAZUtCak+HmtyDNLP8E76AiGjk8fZXMwE/ivTSUBW
YA2fEnM+O9aFn9t7WLETCl+kqJf3BQFcYBoDT43CUYBmJPqrHVMWqpxhRWYnI9T+bohE2oZCQ5NN
dAsEjax0GmJ6zqO9S6j0BLtQnGEnzIAJ1rQyFQva6FEdxjpMOohI3ABIPtMEoduNtJ2/8rFX9jl8
i2Cf7E++37A4MM51bteJ0/53EnvkvK97ZefWEXgu5jyK17rJXxoBQqY4t0pp6lAeT3pEBBhGWOZF
KsxS8gVXwhEFRsNKsK9ysJxp6WAjBmDor/59OG/r6c2gq5fMMRScNm2jqFt9NAwLucfjd1bLip4E
JxQMMiedyTQBoI4E/VvTJUU2ZkoFgej36ht1IWGQf2eLnETsZBdp2zNHDzh+HRnzSgBUS6GvIwgv
32/N7rBshFVC0B87B/hzQd0L2fx2GLFxshpwx853m7sUq26iOMwhFlilQQQpoBX9fVNU8uDhjvzD
eNohyebQWbUJyurNnziMLyxL1fcR6nUgSLxkKqDBQFWwBQC+CGZ86P7OZdM5wCgH1wMCSzAJFjrn
6pjggRwbSZab/bYzdIxCo0DOvpt6rWuFaCbjbJPFoyZ9FhUMLJ07yIInfvrBBLnhAEpN+zo+RW+1
bpQHGNqynHmM/DJfiq4ovWeuwixFbNUrTLZv9l39sngKxMP1Kga6goe3UVrXHQ8SRijNlC08gzJZ
iKckb+9hAR91UzbzlWAK//MMuV57BikjGRJdASXJf9skOUeFsPNRyv4OiPlodf7W8HLeNiXn2vbA
Irn22hBmC4P/J0vcfMYFGQK83s8edYV1yBkBDHwRuOu5b3xC6YBcq2MKrk5tintqgP+et6p9mf1K
zw8yxZWyQjvWSMClnayDxCHs5Q+opcn5Hb1/sqAxNCp7rKLP0nTPhOF+uF/RlipTUikIGBWINJ9J
QtTHM6kxltUMJ0IUdkTMLmlW9E4YMkDDdpUmvh+uuuKB0ujjXWoOEgWqOBQvto5rC4d0o2gDwQYk
WqyjFzGupu7qCy+gOIgtBprI0+1zlOg0+QGssRTCEu2mNxHPTbN0wdoUJMVMke/G/OmJvYeJ4ORW
JzLDH0/CnpI6R1eLczXCwaz+s3CS3kcC0r8S6GEvWBQ0srTksfazScbjCZUkzKUXUSiHE0J+dLMn
1PtSvK+rWStPGtbhUiMvL42Mdwyq6Srs5juF8irfPplLYosiutbLkOL4SKp053a3RaphvhquGPsa
BXiuz2RRHzs6zS7Y1DbkN1bI2FubMiV0oiJ4Ry8cdfwbugscO0/DjzYzRMqm6yoLixpjpml79wiW
TmNhjLJrAQ8/ljAs7znMiD6T3WAnBeD39FgomBhFfitWolxUoym4YxyoHV5TsVGQWWY4+oZvNWsH
1zJQi6Vw06pBtKxIi4iJ9hZQKpgEItCmp0TQen9w6izqxZ216LEJao9n7mQ99LoQ9C62xStrhexh
w7+EWZ/DmWTTdqrEsZ4EC3+k95NVtCcjN89otWup+6I+YEuCwUGQRYlNJQuNUR1HhUWGyOZdIfUS
WNZT/NQiEoca8AbU4XI1qJ44GJ2cwNneCsOPYtRuvU8os3DCEfSXvcwqTR1flU6PevP9qYdsAFyp
4xE/EH8GHoXEgAFBKXD0/43XnGFzeY1ZqZbAz12yb9974yAAgnNR2dEBl9DJUChsnRVdLNH9f1zi
6hYeGGYn4198AjRMLXUN2G+VjmNqVvG/ze52ovXhNHybwiQy3fuVN2Du6jn4v2077HY7a0Dwcb74
z+qW1Q+m4g6sginDGBJy2jPRERnvC1lKnwdgEyGOl2MxC+JalX2fjuquIxGA3BCke7V17tQctJdE
fm3VbT9pmUOLNLHHKhVTc+mVQyHhZx1mdJI6xIKNuERvtjMY4ijhnxdl6cPb1SAdoxqBVNVWtyEW
j5UjAQtfq78+wN8RJCC4ba10eOb/Ox4EbN7pwQvuc0J5XIWb9/Z92rQtMAZ2Y50vd5dF3BkFmAom
nEjbtacHpD8LCOHShHSoOElpJwb5py7o1h8tMYMOnIWMO8aU0Z4iL+6Pz+KN+Ee3MsEmgrc2AOBs
fv7c/hpf2fFNB5lLUu+yxXW7I3gEE94+1QB1BNYOQmbsoyY2UC1oPDS3wr/ybKYyHYgptGImtr8C
BFFBJ8pgD9KZfHWTtMy23h7sycDIGugJEtAICmVHy2Vqksluyjc9tfRtCtQXbfXis+vFU4fzT/vn
FMzcja93feHqaOxEikUXaACiZrX68yTksuR5X78L1XJntiTMWfLBd3ZocwPpNp+TV7qFQOupVVP/
KlpInNmLJQusN/bJ3PyzAojoXlHLUGCAbDU/YLRF5fQtcC2oVtXungoY+iKg1gP4U0hPyhBg3cgd
EyEAMX+n5V+CSHrB+yHv9ozqsnl8eDYd/qiTQHz2fk7FgbL+96fKCk1zUvT7rVmFeX8Lv4m4LXdK
ENMTSMFiscDJeXAxu/aMJiJWGELCdYd9wgIdNqcwoKBZHzRoaAcbTGlbn2atjYn9C6WaAUOCcq7o
tlzhBLY/8YChE9RZf8oiGlukcj6PeF+rxeL6hRQVcLig88VKe+biUtZoLs5SnHJjmPtm4ZYP9xG9
exhIPTBHBSh8eGNqPuDFLpkTX39dtKlOaV6ToSdhiM4yMoUk+e4n3ZihM2I/QDpzq6MsjNTttDCX
h+HO2pkndauyQzQq/e8cXdBu5AYbLH4j6liHKkcjr9W8fnVcEEQw2sGhmP40JZDKpUwRkMrVq0lq
VRWTmvKaM4Eay5UchZDGjK1GBMt+minEcPxTQRLbcmp14iodbOP8NZOOHEgAlYjYlSi1wMhuh/t0
sAaeR6QtP0tx8NOs83T3PHBc8qz0TEBhwS40baIdo2j/fE+hTqUIPCXZHxFHmAZG7DwQqmu+/L2P
opDEVud1bfqhJGRdWXIMm6qwgIP7XqSKIO/UmgLdxBugXusfGLyKlI4HNXDPlprEMW79bjDmEgEz
a02HX8srSLd1pfFuIdyLnRcuP6TIk2LojXkazTLR70m5h3rVFcQiG72ZgafuqR8c9njfkxhPMV0W
BayjQLzj0ZnalDCZw2DrDGNiHYI/28vyKn53lQ9zeflF4gT2YlkgSGT72VruYPH45Stpd3ngax0U
xP1tiDUXRWZDAimUTi8AFHA7lGXsQhZp1kQPBFNKnAQgvJNZgBeK0KHbAv8SaeF4YtXOZivkl3+F
J5PDV89wfUPM+ezGMwNn7FmWdnI59jxlBZg1GGwY9P78G0I/s1HDDue90Xj+9SfltF5wMVlk5Nsi
P8pvgUscCZwzILlUuaOLvmLrngUh4WtaKWC6cB75EvUFB+roRHDGah6SClLYZx7bMypb1ipKETWp
vJANLmMUzD0glMVt7vNJZEs4z1HDUBhtGCTURIoJG1cGBpraKW5CqQ6a1W36FsX9suufc2GSwS/c
Tgvf0eKeft00iRIlm9EcMz3E/26tvvBQBOpfb1Ldb58NMLtnfrWbBDYmd4DheegmZPwN3fwU5x2J
eebOQysI+JiQQMv+v3eJr3i+yKKjxsuTM0/SRiwoorJ5XRVRkXuvq2Zy4uEZr6XspDA5lMtEqArK
8Kmn1haCUWte8jn9Zx4OkL/HrkBeYhtmiLzvLIv/vFKKzK+U4eouqyPwj5IHgUqxXhaH4Z3+4hMy
XDhWcKsdO0TaMs4df0pEDgMvF+pWWZsbYglDp/zy+jwBBVUiK1hv50s1hJxEgVRNdIyOoxutV3pA
bSbM/oP4VmvLq3aHr/IzMB33vWPFI1GrqpocDMF2u6syHXmPfsdlczLf5ZG7HrHiUi3PhWKKt0Ar
ObWNsPhQjGpLoc5OvWB6yFjBoJ2GLEGeILy+XFd7rdxAUsUc3PVpHQ67WeUFqu1xqeeBXr7mKTY/
+RbFAbJYNKEX/MGgaaZZUF9eibommrlfKHXh3AXF3RVmsJ1oqV17cyieElZ/cFUh3KhEkP4/O7F9
h0DWjLFs6TJdgihuzsKqD+DY7dLW9S/qR4H1RUflsBiw0feJYbcuH9hIZ38pEa4k0WD/pqi7F0Kr
+mGbdQYZsTdCLtSsMhNzzQ6MHEQasysWw7ezBgTYjYKnx3VJYP8hiKbcnQsgWZO0rf5UhH8OAvZz
5xXxknG4cEm39S1JR4nJ35AzlXb+TtAS3j2cvjjnxwH17GsLgYMFasIWPwD37yDMgEwKVQv/SVrz
HP12hj27R5J1vLvWErSILvNOeBWsQ8PAPWTSyZopAxUTK3sN9uhZGiFuL28U50oN9r0D3L7AyLbv
KHoZqvWAbq6TvLVO3QSEBMNvAuXV1Noa3g3IlW96lozRquN1/JfRp2k1LZua4tGfR6cMk+iKhRUy
ksALTaOXuuzEhv1WGEPT0JF9lGZUsp8xXUzmbQmQKoDEtiDzTjxpZU39uBIO3NN8aS1pu9gPBh6k
xQuFbGqLbOcgqxthpw/40n6cu0xvrUaVZXU5hPwST7hao5oX2zltxsd9u5eOXSRrgDislHhLUPoc
yhiMd3jJT46tiwv2d1koQojwrqWh0VswykZ27YeTDSXXtCaTPO+yE35lA/mtr4/2ytsIGA4MIUB1
ReAgJK8KnoeXRqtmiKGIKq9V3nP04I5m2jeuchXA/Z4PDk1cTcki914PcFElcZIq19ZTwy/1ducW
dqMCIGBrdp+s1MME8GtRUNLY7hkpIFWIuspwgiGrblz04qOxd+XIzhb8SaoGmf9/g4vHdghWa8+6
Qjq8vQc0UBGKvlfdoWGNTXKZq2oPDpENReCFo3sXe7WtjO8OvI+dZLgKIqrew/ckaZoh0CWj1FZe
euosXAf6I+71N0MR7Zozn7H+obeEwWLBVGTCf2m/WasuhWOpGGd6UmkTxKccon3fXfygEjYHlP8Q
BCWmSP4YxK6AxPlc/pGxNJhHeQbQ+R75BrgNY7oqcq9TlHTRuA/3QrHc8F2e31RBnuGnn2FciLit
90U93mBmPJWY1qwPT7DLQENdowqKNSVkFXyqjO/NuY8mylVbx1CI3hnAr1j0Pe04wy4e6rOrAGJA
iVa+PTWe4sjECv64AVqSqXcm8JTOAH58FqaTh9MjGBzMuhIqih5lVcccBt1FhYtZW4yLA2xeEC9e
UP4o35cI1lLKnPUFB++3ndUXj3n+OWXn9BtgaoJqPd4CThrwr1bOQCWnbm1BKd4PSAkEUVP+uEk0
U2Gnn7RODW3K+WiQb0NBw3ZgIvy7rnOy4BFmlrmOt7EW+N8KIZrRfr1QUzCpe3a6SdRJfhiCC8cN
/lyWtlA8FYtT+vDLAH1DWowBtmTHpVrKfhcDihsK/9SMSKoP1IBKPm2Ah+3NDafgaMKTsD+VBVGN
rtgDxmSN7imm16c3vhjnuMtzgoh4+dMD+Nl05Nomk4hakryh5W3WYbXlNBmYNScaEZKX5VXtyT/N
T0aNThmWL6NwG8rSh3xE5oyS9LULKbmcGvpJbNprXOFflKrGqv4pMXh5CQ/3UJ8OoRmURf0CYS6Q
/hfqgW0Tanqdh5IqtvxRm1UlVPPTA+aJG0+gyXaM5m/fD9UIEZAYf3Ay5JaaCfZCScuGqZ+XJFbo
azD9Zataq9Qw+FOOC6lIQD8sJXIcH/npPU0DXC1UNn/7QP/63nlSUPg55TDMy0aeE18EVTFgxLGh
1CJ4yPJrUANwv4Fu/R97rQzD8oS3okwmy6LPiHo0tVm+IUrAuJ+tLrDZrwCMzErlFQldiJ1xYFSF
c7movhOhzQDb51BfMISzlmtLPgUdFEOmzVqpXjkXzqeLzqcjZKNGHC44FsD4AhuUzgrf7rFy76t/
o3JY4Ms5jWDiIFQSKgx5HoBsW5VPpID7DdwKK4g2CHhUzXojqyANaJ2yGFxnie4Po6pqBFkp/WMN
Y5XxPR6bf10dulFL+MXQzWI7OxXGtty0fQO7PW5kaqrgnvKyHowUvjYAUfQXhkHjQ9ZwbTlGnfqd
gGos6sXTR4FiCdqerhUTmyLjJPEiRcYWSnr/71x7KIlJSSg3xqPqdKiasruyYoRVExVKyzOnqfQk
QYcMTjlMeesJiIwrrTK137wL0ZlcwL5fJt7FjMzogK/ibFxYGkNci4QlNNIV98fjFo1cypmZAaUm
pDEuQ2Q8A48/sqbBGZhCzuKhN5p4J6qEuJmEH0RVu7ncCr9LWlbxYJKuCuvDmxj6tBOO6VqrV1iu
3Yhmikmj8+4El9AN5ZkykEeiMZ5tTHDa9hFdpwKLdc5b+e17kx4hB2fVR6bflkkU/jzLePHQpL/2
/CASl8v/5z6bg5781ZXurxvcDtq26SDaC0RTsAjQVIILSKgXzHJISf9OqGS9IXMI6U/qBSRn1gQc
A2zKE9NTF1+GjWSX9pGhH5gzouLRhlhgh0NArWrft8seYLINbUMeqrYhCSO7u8qKuo9CxQlZM36N
ooV7mQaIhtQO8kCRSNJM+Hl8p/Dp6gsd9EgrWWbqLxd8jttaR6HzQo4zFsjf2xD8UuneLs91nWfY
tydvLibCUXiQGPommXoABv0iKzEBDpkMeb8H7HQV9tE9d7NyBalwqBWkQkV0Vk2FGiPB8wCh79jR
6d6KjRta+QLsSlc7ID0sLWrHEpozaQUijpyuIr3cBGIQ+G9LRGg/lqsHj99iXJ66ppluNoA5lpW5
Vemd+X0QuR5JTWjKi5qY4hzqagA0Cevz5UXRW9yjMRf06zKnSl15xrgHmyFGOkYw3TAiyhLmp1mR
v4PCqFRF2zSsTcEUr0uYAvcQx0OKuzrdDzs61dt1EEVeeS1aFEySxW72R6hJSgMyyxqvp7O4ifdz
1dHeAHVNIdcnwLUP+6GFN/u25IN61t07D1aalJruHwuS06xrBl9j1dseP8fKluZznEgm0s/QjNwV
+gH5Q1pUhBhksNY78kj3eK2iTBTsVe+oTlgukSfyzr2vBPJzwrf4yIcu+v+G8LaxDHYlTln2cnqG
pyydd98hEGrWXKNo8hUGm+WqzqAIy/y5dVvnv2QncVvOI2ZXPt6tHndFNqafPEbezEOaneJVQzCA
H/wSv9OzM3AjTRZ9ihCsTVXt81Y+Je1273SG+vfOy7Q7bafY1KzBy66BEX9BCcYXhPhM697aPVDa
KNr5TJM2iZOocgGvh1D6kUj6p/XOhk/EYrVNiV0NtAW7ZNP2hO4RV6m6xDZN204rvMYKwQq0N8Oa
xRXESirgrreHazIFm1YkhQSF9JTDv8PAw1dUsjL0I5+1yJeZ0exvfw07YAuiKmnuJT/fFfNHsti/
pcbB7UHjwlZdHWIkQ5hGytS0Jm1SCV+6OYEvc82rbjSwx44pAHebp9IR1CGe5M/KOECHDIITyK4z
oJAxXIE8D3TzPSAHVg==
`protect end_protected
