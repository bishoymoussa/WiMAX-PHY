��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$Rx�y�<��wA�*;�x���@�̦�W�X�fa�M-$u����n~�%���P�$��W��kYَ���P7�?UMfT��q�6�U��k�>����~�\N�(�����X�e���/6U|)�X2pF�]$h���d.���9Ecb�%���ow�Z�}�;D^k~'	�c�'�ɺ����&���%P�h�&Fb�]�e����榋�y*�%�q�����Ѐ���!�B��$]/���kc;�V����պ�3_�v����;��e��嶰��'xuZ'�+��3@w$��
����O��o�45U�4l���ׇ0Z#�o�D��<���N*��}����p<�#黳#�I��ן��)��0�Sѣ��a�!���ߨE:��RIU�c��˰�֨����`l`g9c5��D ��?�xm��,at��{s- f^�e�7��<%�Y@�x���m��z`L;G�{vR�,
 �����~��'�J9�zҲo� ��.r��B���H��o����k�<�i`���@�a���4 ��_�X�j�]��8���DO<{�c�t�Eq�2<��38���M%S��8Nd�Ҫw�������)��VH�sI�1�K��6�f��"���ʝ��Y�����V�=�/Ļ�M(���]h���H=�.XɓQ/�)c�"��R�M~��9)��8*�7lm�^��3���$�҂�.Z+�$�r�n�w"q�=��e���7n3��Y}2��� {k</q�n��sQ�6�!��³x�
��6J���(�c�75��g�����@���B�nU.xb��X�Jɴ��w.�q.���i*c�@�p.�&��@(�3Y�P��O,�c�s Y)=ҡh�N�n��;Hq�W�U7��k����f�R��4fc�_��^o����SG[g��kk����]� ?!3 �����MTW����j�&�j��N˺d�A`��7	�V����#�fQ��-��ԑ����f�y��"��P�j���&��%��/Ӻ^��ڲ>q>U1G�=��G�|"~��ܧ��1'߱9�<�	�O�C��mBku��:a5�O'��<>�p	nLM&KҖ�nO%�����*�c{V��6�_�'8��73�?Tx�k��H8��L<+8�f��	j����3F��Ǿ���ͧ(, ��S�A�5�I�斘9�ճΘ�Hn0olK�ÆKȿ)>G������Er��-����]��S�8c̠��!�:����J���8f�|�� 𭄎�q��p���B�-��J��[h��x����ߐ"��P��tم T}{���D���mmg6�k��M>QJ]��o�J�!�9�
�]M�ڧer��1�0�jv�A�Q�2Q��u5.0���`Y��AK�A�d(��٢�����Oc������ҷw�r�j���r	�_���!�gz|��!'��jܐFKi�޳I"D�+)��_���>��WI�7��Oy
���0g͔��-�Ws��Cad缡\F^��ԲNiN}V�G��a d0���hm�#מ��@Un��	}
B��դL�W�`����	�+YX?�2�����yoJ�K�
��U`�8<�hՖyZ�p[�T��P B������w$�6m{8�B6��K��k̂|2���f� )/:/~�5q��|D��9�>��[čQ0����h�3e}�K_)������.���C�D��?3�jq��s�V�le_X����;�<��L������ii�x���:�,�ݕ���3G��v.�p����^s{}߫[l�r�,T�T2�g���B2P�dVձ�2&����+9Wx��O���8Uߺ��-�8�j����<=̃^�R�#'�xr���$U��@��$��zm�I.�ڤS�#4���p���h�u2x�Q�wy%�o�2�R�!S����H.�����޻J�D����WB�j�J���T� �R k���;O���ui����9��؏����x�_�\�։�>�&*��O�m�]��C��y��7=�I�Z8і���dZ���E	���D1���њ����L�ν�9펜�F}��j~E���-l<f�s�2�8��0����9�#q��V��X��]T�'�֊��o�O7�(��8�u��$/vԀV��	�G��5�[����6��+n8�]m��z� �T��U&J�����sk�[��-a͊�	��f2;�B��lOMZ��(a�+�ÖzR����á[)�Q+�9�	s������\��q*?�/6�D�O]�$����	I2/�4.���L�}
pQ��eb���&V��i��?�����F�M\�kk�(k�Th�$�dmBj>�.�a��?4_�,Ly���w��x̂��C�m.��nOk5d��b�5����(�����;��XP7�V�?YС3��;Ux��7Kz�ܚcU*L>�π_6@dfm.X_�
�*1$�6Rm �R��<��="�(Du��I�i�K�o�g�p�ϒR��l��&G9*��"�:�"�z")/�"a�����TG���x�6>���g[�(.[O�����V�qe���)�r�(���s��JI��ue��浦kca��F�������:�r���>%�ؠ�5A|-���/O/g	D�rJ� A���Y/p4ޖ�F�Gٽ�e؍