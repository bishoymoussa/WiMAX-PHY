��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$Rx�y�<�f��p��}Ԇ��c�Ͷ�Vϛ�6L��q��9fNDjG��E���L���5�\Kk����(7�������y����f7E�Z9^LZ�'��X�E�h���mD�Jر�7'J� �u��u��B��A�^�Ԙ��V1V�-�G��Ɲ�z�������<���Q���/ ����������,�������'��H��ޱ��vՐ
����[�Xs�O�.ݬ�%\�AVf|s:l������e|E���	 ��{��(⹈��:}A�y����zb*�����U����{
?� ~7�����z� h"�\*�B��bo*�����}M�ݯv��doglv�AZav�*���IY'��¾������k�"���*C��M]v������<���hc�Ӟ�ҕjeV�tr�[����ވT얫Y�����R�_�*y�`�H�l./�0V�3����sD�E�G�I��}UB�g`_D�h*$Ǚ<�&�\Z�5�� y���yGd�NC�!T�$Ө�iV�q�9��M��%�3P��0���V�`to"ɳ+��;=��^�3@���*:Cw����>�q���ar��z�y-�#ah+#	�h������D>F��3�&�$F��kp�
?���?�j跷}7
�*�kŐQ�㱳s�	��Gqs���g�eW5Y�*��1̟�wͥ��g���Y��R1@��][@����������Q�G �|Qf��]vy�J���+#�:��b7Y&J���f9lz�Փ�JtK$���?�RC��<�B��L�^p���������DO|�-�ٛ�fۿ�;v �遗�9K9���p�8��-?$�w
�C��k��K� �Di������I��H�ˢ�V<�0���y�g�UgP��m�|7�-�R ��1!i�R���:1ޱ�SC
{�k]n�Z|�����A���m]4��W���6[x(���Rʘ�K����s�q&F���d�6�	D�7ڔ��$n�*5��t�yON
���1��Ӈ)�w���,~��|���Q���v�����N[�H���G��.�
�k䒶7�o�/_O��S���T�ss�p���p�[o�=�=����h��!�7p�e�fq�3�:Kcƨu9Ϟ@�$�?�& ��=O��O3�`4]�d�7�=�x64/Cu�n����W$�ԯK��z�r ׫ �`�#rD�34lU�xiɁ�7Ղ�2`�.P�: ��@�7��@�1���hQ2�_S�#�⇉Hpֱ��Y�x�p�wF^Ն��9�~U�]�8�]�^ʑB��l'0�]�wsBl�3Y��#�,��lX�$S������f!��X��j��W��5��ט�:�Oz�z�d����� ��Rv,"�� ~�-�t�&�I����䔪�*�]n�~��5�&$��L�O���F-�jIj��k��	�!]�lvSd3�D������C��9S��=x�fX�;m:�aV�I�pi��o�w�Wͱ,,`i��]s�b =�<�6�����`�x� ��nb�z�Z��J���4�*����`P�z$�� M�nD�/�Ӣ�v���U|�+�:��Is���`��
�v
+��@H��n�Bۧ9W�Y���T[�$���Zbm�#x�k�`g��/?�x�M�*P3�Ү�����m��ߎ��p�{]顁��V���顪�[e�=^js��PP鈬|������t������,����#6�S���:pu.0�2���q>�s���qߙ1�ү�{�o�,�p�G��$�lwv���'X�[5���F�%��,��g�H�qʹ"Q?GN�
��aCP������Kt�`h$�0��J,l���0��;ol�!f0��yH{�8�A_kj����i�M.j�4ȅ�Α�R�[�Er��D�����D;Z��8u����7z��-�i&Z��ک784�8���[�~�^��|�:0y�=��)�x �*@v�H��*��F�H
����ZӋ�U���i	����vZ{�S�"������D+��|$����2sE섇�e�a��;R�J��2"�UP!�+l�ƺ�K^� ���Kh\hW8����9a)eg&�l?��UN��tK������p6��A�ڿ����h��)�����w���cN�_��u�C�Sԝ* ��7��X��m��H��jq��DZ
����c���+��?���X`Z�"���R؏�����E�"?H��&��5�IW���m%�������ۈ�o�(�� h]i4�Ӭ�3 k�j�D�T�2���N)��/נ�����	#������\xq�5���?x�,�b'��譩���<���L��,��Pi��fR��s��!� ��`'Ed@��0ٛF��s��t��U�6F�S�<�7�-�@1ET���l�F>�~n4w�{�?��\e:,/_�����H<	����2>@�k���ncC.��F��l��kzu���^�kg)���1��mQ�hM�r��e��j���;�?��	n���6�$V��e/hڠklU���m�2��\��\Я��k~l�Q䁛�1;!D�U�~EՏ�T�1x��ݭ��!����H�5�o,7�S�tF�RJL�Y$̆3UC},Շқ�Kl�װd�M@�Z���`��e S�ן�6� N��᭔�ޙ%�/Ȧ��6__�b˅0���8�@�稔��+���_��#L��jy;@���g�j2�/�Ŕ[�7iB�Q։0��Z4���-������1]�<*�})K)��i��DӥSѻ3Fy�9���.B��B���7<HC����$ן
���[�+໇p��pۀ�k�^�6�%<g��3,L!ѡ�k (+HS0m���l���hgԝ��zJ�@=�Q\3��|J�a(r�Q����A�Ü�J��E>U�嶼�̾d!�\����M� ��E)��-u���Ԅ��t8\�^�:�W����Z�j��~��5�\]�!��mx���B�<�>R�kn���,jӖ���蟲T�^�-N^�:���V�[��/�vՙ���Hj	X
eV�f����8 �T���D�0&��_\*0>�~\|�G6�zag���3�DItk.s������<ǿ��y����?�v~ϖ���a���T깘�Lnho��sN.��@'�/��C����� �/�cq�{�c����i�l��1)a�������ٱ.Xa���'�6��H��|��5c�O��������J�#x;͈\�	Uܹ�y����B��_��܈��bX�A�E�U�D�^�:�%������j,���Tl.�-��M�����C�x���0��ï��.��ŋ!׽�[��9���S�W��i�a�5�����l�+9���'�-�RɀtY�P!����gM�[����ߗB����{5Z���-|�_j3�,�ɁG^κ��4�P8D�w�E��TM�x���
+�~lg'DM/��cl���y�W*0�2Ŗh]���D�j��h}D�0�2���6�wd���X�}]ty{�+���F��v����/�ZB.k�"��޳,�y� M'y�'B��%��g����`���=���A������gC�t�B�)��O�]n�%��hI'N��i�.����$e���8��M�+8j;�F'Q)���@H(��
�@��ݗ5ז��,�E{3H��g捶�[����[/!�� �@���b�F�>ctʓq�%ͪ�M{:3oK������~�w�e4�)����
�g�C���Uᗛ�]�k�iw��c�!(@	�������+��.
c_�zz�Xl���dy�Q��2v���e;��xU��llT�3�ă�]�L�j�{��}(��\��䟞��5��U0@jƟBH�YZ%԰��P۞�&u�So� �.ȮI<-
�������P���
~غ���r=ɢzz�玭a/^���� ����G�C���.B��ʌ�*���h�9�΍��+��i�9׌>����,��6�~��srI��Ԝ&q����k�|h�X*+MV�,��Yup��dDBk`N��~��d�2�TJ�r���a�B�p�,]���j�Y6>�~�	)��I�|�Z���������i�����x���<��)����N��AA�X�5�oO?N�o2��Xk���֗