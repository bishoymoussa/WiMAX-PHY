library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity FFT128_tb is
end entity FFT128_tb;

architecture rtl_tb of FFT128_tb is

component FFT128 is
port(Clk : in std_logic;
     Rst : in std_logic);
end component;

signal Clk: std_logic:='1';
signal Rst: std_logic:='1';

constant PERIOD: time := 20 ns;

begin

--clock
 Clk <= not Clk after PERIOD/2;
 
  FFT_ins: FFT128 port map(Clk,Rst);
  
 -- stimulus process
 process begin
 	-- initial values for the inputs
	Rst  <= '0';
    -- deassert reset
	wait for (1*PERIOD);
    Rst    <= '1';
    -- Read data 
	wait for (130*PERIOD);
    wait;
end process;

end architecture rtl_tb;