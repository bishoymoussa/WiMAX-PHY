��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$Rx�y�<��wA�*;�x���@�̦�W�X�fa�M-$u����n~�%���P�$��W��kYَ���P7�?UMfT��q�6�U��k�>����~�\N�(�����X�e���/6U|)�X2pF�]$h���d.���9E��WG��L�X"]�Ad����ľS���8od����e�GT?y	7�������ݵ�^��R�q^]�鍦�����s�ae���h��L��P_���ާ��YЭF���'\��68�b�[����w8�[X��V�F�0͘3����q諵�uW� �h�u\V�?@��_6G�_�*�G���B�絉�f������[�G��U&�����~�F��AׯK1�`c��[<��FY���4I� �#�G��x[X�=�Q1��`��R>(�w����R�O�?����7�,(�H\�#h(W�EH=�������yq��Ѿ��aF����:�U~m<|��.��0=�P/���4ǆ���T(�����Ql�2+N�J��8;<C�g���HRp��`�cW��pk���%�6��f*u�^���l�^υ3�q���tW@��1e��ޙ�B�
�C
P�;�0����"�!����w�%��ڣ��)�MMC�,���羒̇��rG>�H���H��|��q���E�S��">�jg2/�Le6u����Q�U��N�;p�@y�C�$����l�}�_r�~YLX��.8�h���2�罵���,$l�ƚ."$��d����o�66�cu�ׂЬ���'���P�5T�o��d�wsbl��n,^����c`�Լ��P��oD��� E"AÏί��fZ�r����L�6L�y�S��:Y�b�l���C�Jq���֫� s�r��|(�;���Q#�N<����vZuӼܦ��O>G0�Lؠ���)�T5�P�b�k6�?Ct�J������d2J�T2Śy��re �1��T'���B��/(ڂ� �%�U�<�S�h��.�݅G��?,��+��Y籈8��MP+ѩGJ�,�}<�������Bt~��/�
��o[ȁ.��׉[u���B\$�Ǵ�<�q�Q���!нE�����B����I"���8ٙ�D7�n�;Tױ#x9�D��W�z@���a��4H��5Cg��t�n�H�"�U�S���NڡH�j_K��O���=ކr�8�#��֋�	s�pO8�UìN~:"lt8�ġ�� �){W�^K����p����{���_©�a�ic{r�H}R=�`����P`-�f�S��;�R���x�i��Y�{����z-UK ��L:~Cm�T�d����[DT.ڰlkwL�����.Ә�y*4��N�Ȱ++#��D���M�|��b-ڶ�m��`�4�W��Ň�_ʜ�M�m>h�]�Ҟ/</�����҇�ġ�	���[k��.�y��*���\�OhQu':%�Yn�JW_5޿��W����A|uW�����x�ߛ�,�l�(���Jh��aJ��?J����Ǘ�xrØ+���XF:�}����@'��7��n���b�k�3�X"���wT���P8�O�l��H�΄�Z-��3�=w���� t��iR������(�9�q�\7Oe5��2�@UB��A�L�*�^{�}����[�P�gw&��*O�e�{�<X�X��+z�"p	��x_ru�8s����7�����z������M��`�+<��S�e��ƹ��]�؆�u�7`͍��z�*��c�\��k�%t�ǫB��y3�D#�U�a؜NyhZ�,zI�}�'���ܶ&B�?��8����`�	��^!�y�~Qp*Tפ��h"K��0�on�+@�d�d��SOG��ۃ�2��Z�.��0��Ɏg"q�h�����V������<Ю�H��(�ʼ�һ�'�.8�~�iC���i�<�Ց)ѽ��lf�  �QY��J�S�6���/�`h=-�V��B,ԯ�פ��Ox�m>,͓x��tF���JW_X�7m�5���`�U�:�XyT5���-����X�*^��ԲE���	��0� R��ܗ�n����t�	2�B�1�zD��A�*�ȱ(&u�P�H^�~PyC8������6������ṕ̂��	��Lv�L
���q���T��|��9����ܞ;qx�ߘ����
̩��iY"����/�hAD*q�v`��Z���6��^l�����o���e�p�oN:�Y.�'��0d�1���M�+�y;mvvdE�b~�$�Nw�K������C��9�{Ϗ�U�i�;�r;�s>0�#�f*�ߍ�j��ֆ �Օ]��VdP!\�*�'c�e��ʙʨ
�h�Uk�k�[�mĤ���3�-t	�d�����
->�*� B��a�L���QC;خ�U5`��"T͉����^�a|�a	�C�:%ݖ��
3$����׿X��]O{�JW��()c\iW�DW� ��^41�w뉑\xN�/�'~:s�z#U��lo,{�{q1	h��4�)�H6���T#�г�	���Q\o��Z��<�Ο���ispp�,��y��̨C�x?�frby&��໕���Nw���/�M ��	��YB�vO1΀���6Ԟ���~��m�ai���o�J5q��k�b�J ����Ә&��?�E��4H�O�1i�!�B��T��R�� �l�c�����If;���2v;4b�BP���r)��Z��ͣ����+��
�l�W(D�.��$y��൚g��~I9{��?����v<���I�m1I�Е�I�;U�^t�㺓2�ږ�<U#Z�t�Di��»_���NM�=��0'Ρף��\��������0s7C�Z$� ��1�>!1D�7�p��s���3J#<����d��RX��[�%���������C�W���%C2C���z'��R�m}7��Ģ��!�l�1��U��E�p�I�yW��(}��qT���M�t�%^"��o_���a����:e�f�W����_�rN��\3��>w�ʘ�cJ�o3�#`�G��}���c��2F��L�gmE�N�a�w����:���"�Лw�u��/����=�5D/A+��̊$\?��|���W��JFJ�֣�_J�*u�I�:�^8�s�G�|bC�x1�����]��k�4�h��+t�T�h��#�-iT�$�}���D9Hy�}������j̨��9���q�l���Y�5���K��_��\�n�뇎�2�`Hߵ��Lͷ3f�Qy#�`OϷ+�YD��uh(wMf�P��y{��#}".l	�x�:)�h%�_��s�E����A��4�cĢ�8ڹ��ߨ����ػ���i�bD:����3C�Vo�I���e�[����OҾ�҂xB3�i��~���(EasNr�X��,��5�e�9P?h�*U�:�㦾6�(&/Ւ:�wb)�%�y�{Q�q�fFk`�}��~���
�e�Z�;(>��b�5XܿYX�2/稜�1�!m�SʇF�Yy�*���[�zs�B�A����]Q	v��t;�
Y����B|(��
;3�cm��RպSa��~�Y�0���[ú[h�-�	�J�C�����":f��S�u�2w�6��Z����<˂S����D���k��1;��bxj?` �pZ7��_�NU������K�D��!��Z!�uM��SJx�'Z|}��730��G^ݜ�2`�+8�����l�;� 2���L1o\��d����e���X�����,��6,R֤}�?�ÐɎMY�.�� �O@��A 
ư�:Ĩ��f�7�U]��nk�M��>k���>U.�"�t?�/���m?���m^��-�5)�A�!].��8�'
��&p�(_��W�1/�6�E�pD�D�5z���/=��D�ʵ��aO_�O�~f!�rA��M&�7�EdCR��~wO��nC�^���+��7b4u��Ǜ^M�l���<B��W|̿��N<h�󞾓j.�܂�\|���J�\����i�.��Ѧ,���J�x
�c�\�|�?����j��������-(��,T6�}G�}��5�\r���"�������[����c�t�4�K̻���*!Pk����^@f�����.��}�+������Z�h#N�x�G��ռ��=������)"�T�V���HB>���תD� �Y `e�8�8�dq
��SO�:�ׇX"*ɧ֎YZ�	�n8���i&D�%zME��vQ���O���>[7G�E��	�B����5�3��-�wۀ遏y�$4ע|`�.q�Rs��ݳ�;�a�A0Y4n�X�g;�Miw��o����)�[{̜l�tt���@����K��|�q��0�$���M���[J~`u,c�G2�;������DW�Ǥ�C���!p�����@��f��L+��~wus��� r@S4��A90Fjp�W�tzA�� ��6l��$���́!���%�M!�x�`���B*��j�،S��S�^����62�'��?�L�z������G.��w_tn���;b�%ۂ����S��f-s�2�E2Fm�����S�ٲl5��*���);V�R*�Y��2��0�����n?�t ��A֬�eEa�̫
X�r/��g&�O����5���!�PtW�y���oK��s㎖��egބ�(��r���r&��^�> ��I�p�ܱ�N�7��8Ę��(�y�8�}L��\̈���%lx�/��]��m�] ɥ�d[|Lz!��EDo��T��F0v 2[��{P)��,�Jɛm��?��(� �X?3=%����ғ���4~KD��5i��J<fá~�������l��r��~b��YC�=�}�P�HS8s>p�2��9�$O_E��kY���~��D��'#Q
�y��RK���=ci ���6��B�ڬm;Ub�g��j�6��ٓ��hk۰����Cu}��Zq��Oܾٶ�F!��ӟ9~��Ŏ��3��eBТi�K9ލ��)]�:r-��mB>YO��S�`KzG�}���
؜D�6!>B8`�Ǉq��2��îh����K\�٥8Q;�tF�p�D�H��f�0s��%$��O.b[��0��O�����uw��ޡ�pv�zNWk@a�}l%��	M�{\��I8Z%��v���N.�-��3X���>OX�ꞐT�Jy媖����=�Z��_?
��ދ�f��d#'5W��1R�Ia�IXh�^�(P��ĚdX�3z�լ�*'��k���z;�y)%�1fm���wQk�Ct�X�}lM����� � ��f�U��SA�L/#�=�-�Y�#ՇݖV��dbE�f;�>��n������*KS�l�����w+��\����8��`� �Xd˯}%�O�R*%
�*�y4�I�?�� ���}\�� {�irQ����֯b�\��+�$�d�$�
� �rv���~GR��_nWʲ��}h�Z�'u�L}]s�' A�2�!r<k�p+��o jC]��-�I)8,X`��A��fq�h�i�rk�f�-~5��ر�&K�߉kf�f8Q���ͷ_�1'ǹ���
��-š��:����ϻ�PcO?����㣒7�cze�-'ܲHjk m? �sqT��=�2�_q?���ǐ���c
����]��'�NQ-K�c������0W[^�~"N����A$�i��� �]e"�XgQik��(F*欸.�,+.)�2��\qE}�Fj�xa'�;�r�-�S���LV>D�t�&�9�o@L�&�8�B�q���X���C15��J��b%���FA��A�o4#�� ` ~�f&�o�Q���T�[�trP����$:V��|ߧ�� �˷J���Ɋz0V�>^��E��2q�r�<���fć�[���z�-���=6�8
�r�,t}�(݂��7��O|	���{dM��1��g��Vi���%��IH���,)U�L�"���9B���H<iR�tĻ�\A*	���X2=+�����*j1z��@�M�0/*��Ƥ��ΠD�0�����0�qz6�!��q6���ّ(��쾩h���@��$T�ڑK5���7�m�3���*�\`?��������Ri�E�;��C��ʏ�G좶�Ȉr*MQ���b�S������/tӈ��kI�g�-��J�L�S�U�U
������E�3G�[� O�8B@�_�-#�¼=y��T�Dq"���y�9�1٘�X_��ٓX�W�_�}��.�dNu��?-[���BJ/jC3x�+��=��̥�)����mv�g��?ǀP��9�</3{�XH3�hl�
�oN-���p>�� t>P�Q��sg8L_=ѩ���9 �n.�{�aI���L���X|&��s+�ez�C�1LJ/S$o,fN���p�;��������j�ܣhl�Ǣb�^�p*��dGua��Ǯd�l}/�D�5�q���y��D!�iQtp�ñ֠vN������VmT�0�Bï�t�ށ�򛥨g�ZK����׉B8�?��x����ئ�|c��$.��۪ȩdؑ~[���!K@��n�6����"�폦��ύ`P����5��w�_߫q�Bͭ��Ʈl�$.vw
�F��7�D7����bF>rI4���'-�@��v3���b��/v���j��X��_ʥ��o�%,�22�!)���,W�.G��� s)��O��z���1�0�����I�R\S�P�������p)s~W��!P��$F�͊�a�����UK.sYk���V����>8ED�1^�PL+��b>�&��c�WX4�}0!��fh@۫�gY%r���a�5(�Ð	b��k<u2��C�+��LZ*���*n��+>$o�Y6Q?�xҊw����,@V��*�x�|�����i�H!�k�nxu��#�^�o�@�d���0Sלq���<�Rh�4�����#����V�6�3�Y+�S�(��x�<����ٿD\�\��J\Շ�L�y�2c��m1����D\�-!DI���9w
���3�⯵8���(k[��4%P88fH�.����Z!u��Z��*���ƺvv�	�m-��KyZ��-U�J#����bҁB������Ј����<�Neb��i��Wd������|�F��@��.�O�I$�?0�X=0J��:]I�t5�>R�������߶ژ8�Z(�����Ѭk3�]���`��,+�A'���p˿x��pv/�*&�zֳ �&v������b��QӠԊ���޼�����u�󋴺|�����@Y��򖀯}9�R���v3� �����cHُ��R�֬��������q78\�N,�ki�KSj�̏))��$�^��\vgo�z!��w�>�oA8t��_NCʯ:��/ۻ��z�􎪁�"J��������G!��l� ���@&��Yp���P�?ｰ���ҷ�A[��c��h��3Fc�ٔ����'#�k�-b�ǁm���<�>y(m#f��� !ޫm�`���g�F?�<Y	;��W�$����1�����$5�V�*j�ދ 1_(}K���u-�������.Ů�0@�}�8������w�2�.u^N{x��]���s����Lf�v���/��:�}��� m�^V�L7����^�����l��5�r�\P��Uf��P�������b�3H����5`���r�`������[ًv���G΁�����E��n"E���Am� ���`�	�J�=I&<�'�f�a��&�꼘��Xd�OT!9	���$?4�D%4��Z0P�F��
p��?�V�<��e�q��5����1U*��2#m�>�8~\��x��� _DeQ�yQh�C��Z>�d33(K7�R,���;/��Og�Uq���9����շDp�$)�o'Obǂ"�#�Q�{��g7�e��v]$��-Y:!cG�6+P=#��f[�[�q?Fҍ�<�-�&��� ҺK�H�Î��ŗ���s�0��c��_G�����>tx'Z!�j�����i�yl���+쇻us��=բL*aCgq!kO�0��#��T��v@�
|��Hi�A���#0CM���f`,٤pZ��쏦NJ���F|��&��݄�+l�_�3��;�7��	%�����9M���|��H�O0!:_��
tM�{�˕�v�G��Hz����%S�X��/.y �\�6|�f�[~H9HS�al��x ��v0���Mr�U�Ȩ��b��o��*��ѐ��|K�Z��*i�WJ��h!��셍i�Wy��uLD	���m��iR�t�Ġ���+\�cfQt���BxR��ŮFE_��!�"�)sE>���]k���^�b��3�6X i��d�h��.<�j�+�x��Z���y�	�Y�3��+V�#�D�s�**l�8E�[�#0�ңh' ��M3|a@�n@q|֑���:Ȟ���`.b��wU�WYH�/�W�9��� ���r�Q�� h,��B��SU�t�kY]��J�ˁƚ����cd�G_��d�ࡃt�SWWs��LT7��6�6��� �neO��@��e��u�L6��GS���>�F���B�4�����*�yl#��W+=�a��q��g�ߙ��i#Z�Ͷe��\
�����>�4�a?�2���|��<�$��M�0̞rp���A��78�L*f:�u�wڝ�gt��T�5"�=O��.Kl��8%s�:��L���}hRKP��$_'��b�5B:w:��a{5{b1�>(�S�,TT�σmga� ���V�o^��k�
��Z�����^U6���y��I�M}? qG8;̜[4��+�C��泆�dx7���p������E3�+�5 ]�M�$$�Z^D��a�">�+���L��T���g@3�u��`�o��:E��8��&N�4����d��"O������c�O8Ԛ�wR9���Y�����)��+�o�B��fu���ڙJ{d�5t�8�˞Ț�${/trLx�3àJT>����[�� �d�m �R�U��k���8@��q�����&	�r�K�)c��	<u��A�.�9'!ϿJ�w�8K̥S#�Ӫ&��v�0�������͕|b�����@�<�߆d!�xU*k)ʇ3���7�d����3X� {���,�X,գP辣	��&��5^���Y�n�+�#o�Us��Α���?_��$������I�
��D��+]���h�e&��%)���j�ڽ����vn��Op�� a��~ $l����?P!㼭�9�G$��i0A���?}��?������T��N�Io+\�D�@���S�q���$��!�uۧ�\��U-���c����{���qU���#�[�-=�!������/qW㹓�{PW�(%�IKgf�A��#N�&�_Sn�ظ�kw�$�TvG.m?�ƽ�[����8݀|�]�X~H����6��v��	P$2�_Q��� ��
@v(5�@46҉W��,�bv	�����K���]{)͝TH�����P�{���x�}�r}��RC*�/H/ �)Y68��W������_�	��R� a�����\Po��
{>�)0�Q��I|�D�t*��ց�O��Vv�����Q�Cd�r�E~�c��52����s2[ƟKW�H�pC�*�	�.f>P�{,U�Ǐ��ԡ����@ȯ��MUr�+E���r��>A���hw�I�.U��7����7��ώ�Fx��;�P5��k�ߨq�a�JC̀�\!��b�(�������Í4JLOQFwm-c+qǥ�;���� ����0�n��p��]�ۥ7A$	��P;f���4C�ϗĖ3E�t*� ѓ�v��������;J�!�=��*b)#�)D� J�z�;�O���#L����oҎ�[��S�r��y~e�{l�A��.��v 6�!t	Pq��<�)�zk8m�F=�/��8&�R?�F�/B����������l64(�ܖ�d������,����9���<�0����Z�4�$$�o���I��/���;~��5ևF�	=�WJ�!e˄.~5c�Siﭷ��[�D��}8�+�AV.���z�R��cڎ��5��,�5#�yI�3
]3���W��ϸŅN=m��C�}�^,K�̯���E.^�B�,�!�`D�p#��8��>��� �h��S�LA��YdF�Q3�S��"��6ݧ!��Հe=jV�`ANs�d��Qzm���ᖕ����Ri	�ϕ1_D�ݴ��l ��-Z�l^�X�L�=����_� ������*Q�)��>�&��|�"v�O��yJ!:�lω�Xw,��c�!C�Xw�̔pPz������=k{��1m4�m��Y��͉��(�׵��	hW����✛�d�9���=�ȯ�W@�]��B?Ft%)�{�0�BBF.������<�Z��� ƞ|����F�_�����_�[#^@�?���l�|��5xB6!�X���w?B]�pQ��MN��{���>�{}m�`��;���R�B@4�>�_��m�戺&�Ei'�핊��h�!����w;�G4�ط�T,���;��XLZ)�E��C^�����B���N�h(�lN���� �(o��%���l%���y��i�D���&����O��c�8?]�W���`�Lʤ�\�'�ÑYԂ%n�����)��&���ko:�XE8�k���<�,�j4��,_T�N?�w�bh"M����� ��8q���[�JJ�`�,�61A*6�[J8*�+��L�y+���ӣ�_�v8�!��1�YME��l�l: Q�[��i�-��R��D`��9�����u=�ڶ}�Ǜ�����eoY�h	�v�P�dˋ����@�w�h�ik�oJ�].�q=��U��_J��XB��$�-��Ů����� _ܤ���8�6�.����u��1B���7���/^.г��	��ꦲ����-J� �p�i��l��Zd�(�`ֹI����TwT.���G�^��4e�fY��V���|�2��0ü?E����b�X$��P�g��?��lSF��� �a�8���Uw29���0D�K+8�>0�m�čfm����5R-�!��A!��!-��&Ni�՘/�i�$��m��S��r{��l:E��h�;��s}Kғ˅�@���q�b~Ș�TP�}����r#{��RW�T�c�\��v�b��f*�(M��Өh�������BD0P^���ky6�J���+�� l +��w�x@���9��B�Yi���4���it���dŶ�Mש�Nr�6с�[H���26��+*���e� ���ricz)��e�f�M�J1�\��;�G�+�����A3R���߅a'���,o@������ZxG�pM+��.~R�!𕟷B۹P�1W�D����i8Zn^P�z	h��.�[������;q��4�-��%=�Է��Q[�F�Q�.2��V�u����3�9���e{/�K�=F��
�8<���+���~e�U�����r��I\+t��PMu�O��)��C���З;+����iBEz`�v+�������������`1��L��~��J�����G1����h�U��S9^���o'��dD �<�mk|?�b<�`켧�qۗo�8���˘�F-l��7�z�b�h��Tj9�n���D����5iHk�K�������ʱ��/K�ם���j�%8{a	`��l|6�9M���V�)��DJ.�/�y��H ��mvk��"�,�����5�-���"�⋠����=|˞�����Ө�ɉ�M:�WU�ӍФ���ߘ�̃f�]���^���� 8?��LB�~Bݮ �j%Γi3���7�����Ϯ��������C<z�u���XX޴�_�ض��O��)k��Z<1f(5��ya_��o	n� �rP~6�|Q���<ь��{Rw�wU�ex�=�M'�P��F{������%�����h�\�&�D�D�s:�\@��t���h����W*��<��h��lvA]:�V�}n JL�z�X9E:!r����_�3Ѹs[�M�{jH��lU��\��ꎞ��M圊7�foOWe��������9?�#�3F�:�Y@K����C�bdq�g�� ����Y>"�2���{7�ߦ-'��
vG &l@�nlY�c,��2r�?3����l�(S��(���4����[�:�JUِ����L�����S}<Q�6���h���gȭ#n�G��W�6��Ք][�0���~�%�#l�>���ϩS�e� Е�y�ܳ�~�+R�?����m�^�J�����5��R|<���0Etv0�4�ܢ��y���W���:p����XOQƓ����
H�wPy6f�r(��k��<K񗃥w�|#;�ַ&��NC�1�P����?�Po��tL|uR�x�;z�P�T+j~�+���*��s^�:#]���>WJ9;�����{����cq���­�����s�ݿ.��P��<������H2?���\����ctU���˨/
�M��$�6Ǩ�ӌofT�I� K�=�k�l�t�)�{�2�����X��;�	� �EV�%Ԙ�9���E�q���e5��h"��&0�+;x 8!��L��B�I��Ӛ3��*�w�*�S��P1If���0�Xiϥ�6@�(��c�M�o����UI7���r���J�F�͡�	������k�6�7ޞX5����7�@��z<���0� Kr{a.�������.>�A�7���W��\e��2�ƏyRi����]��a�u�Lԗ�C$x�}��:��8Sҍ��'���r���P���'t[ʹ�r����2�٘e'	ıEH0�
�Y�s�P�����}K�x?�:�Fz�tA\t����c�3�_<�pD�	�p�q�iGƟ
�^!�5�Vh_����v*�+����M;B,W�u���0�e�x�?��F{!��V�P��)�)U3ؙ`O�+ktuM=���5b��*n��
�N[��F����&`!8)��9�~	���HY���\�$0�<'N��
Zef{l���ݤ6��U��v�#����xd���Yjþۊ�ܭ��d���1&Ѡ=�T	�%*z�t�>�M�%P�ޚ/��<ڕ˹���fF�����p��+�P�����t?2W\{R�u��-mv�$��D��v%���sΫm�/���@XП7��M$���+����>*�2�W��̈����|��8���j0� ԫ)#P.մګ���:��� ��ql������Z��46��t�F��D�@�PU|>��-�
~C�S��ۺ̘�z�X��NI�Tu`}���pNi����v(^S��	L��-�@W@@T�N����c���������k*�{z��L{4�������i�E#�"��{R�TSV���CFҖ�z`Z+�ٖ}A��4�a^Ζbd�?��SnrD�@*�Oؗ��?������>Zr;�NZ� ��O��a�^'(t�\S0�}9Z�@����R������P����,bC�:�OF5E��WT�9I!Ty_d��6)�뻞�i	|�	`�_�wn2�S��(N_ Yjnb���u�:A�;����E������eŁ���	��vG�%���Ɗ6�/�nG*���Yᆕ�V�O�'\��E�u R�q�j\z���AM�Yٳ��8��g�Rp:\8��mb�m��]� �T�v�-�QeQ���<
����3��M�@9#B��4�dg�/4L>�1��ݧ����a�,�����{��U���s�*�x�`�(t�i����b��d���dIIG%6H.΋��`s��l{0����<3X�2%��������el_ O��k7n��;^(�|(7��b�8G��|�ѧbVl_��
��<w��JE��y9�8S�&�
9��|�b�/H��	!�aҟ���;L���=%�ihk^ڻLt���{��/>�`�' R���_l	%ʰ��M,h��kM3���Lm��cR#?C#�aS�;����s�i���VF��c0��s���Z|���JlFVwf�G	�~;Z-F��RٶVZ�8���b)\w6������ͫZ֚E�ѽ4�2����Y�\�cz��h�2����6�����;��@KB�M�o���"�H��!�;��1-O�fmk����ޔ�&�"X���L��L�����T���{���SG��gze��F���|�ܶ�ey�S!{y���gchqwg����#W���b���QC����^7U@��ࠟ�U����Lpgյ�c��gE��7	�>1�����Ch#:AOH ���ښ�_�?�Ob����o<Yl�3�~2y��1~L4�B����tI$��z�V$S�[� ��ZtIli)�{v�%@}B����R
��&^�m*���S̱����$49��B|��>�� %R���"��W�Fd�6��@�����)�3��@vaE�r$�1��C�c�v?�������!�;~�غ���*���q�|9:���n�3�CWF�Adb{I{D$��҄�V�[sF�b\,Tt�W�$G����bd��gltc�wM����/e�1�B{���4����y�T	�8�%!S�R��]�
�"zM��f/Rh�����<��"��m+�C����mF���|�k��s���;��'lx�j��Z�����*�����Xu�He��iU��7в��8�)�ZUz�6��T����9j�;�2�\HF������K�����,l (�����nPs�oy�B��@�����G�X����:6A*)�ze�7�6?.]lX=f��dH*3��ԧVM_R�Sc�m��C�C��@�0����k��9)ꛥ3��]T�%)�̮��7}�/4���^�����A�ل�p��dC�{^9�op�q�E��g�8A���w��ײ�����D��ÿ�z����[�V�K��������_��#Qz�W/G	�g���=�2�����,m���3 �v�&��(	yEJ�2�}^�{�]h��������ٲ��zS���o�^#����L0X7B���}/���I��/*XQ�	��1K��(B�`'	�֝�iŏ���J�O=�-�r�4�u#�����]^f��E\��)��i7Zz� <�/&2j�4�vFm��2���O8�f�j���}��D�W>�,w�OQj�
j4��8�)�C��H��
i`&v�/C ��6?�ƅ�j�'r���5E|1Vع0�9Z9C,������B�h�}P��m�����Kr{Q�a�<Zz� U�s�2�d�����s�t{%��O��M� 3A+����-e���t=Hd���q��<Z��{�X倶⊛3AhYIwR. 乗i^^�89wp�0�bn�ع��ܜUʣ[Ǜ*OI[�Cm=�)@=��0,=��#����}t���4��a��J�²S{��Jj�IƐ��,�T�#W��]�rR�E���pB��v�?� 3����ٹ��IF�~M{����v�%G����Z�VX�9�-|�)��w�K#��V�������!��p� 1v����'�8�-���doz��GKCVZv����82��bVAZju0����+(.�Q!	.�FEE��~VH7Y�hb!_(�yLZ��\플��L��9nǹ"�m����(��ǀF4{��|Q�Q'�T+[`��.ik^p����T�u���uK�2^u���A^6�*c]�\q����.��".d���|U�6���/ʳ��>U��2�_ue��N�����z%1p�;�tz��m�&g��5Q2��)��e<\�/Y�F ��$úf�R��i��`=��H;��	����.	�h��C�j`��H�t��mA��mCh5���7g���H!b ��B���̂ۥi�T͊�%u�ܳ�����4%���Uo�\�&1	��Y�ۢ?��!�zq�9]0N����`+4N�&�Li��Q❁^3��x���	S*��v��^�ȳŭ��ٹ�B�7�ؘ4Ć+y��tQ;S �/X���X0�SG���4�R:�n�q���o��-0�r�r%#�$�s.�Y�W�i� !��_+��kA4�ԓHS�rl�*e���K�9�K���7�XL�B誮j"����U�2Jw����_@`ir�o�=%�
�� �r5�G��UL���e�i�I��!�,�B��&m#�:�Y�?	��5*"��.*���:	��C��W�6K�K�Ƀ_�J\pX${�ٷ�y��0�݉��RۮR&��;0�$ioD���҄u��������j��2맜J�}Lka&7d��aV��J�l�p+X
T��/������U�Q�ض�R��(l_�oڲ�h�
.�"T��g ���^6;�����C�#~����"2X��	���-�g2x�I�"�.l�ӈ��ĩ�fK�w��e���hYP+��pn��ڄ��M��-m_x��E�F�>b�����F�M#Ӡ�w+�y��s0o�B�Ԁ�Tʿ;�R:`_��5\�?��3�����I�s��6�+���UD���k�܌lM��J���w�U�4�xP`��@=�@'���BvWYT��#C����\��9�EJ-�e?i������")#
��3>G��c���{ܜ�HG�x���Bs�|6� P�4�����3C����Y�\ĉ�ZȼX�ͣ���+�Mrw��jR���o	�ף 1� � ����B�`�o(�<�h��zP�����J9���������1�������tց,�^0��y�33�:]�<�e��,d��q���4�҃����c]��]���~:�،H�A6�y�k�(>Zg��n�Wa���%u������!B�Y1K��I��Cp�ւ��nl]à �#� �,�8�e��q׼�$ O�^^�c���u��bԋ�c��>(}�?Tض��Ȭ[�I�0�	����ɺg���zo�J�� /:�ǉ��Tj�*�E�0Ou?&eU�1�6�ȍ_�>���*8L�����S3+b�^�R ���&Y��3[�K�%2�r����~1��L4=�����yX�ϘZ����4���J4��-����c�[ȹ�ϙ�-�i�^���˹wi�G
7@��ҐɻsN����''W���-��}A�s���K!T}��dT�
r��ѵĕ�^	,w��1���V��edJ�Ӭ�:9�)>�TA��� ��T����4	X��"_�{��c�_W�;�,��]ɳ=Iܬ<(����dt��lkf�/����qA�f����S;,zv�6�s�d��טA�#`��pp��.O�B��)`�X�]t�\	�ִ��E��k�;��P�LL�|���5�M�� h��X�s��d\� �z-6��������񩷡3H[(¼��ڠ^K�H�n^�+$Z�Î�ݷ�SzcM�$�@��Qu�N�K�s���L��`Шۑc�z�w��]Gw<��?}�yG?<t*7θ1��v�}&Tt�u?!�{��hC��E
e,#ƅ�y�%6�Ւ�����c��($���=��Qv���5".,-pi�TU澒�W](��Sa�C%3�Z���{��# ���&�,;0�*`]]7�����&���&�F����b	��TlP���;�@e���g`�Md�!MT5-�L&��1Q�?Xς�&;&j߸t���� ����5�"���+u����E�\E�{;�* 0�a\�-�����˜�պ?�:nW{9۟ŵ���_�!����x������W�v=jQc��YNݜD7�_��v^`��G����%���$v|���(��vi���(^�����څ���h�^	�o����̓G�Bm������6�Lx�x,f��} ����I^]�d�b�
u��Syd���Eg�SQ���#���P�<Ø���X<�Au����]�eK�Gp�����Q�9����|6�M����R���Y��H���2Aחk}ξ��X���e�A �]a��b��2��p*��^�a�Y�Z�Л�͝�^%	�_� �Nwn��D��h�zP
�b�e��:z�����1�JU��t��Ɋ�|���r����5�sC5�LN�_���M^��4�o`�y�ȚvDOp���T�T�JfM�d�t0e�Hr/D�3?#��!YS��J��;/�j�H7(/�X2v�ٶ84������O�qXI�f<凨b�~=�:��wj��e�ǧ�r���F�/��B�y�z�㖎fO��8tXpT�jܮ�Ҥ��jZ�Y��ҬEa<˕�lv--����p��������G��T��g��^+���N�9�G�§S�w�aM"q�Kܩ�HS'�-����7w"���˱۳Ʌ����Ű������LW�\.J��Q���G��U��\�V�v,��<6
�i�mM�R��]g�|v���(-�`P]
X��g�e��&�T�`�e����.�H'�&[�Tb��[gAr����"�3����`W�?��� K�z>�/d���l�Υ�q���8��_��Ea�jj7
&�ƽ�}P�&���|�鐒�"�RF~5�N�y�g��..D�})��F~
��i�3蝛�Y��*F�דy��Q�n����խ���-�h��z�H�d�t�P!���"��a<������lW>��k�)Q�xF���[9JgÕa^�x>���"n�i[���#�(J��R��b/���52z��y	g^�yn6CZ���:;�F�?�����,������B�6z�Wǳ8�w�ن���] �U���-q����T�nvm��
w�L�OO�	�hH~��z�rH��\��	�t��ư�%�=>`�E�b� w�|��Q�z��������fy⁶9'����GS�}����,8�i��Y�ۥ�J�X�c�Ĉk�f>.��[r�0c�ɛ����Z�T�3�vF�%�:�<9�pdT�vt%��c{瀿����٣�%LϮ�����0d�68����7hH(�d����^���Sa�A���8=�hȉ��!���p��Tc|;�d�V���0����O���RL���}V�+�� �$V��(�|w��J������w�9��L��	��lL��.���M��s?��9jQ�nn�(��[�n�q�թ۠<T^��(��!�*ڪ#��>w�Z�v���f����C�m���L+wW�F�):�Y�-y�R9;>FB��?*�r=�cȩ5��?C�32�DΈϫ�Qh9�S���7gM�z����+���-��ȅ@���U6��S)�űy"D0Y�sڔ+�:2��Z��`���Ϧ���/猌'�~lļ�#�M���H�D�'(���
����}�ק�����N)c��M�C�Xx�������P��T��y܃o>�K�仛��q+��)4[�rg��\�`�e|}yv�<���I��uE�T���pW�(��r��.������;�G�v�&��������P��T27V�*de���(�ij�P���yMoI#�����$LBk� ��ΥI]��-�AЀp�B�E�I2����1�*Բ��T:luG�L��=�}�����Ԏ�C��H]�y��l��ƠS���	��Ty\*r���I�X��� `z{�R���e/l|l>_ßL�S"�x��#G���TM�K�d��#�0K��@����s��U��P}s�{w�)@�y���y3�G���U\��[~T8���ek�	��������]\f�i�x04H���"��9�2� 
��'�?��W\�g�si ���фn`89�ridI����v@�V��$���aG;OJ�MA7t>���SV��X[�=$��>����酟 5.���\0PbB�����'��/fx��Ck\��n�I.�q T���S��^�(?�c�M���+]:-�G]Ⱥ�*�^��@�q����7��3�ʟM[�0��o~������v�D�}�v{�MSP��T��.hp�h�t�="����$_�k�jr�Z�-�Å�B���X��iӛ�,*ڰ��K�&�o0C	�ft�+�E/�����ړ��c|N/9[k~֢��y���{�ml���(�������@�� ڧ�t-P-M�U� 1��ʳ��3Y �b�1^7��`N�{�IJf�7�~�7徶��b�F�V�V�N
���^n���#�Ge_H�<���+}��YQ�Ǆ1e��L�N���X  �ѴW�tߏᑞv�!�#�&4�O�_�p�e���~���H���y"��ԃL	/�0�$U}�1l�<�hK8��O��Qy��Ea�1ȼ�\�/�<�B���d����<�"�f���`uu&b�-��μ���2��N�F�]I�m����]�3m��}P�3�ht�yB�؊��B���묉��i�]�I[p׽��b֦����_��UK`��`�Cu�/ C{�~����b;q����G�]�_Zj��N(h�Y`d��fa_���@���Vs)'���&�G���b�i���aq%���ڛgq���"_��(�p��ż��I[X�����GЫY�;!$��d���D��A|�|��,�0�a�*auJX�ί�+z�:2��!d�C;9�tHnL�D(PK�p�O|�Mg<�Wל��%�!�T��*W��hR��9��?L�N���>^uY��	gJl@��Tup��"��3(�Q���D{������9%wi����.��u��cW�ϗ�93[�"-�r�N��K)��\ث����'^Kb������"�&�U�y��ٱ����f�a��b�8\R���6"��9�97��1�Δ���[l���&A�|xT�W��^�k�9칗?>L�� �p�q*�Jjl�'��y�E�g�=���?�h�5A#��
�ƺ��CPf�ޫ�����g�aͫ�F���CD�h�ԃk����X�E�N�����|�)��߭Q ��G�6�z�K������{�~G�����ե�A�!"���hJg���d��:{�>"�bl�J���r��� �Qh5r���` Έa��Kz��������Fa���5����0Х#�{�^Y���8�0�:�*�;��J��̖���h_�t�_���#&!y���Jc�`=��
�(�\Pǝ�j cp�'���h�$��k%�ƌ|��	�hY������(�� Y��Z�4���th1�ޫ�4��)^�j�7�j��4v�W/PR��b��Cf=�}qQ�9��K3D�e�p���/��㤸rN765���;������V��u�I�SuO�Cc�P�:$H|B(U�Ͽ6 >��:�c�3H�-\q����r#�x��e�����X��J�JW���0��A�W�W*@�5�u$�D (�dʁD�A�ul�l��.��=�ܫT�{�U��B �qǐ<gR0?/�⠬!�4�|q_�{i��\*�*-� ���wV=�_��N�ɏ�����X��@Qk�ߤI)���~/�)ay��Jۃ��|��.��9�9�B��A�������9�
�<�PR'��L��
�q$=^��v$��-k7� �/h�,�#i�<f�xO+��yR��Z��	�r��hڊjt�4�p3Fv9�bV����8!6���4��9:2�<�^>u)~D��s!Tn{��������K�V���0u��Q5��HH��p�<,pS��!�Qk��
ǁ9�ͥ�h��)6φ?�*����8*�v
(��c�翗d~���0m�:m �E��J
�0�!G7�\�O,9	ۂ��]�By��yT�W��d2�V+UBa�����2h���ڛWS2��
\�O���#�+\&=H�х��O��^eAE"v�<�����*L�v����iJ+`|�?�[��e���v��E3^�I�F���7�i��&큸��F*QL4�C@P@�{W�|2��RK� ���Q	�`O�PY���jmi#33��9F�#!�}��ݔ^\��E��2�+�rM��#�}ț��@���t��?��U�d��+k���P}5�y5�8�niKs��j���ZY҂���*�"��N@��=��|`kSSI���J�g!�N��p���]�r��{��.��{.G"X$�xd.-�@3�z�]n3B���]�I����{�����.�k5��~BC��=\`�RᲧ��"���8ר"B���:�~1vO+�@�i����R�0􀫱S�]��wQDbr�ɻ���mc��?�*
R��7� ��JS�Q�o�ׯ;b�Z��&��>�%3ʐmrY�� LrF+H����Xfh�dl{����?��m��q?@�^�PBx��ƥ���'>!��cڛ�%����冤A�wN����̃B��.x'i�Τ��h���㦞ͩ�~�e����UۍeF���#��$�+BQu.�
b5	
]�%��$Կ;�4���S�(/}�+@�@-o�U�9Q:"�����Jk���Q��zZжB�k+��.��P�F�!���������L�+��-=@�FV�桡.��U�PJ��@�A��<9���-[�u��(��~ؼ�����Lӯ��L�4R��^���]�(��K=&��r5l��_L%}�u�Hُj���#l��c,��c̼6����/V��ۡ��\�!Ϸ��W�m�U�@\�q� }��������5`�:�=މ��[�P5�^?5$6�9�b3te����x�>���?�,ֵz~f��I!�ԻER�Ȇ�g��Q[�ktPr��	�jlD�S��������Ev�sH� ;��K�Da7sa,F��@��hS=��˾Ծ�]�̹?���v����N9{������{^�0gC�Wq;�5l�����YN�t&��&�ƒ"�	B���M3�G��;��U��0Vɍe%�$���D���g
�K�W7��Q�z]]T-��ӋT�u_ـeSM�?�f��nY�԰k[�-�� \M�u�al�]���Wcd�i9�(U�������<��+x��"3y�3���׈+2��h��I'�T_˥h�dN���[P���6iq8�!��9q��񒨁#N����j*Z�� �Z(�A"�|������5�"Χ(��T�I�P�hv���p!���ԕ��\��NG�LW�6�Z����ɵ��c	�m^W�q�V�`�C��_��l[��ݭ�5�G��ad\�tf�ӭIU��&�Cj-߃ ��y׺�T��Pi��ﰽCB�Q�k$��@��r{�f�������ߩ�\z���3w�m�}j_�2�7������էN|�2�6#P5N^��Lo�\�P)Y+�aw}UO�n�lv���� <)�s�:�$����t����17\ծ�k������,�Xރ�� E�3W�B'x�Rĕ�9�,ΒӴ��_	�A�Ί�[���j�Bm�+^�ke���)�m��Qe�LgY�^���1o�o�g)NNZ n����%͑~��6V��?�%ˁ>t��� �|S��`A	���g޾$�[�f� D�A#޽�o����$�@�;��Yn�/Qt�(�[F3i{��[�~�-��p��n���E'�h����k���_ J�*}e�C=c����X�Cx�&3E*e��t�9μ����9f:FJD&F��lI���1��Y�&��B�$N�j[9�8J��(��lr� 6I�F�{���"���$��.<�A��@xs�OF̰|~D�!�nTx\cA�h��^�0���w����T���aeG�1�g���.ln�YqQL��"��������)�qǕ>�S6���;�Z$pKw �ӌ�6P�"�����h0�{�a�y N��__�f�b-|�,U��2uo�����I�L-ŨHE��^v5W�b�qܮ��-��♢,����2}���wl�/���v�4�?x�BL����/r���uO��_T�i�K������[�*�1Y�HH	c�̃	�t�A�X7/�ˈdI��K5z۷IT��n���R����b� �"E��'�s{����
�*���d�?İ����!Š��p�7���pЕ��/�s��I-A�z-���
���H����8h����~�g���`Ŀ���q ��n�9 ��Ė>�<X��@�^�Tx41�#�����}[�����
IҜ�:�R<���@e�̩�y�����L��uT�����\����ƥ�g�#�5�L9Y!���NҕQ0Pkyy4�6�P�\p��������լ����H�(�:.���)�����j�BWܒ���D�o]�����s�I�Kߩh׻�vlv����?��/��o=KG$�5!�#�tj�i����b�{�2���w�t�6�!��/"�dz����h�7�b͊��I ��ݘn��"�p��6���S�_�s�72�ﺎ��iV'�Te>�+û4�y}�W�X�9�'��Ƿ��Pf3O94:��S�å1�zR�Σ��J�\V�PۣO7�F�'3�AX�j�r�,�4S���}�G� ��RtYp;���p26�7�˃�����s��3�a��P�� �R��{�Lѩ/�˲�e46�퀼(}�S��%}��o<����;=5�ɶR_-U�l�m�{3*dV��� ������w���v��Ο��bF��r������&�5�Z*i0ݝ�܇ �#�)ilßB�a��G]?����dƵ��5��z+�����_ с�*�r� G&9d����K���r�p���1�r�Q�h�z�=!¿7sX�Dŀ��P0��j)�Y��-֟[h>)�H�Xd�br"��!=���6eQ$��(�dǎ�c_Y0�޻��9�L��$���ŝ�b �\�^(, �3����������~���{��JZ��{C�]x�u�=�8�U�j�h�B���P1��\����BCF��i=��N�tF�ClR]���2��8o�MJ�5�P��}����o��Q�ɷ��M���0�2�k�GR�աr.̦�o,B����Ϳ�B����*�mayB��J��_��P��~+s+�/�T�O��w�첣`��LQK���1�d���ؾ��$֎�M��R�#��������.�E^$n�&2�S`z�}�*G�{#��U��R�֪NA�����#��Gxۜ�$���þ�<�-�L~Ԉ.��Z��-����7H���C���%������%X��>YR53hFgP��+60�ɥ�������]�~�s@u���ἲ��������`��<��÷��{U�Mn�)țK�;�	8	�=���ٳ�(��&8�@�/)+�������G�3V�u �;�y�O��ҥ@���9�Ҋ�k�Y �uawjW��p�c��,�O�ȍD�n�/�Qu4T3��7���B\?� @���wC�K�́:|>�������4��~v���!u���j��At)ce�p��
!��^�R��V�'���J;`�`8.�@O,N���H�)�Y�@�J��ս��AH�gH[��F����M`�K1�ߒQx��nPV~ָUk��A-Rd�������	��Q1�K4��*Ǘ��H�ի�E¬�\E���(s��X[�T8�1�a\=�Q��{�*:�����h��R��A٫#�^"�%�iQi@�q��?(��;���:�VeV9��y#@�2��!ՙ�MBߨ;��şC((:>|ʾ
l���1��ڣ�s�Wzd�҃�u���"(����Y�T�9��dڋ2 �{g(� nx��E�4B���sm�L���*r^� ��y8�t!#�&�
�pm�^m�գ��;��w7��Z��wI�~)�Aܔ\=�	Ab��"��N/0��/ƋOb\п|�����bA{H���5k/�g���u�w��~�ث�V��Ͷ�N��w�EJpZt�xH�=�Ag�������T�I#�a<M.2n��v����6MWy��vISxz���6�'��d�YC5�q��Rk�L=550T��z$��_WB�<�����KQ�A��J_�B�W`C#���ϧ�>0�"v�'PM��Ӟ�]�*	�̿���0�#�Q	� ��0�ٍ_��G&��T���6��S�����*{�x]m�=� Z��!����NRt����W!`��t�O�qY�@���H�kk�̺�	�o�.h�fr���~%�!�c���}�
���W�w׻|���$��t5�@�e�n}j���iClg�%��:��C�N�/�U���ϲ6��d��ڸ� G�5fB�������8P�Q1��Z3s�>���Uk���؇����魆R��v۰�hum�0�py�c<J���=
4�EX����H"�h�Nb�GR�� w��VD��Vw�x�P�����Й����p�G�I��l�LP̎����1�HM_PT.���$G�����@
/�mT�} v��kP�ӸH,�7݁��ך����m$2���)0������B-��z���2ظ���E��77���P�4�a�{Zf�
�x�a��Aܚ��<�2�TG���D���|&�>�P]rQ�kvIT�K"!(v��_1%�Ȳ���:��$U�!&��3+���Ӏ`��dJ�/����!��|���2�-*G4�0�m�-�yND1]�G���1ږ#���&�@��Q�
R��#W[�EU�f�<˜u�ay��N��ڟ`�2s�ŭ�¢����yD�I>�,a)V�qG`��(y�8���c��[�}�-;�
�!�'F+֦͟$��md(����P�=�����Cw���?9�2V�L�o}xKN���c	��#�R����gӘ����\hb	�z�����;ՔyWͺ��7�{��	�X�7L��˻�p�q�%ރ)�̷��,�h�FE�h��m��~�)��'@�#d� ��4ڢh�3\W���N� Jf���M����*ĜE�'�6uW=�V�gtl�k�sZ~F���8�=b"�|�n�V�J\(>�
��Փ�N�|�T�9���'Dy�|J�?�G��d�.̀	�Aoz�ol���i�򩬶\�}!�Nb/����u���N0A�$臂g.n�p�5�
��V�}v�����e*(��9����n[ :���Y�+hf����[/�uP��I�	�l��j )T�s<��zn ޚ^@
H���6��1:P�R!�fݎ���Ki�B�z���u����k	�c@��Z��v
�j�/G6�3�k=l9_�G��u�3�WO\�Xe�\]��X#�B-����)�2u���)�c�/~͹}�E�L���LfY�Fz2��&��-�q#F�K��������R+I�΅/�֑;���c��A�_��"15!c:8 q3��{���m�n����������7����
hX"xg�χbq'���hi[z�	j�C~���R�� �]�+O.{���=!2�aO�2u�38� �,*�s�`d���eᏞ�i��u�z�贩���
��s/	1K�Z1�	Ժa���ޙ6L�:5VŜ녿W3_*�F5{u����)�n�Ժ Z��	hhg�y$K��(x@��ӂtgB��T�Q�^���593�ݝ8Z�:y�]���q	If*y��}�WK���J3 �A5n��6����ٽ�9�Zc ��ɡ/�S�Sy�A�k%�����h��������!GaW�qP��7��?�R���e�/B�H}IJ�P�Ǹ��W�r�o1BC��C���M��+�T��~dp��z�v_���U*'����L��w�D�Ĭ=D�sl�+�0��>Ar��go J��k��_3B�ؐ�4��88�Qw�T0�R:O��X��?M\���q�B���UaᓺM00��D4x$-�E���WA���d���KA�'�����1aɌ��՝A���|��oq$e�X�%����:�����E!J�!�#�/+��P����xy���retk]��kℳ ����M�Ls�Q�����>Ƒ�<@�h�%��Y��R5DX�)|�ۦ��G:�ݪ۱3��CBP*c�-��V��|6h"%mi<�4W�qh3�<�BY5�߶T��1��(�X�̚3��]�
�{x�>i�l�+@F��0�dP��&�� �8���"U>����^�?�H�^$�RPR!��H�_���`S��f�7}y~�f��x�Ƹ�����hV7�ġԢ�?�B��D����^y��>�_��C��_��=�S�����)tޯ64�C����ɉ�"�_TMT�>Y&h��3�_�rv�l�{]?MC���hɫ��)26�<gI`F���B��f�+&���&Ge>�-|�������W8�s6`"t"�gHqO�����&h|�p��

N��<�\�W�Χ��C�I��ъ���,$(�y��)c�,�9A���u��u>b]�f�����B�髼��GEk�Z��J0�j�
��>mmCf�؎bx�d�
���pu-u�/�d�����tl�A��h8�1kB�.�?bY���8!8���q���.f@��}�OTsKD�Ҫ�� �VIeo%G�w���O��q.��ZF!�{�^ƾ[׬��S���j��y�(�:;��,a��/����_��D�����j�0&'��0�־��IL��O�����۠�����`�6�{���PL@����m��`����M%�z�yk|����������}B�Vd�d<79{y8�^�-L�E��`�9�$ɨ�53}�8�h[J��L*L�ܣ"�QB?����BC��E�v��>�w�KC1`���$dv���W>�/㩫���7+l{8)��R=2!�qV�ӽx��,��x;5O�Lː�"�VF_���s���)�����M�=VB��V�K�	�����b&��1�r+w�2�<��ML��M��|z|k�ΰ���գ��]|�v��[���=\`Ó)�@[v���޸?�IO�L'�A��=Fx�����$��/�C� ��c� ]m��rN����L��Li���Q�h6p�h��;��%C���/H�IuD��?t����o�>C��^��މN���� �i�߫]��w�" ���(��2��� ŕ�_|�f	^��T�K�fֿ��l�K����_�j�k��%�c��Ym4s<��H:�ЍX�/��C˅��q���4���>J���ht�l�Kb``��:��������oE���p��"��}��9W:sE=>���GY�;�ւ�M�����^��8��Wm�
��e�\nL�S�;�[
r1�1K%-��t4B�J<�*��(�g�320f�g�#	�Lv�b��	t��Kذ �j��f��k+�hڀ�$[�F�	�GM߇�ȱԏ�y�C$��<ׄ����N���:�%f��x `�T�'ܻ$�BTc5vLɝ>���@*"���j��ĥ�f�𦑗����R&���r���{�`u�[��v���/h_�J�fG�O��I�[T�-��jܣn��)����r���y�@&p]����E\E������̌��n.,�K����;��C��]-}�o���g� ��R���vᢣ���<>�s�]�%�[#��47�2B�[��f������~�?N֮p�������$����32��5Ԛ�Ah0��|f/��$K;��]�:�+u|�P����ϯ�����:�@�5qur��W���y��yx�A����p�~��~ȁ�諚����Ʈ�$%|�R�a~�a+���c|�l�8��U}(Gbi<��T*�r��cY�9\ǦB�N'3���)�A|����=�Fk:7�&�s��25��Oc��|TN��إ��Ɠ�nC��VҶ�����Y��$��Kt1Z���4�p��
��FC�|s��Q]��gPҪ����Ǵ�v���C��_�%���WkP���~����_�2׈����u]]7~����{�$n�ecozf���f]���6�=�ec��Ul:+�(��F!� ��
|�c^�;�g�ڍ"p���MQ���G���"2�+; ���|N�z������gDF��#���'%~r��2(C�zt"�|$D\nṖ�C����������2��ܰ@��0(.���п-�^���XH'�=SO<�H�q���~��,~�S�UʴC�}��\C��M�+l܁�lmIHr��,@��k���ᢳ7�Fp�J��F%؍��EkPwW��¥�?,;Q/�T!�Ru>�}��Jr}hF����*�Ww�j�����ޞh���t�c���ý���`�o�Ow����Q{��B������� ���3����M��k,Wr��bX���\ ���P6��y��,�1D�:�X%��"�[�� m91Q 	����a���X�#��i�FӼ�2K��x���*:z�tY;�.A��1�է��*���Jh�W��z/�}t��#��FNTs�=���ꦽ/} � �JB��m��n��9�����U��&�{6	�B�%��??Gm�)��3dF��Q�5��S��k�E�"�N���Ù�H˦G���{#�V˽*-<9CWE<Zͺ��J!���U'$�<�M���Kq
l>�d�"�]|!�?�PI�#5`"K���&��5w3Ũ`9�8�覮+�C����1/�Ylۖ@��k�n�(Pkʍ����a�%iax��X/�g��Q��#�������fC�6�Ζ\�9N�z����,���re?w�oRa� ZK_�P!L��s�tí�vǅi��b!�W���m����*�~�qe�^k�� >�J��r/���؄@��+�ge-/e��	�.� ��=_�v(�0�+y��c!���>�)B�geB.�����|�p�lK"5��ʘ�.��W��%5HY���"�b������A��3=�cS��=��O����;붻�F��êF>?���"�0��`�����Yp��1����v�s@��-M2n��0���>j����܋�'ɠ
��NxVց�ݪ^S:�9�>�u,���wB�D��u}SA��o[=k�u�|��W&l�L��ON6Mou��J]���x|�v���SX��:dC�,�Ct�?�����^��0���B`����4ٟ�fĆ���D)PƜ�W��3�2��I%�-�� ���)��������V�y����	�}i�/�0�n��.g���*,+��V�S;�bLu�ˏG�:�.a#r`��E���\�A��S��wΥ�y0�Y��ӝ�=��� �4�Fj���S�_���e�6��6��..�eNu�d�EƣOb%`��u�h;]̈C�"K������P/t����S�V�[*at:غ>���${����*ƒ�o^���?O��kN���۟K�b���H_���Hƣ�(c61��Ԡ�M��G�-��4����'�ྼ�G�h�W�fI�t��H����g����(&�I����_������A!���M�9:,��5��n��=9ϯS��^�z4�2�qcl��N~�9X7&�b[uDtqa
t|	#��5Q�h�'��M|�2êh>�[աs��I���������C�`.�����l~*\��a���ܾ�]`G���uƢ9�޳�sдcM���>��g�FYdd?Up��+yq�ab'��R�t���:V#`e�ڡ-^�g-�/�� ��ٷhz���Ө����l�^ZO&d�X2?���L�80 +tF�}!�.����B�Wŕ�H<���K׽"�k�*��;:{�G�]�>�1UW��u\�0����W�u�9�=��c�]ό�=2YK�xA�O}�^zW˩��l�Π[�"I^�@~�3���{.�Ve_�]n% -}����^�r2h�+g�'�aF��`����:×���Xv���;�lF������.���{�uoP�׶��@�X���A��ԭus��lj�2�'�HeB�_�ք��9����X�S	���EG �CD|���5��2��j>=��U�b�/{�5*�I��NAd�y����bb�Ujo����7�Mo��DavJOԈ��"jf��m$�Sg'����1v�i��x��� �*GZH��#YY�=V�^�S`=j	D��[E�R�H�(�)�.�
���xk���J����o̘�Ҋ9�d�Ԟ9�zE�Bx,�ef��u�m�'7:����	��\�ysLvu��v�m�Z���3XaSzט ��)N+|��aI�Ε���%�kM.vh���bu:�/3��K;8^�:Km�\��@е�u��l+�����0b�w�w(_c�v_�ԁ� �Vj��8�i����Z��P疯P����������������9�+#P�����7v����IҰu�B�,v0��jx��B�Z�2��ed�+ e�֙b���L� ��
�Ym\Et����l�ⲯ�7�'�Q � =N�E�We\����#4�܍�}1��.%��@�#_�H:���`�W�K���m
����+�1׶���2S�E��p���T�#/Z5W���Af�q�12��o��_�)�-��X�&
nl/����V2I�섗�q6C�0p[��0W.��ԢIﳅ�q�yMg�I����
B�hS�*�3�j�6Շ��-)\ZD�8�" 2Z��$�e��-4�0<��ul�|��U�y0-l�8Y� gS��]�3`{~m�W��Kv�{ѿ���T��E��W��vrRy�_z�&�ASZp_��phR��R8��x���5��줾h�v8k��|D~���GM�Ϥ���ӂ�T�#ò��Z�Lx��V�1Ic������W���Z���F9�2�֚����M�k�Nm��Ũ��:E��S_�����J��~^r����F��l��ُ%<w�Ś�ZZ����%{���c��b��2v�H������w'~��:[�LH�� �j�܆,�:�u�P�E"ti��F�Ao� ����y{���(\����h����;�Ս��ēb<%�S�n���>�����ԙɲ�?R�k$ ԷɒE��Cሬ{���lj�	�]nK}p�|�]aL�O�,I�-[��k�$(2��6@��!J��"��K-�0�5�Q�CUdM�I�/�.����V��Z7�1��C����I,��(�ǣ�,��/h�����\ÿg��#�7�;1�JЌiѣ�T�+|�U|�����6H��&�E�.<��Q�Sʽ�d1�F-Dˣ��PFK�cȄ�C����]���J������o޽Ѵ�J��VS*T7!�(y��������{q[f�r΋LD.���~H��];�١��c:Iӿ�8)����6<��C�����]7�ݮ����J�
Z�5W0��5�l�`H�sf�9�{@\�A�/��BOZ�h�3췩7$�����4�)u�ˇ���6� d��&����_3+�d��1H��������v!�N�9�p�p,ǉl�r�7�A����̄1A�<K�V�?p�C��x���R5�ݥ~7Zƭ�Nc�KV��U��s��|_��6�	�#�R3=�ێ�H�_�w�%�P㓁QF>�3���>��(�ZPq�vߨ^.���k���d���o���$V��_��L&GI5��!s�DX��[����MRgz����Ǚj*,�3W�H.B&+�Lq<�ϛ�`<jJ��6({/��{�^�����J��˻���Le��j�f<5�¹�yԱ��n Z���.u~���$�������q������/P�{��.��A$��,��
�Ty�D��ҙ���Z�T�Jx7��za�� T1G�m�tV��W�Y���[�����{�M���Y��
?��ĉBy��-�Y����4b��j�lqf��4m��F;� AD�m4w��X8w�Z6���&']S�������U��އ:{��x��sox�&��o�k����3���?�_�s���� g�*+2n1}O�	i��y69�:��>u8<�ֱ�9~5I��F8�Z�|�R(D��5��"R�{��x���NZړ��l�/����Ll��Hi�&��&%7���=/�˽�Ȉ��5�x�r'+B�n��ƾŲ�q���9hu��i�&B��Ɉ��g��n���{�w��9�����dZ+
�K��2f���u���ȑL�AZ���S���z��V�" w��
�sy$�a0&s��+���&��=����������e�~�|��V��M:Şxy�k�f�J�*��h,R�1{%�qW�x|�8�i�����iR%��x#FĀG��m ��,��&�x�벼?�M��Po"��O�ى�X諒d�tQ���!>��Η6�	��S��K-�����#J���X�{�m<��_c˸C��FlcJކ��(x.3#�QT�ã����p�Qg�%�5�>��bٔ�URT�P���D,e��˸^4)I�R�������ҰG��b/Q/~R����M�un�m�������@���=�[�hT��qzW�8�B�36nP���Y)��|�!��ٽ�I3;~�rl��^�$lz�a���%�/���i�6yR�y{9	ۖ0�T9
��g�g��(ȩ&sǪMb�Uk&a�ԣv�rQ9�����nF��OR.�z�Y��-���*A8�����U5�����C�b`g15K��8�y7Ų�>��}+eW�����<�ִŸ��:�.v����N�:aP/����w��k���^z�y �bt���-�� 9���g���~�R�M;??*-��#t.X �2��t�YhԀ���u��F��4�:��� T�����p��(�s�Lٲ��fC�@�t��t�����⩣7�����97�:o�E�zn����D0c���Jw�A3�z��c6_=2.�[�.1G@��?G�E:�j��%5����-5l�!Q�N�ac�a)�z&BAࢧ>�SėT=~v��!u�	��L�u��DoF5�>�
*P�T%��[�u=ރD<i2uǴ����0�[�b; �'����%g�j�<��L���F��A�zøV��*X��xÕvJ�n;�w~�����Mj@?���u*.h b�	��� ���ޭ	��]�D����x����]�K� 2��(��'-R]�w[^Bc�@�A$Wb�
���0��a���}ڭ���@�|ݼ\%��g��0�{�B���w���՞#X�XꛡZ�j��KIs֣�g�es��6s��q�!Ks���mr\.���̚� ZJn���Ob����B���(	���+�g�s����>��ƯnB\����3	�����12�A
۴�!��*�Ys`��)���V~S�{\ ���Wm�\�˛����e��{�, -
�#��<\����yY�i���3 �ӭ�	�S�RA�	�R ᇌ8t(���+j7��5u}��;+�����B�2|#�#�z/!�{(Ec� �_e��k3e;�7��ъ�?��ܘ�s6d�����j�?1g��ݭ�_��Ip�����J#�����I�嗮Y���ר-� d-c�Q�z�&��§�0a�1��xG��k�6��Kp�@Oh0�<-�4�;ij~��A��Y��I?��?�'9SF�(._����rH��0k{��zD <
c[eϴ~�q�>b�6̰��8E��A<= Kp������o���D���=�~J"�J�e�s�L�����R����R���4ڤ��n�LTB�9�ړ�z�G_y�����ym���pTBB��JQ��ݮt�;1I��jkztN0��>lj.M�]-<i�j�;B�؎�餺���cKJ,M
L:��*�9�qb�㌇l,~��9)��q��eߌ��2�͉�$��;S���_Eol� �3qe��~���B�Y��Qh=o����7�)?�Ĳc���O���*���s�i��:��_�3�S����٘��w��V�f�r����S3	��#mY�N����Ϲ���s��> k�9���X�ˑ���YšQz�GK��J6I�Z�yXs�N����L�/�Z�^nP*�ᵈſ�Z;_aJ��tq^T-��2�?�d���ֱ�F�;/8��+�)]��������puAq&+�Kw�@3�ϰs�~�#	:yj��� h@\|9�]��0>]u�D�PjHm�|���vqΥ����Ô[F�X��!�ǢŦ_��v���2Y�Y�dsN����.���RMlQ|�)+mZr``��-�I�d�yr���qױ�������^Z� �:��u�q�����ZS�Z��U��/38�P��3�Wۧ�f���mc;�b�Ǐ���o�"��
�y�(Iz�{W�����Ǆ��yM�4�R��{�:'���?c�oH(�s���Ǵh��O/��,H�\���oq�{�����=�8�W���Y�?��kv�kk���Zf< +K(�=��C2��knY��@�1�0���́����ķt��̃ ����}ټ6�㬩�7=U��@y���.h����vi0&�A�Ռ�*�$�^���&���.�Ca �w��7��|�_��f�}�o��"V�����т�ґ'B&٥�ep�1R��@!��@MςMG%���4+3x����v��t�3N�$�X�1���D�ǵ������Q�H|��U;�nPu�(T���{�+n�|��ޱ�[xa�T������jq����pD6�I����\S14`X@��43�@Z�����[�ف(�(� �.���^�&���,w�|_�0��)�����'K	¼~����FP�?Y���%�-+J7);
Q,��Fˊ�0q������.�4�:�c���45��ͻ����ʈ�*�l)�#�;�g�{n��'��;�*��3+���k$_�ֽv�lv��O�k���i-�K��K��cұY�b���&5l�B���H](����{kH!�ج9��1I*j��m�C�*Y�"JM;j�~>�7��#|`"�M;�0ث?���š���ʯ�E���¶g�x�J'�n����˅l�>Q"�Jb�銌D���?���)��)V�kn���M�U����,b�.������LV��� ��Ʌ�LhTk3��U�&YNo-ڌ�SG]�:=�Ąs`��uļ4����!�٫�}�ڋ�o[K�������R�'
��gvg�||1øY��{^�s��������t�W/e��5bw��7�8�X�x�����9�1���0���eBGjGڂ�?K�L���r�J���NRJŅgY���rA2{��G6I�x7�g�0�z$�mj��T�}6t�}K_@;�+$_�IsG��C��i��|��OcE���G�
�k�Ga��S_�8#!���E�ﵶ�-�\Y�A'��A0yl�g���e�7��zQV`���YF9#�<2��<A�cE<'(��r��4l��a	����2iG\A&n.�n5���.
��@\����˺���B,(y������9.|�ٽƱ�~ܲ/e�t+�H�Ҫ�_*g�+�4n�����'�޸��=��(U�cv�
�G�.UӲ[�ѫ�ɋom��85�#ň���|vD!|�˕2XX�~ʋq.��4���ԅ���ŝ��� �2�����3N{hŲ�!�������eYN��x��P/��#J�`]�*���A�����	�m.y3�h����<���f�/k�	's쾝qJI��0�@����e�$'�qS��%ʽ��y�%��r�)	3��o ڵ&�o�^m��-x���Jק�Dր桐�qg�b�k1t7��m�"�T����wi�ڹ K�A����#"�}�������2���O!Q�Z������%P��.�'�҄4CEGL'���R*ܢ��;zy��|�)��e�����tG@��oW�m���h��݆�e,_��}�'��Gɝ�t�����.�U�4v_�qD��ZT�*x4&b�r�l]�Rp�/��\��ԪZ��!i>eS�0�-h��)}�3��*��(�����^��փʜ܃e]� ��[����햗��=y͛����2��h���_`ug�X�������]��614=�Kka<����7مGI�X����XM��������v��m.#䮞�(8LI�j����_P����/�����6����&���S�f�#N:�Jf��p-��z���c�H����8T�49��1k�hѺ���C���G_\P�p4MF)w,把�
���z�S�jtz-A�����얰�i� ��qw#N�d�s�M�v6L����S�0^~U��ojs�y� �%��� �i1\t��5�F�X!��e`�E2V��}Y���*?U4 An!/�g��&�Q���w��v�\���"wJ���BO��[l:_p>��7��٧�ed���l��Wt
w(67�A�ɘƻ3v����A�	���N�����2�?�2+��"�z@M��#�W�5�V؇5|��� ��7���qa�|B����s�N�O�OHl�n�N�xR]�1�u�#�k��)��Σ��L)���Vܗ;M��'�~l��(d�h�H�����^���)��E��"��)1z/�����c��6�aS�/#ӢB�'�w����e�)V ,x:
(�^L���k\>��\�Y�!���З�i7��cS2k�xI�����jʾ�8�����K8I"��H?�SYBʎg)�~F�6�s�^�2�e�R�s!!~-%�_d�v+*�����6�z,�]�Iт1B���]��\�gj1�!a!�s��?&yAi˒��a>�wT��
�"���w驲]Ix`=���*6Y��(�}�WQ��g]FHr������H?҃�h�{Q�58��$���4N�x�T8;�Gy?��7k�����u�\D��]{���������Y��N��5�k7�2��<QZ���Y���4=O_��<��ֿ�#R��\hJ�� b��W��.
�Zy��x�2��4��X�R`�]�0U�F���Gf��,q�;�'���_>%�۪�)���qz�*Kڟ2	���0���n��Δ�4���ڎ�1�����͊n����E��մ�iu��Rf{��^���&>���wd&�"�@\�<�!n�����'r�TA��-ї�l`�1��waY�hs2����C��_��P:	��V����ZկF����Qi���������Y��z?5p�ք{�{�����f�`s��+��(�.�5j~���Ug���A)K�%�FnW�����s��!���(�| ��{�t�;��r�D�ʆ������s_S��`��kF�k������<��9���7*xZ-E�A�{ �R���ٝy��ӵ���|TC�F	��!�ٶ-r�xH��2blU�P���s=�	�ݮ��ýW�����)P�Xr:���]�]b�#G�M �ƐKHw"�/������ꝕ�� �nn�֢��V�H.�7��D ��rU?����L�j[�
s�d�3�X�t�ss�oc��]�D�ș����w@u�nD4��4�C>&'�Z�H��Mދo��|����%��/���@C_��ɡ"�.�M����p��+�:���Ck8T�nj�P��N
��a\��ƀ� ϝI����CE�ȕ��^7C���_���=���M�2��l���~U�^~@V���O� i%�T2Ll�O���:�!��p��wpS�]~�PIt���]���=�[M8����\;~	�^��^���~ I�fʩ��{�L�ql_���>� s/.�U� ���=Y$��"ǣv��w孫�ڷ���}zoUXm�l��fZ����A(�_��>����2�q��7_%�Z��c%`@�ųM����&���'2 ���s�lxh�7?�=�3���;�h���+;��	�_�x^5	��å��[q�`qؔ�t!a=�6�|��;��i�4�s]��W��tϩ�b��}�� �C��g��o|8�Ɵ�d���]p��Q�)�VfZGqܔ�`��'ɭ8=�e�m��6Xb�9,�0�ɇ.HuAF�E.	��1��}�j�K8���3�gu��� ��}�e�mo�����:$�>|�t��,~���Fn�S ��O�ǞI^�G�P�Q�ر8l�\&�)@0NF�IY�R���^,�M@wB����H�0������P��*$u�"�Q�W��J�d� R	��J|���T��it��B�V���;:�&�Ϥ���o�>a�$��Q�!E�Q�f�	���:���3S�k� _Ԫ���v��:�۳��߻@#�hc�5<Z%=�ʄq�{f�_�Ŵg{17�$���B7�u�Oݢ�YYA)���)�3�o�W���B��$�7h,�p&�f�[8
�>��\�Z����悿���d1��Z/TP��n���=����7�\HIݪ��b�]L=V�g�E�	~g���q=�Vxg�=_ݠNAn}ӥqr�#S�WQ{�����i@
PD�&&�|L��Du��;�PE��abMG?�V7pAZ>n��1�I+��d��C\ͺ�99�v����T�C0]Z�����t��]��������	�J���mdl��nԯI=��ˣ�XM�Rx^~��S�����u\ˆ��zS֓���wyK9i�y������xQՔp��6;�b�D��8�-�ߢ	���B8����	�Md��P=�Nj�1ś�輥-�78�O�␲V� J��,{��D�b&�¢Mr�z�q��v<�c�����Kx`�$,���� І��N�̚'�����Ţ�!?�Y�E���!W�r�ed�?�;��!����L���@�:���8T�.��Ĕu˶/�0@�c�wj�Mx�zw�iᲗ�)�i��l!A}�/Q[Dh�m�£ZԒw
�?]���s��Uy'�J�M�;�n���'}��M���5=��bm�6N X=�����@}z���GG�2��8?C��5C�).�2���7�]&�p�������|�7��2.�'������>:EW�cϩK�ϲ�^�;۰�����[�ڛC8X�6;Z�7Jߪ&	��Q�3�7NM�_���*v�\e�Y�� �������u+hp�O��%;�H�鱿�`5��H��8�=[�	ݳ��,F��<��2ܖ��>DuD2[�.�1�au�=�q8��I�~�3�;�8x�w����г��!�-���ӿ�9n�iytW���6�W��@�а� -�Wȁ9��{�K�ޢ ���5y��kb���'�v��)�Fj��/�&�M
�b)4���D��?l����B���+T�ˉ�I�g��}r����Q�O�7�" t�m�D�����L|�S�/l�)@>���p�A����ZuQ�Ğ�����\D�gT�>���7��駨t�`���`���̆�wLB-�C�|�ՂBJ�Y^
��݅mÉ?�+�Ꚍ�w�4	kS8Zi���{]-"s�4�.�AR�au�,H@@�x�����fi�CKw����ߗT�m��M�P�R�|�oB��X�鮆��5�!nٱz[�x귂d����*�[��r��|��A��� B!X$(��dҶ�#[���Z+|�2��9��T؍�خA3~\8L�?X�{������j�'͏�:�����J����7��rC�?H�5�R��MӚ%P��R�f=���`�s�=l>|���,3��q��PS���<T�t��%�Qz��:/�����{q���AY��'9���������>����!For�	�j��(�e���ݨ�%��ZC���iX��)��O9�'[W�&���ؙ��wWN}&�&~��r�j�$0�vv��
F��"D�$n:|ܙ%�<���0�re�U������p޹��V6B>�N�!�!�Y6��r�� b˒�z
���컭x%�T�W����T9Z:2���9�M	���v�K�fz ��P÷g��J�OS�J��r��c��o��}\��s��(���PI��x�$ �O���	�̎��l��c�O�-�Y���$)!h�:���ˆ����t�5wP UxpŻ�9*�e2�'�3M�VH��w~+b�U�>��r�7�@0�>�A��4��د�;ራ�u�n�"�3P���R|�.�W�צ�zp�g�|m�g����n���'��� ��=����ۤ =�(�(�O��(���]k`�qir`�-u8��g|c��W5e�n#| zcB*71��V�I��GHH�*)�W���F�ai[,�t/����r�g"��[X�qX����y�m"�8֏����z�]�T�DS�3>����l���+��\o�d�ї��:��\�ŏ^�}ٴK�M���3�NP��<�m2���;�:��<bH�2�ZФ���Wv(2�}̝����)���;c�c.VH��Y�	�2h��B,T-�$X�X�`�8�7"�[Kk��5<g���D4������Lf�8D���%p�-�kj�
 �!^q�Y�w�A�����#�Zo>�>_�ï#�_O�I=���I&���#C�2��P�t��!����z�%�ٱv�����I%��>�.hy�7fe=W�ȧ��\
J�1��l@ǝ#��}�fE j9�G��p���G5&;�P����� ��uxD�Q��VxK&�ʨ��!�(�)!8�w�2�&.����S�Kp��3�0�)�_���C0�b�g�Z��ɑ�K����]!�>�g]A����u �/�b�G,��/rd/%=�P�ѡt7g�A����t\�e���yh��c0r@ ��w����p��A��#�5�1a���1�\�wBu�?~z�TV �t�	�����4R���xEL�8d8#��&�Y�����2j���^ZX�F.���'7���!w������F���JN�_��R�I��	¤�Awt�gq
:j�;(��͏C��yb-����<��Sa.�t�)�C�a~�w�V_�
9ٖ���}_����@$fy�f&n+���N�3w^H\ϘVYԲNf<ʟ�$�N����F��o���I@�{���Y��} ϟ�����&��Imo�#�^��!��C��
��0G�*g�܀��bv��<N+l��J�%_��W��*=�K��{53ZzbЃ��iV3��a��n������� C)�r(�>�������q�+����εt窡�����g彋W�Ͱ�2�N'���(��3b��O1	��+OU0�����Zj0�d�E6M5����Y����	��L,��(JrvA�{����R�>�-�B	�����ɘ �L�k��S��qu�U��Z���d����W�iD�\:S�:�J>�׾�y�n�.�4}"�N�N��BcDY���o���_�9K��G�HKC�x�d
��Ė���?'�yT�*��HH-E�OM�n��d߱M��!��j y\���P,x�*� �&{�}~��8_�q�հ�C�i6��,v���x7u��B�&��`��5���$���Q�Ʈl�F����U�	�ۯ�㿷���5j�-J]�Hp$N�%=�)���q ��wb%��=�vϿ�;��O���L�/��as�������A�5��{��-w��Q<�L��ҙ"3�.����wˁ��%>�`�8h�p���/
$y�D�>��_^qO���Vn�K�&\\�!���ގ��7��P�4��&�)z4"s TV����&��~�u���7�3'&C�$E�?�}Ժ+�g��9~�k�H�q=��Y�Fez����z�q6]R i�`ǥ���"��ht$'	�4�}�g��jf�n��ow�X���đ-"j�)x�%_���w��.Ӽtܘ�]"���U��H<�|�H�����J�}�+2�;œ �;���قt���<�>g�/�X�V�Q���J��tF7_���A�?72mC6w���L�%)����P�YX!�E�����?z��vhHV���ˬت��ލo5xA���Ů2H�kT�#y:9�q�&�m�iz�O�����&<1�?"�9PRI�ӊ�L�e��U�N=���*���Q��L���Q�y��Z�a���.��J"�D�]�S�bbQ�Ph�>z�;��ҩ�U��w�4�ZA0U�� ג�Y�ګ?��+3J앿
B&3���^�$ ҩWA*��4�c� A��{.m�3�>w[��^��xl��P[C�c�e��	�q�l�pB��5�g�O���2��V<���b���<�0�n�|���jq�B��n��>v��� ��+��<d��_tz@к_�0 B�&t�	��c]$��_�g�Rgl*����wGN�0�׶o�r�4}lA�Q&��4�x(���[�y�G$�ģ��i���<���K�mu��
�@X�\w�Aa��;�=�h$I��z���6~��G:�z̕�p��_�����\�E��&���t5a<	Jl:�{�$�u-�_����,�-�& ��vqr}<�\���R�:��>M�ݷ[����6{�Z���Ȱ�C-�b�V%ޝ��� �����,��d�q�����]l։�^̸�-g~�����k{M�[�J����s�V�둃�A��V���끘��7-�8����񰑙.;�ʥ�9ɩ��i��y�c9�7L;L�݁�#����3)3��x��N���yY�	�	.Gy*�+f�����@R��Z�l��=L�Xʰ,���2|�l�o��K3t��⼧���A��0����9Ltd�#a/艂�;�;M��X5��N^'A�2a���:yJ��a�NJp`�f�u����
��
J[^�Pc7X&�bBn����������5�����$Hl��^�Bi^�h�Q^Ȟ/�����G�<t�j�����u�~�S�$�"�Vma!#v��$�/0(�@'�"ș�v/l>=�>�'�#]l�x�^S������Kg9;���E� G� q�P��E�h5��qH��<儵���E����O��d] ]��pf�dR4�OCV3��z��tK��W�,��K�D���-`k�v�\���Iș:��0�U�P�U��;�VN^������\!3����F:�DBY�6�u�n].o�2\%�*?��kI������&�c<ߘka�=ۚ��}ɨX�Ԟ?U���nt)�m�`�"&%1B���~��[(��I�~iO���5R�gmeF���O�2RԆve[�˫�)�1ً��<e^Cކ���K�5����	s�xi��v���s+���\��T+j ��̴�u����r���*�:z�ΜyĽ'����`���}��A��y샶�sTaA� ���a�yV��*�$��K���ٷ�p�����ݺ����)a�]1tV��Ȳk�W�%�.�;|wu CRf	N]�Et�9Ċ����%[����%Pc�J��;A8{t��˗�j�#�d�x,�9�T��@}|��TnZl�S�7\�e������:��d�*��9[���ؾ�I���e s[���g%Zʼ���({&��*������3]�������O�q~��z(����48>P�'�W�)���H�e
��te�7���. ��� f;�9<ͨ����UX2:�MGye)��Z�C��*��F��[.���Ã'G�Wp�5�WaTil#��t��p�'��+�Ҟ.�0l��Eϛv�����w��!]HelgUD@���TTg��w��?�Q�pn��`FԼ�>%<��ތn�O��oi?g�m�f����&���ꜦP��+6��z�V���hK�+��{Rn�4  �|IzEIK������''��@�&�1��L��
�
�(G���H��ru$J�Z�ƐZ1V@k��I��T���<�w[K?Ɏ����&Q�u�������.|�E��ҕ�1?ݶ��-QK��^+ԢC2@zvg�Rs��&^N���s8���\x��OK��l������a(P;	xY��+�q���a���f��G_�֮��]1�K�m���b�	�4�����ei�2ɐ������g��o����z�m����<
8C=�,�kyNc��n���#+�AV�#�#���7cKR];`�1�ѱ�',� �s"y��6L�=c��B�a���y:nE�V+[A�<�!��k\��2�����\���]�O��i�W��}�����o�y׏]��L����j�b亨��d��Bx%�{���4�I��]�s�O���J4��4̪/�a��{vҽ����V�:�r��v��[X3YT �8X_7P#�K�[w7�����m|^����Q�u�\��$|�Y�9�x��,Zw��/�)�3�si�9L'A�H��<#��LA�Iw���D����n��<qި��$T��W���گ��Q/
MU�V�
f'&Ӆ+j4:,J>Yl�]�+��̸|Z�y!d$S�k�s�n���hgȝ�o�ԣVI5`3��wIO�f��g�r˅�i�S��%�C7�=���?�>e�1�i��闾�|��j��L��T}��(���ön{3�d��C=A�^oᏠ`�mE�F��i~�'c�'5$jF�|%!u��趻r�8��P�� �ئ�b�ul�U�.U9�z��`T)H���X���w����q ���i_���d~doZ�lKc���5�~Z��`" ��(�P��(������)�"c�O�>���y(]bT�B:��,~0N#�=�q"�+�3o�om���iVX�ֻ��R�P&�^j���%�5���r�^ItxfG��5?�j�JA/�MM�:��)�=s��^gX]kOU>Q�4)쓗V�ghM��B��� �R,��O�&��{r=�x�N�5)��1�u�K1�`�B�l�C�hL�5a�ʞ�K
P+�P�qW�;������H  ��l�����A �>�=B�k���d솰�B_�2ӟ�SN��+p{ � �DAG���7,�I�k_e�:�	bM��𝠛��xV��XͯW��{}^���������Z�OѻP���?/Lip�s�/,�M���8H�	�-��Cj� �6�k%��*����(��i_S+Ŧc䱰�>,�yf�8����S�I5���%�@}#��fZ<.��2��,�������<��a��o��ס��ɺ�mؤc���ڐ�W����	�6bl�%5���b��A,g�M}+wŌ��uOL&Hvw�Z�N`熫�7�R�^E7������2(ev0�3V��99�7yF�ޙIϲ�A4��,�#�+#M0��b���8��Å̪�Ӗ-Cf�z����#wB �}(4�,fg���<�����/>t^��Q7�e*;t�&R2�=|�l��=�U)��V�n�O��rB�k�!B��ɦ}���
�ß�Ч��'��'�*�A��;����F�.T+a	�/G��Y��,��^���QdcK-�ͤkܱH�.���#�3~�d+�y�w��Vt�+;2�ҟ�N�>ǡ��!��.-85c������G�f�?�ڳ���6��3�ѕz��.B<{.gl�Qr:β�I��m漌����*5�ɴ�ϔ#MK�£��M�{�C?�I@Ƭ_�ER���!���Bp	A���ۉ�&\qo JQ�E�LS֠���i��1�'�'O���PU��ŞU,���F���7�x ����&��G~� 6���y :�7�S�b�!� �z�,L�{|�<�����σа��A���!TI �v�7���s�Ճ`��}k��2�NZ	�K�����r���U0�NR�v��8�S�r��՘��[��^��1H�8�L	��ڎ>vB�w�`a(������p3Q����򉴄nJ_-J6Ύ��E��Kw�PK��rVEdD��;��ҍ��:��3�P�y8���o�&��v��:V�b�oh7wu��(�17�ܗ��VR�<��fK%���N�]<�3A�0B'¨��x�+��\������≫��rT�	��H�
EM�C)�����E�d���5�ۭԘm��RP�Q*0FS�F�JF"�/��[I(�Zd���Ң�$I�BF"�7�:p}CVA�Q�>�F�O��uD�+��[�ݑn�K�㹶b}c}�+`
��̷��w�{렄"�J�3���\��d�#9n��~��H%��(�8v,�t��u�h�{��J��K��	��@�K	 ���[zv��f�3$'o��Ѻ��	K�M��uARb9�'��J:h��7ج���J���o���9��(zz7��H�r�lS���&cՑ���m��:Ze�����N���JP��5$�`?���%��\�ʽ픒�d޶��?A!?��~YƝ�ۇ�U
y�����~^Zt$jVmmY�f_O�UR��r�G�^���BV�@����Oom߷�a��

C���C���,��d�/��3��e�<W/Io��g3�3<��ׄ��';�X�]��D�a�Ȍfq�<�n*nI�`���$��xW�2C3<�M��qAƽݨ�"�Em"����] j8FN;z���,�$�Y�|X��v�Y���ٺ7�������G5_�c�E�]��;�J�R����
�v�\S��n�2��7̧W|E���s(�e�~�8�!��t�He�p,�н�!8�g{�{d�(' ���nΎ�pݓ��G�Q
MH]���{{;1��~W�mJ���K2�u�"�hƌ9,�wT$�SH�29R$��ܠ'Ӱ������>����(���*����&�Ƚc�Ľ�N��+�
�e���{B���+pnHH��&Ѳ�ԉ�Y�nS�&�����u��@����;E��a���������Y�Z>�j��N3U�XBa��}|�0���r� )�d�
��������q�G+��>V3���:�DC�h�L�T�]ބ,dQ�~3F������A�Hv�6y.N��c��5�a��ׄ��o79��U~���!I�mL��I��~A\�^]�b��J(�x�'Z�<��&�"֎�H;�I���[��S�,��:g&��P���{�N�|9��ee5��h���2c�U'��/x�#��i&���$��4�k�^*�#G��,O{�؊�w�M�6��΅�GN���W��Ӧu�7��dp�:C̖����Z� d�w�E��2Ǒ\B!^.�*C�=j�x����)!�@R�R��U�7�CF�Lv���e)��N�Rj��`5f�ݞq����TĘ��1��ْ_�v�`8*�9��A�!�~ ��:��Μ�J�T�fA�t��2��BKW�ʧ�W;)�kV�VN��Kk�D��E<�IW�?�qj4dXE�
�<5.��3@X��ATQә���SMb՝'#U��P�V/PЋ���)�M画�_��-�^��Ȣ6/��XV�Za�W�ǚ���Y�p�t�0#�D��ݶ��\F��w	���}D���B�U����7��8e�ԷX�WȬϋ�����+C��IQ������A᡻q�e�i�,�lk����@�`u�TYUF�'k"���[W|f�f���K���g	���m�����7�xjC�$�<a�6���<������m�����
������fi4�����v �$>�G�<�p�댅�@U$b�s��;�ү��u<$�{��l2o�5躑a��=��k������ ~��f�N�L9@�7;���S�Ը}J(�����m��؛�F�O<�f ;��+����@�Q8la=��-�����P�~�E;Du���ߍ��33� ���h��S�4���~]Ԃ��fq�0��܏���,.U�b��W��=墆ͳ�ǛK=�SA�T�o���/!��lr��ꞛ��m����V� ː{�f�I��I�Ü����v��f_z����8��g���ī�i3���O��?LP�\�xRo���������'�ϴ����բƔM߯r�Ž�|@v_g{�0�.7���{]��r�n&��q'R�XA
x<�y��Qƌ�7�#����d�+���S�dZ��"PQ��)rMHA9@�ي5�v`(���b�֝=�dr��ST[�0��r?�[32���*�Eܠ���h f�(��9\� #�_�%����s�&(V���L���8@�/P��3�c�����d�(�Kߘ�@�����+ )��U;�b#���t/ jٿ�\���t���@w��S��g�1�]!,�݌���X۪l�\²������w��.��h��@t���)Mn(Fx�=�k���oaK�T:�E�#��H�?���HOe��A:�tԚ,�����T)�x�eD����f�yq;����6�lF �/�c��!��S����������LjE\�0L-!1$!�#-XmA��"Nv'U1� ��~�L�M����G�z���HM�6��[׳Z�(b-B~|Jp���) �ꇞEPf��[��-���;ֽ% u�mH,������l*��?W(X:�g+p�\��E���v?���zOo���|�Xh���t���@�	�4�g����|�4,_���D5(!�i���E�S�M���4��9�>r��H���P:f۹�裧B�>�gߤ()�(ny���IC��,m�G羳�q�xn�r6�t�/}Ӫ86!z���j� |�"��+0��wV�T^m�N�ˡ�����z�uiZ�ĤF�*e��n{3,�TS��H��`|�(�itc�k d���G�f��!��3��IP�Y��d�~����:�"��w�,����[ɂ���΃s..��MkJCj@#��:Q�?b*L�rs+����kx4���2�9��X��s�277č�=>)Ad��xr�c�>���2=RXS�8�;Y�#+�4yi��Ea��N�p�<2���`��HH}F���{��E��K��a��]�G�AZaޅ�W����,�f��ѸI�}۪I~��I�ۧ�HF�ׇ<�/B�]�q$��5��zg���'�xD򻷫t��jPG�IZd�v7[�;��E�O@�o�j������A�Ҥ��83�_�8�&��q�����e^��X�:4�	/�P��
3v ��B'�R��ᮇ4�9ze����4��(��E�b)42hƓ��n�Λ�%�d��@�䒁� �鳭�S����͋��7���o��bj�'�~���	a�Or�An��ӷ�(G(���c�ǊW� ��R����'�h" ��}3�����Joٲ�@�,�F���G'S�|�C��� ������*̡v@$]��L���w�8��TFl���a���3"�L[��i���&Rd*�d�S�<�;i���8,s� ���`y��e�FrX�^OS4�-M�����m������}�?+��d��9$��3ֱd-�p˄1HfЁjӖsE�k����'�o���B�{�����(���c���D��4FYGu����C��O \��:�dK�~�w����Q5�wU_`��)���ry�����H�F�2�N����%pO�t��/2�Nnv�����n�r���!��1N�Y;�i���=5���s��ЗaF�ڞF�}�[�/�j��R��=�o�Z�ĞP�?������%������ڌ��>���%�71Xۣ�[���!.���X��7��0�W���%Q�]W��ѱ�����5�7����R�\�<Aۈ�!�3�IB%�9 ��Q]d���;���_�����*���+���]������R����kr�P��y��ªX?�'9FwG��n���#�KP�sw�C�,��òr�~_Ǟ����� Y���q��J������A#������o^��F�	2���ǽ�\U�����eP0��Vѕ���_�>h�Ns�w��4ӝ�5�Q�c��U�nG}v⪍��h����[���AT��0�0�:YMB�����U�������Z^9�%�N����7#0��r�e���h2�K��^g���N��՗�B�PC�YqtX���>^p��{	�
��П~���gcD�=µ��A֊�_����0�.pz2��W�[si��93�
�ȴ��B_T�g�P���S�ԋ[b��` ��|0�:�&4^i�d��\n`5�}����]*CκWm���!�f�#����Q@m����Ggޭ���ZYz�yxri1�en��y��eu)^�JQecS��a��雧���� 1�����;P n�n�	<�1���qt�4�����u��[�뮼��b8����h�lM�G(����ﯘMՁˠ;�����]�%e���^4-I�K�<��Αv�f2���m!����٧��<������(=[��7�������NE��������L����N����.�@�L=���*h�3�f*,�#�pV<V־�w��ײ���D�ra4��Y^��)z�t�yU�&+�	�A]c���u���L}W�F1��s>W"��q�`��{P�-�k���L5���cPwA�F��Қ�.>ƕ@oiW�|����߅un#��H!d��H�P�C��+��o٪�3�޸E �l���C�<@�m�����w�JO�h3�Ew_�!�*9�/2���䖂�m��1�K��M�эa���j���yF.i�C�P(f�G��:�a�%�Q�4����m���kU���Z�+<myu��r,|>pH�.�b�Z���� �D�v���D����SC�TR%m��z�M�%嬖4�cGp��)_�`Q@>cP���!�<%Tƿ,<��|2k���kz��ԕ�L����5BB"j yU�ґ��Y�h��� �σ��ힸS�D��u�C`��"�ḧ́��^m8����_�9�O�	r �5����yY!Ћ��d��+�G��z�v���A�Pk]�_�Os��j�L�j�:~�c�q'�$�"�S����&^4�{yfh<��pOD�f�sQ*Q��ύ:C��fg�������M*rٶڢTՠ��vX�ǩ���o�n����q�5���#�YۃG�X+ݎ����6�9��O$l���^R���|��2K��B�ֽ7���	��ρmp"_���\�E�i*�+'X�N�32r��7G0&����|�@]� �*����)V� [�GjT�	��,��ч��9����Uq�h$m�[֠y�|��Ȃ��0���Yk�յ��ψ�yfR�_l7`oPPd"5ݴ3e|�D\Щ�FE�׃����ۻ�8�O��A�0�N�u����scy ���o�9��A�г�w��p͉��7L���Oߞ�LU�d�?�|֝��vKb<�̟�l��c���1b����seƑoqz����+!11��$9�c�,�W�[����56-��������г��\h�����J�b�>"[��-�ry>�NϏ�|>���v:T��^�Q�F ���g�F/|�tC6��s 7���K-W����te��I��&�2����P9y̍�rm	%��k�x�P�T���Y��e�A�7�!a:Z�ܡ�Z5:�`#;e�nH#3D�qf�*G��Eqȸ�|u�(���� rp�����V譆�+�<w������r�/f�d���>c�b'��Q5�Ղl��������T�Tk\1G�\��)�0����L~��#��s$t��}d�K6)��w`i_�%̃�ĤJ/'!�3�����@x��/�A���wK1������_ղ��z�xj5��r�:[�PO���	1DE���g�3km�h�`� Sڞ5�lN�������~f^���(�!�Ol�Vb��
r��#x)I�bnЃ�?4Bm}�΢���N,v���Z5�r9��7|���׶9!�*ӆ% �3t}�����6�s��S�������g�R;�Ɩ��+��o�R�~R��ʸ��z�}�P2�{��0�t���I��v�f��I�T-#<�ie\A�:���Ij{�����<�6H��"��{�_���|Y~[-=���>�h����lSp`I��.te��%Ӷy����Ć���ݭ��n������f»f6�Y)�sZc+D@�( �d��<��������RZ6"�I@��x[�l��Ğ�g�oU��QIh@^�w��N�%j��1�Rv�JR�V�&N��L�%��5Ȁ�%�,6�����'e��/Ɣ��ɩ�x�X��T�i|�-K��ÛZ�O�s��C�:���h�
��mޅ�f�%��j��lN���S�A<�����R��͖E��	�8�&Y+Y�?�^岙E�T6���[~�^,�� �dUAYYv-���i��Їj�����)s�	7��.�a�*j�!��W9�̢��a���c�øx�Q-�'��[֤�+E�8��Z�����ʡ�
�l�R�1d���fv-�z� ��V����2}	E��n�%ֹ20Sy�o��fmjye s�ϓ��v=��e@*sr
/���PQ�r���xf�'{�ztrY��;��0#���5�$.��a�I"������g�R8@iUG#m��F�t��'Î���Źh�N=�Yq���_)I�[�ꡌ�tɲ�-B'�K��?(�#�e��!\%�q�]�w}u�K��r1�՟�[H�����@�f����M%1�����8M���7ښ<gm����H�<��xsR*��k��T��O�B��1�֗1��
���z�{�-x��<���I���ue|U^Z�YG2��W����:]��G�휡�fz��O I��w���e(�%��#w�R^��;u���2uI��/�u�������}Q&�B�k�cԊ"[8)����fvde����u�aa�9�i.�iJ0�� ���i�`/�O�{&�_PÃ�M|;̲���zB�����(y�cV�R@9>i�8ؚ8�vȀC�;YC�F?ɀ�+��X�9������5өyA����}��F]Ǖ��p��������e���Nq��x-酇�(F�Ҋ[�m�;d��S��)L�_��Hj��j�
��x�����]"7��-Z�u��p@�.\�b���/-�Q���3���)9�Oir+o�-{.#�+��[�����q�:��*C��Qȕ������붐N�gWa�
n����"f�Y��4X��M�SL��d�����8��]Cӱ���Ojy�Q&$-�$�A2D\IY������5��ט;>]���(3�'�*F�j�='t=p33� z��ͺ��^I�Jc�D�uc]�҄/��Ȭ
r�=B�y*'��K$�)�j�R�[�8�lҘ7.���^;	���X�"���Ѳ{&��\9̥�Q-��=_�8⡾�T���:�m��i#B�u��5�᜔>9�0D>O�L����S\,H�c�@:$�1�G�6�r����+�%%�'�W��=�
���&xb�O���v���?�e}T�E�������i
�'�`Gਇ�+{e�X�3�)��@�9SK�K�["�ɖ*�٘��>����O��{7/b7�bYG̴U7�r~�F`����Ie�)��.�LN��_�,|����7��G�T�V�MZ�5*(���5!�}���Ù�!*��]���wW�|��ǳ�O]��UCЎu/��k���55�y���xNbr1ʭ53u����>�1y�K�Z�ۘ�-B��/Ɨ�&��;OTp������K�
�*��Y�~�IcA�zڇPd��)�!o���4q�Y��E�i2�;��
��������-���c!.f��_yr�!Bb_���[�s���� 'X��Ϩow\Yn�����F��3�j냞�E���C��%�wg������U���_�������e�z���Y��؍-����[-��a:Q삌Ƚ�L�[���#G B��]����.���$�UmlC�ʬj�D���%f�Q�1��₂X>Mp�����de�*���ƿUڇ���gY�0C�=�+�-Q�J���F�Kh�2��\~s�Ŋ 6(��{cLI�\{X�9����_J�"�i��	�f�>��B\��S h�J�V������c���מ��t?�l�MXI\٩�(L��o���+����(�}�Ǭ7I�+L�R���2�"���/�FQ�M#:u6�^�5~WU*�Or��Wj�i&�X9Ș�!Q�ҞB5�_���Z˥�ь���F�S��rOD�x����y�Q��5�����W?ۙ�%�γ�z0!��օ��uP�Q��t�l� ɩ�0;��Q�}�$;��r�*�ޔ&�~ʎj�������lo$�T8K�0��~e��&1���d���4��S���OXu����u�^��q�#�'��(��:q^׀�aF���Q=��9�$q0��Um�n����Q�S�t�������ܬcмZ�c���]5xc?"3]�N�� �=��
�BP�3��k�;BVPc�7�b��V�A�;Áy" ��v��3|yb9K,nm4��X�����g�p�6*}X�������C`4�'bj:_S$ҧ:��{A�[����UpF��?�܅  �	�&�h� ��=e �����HJ~�����FA]��F鵭D�A�:(W��>����<9�L�y������c������e�� ��U�s�&µ[��D)f��a�ԇ�Y��b]Z�Wq0�3%�lgw�Y(����zX��͑±��] ��,���U�'��bh��Ք�73OϾ�,���<���t��:��T˽R��������K�D|���|R���Z�-���]�0t,�O����S0����o��U�}̵W�	��Gd$����V>6B��Vq��Z�����T+(�����w���y�������;[�����A��-��He ��Kԛ~��;���K�] d\R��֩崛C�=��k�a8a�� %Iqpp�){��M�@.���w&!R
�"d�nN�8o��O.K���޽9 0����v�ߛI��?�XI�QB����B$xqq�`"�D��$��l�rUz$<��rv��dVk;�UPI��{2c{��e��n�iR�6kgG:"/PrJ>��$b�n���S�����L���;��	����׽�� ��NU��1;�=�1� I7JDԱ22^� � �Z�"��!@%|���J<��sB�Ml�7LX� A
 92+��x���vN��hS�l �T����V�$��R$�"���t��m%�kb9�X�t��?¼���k�ؤc)��xmͫ��w��>d��JW��މ�G� /&� �m����ϫqm���kg&�t���H�a��/j�S�\(͝T�	�j��tY����r%�@6兩��X��6�t�O��/�Ue��,��&�W�[g�(}�|�t����[���u2Y�^S��u�j>�m��/۰*�l"S9`
f�'�V%W���w����a�g�24�[����p@�M�1x�/5zw��@4���E��D&�P��m�n��������ȋ$��}���4WM�d�.b�#3����͡>|��>�	A����t�%4�V��M��ӎ6ç��UZ�:�b��$)�̱�\�o@����&+�
mj�=���m@s l֖���+�椴�o�{��Px�^��Q��u�9�a�-J:jm���&�l׉�-m����գ�K�N�dh)G�,��=Ob����'4v�,��9�W4؝D��3�$�ɢF��I"M��z�P?r0��C�0�V�S����3�/��(�ʐ�4���s��rZ9��?�,6bt�vEK2aaT��U��Zv��!�8U�Aj̉����\��+�_tS*�\_�mF�{��д�b���/��`�'u��lSMם�k�ٟmG��c�����aª�q��MW��% ��׬qɼ$�Y��j��_P�I/99ke�c?����n
0��c*�9x�8�{� ��4���U)�F��f!�i/a�Wk�z'���^��EZ��]��)����c�e���S�/ɉy�w����&��O�{���8��Nf�󵧌E�]��p���UX1�[�� �f&J�2�c%-)p�9��d ���bs�=b ��O�EC1�y~������'����"`;����Z? ��@�ϏZ^��ۗ�̴tF��rC��oS%�Q�c"�l�+�L��Է�P���7��kDD�2���a �3:�1C��NO5���x�[�{Aw�~�)8_;Nj�#�n�t�H Wkݗ��c���H���I������ܤQ-8�6��D��L4?+���7_�ɇ�şi��&�1��o� �P'7��w�������Ѷ���@�z;JfQ˲N�,��, ��BD�P��Ư�'d��ȿ��ٴ\#--��]��v��b�XaCEE�����d�R9�i���$�&Tgڟ�����]7W�,��t�P��'0�V�{�v�Fj��Ň��Á�90��22��k5LB_�ƀ]��/g]���-j�D��#5�=m�h�c��R��>ˎ�hC��Y)t�w�UwI��)K��x]Tm-*�	�T��YC� �\�	�$�5�)8��h�n��{P��� �1V9
��f��÷C��8Lx���a����J�a�4Z��%������ܔ\HFP���Aʿ+�%9{u��.(�ȪQ���^ˤyy�z��ph�J`�̤j��EQU���%��Y/n�t��ȣ�/;��L��H���S�4�?L#S�=b����=K������!M[�j��3��:h!my���p�/�QmJ8�X�s����'�(	�F��6�1��Sq<z��O����Gr$�ks�0�2�mR��4��q���-�Ml ~ ơr��0 B��g��r	CA��x�6�{��v��K���XZys,%��b���9P�[{��/�z��cR?Ѻ�\�{r[���}�k��x�O�j��!R%<$4l8C��r��� �d;~�l�+�{l�zE�0�����e@�*&��yq'�e��1O��Νq�7��ߡ�| )<Mgb��C��?7޴��OO�SO9� �mq�X�.Y��+�S�X�j��
=�D��d^^kD�hlsm7��:��?-���`(�E���b�1�����>V>� ���\6�e��\K�SķB��-�<{9�����L���Z�N*��,��eh)�L]%3�@�Nd�Pe�<�Dߋ����f�j��^/�^*�p��*���n*S9�:�C'M�|O��f�3�U�jKw�P�acIAP�m>��ėc�O007�RNĻ�����%O���td��:�z�ޛM$'��O�Z��$^vL�K&'-U���$�C�^���K��h!�~2�4&�N|�̖*�qG�>?�7Aŷ�k��	+w}2ȗ����I��#������W�&SՖN���4�� �y��1)��%�J�8!� j��؏�(&8�P����.H͛q��V���Zm*�k�l�p��ژ������)Q&��8�q����T�J��zK��&:�N� #�|���F/^�~�҄J��
S���:C<.~� �]Jr��3	q��. ��Dߊ��8�ht�s����n? J)#�`��5׮�}�!�����39'�7h���#��&"��JJ��n"�'�@��b��[��5��'x��j$����-�MK-��&�Z�"
�A-�S���ʘ�G�D�|`a�br���ݬe�_�ܶy6_Њ7��A5��vƄ}�5�[��\�#5
�P�McB����:�Us��V�v9��Z�!$|~�p���}v#�BE\Dë����'�#����� &h��ó����M@��%�]�a�d��:��N���¦�w=���m�1
�R����Ŝ6�o��s�B6����]��D��w��G�=��N'��G�Å��`�uٜ ��t���'�y?�B����!�܉0�٢���i��<WeR�T������b���ɇ.N�G��%P�i��?�j��Ε����/�$�0
Ԃ^9��O��C�� ZT�5![�3�XAF����I�13B�w����!m�͎6� Vy7(a���Ӥ�+�]�l�u�H�\q�2��	�Q�+��;!`r�(8(�B<m��O��&eI�v�z�q<5�a�O�l7[�q�6����7��C��(�f��7r^��B���6�	������m����X �f�n�Pb�ˤ6w�`7�,5�Z�{;��ұ'�گ&v6�ڂ�W�u�ub��8t%l/���$ERAք�z�!a�n�Ź�/������Z�Y���1��8��Z!gӖ��<X=�a:Mg�� �T���tk��6SbL���D虜
����/"�o�����)�����~=2���m����B1�4u4 7O5Y�$�"Ct]�`{M��'DZķ�# %��~��`����?���@�><2{"O���W�|5���g��-@�-#�W
q��~�'��bX����S��,j�#rͦ��H����G-��eyB�xd^��ҙ��7�8���ʑ$�1��>���ꋲ��s''Q�7�ȩ���95+�9��6�ǔ����lM�f�Im����-[��ifٱb�0f|.�z'Q�L��_�QX'ֳ�D�� ��O���;�G���++YiН��oX�F��aӁ���&��xPH&����X�y^��9���􊰙r\�59�?2���㆝z{��Ė|���x*����s���kr�F�i�0t��8�/,� Hh�×l,�?�,��k�iu����1#�8�~u���k�իm�CE|�g~H�s�f��Ћ�8&�ktQX[F�=24��"V}j�2���f-�C����,m����p���U,��t,�=�׿s��`б�W�RN�eE��{"��L� �h�H��蕩����򑜲/{��tzQl!'p��z��<d"�3֖��uʾ�Z��r7G�C��x�d!  �����]? ?a�q�3CtpW_����bbb7�xc֪�Kd�����a�'�����X����K����9u|���Ў�I�Wl��4Đ�ۄ2�D��U�zQ�A�J#kwj����T��R����"[c�GDiZ��Pzșt+/�I�U�I$t�Vw���'�i������S�V%y6�m�pH��se]^�kr�J�M��A,k竝�ni��v��B�YihI�� ��g��'�|paA��~�]����@���"��7
[T��)q����t��k�-$��|$�"���0�g��3�QQH�7��9FO&�$��wTڊ]�\P�3]m����;�
�R;/��|F��$�!��JJp��Ԉ���,���B�\������l@�dfQ�t�z����F��C�hB�@��{�j����8~����K���+X�a�â�'W�
4�@>L�6h4n]"7���y��w��ʫ�����4�bu��ZũuՌE�E:ʽ�ɦ�4��x��G+��yĠ���i�3��:�3U6��H�����[�W����N�֨2 Ek[5�]P����^=@�r��̣�H�X(dT؞g�M>��?n$.7�+����ȝ��~ʡ���<������W���|2�eP���L����i��z6St���]F�,��r�Iʎ�!��/U�1��|h*���"�e�����q���x��//[{74W�UF=���2"��~ܬz���R��w�zzd����iv<���S���7��W����ŲX8$��<�j�@we�eܻ�EZ���-�'�"�lZ�I������}-,���eł����1�vݻ�?(��Tw׬�h��e&r_�Z���S|��9�o�'���GQH�2��'\\x�0N&��?ܤ�;!�?r
������z8i�����ø� ����n=W-�y័&u�6���+����z �C����p��W%a�{b�1>�v �K׳^��<ބ�9|[�F���q�����J���_������9vO�\O5:�s5�l?�Pb�P22�!W��l�ܣ�r�4{�<����x���)����Z�ݮ_c�e���|�K�U��aqtN�h!�s�'QZИiF�{�5�;���m2
1ǫ�ǎW,��_N�_���)�p!�vUM^���eφn���5dW�-č=����Iֻ<�u����T6o��<�o�T!�F�%U����=�"��[٢����O���rӂ#�@P7W���\JB���4�.�Ȝ�V-ӣ�	]���#�"��a�K!D	Q{�p
�=����AԣY�`��A��5y�q���v�Sb�L�����fV�����L���x~�5UU��$C�V:�.�f
iQ�j�煟��P��0�[[�@x�]���E���\�yU�4�L�`�]
/�|tM��m{����g��P�����o��p՛*�dw@Wu�p�����i��w�4^u'4yZ+�+-�vwt�gW��Bg7g�{�-G�۫��#�H�\��;��2H,��U���z��Zc�G׎o$�$������>L�z�
��G�	�J^cBJ��V����xu���`	��dd�}KG@���[ KI�p�u��^�(�;�>��Ug5m�ĺ�
}���3�+Ig����OUO�&8.� T�U�z"��������ãJ,.�?t=��A}�ō���Zm��u��m8V���T����U���:����Q]6E�/K{�R��@��PD�j�N��|�t��a+�#��G�-���34��������|;�o=+$��I��4�	��D����7��9���g�띔&T��B�4���i	0.BC���N`��P/p�19H��~�מ�ʝ�V�u��Wn���Q����~�σn�����ޱ0,����t�t2�u�(�����dQ �V���W��2e֛� �{YI�����9

��AoLX!���tf�v~+ ػ�R�~̴�g��Yf1#d����o�U�:xݖ,6��{��0�:���|sW:�O\]ѧ�li�c�������5y�y���7J@�d�������L��Ve�}�֍�'x���(��
B�fm��0v@��r�[������_����vd��ƅ�� ɴ�X=[�ʀ��Uj��!���m���i#{��&��^��½8UW�#^����C�r7`�F�D�����-��Sl|�^u�;]E����!L�w�-����&���GB���WN�,��{z�
����B�JC�ʟ����^����ޒ*�~h�9�Y&��Zҹp�O���ĔB��$➿�a�@~����9"�<�??<�md�V `׫�ފ����H}p�k���Uh���%�G�\̣u�ܧvF<�E�2�J�:�صq&��|��p�|�V���G/� �>�ϵ���HC�B��c�4Æ��5'�����Oe�r�}�pm"�x��l������ȟӅ	��ޮ�,9�l�����.��}����0�M`�-��jf2�d����P_7�
�R�����ܲ?F��d�k�L�:��v��ޢ	�������	��]�G$��B�Z7� K2����]ܢ�!+�˛��^�ƃ���&�ij�Ad��H�F��Hs�PN��ׄoџ�.�g��#~C��O����"/�=�u�J�Ge�^�$��W��,+����U��H�ތ��뮮m����O����5�qC��"�'Pt�ܹ�� �*'��B�+�\�o�^4��N���ȡ��$�4�&��[�Z|2����ޅItFm.B���J��b{�'+�X��Wh��{~��9����\	H��3E1��!}��<ɽGd��mcCs��E��D/�"6�)�LϘ�I�R`!�U�jаv9�҃�ՙ��Չ߃�c{���-ۭe>TfX��e�T�%�����<���C48�� T���=2U9��W�eHfh�O�2�F�U�|
�d��Ƈ�NJ/�kL�H2�Ԝ�����/���z<��#�8�lf�;����u���#�Ňþ����δ���n��"20��@�ҪC���I�84�!���荛�&�l�>�1��]��a�e�mz_���N�[+����$��v5�_��Ob���v��/�k�N�P�'No�=���u�8e+y�r�7:�;��A���F�.�vN��xC]�o�@��X�\bի�Cq��NftdpB�-���o�����TT�u�)�Ѿ�W�R�=gٳ�'�C+�}x{2Z��dS�fP�-�dح��E���u�@%�@�p��6]/�6s�f?�k���n���y��x��� �я� ��ڶ�ī��3��4��OƝ���΁ϒ��t�,����MMD�O�IL�8�i/$<��Ly�w�u������`�*?0
m�*f����o�1�d�3�Yz�{�btH�kҬeh0J��V��_fؙ|�q�#���^�Dc��D�N�\���,i��{1��(6u"h�MN�1�ZiCzݐ��9�8uz��W�pۭ�-1��
�� &�	�ڸ�1�7]K��6�ƛ��#������4�����p��V�'�-`~�E�aS@�KtYC����0��z�%�ך=E@ ��F'(�V�Mqə���?����A�oy	��O��N�[(g�-�U�����~�a6��4I``��Z��0��p������D5+���$M���/Q"ޟc
�X��Gq�ƿeJ��A�L����,���_:몍��-�k+��E#=��7�*���2�lH�£ty5����oC�/+��E;'�dzge������h:���� �ጔ�HT��r��Ù�%8�����!���k�؄n���gFOf��ƶ�r�k����0+@�|Ҡߗ|��5![2��tP��ǣE"(_�M�i������籥�z"{_;�*������F%؇H�ar	ڟ&���e�
fu.ЀH)�b�Z�#}�|F���	��W�L�K�I-hW@�b��to���ܖ]�S'u�!	^��ö��0-��5L{�cD�ȌI��I+}a�~���sUf����P��!�̲e�D\"iI�-�=~3p���Z�c>�VbSc��|��e;CY�;����}V�G��"�Y ��nr��Q�?>�f3vX�S�M�Bu���}m�k��U��7C/K9#O�����Q�ec�*��(kv:��tO�#����"�J��~f�����A�/�%cm���_8�����N��g����J� �"�gQ�����Juf�\�K��,?����K�+Y�K����h.��a����5�,v%I��b \3(X�7n�1)�Hֈ!�>�k��V�1�T»D9��5;{�¤[�$�t������d�!&.H�;���G�v6����8����sA�
���` 4ބ�sdю�Ԍك�س\�S�s*d?��yqf�T�>�Ҙr2p� �M�9�W��0~[��˪���{�e��H`a��t�.Tpv��RWszA��	Nf@o��s%R؋/�����B��~9���q��Y�v@=�7��8��Lĥ	�*�쇹�Q�LR���AJ��-� ��D�m,Y�.s[�9̘���r9O\�b|��Ej4��As��g�G{6������#�/�$�q�0ſ���6oT>�n�H{��.��C��6 F|���=�"�a�Ԫ|�j/ad�e�V��	Y�ݻ)k�Rs@��E�sr#�Ó_7�)n��[|��,�R"�1W_�������Dl��Bt~��Th��C�,>�^����Sm���:$ɫ�a�χ�8e(h�i��$��
��
��9x\ �L� �
�݁L{�_wc> ��vΥd�U}[�09������
69�4å�|�/�#��P���N���Q�~ת
�Ɣ�!�-��L�����`�nt�r�m�x��;F����`���!ڤfw��~(�(XB'�O����҆�Tu��j�����yr�����Z�gԶcb�15�1v��+�"l���@�O�⚲�Yڃ#]�2�%��& �1ZD���F��^�	�;���7� ' �d�jg��2��A�>ZM���,|�B�$����r����-�
*��D�aa;cc��qg
G'=�4�͋]ĮH]pq�vf��ǐ�e_o�U��\-���Md��Ԥ�E���/�Q�	���=���3�q���$ǺFs�`�o,��ѻ�e�(��G^��f���|�X�+!f�S�b�=�������$��	���P��%��;�T�{�����ZS��ћ|�J"F����� ;U�����b^1�j�WXKڡ�π�6mZ�I+����2����6��h.�S�����bG��n�+H^ml�58��x���~��6r�F�g�#��������v�B�Ξ�/�E%��`��1J��"�0%ɼP\p+���|�͵^�"5��K�ޚ�Y��H>�+��~]�<���,�:�Xǽ���(��-�ܽ(��G�/�ѻM����1c-+ߚJ/�d�q�"ⲍ#�����~bcbfi`�:�ڼP�',��B֝jQ�����N�:O��ef�x��&(�#(p�U��XZx�6�Y�	6��a��m������9olbϻH��L���(+\���*�D��A�>4��$���7�s�ajx�H ��@��c���!����[V��\�"���b�4K}�����82��Q��۠��=ޥ�8
6r>�N�7(l,d��M�G#���d�&��H?�� Z\Sy�����<-����mh�a����� �>a���%���ߒ����To��H�����(.�G�ß0K�ch�;��o�_���X~ڂ�g�(����d�2���$�x=��0q��b����RD�#�M�|�h8>��W��ˬB�Ѵ�N����M�tl��>���4�-��`��&E�i�&jY���Hq��	�;^8����ϽQ��a��M�`������=�e�Ț�vآ��9bU�ʼ��G���Z�#�ic}�����ࣳ�|��w����.ͳ��胠�����F �`_"�x��08�xc�5~Qq���T��U����h�m9�عV�N8�9d]g��AF���C����8���+�}�%e"�%�n�C'������'Y^<�R:���C��W?�p�<����qz�,�l�WȖ%��k�c���nyJx(����o�����{,I���p*��?�-��C�P�R�$n�w��V6��C��U� ����%��Ή�jz��27M��M�oh�8l�؎�ӌ�DS���/zx�csx�M�B|-xHˀ_L闟�5i�)Ծ��$͆�z�,��u�SN��Ib���st�ļYo2�x�5d�;:�m~�N}�\��sim��=x"��?9�XS������dP��0��BO���6k:���Q'�Ċ��{��5;��i�ٌ3���8g����8��%�Q�&B���qR�����U�(`���A�װϺ�L� ��'zRŽ%B���=�� �R%DBC�y-�ĕ}Y����Tq��!�e*�ߨ�x�R�B$Txу80»�ewY$�i��N�	3L��6b	����E+��,�`�������&  �:��歅zæ�3B?��q6��>����I~K��`�Q*0��	LAl�z��y!v�c[E].b؝M�ꬄeA���i��ڹu)Pn�fM[���d�U|�h����[�{>����H^��xxә��w饪����7.y �d\������ڞ�	����)*d�j[������1<Y��tDݴ�>���^ς�'��^� (!����	Ч��tp����[R�ؠF�;��!�*T�%֘���+	��rQ�D_UE�z^��zy�,d?}���UvvF�D����=�I��^k��A�:�ۂyz�<�r�*�����0Z��)����)_�ǆ� 
���&I��}	�@����]u�%s�Q�������vP�0"<k������`;Vn�&'�������fM9ڬu�~��v>�V��j��]�f�̫YE�a}�=�pWwi5��k%D��T8��=���(*���j"��ܿɕ�&�r�i: ���;��qG�%VJx�h�UW�W`������nt�i����&�����`��>-+xд!��!1Tc���jY���s�j�����v�.0�Pu��p�����'��ZEN�G�c��u��>fdNB.�m�ʭ�����ce&��S^����LֺP�����r��8�]˸�n{0�hD���lq_g9龥��Ж0�DGY�U�>9o�5��E$
I����)��5r�I���J��`P�_(�7B���v�I���k!�S��bE�7Ĭ��A��y�q�{��so�?����6�N��Ⱦ��!���-� ��G�I�Lg�y�v�q�$ޘ���V���9&����#���~iО�b5?�N,a̶um$����w�,W�}����"E~��Z���a���V�~�aǑi���vf��A3�P�QێF���삍KV(�~J��8NT��*T����9sj�k�nC:V�ǋm�B�*�f��6sH�ij��5�V��5wg�~a�q᮵hҥ�n�v�7G� 4E � �
	#�����X>t�ħ'4RX($��H��䍂!l"���@��g��r�ͺ�ż�eY�m@����-�	opC�猬�пX��a|E�JMV˫>R�҅��l�(é����~�I6	�5�Ֆ4l�Y����d?�h�=Ὗ�'?�l���5�����g��s�a�\tǇx�����f�e�xb
�,��p�~��b�eTy�F��*����u�>��?�wzw�pR�c��OQ#�|���!�Fl��3��'�5R�@�=��-�
����E�<Uo"�'i���77��e`�3�P,/�8�x0ٸ���=��^BQa2�{�.EC����#��p oC�J�o8;�J=�< YB��,R��(/�R�u��@`|(H�L�p����WS�p Z��='�8��-��?N����1����F}ꋱ�͊Ǳ�"�$�j2�#!��)��� 4ܩ�TO�W���w��c���Ym�euLy�,&����&�����N���r5�Kڝ��,�b���T[",m����BҤX��??���EA\�X]�ʮ` 3�?�P}W�=b�5hvO��yJ�=�SNOR/̋>K�%i:�A�x��ck]$�o�}og�5�\�Q��'zX*flȭ�V��8;�˱bCs��M�{)o֮\^��`P��<���@���K���0�E<��~��wZ3���&��я�%C�wḯjr��������q�T��ߞ�\�_E&P^5��ފ<��h����9�V~�����b���C��ۤ�����Gs?���U1`�|�A{j�jgyz�@�(�[��b��ƴ"�:��u6�dq!*���B���T���D��en�n�aS�+��F\qԴ��a�f��Z�s~5_�2�MQXH&͒��C�)9�:~��B���vk#�V��Dl��Qu��Ԉ��Ժ�k�S�f�l�3Lre&l=�Y`�h�W#w_����35F&v��p&�>��P%w�����,}�:U�-�pAo��7�Z�y8�-�ݙnl�%1t�"�X���rG#h/�j���K�����5��3�_|���m
�����]!v�h���E�$��0�'mP��>vTQ�
j΂:]<$�B��v���G�uE�|��!Q
D@�F��I�&��i� ww9mV�.�x�ώ�]o����;����l��(�/��-�Fx����M�u@�"$b޽���%�w[v>�QG�V�F���q
��s�EEK���Z�u\���;!�Vn�3lp�aV�S�b����z�xe�L��P�Mb��A���0~���j��|#�WH���$����7����Dz2�߿��M��T;/��\�ز=%��t(R�p���&8�4�����s�EWﯺ���N˩�z���]�Z_�ŀ�rs��uM!�\>��孮�̢;!�*^,���Qqr��|�J$��p7¤���҃D�¢�0���(#vQ�j����,ts8��k�pdh�#? p����������$��xu��I+�Wa~N�<���=s��b>��Q����cJv���D1��$�����~���jS�T?�>����j�KΧzH�OI�w㆝r�ES�u~��u{� �HaE�r��#Q�i�w�x�n}���
�a�xɯ��o(��o!Xy�C-�w�r��zz�hȶ��B  7����7�L!�Q3jpC'�_4�\�5uP�|�valT<!�K����s�`{� �M�Zm,�A�a(�2��i�bt��@hjc�% � � q��ݾ����m%3��5T�8��D�����a���-��S�K��Ju�m�8��d{�vDA<�R��[V/�6?�y��9yT𝬉&�	�h1��=�	���0�Uhe	ͬ۲%�o��.���5�[��6P�os��fy)�A��vz�4:PMHuPk��b��r�"1M��/ӶU��v���9�}7������e�F>���{�*��2�y�;h�<r�Y\�9�z�}��;�)�N���K����1�����F[4NN��^C���Bq����7f��nu��-�����θo��T�)s�h�_���N�S�͆)Gҳj	�*yO��Q\^_'C���S�-ƴ���A4��̍������]��?�*�����;���A�c��ُj�;S�8�W�7ܭ�?�+�Z�[�Z!����QV����{ �� ��q��L_eE!��Wv��k�x�����Y��R
�^
ZC��w��ꊚ�RJ�=��	|�&R�/B1,s�|��`uc*��f�M�Û0���+E��1�v	�FmY�D���
����8�#�XJOE��Bw��OX��L��K�E�������<����q̐W��>��sa��
������I��_�1Ye�DN��]�u��cra�����Z�H�@H�R�H1����W̲�����	���'#kV4ZWDwm$Z�g�q�}>'�D������r.�yF�Dkx�5�W
��ybsy־T���� S+�J�hD�ZE��l[�]�_�C+.���%� �i��t��%��P�e�j���g��;�H4�o�*�{b�i�@�Et
��CM�:%K	!����S�?��/4���PK7-��9B1��y0���R��
@��+�c��!�����F�% ���=J���ǃ��qfq���g�_쎀�4a<д������w(l9jYHE��v���V��}��M���%�:_�oӖ[/D��ad��Ulh�Nl1գ1�7�$�U&4t=}͔��⦘~�/ύ�.5I��/Os;�+��<3XF�&�d�����<�H�4a���^��16y�07I�ф��+M�R=�<;?%��Lq���䙃�:���xũad"�ٱK�Z(v���?�^��M5��T:�h���&0�I�[�[��@		�i4î	]}N�	3D.�F�����,�����#	m;N"ܠ�p��(z����5����j������{9Zu��U#d��:���޻�4���[x�J��-��|�jJÂ*����ܰ�u��Z�n��5���8�#�>}�h=py�1�S�qK�H��q��������'fG�"��|e�I��%��UB�� Ϗ�8L3�Ŗ]����I��MQ՞��Ks.�x�æ��l�-]x��k��~؞���/?|�Ni'=�	7�B�m9�a������]h�b2�q��z�C 'P������
(��$H�ܬX9�/������m�9�<��xW�p�jr����Orj]@A��g��=�{	��R_J8�
Ƥ�Fy��*1���8祺hh�:�5dFЇ�qU�Cd��8e���F�����ilO�J�r�E]���K,b&�������b�e�7�H�G6t���Em'$�om��!�>VGIz}�ϱ�i?��kG"Lu;�0=;F8��� v�C_pf��f��e�����C��P�Ɉa��0��#P� 4X�`y
��= ����q&��������.Ϗ���mբ�B��j���Mw�����C-n�F�5�0��--�)�����~Y���!P��*|��o�80�i�(��Pmrpq/
��5�)1 JB8W�3�� ���IJ*lNv}�����
}��7ECcܐ��E��Wv��K�s�x��P̶PX_�*dv�9�$�?�S5Q��(�?p���30��kR��X��>ҥ�KR���^�yb(�݉�㏵�+�o�4R������G(n��>"pt��r��L�Xu�ܬ�ߥ��Te�"�0BI��<��U����9g1uτ^�=cZ�MD�|"�ZL/���Z�W�кLK��<�y-]���`F����S�-p�ԑ��7lQ��� �wg�8�]��ͨ��J�Um�,*���Ow�>1п�1�V�_:R�7u��H	���/ ��$��X��j)ڃ����2��El�yT
`eƲO��A�R�ݨ�g;NQG�C~�"ö_�"��!$ �-�#���w$��W�FD��mSI�s,�<��U_�`¯>Qv�4p�z0�q�&M�p��'��9���y����j�w��o�]�Q�"�C�-nc��j5ŀ���n|ș��}��3ks���sD����))'��rµ�4�i�BE~c���7�l����i\���}��^*�f���7i��.8������kу�JT����k	hΓ�C�I#/�Z�7��&��͉W�1LXGj�ݮ�<�Z�pb�u�p����\&C#��><O��2.l� k뻫�Ƌw��@)���.��K_&�*Ƌ�܉�-���Iv�AW�t����}�xWݓ�gQB�Ȣ�V�h}�"�0V��93��䇦I*�ԝ>ͅ��3��'���cC�`�n�b�΅��yd���BKY`8�2蕒{�}���џ�r����i�	
��M��u~�s��/w1i��Cmr+�g� ������%"%J����6I�� vV�).Q���p���9D�+އE� ^�#X����8�cH�O��k�[W�ŮH�1����I�<��#�Y9ě�Aep�T�B�����8-��\�҂�"���I!�О�L4�~���q2���D���Ԃ�/\���jP�SRC�ƻA=Z���ԫF�Ѣ����K��z7��R�4KN�G�X�|�OXQ�7%;�볛�(����V�i�5�Om�((ky��������L���8GҘ��T��#����_�����O�=�a��q31�%3�D��|��4�:���M��;�bJ>��EZ���B�ewY�q^&{W`��c��vo' !v՗�����j���(D;熷`P��yd��C�U��W��� [1�bZ��|O+����H��q(�Z([�E��{s�g�hiaF���1�����L�r��Z�|�
�:$o_�B;�@�8���ǯ������[kU�f�P	H�7����h�oĜ��{FC�n[���O������s�U�.-"���8`���T����U��~밬5��D�ߥt�^X�b�l���蔂�Y[�7�]���<u�[���P�nR^ܣi�x)�j�!�?��C_��fYGH��G8�����I��H��so�����y.��ZP3�Z�[��ӛo�<x�%\�H(M�H����M���B��r�Q��'�V9���.��8��b��a	c�Bd,�C*��^--
��[oȁGۡ٬=S���Z�BP���gƸ�-�á���fy���wp��#KJ,�HC�:�2�@�CK�Itj��^�6���5ih�B��*�t���J}�߀��@E�B�fU=�y nnz��G@�d&�@-�W�)�����Y؃��ؿ��	�a������+�h�%��?����X;Z$� �g7�{xL+q��O�LFD1���m�hh��#Q������Y^b���ЍY�M��a��B�V��x�O��5[����"����1t0��Ӷ��.gp5/P5��ֈN�^c�_��l׉R�х4����	���܌ʝUUg@!�� �s��΂�����rõ,/�iq��:"���k� N)'"n����h{DA�Q��8e� 5��Ó˛w5�\��^o�g����O���hf7Z�{�V� y!���ۗ���C87��ݼ�Я94�u��O�MГ��5>F(e*[�A�_Y�;N
����S�U��w��0o��H�c�;oLV���S���U���L�W����8Z����gt�O�C�]�:�
Ħ/~�iq�ZE��'"��|g�UL[�jN�����/,Xq%?\ˌ[ׅ*;^�%ZZ�YR�ܝ]-�^0���牻faxsY�G�����A�����=u�%�f�ȡ���? �y��Fl��̓��#�|�lɠ��bcʱ�b�Ư����D���e��|ZI,5�'8��'N ���"�`:����I&ù_��4�׹��$��s�[��H1.�Yк��(y�Mۗ^`�(��9@�UN����~��.i{o���Z3ͳ��56��d�A������&x�
�z�At���M�BJd��C7� �c����~�B��3�ZH���ϫ�*tA�5[�UO��v����5j�zr�?����9Z���Fۅ��"H6Jd��ب�rR`�7�wԻ]C��6��d	*\�Ұ�mG
ו@G�X������k����k���r�շ��GO�\�����:�7[08 ��������� ��"�B&|8�N�{��&��:n�7Nv���.LvkǸ�bz� v~�~��������U��1r-y��=ױ�Y�&�K�}��h6S�?݊k���%��ւ�B���1�VȰ�c���}�'/G�r��v!��Q0����ľ(ur/�#��\��qŦwq�$�!p��x(<3b�m�݅�-���վ6m�H�mB�cFl�L�y7K���ڒ��K%�pר��E����U���_��OLڡSf ��K�=�	�R(�-ǽ����z�"a����:v�?l�-o�1�5��*m��hW%��S��=���G���x�Ͽ�Ӱ���ƽ	���n{菉�L!R��Y`'��)_�4�Nv]�9��88+���Z7���Eb������Jhx���K�;6���,ډד_�$[�.8�]�pB�3�^��U���`'�i缪�БU|a�}3{Y������_!ge�Y����$��{'�j
�a������=�C��+�fX���������� 
�U�f�\�s���fj��:��p�YW5� zZl�3ɏ�[���D#�c�-����}���kXT���9�O��R��dPjR!��!��}@�U�C��ʺ��J�[/� �?�}��_��v!�%�������� ������8�^(ً��0�QI]�Wp�,����O��_����L�4�Dib�W2C6LI�S�7a{�~*x4�d��\yi���L}�E�֭�K#(^�P�>�V�����39�%O�y.o_�/��I�Z9T�GM���$�Z��'��k0m���
z|�v*����w�Z�_�\��ў��βn�����g/w�2���vSմ�Vh��%q��I臖�9+ ��Y�j����ۯ����U9�6�	T�U���V_[ve?�w:���'��+T��hQ@��k�����,L����4�O�f�w�uY9��R����[��Ϳ��ߑ�"�^��4�~��1_�[l���ԡ�O�=�2=']r��I}��W*q7��b+�A�(��ͻ�{��g��V�\Ȣ���͕�k�k�O�F���3�W7���nVB�+m���!#�,���>��9=�Ζٹ#�a�����Nז�(>��Cq��B-��^'i��B���ل�`V҃3���:�?:���ܮ����w�p����9p&�� O���j�.ǘ���Q�n����������+�(<�}��G�3-��=�w\�O�x.��<!\pe����Z��Kx�"(��p��;P��߯������Uv�i�+s?G{1�Y���q��3�j��_��&x��>�H�0zdN*��?��w�AD!8KxK�� 짙��*)�:��H�؁ku'ÎW�>�T]V�7�`R�vOˈs@�ᰯ>P�w��Ӊt�������n[��b�cH��іoz��\Ϝ}_�Y�i���*"F���RIP��ϕɮ��+�1���A�6��/�҅Wn��h�t9Q@����4���zE(�^r/��?�gJ�fpHs�@}����t�`�#��jh�PN��bdYZ�1��N�J��Jt�I~_�_�H�X�Ԯ��Mrud�a��>?����1[��DjO��ۘ����=�[c%z&�U�D,�͠x���2�YW�୥^c���C���_�.��q��r�/��
O���CGzI��Y@C�̢�]4�Hk�Q,����d�]��3���VU���6^n�:9���^���2ܴ�d1s�)�7P�r����qң�>?�hW�y�(sF�9m�5��f�kLHe��dS2�ɴ.���~	��k��b�fd�5�F���N�<��p����T\�����f�T�p�/����zY���P�O�]�%~/S9~�(EXI xE�o��+�5���b(���Hz��8L��ҭpD�tM4���<Ʌp/�ƿ ��[o�ѓ���C���P|N��U?Uds;*A�)Quꉝ�=�=u�l��S���
ˇh��|q���E�^bH;['��Tjq$��亼o��7�hמ��jN�+�D��H�����Ic˾�5�m����Q�UN���yǉc��qn?9��`�����ë��y�7u9���d�N��I0���m����U�;NH�e�1i:�Q��U֚lv-Pn?�>���CC��.I�țX�n߲�MEce��c�ݑ�X��s�1+Hy����#i���:�T2��!��O���s�4�7�JJJ <_���)���/�5[,(��#[P�C�c۽(���^�ts��Iρd95ll�"��W���X����8x�C�tA� �gm�b/�:��j��?��а���LÍ%�#�'���؜pl�f�T��5���oM:E���*�cV�|j�+"6�[�d�`����p�U@��<�͕r���h��9�_�_
��Օ����n�5Qڷ.<4�{����A�eLZ]�,����݀���и�����V~�ٵ	;$;T�)���6���X+	tt�!7㔞x�Aa0�nE!���&1jAR��G��B�S�ͭ7D�h\:72/��@Q���vv�#@��WK]Ȃ1���z>p�G�V��l���b����N�d$X��Ҽ�����
�:�ol��@N��+6�t�j���go�dT<L�C�y.����C!���_��9���G�dK��qrX|*ܰC�����8�#��#��64��'Z_M��;L��zA���s���K����u��$_��?�X
�����9 z�t�F��R��ko4�s>6��)���1�I{�#�4��$Ba�M�姞�O�DK+܊m�����a��tq0 ���V�Բ�
~Jc�H��`��0���-ޗh
���;a�8|�8H�������(�i}A�48u1��O�[<�������_j� ��՟����DK"Ux�GS>f}�v���࢈([Od� �'��`�r׫�;	��Gx��
�c0�N�)�t�T���M�Z/�[�Jc��B�#�M�v��<�o�c`4j�|�a��D���I��� ]�Z!���ۜ��EUO��'5�=o�`�~ ���9�'5<�������HI���#�����������yBs��I���_�(}�W��FO%ٯϏ`�̀@d���KjO�$����k�+F�j	�7=�䁉��bt�yjW�	''C��1��jp�ObGp��^�G����^��x>r^�k�@O��䕋eYh��tl�K�g�N�O���Z�E�B�h��T	ݫ1�3�ܥ���?(WnU�
��P��s~�&=��e6!�h�aB�}���eT�3��LL��@�Le.��L�wNw W���tg��i���a�t-�*]u�Vy�D3Q���e���vy��I1}��x5�I�(�K!��+��q.+�&AE�1�5^K��8�[7P�7Q�bå�F��B+��/%Hu�|�٪w�@՝:/��t���H���I�X��� !�n[��I�=9�_�7R��W�/��c3�Y{��_O[
Y+�V�{A�CZ� �P&��7�Z���n��MH[*�o���������*=]T˅�}2�L9�T
��5Ujm2�/�8��NR��ͭ�j/s��<S�3����3� �/w��F��Y��,[��+v:S����A����M/�N�'�[�VY�.}/�%AK�Mғ2�\���o�7W����+�KU=�~8U�_xY_,�y�b�;H�Sv��h ��\�yX�τGȔ�)�D��tn�p1QAd��	̏���t�"��Ϣ�K��>Y���s�pq8XM�lD�Fy�AOO���G�)�-�ɞ1R�_�垛����Ny|z���4�E/�D&,'�ҙQ�s��v��HV7�����x�!3-$.��x�ˊ���,�˕9@�.�;���iql��	�H�-��_2=���E��ֻ��{�c:"����%������O1�^f��wԟ�����ᡧ�E�D\�̜qO����j<";Ǹ�9i�1xn>6�����~�܌,��+d<x<�P+�z�K�����o)�ea�r�䂨����ь((�@G�>B���J�O��\�
v����-�F�}e �i0����rƶp'e�M�ݬ~�=�0�$W�-ߢI��;�����O���Y�r�E��a7xU�{
�3���f�������6C��[�:܎=w8<�̴��ݠ�p�&�ֶ#���'�;ʸ�Oב�6���P������(���p�"�G�k��9�	g*S2"���~K�tgr�̓�ٯB���a���>��Ekh������|_j�B����(�Q� c�d6`��wZZ���*�ڥ��E�IG;:�'#�	�H���0���]^����V��jn�?eЄ���Ј�~⍍�d*����Eb��<�;N�ɹ��ʉW`� K�ܺ������!�̚�;v�@��.d!�Y5�:��M�(�`�^HE�-hH�*��.�%�����n�;��c�{�'��g�_�5����^VOI��QfW��D^PB��`��0��:7L��c��\^	ߒ���3-��W����W�ɐ�(@Ӫ,��"
�N�{f�u��,v�X@}%�2/G����j.[���5�;�n�1txfҹ�n��g��6%b��Y-]�����N���;�'WɊ�H��k&��cǪp"��� ��-xNj���Σ^[}���?������)��{�
�|T�hw4�'>�3U�W��2�a�3u+�a�c�Amõ&�@aHSA�UE�{�i� �ix��;�י��dr��妙���}��XS&B�|CE�ԥ�A�<���ԋI�� TI��[����t�[W=�hO�$xE�66Mc;������5嚔�&d,�J�!�+A&l3c�	�#�q���f�X��N��.;G��ߎ����Rz�hgx���D��N���j *���٬�Je��6m"�/~�28����{olA��b@}�����k�]con>VT��*��`����F��̻�ǨL|9W~���VU��:H�Bd+�m�`�OIKΌ�������[�����lw��`�� Z3�q��J��R(}��@k�|k�qG2uƤ*I�^UU�;ot2b��-�Z����DP�@06��7�`��I$ �5�c��2���HNy��B!Yı�]4c����\Ĩ���B������Ϥ�s)�G���c�ݠ6�О)97)�:w~L�@�Ĩd�0��֌K�YdQ�[M)M-�����3<�Ё��o���2�Uc���#���Ij���b}�A߫z^گÆ�Z�����Y)lH�	�����������LJK��}b"��Ew�C�߾��E[�c1���K�k������f�PԂ��u���MH�>~b[���]9��}1\>���c�m��	h��j��hf���%U��ٷ򙏭�jg��<s;���'>3���_L*�3�i4P���,� $K�?M F�� ʺG���q��QY_N{�SNثUz/�Ad">)h�p��9s�?<fY.^�i�5f4����on�
����Ý%A}�'��;�����)~	!nr�+�%RP^����K��癯���=A�
RF-� 7��xԡ�QɕD�J��oL�>J��Ig���8�S�I<g�}���DlW�06����gu���|#�Mj�m�Ăt�q&4`��^�<��e�Ӂ�`��!�M�!k���Y�Z�a(����^Ġ������� %��2k�'%m�ړ��M����G�#�	��"$����%"2�9�X��*�&��1Pv�j9�2dĮFs�ʧBj�(gw�Z�;��	�(7[4�^��!��
��Ҝs�P�`RM��I��E7(˕�\�!"q�S3Eu<D�hђ���Œ�� �X.#,��,���I�S~�s�$%]wa?���UҠR!�����E:�gc D�M�l�I�U��P$�A `���c3:�>��s����n� ?U��b���Bf�G~���7�>G,��d3H��뱓��96�vx'y@f�QE��<̻_�i��<,sd�)G}"u��P><����7�@��_Yl~%�a�S.��̴�
���F--���X��D�y������#��9y`�Kb��緁���?�W��
�J���v\�M|HkL���6CG��!{��f���.�`l�8��[}>��b���I����r���(~��&�*.# ������E��7�My�!��S�I��o��(�TN ��Ef�������j�E'���8��K���XjfS� ��=����QI�ntp]N����O��̊1'ս�^��V�>\3A�3��۱U"l�_��.7;��ʪ]{�M�M�X =<J3�o�щ w�j�^K�� ��uL�B$���_�k;� ��0OL+��hZ�[{��&����H��(�䜡f�=OBˠ�gUn�{e�}��"sE�r���\uݡQ���3�R�~�B��S�?�#��ѯ-A�2���}r�y�S:'���:���a��c	�r����|4ɷ�N.k�W����!Lz����_pR�LC9HX�C/F���y�L��	���i��/��ж~.aV��NVU���\"��駯(������f��X3*�����,�<\7��\e_r�a��l�	�q�ln�4�4�cm&��K�#�͵��aI2y�����݋v]e��z��;b�+>+��<@]*�9͵
8(�kd��A�+U�Z�̱��I&dt�E����O��TD��E�e����	�^Z�g]z/
�c�XK0]�!�UiZ;oՐ#��|�ͨ\V�D>�	���ve�!�"������ ������R�\��;ά�H-S���)Xt�ö<��>�e&�\h�^��^y�ԛ~������ �Q��(�~@��+'�Fk�y�F6��.s���|3����)����I0���@���șv�	����ZSZ�ǿg�!��� �6TX����)[�wT��b����jWۆ�����j���sq.4`��)�5�� �T���*���E��6�2[��;6 q�p��,�7�� X�C�_l����W4�ǭ��^8`�|�J�����"D�/]�x��m�$W�D��G��&I�]E{"�h�����^���0�m�fZq67�;7f�O��B��+�-�݈/v�6S��HP�65�
kd����;tPr�%@�b�#��{eFW[� �KvY�ff�&�3ܝ�g��O�
��~3c�$�ؔ;��gv���&���m�~�/�{�� e��_�������%Of�:[3pS㥇qnd�ߒ�S�a����=��k�&k��W±��F�q�=P�;tLz٦��Zb�SUF�SA�G�lt*��ɀL�g�st���b��c��bb�"^{� 9&���s	}���=���=.�㵇�.u���Q$��`�$��X�zL��ՠM+i�Q����Շ���}�Aol)��nZ0�*�N�?�iM� N��s\��7��{�7oح����/b,��r��)w�<���)�L�4�M3��.� Ag��ϳ���*��ht�r�s�t��%;�6��.X�^��(�-�rȨ_ �q�����4�?⸽)@�~��W�e��~)k'EވN��������=6��p�_̐��Ѿ0>�zn� �Zcʣ���fc�n� � 6n���%xcS��g�6"�4/�U�Yr��sk�%��=�����kq.GmΨ˨�Ȼ��V
R��U9BOי�ئ/���d^�$��dd�v~�;�z�ʄ@��"D������qa�/�D�V�n�I�m����n��*�s��m��8~_��NG��-Q,��J� 7��f$3�y�~s|(b��N[X�婱;(����Sd�o@u�hf�,���),��.����_��`�����E��"��"���@����N "�a�dE��b�#�U�vl8z�b~��s��Bm�9�Ŧ�B�����Ł���<D�ulFZ]���U��{�"�3'�H\��UK ozM�fH���+S�-��7��CP
{�P�:*p����iwDG	�#��������g �����v�S������NN�E_��p:Bj���{>mj�[C�:M.�g�?�!�~~Wt|�Y��V���ہ�.�89ht�S#��]�Ycr@��P\n3�+��]��	�oӋ�<R�Z�ю) �H�J�jW��KȽPgk��}SWFk@]��3��Ka�wl��*��,y�Nw�0�y��{D�ݙ�~�J���]���sx._M|�m�����:8�ۖ �7����<�`�:|g9¾;(Ad�BZ�4�w�1��+�zo���?��(<�O�C3���C���X28#m:�۹�$��c�j��I��Y[F�]q�aBd��Μ��0xľ�Y�{()��9!k��J��A��.]���J��%�$�$�z����̩�n�+3�a��}��'��j^VY\��+=}O�"�H� ����X��
���_�&��	S��P�ɩ�O}谮	��C9&�pw�}Y��-*v1k>b
�T�m̓?�ǫ�;��:VR���)�{�֏��'�����5 �K�:�̨�k��FуiQ����gb���T��T
�/�j�x|����^RG�u�땳� �\{{��:�hӝ/��������I���ӈ�"����Ap�Re��9*h�ӕ�_�I�7���Z��*eT�.��7D�:��׫�[ܩ��
��(���!aČQ��	?�3F�̯���)-RY�9/��9�>�����0J�8FAwi��B?R�c)�G� S�5@�;;�AC�(�
�u�vl�;�	�ڔ#K��ئ��r���l������z��ݖr�&f��qkk|n����Yv�>0��0�`c���|Z�~�!q�s*)R���I?�r��֍�lLqh��g-)	y��������3F�x�����D�����c��d&0G�
̼���h�m��Y�����@�<������{��2�Ġ�S��p�Txb9��{S��`����Y��(s|�k �^�+[��;�e�ɴ��'�l��Y������N�UI��WMթ�)k���a-�It��'�@g���5���l犇GaD>�'�n�	+�����yl���fzr�&���Ϻ�:��X�wؖ�/���t�s��v���e�M�H��?dX�
͛�p����8�D�#�rP�D~y,C]
����؁!����_�t%)}�
���͔$&�Q��*�\�t�_BU9zz���-�Á�m��}ps�M^$�Q8-�8j[5/�W��꧖��n���v?�0������}^��@�E��m��Y�c�[������U��1�t�F��g���~q��0�)�t_P��G�4b t�z��.��J7��R��ȅ����%�p��L!I�B6��eBS��C�R�<S!E��(��������J�����҆�Y�����v���he5�?�v-��qo5T�����}�o۬��R@�����!�.��&g��A����e���Z�L=w�+�-{3"n1��T@���A������x3]�x_.��ըk���пtN=�*y��}��B#�إ=Pso����H�*m3+�x�]֍_b⋖`�!@N��1�E;��-� ���w�)�X���S�>��($LX�#�V+d^�ޥ�겟p2���E肢M��	_x��88��ۇղ�L�?�*o��\����� ?����T���I��^����������Z�G�
�ϐ�������rgW���s��"�ꊪP��H��?j�d�\���D�L��7���\����� ?� ��1�IN���n��_VS4@ؙ?�T��ؠ�5MR2e���pJ_v�a!�T>�QnX�#�<�� ��Ď�~��n�W2g+4��&��ɷ1���R2��T�o����aCx}���^�vh�)!���(im�p�ͦ�Pb�Z��
N�_"H��d����/.I���R*?)=^w����Jk�T���`��lWw�d�b�M���������?J�K�-8҄b�<�ۗ���/�r�0��U͉_���#�U%�)��5Ma	x���q���*Au��~c�˩�)N���1��F��tz&���ؿ��C������G`��7l�ʳ]*�8��� �����4@�m/#�¯�rO��5�8�Gʰ��_
�ɫ�~$�������5�)U�A~���=	��]-'���{d��!��^7>�9H�S(�+QV��[���x���+�xz��u!��{�h�����"U�����;��җ�B����{��w��+�����@�R�u,]�HVL ���/
t��W��=�
6H��0��/ߍ�a�b\��O�O1��rd�W����z�S�̏;�p���cε�+ڈ1z}rG_�^��/n����!dRud��9����Y����l2c�%�������j_<\ъJ
�G+\-@���,ה�1{���W���x��ٍ�'<��eM*ѷz�?���;ޚ���ۿJ��@�3�D"�����>a��s<kg�5`��_������5����p/�z�w�Ď��4K���
����sx�L��	��J��E�['#\3V�<N�B��8DT7����rD06���?�im`u�^��d!�@"L�XՐO��ڇPN�����d���9`N�<�ݭ8[A�Wu*\!�oCCsrQ��}���7G*1�o�L�SnMj.��s�Ǯ�i��P&4;�Ʈ؃6�	J�����6��y�*1�2��y���<�$ML���f�=�Uz	[��1��Z�2
���,�� �PB�~���Zj(r@5;����U�s]��>s�KA�*�=AY�3b��������齻@�pI!y"懶�c�M�S}Z�#�6A9)?���Hq�a8�1�hZ|�_^%?Ҍ�5�L���@�X�����'��m'��f��
Z^��<XL����ܘ����x%+{ы��	6�:��.|DG�E�؀Pk��_���&_��5��K#��)d0wu`�?�8)T�����m�F�����-��Y?��_� ���얀)�� ��r55�PJ�� ��Jm��d�UdC�4���E'uGz	�p��ʜ�,��i��_�:� �ǿ�9+��:�5��p�\s�p����0a���G�OjO9�QgT�/ʓ�����@�B��S��@�������7��]{����<�+n	_c�'k�/m�$�n+��]�-�t,]�s�tt�l;���}�4��t�3,�ZK�����X���2'������
l�&ېC�ك���*�D��F��թxz�v9X��ޒO���_�?_`'�D7R����hFP�=�L�#!1-��t�$��^�L�yx�		��%� ���JO��6[=���ը�{�c�m;fi����{�q�M���Uu�[b8�a�r��~�Aw�D����aj̶g�{.:\�
'z�0�|������Qz�wAh�A�W�/�%u�L��N���������Baﷃ�U�%�u�gb^���d�P����Cb���^p`�@+�y�&�=���i��t�����4&f�Y�����������QQ��'����'��O.��& ���n�8#.�^K��]��p=B{�cU�̃�'L�g�>֙[r^�J:Ð/���k��W�Dd���s{�+��:w��(=�/ښ.iH�6���?��~���u��$�]��20�1��$���TZ���!���ؿY �gh
|!H6����ڸeZ��H��G�
���G���;����CW`@h��y�Cw��0�7��h�1��9�Rt�\����<�����T���<L:���¥�Y����e�v>gJ�6ޣEV�=�FٻA�.�1mH��X) ����L	:����%�{=�a��-(�$�B� $�N��~�j�]�t=��ô:1����>�`C
(�9�c5�sr���nu���;)ޙ�0�3��O�� N^����0�c��27S:��K}Z	�k�׃{g���-�10>b7Dʃid�P ��J`�-H��.&
=��W�;�R���)�1��������P��q%z�vu�x?��#ǽ��,8S�3����d�fR��w����c�����8㾭o��G�TQ�2�x}d�
��v� j�e�r�1�r���3�j�I��̫L�6*@;C#eN�{�]b
ph�R�'8;$��#���n����U��z�d���Ŝ�+�̦�e�����v�0�����?�[X>���$e�t�v)"ȳ=�/5a�<�œi:q��;<���S�qY�כ̹ѷy��ź�g�"@+.w�bn�`c�}侢���R`�����6�
KΓ�I�6竍��}�S���ֆj�UJ9�~�n�xa�鞠p)��*�Mt�Ğd�c�0�g�3s�`|�x��TG�gͽc��i׶�r^�1x�~��c��Uƙ@A�Q��ى����s�1g�2�_E��1�J�YkK�1I���+�d���$�����j���C�d��z�*&�gd�^R��k4����H1/]1b�|�b/5ya�v�s�ק�o��B���k���a�Nj�u������)Mt`/ǢZX���	�M�d�2���&֧�CD�c���>�mR�
�X�n�,�P�w2��"c��T(�m�3̬�(+��`JF���\���Ҁ��
��g�����%�r|���-^���%R���ܲ�
��Ҭ����T*����*��>qz��b&���~�\�E�I�LCl��S�գH5�y,�(��jnS��f;��c�R�p��Slm�dc��5�Au5w�w�̋X@�G��נ�y��>�*��=�5���H	-�_�f�;��T��.�H�����3Cs��BO�ٿ�2P~{��ͫ
7�w��mw��5�д�������]��;��Lɸ�ol>c<@4Q��SvMv4�����a�H��-/����J���73	�c��S�cA(ԃDz6�Z��@�v�u�������}�7��ӟh�n�$���IC�:�b�A��D1����L@y��d�|�qd\�	�0iaT��F���ӏ Q�(���A<D��T����Qg�B�(�:m�d���h��:Y����=�8�)��b�A��P�ẟ@֞Bw|�0����^�����33��
TO�0r4.���]����,�����b���b��7�Fh7���#\{_��K���&������J�7n*j�����������g����Tт�<J8�[	a�H���b휗�"�T�X��Rtl`AP:BWν'#55�	��ھ�T����ȫܩ������SS4T�p�ď�Q=������������v1�6�
L\����)���~L(�h<�Qd����[]��'�4N�'��y�C�~ߎxD��������Q��6�Y�B5�V�wn38��BN�g��m��H7�p�R�8�*�x�6Q��"���x�m���(0�j��{�&�cy�U��2H������������it����T��2��7D?�WQ P�}�]2À��Uy ݃���@�& k�I�5���/tHP1�on������d�Ui���v�Rl�+�N��Ip����c\��t��)�����C�U�[�
w�ec�����
�]��kF�M�;�Ԑi��[��ڒ��%�	$��xγXǀ�^���~�g�:@���4S0D�&\ b0�Mʞ��!���t�±"�80I&p���Cr��L�	��Mp<sR��e�C��}��_ÀsE5��b|���_����f�S�BO�g�n���IZB�M��.��#�uS�q�<����@�3q��L8�ZT�y�����̏!j�D&�7�R�V�ػ�b��6[���bGFcW���6�8飬b3�u��?7���x�7Wm��J��'����Q^����YZ g���*ц@h+{]�{Mliم�������k�ξ��&�b[�c]F����ر�
xT%����b\��� SE����h�E�?�pAz�3��ѯ�C�� ��p%t���h��F����^&6DFM#��r]�-}޾u2��Z&H\�򆶢�F��b�$Ğ���ݵ�QqS"���TC�� ��z6MΠ��wf�ļ���Ṿ�ߒh������u�������Aއ���iR�X>�H<��g3�{B�����`���D�&�It�����P��,A�guZz7��%<鬍U����D�
Җ�0,��^�a��t�Ei�t4?�s4��M��Z�Ĕ����f�3�)��37�s	� 0�Ff/#��'�7Lص�����+�,��u�A�l���hw	'X3>���q���A'�4�AW�S";PP?i��(��D���ńqnK��i7�چB�*���X�>!FyA�ס������O�K�&� ��u}^���r䨛;C�.Quw��?��l~���I�
{I�6����\UD8�W�L�ܪ�b��c	���PC� ��K̑~t��92\-�>�YC��7��7��T!0y~���-�u���3�X��X��M#Td�V���)��&��[�/�L���}K��������O��c��I�U�|nj˼D@c���Ű��u����@�K����I������d��� �q���/u8C��D��C3���y½�\-���-�=�1{�r��9!���¶ê+�r��3R����N�e����X�)쏆���1ט�϶ŗ�6�Zt�ܚ4 ���lhZ��,ӟGM+���7>H�QHsO	��4�32���ceD)V���j�Y����i�Ū�{tJ;��Z!~{k�K$��hs=�0׭?�u�R������k�D�n��'IB�Z��`�(�c����6�^�>Rߧ��`��9!��O�;b@gcC���H��끒��A1���Ɂ��@ٜ�?C`X+�>�PPX)� n�V�ꮾ#�|N0���@k ��&���E�������f��/g{KԀfY=U�!w	�c����A��͚U���	�:��Pf�J�*e����X�~(.̊Ty�n
�WSb�T��m=�త�ꐞ�K�3$%�t��@�zeo9]g�<J�̹(�O�#�[y6̅Lɓ���I�D�]t��o�a���S_W�)L4�y�3��,�����M�W_y��$���Q�[�����'%:�ha�t�_�M����R�#^,��(��%�ST0���L�3l3�.��L��(�zb@8P��a(#�'䐠X��k7X�(rP�&v*����ڡe��∵�l?�P�jmC�²��I��y�u���~?z���Dt|�Q�ͻ=��5���;E����B���di�o~BvC��G~�h�J�~�*�IIf �"�����R+�\2{�7yd���yg����,f���7�����W��as�8��CY%f)�� �F9�Hq�$��6���Ri'�pw<��<^(e�3~�����/��"0�5�*�՝t�� ��u�ĳ643�_� �h��u�Z:�oV���%�&Ѡ�ڙ��1��M�����\a
>��3��͈純O "
��	��@��!!����觎���lּ���AP�]q{{J2�aU�PD�-i���Q�L4����f��!������"��i�d�x19�:{����b�<|.��dw�����I&PYz���mf�V��A������yM�;� �)� �nrmp�7W*B�������ջ1�Ё���s��4�
��wB�W?���8�s��]T�2ոEMV����u�``���4�k:Ȥ<�Ȳd���%���`$Z�a������p��L�S��g&MMG�I���Tz�}n�D|-����Y�c�?L�P17J�W���%�c������=�B����g_���su.�_�G���@"�<��x�f^%�q>#a��q>��k�P%;nt8My�9K pS{m�������E4z�-������h�e0��υ�N���?�T��Vps��X~MkMXG5����������,���5?ʣ �T�|�m��߹���ҁχL]�k�߉�C��_ḷ��89ⴅG�b��!Dw����j=��2x��9z�
E�iG臠V'l���XB�m��AQw&~w�������,m��U4nѤ]�E�Zݲ���]�V8���w)�=�1�?d�@�6@X�ID(�*�۬��r�~!�����ܣ�8z�ߕ�-��E�F�.� u0t�]����59}�h|�T���v���G!K'�*�E�{b¥B��c� `8Z�D�
h��l��#���A��8�O�E��˕��n����k�B�Llg�d����v:�W�F�1�_��;#{1���Dq<�+iZZ\�kh�lA��.�ԃc�����)���dr�ۏE=��]��^!s�����uB,�6��wR��r5�6���)�
�*����`O2ʒ׾���̈ `��?)����n�u(���_�rz�b*/q�'�z��3�4G*��ܾ|�N���5ñ6��dǅ�w3�(�J'�y��}�Tꇹk -���=�G��9�~���A�<��n=?ݥŀLf{�}�r�y�:u���>!4���u�Լ.��ԔM=�k<����a{�,�)ꫢi�j���m\5�pN5��%d��E?�X�c��֞�9�e�)�&�N����|[=t���Ǧ-�\f����2L���a����sz��QB1���Y�z��	c��)��v�ϡ-���>�+p�>��:��۵���Xc�[�hN����"��?��K�igЊ���~c��Ox��c�7�A�y�D��9�^K�N
c�,\����uB�ٝ��u�o�M87�vU;'�2�@Jl�Ya+�k���:��<54�gL�M�V�cL<À�p�J�s�{@2��"�qy�s�P��F�h�a��|1k�>]�IC�����έ	� ��K{u��8B�Ֆ�G븉Ӧm���v�9��F6����6�у��(��9�����l8ě���̸�J�G��C�u%�{����Sl�:��7`��Ϲ-[=�.�����y�UcP�ꔟ��5��	��)B]��*�i��fgB�@��4����%�]��N�8j^�tkD����B/W�e|���|����p5�w��@+xU��*Y]�<��N�V�P}g'���9Yz�e��`s �J(��aq�md���C-{��#����tٛ��6�\>�E�w%�b�Cr��������� R��k�z��b*��Z�J|����q���U*��h��8O3��X۶��-�ůO��%��Q]��_��Z�=�3J(�ꇘ�j��[�?��ύzX�4���9#���gD֐X$7Ϸ��`0E�MxӁR�\f�M��_��bL����	�r�/�w��	�j�B[w�m�K.�}S@��� S��ņ����k�5H��)"_Z�C��}6��?bBt�z�qx�#���{�Q�|	��\%���q�a�<��6\vWԣs�d+�G�z�T�0��-���O��>���,� �X���_�j�{�U' ־O]W���'z����]��E�׻��}�|�|�Lu�4�X[߯"3mk�4`�����ܾ.�ÿ`gcHIJm���wW�>t��]�
M&\�L��j�Y�(_��֣L[l�g]����k'���ͽI��R?1�O5X�����;*��� � R�h��ޣ�BL�3څ�Y���ZA�H����l��L�.jD&��}_����r2�8�.���q��IM�f6S�@�䧎�;oB�h����.��*.כ�F� ���T��� U)�g����.���{���L�8��T�a����y�~��q����	itoq���F>,��kK�Z���"�t
ׯ���`��47X^�{b4.S#�8T Ь�:ƛ'Ҫ`b�i>A���( C�����PL5Yo��Q��@�,�O�:�̥#�����g�2$
��}��i�T:D�F{dU� c0<�}��T^h����B���B7ܔ�g{ �w��^܁/�,�U�|��@m��Q4�2�I�%v�آoъg���QL�a�t�8f���H��6QմTxv����Aid��,���d�Udʿ�S��� �bA��k#���l1X\��4{x@B��؂J�q[I`�,[ �ޗ�?����`�5Ǧ����t���:��NY!/�a�&DnAQy�F����6m�����AЃ-)�ݸ�B�SX��k)CG1�_N���)u�O�����
#��^�K`(�jO�ie����,��� ��ͯ?}/n��ߋiBb{�j��N ~j]�?wI��ި!jdD��yU{@�{��+�/6�[���8�� *m7F���@��Q񰪎2�#Ez��Fc��p�hK��w
�\�ǯ
����N/M�df-wDW� ����@��I�������8��_�`�_��ʤN�� .�.��0cjŪ- ���V؊��E�m1ʊ�& W`��ğtm�3�v�[�(�J�[�02��U�0���	�\�uW�}�E_{Ic���P��QeH@������Y�V��p��%���L�V�Y!�쓚�K'�s�8I����!��f;u
�y.��Ӓ����f�}-�}%,+�Ӯv�f�?k���g��{��|��փ�/�/]㻿�	V
�O���w�����@��֋ˋZ4��z ��Zq�|w�~��n�[��ɣ����%������8�7��6 �kY}S�Z��@Ѯv'��B��
 ��/�1ϱ��E��f�ɻ��uYQ�o�ych]�m�0���8�ɄR���D��NQ�W�o��Xc�<Toaf=� ���3e^����(�u�����y�4/̋�5�>;�̤���������0]���8��(4fml������Q	�����Ԗ�8�W���Q���x���hJS��	��H*$R�K���s��f�]ki�P.z]���ci��	7��oz���[�������Q=��u�}i{��,�r"�K��G���)o��0��+n��Bc���^Ԫ�}�׼S]P��p�]����!�E`))�sI䉣LT�~/kMn/��5��{�i���Pm�TUϼI�чmp����n�mv+h-����Gj�uf���N��r4�.��W��g��`�>�0���x���l5G9CB�uRB�����D'����Jr^�sx��B����g���1������\�F'5[G.�v� {��c|nj�a"r	z!z�m,N&�vÔ_i�
`����\��0���,��_{Ȼ�͚)ǐd��8
�&J�Rv(��r��eFt�g�÷����q�g��)��<����U�
�\a+�a�1�
~s]?��#yi41���S�k;�a�@���+�(G<���G�E�`���BQ�FR�ǆ��u�@%pJ���0%�]�"Bh
������ԂTH&�t*Yȕ4�d�+AwL����K�̖���q��"&���fEz�.弜�/1kSy;��w�9V����{_��	�[�A	�V)�?��p�Sgq�O/��ߕDĉ��]>���eW��s���!��)�ѫ�����s����U�٭���A�QZ���>�so�]��Sˀ����W��.�T���Q�L��ut��#�8E�u����b"�s/�v�u�$1��@�O��>�0C٣呅C"O�� @��劦7+J�HQ��{����@�X#32�T^�;�	��T��>:U���܀��JC����S4<vB���)�7����xzv���W8@�a@b�s��a�H�H�)���n��u�B�e`^< ������X�z��9�
L-	K�Kf�v��#�U�/��^���K��{�*J�����n	,��n�;�ec���Z@����[6�lgM#&Tl��{���J���a�?��r���g�G�,��2r�T����	���]Wd� �DRx{0��g�	ӭ��	Yu�R��R��>�"��Zy@!�@e5�r*Ի��W�@h eU���u�Y��^��o���/��P3�RJ(��3��L��`�Qt�efn^+.�]�!n�:�6��M���Ɠ���F���"��"����}�+�ܥc�ҍM�9�Fe��E	V]��f��
�5Թ=3��K�,M>@Y�k�]G��x�
�� ��_��p�0�v�wأ/�G�v�ʄ�������E��:Y�Z����K\�g.Ya(�����Xs)�u��3��W4��X��8x�S��,��lE�NA.n�!kG��A��Z�5����p�!I�:l4�z���8��'ފa�Z�i|�b���e����M�?��'�-�TL�U/5�1I�z�����������%?��w@����ǝ�&�,��!����W�N�7�*J��pp�:��g�6,��hv���a|	�- ��ɸ>B��'z�	��$����Q ���AƐ�y���юi��gߤ�cp?>�\��n_���|H����<�|�B����&��$1��H���Z"'}���%So,�y��_�n���䜕����{SAhd/r��_���H~)��<ȓ�==�I?$���9YG(�L5P���|���g�G}Z��G:�kӸ�>/�{�d���� �c�S�UR*�CM��.SIy+�T妶��|�9
�1��/&a;�LG������DH�x��t�{ʜ���p|�l=��]�����u���˖ֈR��{�����`rQ�t�~j6�-u�^sznh�_T��F6"�g��c8?�_�F�9�T����LO�=�v���c�$́T.r[���H��E������� s�}|�zia�eCwIx'�s��h�?�ُޙgN�]��~F����_C:M�_jȀ��&���n�2J��=��7���;-9���G@��ُ6A�dD'�bK�V��))A��&��g<9��@iT%�Ӱ�nx�l�5��aP����`�WYaN�j����˩)9��֚�toB���L/�Rw�
靈�K�� XG-���*odt�@"�#q�*K���k7ǳk"��^ًc�O�^������)9��}ZK�P��4���k�Ȭ�����v�q� Ū�O�-K)�+�!��	7��Y k��.��wW�q�a<����ܭ����7.;l�Ӑ��^*��7����b� ����БU&��0NzNk�34�[E�9�C�o(�^�5N*����T��J$�@��*�l��rɎ��_Dv��C�����{��	R�&k�Y�s
���>r���*�q!(�=���&�����e,?O��̡�!NfT!j���,\b�5zC�P�Vz�L��%�Z�G/S���\ �JF���� E� 4�g� 	֎ep�չ)]rn��t����nl��?�uS�-�m�(��6�b(Q�c �}�����f�-��U���L�d �y�ٺ�^��5�D��4׊����^��t��2}%�����ރZm>_e��}&D�RܠQ�Y@T���ͺP�
_�-Y�W����������K��d��c�V$�;���sY5!=4�wM��u_��S�eu�B�qʶ"��Ւ3�~����K�+w0rh�o�8����RY�:�k��yV�4Z3��1I�S!�Fŗw`6N#6���)0���!Ͼ���+7t�.��g@���k���ib���Th����Q~#�k�*�C�&)0p����6����S<&#,��=1��.F~n�t�S�p�M�>��g��Dн��ko����N?5J"f���#�"$|,�};+�V�G��`y2�ۘjz�k;��s�קM�"_�Ű�Q������QD$�꺄-oF6;K\��G���E�ʉ�\���ȋRG�̈́�l��|�"A��ʗ�l�	��g,�Cr�ٲ*2���R���u������P���.�w&���,�\�?��NM*;�L�M�d�ƞD�p:� ��ô�b&�hD��+�\�y��*+sB��գj�=^g�\e~��C���ׄKI��I��8��Ť/$(�:�����A8���q�$��;�d�B�l+�f�4�$a��H�N��������va.���j ��1�m�)d�?��/?�$��6�\'�ht�0:�J@�<UD鴹��2)�����u<�P�A4�-$G˟��8���\��:I�F,�2�~���w��K@c �Ϋ�!_���4�cXe����k�]@�r�ʤ����'��r�i�*�Dy��{=��Vvd�x<��@F����E���o�fS�<=�A[L]C��q�d������b��b��wN����ӹ��N%�ľȄxGK���ў��w�+y����)�?9
F[	m�)����d�k��*'wx��^Nm��~j�x�y�����9f"�KJF�{�JO�����ԆX�p校��j������Q^H�L����W�>�g�b��ݵ_Q5�+Z�QX��r�u"��]�1���Uk�4��s����Y~b�`!9冀�{Q:u�����Y=�U���Ӕ��|c���������ε��������0��P�ߑ��X̡��٩�m����a���wO�I!5���P!��Z��
��'Ȇ�CPJ����LT)���9�ƫ���y;���u��Pb�I��z&�¾�D_L����[+i�����P6��{���,e ����/-4�r:W���Ae�[��\��L��`�r*����79� ��8�M/"����(��N��Ɛ��z��?3=�q ��.nT�h�c��3.��C���o}�Bh[�(#V������H��g:�W޾&o���h��fȥ��T&R@�~��l��e�R��H\�4�^`{Ј��.[ꦑV֐_����vN��'��6{^�v���������Jw�xCv-�	��(Q$��b�ʊH3c�*CPc��Y2�����(f�.���̪k`�Oa�h�p\y+з}"&X����v�k�I~�y,R�����W3Nh/�8��^��$I�	l�'|��C1��q�6�73~��\R#e�����@ ����'�__����b�2�x$r:�U3R ��d!.��_m�����~���;��� ����w������"�ISd䐥H��<�і^B
Xa��"\�eZ�����#9K�d:{ד�	�.�@�ψ��5ҝ����6����%Gk��+���MJ$t���mx���e��� �ZA �Z�_�Q1o�V���ݰtF�� ������`�y�Ko��+�6��1ܓt@���r�q�%�DQH�yF�-������$����м]���C��u�b��P0��ۀ6�W�M�!��*���^�M�Y-Cn�TmK���G���z�_2N�2
�n�[3Zi$^��x�J3y.0��ω�bP�@�z`@�7q(���>�)x�a���Z)�h�<1����\��֌��`pm��5���d�\��-F���;�����E�#:�9&�~�fc�Gp!.��5��V[���c��@�)d��`�k�^� �5b3�*���ѥp����U�!e��'����xj{�>n7ߪ��Y��[=��b����ϳANT����EE�2%VM�I�(�pWkܱ3���:��wT��w.�G5u�dV�$��{�F���w�fB��6�t���?�h�qR�)���65k�)a[!(�1M��^��d7�.SZ%OYIl���R��d�zL�oL��7��ol#:h�M~X�/]h��H=D�#��	�_�e��"�Zul��'q���s�������� �^q�2�Wi'3G�swqQ�z,�ق]m�"Y��V4��D�~���a�jj?g6�nI�6����Z ���;"Ү�zH��X%�|�\ꨯy�p�������A�p%�A#���Yxvӵgw��3���ˣ��mZ��!8/Q���1��Z�b������3��a)�3+�����t1���)l�ls�8/.�
�,А�ƌ�/i(�}:!��	۬ʧ�q���ޔ+�vz`��c�F�Zj�f��Zz�r{�F�VEߗg�D�&����s����y#�h1q3���$p7��L����瓷dC��!+Y!"��'�?S��t|���J���E0��'Zr���\�@-L)���쇧#@��0��B���M ?69�%j��0/������t��kA] 8��d�Zb$I�>�q!t}P2�A�����,!B���-�jD��X�1<ߜ�c8~g+E�y���>58�/��_R��9q)cm��86T����DD�����9��SzTV�x:,�v:��]U+rE����u5��'�6��!��'Y��	u���0۲�ǌ\C�94j�1e��P
>6Xk��P!�i$W
�̃�.6QR��p�Ih�*�����hF�L��"�1��_�4r�����$��yT5�}��+�>�Nm�^0��m+�ՔX���ޭ]I(��R7��|��I&�PTv�p�_��eׯ�O�pD�u<{}�^��@:oH��=����r$h��b��zRl�#r�������T�Z9�;&:�p���2�u�������$*�:�(16@[��D1�煳+>�y?�(ݝ@lw`���Ұm��1@���Ƈ�b�	�ظ\��	�h{	hN��q_H���3������T$���7�S1P5�)�b���6� M�qɕ�������~k ������yRb�H�Xӣ��j�_w��)��%�x�2��J�a*!*�����S� �k�d�p�3� �0�gU��E�-�3��a����h2p��]�N��bٰ�̞�JQ@1���p�9�[QeM��sե�Z��A�\�O���T����^w�ru�`뉟Lss��q�0��.��}�yi@��ڛ�cP�3��N��8��tȊ��!�-	씱b�:8v�#s z���A�L\-�7ny������`��T��nMD��P$��ۗsU����:}���)(�<Y­��Ge�qt�֓"�0����M/�46MQ�Ա�p3�r�E��gwrfa>��;�O�r<Hg����b�y��P�=�v#:J9awU݆���şbrz��<e�n�X�o�%���.���#��-�C�˵6"x�c�60�m��57�����.H�b�$]\y�t�++����\1�|^����l�p��q�.��){�ׇ�h�[�����e�V1OC~Z�+�Z�3_��4a7�w�)��]ww_A��£�3|K��h%`�gTog��~����ή���M������G��4��4}�b5��`�=^�T�[FQ����Ԍ?8EO�g��М��(�R�����1Ɋ�q�]��b���a�}�f���`�d^<]�xl��RN�us|�m�+��������Ӆ}ܻQ�v�Tp�4;Lț�)6�(��bsK? Mh�`�qP�ݺ)%۝S"N5ׅ��~��Wd�*tZ�	��Z9�[�\��t�b��,8�|�k��v�P�e�ťh����⋊�=ۮ~�aQ͛�()U�=�=�gԐ�py;;*~b[r���epB��o��Sw�<O�l���d�%L�\���	a[H�'���'���hSB�]$��C�L�k��>�����
}������pd)Զ���()�R4��7P�n6�I�G�`N$Hڗ��GQY���U?��8[��1qA��@u}xǼ6����M����Ix\�heD����r��y2<�kH3M�D^�|Dj�l�1 ���_��M0n`�Cu���E��B|�]n�X��W�t�
[eӀ�rY�=����v� |����φ�徔f��*�u
F��u�a	12S���V�E{�t �Iv������&$w�>1�v3�8B�pݫ!Ռ�yr}�a|Iu��!Skq�(|/OZa\�D���_�wM�m�:0T,�5����`n�ͭ\�Iv�*�UwE������t����	w��@${[�C�m����Ŭ�	O���uyNS�N��J�uRp*`��)���tL���J�d��%�����Pq��{HX��Sɫ1Ҩ���I>�lZ�D!�]�(��":扁����Zt�b��+��˥v{װ�$T]B��n0�b��h�c��)�fˈ�\k�CY2�"d5k������l�sWI�"I�JJ�}$�M�S�����ߋ��c�WW�>r�
F�Xz�.��
�`���uK����S^V
��-�� ����IB��akx�~}����M��W�p��{�O��8�6��J)~X ����y����5�u�^�5��@������� @�I���)���`�����]��癌US���j[e�dc�x���eUt��Ŋ��f
�c���M
k�6��B:�eΌ�;��y^	����#m"��|4�\��z��u\7���;�^��<�P�L�2:��O)�XO�Ӓ��j(�F,��'�y�Q\q��`L��ö����<
Jа�Ҿ�y^-��"Exm'�~Q�h��e���wW5}DܫF.�,�W�j�
-��Uf�q�w�!T���J]�����]#�V�I�������B2�-ż�&�s����*i�FR�WZ��K[�1�����c�gq�<��_�4�����8���C��LRI-�dS�2��`:���]; ֑z{x�c�Qg�y z���j&1$uC���D�o�%J�	BQ��ҟ��y[��jC7�ɧ}�WJ�^669/���'��$!6�ׅ�TX��ƲDߗ��j��k�	,q{JI%�h�()@E��^����|ެN#���%��>��i\��������-Bį���<�����le9N>�e(�C#���МGwV��t@w�A��/l��U��nALQ��_+�k���E3��"�0������<n�EB7�J��<#�6Zr���SE|��)`������*�;e��>ל���H�T��a��l�W�6z��Sq`�8�� ��j������&[]_+����f2\��@�����Ս?�ˉ嚢W͈�)ƘZ��k3�c ��ga����8���J�sS#�����)�z< ��>��mOc߁��`�GM5�`�?��'�m_>$H��$Tw�k#1M��r��C#�h6�fR��@�U�,i,���NXɂG���\���]�M�j�@o6��R.���W7w�8Qp�B����V°^F׸
�����c�����P-X���n��/0���g�b��]�غ��>���m�2w �3$����H,�K�&*mϾ����6D�M��Q\�{��͡�M��.j��ډ94��qA!$g�j�[/(C���C�r-�f%�\z���yN�t=�u�`�*i���)��$v�����ީ��0-��#J]�~\6mW|�Yr��|���'(�V! >~z0wa�jY�v�r�u"�5��d?��vF��c>F��O�!d�#�#�>�-�P�Qkl�����dl��s�N`���B)xcY�`9#9 �>7�!!Kl�v�����Gk�0Я�ֽn�D�9{�?[$jA��6��~��԰��?K�|�ČJ�s���ْ~��u�>��\�ѺR�A
��6\��V�j2�2�����M���{+�q��}��e��X�u:sΦV���υ�b�k]-�����K�S�0��vaI#�P�̖���L�����G%��m�np���X���CE%Qcj}byX8f\�T��h�?R�^8�V��,4Ge�o��0����yFJ�,u�M���-��{e!�!�2��#1j���+F�>޽qpJXx��n�e'j̸

w>���T��P�{
��b^������\�,2M5���2s�����_bn��,�m�6���� p�G�>C� �C�T���!Ϲ9R2j.
�9�\��P4�0��S�V���7�&%��B^�:�[ÀL-rZ�=!ؕ~UJ�?QR|�T�� �c�]�j¥*[�ڛ�>2Ea�X��n]�&5��ӓhg^�JZ4c�|՞撛Eq��J�W�V�~ib7Yl4�ױV֨Q6ώ���tA�H� H�������$wN� /U�A�_�t%n�u��eN1�BN�ŉ���ݖ���H�Ͼ�z�90�Xz�N|�n��|�R!ӓsC��퓍wh�%��� |#���O���Vy�Ӗ�DO���*N:� ��{.�݂ D�m�+q����iPU�q7�T���aB��L �Y`Do��Q�&U��m�D�k'e�;�ʧY��r��`�:����1��a�J����nO��V/3A���|�7LF���~��{��j��a(Q�gu����9��|�*U@�m���-����%����Z�vZ��7w�,��ze�;�%a�(�Zٝ$�ԁT���p���=������� �ej	_u����O�>
\�l`ܲ"��N��r~��7��@��	ʨs� �[<x����G��%�"ҩ�2���c� �����ؖ��Ȥ&���n̑Ρ�۬nˈպosK�J��C)z\�f�6AC0�2o���C ]?ZR�wׂ�M�d�.�2��?�^�����.��DO���%�r2�(�ST>#R�GZ�#�Q���p?��odym	��jgw���j:~�����w�oֶȒq�.�����ßM�\�-='�pcV�����s����)9����ӯ|��UFB�f�6>��љ����W�)]�>�S�ǵ��GOql<S���F_\�-:.f��(kE7�0v1�[0�"���Y$@�y'^�u�DٙE��c��H�����"��n�6���1C�I��y�Bʹ�
u�]�c8%l5}�S2y�ƙ��OrB��lf排`�-���n�'XU�::�=W�|�B����.����f�c1�����`Y[�T�il{�ԕ,XQ� Y�U@��9q��}_���x*-�9��~ҏ�ֳǴb�ZI\\�p�����l��~b�<�
�����w=��� &#�o"y��	��/&�i)�}���)N3�8��#1�Ni��3t[�1�bK����^�,�C�?���c_:��a�  �����	�,�M6�i���g��˅����r��J�#��xKwq����~�y�F�@���� -J�7lRA㖶�@D@�N/�sC�I��������恆F�R������C"�����n���X6�2�f��5\Z�}֊)ؑq6iƉ�9g8����H+�a��M�Q_���ON�D#�91��:�Q��L�%�Fy��i�j'�|+r
p�R���Y� �������>�YUr����~��A{����-����014F[�������ϭ����(@(��5�Ǉ�t���j�Y1!�>��~���ݿ�Ǳu[��F������AuJ6��ck-^���I;�M�w��D!$
rɕ�tۺ-f(�Xk�
��������ThL�X~s�b�`@�kq��\$J_�Hy&�l�bꨧ�q wb�;L�\&�%�ܝ�
V|��r�3}ȭ�����JRL�ě���,e[���Yfe������Eo�,�n�sR�I&c��z̘���ϖz��p��l����1';�df�c��J�;�M��Y��v0�������0�:pa�*���m��Ȭ�c48�K8�#V��q�+Q��`n#8��[x�Jl�!B�>K={u���<{dPb$�1��Vw��jI��d�{��)��&A �Wb�z�s&K[l�
�SH&^	�e�w��J�U7p��W�%%� ���'_���Ɓ��pSk�ۍ$C����F�*�P)���^y:K��@�e��K_�\�"�{s�Š,mn� ��*�<7���0C]��l���yB�(�|gg��C�>?�����a�S�_����,�â����Z{�k�񔋨|4m�/�7!��=ύ�4��4Ta#<V���}M��wq��Cq�ġo�Y�:�E��XRA��r5�:n 7�]�¿��VO��u��܄.����(��<�'C-�P���yX*�Z�V�S^6�Q��`�0��5��i�{J�d�Y���7�Z�WW�E�h���̽&q���k_*��yi��_=6��.�wq���2 p˽����!���b�S� ��no�h�R=|,�˜^{]��ݯC{���� n���ǣ�W!.�8Y!$��@��J��PV�۽:���Z�|O��u�.�3vR�S:���Y�gPb�,'����;c�Y�X�I|ɃȚL���<
Y�W��&���@�g���8 ��$6 m�#�x>���M�n}1��_I���q�TwD�֦���Y��|��QOFR��8ĺ
)�[��D,���o��؞�TU�V䀩���[ߒ���n�޸PI*���58'Ɖ�l���D/��l%���Z�[Zv�I�τ�\ɾre���XofʁuZ�NzK�6�-K~e3���b$���ۖKA�L�qZ����C�ՕRƹ�LmX}�Ag�K�!=*�z)J�ZH��a�r)$�lMT;�Ȏ,qz�ȝU'�i��3	���h嶈����"O���T俲��Զx����J�:ғo��хljAB��O>BJd�2�iT��)S�~M���:���;|��T�>c�Lr��ǲ��	d����c�+�;ڙu���xҿm��a���pM��a�Z�Ĝ�[�6��NM�j����=ʲ����.�'%�����X�9����Ъ�@$-���*��1K�pi:NS�.ԥ��-cXk��/�a��J� E[ٯς��H��c�zz��?Ё��ၯ��#'L,���?���ɬ7���w	�4�T��v�|��T��R����^��s�Gίl)�R����)��p:G��z�
v�����(�c�f�5�P�Qv���,.��m�Nu�ۗ����?��ҋ��Dd���nW��E��P���H�
߅�Z��9<�'6�M�/4�+�Q=�]Y�Qd�۵~���!��й>�Cޘ���b�65�4���팊݅����
�Aݫ��/��u��O�7�Ц��8�c�F��#cz]�l[d���H�"�(�}5-9M���w`S~���%"FrO�:���}�ǡd����^AM���fUC��93pa+ݐP58�U#����$ ��"F�q#z�?i��iC�k�6'D�'D2Mo)��u,�D�������iZ#=�I!�h�BwL!����Ld������R��E��.�_
����^�YX�����^�W�=��b�>�TF����0
��a���s���\+�/# ���������uB�x����wЭ��V����t��c�łaa����X� �H` �`D�+J)kz"���_����j��m�Cl�\��rÿ�ND�b������C��?g��]V%�A�r0�� ᘁ�����߷���IL�K��Z��niUL�y[��J��><���h��Y���<�5��T�T�ڤĹ�T�P�ں߸i>��t�Q~t5�D����:�SWɜ�B�X�)U��"�ܶ���w{�i�����.�)�r�Z8��Rk� G}Y^�ADZD� ��2Q�"���Dq�*2Hngj8�w~��@<x9�B�w�Qw���]E��	�Co���n�	��ԍ�}��(�����T
�|�kGºxnp�Λ&�~]ZZ���#��ٰ�iSpni��h8�xSi���gzl��-�ᝧdheͮk^����cQZ�+��-��?����	�v|'g�Y�������V�Z��Y�a>�����qn�M��y�*��9r*@�<�N�"T/\j���I<�G���C9 �g3h�v|Y�C��$,C`��n]�Mx�C(��$E]#l�I�5�O�r�A�� k��QVO�b�t�Yt_���3 B���k���TgJ�ƴ��|����7�f\.B�Z��G���fOe�����佩�n�84H��G�8Un`�-��7��А�O��8�l�N�vV�@N0O҄��+٘��t��N_��:s�ƞ�9[zx����ɘ���-������)�|�m&��Hj��G18p���D��T
�_5r�lk�ǽo��_�T��]�i�Ph )��łg$�:
�kS����e�U��i	6�>�X���0��޸׎�~��ƕ�+j@=�^�7UI�%||�Ȅ��g/����*��M��74��ُ�]y�^`y4g��]*~�N�.��e
�D�1;Ϫ����v�
o?,��V�o���(���`?~/Е�H�O�G���nZ.	ݻ*(r%�E��Ekm����UfH��ݱe3u,��kI���J'k.���O-]�F��ў@�U����0�kZu�>���z]��L�*Ma�9����C��\�Mo�v3��'^�lXD��$�������v�8��_���:vގ��b^�IH�?�n[ �2q�b���B"�S��Q0��H��f��Q������]�ٰ6Ww5��@�eW�8e����6�r,}���ȕ�G�r�2��8Y#�4cdú�QR�����U��i`���	�0��N��od�)��;4+�V�e��h�1T��T�&�Q���,�&�j]�0/o�-~\���
����W\���]~*�����S�/,�/�z������<qL�Ь�I�,�[B��]n	��l��D'����M6���3�C�����0�Z�4��g+������&<���$o)����Ix$`6ǋ,M�	�X�7T�\{ﳘr�O��A�4"K��J�쭓�
9s袬��k�j�*VP�z3�@$����?�u�ێ{�j�^�x�Nf�^V�/2�:N"�_/�$Q1ݧc��i��.����Ey��lP�\� +?��:#�����Kz9�g��W�C���_��rW�:�3)��.���@%�Hr�3D���	�:;<�m�z�_�����h�$G>o����j�-�n��}?G��4KN�^�Qnu�f�S'g���#z��;�#4O���j ��z�y����I����iQC�KI�q|��SQ�"Q��aT�+��8\R����3�5e i9`��z�.���<+n����ϙ��6�L������_L2:y,q|R�o�H� $��2��N�G��#�^�5qS�(��Sf�`ӊ�z��'��,�|-V��F�;�?�1>{jn�j
���vD����Ŵ���'6��1Y��cy��]6�gЬ���a(�%�%���#�~�"B^Z���:�`䯞�������ilՒͱ6�
��~�-�2~���E�Hߠ�:�6�p��j	U��4��jW���
�<�&���<�� F� ��C��0�[��a�rǎ��,������W��ԏ��P���q5�*	�ƏJ��%��G��ȾL@4�ǸM�:��A��M�C�$6����`�E�'lOo�D���o���:�mbg�b14/�~
��8�$����ZC��<�}�kMYp�4�bΛ�W���VR���t}���׳b����l6hZu'|�X�������(8��1�[� �pV';dF ��ƀn�c�R��RO*մ��}Y kB{�����d=�G���gBQ�ы'Gq���W�t�L���6���"���(��)�Q�9��R��)S����֒%RHC9O��F��7@�Z'���m���J�Ν���F�8�OTT�k1'�*�`9yjn��n��o����w0�8�%��!O&��\;M�W��G|TF
��C������Y����XC������wj�{��\W�����z4��w]��}{̡��g����	MKj䱂��KFm��Xo�E����ҥW��CqՍ�s���?}��{��S�5�$<�4>����k�/��/q�4u($�oG�s�z�(;S��,Df=��T���K��>P�go�Dx���d�E<	զ8�E��eH�����Mu���;a�Y��^z@�E��zL��nҸ|p�ֶ�	`����%F��S��ؗVK���	q5��'�t����yz����(�-�F'�hk:��$�t�oP�-�qM��rQ��-�[1�����_~`�K�#�~���4';����V����.�����
�����R%��i��ᆏa�L�\�:��{�Nj1��&�5�ŕ���	y7,�u���h�S�PF�Cv4���H��������e�*F���f}���/esJ��Tiv(=]���8T�9x)h�1��ˊ�_n:�hYΞ&�;��PB(�|��0b��3F�hK7��!�;Uk�|��G���f�i�I�~C�s;�h!>�n���~�����#���
u��s��iS1�q�`���_����J����j��L��
6p�ȶ���Q��$t�MV�1���β��_�=�YA|/�L��0z�>��iڷ�.@̃U!ތ~ ��V��xK��>]=�wk*"����*��:����T�uO����WٷGve~�9���C�g}]�c%�m��X5)��{���3�k�oݡ�Y.��Ғ���J�;-lts���y��Y6�U۴V�yo�9nWU������u�dܠQ�E��RR�@+���ԭb'�M��R�[��<�h�r����6�����jsZgkg)*���klc��4���G,i�mp��>k��I�n9�z�:_D��:�ܖܺy�Wcb���b3�.s��ci�SKQs��Lf1�Թ3�}��y�[p~�_���G�{�H0�6&�˩.s4Ft� �{v(�#V�|��G<>�1��L^QR�7Q����C�+�S/�V1'�Ӫy�=k������:�Lp7�ǖ{����3����fS��r�^-��w��-oӦ�)�+�A��Bz{�����P�{����yT