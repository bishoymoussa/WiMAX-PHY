-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
1ntj0IUVb7HYukw17bDHa+E8fXc5cAENcqsz/9BC+cCISSUepeSCdFIHKhYa42UcY2pESt8wpt4N
KzPMtanxZ/9Pvn3obCcl2wj9JPm8D3Q+nYpCQMqPv4NJll91i4LU/iV0dOT6ocyRdeFVimHPuP3b
3E3JZgLXQH29hH4GhU4kt6aDs2kVC82/7gNW4aOIdCzV1bETNAGstxmJ7N+z0NvUaiUxqrvF/2Ff
nJ0dp0KKHTDgCD/eq1HVZDWpXOieXadO1Sq2ctyTj+T4SY3br0VCN2F8PY4LzktW7IVz4Pn5JJnV
7jjc7we0iKWVXNLjrr6c81i7yaOr9Mgx3X3wEg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 114656)
`protect data_block
yZxtTheKgGvC+37HefaL4mw62Q2u0XHWOWnrQjqwl/YdyJCLlYQGIMqmAcRtBtkU/MdKVJ0DVXw5
WgZMfQzG+VoMLvOb6zOpJQsOxoHB8c4Ll78ujZCiiYOwDepGCL12+rw4ncDHEGI3cCotjJNSRFN/
kOJM9UoqqYoITwyhh7+lHvMuF5mzpgzpJ34yan5kNMgn2F6MQf2bFt40ImFsRRtNMGKSkClwMTIN
06lAsq8K4BHvXFc9O8Cw769lkt8OfbtUR1nljQhPsEXu95Vw0Bxqhxim2zfPHNISfz6Yse3KW/Eb
XJth1etm879It7DL+tlQo22JOrvDqXBkmPQ60tByPFKkqHNBLfIQPe2uzDMAFTaocE/KysbNLoVW
V/x5b7ePjZ2N1IfiwbEyFrDbLewk2EcVbFZ+geRmUyrzNUHqB+g9QZ3z46NXCuA4bneyXw+UPI/s
kgDWt/nloNMXrRj/kos8+8BcrC1CxMm3Msy5c9cAUZq2lZkz1HwaQoFsY/4esFaG8LP5PpO7jGFL
Q2fxQFBXpIbdLk+QY09LqXi3hujsOej92TQBbsJe2Roga4sPLNIGEtJr7a9BxisT/bPJ+0sR4VyQ
PIqK5wBEhbWOCB08IAPGKeSdyYPY5zWYq4P2ZgdWwMa1IcPMy0lID010g2GvE9c7KqKKGjjz/kDe
aw9IaNAqqo+e/2+7G/dBE44JI0vyFBzx/KPiyw75wvwBkil01+DKjmLGpmTkrMIZj6cpYKLYs7Dm
Nka2O9ocCgqYNGh6lqdBhwZZVWBTqV0JEoiokxWUTaS8fhJ+yDoNkmxtfl1fVaAL1V42yGaoHOOd
vc0U8etve0Sl0CP5xBG9QgQ4rkPRFkr6HApbe66xzw0DDjNJSg2ikpN3dydrQrU0j0aGmmYO9F+R
tb/Zg2sRBmdAQRJ6BAWAge4bqtIDWMeSccbfI99t1H0mGlymT/Wzk5wSCBCX2KvsjpUdGMdkAd4z
tIvJnUpsWrrp3cXz0fzkOlMH59f7Acj40YdNfvOP99Ydfx+ZaQhR8ef+gOcF/RxgUaCijvUKR6J7
cXKwCAc5YIVKbaK7GGzf/3NWRne4DU8pS1TjtJe9ZAxcN+O/pFtuCjC4gHDuX4StMrRwR9KKkwIx
PRfie4EBK2ah4OfJMqDVP7iDIa/HVJvtYuKKl8GPYYLegbRJ11BChpPiTREks0fHWBdr5/YUe9Lm
9P5sTjvLf27EudIRnx1TMIyWFITUctWixb/qNzeQwrRDi8UV/7gODye4XiWDBRX69DM0DZhD7pDU
gQLRPl+fpGiq7oPpYkOmfvCxeV11808Rje9ulKSg89vReZwy6OpqDLp5fJdmA+JizB02aXcZ086M
Br3tTHiYivInCh6g4PgBVHPUjFDNZtbY767+tJalzEF/K2I+7eMQjZ97zByjtBRFlBmjtDZ015Sz
/fO9TpZjuBPufh+AtI7vdwfiXAdXaE6AR2sjaI7dq88khR0kD3soXLgG13W9kbq2m83J1wnuAxyg
Yaei4MjSAy3Nowf/HlQRsn+8m84hnv9yjqrvW88C3/LRirdFez83HPKSPFsq4W6vfw3Z5Qm54oaC
qi9YCHlsSgC6ZMCYI9X0NY+lcujRhQEu+TAmRohoOhIEvBR48ybpEACpIhXw+9Ye0G19UVc7ok71
3+euLMwkX6UqZQeDkBgJ4VtlHws0aJEaRZGctD+dn8vDwNOd2C02fiDWxxxRyeL1zySewL7M94zn
AStAxdGQH+XnCnRQTxyxgDNk00yI3hV46WOtcuEfd7QzJWSHAx3EkCjqboAZnXvhs3Fg62Zjm9mX
P2PQ7Gx9H4cwWAeUgGtFoZ6UJaxtR897/Tif4nre/HTerjVC3Q5C49DUTjqwz6nxVixWPh1q6Acw
WAwtMJScWBbS0NAX+hTZUSkM0swrgLPEQKZ/TnBUCFGQWHPJmXf4d/3PsZDeGp0f6z/Z8VNumqIr
0/GqWe5UkC/Na7Kucjp1w7D7hs1upyOhL9j1lpbu7HVpdHerNwePehLgr4xDlhrJgVi7yj1zFo5U
iR3g4T80r5s8po9slnRQl237VMqtGhVC5HIlqLsFcafGcwyOc8KeTbv7BvzT4h0RJEOoadziOTYZ
IKaHGxcFN/+NzLVACL00xCCdtyb+uxE/1irMPd7PNdSt1aecBk2EDCClQ2N6pMqKDnaCvverklxt
mJ8GJ7VRYcEG4zOPU+3Z5WRnOHcoiLQdyDjz2GqjQ9RqIAQp04BuYdNS0vKT6/D1L7XxXz/TRjoj
YFaPkwWBTWO1REKgWD5EVF/LiQEnQDzgMifhnMwbO8Qf+0TScqOgBghUJf0ZuOvpgqZQOz0XTVfi
NjnYawnVfHg2JisP3ge6ODOjEeO9nJ1pk+UvyqUkciMlKNnBqL34Ud+gm4gwQ+5sL58MNT5Hw1te
nIIa49wVKCVnL3pSSsLafh0U0zdq/J7irjTAvKrsUQe0CHIzcceFYRn6okrm7hp+cBw9VrwMf3gj
JoF0L/Ml/vF9C3DU6Lf8O2YoHGOedZkgHFHcA1vgdGudnmBVPIMR1zK29MBRjMEyFEVYyZ1SZm6j
Psz0g0upuN/SbPzit6Vl9V/ZSR6VO/jZtvT6xYDTxbXwCRZftEAqNwpVpLYu14qUA3fn+Ty9Iu4c
fTnCwSemAa0LKjZuAfrr+QPZALo6BS0wfo2sm2l/h0vXHuhPWvmKA8NppPjgzRVSfmV8HZVcIm1p
Pxb2K5OllaHqZr3jET0g1IJ8tvA5Vn4EJj/sxhuVwbE+wzqsXwMbDo3k8H15naWJmYjrOlFuC1SO
TkMCswveAj4v7tEmqGoblY86G+8g3VCn+FwMNKIob97qMerMouG6JU6lhR3sY68Fkk8TWW4hcUSQ
+L4cIkdXojZer1TRQpbYzyu4bEth47TueTWWlR2lbl4ARDhRFqf/0hSfNNJRmd64fbzCQMqHt6UZ
hcQ1k6FFNTYTt19agTmYm5ToDBSc1skldlXTvVhf+m4/UrQ3dQEwKZ1Zhunk3GQiZOeVlUIGh3lh
5gZ4LkcbJ5slV45bsJT52Y5O+cssrkgKUyPZbPsQAoVDnEJjnZU6eeNNMi6gW6fvLysEepGVY582
bf60LBl7+nsXm2KJ939YBfyWUYUI73h6G8mOSNe243be4yqxF2nzglq8gv+l3z4vLIg3FTsEEz4F
SF1fcSLUUDLNVLaTvRQlFG7HmS2vbpJUqdiphUdXW6vtH5v13wVyFGSBVZn8znkOvpXF+bzhSC3Q
XLdqibnzG8jzRdIBL3HT7b16um4kICKejkp6F+11IRR1NeMD0PqEbeDezyfZKpjFkCJBcBOz9WvM
kPurB6OeqcDQ7tgx1ikDq6Dr57XF6PUxXHE5c75w/MYIpSUz5d/Rft7PJ96kJGWwGjw5kMlutgTr
gZntxTO3g1AYx9+Up4dfOdxj7BADGHB3bVYNP1MNBpII+Fih4rEy559rSCHEHMOopPHPVquBbVOk
kXeBQ57MzLJIECXGGHqYEBCLJ/D5YZFHYk5j/mn0gMaiBn07RVLp4VEDGqYtluMv+nYtuWTywP+/
mrAPx10KEzXjn+7cAF6wsigNqLvsheMyalppUTrZJubmqSLVyzNaAnWftvBPPpc/5uyL8OcNOiEn
cSWvUpjgyzwKNFFwx8dh5R8M/cGr/QBmifs3K/3nO5JwCCmMdIdA10d4333pfvJsiye77pyf7EKY
TBAlKlyp2mGtH9EnEMALNekNvjn/nHfBNsRYq+a47IOJ6ZKUGJhpR4RCZ0+e1QWsZEr31K8G+lQy
W5PgqJersIU9U4+dgnTMPHLCn+BMKIk3VMypu6aLObYyH4q7SuL25acowKlKZ1QLTAr1egENAXG0
RP/awDvZ49TvJMskU1xCpzZAbhwv3fCN1BnkBwyG6oEIJwbL5e/hpOAqOVQNlqB4VppMsOJ09f+Z
LG4hjJ8JOTeDV0dzLxo1U9Gd0XXBw7yRF3rhD+NMC90x2ZFnG8wOkYTfNHpBahQdoExPpLjCe6ok
67L92846FkTIJVeiHI3HJaS4McaYM4Iib/aSiFSXLwkLWZAKwmyoCDO2vmC1OmVegCrTasfPzvzw
Fqekupnv2hRnQqjgaklQ9K73QWMVIWP8L+1op2lGHm5fvSOc3VUxcKi7Uuw1cz7Yk5V0FCsa0RTm
/L4Ns02Th5TvljRAnouxdvqyJRfVC6wMqXaJQvf5Dh41SpVw0dwTReBplcPlw19/X151MB/2XI70
7JtVSQo0Y1gM+h2QEUDyqOC1Gj84IKoQwDDr26/tGn8zOEktyrXDSZnzW6q0NZ0yb4thvtsDpgY7
3bTn5csewmQ0+/zWcPUZyeP0F4LBAcN70WSKupVepygtBOss2EhzuWWmqkOq3scjQfVLbWewEypC
v9bG2rLYvPYCTnaK9PaHz0mIhA11PFRCmTEwWuk+NM8uia4GIedYQu2UCN0Jz6H0wBVh6FWcq1Lf
VZiIzPk7MuzFWT/ejgs2x2JWLngEd6I/96DxtnGLMXCYAaB53lu0p5bSWrjH0Ba6FY6bOyTF1OjK
zwH+G9UaGk+IIU2rAaR0MPnaTveviqjpZG9Ht/sz1Z8vqnYwHMIwc5zSHcLjZm3EtTizWE0AJGYQ
NDY4Pghm+hWzhGWgleuB/KTmap5CREChwKShylc0w3k5n1+F0lM9ZNr7G5aEj6iXWjfiyUF73Iw3
gPASlJ3R3t0LZzvJHKIrSvNZET8GmcSxAlKglsm6fKW5e86Q8IiBjiG1jW/Q6x4ILWiSYdSiRLq8
eP+LwzX1JtipCCwJb2IJ6QMFZa55H1NzYJq3soCLMftlwxOZzJtwe6ge2MXErocnCbmJgCK5wsPJ
GPr6ltDMoLUOm4SLhXIVdk1CdL9RlukYn/4oWBrnsjCMOSPIq14EnMl0V8k2ywopC0WX7huGDLbl
Q16U6qBqqGxoDmdgSyJbm0RJV2qJXKyBXuzJzMDtjQ3U8ki0BfPoONMHfusiqgZ0d5yP+G9E8v6z
i9MPOKHX2ytD8ECMs09G0oti8owPxc2tSgawes7Lxy3vVnmrB2q11w0UTbCLRgErBhFIlU4oZifk
Y0+HRpYKnBveI/E5nJom3j+g9b8oO/MHK4inelCQLXwBCTLa4UyiFotVuxuLjoRgY3hHneJWRp7t
RXx1zy1JqA9NOswUPoqCJukzprqFDx3GebK4xpNkwmy99C0tsnn1C/u0R/+tniSNJyMeUY/ragyo
pXpd3qUYFkQrxSxbLXkb7I2ZLpGj8AagIIykObRaZ9ApUOwifUooMs78atNzVh2yADVCpri+/eW7
bYOKvcsmy+A/u9j/yk1lNK7BBR/AWbaRzj8wWBJ9isUiFqKVN4oqVe3vSkZYkAI0+BWTa9ZjJGCb
tK/S+S1gMNdEDIaqV9xQ8oWErHzqfegAOYHb5jp9KTXEXVTlM3r/LsSsCgHeXx0pO93KP0LToyKl
M6h//mRIsnpJMPivlvQ/v4jGm0Dgevj8Vg9Jp8bz23SW/iU8pgchgVB43MXv4jEGbwGjkW11C18p
l2MKYNaKdM2bUFUKVLLsEi66vJQfx9vvUZuaUNK4Z3v1tHWcs6dQZjOzfxR3emBh1C32EUXSwMcB
9IOGgXn82Y7dNSYy+wZhzApO7LGCgUQidRSrzPfq+2kvBvqb8lILWiA+X6DUDCevo4F0SHM7AZbR
YsMrrTih+5hRica8DvLq23IdJVLfNhAd0UTHsR56cJWqaQfOMyCxUVmY3viwz+60Itq5zirl1U3X
buaSO1Ap6w7R7WHZ1hlvOMvbmeFJptO9ND6zvJr4I7JJp0ILFFQIHA+6j/SFNdZtsdvN4cngGaMA
KOvUaApWzy8Og22Q0v3inhiiEjLQzO5fCOP29Y0H05NDxY+inIJcC7psywxlof0cXUyRszKpXo0W
icf4/JGjUbX2HrVeXyaKPjPe08ughUvkyO2bIPuMRYLwfpK9eeW3hxaxWegOblX/0gpy3Z2crelh
qz0OIix2pUl1CKBK77YG4dioX4LvlmvczKsAzen78sv1idCbmcRB5dbdMggkxsgZYysHC/XVKVFc
Tku8ALOBCN2rjftFsy/LmkdCQORpxiferePqDwXtfOBMtm2L2I306ZIu1VGJk/066x7nnfVyIISo
gNENBZwP1D2P8aYalQR4f2HHzwQQ0pIg/VjdPSYJymHMxVC8Z8Vp9k/vnph8OjoMAvYkOnaoZVR8
0+cSyPVTrIIBF2jyW4Gr3bkb2is6AFEZE0rsBF0JgNLA9zRSfIJaDM8iYFTbXPKpz/4ePOFywc1N
kbhwtTYKj4/z02lnlVdrp8O1qDpQMV/8CC2V25xYS7FVPLFVpV5wb2yAkBwgn1VGKkVE7a+6hTAM
sydyYSGrIUli5gurdSdXsnzPT/aJ6nTqWAO34xvBiWFutl3efIrC+WnJTWSD9fAOStsEk2TrGmNt
5zfc8Kt0d9dU+tPhos55LEPPk/fg5+FgGJfuW2vFFf7e5zcw8OczxiAiVhmMJSdg+YmRHshMzImN
or0LRPIqSIJb0n3ut7agwv1JxYE26rndUj+9hhTRQcElBedQ05DMeZ+LcPP6/i4nozSIfNWClK2e
93SIIUwI2cUg0iZ/iNopbtm2z3zxSSg5vPfdsibGhOSShG9L0eWVvb/zRd2ZFG9uYXiofpHRQpwf
wMMExCbR61gOhbCCiWYbFKSNGGrdwQFc/Xd+uX5X3N7g3oX0PJrTGVTRwBmdmNf9swEZnA8TrWLB
6C6r+6aiGRGDA8HkPuZ8zT+68got+UQzKTFvy8XFnz8WmteL/9iQ6vyNV9hrkIgK1cAsXY9kUHc/
NMFQs24NaRh/2YUyA4cNtWjRo9x/kfHsECaLcHWBsa/pmod/6oRtWJfYSZbq/zvBeOTFrBHp4M1Z
PkN/zGgSY4UVMtII8qPmlPwZ+irKSHwfXGvUQUQKxyNfiAlsWbyHaNxdVI4jkMRhtZMjXDM/J5Ep
b1nIYg/dLffWv3hO1IYxMJ4UbForlb8CjYwwE1nVJqrapWfLoE6T9oj3DffkJMF3l/kD9vFDgnor
37Gt9vNRcmkNJwUbeOsqd3SFdw86dWbSJ1q8lyW83uNhkreLbb+iTdJRoUaSRdntlZkPL0GAnDjc
rYm+61xa58fhuIpL8OZgQJBEepCTc81eGZ6E+Oxb5jwecwryXEM/U4RVUihzDLNiDWidgxt/+//s
TX9tg+zFHMugjJJu8QsOsQP1+8h46Izkk8NuIEvX+xcyIYBBvTGvRneuYGbRK1cI4Qc8aGFRg84b
inUWQ7jeDxgUHn0CftlL0wZhacoNihFHaE4H4dh6FjHVrxLAo48I0jdAh9iSfnKeWN/Olz6S7zQI
haxtPC6GSuEzUeX/TTmx4MTXs5G6H8Yew0oXlqjiwah1r7k0XUW1OhiGz/KpDX2jZfBucAxTJlgu
gSBh+Rz+WVkGzB/C7or1wSYRWUvgvJ9+Tc90rdTIEev1X+XgBuclLjcJ8oW9kd6PQPn8YY8VhuuU
LG9Lmsn/6bLWEPnzmE7MrdMAvvLM2GsXXykUBNCpJDcMmK+Qo5fso0QafwvXxwTopnFl4YeyXrDI
PtsLosEUiEP6JdGzjy77udHym9d/qVwhpWUZ2MNlDrrUvWUO2SEUsD0WKlGhht4o207fco8Q56G7
JXxTBFekn2+PchpN2fX8MezOnY/Q9zPuR9yW549tUwppKbvduk21Ll92gff59YkbeL7VgTio0rZS
g9yyOl3HfqswBcdlGns5g6ueMChqIKh8wSZh6ToNoX7qEhkI9BvuZ+PhMKWcFWMX5ODbq3wZ0YCG
IFHHPfjn3pAuvfBbd+11B0pgAjaIhnLLICX249e5O5EVPabJI6DAZ40t4D7gLjGyTz8g7RsM+hS9
6wUoVKPFsmi6OF3Bn7bE47p/BczBezVaJ/r9cLfJn1IlqnK2L90Gkxysx0kdViBwxJd1Z94OM67w
34BGxz2LMpJZQ1nuD22TlTTh5Slhz0THsizN0ZnWIAgutbhVIHzy5+NkXjmtnRNudU0EnWN/rdX/
rbaOON+FMmXXTbdjshxwK44udfNT7fDxrYj2z8B1TU1JqFNff0zzow5TBlUBVfCBr2Rc6rwePTJG
z2zCfEqfL2kCRCmBfVPRfzBLOZ1b/H/bgnLFkzDRdJPG2tY8Dl3QGFFXRLPsOGp9F9w3afbTcgRI
6ohHjApl7E+BjqesLeooslMdK1bseAHsXonpA0B5ZRbTIxAryH6jaJB+2rfC9NcOhfXks2x0yE6L
m4G5IRg710nLLHL8hogeZAWMY/kyHh0SSIXW9UMxzfOW3gKrXAoAi3c5wwAcoNGt6uzwN6/G1oPG
vI9tIvLdut/lEaMs/jCP3s9GGkbiQmnuP/Nkm9STQq4SGPi2pYFFstDitk/Xf64LNFNQvD0MAq5M
X5ybZ/SAOox1aUnNPAiZ5qfNXueQpwNnsGageD4PTVMEz1W3OmBOee0Y7K2RMULtNY30gogfaU2q
KBnrKUax/47RSE7OWe3JI3pQarL7Ee3ha/8SOfHVsGLxECNAW5ualCXdGalbNT5EC+OiuTG7ZgVf
NzGQVVVSkNbRfR1k8Xyt8Dht6JOWlEqETeL5a7uYdsH1ewTWYG1a3dnIHOLrvNWdv9y+XaBv7Y5G
djjSqcLhYgtLbX/xgqoqPUhKtPc0KE/pPnr6y8+tNPgl5DDhb68rl7r1DYXG2ZWBVsJ/xbEtqGiV
KUNipJQwBRLVw1SsfjTlxSBtWHH5mtXYx3p6ewWOyVjuvEtG/TvMy/1FnsTetmEPw6e0NRazSr4U
GdkezAAwu9ei/vdkDpr9Ll+nMGySELs0OFb3d0pe+CCvUtR7UhImCkhJ3lSHEmJZwgHpaSf3WMIj
f8V2QGKk8EpSO8D2Dw4IIwr8Ie6IV8XH4/t6qlFtpFjEKpmN49/ihu1vhMGEmo5mKCO+QA7eu7ep
iVw6RXv0Hzb3CfDeFuqj0znBK3WoCtzZCjf6PU9rZGlOJQPlILtsNe711mgHxtKSDiRW+LM9Ivb7
hcqimqZTu155oQKiHKPNMG3pT+dLsYmhLL2lBbcuEN8pRTOeGIOgnmEX+0JEctZJHD/YEl6zsi0l
PN+KN55qwDvEz4nIwAeP/OhEKQh8ddCidp7UZaLNQke+gWSvHHrzdk3mrpK4wpuKlDCYeeY7Bl6h
9Ydb/DI3uJT2Rw523WrKJTeYCYCpgKrpIjkh52RUu+0+eW6BUhRqJ9BKdJyKF9Dbi5DWe5lcZnZB
0+N0WkE1VGL1whcRUGXALd4JZZSD/USMU7Qu+O+ps05fyi4hEaKXoZwLK47MzUuOpPj9yd1yDl4k
Dyx1RsPXjDUDP7BPyeJmLUYvGhnH150M2ee7LoMN0K/ykerDRJRFFHfXVvs1FIjDRPuJ4dg/GDLv
SZXE9mJec6xQJWnyb7MYHSqF4Th+kB37v0k+eyJaTcr+gbRjy5Xv2GXs1zTQVVbOdWwskYThjiUr
oGdt/lBLhdSaCkEAjTPzVnrIFN4m4HiOrAJ0MMRr/pvByaqebpRmmUx/PQw95cSSFxMJkAkL/TIg
oE++eynEBfbQvMH/fyYtGqgpLUKBcdSS2/Ixa58ku0DbmLiiGQby0P2dR/zqY+jtV2vcPlR+ucMn
jivmZJbUryzkiFSRaY8PKCDRz7SBbYh+LJ78TzCbwim0kvUHzhIFkFDhCBy6L5E2q/UfRAc7GqWz
dG/awYgBjaZnX9sPulPDn/F5bAXbccEiiV2YxMKyS48NqqDVKM5Dftf6lg9LLdiSaKHvvI+QO4wH
4+ISn1CbGykHRFt2elymYSGRn2I7XVmY40KaqdkwxDQkZ732ML6nhHAApAeXTtwznJnM11r7tshx
057IYI6pH+js6DRsPG0ZcUXVAIrjuZ3RfhUJjp0oJwIxxugOpqrsRT4LO5uybHuu1uJHBEh8er+g
MzHgPso8wsCvKsrPPxnQIqVubrfUny17ye8m0czM1AuhnM7a2ge/gXh0+WAI37XxDYnBq1vszN4y
7xwT/TrsQT6LODkHpgoJaaqO3fQ2Jm/lpBP5KBdUYQqn8L7qEccwq3lQPawKbplPXzrqO0EaWhIy
SnSH8sD3r9rgRsR/mp8Hh/bZyEeTusQmmx7X+Dl4mD24yr3/2iLiabi4iqy3fVU/T5cI5Y8a2lb6
9pipCFWetOElpZqeEJCLjaf2kpwDu2RA9zZou4kzFCl5E1iIUKLLDNs1hvzd4jMeMMxrM+VJx2lO
0voc7aD4CcyjssASWLY2cB0xhiIhBx6jJZU0XTl0rnoObmNvA2sxIkLxjt9KK9dLYTh0Mqa0UXa+
cUqWqWNNFAwL6i/ByziJB/cG0WVnqPEMRZgJqX9+2+S1UOa+KuyQKvPK8kotFCStIKYEO510IdiW
UI5yfBqwAxtEHwHdRkKDBe0Vbj4AcSzFxX9Cy0I1L9aqHe2zytU71s9IDyPl85bDxNrLrHImgy8i
bOKegL4L7YdUnbs7BUWpvv3trsA4EUIs+BghhfZxkzFjHJW5hp9V3c+mahRowPHwA5O7Z2MayZt1
SgDyEF18ylztMS/9B9Zpo3wvflmpT3wREYSWJ76xrp0pzLKcotQaM68yQ+ja7D4M58tQj7bfEO7G
Ly2Y6gqhqZxECt1RGBDb2yOHWeTfdeYp6mEmIlyePWRKFrNswYV3lIbxpkXeGicyWBo3PHgdT9pc
AIf+W4U2qglHfc8niKdRQP0IoeE+W4LSnGfnYcKRPCV7hAXQ4MK6TcKElmf78hRJZTBfrRXfDpNy
FH2NZy/wt6CaeQYIt2TfUAmtnLB3UpuVHehH2CSeWFLNpOgzVp9XXAoKp3OmOrbr9OeSDUxcx6U6
Ev+MvnNgxYqiWJ/wfEE3ECOqr0Q52MFLRvdUgmVDukFQ2geW+9krOWlO9Pqp0Ry4oP9asG0yt+OS
0QJFS9lcNhzvAgx67D7yWS+BQGWm7imr0la6zl8ZLhN5pTAGMownd722QNo3+AGSPgpd9iFHoSJ3
y8dmN3HEFAwNOWOtgAhywRU2bNVf5+6D+XOJ3gxV2hQzD56cxNQZ0f+hVVkprZhauYNEJAA0c7QV
sv1oKx8Pflw4eDVXWAD6DhY8XeSjCJJv3M7v2ZbX1vVOg0i5fo0l6/kOTDLF6D83Z93siiNKpg81
W0PONhwB8isANnOsXnurpaunQiSu6Ywm6QG5a5mPJ+kkV11KF//0raPVJ/IixPhgBBRXfyBK7L9W
5brv1aQDH9CEJxlbyjbGCorPIWjcQPXM6YP8bxtJLlOITdXroISmFnFaWUcmLly7lI0JOpmv7tFS
rcu55bfm1gS3UJF9PRAcUbFYFXxjWBDqqi71e/LeCH54HA707rU4RbQztmoT0qJBHeYY7U9ZehtO
rEY0sHIH145RFUTeiMxoNPndjApY1ZPcvCLGp1FLh+rJ12rPi1XOeuRPIUhJ6/Zl4Gb/Wycc+bmQ
0dRTe+euPSWoT6SmTaEkn/PrtvH+t7m4lXAqK09FfVn/inVY1Lt5PDprKXwXqAzfO2pv0+MPUNeK
3SORtY/+nnvWkxobslSui2EoP48cuajp3MUgzVE9dAIUZe7j7YZMf8Tw4xpmVq86IJgbLqLADK0s
IKyMXRw/Ox6eRdRhw1qzhgGNpcctieeJ7ImrA8WYn3NYJzZgIH3rDBz0cNxL2VGNeayoh+cnQFa7
Df3hxY0UfPyMLM07pn46iN/dcWh9BpyLbLA9GhfhyVNBh0h84UeshRTWQDrMsalyGjNXlrMKV1ap
jG9k7Gya0Y1JTPHyeeZjFBWwgwc33Jfm8rf7U4tOn8ipyjYnuASgNYGGWdKpKta86PbsXhSSSxVS
qlkxUXVXMOvJz0e1iZbJ7uxG/lqeRnF7Zfajcwxv+IP1o9c3uGbc1ZTNyJ3HVjlDuw+qT2+Qjj2g
oZrwFjn8D2/KymrMsmNlsDP+yOuexubuI1EBf33FMawcg23ex/zahIRYQb380ip+GNJGkljb7fnK
J7qEgSG+uGp6W/0h3LQjOSBppk6rc4lWj46+9lKJP5fvcDiYj6hzQ7BW/bKmvUdNGFBgm6pjuwXW
IlkadHIDEhUFTRiYfjIw6s4fIzOcZo6kkDfzMoq0w+vYrZOYB+6xSezENyadWtCofLNwZWnd0BAA
stIyIWsS6k6UguuAL7ZvGw5JgLUx50Go89QQXfI/AZAMYcQwMEPmHYOl28nh6ap2yJjZp6VGacqy
/exwlM2YyDXnzlTj75DrhzUTycMGTrN0MINCRh0eWFpWI9Khh/z3+Fb5LFDfNAFAWktmzom0/OpZ
GSASoVD9CfJ4C9+bGPhbRc4Ciqtbdg6mnG8Bzi0WXFnushluuOJ4Phb9jEbJ2sSVp1oQ5FP1sv2d
qepvLf/1swn/rYpOz78nXc4vZeaTCKGkcvaLAS55xxnOdr70EPOi16OJPc0Qul48RSB4ps5ucGsj
BJbheOlSBtxQzUmvP19uyR3SGtHwuez154eXNhUGLt0itJoQBuVJ9B55hMgkAcuCC3lhMD2pfUK+
EpN82MM0ch/b7fjySeSNWVaOfXEl27B1LcqRyvurxOFoiiqrFLloRo17x6oIeu9S8E1WqYQxh/jN
DXLXPQhV6ltusRUKPpaXP+Iuhu6MghX/1AxDgCdBMQZEQFhHNpNVU7IsTx455FL8gYf5F1HQpRCC
twaaAOlFtex6FSkrS9QmBXvWL676GIeCNRwg7wuvlaMRvky2DQjJr7CeIz34LSKD8/q2cnr4Ej+P
dX68TjMbx7UwoIZoTZ560AkA5F3f7WH34+uJwuHTwNhZ2J8Fbdwm4SG/ZJ5Ms05DFvA53CoeR48l
viAq0N0l8r20+nGCymNgWek6m2ujI6IMT1NOl67N+94X3C2FR3W0H6r/JVUZ5q2mm35uq7Abp5tF
QIKsg86wLxhM9PLxLE7+A3tWDVrumybYmRh8XV/WkiSAXWJI9GEiF4CKM47Frq4DbWkEfH7BEHdH
IycDi1OBeKeCqsMP656IU9r5TOAXR3wQCz38k2d7bd1fGy4nbx1KDiqSS9o9Vb7wwekhowJC68tp
+Wn3eAjiAxRiJxrpLIEb7KpagDv3DyWRBVnBSJb1kHuEvPcT5FGD79bj3cXi8LtQXWbfJnr/8Olm
SByMd1Fbb7Ryar7JC24T81mcxreoK/KqsKQk6Zx08MjksnNbk/8WyBA5MIJ6QeKoOenGyhl8dVVh
4/LvvLywkWp3+7y3aIriTIQn1x1RL0n4XdA27idcCY5cxxcEoJv4BSRy9qRu25RocS2E3xvcBO5C
l/Z+ul9spJ+qV+Tdn4pYlUPzHovhMT/6Ho29QRD19buo5FXeu7IodL1WfXJX7252DDwYXW+l19bw
+izX/hBSKpY2Gtg+/Y03L5BbljDAJdK5nKx9ZdJ8QqMG2pAt9YpxgbOF6RcD4p5zD45gB2IDSrwr
lulXaXnN4B0MsbYy8S1tU+cTkpTIKXUzwH/o0DXAU5+cZ6AYDd/0hj/tIUk46o2oeYzjJiSjpvBI
A68Y7FCPTvLNb0A/c3DkBIRsD/KeJN399SKbPRIVf1ePppRv/lTmc/MfRNe7hpJwR5v8GEAxDYth
v1iyIeWxJ7Aw8gJVnfXuC0V1B4D9KvmCEgNYYJzRxRGFNhwMvtv1IWADEvwVZtoaO0df4SwAWIF7
6OOb1YQfZUgKs5p+4KhJb+ipVlzznbsLClXvY277a+j+olUP2tKyfnnFhZKROxyDktt8MG3Vc6dw
mYjpR8x/gvn5qIZlFtHQzXC1lbpXXnaok05RXkpFYegkmZGbJinyK+CYBvLlIm44VJaC7DE3pH2V
LM9PK53FHNnTKtNFrhLYG5+ExjbthFBfIKHty3Airc+fXluHoJ6AoSMa94dahGuP71ai3g7iEidl
QW1xbMYGV1MBrj8tlmCcjXG4hJNwPz07qjQRGX9UBk2CQsA54Jv2UxMuH8NgayAn3ZiWwK0oTEDB
jcgESz9ocy8xlt5O5Aq5NvJA7AQ47iH9rZWVPCUDHrbVPgQBz4l3K7Wwoa92mWy9nNOw7Dxk1BFt
XyyOcqtUDJWDbcEfwOmcp35G6vDGWGDIrAexBLWTiG7c0RZ9Q5p2eyVzuIj80y2ikyUWeH0jcWJZ
PkhuXmfUdBPB+Uhlia/hLoXf3EdVijfO5L8mNYNNcHg59e82xCjCyhDg/QELNwrwJDq7Z7TaF7GO
b7rD+DnsPWpuTO85Go1rWICCrL1nrVN2u0sOoaK8ZI+VJiBar7fdKaJUU7AXFDCSBGZEZHhU3Hil
WeqdxqV/l3fBu99+0lHx4gbGeGkNAwJFylNmSXNdNJi/bsjqVIbQmlUPaF1p4pm+hnx9fiZoob4y
d+dWHyVylIKbQy2lViS3/3+fUF9s+snUOE8l+KZcikEWSonwTygtFUiKR7S50VnzT0sMEMYB83ou
YL+g4/aI24+SwSJuUFwGqsrOywsv6RxsRsb7Kd3cn0QYxWiB6jKydxLvi43cpndv/1rD30UfShlV
fNPpsEeOlMV3s55U9De1oxKKKxtd6X7IEhRY8HUr3AAARndA5TSbl5aFt2EtTa8CC90aN3HvzOVW
E2iKbcnfmcJJCVfcZALokm5Z+zB1D6P6EcFBC7+YpsFsxpNpwhrRSjoxmCeewNdKzF1N0mdCVROc
9tGK+sAct4ZJpcF9cCfiXPpGTU2ToeZZpPqrZ0LsdyWN8EnZBuVCfDxL175yUEIsNEcBv05YmP3h
/BvO/GXOf/J2MnaxsdS5Z0W0iEG5M4XixNbxZfOY+53a3rrDBYSGNZsbpLD6cMXoEiNg9HgqSPFO
J47HvIFgkerlr+p0RQdWenAGj3fE1qDhBD84rLByIyhJgIZIRX7eghqsnxXHKEhCA6204bR20Wln
fm22ZJXcokcS5xso8wDLf/YaXHs3T37TDludiDjvK2wTqNk8h/1ibVSfMDK+TYcP6cujc0FTcyyW
g8l42sMe9QJyQaPOvLwxBD9hvQCeqNPYiooIUDeg3DXhc8GK9wsWoXva3ycbNZ+zyxDkKX7mD0Gz
WOLlhElq/+nhgNV09ttpR2HQ6Z3GvpniHS4X7SMdHanioyIipgpisdY5fTdihbbQzdyap3zUDJpJ
6BmIKJ7IukiNwKEOAPrXgd+4VEsH+DlF5I4Z3wSb7zYJDTF47JcD0TJsU/JX611ZmftcJE2oraNk
4Wl0GWc+LB0E1eWMJAPTpNNkiZFoReR981FIr2ZAIPG1VjFybG5tncQtIibAEi4u/jbeQbpmFAjY
9GDRwwIxL1jltv3DNMUQ4h7Uu6QlPqV+CrpACi0wwqawoOCM7zwTL9Kl3Xqg0slZ0FqARoZomBeo
Dk9uuxkUB2zduSeoJyA1quf6PM4wiyjiLypHZK7Z5DcP5UObnMsdwCQooxkPnLR4bJe7AXL0xAIj
MryF1fe3TDESqNTBTLdm90aP45yPcJdpX3kPH+TnPpdt88wP5aP1W4UL4jNEW0S+/tKZRD9KiWyk
riYGHSMXlSTPt3cOx+O5UwCKdbUTpawmL/7He12cC1yKR9kKqw8OHTwatbr7VOuP623t0nSociNK
HdKsjuBDTYFyXHQGqbeevahywvdv0fhup7Zx6pfE7PMmK4TVlyQ7VLZ9N30vfZ3RkfUjkLyvfptP
jMb7aYOw4z0LDKdB39lK3jrg80sGbnPAfEZG2bMximUQ9IdIZiPTnIo0OtrhrUpQeZDyOIusfGaT
GqMewtPbTcJdAtncIQ2Q1cqMseor4RgJzTZFtCZY6SXVHny0AoUgHJ/nUGRHUyp+H5jYUWezIeZC
/dFJZJn7L3pKnJtDqEkOYg7lgOk//HAu1i3DZfamw3uGvEnWZ2dT80iB+1IhOZgxFnYzOGytvIM3
AuSYevC2dq5ibLTz6XTCZm3bJMavrWWelpvJ84PnatDRay/9p1YcDiQzJR/Bh2JRLiMTyb/cKMhS
fat6BSQwsrTj+P9bRjHhbBjNhypHLb2/66X+LPca1xfNb0h3PwcJ8P81aFJxMY6AkWs6w4qkVYjD
xWeV3tjDrjWP6wMjQQ0SM7sfV+TiSpxBRo/jSRrifCzST9sHmJFuq8heBvUa+2fjb6U+OGgnauwI
bfriKWDqrOsQI+SpjQu7RYTkxIIFDsj8kqAyRKyxmrPcbs//sC1uiFJ58Qy5yi1LAHWfy4aH/C4i
iRoxyYShJ/LjquQNPa0MoRyLwwidMBCo3tGghpEzQexmMoyDCOEY+et+lHAkQdgXC1jCj2Nwzn8f
Aur5VBnbBdtNLS6LAzzdBR0ikbowbz87IHJ44sGehQElhPYhU6pNUaityIrHeb2rmum85aLmYhAj
4FxSOCnhSlccCcXFo0m86VEj7bjk/HfOIf3+mc4FNTNyBhoJmi+gXk80b2YB7EMWQxb7IW0mlA21
OmpUzi4pMKa5Ugje7SeiTgS5uCig2MD5ZqRYbMmmU0tpseg7PtTNdCZ6+R1nfsJJEGddkFD3tbf5
iAyR34LKAk/eidi/WVhJE6vYoMuxJGvVoeTjhVTiXCUIdX6dNs6xmZUR2o1ICRTvx6NzHwSyY4Gi
JJfPt7rPIgYARKxlwasgsHqNRywSv1yz73eWEVMQfbtdjTAk2h3TchMgIGIPEECMuB/PS00SSAhA
E2pOl73nM1+ySLwJOZwjA3ik5fmSOp6EmHyVQDzeUWn62mLqCH54OISq9YOK0BWtt6m2n0x+KX2U
ydXQUbp56Opf8mnXxzS2YyinypuzW1XS25uIn5XXZZx9JONj94bbjDxqkxiF47QFE46yIJUuny/8
6zz4lpUD7I+URQ/dBcz2F4QKER6V57c6uxZ2Yv1h5Av6WQs5Mc9orZhKHLc++AV+PinLg1D7FYru
2kAQ8RN77hS948Gt0eyRaVgCQW+cYIYumPeCWzngvin4RFmCRQhCbWw+OJWmUk8aWIKG62Lh8vOV
N5300QG9vi4JnF19tE0G0JjlSkfLnDDt+RrwH9KXnCEBoe8bvVM772TcbeSMO9j6eqzSsTbNAn74
3DHOPQ03WJRExroOstPLtHW++d006eGRgotuybfFU+nPQIbUQ/PGzgeNkSMZR2gRsMwZZMYs+hhp
DzPiXy4PX92v2sxLtt8hYp9UOZxC9TnjKy48A/GPAOrlYn0mY8ZUS7a3uzYwIbFB5H2Rr+jmUao0
nBEFhGKkohpt53xVySiuN1UTMQn1psLsAiqa+/o4bIr1u/DVc8EyBhpKcTIGYiNXr9PkYlHhERt2
1ihpIUS1HJpFNf4iiuDLi/Pg17WAHKR5m0J0EK7s92tQizP/T1sDSnmrdziNXfZd6Y1Iq1ao92Bd
eAmjrMvcR+NCyCGbZv+y70V1Uf2shJml0uaFD0VUQtKA1jke/jyyVWWjtWZs82Dy3Jg3yFJ2hCxO
Wf2SPE6kDkmGC0WlvNcDphfWo9LjHFXuX/xLHgRBV6umpUhlUjyFvvrq8ajgxSJM8hSC9MFaJj78
AT2TyHfCB37D60tbbIF+xar6uIY9gwhq0L16xvOrRD6hGZ0x1BSHdMagTQSIWo3yi5JYHEP2R/wX
QkAwtbi9oPYyuzxn84oM5aRK6iU0XqMPgV2LMlaWEOObWBfHgvszdL9Di35fQWmfprCtgmOLEK7j
zkmX/zKB9YMrbwnE0JHPiaZwISD5w77arSIkT1pkkaW+9Vs9DUHDed3xOpLk0sjAfSwZJXsfDMU7
oJKwUKv7LXlsVKr8TUKW8OLnoHEbmxjE98xQKN++W2dbTbKmbu/xE4vFpu1U9UYn+xyG+V8byZVs
YwWReJG5qpt33VbRj7/PUsbOncC51Nv0Pqbkbotz2V7folQIEA97zENoabEjIQqJuYV7lGH28BIN
QrBcq6S7MmNldJys9Pwqshih1i3iBBT16gxB+pF0lux2cDfmjvJJIWI9mmaeqAV/yE8R/Iu5yo/0
1auzXqvUvcz94Qssnn0r0H1tAMSt/tH7c8KZH22XqJ6iTdwGXypM1CM81EWsxmP/yKomD29/hyHE
R85RgaVvUs5TI2Hd0r+b+z1KkwzZOpGYtb6aN3OgSfMkknXcXFw0TX8SGfxqLwXdHO0Yanx37FHI
ajEL1jGMpe8cg3iiDH0cX1cgWebB4+2qC/XBnYRFQdkr3PcEyTTgGKpMrbIH6ADkV1LWdsj4r4pp
UnKgKCR7FdJ1sp20NZN8P6c5XE6YFDqMlCwsHpFikHm/wPQxkTJ26IqKTbX0JHoxnM5p0Q1hdlY3
WSszNaoKpJX/wHvGP9WMx2CspsFEXf0HnPf2AXwO5Xf/jr06mM20BMMU6BGKAjLBUDm+O79hceK9
ijMQyhUxLlEryIhWL+huOf2zxgZfERuL2JCGfGiol5BCnj2P7+bDHkD9jLUKTKIPBikGEXcZJIw/
Up6b2TkRNtF+39yi3GQRhVEL97AalvH3evfepT6bkFTD6iydNin/CvucR6bVXh5EQroYZKzPEFp5
tG7CA6Hv1YZglouLyfPBDUs3Xmoa9LoNh+BXgYgtZqHASW4I7zM8j/aXIrrwnvezrCepLwI1sGJZ
odQjspFRRcqoKp7zfcbR1SeSjJVJLDpaA96J5h72wLh8n/jk3z0BhnWYD5XR5PXcjadUru5+0Tsm
9J4kzigb/8Va2OSAvlZOR++kD9dbvs8iu4Kzzas4wAxMMvhs42ElOyZ95E5Zj5GyxSa5it6xS7Uv
8/3+qBBJAEEcvsxWGCAM8XvkGxf+Bp+mKB4CJjC4D5UtziOKnR0ki9Wls13EitfpZ8PAIU3t9HAM
kCvofco3ACi0bmXKIJcYBsDm2gxH9n1Cl8OXfGIU1b+W/lQ/8p5HJAU6uLI9UAe1eqxAA+ldg6dR
uSbNTetBJEempnQ9zUFn26FKP8itWqY+hMF+qshlpcZraT7dWSW+S7UHp+IxuyfP7tgsVn161JYa
Jpb6YtQgB+iWf5lisqwpm0Bbx1ZhKxHzBMyMrq8fQ8JsEmz6X/XLeiHCnfDtnDTWP98kwy2pINNY
XG875hDVFUnfIbM/Wx1XEW7j1TWVmxuIFSAQFKW9Z7tKNUZGsqqTX0DI7qyE4VT3+UE+hdf4nRj3
hX17oPaQKBoZkYpdJJ86oyK82u5hQs451aMmJK1oIZZfFovmn1Q+c2Z7fQYJdh03/7+/7Y0eHdlq
bPf0Eg1P4uH51W+Hu00rpDJCwq/6cI2du2RV3LQtccMaGzWJjra1bp9B3m9eZIjNhLDFRjnuc9k3
DWuXIDDWeerDJ3mzo0dSDcDQXysiZqa3vQzw7+RIdOGFHOwj/EPONSXcgXR/u56A12kFW1iDhIvg
emXd9hGaS/pksn3AVQRjnyl3kFR8zpcutWkXBTtSVhOfEBIigvwJ2po2VwcmcUH8P1bWwux5dNDm
qi8vfCx7CUZxIegMFyOBVueiDjdc6DZkzD5KpS176YoXd83PC+p0hyMU4gRND8qlxekGLox3rKz7
mVTM4iIeqRnU6eXHdETgOFfIzYDQyDpd+kcuvTOwOs6Ua1RRr+kXLmqttUet/1VtBjPJqMcwHdCb
t67x+HM/BmcU/uOb36JoK/5NrkFFFbebFyj0IayMAMchnR3wQCAG1DgtEKcSlnDtFU+pEZzpI7ts
0XqyEirJ8FYNFSch3xT3s0RbYNHsAkRiqC2mBGbSnu3MNalaInmOc8M9yuFUo/r/74hTg9psGAYK
JTOp8rZkGqUqP4qZqrYsCrkp8obaftulySGRqrGRzR1crOTMDoDEa5ObIacKJEm+TzPqkTzxwQqn
vk9ap16yZ03X3wo0TyMwutRwXcnItEM4l2S+T40ZYXbTd5YzKv75E+5fwYpLj7mmj0tnNCN+IgxC
z1CnP1RMMh7MuHOKomSNGoMm7h8EbOrSdy1KE4kN7v2BXHJsaemgNvvlzcm8WZPS141WTj6jQIDl
b9KKhTIlBBlr4vNplz+dB1PHJAa3xocvLTpR7bUvgu0hTRwbhp4IWRwAX+babmNCZRYMgAiaoAtY
JJpwErg8VCS8PDsmyMcqo6RYmzhGG34+sK473y27d0snMYmHwh9HtTV/bXSZah8ReTSncn7VS8K9
mj5U2+WgtSUIBR4d1Ob2qz8Zli7KTB+pXKPqmVtSY9KPpZh2wWF4TtMJMoVeh0f2n/hv23K0H/Cs
vums3Qldjsn+fRdKyslWHwuH1kco+cjoUJDSon7WCfiUBr7DQmUR+K2qKkNh9IpQSjtmnDC/o00w
R1uOjZaFuXQB23UVsDwxE8snv1uzEFBN0XZkUvVIHXcAvH+l1YHEGoj4Rjcw/pVxnlxJ1aJezD6p
ci0e33jWUkJahwAO5JZ0Juy5pdgppFt/sCQizDXaWgrYf80cpkrYgO3PkCaelUJJ9aAbOLSgdvVu
EmT2TalQR7JfBLk+s5NfqpytUDXG0hvgyMFlTDAWsE9b3u0LxjSgSu5cAz7GKg99zZGFVysKnnCR
fUTSHptwpBqqzBw7JE4rgO3zqYBKsRzv03+jCZ7XQ0/f04nFQu2oaP6yRWlEQEI7Y9eGFGXHUwyd
FUU1kgfcUbyhw5v4KfNA2e8z+vq6tFFALWEhfvevWjKpnztNvw47x/M5mSGgy9fhEg4qL7JRMJy4
3T6dgd3ck89KScDMEJK8ADslEwNR/9sf7KP8xedJnnk28Znd2HdKVNS4SmrVfWv8KGGKijd4C4M4
YiLGkQpMnlTJokvdN8oIXXU6UKlWvlBpaXI+42s5/2fYUKftqy2qK9QVPK3hqBtUH/57HIQmhNlY
C1YHqsy3LqRk7J33aZrAmA8oSjmDxLP74zOwuD5XSS1B/IsvCMJbcr6dnje+tQF6LRMtKpWMJOta
cx0FfPbld1huOpccqtCfYW9eVdvjd8gJO1RQz1Dr/kTQ1PCx8u0bsq10hTga6STQxo/7rSSIVroS
MxiMDzmreppIDPdeOdOb7obFYGiJ1XgRuLra57svD5WdPNcUuApME2my3rFIBvizQtOV2ibj8SOu
njPdipX0AjZc713NapaKpU7cnwnapP4Q77m9wpL2ZWSegsIQkMbtMsblozhSlnA8XGdUvTswGudp
fXi7BK4ZvxZCPvTPQqC26zKAMZIZBQL5+letYhBoUu3Yr5lKLLTz+iA9lLlZk5FMyr2SzfEPD12x
r5d85cH7tFPN+BQa/soOHwJCy5E2j5MiV6NbvLXAef41sj93kpqBCUpslbbHHWLyZkVtv1TDO9cn
BcwhRM4ct+aag0dXvuz/2p7gGF3eEGOhL1qWxMQdzxS0auAFJxlnHeXfIWhfqe3Dg7cSQn/qrgkU
UQUJWGpV2SG5W0GfARg+6vPEEx/wwzqSCm9qYju6doCXZaAKAz56sHrs6Ys0R5SH4tNoZhx9qS1F
BNPK9b6fAfYO2jkk6wWNuvWWd+Ot3GpDJqiCBVhAaYzrVSoPbwFbE2KRVaKZWi715pAHawABuEFx
rwUC6hnevud3ogWv5NghMJrPzGBn7oB8U+rwVnOitJ+aDKy5qbmbF6HHlJ/nfBcNbEGem1dG0p1E
5aZr+0WLpflPEtiLK246HUXjiHPC+JzNOFEvcBu8OC6FnmqrfF2CWRzANZXXcBhRj0/Z8ptZjhkW
M3q7gTAWloYF/ZsKViUhoGO+wONn/Fvi8BJUIfzz+ND7w0ajQEwojNZwxxIouNiAVFtM2MF2ICvR
CK6Ynqmnd4PUMoh7f/IChYR2/sswlg+Q6hBXSH053yn87hw3fc+vrsYMGm2PMvoJcD+lu9qQi6wy
fnWYQo7dSMuxuFgau3gVZ/hP1Dt3yRcIVYl5I8nkwiocvZ+4e8mcXJcMYVsZQ4pHnJoNSE0XxCnf
xhyDWpsVuJ1rKLsOCr4b0clzupCcWWTepvgVmUnlgP5GcGOZqMbiFle1yBA5pzwR3h9QM+7xV3LX
o3B2LQPJ146b5Q9ZuQpwYcy45FXI/tzEqArJYwTOXyqj86/KHCJ3hndYtwVpSul999oTGcE2+gBt
4LRa4GoUKEwuVFT2GQjFyYFz1oLeX4KtF6xtbbTk/lc2W7GSEHrdshXiumaE+YhxensVNkjiel/P
825v5FQxy+ugsS2hKYF6yYaM2U2yVCGxWfYAvfqgw3NU1xrTayQ1gRHpfSECvJjWPRHW8px8pk0y
tUlTOt7OqDXs0pTaJCctjVkew1jzWShaLWFNY0IWj0BUQ8NJvEjpEBICMkzunw/ngLLYRx+eXR3V
X9S+3JlL/LZyrRg2U1Y/aHn7GCiga1R45UaHa3djzETfwNY2iVcap11xHpVgorfR6iYAG3KJrFpc
zHglWhlRa3Dv8zQFGGY+bnARg4ASnr/XPdxmuyVagizYIW+FMwXdAZ07ONzlNd5AtwVijIkWIwof
a8CwQYDDPuQfEN0qE9MYTD6RLI2G9PL3Mjxp7XDBlsjBNJJhbYgdDUKwMnTcN93WlAVbqcbA0pKK
y3vZmUEuSegFB4bhHj+5sVwBfp1sn6aUZ7h7nmKVbpm7FDYbT0S2JIbA9dDefMukCGFVmvbWNfAi
BCMpHOttW43eAsDznxBS/jguT8001JEEk6vVGi8bBgu5sfey+evVmBpwJDXPlG0xYhYuxxGJZS05
ICGVJpkxJMPpAVNkL9ZSi9G4o7b7MjtU8kALH39jqsFfUbo+MNNvPTfgrmX6pgeWQ5fH7tFZxBKW
34w8jYutRvdbIGDKa7e7Fi6NNvQ6woyq6+veGlqbCutExI4zoFOxDjmefi+Na6GUknsKpjqtR45T
q5Z9Ww/WTFuu+KjAhWV4LHxQVN9i/X76Y8F0KqGgClT3s5GFPIjnX5t41hsktYSxvPFyxih/DF3L
XhRIAhAqhZYBSNk4fn18GwhHJxOmnW7mojwSrYXqfEDeAsy2Vo3syMMC8F/4VtD0uevB1+gn777I
IGYChDGmxk4KYiFINsoGdvU5Kdx+0WTZ8FQeHpOroY/7jYDzn6zQIJbeY4rnzoCZcdqGNhmGVWBd
nV2uXLzYLU+LI+h6oTLBlSYO7kLlHC/B2bRWAYEuj6wOcVPb+ZXLWmUIWf14Lul7Tt6TnQdbNT3v
fTQ7qunBGI3Q7N3S1Yy2N6s6Q/XDXVbyOWJ8Feqv6CFDllG+7EFF0QGvFQGCO8SQEq3b6qBLIwUQ
A6tLsi+yHeR4ml2wNDWPkbIXPqh5UFbsKFS8v8hzJnlCKVuvXzInOiKOBxF/r0xdIm+ygo7Ucc2V
0d4IkyiC/f0ioyFk3LQvEUf0tpp0nhQnC121PvC+CfTlP8dPdezEDRAkD1z5pQQtWp+kp7gozqrZ
WRGWl7rQuwMuTWofiSN/yZZzUVuh9KTuu6ApLDu6tHa1iNnKBxwILO+LNOT1pX5gqlo5f+JEXKXN
iiSpVSVAQdwmYTZIYvzgSg9u49Q4XtgNB133UilPhbvOsIuD9vFllTW8bjO5UxlesDetR9UkSNi6
gioounz6j9wxMji7+fY3xuLVZz4Jj1OqYALDZihEIMemiG182x/Au8agPSrKcMvDdhNTBtMJbgZT
QtMLbB8dCcSQgsUtEq4DnOqcjdRvByPnL0quRgnaDyzxoNiKICdjYDDjcCFX51CF8WuUl44nXR0D
E+tgzdewX985Ot78Co0zWfN/UvBeUeljZkaDaSYRYETZEZStHzstNx1WQsq23CQizMvyKuUZKNe7
Zz/8rcEuDT1t1181z21DpWEXY44IwtQNjjtMDXP9hokISU1oH+h9LlRSDtGQ2//144PYfRIWKRFd
E2giGaEQ5o3a/iZia+0a2fK96BsqVWC57oiPJN97hdsyiLY+qYncpmdoNQV7mFr1J/vZx8JiLX2v
KWpHwxpAZZ89KTMQfKvttAuZPmYFpGsulU71N/GdAQAS+vpJ5CC0poc0QQSadwfZ1r0+G+xE9d1j
Ub52znlPFiLFNqN+AxiInbfO88vQkfCB6Q5PBDXg7eSaWuVvlEKdYjJvVjb6eCLQTUMcGgZKJrsn
kCEya7T9aAyk6UM9dF6W7A0xI3mddzeuN74WlBEGsYTEsz1/FiquTqFB0chduVp9vs2VpjhtzD3Z
j+a0WxfBKf/Tjesbg4RXZeJ7l2xVibTwznMgMEfeVKYi2w+4U4PMpYdqhJXX9k7qy38a4LTfo4eD
tM0xhPyEckS0uJ5yH7NT8VHqoAFw+stNRnBin36Sepc0VacdltpU1eRmF8DWBLpbzYyWCp4NSXeZ
K15nRRnqtiCzrSG7vpH8j+auVcSPBDH0W6mAh8e5lTMeDQeiNZuYeeS3UxmikpCb1vrndQ6QuP60
idbNQ2RaWZwSkU4EfoMgj04BrI10goiOpBWZK5E6IUoiyeAxTxQa3udOHC9NE9Irre7jK6txnhYg
efwVuIrXO/IoeXekIMvZEDIgx1xxwUxHIQSOJ+j501pacrAFhZzMhoz5z0LOVlRrjzsW3U43lgM6
Dtk4okRwXi9/6WVxvkL64zOrr5hbReql5h0/JyueqQ/Ka2lDRNgCdC049vQANJFWuVoF/AkQH6yf
kxWim8Qtq8wnaRetEavrBcg2yMPmf5gjTn9mtb5dnIZOipxDgPYHroG6jObPJh5uh3ro5xrx3MCK
13QyXFjNQtP+zEWmnc3MFD4bSjw+VZKyI88DxnsnozKKsx3uniBpV9A/Shdfzk3QNvuFdnhtuuQy
FI0Xm+ike8Mvj3rFZjNqWz46JQiQwHN/GCppEHr8r4lbzQ9aeA+3jP2Fqp2PsvU84fiC70odhw5y
hYfCjQqDcLMLQZuHw2CE/hHwjpJ/lVn3WnT25U5EvKPbU+Ph2WSzAFZaByFXIIp/5gb/PvwMz/z3
WjTmQ5O4TzYpksr1pmB+Mt8x5LX3Kk2/i9slk9sfNPbPipCTy2/DBqYDuMS4BaKENbzu8/aDd5D2
6izt4LP6Se5eaVmk0QDReoqQ94r58G4l6ETAH9+YJy9qVj/e+NLZaibb7QRPbG70OsdFEYROgg1J
Euene2OAJw+c5JDa52WBPeN57zDfDz/QW+plYn/kgHjrWSz9R1ARGSNAbdU/70e+lso46r4C6mZ6
/YqEE1hMNXXwXseyE2gX14b2gdAeNn3l3PDqHQUTnd6aCIIy/3pFct19l0w9fYRpksoEXx56d8XB
SsBxFhpVhs+jta/6GrGvpLXOfYb1M4j5fy2M0366yXjTsjDJL4bHzZ1M93M8Xm85UkG+IFH+vmtF
A86J9iCUL96hpy3rcxGvotWTXNnqxVCf5OpEQ1pYj81hIwEQhAMJiYfTpNhe/U1lA2VrdYK0F9Hv
EduAtkNQJhk15Cv74bgXP5RQ3V6K4Q0t8EDs2F1aj9NSB4nOdqhH0kvwQuU7VR99O5yZ3s2K7Ss5
iwVg/i/fT9xeKRryc2U4yk7WMpGyDVsoJWifWoxJrCQWTQ0IUwULH/wxRGTFyFPx1HH1E9+wyUlB
cAJTW2CX9gNJoSu/yo7MtOd0M6nBI1k6ZRK/qPuwCwt5SjbTHNHkeE0OrL32Uq1hDoVQIqd9ngtd
65MdqkehNd0U1Y3JlYUk6pLoNwAr1660arxM2TPZeg9Trf4V2iSQx6fByx+U3WWD1FmMzbcLXTks
gvHnncTUKgnK3rzrTc3Buai6vwIec+Mzz8b8+TlgHW0w7F8TqiI+GIHMtEMZ3JzEgN2g67YTPA5l
THi3Gs3oUBLaKT8OvkU0UVnNK6bayK5551PejZ72ZoD7xXV5eX39h6T6KZuOnx7BeIN0SzKEmRI2
l/U5/qVrODvJi5ewzPUty8w4gO3d9HCIxQTVs9ofJoZ924ca8OwPlQyAchDgc+zJKRVQE8/od9l5
PospLgv2RivKkBzaYknllWCnwHZrCUP8C2+QUMlEFVktQKf7yMyJk24m08RmRKFPf5MSJt/zHoND
RLBWbMJC1nE3XGXzQWEJTLREvq9gLp7G9tYToEnPe9D1JtENCgTyrf/PHo5PrynFXyZi4aF2HXjR
7WX2c3daNR2lfiZF3ipa+8oZ+x+/nOXOn4Pjreq7AUI/doh2HpE19sriuHi/zncsvjpWhOVwR+bm
VhN1Xomo/QX3FJSty5vFvloXn7T3M7kUvpVpgJ9DOUCuFRV0Bf5NSH0dCxXBbhgeqjaQ+5g/A4uj
ucCYqcm6WA+yoCzuuKSjA1viUHlGDKuhFrluJvQmSNkPEdLuEb6nZGqNaIhCUYuh7h7Sn8TEi5xQ
4qZ/w1qeqHUvRBziOUOYhe3iKEuCAuQj50Hci+vydgjTwNDsv8rCR4tZi01BNaOMjRTva7GOipOo
pIn1whhNAtEKE93yCoW1W6Gd6gs7s3G9SWG/KC34SV6rH61LbC0KDwYxYiQyt7VelrdcxIxSgj1g
KKJmokgWaSGbsBzmAcBbdd6mf1UkVVLXURA4BBKrN2peiSQDIpXMnuv3zKEMTSoJfK7b66uymcfA
5vx5PW7pykw2qF2z76qmlmxnUxQOhKh1R4sSsSx/mZ83ynkci+c9MCWIrVjFwHZTpppjgC8ciWX8
rXeZYawNaArSSOzxgkl22fmdcMFpMr26JYi5AfWSFvFHsAeKvC8ogNAgxNyVQkZw6YbLgP4H5FC1
yHXhkS2kDIHpxdQO5Ei0MzjWbiRIRe/MIzG7jTAL7FRROF3Ohnl4qPJdqPo6e1FNN9iyNrQ5tL9u
JuWLN+nDyxmQjL5hC1zCcst+KouIEtqLxKDsuSeuK3rOQaNmuOcNcV01LWjnn+XeJGi3Y8nd5g7Q
XoVhr+9nUqgoieA9dP3NQe9XctC5xLn8zCNeZqE3LDKPs6oh+NfyNzTxr7g2BDmR8cBjHXDXTaQb
a58c1QqDRQqz2bD5rUAQHPHdn8slT/6HTMmmthIDnVXs1xORf/vvsORj28fY7NCZXl14GC3hNdaM
gSGWEaq/Yis3z82ovNKmUjMj5wU8JkSe0ZFLUS8rKuz9VGpkCH7k2pQ3/GecVTueZGEvtwJldvLy
DKYvcaYtJy1AGgPZADmCZNPNrQWsItDB5ropIg2vR/mwPUPkR5ellL3GDhVuhFQv/07dDsuGIutl
YVN35lEepiaHAdJ9x2R4HhgUGsNTolIL1bQXL5VRT/q5hOkLe17zOoWxH+RYSpmb9ll7g/zL1QMa
EYIdntyTGELxIdYKjEfyaGUrBZIKOZysjnewOpUD+CvjS3qUprosZfwlqHaQpW9HKuPH+f3azbPX
0TF2czFlj2CRowCxubZs34qkkdhsIDGxJGV7zr8ClK2L/jxkFXSZgTKMyRxztbD+UnR+K1OH2CvJ
XMHBzDNB05d0cdZxTB4jKyRif7eZV4Yvf3xGXSFIB4PX/Besrd2VQCTFulHH9zXJODkNSrljba0R
aLniZO9qgHr13K849VrAMj/tMmBau7ivdu3ZTSg1eT746xX2w9snevgbs17joRK3hGkFvGN/jZIb
zZyWBALr363VpdOJuqSQjeVMClWnSYN27/RjmY6fN0/VpO7RvbHvWFsP70lkUQy0b6BYvikOKDUr
kDrosdWH3VVwo6XyMnhZZTfSTdm3rt1ObjjKUHaeL410qXUqp/dnKi/esACxxlcq4gccclrgT0jq
+9kxllxC+AoBzHhyWXEu+cbqMT3n3sgcOeaLk97FgumCvR8mqlQe3nUt47XhF+Xu32xmnTd9MRGi
DbQ0mIfyNf5AILbyZXCqKogTqonNvTPwgJozXlTgZLJacz1/ryyjZLkrjRzw/NMtP3upE8VATYoB
Cy1g6jO0ARuEjvr80w0rW7eQJJpDjwHv6IoobQaIz53O4c5OPFpEAskQavN9cdUeqML6HMoK//2t
mQJrsTGO8lwlONuBFNZsueFkXedTvhjkKHpoETdXwjMLGquWpio5oyvSoD7lOHG4gGw8cb7E4noI
jwC38MJbr+bya8/NJb5Lfm1iEM0zttkknzhSKTXTlr9LyKHgdbihueJginqXsDttYUd1O3A5bHA7
gemK385QclxK+Gxs94hziFAcveGO5ETlQCB0DTTPggAZ+hC6PGLvadjKwo6jggoiu9yzaxPPFB/f
FMFY0+xIExJupL5Y2vs9hTUJdIkDaUFkSDrW00iL6Xv9lHKGimG2vmVEnLKorHbqQLtHod9Kte3M
lRCNE37/RRv0z/+nSka88kU/CZcEmmQo/ZtIXtA5OJRL4cVZFWfIiauab4T58zvTAusoU6f9Skkb
A4m60mvrxlIKO/3nYjeqnxJzRFn2oXDXKFMk99UotiQSrS/giv+CzQOWUc5a+Gh6b0xnb0mlmdSP
oOQkNuyOi2qSWMIvmu3b8vQkWXXGFZN8RR35LkJpKbKWNUxdLfsKP6L2Lmw54JXOOhGnsev7xtp6
p/jwaWqpFMlqmLA8JazWG/uRaSydjRIusJjs2iCXY4Db2JwUeEAdolcZPbz4BNwzjajDbqmiBMi+
gARHshTvnhX+bKBZWgR41+iRMcCgNh7ARbkqEleL2iz+9OFssgpRT7u/NlLN+zCus6Yp/f4DVyKX
oV2LyWATy/9tENUgeuNLt9adroV/qljMAHBFtLKJlCM7M4II3vAoj6elxZRWgM8VDq5lyKRhPWZE
TCxQSqyHToRQ0++o2A/LsDUxgvnxmAUYHBzHtjXKrzXtjoMj9trZVnd2QtOZgOkdTklqTgZIlKFW
cD2eP4QV3F6Jntm+y1v9kcFOx0a50VAmRyBvYns6nKTTAIl4k2ttveN+VYa84QzPkryCfakDnqdh
Ab+qE7+SleJh9A/ooJdP3M7AFH765ik7JKzDHKYnFwrgaD8/KnJIF1h17w3m67B1lHr3OA04gxKH
szcQ8x1FzAZ+naTu0vDBPJLX+5w/Izzq+yIstSl8wd0mPiMOU1sZy56PVWU5OomI3kyxIjU0poQ9
ShECSGCg01G0WMmsSp1vlF3wwb1nl2O9kpskYrOEm81Z8b6FcYtZOYce1ixuIgFBzJg4d7KNVzCT
Qq7q5O6rMBmObjpLtqSDPlx7/pa7Hn8B84xK4lUoOC77VoFtD94QeYDGJdZn/W4UXb32e52GwjAb
Sh5E2VR6osgVvdbeYknC0Q6CitokLj8D/qTaO7h3UFFJQIailICykAR3OXxmvaHMIMRYXAlPLzAZ
TvSbDuQZqLSPMCBewIQ4/dfdAYc3FHHdppocMqxTvEK9OBIGSjnrkwA30AewzfEuCeUAOEFN9X9r
Yo3NBsWSo4qvjpbAkKcqXI0hsfL43iCrdmkhLpdv3RF/Px6msLkj8X11uX2jc2TBQ+Gbdq1a/es8
AjWGbIi7F36R7UV7tilz2/AeKroAPsxvRIXdm4iZFDHAnYVU87lsHq/5UDgoqxQOGYRMLjP5YzXO
WNCB/lhbOY1oAukzsYNRUFXdF8VNc13C65BwCtPPbsiDVVQbd1dlcRTToGiy2MyqsDQrHc+a6bE2
bTux73Jp8vxmOvHra9lb+RZlp8+plb+XjI+/L7N3zN+UiwnRIPKg7ZRYrgK+ONir7sEvZwMxTYwH
be9nEcs9zigGc9OGOGPhNWCrJ9zvOJ6CuUpMbvFz8PKw3aqks59c4hczjx/WI67uQnWsRJP+pqKL
I3h1Y+FPPy5oSB9Z07oAeZ8GGtjGJaftAbGaqF62Sd3d3XYh9l60Q5UKKzk+6NYTcaJL9XBdY1GN
r79JNBRAb2EEr2AZKRiNT2TD0p9VXOQOjUa/x6J4kKFQT956KchKSApLd1lHECALuwsr/kb21G3Z
9jyNNyCuv94lyfzB9MAZ70Bxmv1hmq//9hi55D1LZVG4V21MSiyv2FU7mCq+POOpluwfim5uUhhV
xDySE0nC6ZJkQAz57HkaY9t97TtalPhJTI9jOKL2wj/WiBiczn+uG+HLm6qx6w+hQ8t5sendOpOz
qzhICnfFTSuPFppDahSqjZVoXFjeNCDpN76p9GXThwjdSh6xSDKxk2ZC1cJuVN8BrNhh1JkpCRgJ
ex0wvp/hOfxW2DRiWhT/GQTj1pazXqmKeSAYxLN1rgfWgzc0d1etOUqm0mhAyOEt7e2vIPWU8XNX
PiszYq21tZ8lvwd5BjNbNXn37x6zbfmuYOVRhII6ssDodP3a4WSMlSDPABzXar9JK3+5KjLv7sdM
BqliR0WLG9tk9XT7r/f4gY0bSDzl3pLKLjgyLs119/x/IHBEDmURhdebQtMg/8KCsMs2FAQXAcyC
eMfYU7mnzS1wZbuFCaO18JddFZBwQPNSRyKydOq4rTp2zM8YeX4oAuazQ6r37QTctUA+65Ezjk7F
mxR94r1v3WGlLCK/ALS1qKriCiJeAVCgzL6OZ9a2ZAbjaM/zb4nv7NWH/2d0xdcmqKmGtS8gFsqw
dWErNIRybOlO3b/JECVh8UKixFfXdo7+oqV6+hNkAvCCyl2AcU01PGLTJC5hC8tgQphUeInMGT/H
7ZLpMxpI8OZNkEVmE90tTPayR9qkZLmL0pEcDRLQb9QcnCjzQpt0dQ8TchTHZovkgFUv82Cy8SBj
DG6I/Tnpc5vlaTyhc6QrJZx2ftpncx/koB9BOw3vV0hl+KnHwhgzVmNJ8cPrRD0SFp4C07JIaVYr
izonobuBHvBwb9xdaMY5Yb4+HFoAecWXNTqg4EPbvFLrpd+06bFEpnjcBmh9JDhHNaxp/TpSvFnY
N6RlVZ50Wr9yarh/icLty1tOtYWNAMg4ZK85n4yfx4vhdRlm40H8GrmCK/c96gzJye+OgSsK0FI7
DMo+XufQqlif+5NBJVzpo5V/p/UJjfPzxOVxSw/5s8hNgb+SZJVeUcECJcU8m0qdh7S9ot9Rafy0
gN7pFHdAS3skbOFWmhaXdRc8QVsORlIDy6dRVIAAbYXEAqyozBslSkZkeH65krGpLww15M4NqWMy
LllVSn55YelIbXh36kFmWqTGvZjs+E4h7PiOJjKiSj3ACFyo/okHVsy2T+2ffStDxwSW+rboRP/6
6ABTeY8IU/m3DdJMNrU2dKJwE1Lzvm+ctoJn5cdklxEauRsbHHt+exJGyOEi9/N84/7H1OFpZ7Lf
pbBil/03ayzS6aWQa1GtGyyB8jMz0IjqK7bxlW7M+7/t3HV1Hh2NZzcJF2GzAO0xXabpskVNzbyd
Q75NuB5kyJkxI1l0s+Gb0c6y/irdNSB4fs854n28Q+fXy2VD700VWtisAFveMopwm6Xyg6cQqYNh
nx9ihQFiOKCY/5Dhq9i4P4TtZCllR94kyDiEeE9Mhi+MJrrBaFlpDBxHMoNoL5HydAjNXG0ZSLeQ
ZgyeX43JVvautFMAYRc9EfMN5Z2z0lAbNtjaYN7xGNeiuSoqLkyh2V4kTT+nH5LlwfeOapB5hq0C
SAhagff3KuwjpH8HyThHlS3U+vLIJCLXdFNPKqmOay5yiLjl4mZq7v271mtoaLjQXNy894vOH2XH
2BHMQmh0FxDJm7nr7Z37m65waEyJT8oENH6vw127noVb6OGRPEVWkGetg1q4PfolP+gQUo1blILP
Z7jxB+Tg8VT5exaemRRJvoA1dPDmZ4cz447aRXFgNsMHvMTDjzqKX/nXwieG4cVa/1O3gou1VICq
DssW618omZrpTNsLwl/e77hO3dA64yks/R3htf8fNgyznQ/32E0AkxEepX+JCyMS8B+D01Lu5YSp
90NMrgs/IttZch+kGROgIPL/2UeuKCgqDw5CxMJoDecAx+QzO2OjD5MXZcHC3sxwqIC/69WA4qsn
mSxceaT8xanQoePIPmIDdM4suQ1DC9W9Y9OwRVbBATMdg+ugv/dD6rTB0kJ/DQNPX44uS0Edu7gB
m5TXcVhQijOOpXQkLpR+z+7R3JaLQN9Db0A1VWfF0AkUPmxOiGBUb/TQWWeYXqv+dNP02ABK8Nd0
vZIDSknOHbPTE2moGfWG4ycIldgNboShfbMQ9vs89SkaB18f+X6xUIUJ5/EaHNw+tLMwxZMQbIyx
ETcIJ8JqFjV1vW2jdreMpazemyjoRXGNQ12yapDAwfE9XxoIQZy1TX5r5lIViXgJg2CIkmckPfPV
Vf7qpesWDny4BIE0MlICWKgDQwtyR6JR1ew4SZS0Brek228oxGLKKJOBqWuS5BYvq3Iu7+CW2Dgq
Da10TubqgdSMqgcmvxeMbpsizUqlng8/Bc0+oTakVOKKXH4Yk62lVGq51jkOtcijof9J6BWjwNqB
O1SblMMrKlfacF8YmV9OYmbDziGZjql3GsdzWyfnRKyunhtKHAuJ1A+KwiKzYPARdQdrimISFz5B
st/vdYUplxYUf25Qv+ZC5TEDtm1a2gK7QyPPippJZB1MJ9E1AvLSwkSB8YR4SiuYkQG/IB0jbwaj
I+/f+rqc4EEcFukr5WYComuDOCRyg9Dejp+acd3co3vpeZeIbXPrT0VSpQSNw51PHvhXmHbrioI7
SxsahHyYBBzZRuHJq8K8dZRZcqpB335ADl8XMJuW36JthtKExvYvMDUcwvYnwd+jdJCBgPv5pSZ2
rKYZj0thD3Cv6L2nlY5nJWXFB18AsFVUQj3YdUM5XkstpRXarZw4iKJ9b2yJPGE+479/fQu2rjUZ
Q/SG5Y77zccr9RaJhAOgn9m2d3eUSspLYe6YYKZdW3X61f+QYsSBSJFRmqaHPWOQ8NdOVvueI1BS
SA0aMcRMTeu869FfP62Jm34Sn7Rxhn79WwvQ7EvkojElBArAcJunipePudkGaXG1DYPXdNMuD91U
0MKJMJDuKGQqc+93cBV6FM0c8LHyK5ZbMn3rVhVNoYpeoEHVoDinIpM0uuJwBPbmH2usztqWUTU1
LnAQfrVsmYCzzdOeeKRNN/kTVOLs+mNXbNejWBcerMmSWFc6qLrOXbaD7DMymDZlxclB3AYlr57S
95i68D/HG0GeyKr2wAg4mly0ic9y/9lA+ICA+zRbFn0g+kz6B3I4dLuabZRbSyXAY3sWN9jc+bOh
3SDRje1ioaud92QTJAqkg7zeIbCgzSg8Qgzgrjc8A7128VFtyM+ePiiIoZpFGyDE+LqiBILFIpWY
ZfAQoE9VdBuXoKtpKLTczDpq9BSJ6oHEWvhOaX+8MKEbMVQV6k09KEVFmfgPUVsPlnKfWig6+dOH
+RqmvLFF8Pts2xWeqjPXlD2DAG0ejlNckkKVB8myHX5lvftJ7C6q9ETLII4jwz2tiMMcWNZrU9GB
ctpSGtceIve1y3ZnRZ0EjndDVsR4cUsVrM1/JtBPrVcDalRNv4dDEDeNp9ORENVgL+n5QQng9nIx
HqcGe4M+Fuz0rZSxMgVrw8EWdDnWaccZF6y4YvpP+ytVjWBp6szSIWvFKsOxAiPbFhyV/OwSY9OU
QbuFrCfKwT+ec7eZcoCYTbvZ9gr8bzuUBH9hWpGGpYv+sFsK/LWx3mn+HHUyv547WavC3Wdv1JMo
XcKvnN7+iC0+9dHzSymbXFVxaIvCsokqHjb6RxcQ/CF3hIPVQJV9Rj22El54ofVtfO1yFasCMWR7
iZSERBkUzzaCeYHCTId+LM7QRsJ+XtrE9cWOUpxf9pIAv3S9TfF4LFae/9a6/inK017ZmmizdvS4
d4m1ehh5AfRLaVAeIUT11j5AGdcH/YXRwB0n5B5Sl5lg8yntD/wKtEscl4zURJc646j5RfMxhJ1B
hitEjEXrMXnXdPpBT7VzorUcoMUTKg6WoBf9BfFNxNBy8/qVSK2VBYyXKOKEWRT2FMctSkCmNqrb
o793v3+PGe1l/TouwyX9OOrM49hV12evnIDVKuyUVls6POAl4605viTbP6WDxHdnfnhxdxP8zBgS
jdNY8A0khJOaoBl7s76pJA9fYvN2l/r5009BxzlBaCgoWRdakk6i3PNKRSQe+q9QZoDbDZukc6r8
UiPsXeBc6O51G1VWoo2+lXMMv1967De6U7EzBW/uZI+ALb9yWO3xvCwHnJgSgiAOdpQ9ppRk08Az
ImiLOWf8QBW5tVVt2copTuAGttN/GtH4g+fGlHnU125QsToG4QfRYBmN2kDXcmOaVTMgNAEp+Kud
6+ZcSHSsBYqGVV7TUbSJUXMNKWo4ieof0tmiSUw1kMN+oL/bppOYMOKCKlXI9bj8tsFgMykZ6a+Q
u7ATgHY41Ysi5jFJLIEtWonq1BmgY7gn5KqTQE+DPjO4wQC6vuINHBT2lCkcfRHT9bxxumr+Osmy
c4k1vLH4JBiEEWpIwo7IWFo9euzg9AUrQo2A70FYoeCjjKPosvUK7VQNLnOXTELwp5vkNJX4B4Qt
2SMn4sbmbM1dH3ihUAVt6TBnd+5nglbuMCux2VrOaX5uY3kGnMsOWR58jWrViu2pj84Ix3RnEqA3
l0QNVifdzpghwiXSwWwdJ/DSeDQ1ClqpmX6AOc6DKBZAaFz18QM/pUNYWyeG5My5z6XNmj6Ap/gN
WSPsy0E18v3ENs5HjJJFiVKAPMOzWtRJMXGRF4qnDdfuMjp8flYmiqbQzUaxpfLb3fGlDi0iB/T6
v71iCKHYfbKr3Wg3pvrxgon3OUHDKaW0x4QSRqn/kree20XYEwDWVGObYKwz6hyA8ggwM7kep2O5
x9PCCl2MYMngATqf4g3wAKDNbtHcBeYAtJNYLg8t09ru+NnaDiJt6d9Emd2mQNTfz5GvGYxmgqs+
TXTU+eSW7YGj9AqS/M2PEHg4TbGhZaaMYX/UUsa1jSWRlnDudL2U8Q/A8lEJZbSWtw6huZID2thx
HPdoib+NWCQBaees8tThc10DGNWjsC/3TZ5y9Hv2vFPxAECqaEyGurGeabGWy+NfmjdXCldHayNJ
yBKZQv7prH80lZDX0jLX97E+XnsbQa4LpZQAsdiXD0sWg+eTvoWIstdAI+64OedjjKg3PU7oxGAN
7xlgM6WzKJyEmg14kOKt3mipTJfTQP3aB79o3VY+WuDFOm8Upi6O1gv/DblgPe/4eWsPnndh7bfc
Ut9XwtxIE4uX95F8EOGDccqHxs+tUxM33p9afR1DqzZOXcOqoKuuAITHFEUinN0FH4LX2CimqkpS
n2Oq5j/YzKu5PrUym12JufuFhvi9F8v8wsKPBzgYbFeNU8bTeEEIwjAclMlNZPco9ttpH0JxgWvf
bch50ZNKswz4frAfVsLv3HuuBlYgOqBQTx7VUlsc0DDv66MjKJUsJylVK+wRtUXyWD56W/YIUW83
/hC6kINjGEH6xMss+ZadrnrxVTTY7WyhJMbEK2658gdfcOWYyMC0ZAM3EpEGer/9OD7Wk86r6mXf
dDT2HHaObBIBfoi72umO+13N7eqRpdodXSC5yDcAtikb1Lpy496q9PTqvPw8eX4Sg4EZs2r/Lj36
H4qaRiBoZe934F4aJ8h+C7BIkitxWMr03YoaJZ/PJ7pYPjUUQpy9EDVTNJrnEniHjYwnmXoeApbj
2RYMZqxObB2HDrnd+W9uKrdCYYbfsCqOE5Ip6E2LgMyu4TPsk6Ny0OfYA27caPz75gA5sypu2RPg
rUzoTa8Qi49drisd4NjGKeGBV3E7kQomF7EYuhQnYdcMhbr3nLinvflLuFPTdgTsaYCRR2L6CMhA
bDrugpo4xquwRVcAVEvMk+Uzz9IMVkN9VMrvDtRP3uUX68RFU9otnGWHP7HEMastZ2hdAoOs3f2o
2i5MJhoxBRuh3Iwy9YnX7R/wZ1G1p1vgkrO1zd0jivIauDqrelQ2nws1PMax4cU9ft6puzmkt5N5
a9kNTZZcCEgtVRWvU07dB+KdCdkCYZohEoDOTus4rdp9d+2tHmsOyt1e5H3jnajbw/dNB+265afS
u2Ygy/Ouxfgr1pEcp4Xphl8gZ1yIa1Yct1NrdR7uJZEHO3n60zERlf8mzxpwFLxin9iljplOTC7I
HfRllQulcQgaZBU7xCvP4Mo44u98Sk4s7pgjw2NOoirFLtoHe1j4TyS4vsOWjGOJc6yemiSqmmBH
vhlCvNyWWgXHLJ05SVXrSZuOBBeqitABpMh7obqyrDjTknHnlNOyc2jQvhSP/ozbjXtIarC5KYQv
lI6wkCs/KdL0ick97ejIz0gxgk9SUTCiWz29E2Y5MyzcEYwD/UiCtq90ljClg/qunUFXRIGMG/GI
RjXyK1K2+W7TibxMahmuGz9CBid/RMaSV1tt2KmQ3hXZHRjj2uGC4o26RVTxduq24NHm2MbQCA8v
8UMx8hONFTklKinfpaoM748Yrs1XfDdGdK68fl7Zpn0/CkIs66UKPZOfdNgHFSILH5sRNTMgAQG6
lYiQRiocWnyV2y8sB3oc6CDhm49Vik0bD/K7mwd4yX/numkKRfskQKtSD4AWfGVTql5zofzkTrRy
WZLeDhGRqQo/AUJ507oM34eU8LGFBPK3g/5o9dPOImcjO2Rm7RzzOOo0a9ioPJhqyjOIqhWHML8K
2Np5+454QrCBnxKP4aSTTyCd8bKzJlBxyBCHrgZEyN4I49W3hXMyxNETXZ1iOXLMHvZEX7h5lmHe
V0xEaQKybsVmw8nQlpCvN9MhEnY5N5ydQjKdAREmuevttiXI3QUyLRWeayRx0mSgg3jt3vG0gMbv
2LwfEacHDxgUNrgn40T0ycEd1oXzS3l1alkkGYcLXncYVXKmJE/0C4NQAXePijMkTJ9sLvPVASdG
jlAP9Tn2iv9v2FuQeFpcM09k9OqBN5dhW+WTSGcZ0K7LhmaWR57M/Clg0oIvp1CSOScljxFcN9qs
ViLK08oV+UQ4icG5dkYsELvLrb6uFv/xMlX08iYqm9oztp5Bg15yYI0IYQmbLkNpCq3hHtK4XQhu
MSXUc7emvh9VqtiZXRleEbtbjTVzy+zGkWSp9zA2b2Lv/EwPGHORCbZkZJOJbY6r7yDQJe5FAWLU
kG9tdLnYscs/lmCvIy1EmUSeuNRONLeZ3F+WQCCV6+WmNjzKVNqLb1t4lHfm4qaQ2G+Cc+B5/6CE
M/Sm1KXxUDFv61Zzm/ks0zb4YysHQ8t4D+6vA1TZXk5j4eazLm2QrxAYTRdbzJlAEVI6FFlnrrQK
jiBUCkCoHK5/SfGDFyL1KVq3uXozAhBxB6FRyZbJgFN0eJO4R3EHrLajfysag6Aw9v9pndqXpzQU
4f56H8bYCCQiK9qvla+yw2IF0/W96PtKGH3XpmL2BAqgyeveCXAMY4Ug9hfadDovmqVBBjWesXPi
3HLNgwGHJHv9ihogiH9EDhr+/LiJHH7oh+QHOj1MbW0voiuRlpwGzxCoVNEzgVQKxHA2U6FYbks1
SNFcOUS3cW4l9fTYd+ARVEZ+gbJ3U5+hfj6U0th7SZ/CKiFinVcZN6rF5+7p4nSVOIMw7cFTV2Fl
pTJvLSvjxmh9qkHICcm9x04zPLJKPVWeV5Vt4TRYIuV1QL+wgNOcORLHiIvgrN0uJPumIjtDVGY/
EfLTS9gneqk0Fj8be0swMbwAsbj7j48tKueq7oExB80LAWLYcsUXGaaeA0KnHgOjPdyIKDc6gSwl
MwVoVcZ1kQcMyhYQCs8gy9Cv1XiIHR1MlTPaRD1vtnn2dTLvj8RxdV1hHFTljYZehD98Wx+WtH4a
bybfUttlk5JEN8EUCtK+eZOFFgcikIq+vNqhP29Xq3eTyHofMe2BsCVWpxrtXU7dDzUb3jINTIx7
6D9gfNQNvG+YE8Kfkhi/iEfZnyBAhnDkl5OmG0kCHzf/p9tkrncYfp+zXcLZfRmcqeyF1hv9HMoW
2/flRIja1+aqnFtewdO/jXs2yROO2qh6l33guJ8txIRTALWD+CJ1utTkaSUhhaYEL28Mu3ihOFy+
Y5W+MfdwkLDoWLeL8UTpYGE2EHm3o10k0t0PSH8wg15bX0O3/YZFkG95Uy1/SUqs7Qs8rPYka4kC
qDox/l/FDYUTmNm7Ke/QsQ16h/6iz1QCS6J+q9D4fGfgFUD7fcEEBrvoT3O9W9sfHUyy6gNl643t
mxafLyfJldEOMHehUu2WDJ3HqlQlgo7eB4Bq8ku/jIHRoDNe53YQVkeGJejf+2SGMzAD/c3HdegX
E/56+UcmPjUWTEQZNAyE7tsuD13tiaQVeK8XhIUln4o3q5hZ7ytzgRgRCAwz8MKUDo8uN1MLdwj9
Vd+wIhLJ+Z4rIWrAQxHnXwoVY2CT5XLYURgdQLr1GxEN6CO6DDkggjOSURWGccxSczd6mqweHMR7
gI8OgUCoJuoz1iCwqQ3h9kwEPX9WTYPRgF8g10EWSwx8dHmM9k1aoqAjq3i7Mu1GgX5SpB6OaUb2
Od/MKL8xZPqXDZJOW6XOQpoiVK5DbJ/aIGqUi6zw7W3pVJorgseBp/xPTwCrRLJF5OHglGM6Wh0s
vcU3akaI4xsKbPgeYSOJeVIxbPNcx08I6iPdLEwi8vEY+/P1nNHKNkN4dT5ED3ycBVOTIrNxBZGj
4FHUQBx3B/eDZ1tzjfwJWt1P5nZSUeWugszicAoqSZnx/PDAVZvLNlllM+4g3H96cLmzmoBp5Pgs
qVKeC2+Xi3IXzgqIWQdFwnB/M9MK+p0fR89T3/pEhbolszcV3snYKRqWOY0ReaFu37R1Tt47E3h+
mTtFw12qN6UcaHeTEEbeLRglRu6w3Oo59SVXtDb6pfVVL56s7BVZx203Jj8o7c8+4oF+JbMpRadC
dFvqi0gtWGDmBE+mByQPt0mJwAf5H6JoD8escevsv2ncg+f2xFOmr+B6yGGOKpEzCv09lqlSddL0
XuUzsvhzYnQOGjklVMKZgszBrZ3yCryqc817XCkqOXeIeaOijLwL5vsOPaI1/rlGX9kk2brTYj/U
6AZ+1xQQ53e7e+E+gbgghLiDUVpkN20d6rdO5aLZk76EkL7kSiu5nGj9QtWRh/b6dVdV5eyoyySa
pCQyT47kcKqrtkyKfmYhsBX4dM8T+jlqE+rv7xDIo209NkGpV5AFbtwtjAMTNjAPIzYUqZ6bG9mQ
f8kTxQPJ30fgd6yBZIqatRfKFndnZJ8IYNOdi9LREVP3k3d3yF/ImzYc7GJ2SBEUYudVmjwtEITt
yM9w+sD5j4Kel2vLDMB/DEbfM770nEB3PYq83cbvLtmB0Qi2GU686m8Yv24+Y9haWpypXuLOPoSv
zS8hY8PRXaVGTpaf5y38nnf6+9/Yey9pJ/4n3lltJSjEFfPUopJ0Nk6K77jmmAag5fu1d7Uh+XNa
juqj9DKlQtADvh0/HjIw0lzoyNWPFMOgcL3b3EgIUh1+C0rGzaf8hdaDs42iBOtOqvgek8edO0pb
HIf1DmSHeiUQ7XuNrvdKiKWreb6sG+pcbMN/OIp4tBJEraj16rKTAqj8D7S4iKG7OtpJmEngoLHb
oANXR/RSHpVeazcpHWp9BNGICImUxU7Jk5kX1Ak1Vn7v13o19GxfiDG+GvyxV3pDDAlVwrthDPyX
up4KXLgEzeUoRjnxpfRloOuv8cabIl/18U8HWOQ1cOfpcmq051o6FufheKsGXSW/pUqqV78A3KmU
YWQhdZ7SkcWUT9a9QFOTvwPyU477AOeyKqKKDOnsz+qkLtf81fUd+Nd6zn+D/opABp1y4H9Of8r+
diZ4ke2McRdKBsb3L6zcb0A0THXLMqe/Zrf8JxwghXuTiv/bNlrMaYouFuWLwVPmllQBiUenQKYu
q+D3oJ9wDDbXJBeCkz+sdzZXerqgJzuJ3jQi+8bGvFN3mVMy67EyBkM4HnD2P4aAZXwHbFQDPjOF
QnOu2BDkv0S01QVqcAWED0WSTVY2UChEKleeBdaB09gJpz0Lj+dhKfM9d5REd2TsH5CXdY3BHYQF
ssTQ3Nv85AED23KcyYV1h4SAreqhfV12/6FW5CXUoRe4UX1sfL34jSy38OvpZJhtzIkV8VOlmunO
Gxac+zH/RUw0LjSxiY/rXDuJgELYiUlqmCmjx3RGT/L+fj0T4Sc/iFCuIV9Wqry3sK0jsb4ernoL
1tOSN4rzYwwN/qTetYMauvyczJJahZk6BOTYC3Gqb8jNHcwOL/wM/pFpU5Di4SDuqa6KcxxiFQQm
SfxJJ/KPN3ruA3+ezFpBTLFSJ3q+r0ncp2z0jxzyf8jOUvymuo03we6IwcABtKEZUUDZQ0PgGyBt
sCD2TiAYpB6dof2zl7dWW7WFhNozzbDesx0yt8yGNdxVb7jGpwk6QF1pUZ3MTf6GDh/iH/WKEdMn
SUVvLlryY0H5RzE6iVt+aNRTObh+Dw3XqIOUAtAVI5GjjNVC4yLY2JYmXxhzF0HwTC08X/ynatri
NtejZE6bxl+1hdmJ/Uk/XVN+fbLt3FbWbN9lyxigfW6griJOi5VKBwBxSZhi8Yh5YinQGcbkqSmB
oUuKqnFHSoWOZYdivetVWJzVKkGDHYFzS/lOOy8OdAOJcGDCJfketv7lTgc1AzqP7jne4ih23Xmn
PSXAaSKOdHgqa2DUwUmxFrGExg+vYakbGWYtcfepy+sGmC9N7FUtQfqrbhogVCg7wIKjZk+v6jd5
lxAo2K97oEVMRhSN0/r4B8hVPOOs9Hbmj9QadWG0rEZ6sk7sfrZnXKpBuQWzlfQncvs+ibEf9FOY
hl4bBSUd2+fiMUu0UOR7hVDt5mYW9EiAhDa3FJcwaQX34j6IVvzByzCwJb+iELdYzwxvCLn3L/tm
XanDX+b78Xg7QwmoIq2+2cKS8pDOOoADpKVkTtNuI/t42mNwb4Bu5XxYhhJDx9OhWDUEg71HX5dH
2DNABEh7tYj3jZ3oIIEqnvsez3q3mI3yedbY5OB6x/d/YzIstylnGVUqH7H0+ntHKdPi/h9m7dv3
4hUbPV+9MKoprIorf02q8oCjHww5Ppn4mhWuNRvpDiX8ZrjFt0b+ifaP6b2ra1h7ZkzebNUDjbx3
2C8RkKg/6XGPMlhuVprTCzzfTpmMsICjPpfh7o8Q63N56xLt2qvg+l16Izzkr105N3Rw7XqKp7tY
cwiRdJghVy22FOottOsEyvYleWrgiCSiBpk1z7XgxlHHzQeF8hkRd6QJCnVEEvWUl7He7SN29mtk
8N59U+JWPVYK/iB1F7PdGmNlGw++DC56KRXA8ErKmRYFOodovy8dd62tnFuQf8fDdp7I8uVQBZ9O
Mx9AbdMYq0xE3kVYawqVICeFWRohk4RWurRkeSCDhoztWFcVd3Snus8ZcDpVwSEhXnaXrt6w2Gtc
8UFxHSSCs2ak8zb3n0RkxALWU3LzSiEdQUERjaCV3liPHyCvCiZ4gt4jDHip2coZg/+MzTNjpXVV
v5+g4nZoxhiNkfpqV5xv3K6AHQTLdRbSCCFrKp9BlWOj31UVXDqu/uRgHPxoXh672SNu+CNQAniL
W/S2C79gIVFxeQDZLd05vUz54hnQb1RWycAl0qsS1ukT7F5WwUC8ynTkktIsZbEOPgPsTIQkd2K5
CBNdOCr+1uCk1BRJSgJd3X7bzLap9Kw/RHrCiJsSLZArCM6OTIdN/Z6uBlCtHDjdMc8bvVjNv6fI
//fRs5byx4NQaWF6FpVXmb9JtrUx1TO51Lt7dzMnOR+joqbLF71jcKXG7eoq2jQ6nQwO+qjKuvqv
7jQuNYarwfVGJOHDsnHQ9TzOCViZrinlUSCgARHpm5uOiucTBbz5rNl9L0nuHD0iShdf+I2+8ugy
UABfzVkN/Wi1lWXlMVwNDCy6iOAwadM87GK3vop1zDjNKdt7CKpNTIGj4k9rx8I2SQbhCo9qtZBu
X1WoFKyh21/lMgjViq0xrXOvEyoNwSZ/SzbqMD2E6J9QC5HveOkSWU4hF6wYAgajyonkbAMvkNTR
xfOv32gv8aQPuY7nvHFrReLe8jOBmYbqAxSX3Yz7UidzRDKTGNQI9LpOrWxVnuFktVWyo/FzXada
pH82qHRHKZpjfbyd4fJiLvheiuwSlwAwTAEk+cqBCEgYIyx5D1Xn48uPJLFAeGiF9OOlLVsIJueT
teR1EmHUDxx8IMvQMc7ULIuUYKj7OqoXz2HQvnplBWysRBMvIGoGJAEZ8DcRbs1FOWOD/+Bv2Lv5
S9+wI3eqeFOwQgQNb/qSc6zFTbtXYbq4mc43ZPe5jRs+DkiAJ0X3BpmVbLkRd+yvESavnUfDrVFd
XWHAJkPcl7w4QQ05sH/ebVNRiopXdZJm+c5HAsJMt8KlG4KzqTDyLWLy78wV3fqZDk0yoDUTJg3t
H5WYebAa0OaGMbuqbWLFRCoSv61X4QWttND3UEGVVN130eilZJanl7caJg/OQcRmH1N6gzobceIk
ZPTcbzsq81PGl01fIVrVuompUnht93qzXwam0JgBW4FV4pgFK6pPt82/427t+WXDAbD1sFBOHSiM
sJ/1vYYCDRCqvmT1cvT1fg/19lIqLV5UkYf9bnCND+cQefnkpX+99bNaZAytuvvzv0DbXWiaR4KF
bjVNPIw4WNgeW2cgOR6Hk889crwxUNhZblUTngfxI9YG86wHcoCD/EuQD88IHSyG4HG2gp/tdZKv
/xxXHHzEGiytNaunlJcCKwQ2yQl/mbVPuhXy4657KCE2C9uG+h4+L0U3pvb/BKj62cIQVQUY+H5w
Ksii/byD5CIJ6DeW/fohzNFBk0kTlgOeZn0qGtNJNvJi93ow9+qfPnC1UvPK/ckcUncEcr745yK1
Kn5I53ZbSXyMy7RHYQG1I8G4noXSyRNXONker1vPfVKbbR/5B8X5b5zTR0V4dc/4WQdwVoGQqArQ
+U8Qc41uQ4okymP9z2ihcCZCsGKXcu4pOCRm8Gi6ytTjWYCte2mLvCqj6r2p0LqUfKW36BN6zq48
SPhXEY2Xv4ckuyhcJ8qws/thVrS5iaNgP96sVs8WoTMBqnJkFFpm37BoCpMcnOmbg0QQVagIMSEK
LEcFgfd8/vnhsa6/1QJMytaeP+5l6mDUma371UJfUJwpMYhoBRlp/fkv32E9AMqAVHljMjOIs/+B
tm6NCgxA6iz8HwX1wqFdQncRp0Gnh40jLjPrYc3BGy1YJ3wKjmsEn7r1yxYJOfIyV62E7PHIpt2u
HCE5q3Z/akushxMrblz98dBwQHDqmeqkAvsgo6iOcEHEsJAiPJVsAlZwO8X31Y0TZ1r2vPVbiFbf
K2o2f1JEyDb+yxNu0JBItAHqnkl/K/2LZealOajw0yIeOblhxDl785k+a4Uukx9RlpljSbobbF0u
UrEtttVcPpdTbiWTr3YhkYqF1IQMIUHZp6L1xaeWBURLQ7zkJ5UyI0dCAc4Bd4SpiywtxKiSnqwk
mlWGV7Hp/djULcO5jpTj8h0R9Qpi93HBCHHr3TjK1uMQB9uRV4ZQ+94zuqNzuGVp1WsWvhaDmEaA
qBbA8nR0bC43D5Yl8pVSmSalTPePUeSi1jkMGQg8VvQbbpCF3lKCF/XJN88Q5zJPZm7tSP1CRhLj
IKmImZsDDudYhHNAE9COtwtByfzQxf+opZOV5viEyIrwGelJNNZfxjTJGkV7Pqpl8hFMHwKk9qTz
unONS/cC9fWvsMpW5EtCAsDJeyumAnKWHC6gNWtFKjMGWTXQqOjNIRoys7qVmz+o2PCC+CBrclE9
U5r2VJSZHclu9aYGgasZ+DHMtJqSKG3wEKrrIU2k54vx32ty8e5RVz2+iwZl8cVQryleAtzMXCcG
XFQq9BrPZhJhOZqKdW5zXx5EV/Xl49NT4jOKO2cN0v2RGRc19FCRLSny9LKlEPY+yFp2IT/GrF7g
6+oa8hb4vNt5Fm0Ucf8G1th6wwzHAqZY9l2IF6Bkhg3uN4jK8rBddfMjCTHkHyGkC3U2E20lVfiH
gG7qN88Xit9XkIWwvSwbo2G9r+uAqCw/Hw4+aPg7S3ct/7mADdfsG9SorqoznGV1FkWY5iQirNvF
n13QwA+xyaAxNbhcwhEobWFRPqbfykEDuNPcv4s4fFG5PhgwqKvKElYb6XeYhF7UmstvLAu6KWZ1
BJoib8NjCgCNGdVnr6FgdzV5ztK5VG8g/7oyEDwKFFZyO4p0Q56hJR8qeUbSCSOPREmibRZKkn51
scFqBpqd6fxBP7ttWDeVACTHZrQebYqYl21tpzpMrl2Jn50OHFqzWMyIHBWG2XyduPEBK0nD62ex
dD3v0cOpFmP1gn0fefWCtBZ0UU2BrPypq9DyI8YF/4+T/SAYpNxceqtDn2AiXtj84V+YHQ2Nc8cs
tLc6ouV+sH+s592dU7p+R+3/xUXSIWoLpOasIMXL8+d01oDVq5yavr28YA+NaJOoCcihwAhJ95qV
lKq48+TuKoVXanHbQo5WU+U8K2EnPZr2CCPy6osPc7TWG8B9vLUlPYNcXwVHPAzHqz3sm0VAEy6y
e1hw08yhAVOCZy3d49PAvcEUu5Lnr5Mu1dz6GCNtWwSXoHUGtYipFS6Qaguut2O5H1qR83wR3jxv
Q1+aGzcMiPkZz0F7X53ZSyywo23qAgM53R/hUdAy2TeIx7cTyeQAz8yP5aV3Bwmx2ocWZPLfeg0P
v4aPOW3q6998LPpifT7zgd9qr/lVrEF13Szzb8wMkw6pVxI4/IWL+GWdCb4oLlk4iateJMaNVZAJ
54TG36fLsm8S/Bj7Dfb9n8dAikXLVUQCOFpG3nHLWMpyuNxDSAv2in2sIrD9Uor2UPc9+Vuha371
ufqOyp6arHO9aVh8e0f2iT6mCU/52nhUmZIs8ZPP6dq53TX3MKENmVMuwDaO2S998aP6b/9y3JhE
S0cu101Ak1tdEwwKd/+XDEk3UX2iL/6g+c9yNHIbxK7i57QD1Hc19azjivlmhFOu9LO83FcZ4rLG
wcOy+TP2P2u7SXYXwS/0InhU8QbHmf/5q8R2wcWs17R8OlzDT92sYcHVuJG/aMKOOoO9RFzBkhHh
nlFXbdKHVHvPqvx9coV2tRstZ3+CfkNROWfEjJ6bJKk9E/0hDGcqRLPNkflDPSXS/sJzFUVZKleO
Ec5BG5ugZQQUY3u6F6JpzCw/f8pmjqzAdkn91eHSY9L3YUC5e1lcz6EVFuJM2G3D0I2LyZ40x+NK
TD7gcQHyF3fZLD5IrxohJEHMzpPqqtxLKXlpnHVpQlzBtk0w2tXbbJHHZkfOzIVzEdMMmAnqhEE9
ohETmJh1vrgQfKwp6o9Z60ZpZiKdurxcy+4sy/5k2O2aZe1UndzQ2c84BBPkuwvstY2zVWVfknGH
vmcB2rm0j0UaOFSSnl8t7uwmOSBfLMa9aAZzlr7Im7YLZ3jeQAsgZHEDzztFT+dNb/rHLRCho3vL
nboc8Ey6U0FOjQPhzlToRtxpVC3n43o+86R56z3BkOcRvewRCZ5n070NqFDU+G+w3q1d+WXoBgbK
A6YniNYel7NccwmfwAfJLfIj3mqdSlI+DWZ2se9IkBviWgfw36uEHXO2//I4cKpjKyx2+JlzcHbF
IrRCZtfr+rWl2yrA9YVQgGI61LBQsNYygAv9T98XyiA2bBlchAf2rX0g7Jggi/iVEm74Uq0lWWMT
3N6xsxhIvDfqDMesVfXV3bfV4b4kdCZN4ulpvauKZcCXsBCqIqinnyja1uFsz7ydUHOkRe9W/MgK
zX4cwJQWu3u3Iu7gduHdhSZphd0XKKXoICV7ONCJJ30JitwI4NcL5HF+a0p+8xsjEuwzKITLRNnp
9d7kB1D/QEj9F+QnklfduTr1/I9/IemMVtI67bzGXWBUs0bq/IF01PJVC7CM9n/QQViLSsO2CaRE
Mb41oDYpguK4AtZ2Lhyw51zj5VW2ZY8KS8NyCkwOnG1MhfZnxgsnjCsmngSm6ZV73zifIGiuPegX
NHlEx5868x9N3foamYHGtB92LAFFsnZd6da3TiasVKLdsXAh7I/+7WTh3vp9MwJERm+ShhgHnZYJ
mh1AjlVoi889wAtQseFgM+4RcSIv/oR2s3SCfC/V4e6IP2jfaGNCqT68QcNLi1Tk/lMaRcPAVLt/
ZSDWwrJ8YNbIxwL3Cx7/abyuZ0bL9VruASbhSQZYRo/CycVITMipAS7QGNJFjmMdbSVwlbuu2HfO
hojbk+2TF2TROEKqoGXskUyPu3SaM3NoMaSQaZccN8NM2gkk13vUIoO0jpZAz6bJUu5vyF2QZgGt
W4xlVDcKodyfxcPTh3JBjFdW94Rjlxmel/yKxDuPu5k6sTXtj2TcljSkc7gOw1IOjfALIVeHO6jr
f6tcruqO7tVvGW5gM4KKg3dslpIG7ncSjwjmVlbgvfoIi1Ik2/90kJdAcv2RK+zmclVqNqvVWPrL
2QEMuaAN3uNZOR7N6MeIuzP/eueZ2HbER19+ySC1pURBb2zDA2o6KXwcFsNGuVtZM0E+il1JMFUB
trHl1eO5BntSmPXfCw3wrMimO3+ztO33IWlUBIdEHTMi0DMQbAQO+kpbk8iuPIx3fX5vKBd96RSa
BH9Io24wQNBhzj+CPl886J0ahVYh2cLww+zvp8MFfPlZyI9bJCOlCXBfhkCFaGnPhM6ENh60xO3y
I0CHtgvj1yF5qrTyETrHYkZWl7Hi0D82cBmtez7+anqi4+jUMLtdVKNONqWqLxgJtzTGmfRR6rB5
OHOR9lEPd/DBo0LtewOa2N6HRR4Id0ozs1RuBI0Czb0DGpyKom/6kiQLKoJjplBgUPS5FQtan3pa
uxagLtl34IY8hWVpDk+cNmQ9modtr2ZG1pImseL7HsmrDcju6lAp2Mn0wMnb1xxrnv7r1St8nMRO
qk9DN+ztfehjbRRYxhnaeduSTVOZvwkRo00FFON4LGcsYo5PR1srE5afOSTtX2N4mhnzqroAGb5J
riaJQqj3+8o0QzCSvpZr7r6XlpHCYbf4hWIOPWt7mg24RSrF+7mmvTxjL3n1ahxRf0OXWHNVNXfl
1wIlktIjdW2E0crfkLlySM/njibJxufqb2Y3x7A+3ctN1JFhR1g3cAQlF7MWXl16nT94IsnHkoAt
/9sIf5I3VEuydK3xSirV24/+MAmrhx16CBfW3H4WRgv4lDRT2fWXYrwBiNDTGRDKNyMvdtb7t5B/
JiV8CrxMi9o/QSBwmZ9hy67IVSWecC2I0YcDK0TIrHVRJzkvmMMHNPvuVtcRpO7j1KeJ2CWypPr9
iUzoquoFCF66VKAuBzhZJP75H8XlkWiiQymf/oldsusAyrLBDwJmIuBOIet9extXAUdYEvwfiQa8
FVYIO8LIws71N5eZhPx0tBDaqFQvPsCDcCBFyDhkscVriKZGElAbljpxIOdsZs6GnsojuJYpFuEa
UOsd6HCkADrRnpNwuoEvFAeNJO209RG+LY0QfQmVjSE0n9Y6RQdX9v9Cez4qFD5vTwO+Qnw1XPKM
TvSU5sREclQIPlkrRs0krexZvRij63zMbPjWCV0NmvdhQAjn5mHIytF6cX3xLsYWUZe00BzUvnne
sULdibcPxTtoobjZKjLC53D+StphuNNJRpqNP6fA0pT08wt9G1FpmYE/soUk98OPo1XV0dDdcyCU
ahnTyUpFrgbDSKhBAc7a+imUDAQk7ONAWWSLkQ1Un/Hq+I+Qt1QSxNPNtY6i8MB1gTURpOXEU2E6
QGN1GMq/oExrDEKQdJ6YWM8Quz5wre5DTEgWvd9KrK4RTkRRws29fsaZemNzM2PHchbEY7nABePU
huCwvpdxPR3A8ceHxPKym3BMvceYtxkuH3/gaBUPjO8uwZLeU/qPaC6HJoFapvJQre5Reomd8/Yz
nY6wJnFMlcGSVJH+ELgSsGJF3gM7rIAfwqye1aboVv15eZRQiPWBmSt1crtpcZHCyCYcP76MuPrL
qFMe3Xq4xu/Jiv6BYbmn1yYOEc9fmYx47Lz0SkAqQxuV6eYlra6RzSRis1jq+2yg8mrFiMMIjJaN
3poqUZ955MG4AX2v+iaKR5vJ87PH0A5f+wpdn4+habdFLbHZ+xqd2JzdjEN6Bj8i3bPjga+AESvP
18vwpQxruMd3frga/ne1fojJ+dpOgP0mKSbNEF5wLk6OCIya5T1VxpnTSYemo+LWVkRY47YtiTor
fxqfGSfooSl6lYsvgHFC4JQvb46/DjF71veav8nezsIiwuwwEkKmzH9gRcbPjm4A+E5A2+aioMwH
q+/LyPZRgZ8pwlharbswdOvCjORIMSAqrDVl8V+SQWHsM9ZLzu6tQoI4p2ZMr8BYV8cn189n3BJM
uSr+3LMadTARMEFLRBz8xZ/7MX0joFKUNPOT2q6iF8kX/UTDvtuiFKObY4AuqRs9pK5bZCeqvNni
8K21LvfNlh5Q/1ozGwZ7xs88vdiHtwCfUWKLWv5sIlqEiOaDdQcN/wFQcRH+BztUkqadVwxJHGk3
pcyF92d0tG/ONalFDgNfR/+DJuglpZRVT2djK8OfalARUb82Kd5wDy/LaUHwyqns3BEd8Fp84Ln4
sPZCrZyo7RPtTFMvb2FkCh8EQT6AwollVg44ifg+haaCyvCHa9mgy/ZyI2BQeYsqOwxC1BkmozE6
w9CRnm8Vnq4JbIunwDnqkSMGx1ZqkTI3KQgmlWnt0XP0ILtBKE1PRTAAAsJGVC8SbSGAI9X4wWTB
R1Hj6d40RW0lhGintXkVo5VA2DvZag6et0oy3ys7zmKr8hJhe6xfmwqapc5/OA3sHtoOCMEP3m2Y
kodfvUkP/HzIDiOael3OcC4PSS8VGdGMZTEC3JVqNL5WgztJxhAzpgXGVV1PjM6BVbzodSc6B3JN
bduDkRN591Dvc6Xk6eIdNgDyi4Jk5givzhUtwpwM39jHAOjBk9JYvp6RJYSM4oHbpbDdOYep+EsY
IorhLfPk6yJ3QnXfW1W2gzokkABWXlDna3uELfgcLo8l5OxGNGXGGlusGEMSqkL+eAr3YyZ7P8E7
d5mpI0RDQXXlt7DTVmPL6aYgauMHEK4+gIBSFUeYHnD89B+/js+FSruiw/UrivJ1YhxPg6rq7JLt
QB6rwsUMxWjffsRpx3BQBXRDhXEhOeU5fhvX02f6ly590I2z5vMBy4RoL8Qw3qfggGf0lJ5kFDyM
V9L7bnAb81cFyrFnBxa7bB4Yl4HotM9VfBxoEgvvYpe354AuvGytjSb5tOZ+6inGRhCQRjtRDegZ
gzqWPsGcaFtAztQ/KnKXK8TmYyjAmB7ofaBRVHbxdMfConU+bsBR59py3eTmMOPQV+oEP8GNXBlV
He2XbA++5G7gAYYid16JAHgVDasYQL2clEBghidx02ebHMhj4QoVjuPLcPD57MZHZWfuRIhdnx+Z
/p5qm3Ug6XEiRHLGfnlmvkm/I/SmSG/vqZc1yJ3Hl4Mua3OO0ukko9VV+/K+aIu4QgnnSR7xqgUx
4f1WfwpFlp9aIqDMAYo9cNQv0nMWKtYgdNiXxmvv7FTsMI6FLKau01f5qdTWs1VpkQWrL4+rjggf
Kp5YYGL14GqM2TO9nFyhcfSGz1TrrP5YUiz2VhWIc0xn3CX2siKtG6H30izNj9NxJBbXTbChlHz1
LZkHoCi1Fdb4IWHwGP7qxqGdRNb+LQCPWpDhhTkPcM9wruX02NfG1dwMMB6K6FhQUnW85zQ6fQJ1
Mat960fSdR99Vk7++8ozpWHoN3If9OOqMPPa/B7jk6MjrSgVXds4crJGRzEK1BAnEfC5HrXHYm5B
CnrweOtbJejuu2klTcmqUB1Qd/lWfwagjcXPEaAXockAOuoDcKgFsuzL9ILoNe81UMGGFBFMtcJ0
mjZxHJbM26dT7d2bAerpUpQZipwh5o+7GZHAZ58Vu7KKs9DYv/Ncsmk5YxPn1fXyD0BwuiovtECN
go2/6Q5+7eyAKwhrUsLo6771MXNQVcnAKPakNIpNfdXFKlsbmnqrqGL0wvVEO/r3lvP2x4i7ZzH9
sY894slidjEXOJST1JOuiPgAutNLmNNk85B3DTGu6r2DZVtA2x4yzTPJagcOWhlYbWoF9APGMT+w
XveV8fTE2tS82tOWKMqhEU3OI4ZAO07GTyD4RuWvoew3OUdWKaxun5JQrFmsV6BdmT/SiQ1QWS0z
WfSxe9M9x8Z5cJN+cHwZq+Edy4PtwRzgITC9VvTvGH6e5rYki+3eSnd0rD/DpgguHErLMW1XyDd3
z/XpX4ZBVyJz9CMP32x0NEwZwEwySkCNDlhVKwh1sOIXawECKYHjLHqkcLl+McgDVe6eH+dvI/zk
75bGJbvVGk2TUT7kGpjw1xO+VzLpZhLDseP6aZ3XZhK+vaiXS4GygxML1L/Yl2QwC3cH+HoXys6p
oJRMvHqsIgMVJaX5qFgzEKJNIhW9c64zOgz/GCURYMly8/a9w5tPhd4xJiyubR4wEolKM1clMGOd
EY15OBTgI5wIkLpsm8UgV1W99UbBn1CNXBVNSX31ssI1BJ0PbNrs70AdSM4pYJizwDruK/Cd72Uc
XRX35yEgOjoPk2IzumifGznVYIAA11mXQerx5f61lI63w7Nh+FMl6MiZ/F4opHhi9nh9TYzgmZ2n
qWDIwbZI+4ryNbDNN+SPpOeLPA+2jWfJcBfnMlxCSrI9F+qIuqw2cEdNoEaI+W4K5O7b0UxzJOsZ
OcFCWg7LtuPucikFFAz14SBcknEuYELxRXNVveu36Wsf7jYGrov9m0ktz5BXYyoc51YA9BprGOeW
Ju+EDHqFZWdXQPxs4IZCiuns2855XkqRYTzlCLDYTIQOoL+VtLANNiTcAEPOP9KAgimntU0TuYYH
FkY2vRVFctfCLqaXSgXmzrO69PcRg8F0EQqwW3U7+8nu0eD2VBSkDTVJLf7slG76lW0CWp+cDaEe
Mn8gpXnrAZiiirSFI3hLDq2ytsgNMBI3YsmhchIZ3kMwuyOTbjWHiA/sOF/4vrUTxkMFV3mxXKI1
UpoAVuXZa73cQLCD/GM2qlZyi0XsUw/PR4RrudfOQHeFel5eXQIXVQn7USgBWJW5w248mN/hF5Oi
8y4JW5BInL68nqgi/kSD4NWo9HD2MWw9qCd3sq95ovxlPqaR2hp7rNVjjfng7ONeV9t8RcOvcJKb
jKsYDxTBwnp+Sui8Uiyh1D8ttPlZa+69pLQXFl4lIjZugXMyB1X/Pb2UY2qVfFBDUDV9kdZRaM3T
HDaK/8ONRe/gDfha+GEeMT+rGtI873QPInmdX2bt9pNC9Tvq7sOnPxUoWJyRKhQdsNuQE1xblToK
eGNZU2wdEQg442eGKN7ha3V0/JwVl1e5aakJ/60z+4B2M3IQxL/0ExSRJG3iIz/xY0CiebuElYVw
6uA6xWWp3OicD/hdsnL1i9jnwRmXU451p/ahZYAK0ZUrVDwmGRSy9wc9aUJKKnusYJDJE3WzaTvu
D+0co+gz7zXGEe+sHUE3BydmMteQWD/I8XEA90PaTkKyrZzQytWEWu2doOPPx6V/ZiEqoCH7Kn1l
gRc/ZHolwhY8GI6sPRtPwIx/Bt9xsEWGhC1IMjughfrA6ESeXgldAOJP5Jk0n+iao9ZC7LBNe6LH
fsTXb1X4r9KhfR5kxSJT1PAlTbp7QVReyFRycqtiYGPMFsT1V1UnUHO7YC3zG1Nbyf/BAoin0j00
EeL32xztyvMKP/7XFPFlf74DmS9R9m8YZtV8nDPGDXfd++aH/ehoqxJ4iL0y4Ii/O2+c+Gv5g5nw
tsPqdR82nuBqvvS+xEyJpz0EJyF+UGIIM+trYoGGgEujUSUNQTqXurOzQyrBYvTEJ/WmFi6kae2Y
hzkwUcmFen+NEk8F3ENyFeGt2XjZYhtoXsFFtbaKA9hVJSTYH34z4z7dYj7NAK5J1bHpHbaqUAPn
OSeMm57SILB0+GVhoD+5/VQ7k5PdptQNLRwobU/OHhtr6uZX2IfulEBao0X0KK0EVJi+/c6eXMJS
jJweQHrhmwseQxjT/czYNn+k14B0bYCPUROyQ8tzxVPDfy/B6xF0dyeCptsCXXRA81k1pX1BAuAb
G8ScBy7siqWapZyStYlAqjPpsAWg0Ch/8+yqSJzc+xHPlYgAcgrjeFI1Tl8uPxclD0JAseoDOt8P
k3fvX17IHIkLvjOoYcUFXK0jTD9VQdKtQK+Rv5skoxxS4m9iLJEwcWLn1KQ7cbTjZp9yYK4oEMNM
N1qSaM9TdcwNkp27Kdlr4RYdxT5vTR8u5z5TFjaMZHVKx0zVMm6zK2yAWjI1w8bQHGM8q+WtusdL
OQtsuj0IkNbjXlE2xDm+Q7SxxcmTlqt6HKU3s4j9wHfDtPUtCmiZ1GouWZv2WWNYHj1hUG5/cbpj
+TpJxeeCAJox4PwkPA+Wxh2OfZBPerc8fsAcS8Xl0DWk1rhAYl+SH4UCNHVdnuFa0Jp4AqXuCcxA
Ci35qfapSeJxs3yYLvoCqAS4VEvEPt3etgadnFZhASJlfz++ri4WeJzaLdoYHQsY83ds9VkA9Bsh
PI2qosAUBHZxnrZNynjTmb1T6cz+ibczzZulZBxUUSRUQywYG0Mga3FEVWIGJT8nY1lf5/DlYhrp
MnOUXM3SKI9SfBEO/rGm850mx65daNqZ+hjJ8845twbXlSQ1cAib/3yZVVE6sAluwyuFn3GG+giv
qbl9+o2kZ0I81pnn/HaEolS9DZaxMVoiyRR5HPqwXA3agE9IUbFYlKfwB+nApsIhpA5z+q+PHycq
9MtDseq82kJRQFsTwu3msxIh4DRVgbpDSs+bQGEkx7BvdCmGH9Rlogy5X92F4mvejYufddMO/fGk
t6bO3UXWnoafoTtj9+L6hGHnhiaHRQsRB1AsE/z4/UrdWvW7YMMU/7z0yWcjJri9JZ1GUdGfA+55
p21CRl6V8Fhmr7wxex2YCSO1thH0FDzELeQH+oc/jR3nWbupe3Vu5vnnJ43mf7Z5VZ01jOJwg/KK
XE5nb+X/MlUkWoWTnlWGl6wGYYTuaGmbB1fJ7eAPTFnMJK1hdL6JrMMImEG3aGifBrx04orqhz/q
TO99xqbZqcjyD5CCWwtXYt3L6EYpPkbuLqIWDtDvBSD1ghn/ebGdPCvBzCtg60gagSr6M2PM7Tkv
4JbQjyxxSJD+zfuJ7bkMd8kxVSNQTT5QwFjwDGKUA2EZ60mApK1LfvCE8uSHnzPNa/ZXPVZRn/zi
K+5wEswV/Lb+6lCHslS2DEPpC1nCBiLTm2dVEmY7vZzUty/AHQwPIP0VcDpuzdFx7J/ckVKJILrW
cZHMq44LeuMi+dC9DbsCiNeOAYyVMyK+HJMNkjRjtSvSfKknQjrDXhHeIyQhdRNIzjJkaYViH9Ip
W5pfqVQnRFI31kKALe/K9a68/cM811zHJapfTMa73slWb4UMxN6Oqh/GTi96GnRnDuzZXhkjw0lW
8J2Hwe5SOe7R68UmDasH7FHLUGJssoQce9qjDtoo3CVzemkkeV9HQdmApJ3Nc9Bl6tLD57VEBG5D
rDFDqI0SahnAxIoYGqXbIc7F1WSZbqe9FxF3sdoYQF+esiUQmVIDmr1VUFzzEptasOoJ8FGp31PH
bu0bZ7FVq3rCtCrkGPZELbps+bRvw8I99pubgo8i1ub3fYXegR6cHigJWDawrYrl/OHBphvkRwV2
gcIlyH5JIGyKFiFguOc2t9R3nQ7SqYp0rDhojc9oKYhInNAgPBLXk53Gg76o7AL7FP6YC1mp6tUA
P5NjwnRWqEBio0jkx0M0KyjenuZo4Y6mcuqvFeMZBcLTQIIKEzEofG8GJFrZQezut2iQpiPoHC7c
X/AFLvKntZNZcLkWdSN7LZ8TQSAD/pyH9HWdxwk7QQs+H4p4L9QE44iTiuG6scxeZmVMnQRfeVvP
Py3lCnHlqmIQmZvGOwYKQXKCw3f5hPn684jYudJKhXx+5NhFfUBSss0sinQRoEumU9KtZbk96ohY
Acgalp3u1osrJTZ5lETdXb0GLa2RwNEADQNkyttcxN34sA/82PZE+YpBgcI7/QKpHQkXlmt00oK4
ZeQTOdsr2Fic2thqeCL/yXfLRH2wdGCjK35SPFnGAy+YSr3KVL3eP8vBFdWuJS71AvmncoHx351p
D83Z5TowNbWcyaJM3P30Glx5GCvv9EXQBxjA6elayipJc+nxfTp4Mg4kbtpm4Tep03rZf21wxylb
AbmHh+d7ii/n0Ojf4t+QbYiUIoW0Bw1sHQ36AjcpGvGzeqTCp6xo7mgslozeF6/kX53mUhUySWpf
XXZpDZR6vDFEhx5ID/irj0X+inqjixTon/vmU01jB3akWkXto9TyYBzJHibo+792MjKUn1uQ7Yp+
UhKsxX+GfhI1XxazcYH+lUeFKAuvT9FJ4eOEnHbV/aIiZlv5OhBsrgoqHArvtcYoSa3M7mPwG7VK
IugaZKY0fBj/8aA6zB3kEYnmaLR/DEFRfZjvbwlifPKtiTNH9dnbU03uW33JjldEJvCl9s8MLXg6
JIahTYmasLAnQBDMuDhANKse8yjg3ZYJMW+LIUrzmYt24roDKa0YSSSPZyryJUjvRiKsqPbpNby5
5TQLSeY0BN8KwtcY1kzdorquWRiumAJq/ax2OTihUN+sAHJ1Fg1b59eroYhexhSqaN+hEWqcgDQ1
z6DxHBugQbq8Shb+NcxV2GHj+X6B8GQWYbQ16L8KLc8CPSxyhvveIsSQoUAqPJYk4wIvC35HocoP
QyR4/S5QVChCeDH2zgvDWyTsgX3KrhybQZIF4W1/WP+cUrntdakPjUav8QdqFwQ7RSv7BJlYnzJJ
ZiNovRPNblMRuxb3IOpwQsdOFn8W/vfKJT6r4KWkn7MId1zPUfxjGSaMlIpHr2aHKKaZPR3jrTDO
CLn0Na3BvbquRb8CuZtjPpH/qtXpeY538qOVzMHCx9el5mf1GU4t/fAsTiBS3UQh04kbZTFyOcQ+
3hWIUuEdI+FsnlQx8U4Tp0q+L6zxljGQOx7i29f0LvVuyxxGhbI/eJQOPkx8izGwmNkxxiZtEZvE
RLhdO0zsPhHgLjq+N+Io3bEI49v2DW/kpNeQV+S0V/m+/RkaybtqCE8ev8AlfrNkR8MpCBXVeQ5j
Q22wQ7CmISxFo/6SvVJb+w7+1YWu7NCHA98xo0iD20342DdARY1zox8L1FLoxUCbJiHkoBqyvDm/
PQ/GqamWuACXaqVJK30eqgbjYr7DmwH+ROOCcQJqqoU7LBBoFkIzHcv7xshlgyfoOMJGudRbps87
gtO6OL/dNGSZDlG+R5mkYryT19bVk/SOHA/vbrGDWOoc5p9R31uCuaw+MUwOaqhiweURDbNFY8oh
rtzADEFIuEPqj8FuXOYaDCMmt2hFFKJd6jxgDTP1hhgA53z6J2dCvKZ2bVN+E6pSO/LcZZ6uVc5/
rmxBtBO+Z1TeDzPLqf5vdrpuAj2qxlNMod9sdB3aCMjMnjeT6jkycy3MvTdKMNFAKGSJHQinfA+s
Y6sbwTGOdIjNJ01iXTPXOm9FamnooKgMUkAR3KunvruHcU15Z+RrwP/EGwxmzfNnixAh68sS6Ftd
6UseRCjLLpdgIkT97qp8y4Vc6CQ4G54W9g3YxbbQWTCaoxfSHQGOKYtAjz51xDyIa1XCmjR6rp7a
OSmmUDmpiWzAT19J5Cad0YxpVNpZZ4wvty2YiKe6t3fUUTw/GK20mM2kS/0yQc/Bu4Q40O2co0T9
SEir1NkeXZwFZ2IPScXP9rKGpe7ZTUrjLJlp0noPWTdt0ptB//C5CNvWVIs6+gnWFQFNEDbW6L+/
K9EUuWsjrK3+AAaXXLd++26OxEItXfSUatq1hMBNc9k39cqVDfzaHPKbDqmcKagY/sSwmsth0Cor
zlMsEWljc7WFnwIUsN3RjYjMEi4z0J8zcLae7u0ZEK7ou1VOaNqWlac7IQiZYpoeXZGTeZkhUSb7
iR8kZV94VQOA5qsIsfPe3c9cG8NnnRCRmZ8x62Sa5ROh7ffqXT4BZQ4ex9QPAHzLwbvJ8sukuD3U
szGngOUGmRDTMsbFrt4EGpN2vlzz6yPzdhVeCBDHkKABwqAXaBOsN4bbExmdtNtD50kKio6rSi6O
4AwwZzGCM+ERciAn2j6hJQnblUfCclDAgP7JhIuN1/wIrJnJI1dBjADFxB5o9JjMh/7j2eSPrM0i
82p3fqnZ9KTOK3o5mlLBycNnle6T+jZEjAnTJmCsYDk6KjQ/eVFz3c8K89B152Cc+R70rEPJIA7d
MansLD0GohW5mA0C6erkdUzphqtr0sLmnjSyH1wY+kUoAN/bsM98uffghZt8Q3FgBzONCAt8Zdtm
7SHxOa9QBqoj5D9XJVd8ZNh5oaAXOwB/LUvyTHeHkDoRYmBa/MvqHM2I7xKwAV/WJ+2V+/jMSA5u
hBodueHzJezsiQunxwMAmI9j3Rwyt9wiTyzgYaeS6spcaWUdtqDKUp4/rEKOiyYrST2oqYu136Ss
fBh10o4z1tk54zglKdK2ngv2gqalZdKfub7DbHs96455rUXKSFUIhNhuGBQgopSyZSKMZyEcPtz6
dyw1/G9Vj5+K89E2DWcdI9WHX/k62cL8//B+l92xjGm2UIycKOAnit45RlJ7679YYz4+jt+FKXs5
TVkbnrQFI/KlzwSgKMYbAOZ5+aYhk3m3lEHkhje0CMmotNsnGZ7TppERBihe6rE+nY7n+SKy0s9T
DWRhqRU9MSeweKUUqArCxdL2mJeE0TVfl3IttshjBJ5YwCTgSSiIr8LQg4Pbb14h5wtX9EWzIq1C
2rPcMfKdvq+EDhrofnvS3WkPAwjgLforETrJDa4oBfPD/oHK7dWDN96B2x0VpokKlaq0hx5YiYta
BF6eBnePsG4EUU2XH9yXzR0zylWrQ+hFKm3CfnghXlDTBM+j75Bjj2I6aSZl9tOymSGMMoGGZ+GG
uzTAb1r/B6YZeZ91tePLBELN8FvbYpxxiS4jvkcDIw32ZX9+TUSn2mlvG2U/jO7u+/1YcQUZe8aE
a+8mit3jxeFx2r4sJcibIq/cvp3lW61NIVeXhK41wWCBi1JecSZjWKx7abTFBvHBzJLoPwiJGyMk
XOmIuEmLoccfx90brFCUCmE8YiipNBgN5fUKR9ZYSwxKidtTfXRzi4KOKWo1057fv0MVaN0JaczK
wVSGtxUsU49dz5MketDs76hGok+5rOtdEXyHMiR2Cq/5YazXtTllU+6RmSgBHIY5sPmXRB1GxNlV
A2o+DqJ+GqQBkSyoRcvfdjBmNs/umhjo+EpjkFBdXeD+H0jYRESbECsZQtDm8NNa9TMAEuQ1f45w
Mw+cZ91DNnY2ihRai894kzjGeFVA0v7Y/PuhBXnHdbpdeiw+kLR6r7DMOvDhYG8Az8Zk42OY0XjW
goNcOoo2yugCyTXax4+ZHpsE/WVIa3cRdxT06rnNbNflNddvyS3QZz8n2Zv/xRSvDpWQvtQPdJ1y
nwSOJiAtBIwMV4Flq+kw6/xQRY1xNmBon0Dpy3k/3fn8leQlFzXaVyuJEmiWy1ORGmG4nbjpdxg6
mgDSCo3lzHLLgK+DbCdu3JCQJFRZs6N4Y3ol6smtxSm3+gB6k/hdUxXnnWnIl+UCN/OR7Hh2phin
IkKykvysSNb1jn/oDQYhSm/bAXCiIOBS4oaeAMkTGE6WQeQcSah7e6+EGhM59m+mbnyIHaY+VctE
hW6Qw/y80yjtx/v6TjRvqmGbcWfjib+eQsV4fTHjqy4I10tTlo3RVa2AuwwlPQTIbva/oMoLZPlD
2gVXPZcsbz1SllodbVdww5Xt4h810FHUvSdueP7T1iGtopPcqPypYYVyPQspwZKwx4C7MYe4hDdw
YTlDTvshCtG0BUJ8pDhPqg33DY+vY/S+HPSq0O4sRVbzYnneVefF+eRmmsleEdE17waE6fSt8dMv
Hmj91pPbWFdqpCxxCkyL8Z+fqFjNYtdyi1AGHzQHoa/xDMCtSVXs/VjYLxTEa1jyrhQ+PY9ARv7N
Jyj0jG40KObZH7+4OsFrkZZSTDOnPv+gbK9vGOOpf5tGhcz3oAk3qH2ML3IY3wdIyYM72ktRAHie
IYujJw1MEZitK9wECH0tkHjFYkJDLDCwFjjcUqOYW9/guZAeINE+S3c9VuOSBaR3gFJR9G1o2ptZ
f6LmGM3pY282xJbtrw9OfDgb5RrOb2Rzdjb/3d3bzjU+qAcicxbapQNIjNiP+UsQ24k3XYM+na/V
uwfXmNU8aFf6RH6SDU54KtEI5yZoJskvpktI6CkHGk4zd/XxmE2WKKtwLZQUfNdsno09vkRPSjcY
pZgu8HfATuYjBZyTbd+netd7bzIiUKfYGfKx/8oGA90yqFaAdTafRovaLUOlyZyrYNJBgOD4Y88x
38mzA1gjx2a34BUhxhhrmY32wntTtDOu2r3LDieO+EupigUx7Umlo2Xj+IcwY65O8QHJaWhL8DDJ
YZ6KGy3DpAyhdsEgnJfDPw084J7n7om+3V2piQuNmmc6h/CGuBBgcdz+0XATx/iphk1ghOy6W8uU
NCjZ7/ILVsU8EgwiZVgavqME6Zq0aeqarRPnVudfBqhv+A1JV/gcmyz1SoDpzhs2CiE4enwW5Nuv
H53KMGBDzOo+DzsVYFSYptqrAImp3lTQonS1oLhRqmOEOLw2NuVeTA+5cb3hpDdWtXO0L+y8BkFB
LreFUOrPiXEwyudw7IwKZlXY3wcw77hnfnvsNr0f5RavLj1YqxQFEaiWi6qrZZo7CQSMTcOqN0yl
rSKqC/REDha1TyErZ5mIF6HcgOdtzvMhzv1ZchUWY/lG4B24XsBZm28xWyGSVfypRO109kzhf+7q
YF5LbducfJCdeaCMTCk1SmhC2zbCaRbjG5rRBGbjxnckEpmhyU23RtHPjlVu4CWX+/JsH2SVr7bn
DVQ8v1/2b+Y3De/xfBNaMJ3XzSwS7nzleEjLQvHaktzcXbKmCQzI7abbz9GMP8//ijR3J5xXanFp
CfiDLEs2LxBzSZ6OrRe6WdvocFnpG4MZo7Dus24d87CdxQApAil2ARBIHDE3e4IlujYICzlUnsNK
L1SsCThpDD7CXNxs0SDc04FJcbxPq3JXNhdzBbj4j1qrOACjKAafcfYN6DryzZsl5N+7EvD6LlMV
qMTohVTQKrpLFCL/V4mBN47GaYrAr7/Rt5fdK5cV5e30HzbsY9A9AEUY0AQRbfoMSavyNeAzhpn/
SIlriIETBHs5AGsm5uD2l4UG0Eieqz3OLygxmavr14uvbGvrzeSXu0oo3m5t8YFxFfBJJju7pLL7
iga1QNvWxxqjCLUeY10EsAOtVtxnti3+ZW4wQGnAbnnANorqv7yv840tgvSsW+12QS3DbNe39+7c
O7jzebJEyIPkkI1wZAB/Ow0n9Q5c3xsCNLZWVbRSgGAJ3AEvLTXXHxbkcWAJdNimEullPZC5f4Mc
sRLJ3F5HmOKLVtNNK3WGYZoBsM6DLnLGfaFKpWjap4N7EYNYIoasykeHMV1X2hDgLa7csZGdcKiv
yoPpwQOlavCApswv8HNN2aY6G0Nvow6PKjJxpop7TuAzwVydHuh9ElOX7zwp6k+gSt1nNVGdB0lX
orbwjxx8x+O6GCG73OTh4CZOOXbVp7XyuPxnDrvPyNdNMaRgXtaOvWHrEYphx6M+tfvM1tvXxoKP
lrWkmlPUXPQ7k8OX6qHtNNK9S5E6KrBguRI+H55gSXXUdKdF3myFtN8ZZCYSsVfPRRsykLE23KPT
sGh9YEHFfLW20iFuAOPwutkQiVahHU6QXVo23OSuRu+d2tdVQjUHlkzp2OqDB4qvrfJBNag987iw
QWWX0vwW9gDL8DE4mdiFN9xp3vtq4IhZ7mZ/FPz/hOiYJS8TIWtSACCSWBu42PBMiSBQVKOxzGTT
4F1z9BzOvt/5tYInUL/I0AGp+F597m3UfVsUivNCft5MitRRdClrNIp6W8dS0Z/duXbHKgAMx4J0
HJwfzbGl9y6bzT1vn0ZqKaI3P+Yrb46BsV1DHAhJoaEnv0a7uHaF6yr/YtjAZ349XOppXrJwn3BT
/2tMF6OHgvYpswfSmRv+ydr9GAjIVucIer3IpOtJGurujQ4ysNhbDTTwY/dO5/ENJEo0oNY+Jw8H
8rlRoY492hQWALHVtxB0Qyhjk8GPqmzssfUJSYXJMGog8FCl+/0rHq5MwaerR3GZBqEXBsLEw6DX
Gmlkut9UyltLicNWwnQV1IOXAp0d/likbpJBtECzG7QgKhWMDc6zMQJSQkeYYdLLAf0MowB/jzxz
9J6hXKrM8ur0FoRd8kAY7vrXMpm+/+rzGVNUyQQzEpqiq3mmrJDyBIk+XcKVp4lEb3p8aYJeQj72
PgIfo8Jou6dmkg35pP7hM6lp+c+rayINspwsjuoFHHYWPEJjkaZwuCNWidf0N+LHS761jIGGfVGD
tYY1OOAN8Ar86WgB0VEkLG1TKLUWG30RWi8T1JfSES98dFaosOfc70QNEiYaZEFZL5h/8oQ3ce0V
r7O434t9Fhren+T0ANQ+w1bRWJ0YKbKW7Azxxdd4jVp9TM5uy17bRiDtAXEYqvOW6QdQQfM2RK3a
vk21/ek0MvyUhSAjGmwd76V2NYCR4OqSvdqPHHAumKYU0CNAXlMnmrNSURP99NDD3g0pwcpP+sal
oSBaCi2ysSqgw0Eh4AuteswdJ09yICj/WkGdEIMg2ctQKNdlBzWtFcwds3Ujgf3eG4JokShT/soq
LvZ5cNj4SSdlMIYx7J6b5HlOvmJq2wFfvOcbJs0fnBc7J/Jzu01QHqaX80FOnqPlAlOoaTzWqsM3
t4zO3moI5alaC6ThEKTyN2dESmorFa0BI5JZWpvc4smPEgHgPaiUAmWZgPaMrp3STFaDvfM7Aol1
nzvdnda8HmJBhlULFNLrw9uBZ2QOtLPlW3C/ZJECh5pS+mxNB0crO5VO7AbNoaTXRqhNgqvHGx9l
3NitkCMcJrNhSyMvFJ/i3L6eZ19Ags73V+v/MGrgd4U74qYX3ScIPxfujxUTn0iYne6iIA9J9J99
42Eidhl+4BijnCVpg8inI41pZaPaMjAWVwlArJT1uEIEdO+py3MDmKm8hYKLzohkD1WCOsm0TzwZ
BXZiIQFyilUDH5jjYnQsaks/V7LYbbJugwKrcLMGPL/WMRGgueLh+TFQR+4eLNprZRebZn87jFHw
0qfxJpL65ijlh4jIrGQNqDsyOmuaRuBIbw9z+6r4jCB9/UQApLq0fuo55G+zO1B8MMAjYcV4jzAh
gjpTk1ExWXkA4e8MEslOEOOnJe8VFXD2XV0iyhevMv504SowvP2q0TbEjupz2K7/3YNYoCMWg/8D
HjIY6JJdpyZcOzx7nEmnMi4f7kw+KSyq56wi/zK9o0uHOgCDyhF/kgetmPwZpfykxbIuS3I0Gacg
eUoeAbbCFJdW6Mz40GIMq832sxzN4fCCK50Weo/fL7g01EwagbUbv89e/ynEiMMzHxdoqi0yn3ho
+3GF4G3PZXduGQMLuJx9J2ajmGXf6eulG79Ngoy5L6JINYhEcMgdg1nupsO3EpcZaM8hg1nam15g
HHcBv0Gtr08+xs90plo1DQ5uhGk+ag37LilWlxcUxvN/nUt4I1Byt/RaFTDJuTldIbfRp8pYuBcC
qu47iknEk5Kerr2fgOMBOL4qAF8OSUy52yrjCKw+Gp/u9LIPPnJEdmdvWBKdcS1Yuiv4IebxpNA/
j+fWANGScbJkY9vBC/TUZ0EfeXe1mBXlST6+bJXfqx37/pRiZfqzVQwdhQcNwAvTdgYi4QGHko7e
izyBU1pNbVgE5+QjnwodMqhApdVk+hzOBqHavE28uoPZB7Z7untrt7hXat8bkwxgHDxE2uydN2EI
k+zz+YRYkPs6084Ou+cLrGTCmjH0df4KKQ8TyGQrsWuMrtwq5bO/N1ECIx+ed/RewA83/SkN4pgr
Kb2FIUqo8e94noCRR9JDXsE483TBsR7duigqB6qDQmOwlqn6//Jjy39JyqUW/b3dOxdNmF5QsUQ3
DMk2+FJVr8PkEQqUvNw3SGczJb9cRni4IeY/gU5bschXctU9M7+70dpJyxcMUD+BmhDX8l+urVAI
iczAnc5gnstxUoQRGblzxtQbEvebUlHjhqYVIo2NrFxxbbonKOEmeTet2PnaWtHldzz+T9YJ4FUX
TSKhijOeZYl9FNLk0VbB6uR9FME4ArfDWkXWeCTWMKi6qBcFHzOxZZYGk1eJY09ezG1pgyu7k2x4
IAmT5PvHP4DKQp8cBlk9YgkeklNpTOdzkXbQEzh7AHT/e5jRv0K/EMTIesakhaeJshC9BE1gzHKQ
4hsASHtRyPHp4UJ9Eo6X+Er+gYD4wI84atMgZHVVa0ZTTb3a4450fjx7zEGDqYNFamSa2K7/XUpB
Ha12nwlsHavZLiH3eqBviZ6mGa0ZxpQHMCASzSme+t2aA8Zp9c2LkRCkOYTyORHX55t4It3LQTIv
XMX31Enh08nRNU2G65Y9bV+Y9PrGGgOMlcPd8R8mOGDpN3tNPPRof7tKBttGbmw0IzT/cuj/9pWC
omuZzRr6dmDVkZCSP+9qWDTfp5U8JkBry8YqmQ3wR/rF5oaR2URNMawoFQVsyR7915HeYxnfM/Cr
QhoOMbHjf0LAWarI4+/WfvisspraT5dw3jxxJHmdujANo5iXgULW4KnAkPAHSlEV2ZUsQQ6PbeOi
bikpG43XS+C/1VlqK91ad6w2nshC08nwGqASAb53hdlOKlknzzmW1Q4r3pTg+IDvAtmmHSQ/BYmC
VLsvZFJRAGglsDk9+W28D44+ePzMG5G/tN008EhIbptffpaY/v+DfQH45Mw9eP1ggHUgyW9dwh7j
tIjk/X3o+UfW15zPLc0IAoN0d4YKw7BKgKhrkFfpHGIfPLujj/Q9g1x2d1zn0jL41ItwHoB0vrgq
yzd8n2ncEx0qpNIEa2qvr03zfz/ExG6IEerR0L7XFNrruGMvB983axvxOR3gMNFy0HI924nORiNa
hUxf6juUFUe80RPXynnXdmIEF4x48jtVDNnZIA8hlzYF7m3qq4z83EIrrgeVx3QKNHUsSDye5lDi
e3u1iwpAgS3bdxLvTAW9Y1gEqyfOTUa4G/85XOPTQhQyXCQkcJDWJXvvuU98dBF0fqdWjvbe7a+G
1UpjLQEpQB9ELS2OAyje2lWRS3Jue5l9kTYkDx5RfK0mEsPlktTmBzeKV6OUuph+KHGXHx9aMpne
PRbGtvOrFTsAfOutiUifj/VCBnAX0fW3JIY+MCcuUs6EqxC2RiXe+VUsTOSPMRWjkL40Ls6tFB3P
5KN7tPybTz4nBeq5TkyMVHeKtXIv3NMNaryt7aWSHTWDtBEcYMxmUC0xNrcUGVORhXrd7o8Ks8Z4
ORUu74f6QROyD92XUBXXxzrH5pUep5FeqOF1WFc1ryVyc9pu9S9XA30zQ+N9WvEBeWPvKswSD6AS
OU2tcLU9ueZ+ifncPStLAV5p1Ja7zyOmANVncMdvm+vQUEjM0/f0cX0BY6eXBuY2RNgMqZa82wy9
6xCIkeYyB75if/w5eSKaPGi3PRq8CWlTkBF9bUGiOn0kI8aEOZbJZtz8cGdIZyj51k9BKkJw35sN
tLZvW0I4c7cZ6/+O17qJutu7cvfeLKnNOAOydt3FE30aJIJ4EDAmIKfZrxT9XGm4Ux3jyx8tb+MO
r1rTBjajoZzMG0T9Gu46bLnr0s6ytWe5aKri9C/s2DU1He++BpfusJBM8Gf9TZEXWozM5rA2etnH
LIdftDM+onB1DJtrkbq5MdVdLuS4+ggfdW7gq0xoR8m5IQSKmPiV3Bn5XM8lP20ONdJIIPW4jZn7
/GD2Q2W56MRDkHr2/yOpdO4sd5RvzZ/SmjGbdTESqaMqQBkvpOdfTlMF5J737qAvjbwnrqdNfIUK
BZATdxkmqk9l0I+eu3Uf5yWG8Nd8kUDpeIduPiPR8QYjxHaVoyjqYfyYIBf70Mtp3cXWbmPM96a9
Bqt3AI/gbNUlwZG4S4bRgb7mXYRbspJRAIs9x/Qv/8UIOl22dGk+WpGGHVo3UMDeT6kkXIS+j/Ci
0+I5cxaP1M8KbvJPjWd6lQLTh04tY49o/GvtsbN0VGGD674kFbPFBxeHHQE9tLRrYDvZmgmd4emq
BsUEedZNKT6cKer3a6he5Bck4W8u0ZCxv/8QjZjOq2KM6AsGsfh0DZ3nyFcXF1VmW/1mndhzZCQF
gO1AjzGlg85oKO08A8EEB+ldK8wk3HV+2va/StpXszPgOLCNM3Vnp0cDe5RI20y9gsxDPBAmxaq/
A61uvlmMGnvvtup5H39npI/ye6UYteW9My7cQXNWdsg5/oyC0eX3eC1mAD5f3UdeqHD2JKQez8YC
YnkuTpWnlu5JaX2ExmpMZ+vBrATtqjgpWeB6goD97tpAF0yMKGEaGqFUI5juhSSTczsyWxpKZKYg
KOTI6gjqzl3k/hyIvLH3Fa7l4tqabjlkVF3/gYD2ba7KXZI/Sgb14Z418PSyO1UOXMFXDIYXhd/B
4YZBmpxdQfRe2M+z0HADvjTKN/03Iqozji+3Ax9asy9k7WUrROLS6y/uvTp+rXgFTomHNnU/fAS3
LLQB/bBeQisiHIhvuzNTVqjKqry6nO5/pUCwISg1QcniGKpOTXCyhw/89AcNQA1VoZwfzWvZP7xk
k3BEVblCCwl/5lMAPZIsihUI3SZEHHyk0U73yShpZX8QhMc1hFEVOwM0T7OxOcrSE8CW7LEhl+YC
T2a8Dq7yyyohWOBjAykk1nivVhJccJTMmzRGMIaUvuscP/3Zn6Mym4+9slgGT6/dsEZ11xaTKwg9
LLRVrqZxA19NTc74lTtge2TEGdznSyYHnIffTK5jV00/ykQpzpTALhmgZQ0AC5CxizTNO0oonv4x
FFwp3gxi//Cdcol7Vugz6EBRnNQRQuZ/oEB8YgGngJHmkcNm6ZfsWlDyiY96HcgcAiiJ/NsDpEaX
S9GiT8dMVz2SygM6BEdW0SNAOmW/gwdp1uQG/hp9rNp/pxowNNHtRPgUdJfIJpePDrF2FFT7z6nR
lyAmPIP//G+P6U6dn5R6lcO8kXTGpW2VEMIMMAuaNaDvRt7guQ73r/Ucdr+8VsbKhF4yvIc6aOzw
HyVcDajNGnjL58IFka2MGHamxkpiPM4pAEU2G0UV+Jjq19BbLfMeVCPC3H1y9rrD5RDqOyHQwexN
c4TEb7WFRogkRJiVmbMHzqhsXlgvjvh5cmw2ALvhKlLtEGbRZ2VCy1fcHRSgRhgdwGw8tOIjhsJ4
E98U/RWCL8ihO7cxhxzsR+vXJp0VRQFcNAc5JHZhJxmQKWml8LUQLOcGrg94o4VER9yC71phvlPt
u2852Q5iWu5w3y8qrSCaxQjluCx9X/WpKlsvpfMBAWOd+2J+Iy7UVCcWFMVORRVAG+Ne0vJu0wn4
A4ZNt4CNjRYRZ1xSn6yWRxJ9EARGc5dcDL9pDDfb4S26YyznLfE82VEDwMFtGyRAEP9a76B75n/P
IJgSgFrjeUtoNC6CdIIOkUQVZHl2hTLr/4Q0XV1DRABXznHayVzBTDXSTJRNlvaAwr37+KeNlPhl
NGHSkYtcyGMgirZMzLdzWYvr4UfNTgUP+2LHE2yLO7uYmFbdV3m1W8GkJKxg5sCAYAzDFldz39tv
9hlHwCHafvLV1cYMzivh3QwHfgnPDLKRA1K+fGXQkntHNhBrxebuJIasan2NaR/bvQW40fpO8QaN
iH0wOWcd624EjLBoVV98In46dGP7U2RrrieJAgGgv99fvdvihiQrNQKafFEcX2S+4PMnFdiXhC5y
9jKiqcOnA88HHle94otLketFNBJkf58m+X6huy+u5gdkoFFJ4zL3pjN70YPjMHQBEtwRm3Xd7wzz
vKqLzIkFogY+GfwUjrHr4rggYR6JttxofqrxBt4D/MhwXFv4uMHtXELkyYqEqwoFeH1BZwqQGPkg
OMZKoXmZerOMU+mmDCN+WeOuRI6IA5aRbwdNy02hMjQbPMXbyeriDL4N/1hFWOO7Ax+tzLbZ/igC
SL4uTCSmUgzV0vLV62+lczw1El7rbE7hG6vEuQ0rCJbW//2M1vGBOqL9QJAX2JSD49P+jrBp/Gko
bZD5RSATE/nP86Gmdx53AIDyuHP1umMpHTYAsc3uCXUFAYb4pOpd44DENjZOrGrqo5TuXKO/7uOk
Pl0io69+b4gfpcMDbXUkCMyudUCFD3sSyWiev1AtEZFY8vthYyCQskMQ+myBvMYcP2Ba0o0nxYvr
kIxEgJaVVtXE59pTzYpGpYNyPCoBUaDUWuIihZfA9bGexolSHQFHu4DRZM3OK4fbYFug3bSq3i2O
CyiotOQEfpnc2DDDWFSYIbyKDicr3okC9lqFluP4xqre8SNYZvx3WWpIPJg4omdF4EgQZjMU3GfU
cZWezmM1eIOt7gkeExXgwTiMiBj+hMac4cLovojMRcZVRf85vePpkWIeMG1+EGitr1tWisqE4Plf
e4FKkIePSzYK+H+Nv34Grqaem2qIMTnC6B2p/Mx0klMltxrayKbiX4TVqmRL6u36Zhh5STllbp0y
0GKSLC247iC+/OzLnRJi6L4+UN8ECGm+M4AOpHDhjWLAR11WS/bb/5gMaVm9HpD/yD9+b8/WneKk
zghP7cyA0s0+d84BQtnGDgHQEuTq6SPE3sBp+GddBzAFRlBLxC1uE9PedOjg+sObXA2UUIndZ8fS
vrTEwDdcIHdpgzV2/fsfI9T+gv1JFEIcPp5I4vjl8dHvwLEeZLYFv8/njTOVLHgr2tYKfHN9ryMh
j5i1W0z3oe5/1KDVvV2NfyGMvvFmY5Tn4pW4x4naY4le0sJ+2MzgE99U+ZX3mYPG1/8fMpQe+4YY
BMThhNPB1VgzqIWeAWGQsqyf+9j31qE/1qZ9EKBzuPZGHJckWs5RQbUqUsf3D8f2KfzXOrBQ1QNw
wj25V3X0A0ZeUpT/P8jfCNPQcTKmebx9cDQqV+UVuiJK3dmLS6kyxqjO7HUlIfd9PBmTzYnztOGH
TV1c07ORVJZNsuE+z1yMrF03hTK5X6wl7Hj2I7zZM0jruyIuVZsY3dtqwzx3IELTlUhutBnSnB8F
ZgKjyb0SdprXBQAvchO1Gcq6jQBJ/N+3TcYhMkIF82LUh2tg8C2uqyf4iZSIGyf12I1vQJkzt9TH
1MgNgs6pU+OGWIRk6xuTg4VSJIEurXPv1Bv9qGCyR+IcN2I2vdxzpu5bTvkao7WaZQdgkMuW99Be
ATfCXMwbTblyUDSStOR7v+9xoEaUroW8b2usEV889pAtwClzU+SDHfWPdk9TeTHVQFrnml2hh6aw
qKVtKks9Z1Mg/ptuPll051jh1Pp2Habzj/K8yz0f6mLRWLvoba9FQhPoWmT90e7PUBdTauMYjBT8
p3ZCG8ICG89sMRKsJHrQxN++YrIc6lGGEvyociLvzicSzi6GIndUSo1eGXPPZLa/OELpXqH6sGD1
5zXIkMOtkaK4aNujAqyGGUP+mQqYjnZXOlaNIaI5W/igz8+wfYQckoxkGnvQNoBvBq0+aShKoCPH
osmm1a3MsG4CD2JgivM+hz7WA3yyCcTV37Ih8XDyb3EkEiEsRLwlfx2Yk7MB2H3uO2ZnBHk3813P
utEqFu7XWARfB6aZC5hQdMUcFl0uDCX8x7LRK0xy+82htXw2YlaVOdq1CxLixxeUpsn2oEEob8zz
moeb8e5etfBNHS67eTWjjD+ipHexGicxhHoU/cHDmzcPEgdj5N21rINWZ/ndnxeYKeIl6kudVmWm
CjL4wGV08uBuSpNBTpLZWrJ8V50+NqBgtxGIJJK8Nx8GIrE9tHRb2xIguo3JozOSWabEv87iV6yp
76RXRltAPXl/XsRBYIrJZGj/Yf5zj2bvsr1WO0Bgx/kbPhxhpvMiUaPAakp96JNJt/0gpXj+KNAn
4zVjpnerGNID5lYNlAFyiO4yKVDsJadD6L+XhHcLLpPsqqLwCXQK9GWK6U9q0omG+AULxhHlNHQq
Z4AAYm9f5R7SkEq8AT7vAO47kUAWFWA38QZM9dxdOT5jPZRROa2g4LrbsKEGcOWq3WatuSMP1vVT
7sY1PtYCo++CvtwPoEqWrRx2VatrfRG3UtgFvVMBbJz9oZTIL/8uAM9qdfQge/7SKUdwcPCdvkCK
4dQyRT7Wp2fOI5xCpNQrS4WnXKHUABLMmQpjiQ63X+64sX9YYNaJJS9GrloGLyiKNJ4LjjNpJbdD
cfeMoierWsYFZSFLx0sHmRhAxB+4fEt7DT2fNUJxsYPj37G6qbco3Z8uG+/Efy9MtlCCRv5JrElV
2II2yqr9AxqyhM4mCoFrJAQcDYvHKV0/L7UbdCfNNPirMLOcyCo+rbxkmyckRMHHrMy45sxHKtur
zElAGqCgOAkJ9sU5NmByLOwbRNno6ZhfF7qyUB56MDnZTUCukjT22mp8nZSXdI6HfPtHV3z49zrc
CEzLIiuMO/ZffVc3mompDOluWfyWNgWE45/+xW+nJ3Vpv91Vbd1V6IvYGDBfFA/YQhq7VRMkY0/X
Lhw6/tm/LAU8WOOm/ASQhzmAjs3lPoLq4c14CFdTpMvSwsVvvmDUlhIt2UrXJxFrJ1qteBsS7RqW
G/NOExX7lSt2LS9OczOiQVUAWkmzvGk43krff5ijy6+NSq6g4+K6yEXLjAlvj7gDxI/9nk/X0Rgz
PRLTbRVK9dPBuZO6lyfO51SsKJr2H9B0yvWux+h+8augApDxPzQUL/LsWYZ4bZgzhyicgSm1PRSV
SOn6EdFvVz0QjYdRILAtpiOa0YkrVx5+wulKFmdwhSos+4bAXNfUyij8B+hR7UgGq7wrDrhX6DaC
9dCz8pqqFRr1JKoP1SgNyL8nQVPmn5lAJYDmGcC4X8yJj3w6kwwm6bbxlCDTAbqIzWyyk5CrCIlL
D+tFpunPBOrYwn/TNACsTuAqcEtgwwFK9iRcn8eiWmyWdHCXyzsaJzznjtw7k+BDzWU/WjOdFA4/
JlngTuW2jOMJ1Q+8OEWlu/5hzdSi1UA0bBihO+99uxhS7lYu2u2E5Fh8uiN/XipUTZESgmfUnPbu
VR4Amq7NrjrPBUC4sG+52NNjZWCDVVASDo7l5liZF+KdFGQ0XUIdkkYw42ub7aoaV0J5d6zbAqhT
/6tRLICkZtAl3JjG3cBbRmH/+cTjfRiIvefdUmS29QGNuzR5KA6uul1iYoS6NqTyWxblqUlTyyJ+
+EANTvUgLd7sdiGcchzwmSBn9Fp8brRhxftktTMhj3CJdlYSF+Cd6UqazDwf2SkgCfiCUjN2M/ov
JN9+CKwiRuIu/jFKpXyiaXF7GbdNGNkRYXEkHtMkartAQoV5CmFTBPA4K2X6ZoPSu3I+QAoAMsgG
dWN2sGOl8tkq7OgCwnYcai8yFEoOZR+8qjh2EtTgR8HiJYS0LIsLdGyp1BHwuyxRhM0H0s/vz2FJ
wbP+wC1DxE2BqOZ6o/zvil/CXvUQ0gvuNoUPtlKggTC5Mfxo5sUg7qa/hBiclM91Xyu4hvoHXcbX
leWhlcorK80Y7Y8kxLOJpq/JFO+rT4hkzxgagq8SgATBhoCYEBNHBoRkBn9TMUL+3xZt2ZmONHXw
s62Zk64bCmxm/QrKdD6hVEcOOTQVSduGbyf2fLDOHWR3vGyhxat8TLB4wBAaZTIDVBewQdveO8PO
T73dwCQm4CpTPTy4KeambX6JlWjQ9nULxsDz13y8nzfL4MWkg7kL/D600qBBAcUI+G1iDpSZJ5ka
8JmaJF+3q6CiiP39iosVPGR23zGYq2k0L7AgbDQkJSy4BPVPcjQzVnxBKRu5OsYmMAzWRXLZVW0h
RX0YOFFKBh2WX5UqRkqJhaiZkmnNQgMIPnoC1ZS/n5Zl86um4nGGT/VKJGPuPmsYhSBg9hFYgkOq
jjgCzk6OKvjyJSvPysZRA6iC7IedRH11qPhbNrwuH5gsDdkevwB9PJ25C2gDXPCPUrkTf38jzwVc
X41FTpxjJCJFSSlmC7I9WYgo/9ARGZ86aGxU7hKQzRK8dGmTvEOPLwbxPn9ZY3k6FsVkCi7Kw0iO
R9FDHPurTg6+Fwa9PteGxwoOJZpLHEMHZiAZzWc2JlI7s1hJKBUw4tsFgZe9idLdCif2cxTvrd0Q
78niJHg0A1XCdL7fPylQeS3HwszG8hKMjLCQ7yzJSxOf6m4fNpXXCYT8h4iYZbS9cRu6C1I+yTGa
Re7htenQ6NXwrwFXLy3s3zF5pDV9o49YoA2l07AA/py60cc9dv0MmS5Oqd58otNnC1LgrWtW2Z70
7wLLFEKkBtd8QrSl7ygFqn+sZW3frihD9T8t7MTXBCAd+X55PRarLiUcaARJ5iisU8bXGduYIoHb
22UTSFWhFFSaQssHFXwh+eF1IIuAvkAW/9se+WgGhR+xhHsidRo+u8teKImsvTympJyLUI36bdQN
sFuc2fs4MXUYPYAQocUM9cLluZNcU9hqKaO15IFxYqyVBt87qBRWRkSCithaIzFOAnE5pFIrBXcj
XgMZPmCQAam74q19JIeDUDGninGEZEAKkU6HDIXMmdwAssAUfXGorHZ5oKU6C1L/QA7vcWGeJhGU
AC6N1iyT2TfvrWGe1E6rTuJiXj1YmVt1+GSo0vwA4nqadGYuDfUPMvCbxg/Ixhto1Pd14DN3YDGV
zSg+8Xeec+8mTsWgPI03w5J7PYOFDF8Y/lLR735BevVlspizEe91geGN8GHHbV0eq3ba2cAFeKqq
iaxlw0a72NHdzHCksuuEq3A1xtq363P338WzivASE14PQ42tNMOvcoGbpvlTolO91bDAXcqWVbXp
3D1M6XwcVHDHwKPqpINcL9RCZv8pnB1hjqH0ai4DajmG/K1gyMi/nio+ZfGesz79YiJTRKfoUjcS
pGd5/JNHzFOG0D/I1YN+Ju3F3JFkINXa9w6ximtGGREZl7uIc2E+PEJn8n+aCb99B4A+lP8TuAD+
jdtIUjkJaL7v2Av3uw57wSh61ZqIzI0hCNu862HAzjehNWdp5LXKBpUPZtnBNd7xEsoEJ5DY/RCW
3X/YgifmaFzbKAjsdmxSWjb7hFhFu0PeNNFJpkdhveFlwXBvdcfEg56JBZsKhghPDWOhbR4Z8568
UdyhZG4wR8cFIlYfvRFzZ6LxfHtfvXuI0iF/kwSEG0fsKovUAqqknK6KrwbQ+a5PuTSkrfEmeLom
4XuSJUVGmkX9HGLzLgCgVfV1UquJ7fApqaWg5QbzNr295nw3TNkNHLhG4+1+5G+QZLViaHS3Hyp3
BdFiZMbYniMNvewM+mwDX3Ge54QkmugoQAgT+KzyszOWgCXvVgS+0V+UgbbXDetvYrtPPpx6bMk7
FQHurmLREeIrJolQrJ3xr8rRf6faMFqwYWAIYCYJeXVB5Ok6HW/N0pkivRrEG2ByzgN8mhKWuhiE
QSBhzJriucKI8nfZTJwmslIzzyCsqVtOkKL1wx4uhlsgptRWqWZjhTjEw5Iuw8hwBE1LWO5Pvr1K
/X6SJAIxwALmPVZcPRxQadAucUBr2YopVmVMF2MCVTM0sQF5vohqv9tNoIVWdb0RbILUu86+OkHC
NbfCTmmsdyqZDdpP59H05Zz0DYBPfov7XAL/w1DnMK96vKdowrO4s3ihKrs5+5Ct+9d44j8K3pJV
MPhEEIqhmem6Ytug5TauATDeW+9tIX+8dbCfUuiPz9yaeoFOOmR3zjRVafl7cTLQDOSIjUY16B72
5cWf0jV7jWEgPGr2TkNYrp1YzAo2X4ewI0wuF9xt9j4v6dDKe4MXnjwZMeZsnIEjviPhRa5kLCof
as6zriJlRb3GikFug12RP6rzN/lREarSJY5pg9bbimVJ8RbIXzg0YW0MpQuo5c1a6WHii69nh+E5
f97vJB1hUHhMt/hAVJi1NGk4UBSPmdhL9S0A+nyAtGrVFI/E85x4PURLffwJkRJ0z+g8vECOAbO/
TiYb8Ify6oyaVCN/ES1jQSLp7bGhWsA8hfKgSnxjkFRAm11KKIRHK5aaeSOP3g+XHvXh7vkHs/gQ
+3Pk5ueur1q+zM50Gp73t8MHUUUf0iJ9jGqKbPLrznsOe9adJEHm8xdp7UFY3JpsUTWtw0FGUjio
P+OEqeL+VB8qWVFKciSvR03i+a0E/OJDENMFi2jmD18qgGqoM7A7QNUkTxIJyb/gMiZCLPGAqucV
PgJlQa6ydYJ/yLSx+nS3OYyklkM2UsIg9hxG/icxzl0VuslckwIgxdA/3cjE6B4r21gHWPmTpK1p
45tND0LgU2GGa9pBeDG8w71ezb8Katvo9I3RgGrCOz/Eh+liohQnauVkieROfYeVlIRP0cWvsAP1
sI4uTJ/WnC1gNafmM9Tys0dnyAcYBKLiinFG9y11fqSvrijlgYiuMU4QuhAGJjXvY77nH/BQklVu
d2GrcB6/B7KfUBECi1ayREBDN2eMHFBTkU5iCj3eIxtnw/Z6+by+M2eB1YNLGj2zpZ1C9PpSHn41
W+m9EVUDOspjLn+a3+L20XOuQiq8YAvsihKPmoVGZCbm8MukEQzDPLa4WdIuQtHvMa+PtMM7+ApG
BYPpuK7bZT8Lt+/kpmTA3DVxjkd7XbI3Q4NbDL0b3zKidYJAq+M0YVlsaakguetl8dYZv0UbxOd7
LLIPjIcC32ZeWV9b1er1NQqHx7cauVb3gIMJDNDQOYnbzWypEZlDDS54/OJ/vlwn7NZ2H2sE2PFt
SwlAI9UnjetCDKGJP7AuYtoKa8GUBoDC2fIYkU0rJkS8gJrRSSOL2tPsdyi4UJzMOF+f/HuN6Xg4
/P386a+nyXa2yZCVEHCZgMF1EGPGXei7i3TmUIzQ1RZ7ss5n1TYhBfvF3FnuqSk2K3j1LNWQH7IQ
QBGS32nIB3x3nhU5TrySh0GTPixIpO8mjZyC1FqbQnKtojzTnU32/6OFmCHWqOWa3++qsviXSX69
dQ3mFX832GpfDomCdqw0TToLOdYX6bpw9bauvQVogplu697ghoVMqSUPqowFlCm/QvsSVHXeGDdO
+JUBwDUG8dc30UmgDpAJjpnb4hZYlLrdOMRvBLVMj96/xIss1RYfjgxbe4Zn4LI7nd2ksMOVWvgA
le1wR3nxxnQxo/bUshfROBrZTVK2znhmxDcu0yM+2P0KxsFp1Y0od+Qfsgl5RoY/EakpGdIeAg6w
RMLAjftHNvGJTxP2/wRHphGF3aYJJ8Kmd36nf0qVcpRO7eU+0S/1dNymOlYToDXf/SyJsFW/eS5M
IqoIazih3VLWO/TumG2UjIAun+BCI1qtkLLuC5cK2naNLfPxK4EfsXQmXC6xFw0z/lxA/QKcThuK
e9hBGvW0xh1FntN39YEs1c+e6o+vtgs93WwF2FynmMxTiC4gqomY88yKw4P9H/kJAPdGBj4mhKhE
uZKQF4oYwyUwD0LrzXDp/yf5rOM0S9MJCimwHd/ZyOqgSIEOWLxN5PBFAYhWU0LYWw37wcOpN1Ef
c9ZD/Hwai7lxauxTS2UdGaupk8aEc52ei2b9tvNyoewtqdAJTjC392RJWrHplpcwfLtkJdXMGVzV
pWhFFhG6dY7TYlNItx2k7mRZQjRRyqCVtuTqQ89hdxppLof3Ny7mIcFNh1snNk3VyIBS7brpsL+3
Xg95hbY/fwKWF+fwrymPFccMGBpRJII+7vJQiwJNz3tcwn08XQow5pheOa75ka2PNuJ5weEUKVc7
kicpX7Pj2NYngrIpp2S4lC+0yi9s/KzFyJ1813Nc93ymnaRBbBFIYKlhOuUC1kEw6tJ9ZesXHWfd
6JyFFOjpvmn/uEkYmKzMZ7+PBfqrMmL+ZU2YiCSyzxibxpeS8tzvpOJ6QVObOTVtUFvgsD568/uq
qou1EA9A2ha0vpKKz6sFlpr/fUTWqQCavomwNCPsRutzMdl1yJcKTO/va9lIGCICR/81jR4TRzHL
cu2f2o9EjJ8NYcu954BqR+suSXzJn2XZF1oYimc+VsvLVG5yQuc+o4wBDYtnbqT3LCP3Edwnc6u5
RITRzG6yBUCMWxIM+dGdD43A8BIzbhCNjhn2zsiPWZeuJXXxRg4E9/rx3N/EpjDD2qzh9+CNxLjV
234+5Vb9/rMX9cAFbHyS2UWGNEKCg7cOs7bn5/7+ZcRnDivdLkpXGQJBig0KFC99GbrmMgewvjL6
gespyKux71PxPYH2RTnV26IcNXoAYBnwaOROfkfIAn/ZSrIAyjNcoiF4Ur8PrH/3lfQbky07pYLA
e92Emhz9pwHYLxJD0vgMhrDk3fUeqsg6U6eeqLbB26vcUktQwbnrrX1QZRT3zMtue0SM/DU9wrPD
Gy5b1R0Jb5xkfVNGRclBpAuU3SsZeps8FlzzTLLB5pVdeTHFbBNYehcE1eJ3G6en2uLYNOShzdaC
jFugdHRwkrpwee2FEJ8Q+F41HSZ0oqNBj/sRtpG8MteneYk4CmZS0pOgFwgx+ktw/VcfsIjwFtc8
uAS5i8d94LVSmL/WI/Cv63USCeZA6u+9wWN0ZS1vJiFLayIiKukU9W3ISum0u3ROASK8SounxpZO
cK9Rr1ebbCfs9v7V4YECHTYVpJXCp9FOoJy/3A0hWxOVXN9fqMSUNgWh6ZilkMrGpXyjNVqiA9uR
z+cLMzhSLP1k7UuVnYyKreWEWUxhI1LHmyky/6G7N8JiORuI91E4k9zfUKEYcT/2W5Y9ZUbobdjJ
iDekkUyQUjBZj6tfPn5EHS2mnCmMsNeZmlLIXA9qEQGXu2ML6o41ex+tCIqM2lP9dHNEiR9qPdaZ
cg9RMgxjLwtyXs6IweuWR9uYYSi+sCx7i2haMgcBLZJvOtaw8UIgKkRlfVOzsvcY4KOtRyHFgibe
Mt6IeNznjPGu6rwXQOMpYSPPlhjs3A/igGWnvRF9iAl90qda/8DqZ6tBjfb8EBtbyq5pGDl/Z8GV
U8xF60zCCUo9zEOLcgfBLIgXUASUYsJx3MtbyQWIjAbscOR8hDKy9Vlylk9YKz0AJyC+NFXdmUgY
vMLmgoCzt0+eVifFVwswO9AeBJN9bMNto8+tE9aojCdGBoghE13XTXrJ2UMt/tkegjcoOgbjQ7+0
9mVSOhjrTXwDnC/h6WjQDDITgmiNz3gAlUt5EVUQvh0A48bccJv4bjlsyPKwvgVWaAkcLXleTHZ+
0DVqJSk1WK0R264aig/v9N0VeT1JBCPNdPD2AsDTyCTfkxflqJ3o52pEmM5x5naEKvG38sRu1PRD
aPB2WPoCA/A2jJT3mp/H2Q+DxO2bWQL+iH24eDajg1/xfoO0erXJRANiHCpH2xR09sxwHr6yYsjm
SeO/Q+17LoOFaq7t8welg5rK2thImdrN9t3aUf6l7DFZL1KXd5y/NUFBenlFcbCljPzs7XOI64qt
DGwimUUBBIkRvVVmPXyPS4bpmuvZ4H8XCEMXnJyfWPio6RAKLl+dZq8TwOHgAwUx49LZpWJ9NZGb
xpQoTgU9rh0PBf7dlxPeCvufzqxgJpCmMVLzfSMjCTK41jqxjt/z1uH6nDYOMZ6Z5rwTb5aNZJ6j
2aCPnaZyVE9nCXzZ51QlkGlVhvCYT6OHGkz/uClSm84VlOnwof/lbPf5hSz7IRb3CPNOq1ag5lRm
g1PvllEPJ8CXJxtn0pmkj34XgLBYKoTvNP9tZJ8R09f2FuQtNwncGHX5QWOGVnCu9Kde8e0BEYaG
ebGEyI64GkTMUMazq/bJWLMggyWRqzibkxsCja3Lg72jRBo6V9TpIq6fSlgRShrvx6gtv9NqntqN
EK+H1qrETzk6WVwhi/YC5AWK95M76DYe8Yp+F/JxD9wP4jPRExpBKS8hV8PT1AI/5buI1nxrxcmA
jVxLWwAUkCiIRuEMkmo9mCOzRsjlWd/ioKA+tUku1eTHqmCfYgGzyLAXEZiqjdQpJnWOdUdZ0xFT
EdhL4h/zsP09mCZyBYfKVANRPpRPTTi57XYj86qWX6ZqChNiup00JpzlV9Xjq0ZRRscnccvuWVj4
9jtJ3HivXORUpU0p+LJtIeuoQE2N74JZq8k9qTqQuLv5Cn4Swk5BrK/jEsGfb6kDZDDtAODIymTe
en4epvxSMUXwnCytc76klh18xTgVBTUJ32HOBqUn4MfoqJodpMnIUuZgKcE1bo0fcrb8hnKX+RoB
bWhNfA0UXrMjzch4Ao4X6yPhFSdkbuEZmWD/zTTq1gjkZWCUd8FWgB70nUjZCOjI/to8WXOBYPZK
vUVzEpImxD7QzhFMQ9uxTsk6qqsJHujoXvSC90rzIbRTxCBn8KTj3PsXQMqgoyjoTXW5i9BJI6Z+
noIHT8k2Q/TwGDrt0qBKcNmWRNv0binDwLP1F3sd/lFzgFsV0Q3gQIMAMAH7isKsB7Tq/4UnzLcH
ZlTuS0pGQuyOZ6vabA6RGHCtY4D9/qnO9j5w2b3u9scsLmIXANj0TMVacXVN73PzpyofdD4TaEKJ
6f1goPPtoEvT2acyZ0oDCEC3I3NMg3ZfsDkishMxj354/R5hGt5MZJGZZff8AfBY1omlsU1lx4vK
FOa1sKxC5a0id+6MXIFoz6Zs5rZmgPDrf9a6sEhbJR0K5MTzwFFiS6yfZeciCCJbxpHgEJiB1pQ5
/Gvc9K2bFAC8gIaHBMdP1phv3opYvyrqBbm1ZtbgI/qdhKT16ETE6ImecJ2Yn4Awlb2jN4Si6PEP
pDXZKXn1XfxREcrNh+pPqCPv/C6NM1HePmw2+FBax9QXBe/KoAQQwGnLea7n+NRGlGHO6X3WjWPS
RszTld1+BF66JJfz1sdyrboE6c2rAV7+1m8Q4zEdzi3gSXcTzMLk5MC+IQV6jdQejxh4Eb74ZvHp
N7u9bXw1MOh+HD16tdjBCIX1Aa5Llg87avlGfRE2ac/JUovn0Be9y9Wdbh4rlYMY8dUFvAOr8jhq
pQA83cJpLVgXFMsckWICdSeIsaeLGA4pj2oJc/5mAyttwDJQqi9U8MkvaqzkftI+nA59oWiN4zp6
5QRPOyj0M/PrAVhcoowUp8m8AaXwQavclEVpWIWkizeofKVe0BOsUhnIeturfpabUzjUtNzv7WgL
JumwrD/bgcg1EJP1dxcQ8Hjd7Cv2J/xaqcjBveXffa14CrSkocXpFC7CGhJeiqvM4CWO1Vax2NSL
pEuuYjJtW5FC/uL85vry6rlC8m/6qdaGfQpSJ5v33NmgZgO89mRkF2+LZ+Ay/lUG8euFN8xn7NUL
uhTRUP/mLQ2ath3/MNmlH7N15nH1MFkdI5Gw6d/ERClx2L/nTBQJTC5AJTCAo54IHoDsPtU9+YwY
JaRKigSZMcfFFLK5S4N7oRg1hpj/p0t9MKLdDyCRNypIm7b6ls0vRZSjfs3jXMcd81Y5+72Q+IZX
OrQaOVl+V9KgJzv1VlpEOj17GLEXQFkL5whtP4GRsCPZ0RXrg7dEMYRdp9RDhK/ZSj0m1Yb7WWdH
841/DWGQDI/8F60AfZ6XGurbbblLAY66BG4pwoZrOsuGoUhz5tIQgtb/rTgU4PhVBJayY7GP32cP
FM20bZ3mW/C/KRCKyT9GNQ5Il/yda+7E8fAtyt99B9zk+6OBuGlDYe0itg7o+pFpevE31l69w5ss
6FoyNYPUEd9gIzg4t8DVAXDslPXoSLU7iVg/ak1qnUIHb8O7/tEwecR6H5SBUxLd03rnYQs/Ei+K
eSMDhNEyovpDvnp6XmLtSjGSm2T4G8aw8qEwl8CeAD4HdWpf3WQ9yZb/BTpU5FTaorbpzsS3kJQO
z0u++fmtyUKu0oLtQtOFERYBr6Ef7jR0DoYo+9X7aGwa7hwJXB8CXsaP6H8i1vdZFAzoeitxVzgW
MB90LWYUKLMUJUeYvWJatIU5puV11GaqJGpzhhL3SD/d9kv9noy2Da/MBcvDMGLtnmNAMllDvhf7
0evEDrkR8OnOaxuNDyKKNMI9P1kO76vG/f0j8G7U4VGmdbDKO7NnqOaEauQBBwaJcKPT6sH26KRs
L/jJJf7yUmvLxcbYGxbykpNNRT+YlLnHb+Ej9zcFxslHM9oCdiNHA9RAuibe5PE7q86Ihn+iB2+d
yGXkBRQpIIxxXbTU86zCR0pU8CuhKZPyFWHTGiaZQYIyJNJtVFTNiuWUAwPahH03slwqsmAe8Y78
SMjLVVASSVOTjoCjRDybBWU7DFJxoBl7fyfWKrKVvj819VVXnzdWh08w3EqHnh0WebX5Wi43EDZS
rtfx4uBZxVs1I9eXpV7jquyNXSikSvI00d0+ACpo5RqGZ34gwveOL2iKe3fZaqm7EdXjuGIELkNJ
bFT4CcfYC0v8IkJ1zfQsGXAZZ1cSk6n0Wxni3kxX4M9DJiK99FLbRKaHGyIUG1G+GAqHHgmH20DL
6H/DhXKhCgl9zwKHih9+DRqcuQJzoiFIsT5Xe+gpu6Biivq9H7eBIdPb7qOdyLzRXCT+FmGTApFI
ZjQsXcC77WnhRk3Ed6zsIMuxAtXKgeJBkymfaUVpEPlLVgSogZVrg+KLW4oLih4pEx0VIwa1MXFf
sMp8Mmu9HQTgcm2406ztuw3Czp6YsSkOwAoSmQCKFYigbAIY0mw9IE5eQiqlpuMXUmAaPJsE+iJv
0ROSZmVrVepdSMUBhsD3wB9X8tLuABKdf+DqFU7puznxXKjZdJCTM67ZMp3pQQW5UWC2x1u4jDXd
3eeN2sm0sjsYDh1WBsCTew7UFzAfkUHUYa7fZJ4wj8jYGzay3gYo/MOveXp7eMtkx6W6sfswugFK
/fdgtA/4ksIsAvltOq3c+c1DipeA5yignR1G4bBtTuoVEz5q0oz2YQ0i4W5IjRr+JKNhh7pBe1Cz
H0RRnrlljErzR6bfkunoKpKqBEi0zKUvHhgM9EsiiLlGdz09U7Losz6jZupCOeWaeqDrolkdzEzt
TAl/HkRd60wTWZlbO2YK8m5s908awWQbLo3W2m95ITFGF6OHi1UnBlUZiJ8RK4hqMG6UXxxJ635U
rifdqBL6lN3G8DUaYPYOBB1jnjnbiWVBCHPWkvgbp71Gs1vvcY/nmh4U1yMdDvS7WPTxL8ypbciY
p+2JvnsTcFHah162eDFViTzQuWWZNJS+BBvqJQ07dZ8CmlOrbL9cKnIPavB0/IjDJo9jpIJa+CDK
LZcvy2SKUAn4QOZe5BhpHyDs9PxI+K91ONjFBc0Rfu1hdxniCfkADUMT4LGPxedOvrX6kuIrjV2D
pbJAK+so8A1PdI+1SyyKYJleCWtIR0DAF4lmUQxLBJVTuuXLy1ctsrm0LJu1ADl+ljArNtWNiNE4
avNjlbIrQERYohXNlsFwQOjUbCSa0E23QYONsNhk+IDoC7RCphpLhRKixv6XtgxoXpBelp6kGcg7
5EG7BqzQ8CRn8xOz/DvyEUH945zhI/bEub4dTfjqnMDQlAdZkm6TX+J5pBwu2TxrSVgKBDKdyREQ
I9upXALGhyk2c4Ah3LOsXLDqHDY5pvG/w85rrmYrWdtn/Gexw/FaCpa5vo2FFguuvfpW2cFtEUjB
jlUm3nwpM4rH80/j1DSmKT+vKFCMLN8iVfPFP4+xgvqZ8IKTvZG8u5E2nQpNCmT5fC8HQfjppORZ
+L0306FoKFbB/EUi83lPA2Us64waCfyTATOk75aqS4ZgfsPNf2T/0ju4vbaH6Mnfr9bhUO9BEsa4
wGAwRAwRtmtDXt/X5Pfb8pjkPsC5eS8XOVedxAB0/jIN6AGguX7M5EtNKiYVrg0010B6doGFKM/w
K97x+Iuzg9A2xQw3Mpc3utIgdPwCMe2hJzvhjK7R0PHLxHmgDag9duE6rSP2BH7s95RDrefv3nnl
pHftD8/xsbQelv4wfUYa8L8EF0JSxNOK1yaKqZAQO7+X7GfZIZG68qHasyiFOt4HitdtxT5/zfDg
SgGMBGgS3PnyJdolKgavuRJhQ872g25JVjvbYdB02JpzgXZAReKRZLCa6DnqDmpmYqzlUSVhLGxk
iVRaISLXC65WUIZKP3BB8OMv36rAoJlTQF/+kqZ3Da/A6zJQuwbKdzEe8uJd4swzY+76P2ScHafF
pEotpdlFEzGWeQ4hBWWimuSk+/jPg7EZN1dHThL1tBN4recGISOX9LWE1hu73m38MleZvRlPnCjG
IFbKqBiF6YQ0KPRv6ysD6RHCPgJydkGjrCmd+Y5aUGyALiT5443sC6Liz22gqHl07GBTgrYHaLYu
z/HfgJAhbtOStdaRW6jojLfUW+EzsCpnXByqgz2zoFftYar0BCMXpHQHTeGwgoe+f5PcSAoOE5sE
m/4NuMAHOh7QY3PUgqHOnm14ozBdw+9h44jfxRPvHlNNsRdi7tHPu9NMPJwixS+Fr6X7mt4mn57n
/FkdltF7whRWzeMQ+R4sAhNou+wop6fP8pAGB4i4z5xljpCpARGLZWzf87l7Bw+J0WV3xhp3bxb2
BDKkmtOeBbIxkOattH+M+u08LZJYZwsg53dd8J30bCkivZgWugPBYpFgJ9zya3Fkb9xGtuon8qao
UdVVkSBVXxPvS2ZLxZ4iYh5QWN5Bb52xN0xADApPUxmKFeruvUkruGC8LkCTSmZ8yvaOX2r3fFUp
le2A2hvDgj1DhC3qMX65w9Kwi4SwcDiXMiAQ8MutrFWcslG5HLaztC/bEmaXRQlp6JIkH7/tJI4U
VUBYCkb94ZnD1hR7cn3PM+h9t6yLlGHlG0IxnoFM3QMC8uLuu+MxlMTMFaX3wegiY7AUeC1e3wC0
DxlvxDC76MwghA0FgxQ9d7xFogwmh5giNErAtd3Tr3f7n9+TBNr3bu+MEfJ9tixdVj9B6FYG4bNY
M/zDRIKztSLFP+Lkj9rqOWtICB0YpFw10lligHz0ICYHvB+0dlIbPlJR2EotVyidai8Oah5dqDgQ
zgWnrJxkHdzuBKJoBk8m21GrZcoExwap1Rbw5gIWnhQOpMg7CeyV9LLtxqn0YpeAIdDU9tTZHuuk
De5dO/qblyX8B6nuRLoJe5XSb+BUXRTToW3l7vXhNg9ygvPfocK//is8vabXj9LAu/cbSQbMm4+6
fWeecGLf+qV6cXtIE75ohJOKl5icHSxgWiIE0W5q3F5qiih1psDxPtTyAzMNUCXrNUvg2wiJ6PJq
cW15GNKMEhQatKaDWWLDHvrZlfsL7WaY6jI9MJxwEO/L8oF5cDSHGVdkkuMRKMR586Pw2kYBwylh
BT+MN2oIlJfmDvJHLfN5BShzV/CyavCpmxz6THsG+WmsjYpqv3Z1y9hG/gg75803BL78urKUUQzP
7zlSdF5HNsXtD077Lg8xml/2JSEYEi5BQp1dSIy4fJLcO9N8l0+ym2c2bbVzxv6YelUj/pM3Lt4m
LiGqToRzlynGenJDu9k9mxNCYPptXwKNP3ex7EegQJW0sRA94Cm0i5okvXmyH2IBqs7d9EOZe/+r
iBjnsrEn6V1JyPBqhedvEPMifihVPVOjPC5O8/hM6j8bEyWzQpGUxu8vdBOeK6WSJqUCJD24ckuL
6D2lilgkBmSGCimB1X0CUbuzrkAt/5Bx6jynVTIikwAsH7scM+KPCRx4XhsSSq2xV4QnFptFcUIw
5eKOl0VnsYqJxvYaXke046AJsjMA3pnW0G6hosBKAmvkUTUjiDMr7AWz89FIkZeQ3O+k4fS99mt7
nL3Oew6ICfFeN+4aXNfyEUA3V3aoHPLbh/nNu+NKZ6bg2qkjmVzCWuwp5G4iC61DFuj9fSQDroP3
tJyRqCLwTVuaoiWT9eAXbjvWxhpvxh4uoOBjT3DTMO1GHFHtSdH85Fkb3ZIemXaKs+xRW8JY5H2k
GumLV0OQcHhCD5OngO2QprR10TGb2oJB0GDZO4YDARLUdM87LZ+9COdSTYJvTAqttg1H+QpRMYa/
8Zjp/AhxBM4/XpSr2HRTx0qwT8mkALlXZ+MqoHKg0rexmVFrpC/ji5cfUPzuuJPtx/3oSN7QoFiH
WQ7VCWOP1jgqHdqE4hrAaqBX1qQwi7Bmu68omkh346QA+3Q+mDpdwE8XKik5JM27v8ugL0otvnmk
LMe6uhFccBYLvi7Z8XpvMULiu1+26oQl70f3yl1KsokQgSkRB7EnNsp9PJikXPBQiaijz+RfGIhg
sQZCPTFtL34kGC5YbsII7k6AZPbrKwF0onArY0cNcDlyTOBFpf0rJDFvq97lxAfzHrRFp3qs2iQT
fogQ5tAftKhIv/Rqa0lmj26AUzLTGOdIxnLLj7+puXSvfDaPAcPSiF+zA8lcT0++wXWpP/cQ0bFR
az4pZ556H7+FaBvYNShWnmZ8yjgX8cCBVihlSVMjhNLSmBwKNI3h8TlR9k+9W6+d6E595Jyk0jJp
p7kGr2ZMd+Q21ddsMKm+u9ZJlzT/y5F8SrdYk5MQGEYKP5JR1A+fKQ/+XULksMjGm0erkZxNJgxf
ejNvmgYBywyViulHgnA+EFjSP3JZ6+359PoRXQ7Ewc1XUZxOy2AwSaf7dS1yMLdnJb/W2DR2owSS
lRMUQqvOPpS8FkNQJ4iHSdZlY1yEj0GoVCJDWo1+ZBvgwrj/OOA2qckj37jDHyngdem1wvspIls1
1lG4wd6Lr5mCoc5Kn9qfsa8VV0tMpaLv3YhvxWrGRBX2xCBxHJYzYSOU95G9ByiSEaAbzQxZBuMf
/MEpcTwX1dkqSoEyCoyz/S6SBl5IY8/cVWKUmRHW/Cmbx7YPtR2X4lNueuMQf1bN0D55scAqldAu
5BSxgvIgEho9Ys9eN1JetQECfgdxxoAxNj7pvKWjQ5iDRKZzJp4om/oqEn34ZYTjazbtS4n7zdyU
tjjyy+eidMKPtY/6PBcekxMm8TmQZUpzW8BJi6ZdfLNX9iQessiRSD83/V9uWollKMrZvk+xoFgU
Xw+0IDPoWMm9YDsW1rmG5Aw4CSUB6JeJPl1IkfXt+5qLCN+utNNRQxtc64YKMZf4HkkbZsnPNbNd
QnF+tm3lJuqrlomz9J4STdBqDXlGQSCAnMP1kDhtyNUOKSq9PAzXt4O9lLIoKx1PwbTNMpxJnxtx
xaJqubQDypXAtap2ZTphZ/rtAwFGcz5Zmo6E8yKIb9TJetUyYQDnH+gituGTbJVli0a3Iu9V79Gk
qd781WhwS36XzhD2uc9zHWJc8Ce/0TDbBN7mYirHYN5eAQdORv9rbcOOTYNmnTcVqb/cxxMLC5En
SdFYf59aYvajgmqGVVijDkPSaqrQHc5XBLo7KX82J1aSV4QRPCfyRmMcXS3uoqi6UqZPH/sDeyvX
xI0rIJP/wzhWUvXN/0K+pYtbC6/LCTJ+H0z1YcIAp/GOvVo5ockbaSTkUnwoqa4Dk4fjQvbsM45Q
FXWamJAONppgN1tX8WvlOSrcmWCp6iNxRx4kw1hucQpowrJU4t5tkjk+C+vBM+L7tZXOoec4IlpP
kTrDahFfhPeGoJz/Iwdute+7pbmLoxO7z7tnWJrrQKwF6AuJdp3zdOtSBXA6+W0qEPcCoc9Vw4sM
dlnSoZtcPZ1hoF9fvESJqu0kTemHlesHUKZgQAGkTpouK2PU5RuI9VVRg0SR+2KghonX9vADNktA
BiXgPXDBkPC+u/uP1btMjR9LCi0a5X5oNW0GY6v2Y2fkLxJ9fVMignuV651nXH4aYzyrYJ/HeN1q
sSir3wYovnloicBnYQnsRr38EVhufzxk+mIzVGRLvLaP4ypGA2HIRFZIjEfTnBLxlMtYQKL6+YGh
n3dh3Jztwl0tltbraGBTPiJY9Gr8yqeN1e6ckdYq2I4XxjYktFNTon6WVsIistzQt5F7/LeUeNsc
sEe/qhBiunPQmTPDb462YhUV227YQ12osC14FPKGdVArXkQI8LU4Uo5iwcfB4k1CZJnEaqMGHpof
1vqWNgWsbysrK/J9m6FDLnwJfLEja2nVQJGBDU5gax/X8nYBEeQH03JRK7B8zG1Nv9ZZx+jgesge
fjvlByhR5w6DRngC5qOqadWYzRaGpC85ZTnQKIKB2S/BwgEqvEgzU3cvEb9f2Quc7YFkmvxE4HDI
7osGU/Lm1YaIc901vZ4oHdoly9HA/0IuZiS02eTtiFi1osy7k/7FQf3vnKV7orT0wfcL/D/gxMwt
lMYqPyE3vj7FpiOAJhkqKcYUVP0bfae37HFc5bYqYo2NFWLg2iX6yWqh50AuURGth7WTYi4Iz3o3
6nByk8WkczZIJGmLbVctVbChrs0drOiHak2RU55TB5usjkZgr3+V8uSBE2jjN2tGgXuLVQmSdnuC
WC+wQSvmcVJ5fmdQYOWaiqrcTy2IDJpqkvS2FJYVd/cSvJUwFiRRUZyP2YGXcH0y/G3td90dJwT+
gFnkAdQhUJ4RjpQBkebMRL1FOdPISDw3+frn5P+FQMXUYHXpSc61bTZ0nNrGGPCPJEUkdnoSiVuz
UHN+cBn2n9zobwYb8XrBVfpsEBRzVyd3bUxviqaKvlnFx+FFTvs9seqgZOkiRqbTv19zVIxM80Qy
l6eQ4H+CPoLUwJY7/Td59PHSj2aZyOKr2YH+iSJIdAYYlEojIYJy5OZPwPjdpR/Dwt6lT6Tyy5uc
SZp1O173Io/z0iZb4+yevBIAPQfnK3nAuo69AkOfxdF2ycwA15aSs9MFsyvNflZ24sz1z7JPe7LV
jpwguDBLWcUbOjS8p4AubZhD8b0o/pm78A8VX5PYZdfek8yUZ2vBphOKijG8qI8Sup7cn28HT9nV
EKitw6KJ95zMJ5kiW2RgfDV4zdj1I8oeQ6pdK/zczE+nwVjR8PnbOpNfSGlPzUC6npRt9EzXIu8D
xZXATzLmeRSFAIkiDgJJntvynMcAjf4vX1C3v13Px4oJdXvSZTtO8qtRQWwjpZ/2Wzm9UoAvrSst
GrUtnQINI631Zql+dvTQ/glZKFuqAuQxqU7DB1NYvFMEfIqGqTFRWySLZiDMPHKLRpsE+CkxwqwD
gdJrqVS/of4f6vsusUWeFioENGoMSsIyZh0j4E3VQZDdjsIIZNIasnknPiPnWx4KwFhxhNCBN8wX
Pe4lH5GbJmZSzRGzIh9fyXiDwYyTu0Yf/J3o9hN5vz8/+M4vbVBxn81i5o+MgUqj0tlK/F3pttTX
+Q1zvUdHfeO9ZBjH1JD2CAR5DRsOQbDrM60UISlSvVc2z9bTjvF3+cAAwqAy28ojJxrs507o4yky
gFS0oeBZ/RVLIed3xG8jFBwIAAXrbM7N+QS0w1IkPo/+vPpssvLuYHjVRPIqD+SPUY7EpC6Ea2Uy
qJpOy+siR4k7A/epSXRUwc3ehXW9+0KDDwbfvt79FH7r11XqrEnL+8hMAgeHdbsAc9+5aIwCR4tS
mu8NHhJwTu+PKqRzZrnuQViQAQT5K3GUX/Rv6qyWMjxXUIjgNxwgIaKOFCrHH0i+7Px73cKZJO+Q
98xrp0edjJRXvt3+w+pKWZFjW+cloMHQeUGxWmDFqpV0KbJy74JC1Vbr4TIeSTwfwFW58ylxn7G1
eYdZjp/qktpMJwo/WcPD9nLjtbWGy2wXDgEQUbAWgwdvehI90kF0MHCx0Qx2ldl5mu4eMvy6EiMz
LXYy0YhyGBuEedZFjuUjQcgPewRVXCWA1f8+N/pIhNK+B14VQpvuZLDiq/OetYLCCmH1nVHg8Ucl
AiMJPHEqeym3SCgI2GAAtiVr6eGbjwEXKm0MPIDhzXOJBR3R9XAl8bNSx1BnxGWzrsWc3kmRLEHz
9XR5M0UwUi3n0DjeL3ovU5ODYpgMU//PFhvS9D3R5ZdfOCPPtcWdeD+OGPHiEk9PfDlat2Fb1R6F
uXyxGPvojtSFX2tSlJcb/vedw4V/ckYOYzZqldCDsoLbI1MtnZ938fZS/pHqGLSOwDfvjYuxZxHa
mfB/GnE0lMBjsXdgNn0sWJd/H79UicjvUSbbvc0o9QOSaoH73UUALWd2MevYxG81XaSvARb0jg5p
ntb9PgJBVHEdHHmtuLRPjGuII8Vk8A17SImOa9sg4s++Ony7guJw+u5aSIUinC39Sbno9oY6AmMP
RLuU+bdHt6+b6QUGewvo2V+qeTGyZIy4iFmodkoYYv7klK8i123LIw7vcF+1ERdSbjNuascmh9/N
rX/vCG7Na/B5hi2IBb2qWxkeo7yu9+ptdRo2AYgblrm1dAkN0U1eUgo5e4a0VYIOkIQZFaq6SVdd
4kLmAdBEJ2mgKBL8FK2pt+h1iEchMytmkevkD+dL9UMRtpEfgyGky7Eck5wvFlFh2PE8Sna2pXFY
A7S/K3xwP7ybrh1Ko/OICXpEmE1CiB6Il4lmyp83xF6Dq/E7KfJ+oVGkmCyn1i5Wwcvq4HkyvHu2
fADmB+nv7xWahvo9Ngx98dQId5ujr4Nm3gDvCkcoULLLqUQ9RYdwUUrs08nwRuydSg81bUlJZafW
DYIPphdDMaESx1V5fDw6UXS4mb2KdJoEm0+9lIZWKY10f0DhnU0WWhB6DO8arp7Q4a5gn88bfyPw
4I+7rnku4os8bmfxSrNVF+JcOZjVkWtJveSPoh1bYrlmgu+3OQoYA2zKaecJf34ecPoE128c6yy3
4F/ELelZJvFPcgwDkYe4z1hvN6981mrYklbTkJlIVSerkcgWipfcShYM7zXf3uO1KPdnZ2LLoJ+y
kgbbevSrVfks4xvhqqJoIBFXS+9nGxqIO0FOEyu8Y9G2ioWvQzU15nURLtbOtUuGvNUctxYQYbDU
qEUTFEk02ViJen10hC5H6gUEl88Q+iJ/0PvCu9eE3LrAnpYjbGVwIcIH7XjFDZ7WWdBv0dSCle5s
FZG6XgVABr4z74WLS3KOt8fwgndhjf/gMTh1TlduUNKyHQGSeIgii1f981WU1r90Zm/EFnaRMStZ
WZj4RxN2a9oUZKYxz+CTU5TBFoK6m/rQMRyuYg54wtszBSbxzdnsObDctRpg2eielgOJpz568V2z
Hk6lxz2iJ8SWReYdcWPFzuAkgDnkQmdM+uECQwDD0RMIMO0M9j0B/y95x2rh8tA57hrv/YKme7sZ
X0rTqUeTZldQvOcH2NWQ1qqI1U6WYIKyE+5WRCuFKrgvs200yrla3LsKzlFZKkLQBhSLRYOOIMCH
nUqBRF46ThRyZ1O1lIbaiNoVIo2ro6QdqUKGhR73QIHa4i9SX6w4+d3Zpaql6rvcITl/a6dqB+uL
Crqoj8GzWgO0IWjuQoXH5hkYSmbawJv4voA95ouRjM6HMgpww6hwKQC6Y8FE6FMlcTHLbbeJ8Fh1
Qj0i01g073b8Ew2wdLqn7AnvP+WlvG9umTI1bv4kV6P8+t9d7lV6nuKcMYPGEbgD4kc15H5lVT7U
8itvqfwXOygnCAxpFniRDD/OCpIvwBa/y8COrzBZgFjj5SKzE/+peJiB9rJWV/fykQRLM6xYnaJK
5D/azUXrpUFgvLnXMrZMOE9ipBhgAvFufiQ+F/hQbl/pkGPD8SHi/dQp7mMFBm9AjXAIPG24WOvZ
+F9CorxW41L0HYZD5lSVe7Mw7LtnK5ROechvhDqPoSNeP4RcErO/3qvmfadeM/B5GBy8VecnJPlc
bhjuQ9xTUQDpHyGrXB614moxFlf6vW98a60CfxDrApwHKlWZEgHp+FHmNYzQir7rgu8IJRSxb7RT
QiKzhXCojHD6INr6a95ptE4IQ5DhiDhAvRs4o/2ToG6T1uuKkMiwQefQhokAepikUHyaHqbyqFEq
8d6oZipROZ7HIJtkUmhQgkrWa5SRTJDCFncGL02iuKjfh3+OM8pBtD/YvDTdYQkmrDY7GVlybge8
MyNLwOQVyASvkHLyG/yjiJ2eCI9sbyuR/r6OamAXeX0j3Yz3g0iwvj0wQcha9Jz7JNT7MehMhHWM
gI55eLfeLv62sr7akhauAs3AXipMF4FBOnk3kqxKnx8GLLPuOJORnsgQczy20cbtKmf4zyu/8PLR
KREA2v+g9r1Ixd3UX1P/COBmSqAiNKsIcundsIYH50NDiBAiVLnR2e92GTLMZBZQlf4yXFwTU1Rt
MQ68I63hPGV0EeWGgYODcbCIyi0rD79lfepU6t2tu7BRr5UyP1ynRhlhSJO/ynL0vjRFOJbBDUef
gpcfWxjEGCxYWgLnDDhzw14wZoTEi5yWZRO0eH6bhLcUq3U+mugFDA92z9JKO6cvBKc7DWlPnUm+
msepdojmSNO2VmQzx1lGGKRMDcV3+zxowjZAAlB9k2ljl3k0oA1YpThYygbQZ3Nrz0FJQpWF1cDu
rG45JT1eG7mBppQRbHKWCBUKumFKT1IWiBFbi/6m8hgxPA3Wf1M6Zb8WCOQzrwMHhYCZSZEjZt/u
zI+4Lp+ntaLBOzgF6bzfN1biCnnirp5PLErf7OITN+OHtlLG+HhdydKTGaf1cGYlOOv001NSMdty
RgOm4iUw8U5EQoUI6TollHkenH/fAphP63MExMdZFnTiMbhry6bJKUg5Q7Lw4OORF9y9e8+Rbxey
aaUTDA9Ktr4/QPO6IVu9USD/HlccqbcW6wBhkrAZm6nMmqpEC72m4A0xishexnpDMi0fsOBK+JxQ
uTp97DLyqLWEz4kL2GqaWD3IUCCWZTgfnga2vI0jo8o0YreaZq6FgnHADKe7bazoAZpx2qWy1Oa1
CCdKjDw776CcoEo3fHjPYdD7BLl/opxghkKhb5gHgFCcax50b7M0rUv28DgXg6FyyCLVQ0CaCJS4
nWoXk3/gCMzJ1dggufDO4alQXyGeajiITtSPhHXBYhDYlGamAqUZtu7kUwB747cDf8CCIeoDCDbg
KOFLurBhnMy3f3CMvYLMlKcbwS7E4TxQVVjfmbZ/BY/fFd/Ol8aOYDFvkcrHNEu1pdEpKp8Vx59m
WKio2nfeVJ0vHMaiXft5zs12e+L4LJDTEpN0SsWUtI5AhKEWkhQzY1cicxRVVrylw0OyTn4Y2S41
lOjg4JwZkVPli+lW9jQieEYfrWFTsMhskOJkkgJEcTj9h/4/T8DPgk/AH3o0zcr6mT7EiCGv/MJ0
trx/ZlDgWJXQd9UzoZ8VyBw/3Q4yL7WglIE6VeSOU3qTgvDnyLDCUoerGx0+UjmSt3tNLFHIAwxe
mMudDCa3GK9Ae4jd15X5AirWV2dTxkTV9DGOmN2Q7Oazv940Un+025tlxgPl+MO/CshF2SpP/pCp
o//8+cQ7cUmKvD9FcRr7BDcWpzpfIxHxDbbL4G9PTs+TusNXKO1Jaw6vB2y+aXUw6wkpaL92poqd
eP8FE8J7RCTbgsxs5iUK/Y8IlYTSVjA2O91C9AaJ4CAeDUX5t+gxUERkQXMp3PnzcUEu36TE7jUV
gM3mwyX1g+C77pdozH0eCUnVBZyxRv7yPxerjcVpJ6dV76u6/V+4G6zqvASPXrWEx7IELiiSYUWG
XfVz2pKCGiSSvHkYm7cLbQvHsHaBmT3/bST4NCHulHfMFJtohgnRnX/Lk2T0JrQikaLGCBLu8o1f
O0B53yXHXfHik+R/4ERpYE9+7PWNZ75BvruafPR2MFsvHOGupwLQxbs3gC44Sddv0AOfjw6+zKiV
KFop7s6TdpANJi48TxrwwemBa00tYL9AClUHUWOBTJQ+tQWy3k0r4rgQtYcgzco4+AAHJ57Rk8if
yuuDmB9sOJ5QXHXDxOf+aHR3LgtKzerxTybuPDLmm+YfmfsDuOjKNCBn9huGW0Yb1keU0Kt/Ygy+
DnA+vA2NphQxfIlWPBqrUlJnw1qioPzq4YRf930gD3A4sO0ZKz/7M3tKbr3JbPDeQ5tKjWiKxZqk
oHr6822qzvzRXGxFdsTvTuSalC5DkBtNIYNdG2/2hTHWGM3kKFhwmac+RcHk7E1wydO7oZHkBNxo
aZmmSWustOKZkuWG4oSJ8Bi3ig17r5UFRN/yHC595eR9UNwbTsvRQnBTHUfqLhURV/4oik/Jj/CM
7+fVxsUCiuesmI+eHk5ENepgtjB6hygv/tlkwNka5dDzEL5GBEkFTaGzVhgQ0LhgU34tgjleGtcJ
Ms7orwqEv6UfTnp79e9rALmfMCI0MIlmgOcX/FhMJ9pJHWmlD/4Tb96z35jU5clb9Cm0TTsdKs4j
CZFp8+cSNHKPSIoUFz7Cq/ppIlbhjU7pAnmhyKOm4R4uT0+DJLkKyCQJuVhPwQjBkJY3QlzWrgik
60cE9mEV6A1gAwca860wX1B179s+gqXHnLMP0JaQ1mT2AMfRhniOcK2f2b4dH9Lh6HW+D2E3uGZI
oEsB8NBC3MRPEv7hS7eyVcCYEUZK0enViKCOzfwwXdegjWSKK+R/aZfcYjXECMJiMrGic36PwNyM
ZKir6r7R64pdGKpKjHiE9n3D9fj4TdDHBKcu8GU03c81gwDbFj1NqJKyJ45Q4ibtQ6ct14HJy38r
Uv3z4IuiW5V0HkQ602gMq566FE3wrEIGw5jBQS8Z6l4+jqKbC56K7sXBxKD2rs6x+pSniH/uNgRf
+yk6PrztpPm7umIpIkLa6/Qw2VeQTko0msCUUAqFf29Rix+DpcGIQmjHUSpQIgjrpmIvplgnyAAf
2FuUjnIUZZgs0/GM9FBUMNk8OyTNUaqfxqXAow+q77Kk7JZLtbG2Gd6vF/Udk82psq/umDVYRBI5
JIgC4J0faM66LuEcyvo5enFfYqxItzTNmm/48UnKSMFMAMPKIWBVAtZLBhJ1aB3DY5pU4JO9drWO
muKl0M7Yk7fFcJfFlwMJfSynRaU2OfzY2JLfWQQ1cukf6XiAM74vWpP5HCUURhopyjbfvbkE/sqU
IqvzNQDHiVIhbKtVDtQRIiYdZiBjQp0SeSttr3IXQtQarPKVhjMPFttobCx+s0RgDwEyHKsg+dxV
a/eZZuvrUKlebPKApFlpcWoHQ9cGgLLEj2F256LnKLy0Fbejud2DiSS4G41MJYvVdXYSLVQY0uy4
2iuhqOkurWAQNQCyH5ac4DB1SZuAc+Ot1R6yPlqwHhUxab6IAkPZGrNAL95qSJfeNcG6S7q6afP+
qngTboVEwoMwxgIjFuhAMxYcnNpk9h8/FeSIA3b4NQFxfP7Yar4TaB86bspGchqhpabYQvCc7Tmq
35gsH5PhQHYEU6DmSGxlIUDLo+EF2KjZpe76jQeV/aNzV3+3v0neSp6CoOaXYix9IEJCzr3z2aZ9
56xzq6ZNY6rfws42G9oJHGjcAAyzI+yNHk064aOq+m74c5jR4OCiBri7laEftnbOnwXNoVjAJAdC
K+VUe60g3hWOme4Ap6BIIBWIjlikUmi0zBL97Rp7rlAzP8aJclp1Tq5BteUs9W+MvbSPpUB1s/pf
RBp9aVgLLmIH+WZEp/5CZg+1ZXLY4VT31NYR4Ku+n/waTEWVj/VnnmZFmyzUjAkLbLHFCPCAS93U
z+O1kgkveF7s6/+yfv4uRzNpp62TG4AaJ+jQ2aQP0TCplVs/35MyMSx8fasJeZsZbC+x2pURqYzv
rmEc+SbebykWOXVEx5n2TiuHDpTzv6wP1zacDJ2LzBqCzVCkXWpBCdN6bJsY/IWIuTtYkbl9J1Y+
hnhVRfyUlsipLVjpHSpcsV4XKATrds6Teu30MuxeLAJKGvMpkgBxKw/SyRpjLhzNn2QkpcKmklXQ
6ah7esnztyoWjbCVs5VlnHWoh/QjY0zd+SMcwN2fxwyE+Q02QxSKD3P/aTWUU32SxZ7iCtSpRf2U
TBNuynJmmNw7q9Zr35KAw92vNRjZLZCUziH1gWWkEl6ZHxNkY3EpW7L425ncuVONtkPIToVhkc5z
RhelcMbRW+mZgX5BbNk+P90+RUo2dJL7fZW6X8aMcmrwgyx+3/0+7g8C6MQ+uOefnbcNtWFoXKWs
/kOMADuNrLdf/9W5BwdENPBMVRaA6b5vlfU66SMGgEVTA6b6eaxkwHLMiCOHtc45XLPV1lO7e4/p
qhTqYCLpNgkJaVFZyO+1+t34W62qNzAYvIje4sVwEhMSJwcrlMRQ/phsbhR6Vevtq+hQlB+OjCwu
ZtpyVjCkuuRsAdmOmM0UESw3uAJYR3RTpmRWysaCaWBgQNl5QBOrhW6YwBsApaGXCRyNrW/xQLp5
cpbO6LmNvYQd4mtZxg1avdsgXLG+QQGXH7ptHZhdbBYORZG9Xz3/QNX0/9Z9ExcX3edc7UaZBpoX
x6nyBfdgXe9VbPTu1SGXqdc5WZ/Mk9WVcOrKqdsuDMj3vx9lea+Cq18lDBiigF/iOPKh+a47/LQv
CQWGcZuCh/IAq9jvk3z0z+q++/xn/v5R2bETfrsfIAlUTuH5/+qcQiueokp6I8MLBESkP7Igrcjn
ig0Ap/MX2iHieo1EBFOQ9otTcbrQC9+GhLRN61caORpedPHd76BpXUNp1NYT9tWoX/W7KLVmPioG
d+liIKYz7KTlPI+7sif17nZk9T9ePprBbSYh56xVBcbWRG2eAs/4jDqB9IGwECNs7fj/+nt9eeq6
txBhtGnyqc8vYCU4sHdDCdW/qNQIMsovBLGNGsI+9dXShpYfHyDioybDD83D4c2SIIRypxmt8VPA
AHzh8K4Ib05TLseNUEDKz9VWvfQArh3uAmtAu5yVKTBnmAsep5W0MJ7opQzq1absYkzrHnA4Z7XD
TONNlZ35E9nJpMzfrHZcy7joaoCNvU7C/UAkIfLrUEncWNYjwLVe05pm/rHtd4p4eGm4LaRlN648
XL0CkuTYa/+9IbnG1vr4DiXjw8rYD4X4iWUhROV9PFFiTYjXGPNaNCO+G/txb++mHdgfLgzWv22T
5izn5ufSj3JPGgi0gTQgAyVRADLSXW2AoOzxzfAecBKeq+Ip0ZgKREQRn7zRskWXznTqzi6x593B
PARvPHDhKVLYDtiSNWUvy6n3rRQiAl+lvdWJjDOJvYOHC/sVgLJslptwAnYHAa6swnrHilTLT4Yj
oBFD8eXvs0XRvewZQ/68yjzrBSTnde5b6Qem9O8nLYTIfsVNF18RqnenwiFUAa22mOq6WT8YF/oH
ydbUkGhCzEc/FjxcSHk4iKAQjd9ppQBhVLfXD3A85hWCHojiK61Nbt0p0nB2Y8AUKbt19VBekKXq
O3FeAn8umNPiGuSa6jZjBq1a/jl2MxQ5/MR00CDBuSceEC2lsRQPGiwfCYxogmQJ6jkDxUlYKhaH
o/07G97cFbheowKmiZ28X01SzUaOXMZVzJEdT/JT43S4giXoiX5GbvmlrJ07N8uMOhkkaqOyCCgm
SqyUwm/+wt0LC5FLeGxnvKBG99IxG1+EXRr7NW192utv/gQ2DbS0bkQAfvF8Y8yt9bi7K8leSfEe
c1/6FPO6fnUUZ9+12iLlS9JtP54Y51Q7wcYxArWu7zcUswWz+0CuvCz1WhO+EwZjPmQe/nwNF1dc
yyOm4OGczGmBSBB+7A9siK3BTpViZyBZgWmtsJ/fK8eX/ooRFNVNpwIXyAIOlApl69b+7QkpZ0im
XpqHuwFAqzodk+vhj3E/5y99hJOuGaDGjl3mPthDEWM7xJ95dWL4nDqXRRpo/Ly4WKwcsZMFMW+p
vfLUbFE5xSp55kQGRfJF2M+9CB2j3CUvzInxQHQJ5fMk1AiM/T6VcpNBTCtS2tuSc2wlJVTCtABW
MBBv8P0zjGJ3rnp31/JqazDtrAQhpBkVujlACG4ezdyKV7+b/nqMai3yO5HECM7kbN6AHG8bpxUE
J1Pnl/d7rvcNT5cxAx9+YX4jcn2gAy3WHNrkQUQKjMHlRQ/KBCijFInUUhTyhQM5XKYcOaxaTnSz
+78qWzKbp/XiR5DKKJthfm4CmpBnuRM8XpC7FDn3Yiu2G9GRXpGQJbmXGSr4LYWUIevj/iBCiHym
HQecRQq67jgh8aH066h4d5VHYYyf5yfvtecN8DkJWuUMF3iefahWdjnZLXUBPqW+WSAx546kmS2j
5zUeiVOse5/PRGIscpl72lMYgHWRcTZwlFpmt4K/W2itv9b1OkBQ2p6f9BuuGzuhs9j1+2VPiSWY
D0l+6SIhfNsJ0RqAGSJ64DnnUKP7NcVooSyD8RV6AXjmAfsYBVTx8YN+W3pwndntt2/KJG5KDmG6
8W0cFOttwLzA3Z1H7vTKbWRs2Z2B5h3hk87DkIBjlr/qm3ommIfshZ8/VXfMDI1kTuxWx3qEMVP2
5s6DPAykUqTpk+D56zqfynNODY/ru6L33vLKrGqm7kHRVUaSt6mZg+/H9TAhS+JT157TjP2mTJBT
ZBEaedYMeL4hPy83QkrRbl5H2K2f0zebBA4rB6P6lo5h5+EZS/9SiBBcZqAvui5UPlohj4r+ocZe
ji31K7Gn9wPtAFz0RwX+eXjzsY9PL+v0Fsu69FmXS2vpohsChD6pzBvDgDlfPF1B9ns/FxXn/UJb
PnX+Fb05Rnz30hfxZtDLZy8n/lFUxkqV+NYCOMKA1oaTo2rgWtH6ScBWdDQ9vtOU/nxTCAJ4siAV
P8xniC43XU2DTCdX2gxzPPJ6CW2K5VmzNMsiGVDh7MGHLEtAJoibGWtqnpGXhtjuC3ln2bUwKROg
/dqpGTDRmjA8NSGlwo4KvIl7WKqaMtqmmRgy9oN6+fGI+GAd59cH0l8hlr3ey4/lGjdT53V0Km75
3jRlIgkfvf8BqeAQ+TIHErYdLKRYxfDvl+6vw6F8ANbj8LpzozTwu0amWHRgGmKVElOZOH569PkH
cchphNJokkl7UwtgnItUv12bF20Tsd+y/TPod1m/shyeSU/97ig4MQ5QANklBc6IA2TMV4nNFwrq
mdR362iF0esVcM+TYIF8ej41bPoGb+gBHqx5MhHwiAZai4hi8qi4eFiqG/DpIUhUBFCM8Wwyb6TS
IIlpU/1BVNliTjK4TbtFpTIE5WiqNphBPhm132Rx3anZnAvX1bjLAjfnCyRBqJ5k9OVeosw5f8Pj
g1r0HhgZrH71kjwfOqmDfJoP380lJQquGikHg86eAmk0iuM4ieEp48ArMKx/FfdM6wn+2Mw1vWfa
67TypbH5QO8NM0mR6eD/+5z1bc1krqI89J2XfsffidYlv4FZpc/sMEudV6Nhd1N/0QK9OLdKR8xv
sciEDrn8U3f/ikMMlGR5XOmmiS6KZA+aeyOCseNw337YV2TTNHOfesz03UGU49XpFjGMvsO3MK3t
yq+ibOtRVKZVZ2boUX8VxuUtvV/9tWO3nZihQuQvzeL2UeW2l8flPljRp1ER6Ct0UdQtkov3Awb/
3zh0Cq+gcVe2biq2Um/Ft0DYlVJ3V5l2udbXdmJFBAaLYfa/BaBwWI6+iG/fap4zXpSJtdoFDGGL
YWx07O6gWjJZkD+g9gZrKWiozwf6gHgMHegEaNJLKcf+FdDOqUN2QgH3ti8Y2//GD5zrPJzVnmOU
EvybaxFpfkYuP777rkt2NdCwqZLwLdNUKiwBhUGJqknN/iiBPEWkjCqc8tftZ5849J6pKQBePpHE
/v5iG3NQhRpBwm3MvtmOlljCp/WrrdIj/YttlewDKW1xs22NmlfoH9iwJkSlUb8s0afgd6wzYidy
2K5nLGfBsgZsmLOhQst+p2ZfCSsJyN6l0WX8yTZH8UMCf4qHb+5Xz7vTX8OF20Km+eZuP3gvgZLU
FQD8cFNMQd8YEsqhYbUUtPlbSUuphcp3sCrM00Tud76iCdfI2pFkRSPiUVD3VtlHFtynI0ZhpdJj
AYOOJsT4tVUTxi/hEeEKEZz19RqnnwHAKvpaEWmFa8qw3iA/hcZOOc5x3hG85k3sZEhm2wl+X1LZ
yMWDACtTy3hiuVqAKd4A7NfQOmrNYq9IicnohF//lQQ2VXwyJWptcLYqXwrPTj5hK9Aj8X+1EXbY
tXmZyHAEU57JSHDJ9vEczX3krukY2dYnKpwzyMima3PQCUEg43UNXULhHcQbI95gJNbKTAGMu+YZ
CEG59WDJkdTm26j0lbGywl3EbHhF4P+L97L4njPMYXfDosyM3MHJkVWUVC8QSww+1trgq1ig71ni
3FDukdrmDcjMUnxppPLIkCJzpX/o7LSn7NJzkEF+usXz/jI8MuePfoZbW0L4aKeX/hqfJMeD31ow
yldHsyLly1gTXbEx3/z6QFacVJ9Pnt3YQka7ViIBpFx5pzWJjoqpXGF7upSGH2G+N5NM7OQAvRv+
7qFN//5KVFpHeyHc8J5aZT12vCdSTbD2eAy/mZNMxTk0xIbZlxU/JJLIx2JE2kKij2mmoNExRhM4
1Z8hZK7m1tt5fYcMmzl5pUUyIQ5iy3OSpZYloMVsQyeFdqInvXMXNvymhrV9bzuze1420IxKm2ol
ISfOErN3F6CWzcTMUlxrCBYOk/Zod+6H4CZbRTNi4SXNLYHeNAaiv7XsKJwdAjVFwsJjef4sAuyg
sgwVtODhl9QVC9S7fLMD+Gy00Z4Rm8lc+SCVRLi1fZ1RHuaoo6owCO4Bjenj5iNDvC3CwWtENAYt
qLMh8H6H+lmxlxujnunxrTLYK+Hg/8WGL2A8Y5PyhSuB47AR+DCT+qfTD1UO8iN0JcSy53J8bt60
Km7DNR7FDthLNlSLp17HWZNp82dNMFjQx4m4FT46eccA/lXKuWMEu1Q1uhCwh8V2r9Dm4Eu8jaBf
l9bq/9VflRB9wdasHEVDjEOsJn4rJzWFMI8bCuCexbwJDlBF1Hc4NNJdkLM0ZfCcposxYoRQyuu+
PK4Siuu+tTbqicp6uTCb0d3gqwuUsrF6JnEo3idMjNUkhEfuV6+Eh8QNBgpvydajSQXCSd0/ws5U
DqiPFIC493qCvUrXGmkxjtgWD7a/FnxYnLsMc/rTgouW8CrRTpX6JkKdWDPinMrbsSRllTvHxMyZ
fUOVWYd6Q1mpaZRJBibpbunEicWJy7ZJPDsmORxY9ZUcdt36wF7B21rhGzBHTRzrx2y5kwjgEKgx
yfJWl8iLd6Xl4x3g49hxCs1hvouiC/B26INnSpsaG9nz3PhJ7r5Ype8QIKT2+mMFjzUAKRgFK+KM
tOsna8ovDyTXaSvsY56QWkcyH6gaw/e/Cw7995C8YjXnWhdJZIsU4+ktEvvYdKscuZ+3lW9TACcs
wEsS2w8lNeXUHTQ8Zlm4gzFmOiXWbQ4zOgGbLK8vKx3pGvE3bYz7bJfPLB6ElR+sZUz6q99dgHyN
OJ80MIaSXcq6HktXSz1LewqyIqIzoWwzMet2ENdI2wPzjf+EcFFLwfoub9Z3Uk8ACqUx8BFKn8Vv
o7BTDzTzgZq4AIg1TiboDyecFwVHxKLFz+r6qc1ON1XiJVCSpqWIafbfGinb61+JrQU/oXEf8O9g
+SSvjjwZleDQF3iacfTilIsFdh/au4K87t4goWFJ0SXF8DVjD46WImmmp/+1TJ60zCUmD2GQ2ZhD
pgxKukweacbSaB6GW8SdLp/CTrYPNYCiLDfgFG4cpFGIHCMIA0UMBvchGA3HoMcTrOfTFSvm1BaR
fD3/EZxWmze6oCXAdWUfp680GJVae5icQsC/yMKlslTxgW8rJvvMGUAASsw52HrNm/b15sqonTbY
+povCZ5e0wAMhJeaVkHuK3nvAdW8Sg7YMjc/FfBt318HAiafcqqiP9A0UIrTNwzOPWk7s2Y3CRMF
PQ4g0JDiIS2QOkY2rW9Exl8oHeG9EHVoP9j31aJrprUtVMJLj47s4ciQmKAYDNuexNdcZUMeU21e
D1mkAesoRBX6513a7TD2cQVJRbqcfAjnnvf9L96dikhF1EPIEW18RaA2T9DMqRct+Z/tFalctCTA
3XFedrf4KOUwAx5sS7yEHyv4eAdv89wW81AP3DUI72SwKoSMy7CYj9MsHGlBiS4/be/WpHI2O3vP
enXvTvf0+KnjRymlHBusMz8f5GKIJGg+l0TGe997iefnDMEZEAO/TGmzaCv308ODUHg1q1Ee4qcE
4/1wBXTieT+ylXX7fgNiM2NhknR9KWmSjhKvVXyeFrmcfFmJLawabAcSs18S5VgybPWJBXQPuMGM
veGfnfDUfWqjvJixPxP+AmVUSqSH91H4SVs9izGaDbS+JGORlMCS8vMHs626Qzr5IoA+5X8D8hKi
qJpCaBP+wVOTwQNGk38kUDwbHRJQXi+UKLf2794mHjSm1DJ2O80HY7dTj56FCSpx6sDcerOQIKi/
6tsw7Z43qGc/rxplaO5QI6LeoSmjFnKlYkE61PLoXVhixaOKgpQlUuJw/McccNirinbTEH/syv1p
2Jifcw4d3diBlTdrzLaNts1Z1A+iVP8fwX/DGd4j5jeVi+tE8iJJ7Khg42Ipp8NzFJlzxeTjVw6Q
SzwiuxLtBGEj2l40dgT8tGtj4ytZLjqgnsuARH7V6P6g1+frxxhzx/rJNTQOA5N98MAJTpp1S7n5
uRS/fHxhdYX8d+S8D4hariBH2bs/q7OropfrJ7yc7H3XMx4fjZUUBIItnc+i0Ke6GpmuS0kOUgPi
s+/N4I+FIMUp+yq6EGDB45qZcL9zNuOHDp5Pnw+yEXkr7zacrz/6PLq80SSIzk0kczj+GC17y+6G
6k7QuI/pRdcg/oLBwdXYbWei8E1TljjTo4SBdjCUAcoViD0pMaNAPLcUKXmC6JtahNpzWShEn33T
kWGyUu1CN58LfKqeSaftbXlwtbrTFVEzWy0ZkPVRVY6mY51ydg6zltvOsugBSvWrywj9G6L6RfP4
g98vdeo79dAAtaD1215en0W2DK8Id8Q+8RlI+FSLzjlEmHXJpRGUYPAGfypSTZvsm92cDiRNr/9s
MyS0oANHt9czGXUg8yvx3jv1YvnRb5vwid/tJsY6XqI3Thb+fBTNsm1QyD7iTd4QEPRmXrt+BvtG
KDYEFeKiE7Nbnqxt/Y2aJKcxNm2mo3h6jF5xJR1A8UFNAxD6orcVOYmerrNL3DOLAl0fQ/LW20/8
2crFdaYuxnLHqNpNCF0hrDYDPoN0Koe2g/KLOQNqHJIm9YDK7HjDQQlmDKAkovPoaxPJwtNt1WbL
d39Ief4Gk1EPkAJpMe1LyxXgj0mprR0TOmSWjo/zJKnG1eEeNHrPTstyDebhVIqAd6t6kRwvn374
dF9Ax2Hc5bmH/AiaNSyRCOSFKrlGzLXMwkghXDXTQD0TQVqbVzD1S/wjRk5on7dyWJDT52WcX6OY
M/C6gFdNEDsYxWldG5gGVm/dpiW2dweSPo/UssGv1mppU/iufqfKUV7C60ufRC2oZxop7fnnYYbk
49eTp9HHkkLB6FH/rcmzsIx6kFejmucDYSpj5WSEL8/wv4NW5PacGLiJJ3XtXon2MJqw9qvnnHqM
PsYtXloOAYt7wXu02STKLh/npj2MK+zUEfZYT95TSq3eq60v2q2Q95scgw1xQVVSiPRKWBUQ/Lal
e00450RStC6WmbIFfZmuo/MGZ2owQe8JfZv3irrJHR8BnSDX5hTwTOMrcVnGsDis517a8cF1Unz9
MEssWwf23A9L1qZ61thqrsB2iWrS4+oDXISXYdFPU+S+DQoYFm3vdqXOIcnQlmWJE7OBid1bTsV1
tYbY0GUuDoEdxe8F3qF1czV2Xgu6h7TcZvzfSLFAakRTqiwA0AAN+PK7WipX4HJ4ID+mc1lup/Hj
CJ2hASKrSe9HB5ZBfi/GQQXSg+obQsFVrMhpEvb0dYL7BtCu4v2zB1uVLEdo5BOtStRr2CxobIOy
y6JY5BM3puwosf2m1BUewUvtxAJbcySPsFHOMRDjBOjDG59rWLp+YUXU3GsXeE5SWKkRwHzAhx8g
OMCicID8/zzlIZoX3xX4f08+od58fcph2QH1h4ag9Vf+B74YxNTCT0w+zEalNmIj8KOyiESlTctH
2DnLu5eiwvn0RdF9WAJL1IwpfSUYqK1iwHKsWaF8oFv4M02Ha+k/Ezqpf5jLrVOmwjvyswRdDvbt
u3TWTlV4FEcuMFy+nor1JADFzlunRmCVvPSfnKupxN6MyEJLedYMkSRCov7vSWNTkQg7r9bvz+3e
Fg3+e18XuhrDQQ4oIOGfBnwdxsc8eGyTd9HACqR4bRg5B309tuR0iXsLks6tDhq8qjqtk4hylWCg
QJVIypLSx1QwLYG6U6weIEbZwUSPrr3QJBGhq+z4JqetuWyTGnwB7QMtw7HqWxDlHo8Mr/DID6Ks
qycPJbs4V+MXZew4XWo4J+4aeHkp5PeTRfmd+c29j7rEYslya7T1hrrzMdOUNN22PsSGr0aZwH6h
HmyXNhFGZItBqDJP3jYiX5oI97VTy/q26VLMOGakCrHJvjXTOHnbHjnEJpdxOFgjKaB9FhLc2Kx6
iO3FRzI8xFimRDws9+Qt6oX4Iws9yZAWQPOFCn0AH2SH+BjsaODKfcFqGNpi8R9r6oJYUoWyahq5
0CJBPz7dELwbdxTUEohGY6APJzOvUeDnMa0Tk6A0CLvO9Jd2xgNE0WufJ/XJ2H+xjheqg76gf4pk
/ZRIUtReajxdUp27KIOjJegyP5qPlan3rgVQrIrk76J6tPyJV1BGmhVkesZfxS/JJ8CKdQzQD8en
I9CMD6dSjr2SM+CwnifBfbb8IWsc9omJPkQhkdoMF6l7+XyCZamJHS6mz2r06LZ0fbDF/BNqk64O
65jyayA8diiXWxS9zAmNX1CMvpYWCeSG8X9U/CI3+ub/zpzr7+XHy/yTPKVTKGVWAbKekEUJIwiY
BpdCG4GPuV26W5+4DXToUEfF52mcd/57gJFt2ZQu8rqwyukuenJBoH6wHW/CSHHQGICOIpDKhLhp
zs4BH6yVaH5GqRlFbg9djOUAo+E/OEffr03mTJ91Bi50wqGMtfL90a85YsQnmvrosQUJDvGogCHC
ncBa+jMPR5qf+rrkqDipS3nc0n+qRvgsvrpKh59sA5/A89ZJkhk5YBx//Bdfsvsm73eoKXdsPlB1
qHWx82lqPGu2Ltm6L4xnGdn2sz5OmULv5yqzuJpLGW9P5netv90AWIJSrj7bm3W3hwxFgYjSwIGX
9JTZkmgdLa0wvRmik8yeS83j2wLS495UrSCMnkxjfhY66w0YsGMzwKAnvF4jzXdrK+aAfCtYR1ze
YUx0sif4PedZIxw5nzljJmOBacAKO76KjY9lJL2rwd+QPwv5cQtkqGLzqeLFwU7gHi6sNlUdJZkN
d2SE26OTpDU/eIUG3v4Qh5VynnRbibxht5Y9s+vVTyhn72Y4Y2GcLT8b600XymGuu+pyRqg4rc9h
P88/DJdHA7yAwA3CDPfgcczAqoMX5fIZlgXZ6B4enwkJTa4aIa31jKMUTFeCrLHXlFsZDllI2mlS
diP3mSf4EQVKRBNVipm4iXztyqZHfuCDM9VnNKQSPQVZWXEWvX5QYtMeRreaRToT9xUl0YmVWU3U
OevVgnPZpQ1EHJycL4OfP8Zxkna4hsElNLUZ1J9WUMOVoyHrspAjMUQXVMO+lQB3O8d/t9fAKlgb
mLkODb1eE5sWesKwype+ns90qh/kn+6PKagxLggkbAWmKE2p2VEXkLOtxD+/2gtf/gadCqCFp/KO
w3EqW9ODYtaaWkd5aUgb+00gWvOCmEuduLb45HGR/KF5x1RRNCH6B0VNq1PBXpkoekBc8kfxGwtj
NERZulwyBBaogkD9VjokR8AD6Gc+gpt5drMQQCH1dFBqjNVmaLa2QGFDhIMqnkcgsXZrg91NmQNX
cuCYujJ7cd4N8rLgMgzCIeYqTS2W20WueUTWp6zw/QQC+aaX2PgbjYyKa9d5V1bygj4kiJ7Rhym3
S9f2LKNRJO18A+7i5J0wCWcX39F6XFNNMZqJNw5Swuryseq10Rdx1EqG0f2MBLIRLBtRik7DlntD
Q/wXza5t1CMNNnjyWRfuG8zgDFh8ggwb1zj9vdNSt3gRQJuaxXP4YnxIoE8hcIuElHfXe8euz3DU
22PGN5uNkRHJhyfIAsNQ3BjCL8uEJnWoVyYYifauTDeQlXmSh9qn4OFlzrDyNbDW0Jvd2xFuzY5O
1qnrya28qErwfp+7vm66m5LT86UQq08ZPNeklU5//hV21oXW29WSH0tmr7ZrycAdBRi+ePSbD8nO
VkhPI/bUB9aew5ZXiqayV5dQxVdzhWWpTOz8wTDsO8hrFBQM49WrSUbLo8b3ueWmygvkMiy4urlu
ol80JSFs7HXYfvBfkyAF7O4quZa3SZnm64Yk8bjKjgfVtVm7s1qH1bEuhxGh6TkJnfal6VjDPRTo
Y6Yxl+HZ2qKHqofLYOSN3EWaB3NN71MhLgNH1qO499QmGAVM8BOSboGW+1ucnDk8JbM47T8mwchS
5MeCq//XDiCG2/H3T0/Di+njRP6JL1pgnLkojhQuM3O/35Go2NvKx1ykFsqwWKmoXQySJhHd333k
/lASMPUgjkL5XMZHeEjBVUCzaStodEIa32MW7KGeEqmtmj0rNAG0QzY4FoiPC+gcxS6qJLBTvuo0
n78MwtGBsb7QIbdTSLVpmTHcKNECKZ0aaBCrm6iVulqxwmevW0bljLs2RqMp81K/fvpLOeKQ50t7
h1ez/ZH52ShG0z5Rjxpy72QnqQbic+k4+lZ5WTmvgGtEWpN7ixjJf6qt6k3eaiAe1er0sZtIK+x8
eBHBtccVt84kw8UAmLvh9NXPTwk9lwEFcpQ3EFL9X8UV8lTHUehmdn41uJnC4TYddBj11AXNS4pR
WbWPM1gSyYaEVhxzW8YS1QgUkelQiS0xDL0ZsMWbFMFFhNqUccEEaFtgXKh4jAXQQgMrlXhS1Q0m
Xvw/Mb9jm6CkHQ0QKzHwBS9FKLkidIhb08kvt0fr6DhUESeHP/ZcvA2XnXcFC0FoaWswCWtS1YPd
TKT+O46Ush60K+tw1ukia2EqbhX9PI65yDqIe4twrrZ6P0CH8iGhu5fL7ZUvNCjyanaGiyba7eib
PEk3/BtKsMjRqb6YFOIQX+lvtJ0EWUzIZPAZaQekl/c5SYf5LkK9e9smnbdIlgdwMLbn4nAow61D
hS+2eaxR8SHEc74s/Vi/K1JJZEpmf/ktfrAR8pRH8de7CWJBdYqG/q0cOLXluAvnUkyY8wOv0R1p
bHINs+AjhAbipDPlgfUBAOFl0APfYfUBwN1s8WQ0C7qZ+N0Y/Nd6KYcv3CpAT/HgYvyKHNkC3q/h
CnSWsp6GHFDMLzWEpk9zHZLL3BbWDg+pCsDpS5gPL5KcSIzPHZ5qP4xssVyE8wymW9zxf45eSxxJ
usU/qrNuTEfsMPxEMWdppPI6cLjCHM71COeebeYVmdsqG/jLM2ubucHCqpbNYpz0uPY42dQruP77
triAQvqpqwblNYltPVPLJ/jLxIIlg6VuczLae6xkTQM5eCqqrco7OJKmsUSzGuBER5F53rL1JokM
T+216lgzqjg4bVhBGqpCFj8tuYw0Qz6Wjsf3N1rco8H4c5jg7NoCJ3BFqYmiOrVVk3XVHyREriSq
RuJ4Jrml439/CRjpepYdgMzxLxGZOKLAozKzvfYKTRsyFwTnAMFiKiBRdz2AYp4vRqwll+h3YRR7
Ipq/OzQckxcIm7oxnQQi7+0N6/W19JOjLj9YphQLXL6qakv9QzhGUEP2yEA1BmdsUuSG2GaXbmjg
nhykeYZi3Z+t0xFVBji9cpbChSYjgeiJiy8NKK62UgYqFwpmaIDpzlAKihpaBiGJtj7IFedlomMf
nspO8g1+Rx2Gl6eQpnDOnKJ0JjyPP0xX8RXCK2FXDqC9MGYx36mZoRhTUG9yaBjETxipHmzst4PJ
prJuhNSP1MWDpXq7api0KA5YDdw9yN8HDYiQTUPGyjiVCX33abWcZW1el4TmU3ynWvZ9ipOeaUMF
SiCe0l98RKQ6CraO0gTxXToPEElI1PzQ8lgUPU/ULHqqMo0kG8mKEeIbIvqiX2omdmtVEF+LTRiL
rK8I4xHlceVM8Qf3Mj5T2+4RfFELQ83PVQkcZR53HeD9kPkX6jnmnEUT7D4/ImY+I4ySiH6eHu3Z
Pkib+lhaMCFADV+ej4/wvzIZIqbbayTMtVwrZ3U3O6RNwyNYcGSTLnSCnVSvmrNnjPcuREM4yqwN
KljhVGTx/ESi1LfG0AmopD7MCXVBAU1JCpOlbgi6DiaFBdfZvEx8nxvP02DMi6BwnTzJUI6JZhcQ
2Zk8sl4t9A3FGDcTTIop9/KsOTEYE+pGz5lDEKDLbw+FKn4te0Ru9YYzJh65IBH8TZaiLKJO+gT+
D0ADw43fCjsPMO6RQolPSeOa9Xl8qgAr+pVwux11UPnIA+Wy0iFZJh0+akL2Z+bAk0F9vjumupLr
P/IfWbeDXkQn3sRLl+b6iGOkLSzPdQumY2QioyvyT1DwdgtuNBK18EiSoTuNfawkRpvITypNSqDO
JvpPzU6IXH03FELJs2ieeSgXn9o7XD6SPimHMWaGY7graL7UOyLSlXtMxe/2ji0GLu7hllnol932
66t8z5Ws0n2emArxNJhMeAV5BB8eq3dqvLtFR9qk2TNTh9Iss2JM2tPZ0VQ62Jw7NnUjhc/0oz37
Uku4lyNE1osrwU66pVdIVBe8u1tIfN7itbUfC/bbi/26qdo8cWTnlich3Td3Vlt8hkOevqPO8eou
tqn2C2HfINVt9q7El0eX4EPauDZhd9Ieb899AYLyny0DzsNJaNhOt8jClJ7W170GnsYr8Ltq6jvW
9iqzvhgIOFPhrH944Ubfs4/SXUjQvTEpc13E4EA9A3AOknE/INuQw1hQvJ5GSBLA9vkyYtMcQZvv
o2+3sEvphTkZk2fJ/+oUUkyViejhPP08mKtEG1jtFOkHrV96ASDa7z9oxq7oZ1UOveWrw40nz65L
EJLsso1Fk30HiCax7wGnRpruidMs4umzFRZl2ciTEm4/nD3CMbsHa4IgTnWeCsFujEWmcqn0c9WZ
zDHCmYCD7h+KoKa95SMzr9pEGIN7stYFOE4Y+JlGef8oD8D6DcyTJfZzt/wOcBasIp7UyQIPuozL
sCVDUuRZD9snZrpTI56uz05eRwkLPC5yfFgiJHaVQn0vKuh60ub3AmXTMPL3Cv6w/l73Kv1zLqX9
Uni7HsFLU0md/PhKs4T5cjHu0jtlHa2ED4GjRNVJ6GdBYm/HBO4z3NzL7B2ZJeQxFkNj4qaRaGFP
p988VHATFNdyJdOqgRWhUkRYUcFFIX7bpxehQncUWDjHCcYoe2m5rEM9fvYydCBDqcuOxbX77TXx
xMYX9jAbdVG0Ec9PSU6wQexlc7uMOcLUsV2bTZoulw2FTqHh8sACjhGSd24tDyzGyVKKvF0OAOID
UoVgEt8NYB2Oyi1OF8WO3Tr+A/FsTbUARPhDoo0OFjKQnm39ghkyss8/DC4G0PQOxbjcYRhBLF+B
C0q/HGTm8HArxobDqHv2qRK8gLsX2Lh1ROsd9NYmGKjZ+OE+5ov3kUt38YfjoSGjWwn2nttLR95t
FlK9N/ihy4RkgVMois1fKVhnWW+ez2OQRy80W5OagpuhqPOxWvJWBBbkR0KIqky/MgRm3WTfiou5
Gghqn6fkK60GWgqt7tp2HkLKd4XqZsYXVDGt/J/AUPQsXKIdKw7nWoXkxfZggC9icDE2exlt9ncN
C2E9jrg3fgez2s14GIW/eG4rK0z96TDzn20ePJG+nyNoxC2U50bXTKGFzCw+LrKgqlL7JkZj3d1U
uKAEAMyPh81j5gmlZMf39OojUS8PA24W6ieuK1ZVCZtn8GhJFjY/eBsbhC9eFUuyOzKR9sdU+pWu
FLN5dXkA962rY7yz5QxMiUYEciiKwzVAq8q21blirdAsEF77dmEN0MTeLYGETqQ7FvUXerZcLXCU
9mx0D9TpP4klr++fHucZbHuIWnHulrrOeQ/G3Z3A2TpyqCHj6/dyv0tA2fBF+Chm5lifO9wXCJMO
XHaxzQN1xOecTej6lS3GRlWU+um5/saqQLh3O4EtYOLXSAX7Ga9ViWS7SUIoAm3GGLEwrI8HNXZ1
MjDlqp42LlsYb8wylYQr/k0GtV8FCznDPYPGlLmj3gsktOtiToiS9bdCjnyQze+2Ec7lOP/IaN7t
Mhmcznq9wY3SzReBpESRnLCVON7htmaKuqf2Gsrqk/jykIwU6Bld1L030Wvt80N0lWfQ+uKjJ3zK
fc0lwdXnp6x65kRQ5SZdnviyOm10LMKJK9leUwcJXxlm45HjCGZ6Ce6KLBtlhewiTEhhxVbF6xbB
37b5nfDD9BG6GrHOa17cMV9+1X8GVaSItbsuLOlMDCZHMnpTJRlaXkbNw6NuI5YGDyfd2Ghslo6B
iQ9eRTPWoox9kVLa3CnTEdvHraaPzDVWEcwpFLYgaBYkl1QKD5giGjRdbs8Q9aX/nuQAKA8Hl3cw
uwGgq7h9VsjL1aKVEn9GUKC7sDzq5jm3H9KTg8uWeex8Iy6xoxiOHyhue7wRbksm7fjPLxngbCAu
S2mePpzzgtNpTzOR6owAle3JWlwCiukgBsVN35d/QuZxOAKMhjTfepMopH+ibCgXUfew8MvJJE5/
4jiHNxFocmjfKkszxTE1e9Zt0SXMuveJYPb/QoPcaDlnWq/ul4QqF+/UaVtplGj4+SVjoIxn6uht
lVGpVzwCum1s7/C8/JmkyTV5pXyKn9FPl35k89keXzXJXP4YN0QzggeCkE6A5LY2/t7owdO/alkL
2TGLX3Lugr10X4RnKOZjAODaNKiaGP6d0jv8tIEeT/lrzzw+34kbfqDR4qJ9Y87qAVEK3sJTzl97
WLyttCl0yRcOZ9OrOjCPvMPsrMJa410IHuonxXBBLyvkbvsN1IqjoLH60ysdChz9FKlAIxezEu7R
LRP36lDh0Qm1uFYCOFIHbwodHdzhlcVYCqcDec6uxE/uaYghiwpYTyRTBCtormqrX/sbzahEjGke
oCHPHFnGWYHOZnW5MyddwyK6fT++/Yk9auObZTfuKsMjHgl92A+232jlE02Vjuj0hamstErna1cK
247wwI/SDuV4QA+TFZAKLzh3NiKowkDZeltL7YZUrcBJJyf3/aEPHhfJaeaiX6B1/LPhixr2RzFE
dtHKY3Dtpwc7/a5yi/7J25417zfD0z0HZEuPyLEcsu7FASWnXtKXvMWx0ZDl7TMVuvkQdXe18Aio
2rvDjOF/g+8osI/hGGS5A8r5w5H8YLpxANxFuu26H5jKCJ6M0B2gDdKLPU7x8roBPo1aSq+4tzZM
Zj85q9ir60o5JfHB3dGH7VmwHdxpKJ0/bOYQyQlHiwHa5mlTrdD+P/Zx9eE9+cH2uK0fWnLie4N+
syBaTOGSWYlFg/G+sfy+A0tVPJm0R7zYg1MNWrSViqP7wxEAI8BY4Es112hf13rhd3rBQ0320+aM
0E7An4FEnGtY9m6pi6ip8SejFipJG0p5vs+5mm5FvCMDtIbp3PPeRfnSKGZd5EhbRR7vliEeZhOF
COqrooJifwevC02PddnrOUtgGidu6nK8ckjaXRUMLuK3EymxLwwuIb9x3EXtoBRKPkqnrHIZQ4uP
S3ln+fAf1sOiJaTLFA1F60j//n8wnS1WEmtJ12tgSGX8YdQ4l3pVNaJDic/e4MGWWRYAwDBP8QK1
Ry1Ttf0KnvbSSed4jZ/xxUbNd9wBWunD4W+rmM0V26pZXPeMLMSc0TwXBOzKIh69mD2JkYN+cBeW
gLPbJPvbwSl1/FzD0Uk4JfZPYVJ6H2l/i5Kw2xg+f9pv44FGoOdEg4JwzpewbsIHjbzMj63cDdl8
HIgQ17k3lLFA46mQ+Lksr31lUkZpLSP9FGGom/Q0deHIcC8K0YiDwM3l4Mcu5gOhS9XqIGI7xkPe
nSMunWs3uQejE+9emAaau/p4JFKruLIjhTZWpQv8aOjwQ34c6uVvfi0nkvGn1SR1dZVjYnUorFtJ
oPWsf0/1OaEbGI0Owzd+/OWv4h2JnEJu40wLTndZGs0ObUtc7SbdhyviH5uDUoW8mhVao9jAPewt
xqi82g6M7kLaR137kZQIDeXOO8rznVoAnftxMiN2tc4Qi12GBsbgEGKiGpE4ErQ64Z0GRxqCzQJ0
8NAYQjgJJdwPSofVqe7dW9nyq/AM0HeW/lT5ZiRDN4uDMJbQ+pQNAIz2MZFCXZHyogaAbSWpS/WJ
kNQ6oMSDU9W++ZJBPEMwIJjhAqC5PlhTJWlR2Vb5TK2Bco/ELuh4PaNNpO9bwG84nCxZjdSDv3od
2sGxE8KfWfV72gkPRXTLk0VWZq7XD5Wibg7Cf1jjNlpQTUn9FkoLwtMcXQcXPJHqW7uHU/XIZYYO
ErnPLWeG58+j1Nv4ZDUtWRSmbMUzdnyMi4uTGu+bvIC+mB476n4vEt46Sl2hwnEJp4jwyfZ/1wHJ
GnNGIDAXQ2NTgwhF01Fi+4RvY/5XKwBZ1JL2AYM9idPaRjSxksnXcXswXA2jAnc2+qcikzEZBgX7
MDGPWRIxVHTm7nZgQPCnAikhFbLjD0/2cjKeW5mmyQJgCQiDxuPOm9/cYKIUu/nLSDrvaU52yKUe
6HOWGlVD/PDQ2V/BhV38OOhk/hzt6tn5eW56wg4w9gJ0+GwwQZYxUofMBLtTh7oYSLp1p68nHBCD
Fcrs7XEBkHduMMg/QJcRqC7OR00I9EJKP9LGkF1MKKYyM9V0wtoiGW2t20S082lUMqwlXMgHg3xg
EWfIpk6utnBs5Xhl0COzqgUNeZg9keLiTktZoekNK+yW0EMLLl6/fMSIL/leUlBmi+TGOj5I3U1z
9/GH6mC8hM/Bmrg3oIvq0Y43EkYHmEdgO5qSV4AvQRiMWO0bNUyQaz8E3Pi632Cn8oo8DyWmgveL
RTbGqQhfWxewZyZvXaSMyRyZHso4aeBGSZB9I6OmusKzKmgLfKsyNP0epu3/mCgdO9BdgynVWLL3
qzUbrej4eu+7FKRUUDMWvGSUuWwENqbf5ibQHjbWdCLAQEkF01PjNL5si1HVO/h1ZTt3H8JZ4M5Q
ji2/j7aHnCNLkWF/xXaiY6H1NBTtkmMZBeGLztNUIKLcfgXuswgJbDxZFkb3AzI0t/bUeqT4+5/G
p4c0eRkk84cC+fKKyzCrhXr/Ipltj2XnoeZkeAk3RtCak8TuByCnPr9qRsz1HcSru/0yLCarJfXs
G0ad5+AWF5mLOytx1IJvMjJ4BoI1k0b54bLKRFrPga5S6+4xo9UVPKf0NQlebgMjPgc7Ebt9mMif
+aWDdQYWXqwcb7RjismD5TSuqQuxfuEG6D5rWMU8lU6UjWuAViJ6gFoftk3kVJY8hUHiDRPlV7Dd
8nIyW8stwgjohlt/NEp6CmFVL51GQN8vK1ODhZQAWRzJNIR+iZFQhKurgZhYIayQAH3VpurgTRlU
aAZ0EEf1abvQHOGXO8N3qgF1JYsOp6NNUmMD3J/E1C8rdkOXT/rZwdHxTYQ775aUtylx7HcNNIst
aoFuE3fB7vlN+26lnOk5BAr4USEcuAa0qAsi0iKa7gYUtcpnOfBodKGz7tlSSRJ58d0Bl8tF8Tl3
wLu6Om2LTuM9pYdf+uKF8oeGXCbh8Ydg5tc1EbhU/khawqrSGETN7bdLR7d9zpuLXeyoe+HDyJqu
Vi4xs2JT2a3GXEk7A1UiLsAV0YXtHwR9Y7A05vT2/5/9QF8DFHW1WkUwQdNzWUPM4jkFmRBpMXTn
ZTXPDT8q7i97586mX3LO9zsG3SXQMaimUj5o6wTjEshwbiUQy2TPravZVWtcnDh3M79zrJrDM82g
7Ap4lI8qfVKthJBAH8Z797Wsrt5yaHywyVT7zFY1qCm3pqxAH1VF9ZiK2c2/ZLVhnq5eb6ua7CWh
OB3vdPu3guwkbfBUq+QhtJEe2X1eexBkYrShyRnv0mK6sIjGIEU148nfZoZfutE5sIt+u7ZWQ32t
xHqxyj71BHkfQ1YBM/O1N1fdOFkS9XlT2btzo5sJaU8mooVeNvyYEz52TKSqwkrT3UFkF6nUWF0j
E67TMaSxBejJuAPxOJsxUDfwX7l+K78zr3am7ZA3HD5UMKJsTjDU+AjbDhBTeEhQYCtRs6ubN/6k
3yvZGH264hUlMEoqj/VgrDm+fvnzD06MX4EaAf7DJ/xAuIuB9uxedNhjYDNQa+KHqsREQec37jFo
i/K+K/V1ze1+HsHKeSgfRfdFi6lvchwMWqY6YOR/ohluCgKrtynUnHBTkbIivFtNWaTqZxHXqTEo
KL19WDPf2irrYOB/5j+rVcOVXgDMv2CLbJuQRC4V1s1iCqMZ8Pr8L1EzQ5s06XbkKDqhH901RKkV
fZ0t7gJokZckwUSbSETNWuqxC8uS2PCcU72lNW1xnwOpIN0HNr7d/wFsb3loTF1HeQPupoi8sLjp
Ri2UkMLkpnI+RJW84hJYEe17usoLIOCBq9Rk5o7tR2ZHsGaxAo5vkHD1/PJzhXuyPqeFWp+gwpA2
RyVAzxSdef5Afk/iLvmbAndh5N276jqGyHODdsAsQTOUS9gc+g7Xk6aGpi2SmTmqKhhNo9hZK5v2
/QOPqHRMxiDqv1J++J1P+61gEwerYAId6/4oRWWEf+0P587l6lJ+FlAIMfw/Xt8c4SOaWRlXg74f
K5pMTMQN7TkebV8d+3BJkD6ykR4jj/49bdmmJrSuUNrQLYUhbm+Xe9EOrDo2TIext7Z1+AVRpJU5
0IcLLrmnVP4jbAPS4V7Ajvg4om8hhaRTyrqG+SJnQwgoBaiqbL2AvLUuek6Gm1cUzPpOiO6194d0
otTt8NgY6AZmYQM9oBWpN16yxstgGx8/OLIimyPTrk6znda+Ce4GbcrF6+8UawO7P+OC4b48fHTU
78vgIZzvCh+nZyo6ZshfgqoaNSNlUmIBFhMxcGvN3lmhaPa4NqAvd785jq4ScIvEu/MgecVfX4CU
6jahAKd2faEYtwla9pU4t2ME2hUfUkXf80bN/2/5g2pPE8Ms+1CmIHkqxgYRPVgDIzzQvO6bvtKn
zypTRleAOmRzva+cwiomPeWX3PW/a3E6sFPUVArzrSSm3rLZsxlW5hpt2Z/xq1JCq2/cCkgQU03k
8G0h7XdFfBFeRmZ7OSdEfKtWS1HIjtkVW+4q6wfVo3b9nj/3iohELEbPg2WbH6wpxNWc+mR8B7Ui
tezvn24KynZoPANDoCZFexPNjWJvPQn8Swr6ZOCOU1lrxRyPk16gpTn53ukcCJtVrmkjkd2NfSfa
vRIC+oB80XWxiNf1nvjWxnDrQ2gN/WMsbOSI8Pmihz7ZU7/ELmSYDIkxNpYsWLZARHdZR7fBCBBL
FVwL9iAIo4X/w5N86SBX1XYYMAAl+87G5Ce0SOXzL+JA5/E4dx/f0XZFLfE44gXkCUXm24AhdcA0
cJ1ziR3RMrXCLiVeASZOZF1XSlinOh5F/cHPPWFoLbOLJ8p3BEQ8leWIdBZbeprkuPusMBjNigUO
i5fVCCPaaPaultrkki+z5wWMVFzV9u17RWT0js5S3EHlsBoB42IQEzftOwIRt6jY3Hwr1NBOzpNV
2Frhx4TXMtoVLm/dPyMi7x1jSVCgcFPrdQmPe/4+56HqN17zkM+RapT1M49SYj3+cBmhTi9k7JOF
Ce+6q4BLmNfpzS5bDn+smked3w21cndhmYgpCWX4SxK0CWZi0/Mz6X82pLPLAx1+fAeNq9FH6OdS
higAV4xKPMk7QRwCMi2h9rBYpsztrmaJdicRoD+uS9cv+5QEsYnCD7g7GCPk3WLCZQPPRDBCJeO7
jYw1z4nYw3QoNP4p1r38W+QLTAUrC75gu7Fx+MWbT+B9eMLnI5gfYYTJON7aozLbdqGmyTB0Wk20
32f9wEtfCnP9NQrEwuuWOsnWUC6jg+eeR5mmGxajf+BH3TMed8LUS0fxl/TY2GbXEAexhhMGOIEi
RLef5V7yq4j5rzL+XsANKvZaYjQhH1YQp11awndhI5ih4DUGRQfyL7N0RlOQAr+xPGI288PHAtpv
C/7gEZPj52a328Rl9YpHgNOai6KCjy289zPTVbh7go+Re67y2EU+8NP3mdgsUr4zlRWidA3FzwGJ
IbDdGjyH1cZzi7d3emviLq3m3Qxu4Yfz1ojDwY6cWL43A884n+Ba97Vl0PmsSxdLU8Q5mi4BphXs
HlMZQGaH8h5s72VwFdZ2Lg6Wr8mI0cAHX2O4R3/jnUhLSWf0EzWcW/k+g49i01884FuqoFW/XXWP
IMC8riLxafOFrkYzs7b9g0vT7svSsg3oM78/cMv0K403PGbaKuBQ5L2lmECPOCWvtkiER3gwmEBm
E3lpL6ylOSRXtt4IntVwEx85AYU7kEBdPP+MOLTqduUfWYip5d1fQ7k2qh8Hul/BqQLtYO+S2QIW
NPAtT3NUrYl+UJEW2JSB3qoGaDZClhVGZv5UW+hh43SQ6bO6B9irJ+/F/PmBv4AAOZBQA4wRaHRp
aPcmqNj2aMGOlGb7ueRMf8dPwLmUoV3ZefbHmdK6ocaDoPE3YdHEFMg51xZSQZmq4YxrS3+wfNWP
WzIcGrQ7YIXMQSZBMqE5GzsQqasWDtuPTkU2nucsS8NEKS4SPgAf96mFAhB1IR7wK0nz8BJyRFZV
XtA5V8FT8wiai+GXB3JFmmLXgMFpvKXtHCho3ynN604Q+F0nwkuuODAc7hhwt0VuRma+9wGsYor+
CLg8hkY2iZjb8Esu7p2B57YRW6DHn0L17GQ4heI3pv2Xvud/CotCtd/GNDgV3GjPevDFA6HxNQsM
b8l4xVMc9ILhuloN61hur10AbSi/hTjBCgnAqDzQIQCn92ebiH13jkbGlSZxfKi1Spwjzrz8WSo/
z8SSKL4G6KWRa33vqeTqGg1fRumL0+PR35pzGajruGtLJkTxVwjluBT6GDCAsNcpfMRyN7LCVAP8
5TMwVeKxCRpAtKomtllgGbjH72DrD+wf4RUz9ycmJPWTRlrQ+H9t4OuGMnAWHu2RGMNlMQxZNPsG
Si4fUrRKUincwl3dxlRYdTqqW9wUvUB6vZ9yBkXu1dvx5A2CdxmK4UAksH4Wiknf1i7NO/zbJXHx
9X0hKr9HZyzikF4LFCwIwcAA+PcWdezuTpryRLN0+dyrRCb9Kvu67xyoCYWI/4MkjrdGJ5BsoA+Z
PPfYW/AZAuP5bg4V3Ze8Fme3FweLSOTEyprNs7LPrC9rWucm7L4CtkBPCpoQj7CPkkx3ZlhWDFOy
oRbC9u/F2YNV9oNY6b+AO35WWvK8fREg8qPmr/498UzWjitYUyq+TUHlwDWNDq/ipW2lHOWsdk36
2dSGW+fCKLJBjqZphYyNBxhbP28d0QCuKzjtW0kAqim94ii2sGccFf4TCxGt0g8CTLRJDTrQnrzn
n3f1g4lXVZVoVqmiLwRLg0DEhMoi8tinvc42KOqOYa9bon6ClGc9vlews23sjPJVhNboUEgp59Dx
NF2FsmmTNRZCfepHNICtaakPUfs1CdixGALjavmGzYJ3NwtgO1nTb6LJeNmiaKcRhizdLcFtWk/j
2nMe333AgDrl3ZPeQYFEPywREBtDaNXtyfEqQM33SXwH4IYHddetXLSD1kYaAFFAkewQAhIec28J
l2WzOWDMVj/HQe9Dz4WiPs9eTY7OiaBKRfNPVN+uYtWf3cM3ubS7wq9Ug2w8mgpVY6xPciOBVxgN
Vu9/HmWv6+oBT82nlVaMr9fMFYy43zSbkUSm9jf8XrNlZzuIf7xVsvA9czFYoH/u10roacD8RO06
SkLzuwdM/dMKm82CnnOuYMpSx65xC4LlkkDyfspZnRDIDRFQpST6Zq9uTBh0InHQ56VkIG7ubAUv
f6OolbrR37kRzN5XBsJsVrw0cOeSsBn7siKEpskKKRwBaUfJC8dNskpSIUf9KeUvrX0z2iYepJi2
5+ryD4Z8h1NhJ3B/X6FkEEeOR2tks8HEsjnnfNmhoM+foqNeb7nCVdmi0pHIB49Uc2r0aklpx5ko
W5a1XcduX+UX0Fkk1NJAGPiE0L2uy5x8Rcbgv4QcDe6eZJgo80qSyfOhE4FzY5jMKseEyQoJHHWR
wiwdRzrfOhfco0nliOUahErcASjK128UsU7vA5sQf9NkBtih9U2JMAE1oFnOyoqeMx7OLHGeZMah
LasuKiWIJU26M4uUicqK4GGokJQ/fvDCkMuJiUPPo7vmMwpkF2qunvzzgBqcPPSfEb1vjoSTJID3
4YJsurpIRn7RgoW08f+72Pwj9PcmYYin3t0fTb6rb64UrTiKOe1dktYeGLwFMolkjhHJYgUT957U
nuPHZm7K99aiL5lp1FBA43GC5OYXkLYwEJgZwI1a82T+6CvUMMIkmJt7Q85dksh0Ezg9XuNk5WUU
X5Gsrq50A9ztrUAz5Q/qTuNtECjVg7XWf6y28uai92V/dSMxKwY008ezHbJuFDB5lFTPlOWpDRGJ
Q3VY/FbFbcCTwuFfTjnPg3NDn4LLpNj0mIeP4S6WDYaXtF9nbQuuaSefd06Iae6May2Bdyqbxr0M
QaJIGQ1wfzB3cNN0pPOQA4afK9jNDkbw/4mxRScet0OmKY/7I4iJfUg+9PLmiJyXnnWTrD1TMeSq
/YB1eRYaePCJMF58sU5mKEH+TZ8ak0NFu57VyM/yifEwsHtXy8jNon4lw43QvQpXi3ss43bkliaH
/TVutA8MTk8unytrNfJ6+T14nvvZU61XKBvQqDw/ZKeqPD6eQrhbQZG1TuYScXRX5Zc3aFHCkb8Q
XfhOvcrmK27yY5ri7VDDIp+Zn8iWOQQshZdMagh7L2/NF7G8JA9kaxQXfWyqt8kAe41whsMoQuE9
S/TMtm6xCLUe7bB+x/gv25RNPtZDoJEZkPUtXfRWn0WB0mDVXbVyZUwP5BkZMuIHQog024KPGAvN
mbkM7Kv7WTYSJnbwoWoUdpSGPh609UjwWl1iy3qsded55Y94XY+RqwyMboelLoxVb9T3TXm4ufcA
l4KUkYV2e5UnW/cq1D2Z0mtNX0DgSk4K92ebhBH3wXiXe45UROk5VfLX8jsVXQPgbItr/N+uMT9t
AqEw8hrt5xU29mum9hgJNbIScWNm1QKsOEC89HSPSePG+UGcXGZRMtgmH0RayLpwOxxD2sNJFDJq
EWtvRk3akE2HeqMxpinvwp+fB1IQ5QZvcqeUCP2YflXICSzw/s1jUOzIIVFXOEQPA4K4A3VdioVx
iKGrGtVwrohmp5kk1Z6ovYXodKeS+guL3OMYeXrGn+cVVT0QCC15byxW1Ogjgar014NqZYZcKhvd
KZaSZNZmWMKbfzuppyNRjo5LBQzYqddl2EacE6VjwnO60cKNGsSvoa/vdr1sneAEciE5/iwDn8Vo
GfU9DKFcwf9evHS47RgvdjCsdpjfF8MwO8zOHysWct5wjtUoTwVUncjWKnhphDEe2VzBFEsQJk04
EcwPCCkPJPFmSr27ujNSCvL/B36J3TnnBFdjkuFI/94hBrSzr3usE2B6E6I1UKyt0HeQPA3ZKssT
871FdhQVbpXSPwYJ4Zu0L/i7rDJmPijrUMuEvsJpFsJ21RaWvN3LohfFD0HXJjagc2iDOifXM0i4
MrfrsmD6Z98wMP8yDTt9GgF/pfWd5fK+/ZFLikbUtlWdRUTeSSg0wnR/bLoA1raN6E/DQ7lnwNhy
1ol2OdqLXlRQI1xRbZP1/ZntSj+6itMMbpZULi3agn65h1RWlTC+xJsPj4bG0YJZgmVjClD8295a
+HuU2qOis8aScISSnvCKc4p/0dZaJUrNGWMhyNStTk9sZt4R0SMB9wwPHjNsiyqdZrz1jaK/x2GZ
9c42CawXPjgDBfy4ymyyRAcqJFDi9pZZsUDnyDoawPNSUzu6CrveWNDkUP2doQJ7QdNcXwEAw6LZ
BP0EBtTkYPdoDsONxPEiLIrJOKiTp/yk77mPUcF5BirLUbBioP/EvRRfB/Tmq7jqHLuOis2U2yDq
uWTIpibsoG9usoeuhjRNwCbn1X3Lin2vT7cjWnTRRF4Nd5SP+XXCbj/ng/KGtbl/KG/zhaU2PzXL
JWsuY13lzF87sseE4687b3zX7heYeEGkJ0nwu06T0quRcVq3iR3L1eYXNw0lGNLoPhLtX/nr9Jxg
eAKrFMpid1SjK54sIfvJBSK1mzAXS+3IQTSNaFv+EV40ivDt2wPwyJkgSJdbpirMiOyHHkPXNGRN
AOq4L/yeZTX8nEhAvxSjG4Teg+mgLjVdtjQsZvx3rnRsy6z+BIp5KPE0UvXjOToi257EVvS2iQvo
GshzfousdorBk6/5gkJ0xnPCF1CDepeWQD9KZxjak+wKQ+Mw08uoZtMi7LbK/o3aoduoneOUSkya
l55yr3M37OsjI4861EgG4rGm1VSEXkO7BBrTEyxXxBaC37KXSfE0KOL1m/+QuubmLWoxLVsVqPpx
KL7CZHnEDoqqULuWO/JCyPV0Ur1tFh8epuprlkX0tPwo/rf9LI1nxSdP4aZ6LOVaqTEQcPw+UBTD
NGR7Wjff9MwC0Mhx9CIHIdZNI0yIRDeafdvWdrlsQj69qIyO8yH8iN6/ePvcBqicst8h/UqLty4U
3G4/Y0Z7I5E5kZhCk+fCsJFcvDf14I6a2xDjZmfyPmgi5sN5gMIoC54RXYr70sbxl4yGeDBBk5qv
4KSDLWqxrhSP6ffQBc5ZoA4zaInrVUI6gzOB1e8ah5mTPgyzaWTtBicK0zs14Un8r1nL3hxhOB8v
jmJ1v4zL/oZroBxgB2zKOSTnZeoiVwkmKaTa79dkOMF+IJbi8OfpqlT9M/YPfUAzFBeH4prZrnqW
PG/XRlStMQVAgaORMKMn0x6FFagdPjmEUHP/CE6NxalgRQQf8GmoF22UpH+q+B7rbhE0tPHNnA2M
gTl8nSrqBWZ0/oMrn7U4iks1X5zHFvd2dhXaUl7Sc5ouMiHFYeToT31VZNYmzOq3QHsimAhpl2RT
qeoDMH6cM2NuSE/6xuMdGKi9lAp/gmzAC5JT14NgyzlD0MfFjQejTIMeXn5qvojDfR4Lm79SrcJi
+6AV8gYUp30oEovHTGoZlPzFy/I0HwIc8/RujX37866LH5+0q6qLBlragLlY91uqvjkMDhcRnE/l
q2iEqFEmIxjJLUH8cj+7qpoWdqBeZJorrcxbQ0A5vezDnyP4rr3fF0lr/stTm7b9ZXg47SC2aMM5
1c1J05PqPZ1K5joMfWzSIO7I7Wl9h94gk+YVnSfpP4oM4uNxNupTGLSyWltU8I8DcDNO5oq48dFE
g5fImxwdp5dPThrYBu4eSYlRIwG7tVQOsHP6ozSRabsuxcqe8pRDVuygnBoWD53IdjP6jgpJGswg
Rfu9kykpUl7T7N9Gk+c+UOvoNkhNIXBYnkB1y18ISd/nyLadZhEl0V3BR4288xtZ6HeDyVBZ0Zow
O6fLGl8nWeOS1aaS7L4uIc18ZrrGyyRRNugS7akKW6DvIejfrNk70QCpocecQ+c5KcbuldynZVn9
4JRDqhC4m6QDMZIeog5u3c0dtJNDFIJCgoa+vWc1LnrnCp5I8G3rLmVF3+PtlmX8etg0uBSwITQY
8UzF3kWcRao7yqCP2zmg0RmKsV+WaCYMGVQJIACMV5M+FpgjN45SrqODYANbCgGe26O6w5c06yY/
Ef9hJHaug1xUS2DIQq6RRJT+AlWWf33P+GWvGK6PoE+F/Gehwil/FuMyCz8z7YxU5+xTCj2SGXw5
JTHESr2MgtE6XkYOQYiI2HYUiuvIriN0RmG4EFbGIkv5au5LUn0LYCnXtxoEhOCUIVk2WfTouJC1
d8oaem7x7lwfpM3YtUjbQ9ErVsoWDLSacvpT4HahZPCbvD+7a2X/r4bSRyf/FOhvG/iFyb72Zleo
Es4cNQFTSTIkJv2Afc9A6OxDVMtc4fiaLPok7ZFctAFhohBL2RmyW07YAxHd2C0TgLAr3Txbt8Ks
xs34FePxAmkvE3+S+0NvCY9P+nNfs+R8txE1PDJpS6KXR2oVMbjg7IvaRP3vDWeqM34s60l0rHEU
g8rVbIgG1abpXIOAtVranj+TRstMS+VITpTKfaAnxrNqBof6GrAzUyS1PoLEQba5eTrogAOf14Zb
pYDJ/aiTrrgWaWljjnnRnvRp9Odi/VNMdbTfY1Q6y/1wJD9izIyRvQiTjkL7Y6KPcE6eOaWLpZvi
xx2tBs3k8YfvglTrmt4f4fYEWH+ksR06vTZ5u3brZPlnW3pSxP+XiI5H1lXDH0D8n1Rd9H9c0ZC9
ijUenwIDwuRoqlf+OsU5JczK7DBV5ylOxVCJg+Cjy4STqTi2UWzKXKhez3do0CrvnA5rnGOaqzYS
jeN0+cORTfO93zy48HfGUMfxCPg13JPCBuNIZ1J1DOCeTSfyG9VzPZJxyq5swzAaH/aPMymHN8MD
Helw8ZUyZjB6po/6XuDPp7BwnDgjB7rdApVimeVRnLaStQfNG025n1pOltyPcoFMpXeL6wSuzW9q
sxnVnwFB5nWaAOGvh/OenOs5PVCyTA93iibr/WTfZ+LdnYKyGf55eakjwokF7ryB4DqUL0J4+WcS
a1d3zzWMC5TmyZAn0WNAX4wSormdSF21qvYWZ3xqUGmGUR9BR4nsOs209zphW3YbJCdYH4P07Sw8
GPQWvICKr3y4k6Kwjc+DoR6QFuFwWmUl30Jm6YB5w8H6P2Zp4sHh4G56QIXBP7aGXBseKL7QTDjY
WO1QH9EI4ZqAq83y7eD/ucEaDGNie9aCLTWxZwqzlbasLQviG251RKpm2Id/YQeZA4Z2Q9hQiIhQ
1D2rXSPsmCV2tKnmN4EP7SS8fDXnHWYKWe8K2lKbn8HpkjqXyBCihuldR3zKaAJrrsV9O2FWugzI
YZbzQKgsYOyhwAxiiy2ox3f4UlkDZIkHKylMb2SZPlSocgsx0uKSPTymg60Jeoow6+lFrm/OCEt1
H0FA/O9NOW3XpgYAagurC3y9eOJA/6F6AM4wM8NJ/aKDejTpaZ6bNFMi/J3acMdm1RGyVuZcEg9i
XrSdOJS3cRhOeygB4mh6Gn0SqjJ6J0gCSrJnjfjHJRZuAENslU8U3xT0aQTiem+/32L4AlR8Stx3
Pz2coI3pzZtUt/JNRLFvM/2E/OteY4ETXLFGfrAyajboT9Ngqfe9Q1p7nOjKr7sjZc7K3PwcRS5F
Zph9ZvP4DFjjvVJVoqtf5vWGpPtOA5FaUXfBzVKs2YIIJ/0/fCvydaMkdGSJkENoor8eZH/AIytc
bclO2hzEam55IUqdYAGtPL0FU+33TOC9Utb3xGBAYaTUpsvuS+p1LekX76kr9R0LiycxMzu7Yo5n
BkWXBSDqJYXAMt825N39DClf/1RLH92cEB0qVBu2un7+DCiJmiITYtjkP6/Kc/21K8Z456q0rhaW
De7E1c/4pDt5DZ+W5Q+uf25b7AQymAGst8CNnlHiwaxNYSoaMPngVOy85bdvvPfj62pjuWMw6gd/
QNvkjR4vOr4zoMr1cwT9sXiOee10S/mcKLMAbBFkVLKIRfMmzwfZdu84O30GNvvMo+B7J+q3YDiV
LOY5MQFCawr3Utqis2kH5EWZAxkgwbxPZdgIbp4t2Q9ram5imccJCWJf9ZClutUrHQK42QZHaO1W
J4UVPnOyXDEs97ppYdkYAl664EA4pu76UeJ4RdDhBP1xMkr3h0oirgHYjdKWAvUX5qh5AdCEtIGm
7nEX5AD17d/IV3Z8uHDhuHQ6LYfbczIpCl8fEE1v+hu9+oWkO/m1jJ1eNBwUU7xku43LKzAA6+rh
pzBWlSyA7hhCyXDjybtw/II6HKpCNCiX7mWicdq4Fi+1nyGaSlMm93bTGMP/3iI1DmTDcvZmI8xW
hwYUvFaytHpSrjoaO0HvLu76jkRC1D5wTocPJZXNIb3MpPv1Cc30YVfs5cAq5+jdSJxt2+uQmfr3
btyYZglQDdrS92/mymR3bZJvxhWZhzQ6NiTr1sl2CcdIZali8upS/A150qglFrw5mhJIAG2Ky8UV
TzI2aErWb9KubPGILmPrBvcVwClMaM8CinxQqC7QLPOahmYxvM380NAyDF75ssx7wqwClMp4+JPz
VRGStOaJVZMacfpTiqmWdxLBhAc2LMIol99Gzba7LB+jS8uD9UuH0SGmw2smhvfQb+1gIfoA10aF
ZlsJCCbRzlyw6s+Wrbc6PZRwp8vToXrLpoyEvyEqfnJLP3rmc+9oTHnkSRIdE74jK+eL9KXOrnda
3d9po46jPyQj2TmgzcYu45l8VnCQL52HYS/tJiR0XSBDMXAKRhYm+NVykEvfcM1Bnv/hx9GrWFml
sjjfQtHNGQAa/TdCtVVGc+IF0FzH6W5RiLCF/G/njenOxSQ9RIAvSyYtjTXxFfVaDC7T9P1oqaU3
eTgaj+XXPX106KOOsa1dc7b3CXP1LU+93Jys5gyufO12sTWBcnVlzjo0SG838EuB/XKfOl2/++bo
OvsEV4TexSrR1x6Z8w5JeATv412meZoKQ5mw//kWEMnvv/h16gaLmu9Qjnv0NufRszQTDX/j9aiq
GPynvCqzUtn1mIRtgf/hPnuOg+tPpCKFvsFETM6TQ0xX9mW6FTzXNSgTNgQSk2dGatRqcqA8jYpf
c9urjMBCfFJbzknHzJMDy1erxdTijBejAprn8pyzZDOR9+qvAbIi9uaeoQI3MFrNqfD1WIPr23V5
buGxq7wI0mtR/AVAe9Pps2m0mF/XxibWCUTwfcnhR79tVTxDloJJoyH2xoXhXWcSFZZDLGIDEJtm
7YmE1uHvh0xZXrG6UGM6Tqv3YMKPXqqbi5Zin/4Y/bYPaRoCVTmTOIW02lDrTsscqQ6NjDnjGAPv
xENMQ7OlNDtvdO335rYDakYrmw4WkNgedO3WmvFvMRubk3J2Q+ORzFcrp/kuT7y7J2mv/DeCcca+
VlAXNfZVsBuVSH7DkGESn+C5hTAW4fFkwGJ2JeuwnZHQbsOySiISO6hKDNLXH+p6YWbKa4Aso0tS
rxloFPqgr764Ya3qkx6DXyXlQN4bfLezoee+SUCxMdXaM3dv4ZKAaX1KFfnlneUlD9Ijy5wwxw7Q
z88tJUYM11zRSK/cAbV63mSqXgGegbAz/MIJv1kweQq79PMqXcO1gzbd7drM7kbc2xIeqa2cAL+E
R6L2r8xCAx0FpAacl34+nmQ1n0emZ67mirp+jvY/ie/ya9V1GWLZ4YKECyC0pof53T1xMAiiF2f/
K1TmEVTYlNBEoFc+QKbJsqc0lifnsgIm07+rauPsdwAtS+HYxVAhLA9VE5s4a3tvLzBh/n1Bxb0k
KSS36l8YWnIRVxcYWCKXAaRk27heIf62kfnLbBNmxkQ9jQow7TTy9cFZ3S/fbgdZ5mNBcKr3XXt/
RA0kFumaiJjpb3bnQsS2ZmcdSavRoYuUq9LqneL2Ny0FPeNAxpnf1qrSZws15hFsVsAiB5uyOS5k
4EgfPY6va2A3o5JUXniuaWcRr7zfQLA0VjNdV+EA3l6Vu5fTy7OqNFjSEMUZczwO1oVqzIn5DHf4
h/BR+EpLsODKBHv03BaJQf/vb4QTmYnXvaNf2ZtoKyB5QcM9XheIZhdqnBJlHe0rdRYP9AKtkPPG
n7DOq0zTTU47h/FfocWMDvJfC+4hzIjtPLZFYnfhYRVPm6BSlmJczbx32nmSWfdav6hdoBzDuZDJ
j1NrA4LqHwIYeFCYX0VSnHfWGCu9JI+OSkZdx+yF3oxfym7m/RpozxA54NRtpNJIMzzrIeeqMaLZ
xJnd5kp77sAwoSf9hREGXExcr3CT/jmQWa37FrIBsoTp9yMjeA0UNJLUMJudexpcAMgL9xzt5yyN
NeCmAQ1RDIEdjgJXizh4wLpAAK5aZ2xznJ9+Rt811pi/cTKM+HFbR8J/5Fcg2l74lt+aePdwIKIV
3i6kxlsbYHCvxbppQJYhnGMr4ZD3D5em0/ZVe4KHXJcNBbPV1ePQGdY36wKxkq53BS8g5w7qg3wb
xHYxTBhbTdRSPQiDeJH67EqMW1Tf7/m5rej0lWBU6VBBwzh3sq6gx0iWw8rDGLV0pXNDSdaae0Dz
a135SQXiyOh27ec5k3PoJa8sw3lqxQnpnxy4kKRA6wLK+X9WM7iCuenQhR5VMGqT1GzNogrbaIZe
yqInC6qHYERUIV7XHTD05tBC/VxOZ0rNxEEE521Z8AEqf48ni9LTRpkDqNA9/pCDqA9PP7AIYs8X
3jeEbub6ASGbieKMXH0WwRo6sdy6fhc3bCwdP7Guvq+oOZbJ4wNNSStBv9y0+eWW9K1JPkz5TeBC
9x6SLyiZQNZEj6JajbLnJECbSnPGcEAEnDXzUA+qBGdOcD4edjAWVl0l0lTBVg7rtVbefPrshTKu
EkNP9cbmkkD5ht4xvT+YK8+ukeb9ZZWNtRtYCZXIkIgEneXtt62L/MfoC5LIMFqvD3IvPHDFVyKF
MIY4kZZdhYTLJhjgthwK+GkEERy79M91J/JkocC+ld4SD+ZsC9EXL08s/hSyxSx1tBrf89doaHnp
/e+V6qoQDOmd3d9ztJ/cY/CBL9kui8ajlDoROBCiiRCjHJksOayauamZy/REmGxQrk22JEdKbTTq
3Xc8vS9N0GQLcoh4vymJdUtDBvP8ZrBcwhIJdHcPjGHgF3wIPTCdqjuLLgpJv4rhGJe99jK+GoYh
FNyNCd+lQlc5rJ3Y9DxRNQs1VSW6UqdT+UgaSN5bKRBXZui+Gi3R/kni2ifyv8zPpWCf2S4sBesv
fZ2tdPy9/U64APF+3ZQaXWa34kd1aU/x69nPj8J72S41ie9+Nxju4FmfnD+nhLawB4JFCbGQ1APt
FD1GXukN2mj1MWX5A14B3+XcNZqEWFBuSHrR/Yr8tiSdVVwhKDElFWPgCxctEWkiwJWRa5GnG7/R
OjvBe7n689u54iiWaZ3ehdfRLCZb9uUO0xU8lqPzAAh6ruYSFTAFLueX629rkdgi6VQDIhktJyQc
oLf0hRl37PLCMpdefeOQnHYdJTXDkp5aKkyFfo7kxL1e57QJMNStkDFb+yRCxecAgQuDe/FfMPCk
0R6Q7nIsNm789hMsHTVKtzF+0x8lpFClvfoMWuulGHU5V/rTF5Fk3HsKIs9nv9bI2OGzxYK0ooWD
dcg+WPucCPonF33BBs743VYeyE8VyRcTno3c6s3SJLYC6pA4D35JWSctICnIvAF/nRlw3GZbfClm
1hFKXz/Ms2w8Ij2P4+TCvc0HqSZqO9/OF0qnHL1GuUQ/f6ZJ/cQYwwykNBOQk4KD78TsQVeSgx2K
5uA7eyBkkvkUrVoBtjn4QfovM2AXKPwLk/VEnMy1nkALpYXkDoWqRvRxjtQOXajMzb077hjVZI+3
cqqI+FFkWHggsEKnNksSyDogzg6SN6epi2xqPmBOkhq8pdc0ErCij+2zILTFKYFSSWI4vEpZ4gFd
SspQ7MXMlfKehjv4TgAP7tq1Z1TwsEgb4boakXmq25UligFOCxBmV7P0fqVdZGQMCsVlLtFZQfK3
XkPknvNx0k84hNmtFYvvTGy8C0wrSlZtcKmUGhTwyuLkIjalVkQL23hxVO+qMxVR9ASdnUCSoo7A
Rcmuk71WDkLMjH0qqaKzuyVpVsEYCJG35k+kgvDbgdlskgHuZo7BsKjruvmQngyQCaReHDCAYb3N
2G4Q59kxAGxsRsVIyEHxTRpKVo6/ONxsZh7dv50V5JJm7DIL+PtEVXP3H/K7TJiFkHKS0MazrOaM
MBlzBXUl/Ir9VRHPWQaV6qqLgPV1RPn5atpr5tuDGKx/shjHXBppWT233oJQnFKclH1Od1F7VEtG
5plp5t733uSSa3T3K3VcAhLJVnj67z0+7l40H3I0VU3YlWJ4Le0Czv5UeebNh0juWWJWW4iMK1w7
gTHF2dnzj+eq7ytCQfDA44EcF/DzuwEmk3ZQkN/RvQ/BXvlpr0gKsnaeF6fcZJ2hC4fijJWBh1fQ
zxh4EYwwQu+3QoTXG8Odu6fcef8ap2djNV+Jg0uMGhuAZSea44GRB4yw+AaUhE9g4uLQ3vwEofkz
zwtSrY138X7Q2o4MqxJrctlfQ0Ms7SifU/0muXG0lt7dGtvddfEUw5PwAtf+RsDriLTIgdFVoNGB
SVToViXarZHT3qMQL+7L7cdeKrHr/qoflN+Wm3UxH42pdDW/q/x+1vns7Q0DaWNyzoA43HzicdJK
kt3ZB1OQckLuIWKMdMs4FfQ5o5h95+pufZvx+4OnVQii4yYtAVNg/cz/+CxYislmUJ2rnc9oMej6
azHe2xvaAndzfSV94gfUbLEX/ZXA/xbPFLCIP6n7CdVpwMMpRWCgnkXA2W5uEAtg2YF6pZh0anwj
MTYBQpFhnFNa2FpK2lz5vd8xil5G9hwsnCeF1yUDt3wAp2LlXJxu9bMJVtbr2C5w+9WUoRYvCIiB
MiSOdau/sJaEPqFTMiiYTAwv1KRZ+OSe65LTEO6TPCV9NGtgKOviHDXjgYWDuQ/+SlPRZAg5peh/
eVLjAB44nc2KT3GB56enu5UAvC8dJxDcmQ5teXUmWfFfDBQx02qFjoYSz6Yn4kYwnBCuTa+ucOaG
sicTQBXqTWkzibQpx+8PkqaVBEFjaCW8HqpnoieOktIR3ofE/4dZidhHBZ3BjXXxD9MWeiSQc7rp
ogJpxn0f7OIPlOnMA9p7eXHgDS7eHr0D+LcK7qwoTAZKlKxAd28f1x3HMWXUyycOpfNgpC/Dzyum
R69aedfsgbhD5Xa7BUt3RQ5WUbC0+A8c1Vtomly5lhh0krv9GS6/1yjxvd9/Jwjb5erkS3NYZ/1q
w0xLlki9XA2RHSlY88DtQSwlQTJDa4czx3tffnFK0ZFBZCxxSFd5MPKEDGXwWwu0T9AAmx0Lv+Ie
MhJUd7FJRtbncpAYi3kOSW53wp7Xivjznhx9jQNCD1+3kY88YUWlu+hVdGjkm2ndGSryFM+LaML+
xs1/AZ2DqiPB4Jilmrl4+70Xn3ncaGttKil6VCXk+/9HdmAhl08eMMwKMWO4B03PJsO1M+XpsRmp
zuZ2mtJLJnbtcaZfg864BopAIhEsn8j9bBWjizGiXj5bd2ceSSdKY6UGq2033H54H/8rAAuKIzE6
UA7fZ/Hw2n6aM59gKlXT7BfgqlWEzXgOasAbIO5UBVubWBJ8igm1Wgk5q/8UkxJN5vvb962jANQs
2jyYy0viPIaECxopSgt/GuaZm6Dorcpp1Yd10iQMQGC3cdLHVE+E/7Fj5/ZGOI8jMeA0tzmuy+hp
isWPEHKQE6OFr0d+cAmeWcQsnGlwHvOUriE8tiy+I5M0wZLJrCsCCqq3Jkj2GOXCkfQrWE3dPaCe
ED/WJrKVXd1dQlthd5lUCbAVYMAqtPXUGk46P9wpZ3I9CbJjvH1NtlJ+qnN3DZXI6anJEgpZjlxw
YDA5HozxsX+oJacpjiUXysl+AmAyijBt/Cfs/IpWCvFHo8xZy9DRM1NW3g6oRd8fcK5vU0EpgIdt
WF98rArAC0SigbTPilaVYrMFoS0gu5ELd+8XuYTFqKvabDMzZ/LEhGdL8ZhlbPf7/1qCv/dQrHyg
arftFoBYCQ8/pKXlKqRglHca7FeacRjyuBRpLbs2ItY0YCJHarbofuQHv/hP6qTeHPtKpahPObYT
/H1Nagaq4HdPFClAXHTjoYQsrbGjW9xBYatTUTh8rYddtT7SrdySIjR3Yq8Oggt7BuMSFJOx9kxH
FvY+9e4x9dEb4ypFMLUouos2eBgYRAfq+D/iI30NbfyGVzHsnePQMjwby7JcUMB1iTImCED6tB0Z
MnG+xhdgVMEQRCaPCksktWELjBum3ewnjtnICMrCdCKf4gLvWOPyl3OUQ1uXSTz9nxb8aTLL4c9Y
MIWOuQfk7P/p1QwhVdKDhQ3/XAloUzbdk/twu1QhbJHFihmyI8x6vWzZv0oN2NUjPnUevewl923G
2I4le4mm6WgL0zPMG6laS5im7G3TSYe4iBHbykc5KWuSUu5neIprBeJxAHEx6FbgNdknmwSXiZke
9hOgAIQP3YNrEcVaUHmxZnZ6wf0cVhKb+6KYu3wOreCXI6DjqTQGUhiwxHc4VCaXVWp4f5E6qPkz
9uCMIC0zZ9bG8iczkhtyRtyciL+veMABAD/7a/QE4KR5OIgtOFYsWLR1anQb8fLW3kvHp/hHC08R
Yyb097er13ruW0z7i56U4KBQwlgmx7M8OaG8SCf4oPHd2mDaKnalVaJ8VEaBIaB1YVGljLRJPx9w
+zi/qbqwz3p0sl4sXFh0WXv9md0hszCc/kHU9TY/ohkwhvzLgODLuVmEMC73xtxNhpL4KftnMkr4
/joZ9ZB9r3c+iaZR74tzWgkmLYgv1FTLCEuCHw4gw+aHHyJAHFLE0vjGBssqTaS8+YRPMt2PxBSb
9//xCJstbhr1TG89JecVKoKdFIVjnCRLPyh4P2o6nEZSV3r5fIEi/mjSJB9QUt0hehNBCqqLsguk
tGdX4lsuPS92zB5TFK3MFWp+Q2Xhz/BZz/vmzXtybwblwWpVXawZjkNVw1sSbgaA1DvBHHjWNaqF
oZF/UZ5SWBodsbw8euioh1A+XMjWnMsGWWGed+xQmom3gFjpjULWBfizMu1fQwALzhsMQxTGqRo4
qR8owR/UxtzWwMJROcZWvatNPYbE7scflloznuNb6XkCNZvmr/jw4gQYBcLqwfhjuiKg/pCZKKhy
GB5jYabwL/5opg6/yHZv2DQKBLT4kyj+vD+B5xXuWhcZoGGjlV1D1nlmq8A7lCwJTZwJLiRtLg+S
KK+sFogbP4PhojXQS+XtjV8OUNATUJ137qSefzLMTZZX3ybyPQzZdsCB/5BasLy/r4gRHbNp/bmT
dATEYTJ2kC79SpYFoiLE/4mIXjMePvjrLY16UYOaeylyF3iU4zdBV5GxOGZDGk9yKOYUCP2buluq
woVtWEWBlJK49Qmavti1diQ9fnObHdnV3JajjsUL4ODx0Z6vGFsV6GioclXZ/ueHtk1u1pnNpcMv
hzVrLQHNo7lLxdp8lCzxpK4+YUQbxyNfxfeTRqacp7iawa79k2Zytzs+3IH8WZKR652dNEUjE0BJ
qRvbULoYYRiOcfCFGPiWF5UuR28QrJykBxRmzhEiWpMfQxT0Q25v+DBkgsj6r6kQc3Ft45dFMODZ
T4Z54sMrvxUYktcNrRhqWeOj7oD+xV5QVCvX2T6bXSksqXmQ+Ab1uKXdFrghz8xC7GNtBFCTs0XQ
3Oj70ljl0v8tMdy1UCBD3A2jPopw4S1St4RnC72erhwh71JtCrXElz+TJXK63hCOLuhdXxw8N7L4
46HSIWDK+PutY2ibSVSPsiHv68814Ze+jBud5V3xy70zekxMwS+12XRZljFC8SM64FCbxDo3CbuA
P/zmiMv+5XIM1OA7xtWmrKOeiDxlThJahtvxnTUmhMfaKd5yC4RfoqkAwnsrE62mHXXYRHO+pfPa
GCAEYVf5NFwkjV5DdRyVUh+0MRUyjMygZAgZLzCvBLv2fTDH5uF+Db1oI1BehReYUTb1mbtHuE0U
BGezovosURe3Nc7mIPJTCodz9o4OwlTbUSLyhjxmhn3aPTleKadFqkeJVX4M+7BJT8naB2mRFrcx
r9bbanwz3LqfVSH01KV1WvxI4X3nrFWVPpahNhGY2cr8pqht/lQvW/9E0JRy5uGiRCBhZzOql4bQ
DIx7Ja8MZcYrvGZKMRNdFcQWsVElV7YVKgrwe/DjecvJ7lYQUS7ORbtH8MVH6EXOUYitl0VqeNIi
3s5dKl1Nas0WXdJev745BttqOB9ZPRbhvLmUJ6oV5AJXe9ZDZktFNx4ktZmOovqdAaL1j6joyKUL
Blk+edvA/tumKU1XBAsheVot5QOrYZRGJevD5eSTj4g2ORIZyhCqzk5ySCHLXah1cjHO2lMchu2I
4QVBX1iCPtVFCvXS6FcT1rzSUXjoYUjWBBXma7QiBBmgT/lfHAtsr8KgEM88L5UwNGuuS/2q6sLu
sr/jxj0sIHGrirIkZOVHkqm3ODqwLVfhbLcryro71LxOsYCuBf4WrlYD2wJYjhOL5v0u46xnjFPG
VfM2O+7FzxFa7IqCDXKGK9NqUXaksW/BVe7CvUg263zAO4zOAMBQRypvdigVLfiyPQ3d38TDjRYm
r/x3/u2MpclWfNGoG+qY1ys9gcEHJt6w6bagY8MdZRc5f8/rZZOxrkKrl2AnuwpA2VU2t+FqL0e0
fYqpDmloUjEwMB0NZ0ocKUxttbSz48MWW1V0TXarMZxMizM/BOphh8uHkDccPjbu0BHHsNh/xAXC
6Vkuq+aTme199PDk3nAsQ69bCbrbGWiF+gSQXIOd8JnDvJwkZ1wK2/bR0TADy6Rj60OaAIUQfA4D
L1uKk9TDHz0aLt1SBy/Xd/c5lwaoYrFbfqJYsWcYjZiuRKi7z+pS4he2Yy4JVjTcVQiWXncbtnTA
8id/mdKh6lu9jKN0uzFqGVzeKyHx6gjr2VyG+PV3CYUyIQ5tcxhbbogFEAq4lUc1YGvHwqVRFLws
gA2KNwx6pNzCBXdvpMBRa/nA2R8nr49CCjJ2nDLitBjOeDKqWdLK9BIjZ4aJdQ7S21k0+6pkk0sv
yQefbSHYURxvSC9MQjxmDdGJZXfdSZCFbVwe2EMC2k5uJRH/QfTk0o9hPEOKit8CvLdr4n/5oxGj
wMmWt6k0xHsKMIehw4fHbbdd0NXUmEXPiGHO1wF692RRABg6wHN+zMdq8Tg7OLOa5NpJEaMCmqh3
5i/p2DFEchIdSlFsLBvZ5RFIt0tK6nIXdUXUsArQpObb8jtVAGkEf4jNT/99ctuI5AOAZLN4NDEL
tzb+/J0/FS03Hy42mS7Ne/+qVJ4d1paoSmSsLKsW0ctzSh+/h7NzB3zq89wvLgRqOLxvnj/FLjpp
uU70n73Z59ruExWRVOYxkofU2gP2EQhGWlKAH6VM/IMjYBKGs6tlyFwdqCQZUTw6MFxsvQjKYsje
lbaZ8S8n/fb838Zy2ftPQKHS6pNUxYgl86L+PDPoxwejHrsM+Of6eqjTD9sdf3csNXZ5fsyq1COy
EzhZNgl/qz/DIfi9RdZsgq9EZFj3TF2U9WqRDNB4g2H2vVzVGaBJyYXBRhi0/3z8sl6JiC3uh8F3
BZhFDXtShe5pM4qz7FqAHgHl+Asf7A1S6eWCFQZz/lt0Kmd74uV70ht7Zwu29rh2C27CIK8Rv7SA
DTbjU+BJpzzPye2qNhyUMZmyIKdtav1/Z6PdgEO1Rjl8JQg+DwNEYncbAZ6oXj2j7I1i9r8F7eh0
fF039mZhDvUYf3Z9se2akZR2/yaUnP8dSJwNYtutEBW6Rs7AkGNgNSisu1/ELlSzusmdMp240ynJ
ISjwoAs0mkf5KqpSybLHd36zfoUVPdxOLBuMgkV5NhQrevGEUO5WUBeE5frnp0aA4LIwAxkTjf3G
gQE/i1R81kULwQHBdc8V5vO9K2zv/6QaIu9fNKyupSMEfTWFX0Qc23kgqnCNpGhLchxEErncV453
j4WM1EypV7oVSNsA9/soa33OURzX+HdOTRmToaorbTpGbbitJqpdIc1dHGnl8lh8vK/DSdS2L0s8
Wr41iKWq8JV/jeQLRKBIuiUlTmyktftnDHgrG6MUFZynRoJNKH+XujNWq/xgdTcFZMZr6UpyLEFi
2ldkG0vo5T5j9P9mTBqcMvbpTAsY/lniPXsKa4gon6suxHhH/kfZNEQHW8GjPpl0jcwk3Bs3cEyL
tHFkbMlA2giYRt5lPQDDWSOY5E0ZBidvK6DaHcwMAhHQ2nMlFk/yYgFCzzPHeDR2QApSqVWlTEH8
wsDAdo1nDXn21MfDKHPgV2n9ObutaAhtnxbvz6QTgwmmPYwBq8TdnhGT9WUhP1iaVQh1I9pe6E0z
E/jzqAOQMyT9R9lP8Ve+WUuYbxG5uelyuu34wp/QPN0zLOoQrZ1ZZ3IN044/NtCA98D0ulQu8p0p
feN4G5QAo2sxN9CSKxjhvo6FxKHFpfyUx9B9nk7McShg/hV6w1M2NgCaf4+mCIH2yDtebGfRRtXc
WR+phAkwDrb9d8bbn1g5jVbzuYIcTZay6DpXGAwT4atEWQwUcU8Kj7TyM3Q/ielulMbZB86aUwqw
oWq/DAeLfrirI+UvFRUUdUC0B/yG3/FGKOxrLgRPrT7aEmqvax/CtkTp3bAwRNuFpc8uokdS6jDd
zPy9mXwtrsnbdyY037QhaJY7Ume7Qtp4zHHoqwpMIMKNnMuhckOyi90kz8lJItxkR6CdzkxmiFUr
JSog4DFi4p31KG9WImeYj3N77A7O16pvS2u8xOaUY3OZc36Ughkm3M+QkJurK52zxfeh34W9KbMw
navQpNTj7RoEQstIMpT2c8N+ko8xOrVjIBXI17gMTZ7emkMbqpZ1PcfQgCt8iXbPnlQBOAiAm2rT
l0rtRpYZqdA8tAoni0+5/w6qr+7xARZDcUKkiRBE3X3/zeJJxV+P7MabGPdCwIUWJnM6c8mNJIKI
IZB0m7xBw1j4jWj+crqp3RLbiXquhxt3nKTKCPU0Dyl/OtZRqhiwfe2LVcLbniJhkqzwg1t6GcLa
OxrsVOEL3O38nRfiNZw30E09ketoVVU77/wF0PwEeAlLPd5+XDRsS+9oY8SqdV72A28zdcYvsTjo
yRx3zBhpzgmdOck/pE5LMAkqGMq6NbyX7Psnmqj/IoWFtAn8/PMOeu4u18oO09CqqzOJZHVs7dC7
3Ncf+PZ6HzxvB4inO+MPVMzAiUmeQ+4GguPQbwWHh8VXLon29Jgiv8LoRW3QpEr8X98X0xefSWPX
9Tf/NQ0UADcC+XeLPvGLfKr9MHuelYZxihhq8XlV/XONKxg1eQHSjWdp5+tdgxbgFVl2tgrVNCwT
AjW33GbGv9UcKIeyLQPJ+/KHcZiPh/etBaNh4Yy2ArSwywHUJPKjaV14Tg5RL+LxcWdMF0ou9Rnl
NQ80FKZsTdXsAF3YMua32AduQnuEDnOVbzD5AUHlazDxYcp+DTzm450lSh1ZWQx/QNXJZu+Xladv
aPXiXV2yoeW7Lb8cRloxHjT7bRenFFWTAwHsIj1/k3NsoYln70O+tV1DrBXGB9nOKxLHsD4X2RtM
FW0ZZ7zZwNWuxoNrl9VHT4vR0maOfV8ylcozTy+ZXCdXkIQSHTsztiXeWkGgYpsHyARWUr6H1E3I
lR7T7gcRW2PWD6KG+gdgQgCq2u9L/tAcX9J950pw5nDzdNBwRnXAgV+YP4NzLYsK/PBziLXRJJ2l
Y9d8XlPJKJSXPIOb30fjzcN7yHpNtLRiqpYFnyava7wQyzXlzr8hJ2pmdMwrPKu1J0G6BMQ+D/GI
z71grIjruxmd1TSB5Z3j3S/tjZdfvBV/Qgs3DhgCvuzAq/O0t+4geWortHDOd9yrlQZlfevt0RGz
ttsdg3+xRLQEyMlctOQs/63Z7LhHGFQQUD40341wpeCjjn6+euPLgH5DfyxT3liz1QJuq0lfIHfG
FiU2XGDT4FC4wAPwr7K2RnYNeWCpe44XtXAeygGneN8gc4A8eJuoR32E5Blp9c1A4boz9384z4fG
Ood6kNZwDkd0hRlUs4V/eFvWPbbRNopeazudslQlS6d1yZj1DefPFbpyiwl2NElNdYq/vl3GGT1v
Xpo1FhlQz6qQjtlT54zNH7wwa0frY3Qgk/CdkBoi2s/14tJ2EvLZTpuVnPZIJCvgAyLQlq6v9Cu8
76uVOLRZs1xyDB3JCh+V8vvQTpZS/l/PjLGVKYqYv6pwPa7zoXP1KS42L2DluzcLgRJHKkm8Hd9a
eK0oLXI5OFyJ5u2LkWqevVC7Ulofts6rjlsyw4tEV5HZgzSz++tzdW3QcOW4X4c0Jw5zzB0QAdi5
0g2UTSNge50q/0zOelP/h6Wk24l1wA2j2fKwe6mnYBT2Zot2bqEpDbSi50ha4dTqdx0DworNit/C
OSR8waD6fNF69yUjuy9Nj1pGrC3+y829aUGdyBN2PC+K0f27e5XSmMevrYBdVKdPYPggrE04Eg/Y
0ui8GW7ARRMJACmo3GNZN53vgATXPFCLwn6E6bUyKT0+5H3bEuTxMKK18s9cxo3Otf7Ir1Siaoca
eM6M4PbbjTy2XjSpsbmK2CVXOTzWwPoUkgXwvca0Kaw1F6ydcVQ+6HvuXpPzV6uGoUgMaNrenjqq
zZU3I3z8/eDPLfw2bG60ZYETPN/zuo40i3+dnmVDHldpczSpBynPziHGB3lbsZ+6QjhBkcP55rOp
c575cHTUtjcdC5YTMoIMpP8U2Iz2luaqGdRtCGjgqCP7HYFMzx21tlilHFWXzdZiryI3v15jHfBa
P/wm8Um9Qkcv3llCdBIR1AgbUrgFCUM08Khdbb8yx6/Rctt+N8AqRYNsaZtY2N1Pu+BlCZyaHKD3
9Pf4qULg8TGrUUVSKtHKY2UoHgNum1KZFSMyDilZ1VyjqUAOAkmNKp6TQpTQg7CLJf9JnBlk7EGk
4qhnaHMKhbJ8jbnnhXcFnhGJfuWMpyo3OQPYdIHLa46iYYVec20sj0ru7d6cogJBC7diFGgWkbD+
PcoTtm2Lw8rG9NHB82KeZ9/+aqRuggkoKp8RWe700FH9c27yTUm6F2nCCvB8ktot1dHEsU76Ou5/
PBGq1YwOqbxoccOKdF27fmJi2Cut2N/0JsX/YSXdZ5hFbKbwhfgJGpGQTMWyVu3EzH1HRii2b40j
pTYFSwJWEMOHG7VsWqAvFb/NJ5M6eyCa/ByzBbfkqJbphLAeuOJ/esLkf4rUxLiEWL1Duvl8I60c
j0s+17+3c8PvS6ipkAV/32U/4wsEL9VSBP6lNpiqfwn+yRBK+RNse33rb7w6upRHHxhhQTIjv+Kl
xJUx5OnckLyGqjWn6r03PPxbAEFhpJlb3TJuKqyXvDEURepsHDu1NNMC5TZiUklyimJ4vrpwfN6I
0YS5Yu0n16U+wpYtsk2i7N7jP/QCaYu4gmMvdVFqndQJR+CDIhxZXZ9/cqv4+1H2ipgc4mC3vEBx
ROFe1jVasITp2EWIjymSNeYfHKUrpQJ0tpB8vyUJnDlOKBcn04VeZlhWrCnVYVHhUtCL7otJ+hOZ
O380EXK7qd7qw7KjWGGAnHKX7MgzTYBMdq6ZmhsLKZ6ER9CR9jWNW8+SJ3RXAVQf+S+th6xZjeM9
48BxBwrjIp3d/VXf78gFnzsFo19e7d2+RGkvtAj7kB/xAqO6fRWTiGZugCJj0jOom0KfEHku8YxA
Ta0ovBDMQ1R4OTvx94NZSrHiptRWFowMspatHLRMiN1O9bXCtYaljf1aejDB+BTcOM11qhNTa2NG
bqiMLw+98q1ORajlHpX0JbA/NLvKZyoIL9FHmDXFZp3gG6WYd2JGpNEIroQfq1grSt5yGPxKglaI
XqHCaTGtlkPxJK/zKREOnRPF54vTkFTctEI2vrrYvDuJhwrva5bu7gvwVm+FXWgckQDO26ZiSEHE
UJYr1BG6l1nGyAJQt8HKK+gs4376YdBUKKX8GAiPIO4r94O6haI7hTRJgU/aW4kQuB+abmRdlaAX
9b0lWmGz9jdJjssCOleYC9msS0reKdSobNvKnFcniqdUJZ9+ryo68FJC3qszgQ2p3Tr0ddZfLV0M
RvlNNS5fyELH0D/u1YrDmWyehoNkc6RVVQ75096TCh0VUqPJeNDS1Q3Y7Q3+Ecuv5wg2v6x7KLiy
ykGaXPcgPKkxvd+XnHIJU8x01FDCiAGeCuJJlCOxxTqNTIoRAcfviJIzdzK+mVDBZDhcmOBPxsmj
iQEjng9rg/gmKvfnEh4s43Nv8rYtx9xFn1soSFmeNFAgNouZip8pj4uarYiBBZHjMHQcJftkH0J3
Ru4VJr07Hxlf8a8sk6FQHqude3BnqZFIqfMdUKkFMrsjxc6zim6JWmmY9tglIeMXT0xlIQSnpKSo
ifZiKJQCnpcBi6QWpb8Ru3Nc27YyNU1krp4ZFR9winWoSqHV/drLfvpukAT1O7P51NtsuVifWDTq
Zasf6G3Ba/g7bIYVHzsqgFDfXP2dyFFWIj41CSeEyyICZiYZV+Won2gvda7XN3uq5OxAiWI9WZHw
FX+7YdtGizzJyf0NqEFlA9w/qsDZNaoKfBpIOuCGyDLoe85krsTR9TEkAsMHHwQHL0QwYsOBEH3i
3dgIZG9Bm9QV/ebKeMoOeWioQCW2n28GynyYxSl9RM9P0g+eb61qlcuzim+fjtYjTxOc8ruJhhGI
yWrgSf1NtXUhg2ZQ1ZQjg8G7zcXYCyxHke9EQkVqhtDCBKBBM+T9jX1tcP5fwCsxONA84V+2zMJI
7N2FQ9UcTsdIvlSeC+VZnP6hsg4VdpMxzUYZmaumAvDp1XQckGBeGsbxfyxZEvU9x9cdjVz85w1e
O/PkcIJ7VKd8XCAIgHH+ZqNGbVaI9LyjC1ruSTKhv+vt8LnxnDflIhiTDRqXyqYFe2dYQf6ABpPW
E+j7vNdSrBjm8lCaAf6JvvyyZjbsum2mVbQK89dfiOyjSCiFLEhFzRBaTmB1ZPu4KFPIOisPRGWs
wZ+ob4FyICKG2RA7auNroqJUp3EMt+/xhWYymbWoak521ooKmDGMyBxuH4QP7pe+EY3/P0wudiRm
WXOAlxHYAQXviYapo1sHE0BdfK3994K8+PPXt75a1TNUan/bbhWigZVhO4NwfMW9tCgAkRARa7ot
+W84wVy1tufjo52KEKUiUJFAdAGTuUdRRwkVBEhoN2UeqQr20FRzy+bv8hC0htfa78OSNXZkeB6G
yFHflCckkHn73XrefGLWaoWiSIxp4hu/9y3cAG6LpRf1HdUf+FewXXihYxlFIgPWfSymvSgYv95o
TvXRT+DT5Cg3IkFXcvZ81RFuOWJT6ws2AX5AjZvUmU4ScfwOT8z9S1a/vlTpn3GlsKMY6xGPCxr8
fX2xwxR0Ub74NtIZovUqC/fPv+DOJJ6xZC6j9uHO/Cz6skK1RjygW74PyorRba0YUHoP0oHdBcV+
SOo8o8tIqXbYecBzoMZSeeP9KgC3TIEmhBN8tFAGIfPgKln1ytTF6CKvuumquP//LtwXSp/CfK7p
tm9PCqLxdVUI789ID3zQqSBZMqM3Mps76NqUAE7SAgEDZyEBtq0yXyPDyx7u6ISNBpM3HbNc49rL
jri33SAOipbx4IU42ED8PIx6ZT6WQRN0RTb1CPcIcaxIC9L0uKeAWbrtY73A1XP7hAUf0FjXmn/y
Wr7+Kvf0lgrnZCpMkMJe2FKvqTyixhl3Z8Rv5brqFlGZiKYsJs0Yvj/gujBUFrtXuIgaLJR58AtN
Q5DlTOU0Ic7MnSzC7e96Z44fEr9C7Hz5kbVb89o02ZV8U7zmbsIrNofP0NaQhzFX0tYDX+I6PUZD
WWlGaZBxMxiOkKNpOm2SjDaiJ9vdOu2hN5wUSvtidHJddaJdQcaqcarjDhj0DDBB3mVzrKDnhhRG
TFp8awKrU4saesUqTPrrGWBQqlM1i9c5yTtleXo4qxhGW0nWCX4yGOFFKpSpnsbNJmSI0BoBUjh+
fprUnx9qnNfEntjmrbF4xCtuXVWW9riq6OrZWMcb2agTVwhiBb0gGXvLPEjd53Ks3g3bF/756rwI
XLthaO2ciF20ALqpf0+MS+Z5kNHH/AFhqclPDlZhQs/zcIyS4ogq46Y9jIDH+xyCijV/QhxYaMjm
G10xWrzeLyP6lpiQ6X7RZ/Z8ZS9RXNz5kEBOCHFk3Gmc3kQr63+rEK1yYhyCOrjdd42MjCYRQNqu
VLeGRj4KRjytR9eIBVV8kPsMl+bbLZhborioHoPXfabCv+BExP1aeeIi+spCFSnIEYp5T9K6qkUO
iLNh15epkwumqrF0utHf5Htemdq6BajGJlD15l0nEzFyOIKrIvH3h4ApY7Np2YEj9Gtj2wo9P/T7
mO63O+cxe7cDuyA1cUCTUxueBJrkMPrmBu+TKXZsJwyq4axUryBJ5i61wuGh2DyAZB0z6Mb9myll
N7StSNEe7jcgw8HgwaLuHhnT7QfdeZHWug/u+/WBxkNQ/oEiMieKh0cHnPhUROnLm9MRfgkgD6IV
bTtI+RP/l6XdNx0amN33CH5sO8fwLk0poZsMMeSaQyzdNdF7ldDOHr79WESJroSUs+FwMgUVg4eD
3pyssezD1DUUbD1P4WH4INU/SNmQCh074dXSIUaC2THDm423ZUWMyn2kmIipCf2iqijjNOn/viYd
RLpOxEumfLeL59fR2um284RW95R6D/z0cTuCTdBbmkPL+k+zZcgpWOBo4MXWIEll9G+/5rbTM4eQ
WEVb33RDb70ZMCqFDFwFXAq91DQQwXGibfVgxtx6GABhb1W7QeW8jibOtDuIBU+Dyll6ji1B3yGR
FnYZDYJl491OP0pvqxvU1qF1ekAMjPFEd0Z2Cwpw1hmJPosxLT/CGLbQu5ptL0cX+/oVaSx+Js8E
LL92RbTyzjcok19cC8qIy9dc24Wg+cycBFwDzFwQ0MpdEo+oGP7EaJdvCpUSs6m04ZG72ydiXvVK
KRrzF3aV2+GCwzX8J2dZu3jGlkEF7Co+9sUFGevr2LQRFnvBufl7MqDMjPctDs1y/pK/5tFCm8FI
daquzwlnSuYcgmtj1GHUFcW4isuS9bvFPbOhyo9lurh6uj6rTc22iu61GO8D55MwL6WpPkfjp31b
qWgr6QVEOWxbk2JLqxPoBOuzeeAxavk6gDeq2WC1PyvRJTTnWvpn8cyol+3RXsDiXoklvQt/KMqn
HEZ2f5LWhXlwPXsMZ0ZDNyUGwuqwSoGEaOUfqXcLI5csyOuCygeSi+kTjmkDvC8HEenMmy65lDCp
dp7nJbXsm2Jp1ZhWMPPCguxBZ4WqhWmbYJJZpP4UQzjS0L9+llFdjoUqacgW+KknMqOpOWNWICD+
8M9oElrE1bxlHDLdecVyH6eUIwwAriTSf9FtfcGngPtLTTlokjw8zyn0UTxB/vz23CLwTpc4b+2v
WFUa085iyhEilrlYCHp2m0oGMMBAVrO7tAFcwWA81wBObNPzkce8L+FrXliHgSHLRjKR9ZNhVBwZ
zVTFf2vqCeXz21Ic/MuPXTI4qzpFT8/g8dU+eEQJMhhNUkatnaGBJzaKarjg9Lmv4Rsd61Hgb3qb
rWMta+FrBaZkqJsfqqFxjHLzfwmt+Z3SVZBfpIn7bEnATLAbDgdZWrwOOCDBTK1v0VSmemx9BkH7
TlJDoHJ01uj08BHGZMC+6e6+oDFC1H7Kk4RNNpkjnh4EjAZ2fUqaI/DYF05ZotKDqd2eH8hoSIMt
FsU7qH8N1q4//GUmuAlUScTLDdjjTC+iff5G+lbVGoD4MuadbeUOPKnNoZBJcdDUdstAEEtHvQin
AWXYmCPUCKAXVm36ho5Y7/WE+HOgIjakFxccbBxs+4ZFwzivzA5OvjFijSxHAjBz1vz43EZj1PQB
X5f0yAixdzkEQ69UG9PIED/nOnk7rG/iqimARBXvdnPOliG+t8SBvJkrKOQ9PvjjuOEDewqOEd2p
ZFE0PfPRZDbjnjeA4xopIs9rDAT/yWQsyfn1teRvC6HWQj8BmCDem/t4zwD6+hcl4pUfGESIyy2m
PvrPYvTkm5pz2umEkN6nfM9Q7BFkz4GVlMadq8QAn0wMCxN07dqRLBpevuar9fvPBTh1xiVxnmIj
LiA3xUCkI7A3rDZhjFRb5+i3In1wq+Bd3e6nYGhDYh4vvVW5XmlaZq7IAH/vAPWipdN7Cd6sIcYO
gT7mlhXcwRUL7QM7Fyxa1cp67macGwzAgZPTI54HY7P1+a5/DUMB3vLC8HuHwtS5+26y/jO524nd
wj/FaxKDVZrWSMAZFRcIDf9HZPW1WOOvRnO71IySr5fD75k/n5tPr7kaEM281Bz86bwf7oD8nU8c
FXMLMH/hltzbgDnGVBRwzCr4S972M9R3MXCIn92/s4PEopciosNuAjyctMKY1MDb34P5tZVsDbPL
6lrYDN4tiy5SsqKJeWSAcdTL1mMP1V3EmO2RwmF8D4y52O1S7STfU98vRGfNcc/65gxmHFLiYekM
fR81Fz7RQChHYf+GdZDuz3OyCgWNPZvB/bX6L+djkz1gvXckkR8CHcqc6rFKPz58JTL5ioBqK54W
7x4IKm/1nXp2QPdxGXYr/s0hBbHjcI7I5CpKHE1gOshU/ee1LB2HVqR5mnFIiizs7amjwoPeekox
PMXhME6neAdxJi/gfK4dA80MxaSA+ObUEZMFnS5CR2nWIRupcGkDzGaEy59Q6ep3SOPNhXSf/iMO
8RHP/QC9v5Hlw04j3A5Sf9f+OzPx0gU5JH19EgYTpt55Oz1avl32SR+RsQa5Z1rFrIsYGyg915Xx
ANwAD2VbiHKqiNCsHHKazWysneKG6svzTXnVWElfMT4lMXlns/sIsMGYlMe5k2dSQp5lMdnvL25O
dwhyez3VPg5ts8yjoIwi6BTKN4AIyTRWyMPJDOb12bmWLIZAZI2xiaHTazLJgicV0jtKNHqx8etP
FVBJvSQeGnHbRg64oMgs5O9Sre48JhzR0qdDKdqd3qaQaZRnZKqSnQ9tuSGWLxt6GukEvXo+pObj
K8KXPm2w2D/T4g1O7kI0YtpChimqGyq5xfWEBFnEljRR425cKQC988SHd26qRx8dYE+MfZVyjZbX
/MyatU9lEwktUbn2Zu9S+izemd3105J5H2T/h6XDf641eakR0Zj18Y4gEkpWNzCkb6GL2j2kxF9p
6OOMO0+MJzVmZ8578lSbauTx7cgrvcloNuoV3enMznWSSHlugmFy4v63XcyY4E+64TXHXxUofUBX
GnlgodwBkTOGWYwDitG+8Xr73uXbOk9B7xNNLolntntHLXDLk2PnNv7H8svwK8osiNocKAYZce4W
J1d80klnGp0Io3pSxOcy24m7h1vQM3BpucFi+SMCamEJgnJETQPAlL7Mzyq7EjbJIM/g3g/STdae
DNsXRa8m278lrFvK7Fv0SujQCxDZZf84TN97GncH9Il80pZlFn5V1uMcJbjxACaB+PGNXgbFnukT
QtfFFGXGKWAHZkx5EKYSGzbLPPVGB2rUQrdyeyc9BgQ/EFBV96xJXduCIbCyt7XnqSUVkkSbqqCN
Qxh0nRmpvtSvPe+xfxxSRxVyCNl0fZ/Ih7NKQL9G5jYeAHLVyxVP6yM2ZBHyYkHOlCu3VZxBT/BL
DnO4a/qlPLm8L9uIN7NXLV3Zpsx4MVEyPn6Tv6YAKYotzmSUBZvBT7R8Lq9KFYQTsMn92oLk1tPr
j61nAIL92U30XlBt0SDcKThjWCfYsVdxwd/C+PLNP8HB1ApMsFImm9zZLHgacg7LIL8UGuAP2IYp
WD99nGwiuyMJwZHpbJTVF73mgz6NkiHF9TxPXTzWh31ZIDknlNv6pUN36/3V6I1fRQJbjvxXd3kB
8BilhEge51LF/80o6PbpIIeb/6N8UEkTF29ooEMzygBrUGDbn19/XRMN1ndugyecLSwIAMHsO1DW
Oo6A1r2zLNKZcOuiqSkOAqjNxHEjfEns7esduM9I7qfQ0a3k6emkCycfaXTq3tRvn4lMR07uHwbG
BllZxAEpPF8lFAf9hJkbujUfsXMd22XrWdB1wEoVSbBE6J+OPTt2Ax647OOlt+Lb8HR4nt6HB0ph
dhXP+tMITD7VhDGgiDrn/JJWnsMRdQ6kcY+UuVLzvA9u1uA+MU4+pSppXCuJcQCyol02YVbdasLT
t4bhIX1Rz0wqecL/2E4k31Zq5TnfD3+Gy5ERTqvYYwcuejFYf1+xOtPE/ebY4ceBfija1LT5PbNU
GCq14oVNjVFVUi8AtnF652Jk1ED3lNiDx1ZxYNCEswCDD0iD8fGhu4R3NhIzKOaoEVWcVkFjukfp
/N3C294Ya+9xuTxSn0T+tlTfS6MF6hHsCEraMQL/1pbQ03fDbyuwAhKp88VW8RDHqM3uqStEpEMc
v9UYwl4dSe9ZGMXR5pkZW1yxtflsfl4PaVgMNfI0Ar6BGRKRGCjbd6ngCmNCdKdJ4KRnu9QBpuuD
u/eOjKvIW71a/8/wZDq7Z8lcwh7xJgwOBr3QpMBwrGtDotaXqSl79aVq9nNZAF/C4HJo2u3b9pnc
vK0ETh6lLaze6fF+iD8iZgaCDkY25rjtFz6n3M/jfmCj8DV1VbcK01MZH1kVnuZs3tOTeCylFN+N
RzHeAJGOMtleFNpdpuJiaolbPZtz31xsrENONmEiLq6sp9Jsyq4Qf991Y2ZVF8+Qi6LRor25yiF2
oBHmYUee2ChCGv99/2UAMDR05ImEOxzxQdJY2YfI8W+5z8RV9Ru/CiB4yxQwFCeAsAJE4SmTFoTt
xPLEJuAvcKBfkWB77j/qmg4xor4oEUByTSxgHLJl1tl6QuCFH2zvEGbFPYRMNOHvCF5RlgW2jEzI
iSqKsMWnw0dfsaIvagPjykBqd4ThJ5n4GKVofIQA1p+fztHdU8e4pme3sVaJ7dhcEvjSUNksFK1L
zikAg8NQeMlylJPb+mcHDf+BNCcM88TF6XfO1XyMfBTyrSRpZxKj9NchaFsx/45yQxi+8JhqRMoR
PAHxXdZZCTPATIh0yN3oUL3jiIwBF1CASAi13dZC1CvW2mvHpT6WkD+XFJAikgcB8Smjs2lVYaL1
LXMGqhvr6dwNYCwCDxs0lH7s9EHfDky8MXtiuEXGKCiERG7mK6cCQeCzJ4dVKj2Q9xyM3bCw02iS
M/J5zTR/y9KesMNeqDJ0jrjIZqTTz5/cEx9zZ7D9JeYnzx0Ndnef44xIc2yPe2adRCgFyDU3eEIN
5Cb4dMBMEHC1AghcJr07bCvwgAdKSyjl1aeAkrDAVFR5KfNoVq1PSiDjHzBsxxMHsRID62KpfA+T
vvSp9Yply7OmUX5Jlcl8QHiQRoDBhhc44QK02mJVU54Mpu5VkIo5AzlNMRPJKG+FQ5lzC4uHWEXr
sToxE4HQA/3yt/vlYmAwnqYeeKCRuQY5DKHpOXzOQGymZq/PrYfmJMwNxd6Q6G76mJrZrNSJp9NY
ly9WqaDizJIZA/oFcojSaN4cpHLpp0LXO9sEGaeFeF1jIFXZIsMYk6nDqdlOf5aWK+ystGOvyHaP
CAqcw2uMFtxgleOxSVhpIKznPhhzT+GqfLhOoPE8AnCqkRTguc+8fCcopw0b3wFIDDiL5FjfjkZW
+cmvZ04YJT7zGKvOb3uCQ0gQZd8Fydiwug+1QrGPCQupnWuV/PZmA/JE2m/tz65hFs5l1vsaPR7f
/t/v6NYqtLNakwXPAI/O0HEx15eNbCthkVQVJjCNwyb/Nz0sJkoAZo7EELBmILd1YLjuSSu87uoS
Fzfbvzjp8TcEhvpA96xJX8lU0zJvE8aKz+wZbbK83PBq+M80og8M43QOPEnq+vrDooVTHkZ/N4oe
p2968mUF+LaMQvjrR5o5sPQe0nEkkYPvB9n6sxvC4Z01xEAjMhDmhm7pthTu723eKjiqbVMkZflx
GM9wgxolirrwR3kWk69yyDzZvb3PPCuGSfyLP0zX89+GTAROELsYCtKk4Eyur4DvioGmuRj5t0wt
+c5J4Pvdu39J9oNCnlf/H6/r1+rV2xSCIpNA9QyQSUhkwedFuj2aASNshCUn3C9yPwycHKvHG/NC
CEO0ljx2roWqT/P6tdMdcZaPcOyxOYoTqNiJdQgdl4QwZux8H8e95CRyfrlkMtOrgTd3Cuk4jvZ7
De9Bq/q0JaKrZU75Odl2WmyumlZJgDmlXU0dxgdv7OjnoX5kW9HcXOcF4TLiXCsvb3HDGvYFUSAL
E3mdrgMkpKjn0NjnDGawmg40jm8sHhAqzAAbNZysCPjR0t9fI7zClFNBmQ1UQhtdYsxl8tAi7GXv
JIatkRNBT2T+PDgeSpVusRk1U1pTBTGwwEaC4Lg4qtTIrckRfMenzP5jLfQlrYOn9TB1Qg3CjeRb
14E/8Hb8H69tb4oI1lIBm4AtL/R26NhnGt9OiXfXuWrs2H65CTvIH7smeLYplH5PjSAL/oK0W7Gd
zQI6zZ6IdHgMsjx4cLJsWgaXBlbmDWtPJFx5lXzJQCrJK04dA8Wf+jufxZLPqyIwhAb6UX5UkxQh
wJoU89Q3mF1kwLnBkL4yp7O2KaV8dfxiDJlyK41S/Ec5/fMN0175FygckOzDDpJMrMBibURpihGo
9XG0CkPeqNy/0by6zyY+JDYviJt8SfN6hmKYvnY7wy+dTaRGbE/TK0K6BSZxGBcr/FZCXl84Kzh6
eLCWcM7Rv4iFmZelqe73bSGT7OMMQUMxnVidsWnAC0LxL4EnGJHoZfQFQuqKzqdFPpQodikgm+N0
d0BzaA2oVwTkaUterLeAyqUTJ+CgVtExwBLk/bUe7mos4VDgjVdHqQ/fKZ7grcwVZPXg7NKKmK48
ZQpRwbL1aUnsmRuprVEPNgKft7Lv1GzUxmC3WOWRsYqKcV68/C/Ij7RsGdFkUDtABtx4ExwxF8F7
wiqy+lLZXWCtNYLy3jOf/TpCXxajEsFuCB9cH34QhnEawdwbwO2PnkbYhHgU/Umj3PY1OIMi/PlH
2IwYnTXJaaJEZvX+dsNbSOqAeNe8/LAPhqT0dpRNMtq/2paWvu7trAzCDIVVsMW6A6ga0NRUkoHE
kHUgmx9oSq2OXx8pfqqRbsuCwcaWSaQpqcT6irEMpXtfeTddfOUabV12Wboy7un5A44VppqUe4gC
SSL+sEHgnYHBVawIrysYc+1s8JMD8mh7ypG7Dayim3mrsi5nMiXxYA6hZSelLQYSFUBVNAukbjna
ZAF3JYfeGPz2OMNVN34PN5pGfXflUoMNCJRYIEof4LsV5toPvU3it0+5X2jLIWhIuvT28qJOEC83
YhO1dmrTfUfeQwAFjpZkYzrNVtY0ROUfOtXhcVoD1qvCaljrKswo5ZAfQbZhBXez72db5veuTI4p
pyugDLCS9N7BMm2ji59frL71N/WOfjCVOXf1hI4rdXbFbIyx6LWemUUUjLdZyzigYn+DGRUii0G6
xK1kKthZolqDEmF0VO4Wiq/XXtdQ2CazftiHYjrFuwWmS+XwnVEuvOnAwB7V/h1cLSqs4PyUHibU
PgLZI4dxSGq1lkaw//2Ly/Rnkl8h3IDJia6k+LRFnhL7PylI80H62gGbPA1M0MUj7qHr4rhf+OoK
5jZupPmyBHvZGq2e/Q5DtewMX0lht75wTYj91Tg18drfinUSc/FGh2RSKCE4m3n3lLNqqlt/ho1p
bu++Y5K7g/4axyoDFMtzxnaOUNSBTClN3WSZFuDX9WNgz0iYTFBN+9cyxfMLvWp8yWQFcHb8mX7T
uhOyEChbsarQhwfpcLeO9ZyXJaxmKyrB3b2pLYaYr/Clbtvs1VayJ/O2Olm+6xFny+0VzojsK9jW
3GvwYFW5pe7sisScuQ0cJYq5vryYCY63jjLZEdiKelE7Cz2xZv3os/TIkdyiEqtFS8aWPk0fVh63
dvwF8zVsrdOGHvCDOnqGXbP1D33W+hcDjmNgCJX9k+xdPK5cYiVogi9SJlO1AVFysDQhgUSL7uho
ye0uNd6EQq/sb0ARxr+Uf6RYxhD0ijX5nvCWL9ApNddjCq+MknIWWDF7qajnefv5ueMFd12godhO
AqYEbGMgzAiEEXQibu/L4v96gAB1uKJcioa/yG/lMOJtF3MvzLsRYDq6/ed0UYjGiCzOJEibV1j3
+6FtShpi2dZkfSsaBx5xGU/7h8Rq0x3SRsG2UYIAlMroJo6168Z3p8Lkrg3wxLE1yYfqYewNUVmn
/XWRYPfcs7gt5nHK1Kl5Mwqz4YAFsSqzDKG8VKwzpEVUW3Mwtr1JBFFajrSKKUbHJisSIgyhrIdL
yMevs6FO8mlYw6MWBJfVV0i/ALwvmXFjjZjTbxpSbO6631e3xYpuAmx1u0GNNt4ZnMe7w+USB2uM
o9dN6z1YXNUdN9GPKBxQxIt4DGJ+cUIBfVhd48HxIwv3qHb1op7tqupcTto3H20B5U7Ybi04NGY3
DFFB5jeXM3ISzmo9gbvedS0/hIz/+4j/IuAhnGKYLVHbB+5PSDzMr1Yz7FpEfwTHleU05vez4Ihg
gJPpfa10ipzJ9sfQdUvheoD1UL5rg0RQFyIR8WwTg9qEufXD6/qmHbaHfjc1aIrNiCjfntUAsWSC
tvQJW3OGVXU6ue249Cl0r73hdnsUMfrSPnnSlEehomfahA4luJLshzymn9ebwYs1e7PTwpMNNKR2
Enlxh0q4aiaU0/eWtzIFRoW5icsB/5donxOJ3lXRWMRURt11YSWn8iYRfh0+ijPWC0SO3RNH9zRZ
nF2KronAxvZMh7+RJSAszmipyBcDVo1T2y4IY4tOouXMdquy+LkWpyxwCr6wKUUTD3LgRgRzBB69
s72k9sc2ud+/uiE1mxMmMapDX7kJkQ9EVTTDDz5Aqo61C1IYNsVZctqmvs8VLvRNAkEP9oeZJDpE
dFWY0xc1vzXDZrDTyNTITmfu7U57SqxOctcj8TilOq3tdT9MN6nJiJAclsKsUQg6gXdeU8ZpdEkm
j4Hj0+jBaP1/susgw3vgI0TmkNFoW1XX0HFDDiYe4tKjqM2ciodm7fU084CxjRStMJQL1P4o+HTo
XI0wOAPZLWe0Y+Q50Te44/UB+W7tjNYr0McBZyHWB7lWMqzIbq7VlPG8qfLUl4WXF3nAHupUZ1zW
2t9HcyLaTOMK+t4JLN03m7Tq+/LSurV7FQ2gPUNwVlLNcxUQjrpg842Ztq/Y+59L9nkTIhWl6Oxn
8lRf9Z/JvXGKUMNeZqTGHtfkXL8W2Xfm2cqO+iOhk+/CKjyYjNX0U2WaR2sCvUDV9QZtiRVJ1mAM
IiVNg86cKcTeCno9Rts9zUIeBM8KL/yzZx4kRwDDG69Teawx9pJ9jttZzm1FCbjFf+xVNWLJp4PC
7MrUFSSgsss6ZG0g7Z3O3dGd5+kTC21H5UYlhgOoEnd+gt1ZW/EMUHVfkN21mZTgsMCNBEDihquf
yF2E544r4czpvKaHZJ/mL6cLXpeILw55SkqTPaK7hA9CdFC4PRHeCKovc1Y8QtcCylQhDIfr1ODE
09WozqmaVIOSTF1Pj67Ni5DJtegPlcQ+QWrpFFVDLBF2yhXzvjDgVx4rtoUvOIDiwq0WhjjQBO0E
xEEr+3j/Uy+VqMC4C3sJw7yb+ON1oIaJ7UVDfLXnquZYejoOmslsO6odEQufJDH9UGtAVMmF16Ru
RIgOk0JfvM7RIXlQl4Xle6WPPs+R0AuwY72JoTELVlX8C25rbCMNp6rkR5P5untpWRaXH+3I4XCV
gW1q/V6fUvr2e4a4jQjMUPJFbbNKalZRgPCr8Sz876VRM/APt0hjNdkP++cZngY7OOKRaHn/I4Hl
qprzLLg/p+DHw2CLxjpekBYpShyiI1XQlMbCR1w3IvmZbqXQkJWUqUU0RxeeqMaOpmJw85C3wBOT
ahBkxcgc6Xx8/9xHmqmZj7opxs4csZjtR9IfgjCWouBwtY+w8UYHKUAx9G4eilzdkOG0bM2LSzbk
x2j5ob3n5pNN3pL1DObX1jhgJSl/n8al4TGpwyA/xK4rU83p8VY8rRqSu79c330tjIkROM6sZtUP
AAHTnHVeW+7+6I7KCnss+y363E5ubia/oQFf3fEXwoxlO/HE/ZksLVEAS02haG65pXlRH4uUwX+M
Fh9TUJQ9PH9wFX8i7pGzyTgf71xf33bXkgB312Xr/VMp28wnNr8HcuTS7BAjPbgheX3U7SllNOYj
Odg1kFXmYLA+L/9YeRoWlqFznSUPoCoIbEZrMznhX5JMbCmx0u2z4vQQaLSJaBCEUOcMWB72HZ58
uRmtYmzU9KreozEWBrhwyvJZqsbsqLbQvdBu5nqp+GqAPUpLMQ5TqCTtEQzhLGXbjIN+kGgsPL5S
yGeum+Yd59R3v0H7+ygwZPONtRP5yqnTij0Qq/cAHrTFQyDdfStpBJUopVMdaMwYtzLfonTLYVYB
h1X3/kndI1tKUCo5CxZNqdQK/yhHQVT1H8+etqUVIlFGrRJyjmL3mmNIBhYQ8CteGu2+rWNX5Vrh
zohUukN1PNaqKVMTXFy4P5SXZ5Evv8eYBQhD8h3A/QyDPPQjWIzOfHvyf52ckgnjOtQzZLeQJCaK
5rItZMSWZlg9CbwGd/3TsdmB9xoFpfPUYdOh+C93O9yBGp659UTPor0J8IEh3/oVUoczXlro3AM5
+t1yg8TwaGwWDzOgrvSFk1yEM0WMsK66p8HrVDXi/LVqCgwP6nIVj+T+23eQ0CkdmWgkkzahgxmS
Z9k0q8lVtv9KH379gDdt31OX+bbRuYwRguYVZepwZVixDCzNf8Rh1AsHcUrG35ZvqORhE7f+fC7Q
QOWqEn/H3EXroifxVOfljiR1Mw2Lx2D/rxY8smdqFUih6JY3UZx8xVwarEmIRTW71yZI03c3HYDM
WmO79J1+QC5uKuT5j//WojrOUzJuK1k9VK1c2M/zihN5wmCInxJUTp1PAdZy8ogSU+OeAsPuXmp4
puEzhqBqi3eQ9Z7BhZisCysJ2YVf5p/8BvXcFhwpQVEv/guHT7fH9DQVCNDI8IUt1+aVphsfo2A/
kdZ5rcFfu6tTP3XYak11h3mSp0xR+Sjbzzp8uTEm4VI6DD1wTZ+JRhEAgDqzG4UKqmgCPCoXTZGO
ucYrnAEKBQSM3H0w50arRzRXeFrehQpYQVdEgQzo8cmB4iVqRrAkj0aonTOljZpSNPzoDWkhOYvM
7V4DqHYMtmBeKxbA+bBQaqfaxO89ari+E7h4fNmhT6zEPlrZWNqxz+vEqu0hai5hkmfMsJy9zjmP
Saxm3DLwYTJheNNUwGxjEqlRWj7jvJXVAislSxaSflt1LMvfH6VRzMXTjIa8G8FPHVFxcrC/0Q/j
bz45TGKwuCyK4rlk4hcZGEobyGy9kp//4Y5LWJDG7aKGY+zlCdoxpZP05tGjjK5jGjd8l3fMrM5X
rBCJ64CwY7OJD3mWA+OfrrB6AmY54rQfqn0dTE1Ki6F+Jl94aAP5UIZ+1GymOqOZJ7lHYzX+X9OH
QIbs+9kcD0nuTOkM1i93p8L2GIaP+5qTJ3MDhQcKrXV2U8rHLnny1t/+AENy7Sr9wvHc+otoYL7A
wuLoMVmf4dGLRfij/II4VBpGct0vKOrHjzP93P7Z4XiUOzVBwmVg0X8n35fr4/47MDxJ5XjgQLkO
v4zOxAVr6IANGfnPTK9MhrULqRbL+hVSXJVS5dv+t9dpT8t8fAYT2/9okNcuVThVNqVpjNza+wQm
jB2b5zEUuXOERZ4GJ9h/4F1z2YZ9iHOTD07AKFsXWMGiyLmjx7c+ilaorhTCY4YPfy3km8U4T+DI
JOK+uFOr0nv0efkaO9LY/PNlTpxiRFkolol+aHkLJf6WcZr+jSk1v7J6YrqP5M+Zmy8ocoLdVWfn
WEDfX98Oe6o9ckCC8spuTif0cvAe375uZm84a+JDv1Sl6dEpNCkfRuziuwsQHyYJ7Y14Gf3J9YAR
1cIEY5rz1HMg6+2eOiMsV1zjOAWg+wyf8PbiXGsGeht4UCEH+DkIL+pJ/KCjt0Or+mOD7oDNihoA
Pw22HKpPk8h3IEF+3Pg4kmZ3u7OTqL3Fqzvl+OBdrZP7CpfHtzcg35rS2vxLkyv7cKKwK1cEuNmN
9Ng+BJR2RdOTC4vM9EDObA6jD+SAHHyqa0mtE62aLOPG235cGhinF55ULBlNSwE8+lPJsEJKEqre
t194Nrh8RQYsTWaNHhkhyxvUvd+72T4Q8M+L7U4YDdXwXDni0ITEql3GLi/G4FwIIYBLMvbbhuar
zc6f0padnbzCOvxQUxLrOJqhoG1EyBmGeS+kJATaEt150HNEZv4cD2v3oN3rpx/6INcqEtdrH4LS
97zsWxp4tEb3uwhmXGp2/6t2ploY79WBZk4NYuUTGrJzBc80WeBQZIHnBwWKi3ZB/WB+15nODDpD
ELvGic8CnJnu45TjI3rEazJkmHAHBDaU47RI564T/UftCSfnhaOdYHXYf0hdGkQxFa3KaPsTU+pK
0wXHE36R8fD+awOVfKRKzaMiOuyWkG4JDbHe6zAOKVjoE5T6od5aztsuouIQSncpV4AXCevBHe4g
ZQKQgEmWXC6Rgpbc9UGy8CzOKWPjm/U4rU1VobM5/UUKGy/mcmq7pBmx9SXurI5Oj6GsT9busDy9
aXdgK92ONgdJYVVyID0xH0jF8n0nU2bQfnZMVz7MKtWPUcZgDKlbP4SUnHMd+K9oARQ1fzJeNpD+
AN1nbMXfj5IGMJd/BvUvxvOa/Zvla9Gfuk5a9/cozDqqCFZ6S62SDi/ymJPYIwwdpk5AaCqH0ChV
kwYuNwJhQ7E6Tfc/luvTeXComxOwFR8szVFLAaxqB8TsHh2oWm9EfQSzOKg04+DpJ5UL7jkFzi0U
skpPMluO3NlZC9Ovrc8/V4OdugoLYIgcv9N9xiYe2mEdu08f8KycYIvyo3KgTG+W+EMLf1gfaskx
GVcpGluj9a+pxAsUFx/eUR7YdPvAKXOBSgYpUIGkl3aDMKbmYHHQsR51DH1q0V6Xov+OSAvgBKa8
js1vqbKXr96pb00AUeoLKpMIZn5RIPJD/S/J4WFZKLC0/2fq9IYWZpO+2Fcq84saXv8uSJKM01gG
S6GSk7ZySTg588WvmTjn+vT2qc+yDZs2K1As5QGN8igWuqlQnlLCW4sHgonnij/nO/mz/yETQhz/
zyBFflVSmjyc8i/CB5CaIyARv3utaUQzcSpYCwYw3r31afQWFRkQj7vIBD1DsftitK6cpxYK9Fog
9c7F0TwMneBGfF+CdYHr1YPr4fpbSnh6oYX6bySe7aJZqpmdORYGbAak7WiqWCmo3FcImJXSYSm7
vwy9nE9KLq6cweoCHJdO9HOHvTj2vIqoX7bd+iAtrKmsL5El2XfmYD/0mkOYB1QbvH28jwmwMG5Q
SvgPtutRFgyQoVtB+ieU8Rct35pZFl1wbrX1TjLCTzZurHA9/3/e9XogNSF50sZDPhftJJ5o91Jd
F4TUMMWgqNbNUFkCJSpc+cH3WwH/+vx1+26dJiNgo6ZDBi0aadKLESMte2tSitYRfEoOliy9OF2x
XSaHXcIPauf7WOnBmDgWmvbAqavWaoUeg/Bk0C1VkAa0PCu+q3uN4kCHJHZtxKkC3mhzunvj35W1
C39a5wm5Rs57zN13DUDALtFEXkB4NisjznZq/ZBUM/yPQm9wv1l+DGeYT/97QCX1Tjfpn/CHQr78
3byA1D/TXHOtbYC1CmGEPBgVIkq876XHuAJy4Wd9QI/EYVh+1GJfwodUQt9Z7zORKV1i8saidmQH
QzyZkca4A0FQAqoAikdlMzjDUw6IJp55EAguhtEImo3VgmfaX8UfXY2bEB9h9v1uJFVfufAGWaQR
vOSP89kIYNo/MXRnfW0mRTk1sQF+A/K2jKjZhAXrvVBIokuqDGbql70Gdel3YFHj5kJHCXApUzc8
qQ9TgaiPgziiLsoLc78utAUfjh72NWWxNlTEyybQdkMyMLJ6v6ywPy9fSLpTLBmMFkPIh7WSsTi3
EvmEgDoC710z0XUFhVZqpRDdvFEpN1ukHojipAZhAUcLah7a63W0wUlLqAyULqHtpjYxquLKHaE3
MaWLL+AAf+gJAZKcI7z889sbd/XAwvHHsZJLmcV14cv1b40TgzwROH+I8i64vJQx1RU7EYkhKGhV
2Zb0ZEYo4Q5pnDcjmVHIVz5JBjmIZNe2L4QDxU1B7NAoJQzdd7xFQ35URemJWK1vGjISvb11prQM
mOGjnl74WsWWa5SudjMT9e49lQbgyuwWKaQ3pLGRJX8JpKrhZfI7ZHnxQg68eLaSYin0UxMKu/i8
VVyxcYPZ6YoMWK8NgzO8L8iricdvzr1q9FnoqPOqwgpOgeKsSCFFutBX/gLyp6rx3tWE7lFGFZK6
iJ8SH6yztwr+ou7vbG7SS+xSffysh4uqVhTlMEE2G01YS4JyIBVWvpKGzCMWXqodLMFczSgg2Lyo
NodcyL4QUwcESvC50aWQsRVcSzcnE9JZ9ViHjHQ2D71gY3B/Q7fvMYfV4PcBNQzJUcmwsHVla6+2
2Wuu8yPAUdcJqunGv47sWBVakHq1ODx/FKZqbN862wVJ8z1AY9Mljeic8MagL61OFeeelskTFGh4
R21j5ufUzSl9kzRAQNGyTSxQbulGek74azCpUsmblUqlYcXFtzhldkESfvns6M5nBAMnAqrwTdl5
sjWeraZs1wGD8h8e97I1yMd/jJnXx2yfrGfdrR0e/2renYJbJ7VYemQ2OWxKjr66yDX+grogUyPX
ddVZC1pQ2+k6djbsUyAudgbwpqiHz68FFRObDeEZ4/es5p8U/BXT2CN+ynFMzoRjHZKknHfU1vcZ
Ml1wk4AAJIRAXoB8z9JTIf/qhvZxBujPXjSpv7hhZyE+cu7KoFmDfa8B0eFg0YiXtZJoMJJdg5ye
NSn33IiIwAc9LUHvUQQIcXGenCctNOdZQpyImJwhVcy1pCeeHySY1C9I09SkZz5d+A+cRvNyWrxi
ysoXwYk/Fv9TvCTkCljkbZ7GQQbwbQh3XNGLNZvK08xZ12B+HoVaVYhNYBL19/icY2FArr0bRdNC
/p9RUBJEzMDonkgdMsOm1UGE8Rq0EmB7kYxnWZH9XSBTKeUFKwDuHJHvaq03N72OFVKmHgFHsBBR
n+B/OI+pgu8h/ORjaZDCMxTCW9CtyL/AKBz6FjzkeDt62WQOn38sm0cWArFl2jQduuJtImH7kyNA
MJEE4wRYj2Y/UfOMHs32vurrDw3NbeMD0WzVfx7/byQeKaATLVcCzr1mDtFg6lPbG4PE40nNDqG9
BwUrmnAuljc+Kjq8BhYh91wDsgH0P8uULw04nJczg9KpJod/UAxykLDT6DrihGloVAbyb2cBTmAJ
pRbmg7f2pSgfnzWbvN+Dymhvu5xgR7Tu40fLiZepEuS1z8Kkslz9jSmmU41QJA64IfC4la7ThmkS
aiJn0Lert3ZIBYbMnpcTK3Eti3gzFalqXqMdT8gWSrOZG6hjkJmm5tJuR3V7eGStxlcZ0v14H62m
tigI0Y3xAtODFMwCdSI0+3HK2bgK2TUOkdrxsqUW7uOZIeAEOJBfrXG3/47tyxvckPKhDMUelVnA
cBTUXg6xOnqxmYl55Ugp/OfBPd9nbOp5tbRhOqB/gX5NQcHjRg3qtFmCwOv2UWBSOeJ3K1vkgClx
g+po82r8iMhV8mspehhYSCkHJ/NI5946Iqo+DxVbz4pe+BT7+BYN+URuOgmDOo666MuLOVPLf1ra
ewXaApPl3Y+9ygOijsm0eJalxPxZi5eifIDo89oRYDPSJgQo/e29E5s6FYx7GOF/awDrmOPrxqWX
5Ab133OZ2KH7l/6VxsO8ryk1eiaReOFehXs3tisE0f8/YkJcXTAcLBfs3L3jJXALvWSX/5fEoST+
Zl8O+dtoX7Fo88VC6r2OLkW3cDBYM2d3UgRQikjg+VQgETLfgeO19yxP2QLmCwssT8DloNck+a4w
B4cAbi+fkv5vOCwKHnE+oUSLxwNAf9BdCxNZ7alUQ7h2i4dzJ4fyvVm1loFClWZOmOL+2rjccgu9
VSPJuz4OhxaBBgTKSc/sx42tdEbQZhGd4CPpdmmKQ+kZGFHBABH8y6S5Q0j1Cg5JRrgXUEpmJcV7
+EIRVZSI9+MTAmv3d8ufRFtu/AQUy5MJGdaMuKBtyQ2x4R0t8WeLSXiEB+cpFLkB772XHgXTRFpp
TrMtAlaKgQeY6GFfu/7IVJCrTLuKtNzlXyfGOxDo7sdMLHYQzGJZYJlW01KSlr6B5BUCDcVDJ76l
cBhKz0KAHib+yEJjlp3hRm34/rNSkjGFjCidrb26K8Gxd2Li7Sz/4dngudIKYX/77ER4auXVXk43
/i0GDWLcsIVMm5tWwnLvj4kO7+X8RmIqPU0cmTcIpteBSWpMzhkyTpPJBRP3FTAmE7x/7guuevIm
TGF31sNWEJFomzLAXAv+vzTQ8p0ZTyb2gacRTRWBvAFISu/tDLvlzXrRh2WKkvpj5uDvCVmSCRtv
s37fpg/Ua5Ul5JrMjQSnUz6vq3f5Fzk2286I8e0tGXtgK2wuLDynECsydn2oBOAD/L/7+vW+egop
8sIIhJ5Pwi4IdC4KWD4wns+wNLiJpIUVoW8ejBaUnI0vDLuGozwc5vygwGv7fIiUy+4RGVhKr9PR
hPl+e2BvVwlKkC48oNeXJndYum2YGKNFT1CN6urS6MGoy5JHilLHCg8D27HOpEumiqw0OdE8MMep
bbBnNKAy9Ml77xdbw794kYsTZ/InwOJAZnrnKxkqnuQtamc+8Seiyh3naxvyZn48r9q6WCIfngWx
d8t8Fv3d3rIAfIc9oqDTqIOAuzFcf1NEOXkISNkXtCQwCtrG7c002V8iCJ0qV46fQjaam3god0dW
IuNJRdVD+2eHQVgEwhvq4VlbPWFt301uuzksvHQSBRMxREDuD1KcnVQgk+3hUG6Gf//RiU0niXJz
Eh4U/bsnYQyCUSjeV9ZikCC9vl3DV0KX/AwE6NS9LLwyZZrGyVKNwKMPlhY8ToJ7gVl4s1kgPXZP
GIB9adm094z/UpqpEylKfb4ACOmcJyHyX3Baz9kw2LUqWhdBuVeSFDHMUDi9BTEfX9upGd/byWWg
MPO8uj9VMtaqgrebmtQ2QxN77T3kVbIKgyNGm4Z0UDJL0S0fxcAmJepKCCZ+T8cL8DIipM0D4w9b
A9UXN2DM6yOIMGOMHbPXEyrTudKCWRLskZGKGtfeV1BSqaZ+8jjO7D3XTRan/qONmoO7QEAW8Ft/
kPyVV+AAmrJUXYeogeUkS0hsNY30dsiDPxnti0bMsCp7zPWj+affAVxXzEEcflAw4IWBYh0jSMNc
TzaSjnQdWOOSUQru4rzsKZ7lru++W7dIHn3RGprxRazJvMWQxtT+qS4mRQhPCVa9Lsvqz0Begfz+
aawe2gLqNAcEA8LE8YE97mkVTwk24ufm4cId0rxoxt/i1DFBWrW6rhOpN8b44LpyqX4JOVNjP9+I
WFwHC/1mMm9cPQusO4n5DfLzneIK4q+LEJkKXaLFUNmibNbb1rIer54NCqLlA4iPGrSsu3d7w+Nt
8jSjYbGrzPPgTsEl/sZMNtFFvlFlxQefjs3tI+DLYMzkO6w+tHChxqbWQZUHJB0QriHiVJweJ7Ao
UBMussWI5WmJgU9ZcWUKOR9M04rAVFXaRPPx9QVGczzUMZH8LTp4Xe8Zh+YCE0EfBgPmtTclHBxN
aTHP/zcxxxxs1jbOb+cOidxZ3l6hoXK5Vzt4FSFcp/wcu2DFGqBPucoSwgPmqChTO5OSDvmxlGiP
ude/AgzEbRGD6Uaw8XXPxH9VAnxf0hO6TW+88B+1mJqtn17iokbv0ECotw5RcxipYjRb9YcIjpoV
D+RY7xqPt7S+fX23TJjcJVCLEGAhF6c8e+pa6e9dHZcqqG2QucdPSWGUf6Y3Vt/g+exeGn3vU7wU
Sl25SNhh37fTN7f4C4oljYLeKjT+vIBQ1ho9wPp9C15/jcZBXKoI2GHZg3McJ5FuCsQxNEc8Je4C
nAq2xzHpRxGZU8osoBplVOVaD0zVPfLszh8YOQlX3s/1XLObJUjCgb4g0Y5l4gRLawU49YvucRVZ
H/BzM/1k6Yg4XD5TtOXRgVc8Tg/AHHjGBhN/Xf2yRCWtNq973MyLeBazO1M3Dg0hzxvUErdG/Bq6
6tRlVSJ0Oxr4cGZQ9Ac/HYsi6a3XaUEjaf/jyjE=
`protect end_protected
