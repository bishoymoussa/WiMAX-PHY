��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$Rx�y�<��wA�*;�x���@�̦�W�X�fa�M-$u����n~�%���P�$��W��kYَ���P7�?UMfT��q�6�U��k�>����~�\N�(�����X�e���/6U|)�X2pF�]$h���d.���9E��WG��L�X"]�Ad����ľS���8od����e�GT?y	7�������ݵ�^��R�q^]�鍦�����s�ae���h��L��P_���ާ��YЭF���'\��68�b�[����w8�[X��V�F�0͘3����q諵�uW� �h�u\V�?@��_6G�_�*�G���B�絉�f������[�G��U&�����~�F��AׯK1�`c��[<��FY���4I� �#�G��x[X�=�Q1��`��R>(�w����R�O�?����7�,(�H\�#h(W�EH=�������yq��Ѿ��aF����:�U~m<|��.��0=�P/���4ǆ���T(�����3�{r�_�SK3�\U����a�����-�SiB�tv"�f��&Rq0qFi{�}�Qpv��M��M��C��ʻY?�<Y��M-$�O���f8�Uk"�9BUS�o�62��g�L�s��f.R�_�U�� R��m�ߗ��Q����@ .��G�sZ�K� Y�C ��`�lU�f��ѥ�D�!��58 �v���-;*�ʛ�M�~�l��˽�/)Qx�q֏bxWY���L4�p�Yvq���]cC�=P1��=�a �ĝ�(��+i㣆J��\��(�C�Җ���R�YQ�v�.�����O�I�8N��DoK�}<����%K���]4���p�14C=$	Z����XE�|]M##�A�@.�ƾ7{��ه_��dh�b-eYJ�[��E�\����҄=g��T�2z��'� ��)�ض���İ���!27Uv��3�.�T� �/hh��/��� �'�w9,5�o*C���B�N���M~
vu�ױ$p{�$,}f�f�>���<����HcXӝz�C�4��2��=.��h!�3�)�qn���o�֔�(���q��9��$�U��Fq����e��c&m�9E�_�5�_�3B�Y_9�^�mVɑ�Eq�(���	��-Gb��C���Xx�Q���fTSy�r�ErKz���ڰq�x����iAM�����WȺ#=��rn���s�8�u2<m��򛶪���$2��9U}Ňa!�`����"k���+���K%B���H��Cd�Fr�u�-��Fǈc�:h��/���L*��ѰC�Q�@3[�7ٷa�W.k�̆�<l��)��Dˑ��r'��:�Rm�W�\�^���%�漖�~c�-�07��fl����\.d*5�I���A����wnC[�Q8.�{�W�`��Y��X!�%���T7
��b2�e�90V��
z\X�6E�ci�?6 �[��<1�źA�0|��?_�'߆�H�#B�wgqlؾ3���O�����$�.K��XL�2�Ի�ۑݽ{6�Z�&��O�9��锜�?`����!�)��To|4ih4B���]m����a�o�?{��mյ�;h��.<d�DT��>�JQi8�UD���	0��2L@A��=3f0O�m�+n���W~��6�a:%<���uO��C���We���2�jȴF��_�s�ϣC9	�����sĕi?J��1�'��u%?� �K�O�h�0���PZ�����#��O/(vE\kZ@��(n�r()W~�K]eJ�mse���R��n@�o��L�n΁Pt�Km��ar�<G»,�m��4aޮ�}��%YcR�43e�<�XN�=?��}�s��ԍ�\��'�f@Z��M�x�S�m�\�R�G�v�����n_+�}� �KIaU������7-�P�s;�5�	L���/���Q)�oi�~�f?)%�aá��ڮ�r\��6bW.��Ve�pW�kZ��Ϊ�_C�9I�㬼Q�C��5ߙ�3['��tԲђ,�����	���1A�9�%�-N r⼋���,�F/]�~+F�<�NȬ-������dмQc>o�튤	�ߴv��^I�k���̆* ��i�&����d�jiM���g^ yR��8o���r"�@'p[���	"�
�s�҃�8���&��24Nը��jf��C{Vf.8~?μ@M��%�[t�1�bB*�/�:\`�ŗ{�|����p6Y���P�֒8:kDּ�2L�#��֎�Qa��ݦ}�͗;��h�J�����C'�8����/�C����P�^n�U͢���ܴ�.f�9cR�Q��3ժR3i�\,?�n^����]���n��<<�=�2�� ��k�	�9��-���v3Fv@-k�I��[�Y���Аw�?HJ��/q�MPswv�wH��L`�>S"���p�V�c�hso�d}ٝ��]�3����yUfI����K	����k�u�y�(4}*�-W���<.�=%q|�1�Ѭ����F���d�*��Z�3y�[�Y��s	�VN�E�yL6��C.ޥx��
0ab��JB��]��������F��hj�E*�,���A����C��ǣ�i}Y&�l׹5=3��%h�zz.�_(Z?~O��E'R�O�>�:P���N��ή���x��3���T�۳�����9��;��
$L�/�,�ޘ�c���i�h1a���~G�]��/���Y�;��$d�#|9�A1��4�D+<�4Mқ�~��sl��Xm�r�K�F3<v͹�816��$�	o�%��uh4�{<�Yٜ*�觫T��WƯo�/�����m�n�4��[��4�ԏܕ(��$�j��`O�/\N�64 ��]��sN�O<|uS�nO�V���*}+r��vO��7��;���>
1/� )���_�&�')�*ŗĳs Ê�)��6<�j5n�;�����1��[�K�H�BM�-\��-j���p�Od���m|MӜ[+}�J��M���,:�-�\8�V~���Ǡӫ�Rq�	Ɣ@j	�=��lP��Xqlm�1����LR-��ύt����������peb���c�;HG�B^;lOMz�S8Z�gy���m�8�$o��=��^�j�m��2����|xrE����Lo��
�62�Ѻ �[.��Q�0V�w�<��� �p���M�������Bx����	�k�Z�t�~�V�UZ��A*k���c �O�!�1�J�do#��}W�[�!0j*��~�������NO^����#6�:5h�X�W�sV^a�@���\3se�����{����#Je`������nͩB;�̪h5ɜ�F)��u�����(��$�u�o/5/���k���ڏ���b��?����U��\#��R8����c�UP4i�}�:���$0��b/낥�@��:)$8&Z��0���u��]��@�J6Fz'KD���:l��U*y2�3�3\JD�gQz_\�rJN��zD���H�����U3U<=[�Ih���f8PANC�n���p�Z}���>�R�F�Z��l���(����Z���<Q��������({��㘤��g��|��+x�_��εi9��t��g:f.p�[K�ǭ�LD�,x�FmN�avs�#"��ɩ �=&ˏ�ޣ�H�ʂI
��2,ӥ��C/���.�@41,�2�
�U=�5b���W�EA1(��Abe�vn[���d�s�~���h1uB
2�I�3cG
�?��w�ys��ZW�ck�
}����|�`8�6ods�-h���<v���j�-Eן�Z&�ؼ'u���w��]��*�ABt��f�s����C[K6]���{����&��L�r�?�F�xƅ-�.���<�1����&z�����B"�'˞a,)e��7ܕ*�ı����f+�~<��)�u�A�l���>i��ޣ �l�n�7έ�o���<�7�J���ie�j��Rzע�4��'ˏ�tG����4FE\P�>b9{"��J��V��z��U�j�y��S��-��������<�3d�]�1��4{a�-�u&�]���B �<�C����� +��vq\�ڋF����W3:6�tF-6������j@ġaf���7�K��6��қ�D������c���YJ��� x�6�f4�&���N�����R�����/��\%~t�:�ڏY�\�E��YI��Q�mč���1�ڛ���a�ٞ��
����6(�޵o�'驾S�ڒ�cz-(R:�>�u�%o� ~�!	F��Dh�nQ��L�'���Z�����{�
/88O��{��"�܊��]�>�g-_��x��-PV���ys�Ǯ_b��kÑ~��O�jV��TZg��T��6p�>2ʵ+���4�^5�n�X��NU���ЯÞ����ང*fS	d�ć�Or�jc��e�'в<�&�����T�ߖ�?Y;�
92���%qL�R.88t-�7{j�	�{Ȯ� <qH���B������E{wt�]��|���/�-A5G �=�/�����SYF�t�+^�ς��y�@b�[N�4A��;�.�Q�M{����J���`D�$���@[�p_�O�ͷt0W���,1j2�8���֌u܈/��5�����8F�GsM�;��o�7#^�}�L�ȧ�c{�K�\�~kT˟��{c)�)m��H[�S=1������XeS�g���د[�M4�K�ce�z��L��U�R���I���ѹ_6d�m#s)�mU$#j"rC �ջ́@��5�LTTN�/<�:7d=�<p��W}��#��^�w6��dK6h��f�"/��wI�����!E1�s[��[ې}D��m�LG�f4쯱����p3^������4p�_������{1�䄹��.H.^���5��ڐܤe$�FI�~NˢT���I����>a6���+γ��c��:J(�?�X�C"���;F	�wD���re5�[p7�T�����Z[�ұ�3�'Bn�^[}g���q���5;�'[	<�Z�V�ٴsa�z�$J�F��S8���9f�
b׿z���͵8�tU�ޕY���ϊ�u+2�Prjm?ۯ�lμI���I|�gj�:�%����'7�$\=FZ�ńN���t7��9e�1��xd�:�z��Yq���� �.�%��I� E_��mr:���_-��^�-n5kbs�*
VюOep�s[��Q�psɆ���1�9s&��%��v�s:h:H�У�M�O�j����2�@�(��^�.ֵ;�����\�t�rӁ*��lF�,-Jo��Ixx*�^�^@�er��V���ݓ��.�]�)B�>�S���~��n�m?п�L��ZOĬN������S�SW�&�Iz�����t��$��UV��M�Ү���C4-��\����~�&lǍ)����h��R>�՟��#���-�z��7�B
lO�Ď�hcEg��}N&P.#9�	�Ť����)A"����	��IAw��.��s�*�.Y�=D
����'Nq�Y��l9`��'I5܎����"�A��*a�2,!����s�Q��WY0,�n��H��Sbc``�Dޓ�����9b![C@��2u�4M�1]��ڶ?�Tw�ݰ����u��(��I�����{�>���PU�P�hv��V*���>G�6O�����ƽ���b���
���X�v����p/�� H�a��nME����G5}fQ�1���$.Q0h{	���żH0��V�x��
/r�+_���^SS(qV�y�8�iTzZ/���m�}$�wc �3����X����I�˪˒p���+�d��¥�pG���%��܋�Ջȼۗ���B��.��m8���5{�:Jp�)�2�q�Q�13ɵ� 0B�K�"�?���$��7��]�R�m�6����6�_��Ӵʻ<�m�epc�>�*�\C��]H����������� Z$� ��➉Ht$�|v]o>�X�SJ���xk�^"|�3+�����1,�@�u���"�z�� H��M�!�5Ϫ���\�<3��4�M���t�B~d}���A�/�Yq�Y��iy	 �&$�=���+���Cp�(�S�6.�)B���C�i��M�8����Gf��m����i	H{�3&~�
	����굱�Zl��r$���li5~���6�=j9��O�y.�-BW��b�$�v�:��.�(G��"�7��3��[p�v ��
�Ր&�2.�f���٠3�)YQQΛ&~�NfE���5p^:�tڴ�O��x���d6����=[
=@�g0[SX ��(W��h��񂅑�0(v�)H���M$��"ݩ
����p�\p_˶�w�h�$�4���H�r����5�8�9�A�1�,�W�P �xa|=`�6DS�+k 8���*�����e���$t���<%D�i�.|b��ntB?xyJ�P;+H����K�D�C�����,���tPk�o�	�koC�!��R��R��9�j���zm	D[�,._��-���[�1"��]�+�"Ϳy�w���l����|���e�y�_�	����ɫ��a�=���~x6.O.�v�8mIȥ~W����4�7iq�:h1ڛAI�o)�K�*|���7�weB��%��{�b\Q��MM#|]U��dׅ�ߩ�ɹ�0���o�!���P/�'C9"�dk��,g��H�e#�%"9�0ߺ�Ƕ5��}��t4E�tb��uP��Pv�Hq�!.��O��(/�PcJhU�-�jZ
`�S8qc��g�0Jy��J*��}I�nq'���7��B�A��AW�in|g�B[LK�3�}�S��_(���--t�t��$Vom�/�W8��jG\w�	14"֥�l��]=�fu-SA�e�k�|긿lS0�6TU
����
�S�g�C�Mx����}%��O*�U-��u�y�M������X(�c��z �@�LS�`�g,PQ���u�"�x.�A��y�
J��0v�!�˪ Nh[��ٳ�ߢ���T�{�5�:@�T���=p`-% ��M��]۶��`\��ǥ6�g	+��5�;��[)��Y���^Ϟ�G&S7X��s,o;> �@'��Ʃ��5�t_4Y��%��ɏ̹l���X��!��fNKׯ?B?(�[��Y۱�y��B[
�����j��ε���9h���t6!(~ˏ�����|�b�]��k������H	��e��I�@rR5x��Sx��A�rW���!4M �s�����82��ѿ���P�es��Z��(�Sg�n�4���E��q�<��F���,�"��f�̅kd�Ch%��._�t�a��2j���B��2~6U�Q�SԿ�0���G���s�A: D|�� ����@DVG�5�"Jͭ�ʼ�R�3��ڜ֏�[�4������e��o��!�)wԕ�'�v�s�y�e�9��<�:��i���o��#��J��۱MOˁ"6H�k�_�5+�+��]����>���L�4��"8dj?�+��b���:��9��@����&�`�!��~��D#_���=�ŕ�V�LW��dhL��j$�'���w��`k�$�׎�93 O�u����8�ه����M!�_ ����Snp1����$�]��'�n0;�Ѱ˾��q�K���ؘЧ�
-s�eyө������|�$R�˩k���J;�K��Z�w�w�������;���P��_�QS��A�~�I�5�n-<1�+�K3�B���Q3:~�yk��o�����2+��! �x��!\�� ��&�	��������i�d˗R>z��;+B�_�9B�[K��m�g��CЁ�<��6��|yX�(i<7����|��m�4E��Y�g*T�H���s�b�į�
���k@��\ҙwr<��f5$�o��񤵧p<B.��t�V� �����t�;�3��[as1�1����)�#2:8��5e>D�(r���(OM���xj�����H Sqe|�G�c�O�y�tCz�)��������L�W&g��iF6�Nk���
����_���ϚC$_Bw�0B������("�,��k���)����Y�C�շ��6y߰��A�L�:�h�j�	@��܎of���,�0�ijѱ �)d\q��6\��^`��� r ?��WlCk��r�P�8�� СƮv=������fn��"j�$X���j�*�+|V��S��W�5gF.��g�(��z�/S�?��ΣD�h��'nc؏(L��×a�z�2��Yh}ߑJ:P1cK&��ˍ�"vlez�h��;T���8�aX�%?m�Q�}γ���5^��>D-�"zI�r���}�Ϻ��ڰX?v9G%Q���<�ijD��_�D8Yah
RC��
�L��N:Ϧ��ը�EL�����47�'��`�~�H�[2R��{��i0l��rYh������3��W�Dİx*,���Vud(`��w�����\��Gm��5���s�9k�:�E;�Qn�!vk�F���cjhA9z��0%��z	?$-	�	
�L�G t�Bp���}'�>YYX�fG�J���z�#��쾼�l�����ԔF�Ls� �mny�Z�V�7H	 ��6��ؙ�|i�N��� ��`=B`|/]�Yby+4�̏�t<�Y�z����۬=_���pq	��5%	F2��UFGBb��ت����oa�+���N�|k�/�ׯ��'�q:a��U�`���I����k�Q�3��\�]c����>�Z��ݐ�`t0z Փ��0p�|_�����.~q�.�i���X9��~��L8�{�9U��O�R ҵ��3
��&�)W☜�B��u��p/���~��B+I��Gh *,���f�����)�;��%W�FZ�[m��9�2]��q�or]K,(��j�����!\V�
��!��� #W�5w����0�,Y�b�BԴD�p\�����D�X�r������s��p�چB�Y;p��M*U�-!�5|���%J�V��l�]��q�g�i��g�����ěu����(߃�쯄�y��`�iVe�3˭�x+8-�)gF�������1�Z��.qs����>���o���y��c��W.>�f�]����_��0NT2�#x�9bq�Ɏ1+�=W*���o\�N�r�.�o���3�=��j�.�\2�j�#8Y��QW� evex�C�*����Z}��iG<E��?��w�<�?A���9��9*�&C�Z*No�$1��o|)�>�y�������]�[y2P��6YN�;@�]�Em��^hgH [���Ba�p]�9�;S��R�Q|Ʌ�qP٥��iԥ�P��N8ᴪh %�r=m��R��E&�6*�z��D��r>H`eq?��%s��k����R��DO��~�ʑ�U�Y�p�%V�Ju���u�d(b���ׇ�te�E�\-�w&T�g�C�΂�8�K��HxM�.�&R�7�@Hq�3�`���'������X��j��s�Ӕ�#T�����yV�T<Uf��]B$�JyFm:�DZ�Zh�#��94������{K��e�ϸ?��=�y�W+���>����Ӭ�8�7�������@�ǎ'�rl���3�ǎ����{^�������JE�;g��Wwc��>���$�6 e�	vs���WB���S��`|��[��`�x$�<cX���~ܧ�]���*B��M�ߝvF4h���=#��Ä�1{�"[0	Jt�]}Ϲ�^�ʍ|y8�[_Ni��ܦ��h��@�^g	���f5��0SH�2@��/p��/Hn��֨k�[�zJv�'��pc�K���+��E�ݩ����ῧ޹ϋ�'�M`p��U'��F�hˤ�tW�E���E�#(Pw���,R�.L���< ֓a����d�u�'�Fu�K����P��u٘2W��S���6�|�c�v��
|C�p�57x���H�Vv�����^�9��~_[$���^N:�#W+�b�a�;m&����aU�g�t��^�uZ�0�j�i�="���U^� ����^�g�|�	?��2e3��8aT//����AAE�ԩhe��o�[˭=i��z��/?)��VQ�7�t|�\D���l�32��U~_�Q��w� �{�'4q�Aʞ��n�J2� 5��攥����d�����bC6o�A��:�ğt�$ �5�"�+	��^5����q��ZƼ����a�By�R���/�%��m�S;�
Q>��?A���񧧳:��	���.�I��1+��ջ��qy%�"�譏�([>���Q
�eE��O�E���b������Ld~�H�º�#�uL	s^�L[݄ܦ��"`ehI?t�|�zmY�k0�;�E)�w$��Rѯ):\�i˄]�#\2���L���<��yɟ���ka�rHD"b,� ��1J�rQ.z�Y�*.u%AC�}/�ّ��o���T�ݜ9\��R-d�}� Wq�a$��$	���4����}�Eqq��bM���>�>�$���G]��>.Č�����< ı�������P��l�5jx����k��#)�@��r�.�ܖ���6fՌ^<�g�o���c�%j\�f\�cЦ�1��t����Kl��/rF�?�Q���*ȹǔ5�d8�\�)���bx�P r�3�jaK%���E>e�������pٮd�#�����z���$xl�t(�-�J�"�\���eN?M�Ҳ� q��c��y�#�~�u+�i:OU�g����q�v֛#�+j��w�m��ˣ�d+���C*a��&���b��2C�{)�O��������oٯ'�z	DPs)��}	t�U��}ߘ�>D%_TM%��@�Z
nـ[mG�x�`MPO�C��QM��Y�^Ө�gvJ��Ob�����ս�Q��+�J�cqs����\"��8õ�#X��=��?�]��g�]���o�X��
篚�H�dC�`�b��'0�e1���j�-Οߺ��!5��sd�tã���r�5@��pG4�	��x ���m�2?������jgw6�P��g~o�%_�Q;f_ ����4B)�r��m�=2���!'�y�E�~�"(:��W��ò�!��r ��J[q���v(d)�i�4��l��خ�����ʬ{�Qа`P����!����W��� ���Z�x<��m�T���0�z9M�e���,
�WlZxk�?��w3m}� ;ί׃��b���ܛ��d���roQ���-��9cE�.TEa�m{������wY���t����\w��;�����7)��r�M��y���A���2Q���	�6_X1RY7��G���胾���B'23؋�!	�ㅸZJI�!�/���.3ǽy`���}qE	߃�|X�,_�`d`OY��-���t��@қ���V�4�D��ܾ
�fgEp��7