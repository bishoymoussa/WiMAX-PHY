��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$Rx�y�<��wA�*;�x���@�̦�W�X�fa�M-$u����n~�%���P�$��W��kYَ���P7�?UMfT��q�6�U��k�>����~�\N�(�����X�e���/6U|)�X2pF�]$h���d.���9E��WG��L�X"]�Ad����ľS���8od����e�GT?y	7�������ݵ�^��R�q^]�鍦�����s�ae���h��L��P_���ާ��YЭF���'\��68�b�[����w8�[X��V�F�0͘3����q諵�uW� �h�u\V�?@��_6G�_�*�G���B�絉�f������[�G��U&�����~�F��AׯK1�`c��[<��FY���4I� �#�G��x[X�=�Q1��`��R>(�w����R�O�?����7�,(�H\�#h(W�EH=�������yq��Ѿ��aF����:�U~m<|��.��0=�P/���4ǆ�ZG��
Qb�KI� 	(lۍ0-�*�����z�
�Z�I��߇��-�G�x�<��v�"����1��p����r��V�Ͳ���$��Ӽ/IG3n��G 
��W�d/��ۮ,B�ni�-�HY�L"k��H"R�y@�Ջ���D�g�ɵqg� I�W#Z���p�DJU[RB��7�Dz+I�`dc��9p�dT��p,:��\94:Rtv.0ݱ�}RmHO�6QÜRx�y� 2���&omA[/J�+�I����6�M���<���j��F�����z3�>+C�1����J���X$��o��	[jUhB��l���a��%X�Tq�z �f�7����Y��:@��	V���6Y�%���p���r���W&��:-4P w�=�b����	8d�H2Gq",C��9��C�l��F�{�̕����'�)֪���kL8�>c3��cd�ݶq;��ͧw,@3���}S�$fYލ��{{Y���9�E6�@�Mqj��->�zLF$�X��n/Q3$�;������jo�,1���$*�Q��%�r�H��\=L� ��w}�� ޳>^����>��۞��i�W�G�ϔ	��Z�!8Q����Cy~Ӌ�GY1�1B��Q��I���72�|���{�NS�jXJ.��X�oȬ�� &�r&c/0�˾
:�� nʕ�D�'!fq ������pj��`W�.-g��Y��Q�֖���L�`��ꏿt�ƿ�^�m���K�;h@b��X�>��|�����`�J�����b�]K[SW���X�2����[���vG��XV���r_��EޘR^�W�jWz����r-�;6Y�iÏ�A<�F���G�t�����.$��?ݐ�w�����a�Ɨ����#�t<�U"��T�V����⑤��X%	��db���0F�̘�6��_mS�B��F@�.�_�WPSci��������`pq�&����<0���g�D�W�b���\j uWܼ�X%4�T��9�k�P�^���Y(a"��M�r�
�Z �|r��vʳ�~�5�)�\�2ϑ]��!����B̌Wh�7)��~�q���E�B@Y�`C�d!�{�� �=�$Y�[�K+����6�m���=��fߺ>
ǳ ������P��
��I�*P��3�B#i���}��F���n>X3pځJ�~��(�L&�ӷq����ύ���B��ݥ�(E��1@(��B����4 l`���9b�#�lPJb���0��A̡+�b~�0`58��N�z���MlD�K-���/�ܥ���a��E}�1�B` -e��n>ۓ��=�ړ��=|�nS�.�*ص��)�#|�uD�z��S^Ŗ�Q�rA=g�+ x7�k�՟��uȒoT�������
���5���aH��gG['��������00 �V�-�"}���C�\�q�Q��!"�C��z�$M�RAQ��r�������-"仏��}�ݑ�@(O��̪��"��𷼱��H'p�_ �G�j������@�����=�!RUm���Q##E��������2��$,T�ήfuIn7Av�`h�/��t[t��f��s�{au�{|��Q(����xl���#�DH����1�A����W����`l�{��
q9�ܥZ��2V��l%7cb�ޮ�,߇�;(��*���y��_Pe����)�@q������w�?;�fO3�ON��ޏ6J��M�>
��n����.L�A�c̮B��"�[��Y���J%۫�W�Hx��Y�L�^:��[�2_	������5G�S��c��'��=Mu#��Qk�"��;nQHL�.�F�u�k�ѫ:��r�1ѹ>X�"��D�S�ֈ���Ξ��zY������i�a~�Ց����s�#<۬@A	�8�^^KQU�$0�
Ũq�t��g\z
p̗���K=�2,��)Х}��AF�
4�KW9�F�<X�[۳��PE��jf�]4 �q���f#��H�մ��{����~R�/��*�����o��F"�[��B�E�i��:��͐��g^�S��<{k�2~�y��X���Z ����5��[9�/d��ѩ��C�#?��c諡L�9�1Q#O��g�̶/�@[ŧ�k��i�pA ے2H�te�3��l�P6�x�ޠ������Iyɠ
�l"���)M?� H/W�AX�9�no��k��p��y9�<d``� �ɗ ��֛��[�ޏ�5U\HV'�՝����2nX��mx��+qo5
�D1Gwjӭu���y٥����(1}�u ��eև\_�3532�$}�A�)�j�����K��O��lI�@¸8y�5�Q��؎�QV{�;�nUe��c˪oM���?D�]cu!J�*[
b��IR�EW�����hq�4���zf��N$x��,ڷ�c���7#ml��WL���P�c�;3�����A��! m���yT;zh*�mؕ���tR�� Z�7�!Y�D��ĆZ��KZ6��Z�⃺��GW���t�V�,��U"�[��E �~MB6������+�c��p�+���wn�L�uZ� 2�dJ���xb��%B�S',}$��쐏����R��#_S'`ܟ^�@_$��P��j�x;��&mF�[#�?Q�Z�V#�WP�*t&fwk疕?�mɈvܦ�����»�=.�(	X��a��W�Ǝ�Ź=�B��l3cm� �h��w��Q�X�[{ƕ��Z8��'�O���*�e�Ί¡��b?��:Ne	��X��
���v��z`�+�ݐ�&���~�l�b/S�86
W���&H9K���- ;�`��Ν_���˖*s���a\�h8�ԁ��\��85~=�|�fm��w�u��%�Y�_����>�bMz˦G`pT<�D�%�~;d;��5����AQ�E�ՑBGlsa}�����l�.B3Vx�n2k0�l�I�N(^���U���ɗf+���W���Qv�O-��ؤ����^�H.ѭ�q���6�
�1��ҧ����m����-��������Y~��Klݭ��~�+����+���~����!���ľ`�����-��h�6�J��{���J�bq�� ��]o��F� A�>So8�|���͑�㎡�q�d$V�6�#��*&?=xX�!g�a:�&����DG-@S�V>�x��$0�d�����9��+�/5)���r�����$`�����7���s7#��%��WI��*���|B^���u��B>=�1y��o|��#(�qU
��:�;���aO��JP,>��؞� I���{�Q��~�'��$�-���_�-�Z�t�3����M�ֺ�}��	G�γ~�c������6J*��V�0�z�D���<�	�t��'4d'T���MF���{/C�����D]�z�-i!��83���f�D�:�����Foo3�а�Q81��s~��l,B��A2z�Lp�S"3!@0t��L%�ǓS!���`M��>������
��� �b�Ǥ�n��-���A�h��)���zHZ3@4-e����*ɯ��(�b����8 Ռa�/sɰ�Kn�ݲg�e:�,)*[o1�>���_���t��G�:O����`�(B��̅Uר��6N��h���f7[�{���튞԰�o�oCt>sp]Ɓ��}:4_�K{�fkg���1����.��M��L��Y�7�kv�����j>��A�&�;?�Uh�tH�q��#�E���'  �$��e�	fl��m}@Z-h<{QF�^�O��Va�t�r�@ա��8}7G��e:KH��[L��uw���-}�����P��W`%F�Ԩw V�GrG���_pf\d
���e=��]�cb���=�/�:��8�G;6ͅ!.l�F�af�7۽�I�Ґ���ف�Fx��e�z�x��F��>M�w<�4��k�.� vaA^��Z��Rذ͙z�����mQe�Sxx���1��(_��$ca�z�Ľ<YF��,�E� ��Opp+�n
��(Ϯn���ø�4F,���_Q�UM��̫��#Q WA����-n;����o����(�����F��9�F{3x��#�(��t���#n�?�C�3L�+4�k��i5�����&-)<` �O���#�@k�w�+{w���B�����	���${�IW�N\��-v��soӖ�#�<I�0x_�,ugRA��WY��f>�a\E�I9�]��k�,�U�5��	��3>�o��<d��N�1jv-C�/��}��^�i|W�^�J�NnMı�L`M>��A%�*�i��Ps2�ƛT<VP���8��W=��D��u�+�v�g��By0Ȇ�p����dx�~$A�L��2����� ބ��)��au�h�u&>m��Pzӏ�bgpa����yD�,ݾ�ֿ���FW�崚�N�Z#ԬVV/�@Fʲ@�jy!xϬ+6�!����
������w~S�ܚ�Z�E��*axZ��͗1�^�+�Z����UMbOb�O���(�1�R ���	��ٟ���$q�sZ'`�;ur*�qAE'��X�d@�b����w8dE�����d�l��Yg�)��.�'�$�cu�>�>�@}��&��Q��&�~l�Bfs$���Fņ�m�Y��ߛ�%"��������x�������-|�$ڗ�꡴��h�����R��������+O�ɡE�E2$��ßY0�=���o�%��cT���8Չ��yƵg����jקB�������u<+� Ɨ=��<P���� ��|Q�y��5�L8^��k�%�u�aR����K� Z4`[�J�dM-O�rj��Sx%�(_%d}���	i�;�����[{�-����R7$���x����!L�(��!���m$�`:�pw'yi�=�]^O5J��rd��NumE˹U6lU���T�(u��(�"x�&6�I�#�o)Q�p�u�= �	�{j��)Ue�x����u��N��)��^G�0�38:��L�������ht���CG����#�qV�����m�:�����H�?��	3�-�c.�vɞ����Z�P���i���r��������kL�<#�4��)���z�����AE��:�Ҧ˧~�`�6���vpl,�o:��-�/҉#����OA�~��2v߆��K��F;ʠ��(�W����2�"�.�Yz IjM��J�ѻۿ���������#�&x��QbЬ�h��8D�g|.�U:���
=��m�^��d}g#�UȰ�H*Q��@��	�K�LD`�b�)	yG����e��a��o�r�����R�MM���Y�ײ���u
G�!r	��洒0��r��,�����LG	����(�Py��A!ʏ�lZ�=�x��OiY�-зMN;�P��:� W�vV�����KO?�%�|��>��m�P��4wDƽ|@��"T����1be��U�d�\�����/�&�~����B��͢��o���b����*c2��ΐ1����nZGT(l��]�U+����y6��Sy�K��sf㍫u�4�����G��3ٽS�cȥ�дjr��	�v�N3l�~Bӥ3F6A��gP��?_��k��lZJ��?�V�:�k�0N��}�2z�)�mOB�{�d��^���Wɰ�p���D�?�Ҥ�J��6�+���#O�����KBs�4sG�\�1�[*������5bfZĝ�n|c�I��s�>k�=�収LZ(T{K�S��@�"������W����2�u���ڨp}{B�=����0;YL�p��^���[+��#:�z��bm�|��hw�g�(-�v���GK���F lNK���~
"&��w�"�W�&��p��p�9��˲�4m=G�R��H�6tz�;MYut��Q�����!ԙ`1�N� ja�Ql6!w_��wi^�vD#�;��b��A�Ca��Y�З�mT��׵k�c'�G-Gx�T��0�. �<ɒ�����L�5�A~��Ġ��`��0�=o��[�B{��h�!���''����;j uB��a\�jC�j�ü#o����,�stY��U�i7�>��3��C�݀�K�\y"_~�u��޸$@b��� 
�;W�e�W���ŧ
O�;N�[�z�'�|J��������CՌ�G{%Q��Ao��{�L�c�p7AB"J ݫqrS `���l������S�I�p��"&�gD�[��,n���_M�͏��d���(�ɹ�S\5�tM:���W�����?�B� *P�f�	&���dmPZ�bt),�����Y^��ۺ���B������j򍸾�s��б�>U�h�����@�:�����$��7OE�R}�G�37A�U�r�6��r�k��d��=�8Y�μ����ufʶ�����X��>��&ٞF�	2-�D�Y���m����N*���I/���?������{�)b������b�X7��:�v6��@)h�������M�̰��J[[x��c��H�v(�	Q���I�0J¶߂Vhci������&��1k'������;Ҡ� 0��mZ�����-rP��o�.>'��#�.�|���j׽�Ew�EEa,Gq�yL5
�ww~���D?�ۀ�������
g����j�����
I�:�RyI��A����	��Ρ�V�?,m?
��Vu�����X��@}��TUI�N������FQ�h�K[�g����y�q�0k�w�Sc���f�`�p��t�(�2������0����\v���������R?W�K
^z���r�>����-�Vi�������cDbE4d�����n��R����;oÒ��!��rn�t�t���I����S�S�(O�/����'2 �.�y�j&��j��=�T_�ܸC�Nr?��O����]3ٗ�TW*�}�POn<�UﰚJ�_O��j=��!���Lgl�Iҳ�(�}���n�(TWHUڝ����l=��7f>��&jYq��a<��A+lM�.|��%NN]��.W�|Yy��Y�/��)UEw��=�CU3�/��/�*p�9il5�(դ�Y��ܻ`˥����`L���V�����ȩP	�CTX�]��@d�I\���j�%�|����%&�#'�"ۣh\:�.��t��$2;K<X������v��O��FŠ��[9x1��׮��5?�&����&GG1�E�U�L u7;>���>�X�W���`\jO�u(p|-�5B�#;�JG�v`�wG��H���RdY{��Ы�JICZk�����gg��~{ ,�����P��>:*>��83^'Zy��r���r��:�?[j�Z�0�Z�Y�÷��tU=8oxjL�J
N�t������7�k�B HL1[���������To��*AD�Cٳ�Z���o����ޮE�PK��5�d���`9н�Bs]L2<r�q���
�(�&�x}����y��I�)}�J���m<�+��(�'Q�i~'�ܧ����]h�n��k�)D����3�-��Wt�c�y�IS)��������djm	޷��F)�لPF�L��h^
A�^���#0�X0�U_��k�w���B����[R+U�I�f���'���sF&q�(o�V1�1�d�̷V��%������O/2V�:(W:Q~נW�����Mw¼w�FƓ����j�ru��BW�]�+��ω� [��'�wS[C���W��Ss�ɻD3��@�����c���ͺ��Z" o}�:N�E^ޯi��S�d� ?��g���$0�iq�*�!�Bz۩1�_e+��2�eQgTDC�����u�&���%��t���|��6s���
�?�FEW�)Z�� v1�����v%�;��$�2��~X��_HE�(�֧���H�$]�Ï;c�u�x�m�2����΋���*t�{0�z)���!:�E%�f��	�� u��+���%FB�Z�?^���9�-�nS6�#�&��t�EL�4|���0E�rޯ1|�rF���6Ti�a�x�' �ŌKe�s�\�@~�<�.X>p�҉���.�}g찼����^PM޷�pzKt3�2�~Z�#�,��p\�톷����!��c<4���Z�Vae�8��c{�H���`,A��-O-�ɾn�� U��c��n �|�fѻ�E�
h�`���S����#�x�%�_X5�Z)�%"���b_�(cq�q��QXw�<
�s�M2E�������I��l�{1�Q:ݭ�J�D���ُ�?��t�Y:��H����?��Y�<��fP ������
^��_�D2�jS3�p'����B����`!5��ꭠ�@S��º,{�:�[#�������t��H5+���<��DG��ȣ�Ӓs�y� ��@.	�����0ia�rE�m�`��4�rnHB������
~��/� �m�=��(!=�>�h�k�y��}�V�[�}��7�G�7ĵ��#6��,N��-	�Ϡء՟���d�(�/��M�t?3�k�<��xH��{��iQ^ى{dU�M�B�Z?uqZSö�%H����Bϱ��a��oR�>��&���J�-`L'���M^�'��z����nz���y�d�S3Lz3�.���.d,�WEv3��%�0xN�ܫ������]�g%�a���c�W��!�i_8�D������D��#"�g�P����0�r�ݣfc( �� y������!�����#t��E���4���B�bo1~}'�+��T�0zyS�� ��NQ�FO�ïo��u)Ŭ
���J3���09����6���L�ze��@8��ƹ���m��A��y~��.�vªƫw��v��o��S����@�Ԧ��6MiƂ�{��r�b:6�q��b�[րu��ɎIy�cG��B�q�ɝ"N����D֮I��%f&�HVj���<d c��X]�/�D.$���ˣS�_��+�
�lG�������sؒ��n�(ۘ��f�v�t`�s�Dm҆ШS8�=nu���%\OQC
�	��{�P��Mk%$C�J�l�O��������/����,_lp����%�bu���K� ��/6K����j	ӭڛ�r١~�~�h�;;:+� ��Q��,72G��X������*�e���1��;OD+�P/&�g������&��{<�7��W&��?�q<�%v�!U�u�0Iϼ�7�:6˓���l�a���O�����v�a1�f�ض��Ho��
�4���O^y�9�j��Lt�)	�r���eZ����R�TIb�1���q3�<�I�aG#	6�(�ʜmPZ��\�5N�龆8��9��)5/>A��m̌پ�:��S�K�x$?�F��X����^6��{o_O�4/�$����$|��l ��8K>��x��=X�ꗆ��0 �(nz����4�����%;"��l��I>Ȇ�4�<	������t�:�Ey����1�*���(i�6�x�Z�=�!4<R�EV��"�+��Ԍ�$��߂^^�Qp���"�Y��5}�ʾy*9���h��E�qP�jc(E����4�;����t��ݑ�ua���4~��tj[	a<gRŜ��=Ko3�3[�1=���@�>
^�J[�N��[��R)U���A�s��X
N�[��DF&@vhM�P���
�3C�� �H���]��7^����m'�3�ߐ����qz0+<�D���.L%a��<��%����e��2����Wl��W޺� Rz%��N}hfh�xY�%�tź�>C�7�3��2������������&ͻL�Ɍ�pϼr���%lP���aN���OVa(�˻��>�`\�qc�3e,|X����#�T0��124�w��cB����L�C�k�][���e�:���Օ��@�~"[���J����Z��5ڹC�"����N=%����y�͖��Sh�aa4�� K����~r<�Z_�T�}	Ays��EutԬQ�䜡і�CgB�����/h�<�]�-�t��,h��| ���}����{7�d}��V@�g\��Tg�n�=d��R�T5��*a>x�!�hI r�5B�U"�V׭`�� ���j��f�,����< �[/�.��4�q��X�I>��<x�������Q�	�GU,n���
��^��#R�0���N����hV�:�сX}l
Z�1îu�fNh�ex9�s���c3�ܔ�@
�.O�盄�m�سgI\��D$
�e��I�6��N����EŔĉʙu9yl�J��^���%�z!y$+d��sfO�h�����j��	�1��נ9��A�-Z���r��%�z�00T�IN��(�;
f�T'��1���ٛ/C����.�1BG7*��9�`���]��\�$�]�ՙ=̉'i���*ZbI�I���1?���d$�+ŷ�'�����n7 X�ϭgd7д�hl5J�ė(��?\��{�'���Y��}�9`�����+�;I��+��F�L�EM�$�ˊ�C�uv�5���~ī��	�|�m�Ř�Xcƨ��×^̭�J)��1ˍݱ�|h�9��鶕�By��AJ�p5zA��/μ5���-
?u�O�kEU;�?�	��7~D���>�ӱ]�4��6<��n?"QoS��*nG��5z��Ǌ�R�A�[�zZ�����#�X-���o��1�d5�ƿk�GR��	Jgj�{����fI$�k�m �\�<O�ˋة����H�F���/�x�=�C����K~�Gu��=S:��k�V�bP�gF�~D�����l����c�i]��8�Up��1�� ��R?�%-{Hbw܄�dg7[���9T�(9ud�����?��5~�0
:�=q��E���Ds����0���ԜE@�*�|<}RH����ۏ����.7Y��	*��Wy2�~oVH��/;Z^{��
;4v$}=��c�c`�U�����<��r���l����<�[2r�҄>>���}Ā~{llW����EoQ��7�F�]"W�����7p��ڵ5H�5��q��Q)P�6�q5�UD
��;�^<�>$������z����-��J�kV/ŭ�n888�,j��q���% IP�� �f^g5�T���G��Yw�<S�v�,'h��]恃n>O�C��X�R�P#>"?����^fW
���H��r� _��9Su�}.����`�#����w/��y�2��H�w�L��9{V��/9�)�p��^�*k�tv�y��mO���z�2��q�g�O#`�J����H]3��n'�MR�_��#%������
�����n���._n` )[�'P��S�{����x�r���a�a�;�O�����D�gĶ@U@�9���*�_~0틪&�+/2��i�2Fs�i�$�QI�I���������GLa*�kH�=������h�,�'�h�EbdJZ�9q�X1�Ѿ�⧤�ժT	Sn�YZ^����R���9u����d���ߚ،L���v\�k�qJ�^�ě��Pk�BH�.v���$�,$��CT�lfs�I��-j��un|5sùg1QܴP�tt�D9UP���%���4� �)�=L;#�d���6��st��X��_�TZd�W�=�$4h�O��*�u���13O�Q������؅v�憌!�U�^���v7��</Y[�����xO�o���ՕIko�Oڔ���e_Ẕ����`�oq���O3�T�i��ϧ�`i/���K�0���g9H��O`0|���PY2V�i9�g(�P���$q��A�Z����;d�7�HY���8l`d��{�E���.|�U�^ �.�WS��8`j�D7PB�k(�i�E���⾶�{j���R��y��L,4Ư�q�|kj��nE�N�Г�E킵��8�"� -��u�� ���0�h���:��a@�n(G���$�0g�����:Y�����B_��w|��S�t\{ �²�/�f��S+@����Ǵ�G�"�p��P�@��
�� 9j�hČ)[���F��s��	T�����[�S,�sD�n��>��\oԟ��0m�l�4���ݨ�~��l4�er�@֤7�~�a�oL����|��d�Ց�e�$QK�d+���b3^ٚ���8Z*@�����2l���D�'����l]9XS)��
- �����ͷ|�L���1rF�$�#/���>�I��V��4�Cd�"�1���i�<��k\�ұ�bO"b�|�yҡ��O+�:��S��o�FT�E���4I$z,6�&"F�Y���i���7�q,��Sre�l�Q�N+�j�A�觩�D��S��k=���Ǧ�4lc;�g�yI�%{�h�*!�=N9�n�(���
����SYm��u�p폠R�F�A�a��e���̳C�X��'T�Ƥ��U0��1��ꃢ���t���l�W�'���^���Ri/��>�F�g,�@�O{j^��r]9�X����X0!n,y����#C,zعQ~��(Sq�V[J�Y{��W8!3���l�H����&�W�~v�.�j�{��M�*_{w��Hc"0���t���k���v���4vzStu4�ϊ�*N�4�떳\��W�P��}>���K#C�%g��{��UE�B1������-F2�>���s5��ƌغǲw�3���?�=p��T��huJ� ף��;N����1���P$��>8�x2610}d�Z��r�:��A��gw7�p��_}�?G��.�F3��<�ݡ� �Ε@k� t�W��D:c��kG��1�qt�Z�v��L�q�l
HGxZh�<�:U$���7Z<��N��p��"N��c� =�~hQ&�Y�/�fo�#��QC,u�l�s�n� �Ę]��t:kV�t@�k'���� G�~��@$�^�#4��sOָ�2�x����!�R?E�����ъ�s`�ef<��܊1�j�}�ê��峩�h��X	G��'��H�(y�����ЧD�sWR\Fp�	3�홃��B�I$�M�X�h�q��\�Zq����_X{&d��$��Ѷ�)lgS\��`���T/�����l�j  ������6"P���$�S��u��k�qi��}��]��č�SB����NY<Z�>�v?���a ����,��5N	����H�v����b�uY��ːa'Ju7����z���P�fּ}�h7��:�Ռ�%b�Jzi	�
0S�2m��+q���F�:��3uY#��&c{��qį�:�����T�����T#���VǄ*���/�+x#Pۢ~�%n
*�1TѣQ�TU�N��9&�� @[M�ѺT!�~���+z��;Q6�F]����0�*|�s8�V�*э+�x�]tKj�����~���Ù���a>,�T�uρұ��7�T��_��3FO�����j��&?'��Ѷ�a4�C�t9���1��:�q8l2��Bz2pn���ݨ�S+�s�R79�4D�J -5�o�[0�>/k�ۯ�(K��(hZ�mOrA)>)F�����'~�X��`������u�X���˂�w��y�:$����Ia�h��̿ey ���6���&�Ϩ��~����[�s
�tW�;,(�p!�H;���J�|'R3#o�����d���y�<��l�*��W�^RP����'�&�_��Z�}���"o�\�M|�F�X���iagi�g�m��"*���[�d8[9�ߞ`��b�@g��Η�eD	T��6d�<ñ�Msmtܼ����� ����7M7 u\���\��wn�jߋ��w���O���>Dt��i�݅�>]�P�I�:��ϴ	�ʂ�3[��EƬe�b��:F�ǀ�n5�s:K\��؁��x��2�S*��91k�NS9J:׏CҮ���s���%�s,܏X*�%˟�&��"�L�j�貤����f�SnE����|̽Np�Z�wS��82����џD!&��EYbpǦ*q][�9f��nT�8����bM�Ba�����M� <�8�v����Y�'��_�7��[�P2�p5���R
���� (� �� ���hU}�$lg�h�^z�B���v���l=N-�r�r��7�cR��T��s���xO!���Վ���9����L�=5���R�A��5'��8���`�S�u9 �j�E���Rļ�t�X�NR�Mi�@�i�D��k��e�M��l�g7p�z�^����oe�T�k$�d{h
>��|���͍����% ��ڿ��KY3��a�p�݂��>�֎N���!�P�P�"��ڣ��<��h��>�9"x)p���4O�7H��[��j�Я��i���#�Q,4�M �<�ܴ���?XnRb�V��1�$im�� �
�s`�?4 �������`^�vT=Y!�������>n��JN��W8�<�Zϧ�J�����gw�!n}��|�q�� 8���d�ǰ�诉e�/���QJW��{�_&����s���Y�zK����G��G/y.�p��3l��T�o��������j[s�0\��{튟ѕf�D���66�h� �g:�k�#����9�E��>r����v�5���tq֘#RL����>P>���8I�#��ɼ��y[��2؂��(�͐��>L�K���/@[�~	F��R���C�1¯z�?H� 2�b0ɂm")�S�����JV1S�?���� wç�m����f�iCL���3W,�z��bz��!���p
��.��n�9^�s�<�@�gr^F�x=ʗv�x�^l��}Hb��f���¿���^e���m�>՛Zϑ@�l����u0���'�4�dr�F��S�؜���QT��EU�FF�﷌#-|ݟ ��x��|Ho��e)�G���������@�>���h"�h�a)�g��f�1�p��Fa>�q>Q�@���T\��#��|!���k#?ќ�Y����WND��ƛ�!1��:\z��]8��:�ſ�Y��u�e�6���7�
Z!��7� h��6����2��9�a ?�A�tm'$n��&>�B] V/%k�Z�;�Y�0?t�j��\�>G���A=A��F;�8�ᨲt�^3��/J1��y���,=�=�=���I�ҳLg��#��&x�Պ��S@_q�N�'n�$ݦ5){�1��@���������_Uk��(a����p�p�(�iW�Z��Y)n<�O�]�&Ew���9������W�*F}�ŗN!�u��B_��E�a*X��oz$�_}[� �X	�QW(@K���(	�&#.b��L,}!����[gW���vJ��:A��	m:���O�o,�ibW�����ЁaV��l�_T�U�F\E�~]���+c�e�ֳ��o�X�'����'�hh	��U�mZ7�䉰��h�gy�����?:.���*�Cp�ki�b�$:/��&�J
�D�����Wj��p��c,�D�!���h�1���F&���1��)@W(�uѿύ��2%�K�yi4v{����h��!I�?�k��<Ԁ��p�D���:�f�s���ݕV]�a�[Ǉ aǗ-J��
m�v�x�An�_a�v �_��ܼZn�q �S��P[��;����>Γ�_�ߐ��(9LHi���Z�Q_ʡ&�y�B<���)��Fk	�[��@z<��[���w�|����a���X��#�#�G�� �z��ХUQ�$:���D�_�|�Jʿ_1^���3*�K	�v����Y��cN�?X���.b&cw��R�B���<����k 44U\���N�1�`=�̜�!���y���
�,K.�n'0zo��P��|����$� X�7tå��p�d$��-�������7trOD�ivګ��^�G:�1�5��2�pS�4bOuݽTk��Rk�hf�7�=��*Um/�� a!�U5��p�o�i}Q�Cc�H=`��� ���z6�x-I˯��yW��0TTT|��R����Y���洘o�G��*2o:��H�*���5��{2��� �i�b�!�T�A^I��a�yo"��!��;хU���4�"����Ω�����W�	�:�as���z�5�]�imgP.cR�1c)�'lA$�<D�]l��+�g��򋁘P�e�"�@�;��e�%�V� P�e��i4\8���|҆\�%ʡaβ���
���B{Q`����3��gz�T���}۟��	#v:����)���2��d��[`P/T�IziXy�;��09�����@��O:p����~����bL��;��.����c���`�0ߚ��g��Ǿ[sE����m�����GUKo�7H�w3H���yD�ڸ���������u�Ԣ�o�����%�{7����~�̬uP�	�xc��(�������`\���@ӯ�3P��{KՁ�ߓ]{����r�6�x�ۗ�7p>,�56�dXܖ�ָ2�������/ *�A��Õ�OJ����#�ө��7�
��06�	���/��>��8Z��N�N��)�DjS��6�	��l��r�����,cqʮ<�5�=&f�p���W�^E���8{A��L^2bp�������O,����sw�7z�,��Z��mԌjI��k#o��6Q(�15-I -4�r!�,[�J�z���L0d���Zd�p�� S��w>^�o�|��ޙ0�8М>v*�j�a.w�XuW�_,S6W�w!��Cf�n~�M����TnƩ: :���ڎ�%X�_kx�D�%�oĞ�����}�2��5�+� +�b%�IGZ%�UMw?���D� �y����%0�^�,�컂J����_��N�����6E�-��?ҟ~WJ�QoC�}@�X�2�D�F�S/�/���B�:w��dJ'#�J���x��!��!|"��&̰Z���	:G��B��C�NjW�-K��0Ǥi�1�½���R��YЇ���%+�6K̤7V$��"�Ȼ��*1۵.�>5%���:�T�Lư��4�]p	.Ɣ�<����yJc'?a�R-�1)C�V��4�h_�:�4�z	>����J#�ڝZ2��T~UӰGHM3y�g)#�(~�8L�_g��Ҹ`�������C����q�8��T%�nwap��%�X t�r18�o����'�c3Uо��x)ds�9�$�k��8�^b�u��N���4iY�p19���F>��`ރj%�?J���$o�pt�±��m<��G4��3���Q��6��:��`��?n�j�@K��W��.~����u���C�7�WM�*2��?�f5X�$S+_C����S����OfA@���p��5�{z�q5�����_~ND�C��=��GPnK��3fC�~�e
�⻎�~Vu'<zbT[#�l�1!AH�C� D��\��z}�2�'�(rb��z�e�-8`�T�ŏ��I�MtgU�%��@�|��|5���Ye�b�H.�k1��*8!#�7FE�%`�r����vqK�P6?��vb���Jt�n�p
�T���A���w����J��Xݸ;��OT"p�3������{���u��,d�da��r<�{b֧L��%�-qZDw������+�"�8�ͅ�:�:����� ���ˋ�2�i?���ޫt�FHK��-�FUa1 �+��#���q��=-���VM��!9�Zm�b �9�v�����s� \�����n�ҭ0go��l�����/7�E�rzfw�r�s����z��3K�ќ⤀�"m2�^����2�kPӋ�t�_��7-[��N�
w=n�~��������c�������i�<ޒwT,c�.fK�4��y�`�M��h|a4�fd���$G:'��)�t��a�Å_9ߒ�����i�Ɇ0}4:�gen����ޙ'fiU{J������q�H �rHQ+\�la�_��w�fD%GV� M��3I�0�Es0�,����	�?]�X��M��L(6)�z'�T�����Q�J3�����3��E^��	�I|R@�H5LD��{Q��^��{��H(d ��Ö�8s�O�!���q.%s��P��w�A�7��%Ƈ
���w�t���e��	�U�,&dZK��I�4�\��߾7�=�IF�9G��,����ɚ[oH�~�*f�:_���vE�ڬ&ۢ���r�_p��~+(�D�O��v*k�2s�X�	Iʪ����$I�]!�jdF�F��U��7j�T��H���(K^��'fg��I���m�VE��r�;�fF�, :�	�86�O�u��s�(�i$ �>{�a��r*E/{�/RE�k#�4%���y���m]�mP\�����Sy_*;��*{i�4�7�gW�Y�	��*�^�N�P&X!>v�]j��zY��<,��G���T�ty� �}OB�T����k8^��gy�Gh��I7��CAs"/
|�������2�{e�nY�ݙ�l���u@	' L7�?
���S� ˥`ױ�Vn�b-�JxƉ�=m�	��Ku�`�*�p�̡��ٽ���{�����Q
�ҽ�.G/�`��s��v�!B�Sn���(i��)��i�3��ʛ����5˲;N:m�]�ۥ��6�2��H��ٔlK
�YDp� H9���s-��Q�'RT���HW������	S��~Q�\jS�0m���؇��M����\��3�R��X$�˖J1N��J����c��0MVwmo���Yk�
m���l4�4AvB��Hm#�����s�|v�	�nc��P�;�د�Fu��|Z��l�V�9p��}.��y����j� V͔2�cO#�I��'h��N��*|PH�A:״���N�O�h$U�����P��6��c.�^99�5�$*;�6�n?<6�vӌ���{L���;q/�Z���`�������l~��+��{�;�o�	��FM�<re:.Ҫd�#S�0��#�\�,9J2��)�y3�����ʥ3��[\
k�mŠ_�BQ���h�3�'��r,�PNٙAW��a����b5�O@��vfP��:鬢���5p����I��A"���1�����M�	2�z`�Pa�S�)*�"̯������c?�����6!e����K[.%M��ց���b�k�%,�?�4@��qL��gBXY�e����1 ��ʽ�.6k���t�Dm��|p	�v=�T���z~�o�2�ϸ����v�9Ҩ�[�	�Jc�b�`��i+����iI~b4�P(ȫ��'��( l69ݽ@�rUA�?*���V&�����>V���������C�����w�g��$Y.�b���'�)O���%l�3-�i
�E~a��"��O�C�K"���e�yT��QE�:��)>{ڷ2�b�B5��k\H�,H�SLL�@��y)��M��0�Q��䖞I���^��=�:����MK6���7����P��|�ʖ�������q��-?L�ڈ� �۸��78�;���r�J�#�;rRM�W�H�w�ʙ{��D�x�.?�h��CDN�EJ�ҝ;Gf��偟�hE��c�x\~������1�}�%���Y��1�������Z��`p;ڭ&7|���U@uR�]����J�q���[� 5Tմ7)��L�}m2:v�OH����*Mn� ݵ:��J9]��+k��oƾҔk�	�n�v!\�I֚�;�H�D�QXΜ3<�f��h~ַ=<͡�@��]�5׳�y1��ꪵ���~�of�A	g�:NN�ɺf.k�[����m�A���Հ�e���,m�m���8�Z�F-���:E����g��f�<zW|�!��7��tRi{;���FU�x�h7������Xj�=�"��-Bm����6{8�aċ(��|U�>G����+ے' ����w��|6C�E��o<��Ӝ�w_x��pX�]�}�q��zS�q�2�dn�J�[_y�/3�L���UIX,qŝ5Y��gw� �{<�jT��Yy��x�Յsͦfc6��1��on9x	�+%A�n���"!ܓ+{�o�<��CJϚ>��ģ�䚹v�t�$��ݏ���FD����*N��D��{.�V����7�ُ���|��-�U)=����|r��d} I��qk949&ϒd�́�c��2�9;W��x����)��{���䨃U)�ҧ�g,�Z��g8CGc�g%E9P}��_�ӈK��j�)td�ٺ�Xx�DxL	�^v�6�
�~�֔K�3q+���3V��-�n^�'��#���&�#�t�\?������C�*�����'\��0Zc-Y�$i����l�5!f}㎜����J0�*ķ����	���S��|¨A�,��]��=�D:P>�.�-$U�j����)��& ;�D�;����>�e!բ�,K�0����fG���ߥxȍ(�G6��l�x�oq�O��:D�-��G^t�1o�����5���%�"�� 	3��qzQ�,A� w�S:���W�+�i!���F�RJ5���εkR}}s��_M�H.ӑ1�����b�VR�y������B/�O���������cc�(�<Y�%L����.������LT&>'ߍK�ݩ���9q�na�O��m��)��9Q��:��ڃ0�5��&s�h�'�@D�(ĕ�6���H�B����T�GUM㿈�J��U°��i�1������T�1�x=��K��Xkwt���Ă�T�Z�]t�f>!����/�Al�0x�Ț�/J��y)D�!P��!#�}X�wgU��`�~�1�mǇ�S�H{���@�=�����G	l/*�=xXf2�Z�$��p�U�e���j����(��4b�l�(Q�A+�)S�4��
d_ �N��<�b!�#.��4q�$�UBx'���g\;[�~��zK��$+k�I^l�C{,����3��H�{i�{��A��B5�U�g�6�%�>YrvPdV�4�����]�d'��Z�Э�
/�����B�Nb��-.��4��[�ا��6. h���d����$W#�š%_�Gn���yQ���"����:���1Ӗh���j,�����F�G}k^G��AFTêw�`���iԂ��ǉ���� u��Aq}^�JIz��.���*�\l%	n����dE@=�w��5�b
�Q pЋ���a���g�?�{#=$F�
@,��WbU��$h !�Hm�X�qj��W�;*>ҍ�u{����bkk��Nݼ~j���{e��-� �Ff�9a;��Y��'�RM�PxH�����a�b��s4����d�o��pN(M�C�X ��Ϡ����{�8V83��
���	1��R����#	GH�Lg�"�m�cI���5o������8�vE�ۨ�^f6����9 ���g����}q��g"�]�Z���)~ʛ�:�(��h'��7Jߦ��NXRFP�<�&�f��Q�{P(���.��bt�����������R8qq5K���^,���»�(���I�M�_���2/c�.9��D��v��{Kn��[h�N=;�)
!���|g�g�R�����MP4�ܬ����W8�M@�Q�h����R��E�G-G�����V�ʲ2"��]��_��̓�-^wA[ES���G�0�4�&~'H��j���y?�(?S�u�C�»e]�����U4�7��&�O:~=�/+ ��T	j ���	��_�~K�x�o�<е��a@��S�n��N=9A�����)�%)�2S :��jE�̤�i{��������}��MH�³���"Q��;d� �~!@F�nTr4�
�h�Ѿ
VC��^mf�]�� g���'P��V�$L��.�����T��w���7����a��╾�C��Hf�,0g���Do��f"���5M~A��jXA�Q��
�	�x(��u�%�}l�;$�»�G��{1��&E��5_�u�JL,�PG������>}���9��0�W<MK.�+ȩ{
�-%�D�T
��'���a�9n��j덏�aI��6�"[��J-�k�g��+-M9D�c�k�&�R��6�WX�w�Pi���S&���
p��0�k%�;�v2Y~!���Պ�g홪2r� ��B�^��
L��0g#��Zu� 60�!����B�$@ k��'Y�8X���Km�O�jc�7��ehY�j1 f�5���&"�%"��:S}��������E��:�Ӵܤ��x�>ͣ�d�Uq7��Q�����{��0k�.+Km\3���c�}F��i�3B�窸̶q?�����4nЈ�V����M]�s��,�?S�x^��SQ�v_a�3����+����b�0��FerJ������8�̆ �����A���t�T��Y-Ӆ7ﲉ�<���x��-kC�;��F懩9�rY\�ڙ�6��������.�s���B6�@Y���h�J����9��gΆ�qFjV���i�͌b�/�ɿ^*��kA!q�5uE�ko���@��u�g6u�5#v�ʧD��C���xD�����(-���WŌEP�����d+>1�R�������=�3�0�j{�\|�E\ LU����p���P�l����h[D�Q><��/ j��ݎ�6R�#]"�x���^�B��.��&�3h�� ��������w6VC�������]S����/p�ss�p��T���H�k����j�d��̢Q	z&H�x�䥲�P�=�>x���o�P�=�Y�0N&;&:L!��������T٤�����ڮ��e��*�D��Т<���E�	I�E������(~��q�H�Q[^Ծޯ�9�ZJ&a[��Q�n�x�mE����-��P�"�
##�Gf@
'_Yu��?5Z�G0>C��'�Y�g�輝hN����	O�[;HT��B�YgJ�H�-.�w��1n�v���p�|�R�{v$�Nz��'s��0QuuZ ת�u�R� -��D������D��#����t{o\Z���o�T9M�sg?�J�</e~�����٬U��)���t L�o�A_B^`�5�~�&WI��Wl��/����X';\i"B�h;�qj�!�d)�I����]b �X<7�[y[�f�+t�ހ~��!�;3��mY���j9���H�j�<��9m�4'@F{Ѹ< �P
�3�"2,�z��U��܆]qdU=�B���l�A�U���27c��dA:>Q��J?�Ͱ�Fގ��n+x ��dv֮�O�=Xj`9P����͢EgM����cFY{_�Η0Fd[�\8�u�����Eo����BP��p��{���4����cn���<��{2!�����;]#��̏�~�a&Óԓ=�\��*���5g���oo�룙+d=k����c�[<��,�ѧ�Ki�a��ٗ��*�������]��g����%K��J���/�Q�=�߈���.�jL�J�;����Y�3� U�̬:+�岄���*O�_z�HMC��5�P�s�[jf��.c��&����	�c�8��_��N��ղE_ �j�1�����K�f�,S�}|�����555����W|F�Y���Tm��#�f܁�2J[$ɿfK���ฝx�]����(o�˄7�]Ǿ��[�Ճ�DҀb���,W8'������� ��uk�X %.�ސ�EӒ�{Ѧ� [\���@F��N�e�|H(�WmY�q���;G�MNY��"����V
MĪ�IJ���
o���h����Q��t�*�:km�a�0�\j��3�sTW�݊���L�T.4 g�1xx��$�N)���Y9\ŲV��|3f�_BJUS�"���� Y1~��jEe? �m7�Q��6VTͯ7`-�MF�!���z��L��cvfI�t��?�A��3��`��蕪��^y\U����?vo���&|�h��[|�
�~cU 3��vp��щ�Qfm�kw0� ��&�Im]�m���/h=+A~�ˮDg��8x��ZҪU��1Lh�7����ݢ���G�6{V'U*x��i;R���GI�B�7�5d���CO�݌��Y�ʱT0��ø+��!\-M?`k�{��i���%^|׋,�}s�:��U��$uA�f�x)k+d�!zy���a%:{��b��j��Eh$!��J�Q��3̪V��x)Z���pt��3�Ğ�b��¯��}�������d���g�j��Ð}жv�jsn�o��R���)��?��r.�i�qF�2��@�K����{g�#��<�������y(n�����ý��}4��sѱ�i��~Q�д��qFО\�J]�;�νnv-����F��� ��{�B�^'sQ��i��e�z̭	.�A�R,>�EB{H����D_0�\�J��>��|D���0Ћ#0���@�i�[c�|�x�iϧ��Rj��v���|��V2��(�n`L3u�T �6{�{WT�(��cӕ�u�很�P�G�XG�ݜ�,�ob�4n�x����લ��B�8Dw݌�&��m����֕�u�����k�8SM�pg�]#�옽��R��p��=�~������8V�d4��\��T�'d���i�|�p��A�S�c!�#xb��gW.r��[�ŠzY�a��<.00Ҁ+a�ʹ���m�l.��ȯsEvkِQt�i�@Yt����
�o�޾���{ץfЄ%�v��th[e�d�X��L!�Rt;x��[٦y.��p�hI���x����"]ei#8L|e,%9������q(nZ���4vl��a���p�*H�k/��y�xܱ��͂Y��re�� ���5%l��˷���w�Ȁ�Z�|�5�����K6���TY�C~jejQ����3�G38c�)�A� Dt������z���l�}k�M�N���	.��K��밞|���OM�^�X)��A��ȅ��0u#�ᦋh�B���!:ϊ��z�io�B6χ6H�C���NtB���\��d�#��*z 7���AA�w&�(���n�RyC8�Lll@��И�	!��ܮVC~QA羚]�蘡z��h��qZSBs�>S��Y�I��$��׹p\�e�=%4pI0_9C9�k�W�];@�<鲆��v�Ac��7�m�Ԥ��. �No��Es�d�%�;o�̽�,>.����`��<^6F��&���}�eZ������/�����)E*_c:�s��"��9y&h6��!8_�(�GC�2��3�u���Wȕ����Ws[�nc���Ͼ��Kb����;se�� M<��0���yH�ް~�s�j��yg�ȺdH��7.n�M���h�먏^���B�Z*my@�f��"�8�x��l�S<���R'�!�a-�=��|��=��p7&� �t-HVp�ARy�m����7B�^-z��D��w��YY��a�����\��ϱ���Pb��?(��`���Аi���6yjQ/(ϫ+(&bhj����&���yF��=d~��~&��җC
�mB�[Xv�t��չ�=l�q�rk�qY,P�!/�e�ёm�m�K4/oh�q��}xE�Ω!  IT���}�ՠ@��S��]��bZ��v$1���}[$Cg�e�����G��:�~���B�w?���C���o����e����;�v��m�$S�F]W���F�����l]�XZ�ڮ���C ��RC:e����[RNT"<�����K�0&dY�?eu1J4���=��=X��=�ғ����XːL�$������F���c0%���6?ʣ
�)�.�_�K �_��C���>�|�P���1$Ù��y��Z�:Up��׆x���T����U�ޮ����i� �N��~oZO�IE^͋�&���������k����(p�®S�ݾ|I
�IG���}}�w����?"/Uܼx��9�oD�w;��K��qH�|������DK(gE����(j��_��H�l����c`#<3l�N	�t�$�{���~�x�Os���dX=�lrGJ��1X=dk�{�3�cc�~\�Ȥ $�-_�h$3�X��v�T��P��6)����2�ƚA�g]�F�7�"Ѧ5�Eƞr�H����7������L�Yx�#�8e�:D��3���t$EX�[K�œl�-t���A��d}a+ֿ���5ލ���~Py6a����c'�@��Q�ߘf*ͣz�a.o�;S�2�:��H�~�%^�Y��BU�h�e�L5��w�$&��ΫPP^d�>����"����Tt�_��đe��J��,k�1���5ڂ�c��Ϭ�`�3fAv57_@7�)�ψќ5��DX��=!6i1떂������2�"�{�(����r���n Q��ɇnd�F���z�g:d��GeiH�%]�t�l8���R4s\��\��S�`���������{��30�n�!k�s*� ���L�AZ::�HY�)��[�k�(��3���]>5P)�ˎ���1�v�p_��#-j�P��'X��zW���xW[v�nq7��V�䈦5��5��bX@���� [^���a�Lю����HF��ʿyU߱*���M/ҠR�t�S�F��nhl����Bp�����<���y�-A��Y�V4�K��+90�s���(F�L��vDۯ45���R�pD/?[4x0PUٺ�7k�9 A��3�̉0:����M��_�O&���B1P0)���t�}�����2�A��8e�OY��O��,_'l���|V	,��ٸV��C�5�_� $6��=ޙq<��A7�4��лn�8�}����p�r�$)R� ��G�v~���L�Rt5~�S�&�Ŭ�r
����VMI�?�K=��Aռ����QB�:�q��^�[d��́<�q��Y]����8��Jt�40��R��wrz���yKe�Pأ�j߄=���}yVft��&-�X��M�m�;���>)fw�4B�d_�Xr�������j1H��Cڗ�0?���H�u�o��ˋ�H�o��F2h� �]��O��!�?5�*$7���:x)G�������<V��v�9xǺݬ�r}Xh�Ɵ����rk��Q���8_��m������������(���=�V�'qz�oOK�:�������S�z��å��Goax4�`����I�V��,���/}�*#?�1u0���^5��&�b5��� )�������/�#�t��{���wV���v0؏ckX�y�=�ul�5��$*�f��:�����4z�znc
��?�(�Q놝�F9*�Z���	f���&��y���O3	,৖?����d}WI�,��S���t(Ǌy�����Ya����r��{rXs����,��(R�,-F�#:���M�֫� ��2���KR��=�R.fa�vE�ĲC��&P�\0�\(0Z��9C�&e��Kǌ���	�ıP|��°+��F4��H>I|qݥr"	�\���laW�P\�l-Jz^���
�I���+�,k��b�洢j�ض�:�N3��iſ�w�Y��+���#7w&�&�F���YA��`lܼ�Ow���G���'�?�Dh#���;�6
�������$v(2�>���[[!>;�,��ZE����#�(Nӥ��E �9�u�1[*�����>ۄ��4F��P�l|���C�2����p�:�[����
��
�u��"֒n��{�@�	�.�����4P�	�fHA��n�%{��HՑԐ���QF�>"HD��yԔ��(X�� ���h��[�?��2�����A[��r�]J�+<k�
>�}_N��=.���o!���u)�O��֜�'��~t���&��o�g%,�hk�8�ٺ8�;�3�P�O�W���4�/��N���ē�@a��S!w�(���^�ɲ����*N�r���1=?0��J��(W7��Mo�S�yh#@j�Q_�G�n���1����*���B8����B)Y|�>~������^1N�P���7���O�~��9��`Ԥ�4���;i��Č'I�$.��(o\n��`�.��?֔�9�l��1H	M������@9�BA�]@(}'�(ѯ��TCf���e`�å��x��k
�������$/�:5!�vQ��0�1�����]����؅���אt/ZG�����Id)�+�SU���&G,�j��C�wQ��oO�h��f�Jr�Z�9ًz������&���6o��c���PJe�(��8R@K�q�"(x)u��G�Jq��|C��g��֣+�釪��b��oن��j�Yo��7����T5H�P��k�%�7�l��i�ٲ�"�]��[0Y��ƫ���\~��}/(-R�38yi+j�`5���W��d\�Ik��M�E�'т���N�+��L5��������C�_��w���B�h���`���s�PC,o�	*��d�S�v
i V�"�?Ʉ&�I��3��:�H"��T��CoK�p��p~Mi�w���<M:��:��D�=��C��B�$=�����S�� -RS��3�*��:[h��ni�ay�� Y	�"�Nv\[�߄޹uM�)��1�[�X�}�ڛ�D�U0<@�� Ѽq �:��M��@{�u�s$*qAk���vW��\s���(�H�MA'�񰬤�I�{<������5|_ �� �ѰE��:�&qP��ձgH�i�2����E�ޤ�D.=Ҥ��*�<����\�$ku��S���vűQ��p�������{���p�T�y?]�AXy>7�WU�/���W��&�|�f��ln�/�F�PV'��VU�R!�q�`��v�0žy'<RE��7�N�j�\��)N�LЊy~�8�+�T1�1xڅg@5��/d�m#<�����)h�}ᑬJV<*��{wn��9���e��C���#Y<���E��\Qe��(�E�ؽ�}�T�i�'�75tz,+�?IiܳA�v�`Pi����3�.�p+H��U���-zb�?
�F�TR��p�Hf9ض�N�L�I$sG��y��G��f�5�ω����Q��pV�[Gr4� �B�I�1o�*���"��T~�Gi
tK'���p�*�t�]�d	�hM�km,�z��=i���Ϩ���;l3��M/~,ӡ�h�E1�m&�)]fP[��p8��őӒ���ǖ�N.� ��6[?Ӝ h�M�G�-�o�`��n�T���qƅ�U0xRPf�'�
a-\{��hM�Q=�r��)��L7�v�a��b@_��2���a�G��+s��Ԗ�^k���VkS�|u[ط �-n����'�
jxHU��&���
Qz�k%��o�H|�_/�앇x
�^/O�c:.|C����%v	֤͠e��Sпs�@g�$�I�n������+��;{���&:ѽzg�����2@���C����5c$nY7�Ձ4J-F퀝��}v�L���J��vjH�Ǻ���6� ̩T�Oi��w(^wT�$9'UǸ��B�������e��������WĨ�|P��,�df)v��l=�Fg�3�)6��
t�'C�̘1}yR9��28� ���LJudQ�ք�H2��;�A��g`��ָ--�|0�V%�� ˢ!�I��t�c��h���uP���=�
,n^� �]`^���2O�#8��}�iS�)���ƥ�KY�C���%Mh���%^_HM����d$A%K����N��M�mF~OT���ܰI��o�_�ݱݽɹ��<{=�G8�] R<�i���+ȣ>=����1�8� �����hk��?\i{ڒ�=��W� �+
Qk��"�1��{����<��Q���)Ҙ1��1��\�:��;`^��hC������R�y�0��"�z*ύR�Sͥ�k^��n�(�G  F^Bi3-���J,�P��fp��-AH'ϔtg
�@�D�����P堟��u��,�	��ZA[��,�ʂ��#��xՅ�.�>*�tEG߾@G�m.���g�f�jjV��+��dO4]��-��akl�<v��ax�e��^���%��ԋ�R[���Ŭu��H��r�V�Q'�i�eLuvd���p8�W&�t�����B?T	��<�2���-��e�L1R�B�럈�!~--��M����!�?gA�Q�^=���S[	�K��H&�3����7���~Px}�����ͽ�0�)������WCЃ�hi🏽�k��q��"|�8�*ȅ�w[�Wu�'����dV\��^H(S(�ɔ��|FP�~����!�b
��+/I�W�_���y����5mt���Eǜ^ӧ̵[;㼄������<�����%�i����/�g����X���i?���D�ȗ����ya	OH���_���R�%�F_|�TE5�"�j��n��TaU�(�y��u�@vi�gx�$\���\=�qFo��:gYpCM���]&nr�ި�4wz����\�'=K���l�5��6)�.{�ɤ�&���ߣ�	�'>65�裌'�����6�tKh1��JU�Js�];���������by�
�ڇ{q&ߧ�M��F�ϋ�_E��?�W[9�^��o0F{�Q,�a��N����Ge7�@$dݴ%{�N�R�O�<�K�(�u��c�}�Af��˗��G�?�b�����l���#�B�ˮ�蹪����kt�r�D��˺�g'�'�3H��moJ��A	�RE�'��D�ib���40��1���(��V�Wї4$��e���%U����?�;J@���p	_�d֕�b��=�$��Kj���ͥ���fG:i��TߺO�Ai��a����f2�泧5�*��7�|��S�L�H�u���J9W�>����V�z�`R��c��m�̄�p)���l-_����oT�DQ��r���/J$��g80Ԯ��p��hf�����ap����CEş�Z���G;�'�w}��g��K�D�2�IoW R���k�U�%��|[�0��n��ُ)p�g���{�1&8�!�R�v:!r�A�2&u8N�X=�����R����Z�D*��Kgw��Z�[c$�6cӛ6܁H���`�(���y`"R�n�ړG��(%Ѫ~�ǣ�X�U]gQM4����u������
����}�+-�YR���QȊ�<��M�q~�i`&�	p��皈�����¦I����\=[ǚ��� ��t�+W�E3 7�b��\�Mw{_����H��P�R�����"2^�!{�lWk�щ�ݧ�
�q���1<_n� ��Mi}�Ѵ�r�L�ȝ)��EI���+(0=Q����p�ga���a�|��a�ooCZ)�k��/&/{w
,��7A�J���̾��C���7����I���	�B�[X=7�����G虵���'�����1�$�J"j�����㣇nV m�C��9�8a���tj/#Z��@�6i����b�!g�3}I"��ޚfW:3��M�Y�N�����^?�ƃJf��F����L:�mb������d,e�6�|�e�w̋v���O�a���պ��\�U\}���JT���P"8薃��ɐd�p-)VqiR��W%(��1����j݅�e/����Z:I9.���y7�֛�u�V�>C���ٚ���@���S
qQ�O�ʀ����z�x����E���Y�^ߙ�v��pFЫ��
��Zb1)��Zޛ �(3P�lu��~��G2P�8��U&�z~Z�;I�JX7Kd���A��G)�4l]0�{h/�Wx稩������tX�V�:=>j1�5���ٮW��~���h��	��Ǉ �2h��8-5���
Wת���4$�Q��m�#��[z�Py��������][D�{˵p��.RꊔSt����	�qkf�����M������5�`�~&j><Z��:��@Uaj���v�o���XD��
�Nn���l���*�����KA���B��֜���^��9q�m�Ǉf(��()0�W�_4�������VWII_4Kv`��~���]+bP���{���r\Ő��S��Y<V0$ �#T���w
�w|�C���gV���l}�n�� ��@�Z�@��_���-6j�˦�3��)=�+�nk*K���]��A�n�q�ñA������O��Y��Y����ڹ�˶L�����N�o`��5��%����|]n�8���F��˝�k�}��u%C������<!|��l��N�qؕN�\R;�h�5��ς4�^Z���L4Jb�}�B����>���ܻ4����
����*�;�G�7km8i�(�}�Na0f�N2|�����r$]u+r׸AaŪZ�������@2Pr*w�t��g�]�Y�B3.���I,�r�i�J�(0�ϯ�"�,�.��Z4��9={��4�w������	X�!���#7�Z��~S��G����9-q���!9n��~���1���b&��+k���^Z�s:	�t�?4g�k"\ek
�F7���*���tlM��#�4{�?�����s�<������Yl�a�o�ڕR��IR�����J���e�u܀�l�L��m�G��8*�ٙv�L����
����S�W.���o,�4�ĭ���c���x`.��l	=\�2gL��^K�h�<��d�v_��޴�z6�3����"0���/�F,�T����(W%X����k��|aHr7�N��[.��&�1��GkI�]un:�u��s�u��*��iΏ��6�h-8�FH"GX �l��o�闿���	��Ǭ� Ig�����t�_d�7�����xC� �v��	4i�����Mf�S� ��dh���%��a� 
��L�Sc��Z��nQ�e�� �
@��e�-ۻ��It����29��=����]e:��Yn�xn���~�����J��H/�+��AX��)y��.쁬�G>��"<�6�Ӽ�ک�Ք#�BVL���ܼ;��\�(Iz�^�V{��j����bV�(��/�uo���Y{'����1�J��~�|�E[T��hR�\����~:���cB��e����/� ��Y�w��[��ڿ��!ln4��{Ҡ��i��S�$�:�"r���v7��3�T�R�-[����L�|�ǈ��N
�gY-��{N��%@d�b"_i�������m+1{#�rn�Pc�8qq���\ܾ��X	^�ϓ���ALQ>�N�c�!�,��囥�%�Itgd~�}/>�}����`���;ҋ�̖�y�rnJB ��< c���i	����ƯH�I�e`&�j�+Ǿ]� �N'��0�9�k����h�nI&s���ePZ���^��^�w�y���V�u�?nx��g���%�+r��i�(H�0\1L!G���ϯqw���B[����#{c���{ԡ����)	kz�� �"���@4'�~�E"�}GOȀ(��D�q=h�W�\}3�os��>��(t ���`Z�sj���⿀Kry�l�慌�E9M�ً^J��ۑ�^9�>�nפ�>�b��eb�׮Xs�~�+&�	�K����矱������E��e�⁜W������g�斆
)��=��8��Ic����N(w4(f�D��P�k��ʑħ����g�#eг���+�v��j~u?��.������=&W�߹�_��Qp.��{bo��LA�����a���!���������R�3x.��QM�?�n��ٰJ�V��YFk��ƴ������HII:�[PB�ȧ��*��3�i5�ZH�����`w`e�8Ζ��6y��o��o���0ۦ<��Ɔy<%���α��79�x�O B'S����Gɮ-_l���ړ+�h7*�z{�����G�X	|�b6��T�d�?ϐ^���R�欷9
���U*R���ofV��M�����Y��X�M$��J�(�癃��z�!�%��d)Ŭ�CR�w%ӽ�$G�����͡��m��C�b=��0~)��	�ɋL��S��R�V'���?
�D�dt����2f���5��q�����?�ۇ�1W^/��b�Ax��1�T���d�e�E�~��h����ߚ�y,y�>a��P�dz�\�[�VW�n��!�wb��PRB���0$n�y�kqR�/�Xax.'�<X����qJ�'��������� �I�jYKv�a�K\(��ޫ�'l��G�`d��7�H>�C�a�_�i;1�C��9 �Ks���ׄ2?���ELC6�;�]D�b��&]�Q'=�/�nj���+�<��ESLϤ�O�]3B�Y�g^$�=���5��2��*��r�k%�:�	AO�[0@Q4-�ܴr ��:�_��6��y�f��C�>,O0�|/����x�jB�pa��2���'�#��(�u�2�Q���������F.����'��8�a9]��Bߤ������Gs��]�e�/N]P8�au�Q�B^N�v���}�����u�� <�ef:�C�NIG����x���ɳS@��/�#����Z��|%�ս%��q�B���m{��5@=P�A�2'j������]2��5W��eXٟ�����t�@��i��wJݺA��"�e=?��@L�A�n��p�_�[��K��?�atk��q�̜�G�˙ݽ`B�v~�1#��|t}XV����f,,w�w!�zm�L�Ϋ��*q>�*蚮O���,�l�ʥ �B�R�$���b�Y�T���6���j�h��9O�puć��		�U��&�Uk����]�������8\��Uz-�����*�3C�����2�?O��zfh�H���=��v�1��
􇛰��8��ѻ����2&�|\�r�o��U��1S��0F�mő~�m@`��g[s��.~�C�x�m���F?�˄Jqb���T���r���-C��R�u���u�#����_߬&�1�.�S��ò��
����y�k�[�!��m*K�05�r����yIwCi�E��z���	�ͥ�1m���>��t�W����C=KiJ�}J�ؖ��*A��t��c.��;���:��7�'��7���*��>e����R�f`��?�B��6�b�#�,��n�ͻ�{Q�ԋ�̖����N�
}��#����up�{���W���{B���l\����R� %���FG��`$rZ�9T`��Z�j[O����܈��u�3���GB���IU�-�L6c�ΑS:�(�,q��ax�6�6�`!�^D�ʣ�8ݽ�2��{��y�[+)��P��#ݵ���6K�K�$'��ù|1�al��Kc�ϗ�e����$���l+kp��,�`�a]�Brȉs/n6��ln���Q�Jհo��G+C?�#��8�����&0�W�%B�/��>�}��M��sE���#��3����t��Ь�P�wr���61���0c0n��1?�oa+
N��g[kq�󞻧�Zװ�G��Kj���j���'�9^�5$�����.G���DL셿�W����զ����D;5�?<��[��$#�@a��ɭ���d�U�Sm��ۚ��4fQ����:3�YV��m+�DDY���vQ�c޾<�՚�?�H�@��7���oZ_CCͣ�x��N����o�$�0(��c�tfAoŶl�l��l�ג�h�,"�?��ɍUu0���K@����/P��2��?�H�1�,V�{����v���ؾ{�W�:�M���˓j��#!�^��g�_�H� l�z�!����^�콐Z��̪���K��XR��tj��j5��Y���G�o�~�7 ��;< *ψ�I����8�|��Z���e��v%��}��	)é� s�j皵���5ܚk�,�����9���G�vqX�M�F��R	U5M���U���stXH�T��g@��[2K���ҀAe����ہ?�[[��YŠ�'����t�7E����$�`~`[����W/��;oy}�)6N��{;���h��5[o�̅/��붢�#�������(�����<�H��h3��Е`�Z�_"J�!�*���w&P�x�˞�T4�9s��Q�'!��?SV(�-_/ˍ��灈��l�7+�,�UL�1jg��G�:��0�r�ؠ�ɿ���W�'��O���mqY}��"���z�u�@R��\�ʹJ#;�B�M��WJ��kc��_�#�=�&�>���6i���$Q/{Ϗ��K�@�]���6��]#��b�*'m7(,h)j�*�o��.�l%�+A̻7��C��[�H��3a�`3[x<4k�2�/��X�U6CG9أ�k<�������DΡ#����M��;���M���� ^y�sy��A�PUx'y_���*�9�n쩬����q���CQLjZ=�QQ�{�[2M��3� eT;�{�����_&�[O�������{%��n"�(I�.��kY8�ڧ���0��гU��;�A�V�hF��m�qI\����p�^{�k�sj��'f��'�5�n8��b�M����oT܍À_7����~o��ƫ�r�����L|J�#:!��&KW�^������7f[m=k��c��b��]B����4��a*���^i��L�pJ�N���ě۪�B��?� m	}����v�S��<�Y(t9����oq6&[��/�P�4�Zl���Oʹ05e6+  �C j�Y�ݿ���/��|�����<� Z��K+5���U�M}�E�C���j,�e��9-���D�����z�JG��Mr�QȜ�_na��p�ȥ�N��\O�
���])V;5,B~��Q/��H0:�Qׇ��r��$���d!S\�~���	���F��|�
Z��� �T/�gL0f����cT��)�����Z��u)�NWs.0�Do�$j�L#f�C���`���Ľ��d�6# +�D�S�D-{��ՑR�|;i���p�3;�'
nE���+	�H�)�3[�C�����^��?�����A�s��s�>�>�O�Q��ǉַ�~+>/���ǂZ����P0���N�����en�\�W=�w��#�t�/���C._k�)BY:��S���`��a�X2��]ʪ��BIA�2�7�9���a����v�����
���}�Q�d���H��7���*}6�����E�:1��������}Y6
-�|C�#+5�rlǠ�,�o�cs�^�P�:a�D����� 7�o]^�tn�''��E��Pl&f��� �I���=��p���-jr��_=�"6x�h� �g*_kV�m$4-f�y�'�:YQ�-7�(����32��_:�kp�ܟwIx���� �Ǜ���2 �Y�3a���( С:�/��0�&�	ٵ�a�]ߪ���t�=�yRN'�n��0����*���/}�<cX"����c��ů���>�)".����E`��{p�ϙ�dչOɁAzd��O�3�I��!�z�������D���|y��,��	Ҕ�}Y�c��٢�@*U8?UK�����GNu�"�m���an��Q+�m4�# ���t�w��*Nv¤�YF�O���BѰ}��[0��3-���iQ&�8eK��XgG�ƕeY�D�9[����*�(���2g��^	F1��qb}�������%n�_��8g�G붜�S3M\TG��NT��k�a;8/�E�ĊT���0�V�.Ur-����/U=���΄��I����;���^�p��L�� ]�,Sdځ*�`�B[K��AQ8�aakr���-:"=�����x]�^�&����	XI9�4(=t��(��PZe��I�~��l� ��A�-�ݢa��y�Y��j�!�76��w����_,�R��p��d��%ĸl:�	�u��h�s������>D�SJ蝟}�fN���	��6�����=�V���`�* 9,,�\�)M�	�lͣi��rN�}`����]ү�CM]�j��+�8�����@�[ج�=�MS�D#vB�I�B�v�+�ׅ�-saѷ6m���?�6���Y��$!�\D�K#���D�,��v���[�^Έ9����FI<����m����)���?>���}SK��4�x�
�>���Ҿ7r	x�&��l�q�j  �v�S=�k����mL��|��o.���P��uY#Rh����*O���i��0`XS�� �S!�������4qG
BnJ�B��t��gǬ|o$����/�`��:>0ݟ�w�Ш��f�ߎ��M��3ϊ��������u /��{2��A�&:���M�r����ȧ�����kkd�9��y��ې��HA�P?��_�s�i��\'�aC�)p��m�E��k��OW
�Uڃ�_�K�)�3�S�;�ȫ`D�N.8�tánw� w@����0��o�c%{$yxU5q�g{x�M�1?$'�_����/K�	W<P�{�|L��0�����$� 4�k�θ��c
��N��b�C��g�oYr���D��l��2�����3#�H~۷þ%�ǳú�<�O�e��	SyN��7�6l����s��������i�Թiݗ�	]����<vO�ڢ�!�
��-~�L�H 	�H<� �؆� DuL�8t��c��D�5�vY3�uH��/�z;���:j9�ؠ�r��c���{��v_����G�	ַX�G@J���L�����X((���EcI�P�շ�i0.C�od�D�����{�n��� �v'/����,��tCf9����g1�-�1��D�Y��mA�P���w2fx�!����wT
��L����>$̤�X]> �Giut�X@�yy|*b*���/Y9-Hy��K�_b3s&�`ȶ�)��M)����!�n�ẋ��Z8�GJ��`�6QY;@�}Ǧ��	��|n�K����H�v�1�S��J���h�b�Rҷ8��	\�D7������g!��DIVt|�M����|ds�~8�QG��RU$�})*��K���
��J��[r̼.�j�ʪ��]�e����Sa�(Rx�g���͢	H
�$��tEo(+�����`O>be�y�'�#����X�ɳ�_4M=ۣ$7�7Pn�9�li ���RЃ
D�jm��Ǆ�_����}B��[���"^8/��:�P�����ө���g9T��g����_�����x�z*��yM��f���"J���.�����,Ƌ��J�Us�}r�����p�~ ��M֔)�s_|�`Uj��c�}4��!dM �Y�.�}F�����t�삩-Sa�B�`#�Ш����\-��!h�a�"�����+����P��ͼK���jwg�(^���f��K�C�������Ph7�6L�joe���5�D�$��3:��o�(R"�d5D�&J�-1�88Z�U�'��Ұ(CC����X ���j'����	r���謱�v��<��c�<b�5�+9wH����
1ia��Im�RJB��O��vY^���<��ޟ��ݣRb��]���G�c�x�Md�<�\�wn�1�=0|n���̀f��a��3cMs�7����p�9O����2M&A���*.��C� 1�ǐ��a.�|�X%�x<,���s\���m҇� �Ow�b���D�OH] �8ߐv̶P���R�����͆~��X����X�����dQnF��"��lS�����QM���R�w�`~-��[�jl5z��H�j"t����-�c��؀ӡ��f���u���6���I�4�e}8w+i�Ib��$ܨ��O�$
+9N\��(:@;�V�i�C��Ww�Kc9n఼��i C캸14��q4��2��ՅHd������A�٩,����	G���;_�!:���i��R(;L��	fm��ͶA�3̞Pp�x�L��sK%|g �pOo��ۄ̭��Zi��|�NbN(������N�M{����H)���#F`"���;#0׷�9�5yU� l��n����r��y�:�$��4�h�����F8�N OP�2\��q+�P8��φ�����>mL:#��|��(����k}_������.o-�C�(�*e?�Og�����(*�e�bs0�O�⨆>��1��$=�-�{�q,B$|J����S ؾՋ���B���TX�":���t&B�ը9w��S��3jBP�S�hѧϿ�:�<��)j�gk?�\����n�H�_dSB���C#�W��j#Z4�1"���tc���Z���:M#t>�,*�6��`��U 'Z����,/.���Ȁ��b�Ԫ��-<�2]f����h��ь��լ>�Nz��g�M��6��6��<�j9���q�ӸONj�n �3��KJ�RQ2�_p�)�����K�n�ަ� ����鳘n�Ld�CWD$#-�-�{-��^��f#`�\1p�p���NFW�`�TE�f]'����y��?:�t�N�j)�[B;��{�y�4q?�-O7=�߶(}9�'*�����a;4�5�SX���DI�'�91>�e*��	B�\3x�a�9��dh6��P��A�����J;�5R�e���24�M7FuQke����8U.F,d����q�')xX��j������v.vP-�b��i`�~yg���oٌ}%���}�֚����i:.'�x[0D��XJ��}��wb��ĿgA|庸�X�S�$Hݜ|��x�����,�^�¼vE�7��6�����pq��5u�A��9fی=,h	�����9g[�,^,��X�Z�kO����*j;Z����Z52����_� t�#OM6QC�ؠ�X3�1�:����G�*����|Os��D!�~$0@l�8�+=IZ���>ͅ(�:�|j��h�#�Η�,a~�'�N��ܛT���B*\+�0y��U�m�x���EF�	�ϥj2����D�1�$:�PDu�O"�o֘M�]x�A ^q��m)��򏖖�Аr_ª���gy��~��(���3�f��K�&C�|1Aj~8�zb����>0r8ot'�������$쭄�B :	��R���)0D,�V��M�ꝧ�<�*����mb��ۣff�G��B���R:@�C�V���WJ#/VO�N�/$�ի'��H�͉�eW��D�k���JV������.4��# E(^�ޠKx���o���`�TDC��},��OܫR�bAO��"��������Vͽ��p��!����s[ߓ�ip��I{w���I�A�Ē�IL��ؼ���8Q���\��w�|�g��|�<��L�w�B|Ox�:�v�2�R�(>@=�FP8�a�6��n���Q�`3�z9�^�B��c*���߁}�y��I����j&��L�/77o����lP 5t-.��mx����>����5u�,ڕD��_T�U�ۑ'BN��,�7�� f�:��#
f���7����Y`���dզ�����)h
6ߤ��$��VJ��V0K��_��#�V�>�e6��NC�\I��Hk6�'��M�����T���SM�Vq�p3pS��sS"q,g>_�Yd���&V��l����	�s4�&!������!)�ƒ5��:w#Bò���\ܿ��ڌ�]Rk��:-6���N�j�\{ڷw���[kF�FHڭS^�V��YW���y>o����%˺,u�C�*;��9V=9�Č����I��=�v�.��ȁs��W�'~Y�b�MK��4���:+���G�e��A��H��#�<c�1H�������P܆S��{�D��(f���wcA���ӗ7��)�=x3NhW8�vg��j�.6;� �"�&զ��XMW#:�����ȱ,��u�/�|�fv�7� �ق@8T9���	2 �k�6�xpl�����d���v��n��b�!�ֳI��O�l���.ڝ���E����7�f!P��M�a�1��l�FM]~�����|�=b����ז�T���h<t��+^��"��?]5���n��]-���5�`J�K�jC�i�^1w�'�:\$h�v|>Ԇ�2�|d<E�ѬȰ��CG=��`���?��j�BovWษ4w��=�>m+Q/���(���VK+�a�ꉅ�t'�I�8U%��~#ZD6��!�`�3p�U��v�?�D��ӈy� ���G{�$7�C��ʸ�_D݋���v���b��ߟ���\]7�gYS�!�q�cCj�OA�cmOjHMg֢�c7�o�0d�`�+���B����d2k��G����E��Y���6�Ef;��(��܃z�S3�7�/<��D��9�v�-����7hMA�p�J�����3��!����+��_�`�M�!1b�^�3���gG+�$�WP}�Ӊ�⢊B{�Y($s��0�!�;�/�*��'��W��֖(���d������X��{����H4�X6v��!_���8��΀v�Κ^�0:�a�&�����Q��6�+"#"��^:Z�_�es[��Y\�{H�j����V��DG��0|G�헴��������	�i�mL��m:2����KU��߫�j�X��냪O��풓����L�����m�� ^8��g'g������ڳ6��YѠuOP�?���P�j8�F*Fv�L�/y�|Ҁ�W�e.�mė�ȸ��y(v����z� pJ��#�;�,C��~߳�P�g��Ēq��o���Z�iJк,�#7Y߳_5���Ɣ��O�u�l�½��(����
+Z���نm�����}'�9H��jy�F�Ϥ���MZ]!��r������rl����v�|���V>�9:�:��H��<63( ��S�ʷu`r����C��ag�-S�3� j.\�˴�ZeC�yn�]�(��&=ak����~D_�E��(W��N�Xv8��.�9�W�TFI�{�@=��+jI��@�g��%���O�|"���>�`ၪA��D�C�&���v�~�7�����j�P�K@��٧�����~l�>�UT ��C�A0�+yQ���=����vP���DLcE�gT��������R�G.5�t�#��I��iD����~73�C۶�����rĊ�R o�GDx��rX�E��{�a6[�>Z���X^�g{��Z|�"�ݖ*��s{��	Ϯ��~WO�Cw� ��24rz�09j���.�J�"�a?�6{�|ч?�E5���6 Ɨ�@e���P�:�@��V���ԗ��OM9+��0�f6���^�p�D����������ۑ��.��h���|����S�F�ۢ�%b��o��}8�#�Ѱ	��`\fMe�ȶ�]-DT>�eso����ô�T�C����y�e�N���Mj�Sj�P�Bh��2��a��2n�ע�[��i�AD��yˇ���dj%�]�	F׉L\j�&B���oo�rp�8�hE�л3�4�Y��Ǔj&�D�К��9)Oas�^�Г�o'��8)[f�mMr�
\L�����/%%�����4%Wo��StjX�K����T"�j:0�9�92=�$��Z�-EҰ�3��qI�*T��	�e_�b�%���B��ex @�el'�5�?RS�z�Ym!�"@���T��Tԑ���`[�ѷ�����M�������O�2�q�Qa�fUE�nyJ�EiP �J������i8���Lf򵍗����z ��?�Zƿ��b��
�C{y���ZI�d����i����"��fS�:�!�G�p:�@"�hq��8��_@
�i�7?vBeu�ۡ����v���ۚMig��7��(�C�o�#��2�z\�H#�yi�g�X%o�O�$·U�D��N.yD��	B�3i<�ZYfgO��޲�Y�λ�[�j����y,��Y3o�Y�O:���x5���y�:����"'_�\������VI�~Q�G1T�X��B�J��M>���0�!��'�IĨ��Y�̤�IA�=�BA����4u���$`O7��CL=�dws���g���L�&|�l$�@Ʌ�:$ih��͉�T�d��Ӛ���Z��B|�kB��"�jW:���g��Ͳ
����VPɮ2�0�ߦ��e9�ܝ���.�ӣ:����j�>v�>7}������!*=�k��X��9�0��2�a�출n��O�E@����XE"U`�b����1��՘w?l��F*����7űNDC��C8�_-��¡�U_~;���#ܸK�f��a�&�aZ1�6Uw��G�E�O�-�|{ҔD�k����T_���7w6���5�$���Q�YUַ�0G�|�44
�/2��נ�BG� X��y`&욝�8��// q�"��D+�y9��s�'�;>��F��DH{����Zv 
vS]�YI��R����.�`�����f�ǃx[w+�[]�c��eF��x�\����/�i�_�N̅�e�0������z����à�ӎ6��強$&�+'N������L��;��G�:9�,�g�A�����"�E�4,n	K8ƥ��hU��o۾�$E�� yV����n��)�XC`0��_�����)���r���y�;*W����_���@=�-y!�_Ć1�jcz�8����:<�j�W�s�����K�.JGN���~���%N�c�	@_�d��40�KCB:�tN� �֟�~R����_�TEۮ��	y�Le�1M�v	{��ZzJ��Z'�eIHQ'�i���%�l�]$��F����(؝k���͊1�?c3YL~L�=����OL=f�Z�2$�~뿿,P�G?��g��������1_�t'k�4)i�3�NO��4�K$�7Z�L��20M(5c��I��G��(ߍt�e���+�h];0�Rq��GV��)����Dl�{#Ԫ[U ���v�ؤ���s�(0t��ޡ-Z�rOAZ>P�����ra�����*X�Ii��(���
%,������!���3Fu�_Eo���B��Z�������k��:�يKh��?SQ+
�����X����#6��5�"lL6̘gH�G���\_h��,}L�b��Z��~
�H��N�,��6�!D�r�'�	�-��_�"�t��v|���0s�|��͝<�O��:��4�T�Tv���l�AwR�$y�L8��ي�?��}�cƁg���d��&mڈ��\��A-}�f'^ŋ[�~$�9C�\�cQu�X{�}ڷ�=��{���_T6�(�p{����ă���ݮ`8�6i�"�Jk$c���'�ß1��#*FĴ���ֺ0bʃ�ƥPs�hBQ�mWO�4Ajq�B�.��N�>�W%G�v��$�����'Aa�F��C	�	����:׈��M@��+"��׋d��W���q��٩Z�|��Aj������Kv�����2�\�,_���~Qb@T��X2v/d��Z�Yg��}%?r��Z�<0/k��Z�*����%�*ϻUp�:%L�z���h��n<}��)L�Q���c�F�R�RMo��'imiF�)�mX��6�C�G�R��/���1i��3aѻ�
�u�N������+p7��]g�}k>Y����K��`J�攟1Eg#~�;����g�Dm���:B����&�n��O���� �8��e�Աh{�8�ͬ�ެ�mj��o�-�~�ָVs�����u�����*���\��8��B��p���nsa�<c��n�χjIYwT�j>��Oi�BA�h�MXzMӁ��0�S	�+Qs~�V�A��8!ڿm_`f.!~��`���ݠ�Rp���-	��hY`&�aH6[��`�[�e�L.�lZ�����/v����C�x�z�Q\�[��a/�H3����~L���������T�!��M-�F(V��nKW�}�PD�w�cq�q�Gv3v��a���gS�����q�!�b�UW,C�e��(�F��ё?X=�λY�Lļ |�(59�ѝ�PC�lߏħ�`���m`KR	#w�nۡ�ѕJ̐5�!��&��PR�_��>��k
iN�o*�y�yQ�ϭ�0bQd�*[xfՖusТ.v����)f\�����x���ӟ��<]P�Y9K���9/2�Z�����nҺ4�jk��
�\�����Q,��޴�	�/7��Վf��e�-~#�����J��U7g�4IHskGy�1�FYV��g�$�go`��@>M���	D�~�MR}�Y�� �h�I��lF����ڰ�T�1�?F%����ͣ�E=�����eߪ��I��>&����Ɵ�fx��r϶ϓf�?d�6߃Б��!j���R,�-*�**!3���N�yA�j}`�}f��o��-L�7��/��KyPmZ%^"�����Y�<�[
��v�#@u�C�h=*&U������](3%ד��^+C`.�@�)+��+aG
:]�5��ss�����\�s� 7OZ�[�'�Gd�Bt��Ļh�F�]�CN��it�%s14��õԅ!���ݽ�S e$e�c�q��5��&��l榍��^o�4�P�i���hg߬X�q����;�-_�:t��a�	#�tG�����{��]f�WO���K�@WP��[�Q����P�hweX�&��]�lhD�I�H�U�5�8� �ٔ1JN���QG0!+y�3o{������C6�� Q:�U���kT�A"�4��i�l�Hu��,��&��Vn��pl�f����N&�5*¤�`����U+#����קJb�D7=���:��O�)���M$O�z�_�2Խ=@lݹ���ߛg��O�+���3]^���a��Ja��
��1�����x����RQ.3	�Ҕ���1��4�5�]=T 
�,��m����:��(�ƭ|�}�=�f"_���ܮ<^m�ȡ��mV&�O���4Z��<i�̳N᧿�
x���=~;
��˘<8���`֋���.�ʰ)B�`?�g1|�E&�y���z��a�� F��㑮<��[O������ g��E����e���[�v� �|<�5�iʮ��!5Nо��r�JV?}��9s#q!7DC����3���Ē�8�J?�u5��b�0P�1��َP����5m��1�O	�m�r�w=v���y���F<3�\�d-�3��U��9��z F.�	��|5��p�{���â���yU^��*$��-=�U��#��E�n}�W[oYߐl
1�����w,g��'��~bU��m"wn>��󤫐����2�������^ ��%O"<_K	������8�-�>eQJ"��5t�1��-��xҾ:�E�"���/�~�
~&�9��N%�vw�R�^R�T:j"O�y1n�噢{�U(�d�RE*^Q��)E-�o�o�ݍ��^�]~�����%�p����'���3s[5Z��|��`�0U�՞$Y�*K���`*	�[3���n�I�m8ި};
�ճ�WT���,R��i^���̦L��N-$���Zv������)���9���mgx��\(���Q5b��O
_Ȍ�˰�}�ڟ�y�����#���Kk�`��]�O�*s�r��c����[~W�Vo�{��O�H��1��ID~_�;>�*cs�����:l+`j�K�9� �ƙlmĘȵ��ͣ�*ƛG��7�0	�F�L��bh~���2�5Ϸ@�8F�_䁴����%q�9�,��!����Wy�m6�5r���Iـ�{f�CϢ����Ņ�Ox�����b�{1ޘ��nV."�K�W车���<%V�=8���5#�<i��C[�$F[�SGݙ3�ܗξ�&���LIX� 9�p�6��!"*�Sh�Ƕ�X|����zY�� ��9v�gԌ�H����������f��u��d����^<����q�4>%|�;�YBc7��F� o�qR dh*�bf�j�Lso&�_���*>dA���"�3վz��J� Qq~؆��^ΉBe�k�Pc��4)�\r��H�i�N(���W���em���Au+~܍s��]2T���Ȓx5bh���� z�����/X�e��0�)��N�;�D�,v�7��q��K�8|W���J�\�4�؄&�R��b�:�S��Ob�+���س��:��^�t
v��4�"i��1��3��֐w3�&���+�V�=OxW��Yw�u��z{��L��|'����ӷ�r�J� �'���(r?Ó%��J�T]��W�(Z�V	��S���>�j��,h|k2X��!z$�����l��%1�
���UU>|��vCs�&ykn�א`�m��������0�I�����)!�X^�\��$���T�Fz }��B$�R>E+8E���۱��6����ݧ2�S:g-��ӄ����,V/�n�(l�W.���\�[�6|��=��F���J��Ll{'��BM�X���\*���`bb<��^@ǰ�"9U���FUXn��6?��B��a7��!W鲠_*�Q�{7&{��"f+�r�j�(��`\����n��ƷF
*��� �?����� �FS@��.��~�"�����0~Bʆ-�Omc�pc���-����%���FgEc�g>�%�
yz��xϏ8��rp(ɯfa('���'�"�2�PT�o�෈`�F�3�Sp�p/����f�1��^�<�����:��3$�l6��Ǖwx-���mn��Fet*t[�.����eO��S��k��}�V]c�v��x�-GAC��љ�w���:̧�W�퍔���kQg����	Ď�f���X�6��=�@5�U&����m=�sR��i,�`�6�C\T�J�y�=F��S� 7���g0�2OR����e׶�qҎ7qD�K�Kߺ��y�?x	�(RC��R9�:d��{�x����K�$�Bt�0Ǡ �=$�m�#e�0K�J�>S�p��|�6h-�C�%;*o���8J'��e1�i�/�\/f�dFH�%K$���Q�����Omjt�R�u���W��AL���Iu��[΁R��O��M����Y$�<��ۃ��T7[�����э�*6���*�ҕt�)/9ʭj��ؗ�	�Wa��QuK|bz��A��%�^�p�����	�a^Ԙ�=:tW<LT���2�U��Ţ��N��h{N���>A�{���������2T�������2H�9ۿT+ �q`e`����-7${�J1B4}��J�mb3��q�7<$�l����zh�Q��h�G�vq4��g�
]��]Ki���N��</,Xs����4K�!�k��� o��y_}�#��đ�`��0�-&Ȼ���(Q��g?��C��/{�M�7���dMd"�>��I���[Ī9�\]E����( � (T l��yQ��
&P"�=�Z�2_cb��.EQh/hz��՗�)T�n��YV:D-={%���,�����)�$�雋�^��v�������'�7�6��<_�z��9�qb$תeY���ӏ�`|�����QZN�
aK6�0?Bb`�$@�ߜNz3��Iu��F��ΰlS"�T�_�6{��(�M�u��Y� ��$�,��r��V�����Ss��j2��!"7�<D�/��D���_�|ѫ���y{���(��������·��Ǎc ~�}�����RN_ZV��eH}HZ��shI�_�]��x�)���#'�Q�H�r���E�Z4b��0n�6eDxUk��!�Z�j��uaß�*U_�-S}�+]���x������-����<s�hݭi-/fӾ����{�7���w�~e��~Tx0�3��z��i�$G��(�j�π��	,�¼k1�I���3��}f�T�ּQ��o�D�٭�o�׈���i���3}���	H�W����H�?*��^Ԝi�x�'�%Bf9��L�Ъ /���D��x�� F�E�*4�5���@A��o��b���k�Aתy:��~jk�8=�{�e��Ȭ�^D���%}�h�6�(>�D��Ӊ?,��z���&X��=�-ڏ#}�?ݩ5�в쪙!�/uz�YeM[���s��,e�|(�R�|z�]���ƪ|?~�]e�	3�\F� ��.�Xq^g��O�^o��!��V����{f�2�m5�w޻YI�Ъ>���T�֖��3�P� �N73������vy�-��%�Uڌ^�ٽ���Cz9(Y�ߢ����-s��	`�|��$T<�u%�F��%��D�*�T��^{�9ֲ�\����U�C@nc�yـZP���X�>����5^��C�ɹ�L`������(�f���y���r.�C慕kz�ւS�Ppeu׻M\%�m0�����`+"���� ɜV��U[��f����z���-�+�U��t|�v^�"�-�{� )��ǋ%�N�K�Mu��i�G�e��o�YH	@H��S�xj?��ӎ��ȏH�����.�A�*9m�2j��j��T9_�a�g LO@�O�nL׫C�ݽ��)Wt��k)H�t���nhw�&���DX2﯁Ԁ~�} ���&#�ByK�>��� 9�����,��K1�n���Y��W��h��cǇsD�)��8���ݠΗ���q���7����X�u,@��g�������:O�ۺ��Y����{5 �tz��Xe�����7B	?��p�m�9��$�7yC�.p*��X�=�T�Y�Ը!��L�8��#� sDH[j��#nj�k��	h6~a(�g
2���9��?�T��R�TlA��$��\�{]>%le��Do�d+�����*>�2m���Ճ��kJ�$��;z�C��7+���N�8Hl�\C=y~ь��-�"ys3niUх����^'�YD��C]�����,6�� �	�*���42���UЇ"u�D+��c >�AH'����_r�gx��͹���{�/w'W��G��5�A��_���ɂEZ�[q���$�gS�I?�ah��F軙��~Y�!����[�%��̢���&:�+�	$���Z��t�f���ߔӳ�V }m&eg̀��:
��l4�u�:s7�w{UW��Hr0��e<5/-!�ͪ�ub�9:��H�	^�$�s�;�
��O�/$��P�p����~SL`��VK���&�o��	P9�)�GO
��:���v�`J$D�.ԋ���R s,��AF����kɊ�Z�ڤS����g̵���|(�-��ߢ�(z�f��?�/B!�	�����s��
� �cؔiE�$[�_1`�F-+��4|?�o`xd��'�a����@�X{x@�d��uj����xԡ�th#�$ڝ�a=+S��kV�k"F��CF�������b��J�{��n8J�R@�)�åf[[Z�v�f7�8�k��d"����9_��k�~l���4$��ۥ]��c���U��s����Hql(2��;ō(aQ{�V����36���jB���C��*@�u)�3��d�Vm�k9�X]�Q��4O�Q�[M'�1������`�^ �?�uU���?&{%�Ao�Bh�I�(b&���Hߤ1�����AC��Q��`��屫�7c���dM�֕zY�����&<���(�4���%�Ίa�_�ٻ����7ϩ颦�6Il]�$��S63�xSx��tt`)&�lXƉ�{�+=�N
3-�w��@V(4i�*����qk2W1�챤�L�R�a����*&H��ߓJY'�0���|<������^�)������d�91D0J=������
�*�Z�R��c���ᷔWI_�e0������B^,������I�$"��6�2t1)���5���gmV�C�	���M�}?F�@MM45�D������|�_Z����}�1��ɹ������~S��t�������������\T��9aaj�������N��Τ{4���X�t��]_I'�	z�9W�yVmOc�s&���<Gp�� ȟQU�KQV!��'��|U�ԫ�n�ԃ*��+w�3�z1*��o�q4t�hH���� ��5ٙ�?�ە�-8��CF�\�p�¥e���k7������i���n�|||�s�L����|�J�;�xL�o)��xӝB���ڍK�K��Qx���ʍ&�=8��l2*�FB�0	�4�I�/֋�~']�:���w�V��*B��=��)�]���"s��sU�"!k��j�c�m�,�C�14�.�2�gZ�?%]x�"S��yL�ؼD�ˆ�������;�
�*Y����:~���P�¾�r��	[��KR�h�Y���|ͤ�L
L{I��$)%RgEa�/W��%�RFag�M����rc�D(�L0s�oA�'�uX�*�
�A���m_��Uo"(8�p��b��0�<�+��MzZ[�/���ī��Ӡ�sd^.4�`�����gEf��B]w��X��������t���1|J�,%�@c�M�s����R��5�������Z]������΀��Nj���#�"��D��]Qz�cd�U��I���6���z:�k$�	��q���CCs�xȓ�G�$�$��T6櫢�}w^��<�[60��#�I5���
Qbˠ��oүE�O)7G��>�=����4�H��r���ͩ��H�[HVK}2.����� ��
_n
~�k�!&Zy���چC��̘� /:�¬7��12f8-�=}
A�<ZE��Ż�+��:qod%i$X�S}��9��O�KY�hnO�N3�V�T�A��{;uc�kղ�����ڂ2_��S�j$��!�5��*f���e�����-�ÒǦ?���c鏀�r}��4�um?�УnDhC�?4"`����K�~�m��'����״�ߍ3�#󇦰FL��Z�1���]ޫ \kv�"Eʨ%��BT{��d(g)E�D%����.[���_����=�q��&���ݥ�ή�@�B'�I��o��hIϞ}.�=�*Fl�֦�ϖ%��U$4cd>�t`���S�,wb�F����*��)���MB*7=�8ǲ�n��p��q:e*Q�6|T�T�G��)��&%a�f��̪Ǯ�;�������s�4��zj��lë�pH� -�hR���(���Rζ��@!i���h�]bei�f?x:���ǽj
!�\��`��$.֘=���T����H�䆶��	vW��7��:�r����xO�!��R�(8��
Պ~��S?}ˣq!�q$��E���<~xz����~Ԟ����2�tS\��V�����cN��$�M��1�N��xL>�X�$p�/��)�!>x�o,5J��zX�
��ꘟb�|���A�D��]��|w��V���h�!F�l塑 Kg�%C@E)[��!
4}ݛD��6լ+,�ēɰwPÔ���#~&G���b���H�����Ē�WW�{m�ؤV��֙k�q�*CG]�V5S�Q�ڿ|�qӐ	�p�<V{����2���'�r��?r^v���OO+E˘�m�K���B���Q��}0��}�B+r��7�s��yq������ ������3��-I��~w�+ʇ�:�[_kہ��)��D���CU����.ĳ��eƟ-�Y�lq��r�f�؄ь�)���Pt�d"Yz��, 5�ţ����U���EʯW�'�2t}�
9��x�YsP�:H%��E�t�'aD �sݝg`��\������
M���k�0RZ�-j�rm��%'L�)�X�!B&�[�L2�2VI����WsףkK���ϊ{�ǳ�~�Fdm��E3�cp-i��3Z��v甘�S�JHq�~'J~����Sn�XwC��^�҅u�Bk�y��|�6X|4�&#��KV*��8�*�4����g\�
��;��!�E����� Z#����~�C¼�g�䠝jWB�O�o��K#l�F����ϑ�ΠhT��qў�����w��B�z�=�^���tծ Z��M���-B �31߲���X�t���7��7N��!&φ���ER�Uͅѧ}�x0h,�C�?�������KK�c7X�H�vR��P�-8�Q��!z߫���\���t�P ��ꔇ�i���x	W{9Yg�!���?��?�㇥���{�d
(YV�X&L����nL�&�E�H"*��mH�v#E�fs�>f5��2C�0����I���?�@�W�u��Y;���P^���k��b0�b�w�tV믅f��6CG�G�!�B�'*�a�w�_:*h�rb\��]Y�&�I����ʘGʏ��kD��Bn>� Y�����<��5�����W.i�>��'��C�^�y3JÓL��g��%�n��Y�J���]��j\q#EpUtxm���CGNߞ(�1�A�ב=������6p�@��.��uU���M��A�i�և�k���.�#t�]����^�1Q-��'�J�b�*{'�T�8����آ�g$no�3�9��b�^�|��ɞct2KK�4�a�N���� �'v�=�;Jb;|�lR�<R���Z�ŎC�ct�9�B�`��������J��0�.�?J_�/�;ڱ�Y�I�c4W��kPF&�YY	K2�2����o�ҠO��ly��b�NS��/�Q��_ghJ>z`�o[d�Z��soL�%ƣH������-54��n[�d=�5�*�Mٹ�0D������$����b{�C3�����{���c���:s��������o�t��Am���8E����;+o��$׻���+�ܒ�)��X����=&�P���m���n���s��FZ\�cEY�QQo��G��Gz� �3�]��ΙZ��,�>���f:$L���Uƾ��Hr���\H���d��)�g0��	�aV7bH�aq��°��q��� �P�̓m�"퉳�|�����q��4��x��Ŀ�^��w0�梵LY�^�����Y~�RÁ���Ɋ�H�r�]���FR	�����=b�k�>�2�S4��3�kQ#�^%=%]�$s�������pՓ�5�[u���|'G�m>VF�©�!?�;�Q�N[x��ٗB��설�
%�P-@�i�L�"N��F�����Ld��xJ�Z��63
�yE{��In�j�$��m��Xa��X�N��vW����W�%�.��{�W6��X����r����W�y폮]3���ZL�0nf�j�D[��kw�J��8d�ʈ�>�Y�����C����w���vC(U	���=s�a�,���;�קD:�g�ۊ��� z��RA�0�Q��p�i-�t��gL�?���{md.�Չ'��8\�d�X��HR	|r;�nK��M�cD�l>*�Aɶ\= E8��b$-V�9/������ܘ����U�>���҅"����ЯDa7f���(�r��@��e�JۓΚ�����	+����cl�7@�1հ� >�mU�2����&
j�3⤹'�
`7�|ky*�+� p�MwW@���h$ѯ����k�,,V��`@���~5��h�e3�_oы�߁��⵼�X֊X*4��}}�W��\jphJ"��.�y�Ei�huΔL�j;F2�t#-������߯�PdV�k_jt��VW�yC�u9e���~�'G��.��:��G�o	��z'n��V�X%�Ƌ��R\��7:�d0'q�4䓨-P�?Kz���u���������鄃�_��0,��N������I���
�"U� ��Iy���md�����cG$P�� �݄t�oy4��t��q`�{*��EOc�;6��y-@�\+�od��5��5O��n�,*s=K3�/zxމ�r0��*�x���|֑��-��%g��	N7�D�a6w�8z��+�5:^č��3�P�f�V��ڑ#dR�x��[Z�,O4�⒍�2��;Es0�9�V�DyE�o����|���$z����w��S`�q�]1<���]?d�W4&����X�L8tɞ�PU<#���fXXi�iUۅM�h��Z�М������k�n��n.��gT{m7�
�[7��K^-e'�G(� �|;R�w��ͥ���42�Dj�b4��ՠ'���J�}���]��K>Ϊ_���Ly] f*���hc�OAї��w��%e�ޟ�'���'�(�΢��s$�YCĖ�n��p:���R�}���Npe�L�&�e	�62�wgO��ފw�\�B�J��*&x���D�3|��ɸ�V�f=�}G�9�k��+�6�<���v��d��!^�v�-M-��利�m���r�q��pK�+�ƅ��ZsO�� �o1�|�/)��%�9�bZ���@l�1��!$;�v�h5,�;����WW�J&y�".��#kjDյ�ϙ��WS��!^X��}���}T��*jiA	���1.+d�s���N�!�Ր����̞���z��������g;&�Ѯ�V����z,�������b}��l�v�刅��+;9t�א_���.�{L ���[���p!����X��-�� 7h�e���mP���j{�z`�%A�OGQ6Ul�:�vwGQ�^jnz�A�G
�E�e��	�]��?~��И��uñ�В7�����Lt��&�C/MMQ; TPzHP��w(�����+Bya&v�A��PJ��`��)3�>�جs5�C�����l�T�&�^�Ԕ}�b�1�;�Kn�>����m>%}x� P�����$.#F���!
��6~-��|K�c�,����eX��	� �;&��r����gڔ�8cE�̫ʑ0���%Wx�{����W�C[=;�W�5���V_mjk�W�_�C�4����tJ�2)0<�J��K*g���Q:QVS		���
^��[�*�f�KZOW%o���QN@@|����A�����|�+�X��Ʒ�VE�⹒lL�iT�:u'̎���W��Td�\5FN�;O7�G
�

�'py�<�:�g�nj�6q��t1J�C�4Ӌ��IV���j���+�Q�E��,+[>V���eFg5�	jI_�n���D
����2�Q�P�_�nXy�=�4[u�oݺL`D0�����]�]���=Y"*Zr�Ez�ɪ%%p=.�D�ݽD�aHD.��[9$x{l9Jf�x0+�F77���fH�<<R���\d[ �m�AL$�VJ��~�md���@_b��%�!���T�A-�b��FE" *�0��|��Wڋ���"&�+�3]ӷ�;��+�Ё�k�)��d�~���X�?�H��״���'(�i�pѺ��zo�!�y���Ќ�a����?:ո�2H��0��-��;�D`6��{	�:9�ו�_Fm�+l�H�k�r�N���8�z��`g(�hmmpPdJ|��N6����%Ⱥ���;�ր0�|�c%.	í�jo\�A���X��%����|����������㭓o�I���\W-."]�Zw��:�`�*I̹���p����+�P��_[i3�m2�� �|sd�k%^�>���G!|)I�I�f��5 �(�0��TE~!!���x3O��ՁI�~�����8��E8�Zn%�G�3dQ����A�{W�jBB�������XEQ(.�NC L��bNh�X2_��l���2�L�Hf�{��d\�[��h(��w������VPZ."6�y�-�Bp?�%K0LK��SI�*�=ٳ� y�v 2׭W�y3��i��K6�F������:6�N���FiA��v��2�"��h�o���� �.J>��3����N�S��Z��p�u�S"�m�s� �-o&��x��QI60D�j#�l�K�	��f:�\Os1�&j�xꭽ����"�?d�F�
5�=��@q�==\�Xx{�^đ}>��������`��N�Q�	đ _�:���.���5�A���2|i�p
�0��y�@@���y4���G�!���V�Ҿ�En��x����](�����|ֱI��!`%�qJ
�˳ ��^cn����CGK����=ZY|�f����<���M2$��b�����DM� ��"��KI�9��j����s|��c�#f��{Gd4W�dk"��
Y+w��8J������{����H-��2�<��&�(=��arF��U�LȶA:��:"B��H>H"��.J�&@m�N�����0�I?y5x�@�kڊI��Г��`0���\�Q�d��1���d�za�;���?6gb��d�� �6�Gҭ��F�K2SϷcjt
\qIn��>�ķ�UYi�"�A�zծ�����#6��H�����0�=~�����!�w ����)�gNq�<j��sK�t�v�P9�q�J�UTW�L����#�w��0���L��F�ͮ�eT�~zU���>�b�#��!��4�V3����kq���{)Ĩy���$4���u��z�Bm Ք}|}F&���!4�a�36Dj҄��p��n�X��i�w��d����+Q�e�k�F���_����G�3�H�y��B�+�ޤ�d?��Zu��W�T���y7�����K4��*7��.�[�ľ����QMP�(ܓ��x�ː,5vc�\;�LD���C2����E�_ݛ�Zǳi4C�䕃.M�~���Cc~p�����`�)*e���o��]1�-��?A�s�wӳAM1�����Ѩ���gF)<^�"4+=9�n������*�9�!���0�λG���ҡc?J.�x�-��>�a�ē�`�H4KX��m�����_3�F����A�8�E��@�Ǯ��i��L��ͦ"��#T�֛LLB�WJ�T���_��2�G��HZ��tiQ��Vv�`B��Ġ��
J�D���L�����ϧ�ߜb�POP�vQ�1��Sb�Ǐa���Q����ג�ȉ&o��MNA�sJ��ϣp�qh;|7MB�jH땱�Y;�?2����Y���VKtX,�G��(&4�K������8l�a�vp��JyJ��(#�%�!�P���q���/k~�x^5"L�|�G�t��Ƥ=kO�۰=��A�ꦤ�MI��<g�ff�P
ˢ�vRö�  ��ʜ���t�Vâ��O�UY�n�_�0�)f�i��v9{�i򩬴��
�������]��������)ڀ��wX�U�U�ӫsYjS�ӧ*�7s���?��g}o�Á-�}��e-s| �I ;�y`~��I0�;�$��fn{ϻ!-/���?|x�07�S?/��+q�E�㒢C\1���>N��V�>��#"���ݙ61|\��2��q��I�]G%��E�z (e����Č��G��j�Vጓ�w�E�9�3�@l�'�:bE;�!��s���;0��vd�p�P8��΃�߁ߤUk�;�uHs�N�l�l�u��3������g9.?0`�������W��
{��v�Z�(�-���O���\5�*�[3�^@��Y״���YXo�f�ǟm#,�&Ɂq�FK��?�ah�e���&�U�1��O���3���_`,�w����auI|Q%�Jp� ��H�o�o\�튶�)2}�p>r�gM�wv�9;Tҧ,�"OH�IT�1Q)�C7j�+����'{���1�p3B��bXF�D�q�)�ރ e���oAP����H}�#<E'c�,@?�旋|K����?wv8��k|ȅ`�����M��j�@�z��Xس�[�Z� -&n����H���K�����/��Z��m��	���^��-�+��>سS��t�EU;��j9��
��қi�����3��ٜ����i�5����l9(굑~'�1E� >k�'n� ;7�n����	�T���P{'Q�)�`Frs�*��xN�f�P)#��[��8������@�l�`�H�^m;����F�$���*ZA�Yp �R����o���><=� k��gf�6��g��'�[M�7�� �����A�ӸeM� �\�>�����gu��^��L�3�13�Vg�;������E%�yL%�W%{�`E��k���1$�r�� )���њ��B� ��e�����f�S�|o:pшM��A��G���X�|o�!�����*N<���}m�l�K�� :��v����aج�0�0�,�]��J2���qFEjG2����=f��z��	/�(������Ƞ���A�'��Sy�KA�p���6:�%{s4�0b�Kl���Z�����1*�N�9ګQ�7����7Qg������������+1���<�!(���	�2����@�6�����O��$>���KV���`=��ٷ�B�����Rp�W��(T�c�������#J7�����i�En;I�9om�L�{�h��iZ����.��ϧ^��&�K��oܘ���&>}����M�f,���؞IؗxрTw����3����g���C?��Ka��ے��ڌ���{s����nщ���dI��Z�΁�x6��G2u�~^�7 ���{�x���v?mn��^�
JRf)�;n��R"o� �W7�7�d�|,J��_�!4��䬷g2��%�ͺ�g�N�B��_r�����oI8t_Aj)�?�$������"���^�ꩨ��ĺ�J~�v���m_�P1�EM[��H�1�t,r�M���	��W�?&;�m���>�+��j�?�ݝ����sa4�l�q��Gj_Hډ�v��)޵��S�*�/��7�ޝ����a�l�8f-'��`.�B���!DhW��m�_�(��'�(M&���lhc������B>5=v�j�~S����Ad������諷@��d�I�C�f-�VS���i(�'r<ЏF���|�^�MJJ��h�ۭ� �1�^k�o�����ϭu�"u�E$��3Lu��l޺$��a��u���` cn��99�"ۭ��������k�+"9��d�Q�b,�XQ�����YU�7Bu���PM�����$��x��)%D�oo9�����0�@)I*�[뢟h���ĒT:�!��q!�g�`�����|q}��mh��ka���(*D�Fj%Ҳ�F��Xggs6�	�L�!��݆��	lW�N/�q.��j���2,��dhB�&�l7�_���OjVHJ~Inr��[���ϴٚ���R�3%Y��㞋�I��W��������:��U��O�azFr���K�w�ōs��1�J�'1��|�*�߯��O�̀�}� k�jcD��8ۏ$�h����YLu����`;.�oJL�#@I�֢.�rYvd
�9����(�2h�顤D�5�����& _��wZ�@����K�	�sK�?��w��������]���I+*�EB@�� �#-4�ǈ��L[Y�/¦��}��1d������}N�c y�a�B3�	]�@p�E�����}Nk'�lVpa0����ĐB+��٬ ]Z�ʝ��c<�o���<�!�Q���uS�:�+ڪvK�D���}|�ʈP�,�;���VG{��k���7������zf�h4v�<���Z�	���}Z�QM7_'�^���k��Y�u�Iy�Q[����kIP�u����� P�̲괜iCKQ���H[Vt�=��tF�9�P&U����H���RasQ��M���u��맮(,��R�0zҴ��kBR�>EPaz��~������|��������PCD�6�|�#2'1�5�x�������<�M��~�4C���];	ܩ�T�a�e6��ϓ�ݼE�0���C��T��:ٜ��3�!P���mM��
�$�j0�Y�A�Wj�C��<h�_� ����F��!��˨dW�	m�"�"D
LE�Vhb�/y��+bIۋ�����@�}��:�R�&�ž��L�ٜ�lkI�V�i���վ2��Ƨ9�$
Bm�R��S�.Al�eq�&5iE�v�ԉ��w5�V�hT `�[=?T����'}![
�`�ĘȘ��Ө�*�!��_¤������H�z~��;?���2#?�-�Zʄ����*nd���\��{Y��Pdh�'���M��;�/S�}��*/�n���>k!��/��}a�q3�g��_8�H.W|�EX�G���5�  tή��sg�~Y nחIz&z���8���g�޾�r{��.�w!{�ãȄ��H�Xc����y�q�� R8� o��~|���������CPwc��-��T�����e&���F�?�j���.�tpO���Q�,�����B���� w*�l\7[[U(�����\t(f[@��m�c�-=�kS��� R���)��&�^�|����<.t��ԌmPd�hJ��\��i$g�x�]�:�&w�D�z���� S�������Ӫ��TB��ų���[��󰇨}�:����4]~�+����/$y����/�Sle��9w�(�DmW�91m��o3�NRb��{ۣl����i��`�/��0n�&%纐촗�"����"v��j�Wcfm�W�M�.�s	YK�w�X=��`�4��^�EɋT��!�J[ܭĎ��+Zڮ��⺴�0Z�J§�(��*���E�
e%0^��i*���d/j��ҫf�e;Y������։I��֬�ؿ
6��0ܢ�E
��ކ�mڐ���Yy�7Jt�^��~o�{�\�eܡ���;�/H6hG��/YW�'��ڥ�����w�c딶��-g\���f����rQR����Ϗ&��"��F���p.��g`Z����ǲ>@UsQ�Y�t��r[�8��n'�^L%���F3�(M4��9>�C�O�Y����0�J뗍�쑭XʲҾ��t?}1�Y.���>:�� �`��.�~�D+9����=��W��G��M��	���8<O���k�R7p�jQ#Q�3�"|�P�����s%�o'RŪo�&�T��0
M�g��ep�n[%mi���vBV�<���,m�)HDx��D�{n0ul16��^j_M�ֆ9�Y��G�u�DE���}�vWX�Y_�{�
��wR������G�r޸��š�4�m���%D����~P�X%�h���m����ؗ�]��˻�:���EI2�y@��qh�0i��Ư'X_+B�aʝ��,���<�G�k^- k�ͼ�	O��D��x!2OW�-���O �HXo�#gF����,����Fl�2Fp5��TKۛ܏9��$�S�ۃ�M�����wqU&t:����ɂ3��ͮg�up�ED��[��R \��:0���[|	���~��>'���o��r8@�g�*p\��eGq�.=���LP%ŵ�6\8|�N�n�/��Y�*��y�
���{�P8I����1�@�E'�\�I������g��s�Fg�=4��7�!�zE�O8ֈ�ځ�H}�p���qUZ�6�����q��ƨ�S������@�>xh�ǅ��1	Ƀo<��^눣b����n�{m�怦�O*����i����;���8�M����=�K�}q�w~7���<R�p��	��+z��n|��h`6�!�w�U��� �I��e7Ng���n,�#�'�HG�В�B��+�ϣlCJ�����'�*�����# �W���)�Xt��m�N�Q���I�2&xNT�w`c��pQ��� G�9h��%����{����Iwݑ�(���<��P(邲���4c���JG-"�bH�f����`,�U*S"��]�&+V��`4�.����@����C�=��际%2F���F����+��ܸK�f��SrC-a�'���3CY� �i�grf��fI��^E�!�����d�Y%���D��R��H8�=�g;�9Z}~�`c��{䁫B�Qa��ɘ�T����㎰E�7~�ݨ��!hV�C�]q�lg���x�_(�A��0*���q�ݛ�c��6�ld+o>Dr�kt~��r3����>	�p�����Ԕ�d���%R<1l�o��8�uҬ;�ۃS��{����l6�{M����1r�d�3l1E�����,��,,=�;L��u�b՜vx�D�k�H'�紞��h��2�Ȩ=,}���l�`�6�E#d�T��2��Jzs����ɩ��ʌ��Fm�ֈ��LnΉ�8��n|P�*������2x͈V�p�Y�V�j��TeK���X�ނ����j͂z�=L�["�I�pͩ����1���MlU$SFK�;��N����PK���l����A�\��Ek#��ؓA���L�z��ߘ���P��_�O*(Ȅ�e@-;��S�-�q��:Rt�r�2�0�#�A��ݮyh^>2��A3�͹`�/.��&*tÉEt?W�3���1�^�B"�O&��yxu�Ų]�<o>�JC�ɏӆ\���i=M�n)��޸��e�-L�p���73)�l�#ݑɣ]y�{����$d�̈́|����$�υQ�rM(Ɠ��D
Z;ֈ� IB��,�H�Vݰ�(��+�c�s���{�=�\��F�f7�0��vJ�Bt~iCF���	[�A۳�Gĵ�h�Rc߻�܃�\��H��gN�yb-��Ӈ��j^̥�6�G�QIF�"�%U���6���7�|_݆R����1	���3k*w�gYܸ��\�sC�%���%U�������2{��e��W����<!�����j�N,�[�q� Vhа_0*�Of8MP��t��=Q�Ő���b��H����������:��X2�v�AԊB��!:wB!4������J;�Ɨt�f�5����bi��8p�2P9G���E�g�1Q�[�j�����k��+z]i��6An��=��h�c�V�F���QiQ2��������J!ͻ�Y�pD��V��\���ކ��O�+�l���(�ܓВ��0통"��,�Ƭ��}?��I$"�Bmc��J��E�~�[!W���kr)�� ��#c��Ʋ�߾�4��s�*h�r��ni�X���?F?�k���	��Y���q�ӄ��[�rg*��R�h�aSO����x � (E�J�>�mЁoV��T��s"J{�ԅ����5]���?��K�5���JO��c?�`5�;�5#����՝bX��Ѫ��-)*
 H�7�9�?��ύ7��-0��-�ߕ�1�X�,����L��i��rN�%,�E�?����k3pL�ŧJ=+�ɸ�P�� `mؒ��{�hU��ĩrA��OL���� �I�E�8p�^	l5\����X�m�s�2��-���{���E����c�ʻ䮪a���0=s,�C�e�7�
��\*��Ōd#��	��(��&-�V07��=�L���BU���e�����(��e1���n��=QG�}�����M� ���tJ8���Q�>@D3'N��N��h���X��0�U�`: � ͖ }����ݮ����隽Nc���~L���1�n�<�e^��
�n�	���,:�ƹD��������:Bh��h�pҒG�2��@� �	���|����M@�PճϮ7{��<E�w�9z�OV��5F{��k�F��+�i|��7�;ޗX�73 �1�i!iF�ҥ����'�I A����3t�_�&fdB�P��fl%`��j#��!�Lv������dx֋$�t��Z����ߪhb|�{�C���Fc��ӭ9G�0�F)@����X}��;Ne���;�Ր�(�������C�_#���l�aIX��|��ّ�O��W�8�vH��="��@cd�λ����0)/P�O�	E��4��p���Bb5�V�K�qs��,����[k4(���GD^U�q~?�kI��� e��i�$c�O/��x�K�]��im� C�V�"�WF�P�6CT��i~t���`��$A���Pƀ2��9���s�)\�HtqЃ�IUV=�U�vp|��yd{qM��D"N[��/����Tٴ���Yy!�(Z@����*<�0iS�����X_t؛$���=�N�Ö���c5�h���B{�E�+f�ڟA��,�
Pv��������v������@J��J8l�OZׄ�;��;f�ӘH}I�Q��0��-hp+);Z%���F?����D'N0^Aot�iF��4��� N͵l.OmJ��ݐk�#����tZ#.��潂�������Y���Qt)����j3�K�J������Ug$��D��dY�h��c2	���t�� \�r�?[��E���PO8��r��h fcV�^��rI�FKo���y�"։J�.��XL�P@f� �3��dr��R�(f��d��N��j&�6�cڅ
�B��m�\O������~4X��Ձ�=CS	j�
(oyw�װH!���@Fa0��&��S��y��hcP	�B��L:FĶ�a�$q��Bہs~��V� ��B?�qq���-ܓE<;NIag4 ��1A�D�M'�A�,#���&�y_�/�ei�N^�I��
��j�(r����m@�e�aB��F!������i��fh������MĘ�O���D�8�Rג�AX1�L#vA�z��D�h�R�y%����-F��qf")���?�����2����+w�\�7QI@��5O�ܿ�����,5��?��κ��ʰ�N�*�B�ID���1�3kCF9�L��bga2��M��7#˺H���R��A&���ϡm-�X�'c�.Ӑ�`j������%m�ڛ{9s��W�3|�`!�;�j�6��dRS{���q�i;f�VX�{���('�g���  śރ7�mѝɱ����g��U� ŻM�l��{B�J�rϧ�!�̞5t�H��n׿b��jmF�"�r�F��M�������Sܰ`ǐ��ᇩN˹wqu[�u>]��ЈT��LU��!`�֠it��w��PA����0H)]棿[X�c�r#��[T>�)@z=,�n	�p�R���8��W�#������hᄎ2����O��gw�lT�/_�%D����"�;�$!��yѣ!ïW�]�IY�g���yN�`\�R�*�-��̼(iM爢M}��Jr~�x*���^1�X9���938��֞�5��N�̐���j�$2$^��\�S<&e4�������!=�Ǥk�'6+�:	<�s�1�,������U�����$�/�VV�FN�׼<Q�ǯ5p��@:���@&	y;M�v�;�x|qǓ��՚�"s������&�\+$s�x뤅M���pj��j���k{�a���Ώ+���ǥ�,�lP��N��`����{xh������oN(�^��g��$Ң�5� �F�� z���B��e���K��tZ�8��d�(�7a���mɯSxv�[S6s�-i���.��Y�f��,:����р�SO�rsDv�����#�Ap�Zx� �!�5Oێ'>q=��]{/������6mJ�l�WvllL�yͅ�{�'V]]�+�Y+H�����1}/p���5gŏ1��8Fkv~&�D�[�%�S��V��S��l ���h�h���k|nm��ŤvYL��m����rY詏O&vy�w3x�@8.���z�3t�t�;_^↉R�Tc�8��X�!�)�w�4oK�r���0����9U�M�PJ8>_��������J�+�K�x������c��b4e��8~�X�UEh�6,��?�B��H��R_�a��h�V�k��MKA4��4� ���1�U1���Jj�X�O�zA�O�-��5� ���{-c��2�	�>G&&���v������T�Dޖ��$��"�!�<|�P ��P��aѺ�%�ٌ�3���?����p"=_���7!�欷/"�B���텺f9���_�y2~<q�b�8�G����Py�cwc�`�{6xF��p
0�̝��LK]r.�z+��$�����~Uwn�=a���t��n��(����5���<�����X"���0J���q�kU~7�d	b�v��p;�����c5�Ɔ[�Ҙ��灸�g��m��	������&���B��Ԗ�,8\�:,�.@R`���D
5W9�p�B�#�����@Bi��o�R�,f)����-:oט���ŋbu�G��/(�D�x'g_��[��Yc�!P3#���O$���H\��๫h�27�Z�bU�d�$���4-��=�BS��-E��	�I�?f۰m��1�cd�(E��2��iú�=�5s*�,��4L=%�#<���W�a9�l0�[9���LۓT���S���-A�@P�ֻN2�m-j��z���_���q3۸�g�g��~���4�<}ʝd����2�4 �w2w�p�fzA� :jQ�<qBpi�X�j�jϞ� rX�8�@��d�Y������m�}3�?�W�:įq?�`o���q�u���:!�=�]q��-����z	����垙"����!&� �	\Y;I���ZT�ffЂ�I�xc:J�D|����R[�q頛7�Z�>��ǆ�qH�Yn��Y+����Y=���$�QN,U�*�̅���)�����������P��~���O�P*Qʨ�`����c����s(�>(n2c|e��O��t���0z���LL�5�����H"��X���TJ���U_��\S�ϗ�h,������:hl2T z��N��F���Nk\/��G�j��
f|���V�F/�ui�2F^�1z��f�e ��)���;Y���Nmf�����_I�7j���3����E�rz[��i�4HV^{ ΀)`"��߶����C�-Y���^�d���.���H��m�����J��!MP✘Bk�!�X��{�ͺ�7ݣ�#I)(Tw�m�GEe���m��3���Siv��!y̦N���mY���2Dp�{*Ue�pQ���sʆ9{�|,�2������R�E��k6�& ���.���iʾ���v*�c�z�H)r���bY�:г�1�F_��¼!i4H��ZҚ�6��A�Fa�ʈ-=3#���m8�m�[w����t���#�2�z�,fft��yf�CU�R�Ws�Ht�|9��zH�H*-YE@{zj(JS���m�(h>��[ UM�NFW?��ג�H� W���,�p�X�������;��P���֬6�O�{���vW�����̷�8}�
�DM;'���8E�$Fu��ūV-���W��Ge��q�1G7����;��Hj$&�����/�*��ν(I�n_��{�],'돉˪�y�@����2�_F��F4��3��=�91���K�>������߅~��՘$�S�ܹ3�6.�Ӈ���8�F�jW�9$?�PAaO��e��9�_�~��-$	�^����K_c|n���Rr����^x%@/	�K�1�bq�MNz����G|}*/O���>L^T(I�e�(��9�!��`r�n<{o�ky�e 	,1�xa���`3����:��<Dׁi�&�E��c�o)C\�p
����H�|t]N�]�J��~���7�v��VI���|��\*�m�}��!��JMhH�S�����a�42��;+�<����[�Y�m)P��|�"�ZH\��]a/C]���x�W�I�[�х�� 7�:�]#Bml���s���=hY�E��*��EǢExi&�է	ą� ���|���Kߗu|5��5s��V�Խ���<�aݷ~�)�W�r�����|�K��f�F^5�i]�3�:��	!���;Oh��\�H��J�����< �P͗�Fv��\d���{�_�̨ߴϴ��������v{@�ю��MD'aK%��q�Xf�%nN�����5јU��&;���xZ&�%�_��F-��6^$V�yb���ony�a��-� �&�DiCo�j"��dՒL�m����.�~���	b��b
���Ĳ	��p�N��ᘘ�!�O�f�S���A�Ϟߒ��(Z�|?p�Q��T��Ic�
��1��O�#�&���j@�m���R�b� OC}���Z����[�b��3�B��c0pνK���-� ��1A�R#��`�����"�]��!��h` ��]���v�qt]8��d"�!7OX���ܱ��B;���{�#w�@��_�Eه������6W����:���͚�X4~o��v�/�w�<r����)��4��c�x�hM�d່
�vor�B_�A���ChuO�h���τ2TG��R�"!tĺ�����Ґ�#Jp������#�����g�o�Xa]O�pag�(K48\�-��K���{�	���8�H�a~����x�݋\�£'\�ʆjv�M�Z~��5���2�yg~ �<�!��u�/�+�Ku��L�D���Q� �m�~��1}�Mb�Q8���I��K8z�2�-pVK߈V1֯`���q=�5��LH��ɷ�U;�e�9�B��h�3"��G��ѣ�ۑ���>�R���<�6_+�nc߃�h�f$ތ��F�:����Kv�{�FD�N�EY�o.p��u�,L�܀߬�y�Cj%QN�6k]a���'��GF#�W�:��ld�Y�T8�Z\����.�rψS���J�?�Z�XG�?����8���u����]�E��7��v�Kw⶟� _�9�)=|�nEFT*����|��� ����4p��QlQ9O�*�����Y@u�����_m?���~<e
KJ*�D\�d��'YEZ�z?��B���C���E8���׼�R�b�'���(m!ZI ߈���- ��	C���?���n6>K2��[3��BT¹��p�����;b�P���Z��8�"�C8B�������-6�3pZe�|h(�		�B��	�=/��
u�������$����
�!�3?���ƴ�X�!�ʍ��c}}qܟH^]<�m"Q���*�<�j���*�|/�Ⱦ�?k��J�����V�a�j��9����bn��{���r;S��&�O���` ���c���y�%%���t(�ݙRQ�6�F�m�ﺙ^\�j��Es/<O�&¤����� �$S�V�T�r�};�]m��}@��"5]�2����t��������I) *i����e�Q������&���=���0��;^o����L���_J"�;�%��u�7���z3�M�hh�஡j��H�b�f�П�]*'I�&Է��"9Z�4�œ� �������6.�إ���&��T&	�� q#&S�_�>�UA�U��9}�]f}�I�x\���p���O��M�I��w%Hl!c�G�ڮ��������w�e����Z��2�aa��mf�K��a���D_���8j���(�V1P�Q3��������c�6���4غ�k _,�(8
� �a��_њjpp���g��J1� �þ+`��܄��\<���z���� ->�_�&M�/�]���������u��x�`h�	�缰RԻ{f�YP%��ר�QV��x��qL�Y��:��������O��:M���j�/F����o�Yʢϵ��;�~�0agW]}R�,2�}18�)�#���s�*)���w2��C)ě�i�r� cl%��GU�z�L����<7���<.y�H��
j��lH�*s�]y�^6�� ���o�0��t2�sd+c�ps~���� �7E��e4f�taT��0��ŠVZ�ds��rS�1)��P�ǟ�3n)���e�4���Kz���K��v�S@|��m)��ct���,||����4���*�C��	����J׺]Ƌ2Z��$Vqׂt��'m<Ԃ��Y3������dlA6�$T(p���;2]���7a������i'(���c����܄ף��U��l*.�/cK�,>۪���3c-@�x���uk������\z������J-؍��3ض�.�B���L	�+ڑ����,h@��1RgwU$�>i�1��M}�nHB�]����%�h�g�Q�(��YD����Y�d��7ex?ګV�-�Ar ��C�$��'���n��%�d,1������O��=�T�tk鼈A�{�%D0��NLN=$�8:��K�� .�N�z��r��j:ݽ��oL�.Ssk ƹ�̼g؍&��}!�^��]X�e�oƁ��!�Er�|`��~�:����f��C<4�� S!���⯽��C���E�B!U�G�C�̘������G�gղ�[��S�V�:�EE����{ځ;�c�J펥Z���H|��KҾ%8=�zQ�{�pˣ3��SzGz�$}�,$SYd5���*��9��dZ���^ϫ��IK�"Mu��/^-%P2�^�3�k.o�ա�i[8ȸ;[�����T�:kΙ����J��b����:ǲ�bm����`�r�!�#�|��:V�N%��͉�t��܏�t+����kO�">�hX�#���qi�`�s5��%8��*(�ޤ+o58��[�����/�C疺�`����$�����@!A��<1�nj�2�D��۴���ဧ�*|>qH�D��!d����	\����2�k�V���d�Md�o��N�R����TNE
���.iu�j�/s�pq��G\�~`;J��S���w���޵} �Ge�����d;���Ŀݞ6�E�3�:��(�����
��g��NJ��/)t��L��iT�g��s����T���������<���nm�m:��z�� ��j�����B��1e�*���9�-!��+��11a���������J���C���]�ݿ?i�<����DɁxC�Γ���>:1�PzJ	����Յa;t�.C��]�����Y�ua��[�1A6� R
9��4�X$��LR8�`��4U�?ߖ&��*��fQ_]���r�L��j��� �k/���T\�kv��O?�}M�en���P�0K�̟򒫯��O�๖a%�lM��>��5Ả)�e�oU�X����B����}o���Պ'�sz��<i"���!�/=���ƣ�F�����:�M�������1ѓ�l�BՕ~d܅W��'���wL�D(���WayL~�q�W5���3Q}ҋ�QG]�Z�L����C�Ї��o���d�D�a�,g��������T¼�m����P%PS��,�$������܄iz��
9=�T�"����͉T�A�6����n6�����G� ��ΐ��UH�]���M�'�L�A��:	�1�˕ !!�`4�z����c��Oe7������oA%�
���;�,�s���na��n�N�O����3-/K.�P�5"m��'��fB�}>Q3&����~:mϽ����}x�άb�p���b����ц������MʯaM�'1��L�5��A����m�+z��X39�rH�Vı	9�N�ƪ&2�`k�O�J["�0H�x����//l��0�:Y�lY�9�G��/Y�}�[��d���Պ.�J0)�\r�"��y:;�<�M��MzU�w�ᇡ��\�٩��/��x���O�/�J��k9�f�1���3��$`����G��fрu!?�O�&/GOj;R����z��zY�i����ow�0z\!<�,��U͡;��
U䐥DC6Nc������c��Eg(�G�N��F�m�i��������G�N��r-�ZC���EM̒�(H�뗐M�c���4�`�!�������V��X"��xJd�M��t[�)�} n{����2<12#���!Κs�A��Z�z��b ��G�`���k��s�I2S�b�����$�ps�q�z�y�x&��[��!�Ϩ���}8R���������]:�ձ	��?���Ԗ��]䫙@�����'� *���Ld����|cnJ���A��x}�&� �MY�}�p�;b1�D�7������^�F� =<��?Հ��0�l,�	��1H�(Al�zz��$�e3�0�\�ϊ��c���-AC��Si&h����7�Q�n�=T���v��|@t����!/�sFψh���o���8W��!���]�n�3;����P�gBp?�Zؖr�@��*  �Bu!�:�O@����TG[���s�'�������p��<�<�y�/N�-JEu;�F5t�N2˅|���/��$]6���\��^��H.r}�`Ѵ��s�_�d�Ҵ���� *>���дο�*C^�3T0Yw����@�Tw�3�i���G~���&�1�����,������`�I탘���(˲ـb��SA��5f_nPfP;���S�,%��ų�iGg�Fo���=��m�v�j������P܋�H몍���T��/g(��1��1r�Օ-�Z��,R��Dʅ^�=��ӝ{��Ψo�B�L�ե�"kn���6ߗ�3uUr�,�� b�[���ⴆ9+��ա��<� ��t�bKQU.�:�e{�;�"(�8P���M#4#A6Y�w�:r�vd[�n*�[��`��W*������7��Mi�q"w����N孿-M�$گ��6�OD���9�cQ�3�]W��?�U,���T��Ҙ�q�;'I$jj>Frzۨ�%�-�)'��`*��i�Z��p�!]%�7��0||ݮ=�i�&���i8M�0����!}�����F��.{��BP��|����Н��c��]�F�I���0�����ZqX��yn�P�cQ�|���s@�݈S\���b�
rx�I,K�3G-�d�"��;:w 8�na`w�?z��s������"��U��� f�F� ����N��L�S�G&�l�Į5[.���+��"�엲 4C$B�Yf,�������x��~��0^�P�:�y�ȩMk�����,�$�C/� ��^듳[^py{
s�ç��Y�T�Q�ҷ=9�-�~ (׫�l�=����ZУ�Jrݿr�P/��o�	���<�llЕ�*l�7���|}so���f�*R��c�q����1��zsS���4���� �s�.���������ޕ|{,$Y�T�5#��~�u/lc�D���G�k�����!��Ί�A`��J��Ȭ����Gj0&���0j�wߌ=V���.�>�O��Ǘ������3��m����UDz�:t���oC�5�m���jү��d��2���m|��J�#�Q��Uz۳�ќN`��q�b�1���5��I����Y��HT�xq��e2?������ ,#��áx^X����]�g�[�
�R�g�a�KeS�������F���(q�����P�=�)��z��8�mW��=7�l���.�u,=��KT�{�3~��-Wn${�
��nU-�65�ѷZ}tӰӬ�k����+NC�aZ��ܛ�?A��� ��x�)P��3=�O�6�Z�bXd�@��c���q���m���d�D�kT����^���z>^l����;%@ϟ��*����M<�h��q�K������@:�+q��D��h���cǓ]3D�B�MsgR�d�)L������h�eF��H:yZ�H��{$�M�J2��������p�>6�)���Z�p1FEC� cԋJ� ��/�� O��Y��O e��V\{}��3��J��)>H��!�R���@DM�z7?6#r`"0��c��@��C��8 �D���,7pr�c(	{�?�{6s�e�G<ې�����>O��E��Ot�%��q[���;'*7%6ܹ��PY����W>�#��޲8��&]x(�b�*����8��9��a��o��ņg�
j.X��-O$ ^���l�<��^j�W���u����~�a凧<q
�`���|�(X6}q���]$ܢ��蚪 �o���u'l'b?ho��˥[��߮�'fO1x"	v�w�%^��M�Us�������l^m`��%	=������{l�2���露�n��-�n��8�����~�ɢ�]�y��{���]Ϛ�{�_���n��n����&�����i�����{�[S��� ��\��oF���zi�V0�#�V�D��E���@�N�;a6^�]x�1;�{��"S>�B�C�< n��B7��T�mm������e�R��9�x��.��o&PN����_��j��`��rN�O}|�S%���~U�����:TʝG��;�RO���7>�$9�kf����n�E�XD��~f�N/��I9nP�Ʈcn�c��e/���0<�Mh��;QwB�R�fR������:,u�Bv^��R�v�|�/�-dЯ�-�������<�S��
�����+�bw�onI���cȯ?�@#�^7Fv�|{O���FvȽ��Ah<�A��PK3����ڎ��F��oT�"2�?Kvw��V	�ۤ�+�JJ����3�,�P ����iz�i-��ܽ��%��)��mvP)i(�d���3��^Bzg����$<A9�Q�%T��HOE0��W�[9�������t(Ԑ��%��1xe���=ݸ�W{��0V�[�y뙛T��b޻r��nO�H��
ܕ}c�N'"��e>�����\4�L�oh�+����P!%�d��I����$f��@�_�}+�<��T�� ��|���>qo���0���p�r���A'�V8A`E��}�X�Cÿ�*A>s�x��0��\?ej���4�H�F�3�=ev=���\;ۈ���+�h�B���ssmI:�Ty)cO`Yw�>�n�m?�*e�����r��C�H�~G]�N"}��,�a�&Fz4�&u݉:+*�$�W�H�@}��,X8�h��|�QEmd�R}��a=�Ϊ�D�ê㊑4���v��e�a���������{��Љ� �3܈�V��	�#��X -�D*g�x�)ߧ�锰�T><�E�Y��;�v�Z����Y��ʷ(��.�<$:Bl���X��ǋȦ��ԥ���)�@6!x5휁a~HY*����μ<d
�N���p�\+�3��ܲ��l���B'{��Үg��e�6��k��C���,�D�Tr��6�|�^SN'Mfӯ �.l2)�8a��e��f�q��O6Y%�{��o��83��>�x���C�����эK�C���	�H����ZwFSI`>� N�� �h�h)�~�"���:�C����lk�m��SRo�×�yN̅�+ώ�k�)�f��
����|^��'��f�O������u���n���0ʒ%z6y��bWU�����5\��?ɹ�Z�WƆA2�ҝ�(�˺K�V��ඏODɯm(�!��(�YZLF��P�w��|_L�5�Z&ZX�P�����}B���ڑ>~���V�4�G`#��5*I��}?5N_r�����,�;����P��C��Q�������>�񏒠Y?�����et������?R�"�C�h3���X�3xێҌ���&�	�J�K�}�b�y�����Z,�e�d�0��{?�wK_�`0R���!��Z(k���*>$�s���N�i����@�mJfN�&gߺ���轙�D�-�����˳��ww.�w�5w���s�2�	����ڈ����j�VXIA}���)��/�(�����|�!U����@�"�C�S/��gF�n�K��U�a'�N3���a3���'�d��*t�FS�N����<;�C�J�1i1��z��8����^��Z<��t� �﷬*\F+�u!��i���w��
ۉ^0g�<A��-]�f�`+��LG�{d��_�"~(�Lt��m8��
ڍj�-ZFǚg����c��	��s�y���5�^S~��L�߼x��!,���b4�+��� e\=�qi*����h��7�Ǯܘ^jlx-��8ItW�C*��@�|��Y�j�1��u���ޢ�a�-[�#��4eT�[��:�Zz1�ëΊccFE���G|��Q�gD�.K���9��tp��,-���~��V�XΫY#q�/*ZEsV�9��6>ݍn'hZ�xi�����C�*�w%���I�
�Ж�d���s�%F�	l�Ȧ�+��[�U���&rn-A��W���ħ�B|���`4(�J��[=�1G�A�9�)v�c壛�<����j���KW�j����E��Ø��Q�Z�	����e�mO��$� M�G�uߧd��
�
,M��g��l ���A�+��uC^ O�)>��u���ѷ�C�iWJF��9��_�5_�
�g�b*Z6�7����`��Y'��8�'�ԃB[Ȁ���ea�]7!�SR�$h:h�����@��i��@�$��wC��������h���c#[���z��A�=�"~2��/�r�7�A�6b�F�3�s4ቲx�.ِ2��yH?iô�ہ%ۮi u��\/C~��<�,��oSu��y�c(>X½ZM�˜'6��A���j
��@�[C�z��\J,��oU�l����A1�IJ�`_�w�C*ĬwFH��f�L�MY���8�+ {�Y��pD������oL�2����׽S��nT���B j1��R�LS���t��Ё�Hσ�'s��_�1�y�]����R�.�M�����*���J�dL�����q�'�&'����S#>g���{κ�/ۢZ���a�Fy�m�PC��#��>�;%�<Ÿ�R�x��[`N��}�0�8�|É� �2.Vg���h:�W��} v`���=�>H�brW)��M��0�D-�hYw�^�D(�N)2�A��n�[,̂%p�I���M���YQs�R��k^���F>����鲕�'����k�k��w1e����W�vHKgџџ��cT�"��v��p�4A���(�������M����9~H�i9��&WlJ3�ڋu��l )
�; ���5� x Y{u��b)�ڢ�x}�g-�{KMq�Dm�c
�J��{�p�_�Ƞ��ËS���O�17�Ac|�c��p:�2����k�5�&�))Y���*GD�P8Re�ܧ��0��D�Uzv�L��Ʀ!������0S~	����<0M�ƭ9�0���9���}W?�Ƹ/����lkڴsT���lAE��r?�4�]�H�$B![Nn��g�W����z]����=LGi5H�nF��>T� ~~�Y1هRo����.\2xk�֯��
��Hΐ�69���,�Z=&?n�&��yoMN5/io���u�uk���ni��cf�q���n����%3�҇|c/���kQx]'�M)?���ۏ��'�&Ԓ>(ݖ	�����N���#Sf`)�2O�x��v퟼<lU6I{	�A@X<'�w�"2%�P������6h_�o�<���͂�ɫ]�<�}ܲ� -�A�X+Xq��V_��`7e\��񝬦�>��ɽ�����]�_,��| 9��;~��.��q1�7��=`>�lȨa���$v�B/F���_ Xt`fǎ��{�%�J�����y�,�l�(�>��	�W&*;����A�:���𺮙�Z�+�rN#&��{e���{P�媤=�zVP�#Z�A���Ӳ"K/�J�L���������f���/���R����B��p-uD�%G�&�e����C��ft�.��y��`5��C�
aPݒ��?�Im}@�u�n�0��
{��"�}�id3���5.���k4��55� z��W�CN��h⃪���1�ተ%�B;΄�r����y؏�%�M�?jQ��y��K��e�# ��k�����X�n���;o��*(�{}q��J�����|,�A�~�����O�C,��N�������4�DB��}q)�� \̙��hk������K
I�,���B�;D��}����ŋ�WZU��}��[�d*�� ,���K`���,�_Y� 3�md+�����̍��\��K6�#V����a�������>���:֙�Nܼ�6!����;�;K��%> `�T �ᒿpb��ܓ"�5Z�9�A��(�@�ӏ6�_��B#os�o�G���&�2���ص�?����lf�`��$��GBܥuH7:3���5�@Q.e�7��~�Q���%U񦫛� m�g�}6/��)�RTN�i�I��V;�����1���?l��DV�w/�@��!hñHFq։�)M7h031J�60Hcjk�(�!ԁ �`~t���Pƣ�ruMK7pQ�B�	��m-^�ᖍG�Y��Swј��~�
Z�6���Z��Ȧur���ƾSk_V�D���Ϧ���H�~�jr�+S��q ��`T��I�5=�~-T���
�&�XQ"������f�*�#J6��UJ�۾�k�[�^�8~��L������������Bs��=�r�3����j,Hڢ"	���TJ|$:y�۰>8����:N	�Y��}��^#�gM������k�����96	�5�?ymgG*�A�cg�16��z�q:А�ǲW���&*�7I��|!+&���2�Q��GD�ztt�2�v��8@���L�n�l���F6�{yu�Hq��l}#'wY���f�M�#�Q~�[�]q�EL�ԦaЯ���Y�b����qח���CE峺�}f��[�Vr�]�Kb��f42�"���B��[k6jϐ��Jf��K�A�Np׻��o�1X���JM���e�K9w�&��ISE����r������^O�6�=��aǙg*̅���/���'�M��P���FY ���1Oz���=�B4���7����˝�q�F��eך�̮�
yxj�j�"���v������0oJ"��a�Sd�!�0d�3���>;�j����3�]���%�= (���k~��42l��	}I`.W,�m�ijA��n�\>GO�lш@N�H*5��פ�S��|��5���J�r���w�~؊b�9οk��� T�����1-�q�y�LUSE� P����s[oϬ���O�	k�Q�Ǩ쓃ϓ$���ϓGc��r�!���UP��ɋYJϏo�c��2������}-�'S����a�
��;��ދ႑�IS)V�a�U��KS����>	%���H�@�+����	y�v�p�m|���3Ѯ/�Xrc9���lN���^72��0m�c4G&��T�^�<��5E"���Ig�P���<|�ٛ���Yi��/�7hě����`�j�څ�n��Q7=@*|T����X�ZG*�#;v!X�$����<rsa��ލ�	�m�}���:�/�+2��]D�C}���J@R��o��x~ Lq��;�d�l�
�t3� ��^$Rq(]�-܌߄�(,3�BϹ�M/ac�#�~�LSٌ��)����/e�|$�u��j08҂4�:�H��<��)�ە�AH�nE+·�F� ��x�r�bm����5��zJ�>C<ȳ�w/�9�RcF�^�|���A���n7q5�h�7~�γ��G�u�Rj��9f5�_�<W��}�*<(�}�P�5��ʀ{�:������	祪2-��.�d��]����g���g��p�5����~��<���R�%%���Xt�W[�ȁف��)�	�l �[vC��̆�C��J��������c hd�d��٥Ft�h��J���ޛ͸ڍ�0!S��eP�}%G/� r!�<�_���� C�^`��9Ν����
k��}�U���b��V
���n���qؕoi%��s�n��vt��,c�|Ly6.)ã�L����6��v�{{Gn��M{%��Ea��2�6ʖ1ja���o,�*�c��%l�]�c��~ߝ ��TSi��n+l@aA�v��ձ���L�~L]��n=�׀��e�(��m��7H�i?�,�F��g���wc �f�SL�B�?�b�~���3m�l�����Z�y���s��d�p �)��D����.x��s,�{���0z���I +5�I���!h7�P��_"�J��M�f�(�졸o�Ş?��~���o����ta.�!�؇s=����[RE�+���9��@���ۺo}��0x�^7�T0�d:�Z� N�n�rC��=��M5K2�������^D�F5�$�8柟ޫ�w����6����ud �O�
�Z#zx��yֲ�����=�W�-"S-��f;�~�"]�fr���>h�L��3��˗��}�`jߐ������PU=T� wI��1���ꐜ:�A��((�)1%u�`uo�AJ��А��) 㤧��X���]�m��TiA��� ��)�����h�ΥWq��'yc�a��9�Χ_�2����uB^x�W�6��~�v޼%��j������b�M��O��W��(z��z����F�o�|����L�	H�U�W�jˤH���[YT0`���Zut�!a< ��A2�����_�蜥��yT�C��$��z ���%	�\>B� gY�,�U$��7��@�N4i���S�����2I(J����2?Krl�4�v</�����m]��2�mP��)�B�1�^֚�Y�O�X�Q��W�k4�-������G؜��{,��!@��-��E��[c�D�����Q�ha�Q�l�w:OS�����i5&lF��]��UJ�O�.�&R�Ο�����.��Voٮ`HW�[e@/���DUw��LwL�X�<	%���2�b�P��1�Ϡr@@�|�k��D.[eX0���N��l����:�$,P:�
8}\��%�BY�c@GZDb�ƅ��?�R+m���m�o��)Ƹ$S����S����v_]pa��<�3GE� �v3U��Y�V���Ui�]�jZ�P�?u��<zm�Q��V'6 M��u� �$�����4�F�%iK�h�vP	���\�`@0b��K7�Q/�!W	N(fz���[�m�+]�9>^�Ԏ������"�>'������=G�L*�������Y7J<W�}Sw÷�B������$V�{��6�IO���Y�T��1��s��[LF���	Yq�C�p�8���`�0C��=�v��|��u�����Zu��6��m��H�&���#���ԅVf0�9¨'�������Z���� ~�F��R�5�!J�A��.,���a,��{�R��ȖX�2(zX��t՞�rO�����u,��Tg���:|N���If2������E���b�c4���#���_D�m�v;�g�R3i-E��\�K�02�q�\�9����+|��(R�׷��ޅ8F�u&�HZ��K�[��
]�x'y�;������ʰ}��j�:`�!j �����C��\��Obm�	4�=��>=s�Ɓf����aG��r\���w#�3Q#���uc6?�.\�Q�^$��	b�y}R�>�����8Y#2h��9V$����L�����N5��.�Q'���=�����6��|¡1r3��2�76(����>7�1���BQ�1���s�:�%��}���{��ZU��<MZ�=���g��b��1��E�~��Ē(kW�Zo��j���Ai>�+4�*�ϩd!E~B��X�3��2�xJ����w���q���Zug'W�-EjY�М�7G�\ÈX"x�7���<�M��D�S��2n��M�N��y-4�Qw$�K�Q�E�cw%� ��-n��י���q��7����L�v�����y�O�{�(Oy��QĻ"�4��	�5k̆�c����硘�:'�ИX#�^oo�VS���d9���D���!$������f_A����tE6g���D����6'G���?����Y�r�f���y�ƠQ���J�7u�ܓ��6�J�|cK6S�F7M~��@�e�y�ú�1)�#yq�Ȅ�ݔ�<^�I	z�M)(� yq�9~n&SP�{Mߠ0֯>Z�x��U_���\\���~ ��DQS�H��U2O`�.f�3&�dFK���Ĺ6����5@�."J�-~o^]%(��Q:f?c���BN���O[�R�?'���X�>Dئ�B/r�4��W�0E���y�Ќ�xsKͷ�E!�Ƣ��Ny�LHRC� ����^�P������z2�Yk�	� �d�|I��Y=A��`?���=�'��d��FK���O3���f��o�suA'䙝�aܚ��lY�܌;Lx��U�S�l*���i�|�Y	@��F��	���v$���R�q��9�̵�k���� T|�'���&k��W��a��}��k�].,F�����K��r�(�GZ{��%$���&���F�ozGWR�r�r�hE@qK�}[ u@���� @嚅M�a�[5�ӏ�G/糥�+fC/;�n���}5����ꛃ7�8��T���Q�TSyPv��#;zc�-�̫k�9�rZ�}�M/Mt��r�e�z�2bߝ;�O��f�PP���%k�3"C�Ή�ga�^���r5rٮ���6���*��@뛸�n�vR.5��	�@Q��߭	��*���9@��7ϙ|���=%�g\Q7�yi�slF��] ��\&��y��-��"�������E&:� b�Vf�q���P�b_ !��/��R��>��E��=��,(���<��"�%2����-wa�����9j��x�k*����(���i�\�ϵ��m���CU�c�w=iZ��	 ��<����S��36};A��0�&2���x8^���#q�^�w֗DPd�P�i8FC�͝�G�"����d�$��W->%i@���� ��X<*�:(۽��y�T�:x�ǉ�LKJ��o!��{�b�t�	��0:tPDpe��{���/W��������V��F���H�;V��1��}��4|Wz|�F�0�oY7P_!Ǔ2����m%��q���?ʷ�#�)=�+�S��ҝ�Cm�6�6'�;��vP߾^��*�ww�O���u�G9�-���d�Y������'&1�K�!z��	Ʒ����O,��	��j�(���r&��|�k$�{HM�K4��eԐW����G����*h�y�4&W���� T&��$�Mݯ�6e����8�B�����)@��ݿ����U���[��:9_��~��C�ٖ���d��ѷ״�a��A�<��qPAH�;�.l��z:�[1��$�կ�R�:��R�I��l0X�o%2zp�5❜�Km�'ws-���h���U�<	����Uh֙��}cK3_St����#˩/�![
�C�#K���ۗo�E��(�E�4��ZH�_���6[V�`��A��+s��_K]�S�'r��C�)IT«�l	���l]Ī"(�$��  ��]����>k�Y"�v�����8�,O��!NY
��xI����C�J��3=6Y���^����� ��@8s��Xպ	e3�Z��ou���y�͘�.��s��=���k�����,e��`?!�F�L�R�z?�[���c<Q��CDk��QL~����M|�=�A݃|�GF�Ð�-�f�(7�N��"eU~�n0J�(��r��b}!=:�;�|ː����Ǚ�A�Zgħ;G�b4j���Y�h�`��G�rw#Hp�!���%�w�]VYX��߽�����8���.	�B<B�d��ćϣ#�.M�})�P�ξMb�<�H�-!jӧ^�t�xϫ0��\l�y.$�:!�Z��Y@�y�j&M���2S�&�v`D\�T��cq*�5��lC��vZ�U��xξ0�[g��~��+�_Ȓ'@R!99�`�����>Q�~쟖LX��`���%P�7�-�ymeR�*�����E �a��e`�核5�o*Ճb�K�>���6kV��d�G��Yᒘ}i�K'r��F�_hЅ�z�p��߮o&�w�RB�V��^'���[^�qhXҙ��h�����u�t�X������B�����v;��G$��?����QW�gb[w�j��0�l�^,4ܤ���*T\��'�C�ȅ���2�C�>���3�R�c�r#�-��V<���/�b ����ߝ�黒�wa���W��2�x�A�]��Nȧ�#����來�=�M�%������
�i�n)�Cyv�Ӆ������Z��ss3V6��<�������2Zc^�}@@S���Ӿ�n*˱s`�0+|��>a�S+A�/3)��c�йT��~�f��c��1��
��J<�t�A8�8ޣ�8�+�؀��_Ԓd�Ndw�|v$v
e�?�cl|���)�f<��w�s%��Ջ{w�/�X%������J��Ik�R���g{	���0��ᤗ��?ޜa�O׹��B��h��ߵP��Zk{8�	�e{z��aA�"C�/
�Z-������\��PnGpPE� �
��ŢP� u�~�@E� }���\Ҭ�2~Ѱ�Ϛ��<���"_�-&�쭹�}���6��n�}���N1���|ض<6!g�<3���^Q���:��>	���+7��K��g��Jsp֩���QH:���SI�Z~��|B�N�u��%�p�'��0��"U���T6�KD�7�3��&XsB�꼱x�����:Y���xԹdQ&=IP;0�o~[{�wTY�1}m�W�w���O�7�D����O\�Or#BX�6��Ԇ����`C	2�b�o���[��)��*��|f��Ḷw�/L!8"��J9�M������9�Z��d�	� ���\j���N���p��c9���3$�?{��,��o[$M�5e���L�K>�=@h���8��"K!MU�7���H�I-)�����B�ƈM�3\���e�n]�5��oS>D�I���iSV�q#���%���e����y>x��+6 #rf ���-;�d���'l��C$,,*v���]N�����˛�&5�s��+{��[