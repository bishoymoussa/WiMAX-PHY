-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Hwnb1V6OkVjqXSt6aUlrYNWhTMgv2irVy9bYgNn2VtuT+82x19vxfnTRGs97mVK+WzSlGBfzlWMx
cr2R4Dd4aT486j6jatUDbZIZ0EV89F9c946Om6JnVM8bf0VpOjIGpzSkLBC1TLXva2Bkh0OuRhgB
/LSSVDdzBv5AHaOKmbcDtnGcDaVseNugvHdnutiiAX8Tsd5JBCg3G52Yq+g89a2sBJD/Ltfi7KJu
osFAWICMlW87mpKPCBcu9DRBftlGFqgRGJfiplI7OYZgPBK/rhnrtqoI9jThNyrQMZLpj23cYsVd
EKRuQ5MKO6lidbLvdtubzhQ9ADyuuuIn65FImQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 51088)
`protect data_block
vubeyEZbyhKYW9PhU5RuO7bmIuJoXLPbBMW2wON/xF1s7uxEe4TYR+nZE84+8Go1YuV4LPVa5Fwj
j74H6KDOPdGttOFw21oZ5K75kpcfcs3GMx9zkg1Anz6dRUj8JT1wwRsqglj9r3v3DxiuCVztdsc4
rSOZeIBgwsAfln4mp/BnDJx27OF9ltDx02G6/F9ROwGRGmugFVodwL9o/vpaMryT+rgkH1FfxKLB
or7F4ykzwz537BG6cg6cEct3AWYECdhpIETG2CUUSTQBUvJ0Imc8xbxJLZC+q9oKV0PwEr9dOgnu
405Z3ihyulAEc2NAE1D9pogqtMdqYNODox8UKf8hdj3uMgN5wXtuJRa17BTFei0KVpbxA87L6asr
XfDtzOHWV6KZEPV+2KbpqrcYUkIwG8vPNOLZRk3K9ul6fQ43lwryJvBmRPr2SeBbTHIsc9iP4meh
uAfaBgolsnpqZ3VjHaDbU5AiIA5/1mlp7skmpk8VfdDYcyeKehRyvgC59Tqoht63teKw+56JBx/r
yEIvCQYjwjAysCWDXQ0Dh/q6CAc0FPz4lEswsy8PsnWfWjHEHolX60a9Qs0lZfvh885Pba5WPPiC
vC03QnYSweIi6Gw1K6l8B6H6d1auMt06Z7mEQgojzMGeP28mhTu2ZOXjBkxtCJnnLrdZCauP432W
+m6ClHuJbMgOTi710bcUf7Pg2BcfUqoMb/ln24LPS7XgRH+VyQflnXKkyBxbOpN+oyM9ySU7pquI
EqJizKNU9YrZjGj7OhWvGZLKNZSAnyusIRGQzwRYzO7xeH5EuGAf52fz/+oKMyu8g5inXQlEUNfB
e3g5QKDk7u4HpZTzcWXIMElRzTYmsC3xhqXIMEmnyTUWalDPmYS/oGBXPlzV753hwcYv2uTvpzIx
KQZcVamqKkcuwjgSdOlgji1Ac2avmxFvUAfl1quExH0E8ciOz8qAuQVC5WFeh6Mx355g5ysYMsy/
0X/9O58kCQcbqxcxReu4TpCkGwH1/9ZLkfc/waQoim94znM4mrQyOwO019yXtLx0Evov9eLbfJcC
RmbwkMOFNId9DgH3v0Xq90eDkZp5gsn1YvFDaqgOjIehw/+1p+Ey0TsoGvPBTwg2fnsOLQtuKIA9
5z/S4qt/iU345ccGp2niV4/WMY6fPmegruxDAjYMlGoaximgHcpfRzU2Lju5oMml4MgauKdnnfni
dvu5ifrQ65ggd6PYWkWFNxi/e5PzIG7k0hadoh2WXFp56SuJoS7QSPU8uALOVqF2slKA8Z2K/YdL
MtG6NRno2JCtIJBuqq+1fEs2debP92s6u+eiUcBznHlLxY7WvEmMRTdxjbGifxs/xE1X14nFLQoU
fTxtoBVURB+Gfb9oCmnB898mhc5Ge3Wti1H7JvkZGypMCJVsgOjmHF/BQLAykqj3ENBZbeasNPVf
cjSouwT8mowN4hd61hkdsLcmUqA9+xAqrLt1/cLTX8JgfVN6o14XqHUAVy4iE+41ftV+rrexbAk6
gEb9vn5/kOAN0EIlXFLjLr2iOv+0vSFHCBCxcZmMAFMRDXLogZy1fR8YCChAO3BGRIxzRugHeioR
tMVAMyP8ZdljD0T4G2ZyK7u6oEa1AkvYcz0Cf+RJcLynL1WkknU2+pNuGWYP5Z7gK01EGOFi9gUl
PqkuzP8sxCU8e5FdQrjaQxQHPkao559idlTinfHyIR135Csjxm6k6QmI69QBePW77QUVlB1DVyIV
Wjh4PfIf687zCQZjarq0hfgbOZlAY/M03CHilmHAbHhWm0VRe7ShgXS1Yn4MfcTr01/Ixkcjf0kF
JZgxpU6AWmqii+eP+/s6PTb8G98+7V3IdFS+w4j78K1CvE7DouGCC7jkEIlnFgxdAR2FBah7Z0wl
GrqIkwTXbhJYvMKHl8fDUPzmkAHRAjy2jiko8JNeJd3JyvohiZHhA5tt3C6NZy3+dPE5j3f3zClG
NmvN2Mp9g2i84JlxYwnDUqiWU8ZlV3OpQ7fg3/ZlrU72L5rrNaAmc/pr5w4kBV4lEGWisGPpd+FK
VnToVyOepLbPuGt/k5KTkoP+bLfmH2jx/cU86wCu4Lbwd1WQYP8LzfaSS+v1tzIqZ10xsgpCta4X
lySMZDR9yFUYbEy+r+6zP31iX0gb6xcWBsuqmSDQgjIQxpcIgWgHId5Kf2XxxB8vuv00Ud/GyGf3
Uyl+ORwpxgKIQS7rpjasGygnY+as2UbaZ5pOKlndwck3/8fEDWM5LsHqNwwyb28F3lzktAVklGhK
8q/xtD+gGjWgHdf1rVwlfn7DVE+2CCCLQUTgQc4xcE7/LHRKQcEm4lKwX+z46CEJU3gK7+ifnPYz
YgXx7Hu6DpugoQ4pQhSJ16duebOLm0WUgEFmEF8fSMGxB8N87NVm4FwUiQV65EpjTViO0C2fMusO
9Z5z+kM+RxQ6Hgzt24kNZ2E4bo49cMB23e2OZDVZUnrqsbBO9PvjyLGCIX0RdHFpjBE97zulEepS
dMnHWMtGfignK19F/oM+1sZiL9GQHKoeY+gsJv0CMHoBMNSccyp7ABtTA9KapFyn7ARcxPRBO26G
BIOoDeRU3lzE0QZOPDLoK67AISEHKRDMWcWuXLV0DB+S9wU4ZcEK1OteR5B6IOEhCo917es3gb+H
IZXw+MyVC6K1W/f8ozvuUlrzk8ui8peXKGcd0HAT+bfRWF0aIn9RS1XN3H+VKX6mN0Nd2Ip48e08
HwBjIwPjE41Su9DezXCqNA0QL7hViknJaekpWBTV1Uli6a2juOyF/3tfG23ggvB2V/XegWpP/CTm
YXse7bVnkAlQUaH1/sxa6OKNZ7BCscpMMzZD/+VhpEVqQePrwydIonC+4EqS/O3ijlE+zBOAfX1J
uPL1oYptZvfR4XEvsPraAuO+y9c3pQ0QBA1rMD1FmvUglhLCsQDLHRA284p2g5jQWwavZlxN0Z2K
nrWGLSFmGXFFZvnUoCLrI+Ogwgz3LXjKjDBQJY0kbTwWNHQrgJXCviA8o0bI7myBftvQ3nYEcm36
+1q9xG7hMhlK43AKE5a2gJChleIUq8odZBQ1rAvAfkyytRbPPaEKcv2FgYKuBKKaaEDoeextepDv
FAJ7pKWQhOr5Isv0u2bkAzt/HV790ud9seSeyROufTrGN9tO4hLA9EPBkvs7AmaDDmY6/P1gbwBY
2uENpkaFF6oCKywAaoFIYYA8BCyod3c6NyXSn00zY+Sg2AW+QXDm4L+w7XUdltaFJvlaFPe0pZT1
3KvHJBNWQZXLSGe59GL3dRLVnW3rGI7/3g0Sn6HrmkAYMf4dFHvvs/W+PK6gRsfmS922QurTScX8
xs9QjnZ3dDRONRulwtsIE5GrHd447XmstVR9evWqNrp22FsfNy7KDPMa4S/9zbib4Bn+eEKtO25I
7mP7HUJjDUZGLMHHz0nrcQIfvu9COjgpEAFgaOV/XqDrSnAw9XWI+OX56NwSyhTbdo/xIQK+HaG3
mxlT8GAgCAhj7Yh6YGpMwEYPHz1mcVNwn0q5JLyYOxiLeUwBLQShl/aUGD6571b//NKRdZn/Lr2V
Kj4m+CvmqMzP6G+oCURMPoAkJ1Rkcf1/8N+WGx1RVPSyxCB/2xru9VUXZoLsH+DNJYDvKGidt6XO
dc6zLt+VjTvMdF6OuD0pwkn/IQMWi6hq+i1MqDe6kztbwTu64pd+iuBHN5JM8FZ4rRbNvOGQZyk7
Wy5dtqMudhC9nhJMvy31i8vzLCdTRhW6yP+Tm6xedGxwxnbtL8c5mUOaIdELzNhTU3PF0y9lY5xS
GdGZQj5uP/bAkTa5dT49rOytD/85l8SXrQElvM2gJXLxMO7E256o9fMIkYJqGqdUvTsITq63iXOZ
QTmMpSQxcmkKy+INjf/CSbxOWIUQhra7UmZZm3p9yHdSunB9EYwlr44dN5oWGPNSgTypbqJkMGBY
KzTRirJVBxJgD5d+fjST/+35ZgNbvh/OdWeJ7cGSs8Dr4XStbIHyXTwElPH+LlgdYGPl7DX54qRw
1fPeP7BPoydJyzAf/hDvLRdGrZFj9S8zOoi9WtImuSKv0/fSopxJhDSh79+l1Qfe5juW0AOKNFUK
PaGvEwSu1hXj8P+dnTvIfV57W3kOFmNrAyeEB0eK2U5kyniDSeePJr/57Q9aiIUaUzu7EiMiF9XZ
0+Vt7zT9g2XzbFOdjasSOsSlCKbZlWfn5UXiacP7VxlFTrKSivKj4n6zVnlvjS7DEbMqlS3lkSyd
QqOz0GuAhLoaQ8ynsGlwlYWoT8ITY+8QJH3F2kdcpYtJCfi3VTRJBFW5tKgv1ZEafKagszBOIKbH
X+XAaKLsZxyi3xJc4q2thnLMeuNRXuACK2MEohbjSLI4xKnSOmw4lRt080g9z4kYNl5XOhpHLgdG
oZFFPWhNKgYs4oF4NVlO/I5/Euwi3AHswaCwwez/nrJ8Zk6up2Mkq/mQA8jRTRlnYgU+pQJdJp+3
A0N5kVMGCWFbEH+x9IXo7DhyGPmUgU5gEpaBGOQkYSdpNa/RnJ86vRdr3agADlKUitTNF+9vziVp
g+LKWgR7Jwy+7UP+//IzCXt4uPNRhK+BCqEpkNXvJCto9MeHaHlX2+DpAA7PpBxvLQDT4eChFtCf
z1H/uX02Dp8SrZ3oxOayCT+Opbq1tL0pfDtAvBnS9Mt9onsv93hx9LYEJiGsAFdUQgyU7AyLJOEp
FVGlYm6/aDjooox4OjHIWxyXGhm7sFPCYhPQ4mlW7OYfnKlTxf1P5aodGXhMvDpf4Ce1DVQobVCo
amMJY4sX2lls7zMF7IneJea3rXwDFA4/yvhPQ12hrwLRQlJUFDYPAxfKxJQPCPpzsREaYYUpSl0b
nnIk+n7/wUDl+6q2bi3LQVsTV0j51URoI+mAT6G6a8NW/74HrZ0m4lncj3hXjM8zDcS/s+ug9avG
rFurFvaObZSyc6daK0P0QXxQLW5sF7XTL1k8oHW1bz7cO/bv4Jll+11NiAEtANCuevEjVqpUoaSa
O/FhEJXnHcuFovb06O5LVSvyRYpJwkU5Dxe2mrMUfj6NWCSYZuexqDuOZ37nJyAR/zzJ1CEF8oUs
gZepkW7/YSjw4lmXrVoNxtxKSpvkdfqmOv3ynmSBt9JQpb0dqLgqktdLH71mM6ij/FGJ38HHwKyX
DA5jc3oERiBkQiXstLBGW9GEe8x35C7l3AxaSCjGIy7eYAPkPEnAxSyMcmPLh07UaUy6s1vByPHf
ceUf9gC+xxgjet/sURg+s5/nU0Zp1Nd4Mx/d1C+HSu3s5B+XASoqSh7t5vrRgwQMQA78uRcmEI16
NEZO+/Nt2hVwO+E+mQb8aCbJgjjuqx6m2RS6qre2F6kUgS1m9RBRqdXjtg32eGnyXc0PJeRpDX6x
5GfD1iaHU7Ev4VQhvh2ByyjT0reTQ+aDS5qcwiJ/o/27lNUHFlRZyiPbAuh7n/IduiPkAimXuYPq
+jAN5Jx2HPBc3SHD9tC4T6BH+kIZbqhpg1oDD3dqU3ak9X8Q11OEkO8Ndu11/8vyF4nfGiFLoWBx
b5dnDFA2cRtRKEf4wIPZok/Grvis7SZ7IymO0GGb+u0R5uQpLgxlyRQmu7jWORV92/hWtidlo5Pq
KRdeEQQwcDjpOIhQoD7q0hr1iGgg/Ux6nyjOgmqZl7B+PDeYzQpuRmEvo7DQOIu45NkhgQ1QBn9e
UfBnbxVsHlo8sRb2hoU2brIyv4cw7JQmk1OeIfvTzP00M3ZdsE/Swsv8vPO/tQI2fp88SIINg8hQ
ZEy2lRfaf2vV9onPjHIFcadAwu0pxnde1OqOlDLy/5xR++KTbxdhSLzSONL6V6wPTIwQoGKT3vVe
imjuDAdSy4xiX6M9BrzRsUEMc3RSU5mZ4++Fr6qqS5PHiauxaHAqgJjperRidMKA2mEp6c2JO9qp
oTVVGztpIBfWjbWRdnUKO9o238h72cA6OqUdSO7Odx5JlatIAGCrSOfEAMpP2M2ZmNc+j6SmN2EF
3EZDQiQ98TciGOK2IgbkeRPWXLsVS0jOo3lDSqAlvrUFS54g1fLUq5OjhMi4++EsX9aOg86nPbj7
Y6DhChwPeXouW5T+/ZJVXp52vNhD6XKgu7ynzLM3pEqnj+3VIykNIWDmle+v3Zmm93vgBwONm8vP
YHMEyfcW6Og89UGSzA6yeB3ZNuWXdJyFaew6fAG8E/kE7Klo5pBpTvkdt5WoTL0z0p4VBNIo/dYp
t+Gax6Wf0GL03JrGxLVbutWn7FDpPuP9a7n/6Bqk0r4MnwTOKrvIjmhn7G1u9BRrh8agTpo+XOwO
+6RFqB0VtH92KgcH6czd2M4YOySAsTgy3jR4I2CUr4qP7oJcSSSdrAOsP7a8J1mNmOLJD7WtSHaI
loE7Arc25NelsEU/h4Fw8fPL7CwLmoWuMHhsTlhmd7D7LKmXKBzemstBGBd1mLxSw1DQbL8dSIpo
p27WJtD86BwKLcq4Dyq0hy8hHZGGX2Xi+Trf4YH7J86DpzWvwLpwsZo42j55KJNV2Hyyy+xmtmEv
gJqhdm93QLi0QAxssmhlAjGiGfQYmEBk5qNJswfRC03Ka4cXdb4bHUZs5FR56l+C3FLONyIoEOZ2
A77yI2Q/OKV9hv1B1JSAWCqhvvS/AJx8BQOSFY5n0uudRqOIEyG9Rm0jXBNQypGI08a4ailBM4qd
2ySZt2mDDuTfaezYdEAoXqf1K67erXXPEIrbXRD4U9ybVBzalREzX+Gz9VgEWW1MYfL1Qc7i6vH5
SlLdHUvZh+53XaLxUNKo09929jhOFK9KKADUB3tphbLmRJX41aXtqosj2cqpt7LKRMiPHsS1pfI1
YWqPuSu8fypPkeYFF7qt3RYfUtZfDal4F2f/nSTkNGbbRubPL+D62lNiitXQf8rk5KDckKCN6a5c
c/GZFJLsNcyPSmMt02n9TCUDNzzISJND9hp8bfD33YUiCqoU8y5alwtdUmBOdjL1F4SK0D4KQIde
j3ZhUbsJxyHMwearJWp6HJLUx6Ypsl6gv7H9h/irQ/K2EZ4m6phEBvojEWKHIUsRAqbZuQfreH6h
TC8+9lmViNtkAHGUIZqDwdhk7hkph8R68znHLRXlh/yNqudGcHftgGTc63c3KBgJDxMX+Qn6zIqG
l98eUSJmyYsbX0WT4jDlhO3y8acBUBqsJFNr/IBCgK37sCgBsDvy0bzZ4WnMsCVqpWlp8xelO62o
XgN0NQflHQ7rZOF06+S0mFq1fzcuLrNrEpvxsxJ5zjwrGC0v4hsJoSYis3dwQo6j/pTN+ZgqyvTt
YzsjN5SgWVmzsTQ2fmSwQ8o8oCjERWBHifsEvFoySNd4aEXiQFao/ueWdhm1brAx8BznwRXUnrA8
jjq90TcvSjfuoRJGpNvYCxRB9RJR/TfgY0bbvMNZW0Q5rBwZynZohv1tQG6mqDG54jjJv3hmEcsP
/rYwyJXrZuNJKPa//mawqC34WxDKdY2zGVs6N+sqrpvJurL8/9XEi2JDTuBbPiQSb8kI9/mj7LGT
jTzV8AZoxesWwM7+AgmReWoOYk1omSbrPmaJGZn/5ozyEGv+WeeShQV320BJuJipxg7xcszFsdYp
F2Eqn00B7fWy6dRAYsFxETnm+LVpRKO4AV/DrStm4nXv0QCt3dAlD52xeUXx+h87NDsmVUm7dROl
BYqhbkno8/3O/klvt1BkEvUl50xt4ocYWXlMrTos7vnuf8/tl2hSYcrzgPhGwIq0I6PIIxwr1Mh3
MjHrSX6m/+/bhtnIeFV7UJjRYLQMZg4D8qZKcF/wgJ9uanBErZmPwn631Q0mSFWOdDl+4GHa0YcI
KpJky9Xh7EochLFs2XeEn0DNNrt1K8cgnXlFdI8wB0U0r/PvX5z/FqEOq4AVgjXNN2aMEm3ypwCG
IIjLDgeJdMB3l7z/+VUThZcUdfPo5BsH2505ia5jjpZbDm0MjGn07uW5RnP19i/a36gR2asT6So2
URyrODT9YKsYGXKREFsReW4PrJvhvIbuY+fbLG9bfeYygyVqeFPhHrwPgAIt6ewFKkCSHqT1caiG
AhHp9F5aOfA9feG4oCT31DQxmvklZw0BjWMXhiSculbQhZ2vZWcIuxMkITQ3+Ao27eTokSCGGbGu
nPcIzABYH13CY4e4YpSMiVFv45D6nhOi87Tdxsjld7/ETNNkvRAQH04qZns8u82uKzhqxHvHtTvp
7tvYcXPiF2d5P2FupGtyhI+lYpGll0oNNcweqDSHT8C7VHM4o3g3UNUjOrJoeyIvO4dCziECmsB8
hdMNKoSX+QPqMMKgsxSD7krqC5Nu5UlSevHX+pWqomfDLzKpB089H9ARLMujHCFn7TrYtnS/aSUf
Rv2eCnC+uqHZvv9OBMxwBvDV5FBH1ekR1RXHgcZWE5aJU+n6F32lqG1snhiESFh69JZ0EsNtVJgy
jGA9SMtOq0X10kMHGp+YXm2HYhJ930k0ITaYjeVQ1wnd/kNlaceS+DvkRRffWHeueBcxnNAWRF/O
n+wE8mguSMbyCidxYPKKV+lJ+bPBZiSiJiGSEcEuxU3zKZdlmvmZmlBvML/GLMAImMPA1ZRgr+Dz
sMCTTPpIKmUybObWv9Bn6YGkMyT2tLX9wIx5HTbfd31NHD/94VNvJzoBmvPn52aRy0LI/DIidldv
SW2/jxg7zDwyVPm4SCIWqk29NG89Cde0Zvv3e1DUO7dLhwZCGWEV1p2liQKL0cnQYXUlxk3WDDZz
YV+8MSLTLlItM5Yg324/fflTWhVS+U0KT+6RFYv94gni5DDKXf0v60vqVYKyhhdl0jx8nkqQZN6P
9EAX8s+A7TKsOzt7Qdn5YZRrktLlDcawEO2gVHVCvzvyIWKhjh2ZwpO/gtl5CPSzB30tZ9emLsOL
6oO/fHgU/g9z9Sq8WVV+FhH2JnzBcMtELlZoeiPRFabDcRhsoJgLDzjLldTGa3PmWweCnEvs5PK/
JSO6AwY9rQGAECuKZMM2sky0WWBVn6AnDvxfYmqT4hcLkRoFwVD5G6Lo0ej+BQjXil+d61xQx4SQ
DRSTVTleeZuoou/GA+8L6jxlQVULnO+3DSo7XDA05QU2KZ7A1beHLmYYlhV/HAq3gmg1IGpVQybj
9840L3zqils+x7MtXNo5Py1HmswXQon9kfWgXbr88IgUs1LhdqJNVVqAj1eOLvUP56VlajT55Plb
n59uwCqKv6RDpDlneNlfN7Ueb58qmmut50cJ/bEXLFtV27p5CUjaZfWrH8gLnkj/lbyR8yddCWM2
XHhA+1Neb+M+yF4jdzwiCGUP1vfCZOu94BP3loofGrBQcsGtykOtyjJtGkCYmhIEE/YrwvlCH2zo
gXl81sLTjFHAEpl6KjgFV0qkGjtOjRT0gdFW9x2gnha7v9LAWmg9FZPhdrrzrJRcvZCn4FmPJ/9l
lLZOIbw5/CrV1rf2Az1k0ZUdl/HqlZBS7kW3A2YhSFRGIOaC2QXTlZdZEYJuaPsP8LMVoH4zWdz5
V5Eaa/SEC/hLa0CzXgxznBaAzII+jUAv+S90519GB7y+aJ3B9cYJsxmrYH3T0PWhAlBvNKV6QFGb
+7JPSMwNfDzg6ezhwRrHNGJz4tNmKz1MZzHI9rmk1zOgJpEiZT0Tif147wtRNN3H66eXL/Dw0Z/t
vP9dnE0A8ruvqTNTsUIkN1+m+z+rIZm8o/lDHwOFC34JiZXb+jHRvZ80zoeQs5TzNyXv2C9PMpDd
QCFHJ7e+75Mttiuede4FkfQRtgFwV6j2O1tmF0QVmfgLMHaFMQmRkBBk3u4MppOGtmJpmYkRZ+le
wapTkryB9F7x3UpvjLGd8tnJSE8u4d1TEmQWP3RwTKmgp6hL6JcWkdSv7Tg8TI8Lced+YVE0SwKo
rORU3SkBgseFJxIna7gqTS4UIja2x5q3gAtaOoHZ0+GfS9tt6mFmF8nk29Nf1h6eNrbxuuh24X1K
RrSfxcoDjbCTUa23DlhYqW7chTuM/fcmSX1Xi0mp1fZaJa4m0Xi1JSBtkg2PhwNr8SFbevprzTV6
uNj8qzqAxMC5gKd3hZPCfGshWdSbvxqrgmZ0LtXjcWLDbgb+a8nSplY35PAgpYnC126jZlJ+Yage
osXXb42ZAxA2NHmQ/VG5esXjJXNApFK/XT0Ngl+Yx4Qn6fWmWuDeVrVlChnjq/F4JttAvjGkOEeM
u+SRxGcltTK9JMtF1salxWvtCg8y7kqyzoJlAQiQMZfXv2fnUMHtRcF6Wn8wY8wpqSNZZw6PqNpR
MsCDwdI+qSCDbn1d5wtezS6kkGqKjkNPgBUNr8eixjuaB+iBdxfiuSePgK1cnHI8uNIyVWXQWLH0
tPjngmztQZYe935HVoIheBTsjD8uzHc9aE3C4RGVCvt6b70KGYxUOTgm/T75NwyqVN7H9hxVUB5u
LX727YQlhsmTTJYsiUZmp9PwVNe5sLiIYZ2VF4GbgQOZ3/M5GQa9B7yrjumoQM+iy+JHosciTKdt
4H4N/pcq+VllgkglD16iL2LCWFaK3GUl1N+6scalCVWP6LMPaqbaFJOFIYEz0YcK4b+2zqzegQP2
Bl6vggtT6Gtq19UFSfLs94gUFcrayT+cxAC/rkobbOAHa7AC1EnEE1qL8whojM7suu4c169NdwRs
dzxEedGGomoKuYnVfftXOsGpL6YSIxFDCuxz3UflJ6Chru+GaadwTyPYoovm4a8bOQUn/L2lN9R7
6uMH2rkF+i8vxpQxT7dB1owMao5CNdSProis448lGjWuPxmvmZ3CGkIWUIH6qnKUngndeoQXQvj0
bM/64T7qOq4XO9thjyIo3NRK0LSajCad9kP0LswS0fNefihZnj1COGdUKUu8LTpgzuQouVHfgiBA
hz0j5dj5AqjQy3mWQu/Zgt8798U/uFd5+TvepVQlOnKohOy5yBLkef7TquSNAc6wUqL3VK+7x4eC
iEflUJdDHl4YCRvGJ/kfvLfBy+PS+rnL3tN9v6UyyGTt8L4DnN5ZepBD9yNK15vEUD362Zv5LC1g
FP1X1gfCLgiSCLfih4cFEhP6TWwRycPZGse6XdFNW20FTEo9krJALs9N33XfXfyWAWEe2rm4xAq1
xKJuGRxxuUa2tBOLzw9kg1EgAF1EefmrwRxlnTUf+qRiQKuFoyjyZzR7LQ9xC6H8Ul6sq910oc+3
xS1QaLmLs9bGko9tHkXc8qZX01c9quh+t/cjrLMo7QOlUH7TO7qmN7eAkOzGf5OFb993WS91kFmw
inwz3XoHmYRCRTtIz89AQuJ3hBdSkmnWFN08JdNxzuzLm+HejG6yjmn0M9UguaSGxWHssEYZ2FUQ
VrzyFAFm7ZFVyj9GCsgwj7NLuaXWrOYpCYCaUH1hwj89NXoi4ruMmZyiytdBsqemytSJHu4WAdGZ
lATXEnFPESo3Yg4iHepqpvsccBpnxdS3tYsvlBc/vkVDeR0CzB+rGQ3BtPVLpdC2tURBOZ6cHyBX
fHJWFcSxfow/1tg/cZn5T7OUhOa4S1pk2H4rzATiTcXAXNvqz7/QIV9f1gVxbPQJNcAm6TeIGgBS
uKc/ezgnH+Lde9MfIajQ+l9ALCkq9bBib/7JG/m4/3UgVOQYwv83Ul4Z6kaOwUL+LqdJBvMWBWEQ
q0sFcetMBIXqOGpvn9zYinwaJQaWGCiV0k+z222zOo3tcf+Jb9nJWKeGTD6VVq5uykHwt5Li1EUR
8KVkhz+6lDQk7Pc0/WoI427ORaYaewep2yTcC3Kzp3QS2nt4/4EOH9Xg0KfOoyloLNww5r3nyDE3
lf9q90pTaT/+kJCbYBGaIVXks1G/Znx1e8RiA/paBuHOiIElqsYcmaU+nF3dq90/s7sBuD/0b2GL
Q4KJVbQy0WOHaoqSWY008buqsXe6xHvFFWmjURlYPfHJVV+gXir3JPN8veyimHqIiM/MPyacSW/4
zIhjPvK8EbnAKVKdwnmki1fbf5vqbRDhGF1MOlEdrBvUSDZyy0U2rQnuGiccqeyoUNqBKG/C2Ncq
EJUobGo+8NEUQEQtf9VASqTUcpI3CMqUy2IzFOSG3Trp1WaVadudIkJblHsx+D3HaTYge3gIjOlQ
JSiAxV7mJE5voXjSnrGUcC9xt4a9ivRDEoEMY8kELghYZvm2eqbDDvS9N9h/vIjQX/V/pDBS2nr0
BVOT0IVCUXsfeBbyiZrwAU6nRoOuqkKVaPplkTRD0bgZfJa4pX4ZFDS6bO+zgTYbs3a5nLwSxXkr
33wPZEhnYWlIzpRxSNSQoIYJxm3RBgRgjkuXg8nxQBhJrj+fJhvAxk0bCoFxJwbBTcmL3+u6BCKj
SRrYBjViOwdbuApUv4kjqNSXToGVMDSxtpmmr+iH7HoKpGvmFqea9a8uSGOPtEswuASFHnHHkKog
y6smhaBGQoi+iAeHUQ3BP0OfL6LTFwWxBNRjXCoZKe9YG0mNnXHZYCuaQJJibqku28BWWIgvTH4D
PskQ2Vl1vjJMo9FxDkE+nQTKuI5gnqHb30jiJiRR8579mptmaQU4Yl9JQ0gOWePF0+LnSPiVw9rG
cIwEY6gqyysa7mXyQUtSU2SbnDbpuZe+fS3ui94Xxb9KHlmyeD5v6vHzK8eguaIajaYb158Y5ZMo
4Wq2k+fPcLEMuBDN7CRRRQ2ly+sI4KNpFUIx0cWWA7S4Z0mg+iWu8eJjgooDIGGHBMwFPzKt1MeT
B+yX8ZVwqP1JeiPlpsTKvMzFQixKZvUGYUJv4PBnYRHzCFfpBesVbEERORXPeWhQKr1sE1IzmuwY
D+443G/cXwsrGD5LX6uom+vC3Ub6lr4ij4XuYVW9Ph12HckvoIhcrz/l4pDPFx4l6feBxeoFiNSI
xAFbksVvRq+IfZd8j1IeWLW9AYzSD3TViEwBaUQ1DkzAQNjfZIHNlVB/+3PRR/JQGJa3D0rKRYGe
hAfE4c+zSBxrgDLkY1mV02eGhyVsL5rvGHo7lalx28Nz2lABL3Vr7qNNvbrWpK21Su9PrO/KqTFC
zvqRetglUwk/FGSwRlMuKDNDTOc8jnXQpV8WVQZBLWgbWiv1AScpVNm+PrKa8jztNiuLI6e6zgV8
VlkIk4w576lyIArG8Mu5qUYfQxd0CHYqZEuHW/da5ZwSgBB0TioilUHODplEuatiLPdAdp6oZyqk
L1xhbmcqHLhRhfx1MUYBkpxt4Xr+AeS3qizpbMyxZ/igJsWwNh373BxUduj9dGE1izCxTe0Wh4Dc
gM6SPJYDBhYRBvG+ICr43CLlgR/50HfMKNycZyta0yem4gAf+Pta+oq0aP3MuqCoHRNg5cJ2E//9
Yoqi76vVDxexJLnC9cVxrxpUAvd6FP5kEfbvS66VLJ45S67K9/Wum1gu/SA+7//PFPXvveIWYPGf
yTLCSARFViX1MsVw4bvtqklkjMFw0HPkKexFm67VQWyPQ7DDLM/m4NLghV07S01pXgYlnm2c40LV
tnGPv0D78Z93X8/WgU7mahyVKC5G9Mot41yvnOCpE/qRv6N9VibDL4YfttJwOEmm7ydtTT0oCeAL
3tFnEV4jyfvCrd0ywg3ZXyEUdbxXDRdyDw3gn12q5H41bSeQy9r9+78K0fSY9DOrPb9xzrKGAL5j
PeKwqXt0mvvmoje6kOp+WEXS7EZUwe19YgcsptXDQSyIN1dWzGtr+j3FZL4OWpjRUvP4PquIAqaE
929Wcbvg4GF2HU+MSOBP+H6WsUflOeiSs74Ab0PFN67T68NTNUaxqOA1TwDlFJ7Qc2u7qJNuGqn+
VAu5v5eaO87EVtyavyAVeu8qEsm0OQ0hhsgxO0eWzbzeYKPjlLvdhUibM94XvjMViwkidU5vhETP
ApsrM89ESmkvvGwf7dxnnPYP9kUkyy3K/eSOBIq6xKFzLaixbvZT83dTEMJIi6KUpCvBf3GOz9ki
mEpI2ZsVTKR8jzjemcVVEC+t4kARwuHkhRGWMvVVzcsR7QyZ//pVjZFecsf4Okq1f0SdxUu1ano4
x1xlvauvILRovIXiX4B0pL3PT1katZMR9jt4kMfvDgUFwmzUQbALdlsfGmCewClALZbgXqr59aO5
RauMz9bwC5IpmXRY+p1PjHYF657jYbP+YdLXjbTInBX7FJWWVgXld+AcNR8qwvjDPAJTn3YVV2/P
V+FUc+SUHozqkrDQd0yw2aSTb5hQLilT2zNIY4Bss5NokdTMeG4ItIPEW2A14RGwO8mjm5wLDOm8
MjvdWEqIaW4aL2/h4WbTyLGFRynGTatNhxhBK6icUhUwpIUBMhtkloGRO8Z/cngpWm8PGR/JFBrb
dZuprjR34xvtw77oguPlibON25wd8W7U4aTKJj6hrTQkHuNpi76l3F+PppI9+i+2UvQwxUIY0C3D
asnV+1YrvFpAC84ctb7Hw7+dRtKZl9yPp8FJHeJPwVis0YuujoMOCt11/q1dUa8sys6qp6+0rOMi
h51Lx4kYloi2IKzIhUjyJ5OQyjJxepXjnjs5oN3+knPvaAsOeMhjPFgHb55sieLfBwQoUp6MFwg9
0e9umdkfNRrMQIULQwfeg6VGxPR3BoGny1rfmdVW2iPEoxU/W4vKd6ZhNTUCGIcyrjlUYdj/z/m3
mA/g7L505yy/QrXok9vk+HYLwHfwmFN995CLXUNjXEmnpN7jJL/snrXSUsO7Q9hhhHj0ZSRXdOBn
FIulPnppb2XbOGX9o/5ak0J7Y2rmI5eEAFNT/91Msl1DDl1n0Ef1DAlGWDB+N8wH5+aAlBNh0DZa
E8Y9Ke3sozA7YitceDoq3QC6wotg8CFc2Q4U/VZktso0pKtjsn2GLIA41VWM7BpvRUvIvSzvJNT1
1z+KlDpUvhutRB7fT3aSEvebOiotb5MZTDYQMmcqYaP5uJwMPzg5cscqVw3ThhKgPQnLQ93BiMZW
RuCH0xOFWaHq0cuqsNXp5kr/kZNhYYDNpEhCThlBt4TjEw6pc5Tnu3cfxRVEASjMTX8bP18BiR1K
5jledms5dAlE970QpuFrqHcjKBMekbOAISdIx6DMWV/SBaqtn3PKM8cYNyWcxaegr/yhQt5z+a5i
MxXmS0oP+v0bvtfBf9JQgZCIzNuc03Fa+OHjZY0XQGsUh27pBpJE+PqsZTuIWtltL44LrzoIsyXb
YG/Bwd3J3WrkaaAli28fHtG3MoXCRL6SOX6R3jNYOcjDgvQ9TCtT54uo/AV58X8jQUzjP0nXLRYM
+phYjVnBgDqP1Z5T1KgIgto6kVkZJA+XDg9VVviuXD5bi+/OCdC9ouew9YSx1hBXDxybh3DgMT0W
iStXPfebchiajuymvmJl/h/Ani8KVSNFTFMMGObNCmsbQpb6rQQxaOZOj6aRdtiOQOlOEOLN/II5
jspU7wU0ENa7RuM3yCbLd1ENQK1yBlgFlc0kD/Nea503LXSYzVRVG0oPTbdV02RBPvjpr8+tq6Pa
pIR3xroyXBkr+OeZ+rCefc21Yd4APALmO6uipJt4XRxSjLzDDX7YReVcn2TnZMjB/UBrSI7rUXrE
/a/DtwUXxfTOPBbnYy4NGoNLWLa6a/uwYSSlmklZYr25i2r2DbkuGWfiayc8gp0+F0QFXNFQ/OMm
M2dmzaQghOjaL+bth04pfw5ATgdobRmEWbzXE/XtPKb+e3TajNzSC40Eko87RRqgmfllf0+URX8E
XEoM4arq35lE+DHMd7E3ioKpvT1Rs9isnKb6JWJExDYNnMetggo4zshASNizTz3uSpNplvrQeWRI
dPwZLeydE80dqqoQuAtAcD8giqtoVOgkKxoR6xUurTVciNdF5go08PnzgYx5jwpo2cCOsH5/xng6
Vvl22uBg6A1U6vZoLzb7vI96XNXOMBbqTqquXleH3t7z1+JoQSXWbr6qqQeezPpoc7hoj14fQzUt
UxnZ3UKA7NKaRYq/aVISBF7TLTAH5SIKxEsgh0mmMLCC31vdNlAfzX7DqgEju+cU5gViY9z9dgGj
A4NZnvRsmnfP5ST6i4w5FcIey9mlBhLGT5MdXpuWNufGOOSI3OQkzgh9e0Qng6AbCi4RN/dweoa7
rtrr2FSi3A3+Uo7QxqXDy0Ym28xNb95dG6HwdV7s2TtcPCymFL+cF8Gv73aC2FCb2IpRdg6szAYu
rIaovnJRWUrXEjapW08E045G8m9nnbZjN8zCngSmGWRZXlvf2olM5i/LEGJkIWG3dd5NSox1tsJi
oEmJ5rDqMTP8k4UZHFzFWGXO6V6nqT+Obl6eYqhDX/U6TITegB6mQjffjXFN9H3UIsKlHoZtjz18
o53OFpVrVdfqdfweLBORp+R3+Vwt0xkayI02K4YTv/9BwUX1GQaQjpbewhaWyeanh5FEZ6qEQR8S
LVE/Vde/NgzK7P/I0mh6erj+yJ1gkE0sDQ/wlAIlHmgoPY/AWw5JDq6K95KN9QeJeceoJooAmVlr
9BqiyhgV3BGrQM9EMAQW/yKimpScOSbykpt4tUJK9b2Y2cr7mJCNFHnjod62mjEJN4vGFIhTZuYa
8lYCqpyfu9UHvOmiOYMTxrTEm0ixpqazvFDZfL7OPHZ8JDRDP89kesCNmJHvS6TP5IwWFTwGXN4d
gI3th0uj6LF6NEZYNN/UozHpA5QYr69LPlZaIS4EqZFnyHr3ilRdtzE+XodgPUnW54fw5Ft3SxJG
EjiqDmWv4qto3Vk8nsfM8ILUa5NLxCb81xy+6LM4Ft+e98W3mGe5lzDvpz0j5lIIhPO8jBTPphTE
zVN5ga20ytkkUefHhh93qFlw1zutIU4RBUEYkQzSta/ICoa7h3QKdtOMNWwDJVcvWVmAtOAZwLye
yiBQ/hAnzy6a7/5otrZeaZw2VBWGFvQODWGN8kCw1v86eWjK9/U4J6Zfv3+JW7E3HBcpajBQRj1t
GABkz7xR12cxUkoMh24Y5lihae67ZAISsD9en/uaSwRjO3lpLigIX86Ahwq41LmuALXEO9RxRmhL
EtdYyrWOL1Idt2nKRGWIcwQew+6F1eov9suG828QrQwjMEItdeCjTEu/7XKmlULDJlvboqLYf6zr
NeLk0zzjZi1Sr/CRAhKD4xxW3GtGzTbYRHegpJ1Vsw9IVo2qkQyGxEBPiodXWzZCgZ5EXZsEZj3n
CdzoYu25/VXINtmSBNMGwUbkPynrnnJQSS4gLuaI6IPLGF7WdtLK9VF9/JP5n++hjH0qDLm/TqCv
keTDYz/iZ4AnKIov8r6KYadtzw4Yr/7A55epKsOdDb/P2a+JgYXHog7kupcZOuag7qf3lbyOAk6H
58xrIPAsesXUIMHm6mcm+La5Nprf4KEtKe4OXRPvyX26JjsIEal9oR0vTTI5/bdd6E6gd2pnZEK4
jaJEDdX3HHCGkgQwCGuLzYu8TFwU/zKT+wPDHGqer23PxcB58nqVLVEDj5iw2lRzSZrVl2Gzmbkv
d1HoJ5s46v8kheOxJ8j65bZsC/Ug3TBr/Fc34rymsf7HulIruNJBYSIvRpNlqmDIqbUWH9FqQm6F
GNoJ4nztn2NfQEUFg6wDjb9l/8WpUjONuqJGa1Y8+3I3OL50mrRp/oFM5UUgLweQ80Q9fVJjEwM/
NrwCYPTJZ2V/6xlRoBlYuQ++38ABYWc1GSSDFu3T0DMxX2gkH7iJxkbQ9C3cddo5+wg7q/XKC/wY
G9pc/RFGpGG8rb0mxMkWLGN+2by4kZsjoBhYtEAfMBureqUm6/vQsqAApHKFIA9cTgqeKvUgwAeN
NwQ/SFkmnbwQYrN+fUHpFB7pVrxPDUYuQVWmgBNIYQQ5iYJSbkWPw2YhYxJhGLqBKoCQhLGTAiIh
bwl1C0nt/UOOT5YuGi3iSf520FZUUUUearPt9S59ix1eXRtvd7yWuRJtCtUEY48S6oB6jG23QkVK
lg19BulQrn88SBPg8hrmqKx8OGW0FJHbuOy1vmkhFufs4IULZ9Hv1PAZ7iWshNsWQ432uuVOOEss
KTMKFm2CTWpgu94owWoivPZCBoW3usjLpqe6xZDhclCvU24YAOG4S+Lh5rm7cTXAq7mDhYpN7YYz
6lIx9D/UCJdmMEZ4nCqT5azK0QZ0O79GzFlG5l843AJUR/5KCpjPJ7oaAnSxdnaIK9qlVmd6RzNI
t9RP3kZPvle5pY9TGfoYTLo4SLUO9xbQKrRVhNBTyaP8jAS1T9oWdGV/pjTJAx5brxGJ84wkyzVk
3mJL36p1EH0h+AWONfLhRNpTlk/9c4lz8SYr5JZEQJZoGyqWtJp1oZzBmwmMsg+O5XisURye7u0p
VZb3jZ8Ak3CbWRVI/zLRjDBO4em6ltcaGwMXmIky+igM5QUAncfoOTF3V+rm5KMUlw3KIt308Ys0
2JOQ63wINtWDt6xYjtE9uu/TvTvQ61U/TpkPIoWmYdViyGeS9YY9NZ0ABceblE2W/l2knZ3Oy1Tw
ygaJimnPBg7RMay5/wcV5gjyNqmMsURCE7qF3Jr0Gh5wVE1++XwUXmYTVV5iFc2/PzzLAPdnklfw
20omwG1TDmbDrYdBM9zY0NYc0SyttOk3G/wf1pHAQa5LwqjjXWRIEZL81nbU4p9ayDsn26PPHz55
NgfCo6GkbYpIhpqOAAPitkcjflTmagmS/DiOPQ3KgaLbDVyAStkR0dezwL8ug0SjVCZIzK4Gy5Fb
E5kohNs1LfbZ3lQq6nAUz4EmQUeuCuZYdpzWeLcvNVMMnSjE2gYNTi2yuy9CkVBCagD5/PWGuMgg
9RXzDfjBydJTslas1u2AUgAlvwipMwmnQzrto6Yh/8T6j0gRVMtRcgftdxMK9YJQRaEj/48HM4Fw
nb40jT1ni3IA7k/UqbQFNOkwLX1h41cpedEYdhHC+RcmUSf9/NXTZgi+uzURgZ92RuNLvefZPMZS
hQ9w56mCjXub/oIs0c13Z8VuP9oOwTtSEcpiPtUxfzxtFqQg4IKPnXhszmI/VMRDYzcIwXLOjXdl
pSUP6kEjtUg83V1+YysIp8yn/VigzKCZ+3WraLP8X6zuBfNlAJeA0Er9Rs7PjUD14gxq851SlVRm
QZo17cCKcWgrA7v/t++0JRHLyyx0W5L4YO5wGM1VnYUkn7etkOjpZo5p0JiBRAGawgy7U5qCzQHO
xmd2Ka3HjXC/hcXc9xw/keS7upryB05Hq2IfDf+Hcxfu18x2IU1jPG32NY0kmivOWL6S41qJlwp3
1N/XoRocPcFRBrONcXH8k0L8u7dLUzXeoDNo9xr4j+Ri1H2TQ0kga3pnvzaBw4vSSLC/g1zN+l6N
ulmCcrEU0ItFn0b2liPzDgK8o+I93h1chq4rccnNxvzjqRBjPldV9dIYIFv48mfskAi077d4wIZA
J6YOV5d1jRjB8pnTRoYNvQS5PWCsl3g4lDGOJDTD/jQmlQcc9Ni3eO23MHjoC3molCPDz3vzTCNv
OKCB33qRN07zmoh6Fw5E4YZT8mxkj+UEkAyIykfSjy8tqsQpc8boPGckUM3F5g35EIRK3RmICGVa
PgZFxCA8vv5Ke6w0cVuweWCMjfJSUXeLxIHC7SPKXe1HIBtIMBpNX0pa6hBmDBH7w+Ov8MKu3U6f
+sfoPByBLmWUJ8rORluOligtqENroUpUqCpHMxGDW+VxHVK57boKdwzIsvNymfaD416BopfMrKHQ
bObEiWYUYVxjwKeoF4L3Npu76HSaWF0ZhVmTrQVD1+Zty7GI5/cC+fKbvk+JHjZTow37BeoHUO+i
wtYGy7/b725pN7/BGJcKetgIxhA48Krhn7VJ5WFWJIa9tjyzBypMksp/2WOuEwf+Yhwqoro0gu0i
vGVP05EIsODcZYc4eZZXEwhOT0VExj6yMxFtJvWZS0xbi2V+v/SkgCk+NanDoYMqDWmU4CA8Tcqa
KKlTe54hG/Gs+stMuebXxe8kwL/C772eXgpoOo/PlKh2vQijlwjZjShzJYBooTyGjDbao8JYmj2o
x2bCAHdAkOBLM84i8F9dxqRwtUXH+2JG/pgxehfEBTV2GeFAdqi3xglpn8jpiAomAX4V6+tJj7aN
/GMZJS/xsV0k/6l7t2HD5GjJO+hjrxkhq7E6n2rQ2QTKYiSIzt7oiDQKpBNgza547CmyHmqlyoJX
kaBfzlHqac9F+QAH6pTkW2JYxZdKAmg1f7JVwPrsSzqGBMTOMZjaNcM0XtXAPu2xFn2WG57kt+5E
1IS7NG6L+qarxbys7bbmpdojMTeSBosfuVrLHzhNDzE5sJZTkDzW/exMdUa+HsEY3uz9llXmH296
fUxiAWrK50R7pLk5BmXBSI+zwuWTVp04uyB1XJ8l5phyEh6zQLLjgf3iiotzhlnuWP+ex9M2wzVS
YqubpYAoLAyfFx3aboszsTGuAd5sUIKAnsNgRSeKFjv2hU0VpOZX4o5DrLP9qDS1Na1Y/ndwMTpb
z/2ZIxJUbyKaPFATsxovYU2hVGjtzLVdwI8piR0JXvVZnYuM37jO6OWv5X8Ml7CWhDVYqBq8RMmU
p+4OI9pfMYz+alp3kUtXQHM9chhZJ7/nyqAKQaVNeuF7Yi8Ns5qxYiEXjzQHc5h7ay8lqoj5zIhK
R9VLBIVbsWFlE6PBzCz/ZUdumt6ir0CwHmlSjx3VaHY5DV5R7vhMEuOsYf5cR8+SHyywJHNOMrXZ
JnRO92DYXMNwMZRm3VniFfT2NxkTNf/UemjMF0uQTp23rpQp0MGJ+erD6E9PpZ+4KUitpS66aglI
wi5B8/tp2pxWdHD630hNlRS7a+EHtXtHL7KYnK4ztzILfxJBXpAWvI+DAjVQ7sXXdVaz0vL+mN/3
J73doBer2wyfaIdYsEZ+cfFY3Dh2/1AwMkZ6pVsgQJ9n+f83CIBBs31uHaQuE2LEru8REz3Cuslw
fc46uVlEh0MGkRb2RYhBEut6YOFG9gipQCk5anV36hYm4m6RuFgnvCZKAVCMXf9O09erRT3zw5+C
6mFJJ5kczGO3ZLce7d+nNQvUiIkfXl+aqwksvQNjFNmYFwOadIhLpsPe4Q5LdVDP/pdOAKvHyN6j
S1e78Mp767IcDerX7DYdEfbAoOC1wZzOQBxgtmjp1MqkNBn7+FggLK0h1k2fRDC6MPQGT7a6PGBe
HGTZxgQh8x8AIIGCMNE2D3HKcZP/BQP3IGq0G8vjysHNE7YL9Fss77WzoVz1LtfjpIingsoFKjCT
+Ul9Ijmi4rUrNq0VWUIp94aTjjF0UwVWFIAKcu6T9S7OTJW1HWm+9WieQ6vEplsiNdLBf2Q0dv0n
WTjTtiLUToVLuFIJnLerg8ByNgX8cQdxvXuwe2q8ELfPNrKvWDMCDTA02cUABscmBEGylWV3J9Or
aGW+kl1YpGhBBybUWxdmFBhMY7h7oGZJT3cfskDR0VoGr4mualXfUHS3XeMBf9M7JsKzhr3DL++5
1A0A+xfvbT7s1+l6RLuHSYf5ZcyeKOZerxoGHa/td0Sq2Sg7JwedaYMfMgS9ektABgX7OBGtq3cp
u5bL8e7sgIgQyWZKg1OSYIFkwU07GR92oy6c9kAFIG7d9eddjRkGKwtgsd5oZzttK7vxu+RgyZKI
pPNWuJvBVtYClKK5sclc1wsrmFdFivCNeab/8hbFv32vOc6mEZIVR5f6OOyR2dpUco0reSKpRIQf
OH7+xfp64Xsi1/iAsRwBCfIGQz5RnQUn2iAXKXeNAWIGZPE2xLiwDLid1aI90FVkJnxgSAcyFNAB
ywrrKaekQNfcOLMad+I4IVkrnlM+jj+2w4pqSZHCyzB75uKitW9SjQavier1JB3aAZLxni+IYqC8
VSkeAF6gWTP0Iud1lWIRdXBFfz9s57YqhOUUaX5f/jvnpap6dGDPU57+vsYL0PMSD8ftl9l6FCdg
rggDEUtuRbN8Kr+E6OLpCt8bzTZk73hO3Q6yDCamjpYPDK1asUNbTe2h6adGZAYD64J4GFXZIAma
gX2fHZ0axdnVzPtyXCs7TZ16lcKtrrwxovfx74WvMnQOVoGaZ25BLWjYp6J/0LWlH+Z3qixhZaep
vPYVld6oUMCaQ4QsWClHJrqoUwKWuMZNpB3OrODqRA6kG7PQbSKBdw4fe6S9UxnuO2ZxZc2IHhWb
a2KgUrEA7gSmqgQtqDzxZLd1837iAY3pdrtpR8goJwqx33A8HZUdR0f8HmNsEqHexlX2KRrf2L03
mqaqt8VAme8v40YEq9WKueaPW2K3MeK6BFmexAhGgWtlks4DBYoLjIkXcKv3igPNIZtmMM9NUYSz
3yFGUt6v4UV53QUJshucVj0MHmjyss0GY3ao10/6B+a8T8bcnWz08ZtrJs93BVkTL8JTm7vWvR5N
scNAmh8wqEhZh+E04zak1krec6XCgF+NcRcvfkm+MNehXMWeSHYpvdn63NKdEfdDItLzxYmz9JHa
g/+/kKG4q3tBknrKv+sIGpkfRrkWLgECHxsVcOQAzR7K+AJAIL6ZN3dwpM8Ai7xYdmRHTe2pkJ1i
0SHdhX4JAjqloPespUpK0tvhBpyS5V4srvG6jf960rR2OWFSOF0GXmByHsE3kj81OH5Y46yuFlq2
KPoswhXZF03uFikF3lkj/at9Bwh2lBnn3lGMjkyEPDgmEulY6NdlziRalpT4lGQGtYR8VP/CxnT/
rl59p34GXT6ahumMhJnil3rKbsn0eQVe2YHQ0q74ZgKeobCAKxIZgnG9X7qaDpyMBxfwPF75SrKR
R6QI2e+PrOcccrhujn/+IMBBDvH2oRuwJzKW7xTnH07/PHJj/Cj227RrgmsSm53EsD2w8QKK3/Fg
haVGyRD7jT6Ht+6Azh1VjT1k3oYBki+10Fz7NUeGE5ZTw5TfdoTPizcwNAR+ASHtL19dNH31SNcE
8rkyj3+qIcR9N/UpqFL91OJfR1sRhuEthw6oiyIaePUIp21vRr11qc7kgHSQztKp4ctHwr0PfFUe
sd9x8bCOaEGv3BVmvKDA8njXHek6+gRQkSAlxkcC2OBeXyIn85o7CcTJ0Q18lH9Jvr5f3TI2FWZV
rPhWc19c/xR2VaaPlPSIb5veCaEboCFL2sABst94agnE/xGD+fT3F0Q6znwxjGqoy/adeyX8+WT1
0jn7wW63AHSf1wdfD5M6TBjhjjhsNXV6ASwZaHZHe6giDw/Lcj2NlgN9MQQpOH/cp8fXRIxpfxPN
TBQ5Y9HgceXIdQYH4Af3QQlg0xU21XYyk3uJzLld4zZyN6+e3pgLkkJDQpn6ZAUv2vhcsNPc8aO8
fMa2UQ1CDacUPxyYpP5kO4sB/pRXu+PKM4xd5pQ71IS33FUYJP6a9mCX0ovmuywW44Yl1iktr7GV
ud2azWLCb2eiCX0C5s08lejKM0qPgAvp3WLjBx1HZwBEpn3VU/PPvO2uabL05mhyHzod3iYBtxNh
Vf7LdbiF2DBnfch5McrMABiiY7kCKDZvfQT/B63XukD3DJLkZffuKVvZ0H+NH0sgzAlv9wtf+DJ8
JBPCyiZdi1B5mPqRiAR/hEv5wJS6AU+6NpDjgHMV76RJF2g7QYLTE8CwDzHyqpIbdLV2AyfnIny1
1z7EZV5I9y5UGwNC3xobLWfUqGsouvVbgPw+gCRwLrzeoxFLvT++J6ZCVvDbpeB073C+ROjn/PlX
5mtIQTzCQqmlsQDTRElvQlKCJPUUHDX/nxWkz+h2Ya4qulMVqbyfwqZbOJ6pP/DBE3SfV+6aSwwJ
0sW+DixAyfkyPbtY/sGeXBQwMWTxtPkJYxgYaFrQNrzJYUGlXXlL2gMwxhWGNFAOEZAwUoChzG+Y
andlHMeyd5iNlzXId0XHW2t8+Xfxz/D1eYY+KjP7XL8mNOANmm9VMHhHv3B9z8SB7qTpl8OPgchO
gffrCcjj5VEKa9ZtFqwND8UD1Do2aiWMS31ShbGKBC81+MjZQ8GyXFkBicm5yvyU0Z2ugullI0HM
K1Asdx+IhguEKMGMWX/OQGNiCw2GYdxAdhcUJEaQ/Zf7m1o0o2AisTmeI8iVJwZH6gvJaAW0/xNw
FiM0HjYmwpIF8lVgaqll2dyI4J1iURGrT/UKXmvZffvwak82jmcRLRcn1TC+19zc0fAIAQB1sgJq
e+/AjHRmSvQ9WTZVAYgQTqmD1G9Azcqkq8vKNCADmOGibqNDg1v+C93H1Kej0pGqTXrw7bGYZ75e
vs5UzwwCqvpx3uqczv1SOPAim6lCFRX1Y3RM1h1Z7ump3knnRdUAP/ojrFKR/p11upOfgZhfo1hE
+NjiC4IZVZpk7frNqob9CYnY0+OKxy+9x7qZ+5lKVLno1kzCRbC3i3Rw1qDdBdmR3oFh9j/h7vHT
tYf+uLbnV6CvZXMPgbcnx2HUrLj0cINV87wiAPxGs5zlRLBgcUTUQftA8z1ZpkXSOKbb9hjajNF/
egRsry+DTqC2dvN6KXnZa9aL/1rYOk+yW8a0SGsAS8l3l88a/QeP0j5aI7xo/yLQCNXB33ZoXPEb
ys92VezBY+JGI9QL3s+mfb1IjIMChKw95R4hcKG+eu8yUgz3ZEdIEof0s1sKL72p9bZgO7ytD4AJ
F7tsGK30hn9YGNW4jznsARwullVu2RdFi/2LT504ZcxWZ888QLTAzxwmADsznERNDjtFnyhTt6Mo
83rtEk3BGih5X4D4LWxgKnyVMyceMMj8ZVL8+iE4bHOg144X93DvaG+7lzZ3m5mLG3sQozOOmrXB
a2Aoahx0AdvCeQZyuDJHuoJsdaFRoVdusZKnjsvxu/fjV5W4dwVd5BNYet3/RHBDwQ4gedBEpaQ8
f0EfTIMqmHWHqBrXrLsjmbqOZ03hZhEtrReb/ps+YoBzme6Zi5fnmIyCsNGJVcomw0048WcJi2sy
YhjzlzBJrRol9lQKDNE+1zQFdBbPx26slIlcfJwoFg2K+PMKsUcCBG/6caunsixVKoqWvz1kkbOM
wp0fT7fY5Fj5AJPRQig7jLmnVKRWt7h+cC3PPO3WiLUgn3Objyr2wiF+5Bn0/D8IcXxB/ePHloqK
LxUKKXml7N2DITah1R2d+hQk+Ay0r6AU/AhdSm/gdqX8lCC1cOUznPMTZLVrv721IeRqy+NkSV7Z
8P2DmoO0hGWxEyAGiyuDUKDBYYLKihULX848H6Ggspu7amlerfDRtZpA0YSEWxvg+qSPfGjDSqwh
074QGxIaCRRfE9z/kliBpRDxyKRlr/08iY0++7slt+bsd62HvEjN1cAtW4Qj70+c4DfXPxVpR0L/
biV1MHlGLQ4w7N+CEHYl3bpulr8Et55PteFhvBLDkefvTHoF0e24ch7h5MW3shp/bjrSbOUYAgEW
C5I4lmG7QIoeQ0bwaMRZ+apDyO9VYuMCiKdTUxoT070OU1NaAvAf9qOTv4mFXNbNnFTcWMZ8xcD/
RkRHyElVwVwzOJ3gma2oEQ2UqrBqgRKGuuwZyDwYllLriyI67CisbVV35UCbILUme2zGqE2Kejie
jJU9wSLoEHxOq7ox9eotp5iE0yAM0i5nh++DKjYUjc9+JBTC84Fefksn9X9KfmlhgYUzIgF3yJtE
wymqqXIUUWYKCnvj5nt9Uw3Rs9CCqsAMwzYJrr5HNFw6YUCXda4x5CyocwMXRpjiHHEQl+ECdKR6
KCDldy4LFc6PNkeXg68fZ6ZzEOQBDHtG5NlzKw4CBmvGZRUAGRtF8timFLZWGn81QSk51KCtz5Ib
kC4/JqhM8IxawNteoKCpvP6heOAWQEB9oTG+TdEHM+7dTD117l1Al0tepFYQ+efKiuMWws94J7Bg
7mt4/g8E3Y4O3S63BrlIS5sKHSadq6fKUWGyPFVHnhMdaD7bCoGzx/wbnUfErXr6NJxsPQgXzqiy
z7gmgPrXntm6REh73bbsfo8CE9xzobDCC2BTY1PugqM4tTqTEeVzW+HiU1scj3Ja2bo4qsbTxAie
ui8S2+8MkIR/3FCtQYIffBbKxNhBHbyIbXkLIGpBZORWA2q9qiz3QZhTjSAy0ECf0vGdQFSMsj29
W+HlMmZW5UycwGXxYJwJ1NB+yy+TBoLErXWDbpjzScvhCaAnyecckWVq3TZwjKHN7rB3w3oa05LT
sSKub2cQ1hVzpwYWagGKt1+N1JFFJxAhnNaKXrYj372wD78ZZ1CdU5pd5LfI5FcQphVNpQpxMkQw
WjtpTpNOuVqEXELKaTY7VcyDYSnmt886CiPsf+0nwZCVWGmF5bHoEhcXjScR72kU4+JDy5jdrmMI
wAUSD4s+wLfYL59NR1krWXzGVgZ/xclmEJpeQF8g1MVRK0WBfY55EGAuztY5cezWHLLnEEEbupiC
1+LhYxCpLqfCjF2NeRBXnptRm5yJJ63H3X+gN/lUlbzKXU4HhCf5mBNONm5jyiXt9TzZd1mDt7s2
OWdZNF2XzNI+pCkGF7bj+mHSUmMQD3T1KvDqvYFylxvz3ZB9WbkURNAZp+XJ13ppLe9goQvg1YeG
xAGFWM/zgYuq/W13d5IeZ6XU2fW+vvaZKR9DifkrYdahPi2eYcXCOx23xjizstZzaR0QGxe7tAoe
4klyOZI0GWzoleHXtwYNxZC8IdnRzlummJYzW4CtXpr8+gVRckLUTOyl/rWGS0EsRIg98SqHtFam
rTqePfB0A3g0PQ8SZGCv7K5gIlpYxccytlc8Byi45N9DbAwQpahurBXX6s3Kp9ul0Pqc5Rng+Hn4
pZIbc/ZMG6Q0QPjHiChqYa0sDcM2FL1MZSwRSzZCSr2Vo507AZXn23eb7Fl9liXOHJI1+UxhhrXN
Ai36mgwmckTnuuSqPviQutqKR0ny9BI1hNXVlFjnfObrExOqYU3nvy5ag1jtFW5GTTF1DISmg+kV
nvO8iLSA8DgRh9h+8pf7bqVkA1JXitMf1cg6kSeS0MviwNweDyDv7zl2ajumoOJZ7YH3cr2P8DnU
12HUMtWB+d/tKjfQiFDW7eNazw6FkHn8SfUOco/czc3er435i0KFpT8zYKXDvA82e73IWIUGcGV9
33R4/uzEYTG7eQqmI0CJTPBwjhKyB9D0f1WNz+ZCsxzYTuhiyHdKfCG31VDYHGDHm/qD5moCWj9R
FEqON/DXizH/j2IsOs29CaIrKnnW6Q56aZqoBSVSd6imYpWQdc9n3jwUkI6dY+2Ao8pDvytRrq5H
HgCYwUN9jdziI9uzCwUlZlecxzGgcpiSCQmoGfMPws/XWQA9Kjigjp4JTnMquPNSsXygfX/gEM3v
iloAjJFcdU30oUAvNU4qdXi3WAEKuHJYnGzSJy/PIBY72bFiQPlnkvCYnRDJB/b/y7zUa3Lj1dNI
R1zbFWqJj++3weuNymt9SabS5/v9LAwz65RWqfkdoF4wvCVKFVO3nEBvwOb2xvxXfBDTnQ0Njfik
z7nCZe3tXVoVl+4K8y4fwX0XUhLK9+CaGihLk1ilp2hrwHdQNXs4vLfgapB/54rcg2LY/qJxq4e3
i7AM3Br9yOmJDUWnPcW5AVGrlbWUd3WcsyZkNOMJ9gERHL097hh62jnkpfQf27aBh/6ouwb5uMoK
vjFCPvRiRvmFniUGrAQQdUTcZI+rCjxYdicrDdbr1Vm/zZ9tWpu6EHMsOVrzTy9PuuS3blLKk9B0
AcLGHoPYTcs6NvedaobDfs8vf+HhDfgz4F3SmzbdXm2H16kKVn4+VpgNnXBEVhuMSQQC8165aEOO
52XYHvV7pa2oalcNudLW2PyACFXn/Z2AJyHkCPS3EGmvvl3nyLk/gQlfGSibqUdQZWH3BH0ad3wv
vjSyXWmBCmZTv9DieK1G1+5fmB4R26dFRdSkR4380jke05li0gPCGide5sqMFw1MGLqVlVIOwVU1
EmirwC4EDYAUg0ov4E+tyqJnBcJnO2/mcH51w8I/drN29bRnNmRFG2NO+xh6WqAWQ0IipCaJIXb2
COfYNwnp5Jgf6WQqaSwSN92CeILFqQADzYDbbjXrIdluoqCtfFnPfgzgORyKWEQy5j50/nGJHHeY
qqA69ah6a5AXgz/KRSJhBBwHjmpXxEfMOcBjplNvSwaPiWVKljkS2w/s/zkbnuXeEoAF8hvjbTgs
VBLHzeg9X2nytG/AQa+306/LbuOquGxAqNeBHRSho9xteGi9cAY2czYK8rIRilnNM9o0S/eFVx9k
5iHMbcvDvkqhKzklon68QtXXY1HYlZHegmgjtBuRqu51QJlpGbjeGT95FbIQGS/TfQ+MmnfkYX/A
pfC9F2lhHLMV/Yo7MtzWkTLEmePmvx60h2K1CfPbMcwjUgbHDkzAseF9HY8bZZ2h5kJjmvNEJgFK
BACLPiwmchkByUmjA/artaB2P0X/VVFUOZTI8YeKTT6plZrYh4HFdPvwQTQhh7AO/93OI+fxnzo6
AhdQ4NM/pDapJtqGm6zVFSOPwUVfMHM5dZy/fh0ccf+URZz2FyL2I4WIYqWqh7BzHSb3dRCNefVG
d6yryqE1XOiHCrcxYutiz6fBEKEQ2g/eJQ7QiFLho0g1h9QdAUnpo4FnGle/NNzyXPN5rQ6Encw2
Xinrmx9CGFwlZjLYHpcOHdxuJtVM2+VS5epeAGOHhgBGxho1AjUkMgUDioCd2t0YluvQ5Bll7uuD
TXJl+CIa3ipSNQrZycMjzOrmKCD6g1bNtJtYYRikJXFMXDrukms4D2LOumv8a9ljgvsirKHWuzYa
QaTi1SbcwjdxGUn9QZ6pItjeXN+xyul8zMlLMaulxozBE37nk1euc9a87ju0c66tgMHlRBSCn+Uz
qD2AsiZh4+EtoC2x8zWgDViCeIseCmyIZBbHBGb+1LVwIuWpSTZtRsx6XldCmUF53+zTTp1PnPMf
cj+IqbaJxecEx/+BRbx6xv7E+SarqdwbqOUkguaZFY8yF1/J+0dNuruIi5HKYFJj7S5VbIu+XjIQ
i5rcAhtBaf411ZCrwXF6Wvulq60fM5EewSDFgNItGy3Bq970vhoR1sCTm3nFaAGhmQUwy8rUjI3W
/eaWzxFbuYZph0avTD68avqRNNVb4ANZ8w0qiU2bmXbko5zDAYuxR7Sh46Za7Ow/mG6skofe4eFr
cCgg5xNG8gzu3RARK2mb8p1jXecVeKaV0iaBORL2H8nP33KvhHcXcShJjPUB7efG2LBrcNqJMeWt
YetR3uV0fJSJy70mRcrLKI3EVC/2WYfSmblfu0f3xAQkFVH8kqm446SlUfYfv1Pt6hS0X1u2Hsjd
lwTuATw0YqW9ZadXWOKYoWFO0uU9A3rhJcvmVCfG/68lhHd00R/I9GBjQT9lgQ3Nv4+dpLMNbJ0C
uyvFEwHbYHKppB2cAjOgph5Ydw+J40j9oEoUX9R3aZ6cmQXP0lzxSE/hdkk31CVlp/2Vu2+nXl/u
C1F7nhbF+ZBP7JENik2s9h6uVZl47uFZKttlSc4wze4deeGDcCLVPGv1XSI86seEKudlXKChxtFv
ajLL8NAvC8QMCq/sUkoKOBm+DR6wgg0nrGEhsiuyk0Qvn2WjHx3Xqaaan+m5XZFd3tOS7vHr4RaO
fcKl2b4WRqimNF872YAflWqK9hdMGngi5AO22qH46EeCRkbZnSjVPtKv1zZPdA6YdbbxVtnj6ge1
BhFJqtpg6oDD2Fiw8aFZFDcDQeQS8+M9JQUPAHHvufEBXcTFXbChtmNF9tx/cpBbIsxcbvhGtv+W
U9JNhK7t9wa8itrjgSGoq8ZSGvbFObgicR4c4H/JmuokLVXzJAU+U0XSGc+1VVQT68gs2+I6E+S3
5p6k4bkmi7Cw5mdPk5EiwFmTWOnFx4RKbxJoNOvmTOtRDXWdUW+0Ok7YGTXO4UqIhjIf+f5DoguD
l8gN7xKVXMkC1655r7+o1EMOzubB90SrgjpRQ/+ZNjray5JkuKX66Y/CdSUMTGIujklC9JXUZXhQ
4CYXFKMvSuGpzuvWiAayAnMVByondlSTgegt6U+IUlPnRENKG+jrE+zMJ+BrBU/aoCis8NKUpKH8
7W6Cp0fTDFCC644LkAcx9Mtzn37NbUhvpdcLuZFdDQpUEL5SMn02rTUJI3tkBy8hycohM+KoZOg8
Y4rPlK2bG+lCythwnmAiDR8vczKfg7GhDtW7ZnlMv9jfgkiKd/s7+2KosLWWHFn9/C3HySLWzghe
3xPsFPw3mrUECQPdpVVWDnNE2kYeC4qb5ghlT6BjuWmn7qlkcPDTOWpbEVKiTg0EUfpAqnf+TOON
jKvUVRYaOsWzvuU8YgN8044TEYpOTH+FgOkPVetpJ/lxqWm1p40/1AH0BFrrPLeF1L/X5QruUkDh
XR4Bw4AkPb6qpitDPXU/yH3yB9kW+6l37W3lS070I6VUWHSMDhL7w+Cllh2gVddvUwLTFuQ106YE
BksT5XxATNk0+1sa3qnXGdG0AXn/CCdPcPNIby+qDjYx1ebB4rGEnJ95QB/mmvEwDgoQK4BHhUof
b79u/USz+m/Uoc+NX0jcuCZZxbtJ1rWfP/kKOKXB3/II7SN5IeErXX7WlYgAr+eJAlQWf7RAzO68
sqlA0LplSCWkfZg4j2N9FPn3DVPoOcmwZxxCD95p0rypf74SiKslQZ9mAmh5b5k+Yv/SqtgctqU6
UBmlBayjYJsMLArxE2ktwoqd88pxXkbybUAva5qJwzaTjU5MNcuWKaVhwKfBMbBnMLg/CU4XsRwG
8lMAf0h3nBKDO95VTDQ0Ip2C8F5bNLjHhkWWM40MQw93XwHgTkCZxnJAClPtsw9f4R/kUqkhZVXU
JtU99nO3atwEsnEfkWxrStmx0uuvoosq2NJR9FOdx7UbGZLE2aEx4gYayQO9nyoHoZYBc+yI/he1
2CR04rb6FxPyYgt0KKcsqT8f+LjtBcgmPKrIEotjJOSTnTwGiQSdzRojAoAZfQgZR64B7+uAW2cT
DGZe2VOq1BDv4NsgFsjGpirUJwAOpsXWpQSMSq13pAOL7aFhS78yRebIPH8J4jjN+nLTQpxT19X4
ri8QWkI36+8+KQsObyvsWeFnNPpZa4ICEx9rjOGzrB253wrnybMaGXCxfAn3nWQAc9vkF19zTEZM
MbU3RbaxtAf05CggXWlJOnHS9UcYdY26yb/N6rIIKL9qc+mIXnWzARDhtFnLB4gw+OL/avIiiuJr
gipVYgAp6rwcp1HiPwhLZp9T9RgU9axGJSsbCDqwibnHHI1YjO6RVGrdoQ2i0p2x2UMSR/asAIWT
zlnl/iE1K2U54sJiejizXWmfMiCIZz16fmHqUDFIR1iHXicL8Vb7qJr8pfG+vj2Ys+8Q0bnNqSRv
D6iY6g49CgNk2FYvheAVm/jnFY1INMOZ8J1BG+WJ7qzZ1Jbx9kxQK+soLMGNFGrtjEFebnNa4sKC
/XgUSugC51ewCeCgrq53t6seZ/dZXrWnpCbHOcwXZyRBF7BSenTmLkUxwDvdlsWuayoSQ5HhMctp
7A1OInqHwIzPmWX1s93802MU/vBmQCpRMKscR/ZZDpLqe3ffcd78s51BpQu2xoYxpPfddPbJbsvX
IdGvM4XjksA9cE4zZl0Lk7sWhDDyWNjLTlmuHiDwnsM42v22DVdVY7WuEboPg8Exx+XHB0bZ+/NA
ne84J9EcxO2pnOtwR5JHvA7Ig6iKU3ehRY3dTnLKO09nKxVLpb67osqLn+7OF1Ag/GzLiWOb8iU5
5ufk/76fOrQUv/pKylPYOVFEeShSbrs5B5zJ3TWid41uvVhkk+MGCuq+BdcoRMyYaYkmdaNQb4Uq
rsS13UKl/e0Yk5XJ7Js1cuFBziWedpaqQzuiCnY5oGK1s/0ed48Ov0f13KFvrl2h0ozPKC7QPCWy
+EKyUY2kbxixhDip9Bt/aXWsnYNgGLdIOEPH3ydlb0RfItjmHrjUpgghgc0ENvqRJmF92ptKQAPz
XRKIbxRENnBwfr5bdHyWUIoLllqG4nlJ8rmHt+tSOzb+YBXHHtJV3yW+VOcXcknOGA2YyEUdPxa7
bjG2CRm0UcrvYkQu/WbUhDbw6OvIAHEEo/Ip/OGkT0vl8z/HBU5XX6iVOVAoJ6vJn3snfCqHTMBo
5ApkVnmqvFbW/5cB0LQpE4QJwKkTRnXsSyFl1C2gsho3+9P/O246L3kK/KbzNnaB6BczsLbX0HsT
46fo3rUobYJ9yDlVap4hD9sknvBag575CPB46juoUM545IyVo5MQhQcvmHRmV7q3GtWtybqZqJlv
lONTJwTHFxmu1wWUGLwHJVyLBs0QlmlAmNL+ehxM+Zk2LGLbkTL1VezilTzw7h4dzRvQ6X5UPJxD
rhN0jJKY1SbQSXy4h3xu8qB3iCVXtNDtSMmA4aJwvczVQwDSm2nM8Bfq62KrxAY/XMxvNKVsaW+l
9UDmg1CIceLLH8Ejoi7ALBLYw7QFARlbS66NHB7REWAvi5SsFNeahaRFNvlYkM3EX37yR2CjfOk5
us4/1Rx9VFOMQfDcViYjeNweWWPLAhYMZJ532hTZSJp3N1O3OtCzdAXXLhRLGiIDbRGE6IeT4ZEK
7k3cEp2O2Vkb/eWobdAYYTKVhOmEdDQbFnpcy7amOl3VfnVv6syIMcK8/AGHPMki9WWyQXAE/haf
2R/Mvb4PYys5K0Tt4DfaqYhrufWYo+JCHGcj7hUWIvs6Mqfw/uuxKy+fe8so5wIoQ6cgxHLKP4PS
12LiA6q4EezbkaTdVx59r7qds/1GeEqv2Yio5T6gzRPDc/rA6r02ymDLK+WjbC7mBMUsNoSsAn8A
x8gCML9UNH7dZWzgEfWI1j8VG4FdDwa/R0UuW2KDz0CCNmqO2p27e1yetaK8dHJ/MO6g83GJGDwN
o8lR/GlQQgXyY54oCYOSvqlb78Z6Yo+o1MaZ2EwKzfhYjwkgJH/D7ZFW/h4bOfMAbLgKuNeSq97m
t7tHF4SN2dS2QzGJ/4En1tTTuGyCZMtQRKhhdYnRK8BtyXhpS5IHVJXEytfqjBS0KmVkhoxD4b6y
zcafLPoVNageGAbe6kbWbdebyGLEIjxd8Gj72IXg9CUU3X8Bij1v6B8mYsJUMlPn2x24peRgERJN
PtFu5flN3HUM6pAPe2z7YpXLTWw6s8b31zh+Io3Che9TxFOnntGHZVujARWbUmrkTi/aZapyUkVI
E39jlQOpOgzIPYHvOW86t7/Cxl8TV2DJn96H87y5OFAhIXTcmZkIzyH/mN4zEp6NMAxhHnd/zehZ
A5HVocpl/bmRs+TJvIF+zSCVPf/ShJB8yOob8WgyGhuKtL6UEv09e0JaW9dQKJvmcCpp9A3MhSRd
SW4Zv/DUEMXiZnoMOmvw29WWXJcurHgTkP2/DbjQrsrZtKlm4bzVCe//Bu4qGJCfcvEV6Nfuxsgl
FTOfPfKirWtbD7rwJYW6lKMGiKQLgVdHDvMTGio8ZBZb/XNPsz9luuq7Z60intmsNOHofsUWjyPz
E48Yur1BSK0NWy/dxNLU2GUnpa2eUgCk5HF27mrstSdnyGJamb0IN7373UQnAkkRHRzsXoDGcAMt
VZGAgabRrY8hnwheiBTgwD6eiVFxBgqAYbZYVdFMj0rTrBzmUsODH5UTdH9hzdAzdKhA5z4qptUe
gOMh82E/FKM91BvG9iNegdnLGtcdsc7ZEbA6mm32NUFeeFLQZGef5rQ/lx+TxskpZ68g5zINYmZu
hXUw7Q/Z6ubkvB14DgpNw091ou7RvifVUizWddf1eCu8JHIx0CDzpJyAVrDAlF1ao7DVFAgqqAIC
oTULVpjJ4P6BShxSmOB4Q3yfQVn3bDb/GjuLXZgZ1O4wrDyxt5UiV+PUeRP6H8GnYtz3Rd6P7BNE
BTjJvg8taXhLHuKWprSGbxPwjJUreBo919qvYqCtCb2mByts+vuRNjeYxWd1YsgQnLS67u8U4w2b
rvcv8KrkjnWZDvtH0yF0saU+pMKzu1yLiHJZgO0TEZGwS3Nz4IH4cN/RsvJ+nGy5SkSclUnbVFAk
Tn3xtatSQ9qaBU5h3/Kdc94mBGK2kN9wrNwzYLdLYxvQ1vRpVl7IJFL7LmGDsuDpEqGCT7qR1qXc
HAtLgGcZi9ReJMgFv8yBO8aeRjpeNtHDjuGeAxmd8LgeOjYiP4aBwKl2Df22g2gtpAWqO6kIiL2d
P1jog+q0j3MzXqaznJeQB6zd9xYjJ2K1DeXaNMyki/u3ESNW+ICp40rkXqyuyeA9sGms7v0mS5uK
S4pAtpPVmtsBOC1i0Q878Qib5g1CzVoF8uehdukr9b3ylS68tI/gRCfy1w5nCHF+rYkx1m5bJ9E6
GYc4hBJ1OySFECauw///gCiXEAM6rrox0konUfPtgZLpNMp98cHa5wt+RUSLFPUAZ5h4fY8eATry
pzc/8Hsvnlt61EpM+naubeHFjMEPZq2PlKP3OAnJdfq920IyY87fkdvVCf1octs3jDk/Ta3Clku5
Kt1/V16ukmxHf6GYeMZasqag44V33m6Kp7Agta5RE2JXiarbFs5UBJRETCpuVbJKSkDdrjtWdFC8
aGTPoGea759kMjWt7Le/Y3XDSW7VUAu3EzjV+VYjaB6Afc9IubScpxnIOY6GgqHshUkEsSpdySnf
C6xRqgb1gKwowRcqcLvjFpYIG8b061dZOqCBNzpexZNW9UKdTUZqJnmiHF97cQ7VuOCxFgInb4m+
89TtCxAoyG40UxvzFxXEk6AtJLpI87Bv1kd6Pyqp6KJCQcn4DTUTh7xLo5k1UtGLx/POAG8PFqUY
VFlrDWsTGzNMYChhSfZfAQ6g730YSxCoBAE+yGHXv3QNGqSGQWNbzw/Al07WiNJIh0N1exqyE4UV
0IckMgXy4ST4qRRyzIZ5bLY8DfaXf0wqX9ffYYB2hMBdrOj8aPJsv0AuSXtrrMmE0dBLPt5vnlx0
4586QYI4GKxg6dhkOmKY03K35C0H1F/fpwEB6zjRzFE65+t3mjoRjxqwG48UfQniITekIUYuHxf5
o5Mhe04iLBCgK+5GwGDt56mr93g8r3v/ijGxytMuBRQ3uSHJI5YRcIUztmu7wXbGwEXzEI/n+aiF
FjpLruKXWJU8uNTgYfgo5/vuW49ybWXExHe0Fdt4ijnuMYmRyCFao9ghkByMSyn7AzcME4+LvhIL
hyZbKS58r6Dw2F6RO63Zuv1eWEYMeYqFhcG0rA40zvJDpgec/6lv2Vx2Ofku9OklyEGnzWhGLXaC
eSH6aUEpXEd+MXSbtK7yZwKB2clhGhcRHVf8BuLILPrjD6e36fFC+mYqlkAiUgNzP6XDEmbXey7u
VFRklkirMzwlteZxMAA+FW+fIsgJxPgdJhg1wQdbtiJbf/HPmLC9eZL/pA/CKQMno7QnRNT1F/4/
3KPY4GqWG+3iekjwH9fsG2FaWqco0Cwzp4j19c/3tRhfkdwlclJeWXkCrWdgmTpRlG955VAZV58m
YQx7aiunwvHF02dN2e4SIvPJw8VPKjAk1Q6DffFBefbZ7Bk8u5aY4xowzDsXJKJbg7DZMb5QTElE
kK3OS8N2qxXnKtwvsj88wIoaiFbUHSDF/iwCPTDi788jKhoEoPfcVyh59lWJ4VTG110jRzBs+hxy
3brQwLA039rGmGG+tXF5rXdFFmQ5Kh3F0Xn2MkefabA422+nWiUrZEx/K7HNJSdzsKHZDPItzCPj
fTAKH8YXUG97v+c7iTtKQSyaP4EjflvNlyxpGsTIYQBbJErSEdD67AqdIQog0VjQvHpsas3Kh9u3
DfhDJzmx8vwBZzPKw3GcczRn8lmI/y7cZceUPQL49f9DCFin44jduFrQwyxltAcLw0Ef688nQVGk
nF9gphNa9OH9n6aXEN2XWG2WJmLLGXFifZ2qXAmFZYi83FLGuOUBbKtvmpul+7CF7OqZjLewm5Gr
WaCpRTKuJdW/sxJnJqyKvCu8luLuT1/1Scp8353a1F/xiSZ2Rq243iVJAVGsqzp4TtwOhYUkvcpe
8BnMG4jkhMfAlHawBBL1zDCv0g2BnrU3/oA1Dr7J6KXnChjf5ctMPNHt1iuS+2WrX9rarnqFpaEi
e5TVPZBsLT+pUWjT/t+WelBBaIMrz/K+SBxj+26b0u10F9sAhF9ZGG2r470SROKtYMp3ezzAPo+Y
wDGo/Cjy74qNJWl2fWFudwDsObkQy44I/XYf8qGbhbCBWI3lXWbFC4yKFbEwhXeRG92gdJJjeDKW
f3kooOit5+wAQE0naYsxtSb/rdvF7p+KArfVMEG6Kd/qYva55fE2YFbcCDKYOkM21Awh5bft+4/z
DxwuuJ5VzJti3rYqp+9koQnr6lG1LsO1XDf0KTW+iZoxdqPVXAdA6kzlXEZRGeVXhplb3dUbnm0+
2FjohHAygdMRuVGO0uAPIo8KQEml+pNLMzjC1NZIExyW+riVscWRjqe0NUM9U37jH8Rg2d/P79D2
Lb7xsbqHKAfogE5vXy/Z1paH/ghejBx58q+ZRFigEFSwM889P1mpRf1MvvEYE8p6/6SW3yL1aJun
gvvqyAuULMfbtABbnvRohhec3pkLYYBoVwNXsIJ4BJ1Gv51a3k3ZtgUVFU4bsWTbD0XrDd5sMWc/
I2QsCb6nM6L3eIhyy/p0F3A/3ygjm0iTt5wRjGfk8hiYm5vQEB9m3i6XtR7CgGWeyYhxyTtKgiQc
vIz9kx4QPev87IOKgx7jdQ95f0IJFRMXAykDxVTAfOZpwT8gTCGIIX4I4ePuqp9aH5kXtXnc8PW+
4Zwuywvh4dlqOpnm8BNwYUaUJXv5ZdBcpbkhlL5W7jIQopN2Ef4SEQwXxD7aKujwPMcRxXcZTqsm
Wpr/FXG79YJh/H7dv5LY5H+YAA3Wz6Xm69lcmxFZCkdyD5UCM6t+O/K5ybnQq1W++ibsRvvJvtsR
KZwSrfDvnf/Yosu94gedwXe/VDKxkqzMh/ktFnTNi+7vUu8bJISPnI+0vmqH8mg67wjHpFYP7VO5
ite//et9YGUCRTinYqeXH2xpv3NdBTPCKRH4gV0oUkKVI71Chq28O/SsH1o1A5NbONqosoicZOhi
j+wsw4QsGYQam5praprMJq8A0i8r+FQ1EvHXOr4ngCMnnulY/3ouJQtQ3S/zwTgLATKlHU6/GyGF
U8qqAqqhQYUKHDuemgnvCpZ/4RYtYyZoMzPjnnqS3U0tpo5C4dR4G9VoluwpnGoyiEaWYs9a3QrN
EpaejQeqDNPPObDSyYEXgDLDaob/tt9TDfEHcjSCio+c0dciO4WvcOJzmUiz9ep8jeOuNtVbh9/6
0EQnkce4FZyNWbfeIf/ej+c2p1bqFc4zsGOZUlz0f0OxlI9dLN/7eWGaeV8hTuUVDgM/XSQ7W3gx
Ywvoh++G2Z1TsR8DEEX0HXsV/VAUTkYjidSiVs7qr/fSJH0dp4uTviUrzjj42z1uTYVoUBgFhxsP
G8ntxwS5bD6QAAeJ8HoYvzRUEYsPbSe4J0ec9Vm/Dmvce3GhQrdhZ4EpYSZWshvagkypFzsF2reW
F38Zy27uNlYGhssJZg8gVe9tuueXvsr+buDvGNiMuqraPIhLvcojOCPmmu897ml9U3txk+icksTB
4jcCrS7JcEc9tsYp/7epPMsIXL3MgmpE1CEjIx+dJHgw+qRsyBBFXl2meVSJMlVRPmnsxet4ynJ1
tWU6zKyUEmSNEhtCGltmJJEuKrkxDd8KV6UzuqJkl51JcHwNoDIUfpUinJvRhy5LOz3RwtxR43vM
h+cqahMXV1ZZXaeWT4cx5z9yeFJTjy4WgLS0CYY9tlRRA1h1DEhPDjxZGXMSowHsDKgn6l3Ntc/C
GApsVg811w2I2qQCyOzwKY12oqp2HHpAG1MaT+fcXsYHgdiRBtAi3qsqEoeMWHOVBGh1YQT6cjCX
o3AIJDCY062dk9QiO5VPWR79bCB3bK5yPtidRigFA2H+sUQFWi5VBFbB06j3AtluNjCe1JJEjhNE
FD7JRklzCbydtsgxS3uZ4BQwWokUe6IylB3qCn5yT18bhcvOQFZT45nWmkTo8TsCrqEOOG0EHTIV
bZ82eSF2tQgU7nmhWDmYz/JKkZNtUO3ZkHdxc6DxT4auTdTNsbDwJiZ0LmZrrZYOkZFFebv3sg2D
oVLH0Tsg+klnaPzpu+qubo4b3qGhcV4MLRMwmu9Ge2abvbn20jGT9ey5jkCaPVlBZdkmvMsXpLVa
OKvHk4/DIECJVGfkA+7btL7v+tlxBmU6AGsF2LvjNfqa5hzKUAuHSOvBODLI5oTvvEWsbnMQLsNu
8/cj2C/xDbqVmGpnKsYSmdxzP0+v+cwlSXGI+NlDpZZzbcPFdT4uzYYnu3h02O+xS7g//mpLelUE
1Q8kYiRj8m2DHGSb3NIUWW2PS3x0sKebxYHSoADw+lZWDs9KbRaYm2tky/2HT2boNxkAFVtWQbKB
qW8K9q96snUnegMryMkxeenQI3SmZDsuKvMu1NXBEBsZiFRFyNkVTLCqIH5AWgiqF3wRfAFgFtzC
FktKxX0KdxZstJmmjTYOQ2Gm0n9f6aeZPJzr4mJVUml1weZwM1b1skfb8sIbN6xObwJnVTiL0uQs
TPM6EOfOv9lbLolERYNFNOstCfxfduZUfuO+wh76qgt+5FPBRPGq/BZN3esvcZFAy32EHIc9rcUr
NZ2bB4f/+vstN75odncgiORYzGucfyYWtLl5fagM57eOAM47Jt5+v3myS3qYtiiVqpz/QTLwWaK0
cAAZTCOyshOwggsqQhx6o+sZUo4B8h32Wwgr28H3nyAGYAuTx7xoGy2mSgmIjaUGByrOUEuN0JY6
siU0SGXCKCoPkdVzh6lbs8L4RA4ZmYKxewCfJRv5L7TaxAw6AnJkyNZBvluO3XyLXV4bKWa3tqbn
eIZbmBfrZWZdY5cud7XssUSocNpYtWeUkvLIroko7kYSmyRU0B/6OsU0QrK3L+xsdLEVPoDvsgZP
eE1iQBTKECnDWrLpRDJWfc5ZyRtlNhkjBZkdTE2B7Mnb/wDceyYNDWPzwaj04MZS5NqpTOnT5kMr
b9/88MNDtkqH3u1lDWQXeMk3vOYaKCRfKwCyR0lCtnFccgBGqAeHTa5wlELFqNSJt2BQOZsQE1jY
7w86ojWtARqleJbtY3Jb4g0jB8hkdx9ZH3QHdzRI2T/66sjl1OQzX2AsIlYVGyV88iAS3Ih2dEY1
7MjKrJs1q7hjE99CrmU34QCSoqdGQgyXdA+R4h9YZc1Pmlp08z7gtj2C6ZfY5RZzHSVTP8HT/4OB
bK5w5Q5TNFyzl14lNu/ILbU98Xk2eURB173pRv9SlKNTOeH0k4aJ7ZK4OHZQ+gAlALx96Li1t7+p
ypg3fyGiCqpV9353q6bG6SiTF1hohz34bTp/xPar9MFisILj6lHUS0rVXtVgCM57l/S4R+ThD4C8
MLpIfXxTpmF3jQYMz7iFUmF7rFjudr4dEM0POWF6ERtroT+6M4DwzvRVvT8RNvmehld2dVDMBZ5x
sR3bbz1povrDkiFO+tT8NfH99buzrbKPVLsNn/inf6HkCtausH8v90y/47UiBeCk8Z6ygCRfYljq
DDycbxJEtBjfB186G7CiQY9edPG+5P7e7QcgxBZzhuS47AQa2xJIYd0scg/vmw/0/HCqcWCzSPBW
ZVWP0G7Jy7Mi+zD5G3cBKsV8kf2Rh4Pm+6/fZWFMGgGAWBNLpXCfhEn1VVYkZcHBXAFSVbJ+cSV2
uUMBMRWZva2EdeVOEywn2bAeHt5DSW9jsL9cM2NOM4LDSnn+xFABDSesrl4cd3a1OSdW8qDfSGhR
U0pnv1Bqw1gf8ONXEeITVPu+TvQxEjM3LlC67etEjRN5qvPLP4ZgLmJdmzkopaELoamLdmoZxsJm
0OJkd6tlumYMa5bJG+zmG5847JhphNLyISogNb/742mOkFh1s6YfnWczHmJ3/w34mdjC61xuaOjQ
COASrnUU9OOT37/0ECeBgE8fxnNzVrie+nktUp0P81Pe38uPP4x+CPCK528prxI2Vxc6esbeaCMw
mQggBBukrt3itzuHy/S1frGjUKdfCIbYuh8am+TPdMIbUJ3GiBdn/9/3/KapSxRUAtTr/NUxkfqs
BjaytDKAVdsMEmpJJi8vQhZZLfUVsFIlEBylf4rPEpcmwGEQQ4UCcvFQvn17/mN18NjTi5V8pLah
2IdNWCM2T58ut2Vu3R/AMJlWVY0doRcgb4M1QNJ23yj2ckGgPnKdYc4sy7q92kd0eNkQFMF5bvFo
8SkH78GIrYrod4pog9UEmSYi02n7427uOPUw5LQYoXSDEbF9Dco5XCXSPn4dgkpKsAydx8z6f+Gw
U3skoJi0cb+laYcO9kjfcxMR8fZ4LSbVIX3wUtPqxPDrU/IZ7x4lW2hXQdVHnKksiW/uDS2N4tmV
hhRbwwF+XJBaI6S/BJ96GlUeCAM8iXNDqlWdJ+XnGfe/yDoLtoAzMWxy4SOg2i97aFUa7cBnognt
69SflUtMy0dFtPpQIfifl46Tl/08VBKZFf2dWgW/pRPixHgLSotmfu7VzXxbopXjogqunYzeovwB
88ieXFKOGL/T3rOaMKA9BICJshhqAyMJAIpoV9Ia7eJu2F6vmpGa5q5+TrhR7W8jIBZ5+UlfRD/N
ReVp6XQ9OPoYTnRW6NGFw0TuK0OE4b110a7gsQnSBi0M46ORLTtR5ymoljLPSBOeWks5KH2O9l+G
NERt4j9xMpM1USqiz+Qe4gkSBXuqvMM1MM9SU99iWNSllBkouFCZTFKp8O7TiDwDq+ojtiMTJOUc
LGMslPDoLyNlibG43O46eAa4gqo8axqgzIjkBleId1wSAZQLKlqhM9/e5pwaVhGmqYJaJmzZ7kqv
ijGyxVzcUCwD2IkkwzytO07gns/PAlpCXo52Y7sR55vdP1MWkjoQLruF7CJwawNAQZhgib1Y6Tij
ki0IXxwh8+QH5mCV8EWnxTEM85m4A3bQDxNMjrVcGw3UhPF4HCy11Da6ogcGn3jPr7yy2IpREVuK
3qpfl0O4sTL5d+Ooj++pRtSP+0c+3FjrdqA9gNfhg6LdJDk1mPJRmgcT6pUtp2FEoy1kJmBINKoh
9ZfzIWFyHmCxk7tR3ElljTuvOzOEUQMQa8FA0DBpCrymBax1mtoh9o3tKGvBL6wPiqsCtbAll1yH
bUME3T4J2DdDetFpOGSextcefnDRgoDdbpx6749A9JIQUXPKsYy4ZHEUd3N53Sy9d9fe6RRKqXGj
grxwMKy6mcz1X+ujHZHiI4K+mrRKltreLXsrCZnaNJr8xw3W4abnfXJ4yhxHKd+95wUo+ZO6sOoz
C9GjdeyNXySyB6dwC02gkKUmC9US6pDkgLty6Kw1HYszZDBtRObOMI4MSxWKDsOOKw9tlHyb+KQF
DXZgNMNZGFiiTYT2DVaoQAY23HXAuY7FNLnSxL2Vk2CQAVefOeiKRgRVOlIpw3Q4rFQqpI7XaUxQ
bxoWmP8ttMc/P7F7SYQqJKSVLORnpJw99QVntxcrPpwdbTxC1eTuXptU42aBHSkeU5QH8k5wNArd
DIW+BJaE47Gt6iDTTSou5HRfMRO6FCjIUh1vL/tehuNkbzVuur5BWh7OwZp7bvOf3ig935ZryshL
ONz6GrfEYZE7b4A6FMHVQciQMLJDU3djoQOCBYIRB83RBoMU7YKO/8EiW/xhFroWO2F4giVzoL2U
m5J2wlrR4UyycjuiwmXxPR6+I0LTnnP7YKsGMqGefqLthhGpx23vgpdWruA5oqDidIV917TogLJT
rFdgmg6Ihc9M3FstUu7pGilc31I++/unLHS39s4pEd1jt24r+yLTxHoh638eKYFf7MZ0AmUaNPlQ
yS/x/iXHeRV+8/D/VCpvjvsgRrtqOrICiWBWlGf71QdBx0UD0ttyF/4y53rI648rtN4zVCCMwg6n
4vgrLQLvhpZ/Zo1ALi3lhQQNNPorzUVBQjKXui+EUXMmtLQbz8E5pOxyxxvD9GbsEMkDbWwaBOhA
83QY7SaSHZdqTkQVWmvWGopv07j6wMk5IJAO8Ckp1Ot4T3Kiz3dG5L4DlFJdF4gQlWR56sSsq6xV
XUU+Ap5k3mPS00T7Yy+cDuMcLX4yblUKrPEEqDAQiBMb6HUrM6ThsNqz6SAyKplBAQGlEKqenAjg
Jrw82Jt4C4N0OO9RZSGSQnxlzHytQD3eypjJkiDSO2Sn0+AR27wHLXDpGqUa6LH8JE8nBY3OUEoE
PcUYpf1Ze3PuF9qkC9eYCZN626tQ9NvleAt1xp2oTtS66wKhn2qHFkEQpJTxvj1uNmS56Edw1D4b
96P8CYxfekyXwMZZ0dhJUewxUxmga5Y+SR1sj3M34u1Y4lZsW8kh0PCEZ5tqGNn2t62Uu0wyge5g
66EMq5eqJNul2ygLku3uSeyxAVN4WtM7icRbdFn5ldOh7AxBcuqfx0HoaT/uXxYakRCt96f/tWMz
LLgijtCOYlzrYBLCUhqAGs2bsLWgsI1aOMFAFE7usHWjOC5vhNk8y8gEWqj2A8gyp+mlhNrzif8g
jnCasHcoXJHKa5yz4+f3ItSpDYL3OCtWJsY7oKFjmNc9YR5hr4tOx4biepWMiQv09loYnpSX8Jma
oH9iNZgdd627s4s+ZbUo+6xhcMWaPa6CzGEqMJZ3/p84n2I50sKr1t2FD78DBJAQc7llctdmD5Zn
l+CxxduToVnudDRLoasphxzc/wivTZVAoM8SDMNdJA8d534hIo7+2ccCw8uNaYcP0mkHv5AtJB/z
L+Vpve/s5lizYwcE2yLDoVCtZK3cxKsuJm1ZJyDpa1e3eCSmV2dmXDWVs/trvROs3cPJI72O4iAo
0PWaCE2flEa7IH3GfASdeu9XwqmzctJF6cW14qFVYvwRIoJll2tbfYf8u9LqHrXpJNhBijE1g3eT
YYrA3YBLovIyaZRCinANc0wQUw9SgNADAe2T4xHBvrpQ7oFEp6k859lwwrdD6rrcDqEaINxWimo8
zd6uAQBDAtzZsEi5pAOB6h+Lchqx7qjFZs2/ie80Hs1Fg/uLCmjMBt7K9cDkELneGDn3hd7SXsh+
r7sGqzhWBWRJtgWspaCedyl5gWrrKCsALAuON4VSfUusSwJ51ygQZDCk658xba1/N66XOXwVu3gP
Gv0uvBOUsX6JOMzQuBuCxfFNmWJz5Ii+V0bcIm05fhQGnrq1oYAL/qbIC+xtarmHRTVpPhxC6lOF
TXwATwcDCV5h+G4mtHthjEWAEdFXIK0yYcelXA3jymIAATy+D+qVpuRuJoEfreOMc5wLOqaZmqDf
cSsJOYnjLIuSVfcZZQuSdOpprtoW8ArirgskZF5GjYYQDfWieKgiUmHmSIq53ujxFpJf+1iXPuM6
7n6HW3eihEvLWb0SF+1CbObXjBkMjFgBiA3rIBo0pIzKHEOmb1woWti5nUGozQyrSUfFF6n9925z
KfFpSQTpHIdBaq1N0D96IbIO8SAYLGQAYqL5u29iMNxzpwpXgBZC5L7Ge3+qjyTGj64McGu+jirY
yarBq9fkB+Rzjf3/KBKL/CfsKSv/Z8BT9XJnq3mdA3cNW5wWIEJQldRremxccMlz4EcqUaohe39t
CJ6NJyDoGjH8HIeBesx21RoDVhb3uWRfyCIiFNFRWzbP4nbIRnWDlPu0+z13EkFvs5pdV9zYYkok
CDfesBjEnr+7RBPOUwOw7PLTCriKcDoqrCAgoCTP5+ByCNCLEz30I75Uazu27AGPUyxbTXuhhAA/
vSW2dfQxah40c5qLBiLuSvKvS5j83B2lkft9x9R/RrHTA4TSOBK0alv8pASn4zGdhuXJlr3F/Yg/
tzHNLnHsZ3R09ConzhwJ7BPtYhME/q1ItZsJ4CYUN55Z+ES8oSKmW6fypt3ie6YtglqmsDRxieso
LtWO56sYm7yuuoKOih4lgq2f9bT32XfEzfipC3JkvXuDTaTtUNUoaBmL0Wn5Mfh6y4MDE644ibSm
waQTNQMXH3xJmQaL8IzdKSEdnGvD8DdWN3mY7yD/F1QY9D4F+hGjktjMx2lHmv6nTPFJgCZoPUzg
T8krSJQJBW/l3ICWQJnklwTWhckPIBxTtkj/+2cDmRC04ytqVsi4CGi+lS4HcRnWx33Lxbf7Xcyr
UN7Ve+4vhhwG3AZnX++d8hVndSwXOaSp37rBn46TdFCBdXGZo2idraUF7je1LzvCrmMh7HNtF1Ex
xc1Uy7vjrgPjfbxGZvzGsqXYJIUWbpSQUNP1z4C7VhJuca3jZIFQDnXJzIhzljpB8Ey3Kd5EG9J3
bw/GxiQj8nZmO+lbLtHXHxfy69yf4Ap4Lc3AgybESMYdgiOblaxaIkukpbNJL+BT5kdNQ5HZlgIP
9NJOPYmaF57ZF8QaHkYM0xfWsLTXt+qXDaY86e46ZysUyW4jrr6uHh6iSdKmA5k3MeJOI0N7Qtt8
CUc5w+3cxPZOcpto4fkRcmPIQjKstNjzMWDZgyiIdc19fIDb+8Hc0TIJFgWX8lzJLFBWQw9OjBAE
NfJKfeSDoJr/DIlQl9/YMDwAiHLVJty3pyPBGniK16b6pDKeKyPCLLqMKytXiwv5yUoNXBnLukJo
zYodZwUwTTkNCsW+pQkCeFc9YvKMz0ioig3NOuui5vVjGXtmZN7DPX3xQazkOnMjrAVoUxB33mh9
FVW5c4PoYwaJa8dMkvia5JLqZgNxFqQXg3hs2sZomHURFAb3qAwGqCYvxJEtid64z8ZWuIpP3R9X
L5CmO6SZMfVfenA6rd5B36ZgkAMHkJgpRLDarMq9NGCzP1PXi7OOy4J16XBQv8O2pa4o48ETGuJL
0IC8CTkdLF05MC/+/grIC+CEtwje9Z4tUHbC2VopXjA0bKCtzcrjQhh7lxpS6plrqKUx2ngyilUs
4rIYlXbFfa47jcPmeiiCOqHIzcmtQ4Q/wdvuskD3gwFKGupAI8MVXA8lItWd0RwdsgRzCV1gqhFf
gBdSG0Jo10CC7N2C1gvKoKg1qUJLDKUU4A3AfOmYr18ufPYjuLkbkC8E61zmstOE/1KLZKmFKtAj
7Zg8dPodU+suHDZ5mua4Mk7ACbHWPp30/j+ETxnd9bNEYL3oYxVmTGCVZO3s/Zrj1XSlMQ7mbk4x
9YZFM+3DvtSEXVFZWNA2i3e6932oR32lztuL3vmZQJ+d66KvDfmdi073KR84n1VsFmIIfToEi6LM
IhBUeIK8wmzl2K08J6eFX3QJ5xnoC/Jz727IJFxR1w9Lg7ya4pngYBgpFdkeVkc3nqrOHg7m8UvB
NOhsLPuA5hUCYoe9VdChkmvGnUrekTXZfUlFsUbRDR9k/TFViJcxfnz5vvTLMlMa1es0S+ve3Ngr
YyxmQ2UpJn3nknCwgoT4D+njMwchGljzd9rC4kQwsj6fOwiXJSJBaqY2o8mzKuq2gOAxeZcJ1LRR
0TllbL3cx2HY7ZaTPqJxQT28Z9sHSpsfhOCo1pgHcdvjseWEsiZD6Tt4qOKWBz+rbb0QLr4u8e6D
GFty5/JK10ZvgY6VCz0E9ft0rt28SjUng82vFSEg76r1FoHzlTuM3KoYv/cmRrdbijp5cGjZmqS6
0gfW9fRnbna7aWyOVDDug2iFdAtDPpvrxoJJqdyj2Nq3Mcdi4xfxXKzjJJQkWTI21TSkRjMdI8Z+
dO1bpUWIy2A8dHM2oj0BrY8gBCvyNkVXc3E/Lx0bMPj//W4MjVHOenlBKcCSpa/BNN3NNQdFANbU
yhSUVxTGgweJ/Y4HYbZsI1MG0pORmAG9UtnVf1hRUSayrAeC71K5A+pa4vD8JBmTYEYTtw9toAv5
UUJZiGX4DdnvrlR6kOET8daftUtQ32RXInWJGLuJR4MsnjrJk8pfJzcMDUuWRBJNPqXoTwzm8MY/
ZH1G+rw9DA/CiB9s05REbLWxOuZnB2DtjcMZHDwN6Mf8fWtBScTWCeLKDnZnXwIJO86vPsQVubcJ
/LgXbixo00wqvoIPvDFCC1Oj+P/U2i7KJgdSA2whf+ZFlQS+FxCVS67NptDu2mLFJvwweOlUxIrd
QDqSH+QbbDe31R+x3W77cUUUOSCZRQp4eqzTXnrrGNx1lVfM3rFYHXRyeKqegeTVUAsD4G2TyI7S
972sEJMBI9XpsVyU9a+fv7aRf9TKPTQ6fCoGlIE05fNMOGAjrcwFwHiIS4WWu2S8YiyuPCyw4HVd
bSwxWFCVhdNvRghoy5+jbPcxiNcSUdpK7Nk5naEXXhAIegwqgqKal2SRRI51Iix26TvdYwydKHj8
g2rlN1fRusicpalUP4A/2a24h1qE6NY0ECnoO5eTHrid8rPjCEPWoZs+SANUqFCmorfgqhitCpRF
crl+9/rBctHpb8fl1MXSyLntdTGe4MzzTCdfSB35JKBQ1T4qxrZtWmosz64OCMOtVcl0ByQ/FFLk
hc8k49S16XFEGxQ3EPKtGD6ujBNFTAfOVwZs2FDNIjfYb2UePQ0YD2gkvdkfDW2COJUxLsDCF1nc
+9dK0gRkvrhHoHoaLu2QMl3CZXV6HLiXttbc9YhTYmp9AkQoC1nKeWavN5414Xj1M+QAq+ROtG+g
lL6f9FKWGBdf+hEPNUktj+OBAaKkIxEUjeH+v8GjtIzMdCvAyhjPRTFHmrTBMhaLVqa82fAWtkRS
F9SJsHmY1bAELmFbb3Rsy+AgVwrsfgSG0dxpj6lZIONHWKTXZt+FDqgOCRWm0H7pJSR/wp9zfAbS
FkIQ2vLQHtDQwUPATOBwVfS0FCljV4Ip7Lh6Q2Q074goaTvOVAXHmCnC/80BmYF5Qd34L7QKU04o
8pwZFmU70RODtvqCzclMYxVcMlhc204qsudvLhmwRN3wGFAfEEolD+qD0A3fX0YctBtPjHq5GCOr
K0fgJMx4J1AdHATV+a99yO6RW2jbYgbosPSqLcckScSQXq6q5QsLMlHWCX2zJiLTsc9mJQaVJwnr
TOEFUmPna/pZ03CMfkt1qRNNcjqGDXs3Oh9IkTHt0drMPJg1c2l75wf0O4JR6FcBhz+6uqU2RzyJ
BxUs9mJZeCeF5m3KA3Xo81h4+z22CPQTX5P4U94UrxtY5e/KR/BIvfI5Hv5LTInEOF0SZA48hg2Q
GJ4YCNhC3DvmXJ70HPKqK/UP1ENvis8fi8kd2QhOhnb9qaM9U9Cyb2512PRtudY8VD7pmMgYXa9a
JO44HprnB9HkYe5elU3x8JQF9h6lfRwk7FcExSRhTSRaKWBhxjAzKeMiJWKqnuAmgKacEGEJtk1H
SqjPbYq6IPqS8RpsQd5E9mUniCoXX9SzZqb12WCcHSmN3pVXdEz7xHiLeS5azzLYnU67xDHtdvzo
DIjlrnIqaxPbcFIX3f0PDleB0ZTgQcFufpC0pIfeqbM8GVuzb52swChlJ+qVrC8B25ccL81PALet
uOX1g1FtyOHvK0TfbEbfOPFHD8xIXys4d5XXTT3REj26xObT6/Ejawk1IBCdz8XsFam4AYfXhMmq
kOjz9ywSHSlfFyrn17lN2iXi08RovasmG4LXxPF9F6HifOtE18J9ryoLAfPwbenc1Cwq6aRVn5gk
0+FkMOu5y2/YPBAEFbGrnSLd6/jQbkl8Rwea0WBPu5EFhzxnN0BCI3Jqa+MMOOJ5mf8z3oEfDXTs
AJRqK3bXR2mwzD1e62MnXAyB8ok4ypuJnUOdWpiATqwRXjB3Fw6HmD6m5au+onbTf/2kTZ+cd3wX
u4X3POmOyi4Z8wOuwt55k+BMnZ5UT2u1mlTh1I+HfP+xRqfcchIvnYuekCDhRXdo51U+oHNq7Nso
Isbs8SnYW7KVYUfG0Ad0yNFZtGA9EpYMIAr6AOi9zvwADm5GRcPclDbQPJOP4Ebz0G2KcpPilb+t
vYWngKJgU5PMLcudZUtdRMdzgR6+mxIzcW5jQyYdy5UQAb0wCpiIaAJ7NqGGhuYtTpdcKfxCdFfP
aHBdR+AifCIhEFgMHB3RmwiPSW9f147uHGP3RcGlwqjcWiYNO/IX8USIXYYklRpRW9jim5HS7Vm5
08otmyXFGy7yaGOQXCLSEfQVYRTDVCXqc5zUYq7qXrdtQmG05GLbMs2WOPY3UkWtUVZgxHksAC21
C0oAFtfjgBYkhp+lCeLD2vZmR74w788/WtUEtGp6/iBP2jphjPfYj+IF99AycMGhDHtrYTQGjNeL
CcQjPnpr53DabJOPPaqQin0nG9rg3a8FnPNlK/V3jn3SKBi9MPnzveWhHKMe/Un/D6ul3MDqVSUz
KEESXZmBYl+dFnc+fLd/I3eP5TDaxLFWMSnTTIrFMRVfki1+T5yJ/bbyVlJ+I+c+CUw115YurR7M
nSydC1g/q/3EAmHEOJpkxaNCf25aN9O1V9w0XZ/XsKwQcCLJJsdRALsJe7VnIYYetYy2r7t/HDPx
754Bv16Up2Vdr02/4stzkK/2+CjE6BEZVUP2T9HSbjkDNZUqZgHHOguOKqn+uqFYiQylKyk29aKf
Wh+4V8qHsfVT7977kRfqFFKnm2K7R6WgEPJpNGj29EjDGzjAzEKt+1lzZ3vsz3PjfeEde4Pb1knL
sMeFGdUU/yw5cgWQhvdhJki9Rueq44z/J52TojFAvcLaq+5ZLJzVqoTZb9yKIaONPpvY0UEhfP3X
NfObywaqX9uWIPL2VyGOpfN39G14LfXQu3qk6q7nlSWYb+5gpYlP8/ENYHLYV4gwLEM7Iokl1LDu
C3vNLKdH7Y4nWZsfjw42/2SlvUiByrl83RLZSYFW/BZ4NTGojF2xswjfC5MgefJZtP0hmyD7XokR
i7ok+MI+qUYwhfZAAq6j2TmznVYc1eSq6XHZM8dmL8P92+rrllVg+FoKrtLEDYuJ5T8PSG1foO/q
lwM+n3N7dblwUHAM4siGeNad26MzP9cIeqThSHP/4CLZbXY5Nv+nUSHfgYOhVpxiCub5c51v0gw6
gQX03vNpGsELeaM1NIa8M8rJ4pxInqSXDXO/DOrGRSJy5WKqJqlAPz3XF53cW0zRjGajMe+3oflB
Qq7fJWj5vEEYRZzcjrc3JhAah/AahGvONlZXO5T21crTKH8zy/LqeSsCcMaid62OpuTvn0tcM4Kk
5veM1s1r1cxPx9M4VLKVlLIeVeOgThAah3ELirppL6itwrjFRjx9gx2/d+3auhTPqG+bh9Zm+p6O
5gDjvYabK3/G/cpedOyC+hlhIXdN13+13aQNyPKf06On62eI5cyZHjeBIZCXw2anCMpCK2arzlIW
6EmRp3DuRza0oe6cFNRq95DvhA4yQmeCc9OTg9uQDehQ9eUtehz8CdHLFrGw7sbCXa16hU6Kk0pE
grsEnVXx7d7yATw8C2wAklmGicMqAE5CezK6fCLUBBVlJM/OnbRjcFYOI05jQipkaV5mevhw4kaH
ArS5L4TJ8ie4RX6BTHqyo+nw3WvZFx9Pa61K6MKmHXU29G/rD3q+gWES9O4yMtNeZn6LYbYFidhP
OjGCQwR0OvjKcRhHQeJWaxHnbauZU796X4OK54Mm/z9VrEm2eWtf96xdecyfV67GPVSnsHPV8G9P
t1daa9R0UbzugUKOmYjKZKQscWmmVodDabouEVLzQeQH2IqwvAvvXYAOBDcVaFSeh1P2/f5povf8
hXTO2AqWKH0O0fyDcCGAGBNP2xzvqfo0ksoD5vnmw6xpsWzTAgnjKyVR4Y0W6PMrEVpAxaWtSXzp
M3fl7suG3sA42FD2qG+a00S9uOQa32+Nr8lGb2ZYf4U1mzNvfp3LBKzBExmDxc2IaSp/Pvp3XWhC
SHHbf/hpsPegZh0OqRcIsoUDWZJp+qdm/JRPbKVeG9vKQT0wHQG3QjY1cz06AP3zz9uVITkH+k64
MHyR2ipwV7Vx9W0mimr5iADM+biyyaCA9/3C9LfUSSawwcIfPSm5fYIZ0lzMZr06iBhXPavZkIRW
MNRiqeWjRUlFG+E+Eh8RYoHqNJjT2JKs/jRy76y7k99DZRi4KsJSgllyhN0ZQi4Of1JsikwZ1dF3
pgbfSeHYHbniZqAUyOgMnIqd8/S5hcEEgJDkqeyT6iUIRrGp0F70j4MhXmpQyG2T90DJowSBG5KR
xugfdqd5PQ2NSrF8VR8s6a3f6ldtPYWJii8cLDaI/JBafnPbON4DpWiAsAHkOrdQkxlQvQsK7yLl
XZ1D1i3JpLPnbBkqkTWHZlh0zysavsggLRbcGjb3eDkF6Ky4IgyzhcjDD7brbaeL9QaAWoserjzP
jk1CpK+RjSHK0znG8X10ynELXROVOSG0EQlChov1/co/SCds6xJZxbFetF+4EatJaVsUApu++5rC
djedq+vyUs1icz1rXqzSOjPrUFEXN2PAO4FxmIKjBaZ5uXPTIha6HCleNpAgxYVNCEpRr5U+zXoP
2sd40yWpugJLwmx83cZhzi/2luu3L8o9PteAt/oyiAE8MTutxJB79ygvJPkOjuMWUcYUsuKl7Z3p
/wIEWKCswdCa6WiTVav+NJOcGK9WMImzpSpFgNhdW1XGC8TNpW4mKL4CpQe/2tregifsbJ7bRdRX
zSb36Mh07I7uPrY2a8NUtQ1X2rAlPI+YiwoL1s4b/4lbhpBgh8zDd0zogyxO04HF6JeR86nwUuKp
fgwjj+S/5s673ZQmEiEajTqOuLVjyKp29iyU9tFLmYmn5vuaEC+a54EYHGvJpgRXbAG3WWyzncL4
5tsRk8rXbI9PGIRxhB9nAtcn4g7oPAjBdrWIG8gBG9J+9Lhx2ninu/FcQUwTkWsmqMON5s4hva3Y
Asa3GPF+K85hs9Y5agBMpriEOAeoP2hoZ94col47Zufy8Z/ZBE7Z2cn7gSn4+KZvZRY15fBVS8mD
I5t/kL9Xm3z2EBtmlx6ZstPSEogURkA/uCSFixWOtoEXozhSXexVakwz/GSx8Iijd7AT1oos/zLr
H41h8KoEANWtTTN+fs7cbFRJ8iyfQOlZkr09LelwG8Ne95WfHhQBLDajzM4B9GAaDR46edxf4XE1
V8Bpdo8vtzZqzDJ+8ol36MYt0OEHHtbNtY0S3ZXScGu+9VwyeFR7BAPG77yrwpmRhuZIoXLiHlO1
Nwv+4Fx37MzoI1WFIUgt1tFGCOewUNz2KYUMg0AAJggBw94+Ss6Ktw7jUVUJ8D1B76lrd9txBB1C
1Fp9Ec2KrmhLtJNq9QVMuOwd2SCUc2by2Ja7yzkW6mhKkuTFXeISl5r2dqyne3+jZc0Rfw5n/Jl6
sDXMCgW110ws8Z59OJFSmz2PYwjwrOXvMRt7mk88LQp/8eya0vdYonGvrtcydK8PiePBXbwKGTbN
mCx7+yEwygbanqwAsz+cq9l7X8zBedsqih8ZOOk8R4471ikX34ciAmJHYILwhNu8CXuTsjLo4wT7
qO95Hak1SdwkjtMnZtoACb2y9sPqTpuIHW6Z5JzRgm81MLpFn56yayrhMT7yO2vRA/FBeoDn3bXb
uWUwbmnoht1mRRODyZjFkbuAT6A+BA4B0x5O5cu54IrSpHjepEmV6tMK3BAuCVxldIlX9OzIayGo
hQ7EyaTTUGSu+d49NP2YH+xL9FAfzwMakW1AwXP/osGdPWsx8BcMUY4JEmLivkmXMM2aoLYLrIBR
QcjYauPYkO9K8Mt7IAZflCg7+7G2XMGy+HZ4n/mKWXNUwxdNpfJvZNWp9mEtGKX69CdtjELSSMMF
AjPsUJ5ryyao1thKWotGmHyWa5zYuK4GwDZJFbbE/v+GBJwSV/krYX7ETDhWw1B5r55UQt5fU7R5
njR8an8hX7I9rFeTva7sYuvyGAqfkeHHeslwt+6HWQ7SJribXgQw60GYAyyEOZuAiyn6ex0Iv6WV
NKDtG3CS3Ck7kRYZdMJOtSLcBwUr4sEjy6hYnjQ2vY3uOTcBy3fOQCJdDNeBz7pHxWiSiaa5z16c
YbtC3GVj2FrxgbObk3FQIRaDtsquZ3goPxHaEKYtWui1Ax7hkYFECYlLkT8r2zBLHS+DklPxPIAG
l5KGw2uzTCQFMp03s5GLyaiQXRkptUq8NcLsZDG4KaaXAvwCsaAyH+8qehJNGyJgEUPCDYRiOsfe
RcXDx6b9DSSYNBsVCS/HJ+Q7ZNFZKrcE23T2CnwYAbTBTNO1d4EUZOUiCvf7bZgldUgZamVlmHdT
Fi4vehfdVLR+meCoaPRWZcgHSnj5fi80fWRte1Dd5tfB++X1nmKOBE9H9JRcQW8fq8TaT0i31lN9
0Du45VeacEp7D+2SeBLxUppzliwuESbPoSJ1WlTz3NPbt6PZuXMCNr5xFMzhDLnN0Pb2+JodAxQq
Qwp2f9TsURXy+mSGzP4hbeCy86dBg+Oii+ltwJAKaAosow8NFzsMiC1T6BjwdIPyoaM0peu5k6cU
n47fiNhul55+VNRkuT/h+QjlLmbex7B8dn+YruQK24Z9A+b8Ft3xLI6s0Mg9rhhHQIkEhYezmqeW
LCtix4/zkKNQ7nq4pKwP0ipHBnsI1cNUvsQLa1RHnKLeiCW7anJeITwLqb9imQMp7mkzAkHaoQzE
FS4LKYA3PLVL7+gPqGBJoDDfo9CViDsPvn2v629o9YZjX/qUB4bmZTnNUSjVooC6WSVVTbBLVQrM
WDQjPLgW4kFmToC0n5QmcXUV6QPif+NzmkfjN2Q+Lg8gKthYSZTgYszv8qSWGgM5aLAmp+JA+Y76
ApnaU2J4WNuSiFax7rVm5X8LYpcKVn4E7faEj/Mek/9tsuiTC7ERCLhYySNK9n7VSEW5B1Sd13gY
7XoILtTP6RYL7oyPClA51mddb3h96g6yxUmZt0BSEL17NZLldmmUcrkUuMcDVEYBhnbf/vOn0TkX
n7AGyw/hvkvBoWFH5XODd277CT4dGZ8dUldE0wJbkbEgGHymdtuB4yYzqFJtIviVDQvkQFXp7hKD
zr3VRE9rDOEH48ouDDPDdquuEOKAe64MOFibUEXN5c1CsR20lXw/iu4uMpAU7+O4fLAEE/TSxx11
BqI+SLsp79vNTnmGSRBc/51Mhu6ozwxQ8Pfc0G6hvfqPN30s40IOw8QdI94Xko9bV9wiAKRVH8Fr
V36yBa6hPVbNtBSGmOUjy8k0icsb4cbj+vtJOk1qslcNZxGsf/wGQTdSteHazKYV0wdGBFcW1qVT
vMpjL8421A/WsYOWb7twNS2kyrokgGpY+YmKJ6mH9wwKm+38yIy1xbQSSXsIaTMs3rhUSKaw85YW
kKkk9qFiTwauJjzSa59n8TqI819wBjmEkZbOY3RUWeYr0vwCVogJ/BEMiWGg2iRavE+c1q2uRvQn
h6kWk7iYWqWBavlpOoEeIwt8O9MeOeJxI+jmwR3iO6lQD5g7qY7I6JyltynA55UcNLN3y0UVbFNO
+JMlifqVDmO58lBF6CHU9zpxyTidnpuMPWB60j3rtJIuIHi2uf+U4i5YjLgrVUa2/e24UQ6ht5Yi
gecetxB68TK7KQChRsPehtun/qHi3L+Xb+Poh7NaJq1ofAo9m4c1cOSQRdA10msYchlj+P7+5mRo
VXcjKgKYXduwopG24uLZdZzPrbypkmciCaruPIrIZw2bKJJCTd5LcSK30++r98uP2YgqrbJMMTnp
IOvywW8wT5n6xJ+896JKTuk91t8ESOz82EStIP5Rs2yfQFuANNTljmm4rR5Shm3re4dOyWwj2+bS
kjioaCP7pmVCZvv/xl7tCp1UBHYOBBNM7DFRMW0k3UDgxt8ES+/Y2qTfIiLP9rAQQDcQglEWo4Gz
x/DumeB7khFkTr9ABzja5m7rmCj8B+EfZ0Ku5/Ym+XcFITO3IXpVMl4JJs93CXtn0lQIL000Pl2h
aT4T5vjiXpokg/CJjrCeK3l3HJnOtXaaYT8eEJZ2VqmCzVKHQq87TdjpjAj5yzkrHg+GOUvozDY9
X7jWdbZKie8/dIpGJxv1185IWOK9d96XAre0h7XR7cXArNtjBfgSyfZ4EU4mXXMY9I2kUuldfclz
ECTZmhRym1oXEoSmgSmCp+fyw27pWnvLDieNOWsM9lt1xqMSCGLim6z44C2yiNfYdhSOZ+NLxoo6
pXpLYqFsbGoH/ilQGIT9HSDhnvSWl99aC2K3+M0nYLrxO/zUjfB9eCv2XcmS6so5rXh6otAAqoxG
PfXY28BhzZQLOQHRIQyqW6D4auB7KDyL0SpVzhsPQAd2yyA6m+pgkOABdZThox4K4R0sPNyz0Ovz
1Ys1rzG5kC5dkdVNB82wWX8AaPWn2l522LM/BLzmihtH9rWODSNrPeEyPVP8lFdeqTx1rJd3hJs9
gNzsSR4olPYF7RqbRgzhHTSrRr4NDHqaI2RI6PpsXFAIap2d8+OnqoDnPRIz9t89XE+rQxbGUqBH
8EM22rE7k+FTnNswXAwu+ZhC0X5KpsQZRO6H78sA0dk/EwspNDIJbudyKiB1Qy/UBOi2Lsb4Y9It
YaShmIZqFM92w8TAUHqrG6Iao4T6s/JK/2ibq7cd7aDr7bxVlTYYFem6LQqq5QAVG/V+FVGbLDxt
Gk6fz6msgKNR2Y9iWCKrJVAwpIJn8tdlUIL1KHQEGOue+CdF2XTVb5yDO9PEgeQ1XYwJ4XeDhXVS
bswpvBvarwB+cWVKtlziO8KjqM7sfbKzufQrs2L2viJbfwNyxmbdLEtBlV+ivl99ahOMwEAh5spi
ZTkG3pFckEug6gNrdmb2hzu07gyxvUPzBA19wLi/DxwoZFLGaPKj+HVHdHEzoqYOgL++HvH+w8gu
80dHa0CiUFNuGegb5ngynGjnrfuP6WZv1X4ez3ReWLnTNBX8cV1DhfQxI1KwRtp1Nm6HiqlRgzG3
jLj5viTPEk2l06cNeUzk31Iedl2EytscGEDhdfLdYtTKBMl84njVjUBXzzloxHNKusvhevdfz25K
Ios3xEa1ffWoswwrcv1OLNZi0NcthNPcsmvb/4VdQIGmLxKIFbTFEGqripj6k3VWFdv/O5E+P8Dm
8MUXh4PXnzXTn6k/lUu93GXLfjY6Rf+72/hXpfWN2S1H8cFaDBSLmgKiG06K4YuoPKN+lFBGH8Eq
iPQRqMmbJlNXGbtTdV7Ldr1MvgyM1dclZeLKlJhau0IegGKOH4PRmGRAD6DQaPxQTSnJz+tpy4Ep
Jf+L0w6FHhVjRgPDIbL60G8JTNP2MOTyJT2N8z/+g8JLF2/KeqdgWSZJYwVTYKlg+AUOZHjSOe9O
Jz/LrrEgZQpPzXqRSxBjECCTRHdhgLiMCyN/ozaIFlm00V6bJkb0H+hocOFdNVlX3gMYVovLLJiI
u0ZvSU/LHaok4h6NQO6ii4ytkODzXYWbZfE+0hlnwl8whCmmn2YPvTvQr9UvvIzeTh2T8S4/SRhZ
3x+8F0VP/2+Qozhu2yy6h43fGFtwttEFCoD8RW/8U9S/W47pXzSnAo1x2wVt3N0xuws6ip9GCA6P
Owki1MmwBh0duZlMG9hI5LJTowfGNRQ/H2c9tnSOxW8Xt11fxSF3qWaQmine25gN9rQSTqWf6tMb
AQxWbT/q/SHHyJ5dcWRvg66jQAYKxjsDzXLKp6zIQaqt0psizMms6T048SGmCWeLPgAKCabXsrp5
HIMRJSW6lCWfIkGjOKzwE0MC4PbvDtaEjZBUl4gXOGqBI0ONQZKlHE8u+vPuDBDsVgTTDGdZ35tB
w6ycOZOEiC+u5nC5/9LlsiQD5SHB2lNBuAXWSHRakHGmKNQRymBGo8wnYcaYTS4nEUQ7sV4s+pSW
LG4IZdkxp0KuDk7tScAjTAJqZtuf2eBtD8cHYs2uNL5N2jB/a26/+Oq9EuhERxnBYDSD+1DTec61
0+GybqblTidzA1M2kJ4X8RqRoKhxRVFSYWQjvLdIgE9v2ZnWmPNEu+LqXly61FxMUK4FMiK29XG+
r/RqL5TCQX0YEW/pWtRj/PPJFfAgFg+QvWUPcUkepg8v30ROw4Y/UH074rV0FcFsqS35j/lIk9O9
4dMntZX/wuBh3JsrMSpKRQsYyesz70Bkipmi24opcRg2xDD56K+4Ai+CIaJs96tV9Vq0jGCRPCtb
lLy3AoC5PN70gyUZ8TAGt3rqX7yBZlAcRWXeGiatREqb4TgwTZnXdEk9TodXEBLqC5q63mOXyV8e
X6n/RNyObzFGi1vflgzBplJWP+JUtBGGk/TLB4amG7PZqtAl2Hg+hIP77wbBYdlT4iULcca+CUHX
B++pygo9AcTK3BT98FMesIqSNilFL7zbAy0LsASAGwSBfezb9qRN2fdbmR7CcAWAEW0S+s8Bjbdy
ynrf0vHa8UVHFkW5nE7RZCH4zlMZPA4KLAeMuG752rx4WnrKw8xt4Mna9o+/PYPsAp6gKLqu/uPP
IpGEkyTo1xcuwCQZYiyJeyhKyPxSXux0qUtpR4wIKap+SFw395R3Ys0J7lToe32HXrm0ZUEopGia
shP2H5bWQU1/wZn5o83/mt5hkS2kuJgqVmXWcGk6naevYxE5Xdc/Av0bxu3f2ZOkeVuPsuTSRfkF
EYqgAFnYvk0X4wD8ZhKUXhZrlCQmixoRrRWFBtiMTyAdpP3f+oYmrfLOTy4jDSJuWLABWoUaLc7o
0cI72ERX29Xz9+QDZa7RnRq5zN6JYXCf9Kiy+YY/YoPNdENOm94c+kCT77Fi2+C779SgMKJbhw6q
IvncMHkcn2r+wENUC6bGcTFCqy7WaiPos10ZbsK5+4ycYw6BFG8QbKPnZXcfknufV0gT2uSQ0Yvx
bLO6FcjQflUwJf35xxxuYdsK+XpwKqI5zKC3vFAdZjQRiNRMMUyCyiu2xJ+b+FyBUK5ZkcL+b27y
rMoV4dV4q21IPtwijdkbF3tDwUjzd0TV0zAHwfkBtnU1KauwNpk1HjGpsIJrabJ8rTAhMcUlmC/S
2eRYNZY9iIinLKl0SOAq+pEKvPaBl0GQGM3GTySksU4AVznwm4NjFUel34HOEyF5QP2tI3hBgg9J
3IHF1Z3RQzk6Mm5kaSCyqVXXSfYE/7/pggUyml1AhLc9uRCXtI6NXhxc9PkkgX+kDOsGvNTDe1hy
PGogxgwVK1WS1hcJBGadDkgFgt9TCxw/5cprjPGau10nmIDowm8lkJfojxYtq75Hge++5szABzbS
R+5PlLvvcB6jypyV/K2gH9pKRwyjUnPN+AfijGCSzudTZzBNqsf9F3mDaAhgWI4awxbiao9x4Yrx
TV0XUgSjPPrXBseyXp+ZHrK8y3iDg0OoayCFf7GonNb4kyXtOL+EAtgHM54IQqhCKa4Hc4IbzhU1
5YIY9oUHwg3cBWYqzao6iI1nnkKwMxjmS3IgZ7Lm9NRM5Wxxq46r14VUjmdnlat74e0cRRrriXPD
v1haFAgKqnxdjLZk6SMiw7rU5t8sDffKs+/rVgVuG3/nJKtFb1C2MZU1p0kmC7RI8M9ldZaSjUBC
hUWljWLRKG3jrRky0oea65hcuKuiyNrPojKQJb/pUyIRmKaDzCFyMcO0ZPH62b7T58HRJRF3SGnd
N382PEuNjkLHdh2qO9HQOOnvWdKSk9hkYgg+rHD9mZgalpU+MjpwfRqddr1uWrP/lD2sHAy3l/4E
KVJSCZyA9wwm9UTyc795WhoissAUSHZaJarNIIX8iFNBvRJBWeZXl5w5Avv8snj5p0qEp7GVtZFw
ZwCwIs2ZvAfURcbTh1jF9q3neeg5AKwF3ZmwlHIeLpUYgsrmcSL/fiSmqpAQ9tcPBMfCrlNzOO7S
D/hep6wisvcLHCvhH9nMJ2FpUSLTGNdp+UMZoKGkjUfPTS0ZbQckiAVBp+jOaIQqLxvO7aGFIlfe
/CNa49IW0FsnoV1856TE6NDZ57q4/YaX68o4F23X9kV/jWGH8vj4BIfNecdNjkG18eHwvhRkNGbf
GSjsOvKyJIZE3t4EQlNiN3oF08DmH0OII3UXa6Ti9gptduiD7inQx7N6l2bd3oToDEwPomXIyCz+
DrzVA4H3aeyCa/wpdu58yLiOztk7CFtBZ5aPjfjNj9C43oBk/qb6U966oNu4NRa0697ecxjDLBcc
7T7sd59kA1RS1my8lpiZyVoYh2cG/ZujEWZIgbOEi+TfikBaGRDxjrEU/JksrDajPtdgnlKG6s1S
Pg/eh3wxyhnkZ31wX1u+29JnXKpB6ZZo47MI1wrKtFRFbNhpZj1AMH4MHR0Vv1vTCIr0aAsp0LGi
TBWaTIDp8CO89Xq6DtRmQCs51I6BRcy53T2u/GmakW/WfpulMZ1fUGbyldHHPecYH0mpjMrJRSt6
M2gLTEnS6qLSc/UkXQfLmA4stPcq6yG423A4cNPjoJcYFP/rKS9b601IhayttA7OZyAQghxWTtaX
cGut6NFbp7cTaCmsgD6xSZcx1Olpv8m89Um5eIfXSvFALOhotbeFY6+qce6UAv5fmD90yGWwhXKB
lH3w5pXGi4/LhzRUcWaQjr8cKKawRHjuSrNRR73YzRuDN3WXqUiUI50SVS9TRzS7H+06uh9H6a9H
OJLLzfYhpzUK87dSP+Igwde/R2DZEJLKnmS/vikirn+4t9e4A8MXrELEZaGZAR040hPKTzAYuge9
GyBccmxAHifBu335fCdYFofBpc6WmLTOBh7kB+8aJfcBYQUV/jEc6Rg0FY+Xy9PJRD76htU43+n3
QFgm2Th+KseUV+rKKt/ljyW3WaZu9wH95THV93Hh//xAjKG3jpJxaNChwpLEn8TvMG81HpaaZ5SP
phd4ajiITD5ZfX61q7MbGL5XeeFmlSg0WIkrPWev2dIu0MR/aP+9ZSqY0SlXvZzjHsjbwEDktzgV
C8hkCrmWii3/qCVAcI3oH/DyUOMcXY9gb7AlWlnXOx7FuyklAGD7vug1vAH+bEu+hxzyWv5sj4qi
iPjiW2PnfT6tkdYtimEWT1rlDEUEOWBBW4EWVR4eIwBQlY8GVUH2nf2tvgjOCQ18fTQCFM9SxZRT
RzYPRoyjbY3ZD0d6dPNe4vA2+upYkOhiDejY6FXKcviWw7vV3mJis3FK77hVrmgpCHhfAZKrYb65
PITRRavGyketslodAIOcOlgmoWl0kjJ0npPUF4iTB7ztUhEy9EqkHMkdiUAB7xCfNx+df+cKczmr
1JYcHQRAmufNm3xmSE1+UMhjna7idK058V3WW8fMlv3wnIFK+2Fi1LXwtV73ivDfS+wa5uVSSnPp
DZ3N+VSnajZODJ45yh8AlRoeydsKn99TcsyctkTRkyikc/8263VTeQxHSAY3HGMIB7SJYU8i5LaO
wyjedqKD0lXG5oOGiuwX4WiRs9l4MJk+BIfYIgIueQN27gTQ0zdNMIU8OM0AEIzU5cPRgcugAo93
S/8WmCOG8ZoqmGcJEGkuYEoiF6h/o1oYM639b7fyXUZo1yk3D9yhijL6vxmgfnR1h8gkYmInkIe7
Q8pHmH7ft5dFXlWmt+e/MN2BhynNPYh8UG7ui1ZEO4vaFzggHCjxUvvR/uP+8duz4Fyp46RRKBOW
61X9Ny0y4PcU0nDTy6Ak0rZ8aF+IK+K+vbbSfABvVd2tXQSyo4reaLVAtkkDLnxZQH3sJYTZUoNk
0K3RPKOni6r2MxWR0RGqnQ+OzUnFxnxxaSqi3iHjYmbYdL8xaQhL8djdN+Pvgd7oePJHn+BGf+pd
vfe9sYacPp/FhKz/GL+RE5UlPmgiduCMBxuxhtHxlWjN6wpuAjD9W+A2HpWwoaTZnagoQDmki3Ob
m/x42JVGKvFyljSB0ZmtQ9xDaJ//h/EHRhRHSRymrLP2Ak5kwYg6A4jjFJeY0Y8EISc0jB/dzj81
D+NhlA6qIyzO8+5MAevsAPm8iFrJglqLpIIHFz0mOwfkBNRA5Ip4mQBKax5DruJvUwBmflLS77uE
iyw+k8rGLGEGfAB6+P0akYiYBssQBhMswtposW68WQKa0T4GpsJF89WB+6WZnB50sQDWrh4w5Jp8
OqdXkdoX9EyOaRNejNb/h//0WyeoYLk/L5wvjw/y8o1RzeRslpWoPJlpigdAW7YY59QOfutC9u1m
oa0LBYaWfaYdQQYx8nCa6iw5Dl9xFCXBHKw60/YMUyQs9kAy/1ImBJm13fz9F+Su5kt3PIkcvVaa
Hbkxr7F2dGSQBfkTQIlu0t9CEyjtVZrf9oXk5pQm48Vutq1b0YZq8A5jPOR7QrUpXEMlgTXCjFlQ
Y5H1OwLWTacRkhmq9mjDENN27Dty3ClnnD5y4vpzGKq3gd3hpWihx/KV7ZGZCBXKkUA7shrF5Ze1
iAE6NZzFVWOSXi2+QSBCqBspopeXJPKLz9yxu17p0mKQuOcxeEoXvGzFTmHltrcTtEYwTXqH7GxM
uM551RFPL2Upc9oNgYqiTV9AH4PoNtmB5WnpgxAa+jb4gUlbzrhB5gp2XdUr4myfEeMKXPqFw7Eg
oE+yujKaVRxhXWfQ6QcGMssX1oZ6O36dO1b5SR9h5QeV7lmJjciUC1eUI5XraLuhuhd+rY/Pv9z7
duZ3AdyJScH+Y5TMwZBO3WRMhfMARvDAWGdozmGNoxKVQYT5j/QWCJpGhCKIpRSHLPxpVOTTGroQ
RjPIPUG/EAH4Sra+SSM392AUYY84OEFW4AHMCQf4n9VwW2WBbS3lMzPXqMWlMYlpEWsOJu7Kfpd8
llaqJCnPfK8Ee31seRybDpgh3S/3uulM+DqFVvo0g35EHyKxUuEDJY7pQ7SQmueGSGg2vXwXjWvx
z23xZ9Q5A4FriDf3uchfRawqZBAWxIYyq4asQseQKqjrbzXb+gUTd3n7pWhnS8yfz2Ewe6bkuImu
jUAZVNk+c1A5BdeAYKRr1/QxqLiNCChRlYzfH7Bv2oo+VmilTPqSd/+v8dMswyNmeeO1ZvyNEMw4
6GHUhScXDCpG+W6e1GfGSCV6cQnyVO+BOuuQf7TSUIiyHXl/YxrujVBcpVE/MjF222v4yiDCTLKM
OCVku4sGaRS+9Dmo8AKpAukzmnq97tCpcGSq1UWm7e/z4pyvfEbVRS+BhnC4qHkPCQ6/0gvlRTG7
EVtrodcCgXUXReSfUx41J/ra4reYoO+rkzae8XS6UV2oOeY4oPwwl0MYU8pKXrnpQlT72Rpj8YmZ
kfnMqUsUSAZ3j3YcWDmyBmxRdQNgUaT1FIDbv730ia/5io+4uusL4fCVd64+44Lm2+UgF+33Ac4G
O3zV3uh/SVRvzgIW9N3OyJLCgFITfExQyRPyluFEKRJ4rDqxJ7bVNf0r7TM2sKbPBco3J9czn2BY
WDVDxkO7kpzkdatlG2OuJRm1sPxYzL8MgoH5qkgkw8sEYgoFUGhSCw1lqIkBFlfbZaaHwHz5oi7k
pvLf8CLhcIHGeFfXzT7GudALTJU4hyIfqIIirRgxms4GzrfvWU6KT5WCcIhAENGGUf4558c8V8fi
NK+wYZ84K6bQK2J54PGOACeOhan3WSSidLPq9SRdyVx97PBWloouvOedWqN3eNghNtthJ2NfWDRC
+zCDCIWHSQ4e8L0zwPx8rgSVyVjHLOnLg7eJehrw0i+47hgcEtNuP4RHxtlFHYJes5FX089Tyr0X
G1sJR5hhznLY+ail4bBcSXUHDIk5yPEVlhMwgZtLLuCkVgBwzUXyVI0ok+NCg5hHYjZuLJTefj98
G56oFvkalJlM/STJT3rdATL9yx5TfWcpyLR4fYH0orq4FkuTDqWi5CKEoiy0dJ1jZe6SIK/VakX9
ckHLPqMLjv5QtQSNJZ/H7pytkmUDqyc0px6V6lfdPSfCY8VMYTkeCvsKp7uStevAlL6TG7AMZMa3
QlWIou86gY2S3TJcYE86SXc2SGwr323B8ppxwot1xIxRCnkuqdHH2ez1t0/1F7Xoo9grJ2B+o8m2
4h/OEkwqyMyr23Wcmk6CrqrBBkNfURdM2nYhKpby9BkdNhZpfp675m6AF5H8X+ySG6brxYKIrP2b
3j9qD6HrlSeTHQuH4rthlf7BSm8UoNLrEQHX2XJExL66pqmTo7K0DGLrycQOE23ZcDCBRRg0Dd/T
gUWiY4dQGKiyLqPEyy66FnBmkcqBfztZ/9UIpAs4TnmnnyvrOImDDvPmK4mwZMh/efH4neMLHTpT
2HV0loNxk52n8719uVNxDj8mRvzyX+dX3rjvwQu/xe8k3pAVkpaSP6VdxP64Umz+zm26eFe/omaW
qeFaUH+PLgPAmZLvjJiK5YCmLwyTaj+D1WWGNCYZSnLyc3R9Xm33Lnt8DzwScUFd9PLXWwIDJ7fx
ef9X015bFUIxtDJU7Y8jpuSxRaGyXQRihTnqtkJ8xse6H8KuSnrjksJ0QwiNKrCGGbOu7luCRSt6
fQwBJXj3Gi41WYdAOnbPCxK7gdJl9VAWvFhKwmPDOkHBwy0JRB/0/0q7NKA/ZtQd6w741ZQBnzRU
g5ZD/bwOvEcRH3EwvPJxqIWcgsKa5qw6/lNKF54IAxp5Jfr4CYKa95v9Qxeh6XYSNSscuuuzItXV
AQFHrKwIJfDIak2DQxJyRxjQR0c8nx0a9my3kn8e9+wmhedAph5w+Kl81+UYdKdfgE3SWYxhz/Eg
MS/tTxstbFKXuxvyKD5HEObdOcm0UMpK9m3M9464YwyE3dS0n7WC9goQYF6bFcXZ0/Kjle5yvDS9
gDREOzoeELjkAYoEBBuwnY4A4NLfsV7U+09ehPc7jGwe16m8iWGUw/Hn4KYXR0h22qlMQQdDSouR
Bz8dJL5Gb70PKHh+wfAqHTLmjZiqLXSnoVkjhm6gyiEYYlR+q5rYM74hdJ2G7/ufp/G6B9JVwDOR
jdI7r+areWS3LUn2GVdeD44TmPdiUeYQlqLIa7poiOUjy3dKNLg39gjR04g41mL9yCSjbFkIX0eC
3kmIitOyEuO1RjJDIwg0KJjaraRMYRBHLSway6s0ekALgPgkiFbW8qjDX4C29O/UN7cwnSSofJZH
bU6cooYLLkH/clzMhPBacWxwjZHsm8/XomtOY1xJHqoX5mwBA7CdT2reTG19KQPyq+tW5uVTFpVp
hNI28o+NZhlstA9pW0JQlkaAdJgZM9m4VDqGqbZc53Zw5QH37sLyT8fu8GFmNSvHvefWgiRR8fpM
4GqHM6H88h+KMReOZT98voqujKpW+6pNA+HkgurFhj9a4hGhJ1ltaWBPAHmBJ5QFR0fVmluDkXhk
U/Cx7GjHtIqWzXegDcD58K1vukJfjaws0w2hiaf9QLZ6iqcnQ51ysNT1MN2F0q0W11DQ2MIvvI8d
TvNlTcvAVwzBwEa8o9RuJSP3kjL0pNCooDAUMC2oT4eBlDakICPKlC/+WU6bO2M6bYs1L00QdVhI
QPB7+Q+r2ZyIILz5Lys5c8xR1GdWC3ozasB6GdZTKyOcZIeatgRyovw+rfjA2w9sTU9Ws/Px+170
au922sFM7Q0N8+L12HSKrBvZnj+AraEL6YA0nCAisDMD0wJw8IWysp0w0jWIt+c8zy09RYkrPZyZ
0veSEjXv0KPK7FKHPHHI0I5x+XDgRLaiIQhBN+aRGOx5qk2mg79RTdqMbhbj1AX/HBwJVH4T/C4s
kTb7Vt7VlbBPzOLVQlwy38P3tEjyR0n0WKGMoVhnPykFM3GbZcYEL986yBYMSMkDZJUvWW7opmPz
bQHrwUci2VTq2mSJIfMlYVIaaeZBLi788lfJVXJ4+1/7JBlKj7eFxshjXNCpgHn/K0KRekj1E8h5
ZgoJPT4zBUaoWOSNGLd9KPH3FUp9NN9DTbaf5RlMbRkSf97rePm1Ues3C+GEkCgmbGXO60MplzVJ
/maCPTBQhKIRbNr/q4HEqNpgMD7HpSrWydAsV8tTx0tcXhMJhz8dUUbZ38a696HVaddhQoveJ0bm
syAl4SfYxz2CUaUvaiBkK/cbB5qNz0MpCSqMz8Ul+e7pPXCHSbRrWawylyBZgM0Z5ldsgub41Pmn
0YCfmtXqioIzVLw/tNd/NRGWfvLmqdLuGwaVkCOSMTz87Ek3454bxkbi+Io8JMxEyIdXfh1cSSmF
/FE5b674pMgrcP67F0tTSWNPQIgsP8GvgXyUAebISdlKTbWkuFpG0zp2NPBbmo0cFe1CVewOlqG2
gwLkhKxg9TgWPOXQe7hRCFqo85mIGNmMawomOoSpfSQjrM9JD5F21Mz5uuzC62yD16hDqpcbW7lH
6V1ziRzIWfB/CLRgO6A6A/cD8Asey7RuX+me8zy0HfSjgz1UXTzLCczGf/nyG+QT4P/yQ+pVWuo1
2jhqP8ad8X65DurY4YbuexIF5qNbmbFw54I3GZSmNqZBa/lyWD8RoUfS8BR0AWbfAyPJEl6Jj0vA
8kIKAP2Ha0D4odUUHPghyfma8JGdRhsycvgtgndwYJsFsNcMoPY/1v5s2BTBnIjwFEW976cnoHpQ
ja2tkc7hXMbRk5wlVqA5SLGnF8FL3HU+DCtQ0mGTRJF5aHU7lq1O9yChN3NEjh2y/n/QHNgMaORk
6yJgdDPIbyVm/ry0sRL5t2es06o6ruzOya7iXi2wgojsVmlvL01jneFjAWnfdChcY6wu0oiBoIPz
qBQT1YnMGwgomKRGJOSV3KRS7yxNARG2LAT6VukRD3wL6HCyqJ7J4Q45DkVQXEp+jzIvPFmlJbqV
Pwopom8Zjmy3bPBxOj8qqvZqkYRXIm28NsQi1GjUnkfV5ZslB/KLbJ8Utv+jiAMhZNRZCwhraCNL
RD5vWdO8k1BsgLgYrz8gg7GlJ37Rg2erZ0ZTISxPQa0bqKUp0GqJo0nk2nh3z9VWvQjC+sE6o+6Q
7Hw+9ia5xCQ4i0tbi/nLJSUdwJ4hBgkKeZz2B/cpj8NxCfaOB7nfhhfBLS35nPUGWB6sN840IiKs
OhBZYBAA7fLRaAO8s+eGyDUkSAu3cGr9zDseL6DF8aiY/tROE4y3t7qU64NwB7m0qWPUjEKv8K16
RRvmuTFyHwRiH4ArKQROOk91/YcOZhiokHYEf6kWseGFbcuLahBZSC2uBPdM3luTvp88/yBIEN/F
AWatmhpSXzH/Ha4QZEwVCgAqn2P9/gwyEFaRGzQB8pI+q1HZ8mAIGoPd3ABQ0O9zlNktSo8Lz6qK
m9hi9/HkTDqaxXN8tdnjUgoiYiYWQ5A7+njWqQqgbxgOz82/OJ8EtjC0wbmIt5V+psjrSuvpdwaC
vFVus1t2jUiye3EwK6uUJfqI50WqbEddhSo11pXr/u4fxouc4NBNqGFwnv5zg+ytuBGMMUQZveo9
mnLJZ8uE9lQ2mYTvQ49+vcMZdIGwVMhxgQbIYRnA+CexxISSViwKwl0yzwfpIqEvKkxoiXosjUxQ
S2p4uCqUTHnUGQ6fJ5W0d1YIoMZiWytS/f5dWer9UJ5CP2r7jcQ7vxdOo1kK1W4BtvcW5YUc7lYL
F6GLerFyZ3dbv6ftqVTbcwmn2TOGqo4flNmePoGStbIsoIS4hrWllRBjd7Z9NRxbCpvdp+s24i6o
iQMNW2xwcR8Ote+l+/9zuGiRGmpe0u1vydDfdh1WiCs6Yg8IihhOmTiR+ST1K3hlKWviJSqn/ecV
YCe2LeWaAjGQZs+77U+hjAZhjXRwK+Ig4kxiUNdsbRbShEsD3wJ8Te1b99Vd/3m4zCNDWI9ebRjk
pvtPZFkk27t6DN0uSBEe2JyqaHpyHflJFUd0GoKj3jCZo3ClO/dEH3WG08z/fXGAp3jvZ7g7CxOL
05PumH7Eo+b+xFLtN7JjARdbP6+tLsjsiTHRpzGj9lRQugpm7P5dfGZNWPci/czx9I5y+ch/4OQ/
pFvL5QzuPXXJrNT/oFoSCFXcVBmKd3MEdXd6fbNpFjfE17SLdEIijaeKnxqO3Ui1mQ8DMLmgVxHe
blISlzIJttXL6eeTmM9jJbmgDTLLUWe800jxRXfb93cskekgyf6P03rWIUaHnOjA5Cie0Zp0/uoY
+w1Q1P4VbyvEFaGfCUfDX9pDuXkrFD3+5APA9CrcvtYh3H9CKuCi5ojf5kmyskkn6UrAlvKO2x/o
FI0joMJlLwaD6acmPRyLujs/NtrIkiJRJA9ymKq5vxI30NOLbvd1mfCXwm+By3Xs0MY2CC1VCuw4
L9XFOeoekapzAp9Ryomj2dpojFFu/wjhdc22DWC3RrbMKx69SB6URKGJVJ5sr0okh5X1aOABAa9G
3r4qMx7euU3UcOsKh0DpVNYu+zr2x/+VsLTgneBHJr+BdU3KsYJ6oj1d7eOx8yGJbe9PeixsRDZP
e+6PC6atmsLiZRxvJeK756qqxbifZuz/pW9EaTiH8wUBUBFhBDnvIdhbjtBxjCA8tkTVmtmZDrKH
eXfXimvhmiRZyLrX6n153EumVUIgZsW64AiHTGb8hb91bCoDFRvqsrgjsJ+8dtDB7/75gE5BLI7a
1JMYFer5qvA2eeNHNvArXOJBl5ZBGSwEUZia7LPZ9P58s843kzZj66zeK5zcYgkZSg0vhvmtIFYs
13uyqWLrP31DbDvWnPMNquT4KhbXpCdPVoVGxpiY6sZYPLA2tPDDiy6FvvfRGLMGn9STvdVKJ5DY
8awtqxfnn0r+hshUX45iQy4o47cJ+wcLQrAls8HdsgjFgdrtLh5VGj0vh8UZY1+WwYn/jfGWGq2u
6Loo6pDKqn3ZLHyWAVAMSr2KZfY2FuucMqWhQINuoNX16+Nhb6cjAucFpNyNlUeoe3SA2yYEKyga
hWE4hHXpwIqQaJyH6DxUh99LgPB8rfASZaWYmT8vRLZDuyscsgqgw3edqgOdNtwWvp4DC9jejD3g
eW3zLHuCvn4hR/GYtQCNH4PlGC8v691xuOXG8/MK4uW9kqE9oPJuUqSJoUIje30PgRj5za8Fo9aA
eJaHg77C8sufUhacZ45Hzpj4t/1mgadluvawOoiKy4SAVK/QaCEIvyzLrCUD8egESVGEZWDcRIBc
IMxdTVTw5KASI60Fft3RYcA2MzKS5xqdL/b442H3IwP0JvXAp3MQ7m722qYn8zhhJs/EwAOZReet
0FNU7TkCJHEd0rvXFSL5jJda5h0wH6bMWLxglu3sNbqo232GxAIAkW9cvP5+ay+K/1hl2Md3F8sH
/8Q7dpTXBzIe5y0vuZFAXowqE6+SZEcFNFw8YhR27vNiSvhimoJUzdf6uTCp5SR1v3rRkfdFePVE
BlBsFEc7UoY4Df1jHH6gOgP/FXJlIr5TVw1brwY6fGOfKk7OjsfyNUDsKcnJLV9RoTSowi6vHzSn
1X3zWsJJMqehqKVGdQPJjgH6ovH559MY0wuWW2BLYVGc6HOgjQMdLD9Jt+SAXai1Fw8MKlRJkyUL
+SmJK9HWgW9zXEnk2mEQJU7BM0MjCWMTw8ADtMLlShS9JnbSrk7drkJ7QNoEHn4u8L6R9bOSmazi
VHaMOnd22w/k+UYnMCj11YFB0Wue/zL+ZwKP1Ae3sEvqbnRL9epjzQKP3WcPxqAACOgc65wwyjnK
Gh6sWOnax3U2KkcQEqo/3ZxOmD3RHhQnikvvbHIUgKqKQZcqnrC0K5NtenUdubWLb59fl6IYMbKF
KCg+iw99nvjsy5u20cfacki7lhfobC7KFntMrY68BgE0Ui09NUaymDBK0P9sSR9P4BmKWLcLxqln
UHxl+nnin3SsojzJYv2/lkgwj5MDL4NKSr2UYIVu7KrBFh7yrA28aNaW06KvqJ0b1vvIpzewENum
05Hpo14anZnn2PpEmVCmI9WJ3T4LAiJ0mrR/rjobRZoZF/Idtz2qGJVfjDL7nNVYPc8wYZFCvycm
ciCwI2Jo5qhWuPS960mxKzThnX1GfAMjQR548uKC2ELadBwRAmiG6FrZdV/m88ETDv+3tmwN2exf
7+m8oMvDMtDxEtY4ZJEFYWRN+8WN5LzQZuKYR6jFZzZZl6CnG3tILa7YlosiWa2ztCBgX+AhpYxz
08ZCOAY9nTZOhdlCOITm1+hz/qafw8++8tmCBkp4tepxSrBbcfHhqknOA+1RrNwmFyqgEibWF6AG
4s9jRbIJsKps1TrwRn3JA/Qxp+UTt9cIpBrwqAq32Rw7Id/IKHYo5d2LsgKGq3lND0cR5MWs+/Ro
fn6Kq+iNofNhycHUq4hCF2uyJ59RZ1S97HmGTKttYS9+CQxyPXwaOlIPlEA9b19j+F89tozEFOdV
py9cBn2tQyATh+rg7fXCgKsljch+dL94fuyJHxVS1sA3QUJ3f3OyIQVbHkAnmpY3DlJhnC8VgQMD
z4zmQOvXANh0D8Bm49Wn2EDljZgYr0jiGXbcjgDHAYwEj4NQz2yhN7ZZe74pYZVXmWTgUDKTnttQ
UeOSF+x4GdvmOxfrLIOxmgUIesadstaSCvKOVHs3c3A5eVsEVD1S/kicV7Bp26iabFTBNOM1NmiL
UODoooqd/vBwi0epa5vBqFjqxSUn8ogNYTsd790kqpUpVvcZC6AmbDeql9nbDuFEiDbRL+K1mLwz
DfjZDOdMA72FcdNSwtfLvw==
`protect end_protected
