-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Ae1N+btiwY1VrY31mgYyO+8rHcdTRS70C5VRzTOlHgSnP177yLfw9y07DnZgjWJlQm3TOGX+Ag5Q
bQkz8/k82MuoVNHgbgvFfzxnj3c33F95vI2AHa53Q57wGWFnvY84jrdyM77HtKOPKcgiZwWD5r/X
hGvbnQ6yh9nUFVpCr+K7qHamgbUlH43OMSKNCfmforNfuE/4eDhl0a4lJWGGSqmGu37iQB332XTA
KncSVY2f4+dGBya973Mo/tV3tFH+gx8K49CQLJ0hAo31pCVK6oEI38jUTSRahupIsAiR/jjwwjlP
o85iRfE2rxEWFVk2nGP4YGABZbJ2ZlXcshez8A==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6256)
`protect data_block
sp3fa73zl7qX058OTPFPwUSR8/5a8EAR0n/8k8bkoPYl0vO4vbsulQklTmji8Omn7QToSlcGycb+
b1s6My24vXuL/0KzyctgLijLoINhrzM/rsEu2TzCxMs05N27WnDy5H1EB0DjHyHViIQfn8f9rkdZ
at7fDhtcAhAxa7EfS53WDwRbRR7GtyF4cZJMQ7P2C85vK8OLY6g61uY1uqSWX/JKqvVPQqDk5LNh
vvASvgR+Ol9ES59SymkHqYYrcIQIW59+KBQ+agmUjTRZuX+Jl5aojkG8igOXNNklCUM9YtWSS4ER
QrYmheDwMlJaF7U23KZhFHOgoW85VYMOxL8Pr/rFQRsqShfKolzpi9h9gbzJ5qolcPvu4gAM3wz0
c09ozw31VQE+ETuABAfvE82Gtet5GP76R4CnQbM54t7aXGXeh9VPg0lyk01qAJ+DolCDW+0M1Kjp
isVBHn47sZFZMKBqxr///DX5cjAj4Eje2V8gjaxIcSUyNBInGzGlgm6DnYLcRdkeV4yoNXcZamP3
MzCmKYogazLA0vqFyhkuexUSkGXNtc/98MmoCIeBGDR/gqIWtJf7NuXXC1ZEuAjCS6sDIR8ft/4d
XNsggLIsV8ox37Q/u2d2BYevwPzPM9KytGu6xAR5nuAfiI2zKRZ5c3trP4URJUoOPsBPrcSVrD/8
OBXrYHa5n712di/ubPikU89FVDIkNOiI6kCogXFr7oLBuPGZGVfi8JjuvH5XIdt23mcCtGV5puWX
c5gf0j35bN8wSce+cur6Azo56wdvjUY+DNBx9fzL2yc5wkgkRivWgJzh+ZJwhffoKgZd5ht1hJIT
+l/nKI04WTFgaE3F5bzrD3YigghvFfOHBDVQevcBPLXrQXePJhpWnCwXpZuJ6uOuI8saoywQ0h3c
Aj00FRQcD6pfYzQJrIh6xFkFNgaFpZovsUdip1X4FssG4xVxFV68gVVBQiodqX/+ict9N7DZCBsT
qSAObSMfTuv6vgeA4whHgcZx++zJyN8DBQIPwluxGBnI170IVQf0Cjy42p8xR8+Vn619AdRGRcjj
XG+x7du9HtQURr3kgatv0gnz782BvqeoH0mUe8JnZqI9kYrzcDZyj7lZ2kxP/bWF1CwIrT4iqmed
RsinUn7vwcpPe++9GGf9MFTwtY2nHY2DlAYprpNvDaMe1cqYk4Cj2QPAxLm3R8EpqmhxrXfH3Zki
LVknhPdK2Pr+omTjxdHIG/nUhMOHbSDpQ/7l2lhAtQr/g8dI7GXcQpUWyD9c7H2p+ApafwypUfTD
2D/ZTq2dGpVRdD4e7VKHPia6OdexFQXp4QrMJz0Rp4ybL+tu4zo6s+Sie2rqblKofSLwYV0MmkQm
5BtEobMJMkVFIi3vC+MQTaF2YR9J5C9cjCh1S7oBt/HgFKO6/xAcHMtx80L5pJYJs8V7z8Cv5fxn
iuryh6pFvN/+OR4D5wbdenFsT/MSdeX11kVfxN+OH5TcuRBHWBLOXTqm4T3xxajyjH6n8riApWaK
FHGMVKtcoTOSMNc7LdB605VK0foMC3pqiolHpwrh/dNBkHfvHhrYYRft9qNpzpWlmZo1KPAt9jhI
uFiwRt2LiFslH9CAo5onlep7WmAvgtW8j/33qKwl6e5Thn11k2Fw78jl1/tNeSMYeaFpaSgdinfx
FzWhBXRxRhxBCDzbVUPtDhNapfkBpFPmyo6zJnYCDHLzkQSW4hhJExS9G+oyU+e5epqh+u5lT2Td
dokR3YrceHrT/Yu5m2adVjEEh4m0F5QP3tI3kZNm+fLr37h6E458lBdquqduOLHyir4AAeBYyzit
EHGDE0JnV8GudYGmyxSn/4DJ37Z9u/kFR6hMhvx9K2mnmN7nBQX30vHcIaZ/ZDg1q/oHPxDcc+NW
B6v1BG3SADtAf9StqKMRc5y8Th2YS4v32iEYDR5uRX185N4b8oceePSujERUUF06kgC5UJpyOV8Z
vaKodTNdsVRu63sBVWhV4CB4089VP68YGwAU7i5Xje7i+/rhXAeQ4tYvvEeGTxrHZNatQnNaGy1L
Q5QnRokZIEx3sC2DijX4fqo3iJdDr7HZOHAvgKlU0quyS3zBgoq5K9s1S/1+7ZLZuZTTJXBqX7B8
tpuY9tna0st2IuMR7lDd1TC73yat9ohtmPpcJ0roFNY65lj+UsN8F0aFXUxuks+y5hmRPAnjQ7Is
ysVmy3b/XntsGiNMT8jACYfhflaxVe9SsaILQx6gpkbfpuj1Zez6gCgLmCFnUgYlIivrqW+8KQek
nuHz/UA87y7tt7aQF5tuHXvZ8HTV4pfNezELsilHH054nTWj7ZW/LLDQHKI5YtR4Bdmoutq3n8zh
DuBH1JP/xA7CQRo/nk59GjhQDf8izWHtMa4krBUpNXviuaGnQbX8yOt+GEe+7e5Z2vnEao/xbyP2
YVct3YlhM8wb1hFL3KLL7cXdn9jsUBjhOberIvGQCnxRHqJ0IqRY6OHBgZDa7vUuL2aLan5UcBL6
ICqzdSPfYspL1ZBts8gEV7omtP/J6do1EsvV0RVu+m2qFAyv9w/9mUI41stQ+hnH1gIzAS+YO9qP
1mMciELRA6EgFIw/1KcY93oor5JQzfnMb0LhIQg3eN9a+ynGilKfdf4mvQASzu9sbspPp49l5I0W
j42nB9xsMWM3tWvlh/gKbek9oK7VtnAgeLbN6/z22vvhJVtuOzNTVEhzqvTRcYVNhUD7ryuSfTIl
jGKSAzXf+5eJN9AzACWJxHBeKb/Gzoo2QNywX5Gfgm4226ZaS+WiP4hpX9oLKSjDpoT4cRbc8gxM
9eKOj2cSOca8zDZwMXN1fyMSkVcqkBWMoLwVvLBXMv9ma0tfC9dn/xeH0aj1MvmLv06G+UR7fLe1
Ab4hdIBljNJMoNQO8a98UqkvX+rrE3PSWSii0BKoVH5zDcA8fQjfex5xMJeogF/m+OHRtmEgkbZI
fs5zFa8NZLLgLHP3Ei2dv7x3hY1Ov2vastpgdZEmXsQ7o1uiLrxBfbG6NCJwrJEuzkPo5L0iWs9b
Hra3dRVrsSIx67IwsKc+f/viJarQEiq2T0W61DFy4/4l1xlT9BL4FvXGTVNCDP6bYXxDyQEwZV3z
6/WuhW7ewmWZUfFswaipIps7pNGIOwzftuN5n4DujXdMA9cVpeYupOtMOfiRR1hLB4Yo5pWrQHpF
qsI43NYRDPmxygIbXAie2gKGYDdbLSUXTGBhuxmYlqN4crDByYbpcyDgQFHqNfHeuBjNBDRJpWL5
Kmr4xku90+r7rLISH6IS4CHABLd++/b8UdQZWC/D4xLe57USx3mWdHlvLSOp1XX01xTMmqOMEctg
AfGblO5RXcyTXMRg63KMmfy8cxLELL9wWcxvPUzIJowTRKvGY6+A46YbYtTH1jdYzW+WsNK01fgV
Coo/kfnziuEAZhZSpWSkDKmntwrES2n5HXp3KLq8XFZeEqXBHdN49eiGWqzjg64OkAO5Jax6kgvl
SFhNDgqKiZtZUOAURqgtWmcWC7sorhVvMM3bsCalTVhu1fPTM5Rr+VPrISUUvZuCmUW6zU/+2ohB
ck7v0nJUzGz76WE9rQZ8289aKCIBAbIvvfp7ipFaQaclgY06OYe/W7sbLTPzH+t/WNLH2bvtZy3Z
eEcnTJmv5ubfUA47x3/QP2QLg6DOexqX2lkTHunheyU688WhDb/nRWR982TA383++1ZcvgNv7r6G
zLyeNPUbOHj7YfGCtod+jwpK7S9g/9QDHo/A9ijXVtvo3SxTue4Ufn2QPIZWIAVtUGxbXIniRsPJ
ARdDPhZOvcnwJzUQz5zZOqOZUOlAgZiXbe4GyNKFWrKfmBZ09jvXDVIlwGXztfQKk0ySWbsLjadf
YLTAXn2u1FASxePeWnuxp7TOlfFrFSGCdidNk/oMg5FYJRvvrcOpFcG/H8DJeQ/znzkdkVC9Qspj
khaXeWpV8UmwS7WHB0pPI2QfBvO5DUazpoTkf6ZSQYMcdBrY391ln2xACLB+xDMnTKOaQ7zW0N+y
p3/8STekCAqrwuh1Zn3QFujJHiOEptvAdtrv6EjD4HQLZaAEuJX3GIrAoe4mHwvB2ItviVlephYu
1S2U1joEDDNJIAeEbjmHRicOrk+MAeDo6A9DkN4GLc25r8TMtvFlGeSXS9AEENtmeJwi/ntZghSU
7EHqrXNWuInRI06UUVZ9dcBeZD6WfibQe1kt+JWxJYOp8e09ltCBRlddA2r6ftVXf950AVJ/VC9J
h2dPNbmcaNZwOpSFwXciPaXR/9t9M6xptbp1SaISRX0yUmedAj60mYlK676hbS2A67+VGGFXbErq
t76o9aIv/qGH1wrQqc/KQ/ylff2YmSmtr8DyZWzfIxdMiHNjG+uhFZiznwBSc7oQZMe6GMt3f0E9
9A4lHO/E2pen1vrlccec7dlBo/FVgG24RdQtrJxicVtZEk1kK47DF2/UP6DLZJNO+nctz8+lmRNj
ewb4zJ8mH6lCBaDrrI/w0LZVEJWPDlUq7/rUI12QMzutJ0k2pinwbtJ5/Q8Tn0gTEfDVlUd2Ob9R
7l1/8tbfKL+bsEwmXUt9vjtlJFg1VeWOJZN5bD6lKO9Tr/XYaW8cdX+OOW7ulu58MSNm+60wkJF8
PWGDqmo2G8Tu3NoW5Hpe1e8zWyOyvGIZTkjBwxkX+9YCUBn5ejRVT3rJkLkDq54Op8lIvI/PeL7q
gHVqbyKHACSs7FQsa0dFRtGaDcCuW50cXW2liK6h+Rs/ARnxXuXziCBRqgnmwu/u8JCmG9AFwFd+
N1IpGpQt6SsbUqtOph1h2+4QGE418bgUaavkTgIQ/V0e6iggrYI57nF2mlCZOfyBCBwevkuUANDv
zzVrxvWGvndIi7LaXwOfxmk2d5iV9+fe7Tl9v7gJC0QUqhUg35IxhFmTCrhwr94HLT3mD1kak2H2
i7Sg9lj9CP0dbrmm5DX93+gafZUFB5FGeiRfshlgRKWJHjioEhswq/W/FB2qDHJDHGxMuhx926iG
SmBr1AOy5glHDD2VmhW7aBVhFdLd/bX4udtE/SSBKpYO0fok5i6LGU2/10VfZH98W3yOoVb2Dljh
jXJLQC4wrFwf6ZsMzJUGAg9mm6voEKQFKw3UbsAmn3js34HUlk7MsWMOYryDGdcZg2Te40aQOblc
NFe57jBX0aocUuP/DZLr7xxtl0D0UCtPy2L5nIkiYD28cX1KLT5d0NJdniXFlQgs9hyjlh7EJPUJ
K/6pDFnTOcVGxRcnV6PIdt3WUqtIet3cf00s+ppe2y2HVJduL1f2kglT9Pmzs79WpAfO00+pN3nq
gcikNbj1+ZdMyCToRLGy3B/6SyoU4cD1Zqlzs4GthTXk/AbiVO8lj4R/5dlMQeEtwcBzyMvy1AXo
zRYabZmu4SpOpC/abQMW1w1ajd/T/ObCS1gDTBHT7cMK8XVd0p2twFs3E7aPRY3I3+ukpA4enFHx
5UixTLTqPEs9apl8fSlBL7+Y7lubADNWU1WSPRvZHPAgxifZnl04tPjQrGZMOHGIAo0AxNqlxB3W
hZ2RMdv1zHs/VbJ6Hv8mQc/fRgvaAc8JzX+5b1gflBTrpvA3GG1cTQQtJIl+KPMDIPslciY27abr
PC2OMRpErr4X9/JZAc0OagkyDBNLVeI71dXHK/xvrDNxuA7+dNLt78LtF8aA1cCjqyumUR97kIHy
0tNcE+4dH8iztXFZvC3XQC3cDpn//MWJPq/r9BASc30FUlDsNRYiCclFJjOS/JWDP3PbmXWs3DNy
h2Xf5Em0+7CA5PGae5TH8pxETCgK+Oeks5ZIwnIGB7unNdG1rnJW/49AoSD040mZSwnD+72FtkJq
fwfLm2xYjnNQM6eJcKvgkeur/ja0rnN2s4UMOEzfoQkmzRARBZvOHw+hj88hN+Ph7WtJk8wCgmKk
RAVhmbzo4dGHv2tXAbzPM0eaxVdUTHU42uatKcHGTJMTB+l9UrJfXT0FTDE4sNX8LR+vO5dc7eZ0
sOT8dOgwcD1uVaPmTmlZa6ovPFn35twUgcwgHP40h14JOIYV752EjAq7QnyWiOOMX4Ulyi0PznJQ
spTiiAw7b7Jcr+4WyEqOopVDWPBMdTrResXp40i7TcBCTgTdVcfbqAal4cCdpzzzGDvPl7w4y5qY
Ixoet2b+YNsGg+iq/0Q+jIs8y61ryvR85nrY4k+XGg+g856/MMguxKXe60e9RydjaFVXoLDFJHN0
CzRoZHGtuIX0e2MZ7vLq4g0BHNCRWrBqugiqHZsBpqns9wViAz0TtzBGavE0i+8A1EudT8SvBeXZ
wWhPlxOFqaDdLt/o9ZeWpxIxWVRlf/tBcdFTWN1yh5pgdhHTpf0jWkxRVlL6IlmJSQL8ItYGFAgI
c/0CXqgUVGdV8gvPIymYw488JlTxVqvtozeNgCp00Hkv8orSfySP95bz+t3Qk7WmPD+WIkNz58L+
LAmhGFm6LSaGO7K7r7rlyy8FeRYLMQ+2e3H7kA4zTQI4aoEvNvor+gj+jZEZ3L13LKG6GzmnOUWj
wNalPY1+xebCXW4O9+0SbGKGk578xrzlyZkWJdLbUWmC00FS5LNxoaHRtcazGTNxzxUHVgl5ZlgQ
aKBuHwCnz7YxnidZvljIqM8GQAcC/YVsSj/EZWSt4/2p1+gTEmKWrbIrU4MtraMQARMzVr0xNrRr
yD53ujY5to2QHjNNr37u+iQN7HHoflpbcqIE5icWv57HFtHdanNv1+6EmgEqEO0Ta7jjrIA4YORw
9JgJOvB2g0b3oHkggsC++AoA2A5/j6tTOLB8QHYg65w1s7s60DoLLOIViKrpQIApblxpzhzAOD4H
zSyMOW3kz7gWgAZMTJr4cFdg4viol/fS5shjP/M57Yj8ZakZBZjXdcKGOrpEVftpbjT9CJE7Q/AL
IVg1fqxZKpAVkanUPhumqrVerJvGda8wzvIgC1GWaCnrNtM2Q+vNnb4yIZt9q82HcL5KerS1hUm8
JGixnELveIhjapACNI4ispdFyVz+6t2bqBzJz/Qjt2chUhco14r8+Z2J6mr16s1+1HnThaloqS70
HYpnWx2z9ettnYmHI3QWIcUlv8jjyttbseCTV+CpiOOgLtE/febng/28B1k5EZRjYZV6QLFkmFS/
kvcINEetuoL1p4nRYgOrGtBoMWbzvZKVB11rndeWKQgEdYq8JevuH4QFTt+pJusn55RG//fpzT9r
ojnoospcb+NxxddsOpi3ktVxmVcolmtPLbX78f/gfqY7OiNdLvT3dCbTtxNaAqddvCyfNsm8+E1W
wW4Z9dmn5+VJbTYWPZDgMeOIncHOuDSDZp3rrAm+ZQRNDnSXaMOXBA6DPst7A2hwt51Q1+engP2C
AsCARbUCuVzXHAAZC+0NAveKAwjVES6i70VywxSGyNn0xlyog9bLFH59rWLxWx0F2K8gXhMAPGnZ
sH1T1OCGXl5GPv1UF9r4XZl9vOU73W5aN9VBMmyvcyMBJu4OcM3tvEpg9fp4XaoBcrQNlJAhHBdO
n+mfZHzXr47M/pCxzdSda6cUshQlSWU5nRD/kGCVEQL5WmhvtozSK6cvFLGNy3eeDhJh6aTt6kzj
8Ayjx6bCm6vbKFrTLAWP77/eUvC05pPrc/Fq8zRgRGFzhnFq/ZnwNHf7c+gsK+jtyyzoSKfeaTZ/
cQasg7gjXfyTZyVDugQS4fmjP7YZClYfq1dYVW4xTCMLYJ+tOVTBOgsVfRm2D4vLAluAIQav7Jpt
kuKQd3oFAL2ssxQJ6uhIWtVtwRBagNIL5ihkNTn7A6LsXA8a0dt0OPYbpZLZn/TCrD8mnywr3uAf
rOkPjNPEsrMXEcNfOXN3JgAjKd9vzzE2QiEDpUPAxvNZ0zNO21u44r06okztzkQGF9O35ueweUue
tPZhmMJqEIGWhgggNmJ1z0zL62XDCgZWaJcxOwuXCW7MQPE+bR6x8b+V/WbGm2/S7FV7LwUkJmAr
HSUG4z+4Tri2y/rZ2Hj0qV27m7k6r/r140GjAThuihb3upMcdH/DDWmukSH1BhSnigjE242USMsV
tvBggFhTm6yCACSKBy0ywWTrhK1/l0hrBHPj5ihYeHC1OMeRc0SkQ7Bvxk3u8VhjuIXJFtgsiWAp
D5mZF/o0uCdKTqb8RFkGGBEEFkPyXfCB4EaoMKXsUSoXOhhlBJ4D3iCV6eZkf53RMdkTSf9mfGqI
+ql1j0plHypbdNS+SzqT2zMw8JC5JLjVJxb9SubnoInEnakMl3Vksdb8eae0gyRuFt1vchWD8ohH
str2z6y/KSbTG64qDSsneLk0sfiZx4DnHdtHohZJJYv+YJ0Nq/7WZ5o0CQ==
`protect end_protected
