��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$Rx�y�<��wA�*;�x���@�̦�W�X�fa�M-$u����n~�%���P�$��W��kYَ���P7�?UMfT��q�6�U��k�>����~�\N�(�����X�e���/6U|)�X2pF�]$h���d.���9E��WG��L�X"]�Ad����ľS���8od����e�GT?y	7�������ݵ�^��R�q^]�鍦�����s�ae���h��L��P_���ާ��YЭF���'\��68�b�[����w8�[X��V�F�0͘3����q諵�uW� �h�u\V�?@��_6G�_�*�G���B�絉�f������[�G��U&�����~�F��AׯK1�`c��[<��FY���4I� �#�G��x[X�=�Q1��`��R>(�w����R�O�?����7�,(�H\�#h(W�EH=�������yq��Ѿ��aF����:�U~m<|��.��0=�P/���4ǆ���T(���
�;BC0pF�Qs¹���|��3QU�4�;qA���H���D�l/�;�� ����������(��0���H3N��l9Q6���C�SdGq�V'�̪�5���. IY
�*h�_O�lJ���3��=�9�zh/g[y��$U �)0�Ù����-S ڢ��8I�!s�,.��n�ir&B�� +�-�����-95�	A���Ww��z�����u��\A<,ͫ*�/�Os���DKɾ�u�/��:΋)N�z��kW`9�@T�כ�b�]C1Fy��C�WZx�sd���RQ�����'w���ˋ{iML|���Tˣ�#�!� 3��06襓��4�^Z�Pv[O.�Mi�}9�A
υ�i��/�{mG���ӛ/�l�}/�eU�Ck,�q���R9�C�N��ꥻZ@))f����(�E��%��G/�
峯{����)'f��T�-(0�m�P�� V�>�J�Z\977�֊}d��JC&��{q���N�KJ��n��|�k�VA�y ��}�Ε��[�cRl���"���h�f�:�S���,oI.�^��6x��-q��$K�1")l���a�n(.����n
4
�� ���&'Ԍs,q2�+x���(3=mS�@��2O�[���ߨ�3/D��E�iF��OX�L߶��w�-��tn���u�� VՀ�=�̲�������8���bg@q:�x�}��g>
$���/[�1��l�73c�ћ���4��`�����d3��hb��� �i�Y�,���R����A�Z�)N�M%���gm�hT�@��C������Ź�������������k\��{׬A
�!5���P����;�5�\���&U�]t��T�a�|v�]$��=���0	RX��{�
^Ϧ�~U�e�+���n���p�}g�	_ȅzSd���$"CFkC�b��82�Su�4>z��Q������$�3�����ե��&.kT�]�(J*h�Ā���S��D�T�@���5�v�+��rp�k��B�o�K��M��&�"�oQ0������R��p��͛�/h�P�J���\3B��>��h�<jws҂���b��t;}#���E!�>9�7�XR'�%� ���E����������3%!�mj���g_b�ʮr�����ZU��tH��N_�B�읮�,��U��(��R��c\�J��EjẮ;5F�"�ࡕ��ὠ�p���֮MƐ����rU��{���U�92@JZ��!(���L������:sY�PN�� ?���˦V�F~�Tz��Ż�_�0����{g��wk��/�HF��ͷ�W�eOR�I���;(V��Ԅ�U�jGp��oIdrsx���c��~�h_"ű��=ٲJ*���\��!y�/��ʌ��Mύ<~�4�~����5t�9����@:� ����g!	dϪ�L��/��oG�}�B͔��~	�����i<�	Ǻ'��KD/zk8��� 5:5�oԋ��萆����Lf��1���|�Q�]�	�� �Ү�Uw��g3�Ms��]���O�I{�� �l��DW8�n�]}z�{�'�%�L�_V%��W�i��� �<�g�S�����&��>^�/數�����a풟�L(��Գ�{ZE�}�V�1���qb(�t���"%N.0*�@���>x
�T���D� D�L\�%��jքqG�znc��c�8�#թѪD�X�m��V�ᬶ���8_� 9gt�i����ʶ��E����7�i�:DJ�u~ّII�[��z5|��|&\��J��*'�J^Pڋ��L6��w#�b�e�э�Y���Ϙ���Wf���Ru�5�ߧ�0�a�@[@�l�O�K���E�Z�AF>.`Ud�%���A"c���?Уk�`�B����9/8A5�p�	
FTd�L�?�-�x�(��MX�3�I�ۙT l�:��&+ð���B��5\�rU�\v���v�YM��\࿆���C���E�(�"�7���XR]���<�E����+� �L�݋�m�M�M�]�
��QF!V�+;��NVqD�9\Ta@�U�����B^���L�6][�I5��P�"��_W�T0�>U�Q`0f��d��/[�@70�4����ƒ<I�"l���q�QZ�ժ3o�PΗBJL^{y	�r|�]�r�d��w݂,��4E���ȝ�o�3r�i*�آ�_�ȤFWɩ��b�
z<ե/��g�xk�M����-���:�X�R:谗,9wEI����h� �Y4�Oj��bu")hL��[s���_��k6�(7�}�J�b�?����d�%z������q�l�'�9:�	 j��&��H���(VSڴ�Q�O�0�Ep�ftİ�����y}�,���j�Ypx	��7\,���t�x�倵<KT�7����7�廯fX�ނn��$�yI�?}"p6�h�	.�HC�)c#��	�3�*�@�$�����b��c@'�ַ����kQ���]�Ӭ�S���ܾ��o��O���/<�G3��^�{^ª�3�]�������'zk�0Yb�� 
`�S9g����rk���,�\��ǻL��i��IkM�:)hR�*	̦R��3�A)*����I��u����[�xWP����@���d�)�ѐ�wȩ�î�L�?[��=6�uYIP��+҉8H��-��*�6~���~��j;��q���5�6��ʀ?�c\c�A!���t�$���
��(���P�R�4������b��T��\�ӛ����o�j��T4��S�.�m�ƞ�k��
P�[���-BD�����c����cI(��0���,���H���g6�u�C���J��
�>W�!�Gn~�Ą`���GP��d�:>���l��!rӂ�+�",Q2��^{'os���=�pޟPY� �HLtb��By�U�0��z�݄����
���Js1~$wNNEz,�ZL��Q�Լw7@3�����g_���ny	�a�?��v{Y� ض�xo��_�f�b�E�1��˧2�#���l�����Z���7�`r}z,��If!}v=]��?��L���Zd�$�`Wu�콉.:]�u|g>5��-p�|h�����
�F�7m氜ڧ�coΔ�xz���/q�)�Cxa�Cr�oF[F���ؔ�p�����ݔ�\8tVR��C�}^qJ'��$�u$y �8�~Z��{�����m'�]c�������#�N����_��$�5Q���
ϖ�����Ib�L��ŵm�;C�Q�.�Ry�����K롳*g�Y�-q�r�m�?b�	f�0���ǳ���:r���3��.�l���}rDx���L�I:7��'�u��G@}���"ilǡSq��g�@E���<�%~�����\�:�`���N�v��`������/CʕZ�.�"���#��?�IH_;C>�挗"^�#N�S;��̱Y��QC�h"y���|��A���#S�^X���e�,Ź6t�k
����R.K��L�U����*pPꨃ�����T�ѡg��Is"�w;�q�7�Ȅ~Jl%�)u�#�V�V�x
��D�Jg��U��Rتl�bK�����3m?A���@��R��o�-�w�E��x��H#1��邨�������7�;��!�V���f&\��!eD�@,��`��jV�25�#��q$����z�@_�D�����<��X�H3;�L	9�4�!+�'^$oӪ��d�^�������J&���8�����F[ �ǧ��bH栉k�j%���#c*I8�X�>d�d��X�c�  ��H��F�۽m�U���*�oͩZr�l�R�?g8*������s���8�������b��	� :���@����$uM�r�S���Kd�P�TG�"��å,���(�-ϯ��� F=�Ӯ��2�wx�n�	�2�'�w|ض:����K��ޏҽ�)ذ)B�Jp)��o���Ģ���_0cEֆ��{p�z91X6ta�:��$� \7��}�i�� B��=����L��Z˫�͝�t��7��!�qږ���^[_No�Y�M,Z��;�-���a�/���r�_��
j����\�K�D�f��!�*lXF�Xt��(@M+>��z�py���El/xa��b9�@�a~����f�M�������f0Q%����eZ�����Y�\M}۰#��#ԏ���gȈ�a��|�N,f�(�7��H��o½(R��w�z�u����Ï�;j	���ysϣ7ن�-�Zြ�,����G�Ko�{�l���}b<0��'7��
F��ˊBk�����z���d!G�K|�@��C1Շ��L��}�����6�!|�l�T�v��H�^��*�����{h�"X<��n���(�O�tE�7�r�p}�Eup�L0�gI�F+�K��O>0��l�'&4�p��B�pvp��Xd��X³~���_c�v\�v���ۢPM,@MS����$�E��v$Z� &��n�M9`�W���B��r%~�h����:X����<=)�Zh0� }��Y�dÒnf��'�=Q�C�׫������ceS�a
�|gޭ^C�ؐ����9YF��s_��k�x��v��|��TC��~�܅��}I9{�|W��&;N}_�0�BZ�����'pO]����R��37I
b���~�$�CtuЖ}�^��<w<-�Q�C0B��2_��V6JPfb��O������MC
�Y3�B�dV���y5o�Q?�ۡMP;�jL��r�3���T�˼�G�<{mW��ߴU�u����m�Hd����?��
1��1_Y�a�z�K�1�+���.庳ѓ��X���ܤ#q��m �;M��;��f`䮱<J��!�c�J�4�]�C�%M��^�?C(����(��A��'�j��1�	��[���F�-&��e6XiL���5�96"�EkaGI]�%���6q��Ta�C���b��`ɹ$A�(P٪�����p��%�+� +��],�uE�\w���	���A�RScG-�=�r�u��M��ͩ<͢�u���Q��W:�t��ڇ�"0��ۖ�'m��@+���Nj9���f��#�ӆ�v���Zo:���Aw�{��%X���v&1�����G�S11*�+_W+M/Y��B�%#��S<�$�2���,��%�hH�i�t��L�ņ�s쐇�zu-J�8p1���KQ~�}h�����:9j�ZJ��s�����ѕ>7�M%�0o���D0r1Q[�7Q�Wz�[
�^�,ӓ`�SJ#�z}�T�!�@k���K����%/���p�PQ}ўM���~��wJ����w��-4H8
�58������1��E#�C.�D5�߹�;�!��n-[`IC�NY�Z�1}z�@�m��Z�[�Ov�>���,���O:�\zM2����i��О���6Ȓ�qk���C�T%'��6y�w�X�l�0���,�����mU�Tdjھ�ј����%�����R#H�S!�km��O�Ws4햹؎l�>5�;��/��P��Y�A��,����QSd  �n��R�]�IfQ�[v��K�A-d�X���)k<�zǄ�T�o�T�'9�'���|���j�?!��;�Uč�M�d-Ɠ+����hJ�.�����6#{�'f$q�������"?��b�J�i�Sk��D��_���ւ�������o
���K-���*���&�9�/��g��a�4ѡ(WK�u�:�2�p ��Xo<CNZ1I?��BL�/��?쁆 ��}�ec����a��Fa�;�ہ��j�m��λA��3Ijx��#�l�C�E`�$*�]�)��B�]��nQ��g.��l:�y�"j�Ƹ>��	���_ș��88�H@����n�Ŝ즇.8#H���B_j�ůTigAL����С�nߝ�#ע�تtڅ�;t
��on�r�K`q�D�J�ўy���Zp�d�:.��ڡ�]��d���6�V䣺��A�4!���� �ӫ�WM��u�BJqI��#�B�ۻ���L\޶=+p���1"o�e(~�#F��=z�)����P��GS�k�K��`��n���ۻ�.>( ��x��?�k�b�e���Pv� ʽ�/�bs5�ꔚoHv3ɐ<��l��|�����R�N\�y�;�k��zT>���=���m�lhҏ���cd�I`뤅��m��[��W�
��3���|Qp�O���t/���Z���:6���+8�α�8n��y�lL��58��ğ��A�8���;�1��@�^7��3��K�k8�2�P4a�z���f>���R�&�����U�r��Hٙ�fǱ�<o*}2����sś�����͖N�+�%�Kuw��y���^kX��掺�<�VzN��Lm�ܛ/vy�Z'sW>e�K�������J�*7��*5����5ѳ����~k@������{��? +��p(�2<Ɖ��Xk�{Aު�D�?���I}_�`� b��V��%��O˖Z}+�w���j�r�ɍ7�RشC�%���cG�'�4��0�W���D���jM�.�Fv�_��)UѤ��wr�=-���ez	ط�d ���Ұ��A�z�%��b;$X9�߯�� Z�1��U�Hy$u�$�}rP�K_D2V넫��-&���� 5w��F	x~ū�Ĳ{!Xz'���}�y��bS�*s�F� j���ڪ���c��B�*�S	�;���*��K%�F6"��ʓ*��Z����=!>��CF��rib�[�^�)�ª�e���$�@"��E?�+�с��^@! T�v���� �]g&S@����B��za�����1�F���f��k1����؊-��M��'�=WtKt�>s�B`��$�N�a��2�S0����&m㎓v��-��1�r (J[(�9,��� �å��_�R����gL��;�z]/��~E�f�T�b@�F
<��P[E�^[}�q���FWL�mޤ����5,��X���wvЬ;��<�����җ������_i
@4�!k���to�>����q����3�����l�Kb�P:�`���bs��Q��yO��H|p�$�WL^�鳭 u�b������5�
@"M_�.^��ye���iw=\�l_~Lx���ǁ~�d��!�N4��.�L�|��O�\;������$��o�`�ԯ��$�l���W�m���X$�+lκb��ᶆ��l$gCr:3�=�y�X��lO�E���$�.�@~�)�o����y"�a�{�I���x۝F5o;�f��!��+`�; `+�5P������L{�"�ZD���5���/F�r�p�������_�ݫ �*R�y�+~�]@�r��R��uh�P�<!�ℵ�4�gU�lĝA!��1L�=����Yq����l����-�$�ƚ��Ńy�1�n�I!���\_`���Q*�ol�����3M!AZ�� ,>y�Q�m%Gm`��g��?��3D=I���;�������K��L����?}iIYW1�nh�=Ql����������3�}�>����òLA!�w��;J_ ��w��Cz�
s���Z��S�I2�|�@k��f\�ϕp8�����-u�ʞ%:;��6e����Nm+l��f�B��)�-æ(���_�#8cm&{��v�u�ߜ�j�9x��Ū�D�������~,&/�g?���Zh���,���t%?W�?e���sᢷ*�J?�Udw˘���ݜ�[EO�Ŵ���C M�a�E�q���g��h�ޘ���K���vYxh�\v��[�������2�O��+���8nI.�_�[�~D a�5�ٸ���g�^tv�>x�&��<3١.�΁����MVY��Fl�Jf��a��%&PKO܂年	�8��t.�9<Lc?��9�q2�;�z��<���$;�P�f�ޢ�;z}������1�P*��홾�7��X�Tn�8�b��Ji��o���;����I1��	U�HK܈�f�(OQ�����ۭȘ(�s�j@�>��8]m�4��B,ꪝf-h�ǖ����z��l��W�h�M�/���5�^
��w��b�׫��IZG�8����8��n���:i���Q}�S��1JE'��UG��q�6���K�<X�^Q�"���c�i�&��vu)6����3-q<N4�/#����ٍ�	ay�2�����fM�,�\�U�:�#Fk�YB��)�l�m�	6����)�X'Vc��V�ߨ��@��]i�d����U��}>�j�dSr�e�g����1s�0�6��T�F ��޷��O���Q�x_���q'�����Ú ��1|���
�-���{LN�{��.NPO++�r��Ra�����
����	�8x�iŬ��&X#���GSM	�.�������J���3����q�vr&6lS��Ԅn�h�<�h6pڳ���Ɣ��Fe-7���rA(�l���w�*4X~$��Rg�s憜�A�D���ۻs�:��{l�Z,�\�'�/;̗g��Z���^�AP���g���/������l�aAy$I�Ԓ
2#��L��q&ա����ە��NNML��22wQ��D{��ڶ�Y;�",��W��Z]]���o_�a�[�;�h�Ϫ��[pPT����L�ڎ��*#��0hM��f���sA�vl*~����Nx	��<���qR�����ؙ�T�cr�����'�( �x�x&+,A�����i�@`��ujb
 ��[�h�oJ�Kb�ґKK3��s�Ѝ��m��	�|\�*��/U�a�it�K�BM�8~