-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
xOGI3hZRyRKxFUb5bIAsDVP1aEuzdOtJ0Fh4d1isvCfsfKxVqqg1yZaRxoKiEFMCkc2Q+jIeNSHF
AZPFS5MUvC5WLCdqGBQBMZsoqWBq+LdCAmpIv340+VqHaETLJRVljGVnEPSKgOiM94J+op/kTkpi
V2qOBeHUPbaDzXKXdFvvrO7rKf6YcsTbIZrWtfbx1QwoEGOPNUg18cOzq4oc+qkkiHw/r2stQUKy
nNznV4kfwZOsLQKP4+8WTFOBNx0IWLoLmO27iTNEBDxKAP0eQCJYanEyHoEnHFDNRYxTayealSvZ
Jkw5fiBA5iRsuX61bqDX0vNMJEYowk2T/BCc3w==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 18160)
`protect data_block
7lmS/2M+RqCHQPFGx9RJgmsmVBhtnRhWl5zdySycGuKFKFQxBTMGtR+P78I+cJiW7NHLuviuHaj0
rAm9EYiKhl5j1cdEUXWABjJPk/AStDDcT4ee0Gk44yK5D6IzcUoAiiYA+Zz+3sinF0lWFGhxlB+Y
IwmDJEtR2FBXWNSvrttph9YuVNU2DFjOcz+LgyozH1zHuKmUSBBaflLqn4KUiRDK2rgmM1GCHFnP
wwQcu1cpR4dCm9iCjTemijwAQcGuSgGqrqKNaq3iaNqumaW8Ko3W/tSzvByHQHOamRsSb8cwlAf6
SLTbJbRTN4+AVi4FPi7rliQh76iG31VuPBZTuwZGLVr+WsKUnG8qgBGD4rrX/6qDZJ+FOEoMX109
MM9OfYTr2M6A7G6Um/ZknM09l1XwHE9BCn5gpdCVMMRONXg2jAqejMzPeu1Qnwb9sO+KXWHF3CH3
9/qcok0V6XePoGnjIsPCzE2H/+YtsB192icDvCMvPL9p5inM5AtI1rJ4HdDk9CqOvSKiT1lt5/BE
e+lW/WmZRgKIo/T563Buk+W+iOhktN5ZRDG4kiJM7EXR4xID3uWfnJMr65dnaxE1X+gsZTLbGD7f
Nltd9QH+vn2IbrOu2oWyTHU7OONDL4pOsiOnq/ukXKbTDRawltuCdEsKt6fcpfGWMd5fIQOyTjt4
FVWJ/im4IepW+QnEw/dzfs9aLNzw36VQ1PaA0GgKFBXtbsYCEKE0X8hkxgVRHCvBiPpxv4dm6ehk
0yXEdQD9g/yc+wg0grqMvtgc5NJ36S6ICBJGVPIn3Rj86SQgyWaRT5gbh1cdkgq6prAa8Jo8Y4yY
gXwyqz/bXFreOsu9MUKFNg5zKGy2MM1wzG6XQ/vrEcJUU0Zgs6zEerMKV/d5ieltQj1sgXuEypZP
KiCvfwyjsso5cggTAUPO/Ejf0MKZOBjpNYM/B/Q1cl5ufJWiJSHhSTvNhanpQjAOZt9CgdD/A7Us
JxPA8AI6nY8cdveLZXGBUWNVit15Y43ITMhB9JfxYVFdflGhkVdro0ZJkJKc4lDfwml6B6MACWEI
45HpO6NDB4SOJI40EGxyunJqEV9uRpChTPEGf9EPyahAMjsLo1pYVSW0tJl9OjMstNq2F/U2ESPB
2vGisH6KjK0mlyctV/LLjEC0X5gEsOHA8FDYbvb7ajvO1LMg5doQIv9DDR+//MwQvJMyAbuJEvhc
jZml/Sy5Vlt7fyOj8bVhEwzHfttHTLXAl//1mXbwCVGyhWvEmYGOs61k7k0rey7iW8EWs2Tf6WC/
2DKnHOJEaK4oszwCBxtjrGz6viU/Y817kDTS/0h7EzAKNpMAyw9Yisy0ExUqtuQhy7dlpirkYdVo
A/QnAYqd+suznpZtVLcxlWpQStAf19UGGhQR5uoEaiGstBHY2TPYvGtGMVzT1MBCXOZNWMzMoeub
e7QlpHIKEQE48nDD/xxQY53tmgVuj3hS1Bdpwa3hP2KfuZ5niFVM+qV92v99bJdD6Yo8Z2VQ/3go
0MJwEJ/WqQSapxu5AJumkWlWTaPXYRY+/CeBd5yrstFemIWVtt8OzyC0BVVc38n05H9xmmhVLVyJ
cXg2rzN9aA9r2EJBLSRQL3LsngGekO6j+vM9tnyAc7SE5h4Vq/pnZYhsGmYJq6g11CRCH0VuIZ1P
nTs4bVjRr9voE9jMFczuWVRKZUS3eW/9IgjMme0rnWKjlYjT12RrRNb/BZ2t4yoq/lxbqkqZ8rvq
bms7wrCGGtDuU1ioQqCP0xDyTxLy+K8NeJDQGDEjwkF46TkKP7g2Yedx3ecdgpZt+6WHa2hpoCj3
RkcbGFaeaDI8Y9E6NoDXiqye8t4vYLj+MRapaANzBkqHMhg6vbVoq9A6cL5r427LoNynj33y80I2
KYIQMNxnxcowLczNszeFw++pZNPq+v3REoTuxIW3tYYZSTErXqMLmJEkpHSO77HvMyXpay0ZbayL
usKoYyn5eTsTP/KKRkhDXPKLAXEmGHARwZfGcLATWf0+znWTbRcegfE8gCbdULUG5EYlvGnw0hGu
tzllC3XRPxX7TByppi9LoRWjPVnjVlWQBW92rX543CUAbJ1jv4cH5L0c6KY6DJOTurpoX4fK2KDX
9ujnVxOAK3Rp1US4dQCj4mApcHlq6N/ZSXHaR9d0JoGBqBlq7gktiExb9JtfnUrhGO8n9pSXRUq3
YYYCNvVsefz335xHjZ9gueYwzfsA2vCGgEyUM9fNxNzHV5msKo5Iv+pqFX0r7ApJnSF7Qutkk8GJ
0vQR0y66goEaoVQYEyccygvWY5jXIpOlBdX4Ci47tP6/F6FqLjK/kB4C8939n6GOUXhFEN7i2cvm
ZnfN/vhR25W+WH43ECROj+CaxZiU8yhS8Wd3oS95MXPYDKhSRAGKUQpjYESpBaN6RT1H5DOVGeyo
xh7hPzqt9gscZIeYFClSCWp0OKb7EAPy6NWS35KmKMvIo4aJXml9s8qIllTRTDOZP2eC8VmbKN2b
oEwdwhxea5iwZpsw7XBzoCZj0y2qFybddEb03EoQBUDTU62tQC4NDvIFFUcehy0w/lJqOm7V+tbG
VczBSnrqAnywHKWQBBRn0DYT626zvlxbnCzh9eOGXfDjfu/bZr4cp+prkuGYel65UVKuqAFBT3Np
VQjB5D+nm+wCWDxXTc8dR2XVgQ13dGUIY+KsIuS4Ra4PBGj0Go1EgBtZ+fz54wB2X5al3X+PPzG/
4s6MEqhpqTLOJXlzPguwsJ7QIHjnwHtgFT3gKvm3zG0lp2YYSKFNbWgfQp00nounctnXRlYSQI8d
SED1vOgwP74Y4yIvOWC/jVshcjfFL3RGJ88/ivgxGWVR/8ptVKsJI8tyQZbUFPqRPZhLMpfIDORM
u0IPkaGO3fIuc9cCFR0STavUV//y+uZfLPrDBB0IMsWDokRPQTo/Xn7jA4Fh8qmM6AcO5E23B+F4
+yiFhLh9e4DxsBLxEHj81GAGFjKXlzUwCU9YQEFuHaMTTPRRmxZYfoDYybw0ucrU/Bd8yI+QIfxd
wcaFgH6f1a99wJDkB1scmafSFy1HLODwI23buUMk8XezUZ303uXaew7HJynrAZOuebz8ezFJvZ2h
91O7Y3rPzb1mu+ZyKuC/GhrdVaIoFZ0t89lJh8CKmEoGmrEyKsFjBM3NDm2hXzpulfkesPJPQMtc
uk3ENc0DejARS6nlSAruHeaAAfK3jiNf0XdXQytQd1i7WAZaHNDjpycIYSvp9BHKUMv1srMQu+rj
Z6O1FqwUhgoG1enoxlVWItkgIw7NhP3xV77kExvHkxo4l5yjrFVGJmNITU0AJ8+UUl0gTorAyNhr
R3hZPzBJNbMlG6ODZEnGhulDZxHOlcfKiG5nagaWcacZCDm7Qd3EwG4ASMLC05BM4y05R+hS20K1
9lGTvlOCyjgNH/zffRUWaWr8SIztPG4zCHdLv/dE/ZOtU6eQJ3jN5Fc6nnb7Hv6/MeptIdWjBxNt
Gw9Q4YWeuzwEVcHSAMLOm2yU/aKEMlTBQKTnRWl0krxWOPs0R2W+U9olMClLxIcehSoleJ9uOa3o
ksfUoZdamUeD6L7bPiHFHN0DGycD5IP2SQH0yhr0uIZkuKoKTO335J8excV3A2n3mchw8Nq6Uux9
7W6kiuwQq/09HpzTtM3o1XPv09V1Zw9d+mXhk6YsF6VhN+kmaq+EkZ04nvMXXu/GR+3/64bBfI1B
tXjPphFPsNl51vtNRCP5H8NOYKRlj/JUi8cINVYYZO1PLu3OENKwgA67hghVcqhLPTENbNtywOnk
5lGDVZOeJesdaM+pAP2kcJRuIMES1LTTJbtdHGcoyKjMK8aa11Vsk9p8m+6QzrbLV/QiJYdYourp
bjtHzXy6hzP1NT9IbNQHZGKKVZ4pd/Eqwa0+tUXtBzJd4vAJr6tatIHV6N/MVJDZMC4G1rRTBq8v
SdoqoPYEp0ZSLP8+cUzXaOe3ZxUcZx9lNjMVvd64hmu+ofdqF6+m94oRv/vpdjo/WsxH9vc1GWTG
jnmHgp/HfLWVWoklcLSQI31oXVfF2ka6T7BkYGlrCS/Rgxam7xSUJpRyAQaCJIqLoPL2sD2/LDpJ
/KRx5gENvBiyIcMxfey7wuSjREER2YG+epJAkWpQMnyzlEFAXTaQk3F7mU12Cza8yIsPLM62HjV9
UAI572XuxVLLwDc4Xi7CLu71RcMOhGgxKCTIr47adFzmtUlq9h29Kvq4sDf1OiOxuHvj2Jdn5lal
UcqnSE3kxDS/06OnAJLfHNgBn3jKuYbknj90EZw8oidmqiAgXJVsg8vaf37PUe0Ops4y51cqBRre
8ZDk4AtTp7tFjDf7XShxhQCDS1wDPz6G4Vw12uijc44Mbdd/UC8CHLd9IHGUgc6zgiBNVH6cHpUD
FV4GtSMpSrJVUwx94p6tgb98PzJ5+j5A2q8t18aEap5fpfFgHy1Gyoa4hTFVerPx1nCQtVMAoEbX
lqihQKbJhhmyCq/g3jeLWvBwkcLYaVoFzrctPJTSjCiv6NQtxMOefX0DRMICwlrCGchxEaGj7aqs
A4Aw8gRGiRufUJx7RA6rr/qwD8LgiwijDEYMyvomLTouuKH6XZ8O0mgrpYXIbiyWT74UltMHsX5u
yH0LJSXeCOTrsrfGZiwALDsLeOf4i2GqXSjKSpxPSu93VpNeiEoidptjOJBQl/Gcfx2W7bhyw1OK
zXuoKycLmsYNCYOBcAAJx1LKDuxWdocpqnqLOFdGAMHVdh3cURe6oZKVk4Uca9cA89jvfu8Wl2pU
t59FgDeMw2ZwZuK2OQbdcKDlKJkw640n9Q+ycuKsTf/ffBz1eZlVQJ/9NjtomvRJMT2ZDzE+k+MP
UcWhnnOsPcX5eRA4iudTMTDfyITnWg9PTUfLzCU0k5Zr1PEbkNYo5Rb86JqYVaHNm1cQe03U1hZU
4FOy9zeekOA5iM3QBISDmqjD/+UJuhqzEB5QvBVSNF4JRcKu3JmMDeP15y4jk+r43RhfUHGLo6JO
jV5P0ke9hkRtyG358buCsfFSfuQky1A2EK8NEWscOROqo62lq/lOvb5gICm/ue56D6QdkyuSVCmf
Rd7gcVYA23zSKeEIzfxiE0FvuNi0GUp9Plg+SE+MmIuCSGDdpuWIywpNpU3ZIYR13jGeWsx7BLB0
2t9gz/PCBjTHa7p1NeTIv3dcOiFQNT4IyPToBde8IDqiMMraw1PiIJ8ffi24lYA+5r3Hu2ua8Cdb
837V3KpBysV6ZttIFDdZwNjrmRxvYS7fGvVf80PTUanJtjyQ3m6+9wRcs2nrnzq/jqIpsHaNqHZO
x+gOISGfbUpVs1SdqRl5xpTg93XP6yhqQf1jACgqjwc1w0v2SMXII6CHno2241HLp790l9eIKur3
G/dNxRGgiJ1oKH2Ud5fp6fqA2SFH+RP1qLlUbvTkETt2N4vsImdL5FhTso16ou6RobIVTyF3pu79
o6zJPSXm0AeczDj4nj6VPzWsvrFKSDrdqZWDhxn1ENznZj5wp1Dwo/64NPXZ+0lPmoZ9S0rJzrZg
SajkP9LMw5NgNByi6mIvuP0Z+R6jseiGwlXFNgl5c9oTTHrTxh50XuVGQ/cwe0sWQ/92XWJ6p8+y
UsREUx6+Bt/VG52NXYeBgw8aBclc+Z/oSuYMcsLsslNXDFzQ29wpfJZYnVe2OOfm/xkiRVhQ4lxt
dNghLd4+QbkgfJwWto1ugCHowtAbJdaPbzdzscjyWQnbTeZpUwEBZd4EPs6DA+lD0ETZvnTPKHF2
7bSiidhu4QgEokUawDPu2AoW7Z8+/cE7NU6N6JuLOCBIarHdmxC3Mut5+Qs3HYFIB/cGtmfULrvv
eqlXyzpKHvC1L0KX2kVUlELuEZQc+K3HgJTr9g/QG+ubdqVjxLzLNQuyYeExzkOqGxSqfkY/MYU/
iMfnCoh4dUUvT8go7f3R2eXOsKP6L8kWZpZ4mnp3CdVD7ISe/CDStftJGjDsNH22BT8iu7pIvR4e
LqVbuzlF974gOdDSw8GLNNa0ESJQQRtQ/XIBwmXEZPKE2yHoCooYmmnqlI4xz3fVe7RQFXJUl2ch
2sZE0JKjfq/I8glA5mtUYb30hFtwLUcchNH78PcFzda49FCobJysyxHer5AeHDZLZzCJFM94IGbE
rt08qAd1GqPd4m4K2EEpnTZt4ADxwVNhlDYcxZHPrBMkxFsqTKKfA0R10iKe5D5NVFeuUBD/LBR0
GJmTdWQsDWy/6gKR8Yo5Na8e4a/BKS2uIjp0xqRPD7UBLC4Aqw+GmAoDWKfpuKUpMR+K2e6rHUYf
ApWqY9PWOze93SamIzUnikLYLm6pc8Hhuu353JAZmNVdoYTK7KalcHmBixtUt5BDlL4YK3hgld+c
PnVA65iLK3VJMxyR/R92jS+QooVFBc7L78KCeuXhjPBJN36ph4Tp6OQdQH9q/x4BAibQi5rv2azr
Fqgo1iQM/BbMYF2hmhmXxuWjcghepj9yKZNUwgHAym2+4s3n43zoUTQXgCis32O1wtxqTgW9sbqU
mpdIcnTF52CCoFC1v/cP7MQ4DxcNInGQClTihwloa/CzBO+PVIMp3RjKKYZKvuhfOJZU92AndSvw
LoXdDR3vgOLt6U8PQy7vQC3/SuqqHHbTnGI6bWmRrNfepiTt1f4RUK1OFG+v5M4+ppVxFUbcUHgO
XuIfOThuX+wvWEKjOv6twc7d5OYZqOu2ckhZIDa9145zlCB22pKAfM7VxTkWcy8iu9SqoPcjkHEJ
ZUen16/4NIyuJS4h2JlcoGtzOEUB8FX6U/3f5u7XCAvH1nxf70CU4dkDv3F4D4t8NWQNF19qyENg
PZcG8svAurMNlGZmAM95OMmbnaTxiH4S2M+3V+t/dOm+Jhaf7xHF1fwwU6pMHNYejshwovRjmMbT
WfEnT7Xn+T06iKxI7c9HhBXkrbor+52fs8XxK5YPnforobYjYAQ1qz/mBTxNeVeqOw0IES4b7DT8
ihWR820q+Zv5GKhD46UbYA1XUuY1GEGguuGbLLbdIDcgLp+jgBYeohDJl1A1BtnhnjAiOcm4DySb
SIxI3itnfDLJA6XgQuDrJ5kxyd6RT2zyxvh2M0JM37h/yL2vKHz8lbKxCQoi7F5cyGJbruYMaLBS
hagPPZmETF2yGGE5HaGV+b96/vPF1SuMvpskIbCJ8K3fYGs3IN3pSj9Sdm3RV8+Jeh7tenbPhNUj
QAgDRC3dRbbn5WdZx1UltKLXp2chcrgFivsWlBP3+AiZkk7cjVDPwix4+mrQSVHP8gPQtKGeT3sc
Pk4AKQPHe4kNiRaapdDjB1tD4XsSsal7vWvxM5o6cqoPO4uQiRbjMt8Hbj2ktLdIzVB1SiyZF+Y7
RTploiJx55Uw6TnhtRcZh8p95G9dwb8OW6PVlVlwexP6xa1/NxkqSY2ecHSYDXoyuVL5EPh15TqG
/AeNm+g1y6lrwrTlMSjG4tfPKyEicdBLvhMsfkX920np8HK4Icj0ErxJNRZcboBSsL0A7rvftL6n
wg0SVCh+AEP8H2EuBgB7tfD2zTfG4/NieGIlAAHJILB/qMX9oFFq0+Vb2hxAP3TvqJLbgL5d7xQ9
3VO25kp1VJI1wLae/GVqpbu1DoKKfyp1Sg1SOK12G49+nLsi+wDVKevHctalOtO9oF0uaTwHz59x
5FVT2BMCoTmivlZyU8NGORq5MWxJMc56e/7A8+H2Q8ri2SgyMn6jBF7unh5xmPZVsDjux8Rme3jD
y0EjG8aMS2RPTzOB24Okqirl0NfBidOzKE2LovNzEHyUBTC+i//Q7G4IUm/+pkhXhRkROeM1aEZ+
eXtiF/j2xpbQxlmNhHanZ4zKIv563CRGO/m10IpjtWFVCyJhwzJhBJqzC/rRgrRezLmZ0YvknSZm
r3SXsspO5FVgDB5OgE4s+DB7cP4xtO9lYnmWBAYNbxBblOQZC6sGlW8ElNSU61JW9AAKxxVMW5sp
2NhuHruUFfNcjbXqgs4vKGgvmdSl78i7a1uvEL6wu6hySxBezOfbPdve3OnT5mJxhgMF0hGqNl7r
eebte+7OLRmcMPPGWEanT99UVwH6a/c8FdL9EJxc15mJLGfX6NClOYuBp45kgU0vTrFL1hhBbfD7
VevE5D3tIXNWFSk3Q3y+K6NyM8aDxl416rkUpHBCM8aIvb4TQ6dpBWJ43wnZ1kxqj5f3az5mR2Li
iK+eQeS2kNOzNQLm/pJ7QRKEkjVgChBK5pqDfHlOyXHpILv87/xUVSv4/XtV7PUEy/3JAEVNVsGf
1FN5Mdlly2ubPWCsodEC1EI5hPJSsHOiTJ2WxEhjy+Tgtoocx4ut4sO8JHtYpmgQ8c5WyP1WL1qY
Iy874ray8rhCVdm/1sSeKMXznZqBpYAM7ueytC2zlHl1v9r1mWsNCF9RoslNbS82+lkv9xHarkLL
v3ENrnZKrju8ng59bvB5ewY/FJzU+dq34BNDhtbvTck3GI2Sa6C830Ks9KTofc2RwNc10D8iqC9z
9Tv8CpbxrU2YQjmHLdvqzxJLNV9aHxAktmMvsQd4N/PbHXKfIwSJzASA9a9gBW+eMsDo+FWHj220
X6bgdTsGh7OMXKqjaI9OsT5e/4VHY9Q8FsHNiVOmMB+W9fwREI4S+b+k7ea23iNsGlgaeWArBVTI
hrezr/r9fF9htI3okBe0J9SwPZvPJDL9QeVy7sln3l50AJ2Ede9LXXopTXwdfNp90TmvINrUyPIc
le26+mPtHt0blrMgTWu0bd1PRc7sf3op0GrbGb2RvTCPBtRNkKxhZNVFwRqVvioOXKcx9vau2nvS
pe8m1HkNhFX/L8qgz27usVXUmbf6UoaqzhbzIQlpGYV5gu8V0Scy89Z7pdeTiwTA4aslvL43urMj
ig9XWGu/CLl/MLTiwGYBJgoc0e1BWwb3rRsFy7PFp5odm6QBCbFor9+UIqqefWJKnScyFIKROgEZ
PJzi67H0pdpSARDnGcTiHWfUPRbTr1nGqElfgfFAJFfFM9DLjXmWh9E1I10oh4zs8rqblo8z3D23
b0t0yZtxI7PJKqN4iS9Sbmge7wHbn5wDCXAy2jAw81n4RqcXv0Dp4dUwmuSyHcYJNVGR9uY9EwER
Rf4IRnCTz+aB2pg7mhA1dMPWqilPaLYbcK0T7R5rmEDfgaZ9GqS9QLNej/SiK5Ph6tczY01Tckta
w7grN5N/faawufSM5F3vd9ejqGuocMJy7bs5CGTdAgObpQWYDsiiiQjSnyVT8l719JDsHR5W80Dz
NOzJE5nMPxndnhXDvuhsisz9wD6XhlZ9lsbeDXZjio26gvqxamjB4drmpyFhBVSnWO5S6KtZuW4a
jhV8EPmHJpFddxvdz2RFnBzgNSc+xSiboVl0hSIPg407xRdG8bDczSkiWQXs3IGbT2V7uLeY63so
579bLJ6E2WFGeSze0jdBfXE1CdSZcPeilDfyDKlD72qiXiZNULEb882BQ1eDRPBW1ZnehjxFtlH3
NvmGGQmHVHCA0QvKHeKVA3XkW3JElrwUrjYdddqrD45zRZswc1yPV4E8V7EGhbON94zc6IcdbmUq
WmO3+LLq+86LpzBsRTYT/1eXOddPDustDpFMU/7oHH8xz/DGrA93hYmAlkIfiVm45svfO6BpJPOx
uVUXR7kDV9coYsyR3p52jxdzTsPzH1zh8WQQHpz2SS/U4gf0nzX2/iiFXzmDqUZwZ+P1dBHfctuF
7UfE6MkKnXMy+71HVn5sho43ZIh7eogwS+FLYqhVPcZfanmtt6SxSHHBxwv/Sp7anlrXBY2T7jSF
qL23i7YxnWWNKFw4w/6Bzd2ntTIyadSDeuW/Crz4XkaVA1jl2EQpX1NWj1bUPkKS3TSaWH0alAKk
r6F746LAmxGNxUhTrJeI7idz1DElpkGhXDcbuevH4pquBWzHI1pL0iVdzK90Tf4emmPvOvzlPOj8
LrganTdQaufqO3Dyjv5Ryybf5s1gZIOqNdraaMuPhT2jVlZvDoGNetO/ZdyNN+etvAgHIPrB6ZGs
Kjmn3S4RxpbmoURVSG7LEdra4NdabSXZ9YLxC+T5q3bvqkJMw2E1gxYZo5uVYar/kCbZOe0WuTE4
zupuQKHX0M/L9INopKAMkesLPry+XIM9Whq+5Yc1jonSwbaopHXKogw6t9jjwuMdWVDBhBTXq9eM
sD6pig/4pRx0T0TgRl1rwmDw36ZLYcHMnrDOSoxYgIdRJPFBhNP5utaBVxmgOUL8awTg3TVoIsr6
MIBLZhYwGhLObqqe/dReo4vjfEW6tQbIg+jdF2BdSIIJj4NtCFU6boAyc90k8RDL3rlKU2/EyDlh
hfG8JsckbapQtfPaiF5rcsmzwlzHdTO7bOcQDWq21kV72PGk0k5V7llqFH0ro1A6+wIyuou+OEQ1
mzDexXlJuOBSqZ22by4I9JBAfLl/SmuzROGyC3RokytfGqaHrakNQBdNq6XyWZXiipfCeA3BpBaw
aITQpXzufnPblyIZQi7EgDIjm6FvMNjvrZ0vPU0yYsUrZqKAjEcfoXvVEOGX+xfWGZ2prTsPdA3K
DUNDTFEBuFvSL6N4ybyEAhWq0m+cppOnniNOiiigvjw5i+sTgMsPw5S9tSJgkiMXl4pPKs2r0dhN
rdIXKrGQnpmrSJwlSV7NfLFc1wOJl2giACCUcD2wRnrqpDf24Xb4vKpoF7JgQ4Gg+jQVF3YlDlbB
5LH3Ix730y57qw+SutLTUfIw9tFn72RYqB8jp+FS0DNyH28rukL78L01i04zMl34iurmHU0+8HCh
KH8/DrLCvPc4Dwt3kK07i9rVWt+0wsxiryMa5lWn+trE5rfjOkc5qpZYBLVMTlw7YuBbvQtgcJAM
yCZ/DRtqe10W9s16Uj86w2sPEoE+fIbzw1aAK3Y6jqn7JaDWo8XbaOC2KwSbyESb1IzqnJ3y5Aju
2Yl2Sel4rn/XsNg2yfIG6D1Ra8JB/iSxn/0ZLpIPqx3rWovfbyxlH7P6bGSdm04c/JrTvQa0hpan
zEfMjes8Ls8IdbOyQMmqAUjOP6KsOBN7wKr4lvm1RxLEF0WpEf4NIzOE254foEtAiamYzZ67cXPV
4wSXv4hHGhzIU9E3L0QFjn2Si+r/7goAg5gmmb6UaEHwjxyBtT22mLNQKa2iSc2EhRDDhcbECu00
Cfva5CLqnWAwruLQo7bTKS+EfsSTJJxh5hppEZEBySYRA1y7tS0dCnvUlyuG3/yN88Cgo5DSbUXZ
+48193HkuDA3QG7m1v71pDd99o1YJPs/jlVbhR1Qg6hBnkwzClysING7B04kTAoM+v5gYBaTB0Jm
VS3JOW5CAT1NrbHqfYrdKn6mEI4m+GgYpUkjb1tJEgJAmCXc8nWgp2t3T3wtC2iyJCAd+FMcCVI/
zrKsmHf9PnyEUKy8ek3Lm2iVUXOxwB3K7YXoCYCaIxeHyreks3nc0DjSxcu1WG5UXF32VUozZn/F
RFNNyyKu7tYe9YrFTyB3atPFgxBun50K7OWHaKpxrR/uYg8O1vLOJ2pNSKastQ43taiiGYhvk22k
fKWW9byMQzLJyoGV/I3hWEmm4wQ9qysnv9GhDiqoOul3JKqtBsnMdYLgIB+FfaQnk4z7f5zJb9sO
XlwI9cxLWjHMI+SEKOr5amFTU1h4h5aLxj5H87xRg8OVphMudA0dn5ULLo1M9FWl5WjgsJErcY1v
10puyDLlGdl8ChcshJjri0ZzszgzmGxafEKrXgYtnOgq1UojN8ii/zxGB7dD7SxcHTmWsJMHdKhh
LhsgjbscGibMI+7nmA+4SAuB2acmZbeNlWIvn5bLdAcK1Dny53T6Pw8tvhCQ+3ciMD7ri26DwBFj
V4A0o1TRNN1g0B1S0xd+nr1LIxSERvZACoQrNF+Aj3BY/xzUNFTetCysp8yLWysUNBNTjjU+sm22
Jrc0Ct52JCGe/fq+KfTBo5UhATl1isAVcYdC77QKKrnxad2XALkpN5gTPX777VbMGGkHWWqTea/8
5YkyWPxlFc7TfBuXfeFtMaiv+VRxtWNyzE5WMLaKOgLFcwLrcYzOpcZ5JO+dv31s+APaPphC1Zmt
u2R9UF6iHMze3rOXzHOnYMFQs9SJn26jogyQtmF3HjK0QupJGAJyIe7ZUE+x/sT8/74pLFejEyee
wSvhMF82kAHdOFy2ynMuwD9jpA9cNBFYHhx9T/UPIB6J1R/DeQe4yxRd+bGk8j6uNOcsl+bl4Oor
16/Kh58HEWh9nePOjZfwcwza0uMRScvZmPLRIQxag3siw0Rakr6DsrRWMnRPh8Xy6pKA1i1P34Kl
s3OP4FX2Zk8P+J3lOa8PgCAfSgfprr1dhsIIvUThHUwOzYTtDhD3YoeF7b25X+woFsRshwLPBcbn
CQ/+wQh914rh6shbtDuSOaaZJbZLTbv25rDWgcbunvv3zVssvnTyxvrLxSjpRmAUMIE7R/zZRQNt
HshWsopv5w+QCCxHGntfUEtca2dh7/i1E36KIy+6xINe3RH9BoFD6rUYYsw7fD4Ls/uHqgGOZBAw
7lFl7g3+EHM7PKrw6N3bOUYDVOBnifImjwZaxTGfZG1nZjVReceC8tlpVfMOCjwUpha+5MdUUBSP
aEbyn9sGYWDi6Sdo91TvlPPEz+sqloB6rOO/qO5tH31HVdvt7Gj43C5CLKpFwv1GMU5bNOC+uNwD
9hrS0l7ywQmP9k5Edt3cHZ6ZEVFnUtcJMykS7M/Qqs0FCRmHB7mKKt5EYM5Op/2/Nm6OV2uaIrrh
eQD2AkHPBlDGOPH0eadrWE/a7lpYN3hyjTXkHKrwTBJkk7enED04mwcq/crn0D3hMpC0l4PcLfjY
hyih5YdHxqx/96eQJEtTSp3fdfr1G8uHRBrvZHluPBJHeS6jkEO1ip3C1Q6sw8n6ony+oZqHY8QH
tcB1IayWVHc/MVcpP0ExyTby18xWwFEB628g7JvEYNPsPkRkAJqWAZ39qZTTjV1QyS1YiKzBhs6V
ji5pcZx7Y4AGr37eccR0kZUZvbqfxBesNsnqUe+gXG7tNSXKFgAawY/2WnRhIQjeBb+UUHtGYMGl
HWdrq/h9VzHBiagQh/ff/TmMyx7blt3X/7N56Szcyijbff45Puh4+kNfDRmi2PqgXZPWYP6zzNEP
gWxrMYQI0PyP48D7hQTFKazs8gb/NR/nNDoqRDtu2CPYNdE7+aXpLu0CgP2hFyvYZFfdmxx5rhsR
4INfZL5P2fNrt4WZEKLQY9pJZfrfHzVo55ZInSGV8k/v5FDmltfpEoY2KH+VhDHd6MILLftqJsPq
zcRDwd0PuH5+judevqwZPbE63raa2XIhlLyldlhg4g/DadAhh3F5fO6lTLIOVPBLDyGVqVrGorWZ
oe7cO0kw4Q4nNlWkOZa2Q/wktwFa507XdtAcZY8k35KTiHJ8K5o4wfilUbczotBOKwdXcf5Qf1x1
6K44W1Q3rUgeoY2siqHEte7anZGWbaTHnWcBoXsW9wMY3FvlTJjPO+sE9kl2QCNwCBtcfj6+5yKb
SQGlUBQ8Fd1vY3q4eVJKNQeAfGXA/zTNwyg90pZ05zEXA6Yigx2uM8XCcWn60DaYCOGqh6bZm9Ha
FxQzIGHtHUmM0xPxc8Bw+EG/lJIZNuLZgU4WNXVDQhBtYBlYMYZwFOKQQf0CE83z5gPx3Xj4oQY+
j+77QDJCJW9xDO+pHTMKu21TmCz0fOvxuubykdrG1yWGPwpwGOCXpNLavgShS2DQopL345kB9Bcz
eT4d4eQHuvvaRO3TqTTQ3tdlOy6hdCgLlk8cPqcCnko7NgBtcWn0HAt8ppMC2Wq3OJXWMaOfq2uY
hdBnTFsZLmY6uvuRSZZLf/6ox8qrgQj7rivxy3CoD9Hfd6VMV83Vp7sLgk4Jq5/h0hp1xV05QU//
BCwLvfSSQ+xLqOgwLTK/J1JSfJyp9XxAHqxWObQkNX+QmPrp4mE1xiyB+ibXHQctgWBVQ5q1sLdG
BMZAeRAQOT54+gynUvbQI6Evpb66JVmePUbi07t08qKYnBl0TM3qregWXxYQg314ycG8uJSw0CC3
fhKVDak70TAL2+Rjugk/ozdKBBEmA7ntEfn0Tjva1sSc2nHB12CFz1czwgPTg0L8As8HR3IxfCNH
pU0CmAzU4gfO7MgEUFoq/X4wc1jC9xhOIqB2joDCI6OAKF0V2IziYI6X5i7UpMU7GbH+g/PjNgb2
+rU0f1yb8ER7sh59F6WUfp//3l7qYfk+PFx2FlDn3Fo/qkcpbtjU1c7C0IAvkxLsQ7Wml5MjHOnF
86Lobx0BIt4TIoVnD0v0E6YfyhJfdeQ+7G7Fv1dL6y7R3+0JSOmD08acNfYBgYC+vaCfCuQgj5Mp
ngyvgEWhOdw82iZss1piYxAdKMRMsl7fqr43odSHMqgpAdVunfBA5yq19oTJGKoCM4AaUwdfbz9i
Sn2RQgEMthDrqpd5ORp6QZ1KLK1kz1k6zoA+r/I5JmbFl1AlNza+mglFxDZDeRBh05oZVnhdzkov
lzcvEXwCTQ7eL13jMnS22KcRrqcIYfmpleKg6UMtaAYELqNGGVbYHfNX3zfAk9gD7VIkFjki7kpY
OOyzWSefu4i9vc9wnVgSqcunhCRyhkAg9pnQ6HYA1Xq/2Ie9r5taoranh50NG1zREUeM+KqkCQCS
lKmCyUZ/wxL8mGoaT7VfaLnbayljMwo9XZxPg8L5LwttKbUSyToE59iB+JoOFdNibf1gzWdu3to8
rfd6UNUYYXxPDPaviWBfOV0FSaJKHBUyXOOR6eSXaPVmkQfXCFTamF9imo8GcbEzB/4jPr+j98qP
iL/auB+LwENrPGyHu9MrlBC3lEOZ8NSXuaVrImKqwXlYWWurJozRild/rzW8RU/bKTvGkR/dmEKL
KtiCnNuws6T9413KTOPL3ojw6ElkOeSMwJ+Afr0ZNN4T1sre6sH1oXaD43S5hsR6GUx/B4GsQCaK
qGvtW0ZAg9dpjtX3RBqvW99G5cY8YPcqPP5JEtxLHuYrYsQfzrIV3AMWsPiFWTJhOOxMUVwMXneK
tQvfjcZdvSAqxbeOnRJpG+renfwEVeCoAi2FlTLC0R8zyjDkbA3lTHmlNiOofEorxEb+bGNdKjnY
T27QGhHxYb7Bkh/qdxV4S6kXKmZUm07XJOmb6HflTnNFYjGMbQ9cNfOhyyAuqSVBz2uTrrApA1rK
l8FeNFapkaEOUCPtm5BFXxNoZRxuhn2caC0Uk/J93Ss3QgkvauDSgQ3Qd6S2SJ2tUaZBhLn4Vcfg
+0c2gLs37iWWfCMFPUmt/9m0BAk9jOPdDReG5c4wulrt8O76551lauEetFkuYU1iZLx/UNaBtQu/
1H4qAv28ft7Y8+tLm1bSX01HrdAdjEkmOljQsxCR9puW41lnhoDTcpUpcyyp8qH/r92XosCaYqZV
3sC0R7IZ1Q5zLCfYZd3Ag9pWvZT2D3w3QkTfMRz/lPFX+30BwK8Fjx0C3hSrwuYqYvPU903G1HBl
P/NpxV9T7VUDP2Gme5jfABeTi8fk5ZFSYn8b9e/gaq+lXtQV2DBAqdyXc4lL0yTKEA2Y1NK4GdoW
FHgU8KS/r+9ORt4j5s2ZN+ta2eJcxO0/F+IRtk3cZlSwKJ5t6VYjoO3NqIVbv9zxUOmqgvFHS/CP
5Xoo0lfFk6Q8/3VOkCR3FDSce2RCBn6MLJ8pD/1ILSPXEdeyAYVP8Kw4EaecLVYebWuLVPWli1Ez
Eobn64OLjEMTV0ybppLaYsh7EpWy6lo6ln8dClKf7+OIfYNzIHvDIfuBvr6Qvm6IUxuv1BgWQoT+
6HQ/n/R2JKEskW5AnbawaMKdgq6FlG6nceO7xY25AM03XR/BioFi9FIEE8x9dY/OGAM+Yr0/1wd9
RY2V2j/FhCaZ5+dHu5z6KDh1iQR84ft620gjBMXEsvmbdDzxfvUxR08zFdhb9Gv06c7npW3DKf3r
ObMKsPVhskIg+Br8rIN7uhJHTAqGwouP8h6hcEi3pyLME0zQy9qK57e0kB7uURxk2PLqlGqWeucR
XCzyTQwtGAI6jGosAb/E6ahscj5TChQTK98VCf0PGJd2ubbav0CY7Sdyqv3QVSkx16PliWD7GRel
aJDSNURD/MsEo1ZbZfvCznd+YRqGGes0BMy5Wr9qrweAVzIxSPp/98jwiBdYJMhLpFCRHFMofarE
7DdEVV26axuYDCj5pbt6pfeLF11zJO/G/b/ITdUHK+z2IiF14edF/aYu0yCVNnEsd1vCLZeU7EgH
pgQcRqNv5sIMUznEpQUAGwsYVwCBUjb329jB2KrbKq8oISPhPalxLjLRv3zqZKWZl/veYBlmsjtC
VZkMhd/N5CKdxClF7bHxbCN6ngNIcK7cewKfkgTVkvDe4rcuUh+bVOWVejgdFkuYstiJK3RLLpuK
8mPxOES1Bsa21JMY0b8qwStA09acGjo6vkuMOwncaYj9a4mYc4r0t4oMVwtOvtYuxtKYmYzNMoBK
vjvIyrrpAdYbIWr+ttGBZbPqa1MOLIy9BAFlhT9IdpZ7yV7rglRRvqkNFpTNeQsMZTyhDtFy5tAk
q3A9hH8MM81o0QLw3iOldNoM3ywUtEp8c0R1z3ynV3pzhoeJDWL7kDa6zNTpsZiO1OpHU6Lm/rsx
k+dotaRRK1MAe741oxpW3guMAZYuEzKn35wLC3V7zWtbzzVZPb2VhqUhYEqj9+vm6lWUDXlmErbf
NihtsZr0gmYS/qs6gEbwdyqblmF5pyiwlI8bY97etvBdgyfz34R06yknlSiUqtTHAJ9E9OQ+5u3f
wTi8fViuweZ68NOYmBqDbKZuIOTZwI5lMIib0LH7TE4jriS6PHi/DlSmKldeF7KlodaERAjCTMO5
qP4lPfOlQhMZzO8QLNuR0m0JA3xmJ/vaug42BAks2SO2OsZTNkmArWGaU90V+Wei0u5+yoX9SnOx
H4Sp496zI9wcd4JgTlqyiblqLEC7nzbH/Z2z2CPc86ZOFl1zQ6/Gg/OFj+gT3s/CgLQzUiJw4t0o
6yifpc1uai/CTBO6F8jPF+SnzZOwU/Z8d/jRJQI0TQd3ARR7EQYyapXU9krWwUOIxDdEvC8fbee1
/T8+7duqTra8cRVXKJBDJLzTQiAMkFDPawdvpm60/NCrrl1ImNKovONiW5tBJfCSb5sV4x5JnakC
8RrnFCbD/Ytoet09Y3iKTNmnW5d9qqspmCDyYi/ZaAWFlwNrsKt0L6A8aTSpY/ZnA8JbmrjkcEYc
8sH9t99pWs9Z5H+HEe/RXzhSUJ7+T8foXA0QoAMg6py32yAfVW4rsWkZ9dGM/y3CZw2puOoFjyc6
nJfxhV9o0dfPZv0xkYe3dpXkJXoXJw4yPeGX34B+mc6tB2kdkZGhK6QA7LTq0Ubbb7oD97zD9WjN
Wr13b49WX/l7pLT5GtdWVWyC9XGVRn/Z5CJAIxLA4KfGY4zgu6ol54BA8w+/2A50P8P3o9vkPB5n
zPNIIgfjaN3RUMaHAW4zbtWQoVrb6uz9zLwkj+lQsQzgoMQhcfM0qgG79YobC68FgQ0b4UeHuUQF
q8zR8FkKDj01ul7ZvGyivPUmBbnxMnfG4AMilhwn9Pa7P+kprsl2XlYs8xbgEFhUIMPm/pDeHPTG
wNRpAJlBBAA5UCB7MMAFwvmwPyKRvnkxWK93Gpgnp1UYBSDSTTclDdcV31+O/S3CTbKGCXGudVZb
EDn0EyRdIDgp9siFJF/oR50Nc4U6zRTmFRWxC4KCSO08/9HtkUE/9/vqLv76cd9NTolwNwa0RZJ7
ZG4wtOD2mE26YHKgJNHcQhNQc7KnTRMQDsdlWff12g/+0xConwEIFAfhazObrsbe9RVbJC5sAiI4
MqwPxo5SVSFyUX33lfcVL1NiVVx5fC6FnWGdXMy0Sd2mfy/axsUZti7SbxKX/exkMn6ELyj7dpy0
jMbvNVqDT3wYnsIkI7LugIgrXRgz8KD0gbgxLD2mgJbd2eX48pEzHpdM8WS/m3nQrq5r/ZsHGzLK
yuoxH/gXZscTC1L6ML2QTt5LdoAjbD6OGe3XXYbOSfa6Lt70pwFpSvws8OosLpMH76is4f8QIPxi
tEfOuI9Tp+bVwgsDxlWK7QpY7Z4kEFGYYYpxKmvezEWw+7sQsPyVHkcytaRUGdJ3MFEkjKlPVHFL
ZIbpOTzADPimu4AgGkzgPY0b+HxyNFB6YsAN8ieZrZPIqjtAWZYo1FWc46yG3XjpL8CylGvvgo+y
8evViTeoeGlXc1HR9uMdThh8JBKRJHncbG/B07r/JOsO10g/0mZM+pn7wZdqjG4E0Edo7K3AcbcT
u291lQSUCAMcxJQT+BbpXHkZkYevDfi7OQWV6Euy0FAiEBlrk0TK+Wps8a6miXWuOioguOkWGXQh
h/h7aQ1sG+aEbcafgpnh/GFaMpBflWYYa2g0Rm2IeSapxRocONeA8qHDQjQkg/6CCv/2i0p3v24c
uaOXKyleWf0+DnfSD3jDnadCRtuVAMZCAAdqLPNrNG8aDMOURfrSe/FkQymP63ex2RjwrdtUqHPV
/JLI3iaTOc/tB4BhXQs6stUYm/HYsew3pBMFOEWASE4Io7WJNLTWHoTMvhX9KCO25J6EaHSZwNyT
6HSVTozdMGC5jOdq4b3il31Iqnfo4ktEbFkC8dRb2Y3vKKcdNKZ9jhasjI5WKfwzr1bYcUXW9h+X
SMWMpdfgA3HSM5KCbT79TV/VihLdw59F1UVcntjFjnND7XE7wThdCAo8YImXzLJ3x/ajQWD0n8kI
msKkzv6gi2185cv5GzUyl6LnRWhSNivhtmI3aBZIEyF5r6KgrDU0kVaZoK7+LMz6xyLpQTBVqIuq
3Cqn0BxSsu6IomYlJQ9ZhHof4LCbZwvCIIBeqJu0cXQU97njwBXpiQ8rcyUQV8zWKf/gaqkmoA2Z
qehAu2OH4mq7Z9cn0B/UqOMqJ0UNnpcoQlDiMP++2rGjHEIV6wPvjccj3zXt9+4F7A3DeYQUvU4m
W0yuZm9iDjD9vPxpThVTjJ0ar0xm6JowVxfC29nyB8DK2yfDa4ZprJxxnLtHBbU3Eg9a676IAdJJ
Ydiz4zrtxz8ukxiyDQ4vb14JylnEl3tERITVfp3umvl4OLWMhivsKC1KISQud/vZCd0L5mpDCadC
TD8XX/fTf8Xzuqfsp4ek795pDFvSJ907ZUNQvHYfkTUsa/nKlVPo9ileuPWTMkpMBsATcuzJCO8j
CGmWrFaibxAcRXK+7dkWvP2bYXMLKz+JPazSjS2oztgZnm1gLcpWVNzflHm+WS3Fp+fJ4F5yf3v9
SO5jluRhaxFMVe3JHBNzw5h1SwzBYX23v0RV0kbsYKG7nyLLC8qXFyuqmrSC9AQ9IrzifvDeK+Cu
uvwGvNyn1HuYyhvaVfanePpFn0rYkUR+l9nsxYKyXDzG8aJ6mPexTEGeNQ/9h++9wof0UySSfGtL
mUQfv67KdcxndMkwa19+F3caRtGePb59fb1ea8ndHMJasBJU6bxYtPGgTDd/gPoMR+LbVCY+w54E
SbTc/QKxPvpNl4teZdgZKJXhcvFCjtQdbRhNs7Ogia3CV1itgz6IvZOAdKtvvL0PaHuFn+EaeZ1h
413F27N+wPX29sRCn2DVDHh/DGd8AklYaD7kd0VvHyYF74h8U+PNdq6rTRb2mFhRz/AdTrLEagG5
GJ5kr6HPss4KVWzxyvu17MKIzvWzt+KrmMkVlgKl4qJrcIAJ5QHpURqwl+9Esv7xUDod62YgmrdD
7BpM1wn45qacRqx+tIj+02WIB+i3YFMFPtphu0tVjeJYwCw1Z9JzmJT2yXw2c/b+Zzipwr5OrcFQ
Q9SKRELxI9N8FzceZhNlWURBfY0cMtucxcX7194VhKNHqxaSgo7y2L1XZyWaiJv432IyjPOXc8Tp
BE5DfdLtMH3Wklj9oJiE9GxttGO+bh2eWSHag4+y46vQZK45wyBwouJeCq4AE/+kKWrQ0ecbP7KS
6JwvfpKGoSou6mLPwxO3V4s/i78Ix7L0G6Ghj2Szhz2FVmwyyUPNRcWtSv2jIPDm6c5UXp0AvfFt
LhHv9Chs8+d4loobUSsUMdU0GSv4v4Mv5M1xd31bl2E59UVUKlzfzbBX/oLqjAvQ52SplRQsiox6
XBxK64h+vGr/AtDr1NY1SnFonv2KutEGlBPaHdIr5gSRT6hii2DKSVupERZyvRV8PfW5HY/gO8qs
ZuX42KUpMUAfP7bbO2zYHdmHKijoXM/Y5F6jU+8Lubf3J3PhvvBdvw8LkuDdNJ2St9gA/FojDZA6
p1eLzWFXIUJOnHHmmyWRSySA1gX4W1p9KfVPJqbDThYBrBbfY6BOZjqCaIy3JUZ7JCkwecEZ/Xcd
zFtZVqOD2oPezv9E9bMJ0IkqnV2HbofXQ8lchIv++bNmDvsNKTrDnCX7qcZ+PQXgmnRr0rwCKvBn
jLooGLdqeheothtIawciG/vBhiWSoTVswZpe5XqEx8otlzhUuIj/DBgbkEj463Dr4PrcL/17birg
E702xbuEqGklNui43stdfPg3Z1IRwAKOPoBRtFkBS7yzHTcMR46eiDZeIHXnncD9X2fmjWcSQ5O5
pdooiEgBy4gImQVi1v/h6gczOvZXJhniijlGQt2QKUqzpq3QQTUm21eMvjLotsTFGoMoxbojqtIY
XTdRIT4FofNafc6YEk8RiyDwgIGwWs1SVmQvES5esy97tWTJmYOKK5L3bisLWZjRHWBPxb6ZR65i
CmmBKXuHs0PfMsAX81AFDWxEAIhAhWOXfVcrF0E9kQSs+Ld04hTmjAuisQKdTzjwvzIQHTfuu9dc
M0f31Ay7NrD6AYo7QoE5A8txbm9p7Ht2g/5bcLuZLKigGlmHfYRWjh2u3eD7Y8nQocGphy+RqZUV
RB8eZpQ8WYS/1Clzy4irEkzRNfIC3qMM5XxHkGWo0hsO0NYqPaHok+mCnlFNwpzaFB1MTwaZhC9Q
oeXzdmhaDHOcTl42C7D6T28bk8uvaw3+CUH3pc1foFgVsF2NKAW1jPPgIbeNlN8cCGuKJyQ/K0AQ
4d6uvD+jJF5qjjyfNXV95Kt4GOLKSi2WOIB+2bWsqaKgmsEJNGUcddZ2Mzpd9l4QDv/yFAdQGnRy
dL8y2rtBtXoGIVYPU0aBQKJM627lKXsLfM/iEkYZht1MD0GNt/i8W9nZ4K965Mc/GV3oz6ZNamVs
bw7l1VTwSE3HF9FMY2LH6nPQ/msIOi596niRnQV5Yd1rpowhJ2Y8EhrfQSFWE+5u4/+xipNxDhHQ
6BQlnvcAZD6ZY/gAipxq92Cj+PvJBoNu1yn3mO7KoeiNw2w3R2D/1+40i0ujx5wtXyW0S5h1d1xc
no+kyaUUC9FLa+GA7MDFos5PQU/KE7pVcBVht75mHPNkJ2wwaRoZNT+bV8rFQmeev2ntPs8jW328
uxsK2uszvEypRYEwhE0EetikXM/eb3w4TIDsPIuI+c48v2hGTWU+sOqrpY65TYlNHRRAUwIDl9qo
kQeLdagRAG/xjccVziSkxGuairbqOktIr7Qj6loMzoXqs4iYMtku9MSScq9yZHDtjnLbPxiSMdSV
uHMnD9jHeoLodar4mMB3cwNf7YkhOx0+tWmijgL1alsHBfktwZLBOJIsUr3pK124qWWgAp8EfHbx
uxIEkmg9ZD7Wr4qxZM7KMxb3ffKljtQ8BIlFB7MkxtoWaR63AOoMl//X477V2rStwL344RXrGFc/
4LyyLMUfUNJp4/kJRqeMpqY/MDISsF0cxKHr4Oqd3tbtrcloUJpKhPYCd+aQGcvNc67YvuBf+0ZR
8inh7FlVyR2EMMG4QZcpUI/Y0Wv9inJQW3VOx2Q90jUBv+JD9YldnwXY5pddnaZv9QKAHy4o2y8s
qrcroKzCyMjsgXywboQy5gUBGsCKJ/haPkmTm1AK5Bh2JVySevzatf3F8g2+FdSxlbH/8hcOStmo
Ud9gsNXhcbvTse6cRsDGxMcERsu6U9UeMKTLgtFv78d33KOg0yJpcia6GTHiPMJ49icXjZFTLJDl
EEcwlq39RKD1OeKHNSEK8TvvTiR4aIfRX8MujH8ZoockUdBPyqt1s/GLMk0gtgjHZJ7bxGCeMGtw
ytxUMk5oOTkETtPrN1NfAyh5Uk6D9Zp+me5vrLCZ9vAVhuX2ZBaYz85A59bFgwQDej2noqGQXNdD
VX+hTVsjLQu6R3fmC/YChIKgUW4Hl8gpU0pG6j4rfaVhlFIQt9iDi71fG4l7hER+f1i4UGUaxRKM
3kXHW1+PbAi6sQ6oujAfL/o8FLbymrZPxWFLArZADB2pQd5yVtD2pzjnvG28Upa6F51PA61Y8PkE
wKD0bHR9cq4irsy602rdt3Hcqydp7DdCNEhStMlIMsjpInRCuBDMqXjA8imGil2pUuQep3ZqmwDB
Rcijlgk8KpmjT1bVscfEKaibg6x+mHr4N+GqskRHRAbp24ZWonrwzMSKg943XGrhIZMHkCvH8lCa
QauG80HI8FSud09Ij3L+G5ZVz7/5YYCob+0Axcn0UOPjf4FskRwIMpvQM4Xbeqm7TZVQn61zcEqw
UQSlj71pHdH+E0fX3czNeovM29HKXoxfwlxvipHW88n+x6cSarC1uF+7J2xM4RpJiRpr7S4Gy9J0
OQxBuBlN29L3bkyqvg1LP2BVjRfA6gnHpmo0yhdp2cLNkRXVCvW5p+h84bK/NqFs1y/YGsS9U7Cr
hHnigAIK+Z7XDv6RqT8WbeaCtD/d9lf2Vv8LbHbCW9IHmHP02qOohOkR0c4VKFDsn/fkVeiTnmkg
pTEL+BJx8V3ndgY8xY2KnqsHjpalUPToMciz7Tmi+yMW/Caqt7DMJmfVvUCdFH8V9UaHULgBvAET
aaCccwZLi3nxUfccUTEtF4794V9G4jRGkWyQmcxw3naDwkATb0b0RLiKbW/1ynMoZ+4H2KD3JxmH
Na0KEBCNpmEG1Xlm1B1z6IBIkSUt16rNzbYdVoGz6SsKUc0x/vzwmLX5+hGca+CDiNTDlOnLl4g+
0iq3VVTKKuZuNj1ect6JgejRWjTKTmX4yqC1i3cscc/Uw7ImT3Jj439lhcTmIRLrWgBxTwS4j8x0
7eC2xIFrUqsUajLhMjOgfkCjKlpSR3LFNE2V/CVIaHQbr8JPsdOwof3jL8W4ch7qNbBv6whtPvSW
T8cnzxxqTeUnJVMms6k3wwaRet5+VaFpUCZGg1P+Dglqgoch/rk+kOKvLzOzkzLab/GWmm+IxB4G
QZPurS9vNWUmDZMHn7DJhmzg586e5KCLwvc4zQqBGOsXUhjFFnhC3mJ7hOdXQofwfGTWVFuh+HfI
yRR4d7dZp28hlrXYMy2SOO9UXSoKVbMBKNb8OX3ZaWapr7SgZ9ZjtOSlNdfooZolrAOsj7FEX2he
DAjgZuyf7X1apkOctdYNyBEZo3a0K+0A4ReIhpUAhQO+PIsufY8zJYyBlcMgbvs6+NHQ2oVgktaz
g1gnT5wwd2RN3EgTT7HaAAm5l8gAEWJeKOArmvjwdIcS+nZbl8+Gk4JwhM1OGUFrsPu5Tk3qheK6
8+gBHF4GIB546WBgEJ9J11BebAELUsFBozg231AGpE0dtMtTBFzab/eIkMNnuw1RvOe46hxuWGJ9
wQOiBdp6h99qPWny+rxd7YYSTcab/DaByV2i6dXNLv3VcRM8rKeA327KJfffr48jm0PetEv4I9be
U43T7wJdAV1aOoc2fTxAs2+ZLcWQ/Od7QNuahk83ihRFaVdLoKVAWxZltqzusm2PJRIlvEKR2fW9
7d+wGOn1bbaww3a+dyhjDA9Tt/BcJzidIu7Rli++wAgJwJj2kj7jYf2ZWFjiZEHj2delh4s/3Rzq
BALTMhh7S4uF1Pw8+rweRLyb/LBIlLUAv+pkaLObvp8lzsJOm/2D61ovih+d8SiTMfUoLTzpyWnK
LBi7mYS9CbiKHYayI/fwvVz1YinBPk9/5YZt3fHhe455XNjGGAkhsq7PHKxaGlXOGVxcuY0R5tHz
OxthNYLMP+xdGbARqx4fuZQXMTs5hDsWa4fWKYI+Fc7omFYKf4RDFDVL1Sn2+4YLqsOc6e/bi39B
KLE6ZGADVJ4SWRvKcg/zRT3CMb/kRHr0dnMPQ6C0TRS5+wfZdJ0I54mWmbOyPcmvrLi9pn6zqReK
D8A8W0nBPiHHCddxSg3WQw2fOhVG+jeaCOYe71CilNT/cQ==
`protect end_protected
