��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$Rx�y�<��wA�*;�x���@�̦�W�X�fa�M-$u����n~�%���P�$��W��kYَ���P7�?UMfT��q�6�U��k�>����~�\N�(�����X�e���/6U|)�X2pF�]$h���d.���9E�g�����	bI�g��ȆDE<�篙qU��ٙ�����`�>��
p��Lż�u� �V�s�{E����E�E�wi��(���T�ǿt���܌����Wv��jՌJAI����6ã�I�A��0R=���Sg��CO���Q[ҬU��2eh)v�u�JL�P�;���0ڵ��}�{��� nYd�K3,��  ��m=?@ჵ`���XG5�w�?�p�y�u5�)�4�o�'� ��/�z���:1��p�o���:�]6^����c/!~����V De���@<I�mƮ؃�hj��t��7Q��N\�t������wG�O�W�x�U�����<|/`��b+�8�էr�c��~}�8�n �#�Z�I1�I��르�f�L<ъ� ����?vcn��#{,{���u���1�W�ִ5�-C䒫��d��<*&�(~�]{��_8�D��?-������������^s$�cp�]]�"�f�Vr�RM�4<��D���t�N\=S���i�<��K5(ʂI��z��~I�%��#f/@��o�F��_9��t7�,@��̗�(�Z�����$��;_�������>M�Wc�@i�M�K��2���ˇy�q���Bs�1T{��x~]!��BjD��X�^�y�#g�5��'Y�YͲR��&�R^�hQ2��Y�	�M@{h����U�|QⳄ���)X
�Lg�����w�σ@���0�A>��̌)=Q��� C�h���Ѳ�r�Bn�U\� D.��u�[����+�h]��9��^�s��~l/�Ԫ���D~�K#�$ͯ�BHt����wH���6	�Q2RB����r("F�� +΃���6�6WҎ�Y�7n�5�V^Uu}�|˪�(~�Th��ņ<����!Cy�N�h\�3!���?��w�=L�3Y�'��)�̬J��s��H	�"�B���!j ��!��~��Ͻ���Ӡ5ߥ_�W�^�1��&�t��$��X��+��1�@�vH1�h���]��A�w?�O41�P���8�ޢt���/�U<D	U-hIZR�vGs��Fkj*�����u��=t� \�h�P"�5����B�i	����l�ߴ��=�w�u�P�t��$�q��8x\��qB_{����͓��B� /�p�|+C)�WX��I��K��5�:�\jr=�foE<�����3�lǃ{	U��C���=�;��A��6�)�Q�'$�B��io+�q[�3�b�Q�^!���f�D��� |��Ў�O3���i�ł0��$6�3�>�r�8*��d@lBJԭ�A�:p�����$BrU�U�,r������9�}�)qK�$��K]����v�HmD���u�U��T�@�����Z��&�['�G\fBC;a/OJ���{��nA8v�v�W<.�a����O�%:v�6SP��u�i�<&.���K�7;�1�݆d+��[V����'Jo������x��o
 -ɐ�c�r3l����M�r��	�f�]7�|��5 �#b��| ؈��?*⦅w1�1�*�2�����:nW&����Oz���Z3B�4H�h�޺E��bB��%�g%$�G��䢰�cy|�𠞟�J�}\+��;��9ߍWe��}I޸GvYM���X�D���(�y3�+_\tR�P��>1Xd+Uk����˝M{ִ�b
l�����/C�ي�5�P �u���n~ ����m�D��~�J�������VH�C�G6�fv�����q��Yi +Hmnw�'Pz4�C��[e->!{e#�U�Q�btZ�<��Z�p�:�,��Dl��~ lFm2����W���k���N����}Ζ�ehU7�t��z�A�_�v�*f|�~�f[8�	0זJō���X��µ���3Kb��{�*կ�Z��u����I���C4����'��(�
��������%Db��x ���b��p�-�|a&���>����k��W�^�br���5^�4#5�H�J�ޝ�;Ӑ��r���!��Q,������w`ُ.�D���(���V�D�J�)��m�?����6�y��	ཝ�eb�"�����YIELl�z���kI�U��U�/�f�~�I�4������od���Xķ�\�i��8-����Yy�߫'97/]��#PPIu��ܛ���Dp�,^?����̟�*�;�ZJ�[Ft���N����ܤԊҧy�rM��,H\o�i��i�uq��b�J��Sr.�������X�z�_�n��0��5����q��a����f\�: 9�S�[��l�vŘޯ)2ie����\�#�m5(�:�Ǭ�>��+iP�v/}]�H���f���1��3z6�fw��0���Ǒ�~6k��қG��ʂ��U^h��F��W��@��nK��){�Ղ|��V���N=�7B>RA]�� �'�D�����N
�~�,�|�Xl��zƦ/�&�<�;�
�&�Y�T���$B?��v3&�fSVX��D2ya�"�t'l���z��BE�J�=���%X�
г�_�z02R���R���Кo.E/�o�/�\�Q��c
^�
��������"G����f�ƻ�8�t��T"p���F�����a�F�<Bp2��Wz	{����\4�7��l'}����xw�Z��NG�X�R{ؒ���zӣ�"@�L8
%���J�K\c�fq��_%�	���!���^ׅn�t���l�i ti���h���qX���1N��۽\�󐄹����J�%�����^�4�/�	�`�ݲ��J��2C�[�ñϚS�La��_�9~�Ɉ�"!-rF���QP�R��g�O�a������"h��s+ȓWe�����p��ʎ�b��ʾ�9���q���(��OR�է���$bUFJL�y�@��Q�)��IT�7q��ݹ�ob�;���h?8L	L?��A��h�n}Z�戾J�N^�T���f�E2��o�n��9���{��Ke)bO�q#�I���fO��8YIԎN�ANEK�ԖY!Y��H��ݑ�no��S?\�ϗ�$Χ���eR!�[A�����r�����S��ة�\��6��q�F�T��\�3VxÅ�37�>a;W��?A��}zr�!����"�F�6/g��d7<p�$z9�=���!�T�ۚh@�#w
}ڋ?{���s�!��\7�1RCs v�[����=�2�|�X�БV�"W���?3����ĳ�|��&�5��{]H�߼�-�L�#s�$x���W�dz;��(I C��Ǧq�y�)۷E4�v���%s�\˴��|Cؾ�K�,����_h?y=42��y,Dռ��_lC��-+�~EY,�q~5�,���%�ꟳ\�	 O�SR�#�����\�t��J*~rL�cp�i������ߖ;`�h�����mrڜ�P�~sE-�z��-�>�g���S�]z��kt�cK�������AznZ�y�~-�]ʘxa?~��I˂������a��?��髯I����Xky�E��`	޾W��D:W����@�V�v����;>E�/D���
�G'��c��@��J/"�U#�!>�ܿ�O���Jt��nt����rM�O���)l��	�P��So^'n��JУ(1N����ZW��mZ��oD��͂a՚�3��F&R���K��Q|�_��FE�Tԗ��Q1�d[��l��(e?�52�#}E��v�Ŋw�^�*V��F�r�����@<>fpUq[��A���0����>.�("Cu���+�9k?�	_UՖ���Z�c��[xJ���h�t�U�h'J��.��~�;Ji�)K�� �
ȯ'��t�6���j�5�Oc-�D��]�-/�b�O1>�>/^�u�N����y7��-7�49DF�sG�R�L´�o����ԁɹ�o���s�!��̐O�Bv��7��pvT#�C��&+�xb�܎N�Ǔ�=c\L�o�i@)Y�ŀ�������5Ō党��P/R�g��h����Ì���FU>�@��;M��H�ao���w���m��K�L��+����)���[���,E�N�vT�&��"i�{��c���9
p�l�����'I5A�TCM'� >���R���+��lm\�u ������w�:������Yr`����0���H����vV���z�ر6�G�%�]�k�b�\Fo�!�C����qǐb9���v�1��/�U�#�]0�����ľ�?�x~�U-ؓ���a ���Ax@Z�w�
�9�R����فol�����ѢB}�œ&5�A��>r��}hR������<�Si�и�Kr�6���6܍�3<sb�^�-������h8���w�g$d�Cr�����li�NzQ��֨?�e���3k_���4�,J4�aa�[�Ar밅��scq��Qh5��E���8ϾG;40�7xC����q�	�n"��A>���fS��+�-PM;���'5r����,��J~�ow�(��b���׻tΧU�� ��_�z��P�BV�F>Π���,�5~�?�U +�m�]-K�s�"�`qޖ��R���q�&���d_����-�������A��&
�TpC$
V��^�@ $"N�>f��!�?D1x7mי-K�ڴ�����q�[��?��gI=���N^��ǆ�T���#�N}�G�0��6���eG�E��K_y�F,�v_#l��΃!!
ᴀ�s�t���R]a�U0P��`�cR[���J!���w�0*�R�M3Y�&,�Z�b1j��R�����ly�������YA�:���U)U8��=���ƫ�)M$��}��m�{���	)����3n����<�֐<*����{��D:�֗I���7J�u�k�@x�0?|}[�� v(D�\��$:[2�+�p(�m��w�������Lf8e�a���uI`9��B<"���Bx�W��q���.�as��M���NQ!l�n�)��}?b�Ӊ�q�/�ˮ��o�HO�I��"�T�ݏf��w�ڥ�063����A0\��L�
Ц���kF���-D�<���C���W�*�T�ŵ>)>c|���2��P�gv{�,E�A�?��n�ޢ�(H��ܧ���v�f�=�D�m��s8���\H��V��q�r�XV��*?�5�ٵ�Y\^�_�������9ZE�+hG���s���l�x����D�K�D{J&Z�Q?��U�yY��KЖKͥ�RV�K���{}�q}�LC9���B�yr�Lѡ2�HW���ۏ�
@�gQ_�����UH��m��
mxwi�p�^?�9d0�C��$I��ڻ�<�'��1��ĸjI�����)d[���c�+!�]����'J�tSei��ɼ���;���
J�а}�Z�6^iBWR4ا�v�(��(0�v-�w3B�Zӣ��sꘋ>����4�p��2�m�(�qI�-���Fv��5�6����K�2�[g��I�_��/��gqs�39��d��4m�զ�ܵ�ʩ���4#=[��h�k���FB�>p�jb��%7q��
y�~���u��|��y�Ԑ{騛�PY�8�j�)J%ǩ>�1���]!;{�����Fh�Woj�t{�'&'3��+��q&}�g&�yEނ0�(������%�?e����1Mv�a�f��͡]6��v�vZ_m��!���^-j�b���|�`�Bp��^_b��zL�-�yIG�&ı�F�qZ�v��c��B�̧��"XԳ���Q],$(�{{�Y�R�w��8�xi�/V5�A�i2h�t���,�s}���wt�tlf��q\^D0�����t�޺MS�����z������Ҩ�C���z�d(�¿WkZ�D��$vho��*�xf�Q �QU��0����	��-�(�)�
������,V�&��g[;�w����@�TDS�t�q�e&˴�G�3jih>��W��h��^�²y�{S���-F�F�
}|F<�ٛ��C^3N��C]?/u"ޅ0��R6:X8�K�МU����X���,�f��������
�YW�yL�[�Z��
7)�w��9i��1�ŋ�]���o��J:& gPko@����.�kU Y֢�y���p�m��%	1HCn�_��d�Me��N������XR���XH�=ɚ+?�-��%;��߯��(���� �IHG�c~�p��������1� W�4B���(X��9ަ�>:��D6}?)�����`�V��C�E�߯���=c�<S�ݶf��Y�b̽6/�n�ca�:9)�86�A{�	՛�ڲ��*C��ॢ�|��/������5�	�W:���ճ�\��H�c���ԸgV�_[��H�qS�_��Ϣ"[\$];F�2���������,Em󔆽���clk���}o�jȆ���ټv�#���A��'���������D9�Yʪ��-���l��Om�H!�$�;��mJ;2c���9U}H������M}�$�&-�����M%ȱ[̬��|��N��	�ь[�vpn�TP��Q���o��ֆ�����e`�:�� ��H
H��P�{�{'��g@݀A�Y��n<&^��#~���F����]FդVt�
�7x�t<��� i��6 ��pH+0�4iu��*Ml��y�֍�x�źw�w���A_�#�V��^8���8HeF���T�T]����rs�t�.Z`�a��G�\�2�6;��A[���]$Nq@k_�D��r&�Nպ�V��X��;KQTvӎ�����=�ڀ��">�����7W�F��``߀4��Jj#~�}��.����Fd=wp�}1�K�"���_�|t�#��5�@d~�S�	lm晾�>�����E�F����Չ[:����Uη�n8��{D��ͰnŌ�H�ZߡҴ�����3T�$Litc�d�d�����F�.��Q�����<lw�F�%΁N��3�θUq*��k��S�gO��Ԗݛc3�{p*����j��̝;Q��[SO�Ib=�E<?�5�-��Qv�sѓ�.s�oU#�����>���g^G��z"���U�7��y�s�=	zՋ�.x�U��lˈ/V4E�v��Z���&x�%i�y$S����i�goCts\~��'?�� �?��?ぅ�r�8�Z_��P��F��۾�����3�Ų���<�aB�;<m=t����߮a�T�w�ou:nx�­@�C�� �MNq���cb�d���w$��_�����fn��@(3=_z]E�X/����M�d(^�_�sZtt#�x��*�H�"8>05����_`C���sY��p�X�0L*e$��q� �,>���z���_=�-?%�An5��@񄒫h��D�1���G5����N�!�Ʈi�AM���~�"��@i3b�&xI\������^A\�Ut��T���#��޼�,h�!���#��=��B(甘ܸ��Kz��>�V��kS�hMl|�5e�sN`�(ح�cq�G�{ �!B��,��@� cAG:�7�m:��2*JʫY�*�~S��߂���g3�X "7Y�xrq�}�@�o��ظ�i��=�!I8�AE�g{VO�Q��Ge|�'��:$��Ѹ0G� �<��ad���r<�U|�J�u��3���Y�����!<܋Ǩ�k#0��)�T��Q��DWL��#AB1�#�6�kB��5��!��ޣ�h\׳�m4����i1�`*{���˪(�ĮO%W�CKE����� ���}�h"gE-�U6I��Y��T� ����{ۇ�%��r�1�F;
��DsD��e�Z�������H5CqJ�,�&�3$�9ac�w��E�Z�;�	4�>F��pI�?L�/���s6�#��")4��+9�Eb����g5��n�G��[�ӭ�|�4�;�?��`�I�48�}��5<2
1�}Ѣ2⩍]�$��7]l�D��ՍK���JSp�Y�q�CJo+-1����7�SZm]ӴՊ�?���@y/s��<m���
C��s�v���cE�i��}��������_d� ;SR:i���'�z ���WӭT���w����|UzC����RX1�x��� �}m?�Tm~{/c�*wDD>�y��tԃ��Gm�L�ܥ:3�Lc���i�Q6�ʿ�	����o��Ǚ��2�GP��lՕW�ܙ�����z�%����b+����΀x��5�ķN'�ß�0�S���]�>q^�HRk
���W����?nυ� �k�����?P$�1�u�]���Җ�j��?�o��,RI��#q0o�-WMH�������v	�,A�81坩��\G t��KȾ�͝�iC)�_�L9����Okk��;!��5\ڔve+��4����g�M:�v�j���������!z>�V<Ý��o����H�d��Ǵ�p�Y����\9��S?�d����~�Q M�#��群�
�A�@U��2Ա�-L����|�:�2..Ų�I>|8��*����K��,����q�7�I�bVTm��6�d�(S�??���5�:ٓ��!���TG�F[�	��>�.m9k�߷%����˳)��/�\�`�^��phJ�kx�M2��k�TP���1.��.�U�)�	hҘ,�wrv�\�w0���Y�����w�s�x���|s��qz���]R⫟Z*���Y˞��!�w��B��`���ߣ�\o|K��˸fpձ=�s��[HA�s��i�jd�3Ֆ�D`��g�@�>�k}�r�L���D��Wya��א��B�B�qF�P���"�ᠠ�r��M ����pQ��,����4n�m�Hw���y
���@��\6�s	�`v� W�C�II��p��[zgA�Ƚ��^�e@pp��P�M�3��.I�	�Y	z
C�e��8��hl�l����Ot���Vny^������)|��X�o����� ���aۆ��T����S,}�GP���\�,�W�3)�`����_Wto�:��	��;D$
��U�#zj��l���$q���i��U,걊}Շ�g	�}0�1+��x�[`�A�59��-�F9�l�ps-&�tE�9����Ў{X �[p����L��)��7"�����0�&y��<�����������W��_��ckP�Mkti�I�����'Nt ����(}qEU/�ܝ�'�m���Z�4UC�������\Q-�q���Jp�n������^�+��K�jb�Q6m�x����mW��F���a��`��ᶴ'x�}[�!dDq��ǁ�`t3������6��Ь��,�ݹ�XQ��J�(1���b�.���$<b� �JR��&��hL�^��W��nC���y�)��V�l;|�AK��(���?��6D,�D{�<u�,\CRW~��:��N�)���#H �d1��hAawau@�#i]:yX'{D;㭁�`Yŗ[���W�!p�tޤ+��nG��H��b�B�5�6d�Sm�~LmD<�Oe#,��_O;Q(2���at�.���Y��3��T!��	�>TZ�P�f��{��'Gg�PԔ�e����K_���2w��9�!g4��U�u���3֑�_Y���@y팯�3�#����B9�@���/xRψ�_��Tt�{��5X�~qC��JY�H�?&$�8w���;b��Hģh�	�j��}4̘�rlڂ��y�l�:�թv�f�L
��6(���~��TrO�EնӸ��\�U:,��b��l/%�/�PgȲoǭ���\���}�˘&6�]8��$=(�#+sp���<���v-���t�a��yPL�RC���H �Ct�(�T���A9��SF��$�%4�P�&�d�]��`���ĕ^��"��ii��\�����<��P��)�	�|�L&{��~�p�ۮR��Dۨ�7k(�#�"q HQ�Lv'�e�[��2	����8a�U�7c{JG"X��4�xu>����Ѻ�w�N���V���촰|xۥ9�z��&g�����g���h ��aU�Kp�_�@�@c||2JF`�N����J��\&�MN^t.�U d���4���g@J�«A��`'=��C t"oQ���-O�y �F�f��7ֻ���"�X!���� ���$�#�9K��w(�j�]�zO~��\Q�8EO�i�2|p�b}�1]��[��)�#�&m����j5P`��_,�:0�D���A�=ƣ޸�:���
�l�
�_�_�ai��/m��b��Qe����# �"gGe�՟�t�ML�r1���i�4&�����5�`JHx�9������H�HI� �K��S�\�Ӡ�<�$��17�O]+s�`������ �g��;W��}�&K�3��*�����|��`O�2�曞�[�ԕ.?�0��6�-�c<�RW���}e֯�9�����<�{ԼE�:9hzj&[g�?�s4��<T��}~�kB�k�f�w?��3�I�M�;��aA��(��Ԝjv�m��4�Ϳ!��6�;��P���e��r� �2/^��V0��$����+�Z`�q�Hq���c�%d�)�����
��[��w�u�hk9u�D[��B��+��;M}eX;{��V�z�8Q��vӘI5��gmp�cm�ҳ�YD)�]¹�$�mQ�s!UOO+�򖦺�fM�����ë��%~!���u`�U����,G��D����O@$1�L�17�E���q��q������>�5�՞�xe�1���}[��|��`��he�+�1hn]r�<+���%�Jh��;�q \���rϺ�1J���Tq�rµ(�����I���j� !m%���e�~����%�Ъ�_�/�kL�*qF�7E?y��|V12-��#���y-�nث��{�m�ɞn����-�Ϫ���s�/$�c[
M�Y�b Iwe'dԊ�z��o�{�o��������V��I5eQ���q77#.p�����)��jA8"l|��8H�Nmg���ƃ����!�\^�gd�m��;y�ӌ( -�5��?��0�ܝ&{(�@�)��K�DR�3KY�6�a�w�k/��^�)�R0�g�8�]�L�Z/�;f�$E��#������n���D�Fd�`����*�l6�����	m�UyG�����ޓ�~,�7�V"���.?n������?_�r^����ܫj*�I�2��2DqǢ��
���i ���? f�� �_#��ѪGR�Xr{�l��t�y> �?���9TN����7��&^�B\@�ٽ���DTG�v�r��g �5�1H��50�v����l	*a�Ø%.��B'�*n����,e�N�{�XE���K���^�!I��Y�e����G���~je%2�CDF����O?��7����Y�ol�?�?	�J�89�N��)K[�s�f�T���s������S'α���p_7�^5d�%?Q���UƠ�U=�e�$�/��O�ڶ9�7!�Ώ�>��R�GG;�$����0�#||�&^x4���B�?�n����c`��cK��ڻcS$���f@9�q�D3��=�ti�$s'�R$ۂ���T�T.°J�	���� }�eX��C ��%�S��t��nґ\վ�B��L������8��I6�H�r� d�R��E��$��w�L��C*+ߋA;@����f9=A��O.:�UlBH���ݥ(v�?���s -1�ZE�?ΝԸ�Z;|�c�"�5���A�]��E�9бߟ^�*l��i�'���ߜ!2D��C��J^�#�1�qo��&�)��Oc����`�L|�hC&�+E.�������%����~ln9E��ahe��s�.D�������l����o���_��H�����oR����zq3~"��c�{��\������Eg�,@� V�������wO�f��3\u�
~)����U�C(����V;���E�����"����]Mg'T�U9(������H�nnNj�aFb��=��oR	2N(�Դ�>���� �ؠPR�e(������r���58��W�� Ѣ�������ٛgw�'�H��ؚsG�Ɩ�}��6��¿\W��J($:�Rٔb5��f�A�.�����8��_�sX�ވ}q����o��^
1p�6�\�I�4���W�鏳�eZ������Ҹ8��IE��'���
���:_"y�xf�e��W�͉�
�������&f�X��S{�^P�0�hm��H��˷@�N:��n{wFN�7t?/y��^�7<�Xd/|���T�H����_�;9Dw=�=���n#"�N$��UC�<�ӯ����D�F*V��"���
�0&Q�$mUV,�K�e��o�>�&-xґ@�Y�A��H#����e4{�j�i�Y֙��OU����਎�^aiQ4�Ȏ# �o������}� @*�|V���w�B ��5���PYR#wW��~a|��Q��f���\c��A��s,P�A���e5��*����?u�nw!
��NaF$��c�$~�f,H>3�fO_�C���r�lD�0���r�=���d���w�}m�Ȩd�X颪�h���{7(�ݮ��p'��R�&Y�iR��>hoL�!��%��e�-����ө�(B���wץ.AL����D�c`Q�4k
Y`H�v[J�����(�����Ǟ2�1����8{�J��1meFϐ�Z��{-�g�|�d+#kނe�A��@@HHۿД�j����>8��g��Lէ�߲i^q���i��Q��S%I����B���|VA���W���"�:�"�·�̍����\��9�D���LI%��2���Ro�p��N�_Z�v��2��SC���q��'��(�z����u:�_<��єa\�����4n�~����[g��
�j�QH���v�A%i'
����g�/b�ٗʾ\7tfl�2�ľ(���°��L.�v"�[���{�,k�
9�܊!�P�9Ts'�����`��gk"�I�m1���փݩ�����VQ;���W�?K���Ol.&�O���UmQBmz��^�� p��iiC�,���ޭ�*t#LT���z_��2O���rb�/ڦ�k���«��k�F~A���[qC��~E�BH'b�j����C♼1�WC��p�U\�U��d�9�O�����3�7	q4�8e�����t��C�zxB��½�(���X`��ֻ?/��|��+��X�!����b��՝��"���=~�*1�"q�J�s�T;��ޅ�O��s�2b[�Y�E1�i�����Ur���HE�d��FL>_H=�yk:�jp�
h���pVct�8Vy��U��� ���P�I���1F�[؛�(1��)����:n(���zX�V��k<,rVآZ�:�n�kO���Ѡp6D�oҾ�� ����BD�[�V�(�3��~6M�R�̥}pcZ��}��Ily�S^"���Ҵ�k����dt��u�dS�����;�i�����#k�vt,F�m���X�1'��x�̀���n~V�{��]q��@\4�2�@7��`ݑ>��4kNF`��<���8�Lj8�~?��s@Wk�8�:� ��Z���~�Y�!W��4X K����Cf��E)�l^�V�j�3V^:�EѢ�����"
��Ts��Q%�����K�rJ�#��ikSO3��f��DP���1���U�S��q��<TjK5^Wb���#���������/$y�&A�go7	�>,F���Y#,ƈ@H���@7H������UAͫ@�_���ൌ�2��a/@���y<U "qv?����-����5Ə��ѐ����Mi��>
"q� �?��N������}1��~/(��k{H����8���ƌ#{3��k����$v���֧��C���]K��zF�r�y�^�9��W+�������/>��Zǟ��{��Y��]jZ8C����T�.m]
��獥q�A;��ſWy"l���	�L�����
����1q�8��@{��'p���w�Ӈ<=��2\��a���s=��,��̝������61�����5�'F�?Q=aXF���^n�n�TR��ÀPӨ,ɪ�|Q�q���#�1�Dq	E�ʷ��CĎ�"�p���f�0�1|��K]��k�Ĳ�J�
kD��J߈��+��K�z�Ve��;
�g��!���;����鶑�{�@�|q���>�O+C��:���JD�\.}���!D�2�br2�������|��T� �7��_k�B��G�rk�x���a�����5�F�'Ŧ{���q�35������Ď3��Z!p���Ex1c'd�v:6֤�3�D�����]���lo�����7���e@n?��.�y�M�i�6i�ۗ*)*�S�v/9�3�ҋ�H�\Ip�~�n�(����1���Kf G�U�.#��,뽻�Svb;1�ӢkL~�%�oO��oS�Рw����(��c�sJO�MPqL�+�࿻��ע�w��]�Ϊ0O1� ������bŕب��F�h���7�x�9L�WW"V{���/��~jy���1qV�VX G���g����A�m�Yv2_����X������':�I��b6[,)ڂ+��KL>=��K��o�2�PƳ���H��s���G�ǝ1�LD�}��1S��i�q'�� C �d�0+
}Ke�@���\<*�ۣ��y��h����������(ζS��&��+w ���`��dm���Y���6b@w��I2>
�:ID�լ,�am���ul,ғcl��>�IG3]�Ǆ�-�-�+u������������A�M=�i�H��\�Z�U�7�?T���|���q�hJ���%�9<�w@KZY�����l3;B^v�)������WdCi�5���k��H�w��ϬV�h.�{�:M���" �_��#�����X@ uo��z蘑	|�>��,cY8�R�4ET`��O�\Q�%���Ho�X 0�h�޷7Al�p�} 3�j�l��(�q���Ï3 �������bC`���h�������q�0M���O��
枊���#�v�k[�[n����q�w����#�	��$ԥ�#L���;�mlw�v#���!����'GE7��^����s8���̤�#(�w?��
�O����h�ƭ����e�V�9 G�g-����'��`�X^{���Ę /.K�����$[uL�e�}x>j�O	.L:?�"�P�"3ե��v?��,\gԜ��V:�
ů��w���S��|�-�Y��P���hP�������"0)zӽP85X�hT�d>	�P���n��ߨkfGZ�"��u}Y�L��,���r���L:�3pZ߈�y�� X�H>VB0`.QEg�c]%����yR�7�|�O��i�~��C$�=�\i�U7.D�be��$Q�j�/4���MV_M��!���9�֎�Ya@�w�8��	!h��
�3����"p��R�BQ�xZH3�D�Z��16�[ҏ,�u���@p�"F���B++T�O&��Q�������v�\Y�C���5����=6���6�^�)����wA�-c��16�� �AsF��U'�H��we}W�qNSU���V��ʉ����T�XY5/��PE ��*- �;�� ��ژ��aO��X����
ި���v���_zr\sO�憣]���/���	�㞈a��/���f5�X>�1ż���D��Q\ۍwMn�GA�!B�N�R�1�M�G�e.�v��B^��!�z�[G6����O��/�9�gb��*S�Ou�`m����KO�%xиsiks�q{g�����@�g�L#��l"�>u�ÿ�A����2�v�<�&�R�l�NJ���Q�m�+�`���g�B���l�R�s��0�Y@��z��{� �$�b�U���3� m]�x��ӏJ��j�H7�f�YJ�^U��Y?�m�P�K-��!�d�� ��-�6����"�l� �_B�����xXf���	�pS�
���_������#/�g:"F������9�,/�@��u"��4���I'��!�(�x�����_��rE�(-B��f��d�7�=�:���F�zB$�ʧ��ApF�v�����L(
����.�ӆ�q��Z�����$S�>��0��b���;���(�=v�k�����V��6���;C�S��w�{�$��[���a�{U�U�&:R�H�K�'�5����%;E�}��h\c�H5l�����Ȉ��˖62�����\�J˥���Ԩcew�Dwh(��B�G^9R�6�y��Qh?8�b�e��+�} ���K����Q� qO�eԢ����ԥgҎ�c<k��e#,H*TQ�����܊����@l�ǣ�����t(OT~�o<��$|O!7�F�l�3o�HԽ�H��?�1���$��|]6y9�%DԔ�ٌE�}0�`4�4`C6h���{��&���&!�a��1�3FˠtO�{ e Sz3y����;����4&C�pz�Ԙ�e8X������N�p@�R�3�VpUI����8bV ��$��3�pi�Y���;z��/*��32%r'���F�����`�h�3��Uc�Wp����:"��w��g!�]�����q��J����xH�:��%�����YMۖ��	ᡘ�O��/���H0����\c~5�	Y�چOyܘ@��*��4@�b�ב��e�BNF���C):��Vr�������O��c�9�`3 m/���CM?ȼ���0��y�����=bm�Sw�$�m��u�M�������%GI�	�n�$�<��˕�{�R�����Z��¶
��t���&��V��K@b�T�&[�mZ�{�����wۺ��<$�sS)��K�?���G�� �\�n�N�y]�Ų��AW�D��A<��K&B�ÿvO�*�@���Z��e�0ˎ ��z��d#�j��tS:�h��c�׆�� �&!�5�SM<��E����� v��O��6�hb���%�.E+��z��W,�s�o���!�IOk�w%Oc0�4k�XFe��QZ@i&�f���ϛ��E���g����y!��W\l�����m�"oY` z/L2|��C�#Q�����1�gg�����8����g�@F[���g̲m�hBFB�5Ks�A��E~��>�ߣ����O����G�Z�/�J�����˧ms6��-��=&��f���r����EB.�s@ν~�zĉ��������zj��n񻑍�-կ���ʐG+����R^���%W�u���)\�^?үy��_ӿ���2Z	��������_���X����
��~��)՟ ��V�m	�����Ѯ�9t�M� &&���|,.�D��;��h�FF}�ۍ�^9��S^%JK\��?C���3)b-z,n|p���b� {�c�?�٣�Oɠ�O�cV����fդ	Qy�u�}�SR9s��G�h�I�n������y�b���TSf��[5Lo���(|�ٰ�SYNЁ���+�:�&g0�9��
�?V(���b-��ܴN�7^���.K�}� ��,Te[�Ec��<5�)�+`�e�&�G3���X9��s90����V��fM�yǲ
�p��n�
�������V���6o���Pm�r ՒN���奺Y�Q,J=���r�PK����3(�w�EN�2	H�N2��G�2u^�-�wf��,1�QL����p�e�%
����o��~��i{DC�J���8/4T�v��Ve��]}��"J�h;���ٖtW�3�sO�h�����^"�\����c��^,��4~�fIv<�9}���)����?�R�⢨r��Ö���:dM_���ɕf ���`Z=}1F�w�����<ʹ���;���^L�(�x�>ڨz�]d;|�0�2HǿE�ZX|��%c�����^pj��5���^c���t`��72y��1aBT$�޳�"��2q�x�ƹ!k�*���$Ŋ���l�"Kzikb=ӝ~������Ź��� E�<yf5V7~r~�D��7�_6]%�d$�����S��V�UW4��-";�;��ߧ��5�o�I��%�G����4�k��R��N��`d��A�V�`�W ��d�>���J#�� �$�η��'Lӷ>�9�j�U��_��f$EW���[`
�0A�Ti̱kf�p�	 O�� Urg���+g!�a�bD��9nَpM�Z��r��]�����l�}�B��[P����j.�.�'NJ�ggP��j���ѫvY#ёO��	�2+���&���f?���J稹�Ŋ�3̽���xq?rX��tu�P��e����a)�N��3�~J(� V��9���}�p�zF͋�W��q��'��=��Ro�o�oM2E^$ �+㷮'��ީ�+ѧ�*��0�ĝf,�Vm;�GPQ��n(/� ��FWj;��㯚�`�|��Ř�p�����p�����~�@
^�O'�̉>(�ڠ�?�{j�g�Zx[/�����l��V\�i<�8Ί�:�#�)�C�{Dy8	J�vl �=��_P�Z�霃��>���Rp��#k1��OE��x3u�����m���n�1B��*�f�|.���������O�%��d�X8���������n#���M��}��9�1�N�"߉S ŗ�]�#�՜ M�I��M#%Dz<)zJ���"�!��K�j��s���Ϊ%t�H]��I��eJP�SF�����F5�TmL.��ZEP���R����3Oy���}<NI�"\��^KJn���>�鹭%�z�r����k$	ЍN��9A	���:� ^��濟��>�u&�<�o��_g�h�+$k)$m���x޿w��U����L?���F#�\��˾]�}�ᵆ�m���C[Ҳ�����YC܆��݇��p}AH#a��=���-(H}����Y�;G�x�Xғ/�ք�	,�M�ZZŤ�C-��\���5���Q'����p[ڤ����M���s�rh>*���##�Y������©k(��+�\y��Qw�˾z$^a��l�=>���jܷ�@Hr���H��(��5j�U]�a Xf�s�δ�w�d��J����^�� ���U��GD{�q����C3�)k�:�p��)IecdF�֔��4�Cs�-�����������(��y�F
�mv �4␿ţ)*�K�"̨t�tr�;��"����-�\i始9ڙ��+6����mi��
���~Q!2�D��}f�@��Hi#��H��ń��x�Nq��ߦR����>0r#�/������[0�����P�=�n��]y��A���s��@xä��<������
������[����
MB{�ڑ��^��&��緧�������⾺ F'B��q�H���
C��گ�X0�٨״]���]Q�(!!��\[�2��e�*Q�"���U��s��
���ң9*Zs�=,R{β�3-�?唙��o�
hM?_)X�0pQ�z�OS�W(5 �D�}��F��ŵ��ߡ���~���ⵑfE��`�n� �@��t7Oש��'S��{o��m�WA�� ow� �iMG\sز�v�Y��P�%~ѽ���ᙐR0�`T�2g�gt7����j�/�m��s��ڦ��>�X�2H����Y���+�� ��@\��ODð�.�����՛�Ʀ�%`e�Q�(���>�B���g�پ��?A���~8���q%j�5-L:���5m��4c,�����]t�:ٹ�h�q���潗���o��zd�v���1mw��� l&?��'L�Z�� Tx	D�s\S#�J���Γ�<�n!�]���/������t�z�ZzkC� k2!kN�(���1R�O dQ@� `˓���)�щu=_��d���$O��Z�	z��Ė0��d��0]��a�-���h�jZa�����}��=��ׂ�4��!&�b���=٬C/�YC��uf�~ۀ��������^����7�z���R�2�����O�C�e3�V��-��/I�0�.Ԋ��)��Kd��H���ڤy�51�ZԽʱ�6�E�z���1����[������ ��zs"	�rNX]���5�{렷�s����Ŕ
�x�J�k{����H�8|��)-�B���om���xF�}� ��H2
�E��k�ו��g�I�ڋ�ߔ��	U��jI;76"ϟ6 B�G� i:5$3h�X�
G�@P5D
 hQ�9^�'� R�z�I/�c��([��3�m�X��&B�"��ʼ,x
�{t�/|V�� �&L�E����W��:��F��^�ӌs�* �W���My~�4,�<��`�r����	��;~=���~��箜ͨ.f���=��
ReM-��*�4�R�|��%(HݨVm�w#���%�����2��{���O���/�����4p
��K��Ե}�#���N���q���2V�κ�LOb21}�����X%@���l�G_t}p䩤��|ߖ���1��R��1�eҽM*��Y��|��|��M�O��Jq�C�XS6�\��lG ��q*��3�-�@��C�Aa_"[N��2����:s� ׻������gT�Tӥ�@����z��X޵�����ta_�G�x�[G^_t[�e��+���wV�,4�!$�rM�e��Y�q����r8?�ҹ�|'MeBhF/_R�@1C�\��I�ӓ'�̼�6���˵������em��y=O��ڛkb�,��o�X��:�Vl�"˵�O$��|���pJ��N|J?3��6{d���G��,W�@�u6� R�:iT�N����+?��Ǡ#g ���UO�(�;lH(�w���x8Ӝ����?+�6x�fm�H��7^�J�Dh�/Sf(��L`�	��
`���!�1�%Ljc)���>�!���f����QMT�Afm��� W*�n-�UT�w#�C&��-YC�,��=����0H%	8��|�H�8�Z@;4g��4�q2�Bs2��D���Ƣ�(��b#1�0W����GX&Y!v�Wr�G�-i"�h�W˳*�R ����^
�)+��]0�iO�u9ѻju�Ko�-�xYA�%��5�ё�,�P�"�	\5�T�]���m5�9��m1G#���84۳%\z�ݿ�Z�kb�yw��n��b�U�'Q�>�>��FzScMơ�U�I+��&ixC`�nw�i�=��=��1�3UP,"z�t��XU;��)5�}%8�gZ>;�|�q�mLAY����p� ����;dyP=T���MG.n����u��	����A��|�~�J�������n�š��g���b�����>2���U����.y��o� cru�'�+�l�����`;_�@����_���N�Hc��Ѝ��ۆ�_I�#�F�⮗�|��,�O�����Gw�PS ���$O�I�R�� ӑ�G8J�Jg��us��MN"_9� �r	�C�}��f%�p�4�&)���uf�I��<U�j���kI�i��	�`�\�S�;����c<{�w�ls��2������ħg�\ŝ�h-k/k�>F!{�+���S�j���_N̐kS������X�A�w��R�1��|_���`��jf����xB����+���$���Ł��9��ē�bDw�W�/��+��z�V�nv+c�Pv��C}�,�H�O����w�]&��Tv�����$���$(ȴ�]a�;2�޵0��_r%,��;�5l��������'��Pp�c���
�q�r2*J��cf@h�x����Wp�>����yBHڽ}��z)�9�P̩zY��������K�=�s�w���A�_�p�P��,�d(6��%P�j�5��F��� ��Z(#C��w�MF���[k<*�Y������F�2���:R.gmP��VGS�������>�����\���di��3{E���ݠ�����nV���c�v�`�r�^�W�~�\2L��\��|�µ��k�[KXW���+��Hlx�tJ�B��y��^��U��cx�w$,Q#$[t���	�2fӃ56AS��_�I�v�4.��N�)=����p͵���D�7�(�O�x��>�>����]k��%%��������nM0�.1�'�J|��tO`��G����D�M|�Η�O�[����Ԏ�Ǥh:��܅�-����lmq��M�8���e��r�cؗ�Zu�Ɨ��V)H����˪;�mR~�P��T+M�R{4���	vW�,_F\ָ�����{H(�\����1�v�� ��ZB}<�W��Z�A�n�Iqn��~Q�uk[��� (N ��;H�;̟�hU��$Y�S���+�����������dnߞ��7�w(�]���iR�.r�#��s�C���8�*��F���2T�4�zE^f�k�6�Z���ù���[�.�n*z |i�'����7Ď�R�?B��zo/W�xi�i���I�\_r��.rzFV�Sr���7�i�ST��e��������_B�hʈqo�(+ �@��kC�y8z)(�*Ы��<_nwW/���F�v��)����9�C4?�ol���P'�� �s[O	���ʆW���g���V�����xo@x���ty/A?*� ( '�|t,߶b��t�س><���J��ˆ�Pa�P�&��F����xT�������Cӌ�kK|������.	�	������AsDw����-�������}�^q�j�|x�',�(�s�.�6WN")��$X�=D�%�[`sr���f|}W���O�hr���y��0���GZ�˒o"o�� C�\n�DJQr���	�π�ns�Q�-B�B��C�)���i�A�f�sF�	+�u)O�)vm�Ui��� �aCɣ#���쇕v���fZ��s��z>  ��@I˾��9���>��K�� %�.~����(= F���"��'���9l�pIu|�`fq.9?�+�76�� p�?iP�;����>{��­ٍ;In��u �R1z�z��W��"W�9��Ԍ�AR�|"'�&��a�=ԥ~(��7��ߣMM�m�Zp�/�:Xb}�P`���L��z2��-TH�MRQ��������y	Y���� ����ʉK��潿{ş�'�X_-� ��]d��^�g�gm�U_K�א�����,u��EƵ��ҖU7�u��A:�A=��S颚�Q�i'��(r�@$?�y��$	�8��p0F����t���BSr���e!t�*,&�un�9�gF�ٵ-e=���G@uˡ�~n�,Ia�e�S�����������82�p��v*${�I�jϕ!�g��j��JFE��<�zW���4�1��F*�
����n�Tg���Jѭ~�)ܦ$�%,����LXb���q�+�G��5A��U@���2R���S �F��O$����)MKN/�zkwo�oJ/6cz1G���Ȩ�)c��(d쪉{�l��g�i�b�3#i/��UZ�q3�{ч��tgz����
ߢ�;=�9���e����8q){��������SZ��Ƥ^Z�.�����P�绶���搐/�ª�V��*��ܭN���t��i�����`�L�Q���<t�!l0�.�	����\V�٠PTR� ��v\��,���Ÿ6
dw�M���?��hB�a�VI ���78�nF���%���È�1f{�8� �)ۊ��p�+��O���cqɧ�vc	U�,��������6gڿ�HS+0ķ�ό�GZ��mnϻW�ש�\�e�|���(��҇d�q~��=���ih�[�a�����r���uıh�2�5 gʑOzR�/����+bx�O
�r�I��Y!5��lk(gy4j�?`uf�gX��~��ئ����Op���	�z�}�j �D�������� �0��ל/�o���ހ�]������2S�2{��dGd]@ϧ=�5x�����~�@b!As������q�ʆ�p�ҍ��A/*[�]�����_�d�=�������!���a���T��eDfc*F�Ľ�d`��:֪\!�����$�nO=<�2�\]d�T�Ѡ߆>���Bg|�o����7��)���Y�|�Z��?�Q��PN	G�d� �Y~ \d��y#��� �t�l*b<����r�%}U�\��n�p��:�$�o4��/X	{������,���p�FSq�R I��ĭ�,��&hi��☀�bB �X�mˬ(�^`��[��o���>�ӭ�9������5��N��n�_�����bj*L��t�@v�n�'zh��:?�wВk��hظO�G�.�O՞`j�vW�����3�Gm+��o�r�~�Q*)���h����z�v�0������u�Ɠ�w+���ǐD�aܰKX�g����w���ո���Ȕ�-5��MN�/�+F�����G�F
�B�x����V|?$9g����R��F��\|�5��:����+l��΃��	$Fun�ꜩ���ݱ�i!hs8�;_5L5ʮ�RV�-]��!B�r���,�zY�䍏h�`�be��Q0ٯ�f>x]�l�lF���	�C;�s|(�֖�z��`5���O���o.2Jo��^��ڛ���~�6� ���ۤo?@t��r��zn9�:�ㅒ���OF��ea6����2��W�'��/\� " =K��m��~���ͽ����J:.����QGN�:Q��&��(��oȗБ��� �]tr���M��������X���?W��3Ρa�9���aG��R���r�]�`��+�^X4r���j��IQa�7��z������ȜM�]�I"�l_H$��@���u���)�٢c7Sk�xѽ��*��F�UG�8J�y�/7Q����X���nI�ե��3B�6�lz��ѽ�v�P�E��!f����͠�d�����|�������/k�'�b�sa���N9r�i�v�(3��}ЊA��<�ٲ��ࢃa5s���»��8���v#8��&p9��JW��QM��ڝ`��ځ�q���;��&�!e"!n�*A~�`�ɟ���*�)���QR��,��,������$+8w�l�:a�J�mw�B� �$
�;�&W�Ƅ+���1a��:����$����Tw����,�<�����~�0�rh�e�-w/���Yk[B�ܬ�$��z���}3i�H�%
�`s���j�h�^���j�;rDHJ�"���勜:6(g��=}�sPl(հ?u+!d��O>l��r)5�Ms�o���̍�W8��L�<&Z3*�!��MΧD|r[Ő���^? l�q�n7���EH'�8�@p�W�	�d��L:C�Y	�)9�B�#���c�@1y�d)�~Ë�Tv�ɹ9ۊ� |C՞��B(A���Q`��l�\��L;6/=�37{e� �l���rH���5"�tl�~���Ϝ��%�HRm!
z._�|�,��|��,r/!H��9a������A�ڥc9)P�W�r�HJ(Ĺ���_ȷr������t�ſ��Ǐw��ߤk�I��Xm$������Aaz����}���)��/V���s<,5崺tG�f�3�Wq��e"Ph>�����k�ZyEg�&րG?�� <�0U]�]yG��W�\�]ϲ��n��vk��.�1�Oi�DϞ��
1��l���ػ3�4]f�s�^h�.�,u��Ī�lQ�K�E�?�g!x�eU�)N1������3�H��z
�m�iu� ��p\*ZA���P��m"���_�d��;3��@kg�lÙ��!�}Nɴ�}-ҙ;Q2��U"3����vcb�}��8;��
��M>:_���l>�TIQ3�p���zUG)o���{=��!,���J+�<"�X-�4>�צ���Ai�Ƕͧ(���AM�F:����9�=x�0�5_���軱�y/X�i�r������(ŝ�0�\X�4g&�zq�N��6u���Y���,�tЪ�E�V+��@��^f?e ���\�0��˅��� �=�6D��k �+\B��[�9Exx[@I.�B��������tAy`|�R�;q�e�4}����M����+e+*�"��Dә𿌑e�;����V��\9��� ʢݢ}�z�0�e�T��J��O�y�d�5j��^�Z��5C'��zw���3D�y�a����/$3��.�dh�g�W磄D��:�k	����R�߯�l��4�_`���gl-yW~gb@#J暿�r����_�]X��c	�1�#fB�	&�
�S��_(�jL*QB�����B3��Ki�{s��7�M��ˇ��N�hʲ^k6��,q`nDs�����Yֻ�->�lxY�ƏLm��ԗ���}[�QS��k!�^�h4_eNomڜ���z<����4E��Y��d�,���#?�;����s��0}a����݁�8aΥ�4'�,S��$�@92�|�����k�y��3Q9l�Cm$�|��d���-M)��~{��'i8l�RV�8��y�$�vi&~�!z�_b'�u��-�@lp]��Т�"-\z.�&� ���^�p�$�D�,JF6ؽR�9����K7�@m�5S��_��t�XE���%�{}X��C���aoB���й��ĸ�g�=TdV�B�d�Lm��T��w�o���'�!{y�B��ry2�_!S)x�H�lCv�K���[ߐ=�=�rY�S$G9�0�ѫ���!�a��xP�k�kYǇ��6?T��H����u�" ��ؙ��ZP�h�ȋ�Ψ05���j�~�̑�0<�:��*S1��(�>�Q!Lz�̝��	9iE��rt�-��g6�W�C�Q�!%|��%7�`3��Z.pkCo��bH�ċ��촮PH>yg��i`��ݲ����s+�{�Q�d|<�v�4H�f�r���|/��B��Un��%��E��#�ھ����]�r����B��Ee6�"sY�~�6b����Vn�A�Pw��7��oc��V�Q����b��_�(�~2��_�.��,��G�/�[���7��>��@�^���oXu��.ͅ)��Yݮ6��o��p���ϭ�xܭ�5���+yL�`,�r���dYO#�S6-��-9&��J���b]|f�c�Ӊe�~��M��/�ؾ�Ă]�*Q@/��j���r��_���F4� m��h�f��-��Dt�s��C��V�4��L�g������KF�\5|�ڴ��JZ$�/�,MT�`^E`ʾ'<�|�0�SW�2~	�3�oV3#����R�bHOÂ5Z�����ToxĪ_�޵:V�B 7<�Y��ue|�AW�v����ȣA��2S�2tV� �S	�EsA�@�Rwh��B9{i9�a���~���)e���AJ�-3q�(aJ�Kx��~˚CaM�C@�  ��E�~b}nK�U���M@�w�W?�7+�|~eq�s�8��5��T.:<�D�vptT9��X��F;��
�A�@#T�t ����X��"�Mw9���}����!=�/��0N�/P��\�@g�t�QG7�]n_8��2� ���c�0}}7�%{,��hA�݄�$��l�$6x�v�xBm�@�.{�;��O�d�L��Ʊ���C|�O��S�;�U�$VrP�׈�-�B%�h�]����T͡'�:S<��d��O\pW	���q*;�I�BW�k���湡���]+�\H0��$6ښHț����̅�r��{P� 	~�,6���ɯ�4Ƽ�� �|O��6�6�`
'��!'�B��#e_\��q�LC��N��דrĤ6��sî�������p�̔���'[�K��߼�a}�,ed�U8#`:�^�1[���"4gYm�Z�,��8���� L/����n��ݠB�T�x�I��-y�U�"0���LN��,��)z˒-f�1Y��+��"���S�ї�K"-?��!�ۖOT�Lz�B�]���z��Q^�l�S��γX�I>�P�Ǔ,�!~��$?���cjs���w�{4��{�a6�#,M@+`z����^�J�fRU�p剃W�^2TY�
���?1vϬ���� �!G�Մ�Z�6���Iz@��:$v���0M	�'tz�akY����]%Y��m��/�W�സ$�̂�_Kܱ�Z���PnP�2�!��ѡyڂ{���b���	��{yx$s�+j?Cڬ|�0$�'A��!� F�&���Ø3���S z���n��{��ڃ�!$��@��U}cF�z@ ]E���y�,BI�4�[�ӥ��_�9L39�}N�R��/�ʔ3D�Y�)�L�cLF:��yMf�b��m��g״U�96���>�O#�P7C���X�$��Ȅ)�8�;!hxn��� �pCD��S��j�N�95�7��ߢ©��yH�L2Л�Esi�(����Z&��ZZ���C^����	s�dH��Ν�����Pl��x�z%%B�?+|��"AR��AMăJT;����aq���*�Z��s'h�E�j�h�+!�b��k�A�7�/g �E���%ح�F�#%�%'Q�O�J���ѥ�0��)�y��yvi"���%'�N�hy�j��Y�cFxr3�@�N���)���49Ϛ=gY�6Ҽ^�0���������Aw����k2��y"��I��bx\��X�PľeQ�5�6����Y��t�~u�W��>>H�>V�X|�&�|�2�����hy��5Тf�'��ʒ��@T]� ��yq��k��GO>i�{�����8?�	�dMD`��i䭕͌��?˿9 ۀ�l��˜�<��7AF�L�}I��=��x���o�=ب{�Yh$���Z�z��f��,M*�O�Ck4�8T���~�%@�-�)	c��]�8}(�D����1A:��;�v�?�^��b?[�����擗���2Jy&�{9��.��^/(�0����
�zuq��9Wl^���_��ꚭ�����W��n>��"6s�*�� Qhob+X�g�}���a�$y5SA����2�3�c��;N{64����,(���,�i��z�VJ��
���	#�%Sx�2�5�j)� ��w�Roj(+ӳ�޴#�,�-�k�ё|W�z���a
y+x��Lk��R�y³h��x}(�ʈ��=�Usq{�&ڇ�Mx��c�p��&�u��W^F��_o����3��L�Ip�XU2o��6���A�R��Y�T9I	�W��3�L��>��h��=5�Ď�I�lb�5[�GSr�}6���5.�)���&zV������fg&�_b:"<��_sn����w�4YS��K�%��m���L�a�����w^�`�^�[�o�������B'�N�c���������	�]N�[ "��r�� s t���
�1�X�f흁������=qE�y��G�z|�?_����B��T��ƥ�ߨ�Y���e�F�_�΍2�L,�:�m�7J��	�ə�f`�|�������!��o�B;�x�Ǉ�p��Y�#Bf������%�B)��E��,�@r����憥+4#m��Dh��a�g��x��0B�h0�@�v�4u"n���B$�|����c�@��]��+o�5=d
�d��72E����P%�s���ƍM��ؽ��R�������`�����U&Y+��B�m�Vj�&K�83;�v(	��q�$���+ƃ2),��@Ns��Zg��C(�]3i$���6��z>�K���)��#	[1�mW=&A�W��E�0]z�H�]��Ɲm5�yt��{�T~6�԰�5@�+�]��4=W�]y1�7ko\����GKK���Kݜ�!#
��?�ń
닯~��1U�Ʀ���Ӽy�m��夒@<G�SO�]�( E�CO����vy���4�,@�C��#ߒ���!2.�8�(�3�	�W�[$t�{rA�7�\���3�Ӟ��Zs-��]f�U��O�*��h�2M��o����k���3и��=�l/�8P�Տgџ�E��>��4%^�y���XMe�?J]�@���j&�>������`���,M:^�8�&��5V_I�S����#/s��Q Q�ԇ�HXƂ�4�:�#\��c���Kf?^S�2�0���+�����(|�V4V���IY�T����s�Z�����>�gs����)mK���שH;Z��]�5N�ו�l���N̅{ǭ�]�ۋ��Nh�Wk.�r�k�)]}"E��x��E1liU]�:��К[�ü�r�WQ�!R���ǯ��^����fŊ���)��J�~/���I9�	��a���B,��=M�-G�fi@W���6�Mu��ԩ5uc�G�rk*�����Г�KI>l�Q����@_�9���T>yGB ���y�W��f���Eh��O�^�eI��� ���U�9�WʌB�� o��4�ONM�=1/����z�� ��O3;�ΈQA��� mt&� ܫ̍@ H��}�
�������O�!�_�Z�;Y�z zu��5[��J�d��`S�h�:==��3t:�{됤���S�'4�J2ɲ*�i��D��.��5�6I���頦�}�矴!�s�uo���h�	��A�B!�V!�.�h_�%�8��S�E*�����ʝ�m�Yj�9j�n�g%+���X_g6�H�V�;�[��t�/b*33��T�4y8����L�9�4�:��Y��v��ŴV
IІ��@SSyd�x3�2y�@�eo7�ArP��;G�5�-.�%�"+����(�b `��p�V��7�i���b���"�ѷ����`�燈z�c�nΙ����p��Ї�o�#����ϥ�ڜ�э.}B�]�>���T��'�1JF;�X�%��g�U�E��!d��D0 �\	�V�^U�fU�!�
��)�
z��)V������A����� sk�,n�$>3��	q�+F63<�y:� '��ҹH@�e��w�meSmY9�U!����r͐��y K~
~C-Joo��m^6�΁��O�I���2�{�L�]8](o��4�ܑN�b�c,���&��N�N�S�瀐����G`��v�;h	-�E��ܹb=L-�0����7�w���h�^�/ٝh=��!�R�q��Tu�ת�̉�qj��y1mx�]�",��7��8���G���$�q{�Ǆ��ſ��i�	@����6o�4�Y�� �KNE���~�s�ۺ������<�^D23Y�P{r��� S$zr�S�$.a�	�e<��U&�;�bf�s���o2e_���и~��|�	��W��y��;�����Dΐa-��
!�"�i�&GMI����8:�����X�}��(�S�[��?n���:l��I� Z�lɉ���Љ^�8v�Z�'�:�'�>�U}���g��Ác���R����{MqAŮ�G�l�	n��`�h�2�pH�OR�G�5�i�+5�������յu` NE\�YLcb9=Mߋ�pѤ�w��%�u:��Y҅G�w���RF�~��G����*��/���J�������4Ťu<�:����`�l�������, �"-��tK�D�]��Ш���L���~ފ^�ҫx�-�\0��y�@7����v�찯��Z��VTf����P������2+yh!���F�d���s��m|F2��r`��
�;�G��(��l�;�е��g�����k��ۦ�	_|#$��)����)&�T1���6;N�@=��_����o\a�!1�r���N㼩͠DS�1�f���7-�q��`Z�p�O�]�4@��e�"�92�_ۂ��#�=�{)�gF��lI5c2�,H�3�/?���*�1K3��̴;ɇ�zc����7e$0Ϧ2~�o����u�U(���"�{3�&�-&��K�f^�BR�kxq�T�*EO�_M��1�[�=ý{WCb~?����N~�	5nq?FH�~�'�a�8Xch����Q�h]��<RD7��cPa���N���"�O��b<n
w��煐Q~Qz�gp�����%)�{�p0Qe>`�m��-�~��ß��-dh��j�F�z�[���88]s�0HYMiXJ][�2Rs��dw�"��g���H3[]��o���xm�8�~O"u�I�8u�P�*�!�_E%��@�yÁ?�0��ţP�p�KƊ�Y�� )z>�2޾��&C*������4���Tc���b9�NW � �6n@Ikϥ'�vԩL��e��p�&p�_h����o�;J�:�48oP��Z�lۙQ��K�}�8�{!k�*=�b������Eb%s��A#�ԗ�Z=���(��x*�"��1��Á4��k9��HdA�a�!O�GC�.�kr�p�֥�]l��^���^�f+���.m$ͳQ�M�!0 �	 �@A��JP.^�J����aQ��N@��9�?����,Rj���x��!C9ךP���޲�
����"깈n�D�{Z���Wl�d�����r{�δp�F/Z�U$�7#�n�?%	�쓗��P������3nKV?]ߡf�K ���n��a|%��{���z���m4�Q�
l����=��!��V��a�:���vs9��I��8���^$�㶾-�e��L����}=��PO�M��2�!��Z"0�}�M�qh��o���㯏�k�:���6�4Y���ئ�D�jWa�E�El�Kb"��Y��R�iQگѓFֺc���G��|�=^k��(B_����)\<F�6�|�&���أ
�U1�7w�s�v`�Ϲ�:ǼNP�q���������[�����P|"�_m鐳����aC�zqM	���i��ǟr� (�b@I�LpҦ$�x�޸9O,��t�r�%�Z�н<�K���^��ݨ��м��^nY��cR8��]T��[�t��RK;�7���$��;���^Jǭ?ɧ�Q2i6��C�eA�&F�Z�	�
5��먹<���ޣ0c{F�i�5z�S�)@!l����}uȕ��D�^��]���#*���e�<NUQ����;U���-(�S���"d�w5��8��5�r�֟���[�^�I��S�2��q�BC��(�J������PH�Q�W���6�!�vh$m_j�G-�Rf
x7�n~d���>|*�g6Z	#~*�J����+��yϠ.����&F�Ee#B0�E~��ܭ!4O�G�ذ��mKu �P &;s�TK�32�xr`M�\3[���?$�r}7�SC.�X%�V���{�%�� ���9@�%���h>��<�<k\+@��Jt򎼞�
L��oy�,�}�u=�L��P�&�KkWl�R9v*"���ń�g��!\. Ӥ穙�gg)������]LŲ�>�63o�M�ұ/2}p��pG��K���k֮�s��� h2}/x�������kpf�{��Y��'wٱ��&��gtͺ��G� ��(�������_JiU��C���Pd��a~� 2,�k[�Ck�to�=I ���0���7�l`K���t�>�2Z�Sa�V�"���F��5��	��"O��#3�gƷ�{i�j,�3�h�5�v�>̊����KtHL��!�/Gv�����2���}��M�F<Ձ�(6����İ쟌_SHű�}����9-J��ٖ�3j5����p���ԟGS=�6,1��4~b�t7lgQ��:���D�q��B<��;��m^WY�+(�>n�hRV�m5&�/��sBe��;��}Q Rq-����4Ό)8����D�k.qK��o�����Ʊ�M<�aH�SV����줄U���ԑ����ٴȆ~����i=���@��Q��f~ k�%����jȡ���N�-��a��R�����|��Y�J�p���D�1T��5М���NzYf��Y�&�������?�*��g��&_�q����������NNZ�.���:,Ӭ�����k��=�TP1���*�I���!��VW�n�J��Y_
�����c�����{�e��e-<l9&8޵k-��h���{�n� U"�"� GI����%���H��Py�ǧ��I�ߴa2��b�	��݂�3>����O�` ?�� �1�5\�]Qm�[ӭ������V�	ƟX�N�SURl]��\��<�ot��<�V�ma�C�|��:���5�'��F��_�D���Uv"�|�ݼ+DB1{1��P��^�!�-kT�V��;f���+����<,�x���?F{�C��/��;�8�5_I�'1�Y���!2���拙�[M��97n'6J��EW\�'�Xc���S�-;n�5D��^�5��#��<CWQ��3�e*�����p�i���{���@؛��%.��d~�:����ERm
^n��K�2$�n��~V'���ӎ޽�^�0H�����1��)�c�6�3��J��9D��h?���=Ijwz �k};)����"0��+�鄄���kO56|ىG1jA�.ϏV���a��X�6&ys��L�ꆝ����s�덂�D�XH�w�r92|���V��-�K��g�HSV~����'O�%�����~�3��C�ԑ�U����r�w�Gޔ���??�.[vM�}�g�d�b�%-��b�c�N�� ӆ��3sfL���f��}6=Q���j��[�\ �EH�	Y�®-�W��[�ơ*�ړ+.�a_�ݐ��q�CȈ����0i�~s�&�����R��D����$�G��� ���5+a�`��!P \0����l)�w����9Z�
����L��od���A���[�s~���=���
u�l��;��ÿ5�W@� �`�d��}���#�qP�(�� =
S ��E��܅�㧩��ޞ,��OV�����	1(�b����x�Y�l?�Uد�*h��N��$z����#?nU}�O�RFW�`��t��Sl���#�ނ	G�Z���3t�2k_���T6a1�s����.��
P!�eb*�Z�i���&B���o ]��1^C�uh��w��Q�rp��<��M޳ts����CI�c\`�Nsx��UC�F+%��ьU���O�;]�t�J���D��J-xeol�����f=-��LV�G�<F7�\��{e�v�]�7ė�L)wݳĤ�D%��3�U	��]<6v���Cw���J�����Q\*��fMSSnΏ�Rdn�k�6�#�c�^�W�:qI͍ 5�(��n}��`:��ϺX�K�K�i�*�Q�/D�t��=��%f$���iڇp���g03 &���)�a�;I\{=�v�[�� �$�����tc�����GNk�f���.�k����i����Հ��t͛wy��+�m���5Si"���ٺ�zc:�N'�
�WD���Q/ ����^�~������=Uf��.D�j"�P��D��=��FV)�͗ߥ�y|�4�x^&��G<�	}|��+��b�߉j˲��u��DWE��aH����]U�8#��f"t�����.��v+����x蓚ِs�͝,�9����6΋9^����+˴�:�׏���/��U~Ƥ�V�#b����RkY�ȥmƐ
v|�d�\Λ�i��yO>J0Xs�@���a8c��8pQ�ȼ �;	�m�%������ȷ�1$bw?X�d������]�")~���|�/�~��^���D>�g<�}q&C
�Ժ��tf�����^ծ��^|#ȋ�ȳ���PHJ���rG��=m���W�P�E��>��Դ�w��m���ʦ������#��]^v-LtU ����4m�v�O�ѥ8��H���ȈVh)Q��N���n�"�W_�;8���eI �?U��n#�[P�8|��f� ̡�2�@�5{�ZGZ$��h�b��:�͑ZW|��<�1�dS#�W���N��-�(|��X��ʎ��uf�(�~��c�C,�2:��P��@�Լo�&#�賨���Z���%��<�͵�$Qk��H\kxl$l��y`��=��[a�U�0S~��>�2@k����}��"�?	�����n)�j����W���/���d8���	LC��dlW�zt	�P�Z8�
�W���r��+r.��[>gH���.�𭜃"׸�HR�+��/ذ�C�ߝ��	>�p�~��yC��f�
���p�@_V5S	�aZ0Z<ubw`7��Ş�o�ZL(��;Q�(��3��xs7Q��C�f:���$Р������>1�-9�Ә=GV����������q~w�!n�Wo	�k>�!.��n����]��E��2
7}#�dnu�ڢ�ڨӟ�E�2���X���ueh&Rl��X�W����%0�`��D!Z��\�uA&հ�soٕY�	ά�LᢢP�'��:AE���.�M�b��U�С|�i�v� #P$sl������~bg#�V��,|�L���	��$Ң�S]��0�Oki�_�j~�0���)���S�w���醋��l7���fd��v�:D���A �	|��U���&ĄA�m~"l���SǑ� W@��,���gO�A�p*��A�ˠ��ȔFG32s+��.z�rI�Sp���ǧl�YE��O$,\��յ�<�bb��ȧ!^H�7�����1mC�����=F��-�O�@P~���6����֍J������g�ʃ����{@�!���n����YE�H�fΊd���If�#�xg.�n��1Jb��,2p��$�ٱ́�������5��Q^�D�f@�MZ��Ba(��0��זl�f%��X�X�6�8`���S4���+�I��]/z�)�r�]�lG��q2��v&��xdi�_B�CMN
$g�7#���=��@x*�&��B~թ�.hq�6<�:�L�_����jQ ���|���RiϽD��b���}���~��U,n�q:sP��j�(�\����:]��4a�K����%X��Oɥ�ڲ�Bu
ŝ�usv�V���eƹ4Su������֪�?[�nz���t:
s̟�:Z�]�����V��qO�L���n��B��^��7O���#�v�8����#�ow��I��"A�y.�g��{����-�,��֗]O�w$f���^�@�lm��!.���^���V����71�le�R��K��$�+��֓�/���[�����u�t"�)���z������g��g��w}ҍ-�{�DST�$&6�I�ک��6�h�����O��㩄����P�����q�}X�\(ݲ�[ªZ��動�aQ�����&���L�?h�5aL�1�Xx@ �j�=�@��P����Ifr��Ȗ�k���bU,��!�N����<u�����0OI�_+z�,�M��lu�W�ДS���� S���v�y]\� )mIx:\�l<u���Kz��'��h:����n��2���
R�6hT�:�ۆFvi�ef���t	Dú���0C�jll.3�R7���������^ʒ�-V�W���D�ч8Q��Q �*�5~̨^�"�xF�_k�G�䁎@/_;�TJ�Տ��@�1�0y��qh}��25�����]�P�Bz}�a����4<� �:t^�l�]��L��G��]&��[����C��m��
��'~�����[R�r�6��Y}N��G�*��`���.]������h���l���e�-�Sk=%kT0���?l(o��Sz�.W���ű�l�M�}3�5;�6�6|V����c��4��0"؀�Q=�'9�F�,�4�8�E�qE��̦.��$���
rAD�YI'��v�(Z�����Oڲ��� �]E���zȦ�K�yʏ؆�J��p@�!k����?h�:�滲�,���ѩ1!ODi׾Q�T�\�N����!&ӻሡ�+�XL]{��U�~#�뺀��s�*�#rǭ5�@�#e�Q�v4���G�� �jU�^�'}����	i�������C�k��=hS�F�K� T��p*h���4*gh,pٖ��h�Jş��:�'پ5T[lw#y�ў��Bڠk_�M�(��������)$�SD��2�O��U�hã���C����0�L�X߂��j���s��,b!���C3O�:u�M��/أ�"�Ѝ����|��������;�y1��=���͕��,���x� 4�ɩ����L�ߜ��T�Օs74�G����G�e#���q��`�����=�}'b������\��i ����5&*�4`�ń���[Y��X�fi1 �|��k��t�k�^˷��5���V\�:�Nc���ez��u�M�T��Zr�>� Tf�zO��3��rte328BR�̈́E�P�[��us�)`F���S��~滤+PF]W����E�JE�/��?�H���Wɥ���#\0_��4�����N���sY�EI�KJ�nр�D2�穣ga)[�aN_QVӢ�	xCr�u�����)��C���g%e������{�^I�/� �*�3�ݯ}P�_�<D��}���=p�l��3A�����eD�-����ɸ��5�j����k�9>:̪��yi)Hk�L�q5{ȻIT�����g0�
 ���r[h��t��R�ςݰ� ��6RwcP6�O�rM{/���F�ak����,V챘+�V �?wz�6~�b�������QwK��-��+*m��t�5`Ir�p�l��P%��]=b]��f/h���s��"�H���U^����b8"t�~��@�8>�W���-M5�}�fY��Nd����2'j龀e��Il;u�>X��f��� �p �+5�.�9��,�ٝ��Aë�L��>�1$��0�����Pk�Jg�B�z�B�0+�saH|>3��Aᚸ����ڍ/Ιp�%;|���۵[^YQ��!e�n��pT���1�����}��QԻ�i�opr�E� &�TM�&��^y˞}�RW�t`�����cUT#�Y�ja�4�%�k*�/<��?��������5������&h@?nn#�M�/�)�����r`d�{�	�h�(rm
?w�Т�J�lJ}N�?�tu&�����l�GN��k�p��X�%�ܬH�i��naщ]��I������_�u��]������H�΄1dYbs#29�P�("W�|4��U5���	�C3�dEQ�u-41�F�3�Mq���d�{|0S�XaVh�{����~v6��Lj>w�p�($���1[,�T�ѿ�2�B�zJ� Z]�K��s�dZ�ۼvC��/#�/�6�l��_�����׸�u�~R�?f)${�c��j̽�C��x���3ǂ/�.M��-o%QV
W�#���^eB���#��-#����|B�F�v�Q�g������\�ID֠9N.����.[n�@���������&���k�?�l���κ.�����}W��;Ϲ�U�������CJ���Mz��a�.�ڢ����ip	�s��F�2��:;�RQ����gX��e�AǏ����^1.<*�$1hKMB�Vo܃�ʄ�@0!�@+�~<����wT.Z[l�:��];}%��� �P�>����o���K���A׉W��R�֞5��)1�̨aTY-��=�D4>�$J'������W�-�d�����W�&2ˠ�bx�b#�@YC�G�B��(~k����Y��#[�â~V2o�"<>�(�o��A�pK]J|�*x ���B�a�o�e���dxC/�%<YӒ�}	D�o���x���|��W��w�"�,	׊A_��]�p`��<���/Y�q��@b��ܑm�2J�'߀;����&?�9s�G�����a�[�T���♁/^���~)'p��C܊/ˬ��]�j�{� yk`��I|���ݺ¥ =˞��"���x`��aYDƪ��:�����̾F�f̪w=�����f^|�vJ%Kޥ����6�u��i�|���j��n��5�<[R��T�*���c_�ԉԄ~N�q,=���7�]��c@���Y�w!�x���)��1���*�qX�Y|���45���������߿�K�X'����7�`���[IC�W��o��E��p6�D3ϊ(t�� ��ǾO�w"Z/��vf��W��4�w�r��w���IވL�4ǥ�*����'ʌ⪮��u�{y [&�5ُw������zR����s��`&`�r`g�RIu���b1&���_�Κn�$���׻-��tڨ�T�ڱ���.<�z����Vrs����񙛄�WZEҥ�jA�q>O4�g�x�ŕ��;�\_7s;�B����'ؠ&�ꑑ�+�ƿ�N�a��^^�N�7D��8CZ�����g�0q�cy�0����VLy$�n-Ʀv ��%s�R�e����8\�|ܢ:���H|R��,�(���,��_u�`���y��><`�r#-/Y�҅�ui՟�Z]�޴�E��	���B_���$�HFR�4�f�!�q٪���n��}o�1#A�	e-W^($߹�Y;Yr�-5�K����֞uwvt�9j���}�6���������Z�_�,%R�Lr}WE%:B��P����#�tO�
m��al�qd��^`f�p�#�l�2��f�jh~?Kaɬ_z�owbJ0/7Q}V7������?Y�ܵ汇��1������6�� ��&�&C��+j�Ҫ����# ]�l��%����!r^4?B�VM�-R
�?�S����`�X��6���Z�w���q�놌�4DF촥�ɴ!k(?��c}6��Z�dV1�[��e*���>��	L"��J��W#F\��sE�ˆ��1��
�d�����ˮ(^���ՌX�c��xț��56�9k�����R������%&޿$ 6m(�����Az�^HӒ�8��=T�0<#r�k�B%�^��}}�Nr�W���0���0|kl�X�����<63g��h�*@�`��j��d6>�YK]���K�Z�v��n�8��!�ef:�# e�dX�_��ޱ5%�o�%��&޹�}wtdZϨ�����8�v3E�GN�����:v�5��t�z/l'F�<�K��bxS���.g�)��w^����|�`$KZ,��T6*��eV>t(lQ�g�T�S�6߇��c�Ӳ��f�9ZoE'P*�G�}h����ǣ�~����I3qBfۤ˲���w�;Q/4�t�Ӵh���}�>S�Y�h��sH�M��l�Qk�3 <���sZ�@�F�I�4+.,���KsĎzM��T��y\��^&����<do��|�Ő����|Ŵ,�K���{\s��\���Ns�19?��9\ �y���L	�q�<�g3����
ą(��x��'�͘J@�!b��?��[z&�6���U{ޮ��R5��a{�����$���VIk&��)��*��Р���	H"zo+,���z�\����}BW���0��F��������kﰡ��^*�\�v��S�{gE�i�F&��&�Þ0��*^�t��/,�e�f��i��=AD����C��K���3%B�sw)��Ȝ������-5cd�f��^�DXz��e7���3��5H�Ld�]�v:�n(�~�:��Eh�Pn���wNJȂR���s�ϊ44p��>����:OlP��5��븭���~ӈ�Eو�C��K"�Ec����(W�|^��
�ǫ���R�`�{&l�D
�k�������`�<2\'%eFkO�L��>���+��}��Ѡ/��䑣G6ܚ�v҅R�<zY0���
2=`��������	��.)'�K!��`<��%p�����Zq1��%b��f4�� ٛ-�B��#�f����K����H�N�����X���VY�9����g�������y��� @9��WD������O�B��@�������0w��ː$='��{B.��*A�����d�T]�T��3vc=�} �C� =W�)G4�g��%�?��n�� k��^��\�0����|ڬ��?��!��%p��I�0p��[l����^#D�>�4NC���`D�eu��#TKl:8��#w�
�UÓ :ܬ�n_V�D9"�
�KyZ�1�V�K�	�`�A8\�.�FqV��@���U=� ��KV
�AO�q�C8���G�SV����AGc�ߠpx���;J����3��u��SZ��#5���s�7�U��,Q<��f��˫ӎ��f��ry@�S��A}����i�G��嬖h�C�ļ���Q��aG
�h�Ihd�u(E9����&�A]��� ���}[w���ϋ[�k�Q07������5U��|�j�(��-�� w879LF}�$�WO"�t�N� 4��*sDMj惙�G��@�L��%n���B�̓��������E�������ꆸ��L9�8�j�m������hT��@�p`ő��OV_o�O����(e�xp����P��Y�[seZ��{�V����22č��b4�����#��i���,���)���Yn���`[���ON*t����Z��B���ߊ�$5�F�ɇ䒶rH0���#�aR�t�H�6�>��Fέd��IP�	o	�|�"�3�����d�@�T���{y��[0�VZ�!X�Ip���[&`��0F��M���c0������O��o�s	U�9�̮r$��G8M�N�dF��e�WNx�ʦ�P�Pl��(��xu0@�瘛����Pe<��D�8�}�&�O�6�:Gfi!��
P�w1c��'+9=>�sٯ?�L����������$��|#W��f���]�a(��L�=(0y�~:����=�j��*׶���	c?���q��s���cި�4�@,g�	>͎p�0����Yȁ�����݇�g_��4��n)v�gaOkA�r6QEf��,WO�lP*���;���W�>���[:��D�ƍ5A=�Q�k�OydjH~_5c����4hN�O��yP2#��ƃ����'�$�L�5{��������Y|�䐄W��H5C
80�!�-}@xE�LpW�)�����5Z��G������ʢ�Ku6����P
��9������X�5���Jj��t��89>�m�	�nN��a8���0�4���:Sw9�7=��cc]���F�F�6��jj����ӂ�����J�+gv�?�(r����3��y,���	����>��g��k
����6��3,��U�q;���ο4uB�~��='�=��;??�7}g`�=�6?9�[�����ʏ8�+B�����PuO7�6\oy������`�y�"�3��ӂ��f�|�^QӉb��d��uՅ��-	�F���^���\��T��X�g�8��p��c:��>ȥ���M&��l��@_6%=!��˳�HTQtw֞tћm���w�C��E�.���M� ��&�Ll�&��[)�5`C��Y���g�Qՠ-�g��`��#)�6P)�?����g8g�ѐ�����<4�)�lM�e����@��Oo���ʬ��Ŵ��	���b����jY�{�(༄���RO�K��E(�"�~п�W�,[�
�7���!�G}�_gd���V�U湏e��<����mܭ�������lv�XbӸ��N��Nׯr�BeΣʽa�Hk����S���[0�\;��6C�����e47����q_�kw��l�=���-K[�.�B��:�����\jbX�;7n�6"��Uݬ���}2v��&ܯ
�q��@�A�S;��u��%�򁏡�Z�ȍh�}U�->�@1 �W���+lK0�/�i0�[����e��t��1��lya�VO�m&���p��G��XN󄿛���[M�d~��߇��.��0��)I�U�t����(���'�m�0�L<����i�k��c���*�'��܉Ñ�LD��L>O�_g�LP�j�X���0^R<PWϾ�������۾ǈ���[�^���g��!4�b<�u@�Z �	�R�3�ϩ�P�7�ks+�'*\0^�Z	���G�mZ8��׼;_"��?'����DF,Z����"����(7�uV�\��XH����h�z����;��hT"�Gn�222�c���qn�h��U�@�u�Pd�����a���1�L}��@�%���N0vk�M�i�#�\��x������|�#pi���V'b͗씎h�s*���f���ydEe=~�W�I魨X�m�!�y��c�hI#f�R.B��i�'�M�Bސ�Vq�^���o(�!܊��I�,C�\F�	�B#ȃG���WnVy0�^6�����fW����ٳQ��.V���]*Z-ϳOnT��pՈW7CL�"t�Yڀ+�������	NT2�?+���h0�+&q��+p��<v� ��&�E�lV���Y�_z-{����ɚElZk\�nf��}��1I�,\E�&��uO�kkY��}�9�av�g��t ְi��u��#$��9���I!�n[�D�L�Pp6
M0��뛈�J��~,��9|W�|��+p�{���#/�U�M��"Cg�XfYL�_t��
8λb&5��i��|�F�ͧz�nv�H�$8y��������#7!�I(~أ���^Mi�_U��H���֑֯'��(��?�f���=p��U#?��L�� -K��Ӎa��<:�Q���r^}��J�1����v��O�Ǧ���f��mhꢽ��1{G0��pFH�ek֮�e�A�ܯӧ�bȫb�k��h��_��I:�{�d���<��պ�H�{߂�Hhx ���dV�r�9��jA���}z�8xKe"S*�즑�lU%��a2�L8x�;��n�#�ޚf���-��4��ݞ�8wܱ�x_a�"&V���kji>U��m
�ZZ�G2h
P)B�V���h��?�������.耄���#�	������|1�%Yb� �Tp5g�lY��>yIKlY�a|��봝���B�GA��*�ô�i��AM]�H�񤐫��)��n\2�P�"X�=��*k�v2��).�ĩ ��/(m�.�"�}D��i^,*�	�o^ƒ�����ښR�����'�6u\�tm���;�>dԇlq+bT���,I�"b�"p��>�==�_�d�N2�����������ΰ������ž�h$���}���RK�#wGhTf2#������h<�ݮ�w�(J?zA(�p`X,D���U���~'�rՆN�)ف3�j$��Z�� �&ݟ[]�=��J"��[��vI�jY���1m���Z�����ȿ���c7)]H�����L42��d�WìR	�틀{ٯF���\z�	�b��xm�b�y�4ri�E�A�Vck�ܢ�e�-����O��o�v`�-��(I��|�.�g,$�J(�ꨗ�Q�$nrf���'u��<E`O�+�ɱ��M���R�s��GTheLSԸ^�ks�5w��ݢL���`�ԩX� Oϡ	k����5���eeo1�,�nZ��=2��}�)*���7�;�+�MUd%� ��AWE��܄5j��M5Mۭ~_j��p�Q�?��w��Y��7	��Gx�
��OƗ;s�%�_�٨{h�Πm����(�0�G�=���[�*��lF+A����<���O��N�.�]֔��*�x���7��*[y�!F�W|ȇ{��[��O;�0 �{xM��Hh%�k�}�6�<0,���t�Z���2�Q�����M� 'зͫR
p�$�O���+
$_��U�F��t�8W+���|I�����/��-ɻ��m�o0�L�c��ȧ0��wwd����I�D%�(lD�;���a�����D��0�	�g~#Ij�����2��]�f����G���&�ӧ����Z�.P���$�ƾ{
���}T����%n� RO$����il���kW�_�������nwX�E�ey�ʚw�P����Lw��	m�:n��+�Y[~;�vY`{��4w�]�%\-S�E��ïzA܌�Q���٣���u!�$�~��h�P�]�U>ތ�P�i�Y�9^Dv|<^
� �1.l�d�����,��4c�?�1+��� 
W�p����+$X������E�4�/����3�H�
�*�%���X����(��<e���
���7OY]��B�s��ڐ)��V97\T'���*��[Wg2q��H���ļ#t���k��Tk�`3�̭~��縓�L�N�H��c����9-���L�䬠/���s�d-y�#��8�[�P_ID 0 �Ҏ� ����[-���J#����h����q�<'sN�(����l��T�nY"���L�]�Vak%�&񃖧��`�>EL��|���.��_��u��O���|]��.�7���\��(5�;GQ���Q��T�2=��_&ۗ��5;	�%*���g�R,^��N�Յ��/Eɍ��w��^*s�tAS���5���;�;�$b&ͼ@��~�����^��
����;����wz�M�f�!�(���b�Ýv�ub���=_�-�R�*Qx.H?�Ǫ譩��8��B���KK���?( C��ds�Y.�i��x��}�d
�4/�_𫐨���{�6�/��	��x�λHk
�^�'���eI�T�8�[te=����e{%HTR���{�VZ�Ia��|6�6��Ш�8�`���ha���	��C�et�E�3�5Y_��߶e��P��M1������J���FͲ�D w�o�����^�ù��J4Q�y��L�\���OO�>�c���� �b~[�VVm,E9����ȇ�i���؈��&�XB���1�I+���1K9��Kv�z?��y��J��>��������[�1��q���9����-]x��<+w�=�`1����K�20����L(,��֖�9����K���W�(�$m�r#�׳�bL8��K�k��#�Q-ӹ����2�;X�v�~kZ���wP��!�u��e�G�i]9BkW���F]=e"�;�e��m}�1е�KTM Z���%(S�{Ҟcv��XYG��i�J0��R��:Ml�P�k~� mh@� �ցFo�u\-�s�e�<e7T׌*�8�p(쌥��7���G��s����M1Ox���/aV��|*�A�;_���d�>S+�L6�S1�M��d<չp5�L�'��׸�Z�>��{��8���{��Ϙ����EY�IQ4��W�R���ƞ<��fiz��K~D��x=��;*�րi��KO�kY��'��)c���5��[�I$�x���H ~�#�1�ء���<�I��Qb3GA�h[�?K-}`�%m�o������&��|o���&�����Յ̊ ��Tp� ,�h$�zaG��n�L5*�j��~m��B���<��K�!���S���r�+�z�J��ٰ{��Z���U |���KZ�[Vb���p���n�,����Enm��L->�}g��1o"��f�̡��=�Nֽ �em�Rn˯�w�f���5^BW�&
�tk?DU�t��_�|��{�Q�K�L�	F\t1}nC������*��vn"۽Y��R�-] gih�d� ��(0�A�lś-�0+�g���k�� ͎�#Տ�*|��
�D�GQ�2��H����v%-E����+��7?,�yC:�