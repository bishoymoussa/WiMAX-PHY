��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$Rx�y�<��wA�*;�x���@�̦�W�X�fa�M-$u����n~�%���P�$��W��kYَ���P7�?UMfT��q�6�U��k�>����~�\N�(�����X�e���/6U|)�X2pF�]$h���d.���9E��WG��L�X"]�Ad����ľS���8od����e�GT?y	7�������ݵ�^��R�q^]�鍦�����s�ae���h��L��P_���ާ��YЭF���'\��68�b�[����w8�[X��V�F�0͘3����q諵�uW� �h�u\V�?@��_6G�_�*�G���B�絉�f������[�G��U&�����~�F��AׯK1�`c��[<��FY���4I� �#�G��x[X�=�Q1��`��R>(�w����R�O�?����7�,(�H\�#h(W�EH=�������yq��Ѿ��aF����:�U~m<|��.��0=�P/���4ǆ���T(����T�����)L#G�Ƀ`�;�.I�����<1[���^ï�$p:"c�Mgu�gP!.^��i�jj��͜�e���҂�S��:���$�[��"�9� �Q��+[(�"ᩲXVdTC��i@�H�O�T^aaGǱ�P���RF��(Mk�IY�rA�O��w��F�r�@)�B_U�;�@�w��c,��>D�k֡6+�Xh)�S�hu�3|T�mx��/��8�Q�$�؝&���^D\��etZX��i������y>�:��H�+Qn3�-rm�$a�y�l�>B6������`�T�����z�ɴA����3��P�k�F�>�������������ڟ�f�1�����ē����/aKe6�s���X�K'>m�B�b?�[�
��i3&)��4�l�=-��"�n�H�q���T��>��Vk����aˢ}(�c��q9t�fn`<d2Eĸ��������A(��לe4)�nu\�(f;C�itMd�Vs���0���zSu�O�E�G,�6琯}VH�(֖^Y�e9��b^���{���o�������q�K��{��+ԫ�����Ll���Kk\8ʚ��	���$E�� ��QT2Z
�]*�Ok�G�
��0�Xe��&��+����e�]=C^F.y��O��n�A`�����#]�I��ꞆfYv��M�q��k�>�F���V5L��gڗ��!�V�8��SRAS����d��+�k�����Rp�M�����������+�0ZЦ��3dSzFv�,��T/�K��& l�?�zu'��WC��Bc��#�W?
����K1	;n��(RYC�Z]4D���|�
3K�k�-�7�aCyX�W�[m̔=���T�K0˦��J���/&�cA��)�oH|~Ex�լ��}�O\nX���r<��J���:�x %Fu�e)�jߏ%	|�7s������2
c����p�;Yԁ��ܷ��B�X�[�=����+��b�
��I���{37�/@�B��z 5��@�[�^�M�-%�Z�k��%l2b�O��l�/� �eG@���Tq��Mԝ��;����J��,�q6����^k�#�Y����AQ���s�o�ճ�E�@j��I��\{>wRA85���x��snPf	�1�.�&��L@}���FFNǦKhK��YM���\�P�Z!⼂�~1�S*�}f�?ؾ����lIr8ĥ��X��'�&@��E��fw�@щ���?o�O�<D�4�n�q�&>$�{n&MUG�N�G&����x�#@%t�:�o��ȑ�j�Ķ��A��
�*��2@���z�H2�V����n��%h�'�f+)'����ʁI��p��Q!��݄�s;|���u���8��*�K ��랆������INxR��.�D�j���n XʚV��~�����&ۛD�<|�j�@[����C�KsAb��� dk�n	I d�ʘ���rxv`5��s*Wl�t1.C����ݪ3�Dzn����r�0���%Big� �[�đg��<V�:W4��W��������F�ă��`�K��7�w�w�,ߒ�]��������R���
��)s޲CF�� _m]P�Ek|�XK��;��P�`(��OO���wd0����\������.�o8z`��c��d
}[ۿ�[��</��S��A�R�����@x�̭wh��\�_����]."|��L�ԋ��tig�K�8%�a������9en���ח��%���A�3�-�j�}.�G�6;�
=��.�4A,�����'�0��b�7���F�/��O�GNs�f�y���P�d�ى��S�i�"��S�	�u\�v��(DGx�ifڷ`zR���A��jHT���G�5(�F��u�l>r��˨[�=�<r\�b$<_Y�c��8���FPb���D��}�?o��s�S�����w%����h�V�����cǷ�F�����b�,�ƈ���J��K���6�]i� �E|Z�"/�Ĥ	�8��e��H_M�u���r\h�̏цU��k���HC�Z�j���j�7u��{h��E����I�[i%VnmR�2�S-2�ߖ��(6q,0������p�<z��i�9�����P<��>0H;��u��dwv<��Œ_�j��;,>���9�pm�r��i�?�q}�����z�_���(�Mg��hP@�X��]聢�i�e�F��s���`�Y(�_��p�HZ֧$�X:�'�jQ(��R�<w0�]�Tј개�ZB��3]|h�z�|P���zJ�m�����V��4��
K��:��~@s,�B��B��Ü��/(V<��sݶ6Y��7n����"NzV^�֐�S�PQuI�����;��ۙN.��i���������o�Y�Z��|�������/z��G�H��xXN�͈i��!���ucg�Q�I4`q����X�]������\��4�������DCt�&�C�$vL�yvT�U[��Ydc!f���wu&��Q��s�Un�S@�g�{�)+��J�и�+!�f<7���'o����O~�䍺bg2������d��9'q{�-x(e Z�nfH"�oV2�Xn�q��*dQ�t�.�d�xy�}���AZбRk�2�
g�{�/�*+f �W{��[�������}�܂D/t�"!C������5�k.{��@�Gj�Z��x-���[D,�86����4j�G�k���%H�7�S���ښ+��)�6Y��:21��"y��ڷ�r���dmqc�ߏ	�����5b�a$�yǟ�2�b���K�Y��2[��(�$ ���� o'"�E�	���Q�5����kc�e�P��5�!Mռ�{���h��.�;�	��
l~�Ɂ[�j�-��F2s\��E��̼�\7ܸUM⊟��U,P/CA�����b�%s����[�K��K8���,�15æ.��@����9�<���Z�T�0Dv�>i)��d���� Qf茧ʏ��,.z�$�ڡ�1��[�냍pzx�&����H\�_*����v6���^#��)�
�cT���
��ɝ�>tԴF���h�C-hj�u��E��*]��}�����y^�g��s����T�ME��