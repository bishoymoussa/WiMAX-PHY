��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$Rx�y�<��wA�*;�x���@�̦�W�X�fa�M-$u����n~�%���P�$��W��kYَ���P7�?UMfT��q�6�U��k�>����~�\N�(�����X�e���/6U|)�X2pF�]$h���d.���9E�g�����	bI�g��ȆDE<�篙qU��ٙ�����`�>��
p��Lż�u� �V�s�{E����E�E�wi��(���T�ǿt���܌����Wv��jՌJAI����6ã�I�A��0R=���Sg��CO���Q[ҬU��2eh)v�u�JL�P�;���0ڵ��}�{��� nYd�K3,��  ��m=?@ჵ`���XG5�w�?�p�y�u5�)�4�o�'� ��/�z���:1��p�o���:�]6^����c/!~����V De���@<I�mƮ؃�hj��t��7Q��N\�t������wG�O�W�x�U�����<|/`��b+�8�էr�c��~}�8�n �#�Z�I1�I��르�f�L<ъ� �� ˀa�4��9y��փ' 3|)մV �����P��m�AWo	�J�T_���6E�P�D��V�σ�-2y"Ts��V.W�h�>U���xFj�����/5+�í9m���u��ĉJl� �$@C�ɚ�aea��>���k�t��l柍��!%���VUWq��fIres�0�m�o���i����X8�^��U�]TU�{���v�U\As]o��f~D]�mt���
�q�b1^&4�ڊ�
�[��&Aԑ<	����
W~	(p}��~&	����f���1��Dm]�~,:e���n�2�@k���9����|UcRnzy�:�!�(x���eIBhdN� ��e���cr"�t|�SSt�'�Mh���"�E��Pt����V���f9m���1�08��m2ܷ����rl�Y� b;dsE��kd�Q�3�?Uo�����tD&E��ZI�I�P��!�b,��EU}�.U_����8m��'?q���T�7�:�JF`���6ֻk�-*�Wԑ�a�񷯁���Ⱈ�����Me�k��&���iS�˟�!p�JO�JF�\%N5P�J�ڟ$d�@��^�z:@YbI~�K=K6M�7�� xǊ�*� ��r���G q~�9��hTxT�d��M�E��TF���m4y!��R���桞8��q�"?�E�<� ���:WUu!��qV�_D���鿉N(��!N�ѯ����b��;>X���kf�
�f��[�%��9J׊T��\'��E(L��d��������[: �\VY�a�WX@D�3f%�ø>��k��㠦���[mx��k���DD���m�C��%�s���h�ytoTsZ�^���c����;I�}���!�{8����7_��j�o��À)�lZ΂C������[	���B�ep�Җ�|9�ng�s�A��4�B�پ*&o��*��|N��4�7�A�J.���
^� ��g���еU*}Xٟ������)��ybI���a8���&����;P�LƖND[S;+EB���w���#��J�K{�'�Q���2���MN�Y̟P�NB��@�X%wX�+WD���o��c�N�saqT�4u����Ot�O4�1�T�۩�Y�p�ն�"��_B�Nd�[���nMo�nWk�}�,�4����2&K�5���������y,q!�����k��2S���'ڮ�����lG�C,�؃Z���]w����g�4����67%��+!P�Z��'/��A����ypŉQξF�T��JL�Z"�f8=zz��(cKa��59t[O�.��o��WaYJ���K[Y��g�(GM
��b*!�(gA����7�(R��{���7�9��'�C�R��d�dOe���0���W��R�͉�<��n	�qOl���Y��>�s�>b�;��>q5�a�t!�xS��o��+�z��5�"@�G�N�Wdq"��\�kW&�#R��Yzm�	?�-�,w��5�Vo�ߚ#ΒOG��1a�'�%="<|^L{'��#��j8E�9cg����/�`o�.�7 �J�}�:/1vf�/�]]}�[[�f�Cp1==m�j�bo��jp(���}�v�u��Oz��0�D��`zJ��;�>~H"Y��Iv�����TW\ U뛐7�P�����t��8��� K%�-,�f�M�ϋ��ǘ� �;ͪ$R*��⾛c	�L�$)!��؀<��āM9�{��=�>��9�,��d������Y�/'�xm�%��"9U��S&qCs�ZR������%���_��lƵQ�vrgaV��,^�Vk��I�G��x�1Y݁M.��p�9?�d��Ɖ�B��@�(Vm� ��U�.�8�B.#��
��b�j��\$9�#�@t�����l�π�!Y/��H��{�u) W��'�g����D
��9z*��.d��]��N�	Ωcҭ)�/n)�`�Z�%� '��1�O]1�f����պ��������j���EAv����Y��z&�kƌV�:�0��RЧEp3��w��SAh�1����e�̛�Iɖ$�)b<��3���c������%6�U�s����#�����*� �[e��곣~@��s!}��G��D/W�3UƷ@�$����������0,S�%T��K��<<ԇ72���T��]$���8O*q���
�+��N~��o\<����b[���?ádo��c�6�����M7e�\C6�oLj�w�z)������=?��K���|�<�e3R���i�z�����i�d��tS�^��%N��* ��52}��[��r��۸���Ԍ����1�ט�.O���V�Sgn�dR�0 �z)�����Vb=_?�0��2��.&*P��fYŠfl��)�l�U�0*�K.�kZ	k�Ǧ�⤡���J"���y˻׆��$-�v:	�	�AH�Pڰo� 2H�.^᛾��E����*���~.�C�Q����	���OW�X��6?��\����P����8B���z(Q�r�ʣEyƘ��H8S"c쿋��MGMlg����7�u��~</��˧��/�fِ`�9��T,��{nNQpB�̍u��~����Ț��e��h�]/�S����`�$��-�����%O� &���\�M�mxы.�*}�jiE�B��'��5����@�Z�׸Iy��<���@KΪe�$)�h�x�������3�Vr�s>G��c@P~�N������0h2�����M��)e�g�<���Q�����ga����t��x15��MPN�O�$f��R)69����yh���������5���QcB43
tv�9^ �n�7O����1K�^�>���o<���'i��Ķy�����n���%�Ձ����쯷D�����Σ���YO�n]M����z�$�Q��t��!+>��P!3�������$V�7}NH����E�3(0� ��;��­� ĥ[�+����]��	%��re�^�8�/N��9P�G��hI���<����eUUZT?$7(�-�\���5g�1�V7�X�˧=I�1йnW-�8�B��r�E�	�_/��?��	��c�����!'��c�#\���H��ww'V����]8�S���oΞ{[��'�{�>W���'QS[�=�o4�+�E�p(��� 0��2��hk�`�6w௪�}�O 3/s�t��S@fͩMx�W�*�@��&���\�1f{QJ|L$�He_�`Y���S淀zW�@����>����Ԩ������hz�~��;�T)�:���"é/�j���T_T7���bcӔ��݁O1R�{�G�e"�E�cn��_�(�o����r;8Q[��0^S�'��>k�k0$u� n��ߜr�/��@�y�mWDѠd/[>CY�ZJ�5�1{
�B�p��� ��mn,"v����]���n'~Μ�iNJ��jD��S�o�����,|�ze�����#�k�.���(6mBEEI����.��7����%)o#~N�ʩ��8�ށ�`j]�o&�m�C֌~����
;����5��u�T�v�}T/t�����F�������;�=�=_��B�e�q��������W4�����T,y� ��K�̪�ü��l�/�S���Q4�%�*U�s�bcpw�.?d�Au��z�M"Bsr��
F����-��-� ���~�a����-V����Ç��� 4��ő9&u�W�S����3���!�����4�I��T�ar�aD�2%S��8*ҵ�Άy�^İVQ;�-@?K�}���¼>�Cz7s|�*��ip!�.�n��_�`���J�-$٩��ܿ\��dX��Y<�s)���=Cޓ��4�J��f-�pX�rV���Z��'wc����h�&W T��X����J^�V��Ī�=�N��7��'s@�2\��3y��N�/;� pvأ{������q� �m��ġ�G���\9��3ܝ����#��� �^:NeA,��o���B��*�)��,=WL�;)�kp����U�e	bq>F'�~�]`�Y�}S�����G.<>��1(WQ
���&]�ȝ�~��qj���8��*���q�v#:Q�~t:b
�]��Y� q��#�):V�ױ���i��|�K�:(K����60Yg�V\��t�/2t?>]��|�"���[��8��yx�^�*�e�&��2��AV���zg\/�q�W�+t0��液���A�[%2�u�4�2+لc��=V�wv�3��/��P��[4����v`��Ns9�p�JU\���Iݮ��ۻNp�a�����{���������
b�q�@�Ps�ɶ� =<��Mp�R���q%p9�<��/g��#g�}�sJ�63�?Q1x���L��z�~��ֺ ��(1׷�l���EVŚ��9h��; �8�S����v�z���ID�f�C*�O)M�u���\�����x�1�A��>$���p��abn��ڨ%�[I�d�jVh(�6�А{Mf�VG�_?��T�ww����f��$�&b����}M���_'�}�~~e�d�UV��Z�Z�n-zq`��n]��,�IL]��`ܱb�WqP3}�S�ǣZ���d ��V���b&�X�w���I+��(� h�)<�S��~j�z|#�����!�f^#͇2o=���:�!1�)&R��N�J盦�P��(6�ɲ��/E8��c�H�L# ��k�^�6����G&��m�ռ*��Ĝu�⻴aԬ�3oB��o��,[�?�ַ
�hP`;�U����  s��J��i���z�<P@W�ҿ@䘚��]�lO�B�Ij������BA{�ؐ���<����piw�X� $�޻&��]�h���t�g�Ĺ>�\�h���������q��sj�p�gU|E������T�pf�t�9r "~$)F����&�5�ȦU�S`�"����E�{�����8U��&H��R����Q:�jhyT�2"f�38.�g�Ά�d�����A[�xi��b���Y�ڴ�O6�e����$��j�uX�Ȓ�엹'�����B�p�\p|%<7�(
<Kc�!�ڷ���K^���X�Sn�Z��bhQ�f�ގ�W��BK48t�<����_ww��}�~��x
�&O#��r��U�b�Z�_��́�{��j�yWf�9���qh��V��"o)�Si��
-]`�D�//dOJ1��C3ZE��:�_7��e�G��vQ����>�4�m�<ju�VE�����!�,])�"�^Px���ǡ��j��f`�:0�[�w�S!�z��k�<����D��t���,�GD9j�>PW#nB��"�x�꫶����y�Þ��0`��D��_����81�>!�x���	@��뢤Ѫ��HǍ�o���;m��&JnE�-(U������4��mg`�c�d�2`�[{��l�f�؄�T:�s]��M��^�hC����U�2?t�-��z�J�T�SW�A�4� ��eR\`�c����	��7(��Fl��yL�f.�y o�!�G���r��Z���_\��<Q�/���^�-?���dw)v*D��!�CB���ul6�=���`����e�۷~�3r�,v��p���vz[�+z�e���f��9^�-����gM<zO]eJ^4��b~n!�p�������c&V��lhtj��<�%B�AO��PB��c�C�`���Tk�p�:�Vϣ�]�N�i˘6-��G��ǰ�j���$=�iO�_M�H��+��W�]�\A�H�KV���1�����ʩ�ޔ��ր�c���T�{<y�����iCxň�s���V��dZ���(�_�y5U��2��W��n�ZȻ]5��˪�e�V�(T�0d}��#k�&��X�|`I��mVQG�u��4��G�"�����BPl  �$��/�U�e3�}���c_��;������I�����u���~��ZY��7n���T���1H;��O#{�Ea{{]߈t7+��>�RWv�f'���ä`��X'y�8�ދ0;s���(b�tC$+sB	���n���#���/�X���.h � ��SA���I}��7�b�^�DR���s�YG._�2k��	��=��QB��W̢cqh�l�3�{;)�x��A����d���l�/�^�,��jK�c�[�G�?��7�`���X�8c��/XE�|��ӝ�N�ڕ�p(g����a>�o�E20�w�^�@eLJ��{6;�,缈G��u�j�X8H�Oߞ����7-~�9װ[uuvh��H�K*�y�D%~A��(�^/12�Z!:�E$V�a��"���e-��"!;	g .��L׎R�ք
�e���k����l�'�j`?{�fͨc+�E^OR����B5+[�h@�f�鰄�e�y��L�ܷ�T���j_�̢7
:>���QUl�|.�/���4(�x��,K� ,w88a���wBmJI�� �mK#������U!��4b���b��j�KOmx��VM�B+���V���T��gh���Y$�V��Fdd6��	�~@�Λ��C��XvU"Q�p�ܸ����	,��o���jc~��5��$������U����8e�6E������5M/���Wz��u<�~x��t�w�4�=,;��c:�֛di���6y�!���c�۞�XN&�������=�y8�����M[	bS7	����[a�H%D��1o,���y�0m��O� �V)�R	���ж�����CJ��oA��W������X����Ȑxв���#��:Nk�� ���{R��y2
X���5n�U�T�CU�f݉v�.�7��*�q���<�,��1*Nz@����(��)G'����%:)��^���{�����b�V�q��E.��5�h4�� s���7x��;�(�ϫ�k��N�W@0�|:���l1�d�*���v�lPI����7�@�X�ئ"ʒw�jH�>��MK~������}�*�_f�ʭr�����p���U�HϚ	�Ow}|)�u��[N!y}��������?�R��*ȑ[~�8���O�\Up ���#
`7����Q�<��;�M�ss,ͱEYL���`���lz��}pB��!ԺPǁ	�K�K�%F���=���r�=���p�^xj3����7J�owH���?<���M�&	�A��#�)��~[��V����Y�P�"��|W�>5! ��v��*��㢶�Y��w��}b躸�\9ƝKG��Q���_O>-p!$�#�\rL9m�3��~��V���2��2��,�/�*4)�d��z'Dd���1@e_�&/�l��k��"����=���ZW$ǔKU� ��G���(|QDY�uʔ��t���O��1ґ[酕C֘��Ѫg�'�|�M~�`���\�d� /���^��" ��ґ�@Y�(6�|��i�	��Q���e�'�]hy�U����*�=j�e�`\��9�;�[fR��|��z�0�VYIk
�c;V�Y�ڈ�k #�M�dE�I���ݬ"Q�Q�-��Α�Oq'�dyԊ��/�sp���ZfF+7�ݭ���.4t�q+��ݶ<C��>ᝋ����ۢ,?�t�~b�kh�[�8 �3��z����D�Ɠ�o��W��~"�v�*�"ҹ��E�m�8���W�W��n�YA9��kn�Ѧ�������+��M����k�=���0_jg�k�J�k�v~�@�?�|j�<���OKϑ���^v�^���l�����*�Ҏ9������H�a�M=�������!/9~�;��I�HC�;pq�Yy����9�B�� *�Af��`4eX<��e�׭t�P���߃�E����jS�Y	��N��C�'�Dߩ�.�Lؾ�������|_3�Bm&�I� q$��C
�[���@�d̷h��<��Qm&�5pD�W�np�ȫ�J���!}����Dpm�N��}�P `�6M Ր�:����ML��#ۓ�l�9%�������?ON_�d�+҅����dd�!R&��-�n�P��*.k�mty��әg�28dF>fH.={���))�=5g��(A<ڂW�AL�f�X?)RH��Fj�W��SB�S��F��ε\[��{�⊖Ԗ���c��Nã�Ӗ_�z��zФ*�i����-��dQUՃ:&/�)���m�+�Ɯ����|���S������ʰ0�J�æeF\��zɬ�z�/�咁g)��kȋJ2~SP��R���v�W"Ki�#Q��lɣE��>��'z�  g͝4�w�y{G�8��g�"�H,�^�zE��!q�c=um��o6g,��N������}�!/�uސ�hi����`��;��#�,m�ɔ�)� ,�2u�#���=�G!��CA����|5�.=9/�������x.[�u_��K��r�oHYh�x�2(L�ZU��⣣6_�|�v(LoHȲ��Z���dCf���:��T4�J��B�� �iB��;�)~�'���d�3c�5A�o�hO�-l��f%Ix�������g��n���h:0����|��v&�lYT��4����E��O��6��jX�	�t��/�sۡ�O@nJ{#. �U�M�'mR�4��P�V��@�9�BV�9�9�s7B�a�)��+��5��+���0��2��ۚP�k#d�U���LF�1Y�u�Oc�|���E���!��G�ˍY60���gM�]����"1�p4�!�#���B����e�Z�k��o��\��[T�ВU��W�Rw�:jǽ�̪���������@d���b�p�
k,�!���T�><�^��Am��#Ӛ����7��࿧�P,8���s��S�T��,ה����6
w�%�\Q��AOO36UHXa����=7��?�7�3�A�l��wWO��!�>���J�]�@�o�\���������j�SJv�6�KB+�ۅ�NE�/5���)c
P���T�ϡ,�#^��[��x��Q`��+}�.���6�m����8��x�� �>�G�5���DC�j���Zꯔ*�[��Y|�~:Cɲ>hx���D2��`d)�e/I1,@���Y�?�K��d����QѶ66t{	��gc��i�����C��b���ZDz��ر�a`�_לA�B���T=�)C�d�Y��2�u���S!�p6�H_���$�/F�<0K0a�u�G��B�� ����|� Hy��r��tś�~��D��8V��+����77���U�S˩�1įT�����(�K�S��C:�!CX��')�I��;�̸l���o�|��(�;�Zr�U����+�~�A.��wFq���^Ϭ�Ъh��f�r �e��M�����$��}�w�3g z�9�]3�����)n��m6�(�xVH��T1-�蜈���yO�ܫr���QQO���r�qAbLUc�8�����8��n�"Jnidz'G⁞C̨�>��|Q��C�L:�&�K��^��7��= ^��i����Q0��B�E�?���;"��i`�}3 �})z�F������29ڮ�6�8l��ֶ@���		+��䮛���������� :1ۯU�hȄ���0�u�凉�>���j�NOs��ن:H�J���*'IgD�y�I^��c��0���-�� VY��Q(?��l��}�+��UT �(�Kj:a��y���I�}R]`�XҊZ��;�pׂj'���㡚,ԥ78}Z�2X5#c�S�('X�7VDBQd�
�:l������i�W8С�ZK�+���?���NL�����(�9E�,85�B ��4�1�_�鿦<�5dO(�-u�w|7�x(D�m��|˓v�M"�nT�K0i��P�gt���]fC�h�9XO�T,�)$G�ri�([��葒�a��j�UZ��& R��F|v:y]Z�i�:�D4 �i6��槝�(����Y���-�~)��o n�'�F)�p ���F9�	��� ^q ߀�����>�4J���h �l"F�%�+l��)�p�yK~��f��5�����'����9�C��),�0���G�����u�*�A։�z ���*������~,��9�����j1��n�j�h{t�b��c�G+���!��G��w&Ht��I���x�zۙ�`�X�v��7K�A�t��n@Aj�R��s?H�|��CvR�U=3�s*�+�mE�~�7�/*N�~�����]�74��`�IW�������,�u�aؽ��Zgo����L�JCTg&��R��g�����]���1t~���Pd��1��N�Id�Eܱ��j�m	C�����! QO���{,�^�H&�m/�:b��};I��󲧭���,Qz������w�����b�C���O�`�V<IQ~DY�l<s�K3W���P�4^�&j$�<:�H˚��d�
�#��&n�<�{4$�?��Ƀ���%?�]��cp��2���0��[���5�iXX�8�p���%X��2[~�~7dkJ�uԨ�3w>�X�X�?�8���&n�Spč�\ٛ����*�E�ƺ�Nw�A�3������gӍQ�ݾ�Wx'��"�!5
oݞ�>�z�W����Q̙>�n�^[���SF#q��1w���~䄄O�g���H��w�)*ȗ��	X���L�c�]�Ep� �o�1m�䢡Q��v�=�`;�\;�݇���r��`�֛���I$��C�������s���g��&��&7immFj�x��gX$~�:�����p#%������V; <@���Qr� ���>�l�!*]o]2��2����q{4o�?�²D��e�I�rfXZ}ا ��<ʻ�p})6�8N���J�}`���C�fi���9D8$�0)�&���:xY�r�8ey�$/a�t��j��R��|�O��~n茴k,����(޵Ĝ����ۓ�͚r`b>�`�v���濰s��V;HٮN_ۛ)�!�N��	�l��U���'C׺=&E�T(���m'������es�R� 
9�0�}���{�;X{^��XЉ����'��^e�t*�	�(�c�/��Wx)���:$��a_���)�N�ꤣ)���3R"���Cˆ�c�a.��3�����1��!�v�5�=X�@!�
]y5{�+l�j^��[)�<�K_�ae~�>�{�L&�Vw2�,zV=|�e:�0�9&�h�O{�uF�N��{�Ghq��}}�\�ȑ���d&��D������$V�h+��Q���2K�~����Q�fk��譸=�����
��Q	J©������F�O�.���'p"aeU�!�2Æ���Yx�'�z���z�*<�%�C�~/���,�֓}�@G#1�>$���Z��7�R�q0���_��u�p�nW*O�c�ᩳl�k�4�KxK9S]�	���_R�Ij([#F�O"<M9�~۝Ri�����e#�S�f� Y����D8��ϙeI�'�	Rd7��n�o
�?1h)��C���-�/sN�p�BÍJ�vҀr���{�B���9�a4�DoT�`E[o:@�� ��Ȧ�M����E��  -/[�]6�X��o��uL��^ru���k�ڰ���y�B{4�v����k�BHʜ�Э�#�-eO�s���Xj�K7�`ި�pwV�֩8"�G1��'S�(x�-�9��SFT,�-)�]Q>��ژɰ����X)�����IIgt�"�s'�!gJ��8J1�����P�k�V��8����{�c��g���d����hj0�?�wV�r�+�M�����b+�1C�7܆�^ ������u��F�=8�I�>d����XF�U��"�[E�������z��W�ۏNo��3^a���e6����#��O�܎|	Y���%c�#B�:��u��'�����P���Ԉx��_�W�xr~�>@���j��jq�����;�Qm�5	,(տ|0�0kq�7g!�d�Du��x���T?L�2)���_�7۬�-�m4�����*����<�����ӟ���u�ntC]s���K�3�Z��T+ �Q{����+�NJ�Y�I���aD{J����W�#����|;s6�?3�f�$Q�9�;=5�����P�[�����T�v�����܂b�X��Mcq���G�;�v�����I8	�ȚL�0�m�P/��S��  �C����&Q�&�/6׽���cx~o���Lz���	�>�59��"h��B(�MbR"L/�9��
�F�H�*6��������,9�4SH��=����iMQ�;�/�%�{�.>WGp&��x��z*Dk>���%�|����HO[��dȦRd�g�߃bM��$�N��icr±x+NJ�eC<Pt�*��Q�Ԇ:~�4���V�·���OӘW�2�x|�T:�C��(`�?������:�0�
�O�����,������ؼK�>z]	6�Z��� Jq�;o�ʼaEqH`=�/I��*}��u���	�v��t2�/�T}wK��
��3�􊖅����a�iB���D�{s�pp� ��K~���v�+\\>rG���@�s�ú,�"��sFb[��g����ړq����<}+���A~ ���:�����hԢV�٧ssW��W\�RǑ��+�����t�m)�y�������n�HGb	��N����3��8.<S��n�������^O�"{a����^���pN�<3BF��Л������H�LM�mKms}d�CB^�e����{���:ҬLh��C�D�@���S)�l���\Ce:I5� ���N������g%YOJ�>j���zND���P��uK�6��a��/��	����ʨi@�h���Y�-��Sӧ�'���x��J��,2��(p�b[�n(\�rW�L�(A�����MkW�'_T�
:�𫟦�l���&8PRx6}n�g��[@�G`���f�hĈ7Vѳ(�AQ�y���V����IQ�U�L��v(c��h^CsYV������kx	�G���>2֨AbY������_���ƪ����ɼᾃ"�vڈ�y'[���gdw�2�ݜsl�6��5ٌ�\�(~&r%��ww�j˺�9=5ĢZu���p��Y`���\��,��T�X{r6��^{+�,�,���苩�����n�x91gPY�Ϗ� ��$��
��nE?�P�7;�"�g-,�n_���ͼ����+Nŵ��n��RЎ�=#��P���`蘶v�|�do50�M^ΦiC=M(4�ɍ���w���8�r�)]E��c���(�[�0�~˄ь�]({3�c�����F��p`�� �8U̚�t$1��[$	#�$� 1�2!wV��Lؖ&���U�rn�u����ϱb&M<�����`������7��H9����>�����K��ɨ�낇Ln�<o�7�����So��8q�$���S�am�f�8:$����p�j���(��h?����?ٳz��S��4~�O/�����@�"���
�}
��o�-��풸��.�ݎ�'�n�rS���S�YE���íY���c�RaL(K���(@�</��(��e��q������E�{���	R8Yt�&]��-�	eu�_�j26[l�@M���l�68�H�]THz���Btӿʒ�)��"�+}���)��{��եw|e�@�Û���<��<6��������,ѩ����G��Ǘ2��f�Y��$Bq�L��<ճ�;ZD���>�e�=ޠ2��N�r��m5m��bcx2[���H	��	w]����f(����Oν�+j�-/'�
��7<��F�i�qﬔ��Lm�'�����U !��j\%뗻|,��D�B0����R;��btF᮪D�4���WؙQ�ĺ�.�k�C3A�a��ᘲDp3S�|��e�N�O�<��r�,ǥ�c'����y</�}Ԟ$�\�HNf�U��@p��� Wu{o��,(}՘��F;���r��8@��r+-|����r�V�t�����O6ݥC+:#��
���F����7O���zOiDv1���+�j�G�B�/v|Is��@�s`uA�(��l�<s1ה��z��n��	�>m竸Ч?Yu�"�ju�N���.���s�W��G��&QJyo}P�fxH�g% ]	)b�,)|uy�	����5���W˝ܤ_�i!U��N���ʑ�AR����ܠ�Cvi\�j��"�C��u��yz*�.-�m����l�B��(yxi�À_���t0RB����
���y|ޏ� ��[���Gf	PF���x�:;X�Ixaߨ�>Ѭ��7�QC���?8�/;�����B�����S�LJa��)���l{�p�=rQ�<�C�`��\>+�U����IC��ݡ�f�����hS�
���]5 Es�B�UKR��u��O��+c"������@s������.-W�N�'�@8)��Z��$Ql�V)*X{� �����n�
6��G��R<p��類�Km���|���i�&�|抐��/��b�(���G����FVr?�zl�rC�h��Ce�R��^O_�[Թ��X%�v�X�[gd"�x��W���b�3�W�����iëcR�I\7&d_��\Qjo���6�z�Q��<O��WOj�1�-�A��V�$DG�8�=G݇�EN����&8o�450!�%���H�P]��#��Ì�d�>`C�k����ܪ���Wv;�+�B0!���;�Q��C.7e�k��J��8�	 ^�2��X��\�.����y���S�(��6��s����X���ҹze}�~�c�@P`]�IH����X�������� �eP��6�Tc���Q���t0y��)�����������,W�gh^�ӟ3I6��z�SHb�����T&Rم��"�Kl |5��{� ��ڣT�)������߇� �$��$�;D��A�������!An#@��� �bx�p���a!Uz�/}iFa��.d@*�����Z��T[;��o�(��X�b[]y�����ϣ�As���W��;���d��b��1>��S����a-��?�~��L��S�+g���E��"��T泻�4���Q\o�#N��/��@�u
x3j�6o�h��j�Sa�0w���iQG�q��S2�ح����Vuc����Q@��'Mg���3LC����^�e�Ոx����N��]U~����w������^E���@�[v�i(���yR���͖r� ���㡓˩�L�._j ���|����qJFb��9}�}|����k��s�;�J�����EB�f6��uX�w�SU�x�|d"R�2Q����D��1��i�!�3��Ԇ	G_Y�Z�s���U�ρ��ֿĺ�LF�X����a���!��!Y@k�ȥvk�Q<^�ŕ��=�^3cOE0{rk�D�N��G��mםQb�b�Q��ɫ����w並����Y]�2#�&����9e��.kG��@�Ic�`�mM�+Ki�sTm}��hd�=���Vq�ޣ���f熯&�w�^|!@��AO�!t +��AE�%��p��S��iLs먩l�����K���$؁!|��ڿSJBh}GLĜ�gS�6�e$�%�,a-���$�r;O/����:#38��iub�a7ʘM�Ϊu-V������&�ȅs�����_ԃ�X�4^n8	 qu4�܂)��# ��N�T�7E�
���ٙ��/���i���)��Ӟ��v�^'H3��s�P"g"�������|�<f-�������`���Se�j3+�� �sf�`�ԝ���|hG�w��6D�+2��1��|C��7�t�LŐ+��UJ�����bM9�?�Q�ɡI-�Q��Q�-
&p��k�2o:���8�l�q��,<�*�k��]&H�Oc�6h3r�&��Y����oX/���ְj2�Ue�-�JbT2+p!����f��}
���F=�� ��h��%_�k>�i?�.5*�h|���p�vp���7{�fqqD���Z�z��E�Y/�&�T{c��|���0�E���TAcYt���z��Ząc�՜ٽ�9�l)��ؔi�8]�`� �n�
'{L��9O����T����mo���c#����M�: ��
������}�R?j�j�;9Rm����+ޕ���Y�w�"�ͷ�'T�Ԣ%�.�;f*�Hl����و@7B0�M�e�}��COW״�r�6
7�D��evk7i�$܌~�������E�y�m�����U[������A�jT����F(^ʬ�(�RE�*0��L�������YT *_E��'4�×d�B��{�g��.�S5e)�~Z}�L�J���C�> �kom� ���s�7��"q��Uv˪�t���mn���5�@S"��j��@�����W�mQ/�:������]n-W}*t;�;In�B��d��V���b�_�%��q�T�v��AВ�95��,�{�N�_��Nn��B���%3��puj����j���H �ю�B�O?�,���Lo_T��\e�1J�����@�6�+�|
K�q�;��5�r�<(h��-4e�θ�r�U�i+��sv���B���uGUh�H����o�;�����6=u�#]��-d�^��]3焻H�5�r��5�ЅsF�}�lk���E3�x�Yk�r懪��z�iN�51e�<0��R���~WK%�K��K8�y�Ўћ*�D�P�k�x��Ϧ:�Y^"9<�e��#JQ;SH��f����/��j�8�F�����w��e��
�,�6M���1�^ŧ��pZ�]n	qk���pQ��]c�/DJ�C���U��%xT�H�,y����_�X�߫��Z�����A�˫�օ!+�����6����G���@�4�Ӕa�μb"-��E��Y��1��c���$���uL�	^�j�w��-�%����_��at�h�b&�N,@UW�o��'���*Sa���'��5�Ш��]�x�l�f��ނY�V�:⚪�b�"m"-�EaL�&�� Yd5s�ꁗ^~�� ta��S��L����6c��{r���A,���&8����-nþ5��#/�k�m�=v�
4���k>���M)�'���	q��47�I>\����O�6��Z��'�D��oa��"����((S��}1A(�-V@��_x�V�����d�R��Ő�"T#v
��ږ�3��sV%���l��K$abғ�\���h?zeM����b`SҘ" �¸-�O�����Ҿj����K0"��H�[�#�H,Aq͒gӀ�1Y��bu1w�Hb��s�J!Z��K؝����3d�>�TLxSz���
*H���r��Z�6�D�T���:�x[�t�-��,i�C~�����h��[��t)��wb�"�7 �J��h��i��u�[I���/��!K�%#�*	�fN�i0�v@�0E��	w��˷I����d�J��t�����-<�_a_�aF�'}e��OtǠ�J�8Db�8~����T�	XIc�"����Y����I4f�y�����l��KJ��7H��*m���P0�5����ݳ�dڨ�y|]Ԯ,�K�Q߰����"���@�Z��J�X�8b�ᄱ�݋�]����7�W�w�z[�r������建�-�F���&Һ����%�7d(1ﲲW����TvY�˗'���gy�\Ϛ�h!izz�xrb:�F�b4)�ao�W\kkP�����SԖ��[�~'�-��V�I$|�OBI��L]�K���]�)�5N�<��Ɲ�<zt[�G͵j��D�=Yvb)�J*�����{j�Q�V�i�I���]����#��Quh�"�B�0�����#��1�!]��!�Oga�/��pT�&'���H�����>�x4) 1�3�1x(*�n�t��bG�/�'5��#Wg�fU0W��; ���z!?��r��Sz��}��Z�9���=1g�[�{nI�[�'vR�'�Ʋ|�kJ�bj��L%�k}ހ����~���(���ai����k��i�Z�,^w�Q�WTE.��8-��e9,��~s�� ���I�߈Fc4���R�^X�1'�h?�BqA�-�Kվ>ZjW�q@yVc<���&��
����<	戼rz k�k�.Ư�G�P�����.Bh���e�d�b#sD��;O����tN�\�?D`��	-���EG�?��md���|U8�߆��xm3���M9��������y��9S��q���d�������۪�����Ĝ̈́B�2֍�/W��|�77p��1�%����M!oz'ʑ"<����� 8�'D=�؂�����I�����~jD	�r8�3=���o/��O)��,LbY�;w)G��RV�fb5��H�ӭ�#X*��>�`�*�]#*מ]���`Zy�d�e@'�פ���AlJ|,��}�I�8Xג�A��7�!��Xv�Ҝ ����(�%^mѣf��(.oޞ�{�ƪR)�������ֺ�d��ZD����e�`�h~	^M��Y�I�4������m��q��s�qM�g,�@k��3�C�GD�}?���ܧ�0Q��ʽb��~1W��8W~���JM�.�\&'�$%r��)*��_k�4}ܫ{�-�����$�o���s����%��7�ݗܺ��S�G�U��,V��3{��ky:E�00.�T��#�6ԷH|غ_��f����⌑p�*z���-����7ފVl�|��RR���іO3�~�D��FF��![�2��Z�>S?���0.��R��`����I�X��_��CI�?�y4
��,Q�ނ]Z�9��廘ia�6�}�i)����keI�����E����c��L�"�(n	�S�)@�5���s4_|+��i�䪠�j�f[�����W�kN���<��h�����wΟ����Z���Tz�
!d ��Mr�m���!=��g�����SܮPP~ΎzEhCWZ���8�\�9����H؇4U-G�͍uHS���;��)iN�~ߧ4}##8�UH<���J���f�ݵ2����1q�S�-7���v�=]��M1�;!��e���a ;�EL����# L�^�F����3[��E.��3���P��Z��7��^��?\M/r�����.'���`g�M�̑�,�~C&�a�O������0��w���O=�p25��a���*#���~U�f�.&"� y�#o��Z��O�>���czQp�Ў0$`z�q�[��I�^�:��Q�箾�<5�kY���Vs����X
�%�c).QǢ���%��6x���KyvnP�ʰf9�8c�k��
"gk�uW�R"H�G@���e~ݷ�e�N������P��h^	XAݩ!�0�6pH,)E�WS�:����Y�B��឵r��e���*��������A�H��*8�}@*��ٰ&WP�Wz�>{\�T��B��,*d�^��	�<�q�����ߔ�PV� 2k�m��#��N�2�0-�#����XF�?�S �7��v ��^x+��aF�e�3�ٿ���?��@R��@� �Gb�`B����e��)�ý���ϕ�Rw*�O�s<�|�mL����[V�_�xuy8�'߹��b�d��n2��Ê��oV�y^n��*���N�M��V��]���H�rPq��G�vW��ǀ���W�G�j�~(!3�,T�{%��s����<�T�ӱq/s@ݕ��L�q.�m���zb7��b�p����i5R5����4\���.� 6������;b�{j-"�H_��!h�+0u�J���~��/��ݭ�3^������Rϒn��b����v�H�Մ�Q wB�b9w�K"j�/͓�5�#���~W��P�ndدve�r!;nd������	��lGcE����J�h��ӪF�� >���)�(��_ٵ$��ꔎ�q�x>D���i?0j����zubST0�QUǸ���H*��Uҍ=M�q��o@z�j�e���0���5���]���q�p��^����!�'������9z���/%P��✍2[mn#�����Cy��*u����(�ކ �I		�R(���q ^*�"�ӝ#���ʿ�����tvǷ����	V4�wEn�E.m8״���(�S������c�(���l�t���	˔���q��$��彛�5�&$����2����E���z9��/�oa�5)��!{�]l7��a��b �F"���`J)�����xz[�R�����Z/��r��P��hE�[�^e\�O�Ff�8���ݜk�O߲���K���r7��[�}k��;ɉG����
�lDҎ��L���`%���s���zo�A�p/+���M¡p�G�$%U$���40�AGX�6�P�'� N���jt�@�9�d�$����=r#��
�*��=��x��R�v��_���6�t:���'g��{�'�Z�����Y��C{j�	�qe��I+P#P0���C"��L[�)a�&�k5&�X4����y���i�edF"8�$�o���J�sd��J\u��ʓ��@s��,4 �yBOMQO�q�(��wt���[���*����o�����K�3���3�U�wфC���O���;j�<����
�s���	�m;��s��|�`��������?�Wߏ;��(�>
�c�{�1�������Mg�ܝe�k�v5�Ln]?B꾁� �S�s���
�,�*�%@:3E�0�<>l-MqnWv���>���Ӭ�#b#d�2<r�x�é��Ob�=�[���?˹ޤ��:aq����m�,W��,�yҲ�9����hP=9Q�<�=\�yc˗7ⶹԒa��2���
�Eg�xF�qv�-w������x���|k������R��\o�)���O
AH�D�� �:ܘ5S����J�:�P�G
D�m��)�F��u�ym:��^�Yia�b@�	c�0x�!cH�b4�NQ���gs�?�QD�0!A��_6�+�{a��˛m��U�2�xCm]~�
�h�6tp&�G9��ZyЊX���k�S1�@��u���_)��HoE6P�i9$�s����y�G�=�ᜐ˾�E������XF�j>z�V�_hy�QO�ECyw�>��{.��%[+��|���J�Q��$Q�"�޿��W�8�:�����tew\��������=7,dǉ&=!���S�
W���d~]�$����C�V���Ͱ�T�@2��Q��+W��bq)%�,�!�!$/��y<����O�<С��˻�Θj��59X7i�g8�zg�͍�r�A��g���pQ�/���D�{X�7�^T���X��p0Cq9��x�a���6�~��Z�$����$�v���W�7�C��bp�yK+�i�IU&��i�A��k�q>��<�B7��8!}�Wx$��P[��h���ў����*3�RmTO�9�-�m�I䌭���� W3�
1Y���O�s*A^)-'zߚ�{65UH�L�l�%~��_C�=��?
O��Y�;8��Vq܃T�J�v��v��%�d�:�Ġ]'�*�l�W�U�5�no��#�SWr���W,l�z��.�YV�"����Ye1�����R0G�WZ�:��(�~����YT��5�Gt#=����}2A�3���6��yu��M)�I��|J�մ�h���5lknP�hL�Fe��ȡYڹ|F��M��l�������Uߏ�4Bɮu`T��J5�O�diec0�#��o�{�ȇ�$�wJ ����1��
g�_-��g=���-VUP��c��j1<5�� �-����x�t�:7\m�N�HE��>��-1�N�(�����WI.?+.W�ݑ"E��#��V =F��(+v��qΕ}I侄ľ������!����t4	����z>KBoy��rL�澪������xX}r�l�3̕?���P��f�?}=��
�a�f<cm��Ӟ�?O�E�~��.�����ܭ\���k{vs�L}?�J�NS�_RX�uf��zW��7+�5�U�����[e�U �zI��d��<����'��_s��=�!S��P��x��sƀ@������4�k�%;d.������� �a;w���驝Ü�Yt�\��`���>���NW��S�Fr�"</z;v��J�n#��QX;��plTǒ�#K��0�s�mx��8���O����(jF�d�`��`=�[�	�d퓸<��6�0b:������A�Z���k7�N��f�z�F�Ilz�a"4�D&�e�b�=lZ�Tኰ�{��u���2�fJ ���z�z�(�����-l(!��U����
��V}i%rf>G�y x���}�k���)�Y>|��!��z�d�Z�]��
MCD�
Tr�G�<X�`Fl:|2�"t�E�<�M�.5h|?X( �J�0\����(��jB��cU�yƮ�4��t����,�ӰX�^�k"�
5�Y�7��-��+��7vE�T�u��,�ް4�c�i�'�҇��T�=L(��}�5e��]��oN�a�9�%�o�H,��j%��g6�{��4ae(��#�\�^Wf��ti�I�9��, �,�����0��\�$��pU��[zU�h&�G�v�Q���*�t6�����J�\+B�����0i�m	9����Po���Kϊ��Ñ�sB(.����d�zt����Խ���o�0F�݇	���-5w]��Vj�.���$���j������Z�����F�F�N/�����b4�K�ea%bDE��>����2 tl�f�X$�� ���J��@��%����. 4�MBЃ+ �ȑ��|d����o~Z�O��)�0~�. ��@��H��I8߷���leyT���ze��L��Q�� d@S��.-hHϩ�5����OL����Y��Q���ךd�3�O\px7���K�Y35����r@�	F_:@鰩δ�;l�h"��&�����I����	V�l��kq(j��3��|-4�x��i���d7@3��-��	7������4Ê~`x�w[�����[������EƷ��
��M�>�'b�*4���L����no�(�p�.5����[��
|
$n��Mpa��yV���.#z��[���Ă����p;P�N�3A*��`�5wf����2E� 3ݍW��n��S~��KZd���0�k��@�S�;H�����ԫ8a��������x�X���ZB^p��^����D�Y�]/2<�K�X5��Ix�G�� �S2%�n�8�'��𒐁�>Zx����T@���BJ�X��1��~WY��M=I������׸aa��ᵺ�U|����z�Jz�6�"�*����G�,��*�_����<c��. ]6Õ�KșN���b�".5�3w99*׀��T��OL�y����gݔ�"ޅ�ZΝ�ʞ�zsC��L�d�F'�l�����)�e�!�9L�-���;�]�Kk�Л�"��ޅK��y��z�Kr����Vt)��zRqL�Fn���~�g�Zi*��C�����&��fLJPj��ӟ�<�)�� �$@���N ]���{�x/e"����坤\�̓w��>�#iJ��6�|�IRdR8��$�l��Q�� gL�:��}�����p}s�d�<��D\PӔ�dڡ=jz��/d�xJ?h�R�ƅ��{��r�n�$9Y\ʉG{��c�E!���g.���4���;�D��4��mA��߷����yDT6j�I{G׋���9Eگ�P�I%�w��G�0�~���B��b)�)U6�u=�S�r� (��T��|��έ��E��d�K���{�]���W>�^�52IdXU��C����!��� ���� �TU��z�����?v�Eq�ν`��8n�����>���d�\aP2�&��}�K5�V�%��6P�-��������#��)r��L�O��G��6�D-p �K�B�Ub,�7���1C�ORۚ.Q�j�<�y���8��H��ص��ǎ�Wۅ���S�������=Fj�%`}#���.H��%୕3MMD_*~�5�%�X��%YM�ƪ:g��@��P��Z�{�1��Kz�I��E�!3jHt\iC�T����Asw�f�蛲��:yh�ʏ�G{����P]�n����+qi�U��&?i	D�1j$�c+1�����#MS��)C�2��V����VUb?*�Ō*�CU6mn���GJ��yg?��#�Tֽ�\�E`����n��@���R<�H�X.�K�=*>�nxo�+oF57a~$B�����[(
��5�}��/]�Yp�R�8RΨ�^0���喖�-�e%�]J�;ݚ��������JE�s����+�7��Ֆ�$Μ� 1.dC��L�iA��J��(1�:�nl�$�_�
���o�M�rz�9ޓ�=̬����f�дM2:6�ʪ,�^�q\��0��F�͊u�'9��J'����n6�k9�R�٤�`@>c�:\- h(��.i�)z�:$*�:�^��m�J|#&j�����vK�9X�Q����<��h���B,����n��98},����,q�!¢��AU��kCD�z���|$��fq��w�Fj�%l���Wc�}�r�y�|#�b�1Xr�؏�H��jbw�,|��`Ƌ�;}�a���]�g�իdJ�5l�� 11,P�;f���S\]�c��?)�{�7�Q����� �;,��f����n��,+��m{8��/+Y���c`������z��z�*ܭp�j�� Ƀ�C�f+�Έ�Da�������&P T��]�f;��`m&4P�0�}� �����d��A�K)�#�s!��?@�ӑ��e�h�_��
/�U�2��jz�2t�d�h��p���w�w�F|=|�:�n��W�`9�+"�R�0����P�׸f�A�R<� ���%�$T�ݑnV��^���|j��ش���?q�ev��-Z��e��.o�F�Q�=�=v�|zG��B�W�j�(�ۻV�"���t�~>���#^�����$��nG����(��C�!�Hm�O��ֈ}���݅�������>(7�u2�*0�7嬾���l���A�����=���QL�a��VC��<�>�(���:��E��6�8 P��!_�L�K`\b����UX��QBo|�wo\��}�1�I�-'���8��!�OA���C�66��Bm�i���U���5M^�b���&�f�[���$W��JRD��r��-K����z��e��~��6�ኁ��ؖ��OJ�yj\֔%��kDZ�ˋ����\����,�Ѽ��Np����v�J���H�U�b��k� U"��`����.��#�E �%p9~��8@xjD<G��!<YS�f��d��n��irw��^w�t�e���K�~�� �D��A�̘�U��\�Dd��:�n����LJ�d�@��\�n>ϰ��rͲB��D��(7� ř�h�i�z>X����+�F�P`����3�g!��f���+�ǩ�܅C�����c�4E��4fʽT��o|�=�ErXj��`ΏW�o����:Fe{0E��^�z;��Fa=��f�\���g%���m�\�Ƚ,�]\�Ah-� MX�|��;����^���s�\e�3Db��@��n��:<��r[�yV8��8ƌW~�DQ�,:<���V8�Ŋʽ���i ؉�λL\!�}�:�򵹗:��G<��������7��_��>&\�X�~o�����nL�&���0�=��}IdqH�����ᓳ�Ǘ�D��y����H�|)b�%s��sg�#�Y����u��~�� ^�C5Ƭp5�W
��AZ2�m��5�"ڱi��&�^^�
=�w��5���>��0���	|,����T�Y��Fn�����[ ��7:�����T�pT�|1�]<���y���nũ܄��E�1=�u,�L�{ҕO�j���ִZ1b'���8{�L�����{i�<�U4f��c8���y�2�SFX��Hl]���OG��f�<X&�7�{�P�"+�u�憹Í���%����%����)*�X������K����6��پ,�44�#B���~��aB0oT-\��Ğ�`/>,wzΏ��?"�$w)�[<KP!��z�,���*Tv� ��]����d����u���t��O&C8�����$r����|��i�����`h=���Wi�T��wl&b�&��Ri���l���!ҹ�Şr��=���tݬ��q��B����k#ؗ���Fz�)DC#����n��|�*jl#KF�����%� W��=�M��#ܹ �w|�0D!�}W^TvPyUz�A2�Q�/fՄ .��B|Z?��Cv$�[g������5�vK�� ��dנo~~�(dt����Y�wG����|���P(� StSQ��"]�+y���|���C n�]vo���"��Mit��l��轣2/C���nC�!�ɏ����������G���n�ԟ%^x$�;KIV�����.{d��߷��<��@����e�Iӄ_���B��jUD}e)䄔4g��~I�&�F�fr��!�{FP	Dp�p��}�j�>%%e��\�X(��Z�tg�-T5�E�~h+�ȉ���������}~�2}�t�7��݁5w�a����"fxQ��̱4�<b�`p6ۅ��:�O"�k����IP�{8X"Z�F �܇m�|).�����\�w�n�7Ibc��u*�Tc�/��&k�]F�K��,�p�4֯����`��j˱CӶه�[�	ם��B��ͤ_�ޢ������~�{l�:0��`ׇ�V����������%�7e3��{���IU����?�;�ʒOT�:�PW���N~��Oz�e�ή�D����۟�.��AZ��0�Xf���[�|]����Iva��d2\+b���|��Yn~ƹ�w���8�<}`A�y�N����G�	���qOM���5~�{%��  ���]"�<��Wq� �q%��?�P�F����ϕ��h�=�w=p��QQ��͋�"�3y'�&iM����z�[Y��˄�z�l{cL��$���>T^W�P���=`�! (�nvl�_g3��z�fMKL�<G��Y��i�Kw[D�e%T�*Y���(���;��w����>ť�-�.��^�O`>oqRCy-��� *�Wac�@ꖯ:S�o5#�a��B��h��N��j�`.X�ds���;��Kb���&�a�S�����:�d@�(u�n�48��6�F`dR�0	��0�W4�a�|y1)��7����ʸ���U� ��@а��p�ڨB�⊿Uy4@������p��ďCj�N�;�/� b�my����׾��t{9�Ԕ� E,�	l��Gp>�����.�s��o�e@7ty_�w;��h�Sl����H���&�oެ--/�m�q��2���t���消�o�IZ ���X6���"����yg��9C!(C��v�\��H $M���~�Z���NKq��KZ���}�� `Nm�W�b��Q&&޶���u8���9ld�ۼ��g�?u!�q�Q3��+��A?���-�+�3��1W���>ϝoX2EG`���L)~�7�>2h��1&sm�<Du���OM+���e��%���j���UjH�m�)�G��N�|���CF�O"L(ʼ#L��_�����p����g
�H��̀��)_U��a�#Ȝ�`���0⍦�m������"C�wI����7��+�W�<���Y����k\�׈�)�Ÿ��ٯ y�Q=�5Ҥ�%�����P;.bT���s|>B�}c��pg]�ϓ�z�:}�^��"֕SF*no�a}�(�����B���6g����ۚ#?2kz����7���
��� X�.h��;�v۽��:�j r(� ���g��&ID�m/3��7��t���$C�<�Ոg�"���H���΢�wN�.�Zc�Ė��8�Gu�ܺp�%�3��/t���q?�^��D�N�iJm�U���F�]�(8s⑔��<�wêۣ��c��hR��Q��7?����C���p�R���e�&2���./9�](�;C���12O��μ�4��N�r:^�����ȡJ�3���*,�5�gWM��P��"z��z8^�M~�wx`���]-�rR���f��$��G:��0�8\I{�Y�`�?��|�O���cL�o�ʾe�#��\��Z�
��S���u&g�O�"��,��Y�:�ov��#�f�i��w��2�����ڷ\׸ں 
� �g𢽰�/��-�;im���=d�Q�&��͊�Z���H�2׾"y73��{���Z�tu�j��di���������8�����^:�
��ڧ�@ـ�YM�yY��d5��Ɗ���B����:'� )Ju����/
�n�v��y�}`,D����~++��p�w�q�"2$��^:���&��Q�~<�4
�5�C��!:�)t�h�3L�=�ۃ�+��M�/�9�v�؏�����A%B������|�y�9~�$�?�m��k���
�����8دˑY-���$�'oE��`Dx�\FG��R9�6��\69M���w��쇳ؐPPk1��m�'�1f9��o�_ބ;�����ї`��>�Ȋ��8��i�H�*�ፁ�`�廉�TdX��󣓚�LS����Erzt\*UO��J�T��=�(��3S��Q�W������ܚu��!�9�/�Y]��o@K b���,���㟌��J3�!C����F����5��H�e�b&�{���'����j����l0��U�պ�q�˨������)/����>���.0������,�MSh$�m3��í��\�:�O���<�i����Z퍚��A@�R���R"q4M�W��`_-�\9�T���X�/��96���;Q��d�G)�&C��q]ݞ���9@�Y�`o�������?"z��5ܠ0G�Z���n��:w#��a�h�A]��6�����=��+��%-��=��$Ң��̪��j`]F�{d�di-�&C�(�G1�!N�(rVU;��U�
"/�kL����h��g������y��8���i�TAҞ�a��%dr�Q*𖾫A��eZkk "a.Ss�gj�43Ô{����fVX�9 �	��D���;��D��94O{p�,�����������}���b�u9~�l�<�}f�$�f#Ƶ~�ovo�,�Z�n5 ��m����^/�>+Zb���VS^#�h��.5�2B�N�(��nF/���*0�u�u�9�i�/a�˝p=
x�o�vNΖ�P�������� �E��dd|8{x���J`�'�Q����A@�u~IK��\����7J�n�?f�E?�^�ya�`�'�րS�3�cک(���yRa�w���-y�*��u!m����9l�2x��-l���v�&	��bٞF�ף)N�ٯoD�4p=��f�x�rmv���4":�]��c�nwL=�O'�
����t�f�4�~&Ш�̭e��,�3�1i�RS�*�K�m�Y��/�~����4����?��p������m���d�ЉM� 
2�b��ϧ�^Á��I�ޖJ���6U.�����В�+_�L*��у�Lr�(g$	�ﱵۘ��e��f}�o�Kj�����i��Y7b�s&������PP��&x��h�_�5��oF�<���~i�
	����V�)�>��0��	W�I��K����P���`D�2�"���#�~�b�(�m8u��S��������=�1a3z��S'�~�V�G&����v2�%	E��j�Ӟf|P�eIzi�nϸ��'�guy�
-{�J��c)�e�w\Šb���B)�%�j�O�%y��������9�(p2cn�ֻ�j(8*�!)�I ���x�\�at�<L��O�X@,-����vl!D$o�Z��Eu0[��z%�n�C�o��Dc4��w�#ɩ����TǊ4'�@+��k�3��^�h5�����j���7������ob�g/P�Ԫz����x�E�o�*b>¨l^�����],:9`B$JY���z�bL8'd @�L'a�rR�$����ڃ��|q�Mۍ�R�)����B��*��	�6u��×���~��V���e��VH�?(W"z�u�K2q�5�/E���o2�����S�i�S|��7��ꘚ���t�Xa���0+�F��v�'����׏i�y�Մn��˺��u-�j]�L��PQ�eκ��9�'=�UZ�n�Lv_Gb��;�"~�����l���J>�OS���d����:se����p2�mb�.	�� \kql�v�E��M����7�H4-�'���竉�1O(DzWMPJ�Db|�zt�y@l ����H�r�a��阫j�Y�J 
X�}�|�ǹ��H��������ҬQ=�g����lQz� fkړ�DP2_�BDk4j�`�υ�j�&�����>��a�a��N�+�?lK�6��2�����.���v�����M2�ao�Tu]��O%<��A�lK�B�ۈ[U�d�*��U3lQ�e8��זP��q3�+������z��O^@��O2��e75�+
���<m�P6�,�2�I[�Z�(Z�v$�7����_?�[��ۏ8�t��&j�J�Q��c��2��N2L8s�Ja!����8�˗TE�v3��� H����P�a,�g�RaH����ݓX.qz�f��J���%+F*y	c"iG5�������񚕞0�cg�N���L��$zbB5t�8�DH|ed�/l�4c�����8�NQ';f�9:n�nd�q�}�$To,�7<�Hn�L�%����v>�7"%_|�cg.�Lz���l����ڿ���k�����3'O�;-����.��.�aI�|���������2��H�Xf��m��-�]=ޯ�zi��(����]�\C�@�KuކE���Ⱦ������\9�O5vP�TvX��恉��bBߡ�"���E���$�#|�L���
�������ͷ�Q��X����l]PNo5��D�9a�0��9��6p��ؒ�ʡ�D,gX��bhsH��T�6�qĭ�y1o֫�� ���TspkΑ;j5��紴0d�/fyߏ�Q�W�Θ��1��0�{\�a���Y�JB�eਖ਼�1�!�#s�u[�miH�ٽHe�Vj�ʟ����	�!�j\=鱢�S���O�;�d��& vZ�g��V�s�R1�C�rI`�S�a��A���+�\p�>{�%�)���4�]�$�����OE��_S�lJPA�M-��\�"�_�ǈ�]��0�}��ٮ eiu
����q��U~x�U_g�Cw�@-U���4(���epSd�m?D���x��$��n�/�"���Z~-)�����0��?�L��k&ЎC���wZ! Z�*���ر�X��b+��ݘC�w�����2�c8��7��wX��4��w��I��j%p���~Q���tP �C0��i�-��� ���Ʃ�^K�ƛ�6�Ԕb-��ز40�%.�F���S�b�q$�.��P��7}G�M\���Y�f@��0��;�,�w����^�	���`ap��_�<Nx���B�|�Jp7�;��JeQt#F�~��])aL��i��+��6��3��@/ϙZ�1�
��φ�\.�fZ�Xd�П�2�g
,��M`�n�,�\�#�WT��B�%�O`V�<�Og7����o��dZ's��(,Nk�����C���עe6~7�L����Ӈ�!T��Z���X���K���M5.к�H�ir����jSݻV������w��#dSrQ|cq�z��*H�t�R�ǂ��Yj�n�����7��ʪkv�L�x�b��YL��I��8�����[	��ρq;1��7/7���Ʊ��C�o�i]�!N��*(hL�>
dv�}ȓ�=`;g��`	{�a�@�79x'@8�*�M�t4��Z��l#�S��m-XH^3>�����M3�d��dܬ���|B�8ma��5ͳu�/���,���Ee�60�����ic�S�xbIS7�fV1��r����U&����)�`�CW�]6���y]��9=�X0^ϲ���S>���)Jm��Ĳc���0�G\��4���߂�<��HHhP��f��K�Ŗt��:1�V6Ii*	2�-��a����&s���:�oZ��x�d�ePRo�a���1�.3Olbj/c��W�&/�:r,;���/*fN1tB��GP��c������Sh��5��m���[ɚ���7�����@���Wn��*�§y�A{��7��|0�R'��<QO}<��v<��[j��eC�y�Z_u�D�aw5٠R��?.���2�)^�a34Gۅ�G"o�
{�ȥ�|o�kP���eLQ�,�L�ެ�Lv��޲$�Jؿ�8 G��%F�xhާ�����.I,g4o��-����~�lN� ��	a]B��W�eZ+հUAP�H���Q3�k���@>���e����S.ݲ���^��ޅ���#�4	��-*_��S�މ+�)	wu��P���*w����9^)`"A�1�f����F�W\�s�E�Ɣ�д)֓�U��-hRꮵ{,K�7{����'^��H��`��nkIE��q$bK]R� ��LB�g�t�/�&2|���γJ�?i%�a��}��h�s��[��T��Jk̜�f�	�n$%��ضz���X�I�j��i1���d�4��z�?���6�5̊cG�S�
�
���m��Z�p^���҈g�;� z��d[�XZee��w0�B��2��k�6��Y� 9�w�U���Qm=��JVv �D���Lc~�B��y3;�>�vJW�T�ʄx�lZP��>���9�~��f����Br��:���3��)(��Ү\����K�SH��fbF�s8P��\���I��r�T���q�����J�Q��1��cS�\��� t+巕�W$< u��X�hl�����j�!���Q���Q|lۙ�'ǫL�ZW��-�iz"�I�{��+B��Kah���{ls�z@&.Uj�N���1�Ԏ*�|epG�Γ��󟨑 o9�Nv�g=�T�u��-��k#�͕wk5��&������򤻞A�!��VF��K�C.<_��p[��e��[�FTq"	)Ϛ��=H\�,ɘ��<f����x�,ק�τ�*�'�蝶,��+ߌhz�*��B���t�crZ� �5��'���{ǀƸB}���e�	�ٝa���%�R2��U��h�:ΖL�zz��mIQ��9ϵ馴}��A�Wh�~�9�K�����5 �H���S��j��ϭ�!���G_�/[���hdv�� ^�P�L)��NJ�r	�Çqܛ<�ބ��+�>�z�h�8�	^�C�.�U��H�9a�2���%,@�
� ��.'�M����>�࿲�N�wI8�g�eM�q*˱E�"��	�c��*{
�j��,�`����8��oG�l��U�0��U�,�N-{��$�/����Zpo�^9���
l�W�}|U�C�s��CT45H%>A�9J�9D~�yi�������o�e�+%�!DxmlPmAz��l�`-���:]��]-����"/�7$<\�`�{⫱�9U�?�a8�B�L�� ��VOҀ�m�S{���T�fc�&�1������|̂D�]ev�&�����7AQ#���l啶v���W�ܿ]R�
���W:f��2�ڭ�n�!�P�c���jy_�y�Z�
��q~l��\ǆ6�$�p�}`���2x��1�>`0�l���P�X�f�R�@�>�Xl��Ɛ����U䙁�浵/������vL����$OIv��ܗԱ�����215�.u
�����Y�Z� ��V�@����~��֮�'�K�*+�[�
���n���&5-'�K�P�F��dOy~n����Ēً^�_�щL#dQB$�(�|�����{^}0���S�p�]L��W(�
q�����<�8�m���$��=N�$,K��#+N_'�F��a�O�]�A�=zz��m�X�ax��z�J(|�P<��ق,�})��s9�q�aԣxS���� �G�i�2:�H.F�p񑏘�P�2)6���qc'TZ�Y!�W�A?_��Mo�!�̷5�st��+m6�7X��ϵ�IQ,���`)�V�]L�S6�Im'&9^��τ�w#p%�;b���:��{-�K.��#��G[����s��Ԇ����y_�|S�̦�ů󙽷����39s��]�ʰ?R<��a�q��Z��#l��%�Ͼ�-�k7�ߌ(�*�%�{St����	
 +��:����n����\U�)ʅe�b&�~R��&8�c���[8�=��L�1��5�~0����-�D��6�^!��JG��{c�J�+��a�_6�jJ��:D����i@Y��n��J[��Zdxj[�􄪐������&����;�Z"�[s�o!� �.J$q���0��",Ľ��1O�ɩ�h~�YgBq;Ɓ禡5���|:�a B�`f�aR��4|E뿷 SѸ��|�o`��i�P�y?���[Y����=3� s�z;&�C�Rtָ�����uze�Vs��H�;�=���ϭ��� SL5��0�zvrk�L�^y=�<>ӽ�ySx�B�X�A^���F��I#����;U�0�g�61|R��KJ�����v�Q�5T�J9�L�(�pҼ8-^XX}@G5���r��V}Jިd���Ƥ�����t-����j�ߖ,�2[�v�e'���Roy�x�0��8���ZۉR5���&� '���~��%�}tj�۫��9�����@���PQŸ��5��[n���l�n���4Q�-k�+�v����&×ʦ�.m��Ň�+�Y�=G�J��{��y^�g�htԮ��8G@��cöeՄ@��6���R�,�� ����2�y��\P/#�]!UKO����2�r�~�D������.�+�!Q�_`����TŧE��	��,�B���|2�y:����F5�F�[<3�k,�˰�������[�a;y�{ʾ{T�g-g��K0d�_
�qS���������C͉�!��8昇��l�QT+�H��4�O��L:L�Va��@�Hx���z ����d{H�
��_Sw=p�����͋YWd	���3�d�-��&���W�u��#��n�QB��_+����pd�3�H�	���?輔̿2�_^ y�S=��z[><�x��4G	�YؖG��S�m�se�ὦRLe��!�y�Y�'_-Vt�"k�z��Zt�B	x�b�	�?�U-�s���b��Ձ�3�>N����g�xVc�A��z4g5�Z��no06�_���9����b�_pV<:�HO��@�赓|B�g��D��5�J�8aДE=P�Qg8���zu���"k���\찄���ţ*�*��W�����PU;�YN� �fS}�y!o� �g[M��M���iC<�	$J�����m�j�$����^8�ð��;<��_P�iq��m����y)�LK��f��F&٫���c��\WCQ�S�WL�t��b�9�(�*�.`��&&̠߭qFar1t��z��ק-�@va���~S0�Ih�L����o���k�JI+O�ï���
�pz�lR"ES�>��j�Wg��`��'/SF�x�i�q4�8�QTKO��r��bƚ����qnJ��W,`_*�)W�t&%����*��3���4��rd�Y*��
7������)����Zj���D����4v`ӊt�Y�V��U×�D�|MV�s�����q�|	�BN'_e���+�R7��<ƮU�qa�Mp���X�5�Kq�EK�6�y@�A��ҁs8i��o��_��A����7��R��O����%�ƎÇ�y"Q���} F%e��}?�Ƶ� 0�ĉ�Ș��z���Ta��.�p��F9�X�rq0"�~�^��%�HV����s��<oA���u���v����Y4�tsq��$���������E��j��֊��KZ�>/�;� ���`��}����ko�h�q@��F���%ۮ?�1�����>)�ʊ��ZW@Ł��kL��U8��瞙�I!���V��e���9s�N���/�5dڜ���p�"���-���m��@�-�í��b>���۰���	Bu�빝H:}�$�c��'OO�2AQg�a0�2-�t���$��6�Q̞B��/ bG�q$�53�\��*��)'o)r��D�����"jO�/&!�Q힀��1M�ߖ/K-��"h�6!�qq�g��H��\F��
�x�L�|i�{�$WKJu9ֶ� d`'S�юmdn� ��*]��a�n�+u�GH����;t]���"�9�{Y�����'4���]iЃ*� �	�}��f�㋃�䒨������^�M �쳿��Ör���8����Xyn��r��6�G��
�lF�l��嶄��+����T�֝߲����>��PpK�ݽ�Y/���<ה-�����jM�/;�3�8���{�dE1�}��(��Ae�%���?Z.�![&��3U�w���S�Hu��:hY��\�R�ew �럻�d�krEʨ%��,h4�:��1����O9eF���ˀP��������5�/`܏sS���y(GA�=z�5j�Sn(d���+'�6�'z���~���ƌ��9
���L^��<�N��*�a�ݖ&��,[�|�[���Oj9��bU�!;Ry�'i��F���~�x��YɃk�-�A^^o�[�ϔ(�:l?�#�Msw(����q��aQ����&>a�޻-z��]\��?�s���L��uO�\N�i��@&C?v'��9j�X[��@&UuRz՛���]�@�KT�Ĉdn���9^ć�}�P�]�������G����mM�34�
,�D�Ql�9|-ud�^��C�|;�ݧgaQ_x���1���sA��!�1�?i�&2!Z��9�8;F� 0e9m�0�i��FI ���Յ�q3�!~�2�!\���"�F�����s��7:#� g�b�pп��]��T!"��o��I�0�@>�l�B�������&\�ݬ-�G�#�%�h�b�r�t�x̬� �7yZw{������^w(���n��mu�����*�n�j��g�ϋFsp<�����ԉ[>Å�Dq�!��i�9Iw��،��:��5������*� Ю�̵���	�V̤��낺JiC�/�8}�L޿��ug�7̼X��K$*�ХqC����ꡋ��!̐��<�1�w�h�i<2ʍE�9�^��h�B�GQGa.� ����򟋦��Ӥ+4��OJ�\}s��'U��9+��C�6��l�:&�2-��]��xeg$�R�#ɑ[�E�3��A�ew�Z�욲&hTf��#��>ܪx�6@�양�3�0Y�,���V0,�_�*���=�������c�N4>M,Vό�WH�[vo�]����'t�p	ZUo�,����A}�����.a]7R��?w�BG����7�z�$����e#�Z�gp���x��sV��F:|`iy!P3�j����-{�B���9�]����q�R�1�8�E+\�$&XZM+i���ڳf1(���cvı{F��]�wo�;�mƎw,�)��a@Jk�	�@�� �a�W������o���t�	�b�/[�E�Omp�.Z*����x�T�",�%���h܇���Q�
Y�8�I0�+-"��\�LP��S�VĦ��f��������Cr[������>ڟ{U=��h}�D�RQW�)��
K��n��k.]}�A|!.��ɨS�=4x�����6ݬL{S���n�n��S)n�s�ߜ\@n"�S4	��uTG/J�^M�~F�#s]��Cd+����E����3��Z��8,�g��=�s���Q�$��o��F��R�<�g[:�^;׀J�n�٠z��fY���#�Ĭ	�^��WH�L�pYH�bͩȯ}/��Z �8c`�ԗ���w�t9���(��0�n�����x�"@�o�*=�!�!�*eUy�vH���=s
�|�B
t�jp}ȇ���+�[M�hA?'c�c 1ԉ�o���u�%��jD����k�]����?�q�¤h(����,k�ғ�B�4��i���Ql � ���s�~�F�(����F�k����)�U^�〗����Z`R��D��RË>jõ� ��Mn��+�m��Rq�a�s��5��Kp�������trk�Pbg3��$'������|���	?VC�}jρB½L������9�ti*yi�s�k35���� ��v+f��ԩ��V/�{DK�])��j�������G�p$��(a7zK�n~��BYԘ�~�u�k�^�aYR�g8PT(�\�˸�dEg=c#�t�&��66[%!U)�����sNr�᪾�ځA�X�V�5�Y����:��Q�	h��I����cT�B���&0g�����~ͣZ�3 z����õGIxС��}t��7�y����+�K����BH�{45/t �:��)��mBۿ_��2Bd᝵2�"��uut�|,F-�x\T��^�~�?��ZWK�io��I���C3H��~<(ul5���+,��w8iF���;Lf5�����u���oE���R�:�F� �i�􆠩'��#d�}����i̎��^Ś��+10�z&�bp��4Ze�N=uS���~�?���M��TJY<��r��1��AΙ�A��B�M��!������fU�<��v{jwJw,�X�Mu��fbt�ǿx�*�@hX��sK�2y����?|��H���1�'�%q�R��SA��M1�
}f���x��S��ڷ�xŚ��"8�y��	��uX-��s���D٬lI%���%LB�Xr������@/�$L��Ծ�Э�eB3v�I4�ۂ��W��GE�D�'�xo;���,zҜ%���\�*Q��R�T�ud8�z����s�x��wmRTO@��QP�E�*�Q�����A�7��o�-w NE��=�.:���ѻ��~�׎�E�+�d&+��LV���kTWr�l���sc�^vH3�%�Z��������i�qg�#���h�9Ӄ�J�jq{E ����?��F	~�Y�3�AA�L��=��0e�<��Ƹ��D,���3�����%T ��u�x�w��J���ɡ?��8��\
�������|6 �@z�m��Z��Tm�M5 ��R�e$ �d�Yfid���H5Q��*;���ga�DWg��Ď��V��a�c�B�����8ׄlg�'КY������'����Z�H�ޫ�`���ւn��ڟ��ʀ�Y-���3�J@w-և�M��!�v��v�N<0Q7�徏���DHAZj�p��V�s�_̥}��$��_����	K�1b�ö�w��\��5��?xf�Q�s`W�� z.����(�r"�'���IrqG
�w~� �{0�����a�z���XW�e����aKspb]��F,$t�� ��\�77}��D��$|����U��p`<n��=~�F�~ԫX2WN�y���Veck�Sd��Α~�<K��<o݅C|�s�����w�q�;�C�),��o��M�5yt�i�T}�}U_[��aѺ�=��U42Bi��2i7�tuP��?(D2�,�j�Tr����Ă��~w�CM�)J�~S֍4�����	52t��ԀT��7ʚ�b�~W��d��.����Tib�)�iH�.��585o|E�WG�������s��W��]8U�"<J�4�T����<֞�j���cY$�Z�0>��1$:�w�����E_S�Oί����A��J������	ڄ��I�[gW��K�/���,t���E��I�:�V�q߅�N���?�2�F��?��F���ekw)��7��Z��WΧ��#�F�鄅��I�Co�"8{�ViM��%��
�(��,�S�1Qe ���&M5n�!)�'x�C���R��e�/oǨ���`+�1dH���b\�ii��w��׭<I�؛�ΉV��f��k��������+���z{�E���@�fл�z��j����R'��qr��a�B�qߑ9��u�����4E ���Jc筒_��bf�*�&}����X�����I�j_A�<
	S�H��+s��~�fۄ�Y�P\S��L�V!�?��~�s԰G�PV��$�6������ Ud%�;�҂�Cg&�gzq.D�+ꈃ��C���%$g��6�I,�\�x�dA��Ol0��umG)�������� 	�I�W�rÆw�-פ+�}�QJr��6���v{AF��L�;%
��v����%������"K�Y���F}I0��X�pOcn��\�ɗO��a�c�/塨qG�:9���I��vH��C�|k�V4�Ld���a0�k�m�Zmw�4�|EZyDC��6S[�A6i^;Hg�~��˥� L�(I��dڦJ�3
�ܬ�hr[~9����^��� kר�ɶKL:jo���e�C��R��4����@`�)}�)���Y�P�i���ZR�6�paؾlQ�e�E�q=ENx�d��F}����~�
>O��� �Rb�U�$l3�5�Yd�]j����*(*�'˹������aDɼ�{���g`��=r]�I3��7�(J*�����v�#��By��_�pZ�z+�tݮ�ZTC��g��ۉE�Q]`=�$v�=l_x���y/όY(N�e����g�b�GL��K�(��bL�]1i[��>�s�E�tw"�~�'"3�I	g^4e5df����_?OL��$�{qd�w��JI&I������.�U3ܬ�j�n�\�pa�S��|(~Y}�Zُ�[��2������6�ċ�S�Bf���qH:�N��v)��r/��'va���=�[8��s?���ZO�CW�O%��<PD�ؼ�����y(1{�㸤����Կj��P�xNo�ƾ���,�,���CL`dvZEj6�J#�c�:瀕#��'��Y
�$v��te_���Xu�ER��q~��\Px	W}Y�i��P�M�2qE�Rs���a=;w-�8I�#��f���ޜ�� o-�6�k�2��F3�����/�Fvz�o�xk�A�x'�՚"=�[g�dE2&���6A]�������<^=,W���L��g��V3��&~M D0<j�yt�6����2�w��> ����B�t��|}&���.UY�}ms49��Ԑ��.��N8o��"��^���z&O϶�c̊t��o퍊��^��y���a%tz+�\x.(��r@�bg���eW1�\�>|?�FN��|��	�O�ZO!B*~d�C92p�s����O�R�"�Ӎ�(2��0���۩�S�2?zw.�m��#��������P�3caħ
ܲ��oom�.[�����;�~6fv�`�ծ���gx%�!]N� ���pY��D�n*1�f7խ�x�o��	�8{P:�~�v�ICmXFe��hm����0?�mC�&�YV#=t�v�y��FUN��)��|p� �aE�����`���e�Ǝ�����ŶWw��<��l�-��{`�eҦ	����^;���牔���p~Q\Żh�:���Ϡ� i�aaEu-�(џ>7�p�}�/��^���H*\c�Q�%t=�NG�+���=�/�D��@S� (t�����t����k0}|�p���p�;��� �d-��/� h�&��f
�2��s԰���� ��_
��VN?�0����ު|V�~X@=
��q1�X�>X�� ��r����b�Y�-w;�q�K��d�1�.�W���!w�w@'������`p����#�ǔ�$���0������x��}m)���~���P�c�'F��ad�`� nǋ'�MZ�`���X٨�eǆ\(�	�:iQ�Q
=˭�Y��c��0w#��U��	��;'�bAW�T����#�n�s�&)�.#��~~�q/q�.%���6�sj��f�&���Y�~h���?���Ɛ*	w��Y�i�%����_�|��3��dkh��V��p�Bٕt�ޙL����}�_EѠ�H��|d��ź������'6sgc5��ywj�^�|)�E�;q��p�J�IZA�n�%�E���h�^�-�mb<���2�1��DB�'֩r.	���cj�x/���k��I��fT���T�*��l}���ɭW}�j�U���+�@�Y��J��~4��0�o�s�
]jf�þև��l�Gǟ�K7j�;��q��:��c�˫���S'�� J��,��A��kE��,eVɵPW1��{��K�b����0Ǜ�d�T�	?�n<^��'t�[�R/W�P�)�F����0p��ڝk~H�`���ۣ����J�F�)��}K����peH�zUȶ��C�-�1��I݂'��	ko{ͫ���ύ�DSі|�����w�ѐ%|���f��l�0��x�w�wJ�%c��F`�X�%	��1���Á3��ߺ�Ͱ[C.��t�����0�ȶ`E8�2���oݖ�쨝�Uϭj.~�}̐��jv�A��
���t�ZD��i�����Ӱidg��
/Á�YB����nE4���O�j�^��˃V���p�ڭ(yc���U��������V���Yi���Чk1×�h!����)�1�)�e��)��~R\�
Z>�����b�kG, �X������f|NU_���8�1���'W����W� 	*�q�����t���I8`�FO�8�lٱ���ss��C+C�z����,�}�m �*4Zq7u*Y����D<��� G��s�|��g-�CH��(��������x�����Ub�3���x�%��x��K���WU'�9Pؕ���_�� �mP�&)T�|��u����|J�^�E�	��]۬�s^ʮa���=������ظ�<{��e��[K7�q�b�b�����^L�mznB�4�	Q���_�F�G⊚�f7ԝ.�,`������:�Ԝ���"В#���q-�~1�����gQ���V#E5m���%�=oL�6|��C�e��r�l�g++�}��H�x��l�P��LM����4�IF��e�v2amYစvQv�N��[O�&%E�fw���b��yߣ��A�yB���`_��[�d|�n	1�F�9^�b��̂_�Y��!�#N7P��J^伅"�`E���ao7$Ю�x��u���D�v!"]��VIG|CY&1&�Vyʛ���#�=�W�#�N�G:{��#:MH��&�d�'_@���9��w��W＜RR"���#o��.^vB�7*�vÎ��)�)���V�����>�~�et��)	`�3�ٖ��j�g�,|�gM<��$|�o=�g77;� %x���o�Y��s��]��@�-iw'����^�������{J�XO4���I�u�����ʤ,�k 2���4��>"'����<����/-vll�J�5~f0���ףӃ6K�Z�*F祝=�Y~B=�ǵ��-��7���/F=���;��-֯r�� �[�{��O@�d�T��$��%Z���r1�!^��;(�j@�L
Z��MP؇)t��Su�ݕA�T�WF�T���V0��������S������uf�U������}��n�=�ٽ���Cq�5��C���\VG;4LO��ʐ�$�-!{D͐����$��ֆ���eI�>���8�(w�E��?[��gx�Wo?�Х�GŔ��iʰ3u�F�