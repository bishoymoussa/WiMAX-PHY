-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
ukYYc3CbGo7b9pxJQJNIWDnHa+br8pEZ0/h7wsVI9zWPVm8FtBqlR5yRzLJXX/2xBUVe8Yy0Vg5P
EHHJqTOVss4vIbFCYqCKlrHiLpG/FDTIoe3T4vExSzWkH/AOFRQ0uXRzPkI0us2oKJ0Gn1BFgScJ
dUiaPkLWeG8YTbwCgkDj8pObQ7YvHoWfbk3eQbgJBh5pjNP4+Nkx3p/YipgRyfFiNQYVwY+qrqvd
k9XGd2HcmafyZp554wWeXe9g+xwpi+6GQzGxV+o8sHe/DcjasrH8XMgWiYK9voGuVCbXMCM1aW1p
LK4CWN2R9o1VIt94PNOXcmqjNJQQMdg6Ack5tA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 9920)
`protect data_block
Iu2xx5n2DOsyIum1wND73D6JDTQjXHVVE+vBDaYYFm4o1nOenmchTDVcqzPKKTuxHT8bdV2mnQpd
jfWRLyIZfwscmzw3ra67GoIpgf9dWbTvHdpgSuSetSJ2QscZBmyLPQb4lv/vAlEWDynwypRJsYNh
EHDaSajhXHpcDVlSlavrhUt1iGCJ0J9L0QyGf1k7tYAK8ggT7LDM5z1Ob68/pww/fXcx5HfljcB9
92oes0eCfV2IUNrNT+rkSIxPEsnD2/1yfB5H7DmoXbpsD9twhIUi2TyIvqzJVSram4958zYccgTi
rox/ZJeTxdSDZjsnHmamPtZqJF+Ea85kuV485aXaPuJb9QCyruR8V2R2LArIOpZbp4s/+U/zUvHq
aB6/lI6SAdBlC2kxtVFzyRzjYw9Bi5v3icEBJny9UF0+fGRjmVoaAFIboz0Wn/MEsQcVOd+uxfE7
Epe+E1xfTDsLDGFV1KXENbSrfKJe1Vz1VU7eDhDmaFbCqZiiXwuD7LLQEMTa1Cb7GFVfFiYgyQ7u
ayYib9nHPUBfusGgiOhMuyk+HhZ/9O6JHVMgmXvggNhoE9R9QDwerl562X1o6OlC0uveXAayZnN9
5U/y/rzMoalcFYele1yHremi8HdXtXw8Mvzx6hH2LzR3Dm2HiOLyUw02eMAC3McW24+GB2avLoYc
/R1w7Ck1ktzHLVEw8Q7FZnPdAyUREcG0Ykn46CMjTyqKy9v58o/XpBSS4c3D8cJv1LD9JiiL24Ng
SDF/JdYah1BAOgcQsFtUs9Yzl4k5jCfmBtmAqXJCn6W9+XF8RhLhWRPG2mP6NcRmUHd/3l+ubvvQ
ZL7gD6dD7PCo3DtyeKi03Oq6D27gaz4vQ4gXDtVie49E8TT7lp05OtHcIic6Shhnv5KghKuy7/+A
Px7XBasSf0XKIjMF2IMs0RaADBmTUJu0hCQvb7V4oscqO/WgiiQh8oBothgXqfkkfaQtaS/w+pMz
+JZMvvCE82rw204uwj96fnVeRaLeK99WRd/dX4ae9zwXsrVmd94SnxkHJZxR6fn5B5q8nftGVQxF
8bnclOFgTNMu1yYeZZGgYWEZfsAf9kA+oMxZNFJNCBN5/BnnVCX7J9tCK9s/uabsNzbJMch7TqdI
RVo/7JOKMZh5XTmldQ9iG5yBGFnHRl2rRFkqBB+idU8W4XQXQc6XqIB0eWNWL88DG72sY2SsXqMA
O5VzhufdHvJI1yDs0GDzKE8xGG937EqtIa75kDFYZU781/YifBeiBmA0WQ8lHqspvfOLBkfCXQ7+
LDpzz9Q1ACR3uoqoHIznnSRqBfsWpMAigyl9TvhweLbRMtlnhZrf0l0HsSh1pG2mVhSXkmrywt1Z
QKQJssAq/vvpYKXgzP8ovxpQuARllT0Fj2j9HAwyXfe7Lu4+CSfBD2u6u80/xm/2rCs/i5gyRDPq
97pZQNgBxQu/LqzhDmpE8tF+5qTiIWgMhD6YIR9xmbBzOtsLUraNhpzIanv5Zeo3CeG2XmtCT+jl
FjIYKYPH3IWoHPIDr+N2l047ktuBtzVUuYNd0EQVyp4XKXnsYtejUHImYTpcXyvRGhZSTC9KV9U4
9BEjMrL5aGhuEyzT0pV0vjDv4V7H6A3VKsM14FYZh1UKt6gJD2lFienut7rqLg8HZLamYuTBhCOG
WiBy2xZnQhx+UdmBffHon7qeyonMwuMZ4/E8EdAanGyT09pVi/TzFyAtHPDULgw+DA/mfIZMNbm+
xL5z+y4nN4FUKn+tgokU5wr1mEqyXpQzcRLibaaMJ3MeHzlflrUGc4k50EsAusY1snAeLdlTg+Ll
QYoAafjgHKhQW+XeKisZ/pra6ExCZ3WNo2ifwwph827bxESTV896VnlPP55+hwKVWXYXyw5BmiQu
QcRXfS+PPrbRSFQ3Obbmvl1qg+QKzMyDzWpOG9xinXnV/lLxnc2pLpvsq2IqB108x4lS/AMZiNtw
UefzSB4AI+ve6pzlP9tlIaxBJG+/uuZ2L0IHUGIhei4+uPh8GKOSBcMxsQPZMePmkOr+CtSGZ82+
J6/V2Iv35CvcKhaSmgqsj0YBCnGJ69dpWuYMI0K8Ar8OHXlC8b2kFq7dvLWhBXvs4wT3wSYIOhCi
4tnAed8ftkDZqjv9E72UzgXCotiiGh1ioWSlgliYjzaRqY5RVxp9Bux+gbUoJOeklHfIPe6ztlcH
zFpoVCIZfiiebB6H1yYcqBnoIxHrVgXcCNwRBqjin3lIl1nhSF8wuNofuxrWALwArClKJ8gVYkmP
IiKrTxGLcs3/qbEJnB+8seU432qhKlzBWiwOZxTQ6H2DlnGzEREn04Jd3PewJpTdP1cryMwz0oPl
MtL+dfqQdt3WcSsaF9gzjZVPD0THYzWkayTHOIt2YiAhItSHdJgTchpIgk0y4mNKVXfWmFw+i7rX
IqkqaOYM2s41/gQAHUV+wEYHu7NupdEmm/0myf/y9LcSai8an+Gf+zN2HX21D0tuIL69G0tcKM5m
K/bzT92H6wCwnRnrPthhj1Lem1DXJTubZRjTg2BRkLIqDRSBKTrL1K+eegI4+sZsaAW1iUNnyzKP
nTqp9kPPfmz3Z6wAw69uFsW7MlSN+H9fdexcvUK5daPW4Zo8mb6UCl1PnXFjoZkR4jqkzyrdaxw7
JevdF9wXbaXqbc0fZ9qT+ZGfDkBQATa3ij/8j7pqYVcev6B6SkAsJxdiPieg7DFlHSYwcyovDuzy
LkRdEdS1lOzDO+7HJmWEE/95OlW0FL/q+nPr47OrsIN0L+SkVUKqldtgNk8YHgs3xB1zeaQRcZwe
9hRpL2A2ntsXgYs/Q/Sge3+H4woclBi+BdTFI07AkEm/ipjgIdAH60AK2GjpXMgywfH8lcDPSDpj
oQE1pq3sykwFFe7+ZA2uZUdlBrn+xOyUAMYVGo8+SGhlK8Yx23YnSkweIcnh1ImZt43QessyMf99
jSFnQRbLhC2lHk/L0WT+Ql2o+rXUnvmMjCrcikxmrnYNcM0ZVd+ZlryenBrFlHOXxEv14rdWwo+c
b3c7vXdOomsmVuOo0mvUHGCwPmwa7IeOqDQlSX6PKUh4HyeEeEqvC1KxXmWHyPALfXNi0UlM2oiG
4dzJnWXwFgTd1CVDPsvLkdzZcDo+zXwelusNH2Ps6BbRV94tta9Ms6RqSTP2H9SnCqaUxuCJxbWZ
UC3lON5gNXaf6Xen6cSDReKHEZFq0YZBuJ0Y2r/lkxHkrMcTyZKWjWsMipSceucmeJ5uEg/OzWt9
kf9ShwKUghBDmBKhgF4uCwdLpp9ObgYa5u2Zj+pWq7GxJ7jN/o0UHx/FJO/eOSWN3H6wnfHbF2/H
WrTmZkBd/OEcspDezQ4j5/6CxUCdGMG589fOCi+MoKEKgB3r+LMjFLDcT0Suou3SEF5fB7gM3Caj
XXN0lQ5gCfRDIL4uZRs0X3slF6ZsWiVpEpSfA6lrj7iYAdcKxocIzUC+S8wvnBoC6w7m1oyGtBtc
zNVhDBLF3xWNk8FtVcp5zpuH28+qQUf/ZbcepifZG4+adB1x2wPgJQ2kdsQb4YjWWrc9QK3SpSgY
D3TPqwRKPWHkYli4DK5jB0NwBmYyE0yjtsscE17EJBBcAwzG2gDzLEBr5G9j4jdO+pxrXFkKZc5m
kzo8bB4InTYncL0Fos99zXBQwuCUOxY/7Y1ZISHe8Q07Qbitgk0h+ax63yDSFJOSV4OIGk2eF1jR
k/ZePOlA1VCtWWNATwNOKD0/uBqTIEV+nstuIQ7GNz7bfDr25jLXHFixa2+JWXmqrnXNnW3mzMCh
LkT0m+bXfJSqNjkX+oIGFBk3A99/sHLWQO6KX3auXuJpF5+zwurz9q+TWZP51jjJweruqBQWS5qP
Bil/5PK0xOi1roThLnlup+pCnnAGF2P1UDylsq9MIv022G4jj4jTHqZLUnjmNY4rJVpHQKCFTVlo
2eafr3RPE2fg8rbkyVyCsjui/LxGcqxdKv0GeVo3fltqlJ3EO6kjUYOlXH2r7CWQOA3RLYfpfq1M
SM6k2kyt78zbSEhlcjRQqKT1ckfjP9z+NYikHH5N8EK4vADhw5B/zCFUc4Xsz+MbrBT2MonhwQ96
i8Tp9aBxnp5LaDe3Uj4+bOCfBpSqSlacabnG2leE5zf5P7Asa8l40zKfZ8d93BKpw9Y1WmTOWDE3
pZuUHHHmRXbUyftfDSklabvsGgjHNAJLlNpB4GevX/t4RYeGn/a+ZwCFSDVafe5WyImYiwMRoqvf
q4HSEOTu04otOWnX0pWYnBAwTGPkov1Ge2/XydC44zTpQBVxj1O3cJX2VzsdXdNE/2K1kHo8bgUt
qLN6SU01mLq4gU2HMxHrkqbLuzGrOi/cRTphL9hE7OMYzZ4sspvJ0J4JQiSPBcPpOLZCFrm9Hpp3
caKnzALFR3KPjfuoGx0c4fAicWLug8XLsH1DsV48+1o9IMqlRMc+7asgXVrSIvqUSpXl6pcsA/2R
TtcRc40lzW6olE2fzFuO/dxrqdPS1fKGFlL0TCdXHyoKDvlP1ZsjiD4TMCKovpOuopl3tWdduFeR
ub7Qleg/Yk/QVgUtahLJViRHkDdeWwJB3XNzT9Vy9qZOQ2rZBfg7Uf96Xrgc2tkXTJbsWWRrrsxy
uwGpR2/5Y5v59ism2YLZWpbtS7D/DE8P7Mjbpcvs0jQsUIvIVGTVFYdZB+RSYGwlWBYEXK+jprRy
tbY0saPHOM04Ub1sOultVG8WEjCHWEvNC0156V50ix2sKpqBzedIy2yQ+oVt1WFmP81XDoBpEWiX
n641yyNkZJ+S+fC4AQcuy2HVbag7wj+Y+UjkfHow6TkChNKzV7kk+Xt0W8e0hLv2UW7eRVPjGNVn
+eGzXA61Kdh8wFdFm8Z+2Zc7vEkdb56ChFTZF3jwFJtcU0cSYdqlixMCPM+3G2O5/8llK+8ocE3b
RwBkFG8B2SBGLHMcWMNIFUluttzPlWXgn/bjGu22e4/Gc00snjKYfyuw3+BWPpvG0KwzoTU9uqcL
kZjD7E2lpK4AVw3L8LqfBuP64DnqeDjrhz9IgGW3cOfKJlkzM9qupK2/jqhq0XwvMSh7naMATLpM
9V7NEMg9Tsl4rQP6/h7cYvshVp89ojbRupDVfvMmkx4QlE112OhUpDw9vTBSXjybdiVHTUjx348y
1DzSmNucqpbOx8bbWS4dP/Eeu+AFO3EOuU5v/D1EwLNNizGtMhsmgnn/gga8KZHk8SdKCzTngDEY
TYkjWdlP7olMyS7aWvXufPGtJdgfXb2nMTpIcQ6EsP43PgFdDj90DxoCkPOrqmNWwrbditiQoOpX
n+IsWXR6i+7aL+rgknLyNuBeqBkfIY/tLFPZHQEOdlR52uRWR0RtbASHcVENOTLd3BPKHvgsM1EV
gxa9epzLGe5bE6El50cZR85kCvSWaZi40FzsYfqrUMNVRx5VCUvk8gmFM760yrvGWhu0851xQf0e
h8cKWHKRTLliFUqRtQNu1O2HRNqIlClItMc3OOVxyAg7z154PFUaHX2P2uJaGHL8zzgdOm7/8neY
Ke1KFhJroDROwq1m2U5ty10eYFjdIAkqKjUCkxfjxEZrBwSussyrgV/6+Gs85ZffaNIqhgp5XMzj
li0HdFMApLHfw8bYJ6zxddZBOR2+dEww5QZYQUA8zKjmviYE+gyQYgAAfInIER8e6n5cKrXhE/ax
+QfGwORhNiK8eaPJidTz/N/b0ePXtOvH4Yrzryww6eZ5BmqReUm0aYFnp9wIDjlP+11Qy2GOanGZ
9fAq9K5N88PcbqpfWuHGHUh116q4Fjo4QGSIHwQ541Vm1Sv63mHyM9aXxhMXMlKSJCR1ITwyfYcz
ntHpkyUsQfCOPKSAR0ekfdqC+SGYee6dN+jXpknPIZYtadQ5eRiOJzBAUXVLe4Pcd7ktS0hwk6ag
Y+kmWiezgRRYqpz6ShWnmxwsZiOf8+8LrzT2ySJxG5zCftnrhsxHoTzgdbrBErgAzzcJCW1sO+WO
9zrgwq2MGyMVUcZFkiNEsT7HapD3ms73rRNzPwihuMO6MWFD6NWfyy8u+CgXNAfM2EBjlkbODlep
+ReeDO91YKXykSCc6xuyL7tCELMyYnYZD7JHqgnBHvtZnx+UjDxluJFxcwopzWwtvlJV4lKPtgsC
1960vqks1WFgVpS2ZsM0JYELN9ACr//JDn1hwh2GEl8j6KOCEUS3FxwhXvIsnb9Dudzz5XQvSzTB
er6D3kUnZmlRHWH9w1NepAthfNlK04cdhQF76Q1hUIYNsI+dVYYAqrImjFxzxKajuef+weQGiHgO
h+IUuPmrh0C8wOHBJ9uOn4mi+KW+bO/Ri5qEOrt8UbHrurfuc5sfYbWA96vJvvnsRQzvAH4Ii/uh
gY/zAEwBQaYsI6wWnwIO3FWQZAGr6SuvfOo75iDqGadeDAvWxbVKPpCM5hPBJKAPDWCZxWTw4TGG
QM63b7urlEXs5RWcm5scClJlK44aA88QCBCfwxj+R2cbL0hjHVjEDO7qx6RMqWPWpsnA9Rni3Ozo
qq9WUBtAUu+kYjMqSbm7zZsozQksdxL2rVcWV4nNaA7mqzA/JksMfiYkLCf0iN0CtIFotS/nBQeg
Suj+tDS3Y648o+aJVaELBCMsQQM6Z8z/ziMhVaHidTjhJEn5cDXo8CusIl5mmpQjHvWzk1XkQXY+
8Kd92lQDQB+awF2mZd03FqhsygRSFLa3uPvmBJJx4em7lj7l1gHYEWzfZmSN3tpw+oDtF5MiIWok
agP0YNV23RK83ClenAhFgD8B55jP3XHFajGC+ChhZ456j03YYeir0uQU1jNd6qllhLuucahAh4tO
EXqo7QU4WXJNyLTWSI9oVb4YwM11SxmCxyHzdYhdXS3Wjz5vA5WTa7c7/GGixIvp/0QkTnuQqjjP
Q6vnRwY1czRsSF808H480LV5J8yjSTSkoKkF1sfo7sgRmXXfolN7IUsk53TwNHqV1fdO9Xom2+nV
RgAtThwsD3jSlEe9+8m43H1XMvM1GgBmPHNdLTzQgo3BanvC4ddlzdS4enD51jiPliaF4isJD+zJ
o8HxMxv/J7eVq0BIVG8D33bTYVSgHCCrFYrcj3OlELN8k8hqcIdi+3cLDYSPdX9bD+wqQzdnpOqH
n0+lBGqwaKXhiXRD+4wex8237fKGpY1pu8//CHtE3nyPN7Fxq78QO+7RZutBsIp0E3akBbkgrUti
OeF7C72TlrW9EMbQIBqkZsip1bTG0fPr/QxB+e1pNqkVSEhhjN+HNeRWlxWiaZCKMJt+hT1aYiO7
Yz/KfqtVc3kUV6PKx+MyjuKJLkGBaZ5Ac0GKdL1kYP5aokUuFpiTeZuAUb2I/O4BvIhgEhPi51Fc
m/eJUth7XiEsuGz6c8Zow+x5U2gWSYcGvkkJ6B3X1utzLw+fmakVR5fwOurB64fpGjDjenuplLnV
OXlGeMdy8KEmM+sv09kVNUyMpJD2RfUibZmzl2SO3/oayAcS4KoW7d8G2AIm3UOokgMy6mvyRv9q
7g3c1hP2Zbp70yldp1v4G4/V9VjwTrTZ6PpT9h58jbQjdCGOBl6H5eC68+xCc1OZGhEl974n85/l
/Hy6Wsu4gvVKKlVpPhTznmZAiJbIkg9qZwcCVvumJi8GiwbIOj/NzOGLc9UVl7JPD2oeY5z+LU3T
wgF3QZ3mS2mZkxFl69GUW8B1f4t5u05oZLqWat3MdZ5fNWnnuB8J76FmOHP65MSvDnw9512+PRJH
BjIIkmifFKkDXQs3wo/7S7I2RCKcxJyhI09U4NlDtOmPYDZUz1ed6NNSvgXeIhCQrmP012/e5dkS
UjiweVO5rUZEcMsQiaIZVj+UaVCE5VFnVhjUTE2CrMiVyXFYiOjdlrBJGgyu+LG55pc/ZECA1YZJ
VwVolth5gPch6XbyZKbxuC0v5keVmnhLuVFeyoGFuHhyeAuiVcJ9OZV0A6SRgU7kFPOFHk7hMtVJ
anNKlYy2imZEjyp95BH3Vgzf+rkPu23v1LM5VMs3Q+aJWr4bE6NQUQuxFzL5r8mhyON6WAhQeIHp
uGt/Nmf0CwSavlBOZK2UZMtPu3vgHhvL6dAXVmUm1H0ER1H79ha0V3eQMCoG5bZgUB+D2TR2dTRW
L4nB+suoVVFYhM7umVeAZwOk1YJJYA6bJyCe+cc5UWXSElvsTkz+KLO/ka0uzxDWYzK9033LtV9L
bov0CE7VYFTCpO3W14mScHZ/1PIIFYa21YvkVRjqKo56Qxv9StKNfdWbUWED4b05QZ990lpzqbzJ
OKcM2w8c9MXTUBKon2BOgqn/UiXvlqE5xiLi4+ePII8CGxTlNOYNbdRcxNjWq2IWxdjwdaTu++r4
dhJMauXLKoWGMPB/KwqEWgX0CkYwj1UnK2gyE18mgM6Bs3AJewRO6Y+xta5IZPHoTGWQE/NgYOUG
mIP+SVIVxej61BvC3+IqKJNvfmutG2Au8CppR/40sLee2roH3kMuKgqj+0TvuUeWyfJCOU1qOMNh
MWZpOxsyywYP7OfIhUsnp8d9o/Qp1CzOYLGzFFZdyX3bsZde2VRWf9f2EnBHvmOUdj47pgq2lIWO
Xq5wJ/xRMptuDyOq+QrlmMxIK8c06m5jCCf2KQysjlc2YltF3TDZYGTTPYy+lksAgzb2rKWnQR07
5Awb919ilJM4OWHvb1ibHuC0FHb8rFqlBj1sSDNUqUzAuDOYhiOi8sFFbJOI1+cadpEPxHkUBoPA
nScrGBLBJb1JPOOZWQqlkU+zlqvwUsjKCTFIvWgYzHeDtCxWOF8dj+FHbch92u3wk/8g998Ncb8E
Ca4aDI/9ql+CQ6dcnz0Uu7yP5yYbAswAWEmNCyfKm6/uxmnPSGmRp1TaeThNUWCV6iFKjn+2xPFG
LpD8C/6JOneMsQ/86eSYqAq4ux7U1M3h9lfbCoa4wWmx1BIh+VGl3Pcvzx3E9BdBH7RSjP1mU2fn
Ggwx/eHHPowmg4QSpR2dmGuYv0IvOt+VlxMDNCkWwsQhgvK5alqqRVmWTYhVceDC+iaaeoekLERx
XTEq5HyukSyOPRCsReI8gKE+0ROZi1xrafw4fVyR7KF/006YvLB9SZezhKmjOXsdwdCo+mmlk0Am
JN+6FXvREyiQBNE+jY8TE6YXrrSk2No6xNRBTmu5+gmahEMAsBClMYfYmG3AAHZ372y5u4RD0AQ+
CZLoTddHz3jULaym3c9nFdrWn7t7w/oUh75xkFvRuLIdb5Us/fXYlcyGhBgn2Foj94Y00QKaKPks
GFfC9fo1gQIdl+uSQkoFpZmXZHyIUZo4xtH67IEbLE51Nl/4AU7ucn0JzAgI7ELjlXLkYek896O7
KyOl6i/KXfSwgIE6rfg8yCwPsawULi5pprVF6sNPYJbrMCvbitFpR8yNCQrD4+i2sj7VDjZl3Qtr
cvMLK579hlpDL8qxLlLi3CYjqu1byJ6GgpYKaowJPz08J8BQIVGtUmPo6kx56TPHUYBADNeCi6JW
GFi2tMYEZpXwBqVhrEw1d7PWUazkmxDkNk3I9q3im7Eodj7/0dV1FKOSPCj1YS++Qe0iwkSJwXBw
KjldM1nfC8IbZ7u+H16UvWhrMYyw4soMwjAqqi8ru/9pqpUEzi7RCfG5pKgsCfeGmvn0fcECSEz1
m6OX0J6QN7XhNCbARYQz8L6CDfbvD/2q/zBz8cvhjm1fDQ7RsY5HryRwV9NL2KW8twyl+oN0U/B8
7nSYuNc7FcRg4j5jkvMZ/cW0majJA3KE7Mb543sxF3LcAk96f9GtpDtlmNy/uppkLawKBzdoVCMk
ISvRG0hUQIk10fQ9JpW4bIlDWQql5bFJwLqy2gXppJOgpIWaMNq+320e24W0s0FywCCcrm8g9H0g
vZoohPAKkq9Yr7Jg6fQqcL0aTV6FgNZagkhkhjAD5965R05v/DYwlqOaYj0WdJ+QSAJwfIeHsU5a
/zX8/4xbt2J+zdyuJxEDNQ3YAJGcE9vvxuas1Hj+o5d777XcSd9mAdPFvd6Rp8S2wfWzxTrv7HXU
KK3dnaKGwvruMdyeT7PGI+zqraspnhddwz4/pwjWg/wfJqfsuSgGUilBJOFlWVMok1Qjf8T5qi70
QwboDOmHdvaFC8wMnASfH5qmyufNok4CsQGYRhS9SNVUfL1NqBsHNxWMGmMpSAZQNsoBPz2Z+YDw
MJBIpTFky/RIeMVwSjxW3oAQJVtzCTLkejEXfobdiwqPgxlbci1DZEK9Ya2lt/5B6hGWTf40gKzT
6v+Vu/2L1NO5I8dmFzDgBwEdVwgsgBLnEcCmg8k/sK+tYHwTG3GyR1ZcGCf8VT0GDJC6cIjTQsKt
QShmzg8Dsja9Mnt32SlmiCPD5H4O93+tn+TR4ELHfVFgoxPa7ayFoi8BK0eiPYjD+R54DrFgU9EW
gRv1UKzyYPCPqOKga3KsFmtb5ZQyNyxyvGSeY0xsKCq6J03oLKB9RVzdUf7YO+Jr5Q3g80C4FD1t
7uVLUOsywriNwZh50JPyK9ZWk0sXBXfV/UOvbHNps2Fx1JrUdMs/CKeJDMU2/7NmwKomYOUn37Yf
w2IQKOPSHJJJT4/4njEvkjJFWTCcWSfWfZQFF1UxUKQrQzSFOsK1iAmBsu28or2w9V+sTOyWk8E/
Hd4Ck3S0WB3b7NKRjNuZwVsNmYN4z7hOdqn5aMdXWfXxYFnRAbfkqsQp6nHlz0YELocT5K8SsV8u
v2U6g2lOuCnMMIPg6sbnL81FrcfSjfaTIaXWS8v4uCczxtwqD965SUrjMF/B7tJcge6Vo4oHU4n1
gesR1TGnlmT93bA/YpobR+OYwQ4O/tm+ycNwXbPQXf3ukhkkvi9k013UgQQ88dkoxvLd7PJSP4DL
1XKTd25jJyizwxQmCwI0kVPlvREk1QGwjqKXm11VOyduMC1t1SId/kLVumWMtMIZSbP7TDDRGhaZ
bxeAZVU0m+h++3QZiHmR5nJzfnKvKhTMzpAG9+u9UWunWz1N+2GB3IPbJ9tm6TCyjoV8yclg4KDL
8hHIkc3xgpg2e550iEW1j/rARk50URo36mamAZwQx81MDZ4ekjM3pRbvnF6jNYOmUqeVqvde8CCY
rdRcdm14ERAP6aCX5e4qBi/vjpdjZ62jwGIUKd0x1X17vNcSn3sPp7TgmJwnYt4kvOxi5jEyKF6K
UyxqXe7CpBLKsZDh6bsL/vUqnbU3GvQkIiLMN+AIhdIrQDIBD6I6UIUgyd+cACjarM0x02Tq2fv8
bvtiW3mfk4pPwvz7o5pe53Zne/fBRnWDPoPT58Wv5hD3xybc5jMzgPC2ZLJLrR3GOnzPgy9qFMnI
qdBhkzU7oWJJG4VLGuSaDXJVUCQKtsSPdMJJAIYp6lbzZrTs7jA++Yh4lAbZjCJKNtPMGlM4leKN
tAwBusYg1SKfpSi5FZxPxmH0YQcM1ur6Bw6O55AQBuQwPj6F0B7M441GBrZkiI7UDUPLwvciIVjC
SQ6RM+vA7OXgojEAMCkNcni5EFyvL1iAY9AUyycAkCCJsn411z3hBPetcQFgmL9jFOMEJiQkhHl2
+nWc+wu6ZYL0yFmdOsPt22V1/6UszGjHFCz6fSJLbtKpKoeXKSpdepWhKYv/nwXAOEci4RGltTGG
Kc6Nh49y6Aidm8gYDXXPlC7ADuMTMNgKO6HrmU5qji66x52FRrSvYbY2ceVH82mOhUh3wZGbTJ2m
rAhBWyyOfwgMRBDQQ5cYdvOXwcIuY7MSwZMgVbfbEAcHMgl4dDkt3WdJ8ZQ8qC5YT19yc54BCvfu
UXOGOhqXuSKJNirPoBfoy2OGKj5qVh9hA1wAX5nHNphA0une/YBKG/D12kOaPLx2OvygcXyimgPd
/ghIBcOinaRFteTv0OhL2E7F7W1wSrVG2w+PXjSuX8rCBH1Z1WJioScmxr81y/DpEWKcx/5gMe+v
+PyyTFkzefI5K8Mpppqn3x+AqG3ZZT4pbcC+9W+EeqJPpyb0Im5lZKw48SjrvFf44NCyuQlZHLq1
Uhy7YXpczdi/Y+E/BPWCw4r/ndB/LgbKz7nC/cqV4NuMF4HoOnd0aoyQefSU7UUTGxMwl2U0Gs6g
I6Fwp8MPMVjxuiiGVenZYCPcQGBbGMPaDgc9fkPkVjFMhajaAHWKlQ7/9X/Fhe1Ssm/ptKQItYQe
f9IqMTLs43M3rBjArZKi+hLcSQKhyE3d6gEhNrnGp5XkyEg8NYdp3mE7MSU7GodRpTZUgGdkrF+N
BBALDhYyy18PwKrFcHzeSzW3ihUAersq9nTSW5ol5r8ky3gyLJLQOTydWX5qgt3GWgC5YIUN6vfG
Ojav52KkftxKFU8ghaxy04YGMoUpYO2xdFTSfV1lQZ4GpKIGI5iccaeQ0Si9EK3kvlchRMWjgujg
qaOQxRmYtKfdXkKyWr7XMOUasqOHgS6n6V1R/afNoXzFEHeCqBeCc7LdXcFl+eqNOhIXVi0gYzdR
Vm6WjfK5ule3rrsw9PfsEHc8V3Y1jyZz0E2jtT4Q0zxOEQc24I7cT/8JzXg9IEHuLOEyFHi+N13c
mrt4vuYtR5idpSz6Zp5R2xi6bcup2J5NDQ4SCwsaMRvr2Vs9QkowqqDNeC71QRo4EUquPIKnB/qU
TNd/obKPVO4uIgHrPecIhrhFFzoItSjJjoPqwd3QL6D04C3MBDx81ibohmymZz1zUuKv+AqREGAv
F8YA8Qo1/lPSnLgYkgTW3oljNA/hZqoXfGMYGMM3hN6LeUPNSpSz9d828GxPptf0r5+7inH7aPhr
Ni3kA/T3AhDrTkxh6AS/BhLADmGp4lXyEmavbpEJAIKQ6WXQBfsDFVdSvrXijal8N4IKvrgNwFN9
WHvcP/5ZuXKAUVea8q3cdv9eGemmYbvcGa5uTHJoYAsxob2ZZqPOrFMfPLHGFc7N5l93S++UdwhB
G06ui89CopZ2Y3mL6nWh4nbSjwGbUKS+o28z3zXwA/ESzEgW8Ny6GXHB24gNcXFA4QS8lHqhogNn
e8LFTerxY7ZEXAxwLqqMfeqX42ClLTAm59U3qy70fwPjRlrQN/YE4WmSk3jWZVBWy/+cPlTCIwcw
dt77ONi9dzvG8T0RdIO2YlNoMNrFzu6xxiRrbgFhiowehBUTGA8VeBtTy3MLQahhKJtFq4+2Awou
ccKbSiDrOozI6mf5G/s7ybi8U2M1DwuLlF9GuAQxzMC1F922MsLM/eWgQB2mYNCxF8YQIiNMRbYC
1tU=
`protect end_protected
