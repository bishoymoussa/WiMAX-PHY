-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
k+AZV+529oGOl1fviZ7IE67iWDmjUQ/AqSWiB8Tadu2j0bOGUbT2/zshH6LfnFq0cxCib+28dWUz
z+YK/Mk9KGtUAHkAnjyE5Zc0AD2REXZfLz+nMSDEaWLexdykqJf8SlpwJHH3EbnapHMcNHhLdrlt
6dN2Dcz9yq6cofe2ww9FSWeVWFOfOdGBlwVobfPiXyWImrCDDl2nCTUo8eqcEMS2x7oz0NdQEoac
18Y2WBcfz0kWEV+cqCCIBADrbSIvzu4Uqtf1fDDLJhsjbUyQyN2sL+NzqRzp7M0bKs2r9cyZRUTV
nY8GVrNImI9W6fnSDy7eX0zhy0fydO2Md3nuig==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 102384)
`protect data_block
0Fxhon+dkJPAa2dc2xytNyg6RxNkzp2SwBnNvbzyc3waQWx0dp7vPpCc6FGHE5gZ2lydrh6a3F4t
7LzXRkYxl93u+gKJx/ZYSLeGIXI53anWBNGIEfB00OHmIUVjU8PioX96KYptROFQCddKteJofPCB
rmN/dwSdT26bvHVDacwULkMjELjbNDG8vEQUEouPqXOiz4kfWY9kqd67y1koM+pCjMN95CEvwO9i
f7CgSA5yNrvI5UFol9Z5rGO/fPMGu7t1UJV9eZG5IXbtM1pLcSbWSH9NCSu4Mobb6sDK4+Cb66NA
fZuS2ZDJ2vt9xFfTDxQqtS+rPbGiDGKOYFMhryp/2CYTzn/0GCW9wmzrLxEavmE47+gPdEdbHUOF
f4O3Mp0UUyE7XW+dM98mCK6CCAgTXoKBPIZ4cgW4j1aa+fWDy+Je4mZMrjOYIgcTmQydZK2B1szT
Hxe8il391/bx9iP94/E/NqALHrnssAbGDAzIX/agomxyzb29caVPhC0fVBM/a4jPDkV1NDMI7ADT
2Lp+kTJvt+9uikkDveEBz7ZaiBc261lCfGAuPrLNw8/XxuQRmf2Irm03N9kM7H+le8gTACR7/qir
8A8t9VBjMyIQmUNyZzhKw4zUWV7/bI/V6gZvr5/aNT1P35WsD4Mog9++/C1WA+OH2ec1Zr5+t+Av
co8jBsJLZFWhFttmNnA1Wi1tKnLzXMRPe2Jtb4KKTAYykwGzN5u6FuazMM6d5vkgke/Vxjm/elps
twteN5VwAhz7PKMWygvqGaOS0ncEaWvH5pWXQEEkrEMkExSQ9/cj6zOIW1MqeLlybpRBi0+Ocb2h
ulqdBe1dPZ+YwCsLV+JHPg5NmxvUkmBos5MvzX1pep8pRtVtLua2JLhTPL0NnEm68rQiSL7rFTCh
PYKziJRbW1vuww1atYgHVzYf8V8pgPJZE8T9Kcq3pi5JvEfKj5nQtwH2QD6ht02MEbgfgM2yr8MA
Ev/Qeqn1Xhe5481odxfe31ORZ9ViFn+Sl9DrlZwOjAHSm4vUozIW/ZolWAjR4JCiYrRWtBNNg7u/
cM7+ALtZl6R3rQ6MkI/GtCScBiO3yWA6Xhl+qHbGt8T6KUz/E40HsiPpC0XjnC8vkJW3Rx+E1Frn
XDn3rWCWV+x3VCA7C8kD4t30kcR19/R9H0ld+64wsq7eQD1umwkwO0dzN6cUrq3jEWn22Yf4cx7q
529B83yQOI2YlExlfck62KwPzA9WLrQgLq3inq/oDYpnrPg59WfYL9yHRayFGtnG0XnJT2XuZiF7
Gs7hhtaztIFM6Ix6D+4Wguk4T0OrdlEVG4gMwfPdv5ytdtlXrmp1iPtJDDXCCEVxrOWsWWhiO9PQ
KWpUK8Ez5RH6xQJq9/JhABsGoT19jRGt82eMnjRsUMi65f7/YyPhl8vs4QyMvzpF7jHcVg26hKOe
MClHddm9mPaAuq1RvmCaoG0eG5W7ErLTrsfQwbvDB7r/LBStspfIzGmb8CiNSFgsFzmQ83zFNMQw
cilBOxtq441ZcFjKTESfNb1fSGx2JbY6U5cWo/00njQZlEXXa0ZdDzB7XfgTg37vOz1cLbd0VipZ
IdnLbG+Io0/+QCz8UlZGKACcuQmyJWA3zJh5NDWcGqz1mfH3xtD364lTwFshGKkEoAcXN5Cjr2Tl
aimGUSbgonLrYN3i7pdb6yCZrDAC4WIzKYQAcsAFCXz/UZ+yQRTIvQg1cc9wPZPi8dcEHKWNMUYF
ptUaYE0J9+mvG9/Nx0K8ciT7NJ6IQ9l4vxt3hVJ9nIn7IszccN625Wjii7SL5iGmnBh+0CfGBi1a
s2reDp7YSTMNy+DbEfiKO/LdqraJCIXGF17aZYnZOIno3pZ1WmcOLn+9mcWpL373Dk3zV+t/n+5j
jM1yYklLhFLD7nn1Yf2mejyN0tKS9FOI8TaoFhQzZj8HhdnRRC+zrbGn5/jfRYdnD3eJTqtYuUfv
GMWo57eNwkvZ51cHW171E4usEEoIBS2JT99+7ttzV3iPD+u5bkdAa0RI2y+GvUtZ8lpiRBTmVyog
FhCbbCQgc73PeqwE8N7elDSp06Fv9hLLLxHO7fDcDKeQiPUaIkbv6WLiMGMBtaQBGfk95QQOTysn
QTTviRRrxzHlqY4O/Y9XLs47lwKboXkYc6IjsUo2cHafHiwjTDho8wuz9v2RHCBGE29NjR64NHb9
ExpuNjJSX2cN9kfCFTFUS4K1u874EX1jWvnTzGuZPOX5wa6e1tWxaABekptwCcAk7ZP3wLZLd3Au
qNfhNmDSO2fZgA/qiHY3YAguevDRFgrEAmQs0xKl5rdUBR6RAdNkhlptZd/cR3za8AXEdljoPBtS
su+8cVANIGyU+2B3ywkL6D2bPBRLEKPiAi3/pDB4RaqLYh7etOkBAWYQaK8jKfa07a3RSA3JzvZ2
5cmeqKkksXJd6niPCnN4WQ4YexdYkxFa0nYgbMaqqaLKaJGKDlizEhBtlZNv3HbAhLX+b/jB/Rx5
Bmx9jB9iu96QW1t7potS+HsjZlE9b/MAFmV2nrCYTXr1Ujq6hrlcMS/Z0+hyI+olH9FtgiesVod9
iFzjo1oLJOgwOkSSNyWmJyWGmo5MaqiAW7yJFOLQzEeTeaX/eCDUCsw7xXLe0Zo4yzQ+U+2cM+Rz
+xoVx4ckIe7mffMBJbQNWm9LlD5beNOmC5j2Gk5qc937k5OTnsoxd2Vv0Wq/spZeDq3JO/moQk2X
ZenKal7quKfqVa3FDx3M6b9mtiNKuXRV47NAmrz0lPuyJWSujur6EFQuWgZCE0AXMLEM2AuX2L42
wZW/rWdupZQo4RudGjWby4YHgqX5qRMn1CUSOGqZpQQzW+nVVpSlFnfkI4jQkf1tVFJH4zx1W03a
Tr1tOG2kCMYXLj8j7OoebDj8PCAQ//PsXTIqUFoCgAT8w9Ixc7vh6HmH9xQA4FvU6y2JGEiaWYZI
anXePkAcu1dzhffrgFTH0f3TKK7pagu8F1rtnJcyN1zSt7C5ifrFvvoiXbtVjzhBs5LoRkEGTie4
AdiXXIGjCmSsMQUciuyR9UEuCj78lYGmYdjmi+ZMEG1cRhwuXXQuwMAbClyBE5IiRMazdVhpJc5p
YnWTmQubqdft9T9HfRHxLo2aU8tGs8JxLA6snfWsPWd6lG2Sbl/vEqVi8T16rhic77i1FC77FoA5
eMAGvKF0IA43DjytO77/3vRfST42J9+GYCaeNNkmDcOXG3nJFjAeYcfUlExA1y1Vgzo1zRap6wLf
gCxwF3WIZQxuvBskcCYDc+a1p8ulbl2M15IP4ivBjd1DxWWzI73ADT4W3VKvTFR4qbMZpmC+pls+
Gq1vWzaU/YywI+HEtl4BkpjXC3TKM5gdK5TPtcK00vZGCkaxaSuEkHCotd8xi03m11QlBuRUU5gj
DoPLrY4lC0aagjF3l/JVaMxLTBcc6ACZi74wjR7YPycpxcxc+vig6tQBfAr6mibgSZoClQL03qpS
m0aVSu8w0/OmuLezOD0rjtKBIj+z5mIx9Zd9tbGvL4crdBUAl3TD1VU3hTa1jRJHg8NEX56KYEDk
DBxZDjhnJjgDcyIcgH+vDRNnsk8/gIwq4nBKT+X6z65claVmhSeneQ16DuxE1N9K1Frh1lRjP44F
7o3dk7ZjRWDxVsfH9REURdwMxzqI4LcIjC+3d9N63449SuMwRq/WGfCbEoluwcTeS2OnT+YaZt6C
PhR+jgK8nmGAHTteU1c2GeB/QGvS0d+2KfIg5zT1nH8sE1SV48BlGPdc+1e6DJ3kYH5vawnnYFRW
A4bSH/yskNUKIi4ygwUM9kbkF8ahQgQPf3+NSeG4wj+8JM7Hi2JHjow/Ql7fWGDxrXxJPe/NC4yC
FURxeoO7yQwrYkCVkCxhRZeY8QThZaVR8sLOsHS7Znvtd38goSNuxOHzPh0Lb2YIL6HBgU7eFN8H
AvaFqoFbj9xixdh9Zfm8Wm3L2sJQxKJSEHj3yYfhy4WgrmtOU25uGYU5/KoiZfxvRhU0rr5ofsCR
Qz5/I95Thf3fojphImqkB+ee3W30Yorfz204aELV7jrD8bjpjy3qTdctZo3Slvpg9QR9jUGkGUyF
//iLAK45ihFryeDQbbcjT8tPaO9DWNtV4uEaNfkuNlrC/jauWNC0OJlQHtRnHu/6XrFMpcCodbxl
3ORK+SYXO2OunMgVyNCvPNhByJnY9icucn9UVu/kjkw5KqRmbmrugzAny+U0P+jxBpa0z6r8v8BB
Woxch4iorV7Yo0CsWUqyS91frLH8eBYd3jDoB9Itad8+qW+WfX92CFfIlRaMOFnJ04620wiZhB/n
einaC7lnzyOyZXi090DT2gLlJ5BdBEU2xXj68gaL0qHc6i5JXZNjfFNwNUfTFw+BQYvPdNvOCfz/
hRsRfL8cmOue5ARPu647BtO98qbw7j2KcQPoBXcTBBwkzeTrMFZ77gWKjn7o6w/J+qfSPUcYIHKA
KgDw/vkbfRt9CMAb0QoHfTXAD4iQnt1mpmwll0VlEMT5YkCO7/UDXulbZgj5WMHPp2S8x8drY+i3
TmjkDu1uF2CMZ+O+KhHue4BbjuTBSm/890CCgQrzbrhGLDxwHbzmQ1kAAhEJhlJTTL4TxgDguV0S
pkDlnTVvo5SIyHOgoNXu2TJuUTN9Nr/I7gegRcqMGKjQnBHhsk4CPwIMWoRBJpdWXRyuFQfv5xZP
Ghls5J77/mi4/O+WfYe+re3aBdiDCWWQVw6bQVdPcKRIAQ+X/aLTLkoMCeO80rhrgnAHWS1iMjg1
vZCRlJ8MOACeHMYx2bc55XRV2ekvrrhxfD2MWycSNMi16JfNEbZrTgdnRXQ/ZHAixQMWJTgI48Li
mYMhw1Qu6YAc8af3Ua07D3b4cXdXmkW4R42QMJtAtp+xw9DCim1Vzj/ds3rRX/unqv1jyHOo7DDv
ijo8TWVKbcEsuk+nBubqgauo8Oms2TirzgatIUW6qC+bRwwFjc/s1NN0i/ooxK1g2rosnBZvjkTy
9zK/W1DUXRohN3E8wt7c1u6D17V/z07bg6s7xBLPVGEfhD0GpqtAIizwW6re5N3PyNd7g1XempRN
CgJKsdpihqkT1VBl3wjOzw/Gj/CVc8qOLDk4GF5l8PbfwlIayhGRxhzAoA0jJeKHXHrzd911ejix
44uyhOgAN8np1/LGbMc8+kSXC8bcWN5PdUQS1MZkU5eJMbot8l1Qtq0CG7CgiKZzou/qdxCHe1gA
ZWS/UXKDh4uhXBDa3Dmr7Z1kW+wn7xtkoR2kERQJXV88orI7YCIrRLwm5VP+eJ7Hyuur2luOKuVp
TL/ZHl6nTklYvqaUEEWpiSJnoDBIemsYg7ty6Wqsr2e0IQyHaaVpcW8iKvxsuQpUnoTnf7VzWLE8
OuXDCeARagsQ7sDkV8WGhjEokQUf0K4fDzJdZie0SeEboDUoxqF0/PiwxRdSr8vRaPqN5AlfFLOY
MFJV46+CxqMDjTpGGwiI1MJhinFMVnSaQgjwMBO96nON39DpQHAW8hzQYOjND1cEAP7NCkZOmvwk
E1/4u2/udUB8m/XcOh7oUypOJP28j/OG3g59a7TfPOtQ63lpZvUMt3ypyY9UrgR6xJWXIMQRfo9D
sAlbMCZ5Oi5jG2+SQo90UzlXjpKzQcjqTnN8SpNV2VVdICYdt7da6Z2GwuY31QTkaf33hq8BBMDt
IDopLoZ3bGZI4byzR3C0ur6/OGmrdT1TEVpQkTmXM1HX4WbMxPbY/taS1htw5oaU7PqxoXCXxdxA
ol9GmYAygfy7GR0f4RrWFXKUie0PT86D9mKTcF3btC7TsIBuraloRMj9gDvaLD3llC24055Btqsi
dwZ3gY3sr7H1sO/CAvQxA4rjOgGY1jfyXl5ws29rCUP1xaoeDKslEraBF9wBIRFUzZGjh7PUaT7i
MEG+GlLL3T93Cgnr7UYkCXcq1M6WUKNkAkHM8nBk3Zioy30xPfeQ1Fs8O/PniAbdC77klqzGaoBE
bT/vYA3hljMxTRG61818sh8oGq7GT29+8zwOsBm4vcYIs3xkY/3SUZPg3wdrv0Rn8W5ImQcZezKQ
NrAN+kzfx2AP4EdiaJEJMJBVZLSIfReeNs59Q3xV7R1OGrCsILqCNpS4o/yW5mGvcUvyRzU3Qn8m
KfH895wlAf9AhDjWMt6AJ5PuChE5S10d4wH9j/txz6XF00PYQApdac8K6IIlF3Iq/IlvhJkKy/DA
8OLYeIQ9CN5SwN4s4lc3rN2dVKSAKciVrcVbX3L3JfbIYQSzXaOyBElUYLNvDIYJ6FpTiI5Jv1pO
tIITTSe/TKqPnZSogSkXBzLlvRoy7PYxevlL9KqV3F0gkL8qnmZJibowcD039rpA4OSZNLV6qjXw
ubMmwOCfpgxX/Z50z8arAl8yoLE3Ya7itwfHrhhJLFVJ1z2maUXkTOSLIFnPw2VOlNL4215ki3f3
zCDO5GASIISMvrdmswcCeqB1uhzijcsRPIuwgQ6qsCnfH5r4XTFS4dBf3irYpMnVz5GAZ/KvJzzV
5d39SgDWsuoMz30Fn01zm8nN04/qOZ5C+vhYf8uTNKvbfMPqLa3jzwG8WZXm1MfU023Uh9+VjxMa
oFiFInb2DeFASPljNb924hCD4ri/QiNLwPMxljFQ1hdBbYMzGpbLQnHf5sUy+3xEKMPA/QVVdWXb
inZ61QKi2v/BZcg5dVrIiF8YEYwA2/jjiHHodt96KMnJ/lJzAKVw0dcZ8MEcLyCQ7M4cnDJwHBVq
2QbyulxLzfPstQL5nj6w6VaYTwduZ49Sd+J79DRM5p3nzlv50WqU2OSdnkPJG1vQc2teWn2CDYqL
dsH9sS1kip6sjDrlaONlOF7SkwI56iFxmrIx3ULtl20kBa4UDdJO+4+CBMpnJS9QagKN0DZXBGjl
vE1Hb2KtEJ65AfAR8NsEln4y69S+LC56bz+MvgUJv1/p1P8MQmxjSJ/FuMuWPS61GW5OHHdVQshX
E8TaqCUjjH7DGOQVy23powb3rL2zy8vd6NTERPgrRqc/MwgWiH4krrWAjW5rnGihI+/rK/l/HD8g
Orz/zLJCHPqKuSpEk8I6gv12hgqqWtCxNPA14Z49gfvch/2dJjC2dH5567C5YEMoD+wt032R4o5g
0QJ6dyTXVkbiGFU2dVvzdWzFOLgaaNpqQPFT1ulUQJ5UHmkhj0XBpygVRHHIMMyHGXugTTJnsTEu
GKcYBYc7JG57V8SnPyA4r4Nf3iyrgkl0N8HiG042pfNN3oegwVeGQ8hs3Abh2VSF5MjlvDoImNZS
Wo1R2B0fyUoUvrE1PStxarCg0R6Tit1+MBXApUiAMocr8CetwfUPfHqPMbnt8O9l/GXcblFjb7Fc
TbbNZcjbMUutvnHHNmTPdwngYHrlDHKMCjJgt6GJ1lg+xloga0Kl/c9BFJrhamy+2S9G5HKdeCZf
BMhK5kobh+w83ieAvstgQjnQf7W8JPUQWSBeglEfRJmbUbWL15kxx+nqcsZ+si3aRS0P010Pcjo9
hstEWrw/tXsFbPvVDUtMEHWVY3YDXCFNDz+NaV2xghrxxQg8bFtGlPTfnB4ds+vYvporCxvyfu5n
O15WXvXpZt9edcII/EQfEHJxoGPDui9W8og+UpSfge4nIXGseQSoqQLlR800XC8V58a77VG0iANA
mwm1RS09Q0lKZPxQxRTBxzioXMB8yfiTwq8GT20wp0mU9GG7Lh+J8bB4njeJl0CZzNCLNRoViSjc
j1BGgP6JpSxytjWZ6OR9lLLEwS8uhk8oV63M8rvNeQ4xfj350+9z4J78uaw/QH0YZHKLyw8tWhs3
2srfGuqmJ2d4Rxpc2GtWbZytoIlCa8WQEF2tfVq+jwZzHZcQ30e91OISPoNYAgCEPeKldNDbx+T+
/VR1pOYiQsqbsIhix7b5B/09MYju6yKZop10sd7GVIVJvZ1E9xhGqhKpbPxsmK7zCTnXrS1yKu3P
rFaYkFhV9cbciTU9VtnuGp/oswoCEP6r+MljUrBlet5MrdANfGCQiOM9GU0NTk1OC7euho9c+wEA
a3mfC+gVYU3Y6isHeAnReCuxWZz4ABLZfYTn2EQr1Y0Xy+5unctahOpmOIquBHFA2K9jxHcF98j5
CI93vzegbZkesNzg454ngZpr4zh1nE2K3A7g+j8m84nH0adhYOIkUsBLB4Hdw0fCEkLYe5omHW47
svfjUjonTP7Mg22ehI4eU06dpctxNiZMpuoK8vkRZsr8krvaTKd+k1VO+zFPyXdkM9npOsmGCFza
Xll0ODPEsQnW73aTm6dRdAsmuKCVP+F81L2fFZ75oy/UtZl+uguYYiqXICQegibNh1rp+EY6QNDZ
NbuHfoUdSwqrBZqJJw8sJQA65fFq/q6hgcYQPifvHKtMJqQvlz5E0uHwAQOntrqpvpkRtBYU6c5r
6WbT8Au5iQvZ/L7xpTus1xKguH7G1GLPi1wghYxRRmHgUFyAgyRuf3sF/nyXNzlGav3gV/LElAii
93FjV7x/kAfz/SqUj3c5M9xDV6Dd1TI6nOTLvO0WRUSPSSvCOKYdtlriqBK9hcx4i+NQ0x3Cso3K
rbwzil/qPHmVf/9IXA1sSOvuQdj9wlWe9w2ojyBOllmA34W2zi5EFp3ILobCbTAKLCsgSRgXSZX9
nl/71ECsROo5u4vnzRoetqIYr/zVKQ7PryV8jgzbhIiGa70WLHVTU+j5IXLxhRF9cJpzdCue6fFb
nYbuwUXwD7IesP+eatwnIkdWBY3gByyJXQzHOrmiIm8KW185qYc8yp+cqtCA9gReMrRhnP1R7raP
2ZN57YdDN2MnNfF6N24jaM8eSCUoKhir8pO+B5C0Z5EPdggODJmXfXPtMSch2Pj3Zbu1t8CZtZSA
tJRTlVySXfUlzi0XTGzKZM448SUginghASqXkO8bKwto4OrmsE2X5VAQC7gIdPZ+F8ydlcsaC+SD
Vkai80Ghuh8elj+yVkreCkT1kGPL7CZWldT9fOrhk5JSzLpC7L1mmovVIg41W3dZ7gwi1CqyLnT3
OppWmeda0hGatbaJhlogYIidFWN5zn42QAgIwtJgKR8tcpa2B3CzBu12omxchxR+5XhuIU6IBatb
+aVIMMGsQ2mUiVKThje1k26Sc5HdjDYq1hZZdc3FRM1PQxcXD8JaPv0oizrGMUeYfpFFooEornyp
E+YXkcP2kDNgXt76WgYaBgeUeCNW36UdHf2LxKmloMYmflqJ6w4iBfzuGHRuZzFHi9uBNvx9OeKF
l+4Vx8YkROSSy35R1lPO190wNqG0TW9JnRf0GkSeTEc9ltWmGlzMJmlYynLRElas5PJekDgPkmke
juPja06hqGgj7pWLnGRFJhxDnuV8P1sPrzj/MXqQf8uEa8sztQqJACRHk2h9gDKn6L+h6F2g0x0S
DcbzYVL0rAJMMvrpHfY3MrAXj6ROdcOt1hZMuq9GBoAlW0PXTgyqqmWpyzNo0d1zMBpiH3oCzVPF
hLR8yw295ojfWLsR6Fwo1w45ktlxT8U/47zW4sit7TqyWc/DCWoBth3bKQA1P8NcRR02+LhxDunZ
UWUSvZ78rHa74YwcnyFL+CzXteOKL3Dn6DSm9PK0FNW1rXSACYI3/H1p2ijurLIa7gL89Ei8t5dF
dOofUc04UjYdBeMiSN4MYK/GMk7WhCgmc7SeQxFNnWKY2bzxVW69JI0XvWaprL/HxPO1KKTRcB9E
PU4Ev6ooJvh+Ap+Cfu7whVyanIn0DLsLdAUP7ot0nKGRK+mu+lraULUFtA/1eewKqfr0CbwVr/za
HSPlQWWK7CDo4UDoulilVm9/52624YY1yPx1rNrm8vopPfxPJFZbCL+IrlkchD52qggEozk3fK47
Z+/46PwgzhHMUENT2Nxm1yzAtUUAo8z4+se7Gs8KGIlKcfonfv2wnGV1bA7gKYPWkXdfXTDxwK7I
qR1J2NXXfytfvblsNZ3CsWUAWR8NVAOTudYx02WPGVfYhZlhMYZMTY/9TWg1ste6Y1YMfvC8LfSb
5I6x/BrLLd2TVGtlbhoGkrgLS/6ZicT/4w2n+rJaqORRUHAHLMCHfYBLyIGkovTOIxumGQDLRqS8
JbN9bvGCqQdOM/jGiPQLVMpIFxf4RlLzBahZcXO0pPmV40ol1g/lxt4I2bVpTeeT4wnZGt6aHvRp
VwNUJgfoTAo/90nt/UAtiUwgi+P4YQCAMigyaHGA4AacLjWTv/z8Wies7olxZKfkQ+8/PWPORD3w
1WquYVIytrUqUxY1mXr+u5d5f94dVBwCrVqHtJf3vKCHgI4V3+hh7J/ZSdw0riRZU67N8SMl1OJf
TKEv1Qip2p/4cB70ozJQr29gU85BrTeNVG8lFQpoBwiReMM/PxcUU9fjcYsHsoTDdqnFVahO51r2
n6G+CI9zntbcKhjvwIKUZJyubhpyMGgrnOFkLHTbgroAtzbXOLUyWU6pp/gzOO56YSePNWPPgAuT
lzOC/QtNtmNPJTIWjz6587YNnvhmjPzTMFUBoyGzVImV4l2EDH6L96ds6hCs3RdwvL3bD+WcWtgm
qFOXv9df1rtqXhJCWm0Ph6j/8y9ZbUEqHmVmhz8AMuI6tdELmSOO+ZcU6YLTVk7/zofBmpj9aBIw
UHY+tGpt785SthQYasFhaG3Kr0jbZB80ewi4nj/jw1Bl6XWRQQmCcj6roc+IvTG5LrfWg63kqtwf
uhQiDwPmwbZWMJA0NW6R0CKbW0+eMD5LwZKffY1kuvncCjE38svTUJHSCJ81nIb0VSl1gIpa560b
+ZXjJh/Iq/CKvA55Vh8Zn9DDhNwwE8ajVuKPftHnYzBkSQpLZFgJBmFjmhZZEUx5lb6Dp4AuRHGb
LW+Ed2Vv9ECAj7T2A0uxuV4+cu3RY9v15e7Mi5ER2GVsELgW+jnbKbYLUHm/fahNMpjDVdWjTiM5
tNRFGRs2IotSt697JYwpr7B7V6rgQAkgocVRo77Ary3vL3Fz3y1ZwFwUQBnmPAVAQDPFACc3jrV0
DGMQ0hTBKC8/AgqvbSzqtnrLDjAP8bXIc/xE6uw6Yaln+XefkJkyVyR5Ak/GWWQihhbV88ewlN21
6az/UUpTS+q7gWte3zrNCRgckpbHKjdSuin3Sw1e6XqEq6UwmM3QaHycMAt7Vt7efuMT6lZBiWx2
kJssod7nX9CcjH3/bHPBsTLTC/qyQkAc2spGAEvyhVe5PWYKIGdHRk5ZYE/ZB9uAkBxk3LBdjoyk
WJfI56VVIsrfFWm5V58R5EpHEp5WBEKypvv8bKHua2//FfNJ0rDXWlT6ZSog23JyN1oA06lqsPMr
MlcO49o9XEkyn9qax/rzSlN36NUt3egOW1NkJcCv7E49YJB+HjHJTEmJQx8LWtDsD7Y/GwRObuJS
/kSFf8pjq/JUGA0Qip/1hKkP8waZseoaYXY7s3OCrWglhm8Pd+F6TokHvKqe/Vz2v2d9FXxPvH++
r7FZglAEeX/WaW2doj+v0ZAJb6MnqO7Niyjf1HYstG2grMNi4bDZqEsbwvfC0dKdwSU/5+gQYBb5
FIOpEURumG5uyxT19kaqbP3htTJTguaLj13RbA5pLmlws2r9RJZRuYUWEjT/sxnHLCXs05sUw1DI
VawG6lVGm4BdE/A0ziwmzrd4eyEKESXjcsPQzr6MUPDH6QDZ3/1xOadkcGdt4IX/D4f3Qpt3h0Ct
5qpdqG+gIusmTk21FnIMR22/pPjZaMfWrvKV63fxPtHUCBtgt6Ly96P91PRgw7vwH9ksB6cePCs1
r62SkucMb3RyaEmVoF035fgehV6J2JEdc2fP/OT87hKbUkryi4/ZAxrELKZEm3SnpYq5EGP7KfPl
8GrUW/A5VRkTNWenjtK/JWGJEqwwl4adT/U868nINLZEaTdryuciidjkC9LMp/vdgGV6EnHB7v6h
uNxwb6M/KtV1J8fYU8T7OaoaCNWFz6Oo6rVk1g5JkNcXQtUpjdjBoRx4CUAePz4APMbZHOY9Mfhh
lUufoKuWZ0zTkGjZWxqBwlvqNia+GCi28ilKgDDM1TJVD6+xjlg6lfrsucDlIAUOBMZqxAmwgZb0
zNMYbQJ/aw0FF3UyAXgJFzMRvXV8V90UkSG/50PISJHsOPKWsXB/zqogymetYYZBVEP0SGpXI/LD
lD8CYTxL3GZ7G8gZG0JeaE+nAGVyYp2XF7sH3ubY7ITs9fTWpVvxgYQGy8Dk1nu3GcTj7T/acjL1
geVSyM33JFjNVSLfOQQjBf1IrrZr/CcBaloASaflnHs42ISnYHLUPMlhtf8wFYHnpXcygXV3bUZ+
3a4D3p9U3fodfGoAom6N3aj/M/CoOHyaoJuYBCVXfpZdEWGgslcdhTcCceAiNmThXbz/9RYWI4LI
F3m+O7bgzWWF66UM9gMNfns+14D3og94D1aC13hgcfABq420vlCYZGxSP87rDcqSkz6OYKDoEMFC
ypH6ImRoc5dm68EB2fFYlMJG/kU7jegivzYbntVJeMMtDp70KtYtv+YFeAcLzt08FruAfHfMsYho
Mw7tL31FZloGpZkYNp4rVphAJ4nCtbezR+IqoKb6rMzEznANRrQpYoA8dQbRYE57N64EYJa4WOod
6REPI18W7zJKgfykX2pAU5twEemcJuMtHfCQlmiyCNOFyetHL9wOTlxjOMFusDr4p9/4jR7skZlw
LRJ8CIJnlGKyGnSLMNrQRmcDa9uYt2bqKnbaFQgvDu6IBVbYgyE12ZWxG5OW0dUEqJQl5K59S/8d
7wxeIkWNAviAz29Yda91mDHK38uRKnoHlf46bFfVH6vW8HBYpnyt+7PrYdGyNA0F3Gfwk91NjiL0
hfMm6LVBmUtJNJfc9ZcYrX49HfGy+hp/+3fNxpSexO6263ZrMs42t4x35TOwnd81JjRVFvCy09aP
JzKzLOOT61dzbbTua60VwAoHgI1/qZVIBSYzjuISD5iQY+O35oiDNzvaRhynxHM9cbDNyTeSZ3Np
ooQMHOEyXoQefEHyzb3xiPrt67DJoCCxV7e3U6ggQ2LPeCLHk1O3Lt19YXEqWxZcjo/Jd0GtEv0B
ZV30VlqTXYBJci3UHs3Xq7FnShAiEzT69GrzKlMMCIqijBDvgiMpbuLYMuq0eX+ti8CZ7mtFtOTt
0Nl58UlPC932IpO5snoddDu2Qv9SJ7L6Gtc7qIdQKqv6wJBHwqFV7tRHYt7fCYbs/o388u6pQ8ei
LfbOX9BYrJHdAiHy2p4u0Z8dyEjeUcnb0ZZp2mAoe5QAzhuOBROnLbwoU17rOSlt4z4g7+JjNghB
zVL4vOnU8Me5BvUO45grIAPjKf42lzVstnpXa/f1A9YBoyxe65sM6lGcnUnujPRl7gpvcm8bbRzV
bNOe8wCbUGc4BYaVmg6bXR15E57kIT2JwgIMSSbKlyLpbJu+6ToxsKyKQoVAudX36MTaNhirORB+
ct4lc/3KnKtnK3hA4naPw9bYlx3fmAWPIzVuipr+T1i9nLfl4Xfm44w52H/R0xsSs+3O1dAqfHcX
tTgfAo+RHYK5c8q6sxP26oHv8uBaxgtx9L0VePptQPtNHSIV2KtJMuTrIUqhUBv3npHix1j2f539
kUf0SDV1T3KjPjsGiQC3I4Wko8x11Mq9NWO6REtfM1K3ylg/kmYvDhQnKtSwv+WxVESutBO3ZZq2
wXQ2uUw3fLiNk1N/nYAVM+zDhLfoofrO8XlMCp4HkvqHG2NOzUFF7fBFOV+2VxTTTGh+edKpwptL
t5dTlyjP4GkjJqVGIc3D22Q8iIy7Yr2fm+RC/6jwEz9JzpHo3rMj2V7gG7DQNs+bqsCbe1KJ+sl0
EAV6FQCvkpEVQoSbJYpp6Bz7ptTLvVAzNGSzHdH82NyloCObe/zJyEYK0Bd/6PgEe6CQhlmKWHnx
+75Egwdxpbsb8uV894l3iJrooX+oMNRAnCOMe35YParHn0A2iMDmBGWYnMZi5hGk7af5Hq7AyKQc
BE5yTPOSGRkWQM8caNKst11fa137/YXj9gZAIV/nFKXiPwGknd+XmiF3kbb0pECBxILPXHtCK6SY
q43hmxlyeu74alecg/KKiSJATYM2hZ1ur4VAX/Kk8t+ke0Afs5avMGIBx7VucCwTFmhKe2G7PZnY
VXzeWYHLANAm5LQSSv1XccvYl3tH0af+H+ncEGoUgrnRiuahQqzdUnBCcemroIaBs0H2jHzmxT4q
dbsbm7jywzVQAAFvf0Mi8hkUYBt/K5GzqLQ3FS12DCoPjrmQkkGkbx2UzAn9hhhZKHbJJ2PfSiQB
FCQoeKnTP1XkW3RDguSTHoo9NLNHFuJ+acZ5yTz4PrDddnRfWzwo8dNtx7E+p0bOFXridFYBKQgV
jLnTyBdxLJCW8+ObK9kI7WVf117BupbbC6XJvsIVpVlDZveMARNQlxVgzHg7ENkaCZjWGtGMLeUg
RSWQrwCU/OvWnkSGbJa0bIFZ91Twd/lsDNcVZKzXkVxLLCkyGcUrmjNkAAE5+BI9GmRIivkvxdWE
L03r/tacaJINO3XQtuys7Rx2IHQtcEdmU2QrznCokhAikJbvFsCDUd5+nMcbNFRIAXyllw7TN3p8
98EXwrFLT+ch4Hnkba5NlJXPlRlxeT7nPaYz0MerpqxEWW98TKM5m8tAeqbEwWp0ArJaC2RKwPa9
6lD3tWT3HPKlG9GZlFVp9w71m7+EgFj+R6hDDBaC+z+lYoOVVhzW4aPV+q69szfvhIYbuOZCcXgR
snzWCgPfQX/cG8hxiElnUM0uwpCNsPNNLa2b3FpOgOUlqYKQV35rUGsDplN29uAfUFQy8nBvblz+
C0VO6HVHIIAo8bFyr7eKywIusZiOZPlqiSsayoGbanDhauHFAQ8TkJWgCLD6X36OeQWkkoNWuYiB
4rWXN+7xwE9P77z9SfM5VzFd8mDGWLVgS1AKEXecIHUwj98L89XyRGLXv8FVFNfswtgJ0TGKlObe
rTv4XRAp/TwA1DppmgVM435aghKxhL3v2a37OE0P7JDMajPleQf0SKFHrawAZww1t6fpwq0xy4il
UQMC0G1xDzXKKOnwhnFipRKXEyDQ/SOr6BHf6C0pSQ6mGncRQwpUNtdjVvDdRXx8CoxByJISdhvr
+mIT32+M1aiS8HYWp8yRk3lrymxC8QRYp1Vs7KpbwBznoTnKL/Hu//hBwTZWspdvvYwwkUvH+vMs
RJsxjfCOkgdO0YPNYGT81IZr3wNN0OD9L6GJ/Bl1YXBpE+0rVWiKxwSP/UEv6f8vPBF0ITno09bQ
1IowFGPm98OAv3c8zr5gx801zZL65enFi6zqAe4xlWUR+qTNwd7TVKFmeeVjE333qZo2EsbXnWwm
SrbCMw6gRB1mxyEdCD+EeRwh9cD+wrrUHRnoS6+jEEJBAQ2AMQd6Oo75MhgGTEVa8ZuVzdAvudXW
ZdWtoxy5fZz8aLbaqJXQ5UQCjduRgNHY+ENMovQfneAmhpnR7fsXaGBy9UzDXw8DW2avVR6WHpyB
5Axb4Ul67q8aElQxsjCskhrCKccAYTNQK+vmnn81nseQOWbHitkCpmD04Bho5nS3T5i8S8wqXZmr
FfLhCQpPQHEuoCJZ0j9qMP10mhxx7sa3iJUzHpq8wzSy5sompU2ZyIPm99/vmaVyFyPK0I9SZL67
V/OG64ZWRp3yYzMrp90sN1t8Vc66aFoZEtOFEA6WpW5fYgU4jFdqLMptaNdgrgBQNka0Zs0ScVMo
OPNkLb1BLimE3OorNS7orvdzRK3tFIPRhDjxs2AAAjT6DHblOYpHSMyTwzwiMG/nlfvplDsDlxR8
+cV0co2jAcB6n8hmAhMcZhKO0p2BYOI+0wgfVs9vo+N2H3P9MW+wydRGNWSbYSXT/2fhlLvOeQtW
k6nb1UR1AzKvxaiZdop1U8h2bj1CZZ/LcLvsfa4WAgH1YBwL4HjodfBYmpOPxEmqISJ2kalxMtEr
S+6uGrg9+W82O15Yb+oTDby28GXZeIDcQ3cycODCyZjghiEk8YdnktQ5oZ+Wyx+x57rcE7z+Bi7V
M7TF5ohvGfz2/nxVpas1eoQuSkCdC0apZtgLAJxZpUCCUGMT5zoHPOjhXYYDzVtZAuhCr2n20JWJ
GOLCWG9A985RG6gPJH7ZtdyE47jKhLkMfQsOjPj21ZY6KOmRMSUwcNc3WojkYmaBcmU6kOnfDsQr
9NNhdu6a9BdQL7W9ueE/y1fdfLz7fT1oE+iPHtV9Svf3nZbpBhQEclYj/l4JxRfqKUSTuvjwJhDt
/0FIHZ3/lmREmSgACxyrOOU5qoUNILvZO964FJLBtj3opKTHUMcEKyApjCnDCLiimCVg1l5dKCvh
tcrShHXOMFdzfozRnVZeBS1CX+bkUqqSbkfMhXWPunewQtltazpU0jrbNFI8IvB7JnlCWO3MbNZz
eVC7T5mdpMKTXL1d+h+BAUPk3dUPqYGoMX70C27QYzRT4qwNjdilUIDV5rrwx0uLGtQUu2VC+6wg
M16dQaWI9jTzv3fjDOrWjzas4Wwrlj1nYN5xrgqEwYSR7JXph9mwtMCyVFE8LUyQX+jPcTYVKJlb
FpmTLatvbRI18Zc/Sj07DeT0nL43uNqAQnAzSUDwU+zBa27tnQFKnLgFjDoQQslxKyjgnCUTNtB/
MPEqQaM3hq3GQOhVRwL+EQsY4gxSmg831Hpma0vXW5L6/5PWRbWo/7iSLUN7wObDHqrKW4HMou6Z
8wiVzAxqScI9i1FfzGHV0mqnGaWjWdyPCCvZOKpYbPjAhdSJLEylabo+BHumZSNPsv1fSag6l8p4
JqcGdC11nqXRXfS2emfN+Zk19ge+r/Fj2IqSPXExf3wcqy1ax2x8XiYldAE6AxH054DobpZ0MhkY
RQpo4aUSh9mCdvlEHYepjDDx2NOAqmx/3rdsRl3Ht5Jx5kp0ZLP1F/9zjUkbTKqNmz3WMs7OM2TK
hU7VlqKTdBUntJr6S2MYhY5T8o/r8QK3b+gaqTLn5lA4bXXy4QTv7dgo41SItZwoKqIAMLxcyxdr
0ktL2JyF/B8OpNPMgk33gDeKB84QGvWIu8gJ9ewciLbGVRfnGx/7M98vUuidpM794tu7Cl2pbKsz
w44/ykQ+hIIpZTXSZ3p/Ro1W4zB0wN3FbPs9wqzeIw2+UXBdnKozlaeT8HLsl09BHv809uYo+ch2
b9X6apb5pbDtS/FhZDa9Firuf4RaYtHb3uHfo2QwXjUKW7WvHfhZCRcK6wWA3lAKLa4LutYeOl1V
swL34VPl8h3RkMtDeJU5R9bXroEeN17tz3OYdeeC84Fm7ObVxW+06Pj1zMdGPn3CGSg2e7LubFF/
qiXYExrbYJZvaZgoVReKdNynWmYIUrjjlJm0Pkn2mcPw06/IGx2pHbPH9bRqYNGCj9lD/zl0kaHb
zCMYT8Iy1k9QtlQuRizczqr2SZtJF3ndoTEMASMZ5hDJ62wEO+Gln7Cnfs31hKXNLg2kEH9p0Hg9
L6Wz9RdgZZvpr2zNGZFcuBMFice0z+VtyN3MKOI1aGLgxmjwJFDUFcoVBY8ZiKRQzc15WjBzohe3
7CRRm1HAarN1OqCc7JjQSA2t/hUqE+4n4sXJfmDJKmPsj0W90nuu5pW5AUCwh2YyV2GKbr0iJWCR
aNKR2AKKLuxqy3PITKZNM9BH2N5qYhH7mgiAo5W8sx1Rt05Ug5VuqRUAlORU8Dbb8pEvlPM2ZpHj
OQYYe5+9y+nrZktGz3d3ajEn3WFSyc9KiuJF/1jCojaq2ykIBrBcPZSMQLRD2vrZOEGti3ydTPqP
SmDMGuTtFCS8bRX2tIIoB+qGq0e1Ny9Dv9HEKvLrVfdo66Ij5UAJaL9QhD/ztRtaOXRKyJJ0mCvW
XZPKoI2H6Drn03pA+ipLJPC16+r+Jayfrtrp6VaKlq66znLeMg33/ARnFI4aQQvs+RWjJPheKba2
y55dhS/uxmX4xEHrLv2TxEe+/IfSwcz87yQSJqJm3xv7ZO86xUR7TRidWIb0DcHHH27XaezpCu2G
WuMBHzDBoRrKl26wq6PkmlL0spyUtGRJQOtqeNXrHpuBcnd4AZHl6CPalr8rkLmm2dLJwxXDhZ3R
fdrwk6qmdsDW3VQrBFJNvJYs9uSxwBc9c46dJKbJXXCSDp3aM9rLpXDVMp0q1oSuykzbkscg6OWA
13TbLwpmFVQFpulY9aAg+50O8z3AT7YlCwWudHRo0MqxoX5eAa+fwTQDvFfqMwEn8jJ5CCan8kwT
Fih11OyuWKtey1DgBAYZL1nKZPsNanj2cATUC5H0Ky0/zPUbcJaISRLFXex/FI+yVr+LKJVW3Tml
sY/sWiowRXDgskETF53gCHi2lgjASVQRLOWEisA3+9RcvNKWQPgpaH4FNGBZ0rqBT6OwQJkAZgws
1gx1pUqnQlOvryYEpRSaJta8wcMIvy1R2nr7zzJ9ydnIFQcJQOzRs3bw3yO4g0dStpefbivuASAc
mCiHCLNhNhWrGy+VJ8ii/nPCPak2Sqw+MN3IOIJaR54Y4j6VVAXcH+VloOl2ad8ZLG/8JAKFOFLp
uk8VtMf60v4jSBwzbG9Ykn3xBZSBCec8icf4Nr1vkrLaBVh0QR38mhq5vr0K45sgpGFr9BMm/HKa
UYYt+o0161D8wAv6jtH6TpNLZ+20LF6itBeZKU5EqMF+HbT3GTHu1joYSphCUpwqRz8xkZMPQ7IS
O9GkhLkO6UDZrdl28ThaLT+B9kzRlpr1/QkLr4fpfM91A4rk6z/XdQeFMVjkzOXD53Fpy7mQDnbg
R14vqMRSntoFekWTwMh0/0NkFLVvwICMBcwbk5XAr9FmKBhNiv5d4h9rrRq/o2lL6NGfnEl1d9ZP
4bRPXLW3DKb6FbaMs/pGXW6OVhJAQeEXgrx9+BUxKDmC1NtSYg0IKr0V+Tzms5/cU3NI/3lENvV+
BgVt9btNuzDIXM0hJ/C5fimvs8UIfyJJOqpdi6FzyRHsb+MP2Ry4/Eow3l+lTRI/pkHM97r4OGwe
SEWn+Eui1qYVLJ9TZDqtOG4hIuckvKQt2VXa92+5BAWUZjYaZBPgNRnFCem9QxjTQG3cpBNj23nu
19qnStytEtjVlRQ23y3TQu/HDtgrdiDSHxPq7NSjOtprdLzC1/R5+TKb9JE7kNFA3yc4x2I9RDPk
ZgFPOwKK3OYcdtQdBHW3xf4oCl2k7GiwpI9Rcaepb3pKur6F5Ctsz2/O+fQ41XugEDzoS8mGtP99
M5beoOc82BsnF1GMNutOqMMo0DtQBZUqcz1mbPe5xsUZTcexm+2a+r3Se8ydCwixXo470koVY8tK
z0EVVpLDb5iZhY9yIin3/JKsuYZF57mDpmN0Z3WmFSxkV3puemgPT7YB0MMKkfMv6ImO5ZErE5rJ
SaDb3qK7Uk1Sa+DTX8q0kCDcx31wqdALD3Oc/QX8WkHaXJTKhyKcFmuAGCtJkYotfdWCDWk8cZTf
wLCfrPSQi1IsbIKvwMaazo/B75UZClQ8bgvCyf+X54qMjP3GNceMrxsXauwFXlsoILX4ABbOr3Fd
XG8wexuOlwnsG3Shu/27ygUPJC/RkcjVf49brOOlwsa1eox2VlC2OyOpcv9fmoZadUdpCaMzJS1J
Fx7Osfri6WZmFuMR/ZO/Riauw+/kSAvTQvxuHTs0sKnYDJaZVHltDH5ciQ/4MDltmMa9FzQIfXqm
MDeLaLLg24v5f5WRMNGETLWdjq7kmlX0yyGmJNwzxEb5DMkH1Ia7tOSKxNxiPu3VXvzFuWecje1G
o5+qO+jpUPEiIarAUErMxS+AunMx1t70p9rVC4NSSGE0wE10hsYWkQQnjbac/4Tyoeyef+vuS/VZ
3ESNlCAtqxemYG5Ee4xE/pngGrmLESS7vz0h0wFdHB5ClWlg3GU9ic4nCo4dRGZPXddGukdYAx5x
m1Z9bta6Y3yxr1YN23o4Bjmraw7d7PtLtFzG9qeSwyIlP8zvExcbuymaMZMHf9NYEWKFvm7Cp+mt
Ow90Z8Rg1jxPvwp4gXtYtYdxD0GIJphOVb2Uo6r+9B97wNnuXtOmUC/yF9XEWe+Rbqxy9Fsqf9RJ
z5LhwhebjQrxVUGBFZTHiEiMQSx2JL7zfCLT++ZXu8V0zqyeroTDtAP0VQnkqKP3Qi85Isz2rqBi
BV8v2UkaImfEDG71uGifoReO5Vyl0gVYPuFLKX6P/CUhgnSZ5KFDepxLekDn7eORhxIV9NuC8lez
iA9ViAxVAiDnI+iiZB70ieOSJwCh8LLXiDc21hCoPIFkhSlwUgSuomOpm8TUnmE0sERXpsf+vAiN
3y/X3i/HM17GHQWKcD7ixeWimvRFyjZEAnOhhl0TuJYhavTqXOQCW7cWHPS4EXroGVBcd/U22MmR
pw4MTD3ZRGypEerz1Bzvqq1zXqacZpGTWb9R+7Ib2LX64r/AtYLK58mQfRLJUh+v6A+vw8b95iMw
UEuwZ6AW4P3fnlF556F/O0HHdMrFm4tPhBYeX+Cy7wMWWGFCgeCSj0msLf5bUmweEnbV2ID6X6he
6awI3xTrHe/ZwcpqPw6FtY+lXF+LYkZwJb5I/8xXZUoGYMdE4BqEgGUuMvsgJL1RQut4IupsExLM
VBO6fjVm58mo0fuzPRn8tkt8LNRn9CnYxQCfauICvs1Nn+WegTAMhgk4CUm7tZ4rTYHTuJE/CrZB
oz01VYdVH3FdXqmXrMYtu3LeaU5cItVlfGVZPAbY9L8Bj/U9GaSqjgLiugpV9cXzDPaA447aeAqE
WuAgSASqy438qp+xMHiEItDxbm8lDjZ3yycliMUAHAhHG3ZWVINpYEMeGneK75vGzpmjDPLKA2Bv
wN78u20AKZBPZrxE6XcwSZAnRSIbFJpZzWbzFJDKxk1uRj26wAXIBLrzDOrrah1h5vDK0GqFEZ3i
iYjFuClDdqmXwGeY7N73i5hp2HVnQ9LOl3b1Bv+o5NWVmQpsAMC5ElqKRne6Zn9x+M4s7uBzGtZP
9Y3KMwEPEUoN3FfQkKsXKvy4NUsyLb+nFk57X8Y7UbH/2PiBKLI97RBlrdJ+11FYpsu8D38iTFGe
1kelEuPNeXNuLKsMQk+u+ns7mZAd1j7304EM1IYdaRFplWNXt83j0pIrygQVhW5Yu3gcrUiqNZFr
ktq35ZVBciOWqDtaWuWRaRbjFAtUehahVj92Lp0iDwTcWxqsSVebAdyj6CBX5PxBpEQdnaC+Qzt+
NY+ux5oXEnPQkn1ZX50mvXvialDlHCykD7Y7lwsiKLTobVgHBloIjfi6DZUHuM8VMcbjLdmu3WtM
ja4lc+REMU4ufeDcSP/R9XeJb/VJzZwMXHh9yneonu5+9ujWqABaZjrGQE09gJTJcHtTIQoCRHga
0pbUk72WC78gHyQM7bs2XP4GRR0/eWCghQUwb60dc+pE4pEKSdRTOlx98WIBLInnV5WXGRORLxAy
lTjJG3rqhamZ6fKo5mXRyI60/cCShg0aCm5q+XSl5jjsvJoS48B1bgc65kVNdU7ubD7vfPc94fnP
VJ4ZRJ9sfZvoQnHEMCNaqYlzA+LRx7kiRrUNHI0ey2hFnb5JGkCdzEGmAFgfNJ4E+mjpDGFROkr9
0fzO83ISpPMGZsvOzQ3WKX5PWJheYsQex6o8goa30+Hof4SnkYCIMsrstk20VOZ4J26bEoYhrPiD
RVOhZaEQlnHsGg578MRgRAXppNcSB91seFoIiYEa0k94ZsP6SOEOId1A8Foksfi++95emWvytxqT
65etScPcvrwpnn7T7IhRJZe2IZArNjIkvY5clADF7Oudd6bt8jVeX5yDOeFWwwwnMVa+8688Wb+Q
yN67RjXietkuSoKeP2XDTHAovv98qEWbqSQpUC1wofBcmwA6/1RgkqkTvQ+ygEuGG+s8LazMtPJV
cuUw2FP9tzyRZKAsH84kuWz1a3ahulI7jCWVjtEDd5jDLKy66PachORWr4GYWQN5zO+e8qkd5dd6
Q8YeLBccMauAE+KtO0nyRLp3dYTKBNgUjtAydnUkkqD4SFO9Y0t6C+3Rxrshe7ONGDUwBFpfUvRq
SkefBvm3csgfKJf9ZyW5LDS6AIfrPjzLoRm6h9bKZdxvGw2he5EUUVldCibu7RcOM31WodvrU2nE
rRGieok0IoVRRKWNPhoo1j0nfSkJNe2kr6/oYb0n7r3WDnrzBZ/r6yENaPvxCPmtSbDqJNaoMMfr
LQEYlUO1ma3/5uKu2uQzcHv1IOzIXQbpNgTge90ww0dNyXTefILnM3MM/uXbIpanTnG1EIts3qpr
iRiX6sdUCeI9buV9ErRIfudnnTEBxttCiuD8V0UjqClOg0M3HjgHyvddBUA5Nnnv8YDTBX5Nxztj
l5dJ5QOr50gbI13EscCzDcfryv2ozgavZ7eeJghXUlLuoixdXsfgmm+SerjWwaiSQXXaE85BVFLm
kk83yxvwpLk+pkJ2ofsa7Kaajy6OKqjQwSYNfM0+1kZFhhfl/g4rRhHWE7hreGR2rCM5o9HWdU12
0hgpZXJYe4ZY/y/N3YjvlF2a9m1/+u/37O/+azENLkYbrl77LiFkhSLzHFBEn2b+98iwI6c91DhK
hmHDzY/Br3tNSa4lJLcR8Npmo7o5BSAr23PpSb+Gs9hwhB2MqFhHPU7X4PrjKylv6teZigSM8E2X
V4f+8Z2cyDobe4NXQD2qp2NXI6bU+LbpiLVXy3GFj/VRZ8E9b/vX7J7D/BjbkLiKCiaaE+RMlQal
74lUnF3VcVaaMc1n7Yv/3XWQxBe5qKyVh2udIsGRxNOFEr6kaQ7RQiGLDm80BwGpI7C3H+ICa1R8
8wMMbzLp5dvpy0un2MZoD1n4nw6oibpugzYINc+K7n2SLZWGEoNWOr9Tmmol8IyPBzUl8a9QokOR
0zl+EKDIcBqBzDPxhMjYa6al+Z1GO2VSpdqoShTl4b7n32tluwGsh2IxU9pXvR3VfuknwyuWruVp
sEz79CtCkCrw8PJuaQ6/mL+wQs9heCNHHjE1w8Jk64+vuTVWo/I9kU8TkPuOxSBcqAMdkNZGfY8G
FlIpzbiNt89nAhSxK0GoEBVy1V/3ZhSYbaVpBnjdgYc8PIMz3tNO2qaJOYPFH0wPu6vZe6J0TTJG
V+6SH4QeGYwDMxUWwocn14jokqReI1j6y+SFLBusMDKUyGmCxTRHyzxYqjG1QwooDmLTb+QfRogn
138Y/ZiJT0aKJ50TamOtS6+x/DXapIXm4OKYeW/JPgxHJSnK/guRCSh8maD2IouJTX4yRRNnwPVN
E0xCuwhXENl1VMEHGq2F88sSSWB3AtVhASRPM1WDfxLdt1KTrHVgf4Cx6JKZeQh0cSeIY2nPrdYd
IM7ZeeSwsf72zUPi48OdG4YXDqCWBs7C44genVgyrjnJNrkNPG5+qyVLx5UmE4PHKj9+qRm+4Q5P
cFDPexsgHyilh4YvwoBWiV5/gdmOdhnd3qwf+NDop24Y3+x5FmM5A0KgidQ90PvHz/RE8g8Xy3nm
CI87Txau/Qma+7N49IDWT2vB/pKRZSym0HMb1fyDIInRge0qPNRzeC1+3f/GrJvIqECoazBZEWO3
jOZGGHlrnpIbUrNoYUMNW844KLecobV2tgVVnZKBX6tVWr0SSFAvSbPvV02by48bZfRAMMPZnMA8
h2OmRk3gGN+KeLKnH8ac5GRWNQACuJXqEaG+GFavMikCE4Llr6E6MkgORWxakIfAU4z0f5bJNuYX
aNyPySunpwuF68NtSgZBgF5Wdst/GQEi60WE0R2FUkMzU/obJXu9G2rAMr5hokW8bekYC+lKhxgk
0J/jboNSMXFc9vAC0MowgJgf1uOhOWY2HroG3iEhoqdiz5lfl8+q/NzwuTv+VfMou/qDrIOgdhMw
FGUMLw/xcmiZpDj1FqdwYo9WnC2PeSR9b1bqPk+g63meQ9T8eQ3QyotMZeXYDyrkQ9YloPwAe+0f
UhBk8SGP+DOdF68XYkbxP4KzYTOw4felVAVEb5nRCdXhHaMcE17PZPcn1RvdyoE3wRHmzvWYEWS3
F5xkeMtS6rsDC0Ktf9Axa4ShxRI9jZMMASfjMNG1EPAhnhrckuP1lzYV5ugVRjqr/8IFlzAHHeyO
7xDAXm0Vn0Bjd55a9VT6QYqvFZ77k4hVruiEiQGYZFXx8iLVhwgCXoYQ/AbRF8UAZngAcu9vxiWV
sN/W9EbaQQ5mNEf6KhcFh31JYxO1oS8OGl1QwDCdQPSzrY8BEv9xdmfriR+3r4WmOnw7PJ6aTbeM
h6xypwm1sXnJdgeuxYSrjDM4goU+oc4bM3AASU4rQJu3KXmMi4xqIJGGmzzNEyKX4q35HPnAWWIP
JxH1wBM0hZZueKI8ao8pqdoA+UXaTVrZIJRIaIb6PMfLd69IJuFshkrMB6KlQmOjedoR+EW2vsnL
HH+e3Fw8W1ykHhFSxiXqeh/8rSmVKGUcHGzaYLoAQYdCxvYkOAXhSi03A1zFQ2vwU4oZcTIJcIJD
JlM/36uqNLeWfJYENoGnvRtlGnSe5ce59woGzLCMtm6QiYXP+Lot4hD3DplzA5imJZme+/rOh9qm
ALF5NjLaCskJXp6C9OMxJce9AqiCK2vRjI+okUYPccUvLFSkrdoizn+9HtrArGdJA432H8mqeJ71
B5ZHC6xDKqW7QCo5msfeVPlcw5eGxCWvwDca6Rc27TVULLWTR8krls1QSjxW9nm5Z9YTAGveVrH5
wrgJzthnjZEbKQvsjC826pt8eyz5UuDpO8I1NNwvi6BiazZ2QV9O40opL2aex1Xq2AgcM2E6M3u8
XE3BJoOWRj8ze9j8InM+ejhCP/kD/+cta1VkfJDwzjguWclk6lQ4RPLE334nZlxl4A16Sb4onJQ1
G/NgOpzNhUxGM0Fyxc9jUTucOx/+7I7mppmlpZOtb+aOZCtm3q2nT/C0hFPwGWf1iOKEciimW3OV
HLlOlzeVET6ICC6K+2gaVKOZbT6zTqOoC9wlG6dIedH/CYmh/hhFsVZKmlZ150zgT/ldpJUK7UFp
TBPlLVkW4Qmai1jiYjaJwzIg6hXTF8MwTRhQObUrprLtLo8b/x6n49T/YqdlsCYSHtTiP7pvn42N
ay0rRdfv6zVEIca4eI9gj3GmP4474l0UuJiJngrOB5QWGtkFsiUuBv2KuthDdHOzJEn9Nv+ycSVj
9Zjr9jsMQdbkZhM7XsBAD+I84D+aByFNEiVY2t+RauXel6KWey4QHz2s0cEqWZ8/8QP4m0fvDz22
Et1cGYEjINNEurojf3y9SA4Th5gPMeUVAjykFRTAA5IN4q9Bn4OYh0GQh2ckkO9xq+nalpBPmA6S
xVa2/IzRhcBG0n7tgywJKcD0ePk3BgMReN6baixemPV3sjU8eyAFjJM/GEQEpcXJyA4uJSAuVa4v
WARZKCNyv0PhmByq6VuLqZXQkRNwCV5qwB+R/sBf76JQ6eCfx/QOE6C7ovQ1qLZTft4yM9wgPcAi
qazBbjZwE6Qt/FwZJttJAHp6+QZ0tuGC6d7jaM9oeTfEDyTwMqElLGHnPLPsNOeT1RKK1yxkm+Io
EGOUEb04Klomy6o7N6NLWPWzk/zSVYIKAgL4UEGCUCRU638UGXLry0P3xwRj89T9oswhhjLzcXPC
VHK+Ll9UpgOxVqhDEH4QW0oijEvScWXnKPHQLrZfZ/JN6e4/sRBQG/md+gAMSLWB72cq6HRlpyi7
gEv4fpxbalufxC7cvS2qK6MmA2/iGK3WlpUwmymsBkBLRBth/pSmGugpcOuIZXJ5am34WdeEy9q9
bjFtXavfPcacXKhKEHJj1euaygjN5BFnnsMy3z2BAo15NKWGzAtOfxwGLQ0mcFovex6v1iy1p/ri
E+iSB/e7qtBC3dVSaiFlKKRtid8HSDrA534p/Jez1N1e9YwSPgi2hqW7XBLr8mQxv2f1qOIORvq2
w6i/ofg3dCVud90CYCYvEeb6SqCdTRznnc41HrmW96123Q8bZkycFW6HHuMEhVxrfdi1jSin1vGB
5GO3gQBzdh9v3v561JWmM/BNxCez+szMavYWkwbfRF6cR2PMny3Vy++7+9m+RaznuErdCOGVy93v
EpRW7PR++3tohJaHeIDQKyAjee1ECnKIed4/AtjCFGtapJtNTrX4J1roztlTl9VVqutWfpLtzIhY
NIfv+m6nLsFy2MjzQ3XtdUhM2ryQ6FTgcmOOfDwAQuofBZMRCtSEzowHhaJOGkwN5r94Hg0odSSW
3ub6gi7B1L3rCdBSF2u6DBdZvwU6CqSfrYtivOANUda6I1DsN+1c5AWd1fsMBF6qF39cjKd+hFp7
ea/MqpozEgjlns7Zu4qt3aMax0O4Vfe/rpclFD/y5PHL9V72+ZGId+1F8I/4bxulYLsqJVGXZZ24
pzKNPfvLtBgBYewm2PjcTaqBxq0SbJXSo+BSzNasdO2tAgA4CF5E2lLU+7QNSduLWHemJWuJ2U04
Raa05gJKS45b8tnXCXFHGcaz1uTY+qeRz6tK9lKdk1PAIGTdzknBccR6ke7OgKk4oCO+Lhh9OKUs
twWVVTRpC2IS3mHm2s1cO3TInLnUIRqg9mS5MHgDcW4eX0b6sE+CXmUw0JXFSvvjUBrITwGxM0o0
UrzDS8tFcElqxlFzDcGXth7RcxI+uMS3tM1JtwKOJwAraaqrNJ+vrSakiUnVy5kUEjLDl4TdJB6/
ZGQ0A3qGPA4umJa/l7g59zxC8oJyscr7fDnMK905RQnRCDUSaySt4UdHmqwWKkID2EK41Cm1e9IA
nyB1qN4g4Zlk3iMEesRHWi6WX2TLAFu/wYgAcS6Ma6l+/3BwTy7eM6J2bINvd/NaG5DI85Q6QuDD
HhT9yII0eWx0XQDLs/m5TcUBBAjbZAH+vyLdQHZKmOUQEt8OlqfrPwXjpqeCkflB3f10h8BuWBJ9
PSkD9kWRtfNsl7jNFwpzZgzyI7t4ZdbJRDdN0OZaqbV73KDnPs3oJUJPhDW8XjBs4UPUcAK4uZPA
XqEQPWqqucU4m317omGhmsMAQzWkiz8oePL8KwXpTHax7wNR3+ysZ2IqRpOAOcuA9W4XU2OpLm76
gIwOO2hMyw7+dXv0+LiPC1BoOmh+jUilz3ihci9ZWW6B2xM+e1tWmBM5IDZqpdX9/xQts7cm1ewn
IVKBR3aVa+FU+/eEvjdHPhzNmhhg0auF6QSUq/3EyoIz3upNADL3Sp1CHw4KBMfM2ifBCV2DDM9Z
EhOIMso8ICNAeKAYfMv3PnSCww4w8SDQtPB2TxpH43kFLj91LEr8Krshyl4Q+iIYJPQXMJ4p8VHV
8Wry1EC/HPDgUPceyKyftN+H++9Ul7rwjHSWoEZMmux8UJTWlqd2UX4DFH+ZOeztIOR5mSUGUlmA
dCw51ciOZpYOY/ik/cV6Xl15vTtH2T3HiGPTTdEs43JT9b1K6KQjxyv2Bf7pdMBRttvrRlLbcu/J
kmG6TAp5aeIe3JxWxB6YdKUnXOtIKu50hWvVgFzL1xI16seLgqk711pGtAzYBhABCHok+pG+cyKv
KVWsC0t3JuCjSbHlegcrOnXezycRvZDoPaXIRNYmuAiPvGJ/YYoY3ttRefQPE9Tirzy+C84yhpw5
ocl/vHNANyAJDBhKYWLz2MHAGP00pM5aGsOOaSxdofT04ZnEvy902GHVbPWgRfhP3npKyMbawM+L
/nxG4XclEGgSzltjsuhqBcpUZuEJeXzlKnu4JEY4oIVwJMOheXqsgRl4inrC1PhuTxMBIU/KwdFl
hIcGgHeZPap5WSGaRlO5u3SaE4vb0J9KXFgC1HpumWydiytpNmthx3/skqXIHqbGhUPIJxiOBMjo
WzXMVCmsdGEtmtS60jRFQWgK/WXHo1Ih1zqOjJ1DFYuKz5DxKSrS95nrA4BPi3Aqst+jFOzm2qBY
BbDYTam7efVfNnmN6kIv0W6J6KW/0XP9+eDaCfhNjW04cmzYaSAFOrt6YU3FpaJHay1Tu3sMCmSs
FEnHUarMUcXy0m42R5uEIm2GfHW0p7JjkP96180U2Q4/PxonuFMLlOdobBUxpqa1aeYYK52piTM7
gQ6ey4TkJ3DOVWMWuaIOiSnEpZmZky5c0u7TN3xP+3/jVZx7TfL5IkglrZ83vd0D7vcPfuvjGrhE
zutXEsOJdQdUFMpTHqXk7Yj0jMn/WRUGwtFciFX8Y6gSVlj4Liz5A/M/df/xTivINSiEaBp4b0JH
izxYb4bGgdLQSoKaPuzxTvw9FI4mIQELk1ycws9XmWhUvyw72//ys99HORY7Sg0XodV0JPWF4990
XrLuRzl1G9+CgSW/YKlgtTsUT07owECSwofwo7fsVRIpuB1IrBnRZ3FbBnCOsixuM+UO2F9ocIAL
6Wi71Z1+w7UZ/PxrFudJ8ddFWmT1MgbZMPH9VN7FstT9znAeHVnL/m1nqUT/75TKvdbl1BMvtRvC
YCPgToftce7zlnyybor3lv6msc06nAlEaoAc7Nb+unHWnyWd/yQAqcq1+i1dGalJLtAjKRQ48Aac
THEe/kR5TFaFFzqBxof/8W6XpvvlTTWGitA/+rOcV1Vc+EwwPpuB3eOa49jTr6zuxfkPeNSC/Php
rJIhecc//bFEg2xj0Q62UoNor/BAGQI787XMJCWi7gjv7EctrJRkQDNof7qEGO2KqutdOu284spA
FUXIDx05rZA+V753cKa5uibe40Xwtnhh4q3uCqRaD240ffLpqvZJUaaWvxnkGQ8ZLj9Bjv3BHFDA
YF1+D8dPbCzsZKjQuZgMW1v9yksV3rh2uWk2b042YnFR+RdwDnO8feQ5E6JzVYCydwsGyopzq1za
1URRqcO7AW95JfqKp9abgGF6vnAfKL3+61o8xbVuMCZ6lxqeNar/vznrwoHE5sDqCJUJAOSKL+e9
DeF9K24ihAIkZVrVY0uJcaZkdtBGqONtqIqpHdDHqUIaaNQ7asMicufIvpm8vEYdG0yRu/rgf5xl
WRPu3WOmqiNptgzaHexf3/C4y2I28bk/2Jc5erbSGTexNIpAR2hPvd8+5WOrH0dYknzepb3YaDyn
yW05kE0mtZNcMuHyQFgxxJjRyOLen3JRWX1msjN/XoIAUg0oUr+H0iT0zP3yF7HEPDZ2J1jxfCbu
pYc/auh+P6ESlw8gM54OdQ5BPyIYWLTgHpY0cA1Cr54NfdNorodoCO/Imux6YZPLRjUOyheOa/7u
LgjMPX5wOinVezbLmMEd1GKZFkT0lqmPE+keFiNeYCSvcX1MgrjcXBtYoEUAKehrzG0hbNwVuoGD
OPiB767Tm0pcBQgzI4IPXQs8RJu72VByzCIv9IRlr5uMpjsLmonykgvlnfbyu7XQMIEuwur3FUIZ
plIhSF+yIdxbJngdwGf7tgcKlFrnXuW0EdxQcDKA+Vb6DbDexYshs4xHq7im7RDv4VpfFAhjdnUI
7XBFvPUzhIUOw6Nt4PPXqDSA/0a0tcKj+nUYq6jg9yQgm1tzdAytIVtQ4xD5lHw2NiabHfh8W6jK
+edJlhvJOBcijzZengBZZD1uqw26FLZJxUNhYIs+D/GMAe41ofOPr2ZFtVVt6QKrD/idwYqvWj6Q
nGR4X+cyaeSp3oIionjrHHZS5BSypL3GPZZM9oe3POjgOFiI+kxIcgEE0qbvWT+t74fg7GCVETna
p8LRFhyCwQxgx3gmD7DtBFq9CvGuS7znLSt/3+XJTBQGoTIJ1mtL9tw9afOrfTualh6W3Mq4SXjj
p8jg3RqJo/MHi9ojEG1/JBKoxFsaSJUaJBXai9D3AMIU2DiEixvtcj8eUgRHOPbj1CH77IERi65T
Ucv22bXiop2bm8XetUCWSWWGl0Od/e/OZUi/U9JdJ65LKafy1x63+YeZSu0Ca+3EpsqVS17JPy2S
hoKtmVclDQe0AyYl20+blKfAt9FIVam4iEN2iuAwzd9Fzz7suFoAt1O32ghx5uaLCSbCEkEmbxh0
TfjAUyQVo0AIIBpnjVcGT3MTNllzlmVZ7gvoPDouAa8uBiVbR+7ciKjFXc6ygVHrGQug8BovCoCM
5zj2gXaHya3QL7xuXi76EKuNSgRq0oUZj6rRkXscKLwr9+b/LDmrs48s8FRsSJNJPbDeI8leX3FG
d0fYZvFsI+Q+HDmniYI8P7nvPBdDZopb4Ow9axr76HzdVjNyNRpQVViviRAm4zJwijxudWccm/5k
b6xjgvOyabHlAU1dMDAvgcL1T/CdnQkwi4FF4yO2OicM2rJW5yt3TbXyfvXDlvOl/Fvk4fjyh+ly
tXxyvyvGeVNPzOmfKsx6KcB9ubm3wxKefHq7BFW1fYvVYHB8++aqZstZY3kJU7wVNt60UIKox8jW
4pMIc2VacUfRlXiDibtEYgXIOyr4rNUStdrXDxfERzoM6NZE9u2PWozLxFxtRK0AwgDg2Rx+TWKi
vMLUazv4aR1FpLcqR2jiX8OYIchfXdToug9hmp9lOBnxQpamswxEO5/OIzc9wNfZiQPwh5lR9kNN
hGmym2+8BE52XvCFGndEjC373IofuJz6ieuy4z6Bop5/qaRXMSCNn8b1swXkHgokAe09UvwhORGe
mnpwfdeF2EzDIQhsCmTmIBYhF7BR5k6RXmgTpayuCW60h46VIXnFE3SHoFv4GHwurH/bNitU8SxD
66SpXxe2uJMic0Lo8jk0Q47/+SnRSAP4Tjt4JQ9x0XA8a3jo8zWc6aybU9XNgg12/D9inx7ABAbg
5/I3oBY0WU/inoJniOwPm23nTxYAn64q3pXKAY8zS9udwB9OEdNmh6QaMYK+bCCrpSQ+W+sHayj7
l9gVnOVVgm50DC7k9y9EqvtGd58ArzAPDMCAp7Kr9ZWrO9FD15Yoqkrfnqx9hYV1ggBnMMnOH/Zu
UhMDu4vThLajlxyWPQuXjyl6wsfTovEbAPeW2i435xOLO+OvG8VT63GMUD8d5kHQ+oKGDrhrUI/S
YjTSJMbVbFj7WxVYW5E8+bIR8/a3iUefvptMJq6V1p2MaMaa8d8VymB5OdZidth/05FWPNMAYu5v
tK/nvwcs+EyU7Jh09gyTrzUKMIyw6zuY1NJ26f7xpBHSkjeLbHaf/krlZi8oPc6YMDhzUQhcKiDL
WnoqFgYGy4Wcs7VZjzihEnRb6fAcoEK0hOz9nfo6F2hqXE0+qffmWrsiaW+JcWGYX4YYN4kDU+na
3EReikMVrLqr2XT/XBBGFQdHNuHMSGS6upn26tqivjZZvIoCFpK5yTnaspnYDHtryZYXm1E8rCnr
dQRsBv8bJ688iNgq6QDst57VDUNAVGBc7R0DwFTFFNuB01gZ3tpogLSpfkt8cDqDYVnpboYGiCG/
tid9rJf1UnFCNaQdtz+BD+C6MFT0tuvi8FfVFHNpxb85xIJsRlnNrK5oEeTY9RAerH8OISrg3+5H
7IvA+EqaMANM4OUMbSLmGY4vTzeXfIf3s129c11/S/rzAEerc+Rhi5/VEtcCV0mTGUAYek1de4OU
In307Z/+lDWXU8LqbY2No7/d7BSAjkrW3uSts5QUKC7gOJJ0P31sZYxfj8JpS5qPcPn8SC8KaDIC
kWyVHtVtUZmhC1WQ1jLnrNNOykO9pjX4ezKVrYKcOCQ6BYIsEgvTqeHJuQKKJ5F/gcsRaXmmCPw+
OglWtMkf/Ow6VnITmnqCokf9DKaP7pCSdUTCfec63Wx5TdBm8Ank+7PI7J1ED0tb0URVnCfrqj9d
v/fTcUYbGjVu7Nj9vj9QiA3m/MMQ+md9Com7tv1rL39fnF2XwzfIdoixRm6gbFpUnWeRS3VPtg0X
2eSHN6N+uhOhnKuJmduLY8pcE/R0+Apb8yYB5kTIgZ/vwrsY+Zs554/fTal60E0AOlnWT6r9+t6Y
OZLv0daGftT8rRzlGnTAe38I307Al6FYIB53xyI6S/ikhQBPFYSSn/WoTsltZW1J4UVKqxt8f1Ee
jcyUWmyXDWhO/q/FE56E+IN5mpfylU9LSWRYU8thSMlMXu1hh5P3LFfn7E9MaVWxbf3COXkNHbVI
5DEpsWS3kEf1qKe6ieocTqnDLidbWxcdJFzu23xZAgf0KefNkhYD4VLevem2mXCpQzr+wIsYizK4
Uirk6nTjJ0P7qi1HLk4ithRqgxDXl4VNqm1AbY/e83X5DlcbIrW8H8BKywjWJZvj+Zvp0spr3Fiz
sY/aNONTMEah/pTtJ21DiqrWB6X6a+ZzQ3ou5iWevRL9mLN84xXt6h3XsGcpjK1s95s8UmF+MdIQ
cJbDab4gLla0LOc758AhsKXbLnzZbT2nEVYlwyHI7D9w/Ok2RrmmrNmrjulIdQ1a/qEVAw3E4IVE
2xmNdjqS66gOQd+8RjX+rPHX18pX6LyOd2M7zMCSrDnJHZDVA0GfQFxWnvDzhMQTHQxGaJ8xnqHr
WoynhkSq3o7vMLR1Vdw7BlenESn19WaLdy21Q79ZAWGURHgOXA/0Dew/u0gyn6J6invb01rk8gWt
DZhY058K2zr7G5Bb+tWIphKwWThW3qG8Cek8GdDJmU0KOM6BB1+Yo+vO/FAr5Tlgn+ykb3Yjhd1u
sRcnR5BefiRUnO66gi+1xFNCqQEmLuPH/m1ghvHQsH7nEHwNi7HsfhacL1/eMDkwHk61NByebiTe
vv6KYMeCYe/kxaKAGOOt30ymGJJoZ9TMd3FEQBbVNorT/VLwWs+syuEAajKfqZmikhBj80mcMW9u
Np29HwN/nKhleWQiaaWyNUt3lgb3UHzlElec3K1wNpAzkyli97t4U89Dt1wcOkzTocYmKMTv56+j
9cin+wepofyCmkrpJpFVY2MKnx2ZzCi4B5RzN/lvgT/3UBBGqbvLFvKQlkrfvx0LtbK8f0+B4k78
lWRmHveJz7U5dssGiUPIth30/YXnYK8Ks5Rp9Yk1Z3chY2/8r8atu3iY2D/X6ItK28uOknQyBxIu
Flgc17os23GTVGiFbcOx0wWccv5E7cUYVHjI3A9RFdmWxu0iW20qbQKvwiN3xAKypDqzbRZErCKb
nQSN+E9dTWrTOPFyGKGWVQixI79haKL61kCMdPd/oOecvLJz0kV/wlHouSERafZPjEGRMFf3cSzt
mRO2ID+RhFE7xlrD7qtdQ1Kwafpy9nSyd7Pr6a/3apPjp02T4wamqwSHoii1N+SjIrj802gSLbA4
NgZe0frXgiWjA3y4Za6LezK9C/w7TFXyacIolvOqPd4Tuvbi+Cn3zQcWs5tuUiPfZK3kmbOq/bur
f5tOg5qMPrR1WJSjZ1LVFUHtkYjK7a9INqbd8xOVPixBmtaFgrT5WiJg+T38rBgB6IqnPy6tBvjR
l2FWM+zh916T37ZnS48kSvbPaqtLqFDih+f5Vp1NMYCV/x7tglZ/r8UTC/Y9hr/cygP0UMPFuKwz
61TXwHtFKKVp/34+c2y6RtSRn7XXYxYdzGzL5nucNrl9pCQkh7YVa4Lzo+5192av7rDCb0um4yEk
RVv9jyLCngAgasi2PDPsjas6R0asBSapouy3W8tx9l3ok2ZwX3Nu2v45VOVqNr53dwg8pMl8oUZ2
cSr2n94a/h4b+qQkrRnaRJKmljSnfVH4X1/o6xDqcSg4zbh93uDVXqzYwbXe+jEGDvcUndu+hQps
DcdV9e1FOKJLEudswBxqBXNnccH0+XPIfusBw9jM41PDqdsu8TULQM8GBGksjMl6I7gPkgjZ+0u6
4C1I2l8DkKldORlXaeT3ITQ0+YlGymHhfA04seoHAN1ck4kSX5196GfsaJ2Ls1E79LVdWtKvdTqR
YaMlTLr/7fuTrD60F9Xr0MrNxFiujAJRwbF1Wi4BOZp17II4hHAS//xC70lBIpA+VvaV5OLPzTaK
4K3XqRXMAh8roN2vuOoNhOd5ZnuAe765qtBaTMmy5dUH7AGY+NsXlUCVcgzIxM2SQf3vAJVeBSW7
MjOtCKgUBTqcdGPDfG3PACggv6OD9jCq+Fsa8gkQn9pIq40FSvlU01pGgkGXL+uZxgnUJKglmd4v
fNSHOI/vj8NhJ9Zr9lzCPGYUrjx1nqFiV5JyMHVOs8/JpqdSp7tfV/3jyzOIHcFJb2psKQJGmhgX
lwnrXsEx5tzG5UA3jw0Q58DnppAFtij9UxoYRVIAmCcpe5L90gQySu4Qloa/BHwzjIU1A3hj79s2
/204jO3zwH+PZxdx78WSxvPGPGXCgUQbk8qsAO5nm6UVQm/D+ybAOeojB86gIjM2s73ikOf6FA9y
7nDuMPSyP7GH+pN5VPhj3ynuOziFtK/LppLboYdzhvakV/hUmtF+ZHt9F2KbC/1aBIiRqjifdjpX
4aqYVyDmBY4VmBBiM8h3QefonmAAJhhIdmrq1ofTFGp+FSzDrMxrB8wQfLmzywJh38ad/463sdnC
nHyaM4rYBukGvRmDqBnGw9TTayI8PEqOV4y4xC61e3RMXf6eUcilmLfAff/LeTHPF70F3S5ZwdXZ
/pjFPGJC87fFlsrZejfyIQ5Jnp0l8Gn9cLciPXrX8Pdctuu5fczHXi5XjPVdZNtBOwv0tAzYlXaq
RG6ZPTDQ9IBjzHA+2Cyu3IBwEvyHThxdabR1c8occK4IIHBqjZeDYscZLZ4hiyZ8QDk2KvJMeWQZ
Jkgk6VVIpnGASnjZ2dSwJVtVMRqDax9kbDv5iMzm0BGTt9jWcXkgGrO3oLmhW349Bx51v5DgMU2m
5y9qBmCmRzkYJ4yUxmD9tb3gnDAmM2TmJjBwTybVaGYPsMOwZj3YD7nbkuhCFkyxXvDsIs2Bps/U
f5wGfOzt6QDE0YbuI05i8ElqXAvghGfhA/F2FOqhQQGAcIS+68oim9uQwIJ8t4UQZ58186HVOTAQ
w6ch+Xh60K//l4mmP7PmRq2mRKjXTfqeDk3mQuSwL7ufsOIwHRBfig1ZQh2iU78v95HT6n/gzXeA
0TElMmIl3ty93NDQIS45hOn92wZ1Rl+hgyUjVxmkzGH7ta3h8moZ/6IqpOrXNqV2wv55firo2K3S
5BWHiTyqx+2ZisPv5C54X+fLkmV9IADCsAismiPMNHS+XF6FH1uFXBDiMYogIQ/ALQIAh1YXntc+
J1xMtvGW68TKy6qSYGlKM7WDafXvj3fYIKTc5LL1Z3NwRoDnj2juD71WzovceATa3/iqgG1QMnh8
RoZu7WYK/smXk2w6lmscs+CV2PS607IeGx/vKs0/1EugJiMWK5Rm/dd3PDaU5yrOIfNcxeaQ5WdZ
AxKK9YownN71K2w065cs1Kqr+++YVEyLrFPt614SkRYHn2i4bHvXKi22SLzj7yg3uaktCIA5vKWi
TlS5I1VCqz4P+sRmyJO7FLvfdEp4sSabvezGzwnl40hwlCE2+X+1i4pxh3HmCcProvyjKh8srNPv
rO8nfx2caikcCDbhsM0l6P3jo8uLpXAvo6sZxOsG72kS1To+x28IAPjQ/4wzEq6MuPTeLX33eIc4
9s/bp3WeEfxTFHzlaMA8JakRXxmbDgMqilUO4/6I7dZ5JZpmtgUrqBmu36qTctOZdM7tqIFaU7Vo
xBNf35eNTAQuUFiG/x/SULlwVoxwAnw0yfyyM1rs3f2NYw4M9bxq8nBv2eRr0skIUAv+B0zoCIQZ
AnhNACY/RCwZ6j5aajz7IfMa0BHIFzXqbGzetBFdsttCh6zC/LofUyGIy/2y02pWYtn3zCu2oYwX
RAtNWt4qvNtGgchgABqv9mxEn+znR9PWU9hEQGyfMa67g+efks6ist4bnFtiGlWR/FayPnZgVVCl
gpQ7Z86/sqOqvvvvu3kZYYdti96jGd+9UKZUCIrEj3brXf7D8ikmRWiQvTbx1hWVLw5B37YHpf8/
OIo5L2r/oJ/374Be8wRqD2sWvCVEx9TsF/rUOHWYtHlpHSe7QxKHBNyCRjhphhb+Nw+5hibMOgYq
XtTsDxsk0/JtSTZFph7BEQ7XNHs875pXyMemSmoW3P8wymUFzH3mu0FWI9aaeRUVb6Cl9ArFSD8t
S/GtLL9QrdotzKtuu0qWPTZFgtXxlBTEOG5VIp9VykUNJB0t28uLBC+xVeFzfi3iEjToG6HgQ3/t
JSm6PJXNe20r/Vz2RbBGNOMuGyGxcpzpMakUqRZOIus2KFGqo6AedGtN2ML/7ilvPzmJWo/SY7py
ZANXc59I66LpEQvDEO6PBDqAB4nxd7YfHp+FzEAiSA5QN1AkS2xF8Tyg+P1lH3kxLcofyfws7OyO
aEEMU/qpMo9f0XF5mGc7neVDnFOQt0RI/ADmeffia3tSfmXcRtcyA4UBmuFAobL99cWDZpBuovlg
a5pHyJsXdvP8xCx/pqC89eQB31nVZmHMNXSOM/N8J+xevJ07/h1EesjfqHXZjXYffv7cnr9doFYV
+e4T+4ilBg6p9pI+8PE+L0M+WPMdh4VNnvOaNg8SxTbsvlSgog/JrGrehoLZ5wpIDBpFwrQG+9O7
B7Wmeo0nlnoz2bkCMhuQNLFS8EfgyLMyJ26ju/NA5ugMvz44zHzLglKWaFLB7Cf464gQ+JP3m362
zO8JETwbeMGvQOprNESOEk3iQNYkO871WL2GUE9BsYcX4xP5ZMnXHhu2A19nk6NB9KRCnF2pmS9K
UtVkwnaVNMVoSkeQo3hHzRtQYyoneg4Yo3G4rUWvMJtXNQWgbwj3zDsiakRcqTTodfWgI5Rem3jP
YjdhlBiW/eIUjCgzNzzIR0CsQQVNcPBAE7+PZpdMjNY1WbZWXzdm5nAmTcZ8P9k8TQZZXMKilQYh
HowBr5FE7GpTE1lXPzpzgONGXEbtuSrmX2azC8UPlbhp/Atz7ZRUx0MNU81vMYJB12SmtOA9n4Du
1so2dl/Lds5/VyTm4LPERFT0rqR1cHKnESgCJ+KZJ4Hii9MYnzUXUONRzefrVvu5BB6d3UoeqnqX
ZnEpH47qb0qpFxpvdOq3pGHFuFYgkaWhg9Yft2YlAnf2jZZKdWISkUaaodDermIO0SLRhmVA7vaU
hXggnvQsmLjtyDX9iClkFcYGcp/ecPtdmYn/7cIZ3IBfoe1g9gV936Z/OB8PNCdQ3KbC4a8lelbx
qRkzXZvJqZ/EZyi/77ob0+uSCjNw775WWjQcHUqhQuTTiAaTKSBa+GVT5BLj09bbfPWNM+NbTNyd
kuajILfRQlmTVo50Z030XY3cBSZc1l9KHfbbYI7PxvCuzyB1dO+WPy4L7ehf2WDC5SI7AeUB36mF
KY/TZ7JVIymvTsPyfiaBNKgqqEVG84FA+uUdz3dA00244khOxKMuQOmcOEadlX8GnoMQedPLFkX9
W5evle5j5U57JJa/+Y/k/MTv1wjKlYL4CSS7pciYeTF1AtCxkmQDDbUUZ162vnD7pA6+ut74WkPN
9tC+0C+WuaBf5Ls97Lv9Fp9kstIedztFJLbNBdpFyJTT3S6/SpDFDw+Ygxy3wphvwPT08i1u20Mq
Ij4QvZoVXO24dgTz+PAVTSsvLFogjqoCTCAtEjLY1ZXb+PIZxPjRCL4ZKSa8F3kNOhk3txlpLQFh
RJM62ErlTxorboYhJdJUzHYSJvFomfK/g/aekkC+NuqiDunfF+5ibuNWW11qsooB2s8b2Yu29qih
7uwB1yVYhm6MTtfxohePZelOJz/me1xBH7TshODrdikXKK7zGDMidHhVDczkFQgFdztJc+FHm4NS
8nSyLwh2RRKxDsfI1LuJ5hdULk8k8MdZNGULSZ2gTwvBjssq9eSktSMnZCb96eDFRrKupabTBEte
tYoOX2xYvS9uGpMOqje5WkkWmiLeRU6ZFu1E0HavYkhZBAmnhZcFCUOlIo9uEUVly8r4kuu5WtbV
FvdH9oU1c+5+WItvTJXnnGs25ZZRlptDCn9K8laiM4CqTzouuUzJRucDFZtIRtQdN0zVBXSKIM53
L3eXbsj7qc28EtmFJ/RJxlDzfxKwqUCEWXl4RdGWwWHCP9dpTFBqVa5wDi6rrQCX+896+hxlSgtM
1qkbzNjX/BZ/YBvUCY1TkHVlNByijABWJ1roEdLPHmgNrSR/Rd5o0b7qE23rYasKagBi97yMBEct
zLWoQ4e3iO4n6meY5QA/RXeJUpJoqObQ7lBlJdr+5gr8jAjegmzEds53RpxtxD6R90x6OocInf/n
HFbxw4PDia8/aGr0h1nZpeYsqvU4qvFfRxuXpHPOYRAwmtwozCXl+c+2EXGw+ns+KNJU8lCJEUZC
Zm3tvgsm/xh+6dHVYJgvYf1wICjfjwk5pwrOla76mjYNq2oi3peayss8hVN3foqsMDKpunYok9jO
zTwIvOTp6qvVkQ12qu1XUAEkgtlrybGZKd1icDX5ODlJfW1CKVDCSjlAs20ywYGt7XnFmp8seuiN
gSL+CImFRDP9UwSPx14us/MxvR3EnDncKnyUXG833fVpPWlwfbWyKsgMLdH/Va04XoX8I9rQyO0I
PQHCokfHY5Wm88oQuPx8e5RdomqMZas2bJsV0oUln7O4M+picY/pQP85TpG756CRjFJtyEkFoQ7E
pfhO8p5EAS3p52+GlsSC96jli2d0aMZaLcn8jtmKKZcOW/RPn7fqQilSROxtpos1A+BzL7HW7zWO
git8wmqfKsGGdy/r87ieSLACFrdEtiNujKlDTJ70DERRIz4JJjtvOQTZuMAHbDNGvglQHEnjo2qi
cJSv/ajd4/ARgXi2RwytnYOk+Gcs7JyNqyEPUZMdTixO2Ehy/1OCNn0J00mlHOngmcoBtZq0sCyx
vGOCRJkSdBiXQyAnjaiyJqP0pZHj0F8g4+D9Pk83QKFMNQuvXBkg5+UR14qQpa8DsiXeCAgjP79z
K+WM4WwUfy4Unjf13gg1SNT2HkX6P466xkjymhcJ3FIuVBJwXH0NuteleUQ0OefjME7c4UuSeyrl
vevkI6ffuFPOHo2XDrcGLjLmfFiAqMJ08ftAmbekw5uIuALpr8n2CAylp4rddv7yzZ/iACUZAtsm
eUFbIF8Jb627et+wqRWLCeyfTZSRNzq8ebX+Cl9V//3TdGYZ8IIe9CGoQamqv+cV7E7mmFcgBtFI
Fw0mQGdrl/7s2x5sXD5rp47M1RrAAmE2MNvo7H/fXklHW5QxZaXy7Z8SUiNKU+dxX7B0wwDmsvqR
Tf/WeoHw1uYKUcT185mq46sjX78z+lrb3Wk2l7eaUaG08r1G+AjqLFBvmRcu+GRSS6gG1r6F/XJU
eX/sBEvC+TUDg5RRiuw8BrDK45HYN7YNGvvPd5tly9qH2hDvXub6FqYvCkJAH4mNBBWA9J7Fewy6
q4PwDfwIIoDSStJWkswGFa4u8ZsQy2/8OO+xpEMHRaApqlLwNgigsJlV0Wdgzg4fLcaK3xPAibEB
Gvpccxg5Po5FsEbybbzf7jc44mKRu//hhWsxjJ8xjrZmWea7A2owD86ItvtdKfIOXyPa1SFyJPAF
QzjXItI3i3jdl6CA9SPgWJ/kaP87+wStUr0DNEzXu6hXqFDQkP2X6zCJ+BBb6L0i2hv0iJ5zqt0u
pFivYgcyV6OSo0SMRP/jDQoYoHjHMtMnDqCNbn2rdAdmkLwF8+KFIbfZ0fjQMUp6+JtxV6Qz2iDS
LH1Kk8B3GZqejTCqpzSAJt9mVpESRkuHzCIGVsr3OXRZeQ1lK+eAOl/mtHHrvK/aXVXMvMV9bXmQ
0D3jnWwA+DVvGTH8knR8Jsu5t/Jq+4AV/DNThGx2ikpJOcPr+I1haOUUlML4mZONFF/IPw4ysfmj
P5Yx/SWPGsbku2wKDi7yTX221ZNvhUs7Z5E5VF1Bq8XJOCQ4DOWn7/ByVil7M86Mgh3arRj1Uaf4
L16nX5+wW+geWj3IcIiX6kje8+ybfHubgdRQCLIITF8/HLm/Hc1N0x1hZyLzfTifJyTqFSAgBMEF
paco4PGehun75keH5xya0dLKjop0hEZQa3I1cXIzuZB29IF3gfbg8Da5OcynVPR4d2ATJslji8cq
LOo/3XvayDBHPmKTXsUCq1jXcd1B+Y/bK7dBhuenhZvQdN7+xiKxTjMXjOzPAKPfcp4yoigcoRyh
Kd+Fhe8dQY3ZiM8nMGMECgKAU8fH5AY3B46bTaj4LpTCyVjF1wswSGYQOTy1/3VTqKkba1me3J3k
sBLVXrewy6gYsL0jl+sGppFteJWHd8VtPyhn0FgUh2tKzlsfqliZNYr4sVFWt2K93jDUoDFSNGgQ
DdvIsz9OQvO2hUyBRzjNbwLqJCA5Bauaz4cKDHMtbiHbHASvcjohScj4UNkF/SMHhWln8q1mL5kS
cv5x0e3n82VR1Z8DqlT1QJmOWW70M5QCbWiJakSP9GevKbM5g0x1srWRsKfL6gXxIP0wpjDLyJGj
p6PHxW9dHb5BDPuEQIJMwx9fOElgx5VdpKRGTvlb4Kj3zULTwKAfPvfSDAksmnH6MTCdhKe37KS3
cvEBNlgqqdM5RABdkCmXL2S8drpvNQQuA/RmgpXvvSOEgTIG9j0Oo3q2K0XFAqK5T0/MfpKbBJmE
nAeJElM01sMIB7Pt90anUENGIoLBrgz90h4bd0TuobVT2gzdGgW5Wp0tdx0Jc+f76uOd/3uLaANS
0SPFQ9tYAup9Duz2krXduiX0Ii8lAksac2/PbV/AKNxt/bTmRH2k3tVmgaH7BXxxOp00KvR02JMa
F/n0cPq8raHIZA0O4D46eNASfAnumrPAyJImqt0eRCMnmLHpl7afcj7gUJ7yDY4esfUDXK3rRGCo
2xCXc2DOhfxJoB6vjbGNgUANsrat2qyJgKvBUTTJsyO1flpFtY8EFPmUmH22eEnIoo//fSXaSH3D
nij0gJFOMTjEgYcI2bj0CYCYrnj2RaDUpR+DzLxu2yLFS5+BXU+dLHqrQaZ2rmc3jGz1MjKqUMbe
dQlt6g1eGwjWC+apMxlOtEKLkQh7i1h9M/Rki/7JHpOQrOX5j/k9W9mf+oOXadepM4/BXD46uLe5
72mXISdOyY9zXoCxiRIXvPupq8Kc4gXZlPmeeKLQt7879uwT2qlw/rVuei3UMAQuA3bclr4YRcCd
DrtqUFOryXRWQ33KWmolEvP9hoSdIc3m/NpFxOOHmKtyDjUR0T2hBF0OpYiS/P1Eo1DEQu1sXJn5
cCv2/JliJfGwyEnkrYZoXvdFVElQ68k5pArzonS4vxancH8H8FuhCM75goqkJMLWxB9/cO3u9WvW
WLQRtAHit7ypP6zJgYSzXpVFd6GFcIRjry8Tm+Px6oQeKaPlXMaMnsdgkvXC6SX4JnnwLRuz5+tp
aibMldcbqiRu3DN9sgq29bodM2kzPAzbfbwiWmnJBZyUvTOCQkEN3Mf0yW6azCbELI2LkQ2ExeUh
5GuMkmWkgkYcE2mAB5Lq8eoOZcKXIz9wdsU29mMRdznVnE/YkJFvlJ04rrF5PZGcL5fIOjzAKk6N
QD0bK5bbh/KECe2HwIHHh/CK6wwUmVZ1JYen6x/B3V1EpdMw1CdN1mIf94qtm5anIHGnkTYRbXzh
yR6OcwHFHiM/sP7/iCAQ6+JuTGDom9BCzSRs47NSEs54PgVI/KlR679QwyRtTi2LK0rkT3pPjLxy
kD3lmCfWIcbqCymqxseRi8kOxvfJuS/Tmcxxoz4ANQQHZNzSOPGzSwZNSImVPk1XpUMNTV8XvZep
O4k5Xb5f5XqVtrTGRMbFb0WD6jgf1UFLTm3MDeIASFxSbALaUhiclJPx72+cy662vt/nrBc+FUDj
mMuWAQn8TSuPvwh+PmQ6ijeJ35teZMSRGF0Ntvhfdaftjnfnh2nfi9W35RIVCX4Rz5fbXon1u+LL
DnZjhNA0RrYS29cXeSET6tfgY1NVB4Qs41WIaxWn0fiob7SraUukJPBxsqlIVJ6LB4Fvsv+q2pKy
h/8FL+lnWortAqsfgHshBWZ3tdjemurWIritoQqi5n1TRnqnk86n3kjf0qJ1onhjCOnEDQxsHwCn
EQjoqmJedza2B/PjJAviv1u+i/KrdtKcAHGMupsAmWXqto+D1if1C0UGVaN8oHhj5y+R2oDpSyfF
xhVaylZ1OYMaD5i1MCb8mc/+Pu2ddduUXtTznDeLU2pp6gCFMsYypVzWYFbzm14WE7lF+iubQZ7V
mMCaQDiIGg2UKXQdS4tBPcrN8/T37af5RKj9XAiamRi405waHMPEIGEyZrXr8miFQWukvkqlAC44
QqM/Mu2eLP0dfU2hiLa9YcAULwMZ0Bi3TapzGInu7uR8/r1ge0PmMXHcmfujo6srO24jBUqrjch4
OupZkVLHzzXEx1P5sD890jy/ZrOlr/7JRfBTaccxDC/fsAWlmSq+zvWQcKf5giwpFlWLXtxa3l0+
V4MS6QEV7GRKkB/ROlEfPYUUxD6QG0ex3jYe8LoJkTI/Mzy3s9YXRviXHiSnExi0eAvIzllcoFFH
B4YSDTzgFU/OfCssdC1LGWeUXv9573uaDH9dC49uTc5pIQcgHLQvHT+8NotILMfUI9pXqs60FZNn
5KunHbY0PrdRslrWy1ozFkTNOwWostHA/xGxnv0CBFpfhKeaRzXfqPa+M9U2sZPP+SjEO1DY8jzP
jMLhkIy72XPSw1QZ4R0dxO94nM0ROg3Tswp+hFBPzVTvrr83fBcN/utiLW4B566HXrlC3XBdFRg7
+5zhN/HlQNgEFqnHk4pns/i4p4xQcWlJ6HIqBZytdVZDVCrffiDrhCo6eqU8c6r0vhtfwQd4cwCG
Yobm3ZAkZmAfAN+LvCL7Mrz+IUa2j52XfHhFdMZUvQ7Y24zKoxSTbaHkAnu4qCMb95MC2d8tCaoa
OPa7VVH7vxIWJCsfXaMJOexqW9O5/VTn0Gz8cb2CnyChQZ5tdGD2tViEkZHbbgSXevuYONwqtyPl
fpchpmtno2+IvGtoSKOGk+d1Q+ujMcxDtvNmk7L5NzwV8JUnWtZIdA/PrBYszAli5R9spCoZRN6w
45l5C47cwxf+fImOwGhotkNkpPmu2MfVZzAUItA+t7QOdMLj+zLcp1hPaOhDMmHU/VhGE3fqX4IL
xEYcpIJ7u+nCQQv8s6jwU8/0QD/iU63Mi1RdBVokucwWZ9EndzybNv4fclYEU4cuJrFfGcKRkkvo
q11VnCm6O0+PC60NGxMXOtoRupdPADoW6l0DleQAoggwre70naATLQk88QgXe+XIFGL2h6WKay+s
8c7YFoOaUR+lfa/nAgMqIwmxN0+jCrtOBr2xMQszsnrb3paCYtbV9WERcOZeUSNcZfybi4b+Zdsn
HoHFunWLmQkK969AP7N6VQHv1IMX0/GSGwp09MwXzi2Sv6tPRFnUisJtBBipWXH5VWISDnhmUCk0
PJwDjlKAfZgw5kZFQRo4twA9JFBmCKfN1TYgGRspjCIGa1Zb23/HzMnijUhJIJC360NDyCvu6fdf
3oDmdwRLYbKd6a4ZItB5UyWqio7brsqo+sEaptXS/ltwFRhxLn80XSgJkL2myhQlr41c5wqBkhIU
8c6S+RiEps6SHWjIowt25pUqhIx0iAyqA0R25NrA2jgv99Kd8MMjTLlSKeM7LTSZXwioUUC7xHS8
+4L9n87tkPd+LHC3G7IFQC9uDuqvDRjNggcVWjW7EH6gnbxVFi4ECUypShFBxA/nHVi1T1mkuMY6
cgb+s+ZLRDA1qR0YVxbAQe6vaXJwjQvVU7Tz08oQceK5pZ/CuhqswEYugBis6IeHjJ4xE0eS1lal
SJ8lcBC5X79pQxpmP3Xm1bR/ibezZ5PkAFRvAtlPYkAwjhn51m/lRDrLYNu1IR/P11MosKL3CfXa
qw9kbClueyC+qBsgGznYuIljzu+GUU8obgFqjJVksGV3yZVAgP0Vf916xI8w7FJVpptxXUcSC+4E
sRLeG9FRnWembsfYOvPXP4hCezXz6OOc2IHFYlmARAeuyW1sC0HVWzwjFPUQRTuyoyW8GXuqYacV
6CEKEDbDMYkCOdOESNU+pmfJwK2Grhz0T3lZqthIXHNZwyiR5Jk4oN7CaqrMzU/9fY9UPQbk+Ap1
CWq9MJ032u1yi8G676hTVkqKCbdMR2kMb0IsCkzrmSSOKtEC29DpfgKkzdAIbZyXyUnqKLkQtgPB
A2Fv9CFLj/8qkTp2YpP9hInW4AHENVKX1xQT0lP1hngg/6f7B0vnd7lNqXckqdDJ7EYIk0xpiwto
UbXs8XOEDB/m3cXrF3Dt3/vkbcIwMb9xSQB4c6A1TOVt6hRkZbK/IJvWOVgwa4SIFtVBrjSnYBH7
zbK9Mc/fGftnJ1LYNtSR5sCTb4XjBrBSuVtSHc06dQhzby/5LpcA9Wmv8lFJ7zhNHB84IVG19g+f
aHan+BXM+CwRH2t4vq9sHb0iYOOs3DrtDLOougrKYMFj2bXzUTbglIKmYqRzjJ7oxiDTs+doNorf
R2AmSNHNmowKMAodGZx2CUTOdv9RBv5JQHoB1JcZk3SBe943mJlbekd03Z7E/uI8TEwDf/HwFYhf
ng93SAEHC8uP5NpwRm6C5SbgWKabyFLaYXZ4wj/8ikCROBYS4O/ah5p9dFlhNYZmsOkLKiL10feG
JI3H7VIOhu9jmoO1+4ODFyOGFFUho+5DCbsLZ0eZ1MVwojAnAutEHwBudVCAKBa2jXZmfxCWxaUG
wgKFDjZl+3JrKo0AsFtWljXhu9eLVvoQAUUAAeq+LxnerD4//F/cEUdBvYdepaFf1IdXmyxzsPoZ
//144E3ZC3N1fyDL4HwidHGF33Aj61chN9FULRhImBNFDLl5LW6QQfhUz2IUClywgaT/RYJl5yYU
gQX3TuNLzpVBm5OYbiZQbeu25hvGewMyGK9ab2vW1sf9QHwv8FVtXbQFP0PZQm1SBSpzMO/MAtb4
0RY94BB3TBQTwy1MOHLGTxvu4W8gn3puzf2Zsx7sHm9JoSaLs1ONfXLMznmS/zHxP7KpZ1tgA1De
ENWJYDWTuUxZCZGNwaCznESj/gyZLbQDQrN3t+JcKFqdE4eq8Ucz9AoeI1DCGSSpACVX5oBvbdu5
bxSHV2H7ZY1tLNffSdwhPAl0ISAr2oHZEHaMMq72n+T7nfEe2baRukgQRx8RDdIe/+EEeqPKEQHi
I5n05QUF5MRYgSZHeyO/kJrTua5GauI/zt9ZFPBZ6YzY7RCs+zUx/qcdDBF/GMX6PABECNDHieUb
WbnXqq5v1XT6HfsS/gvudg6D5xnjlBfpYIE+rtK7Io4+PoL3mpk8fABuxyoa8WFUUCovqL711mH0
PZBB2YAqaivR88E2kO9sM1Kcy5+UziBIK5Is544awqhDXGcbgwVkquJjo3NC6ggTXUQtq324yq3D
2g5LQZubzkS5TL/zVmGm0JGgr1CWEBhBwPm+NsjLRLCtTRT0SxjUorNLaMCi2vMNI7G0WKPSmHKl
fLRF3ut7VwM3OCeGo3xWXzCkAlEcGjnKlukBKI2M7eJpEVpJSzWZd+ImLzaLmlsEx/0f2A1XByu/
iao/E7uGJyaYhbkjlbSWmqp+pm5Eb4sfYg386biWxC0K3Aovn7q21MDKAJ9mF2HQ9nfobhaaUnMs
46/oCO4cDrPDUL9fbk8ADf5tbLa9p0Me+MyA6fSumxjPTbutzVpCd1ioeN0SaLsBSGr2qklSYSwx
OKPKFhioF+CJMwdjaIDchSl7OoDbmWZV9m2vpFrOBDdLvDXk58FfxCm2iwE+f032mfLs/43hSV0S
k1TVA/ym2wyAMESLKpvtYwCcofbMK3Cch42ltBjz2E1GA6ScthrUhqnTZRIW7yPhGL++77WRl8BW
VVo6J1LkRRP2bB/RiryZCowOgLgph/zp65q3FjO9VcK962+NDDy7CKYjhgGb834hP8+6wYDAPY2P
WYARlP7hblwdd2tMEoOWjvH7eBk6ogPKI1Lyp6rHFfLYyE9PcZDYb7EAdN1CreTZDQ6itXZFdZeO
GKhhSEmdUmCLam3I28xjQEcSiEpwEMpgAY4kod3beDVP2MhhTs4P+HcnnEzLG8sAr/LCUxRfUhlx
pslLipf/yeGc0HQGsNIx4lKjUq4n7xuNt3Zx5FbSS1T0wtT2t/TROOb6DW+Amho0A2+1VVrqy6EE
6bQLrf7g4g+wH44hhqxN96jmn0/3zrD8GQqudWmTbqF/pe2EplgSaaE6HiozZJACXm4z9j8nhoOJ
FsT68FjJMIgG1mGpRlxW1h01t6JjrYbKicItvv05vBr0/MzUTvRRFXGPuFJS0eCwOro9B2JjR9j9
mktAVh0c6TZKO0OJ1R+AQc3Bt65KH14l2Nyvsv11LPqkvnqBcf4YlfN9K5Bic01LFGmcX2HVy7qC
PuDEx8zyWp4msqjwvK/SxJH871OJvzlYStTpQtP+SmcFtrwp8Bc5dUy5ONQGZSUY9DTe/DavA/YR
GaoOTPaWiZ0lr5lZAJwEe4+0JjoE/H0Q1d/vQHDNjPm/AakDMRhhJh/2PSG5Z79P5aBB/EdeaBkT
Y539s/80+b542TafAcaAjS6bnAA3FctBYd2nLUO/S3m1Bgsqj3CBT95rjqhwWYX9v32MT+I4IX/8
C8ZFmjiSUD8F2s+UjYdpC5ijZphKpY16wvWdng9NUAu5xv61Cmq1Ppjrtdca6uGYNencJ/+pCKhq
ld4d/AlLRDRRFIH3O1o/uGsJvZVNfOcj5reUM+S6yfGxjIPUS1BbjQi+Nt8ODci8nMgxZ8HSP5v7
2jaKQXbwjp7RzLY4wYyY3cOol1dMQz4yK7q9c9qy8oeFEIrO4lfXGqT+HrpXzIVhGoj8eeobz3Jg
ZhLb6yB7jX21wduQttbBu+YdTaLtOXJf2qLo05hRGo0/OAWYVNpdIGWARN0c7c9EAUqnEzos48XM
PfxmETRmHceHMWcuhspRtdlYtzX5jKAGUVTkYA9B+cyizCZE0i6q6xum28HKAcKJclLRK0ZRIil1
G7Ief6PSDuw9jD2u3U6785yvsGedLZmHIfZVYj8Ho9Qj+JU/2AkVMldFcWWjrKf0DAt3/EyA1zQL
6ZBImsaKSX7xVtztAkfX4xpmecr8fSczwDPav4NvpfPo4OpE/tXuybhvKjYRydHvW/iT0E3PeFiB
Km2Ua/KdhJdxj+Di+9nd0M1AsclwT7MEcv0IdBq86wSfap3nC8eGrbqmfuk3sY6vB5CTXkd5erzG
X5uXRwTa8qrBK7jsMILZ9K3hu2S2uGx0TabahTCGeNm1HPcCFS8egAHL8EJZiqIs6bhx9lXPWESS
oU/B0h94oMrLqQpQVWHncnPZhDGC+lBh/6u2JIIbK5DfkAtx5h8+g7s/+1z15tfPHo2EcvmCzlZT
7B9JECAIHQneu971qTw4RorvhOMiobkmhxhrQJIDs0QLXjX5cbQwnFXj8Hy+Y6DRG3U3pjI4Jf/f
pQl0csBwx4ThKf4VI946fFgWa/BmduG6Wb9SskkewEdq6t/xlkFlzLenqSZ6K/UCeDx5+QxNKoRT
jnXIrD4Ak1HJ6sOAs+1C3pSa7EtAzFGLYMW4rrsxyt20EsfgBIF21Rsma/jam+gWr3JwvcgHFoJP
gk+sjU3kA3zs9WjSwZE6DK6XK1yNqnL+NEIh5y+GTQ0gm30o17kBckMDvc2UeFBN4pdUg+6Pe2XV
8M9HWr9Z4QdlUQ+fKtA3SU1sg39oY9rj3BePGx9B+H10qTcbfLbUFq+4evlijHoH+9xM7mWD3i1q
//AQq6nt8fEXjhjfzqM//LtnH6Y2shZ9Q3znHFeXCqaoV17U4FnVWAeQnkzE66+vI3tD6B3GAZen
s7y45COuQWzI3RHyYWqyoWDbXKRIFwDRSqvnCNpoxgk677kO1BGkMzCvXEnV3MoepNKMYMHyxZkB
dKZfFNGF4kQX1NchI7VzoWSt7Lt7C8IbWz/kK6TWkOXqFDMrGsv8vkZlsDCoc2Hys8NpCfSZdeGT
4P6/sg/nNqrE5jQc09RigxSWLdHspAfCQIvxhCdvhpedSLc5FgEn92Bub5t1z/uQfsZ7cmGz9yk9
JJqKSoPY5deQJlv3oGPxD78AZYisThTBnmfJSJj1kDaq+XGKdXnx1K0RZu0dP0PcSHIL8BAzT8yz
lQ1TjQZETCNRfZo4k0ZRyMPEsr1xxkquzTLspeFB5d55Zwlc1gjOdHdTc5BeJG6S06znY8d0ck+r
Vc55FvJt4c9wGNFtHJYfqIiZ3egVAfY7JNLdRt8KVGXQpfz5p906VN6WL9yPKP5naxBYQKjyKA+i
EnCNar2S4EOyA4SzvldmvBxvcXaqXxYehJPs+vWk5h7ruvSpP8nKnONQNX2jl0PN+G6auWSTIVNy
BmQHUpWoeLD3u1vqCJN9GgJBEpsTs/mlnQAWRgJn0rbX08/WqtkoPdLzmjmPrQSL/paB+N7Eq+z0
zFqztK7zYC/I2KDo4IRPLrhNpba+n6PT6azzP6Kxp5cSDNhiyd4jgfVVbFG9Sw32CaLtalyUGJ7t
8D2sw9xaQXPXzbp0T/Sf5ahRQJG6qOxLB+alm3vZu8n0YcGqcx2eZyO7bkMjgyZ/juUDiI29rw6G
7OqxQS39jIY2FWZPnQ5V4leh489jmjW5KpXUAxU5QPl5cq7X+aXep004DSI1k3yxFdEfmvP03TDJ
KqP5wzm1nmLrnsLl3Ge2Mm+YRW/I6nvZKoOU7Vgr4W7JJSa11vM/PzG3m8nESKY4JmbX+hQ/Fbqj
n6exQQOJJPC/kOxWL99oB7JEad+GVS86M4IN+A+K0pJoCzM3EJi3Av/qsVBl47c9YYs2g6fNwUtW
cuf0H9a9zNnoGEaLFsmekHDZUt5vUomTL2ZHd1VZlY9wkN5aaXAi0vJ884949QcpFC66DcAhJ0Y/
kb91xjwhOPNKMepaUF2K+2f+zwgHURE/EN4zzVoH0NWSqBt9KMr7V0fZx3bS6xS4anqUygxD2wye
o1OcC8sMoGU/qb1WiZhIPki036h+s4s4fk32gWvL7RPgEj3AcRshoIU7IDk8NVSIUt2B7yGgAOos
Cip6HoCMiRh77N0vHh1C4hDKpqnLY/sxJnJ0L4zl31MX96rFtx+M8UXtLt0BoCJdo+bmx1RwinbM
0hF0VFc+mCoI+45qm99YELTKkLTWJYxdIUc+o7QzMvjIrqc+5PjEXoSFHsGN9YKHnC2yzcQyb+5t
818LLOdkSF98nOgwf4krcow+Ys5FtZurM4tI8vOqgqtsTKCe3xTi2wMCCnLYK2qTMnbTdZvFbuz8
9TjeXhAT6MVnpONOUqfTLF41nTLoHTjnIog03k9ql9hxpKKUDMnqzc3PWlaBx8flTXzMUKZibQPQ
TrMIQfcnLzeQTKoYVpqLKLFpaWT9oMU1fTQh9hkcdz0PtdWo0pH4NT+rdpv8f22ygalTXrW60hWB
Yc7wTe+PGDATA8/eEpkTeDx64NRc52FdTr+XZsHwz7x4Dg/qGMd7K28z0+fER3zfD8otj9jpBGIe
v6zFLlxax97S3sV76oJbrjH+vsQnn/eqquaDHklWMslO3NeX2ncfIZiDTU+NpnOx3GVIvWe0k9HP
X2LZH+iD1sCxC/HYAuiikBv2O3g2NFkluQJPj5vWNVUetnJVHtr2s43PzoYc4qPF8sRbKssLU4nW
fNufm8AatkC0i6aIvIAH0PMVUX2ypKINIe2zMBCplu7q0TqOvt0hVgsb6kzVMLlLNPYxecQepXpf
P4iASUKvK48pjmDIO5mYeT57NEO+h93TI12l6lyWTSWSwlEbu+3R7Sf/X/aI+rlaN9Tqb8TDIXH/
S8UjHCLEZQiE9dD8BNDqMC7wl6aCKxwBKBSgUXYt9D1Jccv9f1uix+CP8N9BTMrZ4jis7PqCQx6R
L3dZ/wQqivHR0ixE5C7MMqkdIh6m0IjQOELtduB4u+KOOZgQIVxLA36P8aWWjM+8/j+y/AFZDScq
SZhGs2DzbbsgkboAxF7MeSqbbslm+ShU7izVLU99llyhL8xJWf6mFB1NqluUaXXYNRQqKA26u9UJ
DHZG1xnV19jTEtjA26NdWWQdjYZWe9c95FCgvcbxF46Fnd8/bnXKm7GCCDSJiJVM8ABvEyak+918
Lf8x5DJEPwL8rV53bWFYrMueyLRCmFyaF3OGXVctri8wgZ2EYA90eav7MhlG4x6GW3eTCk+6jFqz
RziTK6slSplJGyXxhBktOPAnj7r9GWSbbB/IDTEc+oRE/KdtSWPuxFXs3QLg/1+zYqbEeXnzwiYp
69UAEBFilY9EBM0nJa6S1qGpqv2NOxTIeu3YjpePFA0vrLOTGe0FExAZQ0HzVLrY41k5QdF2hHEQ
3VmMjC+eu3ZZh47Kl9pk9Ypvo6Zu5uQZMODINS7UZmvbvOVfonfIaoSGqKDCWEK+r9edDGTaPydg
iWczehj0B5sEnRnh+ybfFwL01gCnrelOhmfNv/Ws8TZw9V3JAdhlc0ySmW15kRzu3IXoqKGwWcdE
8b3cG8hq+WrX0yOeCs4QbtUq5kiGJtBAk2RaMr2hR3gEasqwsrNazFOO8UIEo9nUkQysJls83UFg
RRAT9cYdexHIGip3jxE+hLH/HLYuExkYEyOYuEAswDFMuZRDm8PpsMhokL5pQ76LTXkUE2LmwMeO
cc6CPP71Q7HdfllP1nkp7Bgl2Q79hrphvqvIv11h249Ui01kmMxvDmrdtAGY4BbLwQoo0e2yh3DT
f+QuBuUMd2uCLMj0eV0WhbTbUD9iSnH4A94rXDRvLt0x8A5q9h5hNEv9FbCXijiZGEyqWuXEJVn+
hrJo+ZNNL7UH7WABKHhyN82s6+tgeMeeuNuE/QijZa67euKOesUqlJGthgpgW9sXIBro7zemteKG
KAySNF4cHBc3Gt35rJk2j8EY829RDFYWrRgnK4jqo2SpwkG0tXECJ54ZTX4U5INVeP05j8cjdfE6
Mq68OwtXmvEjTRUtBK7Zxt16ZF7kc5IlNI+rYrtdvPLHVSrebi35W5mCCB4RGZWvJKe0Xx1ch2ip
0wNLvLUErzBq++oODdPW7Wr3knUZSB1t/GRugM/km0sr8Ule0SQGf82Qq4VrDgQAEam0tjYzL5zm
BU38b99FSemE4VXmInWdh0Bd14bjA5F9QgOXi1JtoVXcR48TBeWJp9P/UXM9QDtLN+aC/RNNKEHN
E8MN8ZVH1VkV/5tQhWFnfYzC4JFrz0btsT1I2l0W/r0dAsJ0XbTfEodV1fzNRrfCqT+4BeclVk6F
WEQOhNAxwZoD/HwdHHmGctUa0kAY9RKSOPNtCPpLPblZsfnHiX7rxk0yjmfd05K3BwsNZi2fVxGo
+2cBNMRCUFNL1HhLWLUct6jC1lU77a8QH6HwqNXLZ31wvttvLg+mWRLKvGgpkNxiTYnPZEFf5A1J
9nX/0c4YjbBKkI0m8276dkrI+oNbK4dR3ieBMh8tQtGfVl8zFDJI0M7vYEf5KKhhvDBkQ61PWU6Q
r0cbO1uQr8g92fzdoQZNj5xThXLe8Pc5L44NC6TtwVI4EKwZCmcndE8YFi6i7GN9KYEzrY/1SFDy
OzVpbF4blnApy++qznQTTifcwgRa6ioVe5Iy3QXenvzFy/aSJ2TMBGQiHjDrEfRi7+0EGm8l+ygi
tr/3h8/pJ8W4qTGqrmbyZtxJR6WzjxsNaYu1fMDtXxFu29IPg9uw6aPgn6nomQD29nhVtO8F0vN2
BRmfQ57fAMfJHgFooZeSB4l8ChOs3xwPtXxk2Ls3ecvaXhf5RIGRIRhp2WXg213vKYS/79c+jc1n
87w1wKHbuvRl/t8Cu5Bf8206Sye5+tqmqe0d1QjPRAgd+hm7eeJlSeaLoyugUa6evjKv7iem53VR
u1wubB6kaLz2gfF1uOsijExH/0jpufk1LbD2qeat6MZEwbRzlisFsNBYDhexH5bHkAKhY7y779hl
5S4kFyhTtnsJXDQFdNTcPeGs9+NJ1PHwVdyHhb90jKae+BaTYqxAgOPbScpRGXENJrhguXOILbrL
INcJGZQ36DURXS6ynQQ6hs/9MqeFU50BcOhdHThlggXt23nt13ieFbgsHEl/CTGYOfqva83kjaDV
iQPvrtA6LVUH06wdEfxV1xuSzTsIn7Zm9ihkMxYZR0ekaUtb99i8ibFF8bPmnqJ3lOXrlS5hqYwx
MpF8i6L20gQeYdPRUn6evmqf4fnaJJoSJLXtSbOoIvAcWAGl1ePoZ5xUZvkAenNtoZooHYKPJ3fe
x/7lJ293kaJrpTZbJwBOjbS8iU8ucqY0rlxmm5ubCWv3DvBojAiYwwuhhZddwZc7kzdeJ6MVqUrQ
UQNHwJH/8a9N4u9MU3CvoLLRswpNpcMIrqr3ccG19v8woB5Qry/FN2lH4BKLv7PhvHYkXCKSBGOs
0YA089J4+owjCKO+0YpHZw5nnek1mdOmr1MxMqhvUSASJtnQVak276tvY815wftvseHZfH1OKmrv
Ja8RqkxPRCvBtqB3nR5j9PdyxEflLlk4aJP0IyNqH/IIQNhZu8QcZvFg+2LiyDqGd3jgo5TXM9bt
xWgOUY7sOWpNC7zBEPPxRbbFaR5si9EEGBnjw44o1bXFXQ9rmhvjKgzBcBIHy+xl5l6tT0HNY4QJ
CUanWCpZke/5DXx+p3gPUbC4T4sj2lQL1ZJqWp/AQnHpV1Ek1KTewGeavy/K+evFGkKiK69PoxuV
sC2ghtOKWhvklGW72MfLmkZqoo7nbqnZfl7FOERlUQFZnh7HuBFfayM7WdiN5MGFs0F2oOXZFW3g
e00MKmagF5dwqeld5duB7gyuj0yCX4rWol+r1TJD1KBgNbIlhxpjnaRVorGQmuAod9+oHNQM6RA9
++qivQxnl80gCA7vYb73TSfJphQFMeo6AH63rOXmsi+KvRtS2rhvl+0jNWb8pSLlciI/0Aq4BPo1
C0IzIsyLhjy6cnpwXcnHR0A1AK3iaKDQH88C3eEUPV4e+lkknPwIl94IGiI+sZDG1Ff/Cl5wxp/6
s2hynZJ+SkvScfj4+IP4/+rEZUGt9pBloPTChWIeosOeoQA0rBzLyNnYiQiiKV9FF3K8siFhyCqw
FnZABbNZpRc1atZB7NZNxg2sCdeKDShN2udNzJJDSx2TGilKbUuRVuv3m7xXgLmDCawP+2HqaHAE
f7f1wUDdPqxU8KgyJxKswqY13rVTkx5QDVrXFD4PXWUBg2e1j0WevWaNCgSqfCQ/SFhp4AjTUc5y
UhTUJ4rWdDV575gtXECGCvsYbf9sdhaCFxDqYL5kkM33nVzfhIbfmwwxwYy9t3wkxt0tFQVgSRCO
fOD5S+9m3m3GbmNXOrK1dQBptznDmVHEhDmcP4oOYqk8+wp4QcncQWLCO8fEAmp9OQ1Yin1ye9wb
7WofTL3DbDJNqVoXAbzeRUODGpzvtGmV4d6O12xoam6G7VAMgKXbVMU/hBQp8v6e/l4mlXxk1Y3j
3/Fp8t5TnbfSYfWe5+bDgIB9ImMdcoaMxt8kqShnJKR6z6fUeh2whPLV/aBGGl9K4DMl4MT4aM+7
+bcXzVNAh5P7PZiTORGF8nDimE7aFjreQAtyXAm9jiFn7kvXpy2BkRx6GezQAkW+YSc/HHbd3dlB
HES7DuouTITn024NEGyuzJ1rJp3meMH17NfiX0F0JZ5XfPOZdTGKKQYRo7Q44teg7/q0X2i/uM5u
fYnuqOXd7pnJb8A/kWkALrPRKT0EBFidpwBf+SqNqx5j5pukT9zXbvM2IeaVmUnliOq4HRsyyNKE
AaqKrntk6a+3ds7XsRvJOolrnwOt790hzNuca1WNOEd2e8UbRjq7CiasikZx00TsK4cVM5baXone
YccLLJKufcrSuKGzuHjvZN8Z4/X7cajO8RR/TTKTjxxyRMnmvqVNL3qTFGgVrPSNwk/nrbKwNYrW
+IBeOK1M8mD/vOxzYqLlD6f7Xj14H4CMQmIcSG1ZYse07HH80uMjXL4Q8H4jowHuAWMKvnu/OxUP
fOBS0zsofZPkDaV4f5587upMx7qxyZMHcYeLiJe9qVYMYPp/ZEO0ttOB4uFA/dL9XN840fNE+wF7
liL8Zyj5GGExATN6R41JWKW318JAfnFYzMcfpbVdR3DmlJzT/qqdvytK+dSHGh0mp9jrQ71lSEKC
VZhVdMwe5G8ajf9MAlbp4dltZ5bavfpYinSaxZGgAXIm/u1ODy6a6N4txm/B1JuPDKpo9nw17ryg
0Jl3AgAOii7STxAGYWeipPGuFLWN25dmzGgDjCIfIIZ3D9z4p74FH5OmIdU/k+OyowrXFaoqEVAY
qqg8U7MPMfcNOKO0LkIaq3xM7y6ORgmdE5tObSYzluAWLlp8AF9CMK16OZKDOR4iD2YHH3ecL3S5
nDmnZmxqStngVMlyCu5U+eqFSacP4NyXCqI3tfL3lODSo8yj+djXi6O6qyBIKaBZbg5yXRduYaQS
mgrqxfirHqpreg2CZgqqUEgecSv06YsMAfRWy8w1l5qjA9QMY1sfl9HKpa/s2yYXT+6WVBxIxuQV
nbWzqGMeuK+M39OvmG9yoyOmk+DJguiFVjdyWY/cWfDKLwYvCrangO5K990ZXALqVsuf3BoILCMH
aQe9N/V0dLsGNnEgv8pxyZ2GuB5h5qTh9Y580ZyyJ4F3cOsUXD5Zt7BptAFkQsNsH6RPiqAtFMsy
gcKzZsyxG8n879StV/gNprb3vmGCYlJXKGHOceiVvl5LolP1WWwTNhW0ZS9nSVLebwCuLmo/w79h
4Izr3itYTLx2/noH5JaFsn9khNeSMEFig135rUhL5ClS3Sa3O2sPUd0spEW/c13VReOcKkBoYRjd
+gOebqOfLUEHMLt0xl8F6KrpgWJvf5p3EN5jKu5jfk7q2OYNAt8U5kxKdlxD3MoHuLwXMbekQ0Lx
bxqrm6Rq5Bj4rlqk7EnDXBBGcwwtl4TjLYtUmpV5IBh+yIwgwKv4pU0yo9BzKI5HS6/VzjGqD5qF
f3ga6Z0X0x/HVQYRtC+TC3kcfig+jfYhDBLRJUEQZThp7iu8s63nM5so977ZQYiDcXIbPSUgU90s
4CQZhSRpJyoxCND0HSKFxD+ZiHKBTXj0afrPCGvjSO+UiivgOcueJJCHKHlf4iiQKHjiGFipyVej
/5Fvdpgp2XuF3n5fGraHwYxmsfu0gtDlkEokDsAENOooVJuuyw/a8DGXmngiAAJNM92kp4AnjMPT
hr0m/p0XVNmnS3vWyIkT+tddkWLsTNGBiXBV2M0H+zwh5Xpl1BWAZO84qfA8uSg2qSCdfwziC2x4
6VoukXvpNg7tqgLMzesqiQl8KNEN2HLYZJeE7g8WU5j60dsDEzgUczOgUB4G/mQ6cvMTKNCNlEbi
2KMkOfdSVTs6Qd34G5CypMUb7Vt+oh/I4J5lo07G1/khZQllc50XE1CYBc2lhLe7lRedTNJYqNlx
EmY2vmeEKj9y9U47t8oA9kV29IJqbzz/e7lRWgsoGfGuX6rkADRBQgtP22JkL95I4lWANwN2PKWA
5W6DWhn2kRHUUCEZ/cYzgEiSrPipEIzptTgEkjQgzVMJq0Bf8qDLd89Te8TueWtHWrTMeeWVFQec
oKnp+SnU/OxObx7zfRaEax7/GSScFJ2POQhlbovldML0To5E8973+kQavxKLMTxwKBxunUv5wiIt
6zTqIs17vBZwf0ri3sySmUOzc8dJgohfv1+ggTNFK01VimZeyju0Ytx+pFbRkiceg2S7SkvM+oMI
e+IRvpnrabYRCkWuAG5X0W/Ii1p/A3XcEeQ4g1qUzYQ+4uImHpPl+fK/yNNCHBKNcBF8HzwdV2uD
vLl9qp9kXcC0hheEEqxw7fnwzdPnYgo3lNqLfb9YnhNHL0PsO4vblsfjWx0/IS9O8hh1YlL9KIvI
UrHD9SJuh/9ZOFelUHQgr/ZcRDQf9vgWBfjOnTq2q2U0YLIBHZz5DsLSbrzkWthK+fSzIXNNpbhk
DvTX2dglr8CV5zXmjjKl6HWFshxyhW/JpGo8h/yzcqLELWxj31qV87FDMam0RyX93JGyQyIouXE/
DjsN962PeCjtVlMao8c/gwwKISoXQqE/B9IjFid6R/YSYvTqf7q09+t7te9pgOs53+67opSMAPTb
8eqpULShodiJHzwwcALsmhTKOhYFpgWe4K+4qZUDnb+dPkmnJBwI8gULPneyMA1RlHBzE1O8piiG
wW5Li0LKQHcGFC5NdSFtsS9xZeXNkDB18XaXqAoPaPP87o70JmpAExss0X9YkKKhVQkeGJ4PgTgA
UFLgUAumPAhM+d3Z5SVtT+FlhQ4BxUWYyRJJdoYvOvfeJGf7y2mTLGz3f40ErNjsPfTUicMdd4jH
jIyIFrSa1e5nzDOBXOrVhTpz3zN6wCjnQVB61/PTRA0b73xt1VSPbMjz2D0T0Rw2oVMiEo9GrKud
1VxtgWLA3wJVfd8X3bTkCSeADPedbR5Ss9tITwAi2aem6TIwL0qfPt4qx2Mf5j31IGS2oJs/5hHH
pln40usNtT42+JN3QVdON6YcOpVByFXE2G0jmB1vyeNqtH+1aoQYK6JxrLNyFTdIeuXZF9zmjWSn
P6tzRegPljsqeQo0qDHWgXCL2XH8l9910/j2otfvCeQNMF4lDXib1Yod7STu9MLsmCMEzDCUj6Cb
U2HSjspxhpUCXX+pKRlgPJPbbTztrS4VwZ2RATTUkdn85A8sGN7J8SfbA0skbF+ieAYzA4PdnFd9
YkD1ps2w5vcjAQWPY/JH873ZIzj0H+f6y+vbVW1tOdzsmDtu7aSQBJis7jYXSAelry9zsIuWGw06
QOirIuVaq0PQVLNGwdHJ4C8Dp+PUx4oni45m9wFVyzMLUbuEMnOOKVSb6rVuIcOnSvWhkDG7x3kn
0MieY5Y2yh2aRSeaj6KtIZovZtYxXtB6ZpK4POnmldmZ9/CJSDwz+ZD2LASEHXy++uPhkWdtxhcw
ZmodSHhF1GLqnvURoBbHEfyYhqZwFgnKPbIi0VAV1zYr/cPMmKSrd2dw6JbqAQygsiAka06qSUCN
/5s4m2Dk55Ok19aCAITw6FOoCTIccY9Px9F6fqrH22z9OTy7jInMWR6noq/eWuLsxrFq+KYma5+h
BazYw4W6JXQYrZJwFtS/9OeB50t3SOIkFmWr+Ev2WItOpKPzCAwrITOssd6XH7n1AoelKlCeGfmZ
nd+4fc3l/+JMC9ZMOxq5/LOIasrWcxIi2bznT6eKh3Lr0qsJ1u8ZhMHZs52F46lmeWjD1Q4fTKxg
3aIU6E2lbM1oePujIrb44L8hl0m10t1rraI2r1Wg1Nq0k9JhGx7eG2xyBGYBlGlZv8v9pjRd/l8a
OND4jjPrT0ES4DGqN0MVq9fYSP+kVXbbXmId1Tqwe+stc6YV1xjbwCJPYRfdLe0swaPvnMM+VzLe
1lgPFKI2Fx713yfF+7dHOWhOX28slZrBJWh2xzKzjs9EX/q/CYje8VHoXXqullXlfj2RtytZL5j1
QTzz6RubMCTH98LgYXUA/Gqy/uv6StQztHr3WY5l9NaYdMMtMA2e1kkNN2MMsZWY7S9w7PBfZjkA
Rg6St2G/sd7XPSFTk8eAAEcf8/DggJ/bWx41b/FB5cfL7olHrpKZxbbqTwX23+krV+G69I73/ikO
Soa4q237lFy53QNyFYeYdARyZOj0Ia2ej/cTsqWp6bY9VDJtAYmWwbn3Lf5zkeno+3VeRhF3JysI
bdv2PJjeAW6/sOZjobWURsHxB2oTho+36mjGF8Qg2WQieTyba+qMf/pYz9HE2OAPvoELBW0QxIXy
to+k0LInc4DoG0tHQniWEhsK3NGeivMiukSqqZ3uutYnoPXiDZ9an1aLmUyqTDaNXSkSc1wGCsUq
SaLRqR4OSQ+XUBkW93EV2SumbSSF5FxSkLCORLUFCQgHrUo1NIfXwGU0wOIgqCdFv2stfeMqwxC/
aW5wbdW00qDxMJdYgEuXRqoNPSdRkyh30vDl/SnVd+Z9Meu1ryykBsJEaBLnwwHqu1yUfudu4Sw7
Z4YmUsJYjHpxIzXmDMuU2WDsIAcLs0y32N9AI/4DYKapEoz7qa203xIzXWSlBrI0Mxuz7Wxtp91I
8IQ/jXyLvDcKAuqzM7mXCrzW+eXqAOiB1VteMMkk9c0mIz9VOdkps7i+JNabs0jUyzK8KE/XLwSP
xAP2q8p8GWKkvmlrNWtyejmv5+eJkgI/WTLt+gbfaQ8azoJBFo4fwvPw9dasN1soMxlxXPZFtJqI
vY0AzWnpeA5l/SCt6YZVKuLdAdI8mtybS/nJ4agco3vnqdff/ZVqf0nCfUbf+FAU6KmdM7qvbu0I
QpMuT/plMWmXKbqmBtuSrckgNdCZk5PeklK9VFaZy4cJut6MuJ6d45oZP9eOduyCLXgvat8V1UAX
IPw3QvXP7J43JWR6/pr2siKM7yd+3U2JX7V9UYh16pc9FWIM7xIpsQtQnFK2Dm3+2HSHan84blv1
NWLpqeVTKOyi1UqAPstnluW1uH2fojG5/Rj0x4GE536o8a50uG3UsE0GxIn3iwQtGjU93aBAzniU
ElO52JT3QYTS1HL0gELvhcAd4EXsj/8P67FbIrxOEVGUqfC/f9INEYl8oG2YlsNy28zf9n7+DA8c
N/yDCgWOBvA4b/af0owC0Lqo98y6Y+AVvQd+DKNqzyNEz/OzB+BvZQEIPoy+1VUYvHFjngnYCtNM
mD3wQN7juht+WYsCYhVhpYdQTTLgp6W4fte1336BctSTpEI3BasiChVdPbguX46Q6pegNMNlHIjK
AHv4X+p9OilkFw5TdmWXOhkdYRjmAmJLVJPxTYpmnjWS8iJgN8O5AmEJu09mEScoc1LO2CfC22T0
JFlOaaW7Kd7/FNUdHaM/Szmzr6u+FEcxblbXsJmOt7BCY4VLg+2tCeAShxMOvdbH0050ibkBhx1j
tBZ3c4Q+cpqR4i8+/arn7BGXnhE3CTOR1ucSs/zSZ8Hy5nDm/PUDCb5j4IcIMyHJY95hQHhThT5O
I7wIC5N6EX4ckZzyPwBLGYhYx+Dz3W55IJEhEyATWx1Y4gLJVqVOossCZd7KCLyrvMVx966Df5jx
oDYoaSKj37nGWMUpCTES0qNu0ndyhtDM1VbNa+398oW/vVL/K4sNLczaBv4nZ9HqD88ZLOp5/XGj
F2OGmJ6SSiI+QSjvzrQsc8TNAX9sUNRxEw6fv8USmQyDf4o8t+PhxzoO0KU7DKty1RkEyv4t/Y7U
zq4rTnOy4nTl0GieaOgtAtSGNYOWL+nLXay3MUm1CI43nwIJtWaiaf/QPDABhkZWCW86gm7fx5a6
ZWVnBwOtoEP8fIWIr+vgcuBc4muDC9pwe3WiJUtNd5Co6H7+RHuUJRZ0dcdkF5pUpKN0HHdBRmgH
z7e1eM8ze1UgTjR0IEUOBqwINV0nUzn6g2N77ugzw3ANWMQEo9qzKQ4JNZif6xHZBau2WIRAMF4r
0cLLLAbi8ernIsXCqyny2o3QzBFyqG1XGnv+j1z3SZGQLTH7DFuz0sv3EBj1hOxfYZTLQ7ANj5P7
2YqHxJ9gQdDh7M/UG25yoa/vvSxrCkrKAHWEib+z8FbGZcBTKbigkoQps1pU37dA4EMTo0KsDqG9
cEVJ4Rpz9BZxLz49tJQ/gntGx4gv2XlSASiFb3Jyg3WwMlXtnIirV+ZMGzP8Zuza1MJhqibu7E14
UtsRX1NVpoHVJiTsK3NqVss21FHOoQC6mWokaMOPSG5S+OcA7yLLXWqQhOc4DF++W8Hp3itn0Ipu
aTm3HNq+hAFVKJK509GHAzjVs3WDwKfEILxsfDXoNYtnMpz0NXxl9iMMUIa1/oDIxrQcqfJYQRD2
N9xUBfRsTNWmCvJ4PhbOQVno+E8aQ3BIsKXLbpEJUV3o9rnlNpv/fW4PCUWTBJVH+0QdKgI50PBV
a62vetqHgtVLEz5qhWf6K4+1wf8Kx1ktXJfYMuUrU4ifNPpoPjC/UX/LW+SIQlhA8A9aaO1jps/d
0Tohy4O7uVFAVDqZ7dhB/XQHKhRQxUauVFKolAZJqCpIPIjGSWdwOQNRVYVYOt4Wdc6COHhXegkI
E9IFMe/GjoG58+1pfABISNjFSUb1Y8OPs3HahqnTdlmh9Rv87DDN1zVG29oTKA4R49kw7lgotv/D
HMlpWpYdDPkY9TOmgf07zA6bck0dVSfG7VetHOuIdIh/j/f7axYkzDWQ4dgE3zBzZBpb+WMYTzyg
tubSlGYn5RC+nkT/B4XMnYv5TAyXwfw91xq06jkCHTcZIoz7zl+bUarwOk5XULZAylUFsGeJQhzY
mFm6fDMC7u/bfqol/TRYxnCrFVCiCZ+NK89sO+H1tU76bpCHz09vRK9vvUW3Soft0Lha/dnlcMpV
25B6KEE+7ZR4EYMfWsDgpBlbyxOfgE0UXBk6//s0GP4Ef6VUzkUc5D5qWsBnPapmr2ielWuDaQRS
R70EmuQI1AEJFUxnkOLmYcRb1nqK7BsDzM2tludxcpGoxFdZebKa/K5soWz1WyDwEqbckluV8ErA
0t6aTlBQJQHUdk+JxVZo47u6b1MhkNSFb8GfKqi3dZ9J/tj+zZNn+7WMS3elue8qWKamKX+8F72z
Su2QZl9pgVaNdUiOia1Apu3VotCpe1s1KKedpHG3xNGF/8YeMrh506rL8EbYZUElhWVpQGo5iXH/
H2ozyBE4EJ1iFrYFwcHO7GTg4feyssJAYx69zPkLXU68FubWc/2K8QR++Nd7O/XxJFHkcC1amG7f
JmHj7xmuIvFbYulie88V4BNm2KgiAIwgce4hhZUla0qTbLr31kvlRAWu2GJSctYmAOZd+9jSAN2p
Yp2kyfhtAuSvQFNryBuTti792oIuJoJ/AGCkPZv786N7eVLAFaSnpncrrcoeaD50d68KOL6I3Z95
9PW/YJz2G6veap7J7bhgLGLtYdo53mDz8P9TBFU1fjsKd2a0M/Tll/8OyXRGMJaGuJaqyDaUBIHY
x0s6cGgyRbnCAk4BFzaXcR95VdByVcj/lYMEqqGKMBv6PFSQNlcSWQelSs83CD43g/WsLGgZQ8Sb
QZbmsNz8rr66YV0D9nAnlROX5CSge6o7ZNuhyrOn00qu1cs3OUSaQhFcsiLbD3EuuGmqnhBWAzCs
Nci0JUoY+5CAh5wEc/F6QCIjRWfq6Zd+1xsBE2DIHVDuF8CDtowalvSRZLLuyQAixwtBsEjXDKf9
zOXfEnf2UGlbuHywhhRQCAPaWvqCfBG2oHa2kw3aHw6j+sETDI68aCXCVQTO/34augjZZlkmf/p+
v0KusztIVl95POtJuSScsDz+x+bWOpIAKisIucTVbVyqJVC3glVMVYAsXjS9t+DGS0BCzc1Ov0bP
h6k9tluxQ5KR6pvuODxu3f/9kUA20SSH4fXt29Y4JGAkujfUu5XOE+PRfkAKKfcFgtC5BWLoZeym
vwWqyKZOfnjmSpP88BPSXI6ij38zRLa8JogUsLKtaWHC7gDrfBAZiOSEADQJUw46+UqDSZnOmFO4
wj+ffGTZF6JpaK55a26knMfKZ0uxTzpxVmd/0zucsWGRdKzy1Q9oe4vNfBfJCSAZPpELI220A2Rb
UGIfQcgrlgGlUm8Lu/Dvfj3d9h+1b/V8rCDIYLEUs2kj68xKt1e94lZBU9h7vNT58fHgWLjchpLi
Et1wocpK+0EyjOJQboo9WeufYxRc/XQdGL7NPyK3DEjMjrp45XJDplZdMPFxbPaV31qXixRtxPjR
HOyYzonDGfbgo2E8Zgc2BcVtg4at1pqIVwOCU0I1R2E9O0uuOtfwv2Y6oZGiJynNNT1PB+EDFrQl
L9UwpQ1ODL0+OLDguAd46CIqyIV4HXSmAqTkNQ/Q7lMbxwyOkiLjiDgUhskK3ZPUcblvCHjTwBQa
qkA0t0+WgaZcVJWnZU8UZJWexfX26GMMY4bwZhh7fhrmCKO/8ue8Z8G1KyBtiNAWF5o3fLtFUvXQ
G+ZD6Vk6bRT7aApcehym776T8wptTsgwcFBnwOWJ6HQCcota+QQtJ8Ii9O4naMsuC5wCDauT6bIY
+bdArs1x14DlTxzQ8EAO3PNkrdnDCKMQl7f9uUsV8MUCcJKAKWjhaoN764ZNV1eFYBgf7CXS1VNK
enG58ngj1WzwJNCGPDDHzYTiZJacNVMieGhj6ofYHGmRCcNYGXDECavHWtKNve8e6p5CIFtKILl8
Ra8PfEyBfsBlylGl38jLza0X1AlX8H+OIQsUgre+puMG8hDj9a5U1ZE6XBOdDvbs1Gz+371pMBQG
s7jMRhYZDlqLy29q9iUh5rXyJAetqRWuMrBg1zZqUo8kAi7OYeBzhA8W4VGaoQidpLXY3OmrpFP5
+NcuuGQfD0ANiA1Ow8Hf1huoe3kf65sbroevvCDW7+mfNoltd9+oECE61efPgZi1DMGcj6wZoA/j
Q8n2JN0hE0WsZkSkXzKA16su24PQIZOJ+Kw1BOtznPAMawh+OIKQKL5d1nh+BNrZccRSzYKvrOoi
yFDqTNstCCUqg1U+MP39INv4X29bmLF5EcrgasyQWEUCgQOe050fn7baJIYI5oTUJ71R9IswNhV0
lBnoKckrd1lIZKSI8XrA8MSUu9STaIYPdEJDQfKGwJN4zb+FF7BIyJ+x6QSJQfy2GaTHm1bPHudE
mBnNQK1iKnORaZXn+jnvEDFJS39QYeL4jXINH9aUkwWk9/Wwut96TJ0K6BxW6okLQISGWP0QYHdV
leCIVjRMiPKawb1Z1ovw7ZJk2olJryskZwQ17fNu+sVwLAtsIwcdwnQgMvgd8N0nISe0KF7UU6+p
e9BOBUklEahOKNgWu5PbYfe/253GEtx0wtSdm8XKoi57Db+jNWiMrMSQb5SvKocxKmycjPhQOwK2
SkhbV1Vwo/8h8nAUWIatyzEh1ujnZ2rMTCWiff4M2lThYhImS9Sah4i8tXXyN+8TRmUXU6l9kB0D
3FIwb3mAdSTn+nvw4sRr2iTXMsWc2xseAPRhccT0RRjZzFgIUWdcd4SNYlxVanqgLoO5DyLlQkmO
MU3mCWVChPUh4l1VELqe1khIk8//vDlMmvBOu6QE0oAzcP3P4QTurt6KKq9lbNveVmevKSAOdLO9
r3hssegXhTkoG6cjwk437gi2tRRm8OoH1keekqbNorx/FnQz9UxX2Og4pZkbgkmQ69lIHPxaJks6
7FNUZCndXmXeGNLhDd9ldH0qBwLAlugjSRb/i9MBOCw6b66ybu8lDnDT0T0NEYHsys+Y7hQ5qSVo
FxS8EpIZ+cvguhR6FnrosjcoFBrWOPwLTemYAibAt3XY+Po0rRnAzhbM0gG6tqoTEMqlNPpgUbX4
W2/mWdWU42cEsU0OjB+pf4dUPLaCKOVDMNzBHYvjHuOazG7SsIB4w929iYD47SbeP3Z3YzMZBWKU
0H9pFyFIae3zgSJrJY4+GF8HBX2H6eoS4GULAoPK0mUlu7GsEs6BXBVxKaEcnPzipElmnCTS4pOr
XCqO3buufO6q0Mw/Z1Er3GrC+/3u5ZKNremNdwzD9jXACwnKO/1sGKa9c82dnK9T8ebsZd1bIt0R
XOtUrXi3gP6jI+Y3Vifn1OmYxq4opOp6WOjVOP8iDEbf1aPxwhZnk8I8hwzfoFCR7zHuaskN7CbF
E+PfZxAt1rIUr97bofUR6Qr6ru78vluKiY+8VgxhGrEo1JcSZjBvSs6QI62MffLGBpasC9r2KX0S
rCwgaxBS59wGC5DDVikLeMhLPZkMey10GDll8qGx/ShlbLYWl7I/GSzPjoOl+A/KmCdOWoO8ZgwR
wEzt6duMrr8kCPIdI4Z4tgud668Ll8CTvFZ/e22/6y+qRncb1gZbZ279Xk2T02eChs4JK9rMiniS
dQYl/wlDtKJvGbrdNTPc/2TNDZ0PaBHwX6b1Xr7F9t5ctYOAgGbOkcXVrMvuweMiRDqel6p2/RqF
KxZVkPLJue6GI3WGgxHbqWMK86rF05n0aSXzP5fA+vyUGN9o68BvSAJ3XW8X1RaRmsiTa8BFFxwM
MMr2ZNkf75gUjVXS4PB5WAK9xnVujgaUhg8ybpPD2Q6N6E27Bl22ISfspbO6A7AzeJ42vUsFcc0g
eYNa4p7aBjjkRXi4I1l0Xbb8VILtIZg8akjapqmZV6OnOTcCvw7dsp0I8ZYXppyR2BnvLse3krXW
0o7Q2hNJSucY6zKkmXH682P/HO9z4lhE+zWWkaIKYyVHki3FKRlPlEKc77bKjAvbASMO4ktiG3k+
vCAMeBpPpZMTJaTQJiK40UpuSOvUPzS63LCXcUi7Mmdo++sfLcjw4xbhCk4APIyKXtTYiltF4Tm2
lI2fBqy4F+N+20JuDBP5B4KBiuN8NolwRoi69xKhMBc2y16OMRI+oqESZ49lLA8JtluC6s/7sBQA
DctbD/aQ2CyOL4tu6MebUDfXuIIwh7zqrjEw5f5qWOcYe8qOJOAd1SmpBzbxT2LtDexHcHXrV1M8
IYzE69IzqyCFA8Jf55jqpoNuc4RTka3TKVNxXk5fjGdR8Xgx2XWQsZ5Jmbrzx0/pImx6E9Ng6d36
czUsJT8rAQ8/1LXid2vESZxaPcNW6OaqXFuX6iQvkgxUem3JJd+totPjm6AiLaNC0Wq5GnhoxOop
zadE/LK0UlPrae0zMTyFz2kOZel8xtluK1LpgD7jP5d+NPjCr/AvZwQ6HM+AwgTxfL8e1yBhzURg
uEJA/cxpCHn7uD0/IBRxK/g7o9oXvhJjRFVXcGBMKEJkNT0BO+8+p8LKui6ULxS/ht6NaIgRq57Z
f0VzUG4asr3OF56jGMkbt7WDODUZFNApegzKyvN9S0nqJyKqRhQ2gRejTK5eBkd/pUiUTv5F1OLj
wQfFR+mrNygR490ZrNCdtU//1B2p/NRWTDROETVd9zqm4/1DOtJiaGPuySI8Yg4Z9KidHNp7a51i
AwEvbto4kdnQmkV3nLEP6DVX05eGgStu9nsQfVsyvGeuEVnsgfSJ7TBtS6GviSukEtIdzuqjjAXx
QjuWfWXxlBrYeAgF4wb2WmecYNNUpqtiQEL6ihHBzdhWMiVGtERRHV1BhSiGgLs/gps0/0d+QI0A
1e+e+QXDHaurz99Enve6G+9LYDd36vBWgW5/Hr4I6e5QzUpMW+By1AQMSIwK4t76g0YLl1IEh6wk
FgnD0LRblQZd7/d5AzqqEmfSmbp/0MmT2J2FRSqLXRInaYuUorg65ASTXEtkv8bQt9/lQG1/0WxP
p2jd2MQKyP2+Q1CIZ/LdUGUlVK6rEuw8zhR69k4b+8lW6dy076NDuuqqHgDs+Oa31d1wqTDy0e/2
1aui1MfKfTgbnM37huHue1huTToH43dTIfjgOGsdHT6APJN+TcemZIlEXdxsJYzdibqXRKS13bIs
NVKWW3A9aBAE+XGymncCUXOho6mXCfwGVkQ5+QRAD/F6YYFfT5+AWSt8UBxV9IPnxVJzvjmgsCWu
QxPzkKekCHYCyXvUFyDYvO82TnwLK4FQTYQvGNdGs1TuNPaAKxxeruQMlOWNCz1tsYsC+KALdsVM
bZXPvFVDawcMuebKJMt+ezF48Ji/DfJ6qUqrwJln89BeuFjdpmYozHgyqKYe2QHh+GY3S2Qd5pXV
f2p/VkUb5oI2Zt0GSEgZ9AkKka6k4tK1Z64cLiHvjDDIOhx4I0L1RW+ZNC6lWvRc5V6zNJDMcYAC
+nd1oeFGO5d+uzi9g1QCm1451+okVBFnB0rs3BvdD3aUNCR9kDi3ooDqwD66C9fBdSB5P0ofef4P
6U7YoQ6ZP6NPqBjgsz3qpVD5X37ZZJvVKpUtSsphFXGjDeWeOphao+arQCs+nPfQUuIconhOetaa
iQAcBf3OyesYon4n6De0l80vAz3ibl+Ja8NY9Jh3yxNMexXnFsAk05WSi6b4leiVOa7Q9SmQ6y0Y
+GqeytaeQOn2BkNYxAw+sZyChJ841y8NZZ/+9bxZyNswWWDbIftWZEk3ucS0bifQNfXC+wskAFE/
y00OkUf2niYxPQxDOWU+MvaWEljHUlpJJBho09RCUqGmVopxvXOGyCc6ekm4K6/26sNQSTF7BdQG
iC2gysVDYPzdn0/Ie/7iF1fII2hDd4bN1cyNjQDRS8tpxfMQAxMq0wryXcGo2/KPvU4Ka40+xnTp
o82PpC90ADCsKgozeVegOLzi2Fu3Vt2wT9FuAJBQaJAMFs8VfNtZ+aBr0f7WtJBWIEjWFddB0CCV
9OHbdBo4ANNjt2uUS77i/n8HABrlEE+znsuauw+3r89TT4G1va6bSBohdl2+Ayqz/IAdtN4FoNrF
r5TWHKuN86JoK8twXo8Fpa04a5mRBWjjNiPLD+4OcH5XZwZlkigOgolEqK1zUqrW2+LsSvYCIA9e
b/QUJQBTyefZudCibN105WWtvVvLGLYATF4bToLhzHIvQKF1ywIc7gG6VzeRL94HXm81FAWDNz7Q
2a2+zBYDZ8a1VzXUcjEf+q42sB3vogPfBK+3g5SxKsCAHpeuz4fO56GIql7nRNlZXLcctSqq/QtZ
+Fq9Z/wFLK7Tqya/kfFXGbsksa3eBZlwkCp9xRRFuh6UmWD7ntZUryMqhMNAPueDPkjoqDdnByjZ
fHROzUz7gxqqiwDnvZYWKr8sfrZK6i0y8CiJxwKIJmXHOx0EC0hkZjiRETkTOvwJivqrQZe7A+87
X88BRPK8NmqiLEUzfNEpJJtqy8W3YF5SZ4inew6LdanNYB++ab6qsvb8m9stDhOxKIehyILSTMpE
+MTle71D4DzMSs5vi4NTMcDNN3gRmMIfejfKRvak/i8lSM6GquP09+9bxWgm+zXAwgs/UoMLzRtH
+cv4vMSa4mADAYRcwxVj5dv0edarzFA4topRCsX93Zw8VamDF2uenls/kX9fAE45hMAqpg0q7nqn
rRlZjgXa2q/tln4ihYi+uZaYScQ4cOp1y7SUCuC0zMmaY3nVcw/FX7KmtVFCpjrXr8gy/4tF0ma+
JEFODq/JhOc75ZZXvBCYWwTzsI8VOL1ei2Hks32GvooZdgH0rVqbIdi3GW7kM5zQA6T33KCCg7K0
1z08J/olrwljMk57t00YkUI80HWmHNPgW4ui1MNNI5sHqo8+mfaeO8zhabf2bkc+m5C00qwJAyCA
WWhqzCESICeQG6synDlBL1RM/E68VPG2lgWdgn8VHNIcln8/5vtzS6DzI4w1N9oInWBcXvfFAWZh
3RxWkTb8OuAzWTGCL4mfEKCpDPNy6zxH+U9+wMqAFTA0epoa2sh1gEXEho7CTtstzdTfSv7y2wKZ
rlYraK09f9DFSFuScfSmco8LpgO5qtUz0bzMytuItBJnzWEBh3w2R2XkI70FStCnVSz1002I44eK
nAYWcpXp74nmetp0d8yLwnzpXZiwNHxybt4wOzqqY9pyqfuDOOGjdKpwjuaKUF6NZ18OxQMZDXKW
1ueqHz70sx4KM3phc28drFQNRxbOtQgyImUTmUGW5AHXIMvmKg29eAj9Fi465mKMT/y2kKL/K7bV
hCA66pw1zMRDDFTEnMlwR+3xwbPPuVbuiVbexMPa8M/lGVyyq/b62AfyXljtHCl9uT/9AqDAlWpk
HXOhni4Jh+CUpQc2/NOvKUT8R0GrG6c88GpEvWErCQc0K+lJnufYsds0mrkc8FMLsCwsKOljE8ju
KSwccY8/N/9OueQJJINXobFjokPJO7WVhHZYtEmPVfVS93/AGuXPTtPay54XNVCFiU5+jOg4tKSv
djQkSBsPdJy9iHy5a4z+rYHKZQE9kD6jkzYNNfYIfdqNvKT2cGLUOqFxXFJdqvfu4bLDuLX9G1yg
d9z+U4ez69AxfASaV/dYPnvDP4I2pxTpru4kGnIVZgMByTgtkljhSqcd2YxfonEg4s0yohhnEr+Z
+1nHjoUzLbv1/V8uUr9MYjdqd2n58yYWoqO36lmmwzLxwIz0E9FGNLE5fHVJcFwmkK0Ad17yvYEg
sM7bvr5hpGcAINFAEasLxJKy1YmD02Xg+r36q5LBllqMm9I69CwY8hjr5lPGh2lKm5TAgXjMx9qi
Ni0tbiCKPr2aPnlh1NSFSssYFGr3F5Dw7Amd+cJp+qDPjAl3OoTI5tGmn4IFF6EMHV80YdCmU2pJ
c+R/72c30xRBDVMLvE48tELGdfIW1iv92qlh2mvNtG51m/eEOjW9LNXjUPRpz36cqYTd8H9i5x12
vj8kKQDLp7hVIXrJ8ac0qtdNeN0Fxo0LWjLtfpodRirO+5K9XuQdUyKVHYdEgg39m2kLLfbM12Qj
GIJ73q8sHOtS1fDCUr244G8aU2/6jjrjgqduIaqpoMaZWMLPsM/jpJmk9Af12dS5rxUhomMSMThv
MobydWhwOgSlV1OrukOW1vbG/NN9M631ss8515Q/EDFo7B/6CQI3R0Q8yJtNaOU1wNZGaCia6aq0
YDJNE42bb8qSEDcLL5pxlFSakEM+8PsB72aTUKnBI6BS4y5Yh0D7y73sCSpMeZJdNyyFgX25ntPG
hssSZDrVmd4jd1u7LN92a/ESrpvBvaHjrEXT2KPkxbSnfIVou0/2kgw5QVNqEcvCobBH65S3YnH+
8H6OgCxgXeLtA784ya7RuA5qUPv/BYw1VybweTYOTwddb9LmwBVgjZ8yhFK02NlhiO6JKs4fwSEt
cn4BcSJo9BIMj6pY1cYHeezTMY+SXCACk3B5xtMuONYk+GCi3P78jzV46F6bF13MVc4Y9ENn2moX
Ksiti1fy6aAeMGC4xjNpeMVqVkywv15zHN+tK9g0o+jdgGXvCwvCnuSlz+vmDKVgy3/m0cJN9hvv
G+Xjghy9K+uLAoYLC8A2/6cKfinNFElIAHvBpfKI7V3YDQHWoOMx7qxqedaSH691SmohrWAxFvkL
GUV17ELLjUuf05nlS7nJ8EstJYXVaCfXTHmk23tDCaZXYeGl0lUtpuODIFLuFoplT9aDPrfWjyYL
vnFNSNFRp7yumi3vCVSER1zt5Dlv+H6kHOYo70qv18y+46EoPgSklGeRODdjHfQh6onm6R8eYLlN
uIb+JwLls1PqbJ1tmXONN4jWbqr/Dx3FwCmAqlwbe5t+EsaMx/qo2TxE7sEny7PZhMIpOtaGtVBh
UULXiZ+rtB3ydMjEVxaaxH1Vz1m2AiHK6acYoW4nyHdApD6E33mymNmCt30/Pi4hZN8XguWpw8Mm
rBmygJkNWHlaCR9FVWZ/6D9BbdNZw+hValDQa4eOk3+8FzNjw/DFdsZnYA747oHN4fBscQnjd4hq
6BBKrhFf5BipPQAxKTJgdsxgfILYzTfZoqfvyXGyZJQIxzZ/0oR7biSh9L1cNWfl1ew7uSZaHwg4
5jn+PpNZ0URIASPAspCIQ9LZUhktTYrrUSg6B6bpvjxKm+4Cy7lcn70GGl7EbPAOPQr7xJUJ0HQx
R3G2O6lPJpZi/mGAmRX8NMbh7Ftug14XfPFItcVxm5C0sBdg3WXEZ8xSyxvI2nHiChfaLcT/VDvT
qCGNCV/6rz3OcT4eJr98OkS8uHoLwLXxc6rBZrA3Hdk9tihaOA1VPvXnDRA6TOimlNJY+v2wtm9v
IoMpENgo8yTaNxfrm+TTKl2rRHpEAiXguHN4Y5/81e5Rw7SVWVH1A4o4dVwkNKqiWukshY7a+1P6
ok47x5sgqQRHMdbQLSNCPRBQ/uKEebY72bBgF7yqxu97DY6AR57f6OpirUrFvaQskQW4eJvak+Uc
HpRggxUcyOtc0/tdm4ur6/gwIKpru7GjRwB+J1v+WMN5NlG4LepINX22uTJJ7GoMA2Z6vQ5DKx+d
2q52klZvNKe/gFfXuAKDIvUhKjTgzDpoTEblCF7g0MeiVI9D+iSj+ASJaU+Pzl5/tMGPy6iENWz+
d8XlSRojtDS1gDj9PnrPViXHrMjjJ8yNItyYThcPE0p+zbBeg58y96RuQmbdfApeCOGMJzlh3prq
ljlGmHhojNPvbJfXRy0pt5dbAjVDgLmOrCmxayQVy0KxmuNgUQA6VdySwee/klMiwOp8efz5w4RQ
3d//iBURr4eSDrVFymn9ATv2/h1ZM/dHxgHJzRQr/Y/EAY/+ofwxeHV6bIVcdrWyUibGPcF/+BCs
+Vu/KTA1oEStgkolL8Jm8LIiGxWKUBIyZXCTe6ABIAiONhvg/XtDuWW1NgCWilBViE35qBvphGNc
kKttGmUD0Lj5tIz7+PWzqwFGuhb6c783iPRFRyOjFUQ+vjEz0Pzkpw/L+X3KD5VnTL/E/Okdiw4W
rMOuDkVkHA2R7r5Qzc5Figtwurv3dcPdNm7imtdMieCb2tTexkboOQ4YnZX/0aVx2qC7Va3BSUwn
GDnWr4fourJqeGhc2t1huCXYCMyrCkpZO4olA7w4ps8pNBWCfxO98QHctsvcXphz1soJn34gxbuL
0E69yiJTRYv1tdVvrgbUFPAKoaxCZhxYiwc1tLGKQKeedw/gEB/kGPkVJVimjRgNh0oYcZ08g0nO
2454PVowc1XFNtvFmbmhgyhvDRpiCZ22TQzy5a/Xx1uvraXm14jVLPVHn8XGE8wChZ7q3fQZQXiP
ol1773kf44dssI2+eBrEeQTGUmCiQLLrSKZtq7Z1gxyC6FvjRt3PDoOfShw3aJo970CMIHZEhtxq
RJSmIFZMSRZPitgQ1v10wx/UVewHWO7Wx3g+wlLVRU3rUExlSHdfXI8eDxGSLXNXrqiuyJXpOISF
Sx0yDElIuIAljOoxPZ2ITaa7S9Gdc8f+YGF0x3u7XBGBbY9QVzYJMzw3RMaVtd0BrCdxcv1SBGKe
6IY4J1fHj7cByPmc0CfC0tnRDi7td7xWvBdDbeEnqqNGBAfO5OZeitjruZFqpMnkVvD4C5R2E+Pi
Big6bWwHVilJ9jXJkGQpQg4LK1qcgHJTjkT9gJzzR7BpR2DL0kr1m1VkKr224IMpkN1nDmJEKIev
d7l/vkCpvRHnCRIZunwzYkx0hzpm11rSplv/tIGgYt9+Yn5Xw+iNfOAksprppbwX7e6gj+0DN0yT
SyG2xdT2Ve3GQ97nEIh0xNNgkhzPLYff6/O5Mj1Fya2aXK14u6GH7qLSi/6QZiI9+5zSne4p4pZq
XPhy1rQA7JiYel1CGIRlOOKWw5YJDrZ+SUOD8G+HdHEWec5gBgiUoAzeARsD31WZBoUcCH1wN12o
XGHEVTh6K2UhGuuqaOATzWbqZGDnKEz7b8QSrEzqHfIpo0hv/HtSRvBbaHV/vj6lQtmLRxaVGZGd
gGvnNoAKbmAYL7pxouUsG3hxhuwCjgUI1YCjHLNe3ByL7bUij394viszTt+Tb1oZVxaErHJEeJvu
rp9AhcQnYJNrg3vc9BPl50i4LGCVhmC3/wA956rhpaXDQYoa3IJzWWQrrsRq45VWVxM9afFFR0JH
bVAf1wgF2XyibK5acn7UvO40bTuvzhhYw1BQ5fh5C4qcUXCCd5ClIq6J/di0XiZSNGfIdILf6hju
BvEb8g/6MhlcNby3r0NzJ1i6K8WScNmEC1G7vr8qOTBh4yjjy34NhsUy00n76UX74mqcjQ9xJdS/
gOwNov6HEDMmcF6uYZUu++LvTHj+B4dNx+OOynA26FPpn83Os+azt9FzTz5KsWGHxLHFSeqJS+d9
3LNe96HrAhz7Elohz0ucK0vnpgs9gXG4rOIS4r6tMcyBNaibyiyQsVZjDGVK/3GGnUvUEiHQsHbP
N5leE6hE2uddyU1XNsMLUn8v2aL6VsDtI5SY8bAF86ylsxUEXhHgRxbu+8dfwrdrNZiIkTlnRS3e
pC/SgNs7yZYePXO2JVZF8zJoRbVhQyQiZsaE1Q05f0chbQoPQs9OLkt9FW/S6a04jf4PyE88fOr+
F1R8qq1yApW2h2gaGszIDt/TpSX0L3e8SGsnOHGzYZ7k3meMzHPHOgIES/uhscdUG0503JK9z/20
Vfp3cvjneO+fx2qbPZdOoStW91c5DplMEwaCykvp5Wus7dKAbI4hQaVMRSVk/Ap7XJqpMifWhWq9
sXbBvFQu6GoHtd3ZCbWBYlXrdeGwbwBC/ginjmqVINVnTNIXocDUNVVTZcFdkMzqMXuYAd76gZQH
4QSYtFzGqox48N3WfpRoIsZtzkZu3uw2m2EWuF5jTTie0d+teC5XcgkdCynFxG6e97ZQ2979qMFm
Yre52/IrR71moUecl7xj+t23Xx/PvimW9rY7MRI4tUJGnah3w2W3M1p/5HwbYPmxoENLlywfN3qs
1h9zHZv9ZDNVJAfiNKwE4Z/WWYBX6ZnU9GNyy7QXBT/uxHWy7NL/xWHPs6WvWB4cOAIL79BPywkz
HpHFPagXAcGSuw27OdIjRLlx9n4OuCSD9mvgELliOaUTAPNmVIuNuXrn5fbD+v+5XkvxsPu09FgL
ckKWeBSVHtMRY/2JObc3rcuLYofCvO2mG1CbJHnvF3udMd8vL8TQtcVeLopzOe9vci9rKavlDLz5
mDEspNBlixg1SrAvpWnU0R/s6BYi7K/s0LvZrHFk+fqrCinax1kxpWLMx1crTXt3W3OYBME976lI
r3Z+w3DkFTvJZKK5r2AOtLKNh9PB6o7aHYIb+RaB+SwMm6Di3Dg3LxjQ/FCyvGtQstYXeV1FYFyQ
DX3YQ1Nc7wU5x9m2dzMiPGJFVMqXiM0i2/WegE10g6WfL0JWXhr6O7vLnx1SoPbTOCnbzfmq8Ie0
FAb3mUZWcafHb4v9pDpAFyKGKBe6Twwl9ycnDcPNTl8Cw6cpTLh3x0V8JNPE5HN4J3F/DARQAfAm
71M/6lpFEHyupthPjMug2XevVXEOuyHMybnqCEZpFv908MIMBpppKo5zoBKTjSJZrzoqcDsARX4B
HO9O9jEg2Djpz7Y6s9x4G+7y0PXhC8wZuqDUnKCHjmxUwD+Qh3zr/G0LOZiwuq0LaG4HjFpqPVnq
yEWQ6NGLniH8vxrmzzkUofSboGFQNFOm7t3ZK4hLF4Nm4e6Emm5034eZEIAu4rIHFSvRcjIvcALq
qgfK7t/RvD76zCFasRH8pBnHMFlXjOuFWA6FBAqobuSKu68lZCozq8Wg9VJDX0sGi6888LONEQQF
YQji8mby+w90yLFGrk7ddH3gcRz7RyELodJh/Xu5rNKjkuSjeA3GlwVdutkXHD/HQ7jdUe0AigxM
QX/cjpuBhVqdYo6vFaYMywPrHgf2gpeVFW743hNKNPTtVScNnJmSQG9Gd3IF1eLi1hPTdvTDOj5d
QpuZzj6wvPSbiwOcrO3JUpdno1aPjC6186dCswqBzHI3vW1QUN7mWMNL2KUthWYRWHbuhbM9oTor
IQWCYBXFMOfJpioSmsYrSrOq7ciZi7XEPaPv3/YX17IyWaN4XVXJ3o0TrD9onai7vfRS0bjBtcqT
8Po+/8EsCi5qt5OsWGj+VzTm4qF8xWJiGkB3y5rCTnrcGIDfLtGMjXoayaLLVjVBG6Bkz4TvqeYj
AHKC5Gi+9Hc6ikAytJgkLE1dlWtOhfNSRxwvpXHQ2r8E9ab2Izpg9p+iOvY9TrCVgFqJOcWRPe3+
9WaxcugJ/wQ5yESNDYmZLtAx4v+fyxHJ7ADxe1qe7ACZb2xQPnUZkHDdCgFKTTdddcm3umCPzMtq
CXgRg4ivor48lEKZ6ZZAJ8Zx0q+Kh/8X/lkMxvqmIin/1P3/Y2BV9ee6l9/3GQQa8kTMhdB/j1X8
pXz1djq0X7a43Eb3cvkayIeZBGAGw0BHEt8qCLPm3kNz4c4LOdI4yYGtQ8hpxbo8ai2XvKmMqNfU
Se0J5uG5CE4zL0EMF5ZtMS+Lvq7Ay89AhjEZK6wEWlg5Zvt5L+YuQfLiop4EIUCTnH7T21xnY/kv
9Az5ARlMNOtcdQXFzl6CdhACxywRbPD5emutEw8H4j7JAMrb8loIvgar5JDdX13bKNQaBtL08Fw2
kBnZEdallAzWkRjRKT9+DF26QUEjmoMxW+Q3/vvqNyNnDcEivpN+/3zx6cC8p+8lvxhXQQW/K8e5
Y+wsuxd6kVThcYM29sDgNcvWaKTX0OGE041LmhUTLX5WJaCEhv8FyyBe7nmHI0oYsH9TebwYnUWo
BJt0trcRGotBl58iWV1DmLlfQ4SMXMhPqA0y6b7QQAj7m2vGRrc+3UY4mCjaHO5cK2/axtECE9Xn
lX3x19n+eS4TS646b7xTexKh3GlJEF603SOWqrXPCUD0T6yqWTwnkMIaEXOibMQE1HK/ko/ciGYo
BEgX1nlNEy2D4yC6WXFDRqnsQfcsS6xMJ4Rp8jVNlA2GLORDvTHa6OjZ0QYE3Qrg81z6+iOioQFa
WNIuUzLQ2X+5BOzKzhCsaA3GjkQPy7h1w/T2d5APs1mYEZzQ41OHIB0CoZnKK76mYzRFM7em2jWx
QN2pMf6HySL3X60UCtIYnseOY3H0uyvGMHe+fd+wzyWAmOBBZZEHSJrOUBCJIvZkAFum/GcNVySe
47g1zeg4ejnfWeW6dX5iJq2SyLT0iwE9qZURgVYBUVws+/t19rI4lnrxQeBQa+n0TjPk58i1qCX9
GRwYHg9B7siy9fqcxYfH064R11y5Kqut2ZLMcU8GjpaNsnsH181giknAtYYYYFQjVegFWWKhibUc
MKY9uPk9hwwgydQwlbKNG1eTG69WFmW/mfbJwiJd0lHvdZG3WkQxm12IaK8AMQv5oZGDtIRq/dPM
p1dhswCVRnzBQ0G9mJWPh6y7Rzvg6M5iLKu2Lnv9Z5PHnFMbdeUO+OA+mCj4KCrgzSHz5TWe6uUV
fo2w/m3GMJoJmEde3/aW4HFCG6aY8R9tTvlwj/0Mj7exIcRIeQHwqib+C7UHrfh5OBGyd4Ci5rjM
I03jKVQ6KTOnkPxE6efK1afhdkj84iXIkeqHB1WFuWhpTZiKmWjlXxvEnQ0e8r3iXcu4Oh7yenK9
Zt/tSkNoQ/Y8NIKKdkH+VvDkEMmyHG1f4dyhIV4eSbkDLF9P4rcjYdGLzmWKn4v5fGu/Ck/0lRh5
b8izOR7hgZ5/0YAfgf9UT9xPzQYzxyGl/V26CaVZToYW86gkEFMKPzPyjnxiajz4mD0tD8ctme7Z
lN9AGVWayE0fHnQs9P1d0lkO4MDn77JJhrHr6BGAXxLiPXl+ufVVKUiobM9JeGhCrBdxVFEiqSFT
Y69F/9eiPkRfCmz6NIWKNNw2oOOnI1+m8oiQOTvxFfOpBSEaMrb0zJvDOup+/eF8zuiMMXnYh8Uy
9MdJhNeB1w1e3FoKYQx75RfmB6T7TbJkJp+mhmtVDUN8Z55fHViMsEWeYCiCdpIdh0/w3MVLyFmm
LPNwoi7vfASmM1q1hn1ioqUiLkt/Z6wWO9H7bQn9M6DIZFM6UIebCTpv8Ysz/GQO1n5Qp1JUecE6
6mZdyWLcbb5PssDiLH0rpiswhCsYWx8nUsUyo+cJDSPrlXMCcR6ZWnkvH20KAt7FH0IY/KzzYMwx
5rc5/riXukmKzqKsdu90pLmdWtYl58lLutsuA4b8gXqAFAn302YOmWV2ubIiC/rje87gYVsPtXSi
gs5NQ2H+tVWbi9ilJUUY/le2BNxJyjds0rpygo28nQMtaRWb4Q2iGtrNQImoYNKG8ETsRziDNh2H
45fluK86+0i8UacauHEbq3JnuhYqLGB6VmeuU/E2JMpKBJ0oES6kDMB5kA6gvsvGe101SGwqdqUp
+j9SpH+ApSuVJKGyyojaq7DGmtmTqwGD1+gvbI1jxzqkHZTCysmfqMBStoIxnWSV81LY4W6+yIE8
10O3dRv3OsoW6/aY0+URWmzEljYq1/IKBwrJR0DqvAOEzR/C92JIqffPDt0aZTW1FFXaDPL8hHUP
MFLuch0oeRZNQhWaxMxg5lU20ZKCc+en4XTSrviYGgukacEXtXkaq4C3JXc5eCr1vo+03fhJk1w/
ohCMOdI32fCpkdFH1zrEfS7Ihwb9+qoUpv5MMKMymKAwhzTMX0/OgIMfGWMRcBDIWWC+ip7ygt7J
tYxIQ8KIeV3ZmDSXkXiXqF3VeIIJvgs0JaFnksM6RqeqwfOYjIHOHEzEWSsuIWVhTZx8B2uwtAbO
OxTvBmM+9LrjWgtFXK8rMHLj9uWjKy+JoZe3O57JiRcta0XamTmxL0tfLcK19xKC8UJXcG7QO4jH
N0AOaf0+kuT7bi0sWqs/np5bjd8hx56EwafbQYs61QeyckbxF6gmRq5XTFUMpO4rcv7J3u9a8w5m
ef/SHnl4sJDYF3J2mIyTtfF2/6jZbJam4po/Zr61C+OlRuZZjeC6z+Ed1+2WLy9UaJxz8QG5A/R2
zjRtOIK4T8hnKM71vwwQZU02V9lGT//34CQbKgBcJBGIPdkFVGEdig0mRCES5I97c2zZsRdse6Tn
feJfWKtCKZpkTU98TJoNb42KY4YipGDhdxMAgPo3edlxBlCm/XEAhWjyj5k2Enhr3enPOtpH4qja
c3B8yMsrTVP0K1Is3iAuIf4mua4FKnT/ouDJtSxE7ppq0+Y0a2AQkjPCgSQ4CDCiKeqCz7bq7q32
MOWUekujdvXTB/cJQ+TNmSFTT6AImsKlqh24V7gcit2psrPavOD577A8LF7tD6+HJ2LwKqMvMMrh
RoNHlUiyQrUCNcwEQBsx/2DuvKpSmlySUwBFj8s8wpA+TqfzEQ523llS7M4DHgkBs7N4oY7PQeXW
JNeDGqI+D8zPKqV6EODgpy7+MXTSdCEGDEn/D0l7sCnVGB0LmPhMQgrociUYqbygty0bbsf2aTN5
3cocR9DDxke7BxZ0xijikIZbIda1B8hzaRLxG9kJUxpiIVB4cHmm8wNs/d9bOT/Z7vPnBE8SmJrq
/kIkDS75trPMox4D++kI3QtKmuV7QryjPFuAsgwocvalwkGianxhmBduS29rBXY7/vE67Q/vbn0b
C5OEmzEteX90s0PJkDgWWU+EY0Krn651NZNRzThJUwBAuqx4tp3ob5jHTQJMJXMr1FEyt4dNOK1b
yjjY7GpZ33X9Apj0JR0A53Wa/bJli8ojLkObOfCOMvhLjFNnITMl2YdN2XYARzao85l7qZ4esMXU
7EV8FxqLiDfztUoDmtYE8m7XClpSIN01KBcx3z0dlkrkH/fzMFRTNgasRQT9HvJOKeHmFCLC0ri3
XSGnjBS7+t4f8tghrk4zxMjuhHosqm3KFhmCNwFXh7UQFPvibEmO8Te3j7EQi+9dz6QBzw2SoFwQ
VzXXlyiTQBQmxnReQZolG6qt7Vy+MV8Eqtd5nkug/Nv9dXyQsLCwPSFHgXBYRiSQ63fHrOobfzOp
ryCEyVxfjDBM8vRQtoe/8RL8Ov37P31mZNzfWG+GUMgYcjF8MXvp9hg5ibZVfqv5bMpg8Q2T87tK
/jZE8YUyti2UwFfVIzdoN9+OGr+wV0HtOOu55lG95782JjmwtqZoKJ4Z9pLFcQ+8xZJzAsDcIUiA
Ded2LIPcskRDvQm16Xyw2FvA6/8qwlIGB5WzTnfQaRCz/Mw0Gw3Pu9YocoE+PmfhU0SGuuPiTzbT
8d4frBk+eGwta/InYBubNR2FUPZ6Wh4kOH+3Q/3c0druf0H7aVgWouXZZZ3PP6OoYE49Gr0tp4cC
fSRyTEH3bFOyEYvyRKaFNIqfxspYRmqwkODWRQEckbzAQELNuI47SZ9f0xeds6Ah2w41qfkOQEbF
NyC14BERm9XV1IUaUUxn9iqA3ky5QwumHH0CBgKU23EKeHqGNXu7cNE8BBskiG2Tj/FtwZohWvFc
ZbG4eanJmgRPCV5kwpxvl+Mke4MypLeuToT1sIRpmZ82Ri8FwKs2FnOgv29pyYOoZkKH0A3WBZ8L
fhcPRcAVBsFslXtwk+slra1zsIGsWbR+JoqzDGWz6gvZj7uWWE1ukB0iDe7T7/issVTxp0BkkvpO
7M2bumSjg3LVWuzdHpcHyLwYUGoV/3PpREmkUcF2W7i7BcsJUVi9FxGJjhsYci9OTbKREf1E7HN9
JMX1j9viWKYjae4kT/ixqfDwKb523NlOOuBYZxtrqgZ9hdeSwvG+3GcxhQnFjaL/Kv4+/RmumkPc
4465Bs35eh5aLdKCYAyc+gtwtPD+OcWAGAMTYlZrklo2eWjXrXtU+n+OAegMY3mW3Q8lfrEr+yXa
3DwiKRIwlhMMTzBEGsilmOOigbQMIdTngbTmbtgrmG6EWpZdJnvEnlH8PhfczZaUEo8IToZwAYRl
1E3M5IFa/rZvtLDejZgUpdYirN/eXZ3dqaZhi1qM6rT1o1eZedS0KDMkw4V/G/oKRmGm5b+WQQlM
V7+/3IgMgIQbYawKiNqP2ZHwHT0nsAxa8rXd3o9RiEynGnBOcLEEO4uZgCiQhOJcK7bz/KMmET/t
G3BSkWjpqXmBhKxlqjLn6yEE250FSf62kCmCjDw6e+BHiZFORdqYeuD3/duwcYIp0c7ojthjfhkk
p4tMylWh27C83PgyT9SXq58BGjLoeeIoziQrYJ5a+49JzJEZpX+QdKXkHO3wgiPJkTIqq578413E
Ou3VYL49bvqyzBnNUzPttryYrQBNZ4RDh4Q0vjHkvOb8WMvOW0+YsP9zadl7Rhcct4d63QcRxoxg
KwHUqqCy09MIK2Sknd34oP9unxVZ3u6pMY8dwSbaFZxECM8D539Hbyry2sNaxfo90eWD3u7fmGAh
6pttA6VjwLk4DReoRTULk5WWQCKxHGm0rDwcYgO+f0Y0XlqkjqoaaRE3fPVdGCNvqYpY/C8TYnsN
/3Myd2MmhgklGarYUXiNigztzLyqqc14mmX3WnYeBnuRjN1Ht7RfTE1+iujG1sxNSFwHCdzXVSI/
hYLXwWkN8u1gXxwHS6nR/ttSIfN6+lAzAbAYHuKTRq2PBchg9JIqm6DNsqi688yqt+eeYymLw72s
/sp3rNwQIypkY1GLKVI0H9Vgo4AwuMKjIt8MwnSTsq1f9o2q5m8OU4fw2/6vNBUkmtB9S1+p+3MA
YzmnKMVgN/c8gTi5smyNIMfKyNrnwz95XAjKyjr5Z1P7un2A8HaEbu+W0UwZoa8IRVbu5rcyWcyN
tDfwwhwbYyYnzKVJUD43C9+iGajNtJwCBUkFj+CVYILUiwDV79zy4zWFsTcI4ZqRxdZkll/g8X1R
oke0tkx3um3GwhPdes9hOQ28wdtzONJVnvfjqdwpmEzdUaxH2HdYRTTJDQ2FNEyul+HmlQvjf2jR
bgxuD5A6Ugtw27VH8b0KqfLlvtFPhXObdU9qTYOVCESlEp9eJLW+URqF+xO8zpEDY/8sEbXFGmpG
mXPv7fxDzRKs2s+fmrS0Q5mzopNccajJu6Pgfz/EzZxslTPPOnpMan66bRqOrQUyzLb27H6UNBHs
PVLgUnqNW0ANOeGcbNgr/Gl3ddaX0xyu37Ls2MvIOSL3k1Nqlyua23uhYXv5nNgx0khLj81SujMI
wOiPxyPiwzNnkNUY9kb7HIFuRplomB4QfAAo4h+VMc2LUz1Q85a9g+/pA/cKhGkbXEXcfRLCDMza
bGLZE6FKAwCsfXIMzJafwN6xk4tEPFEV/PiVOQbgAezsI/rTZt8gmTboutbHzwD3sYlL0f2IwGn3
V+F4VUd5pwYRVFbU8kA8V1PUmTnnkUM9ukKGwDjxXu2yiITP37qMrUbomVrqKOGwpc3hhv4N/IPU
4qtiPO0n/uEL8U72kdOET2ubz2gujFgN0+3WVf1mIpxbVBGvnx/wn9WMgnkdGz8skD3NUgRWnXC/
1xzg95XrGpAY+GwfxkLJLEDFuX3Oh1738Dk35kW1fyxoHO4xs6TqMQsqzOpPHFm/9Dot0BL7V7D+
656Q2Ua9ASeLj4YJkGenp0xoXLx1L3udw3M3+2yp97ya2rkY3VZ/iH3h07+PSO71jYFSBr94Zr7o
JAFPA2a4cCc6xSYJ2/HJq5bWrjjiSzUHZYRRDnN8BW3c1AcQj5wAsDfMLDJFIrB6B/tYzaoemoyb
khi34T+DSiJtMIgs2o/fU0bZk0+V0ovi1aB31DfR5gnLH94p93vR8ZF0xsUxbfdDZTJp8X2NQXyx
zWCP4Euk7XNsuVfrbFlTAWnnqnZnb7xtg9wW+fZvKBhfhfuy0oClPkI0bz1ZizEg/hk2NFeSy/2L
XECpG7ei6uze9jWBEfwBh2gkFUgnbCFm2Oe7l3L1gVK0zA52AumtUzI66y4XU/QbTJgHXD1GuUo3
49AX5QA/6mG4cArS5cbH73bS8QxPeDS01GGvJ/uV/q1Jv4wgfci/NB6rrzfmZ0rNKXnTmCCevIAt
oE9FmDvpo8U1/SnUHiL+D1F1A/rrIGZFMFf1o/+JP4trDx7tll0sjwq9chaZ+7Bcw9nheSYAW11s
bxCXy/0l7wAv2TG6LtoOI27aBamWH9DL9yiqDC7urjgaHEB0y4YeDWg8oLMHcK40TaE1eTzT8mHE
fIF8XDINXAN9IljRRizmy1f8r7bcYg5AMfqV0FvgV82a6/amGhk3biUuIjQUjqAoe8F063DVGgGh
XbOPjLKvJ7sPcY228Ay6pTKoHqUGz42CBGjK60xjQLt1wpziVxJMnMwiSY9VMh05yTIHg5pPfMf6
WlsSpThk7cJml3vo+XCAaZ5ghBRETRReEzZrBBpYyQ5Ax2rFqOz1qB0opB5IUR4nePjh/feNEuXl
RQA5mzySiy6/rmBKOSq1F1E8ht/wbuEXkgu4zMXGl7MWyYQ9WjYXRj8CmJzVeFxr0u38erHqcCNi
XRKhY0lFkwH/GEyAE+ZAzHuDk0K3VUHOABsUo4dk4Tp24sznWciTxoIUy+hvNfThioB+R79BwYk1
PWgsuqqMpkiZvzGxtNr1RuOiccOCt604M+KF1v8uuJ8lYv4VT6XHZqrKS+ykfQ+RPNjFbax/Ogmb
OjqWYqIRpLTw0E9C0kI7mwFRx3uDuqbx/1jvsXI1WIuc6x0VE4lwfcigrTHBxL4WDR0VnelUv3g2
GzwM6jw/oJXZ30JO0TAfl7QYX7UZTUEVhr+7xFUG32vXUOKTvU0kTy6mxTvHs8zv4KJsvG+DtZY/
AqwxP/1ZmtDOsMfPlZfrvHk1NVMjdeuRpzO8/OCQTuqYzhal/SZAYeIzZxYG5wxc634c9TJJswpX
AwfcEcrOzRRUaUHmBLbVLSnWaSh+AF9TMqbK6ijzmqTEKiCr8QgyxU9Sntlt8JH7oetrlBAouJPg
hZfF1fOWaZ/livjvlhylyeyTnDSU9i8OmVQJDzQZQiNp8aiyjmPQNDUz/Wx98cfS3sxAwjxzVJHJ
cFEBv3NgRONb/nzhW3OtdkFqXU32HgnPhsyfcz7lp5xtLJ2ByKUlz4TXdtlWEYBS+4vxy6SSMAXI
f5Q7s/c8Zy2h9x/GGV7IBC1snLBJGOC36dx3nVUgKdsrtr6tkwVMXosx0BDxZNzVgH67Jhx5QECC
b9biClFcmzzjxJFLRrAouI/l12ChMFbAleLi2T7gMVJSlyI0888h68jte0CqXxoRRtwcLk87Az0H
x55ljUI4yhwgfiyM1M3dJBCxHfzWuvZvl1imGzDMcA2ETcKlfFH0FhSiijjlXSSo3/5ugxOSHrfj
kJ/jt0VAzEpbVuCJ7VZ1u7sc+vdfRPU+4LdSj1Sx8rHGcFdq8qKYx/JW4vdtT1ZsQ0zJTzX9oKjt
Vlt6wVr71DYhZoDQ7hh0qaUPLCUKB5/ykhvOR0uPuke076Trai4nVmhhQ525tT6RQ8sUM3tmEAAl
ZTshD/mYL6ZSQOsRqNfs7v97Q/aRIQg3sCzStStTW/uPYPXPDtA3/7ijXK0eYXUZ3J77FNBnBegB
nIQoKm42DaIC7dlz5M86L6KfvLFG/EuA9jhlyUfw5MUgGAKh/HKHXOTlRAwYWvRxsEDv/GAYPeyW
asv9F4j17UkfHa8pG8+wsvyoRM5QkG/NFygVEsF9Y58zhvserNFZ4EGWxGi7U7r//eo4f9OoaIY0
TWruOkT2e6hiADhz8TICxtRrffRtz1jEIl0fZhGrzxJBPNpv/U4J7oZoAifrFr0983ABZXnBO8Ma
LXRNDjmnWMVrFts8llVfIzLiImejQ0ug2EKMHV8bdOdznbS7AtW2ppklbvIZqeFzU4/jj0xCCfDs
4g2oPkn7kLGo6gkcdhdPy55e4y1aw89KbSmPzdNSvR3d8/ra42/b5bvPtFgE8b9xxwSWwpjjIpoa
Tp9gHFk9PmUIn7ucLBaQ10sh6plWcgZI9OnS32cXGt+43XqaZXLuHk2gaFVUsVewjEXxj/P18D4y
Fws/tc9BmZ+MVotKN/Ja62pACBWIfLNIJTWju4yJrqqk0UQB+TXOUVctRNJBBNfPaez3Rem+r1TC
TzexBBlD5trV4bwQzfp5MS0hjD6AFQoS0XCZkg47tNIl742oppSf8VCDxNWIW+fRyoFEMgSuyf4Y
FVf6OS3DM1Bm5KmLda7QwuqSzeHu9zSJ1puAChXe/azBNWFkjm7oNcE3YdfK/1vxmtCdRSGEyUnJ
gKzFVM5k7JVBFPcmXDObdOomCrFe3eL+euCNZytf6RrdQY+kX7lR9V6sb+6rmIyJ6pI9S9LbmyDW
hSPyZTuwCmNlLsWjLoVTFvl390GhsT7SgR9jsaICP3jCwDVr1h7OEE49JGo41beergV8qkJpBUN7
CXtOI+pQGgj1/6GxWHpREVwVsZaBpBfoHUSij78oVI+bXYc5VE4rCtwTtdPC6PfVI53CqecCmCxj
NteJnrUVKAibgowtqwBJhK49GeXo07mgL6i1xSbUyvvRmcdsnZSyydxnwrelsMeTs+5PuqjVilYw
29x0YmnvyDuuw6x0iBXVXmqK1w0ixqHtvPNutAzS5IBv6eZIzSV7DG4KrcWcVLlll04/bo6LAP6A
3J8/GgloOBZx1NilfZ8SJmcrU6N/wqwPdu1SCnPbRCgHfIQk58k5H1RpZ3veEOPCY6Bw2mny/vqa
H7kPkpPyKICi1oRMGqU6Lt59rjPVlGanjJuN6jH/PORSqCQG86kNiR5NQESZZxzY82l/Bo4Y6XNA
TU9Sn0EUGVgsEEe7vZuVS/gkvj2uHEWXWnUrlsmisqchO+S64TIr2pe8I/T20FOrhC+xv437Hr2R
NQ0UqJrgQ0s8FPA9xxX6zOBspNFMZ4nJ0utGjivA/yvmFEJJA9HfTLk6gNxNrk6dBMBFqP92jYO8
IZeceOFAZ36C6cEB3Ppm/b+aohXgpCl0mMEGGon8Da/O7Bd6fIqodBuZbHo6QjktHuDoYwZtZDQK
NQ870yOkRBylFq82GkSCLh6TGa83wK+KXfcRtDibdEGoWikBtHnkCFA2IgC0iXygBAvuHAmsxrKC
wkv+0c6EMA6rO2xJUaicOfIX2cF3e8qyDLm/ZyJCnKemKGb6pABtz+Xl4svcqVa7Vx0wZMx2NXV/
UK2p6aZblZ85B9axsZ2K6pcVPZFWVmUYPgqTGGYzHSw/+V2rROxzqiolJZjE3cgIyNOX31oZRLXk
IRONZbto8IIsd1doGHvfS4L4wm04r7JzvUUatby0j18caXBUCA83rrBMX9AWdTP/0UUxaNPyIqda
FWeGKdBA5W7wPiMvSo70+jB60g2cWiW+CndRyE8Ipt9v4zZnAeucZMtOKWkU6qYr4TpmYwKuAPgM
xQi5ohEy7+hVwHujm6QWN5ahEkcE3S0fSBa8Rdno4MGigSs87+0ugH0tEl+Bh0l0VGk/Gz7qCdcr
4/xVccC64oabF6tY28EhwQ26mIfhnNNtcy7rbLQI1Tz0zTNp7tpHFBE+UOijDUqLPGuuuUpRXGKB
z3IAcEmPcK+z3csIQ0bkEjOXXqqDkGT5sDHQ9vImpcaeoViCx5fjgdFPLCzzTK0grJIpsmJ4VCTJ
N1RBf/MNCRJoJQ7SLoVX6SJjjq2TXLpsACPCj3BLRbu6NaFOKwy+F54ZplqZMXyRyGcWelLWP1ZR
Fi8O44sfCeqVhoNmozLy9gUMEHTWt+ne7eN6xIQOhHIufx615kHIrBD1ptr0514zbAvrylD0iSGl
LCdI+4QUMbgvkVRxflJmWgqsYbJ2rzwEg0TLJE8ofIWwaqeGAIKf0KpGb3X1eFAGbDzHHQTi8qoI
1pIfxTTqhZ+qV6c0cuBS12Hamnr0UIC/gfC3ITMRxq/OZP5zsfd/rgt96gHlME5XipuE+81GWc1v
nd9+iOMxEMx9JeWku6SsxHSlRPoPXtzJTfsXdDzIVSpS0ZbOUZOqp+nQ0yd2rwjAJK7bPMu0Vkwb
eqRsbBOtjN74qU9s1Ob1vGN6yAxUwLIn5oQ0F9v5k6UdS9vplZpuHN1PEqmLAp1Dj3/CNCt7ETqT
atFBya8szXSR9Mmqf1uSwOSHWlLhP95l66aUeP/pIleoWQw23jvxQN6QS/ynwMCI2XwYigNtZa2R
dyeW7uMxV2CaqjyyqaPBRFL4UayrSdYSjti0YwqrKnmQ+q4MUjnQ5oVj71IsDoz2q/CWwc4ZBc7h
Eg/njYPAaPFxApO7L6gYSQG7IGN7XC20QIxF/8Yz89j9hB8o6wNLjR2wznz8IOoV7B+Bkug8ifSZ
JNovLx+pySbyl7sBtw/a1ozzTn/AMZtZv4/jCCwEzZwBgziJhyCUQSEWvUa6blJrXxwGANOuvHlP
zCnqHs12BeJ2HRoIz9LcfKGzc7eN2sznhPL2MfAsF5xwtswFDRGmxPnY4UcNNvolqWaCa1fpr7Wb
ZMl1TruRUM212y8WZj2hMwToVnWOgXcgmC3/PE/EvUzI543MGGfkEkGUvcT8iD0RkAYtr00oiNs7
sogOQWKS+n0t4Z9j928zUaJY7PckhmHXXAYoEhUCuyqseF2vPa7Sb2jMuzvryaC6knUhAPRF1FHQ
1D5cFLHAg7HGKfdEzq4Bfv8CJ0JqiPjQTPSaglhihRpJTC4Sh/wKaQUlI8DIn2TTqhGRx2bnDFl/
T7PeRgiITTX2Zph8tJXQ+91+713JIEhHcT7P7fvow5MS06N+u4hQHNF5IyL7c9C2mij/+QeqPaZD
1NvzJhXp+vQc7A17muNiwsu2xrDMMq+Kjrl9kbqZGeUDiR2nDw4d/1Jq7DL8L/J5qG6/qOurgaz4
6e2ESDFfJ9LWMDWPpS+3KXLwb5ymzVACtivFyn0VMuwl0brjHrE6Z8PUViujax2NP4NoUPftp61s
qbjaYwMk416hCtfQple0vX4tV9YgtCn8t+Abnc+JEyG9V4hRfzbjTkglCQbnuWZzwkX37MJS7rKB
Gl2JYqv+hXX7u7JCMdA4cqBS+miypdLLxVbEuhoZq2JEz8AZOmoSV/raOUTfnhUmdtxfqJlYnIl0
sPXtl8BtQLFwIZDvqa0uxBa/OvmHvM/wPdTUsdYRwYml4R4kDLCoHmpWlld+ltP0wokbZVY1xsRK
i8/7IWTnjMMxKqYQ1umwF/4nzaqWWq7D89U+t7D8UZ5d8lCPqp15UA1BxZnsbAZeC8DmWFLHGQal
WPG6o+MkAKQOAhyeUZowk+heKVVfQ2bCnWF8Sc7HsWseBnPgj5lLPQ/dfB96u80S9tMM4fNc/TI3
YeyIhk02sEdDayjEEL3lpL46VRI0nTxpfOHglBRCXXFMIvSZ/ymXRrarybesa03TfoKOrUyos9Sa
P+m/GGJLsQ26Ck/RwIQyuMwB8Oz7lkH9EfOSeRjMiYHPySVOL0pyPA/LQFxzR54wgwfEqFv1cA0a
2yawAs46y4wvwoKUhu3hg5BRe/UK3cr74RSjpMw++iMwrbkgkMG1vo+Jm7ODRpZg58SriGrrfE1w
0mQcw5bqAHpoQWnLZy4ZRAt0DdgNeFjD/i04KvhXQopCWUMpjZWtZcYNtWtPMCQDW1SLl8CD7Jok
PgXeGkenMQTZNuntLLj0tL+65NczcM57ge285I8+ZWUMgu87pDD3d8bMQIFETZqebcLQAb7gmP71
1moPZkxmdzAhqyVz7rlavcNSBmjOU3qA0ckJIJrBRa44dnTOdhzHoTvhMIdCUwwrSSY9FGJpNhru
NPPkglv65ovdgnZfVHTojgiaAGwXT4/Yw9xzoZU5iaf5aPfb9mZD4xnxmIEaTEwJKiypDUf0o2M3
EJDbcRNx4F480QzKlMQGeByeHXA4VFG15/OZZTSG/kJNYLWRx29LO1+Aw/Aa+/SyhA6lmgWU1QBg
T8d3lKSn2HeWdfivNFdBySZ5jnFRTcSBKGM8J+GXO0RzNZUJ8QE4nfB7T4zyzi3SvZNtOqZTghpy
dbsAVmGIbCQd0JNqlaDanAF++Bt7mT95cGOZAiJfh2Omw3o6xa3UAgnDAdsAOdyWXL5rntyd2z6A
VTYPZB4z+EAMpQFXlDueWg0jPr70eEoFdO1F6ia8IqObXUcW/ZZQNY56XN122G17WwU62oeAmUBd
If2rsyCZ2Jhbo2DdHjwL4576HYjGBhwGVOeCsLxRapueNwoyOHXsQn5K/DEPtPaj5BLGTJwyok6p
szJxiJYO8hCyBcLFQLpjJLrNCwvPczzFo51jewunDO4BYS9lSis8Qwo+DZc2cQe7N8t8u+pcNR1W
5ZNtJBh+cjfQb4PB4ssHQtTNlB7mL2iqo8UEY8NXgK1245fyGOqM9iyfrobrdGYDpZh/R3zk3lYJ
j6lxRM28SVSa4Ayxo6quNUWXG7usOsFdSwkd8hMPy+sXlxrkSb1voDrSCexY05pY1Q7rRSw3ZcUo
8dyOK6XhFfmoEHo1jp3HLT17NBUXawVR0acakb6t+LJXsFAfZ71ehjS8Lk9pGro00R7LU7Nnh4sq
BLVlJCsBKXsr8p7GE1S4GWHMgel08Cr6bncuvXhzKsRYS1bI84rsGsXRwzmGXRmASDzlxnRPPRhI
pFOBeC7tN2H7BIrXv/6ORJHmlJpxanVNby/1utZFN3wFIbG1vH8tllnAxlhVUiiIHVd3QsI03Ouq
9iYJGwT10OLsP0lhpXs9FCqygdamfruyYzlChwP+4VwjQdGuU9L/6Oc9IT6kwUB28o3ZCVgFXJYA
IX/74MBj6M0+J2UpLc/p9ckkweYzvLQiXFUja+yIdDiK36FgqkLrTanvcMjZzxn7tEyNS7aVzWRF
O2PUOtXCAxGwHTNWCnTeZFnv7vBw8izFTq2C2q1BbLh4HOazBDnnI7+QESXBm38HbWuAOlw6ZpOZ
lBsHH2W0DclQICHznnbuQUYR9dL2MSslqzoL+LWyZqu2rGM4/ysNi4xnmdtMiq2o/g9I0D35IhZw
vPRV0pe+fCo6kMB50biEFxiWrFI5CQlGPMZaq6c7EZx5+PCiMBe+kRXN0R/GkjuDr/S+ZNayEMWI
G1vQfzqkM6WRLcvPUS0V5LKzza2V0vsu4yoZ1JRZ7mWjdp8lAj58ZG0aUcUBFYAT7sFyPj5Qi6HK
YMoeDpgeX1/k+czkcH21nd+55UnijivWx8UmGjhzq1GPXyyv/6cjauvvnyy04KCgFfB7XyDsVPh4
bwZc6jEcLWlRWgckTscjIvF/qnWGILkOT1px0qP1prF2IOqnSZtzvex8e8wYQJ8yU8xnFrSrgMvs
X1BkUukBybtMwg/aJRjj85rfzVL+nIfAyTgs9p/bAwhDam7ccmlbDGY7xCovpugF5Hs8AgY6bMp/
0Qbo9eZ+Tp8fEkg0GIE+PDw11Q39hq7v6TW86quEkAcQasV2pJQEGfK9GCNwr9WrgLPENFGtP+e4
+s5GGdWY7X26mLApzZcqu3ifXqPTpoepaBTeTagVeYWEwO2jdBc2Vwn0Nv3M7652w7giB4Vi/tfE
7KZTZaIRq6EHUkMc6VXZl3uF0jyveQtpNXVVaTQAIl5ShkLWA/MDmWaQAqKLk1hVWJ7+mMKd9Pz/
hhDX84dWVShm8jrbISQWUVYwIRw9zn5hpCxrLgkdu7vnt1XNyc4VOMnGsOWOrSXZ2BNDPmbzJGmH
i4m8n4hQlEC6BsLDcWNxae6jCkLMh/bW7+Vls3oHjgiR/ejs/zzS8xPQM2ZsvvU/s7VJKAoQrNQN
U99Q6bbb6tkwykuvp8Jt5MGh6l8nz3uZ/W3ZczltPDifDh9TykzYlBQjSafKpnZJkODJ2RiLJAZB
Wizipcc3hHzpc10/yt8AOjQmZiOzGdzAnmsYFTkgW68YYLQrBbWBx+iNlwPFgdmtW9y9suistUo4
8w1RrKOYUEktde2+sZgO5s/hn/2IM+0Sy6kQq3Hfj7AtdiTxy4Hf45v2OGDQMHweBtz/mknuI0z+
XvI/lqaZge/DKEgHSHpvxrjjf/Vp26KJfr+DCfJVjTV+92m7CVOJiZEz4pAEpyh+d2n9PJEYf5K8
one7MD+gZT7ypbrhydKeuZZUl0GHDMkGDtTEJyxTq5uOxxF9biTwFKXCOb61ASDjGro+64VrY44h
hkv2A3r+eEHLcJWNxShOcE2XBdH0z+DcPx2Qtb355/qkIemJSz4LEJJ4n6go7fgw1dXii+0JwHUH
PnJiJ7q9eoWuEbzQ+jEdAPxFn2s6/nP3DG9XHd7Zi/dZNOF/58cBV8It1V9lGEteyWN+kR0o6Kr3
bfAa0nfUZLQ3IFXFMZltSP1UyC43O3qKdXSat/nsZV0IYvURME4POzyTuz+6934sfV7d2JHqMR1D
NxQJJxcGokbOO78VXun6ZrqWTIvJwkPhU+nvjcg0+CGyKkLq4Qz5r8WcEL3aS4YKFHqEjYTyQ2h9
0zTrfHvDg5y105D7CT8Vhu1rrSqhBUmtsHmLj3z9XKzUPvXvAQMx390AuKC/ixTSaci0r8PtVy8R
nEZnA5iVjM5lNjVnqHuPPYOtUp8gMgDNBFTIcZpfw2I5fBL6aRnHYJQSn2a4HdOVIi1usx5S7/Xp
NHUuX5RDHnqzKyriD8TZgfbdju8y1FI+5kmokDZHK5qLW8ke3x2M+M5TyKrBGXgNWDg1ZEWAqJg/
XZk5VKRBPaXm9jlFLa+xNOKGcdDTYg7LAmBwi1udqxvki+/2aqlQMSCFwKW5vm7lLUCZZeMdHw1P
FdEko80CKUgEZtFiSORc1+PFY+UYjtX3zaVXbeZupTCxZTQqYmyD81hXGxqd4mkJfpsLQN4mHx64
+/UW9khSHclURHgCqLCQX9Izgdb93AAvEmCN/sg9kORRmDs0UM+NUT/2OxpeFE0DnMOZphor5Zsn
pXHU7sVbjOfDO+xxoz7EQmIbeAiMmyffQnrVnK80Vmw9S5W7HxzU9VQt7QoWAxpDqCBuy0t2agj1
AByd6+R8e9KaKI1pbC8Sh7yePQU6LanaFzYpn7sxmt74Mpe0Tq1E6hjXTJfBZ2oDRjebop7XqOBk
UidX5hz/0QI2aglSnMH7iQakYgb4FVHGBOZDBzhKxac/wp+YTT36jjIOIhUrf12p90knmRgZhs4n
BQIJeGl2VIqKw4KyA5RtBa9+3lZoOP8jRHZ3X9ZLH/QjAekNvQCqTDEhPxn+0zl5fXfNksRPDu8y
rWzX5EmLJrOufNb7b4NPiDBDiUJKmqdxtyHKlWhty6ODbJR6I9MvhXXsmiLKjrHeGPPYsyS/G9j0
3iXi15xFt9bYIMtyaPTYBhlTckNgypwxG7vim81GXZ3+w6kzRvyAKDZq3XCtqhWAZkimo7zOWydm
MLzGGFv+9GXr+owlRwMUkumlNh537XXfSiqe5elkIrp4/Cj1+6135m/X9Fvmnq8goyN5bd8wqAvb
j5OGFmgtcDb4vtE4VEJFZaQdp8k5sOtzs/wCsUjGGcJXZ7X24j248ZGfj+rA+rY25sWrTvsOU84w
PAE4fyuij64Aqy6BUX6RA74VC+Q+/w/iOo3b3Bv9wwQwRfU4aeJLekzyhBpuDDtCQfXfE3PN2zDI
DPPn2JGRZppvBztSkjLq8L8pIVpicNkgHfCPN+vIA4vkUqPjhVJZ+7ww/Sgvr7poWi5gNRLYNhOo
yAIO0WCbEO/tidruAEInstWHs0G3FUQ6pxD661FZRAqSckipqYg1JPnO08aIQcS3QLfFHtSlmGhN
BY34RMUCjFEI7bGtKlaA6QuNnnoZ+ppGbI00q+887ZYMdwG/iQj0V1WYGkCItefFf46NqiZs7OhM
a3l1IZwsGGFMo7IT5aEA5/6dy6biQhp/JCueSZYs/k/Mzp0yCXBdNRl/6jWflByx8CIvf9zMycsX
VAYKfNJyloDo/HsoYYxG6ibe5+rgHNu4P4O1PXIiITNKpHAHo65O5jSIX9jEuxNlmNV3rJwqLEMc
y8m/ju4w8xLNaO+cgRkSBmaEwT2qjWpqZJh+QlrfZoXhZIZpr8h3EO62c1+4I74MQGhFCjOhaoXH
XG0jrK/UmyNCUsPxS7Q5AZG+omcAuTJy0O33XiwIRmUzcLsi37TzicdyoViAvTIOmnnYlK3HXw8B
FGGKgOnSvGceJf17BXQ1buOT4cSH2eMgBmS+jNZzMVAJZmJWb2lGXajkfl7Y73DgYdZX5rOp88Ar
nD8p6UlxhLd8KqXb2fNwtMt2PqDo0QbLINyvr67X+SayvlOqtYDPCz44FmoUwIatqCeo3qrLpPyi
nX6EYkIg1W67T6zofRlnjEsDq4hjW7iBHwM7PbiYFcocy4JfYDZHMY7v+kBumJqmOjmzKUYJsfp0
u9PHAaV6aqAKRwBckNdl8jkcKAofX5+5HSgroW+TLvah/GnBo0GlvWbvIVrjwXR88juo+w/tH383
blNVjvq4v2bYkQRJiXhY/3nDrrontZ4OMGz9TBoETK3Vnli3ldFJC1dGl04JLlb6yjtsoGxPpCNP
3uAu3CSNrAlhit09Fq2qcbgY5R4/wrmLZ/4nCczhYjDxcMHTOG3jcv7hGd+Vnp+QD47BPQnruRXI
1eAz+PQsxsnJCz6aWc4dm1VGLCNJ4qM6OfU+xAX5uR0XeAXjJaSZiqOs+wLyKbmMji3E4+chiO++
QygTFTwm7L05RtvI5/nAwJB4+iwlynTzYGMjJ39AyhRvSUnHeas+bVBHO8qiFevbIk+y4M8eiZUK
lY9aH4CUl9GorfzlA3CAw2JCRt+QhUgSHI4qZsDVpv4XAh5c/+7YvbFQ2ld/xaJFb/khTjl0HkAi
o31cfRbfUwZYYTdcLYy56QlLldqQlo+nXcnaTPkUa9mDXTQSEntanQH0+ClpKO1TCup7GFGVyIUq
oYV5sdi7APg35+RzaUZFn9ijDNu32IdqwS/kb3SNmF5JcX/OuF7fDnzcP0EvFuXY0BaFPqMAgaeB
jZQxK2HQamCa6YON2PA2r/Wl8ADV0+rFrtFDVgNBdZc53iITMzu6WOZGZ3SLuUUWVBYiVE5WhYPK
rlWdY9YreXQZJUBYmBilUUUpAPK6pwz/cSbZC5xt6VLMNkgtTDm3YT0hpfs4y86Q6cgP67GhVuwb
oPLVvuRupJ+Oyg8oLD1l3f4VNLObnehvJ3g4xTxJoKTg+a7rzacLi3zIAomPH/5bhQ61irth7Z1q
Ir5FirITEh6oY6pMcqzEI6BjOtEsTyaQZv/7vqQXwq+dYE/AsffCQxCotOJbcmv1x+4e7K01VIfQ
BVUQukbRlYjgsUWK34wwnr+KnS1eOT+qGocIkTQPmx8LCRlX9ymHwzGt2E3j0valHPBVxStuD3bm
UtZ1VicsxEedMX+tOuAsw4jNmKnkSwHfM8U+rQeynOUoAATnUPUzh17tM+G7aNtAXMm9wrTDKXfX
1qTnMZ+vfE9FnrmaXR5e/l4mRjtYldoCFcyiFO4AmZv6eTMi0Sxvh0L6tsNjKDCviA9/iITZYkNV
Heh2djldyYcTCG4ym9U0/XmV8DWaT1e2tXuw7dZzQYtc2BtWxq49L9pSvdIeqEapluLGKzVqDeKC
wb9e8lKsttMJTUIEa6nTNq3vYv4cb9iqG4zULFh5UzBgOuy+Y54+ucdtw6sUnRAmx+F2hMw/4wfa
HxIU6fwNHtpR6hF5qw0xLa1IGwy0qrNQBVbCbBH10anMuRVwNTuFxwcpXIW9thkpWeaYVxtg1imA
7etEvQICNQgeVpquHw5W4Qc93m3wf87LkVo/yBpY07a7r7rCjeaS4R8uMqYT8qhxTnnPZm16lCUs
kZCRZqBSp6RKkQf4AIOqTq2CuG4wFcgQxIQEdUPVJjmLOS/0dePTJHtzKdKkXIU1wMM9mykESA3H
nPQZm2EjBxLeDVPHL/ms9X0+D9VL8LnawdxcaJQMl3sRMIen7FaTB2KUXVewp5Z2C35LqCuLfvYE
eVlXUypt+FK8r0jXJopZ082sGtLbVQsliGdkxmJYvjRnLPrXUtp1uAC32bWuD9/POTtBaWs2lJq0
hnOFJJ2cv7bnj4PxgPgFodFKH94kJGe7PQ2iuDkPP6xhZtJKl56G3ZXstLp5SfIuLb+Z4iJMSlPw
sMwqaw/59/nDGQ/tJOF+z0A/2nKQX1M6imWNIjOGGlB7iA7wFRR7ykDGj8SmTBWEpxH7ZvJqxg+f
mWOlDepPjM6hTO+VkQTl7I+VWkD6v7hyt5IkLxs89pSAQ3r62y00u8NAVHQ7wKea/d9dka3EXW2Z
pNKLhMIl0PdESIKJ4XCVnfEPYTpCSjU4ltqhN8gEZrmyU05UaMF6yfby5nr248A/8xL+GzPGi3Hn
BC4HpnicetdRd9yijksD48ZqcLpVjvwIWacKl9CHyhK2O/6Dv7SvfjrwL0RYm4irkIa9TyY4f7nj
mDA8C5c4s0R/gUmInNlDPf7I7AGE/r7mqipzdY/lwql7cuRPgVQ0cqH+jPwxM79elzPydpDXUGld
fNdbBSshc1j+FcWJjxUJIlYGciK2sTazgsCDev0M+fhamanx1MnYlo8aHro2xQcQmMYkFZRZzE1b
BwkJXBm+oaFrzjYvU+Iz0t92I4ZVIiua8SgTAZCQ+DH6HAk86XnxEkp4sEclgqnNnhPraPP2Bdy4
Eh/bzRrv44g0maqOOHFujZBOGASe4YbYv7eFzFBhsM3O3NirsLvsATN57k/IOmwfwMmmGv4lIrlr
tVEbl8JBUNhZnrKKVuCI+B/2wI/utrNSJqy7BKBxZUUhypAW51JU0uBWPPK/vmO1M5V39oeKkisG
lvMl/RWuxdsN88/f0g+83m/Fevv26qGa8C7TMGMTTBSJmV6QeUVkgkmyv9eAAvecplBd1tE7Q8KG
z1mrMedAhFbNnnOLOg22wbNYj6Brzlmqk1kpPYUi0EYQ4YqLDtmdl6cA5JN0GD6yMGtPnZeP2Wvy
Pn+F3ug4GVI5qt68ZB2vsJTx2BSeJTyT3cEBCms0v3mX3BVXimFhXXaES27NbY3OwHZekskm/ayN
V3YUMe6jcgkcFzkk0X8qtYrR36MxGqMm1iRJK4ahf471g2vBhxCB3vAVr7KXs1G81/IMMNsr6GMP
jsCqKddpyXzFy+3O3n7v3K03rQtGXG0xZAhcWcP7V1qySFFL4lRlk9s4vBMgYmQ9p92pQs/xIehy
T4j+RgB2rWxrFmsnLWs12mMTtzB40Kq06lVsaJg9EYZL6gb+5IU/vAYuvT+sOCm6h/XQY+tCmp6f
sI1/JFBHoDeZsDgBTFjtp+bZox/LaAYuzlUDyOFif8O4vIdMNEgkT5cj8ZC0V/GpjH5/oHmlTWJJ
V3lXGgityCJlhiUeeYIDdMDSmeCc+Y91axRwEn4EGS+G0bOWG4HcK/9DKdMrxt6Nos27eCmN3AJa
e4xC5rFHCIsIuWEoD6202X50EDRV/gtIi7BEikeNQAXlDbM269S79r4PDGKWpIsAXjNE2bLcx5pe
1SV29rFqCIP5C3YHIrrkX9SdTdfC6/YveOncxUNiIBFk1b+Xsn8YMuJJvy/MoP4YlHJm38Uyq0HT
nVnnO8IyH0vV2ynMcXKJzEQlsBPnVkrTqZQbk/fWhgaCLS6QNZEvzgpR8/o94wp67ANEkzG8Mk/E
PMH8TUhZvp7WtVsHhyISScT1NGI2UVAkW/xXkIEnjRhftZCya0X3eeVFRxO7BNoGi6t7b8tlfe8f
x7yk5/Bx9Y/X+aT1WyzhCOJmRDiqgIs9wiFddCIT9lOsWmQuTTGhSUKQlHBTbcXrxdO08EoqGTKW
0iS3uxn/NAJr7hE2U1pqcI9d6m9A8HUfx5f3vXaqoQWZAou1Klk8byHL5FIogtJ/s6kqodydUBNi
9G4m1pdY7xspbitz9wPGbKBSBJLViJtmqfRkGGaf7gRIFxOvVOjhhbxbZvulGO0tHvVedjnT/b5h
67tYo0ayavOz7+2bfjpOCvOzQC7YZNcnWhMyam62/ejc1zBr7dE0HEhcIRN9BzBNUT/EZ5XYJOI3
95oK8LybsB1TyJjsE7rd7pA8D70tj1Mrbs88Xz3ef6vifC832y/nRat+3quHnNP5CjV8FTafD9Ab
k4dPNAUPJt4cWbIHsNrbDfdrwigdqMhE+y309Ax/aHDtkhDpX7UNgbBnb6OAuNTufCtOubLcctaS
Ab8RLQl0Housd02gISFvv3oHkn1E7JuoeebEsubFum4EAf7QmCH5/f3kKzG/4GrW5vBoa/vQbqr8
Rp9r0YaP/ogsJHvdMnnUBPKruimCjXCuUA9efDFTKQpf75l3uqv/sZo5lyxx2ToOCBcAY7y3U1wr
nrW+FCtUXG3uBCX3Dl9K1v+oO8TU98N+ogrtt9URg6TaMv/ROZgHTl66Svo7tPl+V9TdUDQ2D6FT
m8SyhLC6uGHX4eImSIzZ0OXOw+dmCYQB6Ja5bJQfvAcVeDEsMOungwQl08RXghUHQYblJ/KCkiNY
vkFRusVXc0RfxHHrixG9E4g846pJSTBkNplNrayjstpTYa8PIw8TTo4XWqnhvBZhN1cJy37uXKLA
/pRyWan0KiuNmWKLFIXHA3MUC9KEuG+AzUSmBMyH7feELiOj0klqyIFz8aQ+NnFWfMnAJxZgSU+w
HFxuBUuZHxO1W7ogyFcrlY/9/XNHwlXqYBR04hyZJMZibnjV26E9NUMO07DbVnhZt4RRgdFYkdNF
x6gR7Be40wjPH3OIyBKVb9CafD9eUmL6+9aBkJSmSmMhsGRemCuMC+82KJr/DdyYuV3Yjrv++KO0
x9KmVicg9eOLVomJ6pZlyYek37XoFOdoUdlzbLFtddZAK5JewUuwa1OEWVWpN7Gmi6csG7smUYfQ
JkbIJh9u8a/hTSt9nwS14dzOcdlqxA+E7H6dSX7LC/2pmUxuD1iJXgZaAOeELL9kRxYAdw7Mt7pM
CL4ZyyQ4pxRY+H1JomLi9c7kAolEnp84Rwlrf08Tx9f8qNIQgWI/VHaA5IW/wzC3Ig58DWIKsMYp
e3E76fJq6WLBF4KhjYpp3ZreLzXjVcL9+QEL4oldmNhK7jtoKQFFh+T/v/DXcI8jGKWSIKo2OX6h
+26T3yvw3iwXREPq+QNTHvqYd1wg+eLZ9bleUBFKy1Cj4iFOZdCQa5SxVV+Vdnau7kKBMf0Kfp3b
gJEljQsmInQ4rHsNgXFZf3tBBxHzDzzsFhhYOQjVsNjL5D2zyJ1bat93dOvurtq9Q0reWPx+4Y+4
YVajQCP1L/7bG2dSCZB1rxz4nM+ERQ6TW0FI3nYsctPCIE13slFN0hIblliv7XdTu1fw6c5YqRYH
kr82Yi+vc31IBdgl9vwK/pibigaHvF57sPWVhbn+PBNXWvHcB8GYH9OT2McKwAyvM078L7VLu51Y
eJb+oOC7yNdrhzAExxD3ThA7qOKPvp72FTXIwrN+UnbWfahofh7akla8gGehoc+WjOOsK4iNgVvg
gKQCc9zlOm0IADBU7YRup7CerQv26NU2wj0BBlkR0Q/i0xhF7M+hxZDfLr2OLzPEe1zD8PV1hXh2
jfuO31jANhihcGfLFJc/kcG0K2HYJ+vHM9JuaJDuoHEipl2xAu4DQ1g8Klc1ZkiU2vlICUe6ZNll
ckhbCCo+S0oMf4uclNiBZxs+qBfpZAFPm57+ZUd8p+q9h3DwkXKzGN92M+VjCQoLVtPsbNAciEd7
HGTZZHyX8xK2Zas8F1b1zYv3jne21zRuqLSfqkw2EGGx6kQZaB587QSDV/JQmyJRXZKTaM775VDe
SxXMKhDdDRdxuj9H3duF3F2hFs1zrh0NY0RNCl1zIQf7d/sJI7L38SvJbBRVvNlFmKr+mGQeGVgp
d9zvotp3aeDsXRYJKKWhzAuZ+YKoGM507DY9uR57lq03VsYW/G4+pUMHwTUQs5iqArGLofApovte
e59tXQV/ezkbpv1w9XyEel4ZyF+zA3k0kke9M8wjOAMD0NOP8aadTZbeCt2J+alOk9B4uYIaroIH
QNMeiztDIoQH0Potl8jvRFq7uliPYKOM+UuLQikc7k6EUeKhVojcTBZ+AZ0wTIp0rPSGpzkggr8Y
Kzy1REtv8ouV7YrdcjCWloIHr9fNjIVc1EF42Rmm+oq4GOG1dVQcilPtXAzkoSg2AYjx2EnYkN0h
8N083bt0FTjuOdripfTeZ76qoauSIaEoogPYgp22BgtW+FwC/FtDMkeViwoAll4136P1vGWm6i5T
4oyeHQjSzaWYCKY8HWDkEZ9XKf24vZnrOIRptmDoWPOQLF7ShzqhF2Os5a05WjwNyYNYcyg2NXZk
Ze5ZlRM8DxUKDdw+F8gzg4wBRoDep5gmaQYllZhyrcqo6Ni9wI3dqEf3wrbhWSfuqe+lOrJATXJ0
DLiFNHYRT1lj/Svw1ZEqwPs4WIsQUeJ6ZcT0+1kWevZnzRrNMxaKUhm5kNsdZ8Gc3WluLBJKRaZ7
Qg7XHJlWEftw6FvF5HMAWR6iambC2EVduXYadlKmNvLxWPZb34aoCM9uzya4XtLX00UyJ67PQB9H
tclW/HYjAtyrqLwoqnqufMj8RQFEyaS2E8Jj1bd1pU8P6pAUYU4BxPPUSjMjdiphLkDfhEAJzJ8L
RlycxT4x9kepMezABltSCZTBOwLLPUCe+eR2ESyOXtDOsekwbHXqzXzsxTd40s8FARvKMp8QCP6M
zxCv0U2D97gB6RABjRl0DtvLcumHhCxbHTkoMk/mq2wshR7LahHxIUFeP0qTEx3dsfCW0dxdvpWT
Xol/shSpcbwp4YsV9kvema8XFHE8INaP2NJvRh9v2avJ2hz86OC7/DbKTi5fqmPIdHyRAbC+KhPr
Sbw6DXlUoh3QkAr/5yBa9ybDTWaFzTaUS4qcddwocUvmTHnh6/NNcOqZeEsOS7eXFmRjx70E9/Q2
vfbyhiue0oYY2jn9M/Hy077+eSYlbKfwTtDaXCfhFMBJHH1mjwjlq5w0wa+BZBAAazdWHOBV46KD
DJML2wTjn2L2+J7V2yzGGgiAUMF5pU8yWaLhOUoNjbS3JHJC3OuhQwcGTO6JKxJWpZm8gMHUBRog
rR33Xvuv9+AFjZLVBYNB9N3S/Fxq24aU6x+eSqj6+VnUeu61gvY7n1QV4AlBSkrGTWBR2DrySCSE
f0eHMyFshqrfCfRI8HITFTRiXnb5Rfk2sDsel9ww4G07TSc0LEQabnnE6PpDDPcQ/jljHzrWh/Dy
uAhZOJMglPUT9QmxtyBJ47u4hNwR/d/VgDkWOhQCbt6++v6tsG5FJvVoRhdiFqnHjQPXKAkR58/y
ImQfQnv/YobC3zzUlvSVXsYzyQCcpdj6kt0V/mOfF72jo6Sngji4cWFCAiQvLMVDHTyfc0qbzbMC
u05k4vFaq/Em+EjbzEYRGoNu+5V/nJHDpKqUUGYBDuDxesI1ruegVmFnCzC1Jscot/VTFoULzDr/
5XPJIXhAF6NnWQZzIzFAus7gtCBJ3GukQhDJPq28+evKQe5uaFMbJi+bruibLKsGYbBkVGMQOli1
FIDn8hUoKuHewGYKrWM3kaooWCepxxgHXpLdvRrDMrKpHtLraL0I3OW/Oh4wYugCLJvgwpksW2/E
tsQD9rFSoFBp5LeAa4O4zV+TmRtN66z2Ku7z4olykpvWovg2FAnvv3HNVQOtceXVu+SoWeaMMFda
Xzj15t8CiQzU3ObUf8QjtTKVYT63XKXZXiHpEEsX+fp6012X0ThHfYBRTz0Gu2/pPAVqEBLHJ1nt
ec4PdgW5ThJ1o4kufmYI1cdo/mJ7It5Vm8mU/weQJKAljEax/jITlur0JdRyonmsaIAU87nR4y+m
7B5IFEByNF4X+MkrHmnOsMrYqe0T6MoEVKmaUrpK2BpGDNZ8Ee+o5sQtfMMJJaGK29M7dBvCwZDG
6kSOldq2OpSN12kL4nNNMbY7mlMe52s2dTpZGrXXKDxenhqVAWO52Pc+6WW79xwlCeQBXeZN7A6O
4xIYRVxyiwK4AdJBJv3HH9up/uZ4aXnyqau7JHkv50axYn2Avi3ji8SmHDYEikbqNxYfwofPyGzk
kPFgKXtVqExQnyDABx884bxET+mOfD9yyMg9rN3Zn9gscytzLXRQCElTYR/PDQ7dnPBCFHYCrg1S
ZvEvuWnxTW5u9DBJcjeJGCAYPrRjC+sTJZu6i+1BmgN75QK0oWFTuG5CZX6TNfl63juYW7xL36ji
oAWys0o+I7969dJuW+25aJmV4vbrekGmqyxAreGkseSUEvmt05b25kKnnupod+SMt3WK5xP9YZLE
U9pX5hLfVJufHb7KMKlpm8dffGwCiwgUWA2qLNMpm0G3f7jth98XJQsy3A9ZI1rSxedzZmB/2EGz
j+ufBq+HJdxMy5A/vKZbmOCpZuyND5ExzLqeu5bHJ5R19ttMHqAyt63rp4kjEg+gEIUAt37/6saM
hs0uD0yN+sJQFl4tl1BC7dFhAof3svvLMfj+g+FXyke06PAfMS4Ws83PSvy0mxDcfqf/uaGpHhh2
5Sk7eZl9WtXMpdkxrxD2w8oN+rx2qok43frW8sQugPXvyWQvRnWFZsxbx+zESegprH1tZePSkLJO
4G4fiz2L4sRKFQlO6Pdp9NgohEf5vZgjwLhvZc1VroP2HuhuX/SUO8G0dJQ3q0CC0Y75bl97T0Lg
mEVJO5jQmreHdTVS+ijjA+HE9NsHVmeMoLe2IQXBOyXvrwd/ky4uMFN/+5El4ZX3Gmob4wpLALyE
tDzC3N1hH0irlZK3VM+OzA+AQADpNOWvKf8Gzvi3ypwEJP5AQmyi8XhUOVnnjFrJruBFdgyYk/82
HUEImtq3NiXwvhgt7xIlMSGmOl5OtoC5CHjB/kBLiaGmGkZUH0/rBNPBSKr4wM0QPf5icHs4fIGG
kfJ7cIUChaUZLvjAs5brgEAADuiieej/D0CA5ENL+XC9aRDBnDTnHJxyo7obvxCTINJJ+eeNWDkh
vvCdNb8gJd3tbqiHVIWz/QJiOQ4PmxxidiFGfA3nF6fxzGLN2/3GFV9ExpxKSG/LHXM+Q0PxSUPg
v5xNvVDoMTFTVPQX6CBbNgWPvOc2o3oTkwDN2T+I6euxxkfOdWjMciRTK4Mf/XfSc8fplJwaCWYw
XU68kBVVYOZM3WyKqB+5veM8+/LL3X3Sa0OHQDsO+OqGMs+zJbz0+yaaGHvE8+VUg3pzcBXIkIb/
MY50ophLSqL68B80suCRf5Cu3w/LG02elNxTgAv24VQzZB4ZYrRdozCqYRDAttBq5xZbRvheHzQv
c77OJcAEz9j/63AIS6labqPPs8iCeJRa7pJzhlStDE0sn90egHRbG+K3nqdiSOKI3F9/pkhUGOeJ
G2HhhV7L1FE1WMd6sl1ZOJSbX/+/h2zEOWskIV+mW2kP0UXZ4A6eD/TXEtnSZ5S6j2c1XkbsdveF
zLhphk1jZ1f5P5SjiB1eeqbLC5YUOqeCiJQ7owjvzRlgCF05UD48X/zAsjzfTR9C2EOH0RZdfy+8
ikxJ69rRKEbiPd8gW9IeqfPjiaOiKSAQnMT0SVFvMOciEpM0I5BOmaDOu4npDP5ehfvf1fTjeJ2a
VZxzaIFvJkV2G6LvkuV0ZopESw0iH70wIf3yz4bLkk/0u2AzfMLSnV8r+5rHhG47sdf3Te43BPV6
mBruCeqRRSWqq3yEW5mZWwL6ntugu+FLZhOg2KWquxFIALdhhPd5qFNPxum5lyGYm42xMpEoPVWJ
3zTcJMbE9E7q9GqKOkDrO1eyq26N2LNprPIMsM3HgP1vhR/c+E9bBfUCDYTz2fZ5GThuOQDgMNbo
HSVszlMW5yd7nq7kkSlbdJ0jnQdjBOlg3O4Q2sQjkORoKJfTbwnLv4wfb7+/FoSBO5LMcHXur5uE
nbtgK8cHE5ZQq/ZNzw9urogP7YpGDfwbTHACLLKudVURhGkSf4plqvX+y5ir4RPWohnHmuhvDKn0
Q/v4XAB0pJsfh4EMY2J74Qn0hCId3vo8LNAwtQRUOHwb0tGNoLPkvofiM63m8ykJv7KJIz0dV9dj
R8hFvsWy2LLkWFwvPKNkKIFy15HjDMXc7ExjVzVhecIdbt9XIx3p84F4lYatIaZbkNfupJSA4Jw3
IPpflBZbpgyw039W/GPcsJVH4+6dznyMLZs3CtDr0axBdKSUNPXTwViyBM8Irky32hsdCzcseHNA
BXDqteJv+reKCzo2BhX8LNZV8WSiU2MyzBC/mZmTOKRJPGZUtnNsXJrY0NC40qYGMY2jYfXxt/Sy
CfA0+Y4clAykT4EsxRnnBNnspQgb5v/hXdZ4BqJbkDV6y7AM/ShzZ3RD3KMbQKdhxOOmfDfsdIrt
bAyZIQPSboDh1jqQe+onjfpw5iZnnsfQP78I1QXk4mQn4OGFf0U89LtWj44IPQxMRL+tvwyqEayO
K1vSzBaIcbsy1PLSbS+NTH2jTyCV3ScOHVC60opLUNZs5PTjRmATxOU2pNgwPMvnpSwL9/8Y41dT
g+0rAfF8RSXoS9SslzTZB9BBL7mcQEcpCA5Vn3gIBT9X1E735+5rGaUlDUi+Cy3CfNTNguyG4rti
GPFF48SGUx4GN1zeOhZFEgzDuzciqKtSyniaFTOYOAkzstofN0AHexoT5CXhuA/4VZyJ/oAfYjrx
G9TohTvCId7KfvSZ+eukUWJikihbQLdg5VHz+Z4FeO5NBMSr8eOCEebKwDxUo2VA8q5wdVvEkler
PknW3oHvi59aG4yQe3xIrTdXoIbcGpun5/C8ltEbzrcQ6fhmT5iNdku820O0Ti+s7uwJTP/wDBo9
PpYK5TjZawu6qh5DnLe0bfQDjheczOZjCnegAVn7xkHQtph+0AfoIfI7EC25oZUntUrvRLDw94Ph
UQox7YtXYDnxBjRrHAkcuvUV0MoJ3tn35fZvFkjncAa6tq/AniRq3ieQNSu5++uRZywfulXHvs0o
plV0Fwu+D5MJjXULrAjhzk80ovkb4vPF6JsmvD99aS8fDk2wnM/mLNPgcP7tJBlM7nnb2Dte3N4N
HTjYJJnI2u9iVRFj90+ug/pjPqZHhNk3drhLkt6YNq75RXl4Nr9idgN2A3ggfl9AMDSqK+yeuZNX
95kYNnCJQubHKtnz4QvoriQww0PQFGQxbUoBdpRUbSW+8oEALnHBoBe4Jeh196hIYfEw/zTn4D4n
q7FOu1KEjgGU0JbIar6UXp4+8oj0SA62CTeK+6yK3rKQHKqL0H0ddjEF6Vz8uXCDWe3VG9nZgqCN
NqUMBU+DTmQGdaWGeYXSPmcwtKr/ACFZQCne/tFcNaPLBfSI6/5dUzGA0p5t50pp00JHAP1kSvXa
iib11rs/bzHetdmucTa2E8f0wNA7ChW8g6p5TrYD5tZT3nF1r+gA1JC70UYVlbHMe8+pEVWDgpo7
LWov8nDyNfOSYLurxqDJBdZYPP1a0tKVB9YB9gZk6rTWrOqd9tuv8Lu8GMIGQKHOAkbBjf8I4sMc
mSaS5QGLXfSA+jIZe2mA9g6x9lTYd7f1aQJVx+PsWYDsII4smB4CQrQnfzlDoM8GBXDBxHANdBbJ
nTMJqjtrAH/Nvv2WvEersrC3Odc48Y5E5vE/ymeUWe3HVoMT12Pu6KO1tY8Vn6HuPQNrAyimbfQB
KWVGXbOVtliWFtoVjiSbGiw+PSCwHRJ9HYE7/TScPYFQGluw1g5AH3b1+mP3ozv07MIWzU1JPf4b
e4VchO4MmnTFJx4DDQeHXPJp4MjKW/awKu/qVRlnWoUJU4v7eRvWjBGWufP7dwmhjUUzEaij0X8f
OBETjD6684aJJ8beiYbznAYBGhj+VYeICHZWkeIciMEBa3e4C0iwx6sRuhaCandkZaYKtB3d6IUD
rGe71mz5ITg8SKa8yCzBPeczNxfHqO47ry+Fu/qoCziyzWUd6D5u68Uxr4ROUjSO/Ods6D/lE2T6
rgKnf8n/HdYqsIeqbqsYXe5FSayyhbBNgDdI9tifeZewI3BcH59AeePCxJPNyJh4vy4261Z2fXBz
7jJtodkubRU9huPCp2LbeZO7hm/QdTMgrw8ViNWKHhF/jF/YrXBcDfORhkO9jhuI5vYU9CX0ywMg
ZxRdlbNO19EK4xoYsx9nOToxAh0Vse3cchEul8azc+hsVLqYa+lP+1OcbBCilxeUHnTbCTj7M2DK
U1Hw1QTq4rrVhx0ZsOVojKRi7+GaB1hgpi7Y6aPCL0ikkloOrmTatBW7vnR0m0uGbMAfFGMpz5H8
DUVYYljvsSpqIpx/VRYI9vd7wTjj+St4Vra5etFAllFGFk8teu3opP+vu/jqK/Cxx8ktEBaz7J5L
oMriyPUsOvsTZbr/shCSTIAmh0ZiQJM5GgG6rLJFQmmljcpIHapBKpQ2EmffuIo4whjYT+my+lHP
C8C8fa9Qq+GboTSVY4ljwmg1t+ytVMmWarsIp1BzQaF12DpwdJSJoEcU37Qf7xzzoi4ZNT1N69yh
vQb6fFqBJR+hgHIb/Z0JPA2pr5xe20rPmVN+plweLfrbjh5SfARPUW0apZAmEE613cSSJUkinJ0N
0uv9vtueixVhj0KFqJ82rxk7ssjad8lasSyv7KX/Q65fVJ/7e0ZtDWOWJ5sqW9GJOqRmdv9CcZjD
HksicDpxyvycDw21bDe+e4Kh6tp/AQ8XbE7+390H/7FJcvqJF1jvIe1dZVi4pZbb/FH4RgEbVAXM
FeXybDLqAC693LxNBdqh+jsf/5N0FfJ5uzT8BSjGgUoP53b2yQsKEfjATqNMfDD8TXsWKeyhd7uR
k3l7mLkWkDxDqHYEwdu5HiqO54xHXt9VkNcQh+6o3FN+p4Qw2ypY/dro9jzm9WQ7eopLlm04cOwO
dN+JBfjE+OzAx4e+MVggW6tRiFIqr2o0zhjdagKh+3D/HtKLhMesvQoUa224VntmuvMb5pdR3JOz
BEL+/+U9K6gpoR5wqj1zUTguUOEKodG/5wloFunsv3WE2TiUU3sUenkNEJ5pEgIFUc58LHwri+Yw
ufIxdyl5Rhfq4DgfzJMwIn2Q3Ud/T5/udwGhOYR/Ny529cUgbHW7ufIJ4e1QL4//qucIPrM92+yk
oa3G9W9AQKmOLbLc/udw2wdvIkohERLw61gxBkjPlvIaSzAOnsLMSsYrggpenAiOflCwspjmCFBZ
+WmIr4zoMy4NpiBAQqTmAkvub+w9uQMK4HbRjywIeXrTDlmfNL5xwFXqixRmMJcu5H/NRm8bOLWv
XtQqcgHnczAgUt7vQWp3VR7eu+REcvXOHA6psSFDZjvqlQHxsA3PnQu9g8fzmcQIu73hRLZXMOpv
YHCimMQ0s2N18ZVH1HJyMLwot0VbFWc99dY0LKNyAtA6HBDIPnodkOqP3MELvI1NYW/WIL4R3E4u
BZiLZxaFJEUXfSm+i8/QYtWR12k66RBx6ktuANkH1klDz8voIRWOCx09vaBcqN/sWln6QVRyg2SJ
77xZ1h4eZUvxLaS1X1EgS4sKgY1bXV82vBlMrY1jZGzYdbrGBhduypvvJ8kwqIL40+U8Bjd7XRrm
9gPIEkt3CiNRCwqsX50PLc+ayOmPW0ebQ6INLA9+pgsU70zhzPnVG6ckXMKOyhasS7alR8PqS8q3
Nujqk0iT42asDna/Z5rJgJsPSmJ/0sITWQieKHUN460T9Dfy+2t68bLapEk34Mq69TzAMXGTF0n9
1+LQ9CePZ888Ka6SIFQUw8opA9EnP01+lwrk8j6h5IP4PXxQo/ARKCsZ2rDS5Fa/BvNrCHFAvxhu
H7GTy8Hk2zYW+CfSYtTsim1Y5G5AQbKJHHvHaJw6GS1Xj2mNu/uC2OE/SJg2Z5cSqmLR2H8r46J2
Lfnr9o3x7OqF6QAVDsNAghk4/k4SDyI6wE/3rWuDsX/fmpcrK3g7J8wa92RMKXLyfqbYMRRsngzh
HhjPFI2E0vuhKJ9uI/YXM3V+XxstzLqWXY1gFZuimd39aR/FgqbFbX80354edK/m9S2nbN6RDTwz
DGo15aM+ULNA4T/dzAD5M77KHlqSrSWLYddi56aL8Nh5riyigLudS40oREFPk+MqnKPnw2DkVlDN
hJLPfHiBwqy3NUB28hjYqiLKw4dK5DRh7rN4iBi94ncn3KNK/pnfvV2HoovSWE7dSfSJgTGz5oW7
9+3ZBB+2oPr9t7blqI7jfnOWCBl3NxsmIcOtTAVXWjVARAlMcWxq7XFOHCJRr3eU6ofzOp2hv94m
/5mDTY9nMqHY69GzDI1K/Iz0xdMmWfnHGDClJbOjim+zRxXsD9S0gM6HYkrZCMmHRvPWjkjneIBh
DDfUIse969iO56RJfVlFNyFl0owIRhBlGztp6yXG4ruG88kadV6b+vE+PBr0dFvsar794o2y+qe3
nYhDRF3alhHesdUDilhrEBVtC71wk97bIIZhXD1Ru7DgzvJifr2sMWv3dY5jiKyt7NMEUzgp4I7V
JR3QOaUPBC5ecKlom9InP/96gQwab1JL+TEnJFqJM3uJuVRIpxHBKhWE+HJnSwKPHwt1VyY477yl
FJAzf8/Ocz71XIRaynFx/zW9pVCGtSpdmTQtidt60pitLt9Q7yRid9Mi/DdAqh2+gB72yT9tKQ2n
9guq6Tgh4DaGSkOg3kbphjigN1LJOdDQjvLASppJzieCwCVk6LDjOlLAIQv3RWjGHNvRAveep1L0
LMpel63V850nJ5ERRD6Zmk06NFITXworovCcMSNljqjNAXx7yRXrcaf78bZULedHl0Ad2gFjLL4k
Q12z4rcYjFRgfAxu9NxL3CmaIJwn2/SKpeMiuTWPjbThOCNU+mwIhsu1RIPmSk9h12U8JhYUzrDU
Ye1QzStwD5nP6dpyGqHaNyMUH5fStIOm3nwRxN0UO17/IoDaOW7kZzWSh8/315yyIHbxqLv+xg/a
3rTWFUldTXUjMT1NrJfuffIJXiyJDAaM9bQ0e4F/fNSFplDEUbqui8z7c2Qu8JqCW0dtwR1RY5s3
FH7Yhjeqff9iUG1vcHESgVoOgIIcwJMNGu/2F3pFrU2k4yPLb7elyhZTotxrA/A+6AgDegrqTXGe
JSEBStO/HiA6zVRZfU31Qhdy7Ofh6VUBzpt9USf3wFM2DZHZHFWnjwqOBW+RLWRcpkuqclVmiUEB
irsVcekxoWKNRPapMFDpyWzq+TdApuJwZoKfIZiR2RFVrI7Q7M5U9S6aIxGe3m52hbeu+4spRnTl
l1eEkNlWlXgeibB7L4rs40XVQVI+mG73LnSK356o7SKaMk6383bvvu7hapYkRFBOCN1aNktT/8fw
V4PeYIZncB6yJk5WLkRgZlbhLLgtQshH9a5PRf+wU7fsea54S8UKShgSt39DzS7o/yuO72FjFyH4
mzpTuzj8vdJzB+nCeV9jo91F2ItgX8dPXQ3VcSKJVhVSUTFNYAZJ2LaAART1zOUlI2w9FHoegYze
X/M2d52aWeHXxf0s22MDRKIZmzPnWjEJCxHTmUAy7YQfDslAYD4Y4FQrTUHebhQ9pv4i5miBGt3a
kdfOzrklJbsHModzdqblKrLDQwuqK563saM1Dhd80KT/MDNQJiNjLTtocJcAGKR27NYIAOBvbaF3
j1s9QSshGoanJRLMETsAgnV0fVo2TplKysA+TmdmMP0oc38h9u8/17rJyhxWG5+BtJzfimnn3+vP
37UhJXseHoRChtCwoIASLzHcTAOgIHikMV3proj1iOhui1wujb7BFqE0GdimbqGECcHENfQwBNHA
TN36xn2dqpEyy0T5dXYynkEP9DasjzKBjINoBzMC7wcxWPoYgGgrFDrl7kpZqK505yMZ0vawTnWl
R9qgtLis+t4nRiF1PNyVeid8J4mqT9P2Vc5J1dL8o9XixLMQvOTegd7aDnSuIX4OZOkuTl4ST229
uBx/TeO7DMOpJqeI8elYdlo9SGlhbD0nKu8fffGUut4tUSkh7KB1M9va/ENfNlx6tn7jOY3arzRJ
kNBtbyoUNxH/8jppNEOyHuP79OyeRSegfv0ZhecwjMrGTFIXJIZIeIki0rwvB5I8vJILYsHrNTnV
rooTJl17h9zDNBx2aBAInPfQWalCRmICU3f1KSAm0IIXm2CO77Hrla6c3uJYnSMZzskVjwiJ1kWG
a7FJ+ptZWAJ7dy1pgM6nwqaYb22xxAl44iSiS36bCxLd2Y7hJ9Gx5idCZ+0xQMPzj0AKM9LzYRz2
TsY+//xJK0VWHbkPVRsyiLW1/PNVBaprb/PmCzoChzcKm11MeomeUVIqDzD3WWNGhxdqnGvATZCN
/zqo9TVX4Fv8tatfcoYXEnpmVfLDfwKQDixyQUj10fnqwI6y6A6pFzI/mZtFRpM6b936MAFqBrBS
XKom2Shrgy3B/MFFpCU/VeeZAM4jxDc6Q2063ZxMGohgNN7HJMc2pR3SEQxfdDsDPJ9yAp8wHJCY
7NkjrNFRsUKn5rWihiz2zTaBsXP/fkzOA7ZMMVdg4utk4ZFpc9r3Jhd255npCtfMtG5Rn5V2J+8/
A589e94DTvBb6TXa9xtM4BWCY31g1cv+/U3XXeYasjQfp1fWXBihE0nr5hIiM63CpRNMZ+5kJ347
52ko7JzLkQ/evOjnxQ/SEl6yM7pAAf2mGe2CXAMq2emdBZ3BayFx1ytFR7CD5UPxELi1Wi9hZmO0
zUZzlvosKWACIfAl/ISFJsR/pF+mZsIan97mcEDKaSAStkZGW1a2U4yg//p2RYjXnK9aKJFf4b8O
xGftj96FLjMdAKw/IrNfTrkyOfCzSDZVWHM2Ab2ki7TG+7vI6ImSFw1BY8ciC5sXS4IVE2uyEfTB
0wd/ffqDh3vzaawFO5y8Zc4teqntFGktHtg6x2zu8MkGNQVJZA5BOPRFsPU21rAFEHZNxDwAV6/X
P8TOIahR4ClTYmkDbxCO4r8StdQcqfP81+wbLIneuR+brvtuB2U8p321XgqCXvEKaNmOLx7C+HKC
HojeKnEjpSZulRheD+ARUnp9yr2a+SIVjDY/9BJPfMuPsIMr9upf42xOU71zEBWlHxcINuUdW1CG
hiMVwrmFwYAbZL3aOdhu82A8ae61Gg08zETe/XkVSDmeKCv8l4AU8/bKbzThZjFZh5C1UsK4SRnQ
xb/YrqEAtaYD2u+PVRtkrzLZgiKBVDIOODIEgo5HLjneSQ2Vm6RsF3Cc/3F27HlcEvv3CoQKYUKB
ACXUazFd28/YoQjK/bEpUm5OzVXkNObeERLsNPmDUysS9eF/nHDiDXLX/jbfqyhZg/7Yp2MLaP3N
QMVhIzleypbSW/tCTMDHw/Cf9vN+FYw5u1VgiVEe1PMX5H4xL/zT6OXO6Y6RwHJFpeYhERCYKSee
CHG8t7wqxh3ACqP9pGFYLbHG1vkQDiCEuBLdBdeKUUvyetE4qqNl0g0obEZ6s3MJHX4+HUIxHBX6
iAZeHblYbFfftOy/v8aj5kBA2bQakLmvWYZ4J2WzEBTJMtSz8Vz+7ZNNbMNGm3Mb+3HwNbc8+OPU
yQJpyLIFBCHPYl0oKB3yozHYDxNgkS+YOAscFRcUWqRomk7ODvotw/I7k/mVHayx1O0+QC8+mA4h
f2nRqMgrUnRk3nzMIbICFUmNcWl1IkT9PhRlZ5T8fdp886haIdFC+SwA8RUxaxFJPZK2VT0P+F67
qK7GvbhIJWNCRZsOqRwvJ4FBLafkrM0isHJC0k3hYhZuPz1nGP9D4g2T7iaNQ5o0GhSY20Jd7T9H
5UYNhmcxbnKYfPg2tGNZbYYpITIoj8y3Wk8MwAypYtSP6kK4zi4epi/O2Mw5HFVpdHJMFXEznz0g
w0SEyVbjZGva7L0TpCxxhM82wT0qOqFRcvsx1OYO9tERHsAD6Dr/k6yR6MgmWPnYOCM/OkIQ04Dg
dVCd58ZQOmbjLXqEH/NtezqH9SGCnBi2YAxdfbI9EXNmpAwI1Lrbr/CXnINaO6gQvAB0TKSV/bDl
c/n9WFReRdJ7iZ5NQL7fSxQhjpzuHP1ramhUY6Tk+NqQoY8ROi6XF2Vmr8HFPrJhyIJ669gz/MGB
tkKiVFR93aN+UsFY4MBO9tXmpT+yn+vQQqdskZdCfIsSZRaxXXZUIMvG5HSqYYOqGIis1gCunfVR
k7R20Aor0HK63qeFPzWNDuQ/r6F1daixjGJJjl2e6mUTmLqcLsR3FpHbdui+sdkbz0MYFNM/a4xu
u+w1wD9VJYYan3MYGT3Vwyz/TqXhFjsIpLQ9nPPAp2NCZ8X054fspI7PLrzh081tFdJ32cRTMSZT
wtNLHMK2B5B5811wH/rVY0AZ6IHyT0ZP4LreJeWGefZY1loFZc3iYZ5UiX2YBjOf3VXSKCwk+bzY
6QlD+Z8XJNhMd1mSHI6/waXxPO018VJF8fox5IkAbLALYcRgDNUb0VOvr+ICf4Zb6QYeBddpx6AS
DO8+Ud34sYOQdLvF7e+ZB1Rio7OFfkYYYpmacUxM4szzF4V/qB7APhDypyUMv1jImSCMVTO3ErxD
0M0ACKhgxu81AMfGRMFgaUWHRytShQwxnfrnigk1+QVJ/oigm+CoF2UWnJYZQfMb4YDmaAkU/KES
9RpuK2cABrux2sQSOR5cRzJvBVoFkajQh4jd7GKIdxM8cvaQJ+leV/aFAajlmSZUXqp+yvXOHh96
DrWaq/5RktUVyzZwkqvm+wZxwSp4vW3DK7uT9f9uNEbrjYzLr4BRnGmrmF7nt9kEsuBxWq/q5P1l
HWHGQ/HA+BOUEdom8OsaJiejToiqDBaIrhm+yrftVksF0cvHtMFDxqyZvjLfRVfzb4s6qqNzqbh9
N+FTVcLJIygnXKzfm/uSQWue4vVXpSh9krBbZVHjJzpK/zxg/cwBg+A1K3XWyNcuYA03JnXQQjTi
FZaU4BMKnyufWIF/hDiLsqnzcMQiBxFwidSl+Xp+TNEYoyLYbpkGlDkN5ZJ1a9qjxLDpuYXsgQ3R
bGMCmXvUYYacAZkiG5EPx+Uod4cHVSBWyrfPwpWS3sBQpzVCsTqq5fJDLLAi21WwoYJ44Y6146tn
ylADRNdXRgE5+TZfgQNy+qf/ejbYFcXmX9XxYfNmcJ3qrLUebbjB5vJklofy7Wkg3GSuzgDN/qXC
rfleswE9wBbYFZCImn+1jTcIy8ytSlOkHteI4/bofQsBgj8JgZqiMGwwqS8htNoFfaR0QgNYRNPB
X9KCWeufeutq1TSpi3HuH04RFNm+ZM9KSc9u3qTltXH0ANN1s39NQ+J+3hL0xcC56Wu1G1SrpjBv
81DhhvGa/4iwQH9Pkj72hSHe5NQYvIQN2UEC6DlAdF9naglCgBaMjYfeWRB9F5Ti0BzNzJlnstwn
kKxnK2NiPQJl77CscoqFMOu+SKSxvnXLhOIGMsZz1lQNU31ULOnb2VVX/2sWFRDxfDJK5TzP8tHu
MxlICSbNehg1kTSJHktgsS3MLomOVoKxxMouzLqr7quLBo3XybtFVhSlsYjhvsfd0DM3Ja9IQohL
TL2S128z1JKf9rZFhr/LvV+htnEkzDcxoM+Bhk1QfCZ2f1Dl5jePOfcu5d7g9mb6xtqIKyKG/LK3
fC4lT/W841faPs/3bxIcT96gXQrOm+7Kz5XaVSSFgJT6KysYV9VqhDMF5vZ1TsTmBLmrf0+zSDSq
FRtwCT0bN6vuV7AvNJS+1wFpjJws+gCJfJ8xpjh+/LPTza1l87anYmgyqq7cpmhzHq7ZO2l/20Ph
/nQt3Mbr5Fn7fVG7AJ53bo4pmPnOgv7JGOm94B0n7S3RzVq8glZfu4c3scThcftnssRlgBJ4wCWu
AeehUm4jCzbhW/pvKIECaOsZfgw69bMfZmx7W5zn9N5vlaXTa1UTFNsHyWXEoDh+lGQSAgWRQXUm
Mncvg6leEeFz8E1h2Z1bU5gnW043LH0dNioiBGupXngaOGilP0CqP0NGJtm5t97P0ODq6eKSAIEl
l72pGrFPpOafKcbjQVMHJlskxKdJmnCB+BvzqPCEuZ5tcUCb7zh+LQY1gzSSa+50StT3IjjoudZJ
O63prBqOERst98m035JQDlLGsGtOePwddVDFQfCKZxI4hRyGswCtIP+gSPWFaVBXhWsX3cIVt/1X
SgGE+wQGEgf9LjgSYijg9lQGuk0z6fX0icQEUeQdMRiOLk/omwJqCsyjEbYYiCdENciGtQklFQhi
LTCncm96MLaKfMO/Lw/7OtajtpqFq8aWonVMLpw/W9LdPfFLO9x/rb3n7V0eJKSB1IVrkT8n7Sur
KfAPuxynlwS3NUcOEo6LzkUt49rrN5nvPV+ZU4Z+kMlpNnPXZLGZeND0q6C93/vhbHZxIUQWAafa
6crJQ/yeX+G5Rks3N3HCkeANaJom9gDimHhdgXHYcBfO+S2pZo/4IeSl0GOJX58+UffR/oECm4N+
mj2thr9mieVDSLAUbIn/g/75SNGdlMyU200BRf0Ec1Mk94z+n7MirzwN9SI7HVoVFNVEnCpGqywN
VWA+gdH1TbG19flhDhhq5yBgq2WkWjLRy1+4lrcRyWrSHwXWPMg859QWC/oE9XEbDlkPExQ1GFAQ
xWzTnE8XmrJA/KurdZiLV8sbPB2/B0Kzyl0ztPV8A48JFVtb0xftpCwjS0MrsTfJJN2u0H5hk++w
HPf3yq8xswv6TnUHUPiGg80leaKTNdqTSOLN1cQUnNHcV4Da9zNjkArLztIHssbkbebH5DeuInZU
s0a/IxmZUs5RqNkb6WvbexEgN83vA3Q7owb5Slw421GsvIjyvuSidUf5mxTrhTvoi6J7+ad+rj79
7+vfpwk867/c5Pf8B9U3mMGBOxWeCYDgGiLfl5El98CilRj33ur2uzUbNTAu2A+aGT08EDSTOmQQ
EYJjB86XoFMVGYzfwV41ejUguZcZcY+eA4WyvRUdn1vrP3+2BW56xX4/UZQaK5rDnGrFJZ7Y1vqY
4bcB76nxGTQAO0VlWHd4wvRHTJW8OfoFlFvlcZaC/PMoloCsMEcu30IQZoaVDexUzdBGBVYfQ+Jz
p2fGj/8kIdnioALgZ9e3CN/kNr9ZHhMUA7wviHE5sPZQqu3/UcdlJZgN8kYeB33MUK/jHiSsSkHn
HmWFKpVZ46jyt1auI58p+cnI/m7bnzGoR9meEVJNiBmcGoDkSjBZOJCMqsRkDu37F68O5c6eZQjS
rN6lcoSihEaGfVbC3TC+BIOCbYr823WTT1+GhJ7cEDk7BM6ewgKBIecuGsw3VOfr2hBEltDUJwcv
GfDJO6fEuJ4tSoWzMOUwScIm8RMoVUKLMsnABChssxcQppzXVViJU+dvYndWPjTjSJT+loQ3AI5P
aprkcngd9egt2UwvT+gPeSRx3ZyPGgtf4EJMa8koA4g0AeWiVsTASctDTEns3kyI6Np1p/Maqli+
woCtkD4IT7swSY611MUwUfDeeE1+5aWPOk8qy04BAqQn+Eo+Yzj47eL9kiB69prCOGJv0l1TU5nz
an+77PW28f0JGCAq3n3cypKEhOFZgRzHf4swkCqVzXSx2c7M6HFFXa4zT74hUXDSk1JJaS73AG3D
RBEZAaA+v7/g2Lf7OZKecLDgOcCKNmFq3HlgsW4Hdfxkf/Tc1pRA3mHwrRJlHsSg+YOg1WcxW0GJ
WGwMV9GgJxuWx1GDzFUDdxnECepYBSdMaY1QsuWnkpowxe9BhtTL3FKrqmOSn5QTdFVxitLx5/AJ
6WxVX6bynBsymAcaED8WBxX2KpEK51KfOmGpDsX9xhn1b1FhxDSL6Wq8RNRrebUCvx0VRcnIe50n
Q87HD7CW3s6CdB5u8GAxki0lpsa9XMljE6Ew56FhmDypPnebSvZj9GbrMep0qQELib1zxP3nlbPg
wIQi8hGeGmi999N0vl1hwMsf96oF6bFf2EvVvXI029tDXyiH7MvB/UzTpqQgWMhiUXnXfeVh99a7
XD3PoyD4jh3tZMnRFn3MZz0sS0WCrO2CBj8elSMLfyYvH3EtoMbH4AjQtiwbFnTayxGPVJ15g2gm
doVztnKgpFEyUe1NmA6OltD3Huawj43GAU8PK4czMEyBYzTF265+empzN2Uv7G+DaYenBTtjrroJ
BKcSVMj2Pp+VHRme+dit4rM3/3wVohaTLqE378VFgghJn7iOfoF5KvSbJDGzd6hhWxDmZbI3qNYj
MH3C2YS2iSE93nvosrxhVL+It3v5umyfyCHQsi0/+53ZV9vxpi0kc80+V7R3WmAWknswQgM3q8Wz
QCvd6HwiYhV7qzTo6h94gsJmHvs1AgA3vhh4vHhRyeqASAomDeVXlFy3peKILkZ27DYDziZ1sVU0
bxXOd5ps4cDr8daNc1jUTmzim8bjAd4snirD01yISOa/4K5w9zPNf0eGLJsdRMIZZkQyYoUjyuN8
IARCzynHx1+SghnbEMzyxyptup/VgTTUv+RbSGtdNmKepADVvMv/JfouVN9+MZ38ZPtDB0ngz54z
R0gxRs0Uz9JuaGnW0tifm5WBo8KmmISKPSxShWKwZDqCSDZojxns05vZWhe4cmD2QHkhbrKqu7+n
Lj7nRoxRLRPbjyq4vLTR9sqw2BSkAzAJmw1N8AeyKLbn9wxSswVwCAb9jl8YlCBciSaF3Wa8NWHI
SO2yxnkNb1QG4g+SqgT/4byygVPuyDZqYq5rWuzxp7MpBnV/EqQLZu3iGg4zsPkth2sS/EO691dg
FcttMIcmDW+PV7gWe5wFEehR7qQsd3XiBozPQinViLmEEjACaOeSu+Qjh6qGM0JlGlIdFraPgAmj
wGoCMqbiRlhLOuEsJaBjvmqbut8IOESk+7xuWj0gT/pYkZKUXceo8s4T24Yggl8GVnqkXgtK2E9l
TUlZn/QEAiQ3an+7NFBGQ0kLXwZgFSeaUbG6C8EymdOaET82tHYaYQfeh4bNgrDgSsj7sc88ejGE
wAuoE3KHMD/Yp5VeMrtrtFkYVQuY4ByOhtf3mRb/iSUZrMcKYreHXtYGnviAcPkeD9Bg0o9OGxhb
1pvyCQJiOo30vOP2PFUC16dStsiTPW4lhN61rtfGtIWb8WYW3FnVtPU1rjcVp1gANv+DpxtSHd1p
NOr9+qvexlxUe0bm9QqBWa/rwFguH1auEO+0AXnZZxAc+Giw3fjxR8Ja8ZuuJoCEwyq8yluTVh17
u1jwuJow/ay2JepmFArtiGueFNrhNjrP358wwoVY00qm/it6YzODxyU7LFBd2XwVEdCiQc4QBnZl
W+hYn5ANXUiGJ82CN2qUXQA/s4jb0j1YAfn7CiMlmwHbzlLoco4p2mFJSSeGpELjCQwBnqm0042g
uOC+gQm+mooE7/bsU6P5kamRRX1ycpEaryIloElC/v4Lymi3bB96AgPLlPbxAytOjV2cxET5CyEj
+IVir6XZraeIcCNIC6XCRHd/uIID9OH0fB1+2V6TmcEMJm5t5AzyHxhaAQjtJWud1Ge8j7Jlis53
AHz3ag/tqPnrGO70QH7VTJx2+ta+W+NFtSWR8lYc6DsruT8kCu3Aq8Mr6BFNdzOUifizcqZ6qb11
ua+v3Wc3DAJ9cDQsHDzPtei2ra+ene+hxQVXPU6RwDl31/xyb6vtr1aWum04tA2FfaGP7xAdpUrO
fW1qXpYHNP6VD/O4d7o6BG8BRO8yDpFGe9iR72P0K7MB4GpIKbVLwiJw2l8+CckvtGTfNN4lWGUt
F2oEgi+6Bw1aLDpATjSYs/jlZzIQ9p6860qNDNyhZrd+2u0c3olGuYNjW7mqMuUaqCe005ZftJa/
gnTSiwogOJtJXjhYHc+tk/WTeQJtQEMfo7+bH05uo0aQug9vAwvHnwmD3iWMprMKmHzbA2W+7u6G
A8oVrn62KZiy9JQx6HzDWjfys1aaD7cppuYFTJqewQOk50SfYBl4J8JQigMSdYpeM2O6Aze/5EAs
dDfzV2hu76xcMnNoeaCpl1uq1qLmlEXTyCklXI8z2LQHlkQ3bsYcu5AYv4zZPTuqEQnxbDYDyAEa
2Oo8I7j+vs551nD4ddF6OsWLe9eOb9eYf8JV2rglnesJ+ZjMMYtcEPGLGcYTUet7dLCjum7bqPyX
BxTTFpjW29EMLc6a3+js2+jx5pY/t8GPHa9iAKGvwzjmjrzN8wzZe2i/xglX8F0DA2UDa9phi2iw
AxFeU9q099furluYHYu3vVCOvDnjOUSe70llUduKa2+J2tRyrqCWH90EAAjICqp21ZpYt1UnBdLq
WJK56htxo1PR4g+n0jeA2vFLFD3c6YSZyxkdP5ozW6T5Jwj0xWZ8ZIHYuinSDuVtiyGNJNyFZO/h
4IH5Xar9s83P7gKDYVm11P5yMl0qVvBa0O9UJopRf9I73bCabOWa9SEtrcAmgGJkvmqjedUJwE72
2O0+QodV/n8c+i1RKwhwP06Q0AiblSPSQyIvxEfTyxTD8XmuQHEGHEnoZ0eIWdMXMEr6toHCSVlP
lz9aMTs3un4SmI4VPeDHznyJR/QMq2Xljmf8VMu+r/agpnikguwcxDQdMyXtqIjcN4C0rv9CHXqm
zztyPPdt/qwHsfqkiRJ7IpSiOsdjmBU/zRsp2Ey0CKdxkoDqNLAlS5uEJHpF3+ocON9KjsMvNRe4
xlolaWKvl0O6VhZo17Yn894oDNUw7Ag5gsL6BsC50wxZfU4ESKDCxSmMUomsc94r4u2ugfk6rBtk
2WijzTe2McNLwi7UX5RttA7rKaxkZ8hNfCcyTyye6tEs9KueYzB+VPVP9c2LuQVHkI/zNT436mFI
LKGESFmj7G1QN4QPLjJmlzGMH0P39xoSoX4dkL/eOlYLN1Je5mxU7U5Y8c6138eN3AOpvW1BDdT0
ZHI6UQZon/qqK9G7gS3lpeNHCVFsPXgBe/qw2f45fca7MJRY1wQmqAl/fyyCVtwpHhzGCHRi7htQ
ZbefcuApB8ylBAcNGlPnx748SHJTWomEM0ZQW9FEwSa+tc7/0pb15mYjrHVaWltfBZN2qDHKQFOB
coR0y8ageQy8WT0WoPlk9Kw+3XXuS7vIF4xaDpDLyTEDLIQiMduhEEQPFyUJ5wk690bcwUsloSU2
9pQgMw57hgae3beSIYbxhH0ZDasAGaaeKth3MDYfM9C+tzBLqQW6aEEeN5lcH0MxTne7F6JMi+WJ
Vj8aKb1DW3Ayy34ovkh7DyhfMWRfP8Cibo1qglRidUdXOCr0RpwTkqHIbmAMYeUqGNW98s2TOJCa
Vmk6/D+qMuTVPfPWzQTy8/+S1+KqJE2q9y7H3T2oEXHvbOVGoUnQpCpR6sw+rhtZOt4NVilfAO7l
6PyYbfepl31Q0HnB+ZLQzOhkIiSB+GzB+sJT7efb/UFIrvunqHOseohJZq7ZYEwqNJYKsKV0lxX4
ByIl+jQr4nR7AG/HfPJem9FWadUsBIqaLnRdPheLKV1MsDVUuxy2UxOJXY7dczzMOcDUZ1JGNgcf
Wv2LS1cB3w1QcJjeEJjW/y5bMjDTzkiwSmUf35nz3AyaudNO5FGAu2hffTVd3GsyKfWJbwjT2Em0
EqQscoz+JdZ+gJeVm6ewoRLGsJLORlb6Jr83FRMS0RqMG8V8RRPpeM3TashNRNBPx44quiM44mDm
SGfMPbRGj2SMvlD/1lw1Z0Db6Hg8dGpGGFA7/tRhcghJmA+g5jMUPOSspjRpp8cQFLtS0sriUDlX
4oDfJWM3WzV99TtDYc0/2Wj4mxghXlei96YDM4QiNNPXqNuymHDHQlTExx2+GYpZrPkRV51P4wpQ
+JeZFqyEMCUM5dIz2YQi2ZDxQR+7w7CqW/gs8jmsRolzr1ewBhMkJ/zhNA51SJNL5p4eZD4szo9M
8ibJj2VlUDFuMPD13TOPCRoichTVuAh9hnUnJcY+Dv594VsvyQL6cBA+/mRohHFLD4QOvWyu3n+N
Qpzu/kOiSKl9NUeXYHT2VHVKkekm9gm6A7Y34S+324xkZ1dM4O+X3H8tVc36LcyGkSejK+rljXn0
aT4R5JHR+11gYiyENWm5DMFxunpo3GGNE4tA5GwR8vAgfEMwlm9rI6fvKl6ny6hUldkZxpiTQ8lh
YnXBBy//VTr378tBpVsyegP3MZopUhGYRhEOJxpH6dM+gP18RHHbslo6hSemsbT2+vDkAIdsE1ZX
kx+NwRXhjBOfnRCsDavRPqR+D9s62AX4PtI29dSm0AEt/jaq1QsHVz3fFsgiQti1/QqTWQBNEyNG
udmalIr08rZtyfmPZgMdFMhxg77VwIMApN6rUwsAVmzFDhDcqk5Sy+wLnADr5BLE3b+71yxUgMze
4e99Cs6FDQmMHYSd+GgvdXnny2CcLUuMoqTZhTs0XdN5QGpQlZFdlufOoo1EuIW+si7g/qMBGmxA
qJZmNvAw6/ELMYxdFPLxf/UBcPaEgwvvuDOsqEtMcDFL4MvHYEaXHGccuYdoAcjx/jaKXNNN18Dz
9bX8x+EzUrcb1RAnPa8YroEbPnBjPzo7GK5AefDJ25QfTPsii3poIoHEXzs1JoYNlrrT1KknE2Ei
cB/gnerwEZqAIa4YZ84NylMO5Em+bEHbalOLasnBkOPuQ/4Ayqu43Hr6X8lfljemxrvkq3IwxQ9F
XfVAVDDrbacINrs5X6+oBkbrnwONYbtnoX8m9ZyJmxWQZ+WJ9+FdnxYbwFegBENWFaJRvfYcrdkE
vM9c5MvMVFOG9Vh/5gjoJUsQJTQCn3qABTkXijgNl9HEy/gQqsTLSRCkBc8b5HCeRMWl2//IWjzZ
h2+7Ee+7uZfTyyCM1qppli1SMiwSpUGXRHlIVr2KBMg1sCkTFF6Zvwy7qXWJh/vb7g6oZexOMxTK
sXt9S5aCreDA85+dIQE8HBaDUl3eHYHBv4sBGn2/83HGCoQAYMhDVchId68nqpDLw0RmuHqLUIBk
3YZ1OfxpzbOsF9ZIeMnymPIGOWonFD+zNL0go9EaLdRG0BvAPDn/kX3LhS6/71ERmiB4cwMD9paM
s8sV4uyJHPqimNZXr80xHTuCIOsj0e3m+ZaiT92I0itK7IjArDJkLkxUpP8x9Utv1u5lP3EW9snf
2qA/OH6E8Xh0ZtxfU/L4BSR+5bIATB8rdAqxa0hKDfIPVpWJQamcylWGGQBbpmppMWX5mmhT5d5G
3FO1abOGW9MUjR27HmsCOsG7YOXiMLMHz1IztbYrpkG0zhyBxGQQ3qmBTGvShax0mOtkcwp7DA4J
O5nMJXL4lcph9pRawHe9Nm2KjVNqIvSan+K4puN2ZqLE2YeuYJO2ckqudn6p/yXHBoe+d4j1dwNM
XcJGGr3D4cm0pn8IWO12QB6pBn8fZpwvsecWzVEz623wgxqxaRMUiOO4PgK9cPeU3bfPVmZPWBdw
fOoDL/qFaAnbHyjT579yfcXZ319NXW3++mbBg3+sgJ353esL8m6BvL0w1hESkpZOop4MZViE/NJc
Gd655tIPWxBQKtT1z44+aYysEDD1GVA/PUx2WPXZCFumvfkPdnbUCOO/PnLW/x4dKzW7ktm5x1ry
aq1WiSsT9QspDc2EZgmI9tazR5Cl7BYUsBQdY3Iyu7lw50leIwQSGK0dB+fmoeDEaCDJePVi6aEV
cnbO6/p99zYsWyed770KgD9Di/CPd362anevMtdym4w9ruGY21Tu7jc+PQMIAKjI4iTfhkMPOMGL
iWz3WbKIfnW+MJMtpKjMtEce9dGURJATXkScK5UDuDx5d94p1ROIrziph2hkdRAsTKfpbwDzJBbB
PUAyGLuRqhoU9FLHXFDhsufLVCLH1uWX69c0U395HArpZP+8pTl85wLHAVyzOa5n0kuKanu0aIZi
6hs+5Pr/kwYq8xZAbTE30NPUx0Q8K+bmd+A0RiMSt1GDwhaWT/P/vInP7yn4RjHbiepbW6OYdFvd
v4HFghdP6zkwuC9gZwlJWf3Iqqq2Vi3js3dRt7M+zz69LEvJEg2b860zKDP2W31SwG20MI4c3NxF
ZY8C6yGW63g8cFnm418HsgUC2hu0oWGbOOE4k6+ZVy/BhQZCb/pmfejb3epDvORfhltvh23a5bOd
M1OETCWWcLrikljRoGvTPVuL+mHPCJCybUXyJrGHU4IU3dZjtv/5lRrSfJlFybKGKm1Whm9Kuj8K
ji+Q6ewPe777qWyZOUDEDB/DYcmUMg3psxWCUeu5ZhnhMPrDNPLxDQ8wp6C0qOH+Gla+gC/EL/Bj
6iDtb/MJKvNVl5lhsWK50JlLupepKDAsD+FQ43h0h8nrkRptGSUkVQ6tzgUsodFZ8bwV0n7gKLxr
IVd5PIQQS0VxcHDUDQ61j+CNqA5lcEuOTTfHHJIVw+PtIEoD6/TfAgnQgBPn9yzMl1lIbJGPHD75
V/LDVMov2VBDYYzkXBb/oRxXik6KzDD9Hiu346xF3E6Q9YkbArwx/RKkF+x3mShcfpVt49EhuarY
YL8LTBoqDiTkG8LrVRu5uiqs4nmKawLhshq60gePHnawB5JYD6jiJNXNgaJx7xM33RdlX8q5I/3W
n+Da0gClR1bD9QWod22jT8AjFzX9WEVouMRWMFKlyVmU+ocDBPJqbINCNXLNw9a3gtfxasTLd25B
lu2LAmUWTs6nnX6CkUVELfPtIhk3nV3PTt8P2eMasjVRvc5sxnF2HNcgbXjudJwRn1FSHLmhXM1r
Ke9Pb/DDMxdIG0Hi7VktOEOIiBClmpTiyugu4LpNuNpm29VmCkUVuGSc4xtZQNB+8SZqaMU3r/Vs
vhS2yaq9qYpoda2m8qqHxFDJbOkVoMUf/BXueWV8u4eUXFQek0OOB5Au7RNBBBlXcYg/V8p8G4SO
dsG4an1puvkaUy0s4+xe9iYZoBhSFBbfzyW1MnjxluvNwvZERGWeUVgKc4aSdht68vpCrjMbLVcO
MpG2BF7R77pA3f++t9xGf78GVJx7gG4wm9NGpnZCcOIblrZ1+V6o4IOyacMN5/O5OLpWxEjhgeEA
hvjAvlcHST2hg2h+z0q5feW8QqFNJBq7otXOBuUXHQsH4cQ1u+t7R/4eCsHO2n8KnCYkliAMx17O
1gM7txJczA4ymXeILHu5kxM0T69TWEvfvD+Dg1kCJ6cK/dCiQ7JvTt7c2sctddbgkL8SqTWKyTly
AFyKgEDLTkMe8BaeV8H2ipTEikH39xOgj3atKr/L/1hXfRtumhrkLBBxReYC6jPjAGZeKiiHo7Hr
yqvppeAS0J9jrLi3aTO/wGPmDDi3b0mFC/tKfO0U3MGaErj6LazYwyjMzMTAHpegZUDYqZIIs+DN
d3Uc5O65KTbO4RoS2k05vvX47aRSxgIGz4IAC0MfOrPQtQ7OBJ3kPEBdFLu2+cMs4rAfRcg1OKe6
KVPnYMqOopzhRAfilhJR9IWkPoJUm46Nwhr5O9h0AusMoD3Nmr5kC3zq99nnl+TozogJlmG+o/eE
dL5xl9XvgId/QCRCtgyZYPCWuUV0PnVV+SogxiJd5mKl+mtszwKem6zegoyRKjU2PJjfvagWuMVe
uQrCTk1sM1Dks2NS/4aZcWJJO0HlvT30sbPnz0xF43ZevciBR1HZmjEOnTSivRkrow4yZyYX4Wja
Hf/6yHWdWQd27uRRyKV9suYtNiyfflSgLQjFQ0Ioe/6jKCaMRoZkSW7YFsIxy5N/Mi02zdjnH3Ej
VCaN4nqiKtEY8nRdjgFKHapIowTRINO2nsIUaHvXLBlkCKkBrmeJ4MmOAmWZq7GR5xTJ/fQkOMax
HQaWwM9/X0ArkZX8uAGfM00jn2ctkr1V343S7UkOHNNAX6ABl+S5JyuRc3Y02bDiuQs4drZcmqlz
DKS+PddYCQ1M5BKsWDqOsP8A8GNQn6bHOUOA6+27DFcJKWZ9mi2OyrHwa24jaQaSNBY0TAuVKUa3
wIaEBPc8+C/HkOiTSNSCrTJZPglK9wW4B1aclOEoMZoMs0z7TFDRYhLu1kCBIWScps0C3Yax9lUq
OBpuIY9RSEyFO24LdWs3pkGkyx5TK8LtMm7o8FplyhXNXcub2GKo+FFpw9b9kzOSO727/O+DanUj
oDDMawBmw70h83EGSayn2cjWxE6pbTZdzBm8mTKebVXzC7LlVGCHSuA46opO2y6+3fQaHoTBer5S
UWXMppcJ10CuEPsTNaXNsGKwqOcSF5Z1SVuqDvQO8AGWhP5RPJsFro1Ea700EZfcq2zU6OEafOec
7aipfW8abz0wCXyWylRR5edFam7J42zLBbAbloNYiEr5BOxrEC84gGtdpwe1QZVdgxvLmZU4wpme
ZWm8hjIRLGF957rbrSdD9/Wm3LHWu4VksTo4ptl148xLlOB2RAV3dsE/w8e4Nks/ub5Autm4BS4g
c8I18PdCyst2fBnkHq5FPLkhT3awQsui+aII3I3RAlf0lYgZmgQbM05uTUr47ISqAG2lf11Wt565
MsggeJ8Sns7OkUIco1yZXzebTfyZqOh8a3DnjBL+tWLH/WKylSfgBjNY4n3OTqdmeSSrsaNBi7MB
GAaxUskBPtV71oIE+TUKJ06om1DTmivheU+tOI8evMbMWqHjKIkCvbjUfXU49MyLxDiJDeNnTupj
joOQ1KDDobQEUb2z0StddMHE2lB0WtyjW046Lfg0UtnH/5G88qQT9FKXW/S/KzsGNqrA98l3d3Wk
HnljiBf2/ZVLsth+UlAe+S4CYjTTHOWDwHIbBH0jNB0bhpAsIYvu/9NpR5ud5P/Idi3TaSQsB9r5
E9pAd0WvYbsVUC1yAHS1s7zEL8jYcRcmtvNtAZB3mG5P9CL1j6HPAwF+BaAXhACZKQEfWBLr0ZEZ
Nb4Dib1M044H63aj9faImNsjrtLZ5XwdQfj9sT78Epo/mAbCkX7afx3TyPgj0wnR9HZ7Ukw7Qhdq
YANuuJeuTbbFF3CtA3K/JB1ziSRqyT5Lndb5wPzVhQRpFFkvU2sIov2ZSSRephVrUKbL/xHs7Vk0
kQPH916glJk8zaTaWzXLhuGSpMMXew0lexMQ4sIMJvn/ph9ljAmXOIQ+N5JPjrnV8OTHruiCO3ER
Hhfb+vLEfiqnsT0C27H0MnaQfCXvn5syR6ZUUIemWDo5VzyWDlqBMa60u6m+CkHl5l5s/Xxagb+G
t1Zi/Hz2Ibkn5/I0gmXHu9TE2K08Po0WNXr29eXF+kWVz+nPKvMCpSxE8HlI1fnXgNYKXF0fZaTK
GCOFYwJOhnGZGvjSGDMr7e0M7W4ba3C1htnxzDtyNAOJJvnUiHNcbvECKuHYj3ti8xZNhn5rRyvQ
vwmpER25n+Mk1by+haNeILSERpUdXYwsuev+wyZowc6Dahr1eXxB8vE5E7xj34RWyWkdfyMotS5D
elu7AIB326h2JV8Af+tQ0bcmkieZr0eHsjSIc+6AtO3dlfqFme9HO+ORP7iA16mUzueLsJr4GEyE
7DWKMO7QDVt/xkumi34Sbzx803LJ0T5bFu948KhMKVq/LCcrk+y5wkbgsY2RsWV7I65jFyr+I2Ca
anpIYQXhc/6SxiNjn4C1JxPTMk/79qzJMdXkyVrfOXf6Obx5UZXDExSRen91/zkDmNlsOr2nJ73e
2xz+UrbPYja3uuVlV1LOra3Z0szJ9F0Ks9DYSt4r95s+z9chPtHYKotJy0vc3bY16cgMazufQUc/
sj/tqB70o8fT1xwJLGl2toN8zg878LoJy2wdmcZ6Tr4zK5CUFJA6wpMr/6J7uIz3qLYUXW8Re76u
4N75n3uUTDZJZ7AlNSE/6phoxGyLVd637nw1SNJT/koJTr8EqorFDoiVdxN5IKse04shdjk6DYOr
9nxXb2L7gkwB1tImKjuc9NvwmtdPr4q4F+cBjATN6oJ++hCNVdRDER7rXZ/DtVe63QlSqid25Okx
YZgykd3tf95mUh27/K1bQlgN28UMWVLgUKWPU0fbsRT6NHRczYrl6GgFQotaIFdMi1QYL/aYHuWZ
gyQcsYvlRijvz7QX2cXy/dyBaIaTzrYDsPNUh/N1IiUofOGkQ8r4Kr/XEvQtI20z7ZW+m3ReBFW+
g7P1FCZJakiOP1aBACIQgfhU7PPjp5Upv4iFma/4oxORhwyrFNpLT9FbI4xQG2aMTCrHaq6FFenL
tcEJliY19n8/x8LSw69pXXzbYQbRtLEwRtwkuROn6Lr47DAzw9futhXBYFBlTD8jxJrd81Y8LS/V
+haT4gALYRDjeXfap3yIMbWiRNJi2QubP9gwOdwmWNBeBmAc7G41z+og3Pd86NjHa3QcUxh/Gg57
vENNcFkCQYZQjO9emd7WPMT1d3lo1OXyFMxBVMzZGxPC4YvMAXPxUmegYzCVYqqDJCZiZOD8Lw7A
WxPUIlykQV39YfOAY354M/C3Sm+Mw3eT9Ed+e+3uGeDbbfLMN3FenhQeBCC5zr2tKJBm457qkQ5a
W7jSAJ6PvCGRY69YQ2lRMsnOzT4k6n0SySBju7oMD6AN4TJ1FlKMzdeWVGTfbBISxPa94/VVqWF4
uXmLEqrl+KalakhjLuVfYfHb1NEwiP+xAKsvwXsuijHaiYzf+HzN0nrKGDqNBAEF5FZmscJ5xBvq
JwaYxiBo6Bk8XY01qzioXyOSNsTB+PbeHtbq/8niXpdazC4U2eC60sOOPqVrkPcSr/SkiX3VwPAI
LNuM9nph1qG+tyQGv5WUfY6lS4nnhhWx4NZre/ZiEW6ARXQqxy47JzNA+d/8pJo2raPqq2JJX/ZK
WzRIqbIMkMJQsbnhqISdD8/76Hn6OCNMGrJEUSGd9PlR6MFlIksY9JFgJE26QQgDr3ogQlnHhL24
L10hGf0RGOHYXiW8iI/jh+CX8N6DRQEYasN3PBAgpBv2UDb0SbvAYCEY6SewEGRrq+wIAQdGQjHd
nulrYW8DM2NA+JWB29WoaboxLfG9TJHpvepJWZzwjQsI6oPvcLxQKdwEn7RpN4UEis7Y7XC9KI1N
PBU8Yq+urxhvJVnk+XFG3qQClR3pqXmg7tRe95ggfbzK95HXsGT4mHhFGyKuwSO1/AWhBafQ+Nus
NEQPE99F1C7X5Br8z3sheiaIiiIrCakoec1H3GGgYOOuqogxMUUH00xbymyX3BJ1bt7RWwkOt25Z
EAb72ba0/15gpdS72xSYefefxzoAzpho8ABml7ZYlOYg+EWGpvVNG8qTuQGEEiKxI25q0YXPf3yq
/L5ivBxUr8nGSehjaBTSgpSLuer1PvOaCyottQIyWM/WFRLOWegtBJ3IaCOK+WiXj8UeDpf/17Z4
IfDuqi+XbOaz5z7qQjbiAEwmDZpNurSlKqEIbxE3QL0wiXGQD50Rk7Zyx5KgdODrpzY0ezY8JRB4
94OWe9cVtd9YWFPRYKAXpKX/L5oE6Tr4M5T7fSZJg1a9/U1iqd7D6RXFqDEUJnrhsOgpTUAGe4wC
F1kZ/usd2UKfQ47PYx01MuogaSaefUsAxvSJC4wKv4B5CApEEQ6PePPhKHWlAk/E/dC0QguSz9hx
NS0YkotPui6rY5eZSy4fDHjUthoSvCvhgvHXlawCdBHrUAcI+VSBy8fQTtpc4YcMcF37mUrTFk4c
nk5qdQrVsW/r+dH8j9EqF4nwbNbUAfDJ27qWLm9VFkQWM5YqyHPf6wIuI4iJaFR+FGFIW3sTZeuS
romB03TgomuiwoIGSYAx3cwlxKY/d+mWE11CTSWNKtef4h8wdwRYY83V7X7R6nk4C6JTS0d5OfOa
gApQl/QqlPLs6fyHXl9WHFu7dh575fbkpLJ8+3OwIjLTFJK1FYpCUckFnCfkUtLxD4EqTojwkjUw
ZihPqof/Iq+rXmgY1OcyKn5KL+MrRorIWHlmWy62mxIbicqZvbDecBkK2quZm1lIUmup9gWIa1Ya
wm6i23zUEgN6lWtXRfHLZ9bsCI+Fi2SS4BHhJ0DyxO6NPskObeNr6Ttm1ee1cNbwcbnr0hqgUn1e
tT6W6/RS5ih20hOV/jy8tUAe2ZYCWP6FmMuaJ2+uPAiufDuq3IxQ35+E36IK9myOKySjyixj4rF8
WoqED80/xRSNIhqT4h6RZssTh7/DcV5h8GutzpoXU0xpl8HYS5f2BDPiFti6fGnpRQzbXaEgUKdo
caTtHoq5ZZmV11yZPx6bKl+uvEgr+MxuD5xCGKxIq68R9KdXII0+GQvdJT8W88oh9/4/dsZUxK+Q
Bmrg/KwPobLnJtbqI/bvabndqVZuKpjhDmP5tZei+6iHwT7RCJO2bnPoYFanLjzsdFs+Xn2GjpOf
rY+nrlZd3UD6UvYQTTcsmafAlLUWb7ETgBH66zXJh8pNV4+Hz5ElNktV1B4Unn74cDap8nJORsx9
jpthYY7ngdRvBi9x2KYEInSPikWEkMtVmg7UWVTwJvvAfnhce2VxiJFJ2wNEvCsrm6kyxF9TGePt
hQghnBdsmN7XjcsssEm7dG0wdUjCF46u5Xr8dWwbW96b1NEeV8wPPVSWO/sWK9NEQ8c2Cjp55LUA
wjFbc2pOW+6UeH1OI6vctI3jJX8Ke0f4MPsdZJc4l+xJfe4Zp2jiuBefrlJmB53m+tzTpZ5196Ub
nVkhpDxSeJzxfAzqmlovSsAoa99owtiyXSgGUgSFez+vbAPwFGBHUjxMpddzjItDqE0RU+M6GBEW
F0alom0AE7s8yNk/10qNZSmu/jPJ4VLue3R9ryC5KizZO+RBYi+6sayzNy7zp3YCjDMR6JOwWF+4
HEO2/baK9V7POJAk8LTqr+aZcewN9M/RxQJSJk1gdreo9IXhHHA9YCCLhJnLqViQJ/H8GsMi/7/6
AllwK7Hkp2uDkqsd4AxHHLL4VE5Pwtzn4oxzDU3e4LtSletXANyRXGvIPnwX6n2NYf3ukt5IbDlI
NtSNOFg9p4lTyV0+9DC4BwXA6Kh4sdz4fKaxg3Fat7Mre8U0a8VuQ/+kvGM+hO0G5FV13u21702k
pKtlnUcVhf737XOXF32HT/Pi4WDMJz3h5YkRbOMtaPoxjayV3PqbvkI/Lm6hOukEJ1wO6KMbQhLT
nJ1QgGEmkiiwGaE6Z44lx2mFmJRyhnbTPVyXvYPIEHRHE5EpDomUmYeg1RTfmR9O54uiL0mcM4/0
jnmrczSewFdYNLgBNBrteuBexiZHNng+7Z0fdSuH/uS6Lg9nuW/Ci6FFYI+MtvZE4QFbLpaDeqgN
JoN1xcU39VejjbaWNKB6RMnKizL+5CvI+UPWEqXMu1sBe3rNrYXr2qQ2KYPCrzK4ePkfr+4RmrCG
8WiPrFQO7XL6xz6IL47EZY54sOnViRefucG824E6rh5lGja9IC/2t+Ah9gPVHBo4wd1qwv5KRYoT
H7Z5eKGjm+SYX8LRmITrfzMwQY5fNY1Vj1q71MCrqDaQ1Usbo8AJg07yDVocGMWeAJpixH6Z9A+U
AOSd+xh1+3/xchB857WdTqjCxyM3lwjyS9tDBI5OxgWgISQD8Ie/E4drlmamYisI0taMnvtOyPPi
JPiLBi55srKn0M058VT67NjOle/aHG3fZtDT2JV3mHBt+gozX9mpQ/HxcEaHSWjvC+4cDgb2cmDF
44wQTAyakl+cfvmLZxRCC9+rnfJPBJu05e3xtY63ajHR+Zh4bujYjiBD4LG1JBldHZhauOawFb+W
2Z7fb5TFDMCrMazkBkztLdpT0dPL8AWz54G53+bbktnTuZToUgdya11kx6pcMmV0NUiQGGsz9e6z
1lhGdxOroRaPC5CwjzMN0vV/hgnoq4Nv4vnwlAeeg6Doq5LiFv/257GblZpB+r2hyH+1p6fAa0vi
q6LST9SMEJn5d0Sb1cYLF1dJ5WceH33SdYBdkVgQjnJK+jcHjClWo+luN5VzLDygxFvcYXIBtugX
HzLMmSrPraSlMZJOetodTedSFeghCWn6abkW94mjfWa2WW9IS65R/72c8U+W6fFQDmI4fU0p33m9
Pw2oFLPcKzhQWiJpRRHlYe0HAgQ/w7d6h1FjFrCugtG48LDfIQpZtmQ6olNRDf+bLb4/7L/vAmYN
Jq2xcXbaxwikXP/7Rr8D65GXXZFdqLoLFMlUk9v8MvGLB54IWv6IJ5COsiRIzj6fJ20uH/YBBfi8
zQWPyw0gdEqAkSqHLdBD9hyXzQJkMCotfGtCWPWayWs3CPanDJAM7UV+0EuVerDXA4UQXoICIzvz
Duz1R8nIRf3Xg/AwuXLEm81J6LY6bH2HCgCRS1CCRvBL2771upZvwruCKcwTN6W6REhtxLsSWY8f
uod/KjihrFkUdK5Xe3BN0g1pWl34aCSoYgo8JOtEyYJWBTDWsVz6NvOpbY2NtLvW04ieYkSBD6cM
lQKUndaybcJrX42g9OmTxWE4wGgEkFQ3rZ16Cp1MITwcsV03NF0jo7CVRXXtBS+yRTZUUdmz5gCd
UygaDoqYy+K/1JLqMSPKbvM61H1BCtRqqypCNePA8+nofB2OenODmCJqU8kNwMrNrx3ev9f55dUZ
e1wc5ze0ENgbSOSSPC9kPyZeh9bsHF2uz3KC6T02XU3C0730L2hpMlcxP6wJDzBuUfkzMUazfSYd
SLDj9yATmsXbTijhZZNaB+cghXmzcVm0VQgFHjAiWexM59F0eYvWFE+MdV4JGmHzvt7mt/dPwcZH
M57Oz0UDlVaTb4kOOxWUewduWxICevfPR1yBTFJWdgWlPfVXGqsHsPG8KsoAKRZv7zv4FCG4m3Qj
+yx/ED5VnUjV5T2J0GLHtnZDzplxWJ+BgLih7ISynGsc7Y6vMaZpbghT5XuVCsFHBRagQD6OxMnf
ulhV6VD8sEMq9m1PW0mFZTaeLtKoXEFs5Xtwpagf+L/W2BjR0u43Nof0nhHQqeemc3KQzvvy98T6
JgD7iRH6g9RZJAR2voGlJi/nRWkMlllOxLC376D8bwwJEauSD62tL0kk/Zk89s9EIB1WBCieN/hd
3qpefW9rDMmkz2wkQ0V13ANnQuwbtkSVQxyq3nfH3V56bRkKUuNi9HcdFBEDDonRjYZz6pGje5M0
oBIQEqUXZMOfCTlC6JY3DSmB/wj5PsIQ2pON9sbZPXPsRo3CQqDGnrfq8IBWMV5/2Au/7FYD6XSH
B7kZuxsGIv0c3OaHjSzGY1Tnr72mUG1acXIdeFk7cNd9dDNLoM2irdQl/uzER8RPV/Pv+HTcGPgw
TXJ23bU/snETbtmgHRLO4EAoETCXAJsxb5G0uWukNH4IGIZoJclStJugDqwmXa0dKVj+U9gJgY80
EIk4kFA9aLgsuSEbLS4KKVQrY44eLw3rHZbNRRBVlgS3DuCQEOEuxxAIyy2GkoTkAj4hPNsJy7H4
dIED5B6nH9u1dVp7UqleV7hXFr7IzTiPt4CmtY6ttcNHNjkG6e5/j3iqGmxrmY93Va5JXNj5Fdl2
yRSD0ARhBXVChydDyt/PcppOUb58UBmvH4gdF5LbSpSME5B3SKr3M7mm0Y6XuJYVO8AhbJXavPYG
44iUk889jUTbZpr5nHP0IAP9r7FrViay7sB/0jcWrhj9Yc472yR03DR/mOh3F4dwREb+hpvZpkBZ
gwVdXRL/QEejfyJoZewZRGT9dmpXr58ixtGGeqQBDFkDlFtXe83+3JiFbCl3hEx7/xGsV5Z/VOb9
M4mdjBOm1Tl3nwo20ZxMNBSm0PZ1BHgWp3TAaOKO5scMYTvfAjq59Fe2kphMMRuQ3GIpw6InX/3E
ve3mteJqeviPvwzT7Han7F5NUoqMRWbhpRq4BkTs/XIaC+eD8+zulU1gE1ubonKHBFpAVrYCt50J
gc1lX+pLcxT4Bfutvbbc4PvS863xmbLCS5k2KD4gCG6zDB7Bn7mGqKjEQFp2N+IA5fOpwrwM1GvH
SX0nfts18bxU3vngRlSWMSMUKW9kFdjGOpCANDiuGI3OAJbWuYCKvuNjhcCIcFz8Zo9cEPTlNaaQ
q+1WKy2GFBxSIRzrITs43Uok1EpcY3gR5e+CfTdWxUp5EMh/6JI981z6qZwjPjgyGoMK+LrutHBS
tWLPJfOGe8jdp20FhkzgbkdkvcLtmaanQGMCb2DSNEziRXiZN5o5gTZ+FPkerYFLeVwqubvCz4hz
log32lk7G8z88pUyyJaap8dBhLXHEAv5UDSLpqYsFKs3zwqF2jrsTssmIwj0FBzr9q4swiZ1FKl4
pWP8YQjsPttyxPmtb5083TS84la63QmfDYuTIdkm4Jwebqo2lN1wW8Np7/DDUmj7N0BM726OEVbw
G6q1DwN7Sspl6EoYBuFsCABlcc0Sbyku0PRGjMvp1eOvIsdOU0jxpAHw4HfkFzH50JbITx584KVM
v+P0Wf6JzGZAkR60asI81xV6WAEFFsG/GKHwniDTktz3ZD823FNajefSyeALywnTeAt2lnsnq2CI
5ar7+mda8Rkx/OKWZnjEu/gygg+ZrejclVqH/cPim3fb4bygHevtCElIm9g8mARxkxIYmV2UTpd6
cFzVpf6UtVol/GHOXxU4ZSf488SkxaeGfMbaxlBGipMw4zqgPlH1OrrgU4ybUgImsdS1WIIHzANk
mypERez9jLef1pPA2iHsrCSF/vVm51Jb8VcV7u5uV02i7agvvkyn4U9iNQ2blSoZBKLo0NfhpwLE
NI77zQ4k3RKvyXP9bXXBlI6HQ7dU3jd2sXTYwbmrIjZT0HGQwZymMI3prJEMgbRcA/oo4TAy70YN
1SEQV9CxYeoLQmGeZjzFKbY38+esp1DVhoVDaXdRp/eCTUgS82cjFKbO0m6KNgU2YhYofyzjzwIf
tD3b3RPiz30TUfyDKillPC9Gxtkk16722pyx8X4hP7Rm27C4b9IL2c9GAY7OOhKjmNxSJMCXcRen
EV6nhzUDi+KBBlUVsD8yEVpMl5efssLloqIdHiGXoBPLcuQIZA8NT1KMH6S8MZDBn/tMlGrOPyPY
iiVNzakhVu/OPRbdQ/P10ypUa1SxstcP5jLAKVSfNUYZuT30d1Z8j85hHI3pUrJ87zmHWwKRbDJp
tOpxxjF0uZhkAKATdE/qQ+kfd8XD7DLS5Dik+azthCHvLjAeQkAa3PkygUgp4A7yz5MRcAfr3myL
oUIIw0q4b3YDT8SkPfIE6CZ46AoaRAUj+MH1ZPo4Idoj1+k1o1lLSEDIfuNnPbbjgRHGuwNUoYVr
7AMAecB4m0wM3l2E5VC+W96Vcx3m9xaq4hRvQRQ3qmSwhBWtBJPyVTCczUd3dL5buCh2CNLa4La6
qQ08z3KwpjLj+OeT0CUuFFojj1H7ej6x+KGwaAeN8swqB43WbWLC+WMmFUpjgF1AxTF5xXqrKsAu
j53H9rEDPP4WTkg56pMlKGtNWnsFoAYjyI00d0jqN3K3hRrokdUgWzlWWYUkGLyQzRCxT7UIIx48
f3VjmMEPTPC+S1AhckUH+s69tUdN1Z71PgU6sPncW9qWFKMbc6BO+jcQzm+zKxhCpCq2y20F6ldM
foe3OOM0gJirzoXCcJnOGoIwRMmt2MbawjMdaQlIFw9I5XnPLpZl3Oc0kjGwACFvXo2xfmtpvVtS
Kt95Pb8t3lzqMO5PJRGTFV1lq0ygyuATELv5UtC3H342AG1vV2ocUv7uuYV3smePhRWxkiZoNM0R
LU8QL2fwjERgZqVHZeWwMxCQXAHNSR8Cn/zcdc1Zq8Wi7/oKyHH3xHEEM5mlzzaJO6+QmcBprH2y
2W1wxCAv4VQtBdMGEsxV+kL4K0FReSERMr0Gn7ifFmpvFxyXoh7lJrVuWy5LPkUI6YDykIFq23zs
ap6uY/i6FvBGODcIEwmYm29HJrZ3nMuo/YVLEhJefOUHPbgovEM3buFKLOjHolBHdpG6sMUUMXad
KxKJ2FRsl1J6BPfKoHLibLp+mFT/Ktt907JzDdB01i7+roROE28EAoUrJu2dIvoni7YVk1ipiLdj
n/lFR4M2tlywAfRPGBAu1NWv6kC6QhLc0ft4LIDia7JnGIz7BlQoX4dVhX7rXh3ZwH2LBaX/IFFV
87jAqilwlLOMlXU1kOUyqwsWfaYaJlXogs1zi0CW2aeOLdliyyqXcyKirBDGCADwiK94ehek2fDr
T5egwKgzB87WSDXUwuZOrqG2FyExm32RsQo6HrywS0SSE0Uu+a2aV/UKyVmr0EpnQli5GSoTPaHr
H15rOr3RrrBQBq0Xncac1HsZJV18b2Y0jI+y3zvK6F6c81pR34acgT8hbjs7iR6QYp7DXTt5RrJn
LLSj3TWqN3JM8HnWVUp2KLG9gp0opAXnAnebglwiJ/w+N+dx3e74BFK87ak6uWSl6/9lkcPCZSLo
E2XcbmDfHxXsp1ou+YOXtVeC82ZgxezDwCNIoVtZ8LUtx4g4JWlAxU6HaaDmvwjzQOggNFTvpbs5
Kp3AlMgkv83mjEozZlBVxXe34ao6Wi6v10D0frmJ8ISruk1SCT1/gGSoHM0ZhrorOG16QGtXlZIB
cPwOlVHIKSHb9sPSAxrLDSKuSJfQYFEbQwM4fjNAHST1F/oHyG9hq7WkydtA0BU1SQ5Ww6kK1AKC
DoxcQfAoL5ds3KpcqBcf7kUZo6VtJ+poBBFIFEKCx45szBh+f44GFCewSwmulQ85t4SQN5Bp1U9L
fVFFiVtvHNms27WuJCEL+tJJi82Sf0qRzZLtF9TG0VfH86GbTYQygu+dexRK2ifjodTWTPEFGztm
ckD4uL8AGkDQqheX0ewZYuD1biSZu58hCI3pi3hy6BqmKFE79Tr8QdoZTLttRwCFtc1U21lTSDvO
D0Cl/yYA40cK6ANn1H1E/SJs5C2qfoyOazx5EFFm2reu18BOIB8jHbrWQqmFSc1sWfWrJqqpSUG/
pc9+/b9u01MwI42MCtQz9K7M250mruS1WrklN4BQw6vJmTWhUOm+Y0iej+EKuhHIZcKHuzg5m3Z9
IvJW1DqzNK8Zy1brqnnRwCkeNaldPPTPOz3p1WEPlSEuPcQ4R1m+HvDn3h8AmoAFG5iNQ0EshwG6
DnbKJ+FfsX600tdnF53FVyuj+Lx4VO39Er1a7dg4Ao4rDTasm4HguMwi81kySNayxyZx/YQLWcF5
omgnY9ZAKFqC4uYInMV8Xer9XDoOGZ4ulj9Ls3FqjcHk2pwj4/jl5kf/OdEAhpuwds+rgIk73/M0
18lXfJF/4T1zvYBh1Btc7ADjZgy+9f06ibQdOByrdwSRFY/uDcF4tHiwAoxS0hmSLZlffO+SY6sm
SD5HwzhJmuJUva6nfCqTGRw/PlF6tQyF8IksHiz6OibKkAp1Zq/u+PklTD3Q07LqcfYETSZHabva
lfFs8SCg2q0vsIzg1ItbDst+uxTy5fOgEQnGYlroQlzMXgWnaphPxUK/MMtnuZ1i0ruSsOV0gth3
h776ajO3ABImW/Lle8Xa9/jfaIj/5vqJvzVmDvt42RfHN6d2LQvZVQtb+5qtm4XcTLsviF2tq6m/
BJIn4LVirkDsXXgc0C3ENjb85AMRHHtammeSsMghRDLvH6a0AGEgbOdqLqw/C090EIho6XQ6fZob
0l8Z84xv2Nbah2WHlyTvqXEIUOaQGF3oEERTIf/5g0+C6iz4tfrISUpVFjpeH6KH4btK/O04cWy2
0nF8RX6X7yZwy2uk1mAJSsRV6D1erfKOvSopH/2t7GNvwlHnzekJsaw9fCkIctu1VJeZEkf9bIZE
DWwVSlInB4oRSVaziNcsef1IG5QpHLyYlrB+WusRK/mknheS+osIfpBVrO1hJvyRkswe/tnU2npv
9FiOIXsQYfAsgWNkzn5FU/bAZTj8EJXqP/MdPxYo1J65/dUR6OEu44hmLb6Pizh1+KgnqynHz4Jm
O4XSQbYChT/p/OMkS3v83Atairk0sW1086iIEIIgc/PUS508QSJrTrWvw4m2y12vuXu3utlexoS9
Xtium5AeWEINfdK20ymCRPaBLna1CirEla3oyQCGQpLly13GVtZTGFT67jmRW8i5wApTxhDFKGE9
6AmOTP1dOLF7Z/yRLpskwYNahXqU7aUVPVKYA2gdmcA6PCWK3TI6UIWBIf9Y3PEWx2Vg4TX+eT9O
MWX7IKSzcss7OxqB6h0QtZAFoA4XVYbP9HhEiM1VVbFXUbNnN9I9l7e0uGCOx9Qe+UoOpuU8dOAt
5y7oljiCi3kEn/gxZujTrQJKrP0aIQZTTQsnGH5T1qits6KImL5GNbCGmFsHxOrqwY41doF2WRA5
OwZbxEXz4vpXrOC2WVjzzK5rMy3IoMGdGUptIBbBE6cZx3Z0tVxpaMjXqNGJD+b6L6Wc629R8Pq4
xpDhXQ1xeJTijpcgiyPcqmSsMIkTq6XJUFCT1zsUEzvuPAMHlOqd+GVzYs9TBe6xAcgdzYpbjPFj
EuchnY0tL8d/xdofeKvdL3nh0Nv3xeTxPSLc5TrapNwAc+gXv62XfqwPlNoW6b+ubVpQPOtHIAi2
MLiUiva+m+EqQecs1JnnGhQPXs7M/C455rqxsKDlcKVbLkWcSoVJw+IXITZg209i50scErX5UWpO
c1tey3xyLeDgi9E05qpyXovXqhmXAnq0BXyhDCSuuGIxK6Ht5TOr/l7pdIsI00lJvR0vGt5wll5m
BV4IEpNW735GP3jkrpGBLhMW3/8QWzlS+o1/EjWefhma6pevMdpENb6w3pf9dMma5JFyTWQ79iHn
x5iqpUpNTYOt9Ej9SUBY26+zI06Eii7hNRhkUcPtRCsqQ9BR2e6mECUjlJ+S4cpfNzmGLG3UuYnC
rE67ofyhBzg3N8jleKW5sL5r8TAppcH6LJKvHPXu4DmOn32BXJnr3hpKi6AszlQZGiZa210nYh6A
Jn4BGVfKbnXtq9IVBveOiwXHcgetHUdQ6mo15LLSupAQ+c7lAJwXVZt05Bb09j9NErfyA7T7wL7I
YP7u3hl95xBqIPyGk+PRwBQ1Bd9D8oos06y4Ayqi64f8+wVHS0TeIYEGDk5bxeK466LvPGJhvisB
HY7Tya1ydeXZmRu15FQw607D/n+qRo/DWjUbkVpmQpvxyjZFf02ZGF71y75m7TzlEKZ+mPr9Tpjc
xi36qrGREOIX1CWh6tmJDs1f8Sn/r2pvdTFOo/P/c9sP08odUq2ZWfg2NMH7GevNrVynwMYjPoVn
H11InCk41vcn+nShbydwVYwWYi2rXmoKOx4ytKaxOyDbplsAbtI9flUF2inLUreV0cZ+czP1FsMJ
ERMiUuAqJBYU8fEokTyICJJwDeYy9h1+efZfw8MCqFoSUlCU36sM4/TSTtkQ4jMTR98/vbHPwWy6
LGc2JXakzL0o4hlx0RoMcU5vb9AwmQGQNX4dFPNQPiref3pxISwKCXwnydfmfKeRNezUOiQwpSse
RYnEKw+IhqIczNsirItTnEbwzLsdSFoeR37q6EgvvWt4YHFSg44dFU6dyFaFKjyrXwmsbZPCqBEF
97+PZaCCwJXrkrqCvFadgatfqjnG2dkyJxFrSiBWnCYGkN+XE0mJbcTVsvx/cYjC61Vc5zrxnvmM
m7lxS6AteFIqUcXhsBCanoBazOw+4RrmIvTrGoSPzOfg1vH7P8GzgmB4reL+jLuuUHPYiRRFLy5h
UM0ounKTr+HGm4r9cRmhPQkDTzJnpIguvHcP7ZR1lnUHJaCbI4OffSfGrPdJ+r635OQ5NlXMu0OT
A36s7X2Nph3F5m4OD5aLoZrFv1iAsES4k1WcuSfrKGVZX2/zLencUNNIIO4nWeXzzxwHwtGHcc8O
w4TcRaA0T2/BhX/dk3qqU+f6psBI9xa6b/q3zprZWffNq8JnWYbZOBNHgl/Z2wlmg/m9ZgzL/uwE
u8u1gVZy+jEY0cBHcnIWlveWy6hAhjFWsGDA4lECbRDi14w5KpBlfDc8xuHIc//vOVAn0GMLvIoL
SZk7umsRWODfBVdzVQGU7LsyOfrjcNWCnCx3zsIDCNMtrd37btR+gYfDgINlOTyvmTtSkichVO3m
oR2NC2KN81jYJLJJhlujLQbJxz94lr2NCQJLIiyIO7ZbFf3rz2o3vUn0U+IboL7pUswAUPiNS4CD
qTEDljuxUOJ9csOg5/SzHE2ayJ9bxVetGOuAePFH0mP9hf2J1xG8zdWeMtR2r4BoxjqWF3zjGweR
5uj1bANw4s5Dp/dQb9oewHrDdVEfUdsJvmIuJBbEh351L3JanEtJa7xaZURn4KnGrgRQ0jr55Gcn
C/K3ib3afOeFNPmEU2I7VN2vi7nCxOFpE8Q0Zhk9jL9V3KAefPbU/treU5VXXzFz7Adb24WZRp3Q
iw1emNofTLfn9j4IcJyEJkjO6U0i3jpGfKKMw7WrPbrTLjxQOT8JmToyVUmcGKghT+q0zdJHkWQZ
O839VXADqMh/RyxPUtFc8/2v7a62TDnWiFCRTdXa09X3QL9BQ/0jN1VYyC4R1TVgQdw+CHE0jdug
SPnffj+z8t0Xx1FSiyKBm/eK72zvz0kGo8QgxJ0BOPW0mbL4VjvaCBGF1I66f/JCUqFGRiiPpssY
p5MQ/K4/vVwpAlmCD03kxh87BsMUMWx70CIHkZ02bRGhBzXHESRAjpOKZnKdvQgdguJJz/lbd9Ko
8lebFtKuIX2joUW4xn0DHEQfqAlei4xWYxiJz4aXqXXUfGe+fEqBKHBhGpPoE3fM2XOjWL9ifeer
CiKqkeBZeVaVZtNBHNYQ5OUEVimH+lVz/x/XTt0nLJU9mheAh69tjbnGWFY5dl9tifW8tWae4irX
6dAgMXG0Bow2zmtzR/HIMtBhVPwIr4cWxRX/hUdGADeBPXlsb+FV/iGu2By4H1okZUyHQoN203Ck
76AKsTDiWMicSa3rLPKzKq5epMtUe2obeaTgxkyxsrbzm3uikaEGVc2FDLvdALnH9h0r4nQSb+ar
GePof0sEZrIRlPptMUmh3dsxqzqRAKzNy37fkEV9BVz9KzG0EOyj1JEmxcaZ5CZjUNYIW9AR+Lv3
BBDo4DNlF6oliBjIDDWiLonQtDzeJjuljH0cfvDkvfUq4waDc8uzY46AmdxQSctqBoLVXrdeMm8K
ChOpYgh3go0EdlLq4wWtOdzt8zbJt3OmUR0wphemvUuI67iEXcSJlWo1TGLxU7DdNLVvI9pghkVh
+HKAihALXf5v72xff+2L0k5LThwz/sjyRf2vAtwqiNVPO/3jSCWhHiBNQVIw3A4J/3LtWdze3vK3
BWOKpZT+p1uN5xMxiu2ilIqAzG5WtGw4hyoPazRI0DMJnkgF95CmE0x3qeo+oyU/KZdyFwJYehW5
5zKZ4aE4wmesSPEY6uJEe7DXU0yNFqCzr/LkXp+DIWbYxryR+IQA6ECc7gXTAn8dJnc9bqzSbHww
/58zcvXO9CFJYlHbmZVTqnzumGPfqMFc3aFbqX79N1fwCyA9qf8h01MwrE8m5+E3P67+c1D6i/yV
0k5USsFWyuQ23QD/FoZpgmz7ZezQOL5POIJni1MRKPUmlr6UFTLNWieClVa4pHx3zn2yr4NbS+YR
2qDuuHkqRHNBOqaU3TkS/xIZkw7fA8Q5WprQeonVkE83Zopa/v/n+4XqBMpb9jFrf4+XJchTLl21
oZ8VgkoOeFJ79qEKlawJs0SI9pxJM4/zft6vJVS49hmHvohOzMznBQJ7wIMgJRxfZinpI3ZPEUS9
rIABSCoD1+r/+DKKsyJO6K3cBNcEXY32BBF5A15y08FNcfCZ+XdVloh/zhyc+qFMVR3iGT5d2nZu
18+Fdvw0uaTzkTjq8zPqJazGVPg54cYxlzBkU1rvK1R5AgM5wi9gWfoaibuhX0JPMU86logyVNKP
lX4GI8P6iVG2ILn10POXSOnb0CTyy6CrNyq8nuF3wii6FKQhEmzZdqQ+HExN3o7LEXZAMDDGYKYq
4dC0yKez5K2pOWfb9TNVl7V570cWrzDOKtrIXxN4EUCgMLnqOO/NHE9FFVAxJZ8vE3pS8kB/72Tr
DBiZF6Bm8J/JUwzCvaVxAE7b1cKMver9r1nlOg/vfYFZcac5xJFmC4fPhE9mxOC/5BzjAiPO4+Yd
i9DeVhfhCILN3vykZ2vIAr/TLwfTCfzo7S9gWSVZVnBMMZ2tf6Sln+mLlrSmmFeCbF+Wd2uNa1cI
jiYIn/aQFZXQB2iad7E6RpdRJ5Nl4XxI2dxqfz3G+i8sze/EYlWLT7trmz/R16krT3eDzWu4qb9M
szJybQxsYc+DARX2zydegMHIZ8+bJ4mHuTsqUtAnqsOXW9kUDSoe3kTGsuc5R/lQcxcjChsMcuyR
0/Au2qfyn/o6cLX4u666qilZWAIid+3fF7NfybTUZKGdzvlQMTxLNfYmCVsR420y6jPwhAbF3SSu
eVBSJipZ7yj09WDT5oWHo9kVbYOXBCva+aqPG3jE7hnOV3+go8SdPp2bcTdmbuPSumex1WXRKsPY
IW8Cv9B2COMMq85+ZZ/afjRkjVJnGFJ/np+zzl18Fgptp1uW4MgNC1vZbGldeRCxe/Y3Fx+EpZSS
g9aFGAeDfIIVt0i553M02FEgD00912OPhejrLE5HEgZDmWpamM6E7lF/KANfk/GqgOTfUrJ85sbn
5jLSHAzUdIOOjnHTPsoiOPyYoNeaoISyI5dbBPm6DHOTinFMjlevwkWm5H0CMvYXUulFJet3iPjt
ekx16jkgppewzr0+mrdhHz5/eeiSKKMoik0+DDLp+ofZI3Fa3X8HGrFODe6uK9VEk9K7GJkwhw9i
yQRx1yt5jjImGyFFWiWPwjU2dnl/HrSDBzAGPXyHqP+SZ3cie0I51KVCSWXjQwVGhI1sYkqqjRwD
AbgVytLCqGYKbejv
`protect end_protected
