-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
TeemBKho9Y1m8DZF/3ukD+mQ4orbLBfKvfh2FxqDX4axzfUbKI0N6MMQO+ISw76tyN5t2Gjz9HN1
iwPrpOzR/oggZOSN3DZ+iO0euk0uDeLAeJMCYZTbbz362RwN8iza3Ju63fUShNycMVUAPFUqiFtZ
v4fXKeMeOf3CnUnL+UidqMCaVAkWhZ6mkkYqNHeCiwjK3xiA1vHeLiw1ARLIB20LW7TBVLNL5HGv
waKuPXaPXBRnSZKhcEK8nQPpgLLvXrF0CpiKRwVOAxVrwER/vtW9euFNL/xd1Bmgm9DyPt7SMpCJ
Ol9QblEkQCSNFaHdV+lNO2pYPizqsxVuhkNvJg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 2960)
`protect data_block
Lzrec4pzteaojocWPCFShTCt9zxu1ldIfHnqSxh1ml3yZpZTa5wrjNC+SyhvpFI0iPCX2mzYrVat
D4qz3VsfVMpb/kH83S7+OkmP4HUQZxK+WnnFyzsksEZy15UGrHXeIvas1zQCOStxDb3RE3TrjRu6
jhUfmFGhh4JLzwvmWVPLd5FPbsNnntSzA7t/G+YyGogYxsqGkmPNdRRC09t5jCCyaz2GHUIQTuAJ
WR+T42PZ1/a8KfqJLomzjmxJO4mYvOE+eqIb7msxDYr/mGh2k/BaWNXFc/X4UlrNGzAHeVrxZPYv
ROPdzFjZjCPRLQKzxvHq0GWa/iqV4Brsoaa9EVyZlC9xRdfrnRNMHWBAfLkIPWtpUdwY3p4KRCrk
wQv6nHSJsAVvmmLm2gLX5ZwQEv7qkDEChLKneaVJWDgC3YYuSAdpwma3PHEpbIlrbUn7PM91ZqEY
r3TmRJAYUnX+gGvTkc8IhDEQgqe36wUYBXKjtWssTwlT0JNWhVEJHFNmwg9lmCnjsuYli7vE6JVV
avYNCAJtZhpiqtpPPy/NInuJkoFQnmzeti4MloywB6IBeNDC5FD1mi7xlJF3xowHgIhD233GlVkj
T2eZC2Obv91vFmPtvTyswPOshTs1KH70TYraP3BZWiWlWd8Dq90VzOrGLMwEH7PQcY4ueYdaH6Mr
+BoTOPvHxQC8Hq8yvfvVrht20SsOtAaYWt1SE9IjwOpkC4icmcKrpbSf8jtdjejZ7bGtFX4YMkTM
JmEoUIUPEeJ0Gy/d5R3Xzet5mPaSSN/sBFQGLT3ove7eyTMPn3753b7LN362TU/9wg40traRKUIb
3JX2j2loxtFKjKN8ZVu72xW2XyfqEJgHgr3zFaItNLRxieYgBv8QDJTVntE2O5DTnkFV1hjqXctR
h/2WlZr0xfq8vFoKivEVFL/39p5yy3sfJzRgrrEWFUdjXWccIFMFsm7HVpwTy4kHVJAHosZjEpiV
YzHDT5oud9cdRzLM2bPkF1DaH284y78oGcxNUIyRN6XGpRiHn29lWlSq+KcyhR16AQqkVhv7wKrG
zpTqGXB7veky35PJ/d8DEuJPsGE4KVNN/CLruBTrg9waehaFytBkF6mcX1c9zsTYeEbl6tVwmZ0K
EnUxYzjcyjMcPbtZUjECse+qGr0akAR1FhvNIzySYOJQ5V1kTne8lkqtwteWVvx+a78etsf2J+Kz
ElkKlouGE25l8ppjGgriPjjc52+2nVFnn4vU7LJjZ3D7Dl66CoNqTXHgFhL0yycANVx/5yBeYIz3
4hmjRaIuaf+nruCER9LyulXVAznkTNVjco9zEWbKrFHaCVS02YdJwu9L2rKDQ7C/BniWbUwdtKOx
bEo3snX/dYtF8CDSWr7KuRcw4eECs2diCQWWzlD6JbUbPoL7GU3ZkD6MbbGX5ZQG45vF7WuDaOu3
WVTkidACi1AQag63MMc0D05O9WzUDdmgHzguIzQvLZRD5rMoRwTzTJvYk20PnVRwy9YowiiymhNi
HZc4jELLzxHsmUpUPzFvxhnFzxPy+uab9rZjzuJG23Tp7lC0bLyxREEXqeSIeQGLpQRbqvhNiEDx
3ueNtB+2YmjuCDKnBrNSNHIQQlDZQ3cH0hHi5156cKYkboU9H/RNOAXjxx5PzaXhhpP2oBfZDtnP
PG0uKKNZvlDGIZYhaaeMGUSMhGGLeqxP8w8O4HrmbltqLW6aESNySr41PTvw2sE+0TFZf7r7vFo6
CZny1amTJGIzVQN6xX98sy/iCkGbrLmgNlbW/DzSorSckCJGAwmo3CRHNDqXbOpXlA9QDn7E4q5K
e/hzFwOSdRE1vqRsczoGaX3/NFR9l3tlTQ7yryah9DsaqnZvCa3phKL2VpGe90NooOjaP+1U/Stb
Rv3gEOzq3nNCeb56Mr8Se0KhvhhJ0FfCPqF4z3n+DgUedQsm9zfPAVJg/XJ5UuLr6Q0r0H3gErYI
dcExaZGo0ZqA3FnNtud+rReDXAy5LkTmSoLglJMbuDaGP6fwh/d3bmo0G8EtO0eH5i0PFlAYmGAt
RrOzh7X8fvuOJAI+x+y/lot03oYDmvNO10MYyi2E8LjNDrSETUVaqj8akueVJWGQGOAcQZXJ/YYa
sXPdhoZiaVEFzKow+S7DzRnKGg9igxoHoshjk6ZbQN5mRSHzhSH1i9pRkD01SraK32Y9KBudLDvx
qPDKjWr1xITDsmGvxvpBBCi7SK53cPSBn9l1xybegl3gDtRL4H3XF2hWA1uJrzDpAOwrc1p1SVeg
h+S/MLBdcQAPpd6N3hqD8r60FmIxJXtJaD6E1kC1cvQYVnVPJkiivOqdiHjYDCHieiCIgDqarhZ1
j/FgN2EFG2IZn0MMq4Cw/cgpHBkKFl0vqaUn/AwJ5N7RInfiDE3L5JtsDFy+1rXOOqA1sKp0kSNN
xLyRT1EkKuL7krQG+84DIGYAUPTG6AWrDX/IFiGxXY7t03JfphhQqMniuAvHsIuZM+ReCRcl6HKc
PEIDrXFVe2+hmJBLhloFqe0YzsfJyoAAkg9tT0mo6yuN+t3gJM07zGNAdErbBIMwl10AUsYCWKNL
8OmOl87VFreyvgtrnLsugtLYnDP+jW6ULFHCyDc/TNu/ed2ex/3fUrAV7lsKTCTAl7M8471d/TqL
oJw+XiinuF0vXCUg9D1YVDHoGZq4C25E2pXQaYcr31JC+igB9SDTrLlG2SZBvD5LPduVCiOgrOfK
8HitA09w08Vxy1+hEJS0pQBuzxdvfq3pU9WL6pZvItdb4RiwPGp187pt8C8Z5hf3IG2ayI67Qmub
+dZaz3+jqTj843N4CYAfjwL4s8jTSKe5NST/XdjujdG6KlpHxx4+b2dnVDSXxJ5KHLaF3Z+nLc8C
eCO0SwCkDluFOM0nS8W8mXuYL0ALFoa6qMKUSHIcmIlpn26THMZ75U5cpcVohZ5psUpPZwzvQC2q
nw749qiqyYPvTOT/TFN/NZLf6vCblAn1PfDFLGdozWsvJs2UgNMmonqh1nIeQ7dbP0X5q4ZX/bSX
kNk49GSgvjuvWHWTeDEkj1ZD8wAeVTnAQcMiRUE5JCmX+VNTLVqktGxvGRFgNcUf87K+LzJg1y5b
vCFp6Yo8wf2kjbjrGleeuLiJ3SRDBu/jpUvT65u6ORZUemMF5bEGeFvngOF/QuJyLJmkWZQPswz4
3hOpWtbwbzMwM07P6tXKwUHtSrSEccr92SckhawYIRVsRMNsFWhfzBKFOfsI4JwYEuhMrmXyjoLg
q59wPxTLj1FTWY6o38dTkFDzq9OBdblCMTkhCgJhDic2+gNuS74O6CyR77yMDLj8pT2FVAs9d0Ul
bpSPSMNr9H1oulsxV34tmEtlhsoelAvXGggg+kX/CbU8Mkcp8iMwasQUZvBHUM0W6AL1t5taRrob
fUg0JHO1gFbE21fbcNSfcxqf9j3ZeH1wA9sFxA3L8rTOCR4QJAteyYUMPZjJLwUWP7UO51uq4/Kl
mrMOoYRNMmcpOV95d0nK/XGbCVepdcMhFMPU5re6o9Mz4g8cZQr+Y1jD7/DVKDzdgfZG73DZxYr6
IH02QmQeR5uy/wOU3KDAGUFBxpfBfBg9skt1NultsVuguNDje8qAkv7+wo2gDhekolUaAPFUuS/v
yXs09nwHIGR6E0Yqfz7B8yd8ktKePfMrYMSvJSas/ZjCLBQk9i7ca5dZ7GT7stl13j1iOvu7P1YM
JlPxab8lfpxIcSdQv+VnFoIs12wxK672UnUQQCi3Y8eLlVVhPJFbW78PYyr+u4CTSGax4gnduXBI
KoB6BSTAXXnlT9vzdG5BmyTx/kyHvN4nD9UL369Pv3emzE1zbn1cDtLlyY9EXWg4QMUmMyAHLU0V
IlrjsnqL+iZnAjwA3NNEiSneYqyy2Afdd2eW5/OQBbb3YkVmzs8slNisPHTn+Jw5zf5MZPo=
`protect end_protected
