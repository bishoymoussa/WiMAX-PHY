��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$Rx�y�<��wA�*;�x���@�̦�W�X�fa�M-$u����n~�%���P�$��W��kYَ���P7�?UMfT��q�6�U��k�>����~�\N�(�����X�e���/6U|)�X2pF�]$h���d.���9E�	�IN�f"�\��e�z�y�b�����Oo2�?�qˁ'�͜k-�K�P|����y:����3�l�d���bl��ˢ_�d���kx�rq�mh�MذM�`aS�.�DW�mS�9���Y��+�>��!��!�T�uOB���,��\L�7m�O��W���6����'���j)n_�I����2:��$�K�2�Sʫ��l ��!���{�l����.�j4�	��很�̢=�����N��s���s5���_�R�>����ТP .W;������	�"�מԫ�����]�#7@O+?�⡾�Ԫ���e�O�\A�	�ͼ���ƹ�d�	@�nQ˰��E؁Bf���|D_�%au�-�'���w�*%��"AM$w�*'�wY���HAp����E�o���W[��`�>����D�^�}�Ɔ;��`�
)�i6s�=�'H��]ٲy�Q���-�
���P�6Y8Zۗ5րα�9�ZZ۠���t-Ʋ1���?�"��;%�]y6���R�����e���mv3�5�R�99���su�#3qѸ�'�YwɅ��TQ�9��>+�Y��6�E�� tW@��bc��O�@�r�ꛈ�b���4eciU}�T���!	v�п�N?�yY&�h2�V��{��g9��+��_
�94[�\����D��_���N�<��L;�Y��J�pB/�Tr[(���~K����n1��BN����7~bf��j2ߐk(]Z�t�=�����;x��Qd(^�cؑ�K=��Q�8j�6î.����g^��X��uO)��Dz���ϐu�����,�@�Y9T�����Xb�Y��2�����B�h�/�VZMqCB�9J����+9/�9�6y��3�(�:au��=VT|J8?�x��*d[��$���ֈ�i^i�6�N�� [�����OWY�jJ�n�;ȱY��맆H�kyE� ��xT�*n��A(�Pg�Bx�2��,�QQ��uYl-BC�nH�j=��l%*!fB�\<�q�Rs�Tߛ�[���2q��	o?c�Tl+9��Qj�w3����S���Y�gg�p���0dǁq)T~�r[+䜔�>��z�0;�H3�XD�棈�Ѫ����������^8~7����^���O�7c�{�k��J�ߴ\9������k���̑䷷l3�:�c��Z����F�$zr��
3j�Ĳ��N����:��H~<&�@A�3��S@e<03E8u��R6@���i�\�� ֐ux�FQ�����u7Za$��6&��Y�%p4���R��dh����B��߇��zol�>m�X�6�6�!�ݗ�6N�?��[�nN�B��L#��%d�VD��]���ٻ%�T<����%�}����kOΉ2=��\'^F�[g����@]�A6'-
�=����>MKU�P-�30
|�!���a�����'1-�]z�L���8�r�3���
EC&��z�z)I��UK��WF�E(S�L�1�+Qjw��O�V��Ꞥ UI	a�Y�ofl��A �Ф��9k��b�:9�3{�Ox�7���U�$����?���c��xG~���������^�v����Ě�� ���6@|i�^�[��"���r������[��r@�^o;�o� ���PO=�U�@�4�pnb�������2�.�������Z貕�HI2�0X�o�,�2�7�J��*�<�]��(��IB7^q�n�5 2z���XF�(�dӀ���d\`�4</!�ד�*x��w~0*u��SzJ�(jb "����i��ֳ�@�M�.�e���9��-�Ĩ�-�s��4L�V��K\C�PRU�v�:`�ðrÑjќ��N�6���4L��L�(1B�����<p[p�`ĮmO�=�0�<�-Rik��n�1�L50�<x+����+%��Bܲ-��+0O��0]������CKEӝi����Ok�Q�����5@Dp��v�_!�܎��k��jgL�r$�Ӊ��{�)�s;dy�6�Ω�nqC��@WVV	>���%�����ٲ����C���{2�?,_j6�'mI�'����iR[�YQ$�w��\��}�g�rm�e��ˣa�/�g��p#ޙpfͯ�X��@+�;�VS��v1���1K�t>�	�6�o՛��Y����b�T�O=���KK��Z���t�� �����B��݀E�n��F:�%>�>�Z��~���{8������Z#*���N(�n�K���(�=���)2�Ж*1�.(5�sƇa����o��+��}��J �&¶P;Ju`�V.�H�4s��n6���pP4Ok�/�[����N�C��Tp�aG�՜�V�X�� @M
V���-�?Є���{qG��%Q��4[�5����׏�`�����# P:���P�\o�kMF��SE��S
ŋ�`x�{�a�~~�I��l��B*K	�"w(I3W9r2��ۍ��9�N��H�F�-���_����F�j��d��V����O�,>Qf�/q�!-�H`|h�e����jy=�*�[ GCOЧ5; 0�/���C�h�1�5�`�͚���T�;��7�[��0��J�[��	�킊L���%�����g(J�L����l`�+�6������y
�s���&����R��b_{�x��5�����ZbY9�[��d)��+������r5*I[�i3[,.M�U�LӮeL;\�ض1>���{6��s��B�5:K�6�`�<���9�T?m���abڠϿ�C��q�ka=c��;-g�0�ݥ)Z�[m���V#4	Xd�0N��,�;�Ѷ%ƞޗ�c��cXk��Jq�2���*���@�G�8���q[}�l���̉ከ��'���M�@��૬~>=� �o�4�oď�W�ltG�_��.�k�QN��ǋ�Fy���1���K������/�Ϡ]�7(�TZ�U�m<�|�g��b\=X�^�����J(o[����d6�����7ߑ)�{.��K��u]޾���@��sl�E��k�^f1)�J}�L�>�8q�􂉪�
A����H��c1���@�3�X1��l
[5�y+
}�&����?�����T��Y�"���X�j���΂�OQ}�f��,Y�7����Ι�g�mk��E�']�A�P@Y'���9��� ��ЃAl4!�n?�W��S��^0ٔ����X҈��1��n��:����{���F	������,�ca����Hu�2+�A����g�M��{����4f��h�~+��Ǝo�T���vp�K�!P([2��y�n��>��~/���(��"�@�3�����*?���oA'ܴ����}Q�����T�'ey>�i�I2��P4�8vfO�T�����*�lS`^UR7��aX�o�"�ea�V6�N��B�z0t��?eᣚ�c���� �j�����`Dd"�����?$��?��U��u8�V'�xޟ�'Q�{�'.��TYh,�">8U���;7��=�����0D�,H�XO/�Ӌ͈�Z��*pn-���!��[7�E ]BH �������Ɣ���]���+ 	ֽ���K�­LD,;��/y{5�m�G�ˠ���vDϙ˭�k3Vbl��*�p� z�s+1�� ?0C��/X$�uL�m &��⨐�lcfu����i�ʟ�2G��h������%S,L�=f���}�����y�����Rj��f�a���O��?WH -SQȮ�������(��)Bm|#Բ��:Q�>�`Ŗz�B�]���S��1w���gN.ӌן��/���N�Ǡ�5����˜5�2Y��t�xݻ8��Km���$`��:1�n�����_�O�/��0G&Oæ��@��������=��Hl�E(�r�@��# $]o���a��
��V���_��!�L��-̬��aR�=�����t>� ��Vf"8K��R�o2��ˉ�m1{�<a�}A�OKc��`�te�XޏpV�$]*���\��ڷ�~E���A����ZT}n:VI�P�a�#$�8�p�IJ!��K�[gD��Z��W
),��1���s3\S �_��؈����z�I�0��^����I#�Q?���q�f5�Չ�_���g�9�X\N��S�,��±��#Ĭ�@YҐ�7�4 ��vͿ2���:MM���x�c��,`̑0�q�����~�=�� �A�ɟ�'�M��o9MV~�r��l��x4�'�������Ojyyǡ�/��e|�6�W�ұp#��{4ki��{�(E8�[�s�|g�p��3�j�d��):/}$Ƨ��+#�����������[*�Mٌ;�$cx����	}{�N�<C~��p1[�r�w���9�X�Pc�}Пo�1r�ǻU�ߒ�҉^"� N���T%�,a�}IJ��/nU�ʛQO�vz�� �!�*�^5=��ļ�Ǣ�lD��Z"L� �r�Щ��6��J AYd���z��)�a��K@]_�i{V�d��C���&y��wlN�PLn5=�8@Ω�w%*Ve��7D��o�m�J��P�Skк&X�U�v�V_�U!e�Fj`v��,�׬Pʄc��YBDp�i݀mD�l�!�*X�����k��k�E' ���N���Eʹ����Jg��
S���!3� z�vn9F|�]���uSG>:��Z�Iߚ��{�W�Єl�0\��l�<�sYq�"w]�K�>ϟ�xJ�_���Ox7�����*7�m�S�)�}^��nr��!�l�&{�JaNHݡp�$�ֶ��|풡�j�����%!lQ����E�ЮZ����>X�F�q4s|��,�n�M��P2%U_���렛�o��/��]$}�o`��v%?G��\iL�~���ܣ�'l;�%��$�<�N��Q}ܔ�x]�Ş�E�h��l��)uN�+e7�?��s?��̊6��� 1ԁT8��n�b� yz7�*h������_����R^#�{Ђ&��#��i)���Aۿ/-c#�̮��b�t��&�|/�ُjD��9�}���$秈|J��dB����:��y��IN.��T��Ե�仨�|�lZ�ZFu��J{��}���F�ɕA������gu;�d��u��.�/:�:�HRg�M�.�Rn�gK�^�c�3����YH܆�\q��j��6չg���=ek<<�!�����'��q�MieKlK�?� D���6�.�a�0.GH���/���6�\�L`KT>�+�F{%�ٟ{=��(C{gƕ�;xo�|t����j6�z��9ڬ��?M�{�����m�Fj���:t��Q�y����>�m^�	ld"�Kq��{��1�6�X�Mġ@����_�~��Oƒ��Yf�j��֧�_�=EBS�D?'-ʎ���=GH�[ۀ(�r$o:���,ފ����:��Ї��J�K��	���3xqUD�t��K�T$�x��[���O�+�M��Rq���Y8#垃ܭQ�f��j��8�#=I�˨6�+u/���x���5Vp���<���q�-������\���V>�y�'֧�aW�'E/�~�V]������F��U� b�]ʮ�\�}�w�����"�b5��>��4D.�TT=Fΰ�08�\�\{�s�r� u��'�%�'��zƒ_��#�Ku�e��ŉ;�ʽ*J��>J��߀��n_��
+�kT��/�F��������,��[mm93�m���V9t���ݒN6,�xx/ǄVfD̀k�
_�����;WׁOz���!��l���U��({�t;v�˫@�!uS��A�:{{���[^T�8�� =E�5l����ez�5���w��C��f�V)K̔u����`�D�Ha�8~@(Tr�����}�h��9����T�}5k\�(�����=c;;]hQJ@ �(e[���)�E|����!����s	~�P瓔l�76�U0�\'τ��uyqh�!�{`޷П�Mm�&�a0��x�f_�1����|�픮�w/(!�G�����3���f����5wʖ�q�7����5�|1��Z\9�a4��C���!G�b�Fswvl����K��������t(\��X]>o�sdZ�(6w�%���t��d�N����W�@~j9�����7�6������}��5��}[��k��E�h���g���7`:��_��޾��?�v�h����lf16Ho&� ~���
��#��¤�B΅�ꅲ
����O�1^tg٬�߯���#�=�Z%?A���I�_0����a�"��ECNlt��,H"���X�V�%�7�������J�4B@Yw����K%��L'a�;��rX�&ĀZ���W4��QI�c�� jv�V�a�␠+G&����TM�8X�D��w�ޒ�w�+�׵���2G4�T�D{cxy��Oc�^G?�D����(�3�j������ Тe����jQW�N���/���#���y�x}���T�)\e�:��u���)=�Ӹ�a�[����|���I��/�)b�SO���"*yA �IeS�L�����G��h}Dn��ɌL���_�{^1y�"��Z�h���g�l�d����	��-ub��)�����trm��Xh�иO�$A~������G(х�G�0��S������[%����UZ ����'5}F)B�>�*��,��s��8֯��:�|vȜ֝S�z�Ɍ�R�ݭ�r?�N3^��*��")��@�Fp��_��(�AuqAߡ<۵0}�e�lqXX��pA�c/T ~XN���g�@\�_ !,
��l�3�{9���.es�Y?�(j-y`L��:���4��RKy���0]�M]��T0�1΢�[�	z�P���H�-��S%C�c���͞o�9���T�j����c�̗��{a8K��:>���ZS�$�K'��+ 2���L��ՙgi@���G~��H��w$�aMs��]��b}�x�o)oFcU��� RYcbmm�)c��3�3�A��z	��ޔ�.���A���L�?��W�_����;��O��Lp��I�W���㧇��aB��2��XqyȺ����Z��{N�����㊚?׏����g�㱼r��5nRS��:�L�ģK5��Ђ��I0��Rw���d�J�o��]�������]ޅ�ω�bZ/�a�TuIL��x| �V�,��]��n{sKj�	9A���ʓ��f����~���{���h0���Q2������Ej��C���Wq�!�K&��f����V���.�$����� 7��[�yѢ��7i���jYh.-�ݡY�qm�0fNd�`HtBiH��Ո����R�vu<и�)�o�h���ڂh������,Uozא�M�a3<q^M���)b�:䒥�uq)!���$�D7x�	����őR"���ĝ�Vhé	/g��+{8�	���ޔGg�AH求�+�5�1e�_���:�{n���; ��ؒ,ʲ�*-]
щoq���T�R��Ʊ����%8N�����l�fV8�=B�M'�{�ˢ��p���"NK�6��E�I�S�EÅ:�K��Vh-�*s ]MEx']��0���Y��x�{�P�"��Gv�ݔ�� ���7�;/�qՐ��$Ɓd)5��.5X~'q~1ӧ�z����[�T�ݿ�E,S�Sl�����øbu|É(��!�I��zD8��,m�;k�(LhWWgv��r��|�FdB�P��X�D/ĳɴS�j�(ĭ��<�V��#���0=��64��*�~:rj�'�8��x@��M80�6d׷�'F
�4�+��#BA%:�����ANw3�J�#��?���&��_�	�k�f�\R�pv�t�'f�K�T���0+�x5F��+0-Q-�Xֈ�Q��R�_shpQ�]*���>Zt�>��;���Q��<�&-D='54iHVM�R`���H���AJ���و��p/G�*C�s~���)>YT�t(�3<����w�&s����E�B�>��ve�ίiNV]�_�%���������H�Ct����Mn�ǅ ��p@b���wج���sz��X!�_����SԵ������L)�鋢���Pq֒v����7�L��j�̦t.�ظ�|�!��0��q"[�J�F��)�C"؛_���={nu�1����`R@�'�")C~�GG�k:���[l�89���y|HX\��� h��w:��B�Y$�}��+���1�uE�/�V�PJ|j��^��ψ�͉�wu����K�B��&K��h�l�/֠a}��_�1[R�2ȺY����c���7��&t��L�C�$!n����x䘭I��>��D���3OC@���~Z��I���ۉ���W�(m�Ī�'7m�0}�{�R�l�,c0un$?��㦀�h7~t�mn���L5�%���? W	�f����6�a��o0y[��/ݽd�����B�̬_�(0�=Ժ��!˼���}���glP��>�ԭ��C�k�޻S�3��JD�B�#�+M@����e���H��?SH��O]y�zM*����Cѭ���T�摫�W��З��f椂	?U��V��l4<C)�M��*�n�����oʹ�a�	"��3<�؁��:4(懠�
4���Õ�
$vʸ�	b�X?�+�ۮצ�=�9����n'��bJE � ?@���l��6�ȸ(e���V�� ��a��j��sv&#�--���D9ӊ���y�=��������CxV]�/��XF����6Kz�����E)e탓���w}BH�r6�_�'�Wݸ���pH���'�����;�g,��%�$��+��)a��(��"sx&B��-^��
�Y�����I���X(��P�,��cM�OE�v��Fت����4�Xȕw���*�i��"��G���Ѱ�g�_L�<�t8I~� ��;���B�,�n��)oTTظN2�'h����4nK^�����OO�LN���E�πBy�U n���]�6ٴ�QN�ғӍ��A��+�(D�T����F>��p�8����Q�v��G8�x�:!;d��� ��_j)�j(0�EY�h��o"��љn@��5`��������A��H=�ж~"���_�*~2���PT��QW���K�V�䂱4	���.�Ց)�Z��F��R�5��Ř_�ꇜ�7�9��x�nߗ<\� �
�At�DI	�
mՐ�q2p�+����3|�Yݾ�`Yh��3��q����ʹE�P�1^��E��N�(�����/�!��V�8Eo��<�خ���\�G����2���/�&�cQZ�t�8�B�
,F��ܜ>�
�
/y#fF�y���mF�
QL�n6G���dz<1���K��C�{�w5��pn�{��1��2X�Q��o��`=�quixF\+t�I��L��$�``H)��,u��Bpv)0�z�<�_/0��P�<��d���	<Īٛ�I�ȸ���c�k�Hk���H���jK��._�0GmC�� ��aR��0t	� "���T�%ڌ�j��s�ߣ��P�ke��Cf	��i���a�����ֆT��֪舉���!" �3s�`�o
�͚�V/�яĚ9S�`w��j�`�k�p�l�9�EiS��{s���x6Mb�Y�]h��J� U�0+J��9�XN�<``=6�֭����w��sJ%��-��E>���"��1O:����D���K��V/�����ǛI/cJp�\M��|�.��m�+��ED="�D�GX?2^�����=u�GS��T�����O�����Q�c�x���ߦۙۈM�x�{m��~� �#�n�ai��I�����v1{E=;}���Px{g%��*e�v�[������КC���Q��ׅ�F �C�d�y1���]����:�!���ڥ��3�;��@�	�q��
-�>Fvf�|)���o�8g��tB�S NtFqD�tTv�Klz x��U$Ps�r踮�o���,Q�ucڱ���j,�}�ATuV7d6"�򣛧��rV�j5Q�<
�/�3̇�Zy$c�*�pv�^��!p�6�N�������C��XXp�D�^cZ�
�zZ�t�=��*�v��y��*jG��T��� 3L!�1;;Y�s~'�(r�"��}�8�����?���z5T#�t�v���&ȥe���nׄ'�9������|���0��W���b7���$;��D�?�\��I�>O���nFa!ࠆ`'Id��E��*45�4����!�NRh�_z����/1�c�Tn�|�K[Hi�V���M���X�)���� f6%�?/p����YhE�
��@o����j}Ű�	(l��p�XèrL
�x���6��=j[遝����	I��8Rt�Cr��?l��Q��W��J���
�U��'��«��J������b�U2�S`���W����#���V�»�%�5���2�u���gO��3_�Z�^%�Z���N_L�ɡK������^�I��բP\��3���$D'e��~p�j{����Ī��d�&q��V��:l;nH�����(x��g~�:~�!��9�q�%�.�o"�/�rZw���E��>'o.�|�+ǖ2�1���x������&_8�i��G^����ѳ"���x��,���k��~�����Ș4�;�Kyh	�&.fXk�b�p3ޮ�z�� �y=[*�v��s���q�޳x#���p�*S]���}�+�a﬇1Vu�K�N�2�9|�~�UY8��k���8�ˍ:��>vO����|I��X�ɾ������׋��)Q��
��7a0��D�6D�L���t�v��^��u�l��Z�r^���pڃ�����!�p�2��ſ���Pɒ��O����rR'���ܗm2�~8l�=la�������Y���L�mA(YD�����g��Q�>��m-��?ؐ��5�j�w�6��D>��q��4)A�jk7�,����;$�;]I�f�n-����n�!��kR���2�r��Zr�./�w� �<�n�7D�Oo���k������pn�"P���_�;L0��rT�a��V��<<ufI��S����\Ys�ﶘ�@��>��n���ꄳ��nC钮�̈]� ȷ��<jQ
��Z��`��쨄��Y3��%���c|��D'_u��������"��u�-p�C���oO���؟��:�A�9�b>I��5x��E��}���mzy��٧c�i� �����%��^�Tmȋoh� ����lc�ƫ�R�0I����Gf��"'�$���-��S(��dB��d�^�E�♙�M�9�g�(3��Fu76	n&o�5?s�D/�6F�]��b�
ڳ��/x�� �P:�4�QI	T-���~�7��TY��k��\~j�k
���s�&�k�0������W�oeӮSy��AE*ۨ;rxV�*�p~ A�K7��� ��U��8�\c�ڮF9z��';h4vs��� ��Ϗ�x׮B$C��6����վ	�
�2	 ����Ѫ�o`a@Ǹ��.Ż/�}�{�γ��!,H�6����u�B��.ϲ����S�2�Ep�I҈��!���zf�|z�&ƛ���UorҠz���D����Ћ�k�޺B,)}�S� N!�i�l<㪅�;�~��!֑�l�`Eō&��nZ��b����%���sK������8�:A�/�s�?>��-Nb��{�������y��o7 ���e�t�e2�xHt�jT ��DB�vw��I.���N�a��?�q4����9gCY_������lq��Fl|�b��$s����q[�n�E6�h�,�e:�m��U�����˃
���q���?!˨��#3u���P�!��}u
��;eW�ܗ�?����S4{F�:��x�e�,�Bʰ��)\�/��;a1�+=�=R�/c��F�ê�6�?c�pF��M�$S�	'������ �9��RK|�Kn Ƥ�@ tu ӻ8q�1�y�l����x���a�2Ǐ	~B�f��M�-�eFe�]]5�cJ���쏔C]����Mn�s��byo�o��s�}�����V�z��2�g��`��(*�Z���>C�5��²�0���q�R�(C��r�dk��y�1�ý�~;���%�̗T��7!Au�Ӣ5�cDl&��x���6���e�9�<�#P@m�p�5�������[��#��pQ�!�r����RT:0�R�OT�o�
��x����}�6����|S�a���)�DY�7k�g�Ҳ{�"�C��J^�P��5\I��6�� �[���梊�;SP��OR��:&��	6��6�^�J1��E=p��6��n�k�~X�S-���C����z��45�
�Qb	�NS�*��1���!�MM&$������%o������[�i)��H�I���� '��Q��ڞ[���5H? ��<Mm�K�2F����rs
ռ8�KD' �nˍ�k����E�E\�F1I�m����1��ٛ� ׊�+��2��Dv��[�Qf�~�u`i�Mȫ��u9�<ځ��� �J�'�e����$�g��1:��G�sj˝�'���^���x�y`��r�"�Kw�ʹ���e��GֱǊZ6�5�μ��K�%<��u0]��F>��}�ƽ���ګ�Ӈ���|L���%��m��RV55�	�ɴ�?!�%��n*L�)�rJ,{���m����GP��97p�D�a�p	5$���VtB)lBRg��4G}SˣȔh3�S���7� G�'�>�7l�5�쮊�%�C�8���̾�M,Z��AVbke4J�Y���fȐ��ѮD�-�y`T��Dɒ'̾�p7����!9�hqS�w�|�d�|������n�A ��+�OU�:���c/@u#P�(,}�����d�&�����$ ��塀y���K�����j��1
0Q�����y���ȶ����i��8���m7�f6�6�t��֐
���W�C�&ܧ�a��=��Z�w��aԝ��8�YElA�&��Q� �#���FrC��7���Z;�F��2-$��Y�g��d^-�]�����PG�Dٗ��1������QK=�JR�c��A�m_W�w���7�� ��L�~����9�FrM��Gƒ��˩��:�2���Z)J�i��R��Yc��N)�: ���Ű���J@���d���̥�Uړ�����B�<6#���ǹ3�b���
.��T;�B��@ղ�`w�P9z�1�i��+r�����uO�٦��y�>��@&��i�8�y�[(������L%�Y �[���7������ۭ0�
9�ӘL:G�]��g��N�s2�E]o6�T%�.��?�oStPh@Q/v��q -���*��B�B��/ ����K��ؘ�Ѡ�"{�C�x4cc��Xg��t���H��[qV���Monw)<V�G�,�?[]~��;�\��:��6�Y��rm<^!�UK>�����h��5�� !}��~���X�;T爴��
��b!EN��^<{� t�ӦXfb������t����I)_��!����p��߶e:�������v`����i��#�N��#�_��GH�6���p�C�`�-���-;��7��׀�A���3����% �~2�M������4�|��"5+;��7�*�e=����g����ޡ�SB�\C^��Z}}�z�dw�'*]������M�v�*�Ğ9Ƀ6�Ԃ�x�j��gx�Yi�LM67H�+�]��%�v����S�L���zJC$�U!+��4����184a�u�)nM�8�c,��W��>l�j�Ih.i3,W&e����$	C�f�6��MF��r�����~n�ߔ(�%�A �k���[���HJ�d�q9���CA`);5;�2ژ'$U�	s0��/5�'��h�w�z��C��Y�ڊ��_X�`�s�5��H��Z���q�}͏��8�R�z�T	�1fX�{���2�j�m����� ��t'In3���~�#�"e�J�+I�`��T�#���QA
�������`I9�n˖�"�-mESv2��}3 ���t�IRN,������{�����2B��xj�`�k��`��^�|�<�qK�VG��W�!Ԑ�����f_��z�ͅ%J�2�(v[�ø"ٶ3�]rpr�+�� ����({<�ԬN\�/�����hY��8��R�ٯ^��|���mKq���@ǉlal�cn�b�����-�!�����d��$w	�e�(ai��m����� D�&���Q�������-��:o{�I����\��YKߠ��Y�7ְ��mAeIP��8������s�X��)G����,�~��f�4�o��gH�2&S�4 ��è�5��Y�n6=�:Kb�G�0�82�� �Pw�4r<]y^���Xz`�)!\h��}K�l�F��,9��k��!
����
�X-���A�@$Β[BX �у<�I387�	!��]QQ���4��rm�T2#L��ъ'5;�3�\D�ĕ�)�����"p���_�E��}�[�7x��;z�V��P�*O�;�O8��MV�@�r����I*1B�xkh�ΰ^�%$!����`T���,������Ň9��ϩY�%�Lӄ��W��//��h)h�Z�Ԯt|��y ֜M�2�e�����w���1�+���0G������}8z�k�p�r g����ޠ"��R�[c�IA�JTV��AQ�����꞊Z�B��2��"��HY���,��4��c�`�y�B���W���F��A��7����s}t�[%�*H���|)a̓�N4����������g����=��0�!�(/,�7$�ŀ��ih9�hb��ee��D^�3U*���3žDf��嘁N�}U�ݯ%X�۝�D�E	��J㺀���b���|���y)�7G�Sy�����xvJ�Z3?\�x5i�5r��F*�׹ ]���[|���I���}s���MȺ�Q���Dc�q�r�Z{�b#"�mҞp�p�֜�H��e�g?]:���j��VYO�-�x@�^H¨|Y� ��:F]�Ꟛή�	f�t],��S��&ʏ:9o�RG?�ׄ���װ{;z��Q�l9�u6��k
�Pw�ޖ)����AԹd���	�ٍ��[�Q��٣WZr@������<��JC��9���-jO���������Kp1�'lK���-� >�t�iC�^oH}LD-/>bԊ�^Z����*ե�>WBF���`Qn�c���E�7�J�����I;k�b�k`�qI�u�e��6���j����$zH��EsZRŹŇ�)}L��Ň�? �+�&�D`&�&�\�a����7\�{���&��5j�g�IH6��}AX"7L�
�"�y��15�#7Oww(��T�/�p�y�����kx1�Zr�_5֕�aW>� j^{��dRZ�Y�V��8�m٪�em�i�?+����j�_��rn�8̀��<c
rE�-%��7]Fa�#�=*D}��
j���|�C�k���	|�����z:sW���U1S4��h� ���(��cM����T3K(������^.���S��:^kt��SQ��w�ZV�n�Kɷ=���oۿ@
�t�T�!+��w�i�򪽆b��癶����yY{���;XK+,AZy$[�ۓ,Q���������s�;���R2�	�O��9'Ε���d�i�<�g�̙Ǌf�-.�y7o��&ĥ��k�bCk����ۛES9�& �Y_��x��	���ȩ 2'��UpŚ����w��K��I��"���H,��;rx,�f�G� 4tt�!]�-4�����7� t2w�e(��q�>��������[@�+Ǻ��ey�b�J���,N@�/ny� ��-1�O��=ð�r��;x��	L8�����ߖ�݅�X�7y�Z�ܔpgc�H�fF�qh1?�KJ�h
�F.A'�h����9@��m�Mi���P��Y*��M�{n�x F%�G�;�ٺ�҅`����<�x4��G>܏<JY˴E��V�T����=��fƙ�#g~؇��/W���U��e(���ئ��m(}:�<��s�=~�����ՁE݋C��2��KPנ�.�ڦP�0�������A�@��}�ª`�1	@��}�R���8�OD��L9oV��	B5�F$k�C�!��2�c)Ý�z݇<��w�Q�Ez�v7Kp�J@��.�O��J��;��ſتh#^�%��mi�4��� iH�����U���,,�}�B����:��7�߆�R����թ���iDL��Qt�Z��J:����cL���<�KT�����	����n��[�@�~��"f ݻ57�VP�*��p��f��%8��^��@t�
-u:��>˻���4x�ds�\��o���4E��1t, �l�5�����3�]��r�,Y%=��Uzs���%�2����B	Syp�vs��ޡU
F��7LE���}l�bq#�l�3K����T�Bt�a����z@W���y#z;�!�Z�ľ�����΍���؂��hd�p-�����XB&GZ.IqV�	�.hT��M�w[oԯ�)_pz*�=jKr����R��u,�a��
fN�e+s#iOi��3�yXI�Z���
�q\�̛��m�sAk����-'�
���D��&��Z�?9��L t�^nw�X��X*����Zn�\��-�D�/��d�-�+��q�Z,$q�P�:�XG���*-���x��5��7�9�w�[����)�>����}��׆Cf���2���`�H�����J3o=��L���h2�������&cC� 2`�ؐx�H��lO� ���4�����)jWy֡����h��M�g�O�j�Tv:|�g_���R�gX�s�<����ӂ��;͐�:[((~6ｉz���!��>�+-�����ī�l��|����@H]B���>�\��ckҙX�ƾ��:���`*�n��q*����Vȿ��Qr��&0p���)|��v��.ҢyS��-]��5�C��\5���n�F�կ��y%fd�`Y�;���5ѪI�������E��Ż��ϴ*�Rx��>�V��]	urB���i	!��?0x�8��X,܇L/��k�Չ���g[À隤��6V�XN�/�@C�|�]?e�s�.ւ-�J����k =��?)�0�	��dS,�B�f������<,��a�#���8��q��i�pZ��O��ƭ�����5��TXz�U��xq\�ߩN����Cٖȕg/s����˺?�P<Ġ�>ሦ�D���T�'�3h ���O/��˕�p��?�[斉��TX�18j(Wx���l�+:����3eqf�(�E��ꍿ��������}Δ^�\�%����8�rh�k����Mc��c�wH?��r����˵ac��+j���@��XY<���{�@�5x���2(�U���X�^
�)�k�z"xƞZ�Qd�cZ����l�)$�T�,�zAУ�7�����U����2�9���%����������'��b=0<�E�>�->��ߵT| �&��Ò�j����xGE{G�n'������A"��g���T$v\�3��ut��E%d��1����>�C��<�h��n�����Pgt��y��Ll��1"�,r7��0ZhN�	D#~턯>��x��SvR�؅q!�Ě�T��|J�J9��Գ=&e���UJ�	�&~=��8�!�:��7+�po�B����K	�@|��6G��m[��+�Ō2���.)��}x��hrms-�a4�O�"vK7ţ]�=�q�]��Kd6l�q6n���5߃�ٙ��J�9�F��X���3��j�Q���*�]N��Џ�pc��8�l�+=:v�	���(;\��(&Ϣ�~����1��<�-��C�4�)GR��}�{��3��;�h$a��W�6A	�<�|� �7 "ؗ�[���ԂM�3�:u.�A���~>l��v7t�Jʔ%ndԪ۔2r�m�j��X8|��	/���%�^h���ct�2�&�֗8�ڈ��?�z�Q(��K��e%�l�<�,gH�"�W�y��J ��R�<�8U1��@��������@KZ40���:�Pdf��͑��β�����t����U���(7N[�r!�^Nh�C�L�9�i�A��Ͻ�q�!wr����u���K=�����'�]M�.%�����a���Ä��"��.:ծ���2 #���ʐy�r��.7�\��� ��xe�9���L�5�0,>�3A��ߡt��#}+��@kl���m�z/�r�ݟ���g�n��I)X�g���J.���-����|���3�#B�a���6�܌K�z���҈� �Ȯ�>Σ��40�M��j�"�	����/�O��F��'p�
w�^E�B_/7s��a��`|��Z�00��/ f�s[L^P̰PU~�l�&������H�9%��a �iRl0�VZzO��OG�����kE@ [g�#�����ަ9���̚Ο�W.J��I�o\Q� [��6���W�C���'8����Q�¼����Ӌ_O1������:u����Y�b�$k��*�t6X�`DN�5��"�L��R�4�E)��9D��8ilT!}�����f����`�EK˱<�P�]� #&�4�����pp%L������F���3��澺$��'rS��WO(2VV�ذ��V��.���#j"-O�?�����D��"����] �(*#���&dV�e����p�K+{ZR�;�`��ҟH�^�X@�^��.8ϴ[�$<M�˛���[��8�G�o�>��]�*�~�ξ�w2"�rt�@1o���2K�cM�(�!�n-tj�2V�(��^�h2QgJs�8�C�@rT#���6˥��\i�K�J���tM%D%j���&2�6Ŭ�����RJ�������D���q\�8�ʆ����K�R���sP���2^U�=�m�����Ĝ�5�8z�&���X66T�:�[v�7:��Mb�(a*;�b�˓[�L�>�oI�#��E�Ȕ{'���C������C���T]Vt����d1~f�������n��T^H@�q�z�S�^0g�vs�V�����@'�:�
 k6$�T$?4�Sw����D��o��XN�:Vp�׃�4���fr�8F��@'|[E��m{�I�g�F�ì_�cܫ�=e��v��IWP�㑬��]ȕ�m����kd�L�+E؝��j��2���l�-����t��sJM}�#v<��A�p8�c��M� 	����ӱ�yY��� ��A}��ɨ�L�)/�{�2r�6�5Z�kbw� �*���hAH�4�8��0����B�m���tJM�HM���Xn�(��͹�����k%��K`g�S��_jrU�r�*�v{B�<m��x���j�ߊՖ���C�:-z�P�x��[�[�N�n3��G�	��]>�G�
�-�
)}W>V/�W�I�������ACO�R�uVP���.�M�K05�� ��E���*[ج���q�Z�xIs��4�x���0x@��P�����末����z\͚h�V�H ^�SN[q�i��` ��1�g�W�^A�� a��̎t�<�	ai�Zfe}��J�����i2 �o��I�9�z>��Cw�b����e����(�@`�u%H�	[�6����]�5�yZ�.��Σ�����L*��U�[�[���[6G(�i�7ay'���	����_�l�#���<���X�����8�;%�0�t���#�_���s���������W�r̈Y�;���#���D����]	���e�����
K5��1��E��E<Mv��L��	����C�DI����KV{�)О��,�K
�ŵ��gV ���۝x.v�w���@s]Wܻ��m��D�َ��č�������z~r�1���h\���:� Y\��?=��h����TU;�G���I�v�m���X��Ԥ��ύ��n�HSk�� ���Q��3'q��V�\"�b���>�"��{I�i�0�A2#Ԇ�wiJ�mtr�����so��|�}�~@S>�1k�j�vn^O���M���q�YUK�󮴃�:��
Igj_�����㪁��a��Q�H˷��7�y����:�2�cI��� ����$�
�d.$�哤�F��Xn�kIQX�g?qp��t��	ۈ��3�m9�<i,@�h6��!rd��ld���ÁQk� '��SDo5f͒�6Z��^v�'��:G�D#�:%>[P�ro�}�c@f��֒S�r �C&��.9���g�FM7�h}l|y�>�E`�w��q8;�jn�ۡ}��Q!��7^�guu\X����L5T�<��;���vץ��S���=9郶P�}0�����b~��Kj���ٽ�̹���K *D6��`�W���K�Q(:�h~��eI%smo�G[TE���a*�O��?$P1_��������͑��&hև�s0�)��B���F�v뀚i��{��NY@+/釣��\g�Wđ�,sSU<�ý��N9o��G���[={��6��߽:�2.�,Uvn�:a��i�u6�(ge W��J�ѣ��d�'���+��׈隺�eW��й�jx���s.<{7�TFVw�NC�l�t�[T��=	e�i��� 7�86��B����"�<�$�8�}`~��j�vXZ����ȧ�~K}�Ǟ���Kdhp�V#�����/�Fcڝ�:#��S��lud,��_i��]�p6��%-��+KU:�˙ �`s�����l�8�v��T�\dSӒ3�D0OrUGGi���>�4D@�(j�3ԋ&~��"��E�,F���2�Փȅ�IC��ge���K%֓� �+�Fz��'�ͪ-^��������2��_�U̪&�6�);LG:d���[e��v)E?W��s��Ku�dBS#a��o����Ȥ�3:?J��������I(X�eڻ�8��ifn������ ���F����ڱ�ԧ��4���OS���3.�%//�:�,�"5i8�e(�;�>��C�����3^骕�|�5��,u��)ca0h�4��=��Mf����&U�
T?~*�E|5)d��C�8L��.GAE�\G`�+Wtt>��C�r��=^�����<�۾���4�t�w:�������A�8����ȇ�^�[ͫ�e/^tU��&b��:�W� �u$ܕ%�بPtı��A�Y��=x�C3�D�{ޭ�b_�_�NbE��B��HWZ��do����
�*��#���B}x>�dr[��T�%��QA�	*���1cS�m��m2���T��_O�"����6k/�t))��"9#k����iS���l*� Z���ߤV ]�J������&7�����Ԣ���7�A����]7�깚 ��&_��w]�HKh�%�	�4���Ef���M&�J)"�X�uV�&�/?[�4@{Z��,�S�&�e�Y��0h��v�y�FlP��2��Q�޲�U8��E�#8 B�,!��Z��V>+M�bo
[b�:H��c��[�T�VID�N$v[tJ����n�� �&J���'�G�m���&t/,H4�.Tyuz_���D����4a���0Q!*z �";�y)k�`�^�a�� d9U���i�����>;LC�g���$v(+�ltj~9�������Z��|�a��V{��e9#�ը�;�J�7U�1Ԇ܇1o	Y~Ŏ����LA��"h�o2�$�fK�k�UÕ,J��"��ͻ���̩O	$BHA$t�+ƣ�7׺��V���̒[�%+*�ɏď���ldx�4��Ũ"F����=�V`�}:�=�saAQ��oz�M���:�e{eL�����'8E��<��Bە�tU�:`�+��Lb���Ra�A�t�%���ep��&�	[�F}ɻ}i���=U}���!c��?�%����ch�����Ԏ�jE�6�W8X�k\"����w�E!�ɯF5\p���"��.�xĨ��P�,:���%
�@P�sC�l���#�Z�w:}Q2_��D����<ro��Z��O���	�����d��xS��P���/;�	�W��ae��񝜑�8������3y�X5����ʭ`���I�^�H��	�&`f���U��! �(��F{�Ӿ/"֣�{��L�D���y��NVcm,@���l��iH�_� f��W]�F\�ЬI��x�g�<#M���sL��|?���|}[�<4����P�,����C�e�DƮaM9���l���[�ߩ��_�V�� Yr�/].����������Q}n@�*�0"��"{���^�2<�������mA��L�qL.����[?a�?�ꖒ|H�b����lKp�<�Cnz��	ɐ��� ����$;79M�F#������H�6-e,+�KE�	]�++�GL����	A�|�����;�IZ7w�נ*K�W�. ��1jg`Z��m�X|/��v!��^�b�(/�s4hNv���i'i� ڍ6�	�?G?��3���|�/��k������q������"����������H���y5a?:�Rk�,6}n��2KX)֫����h�e���Svy�Z�[��8ք��Zҁ4�����{��;L�5�ed��j�md�P{u&kN��	V/���;7Ie[�g�X��Ќ����2,ۜ��RC�H��pه2�G���G������S޹���55Q��o��sN�,�t�hGv���[T��U[*�QR���!��Oj�?r�ăb��~��o,�/[g#���tД0}��V�Q|�G_��?��ǹ(8�?aһ{`׼2z������� ���,N����"Z�&��U~\�SQ0;��p�'��"�H)�:��1�8W;$n��BEFa�������y錆����ߡFF��D-hӄ�.ء�	X)��U?�����s�P�ј����bEl�'�/�sb�!��`%6�ma���X^���肖#�T�*����}��e���V�xm��%�)hX5S�_m���ag��H#W��GX��UH)��\�L��6BA4��[��ޅ	/@^�(��
��W���j���у�?��J�
�����X�z^~ #��c�������UM�NY'9
�`�=��f���K�"�0��5U�%M|��Y�}w�X�<���%T{�*��	(kc7���Y���|\	`*�/���`��T"�p/��C�� �����G�p�cH����� 
�^������xx�Q�G��p���%՞6�XcOL��+5J��-ډ�
ԎY��ؒ,/+�)��B�w��c�,R�d���Z�r���N��g��>?����=G���#����'��5h|��̜���n7�/��-~X� �4�)��Z�u�c��61艎�:��}]4�I��>ܙ�i� ����G�ޕ"}��U��:Qy�H���I��w'��K��\�|��u�^��1�K��Q� �΀�?�+��������"������Qv;�yZ��N%�G�Ɇ���-�jS+�_�;y����37�Ts�RkL�v�������?�wot�_Y�S:����7#�)��%�l�ugG;�Q�=����o�<���U)$l��`�2��S��������@�L8��A���A*z��`�����5�������B
uo�h'��i����8	���䴤M!0�9Y��*�G7@J�5�����9��Ih6������fXJ��L����N�2uy����J2Mڗc���������X�sNڎ�2�3��x5�@S,�;�J�#��7*
#yM�ŵ� �vHTo�i�N_z�XKk��|���5����3}`�E Ɉ���{;Vkf�Ԏ��O����7g���с�i�mTS7��,0�)�X��Dņ�z�憓0��[��U44/�=�4[g��+���m�L�� �H��U��le��5�2��ð��pl��A�	;N�����j� ˟�mݑ��I�h����񋲏U�� ~|ﴠ�Mhށ�� bJ������?$��ktånHB\��X�5f�c���d:�j:L� ~���b	�1�a���˱�����P��>
��t��2���H�5s���m�P��0I4J�#�1����.*B3P���K�b�VU���P� �x�K����.�2��ۈuK�jE�%ζ��^,�_�`�YB���x6@�Q�R��_,#
�x��t8:��^e��P`s��~��2x�l��0�S~�dO���&�,�wK���w�o��	%ܦw�h'���	�n�)���Ve������Y�,��̷�1��jD�f��T;��o1���Gy�_+"]T��	xn��-^��bե`c��6�����Efd�A��u�R�7:��^�� �tpUlK��L���o]xvݳ�{2�%�=R�b���z1�V�$@�%������{�߀e�z&�R
���Q�%NV�x�u"ڊ��]�����/Nm��,�8S��Q��eDL�1��m}Oc�YM�'gw�v�7�B/� �X��E,�)�A\��2�9$�6|
\���34�`�C��ƈ�!�?�`�)����փX��^|���V�Զ�<��6�e��3*&���U� A�rhu[�%ϰ��r���V�RQ�������yzx�#���?b�Z�ʔ0�sp���^��ޚ�A���=�#xUG1����/Ysq�J��T^˒Z���WX� �8��Lv!�YJ�X��� �y�I�׼DP���^�*��¡����9�Cł��(�7�5�)�va��M�L�G�uN<~�~-���c����)ʓ��(� �E	sl���}��x\c	��g�HQ~K��GA!��?�jR�c��8+���r�Bu�c7k��3v��9_���a���M�
B�ӓBcAC�FΤ��Ձ��������U�y	�@�e{i��3'���hu7�pDM}oգ�������MKO����(�{�F�r�"{SK,S".'Nf�GP�"�*��2ɘ��ʿ�g�	�3���k�>S) ��O��b��C8|!��SU0w��[�/�/ݴ�P`"���ce�Ԟ�����hZ;��FH�>�6��$a������=���&���{���6lAAh�L�� ��5�?K�7��@�fsm�Fٖ�?�BJ�p�y5Sv ǰg�U��E�+;S�NhLv�{��B��%����^@y�nv>���AL�����]ڴ�T^!xo��L���!�w]�_n�e��J��b`b rG?�����V�/�C*U��&0��`����NDM����a|���63]�sش,��p��Ӫa��-�&8ٷ���2H��<jXIC m��KpI��E�t���۫j������F�-���J��~��Hc�5�s�U�83�"\��(�T�����zS��m��Pt�2v���G�7������p��$�+ܽ��ZT^&��Q%�(""�$N�4woB6�žg-J!������oa��C�Z���4�-K5�C�&�YTr��ʊQ��������=������h�J��'���U`*R�Xd6��9A��mȕ�R�
�a]MX�펋�-��0��$PM��A��C+�ł����F��rJx�f�+9q�ݾ|�����2����2�f�����*�_�5��5J�?;�5�4/����eBt�N�L����[�u��.R�2Z�r0��Kd��sO�����l�x?�\cm��������qc��=��]�p�2k�x��������f�(z[]:V�Z�\������d&Ke�$�X�Ps �'n��Lf�=�,i�X{�z�KDC=�(���Ζ���{�
��r��W�q��	�eb�j�̋�����GZ�g�C���������!� ~��q�<�M�?�O�[N�o
�|�[O��1����N֢�եp���3} w�l����Jv�Y!��e#&Ja�e?��w�͹�0p-S���ɠ$��k���S�����å4��ty���},��F/�XfogY���Jђ������t<zݎ�`dz� b#�H�'�� �a ;Cl���.z��e�MP�rI�G�sb}on&�Έ`�u���:��M�K�_�������sޖ[9���c>�v{�]~R�a�~�3ߛ�c���PЁ������B)c�!�U7߁&T�B�����הpp�ER��0�X�e�S�+B���ΗUD��H���L�� 	_��1%*;T��!&�?})�㻶��d��`��������Ȏp����r���mr��t��gu�I�Qk���緋�$�g�̜���%$/��
��U�=&���9����b!��"�|n��.,*9x�%/�xI}�h!vG퀂���h�u|p��O+NF%#�`01q,�a(�p�3O��e7���u�[�囅=a�gD��?2a�g��Ɍ�5I`��D-V� :[�d)�=���;���6�`�suז\D(��������B�yef� �Q$F!neu!�z	S÷H[���"QMea�j�{���(s�}Io�f�����ʿ��76�	���t]��}|�&�Q��)=����()l��N�*�+�$4���?w�8�Dʉ��>���;`�	��Z*�1
�#���݊�`���y✀�`P�S�Uɠ]3]�.=��#������ p�"���Zb�4�tp$As��Jt�Fr�2ga��}󁷬��msQ'��*�]�N���a����@�Cӣ�o5׽=������X)�/�C<q�. l�+�K@H9��ABO��v�E(���yC�Z��3�Z�j8G���s |�A�Hm��4���U��\I�-��t*�0�"�9�n�d�H�,�{�'r����g�P�����%�2]l���vgIT��o����rO��
W2��*�RoX�.c6˵d�+%Q.�BȖu��(�Mh��O��)q0��+�Ws�r]tv�І6������p�+V�����W���,T�G��"ԟ�C+[�$�x�8߇��cZ�~���w�g��tm�Yj9u\=a�]�w��e�q�-zE�3��6��t|ޙ_����}�S5ONkN�|#*Xe�oq�I��t�*J��DK]���q�ʋ_f��L)[?H�;���l�2*�a�W� �;b-���g� ���/%��)�Q�_�)%t��24I�Al�X�#:'���l��Xf(��U
�0�"Nt�����̄�x-���)�V޹v���4��뱉��x�������p�c��	>�������s	��SG#5�[����Jn����T����O$���0��}���|.%~�3g�vEB��{Bc�	����S)�A�v!8�[���3k?�E�c��n���aT�������ɡ��*��U���qj���f6K��������
(0ljF��j�v��y�E�K���O�6or���_+���d}���<���NN�:TH:��1�Ep�ܬw����"樮]jX�(�����g���a����"ʻ�{�g��!8�3R��0#�MU 
����?�Ռ-���Z�rO},�׶��Í�I�u�'m�Dת�����j&.�C�ո�����A��Z��]��}�$Sg�]�ǁ���~��s��'~��X�46C0"����ġ�Ϋ�o����!`����!��e6���}��� _��Id7y�NjC�%�JE�t:Q�<4�E�\�3,)7J�
O�J�X���"k�h��o����cK;FU�J�Z������������1��-�A�`��Ɖ���#��<�ʸod��=�-uפ��ݟ�R��R��B��,�w$5.G���ʚ�Y����]��
i�Mi��&e^��y����5���ɸ+�m��7�G��UK��]d'�06�~+Ѿ���d\�����,�饫42�l� w��u�z�tKR\9h�j� "n~�Aj2Mƅ<��]u�w��V�u㬽�� �Y�i F.����ց��Ǝ#��>�6�o�p���M�@9Z�z�뽯3Ȣ��@�W��JȈ�s4"�̐N6t�I�S�({i�~�8e,�09���B����:�8�X�O,ݍ��K�(ɷa�rh�(u�_i+����t�L�Af2t�(A����N-�Q�Y�
�dI�8�~jذ�6�3�  �b*ȸ�C��A��cp)�A����$8;���F.w�}�0�a*B.vz�.��N��t �"�jx�u'�|���|������%� �-���NY�6��Djz�T�iT3lL�ёޗ 7Wz�Cq����8\[r�!?��\?�� W�_��.��.jR�#���Ǣ}�|��_x	`j����P#�
��W�I$�_\Wmv�	��g���L~lX���w�s��p ��F(�\>��*�T�k��n?�3�7�Z��,�E�.X��۷���R͞�7涳9�F��v��T��"j\L�(�m��.�5S�	�خ���+c� ���A�EZ�b(ǒJLV���oN4��
4us��Y^���{�`NZ� ���zÚ	nA�f	��ܻj5س2����sMoqÄKY��R\��+�^�sR����W��'�]��������#-Aɤ�I��0`}k����U곔��~��fsX������+zR~HP����^�/����q��8-k9��z
=(iXM�-�
�Dw3}���~Aɻ���~��Y��C�m�� Â������]"�>����N�4tp�� v�&��:C��^�_,����㌖�j[�_�T�C$��[xH�IV�}#�I�aˇӱ�n��D�y�stoEa�v
�0����.]���E��8�#hG�:��e�&�HY�{�w�s����?1���ZT��fz�!��L�1�򁩣��+a����#}�� �N�,�9�U�4	��.���Ց������1�B��+G/��_�����-'mn�-����9��55���w�t 8�z��d�����S`+������4���	r+�:��%�&dD�/H�(��f�8h�v�cVAw2/'��ɜl���p���Vw�䑪:��D\L{�R����X�A�e9���ۇ=�C��ӂ���2��[1@�&���!�ɴ�O�3+Ϧ�	C�@�,��1#���>��%�&2�~xR��fB`��W�XN^r�I��9C����������_������k�R���1J���;9�T�tY@ʾ���iv������V�Kᗀ�Y�v��k)�����v�V��c�9�ˤ��,M6�׊�ŭ�Hz���`m(�8�����g�Ab���=��Q���Nu�ڌ�h�w�ZX��9si�ʵw�j|�G����z/${��Q�P�~����o�OAHd��p�t�n�[��V��w��ցGZ7�akTX�#�ϙ��u�8c��Wa1��ؔ�9�o`�lf)����1t��F�ט��&��[?u]��N���BU������&nQ�� �MCח�/lW!^Ģ+�����5E���>���{D]�9��Ȩ��OQ��i�k�:#%�Y����Y�����ڎ�t�30�>��m����P8_nx?
r��?�>�W{�9M?�A�X��}QP�Y���e�(^����ڔ5a�T��7���) ]pd9�@�u{]��m��0�.�+S�t"���H7=N(#��b�3�Oc��J���B��P�=1��m�G�H�>_�P>-�绤��@�xv����~}t�_7�k���(F�L�m58���?�(����Av�\�*1=��:*����[a�%��>�����<��t�v�j�y��
5�b���Zɭj��Z���=��E��(�6:�r4��l�gG���_��R�>Ҕ�K�<���Q}�]�e��/����\�������%�?N��</�i[�Q���|�j��,�7�^��1��\ə-� ���s����FK`W̽��,��9Ь�s:Պ��$j� �6I@��{r_� �rFx>��4�u�������'W��)�VוS82����,:���i��R[�mܷ��2]�Y�s�|��d ��|�L����#bi#Y��:�%^�z�x	Ѧ3(��z-��g�35<�Gd�'.�{��u��_m�Ila�!��C��YOq�R��nAw���M�z��|q���|۔����d%*׿ �CcXM4�ݸ�б��K�잟����n��ॄ�������޷�f��q��3�mw��(�V�/�D��Bk>��[�Y΋A��@�)�D��}3x����Dq�@�7�Y��w�c�p�f�˓��ˢa|U����Vj}dZ��°-öPK���O
$2���B[VXD^g�\�R,_b�)U��eXffPH ���;�Q������(��֪Ufh�P�.�Q��Ev��f#͕���X�͙��/�?y�#@�6�{a�!ҿ߻٧�j��%ں�v�*Ϙ�ǿ$F����K�.���$�|�'ύ �w#�c���S�p��F�<����o�� G�kw]����K�n��3����;��G;$b��� ����V��� �+>��53^8n��������Ȗ�Vn��hK����Ϻ��J4�ds 9n���l�2#���+���Hڧe1>�]n����.�2 ҮK"������o�z�x�/�����`�R�T���}�5Hګe �깾�6���r��3����9��M7DN���f��=�!uX�޸J�����@3�L�(;g��N�Bs�lTo{H�\��1�#d%u�Gb�;D���ᑓK p!�idk��В�g�7��ݧ�L=l��`��xT����d��I6���Q���RG%�%�Of7LA�a2������TӬ��)y�g�GK묱�H��湄���Y9�r��0Y,���ڬ׈sL�\��"~8�)M�NN'Z})ä́�Ė\��L�a�@`�)��4�~������W�F�m��T�M8��^Jw8@M5��B���8�{j �r'��V�*&�)��TؐJH�DՌ.3ġ�S۶P�?o��w��Q��{<j�[��[�M+���j�ߓo�R�vP�Y����b������ il��X��3�׿N栾��| �r�ղ0��Zj�[R|�{>�MY~f	K�r��9�ʩ����2f����}U�[�3�C�a�x_7�d8^[��߼ w޸΂�����3P�oW�sw��-D�������$�Y0���?S���G�N�W���ٹMఀn�t�u�-�lNӊ��]�e��'A�7�L��Ԉះ'Sm������D��\��r^�[���a�� �87�O;Sպ}���j�R@�"���c�~�9��2삩A<�`O�K6�*_P����"(&Z��f����啀��SGA�&ձ��DH�R1�?(\^��o^��7�W-y}��Y�QS�mQkR������>x+�}�Sp��~2���ß�ﬤ䤪tia��7��W���g� /�f��F��֧��Y��&6ocɿ��t��z$���$$m��ǒ?֢�	j4�;�ˬ��{|<+Qt�7c�*�ou��xD���hqP?ᶀ�b�h�aQ+�9f��h]�_���Ğe�)�J*�t �/8]\�L�$\�Ikٕ�Y��F}�®�Ľ�"@!�!�:�a0�j�F:���U:�,��C]pԆ"�F	)����w�ѓӾ��9�a3�`��%��y��mI����aY�L�9a��'��E�Zͺ��t��m���6K>ͷ�$4��̻d@A���?�<���u5��/F�u���ݹ�v*1��Y� �l��j/&��I�f��̕�o�a+���=���;��.�X +�����$�4pR���xxshR��>�n�]���M+i�1��O��K̵1�	��-%P>������Z䟗3��ܦkJ1��C5�C�D>�r5�.���c�^d'듦-�����p�V���$���D��_��襻��L����q#&v�E䑝��rȒj<G� vRGU���6�S���Ǔ��db���|���	�.;%yPJb���K:�7� \���ٿ����^�a�Y��G
�慶<t���cmk�."sm�Eσ����uQ4Z����g�C���Qʫ�b҉�7����u�q/>V��u�PH���l�p=�u��e)6�۳�*(���#>B�ƶ�st*��>Ͻ�"��߂�aOV�5�D��<����1ҧIj;�T0��� zp�t����T����g����=-xI8�O��+�<��J�R~�����_dRԏ�
A�и���B���o�?�wy�)~/$��I��$�_N�Sn4��61't��C^��&�y}:��f�"���:y�U~����X���)����|�ߍݶ�LL{��w�O�-'� �8p�N�����Pq��x�瑩J�T�/xٵ�k������wJ�Ջ�_���=�0��*��L�勜*Ϫm���b���dHS3�Y!\J����_�ᔩ��%��Y����(
w��R�2�;��^��#�>&�;Y���N�86E2}�LV�r���#M��}?�x��x�����SL�9 �A�+�8��(Zn�[�[�g�%�x%��2q��3��Q�.I�{��]Ы�n����=��S�D���GR�����W�0`h�vk0M�DT�m�Ρp��U�P�(��0���)�S����p^E��	b����!�k.��{�@�0M�Э�{��Xu�d���{|���{�j�g��Ȉ�D��gԴ�vu���{c�{,%&����BGv9$?N��Ja����F�y�RTobaBI�e�ߠq�����uJn���2��{�[�qc}��.����g�~Ԧ}E�K=ĄN.�Z��oI���:�t�v�;` ���{�G�N�T2!A�;�������y�[ȣ���LDX�T�֒,�-F��S&�:Y�}d�>W>O����s��:�����_u��L���S�f�u)~��t!���?������͌��/��b���s�F����m�������F`��qA����3Q4�	U6#��#�w��*"��\�<t�z���m٪.n����@X��\@ww�m�m3+�}cJ���Z(MC��Tf����D�똭M��U/�
����zT$�n%=������ГI /�*"ӷ �ְ	�XV�l3:1��p��K;�&����.2���X��;����C){\�Lb����ϋ���S�� d9�,��M����L�'���l�X���6���{L�=W�1�|Ѝ%$�Fa�I�҆F�*�𪫓�/oN}v�����ne��'��Z�n��z箿S��I(�B/X���L��[rN	(�����$��BL��E�k���W&c>�Ф�~N��`��!������ڃKj��5�t![��"P�٬@��+�J���Z��/��$P�B�E� .4������K.�)��uQ���!p)�<	�[
��ȼ� /k�-�i�>J�5�����-�ܸ��.W��@#�t�q4Y76o��i�Ծ��yXXs���>������B����6���>��6�
�{#{�'P���xJQ2pGo:���0�݆x�\�ok�6Mz/��r)?�@�ͬ	�.n�n��[��ի�[�@ډy���l("���C��̃"����M��d81���c�q�w~�+v�m� \pk���z�~B�ĵ�)ג��S#��b"�����PD�ԏՠ��= |��8��	:��:�(��V˪|	3ͨi�n�Fڜ�J�H���n�ͻȃ��d��k�AD�����j�A�.��Ȍ�1��U�D� J������0�P|��ny/�YC1�z��EV��j�`_w��UH<��Vw��ud�O�4 ��P�V�,�i*��L��*n�ɒϱ!�a
J�)o��S�����*��hc��1���6�^����F5��S�.#���v.ˬ[�kO�%O��@q?�c��@2�Sf!���@I�aI:���%�d��u Ҷc��LD?^�9��%���Cr
�F�6i�����ִ.�]���j���+���"�A�=ZL������n��p4^�3�u��p�i��D��o<��	j�?���-�������.���6�^����A�^/��ⷼ�Ke��R�7
N-���ţ({?�\����R�v�&���yFOv�XEG�:j,��25B�3�[�%�Q�sQ�S���=��.)PDC�Y]�P�Z�1c������6�-����1��z7�R�[�Z:�RH'[����LJGȽ`��o��s!?W�P���iV�w"�:K�x�45Q;Tƅ)���XXD��ہ��+t5pp��ô ��`�hP�kd���ʽ����)�Q!s��l<�þ�u�^�i�r�	i)0�!�21da/����a��kϬ��
Cy��{o'@�"p�Q.���Tc�Ȅ�;3R��|�1�<��-e��-��P���l����GRi)>S��Q ,?�׳�],�M�=�q )m���I�T7�_�?!��k)|��U��gC`�`1!t�c�D��������	�1��FGJ#���t���m���	��E�W���n��R����.��v3S����������7�������UP�D]�*� F��d�׶����֛��S�{���Aҥ�g�"�'�X�*�j5�Qw�n��_z�R���tl��=�EWd����d������`}�E�*o#Wk#f`��/VY\&�<ޏBM��f�y]��m*�<���e�{.R����h��j䴶�I� Q�B4N�ʸM���2,5A��P1�x��jg�8�l�8��D=]�Q��y�O�~�}٧wb8I]�}�T=>m+y��KN8�R�L=�RlJ;�����R�  8��A���:���/��$ń�6okd���#�,h��϶�����nj`�-U�ڡ�I�P�q����F�2])���_��BAY��N���?k���UqQ^�C)TC�a�}�י�!� ��R��V�������-�S�j?���]V4^�w}��():��%�*HûRѝ�za+v�	Ze<x"�+u�B�6uEWO����8���x�:�)-�Þ��Q[2��VBVX�2����H��ҫc�E��2R��wHr	��Ֆ�����`*�K�T2�\�|��jG�ga9�����[ݩ���49��H\������wsf}�Ǐ	�M�+�K�H�mr_<__>�\�((�b]�Ұ`u�
�A�r9�')��T)��|V9��L��@�yƘD�wyC/pq��*��J0��ٻ�ū�@��eq�-�{�]BǬ���&�z]vo�Z\ϩ�F��������ޚ�;�%m:��܂st�;
3]6�NԻ8Jt{���0{+E�a������"�.�Q.Pc�(M]������2ͦ@��Z-����1���q�6`�����?��\��p�y?v|���1%%@$m��\m�v2L<-���(>v���
�	c'�㇞���Di�?��v�ߌF�|�1�D$�����YI�����O���1�9���R*�\yw�P)�P.�i��>�qm��F3D<S�	���S։ƓFx��-T�)kP�v�ؔa}�	.�Ss�G�aL�/�lJ�,8�=g���R��a���	�N�8�wUH�d�l-�5��XSa���q��(�Ց��j ��6K'�����B<�&70p�X�h��|��`y!`�q�q���e>;t9��BA��K�h�,�k@o9����
Ƀ���[a�ݍ��׀ Cp�G
w�C�Æg�Ũ�*UM�W��q�]v���͠��`��>��+����m��R ��m��6�G�������潳[�|}��Wk��1���*�n����wl� ���P^����#�v-����I�m ��W����V6|_�᲌0o�ꮐ�����s2�m6� ��g���u-��&��RC�	�oCZ�����p�?�q���;K\�N�a4��X�䙴�2��ȉ�����0�X�M�uį��S���J��a�q�+�!=:���^ؚ}�,����L���[F^�� Q���=�^�́�9߼��4c�b�եz�?M�h�eů�9?��:_C&^`�����Ԫ �̖)z�yr��#�ǈ���H�+��#�8�'p��Q�稭'Q9R�؂>!�缃��� c��La�@ƚ������Ȱ��Ј����Nr��2*D2?0�_���N�d�k��F?K9���"R7Y�,���K'PD�(qu&X;�o����!Y%j��L���6��:��dP�G)ެ��d��(������ؘ�t��f�Q�l����ԉP?J�1��\�,3�zf
¦�|c  
��Ǚ�G��	ݞ��F{cU�U���B>�(5�[}ü��>��W	�˝%���y��5Q�v}�B��0Uh������O���8�S�޴�P� >�_2�ǝ�AD�|q*~lbE� "m\VKҐ��r�h�!��K%<O�q_�R�Z+��{�vQX�{�LL�eW�V����/�[V/���4�.�0����ʱ���k� cx,4��ғ�(i�C��7��4+�p�H'�P�����X����4�0���	���MB.&h�jg���!!j�z&%.���}JO����! 	�u&�=y�G*(��qмY3�F�&��Z`t1_å}��@"3�>�*Ƅ�Ѝ�L�tV@(B�/�C<"�׷�7�n(������E������>.���:T�GZ	.S�\9��G�wxᔓҗ�;�i���2<�CUǜ~�x��yD�-������逥����/4!��ɫ���ʚ�!%�VX\YL�滱��S�-�i�wH�e8���D�Ca��d�lQ�;)�n� w鹳�ԡ[��|���i��l���$Z^���<��G��36�!��踜?y�w�^�pE�i`/�C�� �m�R��r�����s�!-�O�E��|~8V���_/k�,�#� �'y�2I�?��l# x�&C`���C
L���������&�4d$|)�Lr���<�" �l����)P>d\W/�zF�^f�Q� �	��B�f��p�a���'2�B�6FU���9S���g�&�$V��=�b8i�;o��w��R!g�[Rl�p�Sj��)ϗm����D�oP-�ۋ/�.�� ��<�)W�u�I�Ut�׼c����~P޺���Ǖ�Ks"�����y��F��O4�B���VN>� (G�����S�����"�B�΍�<&�r"}~�iP ��؄�	"'���7�ǰ����-}m��*��;u���^�	�#/R�J���q�sA�4��z�"3�M�K��r'Piš�7snY���/�3洚֒�N}��%�b�Y!HTs��<��j\m�x�6&ſ?aF��D���a4ϖ\`�x�Z:�5wZ|+�[i�@���,'��D��f��R~�a� `��aI�#-�32�GC�VoƷ@�"ue&s��C	W�\?[wu�lӆ���]�����ˮ��5ZR��ɟS �GK�(]���q(^�H(�H����T�aÖ�݆��S)���:̇�l���V��#�c	1��tJ׽�A�@p�f�ʔn@�(�ӽￏ�E{��=��?�F(�H���j���*��J�1t�|hv�	���{{���͈m�}���l�k��:�Tw����!#4a��G�l���7��f,j;������Z�lc9p�U١���|�ݕK�teЩ��ƶ \;ٹB���ҲV�.���ɬ�u�jm`���rf��{�J�+�����n��P8��$�,yGUr�?[�U u�z���Fl�����.^�s�� `Z!_�VDH-�*��g���/��&���&��$u�Dؗ����E���58��0��xH���3!����E&,U��WS9�h�6,�	-=��l�`u�q��r��#{��|+��\���4F>2���:h	ƯPX�7�:�Fz�g�7h��0�/]��X�����ܙDk�I?9л��Z�`�HJ�pfŋ���b>��m�oC�L5�5���(��<r\c�'�Cȗ]4�J%��kJ1C�JA��u7�����.�7&KW\fӫ�7I�O�>v�.2Ϲ�]q���&b�Y�v���L��=&�A事��1*d�e*���bKar�gK��%[�	$���)�}�".�����it��s9�O0�#,/;/��,�N�Æ��I�/���*�͗�AJ���|�x]F�w�&�q���%�E���sEb����էj�{T��4�6�tVWl�C��2�k+��/O(��^:�Ӑ���ĥ�O�(Q%N�o��� � �7m�	�]�~?�D;������WY�f�a��k������l����vu��Ή���l��Q��P�.%�9͝���!v���4[9���F "�����7R��1�����%����X�oG��{��ƫ���ߺE���|�|�l`�+���`uܬ&a81��Z?�Ȯ����A���q˰
��'���
lo�o�ZV�؁e�� ������Kh���<���PE�Ad��m�+ [x�8���Nk��Y���2���<?s3*=?�~�:!A*`��W@;�PRi��� ���s���.1�6y3?��,[�I6��H��G9��bSt�L����w��ip�h�]�/��O���|=�����م4����Dx� !��R��6FRO��޳�]��7 �D2'f'�I]�-�ް��)(A}؊�.�[��dvO�2������������b~�vQ�k���*^U:�9�!��)��/t1q1�`��� �k ,��7�H�����w}�}�.�>�#�J������g"9�:���<}�ȃ,�ܧ'Ͳ�Z�c*�{;����*���Ȕ�f��p�MKQ�i>�bh>��I�Fq��D��g��/s�bM��|��ܴv�s`vV���ռWA�p���
�4N�(���,���;I��Èo(�p�⠐Ӻ	Y� Ϟڛ��BYG�V��L����<)&0U9W6��(;�4�K���B�Ϊ�1S�.�������.������nt�vֶ�x�F��^
.}HT�^{��k?�&�<P���I&�F&#��?2��%e��ň|�>�=6u�)~خA|ܜ�%$V��.@�ؘ|MQ��;5q��&Iⓛ�/^�� ��.o��¼2����X���*z�l�p����[G1�L-��f �����cw�/!�q��9/�u����N$9LA�����C��:d�cWkQ܍{ ;�ˆ��/�p\f�93drX��Ȃ]n猗�~��1��e�k��������n�z8�|rit�l��/��R*�_�g�%�S9?�UB.2ڌ�g��x����L�P��luz!��cHKT���������i�r�K^%[�R8�S��*͓^D0GMA�3]�^�>�r�r��|(E�Β}|a�ů_g���[i�~O�~=#G�̾G����%�jL/ZY��Sb�{�+��w
���8�a�~��6�[���:�>rv��桬}��m��u)���N~5HA�r�Y�C�HC,��)N`������G���)j����3ٕ)�����|�2����0�WT�|�Mb/r�5J�=J�D����֣��U��h�?�8��E�����P��3�B�q���S+gS�%5��~��}�m����{�x�^k.�|`G!|$JͧOWo8��h'��f���,�vK��$��"��/���X��ԅ��u 3�-��Y��#��ɐ�O���7�m$�H�3t�R�]»#gJ	�WQn�H�̖���<�"I��i��]�[��/g�����٦��{�>��� ��γ����fce�ýF�
�1�ͣ����N˗+6=y�b��8��n�9�y�ܹ�Ƴ�Z+y���G 2 `%�(u��}�)��	h��bF�rrr� �� ��ل�Gx#B#i������ufS{��� J�i�Vز��c�u���Dh f��c����6�Ν�ȅ���K����B7�O�I8�1i����{�4�� ����d�s��z����8 ��{�A���ޘ����8�R�:�g�*���AYN}몯�e���8�1�uL=��8�~�7��&�����wg�i��'��������\ȮҬ�8�ټ��O��|�I���<�1jz�*���/A�2y�ӊ���ܻ��U����eG����&�����Ns�����$-�y���9��>0��M�윻�a�`��t�qt4Y�hmz�߲,+�*�%-9�Ͻ�Pʱ���nP�U� ���k��f6N/ �n�+AS^i�?�_I`1����&�Z�>�y4��b��8K��v&E����������iR��m��DS�S#S��M�[��N+������v��i�C����& �?๳�K�q˷��J����n7;|Z e��{>�7Ô��a�e�9
�G�`̪/��%W��?�?|d���[�܊��]_�-�fS�̾X�x �kwI���SU��m	ٯ�����ވ�ҧJP�\b�ᐃU!i��yy�ʘ`��l;|˾�;���2\YU�۶D��1o��w��7�NT�y�m��|9V��}���i��?2B�Q��^'���x�`u�Җz\Zƚ	U���<���J�!���b��&��^�3��2�ųX0�D���~���0��7ǁl`��|ט��LO�n�8al�`�*�e� �e*� EMy���H���D�:gs���Z�n�e����@����&�
Ĝ�L��x�\XZ~��?S�PJ����r��Dl�)r d���P�N�o �r��Њ��Ɋn�H�r�2�Q�K{Z�4�=��� �L�Y!����d/F���Q� �"�Do�+�>��4p;�Jc�(�!��ԉܤpPG���K�5��ÑC��A/[l�B<潑����U�z��J�������yoG��#&*������7�3��l{�&�n��0��W�:��_t��o��Su�Q�
�4Q_=�'�`fYX�J��|$a��B���������pxik���r�|zN��5���x��Z����
�5�2ir|d)��E���h�ux�ܿ�n�褔�Z�F4��, $ӵ�U�[Q-#��]���s�OQ�{��1�bK�M�\�z�z؀{(�F��g��a����RQ���+~��~�*�+��{H_�v��xj����K�TV%yf偆	}�&Y��2KӳG3�ͷFq ^P$����9�*-��lge�pL�����U�+u���c�� ��a;J9��.�Y��K� D@*�0
]��ńb$�U���}f*���œo���xr��08���o�%n��Tk���_g��rw����V3���u�ni�S��s���~��Ɩ~u:���.+����+rM��%P�af��>]��OL����W>��°��LG���Da|x).�����aD^��
;������q6?L�$���]�,#K�5����S� �j#U��3@��E�^�c*J��򖃯rE��3���m��^�q��e���,�@��ӇG,�=��)�,IU��t�J�yTG�q~<�2�u�jiumAjJ�O�}s�`��j �bDQW8����(p�X�`j&�g_V�ᡈ��6�jFN?Z���I���y �pk�KѨ�t�����[c7.�0�׋��Ix��R���R$|$����0���-�{�_aZc�ْ�o��r^��%ç����M�.À���|��t�7�Ea��A-��=pX~�kGn� k�� ���3t�g��ˉWj�~f\Z�K!�C �ɧVV��3cH�Ge�&��p
����eڶ��ܥꟘ���i�sjX�R��&��۩�9%G�%���NV��*��B�3{W�)̄.jz�E�+�T��ǝ�i`�5�3M��}n����0x��70U�Q���[������ �/)��N:޿�\��4_��1⊺_��:��Z�-j���B(,�P��u_��N���C�4 ��qvM�E ���y��� o���� i�-ڶ�����`L��l���ŭ��eѸ�*�]SK{�z�y;����5:�p��!��sK�?����V�) ��ڀ��3��	�:>��/�B���2S����Au��`Q��,"��<�Ɍ�<# ��>�>�^����nL>9cG�B�C���B!Ș"v��V3f����� C�̐���Կr�ͦ�z�I�@
Zf����Q�ȸ�~�Kݫ�vqRp_��Gt�\�����aX�k3��\W]�t>��*n�T�2K�Y=�C�ՈӒE����j�}̝~�3���?��SqI�M�X�P{��ũG-�}b������F���"�4����_�h�nZB�8�4P�8>��Zף����=����U��Ms��Ե3��YB�R5��-���tv�'���rK ����UApDMJ&�裉y�D�{����D�᪢*8 WHb�
��ǀY�UDG�;Z�b����it��5��
�a��)z"=��{�Zǖ����t�~���<N\M�.'�f��q�l5sF�K��gn誺�.�ec�G��OFʑ|64��lh�Y�_��%���Zl�BD���u�ޛ�!~~{V=O&�5�W,c"V�8S�=�8^��&�Y	��E�F�,��
��F ��mR�Z+�y2����Z��?�sV��aǹ5S5)L�{�w7���~&��ē-k�@�}Q�!m��L�Y�2j��-9_"^W8i���̫R���B�� �7�q����^��_�hc�߰s��݀���@���3`˿9�����q����
ό�U���1�A^%ن��1��O�v���&�1f�D
Aי ����h�5ry]+�Qr�b<0jĩ�����˽���N)7�X�} ��z6d��l	OcHX�����[ego�-�L���p���B�Ҥe��H�<�0gQ� �3.@�����6�ya���̄���l��V_����6�%��?���_2�<��M�8\���֥�j?���(�ZJ&Om:L3F�$�)��ȟzQ���R�fa�q���a��܂R��d� j�<�N���8?,�l[�я�;�l� ����{��#H?�EN�zi"ocL?#�X�oFJ%n�A.�s����F)�*�H<��&�Ͼ{� g0V�wJ8������tݧ# c"����ʩ3j�v�xs��\h`���vׄJv�X�J�OVw�2�vߋ�T���O��(��� �9]�Xs�a��π����5~F��(a��F"�5=�(Ds�;ص���D���d\S��Q���B�X㯈9B�xaZǻ�g��H�Lm�Րz/vO��Q� �� ���>U�_B�u���i����Ȝ��6-��q[��[Mj�aK�^J!a:Di8��K�1Y��Y$��o��,���kODW��x�Y������!4������H؊�	_��󈋥�]}J}�*�	,������O��:cV�Y���Y���\��Li�0��"��;uM��7º�{f��PҘ��v	>�\���3��=h���b�:�ԑu䘰�����G�̽�Z?���"�<g:�(����s{���c�����j�q=KI������5�!E6�H��Ы~�����i���0t"���g/:�	���ݓCdgH:�T�{Z��*��܁b�>T+֪������?"@]� ��ݷ~r�"��y������mRo���]��O��6#ֿ�=�K����ko�>����9����4�-6�R1��7�����C��m7�Eݗj�����Tѷ�U qc�)DOo��=��=ڎp�C����F�\b��R�NbS����a��׏ݮ�m�f��VY��^��?�nl��e��8�H��0k��@7��5XU�[��[6��}���R���w�9��O�u?9֪�2���1���k�Y;y�CUTdr� ���Y^�v��p�������g#�߸W:�]0|*�i�T��w�z��' �n­u��L֣��
o��mk��Sk|��]`�*�������׶��*�g�J��˔�������G��ej�W8���>6ʒ��G�I]N ����ޮ{�Xӟ9��]�r��W���,*�j��X���5��\ӌ��-G˨鿻:��q� +kդug�6�19]�|�C�w���M���q���?sz��yΆ�[� E����L���a�,�'����>6A�cv��<'�>��ܘ|�>(�����ڼ�D9Ϥ�s��k:�����u�����<yՃC䛩H�j.y�U����_,��9`��3�e({��O7a�cϕ�����ڸ�e��*��[���r��lR����
��`��H������k����x�D�)戕%�:&ɂ�_�u�7
T����^�	Z�n�0��+��n�K�	��}K)jچ}{x	l�eCQ�[��w��0�Jw�w*��.��if�7�� K��=R}��(_٤�Y�C0��-�H��xbmH��m�!5�"�e�`	Y��u\�� �|����<e���Ujc��9Cq��@~dW�K�,o�5xy�+TǛ�KW�׆z(nIg�x�YBR��J� /�Hi��RH{.
���v\��{v�����v���]X���
"5v���2n����2X��a7k�{���u�o�n�QO�^OJ�lS�	J�[ |��N��0ґ��b�
����>ıXIJT���5�o�q�8�@=���+���w��`�r���r���K&>/OR�#����p���,0o�@���3�֒��-"7���6G68�
��z�Nb�;�[q	�O`+���qI�����-P�#�W#�K{a�j��9|�w��Г�$���C����w����*%�@~�b�S��������c� �"����K�J�Qy'���yp	ڟ��D(�j�ȩz~7�k�/ ����UxRw�֋�-��+�Ɉ����5��.��2N�Q��B�/#�q�_���aq�����$�D�?��P�8�sC�>�R3������;�ۚ0���l�8�V;�8_����`8]i�ܥ�8��Uq�{L�`03g��{�xۓ!����<K���OS��, )���L4[��P��g�t���E��z��>!�4��e��s��
e�^��1�{�4� ����.��&�T�g-$��y-|O��՛�������Ѿ��[�9�ks�_��m������rz�a�����]Z��|��cmw�r7G���<��A��P��1��C�a��Sw�f�mb(<�}�B`N%Y�冑!Y�EK?s�L,HԉTS���ּ��[����27��ca
�ޑ��v�:<�M��V���٩��3�U+�-��q̲�9V��g�A�xq��S�lJ�E$x�W����-4�?=]����P۷Ȭ���wf��P�hZ��>]ģ`L������<u�g�7J��Wo�yM�F�3�D��22�'3C��55��Èo�%_�z>y�H���7�9��a�RI�W^TR��-h
��E�<{j=�5��B>y4;��ߨ�� ��f�#��N�@8\�R��3��p�w�d<`�02��PyK&�疲������fT9/��[z��9��%�Q��1�eV���y�l���X�ZTg��i��������O�=mT[�{WSBJ1�䨌����;`oC��^]�e\�kEb�l`iu�jͶ�JT^ ����Tم6�hX�Ҵ�pU�iC��L8!Aoʞ`w�ꘌI��V���f^����^�{(xksn����H����x����w�� }&!a�\ Ʃ��%��3w�C�$���I[�����_B�3�wa,47k�����F*��ɰ	WD����z}�ַճ	�����Pg���M���_+4,�B���]�7C��� �C2m�T�f��:ْ��-�n�+����#�O6éO�gk_�v=0#�A�Z�0�'�Ik�pd�:�
w�����l�;���]�/3����K���+�ߤ�ˌFa�����bﱙ(~�[wT$.p\o3�4r!��1�8�S������csچ�!s0���|�l�j�L]١�w�̃G�u+kt�hf$*���������5#�l$F���uG���0�?Mܘ��);�YZ����S�����E±�(���<	/�k"�~y����Ӱ���b�H%��9�w0�K�
daL���d\xM�!��f���?K��S�ۥ������| 'L�y�"���n�� �_i�j�nj���	��*-��1tҦ'�̟qn�,����N��VV@A�g؈9�xf���`��z���<-`v����g�䴅,�Tx@R���dQztb��c�ҥ�k��U���������(דW�����Z�G��
����I��-��u�,���,M¶sM�).l�,���M1�\��r�ֶ�8D���Vi9z@=��'*""�o�T�Դ�+�Np.�5j�SlS���#/�/I���(wq��[���OE�<xu�T������j
f�/�tag�ݎ����
�� ��<��g���YL+S������POu��g�nW�>�w0��w.���./C�*H�3��z4�n�(a�9yV'��X4΃�ѓ ~7�`MJ�}���Z� ��KeZ�����Q�VM��@��p!�c	����d��W!�*�q�zC�!��}/B������rWPS�2ϟ'�j�K�n����;S=ׯ��b��,�*�S�p4E]���T���<ѴBq�F��/�&`_x9�D�?J�R����ǹ�A�g�'NR]�� Sִ}îO|������.��?�r��;�d�iА�I5?	�d�[Q�BZk�kD³�l��?�_�Τ�VNR�d�{s�T�>��.������vh�jB3��j�ت��rM����,h�ʸ�������K��ٳ@��e02�Emp�OԈ:~��$N��ba0.���'{��B�$v��/ڎ�`��#J�/�d�vL��(�_/[�4���.���J4��F{�YBm�$�8"|�,�Vl..���UB.�-ݏ��X6z�`ĸ�q�{�R/�a�SHήDƗV|J]��{s:��}\
�$ ���ǤD�WK�ښ=�|�i�h>*j�/j>w6������M��q	q�Ŧ}{���i<���Bb�	�ǣy݃C����kl=9��~=��B���0�=���bìU�Ua�Pߐ�^���atAZ�i�E�%�л�uR�{^S~���X�� o!H���@�Z��M��[���%�[��X�Mhnm��l������7�9�����&�ڨsc�K��!�����6գ߂q)�.e��1g�	E�;�8��{�;����2Dj��$���s4щ y�����l_LOB�՝Ծ���u�5I棩[�_9H�H��� W7�|��5�^�s8i8S��F@���,�-�l��BPt��<͐l��-�ݢ�J� hϞH6�H.|�k( ]��u��̆'k��x1�}��p�;���¿��u��/��V����b}�ە�	��O����RD���nۅ3v���Y��
?�*ޣ��.(�y�,k'�h�6m����qy����z1�_����W�-/�4x9pXe��*��r6=k�ny��ٚ�����-�yo񯆶P��@�͗�?o�R�ݑ3f���k��E�
u���Ԕ��T���a��$�"��n|�����P������>[���i�a������������f&��iʯd8�Z�(x$$�nPC�5-�C��'!��P��
1,��}�q�z�sR�H�����	*� B�l2ǰ׆��)LWP���J�񉧗��0��۹��W|
�%�5�� �a~ ����3�K0��7��� �"��M=j	��E�*��+C�O�ʠc����/'�K~�Q�0�����.�5��|������y�U�����ɛ�{ז$`����!��&��Y١g���ΰ�h����E���X�r��c\��.|(��iMT��oA}7�~�99a�����{������:�:�06U��\Y��
�M91�ا�����B��*YkJ[�ۜؕ΄DW7��}o
j�Y�6H�л>���wLMl}��D2�{�C�����w(#l����m�_�**O�YU>�Վ��
Ru5��'�Y��58	\�2S]w�9K��&oG�Q"7�H���� n���`�9j�U£�-��&�^��7��Z(�Hm1G,F�G�ڠ�iw�_�~�܋��SB̳�^"��P�)�h��a&��}G�l��-)��� z�T0�b���=��ռ3km4,��o/��y���=�+�И����U�m��*���W��8���qB�>&Ɔh���
���E��ܰx��s,N[{X]��vO+�2C����~��^D�uE�^��������+���:�}�V�Lcw���]�����t�i>��\.������8'�,����� ��!�C?��������V���U��zl�<��Y���e�^�f�o7˱p�K���C���Ļ8��]���^y����J_��^�i��F
�⳶����Y���+������q�U��xeCfaIڼ�\��'n�ӈy�dU'�/X�I��Aɱ��M�vb����[rψ��î�Q����{c@��[(�DA7����L2�M�WiybO�Gmq��>f$��v��:6|t����k��v��ȷ��b��:�����-�����G'�y�Ta.�� �����WA���9���+�1� �;�#�"�R���oz��y{2}٧�^/r�����	$�,��e��'�7Yh�m����Xۘ5��}ic�>.n��ZP�PW��m������Ra�4q��_�R�Y%_{����DϷ�����4|����2&�bvO��4�ׇn�%V�8��c������N���$7�uۭ�%�lB�*g���*e�������0�*y�	�L���� a�REB �P�$� M�%1��/�PԾ�M~�.T��q�?�Z��|Կ }��LKB��l,�_�M������� |�J?0,�]��,�%h�t�6-�>�Ȳ=4a|����
u��/�ַ�7g����jPך��Y��+�,����XM�1u�e��łtؼ�)7�͊Sh�����I;��I̥�0�-k��=O1��Q��`j�K%@���0�Z�BL��]`�`̲�=��
��O���D�0�4����DC2��v�nKȮ�&?y��D�Ɍ��	 1 eC�Bݛ�ʻZ���r18�$�Nn� +�����8��d�:� ���T�����5wNo*;o\5���0�)vQ!���7���]���	���(����@M<����8<	��<>[~�
����W����"�1���ûx���(�	����a�+�R�_�HL���.V��0o��2Q��Y��E��9Sd�H]	�,�@��O����<�9G��ixK�b>΃D�o
�H��¼;-hs�7|%�V�,�ږ���:'��W��4����`' xx+-sj���L.hӞ�^kx��pcf#,��ܖ�����ћLSM���5�KE_���I�@yF��ye1�0�	���O�E@%� ��ِO�y����%��7�x�M��o�':�����L)���
����ĖR47�@ k��4��D�럘�cd��Y������$/�T�>��P�K���=��J���3yO^8��-��I	%�/�Z�\?@h��ƙN�[�$@�̕
��n*�-j�yj"���K5���!P^}I�#�0���qʽ4�/X����Y���j*W�0A�:G���_���5,$�<��r��W�>=q9��9�:�\y��Q֎������\�G�����33R��N�����[�IA����"&D��Щ�]&G,�VIlS������ƍ��d�!��(��Z f�Hȁ���Q�iW�Ђϛ�Y�I�i��HA^
���ֹ��	�&�O���ī����1�A���ff����r�*=��3a�"�o��u|�&e=���X��H�*�D�L�]6s��@���֮�e�bL~���{$��g��=���K��+�/?�CĂ�cQm����S+��Pwl��B�BJ"�������jI�o&��b�R\K߳��~q�9h��X��n�ȚI SW>�F���	|�r�hڂa�zp/DWd�j���[�.�/Z��U�����"��8�&xQa"ZD��l�����pǬ�� ���O�n@��:�Hw�n�7*�D��ѫ��&%�-�ɖSS��C���8��:b��2kd�y�	�mDktx8.�SZ�LqS�/�;��H�r^�]��&t���,	Q�e��U��((I�7�p�>>'�t-$�}�j�2B��|ų�#���d����ha�l��a�n��
�A~]C�Q� 8��o�}X�@��-�������x�n�(h��*�m�����{���0/&?�Qӯ�3�	B�vZn���aWGy�ӺP�j�Ì�
��\�]1���@Y�y�_:��E�oXU���|kuת8�T�Ap���z@��PPF,!o�!٣�a-b�*ao� ��k.W^&��:#?3`I�˕�5������ՠc��`����F�|�F�+��w?%ٰ\���ʾ��Y�U�oDP�~�=�y�����`�g�'�A��o�!�-��
=�4U�*�Jx���R���M�7�%�W������{��.tZ��8�!�C4�ƛy,*M�d�J֏� �-�D�h�I��{[�HU@�-�9��o.,<��Ϧ�Dj��$��Xn��R��cG,����_�^m� Q��.�Ԙ��9'��<��ʻS��^�����4���9Q�׿.M'u�rw� �z�$�V܊��N"&���qQ���}.�����)�<3��t����m*�]Y�]���eɵ�BE�3/�ˡժx�!����T"1��,�A=���.�(ΣK��8���D �=^-Џ���gU
��i?/]溗eE�C��f9�ǳb�j,�?e
H��XY�A�����s}�>M2EUdc-��b�n�-P+E$JD�P��9z�R2���L�~)AmU�mpp+���}h�e�ɻ,|x҅�=1N���*����N�嵱��y�����ԜBM③_ƅ:�,dpq(��� ����9�t��)���{ī��~��^��V�ũlQ�D�t��Y���E�Ubg[z���NDոo]g����2����P��@'��r`<��y��G�Ò}�r���d�>�㯻?�}�,����s�N����-}�6)����?�h�ד��`%l��K�j�8��aj����?� ��8�J-�ϰ�������7Shj����\�I�F�SRN��1Y�l�������Mmc�˦{G�0,�3$w��U��X��I�z���H�����HyB��1X.C\��py�������G��'+���4�2���$�������\�\���	sY�6 �pe8�%�V�T�H�e�hw�c�h�������lf�S�e����;�M�+�@���ǭ��=N$���V�נ!zN�B�����ס�:X��I�1�$�<������]�4�5ԛf[����u�bOc�w41��y��
��HK4�a׌lp��E��aI4�u�E����ii3�k`�/��
x�-�N{W*�`����W/t9tw3*�G�v��<��2Z�N1�W�E�)�M���A��u���6��H@��YK�S˶�!C����'$�$��[��F4nc��{���G���.H�'F n�GKǸ淏a�>G]O�`���)FM���;��tŬ��`� ����#u����p�?d[�1$0�f���3;7d�����>�z�y#���:as�V�`�g�5:��]�JX).�C�F"t+�R1v4z���
�t��)U}'ߚ�J5�?Ђvc������߳)4Z�ƀ{�}y��	,5�`.��'<o�`;�K�tߺ�*���Og��b���
��P��肕U\y5�#�4~Q���7�+�*�$S�L�����5�'x�ғm�&ϔ:���:��i6.��JD�Z�G.%��wj�.�Ŵ�i5&o�] X�mWH���3(����A�EwU�d��t�ڽ�I��(I�/s[/CSxH�@	�\��b�k�Q��2�lpN�S3L{g�Nk�4Y�J��Hy1+nM���fa��o�ם��b0p�(z9V���N��b����<S�%����3���|��׉�RpjȌɇǔq�Ez��넰�E�����+1���.�KLI���-�w��d��w0KD�yh�;J����eY�9i>�)���7�E��v���(�J�=j����2WP����z*��X�@�'��]�o^����1o�[��?���իƩi��dY�e��0pUtM��G�}11���:�� ������d��<�+�O��^�:1�5J��e�I1d��{F���[BĞi*?�0��=R
ʕ�ޝ��[�4�m>��B%7��G� ���:<��\�a`w�#$MȱtE��]������V�[Ȋ�!�OBy� �}ayU�y]�(���)��[�{f�^E��G6mV��[�zȗ�P�z�W�n�@+�I�n�Z���[�Fy��j{�?}C���:i�����G?��:�b�r�����wp��<���.�i����j�1��8��$�Ok=�KW^�����!  ����`�Կ.�Z�,���,�Ju�t�~';�(t��M��p*��>Z;A�5/.��e�e�2� ���h�	vS�E�I��� �mV�1ѺL�mޣ�.��?�s�"@ae$��p	:���<@EK7���K��v�L5F�N��1Sq0�D��\��2��[��?�e�r���y�z�0�d���as��j��
S��pT�T���
*��� I�vS��d4��
���u�8�oo�LQU��5�6=�j�u��]Fl�M@��S.��쵿��<�@Gfm���ǌ�bS������0T�/9�XA�Y�tVUJ�����r �
�ط&�m�f��ǵ�)���;dC[�' ���?���j�pJ��FkP�}.��8��ǟ(2�^ GN�����q]�N奸*C�o/QHY�!�0�;(�'īf��*t^F�%.U��Nv���,�(���&jGO�LGR	Q�?���ҙ=z�s6n�O�/a�fK=��K��OyWE7~U^g�+��ED
~��\� ���K Y�3׆�_��FD7P��U:4bN�`�z?�U8������1�+� �����3��rg�at�FjI�bx�j��R���C����wGa������S�!vfgs��@�q�V�N��p�4A�8� k�!䬙#���(�Iw��gRǓkT(�S�bhEwpN1�O�8Uh�V���}�/smA�����x1Q�Yy�k~�A'|z��n,��5C��}^M���	󣾍�9)'@�\dcI_�-������q������L�\���e�&Ic��Y,�����ʍ����w�E�9��������3�1`�WY/���¿�� epQ�+^�.y3v�F��JT�8 y��!y���[\`tjM�S2I'|��EDؽHޝ�	<�?�VM~�,�-�*c���K��`�A$��*���a+��rD�*��!$gb4�L��*�/��]+C�r0o[}rڜ��)�j�{H
"^�p�'е�sJ��-�<`��Sn��f��n��.��2Vמ��o3C�mV"߄�s^ۢzj����Ѻ�%V:tBl�u�|1]��B���O�f�m�_���׼i���YOu�m$(���7���S���yC�H�oR}NnK��I\�ˇ
�!|���*�*ZMD�� `1��\:[��
��$z����[�u��exa�,a9A{�:y��4�`_�D�awR~�}�u��&�~q�c�a��f�4�=b�S*l�����r�!$[����&���������'�l��9���t�Ӟ��^�=��7;B���wo��w:��b�[�Z��b5F�� 9@�b|y�_Ƹ~JL���H*��N��[b�w^��L���G��bx��T���{ ��.��y�K�I&+��Y�ڡE~DR�]�!��4�2~�'�]y[�_Kf��W�L��V�q��;�[d8�lݨw�n�:������zM�]qzo����L��o��k�tT:�<�����w#tV�O;�m��yT~]\�P�Ԇ+��K�^�wH'�u2뱿���/
\���W�i�����|��W�7@��4��b�mfu_�_Z8��K#M�]����/ݶa��H�_Q�O]QOdv�H<J��WA��ۗ_YhX�I�u���(��L��wC�,�-Ѡ �U����ԙ�x�b�c��Aj3Q������@a��0�l�E~����!����=��e������@���Pp�!=��rk&ؠ휵dg��x��U���e��M���x-i��ӝx��'�2�y�8:n�c��ԅ�#%�;q��{�d��V����GA�>���uҝ��W&����̩됟<�����9�D�T�J�e��f�G��_
H;���}h4c=4|�l�U�j��]�AX_���78���*�x�Vj�[!�����@�k���4u�]H*'S�����ʚ ?6�ZH�?b�msl$�I�2�.`��F/���j�V�|yzya�r/�F��� w��s+���w�ͅ��=qm�b�#�rxYMQ���h�x&�D����T�n����I�PZ��H����GK��Px�}Y����=�Â��0�*΢Vdw$���LNx~��x;�#%��H���X���|���Qa��Ȓ��r�s�aPv�'"�?�7��8<��l�l�Kv��^�ʃl�_�l�V`�MTr^�����q����C^ꢂ��E�:�Q��<���0���
��3��H�9>���4���@����4/����������ǯ:2ŀ!@�	K���9�Y��* Bv�3�+�>��E6�.My�Ǆ����8��{.�o�w$��Y�S���d��\P����b^�EwR�I���-:0uU���m�tT�ywr�}���^R{��G�Aw�aj6dipye ���(�_>VC���4���6�%"���^��+3m�:�%A��S{�ܙpyN��W��7ư:��u�8�J��LT�.
Q����;���^��Z�V�l�E*{��$<�Q-����k�k��*=%f�+R/%0A\�d�6I��R����dP�V����R�x�y�3��'�,�կ��8���Ol��>0�9�>D�º�"�t��栿>}���L���o�7* <�%D����lS��j×\<Md�{�,���2|d����㉷&��P�3{F$�4�j��2(DHA��o:f2O,C��+�g��C������)��?`jx��s�C-yt�؎��׹ ʙK��F�z �$�����d�)��z��>jI��9G1k��r��U>�t�Jz��>zR�*������@��Ն8g�
I����FY[�����f���ݶE�Fb:%��y�Ֆ�j?�?L��+h�gI�kc��䣢�T֫�q]�����<�~]$Z�o�^?��Q:݊�f���в5�/����thko�P(P�.�s4���ү�H5E���,����F�ԎP������7KRuF㵛�۰X#3�K�6A��Ht���+��v9��1�~��4����TFO�nT�Li��JV��Z!�>8�� ��;����M�x�����jgޣ�Cc�d��L4��}�툴7Į�E���̓+
��u�3K!��W�7���x6#��`��"Hm�MN�1�[���y%��-�$�M�-Ӻkn�No
p�[c��j�-AE�r{����^(;P@7D�^�I8	���R(�Bh�5>��N��/�6���t�~��tG X�"���z)�AX�ͭ�]�W����YM�S+}K�b��Z6scZ��N��X�`N�$m��h"�Ȍ��D�A��'x�歭M^P�z�LS�V��C���kQ��UR3�P�%�D����|8AS���;�/�0RE�W4j,^m�R��:�ũ��}^$��H�:�֋?�%�_C�v�ֻl4�FeR{n^4��kL�£|�*VK���R�b@$ "� e�������VzƔ6����U�|��?�c�%�*�e~����+8"��[	� ��`e�dkE�!���+''�^.��#{; 	��ݥ�[枆,����5!���4',O�^��˪�s�ϧԖ�0�N�lJ}��B�'��U�XI6�Zj�d닚�1W�����(#e�C���v;:�'L���\�t�
[}4��,����%ܭY��T��k{(yk���-��c�oU��R]O����?:273擕�O�n�l���n�
��A��_���o~#j<�R*7&慠�0���][h�l��[��ƄBrp�ӻ�C$�[$d�v�	!�j$gP{sש�	�5н������e����bhx���oQj�����PkL�7
N&]�쏐�?���mcU�zS\�3�襊�".�KI3k�!��I�]b@`ݛk��O� ��WGO�0Rq�k�r��e�����6L��zѱ�S��pK
��c$^�/O�Ґ�8^������>����م�;���8���asɦ�h��C��
n�f��MF"Y]���'�ܽ��Dw'���I��^Bo�������}b�� ����,��f�_�FzG;�x
�z�O\���n���an�$Jw)�+�'�3S)�?���,V�t�����鲖���08u���R+'[��Cӑ(���E׻����SqD�%U�T�����QoM�E)U�tQٕ��YM�[K-�����
��ds}Ѝ��[�g|S��A���E�%����s��=����7!�|��Mv.�:��xx�����-3��%��odV�S����K����gg������L����|s�2T���bw�3�6>Tl�a��k�1p.f���sޅ�Q�|�P`*�}F���Edq����h{�I8�R�xmJ�� ����EN�|����Ǐ��u­�o������(0��T�>c���6�\��6�L(���U�\�A�E�����eYT��U�N[��+��p��m.�E�K3��47Q+�o9�X�*��l.�����1 �=x=�'�%s�F�^���1E��:sR����}f1�N&ϲ�mc�k��\���g�	������B��ܻ���A�a_�4U�����C?��A-T��n*���@h�Ed������h2����ܶƏ��veME;���m�ܸ1��0�R�i�hעY��>����E7`!R
#����X'��\�u,&�F[��v�u��1<X��㗲�~'�o��,������h������Tk@N�#��N���}�nU���]Vj�y�Z��8��S��@��,��Ǩ�Q%9���U^�x�j��^��D<�tA���ٍB�F���M{�g|�e.5^J���,�� �>�Yߢ�t�H>��������b�����9��Gѻֹ���RF��,	?i���[;���%�bKrUjjs�̃�5<�?��}	g� ß��l<�[����fP.f���P�N�.�=!�YU��o�L���?J3�x�*X�{�o����?K��gTE��Re��ɝ�m����(Z^��4��r��+;7ڜ<�3��]Pҧ%�)i��z47t^���\���k�>,�d��%�K��.g����lh���A�� �M�2�OK�td��e��#���A�.༅��a�+�Ӵ�S��2�w0΁E�.&)�2f��B�/��w��c�LW�k�q�D|m��'C���k#r�P��.��r�BQ7&7<�c}�YAV�3����W F;���M,������MV-i9��#1�6!�K�Ȑ쳫LZ�>aV���f�%~�T,��h�����0���K�?���D�K�v, 0l��\�JKY�Љrػ��澗OQ�c��Y��/�6�m� ������Z�^����j���k����Mu�j.�T���	;��9$\�LnU�˯ƽ�u�]"�NK��ѝ�lS�[��6���49�+0�:٢��Ňm ��e���s�+���گ6�jx=�*� u��a�]��CX}^d!�!��/�9���W����v�ǯ1d}�'Xn�������=����:��<R�%'ވ�8�*��wj9�1κ�{���j?�#UZ O�r^E�D@�l��;�x��P3S��)�I����M��m�xes��}�Ĕ���[}OB�������M�3�43��@IAJW�F�<�]��}1��@�r�J��k����������ſ]�y�CE�H�)���H�yd ��+:T�<���'j�	߫�7��>��r��g����\]Q��̗�����^U��ܽ9ј��:�V�H���+뽗��T���( 1�����`�	#�2�
��*%�I�(h鴐��B��]�iʂx}�C�:��Ҕ���7G?��U��k<�3��E�)K���n1:��7C��>�-�6
�ޣ_�L!���׀���>����-Zq�F���t�x��AAs�,��	�z9Y-�2����b��3+%#�"w���������e��� Nei(R�*_��_2�4��`<���Xډ�~�S�s���=J���
۰{��WI�u�s�(�������|�x�R�S��]�Us� ,@i�}�v�@��[Ki�X��B@fN�fgC]�2P՛��\5�uUо���� V|%RU�>��,���F�p�x0E�j۸�����!�Cg��hꕢ��	��X�����Y1��2`uh��2�X����������@!�P�*�^�u��Z���+�O͋�<�C��̯e�hD؅ެ��������Kf�2��Bs�R}�������J�8Ӛ�F�9:�"��y�Àb�Yq��֐"����2b�@�-��0nχ�]��(=� �u�3��~&x3�S���%-���o��tt�R���q�%�3=ZPJR*�85#@�P��vO�BJ�!���G�n�ӭ��,��,V�����.�7��-'�\s}�w���9K���o���˦hV;���	ƍs�ۺ�e�2l}%E��_I��5�w��ۗKSa�!���Կ���Z��a�{	�_yN:6Gw��
�S�`J�JyVe��<�1����Q��$�'��ۮs x{W�����è�����iL8h^��iy@����32���]�&GEu��g'�܁�q!�9a��������AXL'�����.�K���/n�	sW���z���[��r4A���)Q�����K���m�QaO[���;���^� �kj��H�)+d��$�j\�|7�2'���`��s��>�An�d�`;	{�9�0|��(���O���:sO)�u:̘�ڛn'��� x$$=1�61l���)v�2���P/I\Im�O~�i��Φ��m��Gb�aפ�;���V֏m��?#��?�i��,G���P�C]i߆�2���Zzf���3��Ԕ�u'�b��e������2Y�A�	���ߟ�,M��5|_���)�owS�U����H}���3�q/�?Vp2�`���wT^�'�$p�I��c���������v~�f��B����ͺ�E\����N��ۘq#'u2��\X�N�Q�+�/�(4T�=|�>�q,���TS�yd��O�w7t��dCI�Y��b�P,�d=4m��3�!E�K�厤��w��6�C��F�a�%�Y3�V��RV�K�ǁ�cYF9��K	��I���kM��P�E-p�P���<��_���4ڙC��Ý��CzF����8�Pw���b��+��,/B�����C�����E-�9��{�ۣ���q����GhgF���k�^�|��ц^ȣ$_D6�DJ��َ&���
ނ�+ң��7׳��'�7w�\j
���=�}�+�2�ʜ|SX�-�k</Ro�5�)���tI�4*�+\cq�ۼ�c!��s�:T��U}�?�|�X/[cU��i;��Dl>��ჶ���	r|�}P�co��H :�L�V��.� �����2�֤��6bz���%�~Y���*���C�;�JĐ��8�R�a~�7��NTk�$?.�*�
�5���h�;ݦ��M��%�Su��8\M��������Ea��"ذ�����@7�̒6@��M�B7���#��t�N+�)��EﲡB�Gg(C����A;�`�f�S�H���;pD�$�:��K��*�@Θ4���	~��D-R*��_�wʶgzm�v�d�s���cU昀��I?�S=������g��k�P�J>%t��~󂥆Iq����xf7�/��� K5�P�]�&�<��_�<kHИ[�@����ל��l�v����=n�s�ýރt�����=���# ����l9�ew�T}z���{�7�;�Yo5��_��?aNz�Jh�h`��B!r�bp�f��.�7gl��B]L�o�G,�X<fJ�Z�~h������I��m)<����T�T�Ç�Xob�-��#^��sK���\u�9i�e2��<��,�#ͳ\�͏Z<���_��O��"㻕��aP���s-h��^��g�}�"�:|��aTo%�e��M�
;�<5�~���jT�v_у�_9��e�����l�\�c���Ā�_�F�;���2&�+��j��L,���m/ߎ4Ȑd�hڗ�K���6 ?���W_z��l�'iԔq��R�������9��*����S��?�D���1���G���֌��D����2��H׮�&�JAH�"���E#SN�έ��V�b����-��U6��$�Hg|���I�]����k�@�~s��Z֮��N��U�ڿ����z�ܡ���a/'���^>]���)�6�����>�]��J�G����7�$L�z|ur�%oNw;�d�4�d�$�iF�7���+���."�
D����lqlP�lSf��r\þΒT�hJҎǮ�V*��j�E ���Y�E��4�I8S��'�V�^)�ߘ�V0�`��oA��Ü`3��~�؟���=
Z: l��ep�	��U�2�A�ءK�)0���;�*Q�����"`���XK�:�!�{R��?��'��|��k�ٽ-�m�!?a���%������7�)xM#W+�_�]���6��^��Y��Y�/�턩�E�w=V����@p%���C���6�da�-��<cΔ��E��([� ��pt��||�צ~����K&2������d;��� N6]��j�&�B">F��+����C��Ѕ�WK��1�'#F��R��ݭم�8���4�6?���������p*�r�6
����ʮ �
O!��Y���~L�|��H	d2�e_�Բ��e���Y���b�?�U0�eW��9+�x�x\(���/���T6��"?�j��~���f|���E������".)��]\U�`@��uU�.>���q���n0��hh�,�d=bT��~��2uφ⋊_�T����kfp3��J=b�e9��WQ��-�����:�g��9`�^����yc���U_H8�����jU���<�����p)�̠���A�u��;��&J��橝�>Xˏ9��� �@~��Q�?����R����Gi���z݃�~�^ʉ�va3j}ٸo�w���+hя]�s(��2y�A;��$U
��$�t]B�mJ2\��/o٩�}��ӓ-��3Z�!1����&�d��B�X�K(p�/���/��N����n;p�m�$}���K4�@���ŚkA��h�0gY��>���zs���A-D�"��4Q1�M����ǔ��k3��Fc��'�!G�LO~L թ�\Ĝ�����cX�)�pHc� �t�"?6|x�B����|�v='�0�1�6M�ecm�/��T�6�]նB#���F8���sy;[���<�ên�i�s<拉�`\�?ǣb����$4�$	��ryoS��}��Wa^��Ғ>G
��ؚ%�b2t{qR�o�P�
[��dGxSj���T�5f<1&y�޿��pN�[
�Cn��t�T��*���߾E�A�n�{[˿>���p�g�����Nj�dt0�/o!{߷",tA7�G�]oѓ����xE�6.�]�zE�ia��rc{�#k�H�C)�9�ܜ�7�h�]8��迾�FA&��i�1:i�D�-�
j��j��4�����X����K #d"�yZ؁���G5?���Qp��Hp���4�84��%�EJ�� �w; ����������J�kI:��#!"�g{�4��s�3N�F�#���|\kBcǶ'���s.Ԕ�����	��<3�1{:А��
WP1�zya̦�	����f�2�R��;+�L�4S���A��I���"s4�7�&�]��^���v�#�1�F�*J��!��0B
7�7�����К�k�Sct��d��D�2���$/������1~�5��ίϱ�`�AN2bF�r���O�G��c��s)�����;r<:ʪ�(	"|��vXyR`Ru�=��֥Uк�#�)��iZP�o�':>

�n&67��ɕOQl�|.��&΃�L�v�!o��3`�ز�Jj�d�e%�H�z\�Vj̱f8#��)���^���hL�����1�ƈa�(4�Q(��Yq��N�>�9��{Bϑ l�)6��n* n�?���E@�|�&���{����~���/9Fn�Ez�I<��V�#�^@��q�+}�S���`sh �H�������iO!D�!�"�K�J3)=ŵ_M�A�Tk�C<�״�����ѝ��?���%�8���6�������w��-Isd��t�ssj~��u%Po����n��چ� �K\�h�����Bby�����#)�IRr�%�z3s����G�����/NN��3�p��_���]XRܼ/�Ɣ�Q�Q�_#b�6�s��d��A;� �۫��s���������q�����g$@�
�	}��kYl���S�w�-�52��XÚ6'�Q]_0�:F��r�Ф[E��g� P����/������e�Ι���;ߏ(Y����Y��x�~��b��p��WT�E^���)7����0�Ƿ4�B��_\�PK�7�}�1޳bo>
P��6�o�=�x����q�AL$�b:i=ҫ<�x�ޤ���x �s`��܃�+3�^n-�^��Sl{���h�W �����>���y�n )�ܐ�5����qJ�|-��
�3_ak����MW�Y��S�|�W��b�^������븯ƛ�~')�0?�vF�N�X���Nҋ��㛡��ާ��PѼ#oH��,��!|�XN�,�Z�=����ş�C��s�M�`�Q�ͻ3�sx����N��{9�/��6W�ql)���ߛiB�:+��r��x?d��^]dz֣��>vI�ܽ�jU��<�٤{�[�^L8��u�_m+�+�򶨠"�o�{���}�*����DAP1���7�pl�~�Բ����T[x�´�}�8;�{>��AV�������K\O�^��Zz���óт�+~}R�����\������C>Vz�4�����E���Y�9�4��k�d��E�2��`H���ǂ���q6�P�vR�SV*�f:��&gHڋ/
���{䄎5�h�GGc%�]Tp2�_����8�[o�00�}OF"FP��Y��Y���"-Z�nY��_Ze��V�҉
w<�j�QױH΂Ų���6�����S;�MVN��9pT[���;�F5̓������� �4�ٗ�%+��XJ�H0�V�rmZ��J\��Q�Z���'Q�[�TX)8ț��Z�X��4��=�G'���C��h������5��Z��1AY�D�`���cn#������&\1o�	�t�ٗsP�܋A��5M��H�c�^]��a�� �:U y�h_��� ���,���Q��6�0�WÑ�Q�~�.��a�z�p��U�K�鰇~������>G=��Q"���-s�v��M��aX����e��܄���A�j&K�g�~-\�<X}z&��F�|opDô�����,;�7E�[01 ?���W�[~5�N����Q�k��c"-U2D��s�[��k� �Z4��uvb/9y��4��J{B|&~���<k��.^W��B�J�	[^�R��ɤ�V���0�vg ~��N��b��LF)����'Gı�;��(G�7N�ax�`́&�j��.����j�T�|�(�u�7�d[tZ}p����-X����� o��Ō�����f�~�!�$ALSV;�:�����f#�%t���G��Դv�8(�Ɍ���N���ی�(dB�S�e+\�g�+M�ns�	�B�^]�*���E�IJK�~%89H���3|��{/ݭL	6E�,/��?��/��?0]��(���չa�-���ȗ���� _� �����0�s���@���P��� T&
k��1�UΩ@&���:���� &������MfZ��[�	JG�&��W>D��v���,�j�V������A�f���,��H�g��*��8���5��m���ˆ����Π������p�В2Ȥq��ӌ�P
tgCW�����_���/��K�)����ިd�\H@i^��R����%��i�G��ZA�<	���4یI��u9*��A2���n�v�_ʼ���oy��n���#s~
F�/��꼕��Ri�E�liM������`�+�X��F���GN�Y��Yj�vL�j%������1J� 6Qa�`)��5
.�7� B�@5
mZ�F�(�~p�j		SE��g��K.-��0�dB��6������L�c�X�ϔ�'�2�9�	��#��oM�� i�,��\!�Ì���F��n��ك����?͙k����?8��TB�SǋmM����o��k!��Z
�x֊k�0*!�?�-@���PJ��F"��]13�({�Ӎ(oc)��aJfK�pY��L�2<���� �2�{�ݗ(��͂N�0S���=���c)���mRb��0Z|۩��Qz!�-�:K�m�ҝ���tc�u����l �!#�-b%���̺cPkχ�0^l��$ƾ���i^�h��S;L���)���δR�caTi��[�I��.�i�OF�����@\��s��#3O��pVZ:�<�����1TN�#��^��v�SP	Lw�S��b�G�Yp�5�1m� ߽飖��&6tư��苸|�c���Z�K7a:��>P*�Z)^�m�@O������i��K������ۖ�h�Ih�'��c$ܜ��A�O��G�=�l:�s� ���r�Ș�:^׭��p�d�����Vjo�}O�ֶ�����-��ŭX\�yo��a�3�f�n� �d���câ�P{e�Z�(D8��{�Y�y���s����a��lP�m'��f�"�J�T�mZ�ѣ��z�q Xw�ٺ�,�pJ�&��אm�P���ΦҽDj)Q���i��I���|LN����\����b�bb'��2M�@�׊�&�>��9�Y*s'��:���^,qf�VtՖ �D��A'� �|S�P��Ê����>|�"�&9Op.���N|��E�Q;��v�������TU�>�<�_NQ�a��]B R�*�W`�3_�l2�4bDY��ҜJ���4�<�'�����`���9Q�=��7��Tf��O���N��Ό�̯qa��l�����9d��ۄ����dA w�-p�R����6�J�xx4a2�3J�r���E�>��.�R!�:ZT2���j?ʑ~�����#�-~���H ���Cl���.8҉g㕇D�?����d��&���B�(ޖ�0�nE�C���Fen��~��7%,JQ��e<�謓�haI'�P$G3�^
z}�U��z��B��/��s5C�g��tu��M*����=ܻ��|��V�9�D9���t!�98��^��Ӹ:�q��R�;�+TP�����ڋG!��Tw���q!����� NSˌv��|"�;.;��j.�0�'c�m�F
939���~!ǐg+�*�&:���6&�m��Eü���?�&��ų��-��H�2o����o��~Jlҙ�o��@�#:=��*��Qiư��	C�[�fL]L��=���p%����+�T�����t"�
��|���I/���&\�Z�����ÍAb�`ʅ����:}��m>U����ʘ^_4$�Z�徹,�Q]@�o ����SVk&�����~��yQ��n�liQL�T�Hi�$G֗� \��&ӝf�m5 �Tqf-e�o����-l�^��D}`]�O�jT9x��@Ӯv��Fʌp�~|��?M��<LDȲ��Y͍�D�!�)8M��D1N;�Mf��n''ҚcuY�~��:�B^֚�c틴M������O
9�c��o���,�,�*����O�LvTj�S�tu3��EA]T���fQZ���M6@���A�OEU���o	Ƅ��B����d�$�8�y&���[��ݮ~G#7���,�MԌ4��m���EJ��d"._rg�}��GR���b^�F�^���d�x5A�4�$���o��y� @/�
�\�Q����WH������*���y��Us��='v9�0���M[me
emHi�����u@�M>}�m 
z�T}��
%�۶�[��vB��ܗ��|��_��$npЗ�ɉ:+�9.uյ^ܟ��o2mYQ�!�������awq,�j��r���At׬Y��ҷ���G��Rْfb���z�hR�F����!쑵�C
g��mm��8��j����wݱ��"N�X�Y������/��ӐP�j!Z�<��$�ƨJ�4�E����"W��(z&��8$.�w!�և"��p�WƁ�E�:�p���T/@��s�}����P���?��? �3]v��f���`5���قw"���{Pw�;H%�Ѱ`�H��w��M���YN����y�V��Қ�8�P.�$S����QG2q��!�-�(|���ҿ$.�!�eƠ��nC��AKL��:�/���W��!�s��R�����B��6�`�8&�s��U���!�r����b�8*"���-���[�9����b�>OrN�>��\���{t^��W��_1���J����M���s+�*G�SNe��b�/#~+s:\I����=�?����&\�P\��1��	+����zi�\���]:�f:�(�5U��p+ѯ8gx�~��H�p,��@r���ζo����-��a��_�������J��p��1>��Ǳ��x*6�f?��]�EQ�l�', �E�D�ǌ��j��_��ֱ�ήeϜ�O1��/�]L	�#�S9�~�<����`�ܴko��b��_ǆu�a�'=O�%� ;�W���z�,����)t6�g�p� ����I8Og�󨗉�M��I����ͪ��@ơ�O��5�m�t���9���11�:I����Z.=�n�+���#�n�by.�(�t���}�>l߀MA�kB0�y���t�ꉛ���)�޲z5��D�^�0�܂��F�*��-�r�b�%ek�9�h�-���_8��~Z���MfФVC��F)51�7$�K	�zyb�@,c�n	_,V���&Z�߳LJ��@�${���t�W"�%&#-O�|�Ie~��݅N/�o��eIY�U�y�~��tޥ��j}��{��d�9hLJ�mJ�sZgO�^[s�-r_��𮱤���?U������f��bjR��l�0�����='<��f�U�_�q�c�/X%�$]�A��M�O�I���#����P^�m�8�Vu Wܷ3z#7V�Ɏr^�D��w�g;�
Qr빨��3`���{.�T�E麁xwed��1��ٯ��&��U% �?"�����4��m^��{�ە+}F�0,$YL���H͒��O��*�c��d��D�G[r:��>6;�A�5����4Y:�.y�
s�pJ�u��SO��a���a�o���)U�q�3d6(Z����1'��S��;���∑��[� J����]c��w}��R��:������P���o��|2�`R��{n�w�2���O��lD`���V��rؕ�)9)�fÐ2�H��'�݀!Y���}�r�u��5�pl9Ͼ��\6�k%;t"��4�5�Bk5*|a�n'&��QToҫ��a�6I	��m$̦����?M���S$��{C]u��l�
v+hs���u����n��お|O���a�"�@?�U֐kQG���"�D+��%�JF�y[�z�;�Ļ{J_�Zl��գRӹ3p��,�rvM�
Q1Z9�̔�Z���_�gEY*rV^�԰k&{��v]��H�0G6�V����K�E����D6��Ы�J�d�;8�Q��3�Xޖ)}�ς!��䟔�
�xfE�t��o�P�RX�
W'�1��P��e2���.��/P�Zv��:B%�,SK|�ٚ^l[��Ưbs�+D;�s#�bR�Ĉ7�S��
8<��
,�����0���_~>��h
�����JŤE�Q�lI�I�+��96}�-A�D$��jL��>!% إİ��l\Q��"b�A�d~b�z���@��%Z,%��7�DZ�'c�ے��7�������uH��V�5�"'\��T	�&��ot���?��H4<�n��ڮ���Ύ��eE�Iîea/��S}�{�A;nM��Xu�tMG�����h87`{]hh��=�Ӏ�s��2�t;HJR���#�:��J>��o����պ��b�_E'KW6�	$:�[8�����!�p����h�{nlb­���S&��ȪX��P���a� B�<�VZ!/E�V��V�E�"��?��ޒl����ʇH��#�."y���G�Q�xa�@b!��k��5��%U-�4��lB&���WD ���]o�ەX[���UT䨁[߅��Ē���%dQ����,7$NV����3�uj=mpN�p�|Jk	�T�U�����ۈ�x%���!`(��<�0'�|�(|r��e�����s����Q�V-�MI(��j����kwm�[�h��d��L�!���Y��	}�a�]�QOس�]��A��m��	�X��E�
l�[�G�������"��3�s'����<ٹ��lG7�wV�H����cS���uB��m��0�z��YZy#%pL��٣�<_S��-�J���,s�0�;����-�k��u��˷J�*晽a��A��� ��02��aP��\�>�� �A�_տ�����6<X�Gw~Q��^��<:��R�k�A����*�7�6��`<��S+@8�g���(�	 �C��2=��awbyo�Ã�j��)�[��)Ҍ��u��v>e�ʽ[�.�+ԋ��BVȧ��m�S(p�|�)���D]�W:�:tg�&a/���xErt����'@��{Ԋ�ZA7R0���Q��팍*���o
v�33_��(��[��/���V�SߜgTމ��gۤ�Yʲ�D?A��vI��-��sܾ�$���e@7���2IM86�ᅥ�V�y"rC�hG�2�^]�݇�NdE/Gh�M�o	F��.�1��S�������Sm���"s���"O�m,E�� |�=��v�.�Ҋ�9�^�R����Ґ ��A�x�C��@$�a/�I$Rֆ|T��W��K���G�kM��z
�qj��q�����h|��P��I�B҃z�il����3xAi���B`ޓA�n������,)�q]'O������͘�Y�#N��/����ޜ�c��u����NA �>�0%�^ĉ^I�n�7p�tf��5�5$�/�)��ƥ� 4�D�9��qA;��R>G�5�	��Q�i�:ב���dn��X�b@�9�֑q,���J�L�Cz�@1����T�$ӅB&�շ���Lʳ�N:�և�L>�� a2�1l�4�}����9&F�,f�% �5������=QDB޴z�i=s4���o�h��=])��=�@��@��:Ȯq 5���6_e��AN�#���|Lp9$�m}M߶��5`��[)�k�"��t��I �.���%ȗ���0��v����K�N4����|ѿ|Z{��N�$#Cn�w�=���?�G��*���:':p��-]W������,�ד�$�:��}��p>O��\��ھ7�!Sa)��.t33X?U�������M�R��8�7g�+X���lr�L9��w�Wa���2Zˀ,t�(� 7L}#�\l)�ᅊW��ʧ�:D�:Q5-F�B5���/&K�V�ct�lh�_M8�������m��*��]Se���[�ap!��G���*��|lV��a̎�������M��X�t��x8�F���g��aP��M�ө�f���p;$u��D$LO��p4�e9��Xڛw<PDR#����z�{jͷIq��_e�p"��ӂ=�_�#�eÌ�Y�~����{����j5���5nܩs-��'e�$@;6m&wC�V���ٱ�7v	����P���G�zR߫ h�ή�Lé�2���h ���uu���M?V �t���6gV� �������d�5b��Ucu��K"<��&������Y��	[��@X�	���),C�O^B	���/Q�>��B(�m\Ah$L#�EX:>�5����O�~�X̾�i���
�7�Q��B��7��(U�B������A��v]o@��
��b/E¿�)W��{���h�y���]�&iM��'�����D]_U�e���+$=BR��	㰾ǨD�1�sZzނ�$~�Ӯ�l�M$Eg�ww����Fv�H�$�L�_*rCǬ��/�Ժ�DS;(Ks���h��H�N}]���6��Xh��|��ZR]<���5IY�)���Y{��oUS��(�؇�,$ˡ���}����m���+P��u{��k�w�����0��/�xy����S�Yr?٦=�V�^/�����W���&s\ ��8�b���'�+��8�\ ���G�0lo�y����#��)'O ���:�W�i/���
r��I�W����E�E����G�E�b˄�Mr��\mE2�T������y�E5��|��B��M��Z���7��"��T[$K�Dh��%���Sb�Y���5�74jy���K߈�P�ڜ#�� <2�k�¿1�ZM�S� �!�7����Wi�6&t *���<Ha8�l� R��Z��}�mF���Q�f؛JF�zqZY�6���?H���u��=𔍷*Kѕ��Y�p�E�^df۟�pK��G�"^b��{�$mx��E�ͧcV&Pa}������^V�ׯ����V�G�׍l��)���eC{�P�1�0�i� 2�-�tv��͞��[(/�^S����'�1+ʾH"Z4%|���Ky����11zu)]K�_�}�C���9 �'�š�O\_�"�(ɒV��O��ZX�u�L�<�A�3F��dk:i�ö����KmP�?҉|�o��Y������+�2���.)J|���.�U�����dQ�٩Q�5�A|��ծ%_��C����U����ȡ��њ-�[0�d�H��,}��1B�c���s)J�&Q����Y�*�d�}���5���IU�u�ZE���2��4�w�q��\^|f���Ĭ�˂��r&�[�����R^�f���~WR��tL�����D"�|��6� ����ؐ6�C�$"dĢ�·1xܖ�R)A$`@�％5=rQ����7���]9t8l�_�*��:�>9㎧@jR�К�^�音%Y�ޝw���c�9��x�6Gb�-3��%>�<7�#�����=�-@������ ��W���
���| <͊�Ӻ�Bx�r��x��101Ig8%���I��L�g5
�
�P�*�C�#�n]�=��~���|J8�w�q�Yz�;=:�m
�l__w}�i���BL�S��:H�b���YV=����
&�<T_�c˂�f覬��������d>-���}�l�ctL�m��-����1�Θ=�"�ʿEoX%ewo��DA�M��麳F	[I��Q���]������jT�#Y��T���d���AX��A���~��R��4��<5A�d��Cͯ�:�F���W�[.잔�\�ba������yCB�b��ə�js��-1I3[�z��s�Y�����>?/�� 
� ۥi�U�q�1�0�&$�T�K���qӟL�ÅEH����x �����D�+&Y��'�X'v�.)������
�մ���o5�ҒPb�1�EvT"�?yۨ����
:�����E\����'��ǄEK��)�N݄���'+�er�y��S��@���w��	�	������Ւ��QK�߾I~�����%n��^u��f�m���A� ���A-��S1��ܢ��<e�c�g���!�\�<�����х��x�P�Q��Zal�-��@�N��dg�[���!�� ���Y�M���i.��`VPQ�U�e�U��K���[�C�������� ֐�@W�T0|<�7v�`��3R�IB�f�f��+�`%]�lᴓf(p�.�\m3�&їi�'�ǡ�.�V?c��DtȪ�T��F(��s������m5�s�����i�i>(N�8�0��C)����u
�W������n�h��Ox�����PS2z�LL\I���Sd�C����h����B�=>"6����!�ȕ�}ff�v�Iֲͳ�!�ɧݼe/,��f�e+_#����^�ڹ��6�� �<)�Ph����$��@À�`�z��}�]F������'y	�V�q�˵9!�����5�ղ�5�eq�\�`Any��@l�^O>$�4���6 ]�,!�,��N���x���.���fB6�B���ӥ����m����]C�������}0������
D�@�TA_����*ѳ@$��O��G�5���OS��ȍ����W��C���;� ��!���m�K�A:�R��C���ҪC���e��������ߤV!����X�p��cغ�p�;nL t2�N�����!�+��f��w��/��<�x�����y����3�F�e�-���+����'K�i�+1REO�k�~�[e��i%a� ����ɢPlwr��56(uP)�F[uSt�1�F��z��S��:��	��|�b�*�U�|�hщ?������	������}cv}�����~����ݛ�1��Q�?k��,����2�"=nJ.���3��
{�L�(ZE�_U���P^�Z��.�:�t�5o�c�	����[�q��y�Op �U�0�У��*{ki�uH�����Ĉ�$�&�=59�a�>�}�Y��u���\��2yo�G�\0�&���@ײ�.�/��[|:WՂ�.|�s�&�1OܽNc%���ǰ��+���\h-��8�Q�O"�ݿ��v͋;��6Q<��hm�?��
�/T��a#�|�#]k�k�OXa����д)��klf�H������%�<�y�rmHa�3ʗe<eA�_�m� �a�+J���=k5�F�wg��Xe:�P�{�S	���	)t:�� �C0���	1%&)���d��I��C1s���Wo쒷�*j��)X.#�<��&���&�Qp�A�#�J�Cx�����̹f�������dO�>0��vf� ,�]��j㖷�͓k�{fP_��o6<�vp����+j����R	4^��7��g޹�����*#��~����"�|˭H��Y���+A�^�YEs������'��.�qԄ��������6oe)���BN.'�Y`�����~c�o���k=��l�(s��W�������c9"w�֝׻�J����L�(��d�q�㡤���ɐ�Y�()�%�Afk;5����f����P@��	J!�et�����1{�� (#ćw�ʥ�SK+d'���[�g���@��jӿ�G<�St�f�y�̇z��v�(K��,g��p��үdb��EH����V�C����K{-����|K��(�6r*XfW���s�&#�8����^��)$f�f�ܵ��"�Y�������D̦ur>�^�(���(�@V�R���A�xDc#���|@0�1�Ί����w��^���DrVW'h�����S���{ᔎF���[e0��n���1�2Mm{U���7��z�S�@�F�O�p�e��*�S�Ɨ83�~0�K>8^>��w#/��֟�ϣ*1��D�-�0ߐ-��C\&�!̣Ǳ�k�Ԋ�ۥ�f�W�օ��:�g=
�
 ��[Q�p} h�&���&������Ԥ/�3�,$�W��|>�r���e/;`nMTB1 "�4���M�Zޒ�u�;/~C���xK	�ߛ�M��6u��Y?�[�z�������d����3[ϯ���qz�_�khl��<�x�����bV�~\��W�ǲ�*���O�<�H�VNlt�/��iZy�.yXT�40�3�)��h�=	��4�3���h���Q�/��őM�2[S!O��Э��&6i7�H8^�y?�+ %[��3L�pIf4�UX��6��?�*�T����9F�%�Ԟ�wa��?8��Gg��v����@�OC����2���q�%�{��!���.7��_�={c�����wWk
��@\<��s�(���#�����-����/6�qq`�C��o�S�KW���Z8��&��(p�����|.7����ۭd:I%Ǵ�@�l7!���N�S�(��Fa�"�[Sh�~�B����c�����{���C��*K"3p`�sGO���'pZZ'�2}f�̻��f3+�a��@�Ɂ���֮�ϵ��P!iĈC+���F�o���������z��U��\L̛�)��P��P����l�kHd��T�����o��n22t�tD9����P�����|��(� L��Q<���\=%1�d'y�?�dbtW��z�q^~��B�h�b��bhð���7�A��J�2��72���ʐ.#��"����[�5oT���H��_��G�+@�j0"%� 9BE���]���٠P~�ؿ��j&m�^��םז�K�Nn�jd�gN� s������T.1n2V2T`K}o2}p�͈��=�^����5�!'R{/P;/6���6�|�ݟ��������wE�μ�s1'�0eB� 	��?Mi�^���	`k���ӽulEPU�cUH��eV��?���}o�3Xv��n�r��E�T���9�룻�;�ޑ�Ә͐���UR:{�Vn�nNa�^�s�F���	- `��@��5f��G�Q���w�I����$�bO�FA��Dh+3(�랛��W��S*�
�M��^��nY��m��+����J����,ř�Lf�vD��Y�P4�,{�"�c�u�$ |ʬ=��ȥڇװ�p�sИ��/�pԑ�z5q�١�w�2r�}d�|9�M��Y�_:�X�ǂ��R�&���N)�Z�Q��݀9��ȸ�8eS�N5���%ks��ݏ���Vw�W��?�����Ҋ���_��38HW�kSC�(��v�B ��M�zթQ�u���Nj���Y�� �}T�
2M�S�9�5������)�[SoJӀ�!�j���p �m�r��Z�Y;V��?( �Q���F^=� eI���d�D%�	��"@��$; �9}��x����X�YL��n�}�ik���E�G���]�_��CJ8��@Z��B���QU]:��N_�(uI�ZB�X4	θ �3s<�����΁f�aaǬ�6�CQV����*��
fqw*�v9Uh�ϕe�]L�nAm��
`]�S�8�U2����?T� ׻*�>4��L�M�1�#3"/�V���g�+}:K<	<K�i'W�����e��2T�Q���q1`����V�Z�G�)�16���L�ܦ,�:��8˞9O��Y��"��ay?�-\��\_o{_�ƾQ�hܶfp��x1�V�+�ja�zA��f�M �SY@>�D@E�N�]i�?�e�����Pa��� d綖�e��y��pA�t���y��R����7R��0��؃�`>��'X�0�]��bBP�K�q1?@-X+���I��d|,5h�<�D���z�͎��{.�N���Qˀ~��+�:5���4�v��� {XN�S~!4�jPȞ_�3Jm�SoW7�,�`
8K��Iۏ����[��U���[��b�LX�����(Ǝ���b��61��%�;�|>�ҁ��?�߶׌��xٌ��)�@��cc-��jC�q۝E��8��:�4��|SR$����?��T yDOc1���r�%�mF�[�����{T�4ɍX�'?R��[��8�O�S9Ri7������ a�1.��3X�|JPA���Tf����ᄊ I�<��΃O�l��;=iX�R�(n��j�5t�4�����ɋ���aOZ�goW{�3�09Ѥl��?O;��U`�8�3�Q�En��fXp�f��X���o�
3@N����sS
r-\�������Y���ev9Jd�~�H�k�p��4�&��?@eU��/����Z�o��5������0�C/a+m�6�-}-9ޝ���� �KQ�YQ��g�̸��N��mơYN���h��؅Jj5d�&����EM���ȁ����;��(�� �$K�)�1�-� �/��#�v<��'��@��9��kȆ�S�v ��qQ��C7�b�4?�����cI7
,�9��T2���A�RQ�B>w�NʲN8���]�Pr����r��Nt���K)�۱u@��uw�Ww������r�6p��}����+g�I����(��1�0b��LN�H�Gs0/^�w����M[����l�憈
���m龗�1K�VZ�A�f�km�f����a����yRhEY��K�h���OW9Q�:%~��!.ykݘ��uK�;� 1�C3ò��)Wx�+V�5��hRϱ,JX+��u#���P���]C����X u��<Q#�*\��;�$B`�K@�Wt\p ��(�U|���#| O��p�r;����g?�����cG����'���q;�I���Z�:�d�f��tBE�ǃ�eȩ,��Y�9�i/�|�4Pv��B�J�k�uJ ���ר�3��0e@_s1*����~�"����m&N�+��Jd1͌�眕/�C���;��������hn"`�k�cµGOrݤ7Α�����+�ޥ@�?�X��Y7�?��{��-\���Hb�]�ջ*�*����Г곒
P�~Os[RԿD}B6���$<T�g�U�CU����"�AP��-�q#��f��<��bHE���6�h����U�H<��mL������nHnڰ/�]���p�G�Q�È-f�6�͙��=2{�l:{YI��XX�dd� �Y�I�K'�,� �����mοKn�E�U�1��!��� )�`����=D�nGL�� ����F����)�S���D��yB.:֫������"�h.ui%7�RX�a��I�z�`�"F|��=��i�
~2@�.��24�p(V<�%���:M3���_eF��+K��Ϝ�l�~ɝ��(P[�3�s�������,1˒�a�6����&�2��_q�D΄��vt��M����^������x�q����)d�tK��t4�{�Z�`z ��Nv��a�/�[=���2���:l�v%��'�o-*�3��|�i���D(I��1�F��B�a��ؚ���!:�W(�U`�]T6AX�����;,ѐy,ڊ%�ƚ-*��ՋC�"�N��K��ϧd�䇧���1�\�},�K:a2g��%~m����r��j���k�-=k��~�On�x
�r�����}�C�?X�G�>&��N�[HEL�r�%�DDP��o����<@n���\���s
���U���s�m�Ͼ�����<�~!�s9���l%6�b_�V�/j%�WC��]Mu�>er�nUi{+Lp��<r�Y9S�͕b8<qڨX�]�%H����qQ�m���)���'�_��56�e���A��m�1�)D��|Q�CR4o�n���F��΢�7uR8�Hj�4�&
�%J�~g�8�/�(���hK:�͝�o&3��{o��M:4Ī�O[^����sO/2�����}�t{���Ꭴ;'1�����;ۇ�k��m��&���zT=Ȑ�U�b�/_��ϰO1�GHB���XP�*�v g��׷�=[11���{"}A�S^�C&-pIH�K��?x@Kӡ��c�6gtf�Fj��`-kh�+�6����)�;J{����n�?b8	E��T	gA
L]f�i3���8��~��Чn��*,��x����+��Ih[PJC=H 6�p׊�zz�u�0��UpF~�P"��P�dZK~�g/�ۮE�]����u` ZJ�m�� nT���.7E��ʜV������Vi~��
������?c&H~��N���u�`q�<�ԖJl�ڽJ���lU0�q �E���k2��wMx���^�Q��:m	?���j���8�/qJ���o���=L|(��W�Y�c��K�������]2M	�eV��	L���>�0�Jڣ��+���O���B��/]�b�Nk���%GQ!�CZ�)� ��v ʎ��]�Ǻ֒7��-~fqf�j�Y%i[�f��q1ˋWa
�
2I����bj-Q�^2���V�~g|�u�g;�a��g�& �QG_d~(/�h��/l>�9���H���L?�n;{������x�^>�^h�:ߢ�m���٘Wo���C�/8`��:��J������Ȃ�<�@O^8J�b��%류W*�Ak���(���A�3��7���	�B�X���)��_ܹ��ϿdNKu�l.Ba�;!��BڽXwP<��,�C~�2͊O4B~s���1���t\C>wgqz��*��H����&'�)*|#?o~�f �������"}���r�S2zأݸ^��>�B��Hó�ݵ �m^j8�>�Z����1M����lG(�@C��'#Z��x�	z ^�}i�:��_�G���=7��n|.�aV��Z�:1t!�CS��
mnĐ�C݀&H$	�1���T?�p e�%f�u�yxf����J����%��7J��c��5��h�YO�I��=4�K�qK�$���:O�i&#羥eަ ��몊c��|%��D/�m8�0�]
�@�݄��v�b� �4		y�!��p*��*��E�d��[�>ƹ��`���V_�Yq+W����$�)vT�1H��P��|�됉�\G�Q坟uP��܀�1��`�M<�<��i:=��.NJ��u���g�T=��C�T[&���f<P�U)����|c�	U��ZC@���8�qPZ���\Zz��������, &�#��I�d���;���'�*�;��"y7�FHڄ���1ğ��jݤQ}~Y:�{�=j}m���r�I�)�{[2�'��CPc��&�U�YA���~K׏��:�.��P�A�$�M��%�{�&nw�q��1p�'��T��;рq{ʨ���3|4�d�DIel]�b����\�k�I��r����sz�W=����#�3H�j������g�עĺ$ߵ�"���K"�1��(,��G7M�L����.�g�W[��p:sv��ddqc�!J�����Q��K�I�ұ�*��Wɀ50����ؗi؄&\b��%�Ek���e8�tTs�/xp%��h���cnD�((q�u�N:=�^R������MP��׫��&P!�.!�#w�a'i��c���"E��,�Y@�"�	T���î@[�d�@��O���ͷ�b�tޯ���������$H ԋ6�����@��8NVseñ�̵���rCjC��ߐ"Z�-e�x�_/E�ƿ8h�@&�-�l}��Y��q[,�!��UV���59s���n���N<G�
��s
ȫd���3Q�Cb�*��=p��o~^�uR�t��Z��j�����֚|~���3��\��3���g>�������~l�ƴdkw�T�[��x�٦���_C��Zs��;��NT�����~������+�E�X7��I6��9l%*|���ab��#R|��RU�X+��)����>����^�V@��F���Q������V%�n�7�]ã3s�}O2]��*���XB��; ��3��|x��8>��e��̷`��g=2ii��
�ٲZ�����37�p����%���s�C��:�-JgqQ5�G����7��Iˢ��Ea�����5p`>+�Va,#M�X81�

p��ؼ�4����>S�;r�C�V(CV��f��L�Y��ӑ湟�l9������E2���Д��)�[��(���;�kUS�J	�y��a2 K������*3�*	���pXc�Aǡ)��:Z�=����m�����N2��}]��!��6/����k*�6�9��G%pM/���Vh�J����R�k�?]�)���4H�V��bj�U��M�5��N��^�mE$��a 3����diE#���3�0�5�^�|�.'Յ��/��X��g^����%&�9�6j�>v0d!jx<�o���߯�͸�'wͬ����iV�K<4I�֞���T����K����Y��Ŧf� �L��&jRB�b�1M��Ƣ����+a��Qc�z���W���������4#�!d	�϶Z9�d}�����}֛.}�]n,y�[��	��l��wW��)���Dܜ��tPY��
+�F��+4@�E϶1�س���]���(�S(o-�<��tF�&i[��$ �Q�:3�T��w��P�+��`u}��/�u��� w=���z) �֖���c�Y���B�.l���^*CԹ"�b��\�"����G�a~�#��S۟\����1y��Y�����xL�D���j�k�6�1�������t�[�:�=F��l�竞��r!F@'�ǒ�޶�շż��F#Q�Ph�F*�`�
�eT�%�y�[u7������������ïA��h���D��%���)��+8���h�^��.��,��A�ɋ��	��[y̑�R�H�AxQ	�g����& IF����r@
d��*%QS��F�E�ߙf�r=mV�1�R���#Zv���O٣7�[�n�=y��O��eEɽ�`�����0�D���^n���1��O����9�Q����d&&���3�~����y�blE��Xw�Rg�?�?�*HT`�'��T�*���.�d�ttl�����ʞ?\)$Y��|]Ԓ08"��a�Ǵ�|&;��P��j�vy{�Z/�H?�)��9�~"�Z�rΣ����d�Κʮ�p�Hv|b��B��DQ�j�(�<�M�����z"R�N-���P0��<���%U��9��mq�,g�����cһ���G�3��V�����D�j<�і4S栺D�p�3E�����n�rQ���]���QN�{�:	�������L�}��m8&���&;���Ta�p5��\=bS��`N���Mϳ�]鼶���J�����/��T��\S��;Puɨ����x!��c�Y�Y��Qa^����YZ6>X@���N>G����N]m��b�bݑ�9g��{%�����D��΂�ȵ:��ci�S+}�����/�E�/�',��zZ1���oNM�����Vk��[���`�-!"^"�6�1�^�]�H��41W�x����׺�u�hgp������ ��?�n�Ȯ�{�k(�j�f�s�o�����;<+���=_)�/�+�c\U?,f�R���^�;ś��M�[:�����~��8p�K%�	�q��@d�Z��]�s������]'A��,�����_�� X�y���L�R�:=!�T�)��E���\"�A�� ���8�2� ^4�|V$�I�8�"7���
��K[#�T��LQL� Q���O�۶L���a;)����W�ȞU�r2���1s$??��2O���_Aa�ɛ^��h#�U�J��>Þh-��?��1*M)E� �c,�(4ݻDa���ZUk�����fM��bׂ]Zn!������,}i�l��������W�������y�b��<�(gXn:@`��Ώ�֍-7i"]�p�g�3Z8測��ȣm��r��[����s���I�d���:~��t�B��X'�rzS��W��иfr�:�E@#�T(#��P�,�n�f"A����n:��'1�x��z�t.���ԏb���&4��Q؎�k��S"���\�G6w^d.���/��l�[SQ��QNͤ	eEh[�C��r��5T�p����!���]�,H�$�ލ��؃vRU���4�V��,Q�>�:��j^t6�8��(M@E�5�Nx���	�H3�&�W(�ߒ#��I���S�*G 闃sq+H�W%�g<#�R�M�>��I�#M�xI8n�Kk	7��b�-G�L��9����q`S��&����w�%F�]wk�X'F�v��gO���f8S0r�!�i$%�f �x~�\����J�}�1�G}��4���N��0��"�JE ����LS�O�>�F��T��y(�mh��ya_a�����z0�/�!�������!!��3�W�`5�3D��VyR�ӎJ�=r�)킪���LP%�A�@�y�yOc�[@x����CI5A*��G��g�^��p�|z+���WW�؈E�3�<=�+M΅����T���+؁�������u6���A��L�v�W�;i'��Ѐ��屈O@>��iS��G��e���n\�
vcN��7Ax�{"E�)�կ�L�'T�|Ϟ��ꋫ��oS���ņ�;�Ѳ���v���8F���ҠGaI�];���\��{�G���f�w�O���N��X�q֞ğ���й��f�����[sK�w����t���s%�pԤ�vb�b�c��X7t�}.9,�]�J � ~��eC������������\D�dH�)�TU�ՠ��6�鹄�����S�曟���|ij���iS&�6�͌�p�0ߋfi��#�J�K^��(�_f� ч�x��x�������MB�L���4̪.xo�`Z��]:#[.G϶�1G�)������Ŧ4
H2�Ϣu��/g�i vh��,~ �l�(�� �:��+���k"�i�d��F�x����^����kO_
�}k����j�j^hmJo������
�\9r���/�-1o��aWB�3G�l��S�P� mcD�GC8��ics������䖘�ד�#('('>��2���%�����`t`c�U���B��3�d��(F�V�%G�\R?�F
�)���t�&nx��8X��7�c��Õ�f��W��2G���g�P�܀�	�l<��Hg.$�K!`2Q���΅��-�o~J��N�9��!%Hp�pB�Kn�J����2n�)�D�����g)���b &s3�����ܠ�w�%}����A�	!�
��6�6�O&�2�qUxz�AZM^M�\������a�$v��s�� �|���9�z�Sl�����
j�q�����7:�Ƞ*
U�� �t�8q��P&��<�J-��y���ĵ���7&��%�|՝Eex�D�~#�g�V����(�2.m��g�Itꨅ&7�T�V��fY|E�O}�Pj�aF��d�n�k�{��狈V���A���?��R�>lQ���Kg��>�3�2,�@����?:�$��LG%/���H�{�mp��8�q���'���]�
���s:�YUE��sS����h_d�>�xR�%���h=<Uo�|`^��e�����9C��F)کh{�����5�2������܇3Oj�h��Dn4���2�?��Sh�	����_��=Ofu�,�Ց���8��s�UZ�Vu�o��iX��F��Źߐ�W(^�hc6z)�4ڔd��k4�J�N��v���U�Pu��`�7{g���O:iK=ҊI#60���tR�q����PY���2٥��	�l���}2������@�wLT\�f�vyB��^<�rNͲ�kR2�l���22hF�o���M�ܳ��v}(�:۷���yݻ�͎��h��
j�Y-�cW�+p�����`S�D���?�_:���1�G�2	���`m �ԭ'4�(L �݊i�}(b+R�ݦ��6(g���}����I�Y]���e����K���+��m�2! ��h0�΍2������8�Y����c��gR�X��<'�������OG�f�d��j/�GU�Y.��_���9 <���,ȳ���!#���;��,Դ�����6U���~�.��	my%W������l*Y�%�#5�	��R�/:b9B�֙���c2d��B���%��1���Q��
%m��B�D��Ed����<w y�%���/�q3��ϸ�d���uƻ��Ea��2^�3�.n�"���"A)� W��0̓.@]0-/�9�
�Q5L�,�b�l}Q�n����5t�X�Prc�5ؿAX�*rJ�ṧk�
3��n)k�Q�	{���B�w����|۰Wz��~��"׳%�Ҁ�'���?�Rv�-���N�]�n���L����5��
y���/H��x;d�Jt��ב��:S��/����&6�@a�����z�XE�wڴ��xk�E}j�\�MC�׿����زF�EU�����\�1!&�K}3���b@o���c~7���[�3��m:�u
�{� �S��z�7�vq�)��l�2W�XBǸ�\ٌy�Pk>���[�V4�����tU��v4uC�Ɛ�o+h�N=��Ʈ$i�O�
��&�XP�m����1�N�0��)rH��<߬���[���Yu���1+�����JJܺ�r���\�lL��yviF�g�L��ɴ��{��b�~%$�s��,|�"��8	�J�o%�۷�8�ֳ
�bő�r�gJM�EfW���^�gDA�R���w��h���O	[wI|匎H���^��v6�8��Co_�Z����W�E���w�P�Z���{nr���7��ۻ8p
���P)��'���I��tܼ�I'P�i�[���R?:E���T��a K���C�b�h�/��8H����i:G�����Gr�;{}�$���VL���DFƣ�^6�"��0�2���GiÈ��(�\����V��[_�%Տ����^�]�b���O���YSe��t�?�W�^r����˫��`��ׂ�Sr���s�tQ�)z�I�T�������O4��9}x���"��\O�c���̕!mmi1$��b����c[{�/%�U����w�v�1���°�o�\i��n�}�ڊ�]vX������U�۹m�TO��f�1�Q�^�Dy /T;���TY��%=In���mG��q�VT"����@Q�5
�>����l9��D��p�ǃ�F~�ٍ|� `m���JQ��F�t�D�c�\_��W�4���Q�GS����6e`������&:ɺʞ{a/3P4�6h�C�VM��D(���P�^a{F�����*��+O�hcg���K"�p���~����g�����!Y������ueC�J�=
�%ce\��n��a�c�͓I�^<�3H�؃X����wh�l�`c�z�Ğ,�&}��1�0�|
�]�z$����9Ѫ'WE�E����"Vu��e�=+�����ޜ�(o��aMt	AE��$�4u4�,���0ę��F[�2�0k(qL�����7��^+�*a��;�'¶8��gS�-79$�i�;�
[�W*'���̶�_����$%���Qu�x}���Gp��vb�h������lv�+|�6M�3��:�0��\dx�X�?l�k�à�2�Q8�t�g��d��kI�qzI��-a�O�{n�a��r�\F�È'`�AѤL(V���h�^�/k�#[	N���[
�;�b+�>���eߗ�%G��0���Tw�s�AL1�A�V��W��t\��-�lr�A�����������*��T�ve_�D���/9;��m����mZŽÂ���ʶ�����s��4L;�E�6� �C M~�i�
2��[/�����W,�J��?������.����a�`O�ۨT��S_"����~wOo�������ֲ<O?p��,�8QT��[��1��:��)���v��0��̒��o��_$����7�=��Y��1n�;l��yX~Q���)t�H�l����U3�譑��s&#��`OM�Id�E񻽘X kp@�
�˺n*�5������s��B�����JS��d^ +D(��7��$��S�!s87)k-���?׊�r������U���2��=��q�mc�p�*���`4��:��9���d�   ����#������_�Y�C��H�S�(e���?}�yٓO�лC�����}�'1C��V��\�'�ȃ1+INi<�e�+�~����j��k���jf���Vf0��FGy����������$}�r���̑��5X|����J9j'#�xI��Ɋ���za���Ǟ��eo������&Kp������zx$3ĳٶ8F���GA�����b��d����B��8[f7�]�.�[s��bU�mHh�XU3�3��+�x�ʩ,���,\܉R��&r ���/nS����x�S��B��_'}v֔���HE��D��UY���B�	\��j������k����3Ht�:��KF���}D�U�t��Luf�h�N�8��1�J�����jM�6��GcQ���z[3��!y.�K��&n_�e?~	�[�u�7�.s�BHL�dD����o����[��ʆ�#
Z��ey�b=�J �RY�}�m,���qDMJ���_�l����4�������U{2�u/2`�W��>O���/���B��s�KI�5�M������r�w����$N�K���Y�����O3Ƙ���Kq���0�@R+�LEJd�¤�tqp��yW�n}~*�F`��p5��Q�%�ҚL�z;�O���vR̳��.�,�h�r-0}��x�Ss�B;j��ևuV!�=���-�C�V�D�)�6�%�J$�� NU��6-WW7�Xg��0�5�M���E!]��y ��{��̜��V���["������g'�;�g�b5Hձ�N��N���v��S�A�Σ���4�61��%��
Ҁ��k�6�a�t�n�t����|�{��

����v(г��^�I��U���"�L5P�Y�i�^�3F�Z�ְo�le�ÌB(j�|�>��Cd�q�[~T!^ɇ`�Z��\��}���Q´Im��\�'-#���#00���m���o�2����3� �A獔��n��q�ݾ�E��_���ltW���UĔ��,3� �t�� <���Z=�u��i��-o~Ĩ�WG��b����2_��C������F6�ѻ�J���k?O>�祂֗�5b�2����"��d��������H~=l2����I����ύ�^�:≦��������v���)�b��T���?�<X�J@�K�]g� �XD)CriE�����A��(�ZN��W����BW�~1{K�J⛑ǖ
T�2��u��cV���$@�3�E�$WړD���pl���i�-�J)#�OG0��N�{�A��Ł�`����e�`������4,�h���)��n����� A8k�'.B>��+��}�ݡ���3T_#�ǾO��6��Il>j��W`�o�z�ot� =��p�s7��.r��4M>��f>o��g7�t��X��j��1X&0�yV�r7��3�J�N�?���\�����#�c�o���i(�׃����S�m��o�PN|\И*Hk�w�c-�������w���ڶ '%����X������0��G��a�fx�f�l��L��xk�����
�X9��e�"��G��U�Z]���%���J�tͤ�=��:�M��Cw�����(�oS"e�'و#/�_��1S(�C�a�./�B���,��m����3�J�q�6�B�P؟��+qu�<3ؗ����mf�{�y|�j�����8�1K�3u�@K�g�0�������{�jM�A�x�R���mzٱ���F�GHu�}�nA��ԧIAx�#�mW�"��?��*�2����������ݒU����U���l�FL˸-qҘ$��\Rx���Rq@�Y�,��� �<�#(�뉷A����Gĕ "?a�w���
�a�2�M�̨�L�BZ�{�D\WC����Ǥ'-F#*��C���پ#W���B�D0W�q����Z�������W�BC��jj
]N��=d�I���0\ݝ)�C���(d��!�P��;�l��ì������H��/A 9�iM��.C5��Ƴ!mv���QȄ:v��!����n	K�l�m���9; |�+��<���g�9l#�e6���rzɬHjW$�P�ի⩬V��ّ���s�r�u���_���"�$�1^��xCCw�ֱ`2,\ՠ=(^�b�e�ʿ���iO��e1ؔ�%���f��U�`a�o�B�N5�R����lB~�����H�YঠQ��+� m����S���߷M9����v���IGp�yg��0��!��$�v���o��9
C ����G% *��(�!z.p�ELϰ+�H�*5ӓ�aP��6�[��&�x��P��y��'Gv|Gh�ݞ��PiHkK��v��iy���t�:q ΁a����w ��'ru�
������2��ӛ�W�)w�&/��w+!j��{����|�#���-�֘8t�g"��S�>s����!l� H��?�[GSͩ$/L�S�dp�S���}�aM����}X4���!�\s��F�k��/��n^�(���������_���$Y�)�&��@v'�<��27z{�ZG y��)m��䋃g��i� �T�K��79���C�2��Q��'� �,�d���K(~����h���3�d����C�Z�6�}���,6k����|��б��Ԗ!am���ڵl۠��'�\�?E�F�KR%��GM��\������\�%ᚈԞu&ɣS���:�mKQ�0�t���=d�R ՛���Cl{h�ϐ��Z����J)���!���p�"4�<L�1�Z
��^��;��L�E�	Y�^Y�G�Z����*��v�*��A����i	>]\�=�o�Ƞ���&7̋ChD�R�R�����dtҌ+� �����2�u�	),o�!������b�'����ZP#��c���B ڑ�&�~��}��7�q�yPF���ĩ��a�U�E m�	}�SC�qݮ��R�CV��^���91+Bl��1�ٻ���d�.����D:�tۮ�@c�[X���Q�;�Q�_<\�ZC��M?��m� j�+�
6����d��O�r���W������
7u�'*.��4W��ր2hq�-b�I �\ܘR��
[�EC�Y\>Vc���?X1�ӟ�Q?G�`��1��-"���p���䯌��D".�?
KJ��]��#��#�p��>K[�"��9�����oru=hFL�5AX��%3��|���ۈx�;.��2{&z�/�L��ў�˂��1�_,�
ס�l�:8���k�zi�'���<��`n�q�����1� ���v�9gh����+4���f5H?w�`�=��$ڢ��Np�� ����c�!>�n�F�m,�k� �M����u2N��T���{�G���E}nV[r����OZ�2û���,ܧ2�>Ǣ�ny��g����#���I�VH��6/nEiX��y��&�ݳ��7�o1I�+�@�����<��KQw�R��7��P�,2>�Cb�^T3{����
���b�ʛ:�^>X�ڗ�H���U�˵��E��a�
��)Xa&�W-V�����g�z,��}�>_�R�ALv�].%�raN�dpj?帰D�K-a�h�������ܴ�lhƟY6N[�yeV�y���z����|�wN
�Ua�G�H{Z���P��F~2.3����[`�l��i��	,;,��2����anņH1��H¨m� ��[eNM�6��8����k�3v��c�җ�[3�3���o�|���K=�Z�Ų���臝J��xҔS�ul�� �	�x�ͧH�CN �B���ON��[<����u~�4Y�d^��^�*;p%�L�-԰[�%�WΠ�܆�R��YB�x��_�u���0�\�
��Ze։���K^�c�DC8��pW.5\q^�\�Y���~@�!m���s����Th��|^6�0����N3����k���H���֛�$��@JvȦ� �PK���X蹄���9����E�?]|��\�.�J�״��ۛ7ٳ�A�~M�Y?[��)�X��<�*�>N���κ�l7�MNﵜ�d��^���R5=Ҫ
����ƛ �]z��?]����,�G��V��e���R��9��C�$Lz��%�/��y|���TK~�{A�A�1#î,��,;[�� r��`���N"�&��i��9��(�+����ų����B$� �Tk�0���=W	;*�6��	��9��sY(x~U�$l�5sz���\z�<�/q%a�\W-�*g��/�ϡ �� 8�X�H�.wvK��c�&老�I��HO��.�����!xX�xa�NQ�SN�:A<�o{y��� %�^H�N&X���K�����-�Pv~���%��!�G���*�״��7�8 �������^��M�:Y_.��sq��0D�O��	���������������t�k�b�f��p^H��P/�;
���&<{���ƿ���*2�/�Ux`��w�<'��W��޷s�ʭH�yM��4�0�0 D�!�ݰ��	��n��M9�*���(�c~'~�f$�8��6��Ii˽�]A��DO�		��ƛ��v��}gW�X}1��X�Im ����������A������?�H�3=ܜ����i�!Pe<�3��w�C�V����3c�+�i{4��'�
:���HBP̦�ɢ��Q�|�=��4�_�����z3����М�����Ô��q��HK���:�Dw�]�t!Oo��r�@k���L7���0�F� c!�J�tS�+)�*y��iEaR?�,\ px�}vo�B� #��S���aE��p�ԭ�G��}}�NT�,�G�����NM���-�'��Z��~a���Rm�܊��N&�A��N3N�c3�wNu����B��h������y����
T$��ZV+�C�Өsw'�)
��w9mc[�8. ��{W���W8��#r?Z9l�}�����r�]<&a&B�X��%W�99򃒽����=�u&�3�hW�\F�3�ى/�`��bNy3�d&|�d��(��),q��� j����|=d׃H�F�M�~���ʘ=��
_��h�R��1@���Y7Z��H��m���#�6�"���S�sP}w9����Sm$؄��~���'3�=ˎ�L�7sv����cZ���IS�|�8N�6�Ď��a+�QF��ײ×���T� �L���J޽d�~�_�n
ނ!��??_P�F�r)�{��í����t�h����"� x�
���0�����nH�`�W����N��|�s��#^���~���5V�g����\?�;�բn�!m��J+Keu��:?���n�OoR����.��4����#�}�b��4c��W���|f�1�Bc�Ad�ܶT�w��\������'�%`G`�B.��i�8?�j��:���c�����W��J;������`�S˚V�7"����)9\�;|g�d��nT�`��"�si��Vk���w;t`�'�&�*&/[t.��X��jˌ�z-�b�s��H����nNB����,�~j�����|-�}�Xd��D5�$�iF!�t�m����D.u��b���MT)n�0�^3�������'[��z���(M#Q@-`��Ҫ�b���c��6o<{$;�+����~:/I䁕�X��rH���T���:�_���Fr����6�V�%�� z�3	�Y"s�h�?=����(��A�*n�����<k�NdG j{#��5^�{�/��/���r�STѳW��#�}����W��)�N���%�$
B=� ���}�cB؛��뗒�#'�xK�؅25��n����G!U�rr��5�h�Ao��ĥ��q0Y�2e���yR���U/�(����xOCo�7�a�a���;��F{�� f���;\b��A��T{z<�N�s��g<D��Q���o����E�b�)M���$�s9�C��i`_�!n��4'�Aχ&�Y�ƙ�����4���J�ʐ��?.v�%,��8)�p�,�!��� �,g�������'A+���U=�N������%��.4�>����P��F��*-�`0rw�zu��ζ�/آ�n��Ah��!)�i�����7_���Q�}0	0Me��m�k��i�l�PS�e��M�':�#$���<
�v�&�9)6�N��Çx�_ޞ"�����d�a�짧�⸪��6&wRј���W�,h�y��=�L5��$�_�Az2+���QeP)F����Aqa�-20tj��a�Eҩv�����<���B�[�q�c��L��}������p��X�l��vN�Z �;�1&�Ѐsp��E=�Z�RP�f�[}6�i	B������n�;�ڧ��i�м@,��ͻ��#jD��HM<`��~:����2�x�R��A%8�m��2v_4�}��Z�ڸ�	oϬ�LA���ʱh����B�p�����^���E}��ڍ��V�[��C�fCRhd�^�������b�
9H=��P����ZI�AH�4�u�h���'!�@���~��OG�s^�}/���mD���d�[�J�*7|�S�3u�8��A�����i�x3X���ױZ���%�cѠ|�^�Ğ�J��%��۟P0�j���꘻������a�-�C�s������!��l����`�����i����݂�ͻrhH'1�j�U���w��/1'Vz�o�w�z���8^ţ�3��t��k
�l0p���_������8eP{��D�otZ���8����ŠN�[�s��_:%��p7�E=�/��5y%~!�K���b2o�}G�3wZ�����1�00l�5���X��`L�8ӊ�$��WK��zx���ƥ������y��{\�{Y�*E�m�F��)�x�R{���oC�oҫRC��>�'h~���7)�8���f%6D-;�W�8�}�"���#������jxC�inn�y���r��,U��+P���	J؊���ɰ�$���H�Pq�[��ʌ4�\����{���u��D=��0<e�©��"z������D)C&�����g_t�'����|�/}���sۀ!C3h��.�����bDR��}?�^c��g����!bX�er������:����H�������p$ڝpj:eq_#��&��O�_Y�g�f�)�Y��}��D&Ia����F��?1R�@�4sB��ɘ��9.r�%q�[ZgLg�zr��km�Yk�,B������D(�%�ҝ��\nO��^��'�����-Qٿ��3R�-x���a�;
ўr�p���2������=�1Vu]����k���-����3{ф*���n��}D@"�`�DDq�mI���j��g%��
K@����=z�V�y�]*���r����2¦���gp#/PAwIפ�A��#s�` H�8�Y�i�s�����S pi�����gZw�g�v!'\r����9
j%ߵr�.k�g�m��j�93��p-űT|���2��
f}��!)$p�������Hq�'#L�JzJ6�dQ)���h�R��mH��0aYQ�����;iT�#� sp-y!�.Z���с��_Ngelg?bt�D(�>[}J`�x�6=��W�IT���y֪L��c��&ɠ�m#ʈ��O�1ֶm�:�C=�X�&�F�.[t�Ɠ+ʞȼMX��]ӽ�#����2��焝+6V���c=A�~(�.�K�T:Ht�Kbg�f}q�n(X$o+l��&9@����Q����n�D�����o�e�b
��k���� pz�>d�x}~3��-cI���#���^-�э��Y&�Y:�;mq=~��t�R�X|�v(���v�@�+L3�T���.��u��f�@C�G$K�1���o�U��:<(šL��
�~L46U@L���8Sv%Zh�����Mؓcۉ٩�v�ob3�x�p�j�|b�k.zj��j&��*�է�������;��6�R8��٣c���Dt_z����H�9C��cҵt^@��E���Ј����:9�� � ��m��R�)x�K��ϡ
H�_���v)|R��-0����Y�~ۇ�w�`w��;S��fS�-�^�[KZ*m��vn'�S-��RS��g,� �E�X}M�XO�-�tl����c���ԣa�Q���#3r�ކV�Q���777~ k�,��į��M%�����»9sgӨ��g-3�#�C�Ҡ~=<+���qk���Q ����� x�UU� ��(>�X��;Q���!���V��b^�� ��:~�Y���������;F���`�� L�K[��T"ЅE��.d����$whW�]彡�Y��l�'�����M���KE���+�A�Ŏ���V	�iû]������`��ybA�Ь�k+��M<���@�E^m�VzYoƫ, Gd�q���?A�x�/rx�T�؏L7X<��ȦElH��#� ���{E�{��t�������C,&��;5��.L�_�N�Jk�%�>~qWA�^So������J��Nx����m�����Y櫀�4,AEkeEc�������&���U�?�+T�~��Z0�*�i���M�wU<�<� J��E�:CC���<1Ų�L=��ٜ�d�j�4�A;CY&��������C��t��窟������;�C�8��U'�7_�K��1ҷ���z��6��j\pj7����)�2w�,~��f'
d�閮�ZeH�q��M�$�>�<9ұ�D��I��ENd�n�s�\Y�d��}ֹrN��
�`&W��ffW��k������uP���e�]mã��R��δd�F��+��mp������~��H*9��C�S)�( !�#h�;��7���f�&c���4��	�b�ᙧ�K�"�_(v����1�`,P(�����+�s?�>�ү�6Uz�w��#v�����@?a0ԥL�����k���҂z�#��Б�L�?M��L��UT-��Q`aeB�B���c�D�<.�!>���Q������:w�?�2;7kh65 �B�c��E)A�}d����L�'�
 D��E�i#�qec� �񤊏5�*i���u���5��&�^N�*��~��~�M����sһ���=|�X�A�-�2{O��:�mނ�3>Q�?=�h��U2(	��	T[�q�3>4ٗ�!�Lt?�~����K��u`b�z{�R]�|ڬ�<����*͆�'��ai�C��p;T{��.�k#^@.�ׄ[�.�b�6���=C�O{=��I������ �a��й]<�:Z
~b~$�G�I���f:R6����Lw?j��<����PFv	�B�ۇN��ᾓq鳬��Հ�*���^�����D�cq�PM�0��$���p1U�5�>5d���@���ƌ�ʻᛦj���Z��dٜ��YTm~g�y-q��ދ�F�uH��Ϋ_��y���O9|y�D�n��U���"b���F���jRKb��6�õh�0l7��=yy�	(�YY�w%���"B�O�B�n{i���a����+��XR@�~d];�D7W籭�Y��:��S����9N�Ubv�H�!���J�,��PC�i��&6�nG�5�ܻ�"�X�1�)����I��I��	'գ#*�_
�Ha���cf�ƒ�ɏ���o��	�̵�g��ֆ����"{gȖ����2��g�V z���Ңm�6��Y}6�� �_�xB,Y�`x�ρ�Z'\1؅E�F���=nڈ���R�9n���S���Nu�%�q_��f�"��h ���ǳT,���	a1��v�X���
1�~���d]f����t��O�f>��B���Zн���aw{]�%g�>��٢Ԟ]�i <���F;�C$56~#��mJ��r����.Ul�y��\rN��ou}�}�Ȧ3e�ǳ43}f����ΊV�nh��l�$Gl1��Z���L�\�8��6TB�P����+��O��fm��E5m�8�Cܦ`��������W�7������XN�6���d�k���s��<�[u�ڔ��G8��*���	g�����S%G��s���-�29?�F�}a'�/�+:%���f�aLu���x&��:y�j�?��� �ڀ����6���U��*W��x�w�Ձ&7�#���	W�`�YҋS�������� �i����>����>w|PQO*�|�m�-D���i'^&P�+�ܚ>�'����M�x¦�Π!/P�y�}I�t1.L�#ս�F0Y�!����>%���1_k'�EX��ŀ쾯n
��P�a4�gzޗ���J\wX&��P�3r����Υ�}~���n�z\�r����4��u� |$H�b£����A�g��Zr^���L�J�P�S\:쾮˺�x�8?Y�!)�-�uÓ��e�W��nJA7D�$M[�	7W�N���^�!�{�Ю��p�v,wBU�����tX��*5���6g3�ċ�+���޵t����٩-��+�9O8�[Z"���u �>*�ؕ)']�g�,sP���
6�܈OK��+dCk�ύ6���;�e�I��L�-�w֙������Â�&6GVNs̐�����W0�<5�W�J�u�9t*/g�/�j� �W��۰�Dܡ6�̂~Ҙ��w\�<@B�]9=�Լ {��u!(q�G�U�ʹL2!�0Ŝ?�T�'�G���+Ԁ�8����#rf�^��;i_f��&Š���Mb<�rYI"�B��>��c�e&_J��cA��\=�k�;��{cV��!�L/���g4m�&�~���ʮ���=H������"::6�GnL��brX���_�G�m�?�"�#M��p�=��i�a�}*a�O�D&e��ؿBN5l�p�;(踼�H,���"����6���@1������l��*Y�R�7�(Gs�F�3�����M����1�}�1jMZ��"���@�7�"i�f�~��7�P�+[kt�d�c*ءYY�<����$ �QDD4�0'	��������g��Ԧ�D�"����y����Å�L}bK`1���rn'4����U�'�{w+��/ɼ�*"�%����}o}�ViA�J!R[vX�A���1
����x*�T47ϫ�c��$<i��OP�i�;����Urk9�@���_�-�
Qƹ�W0�bc��P�P/B��{��c���a ���ePC�&�]5fC+jpӎx��Մo��b+�bU��������'|&e����Tz�J���+�F���.�w\�T�z:W �`��ˣF�%����G����7�%>�ڻ����E�e2F��(e�$n��﮷N��=��|����n�|���-�$��ׂƹ�x�D�]6�D6�	?U�y�jB��Ҁ�� io.
oxi������j�"}���Ӑ{�ƴٔ0��iO5���z���ټ����f�8fީ8�}f�E��=%�)����oj�J]��\�_�vN{?�dr�Ip��n����	ݙ��5{k��|���U�Sj��]���k2ۍ�Y/�lҸҪ�iC�	�E5�)�a����ra��]]�=�r��+�F����vnYW��m�j`��,8Z�ŵˌ"�{�ԐԱ�����լV�I���2����:V���35�x|y��ŌhޭTQ�Ø��v+�iE�ZB���Y�[��|w5oҽ%;��JY�-��*���I�!k�]8m'���̟��c�L�a�ݻ�t��[����H������_��ז�Usӣ�m�:��hZᅣ���㸺����C��k�'�A�����2E,�v;Z�����b@�U�C���)�{�o�m�'$5���F�^G�������^c,pԴ�׋$��B�hs.{�7�$���n�����T�c!i��=G���p.0�]O�8�va�s�m��9�L��>T�ů=�$�_V2�)[ �P��g!ѧ?���\�������O�G �����'ӆ���Sp70�y�q�I��Zy���7,��ra����R�K"�?�(�U�ډ�&�3��r-P�.Ԕ;�]�m�w1+)[?��)]٩�1�#��O�>�Xg��u�����oY�DTg���35, D�k����yw�z����9"ސ&��~z�(������c��&X;J[�flvF�B����l��g]�LWt1|�$��ɋ��)n�R�J���z|"*�����C��s�W+��(=�?3����V��w��o�j]�ǘ$W�R��QvJ5�Ĉ�@ti��cPG�V��R.�����v��2-Ԗ��#�� ��RTFUj�I�}�V69ⷌj�_"����W�F}��mjps~�+���J$@KI���R��M(ȣ_ϥ櫎�#�Q:Al �	3�so8�;i��/t��'���?��J-]�2?���؝`��^S;>�ež k���2��!����9�L�2�m�gD�oa�NA�T:3]�>���Ӑl�Y���;bWl���Ų�g�OOcwΆPZ I�κ�J��h���&�b�!�H�N�'[���@�hl�/K���.��:��aAc<SA:j�h.�0���x%�\��8���~l�t�'�$Jc��'h�h�r�*ϭ�^.0�)3;B�!�W�l�_A3x�k;�"��2��'(tȟ�l���{�ɸC�b+/g�C3h�*������>�
n�b$��A��x��
�QҜ�6�4��Ì�ci�x˷#+�a����5T�]��_j-ۡ�]���s�4�[/����ycX���3�6���Z��(i�>�7�\��j�g�3k�t4>��|"��g2��2ۺ��W�xfɕ꒢�ݠ�
�B���",܊*D���%tP�/f��7�-t �戉p 9�6�רX/���\b�7�f��-@2j�8�5�7(�UL^�g���8?3�d�z/Ҧ��H� &t1^���΢��R?���s<�wz�u���g<�a�.ʙ���HO��9Fm��O��֏�ȱ��oa��u�CQ�T{	�'o`�O7���9�[Bn(�6��b΀)V��5JF9�,)�I*�86My��M�h����6,�Av�qx�Ap�-��+ƏR�P<	�ł,+���d�Q�G[��M�i��=,���t"���qs��|F'���!�y�d&Z�B3TD����4�&���4,˶�o�]�2oh" n1&�����Ni�m��_hI���o���A�,�0y'�SoڂX{]��;<kkd�L�j���wR���:�"���٥���:�����6۹��g�����e6��fiKx�M�^��j�c�,]�*���9p����Vz(ϕOLm2�o�S�� v�/򩪋@?�<S8�l#�����E�'4_0�Ԣ���s�B�YȊ'/��4(Ώ%qn����\N�c�S~���b������ވ�W��`�	�p^欹ƕ��<�|����ߙz�ZV#�~J��c<�2Fȩǔ���4H�θ���V�y��`p��H.w@�!���0G?-�x��-�`�^'r����P�]S��~b$��l�����ofD�T+�	ݟ��O����2k�J��A����{Ō�m`�ZGF��&ss�3�k�G�Tpp	2H�h�=��K;�N�,�ԕ'��&:ٖe.�� ���l�����D)R���[�0�/�4fYG��:^,��`�����rq^ډy�\�xv�o�j6*'I�D�z�7:���H�͸Ld�腻É�=�&��Nz�u�I���@��}�ԭ�K�p�&��(
���H�W��ǡ68J1
Ҫ4}J��q���`>���n��r8������[C:�(����q\D�*����'��J��4��c�r���?��{����� *¤M�Z;��)��*WX0��z������Z�>9r��T�=�Q�g�t(�=����7���hP|-�����+�ת��I�Q�)j���_�����Υa��r 91��M5�p��I�b� �W�a�y�9���{K*~JN*m��n/ƪ�R���h�}�bbM�����:i�\�u��t���{js#9~�G�MRu:�b��o�
��I��|Y��R[�-̌y[y�Vv�ٲmh�����Yd����n�J�\{2Mqs�����G����!N0�!�V��Ʌ%`f��k��8fq��P��鹛�0�Mۅ?�~��@ >�lx^��4ԥ���`���D��t��~+��v���6���[��||�f��`@�̷� �>�_@��D�m��h�d�_��[Y���g��v�\m>>.�HSі�af>��Bb���#��+���M���Rg_��l��7� _��čP�H��#� qA��Z�Z��&����bS�b&
!ѯ.pٿp{�ʡ�������%P�,��s�sQ�y��١��(~�-\tʊD�E�J�5�s�?��!��*�Ob�CJ�EF�]3���f�L���t��W���m�%��}.D�>n7���5��&�����,�_K�;��K����NCQ�?��i4br�!�O�.ɒ�ΤV����@T�h	-�9�ꚢ"nY�a�&��h6U�<x/ѱ�y~���&��,�X��hn�w��3�Ɠ��7C`]EZM���P?x��/�9?�D�8Y�A�<��@�5��xV��)QJ[@:��@�O��&m2~[���M(�`B�}�	���2�oe~�#��ܨV �ˬi��L �$/��~k>e3�9#�SzBm�@G]ힼ���>C�F��E��Ol��gkdB�(9	Ymn�N-*1�61��z���0;MNd��D|�̵>��5p(��Ԯ��w�x�v��֛:����P�.�M�փ�Q�n��
K���S�0��{�6��Dm} �e��gBr�3f�`���U�G�1WdI�p�b$�wt@��c��?S^"��A�Z��*�}f_��j�w���]�/X�]X��Tdl�bEϊ�Ĭr$N�E��]�'�G��]�ԶK��B��H���4H��Ie��I�.�>[��8W���m�ɒi���
@^���qg�T����Id9�{�24.��q� ܌������H��������s�2��~`�Yxp�a�c80U�͌H��t^g�;[^2���������%m�#V��$gO�O�h����z0��(WƵ���C0c�#TA�[��%঍���D�}uf\S�}O���_w�^d�t��_R�u?�N�B��f�Њa�o��l}�$���d㗚��;��q ���<	U-��軴�7��n�c<{y����iAH�D����s/��W��8���*��3�r�G�l"旯��W��ڴ(+�$��F4����C����G�ڟVf]�Md�Y^.Տ�Rm��>}`�/Y�_.�/�we��(ן8H�&��!DS�{8^1��%��-<���"����c=յ=rn3l
�
��%4l��	�D�n:��[a�f�3��.n�v�!+Y7e�M���5<��/� ��.����IU�]"��xF��co�d���� �kf)+��푍P���%P��Q�7K����fjqd�����0�r��1@�*������t8��UO�o�i�f�˞���`g�����8ڞn=|ʯ�:�N��be����P^��c5cB�q��~E?�:/e�-�夥�	(��v��p�UDBš0�ޯ�{��ytΣ;H��˯ֿ+�=�YqԄm�6I��,@���{V� �3�\���/0Il ݨ���dPE�M!�YZ�c����"�Q,��������E��n��`8�V��ƹ���*\O_��ip�����H ���i���˘r�������ڡ"���������Ê/�_Xȃ�é�ah?b���w����d-;��i������Xz�36N�5r @�P�M,�� �h�ȿ��ql�~�K��H���C;�E�Len�XV]���T����.(��'cQ]��*�َ��oN3�X���*�p�*ϐ��b@{�6=xW-o5kɤÄ��h�P<U+��\񾣳(�֭ؠ�6*9B���.�����=�J'�w@Ѷ�G�ɔ)��(�%��2eP�c������=�|�� w2��hXXh��ds=7'v��\!p&m�u���K�/i)'@�)�x-T���~���z��	m �5Ac��}X>��������5� "�{�W�0N2ū[<�-hgjڥ�I��K>*�Q�Q��}$��v\�o5�&�˟�M/v����eP]0�FJ^=���!�=�ALٞdUg�r
��\����u�5�>A�:��Wl�(d4���
Ԯ���Ej8ˁ����� ����5&�]\G�c��(ƃf�RXz��d?6��Encv�,aV�;�#�[<�R#Ԛ� ��jX�ts�a�8�!z66�Z/`3�"��5u8ߓ��l$��10�x靃����?���6ND�c��Q�r
W
�ŬF�h-g	�t'���KM\�N�̧�£�M��o�)��=v����H�
�K�Lur�5�S 
�=�p�,U��	�<!��3m($[�\!�l�����Щ�����H8��aP�VY�%�ewz!�\�;t>D��W�U����RF��~��;V ,�x`�؎��.�i�E�C4�ݯ腾q�K�%��4�)=�3�ž��?lXB�B�E$N��w����#x�|��39�+��uo��.��� �,�R�X8��PJF��h=蘐��K�]���J�"8;Q���@�����B�3��ZH-��Vk=gOAs7�g�!�_Fx[-gAE�i�.c��ݲ����`tE��l��-��yEby�[ob�F�\m_Z�A��w��J��Ȋ�,��K�h�b$?/D�&^�Ug1(�O����s;�-����ʚЧT��9a"ɳ"�Ŋ2Ur�2��7Zؤ3B��7�?u�� ��9é�8�w��Bw�+�}6\h4��nF�����*�c�ک&���M� e+F�g�Eb��'�Y��؎0���Oq��h��U��Fy	LoX0U�|�
�YRy1�;����ѹm��C�^@u��C�5Y�c��������-�m#I	��]{�[�T�3̸�q����!>$����V����d&>�-����VI����)R*3~(�s�����_k��2O�X��k�|��!����d$��C.���-ʒ��TQ5��`�����3��U���7q��ߡ��"���L��w������IlYtt�M��Ny�ar�4�i��}S&�ЩW�S�S�������`W�I����� ��|��=���q���G��U��`�H��݉��������a�%�a�~
���r�$s�;�����<�,��?�N4�aH��}W39�:ێ)>̴d�6��������ڀ�Ȓ�FY���J.�o4�jiGs�0i���SGA�k@�p���2i���{�sݘ3���K���7�
����7�[A�$7�[T�E���}�_vq�UÅH��[��Hgft|:��<�`L�t��0u	����ZoE~L�2f�+6|1�ŉ�N2_a��y�5�s�B)�Q���t���$��{({Z̀U��{�D���`,	��FG�&q	�dd�Tg�1k� p{`� =
^�"��?���q��oH*��ʸ����=�9�f��6>X����:��Ƣ���%R�*�\6�e�h�k|�l{���3�kj��~Nc�;��������멐DM��x��WO�]��I|�!xj��0	넏���*̱�A_��Zw�9��N�y������L���I�,��B�ƥ�EI�qr���kw�Zn��ִ�׌��0�HNr�d��y�����F��j��Ig/�;S�w�#���Z��Ita��~��(���\�|R����%1��&~�r��~�Xb�o�m���4�bg���%�^�3g��	��Rf�(W�6��,��Ef����-`�:ќ����r��m̵��*`l��Es��p�,~����ra�Ӳ��ȯ8e��#0�y�F�E�`G�r�j�A$��/ �ި3c&�)$m�>������2�Di*&|�¼<��b4+R���ѩ&�f1�R ~D�'I �_'���|C��	�<0�����$g&�"�A� ���Q�r��6+��!lK ���-���ʌϠ��_�2R��/9�k&���4#7��ڞX99-�D$�M�.#E��i,�=���m-�dZ4��_��L4]v�h�5#�EeJ��*d�i}^�4Rx���d'S<TV/M��I���Ķx�/L�yx����!9�b�8[ei`��U�D<�h�.�T�$�d��K��e���i��!z��0/�:��*��r��'E��Μ��O��E�fd�,c�d!ĭ�֕9�ב$z��L�Z&��VB*�^�>��)@�EX�vo���*���?G�u�=��Tu�Ԇ=L������@��_��LU1��9y E�����0ImD��B�����t����46�v"�E/f	Gq�9J���7�I祤b��`�M���"M�2l4���>�����Ss*�X]G!ww���������:�A��uXaޑo�����]x��C%�HR��eUvR�E .�j�wŽ|`�ǋ��ˌ~��+��|�O�5�?)Ï�	IgB���QoW����Y9�A�c^swKT��y�7 DI��֬B�D^��U껏�,E`�:��e�WJ�O��`&bv^m"g��5��5OF��*S�����1E�ZY.ם�b(>����E��~N������g!q��r�Uj8U�i#��Q)��ߜ��xT��c�����	����l�m|Ҙ�����bNv�+X17(��!�F�
O�L>cT��3�+����D)+��G,����	/������
\C�2���c�(.�1ǭ�@MEE &pw/z�r<��>P4b�D��(����q,�i��v�"	K�f%��b��*Ï?f�IP���٢�EԋEn?�GX1�pA�@���n�����
֮5�$�ZJD�{R��=�����!��~����6��2�	�l�n�n�xE���t=A�;]w�2�H�!l��F93ڙ�����;�DK ���ߜA�>�22ȗң6�|�l�mo�U%�Т�,a�K�1�@k+
JN�tۗ;���� ����6h])3"硠2� �	%��+� �0�28^�#�
��0CN��<0˨o�e�E<�����;�E��f�Ǭ5�!O�1����V�Û)
ӵ���Og]�Q�ⴥ[uܿ�\������y���J����s��S|��φ�����d�e4}�Oэ���\�ܛqʠ�N���AJ#��M��NK�&��_F�B������,{q[�!([�<
*�D�1D�� Dg��(��E��ee*��e������^��s5�$�0�s�rr����b��]I֞ ���T-��/�d�@�aW��m�P�6Dud �1���Q�Ė�Ygw�.j�W~�2�2�1DD8���6���F_r�_�I��� <di[�6wy�l�G� ���������z�cJ@ 4Px'Kl4��FV��c�����U�m�k�~0����tZ���+�ʼŹ*Qf�^K��A�k�@J:�_na԰ez�ѴU��up�$�c��Р�8YG�x���@b�dg5n@+�/E+�&�M������o������7Rֶ�7"�sE�u!V���|CL%'�F�DH#���e0��7e1K�?������$wiiw���1����T$���5��]�=��LK��Q��0lneO�&�}���C@��2� ������3���7��mm��.�eH^�y����'�Ҍ�;zn@�,Ӵ����
M�C��bPk"��]�1��d%ū7J@�[��i���6o�n0 (�I�Ejf�����j�z6:n)��+jQ4vA�h&6&�������|,ٰ��Q��~/������dsȈB)m����ƅ�e�Wً����L:�r��j�e-�/U?s`T��fB��`� ���s2�Ro=b�\/8��P���6� �[ٶG;�/'R/oB�AǉN�b��q,g��]��!"9�~��}�0�V�T-<�)��[�Pw��Ƿ����I3fY�Ҡ�@����&����6���3�kO���B`���K�u�q�}�+5���#��.슊�����>�o�.{���fT�㱅��{n��CcJ������x����p`�b��+f�2}�I���^H���Ri5g��>�jDO2�YR���O���W0b���e��L4�:tvx�"���I����K15Ͱ_��S���O`�q[ݐ�����E$�7��9�Ç_��I�H��]�(�pU��C�2f �<PED���H�����o�T�qWy<���Ϭ���kV�gO��J���-Dto�>/S9����e��S�p���&5�%(Rhd�`w!^"-�ȫ�ỶD�Kf�-�p�h�Y���+��݅��+��)���2-��h�)���F���G���.�z5��6(=�R��}��6F�.借)�g��F��e��b��KY܈��Z�_�j{*ʽ߉#��d&h�M�����iI��^�8�(eC�@��Ewe|e��}p�v�x����"̆g��5�4���#�X�[0Kt_�ΎbV����1�ύ��I�?���fp-fY����]��D! �im�Ln�Z
�ڔ��Ո�%�R٠K�.2C�cR}����
]O�y˭O@�eS�ڋt)A:f���V4�J(��K�S�t��!�C���`T^v��ex	��1�6J��#濘Kn��طQ�l��I|TPrx�X����2l^E;d:�%��f���NT�U�,�[!c+�h��p`�m��gYU�����b�is���X<�e�"��=PR}���` (O���78��}5;͌��.�&��6ʌwhQ�3a��Z����퀋���H�ʛ���ڭx�Ai���E�2oI�B��ϴ�M���~'H�hEqԻW�`?
w�����3�w�
V�:��ۚѓ��Gm�hH��@�� >�`��%C��ŋ��ǘ�����?ۯ-�<KAV�Xff��<�4.�m�ǘή
W����t��]��n��#�o�p�\�#�=� ���^4un����^�O��S%:ypc=�
���x�:����XG��T �I6y{�����-#��9�������"�ci�[��n�F�������.eW��R���w�n�zYY�bc	V����t�E����l���}�)���赱ڎ@	��q�zP�:j�oz_/U�'�CɅ��^����{4��/H�8=��ʙ�s�ЕW	_�OMD�k�q��!��[^��v��|���8��',�
��;�߀a����;x�]c�����(�S4����tCSc
.�3)wxُR@�O�dC�h���B`:X�z�$ݑ�(���L-�D*�u�ulǜ��RZn<C��q��	��R�����cފ�&�>J&8�x�c�]�A֯���\s�Q���O��G�߶�	��&�>�N���4J���$g�OG���ut	噞lE[�����˺^5���X9}S���X4� 1���)"�+~��M�W)}�����E�M@�g�+�0�ڶ��릟��/9���V�u����
oў���_iBwإ�g�3�q�~&�I��O]�J��Gܵ�PCjSկ�� ��9'wWd�ɑ!�=\C�yILnq�h_,n��%��JWw�%�<7:&4ʺ��
5����d%�,@�M��}O|2���\��F��N&"�'4ެ*XN�O�TQ$#(���a�M|�t���B')Q`]����P�G�c��E[�斣q:>pܣ.������sߠ�۶؜v�(����8%^_����-aL-�s�>}�N����7h�J)���80Ѭ�(��a��4Ǻ����X����0S��k��ب�Jr��,r�D%)4���iL78�t�r�'�K2	�ܐ\��mi�	k-�u���x{��˃����+��iU���\KٹoN#�I$ (��O�̬�8}��n�ߠY����q�Y�����_����`IF�>�佺Q��#�w�8�`�3��]d�3	���+ 燕��s�� �B:�69�3W��A�*���D}G4�˄��I�m����V���jڙJy��<��6��c��^YRf�T��^4��@��o�?�w�QTc��fd��Mٰ.����f2sԈc����Vo^:�ݫEK�X��h+����u= L����Y�j͑���R}�F�R�����N�ɤ8#d�*���Ȗ
��D!i�iI�7����'�֣
�Jg��.������#���#���$���( X�CT"M{�����Q����f���
����r��b�!��#�X��x�K�A�L���2i+@7CG��2���>����԰��*p���5� gwT:�S���;$<48 �Tr�?���`���s����F��˔"�Q�>��,�[��B�y ��A�]��jY��S��P#d{KZER7�e{�&�ƫ���.�,ɍ��
�͙�^�I�RS��)���e�'1�E`%"��`����P���R�[_�@��-��9Xv��ޕ���!4��]=w���u|�+�!X��ל���>L��3o3Պ)U|�Oj��J �<�@/� U���/lǉ�_G����]���c٭X�����xQ��e�+�5�[%��6�����5�`p4�ŀ(�xYH��L9�3�FN�I}B�S��˺���v��$p;���sR�3�t���ЪH4ը��%wp;H��C��w����tb�N@:[�G(���I��"������r�.l!��"{�!������I4��յ�*��)��|^�x&�1���E,g��S�o����o�3�V�k