-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
MtjuENxjdIkDcXHGpj1+0R10MIAKFBWxULyeZTbKy9ceAJ+AsUWMVeV/IA/y0WyovMwiVmfoPywf
kt/elY93VMXuV8XLNP0TtgU9Igv6l1k8p51dpSSqMtDFsK1coQYpxX8fp1hqDLWDvU+F62KvYdfG
NIu1ohn/amW4AbkdZNmBxZoka72lM9L6CjHYm/CJVjIYwrJ6sxrPMaPSw8fTwagmDJ1t6Wa4d7GH
VDvNtLoowz94dax2ymmpqvM9bZSJQ59zZKzrO7UzA49nq3Or2CSfjyOergzUWkywIx852DH53M17
9sSM23oFBhuoap+UNWU6UhOnG3e+uhGbVWWp9g==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 18160)
`protect data_block
QyE7dUcabdXbSRyKVOxQkq3yF9Sgh9gwzKf25JLsL78JqOJirQ3Q3Bz2334XFSn/5DJ/oVrSe1PC
rtiQy3EtH1oeWr5IFh32/a4N+27Fv3ToJP0LBIsk5CNyx85c7w/wj8JhD5ZtNPhGLlkry6l/tcoB
yOwPNk/ZRc7c5hlNiPG1D2FHW6qT+PH2BcBaPQy5aGaLW9vF34s2xQjzXl0jI43lHCfZj4Dm6vS1
NkwNsP3jMv+ppaFbCePUecvaXb+RoGZoryKcRF9qUiIPTJ3fyESBoRxOZq1NxSgbgGYjExWpJvpm
7HkLuxISAKi/UlmwbzG6QjZKN3YUw0YGyevTRWZp8OOqvmMjv2v3dCAeNW5nR3sP9UkoW7aWCZTI
EvYITNBqo/AHmGam4GRUuGp8G/PuG6zczpc4DWO7iMztjXAF3BHCgsMjpHzt248cWqqwvVqmGWHj
aXTVJjjAI4XkFX2NatUBbyxyaxsDhJ0Gw0EV+nodfDn7cujRhJnkM5nOPQc0L+PPuSXnEbZezCgc
RIrGc01sa/+RJvETK1PC8sLruJqpDMLtEtP0TwXO0YO1ERzkijptVZeOu+6V4uG2mwTXBt+Ss4Ow
XuenABjhyF/WaUHp/VDUp+ic5NlE7Fpwcl/r74+2+aqJ61Ka+Nohm6wqkMSSmMYNJag+1pz5ET+2
czQjrlcodA8WzWViCLXpD6ZYW89JAEc2+NHcof9FU/1avgTMQt+4yQSkeEdJVD3kQJIzYRcKHKT4
78OnfFvPGZaOs8xngeu92mnDhVVilF6VcqizwGWIFSQGajttAfYEI9oXlexkBDTP77LSJYWXbZrd
xRJ8NtjZMwlqbJgipZmQnfPFjE9dST7hUR3qq3L4HW3OVqOVVwQduWB7b1ab4Q/H/rg2x9seif54
pzRihTqKLgaxK6LkN9igsPYFx6bcY1C8Km0CUxZhUBYdM0fet8WLwKrW6IlLLSkPQ8g/WLgrNfpF
SbxWkgBgDLvvEXLEqJgq7Cj14aX8ex6rg67UKr0wOCeEsvhie+zA3Sb0iIZrd7oZ9vEVvizsL1Oa
egXzXU1Iv1tC7U86Aar3afN3zh2xRCCP56zrZlcDG8anQ85VtFgyh2jJ7xuRb/SOQSv1ZAYB3iA2
knLz2c3LH99Gs/1Gr6BJDAP+D5TppIUlCAXkEBVMgRYTeFyJ35IbceSczccsIpAFm/9jSkI8MRUj
2o0lVbDorKmZ4Qx0pc6eXeutHXeMEHJs/hITL6keGr42ukGKcqar+UtYbmoWhb1vO0T6LxEkHzsD
Sg2lC6ZqW7PFk8OOrtJfrdp4+RRtpuaFq7JdWoelpyYFq0NDgF1ZN7Y0w2HaKCU93CyvCdxlpogb
8H8TqNAtPFxgsEFclQO6G+mAVLkBpXDu+ryf07bds1Rf3Rn+E9L+iZUCq/R6SzPpV1Q9YlzNTAgq
kF+P4f6j1vlSDt8bW/bUnrI2ifFkMLKKlDV13I6O6IqkYAFSSx+mGkCF8qKpdJx9Ia5gUEddKnX4
x9XeoXcu1RSbzJBorbN5SQ218FcrNZwkNSnHuHCMJK8K5NWXWOnvgE/vJrwM6l5tdN4gIXQUhFyn
L/A56oBkZJ5t8rzygSUjCJpOoFnQVSMzxtj3eYvenQm6XtsQ+3/DeKmzOdHBVmnsjNyCHxqbwAQO
B+4qKFwolE0KxAZbTg11ipwpsgsDnGDuxavvRfym6rU1pP5YYmXqwIc2hXbMAPnJ3ZuHklQSgAx0
gbqAgC1X5PsVk+2Tog5YtI8Oown346aHJtXMvEczbqYNTB9O2t7/NHxqabK54cvAuezZaLafJie2
U3DoVaJi1DlDUb4diVdtfLyKAdcjOd2YxgHNItvXfkf5AZScRwuwobxmScFGv1n1SI9AFxHYhcC/
oqFYa0Bu3t/FkRGef5p2sdh1K8n7KLE4nputdmTkp3109NliV9JJyDOAwbmlc85CT/D2HAeYefRH
O6x0mAeyTj+A1N2e52xEp8YnicBqNMuV6u7YM1ivJz4Z6x6FQIxfGkbUt3cJaxDtQUyyqVzx1F2r
Y+aOtlQdHwSDWXL/9v7uUJDU5d5P1PxNSCdH0KaJSRG/RJJLRomrqE5/LLnTX/KDokybehZKz4rb
uwl+EIQCoXYMHhj93S9BDcJ46rABfUr6Ue8CI9DSmHm0HBI1vmHfxsgC0g5tczX7Ycu1D2CPkm1Q
4ai4WcwPy2BlcOVYvLEZAZ+CwUKYVLPBZD+XySLXbmW6HZpl8Nof5eTdgBQFUdHhFT2O6vSS8BTh
+vwQ2V2xgS+jAb2RxrpazNiE0Za1IYExr3nKcs+JJgzbYn37FfcqTIjfOxp0GBk8ouLHooeDikl8
R3VP6VOgGqwHKOcbjPVaWO8telWlHmr8BIRvDLCXLYYYPUcRwB0HWzWgQ5m33mdXyk0gMUzUJpdS
X8pQqoIMggLtyHyHmGndtdBSx+c9mPDphTvNnCc1p/E0Z91IQvb7dotm8Jle/LmGxZc9fJEu+Ens
43i2RRBcLNbtgv34BS3voYQwknPV+WMtDLHazqTRJec+kbgvCE9FE95jk/O2fKj9hSg/F+DcnsL3
w9/gb5QSbxMa7dEs2JywYCfqwc2rUO81OIzkK6kbBrreea3kEK73uMaS7VrS+0nQyst6UVOWHeHt
OL18nG5gGX52QG69nRwT4ltuiDcflHphVSKTdx16fWQtjvpn5C+3RLtmCww5Nm6k9AFYd79Vsiwv
23niOqNOL/+fCTsfSNBZvUzZw3287SPRZhzj4qwANwtSBtJqVdTleRp37ca3JxoOHnP7GVpOx9GN
8kU14Q4n9BLvUopQrnhvHs4+1pX4A0Lq3OlnNJgTVhkBrTeJ8Zvj4BQoTOZW7b7cpgsoZIgF+4gC
8XLCVgvuFyxzWevvKnT6XEkOmxOE99wMiYaP+wM+Gv1/WWsDAoYzW0rCNYN3bpnf4iQmhL2IsFQO
73piRkzlzhA4ONciqqIjQjfigJyTMIVxcRDRCUNFjJ0a53B4WKYLZepL6Hoo81q4fpkmmFAPnaEV
brsdl4ACQEvDll/mzT61ja7+0RC/n1jZzc2N0grKJKmkchy+poTha73vCfrng83PSnZ/fQF8zMmT
Rj7onsPDHt9mlOHa7MwfwZJt1LZuXuUHDYW1ojYRtAmHF7vC6s9JMzfPIJVh7KE92ICyIgzzBHMl
65H/fcneZKQK6+cI7+s06TUBYAP2zYEQ6Ha+jKSv50rWeG+363IGiQb3dBch5OkUfkjzoOn1egEx
ShMol9+EMSwJ4rDbiFrHOHd/BNTKk+HnB0vwM1SKupbCTfGXMPe9ZKVCzkSaxoS870zWt2g1on1l
1XFd1yiz1XXSw+NePZFWb2nDEZ3dUQCotWnFMGX3SOn8bAiBlQNIxKZkI3tSSBGP70rGXyG2XUOR
3MF/hdB8x+SszG/pMyXgNH6NC73c1dy6WNm1c+q7lsRr8zd23aEcnnMIOv9I5rsV5qNbbAXPIUKe
gRpmpjKVGtYrG5jhb5FafvhE1EZRg4VCwi8ieW4tl9tMfjR8y0ncSfreFbkEMcItQPerZFDWVnMi
gSZEoxIAIW8ZnjWgYt8Aq/xjzDSfuQCTNK+o/pf6mlL1sj1G7QFDuYl/S/4ItgKtP+i0MLCsTMI+
9IivlnB4X0MV2sQ4Oo8qG8bgE9ASZ4alauwJVdCZs/eueLz7aYce/AtSvYxA6s8m7reIE5kWD3No
+o50otJSuX7HvD6w0mR39eaTH++X08+bY/d6xa3LelsW1GMJON/uaj0A3lCE+XMRX2i70aSc9Imj
4Pt9hoqI3YkooGJGPYknEfSZZxrRqvXDIbZrqliDW5+Sc8KSqBrjoO1ZJOXnsqN4/Axiwx2I/IQ6
Fbq9hrKBHCHIfixKRO0mMmjdwLF0u9Iob3lLP9RTrKF4ZDR60NQEofwKkOtU6gsOzuI1eIY1myhw
7DJdm0M6DfSSdy3OQLMFrFwW1X+FymzN88ZRphQLiOktLoxYCIv9DP2yyOgA9XLW5Y4icNZGOgYN
UXPLmc4Zn7TCV6LsmwE+6U91YtjnP1O7/Bp4+o5hEG3bl2S2N8H6EWBNACoaBMPjq3j7dyo6kF1h
C06n8ywdh3flonFq582EZjiovEjZW7Q5of9bgBiqUA7sl4lJlWdO/HoJsR27mt5qROTZGqfC0In+
J4WnXKZUk5Jg4i/PHZXnmojfQpYnpLoz/lEK9HNZl8JEKyI+taGS3BlnwNi1Q8ZttjyfkhZsIgke
ughaHLlJfKvUUMOHXXPA+Olf05xNZ0hh8AOtkLcBUHEvq8L509d2VMH2qtMlifgA6u4uER9KxPQa
ZFYDodJ9WcuxOnFtk1/5Vt2xkjrMoxH2pj+KwbaYEBBnJ0sPfNntCIWdu9onz2IExY7tbiS4ZLpK
pYIhxpMZVrzZbnh0vShqPhqXmEpsGBzUIaorRvdt+1btRk9P3Jw6g6vFuNVE5082AbeLcbP7CkGT
jDBdEk4NVKQiGdmcHTzuFOAGAKYmXzfTkNGqHo8yjylHslYoBTIumQmiN4qkFY5kSpsGZ1VMuORc
/MxgyB0i3OCRtU9DjrRhORxvlAJJmSMwUCCVKeQXheGXxSXjXeXJeukutkK8TVjbbOrjweR9BTYS
mlgA5rpNS5Oi+QFoGKE9ML/2zOoyvH4E2Bz9Lv1SPSFYMcWHy/emYZuZYTDxYlBWjeymDPjliQB/
V/OEfaOuk9h6egJUW5P5pyBC9bPvMhgNpa6mg+DLOyFyjbFOnd66bSwvBHRhDL0ufEYaEnLqCC8k
JozaDpG2GtcLUNB8sLNvkYY5By1jcaXRz35cd7X7cQKMfJpgqzGbneh+k82NQePaqrJ7Zd3ZPaGO
ALxOVlwS3mFnVj6EeGTYSzfVqstRObupXPKwUYJlg6LpgLoY0MCheBI+NZ2aqWUNWCqeMccaSggr
x/7ozfUS+TyuqZ+fyr059HdhEQ21DiopWCpVJEmWg2naUZ+BpVU+QTkJTZadI5MsEFk/+UG2QRjQ
eYDwmepluBbvSRFDax9hjYiG7gSr4JdZNJe3tFBaa5l9k2tNfK4AUropX4k2FELpIJomZdTliaSB
ZWE+f7eADeyEk0d1Cxz0NcbUWKn5WUjgrPEK2WrYWI3C5UbQgr+dftjyF3R38nnCHyFIqluTdcC7
Z2GzfJh8L7ibsKVB3ERkKl+m0tmKjaVsSuCA7EvbpQQlamYXjj2RV1Kussh0D/JwFxVIi4OtZQHD
Paifly4i8RbI5Ww29yIzekoM9hRlTJymcU3mJjhuxwMFpCw8kiTuFyEFdWqUu2JXyKBsXYDLbCYX
2COEWh9SZRBqbzM3EiPpv+NcxNarZjO/dggfTP6uzauFycJwC1BCQZh4ZVAohOzaFx4bHHaX6iK4
B9mDIWYhSatmryMQSqbbd1ANU21uDwQXicSmZwhGmbQ7H86S0PNg/u99R23oH1gdYQLrlOkO7efu
4lPy1FRZFXCy4H9VkpLrOdpJ8a9O4Uy1hPjC8HMRFWv11gH2D4vUQ0Txy2P+YFvaDqIwHGG0zZOI
NEe5vPNUsH6P6MNe22bHOaFr5H4wBsx4n8LrN/afX0V4B5rQ3dCyEI6pe99baDjFxIrUtTcvZWgY
foaTiWy53RFQaCeabh1q03EhVEjU7qCn2YqYYIdrpOULu9A3raNPGG4lvUCKbh8HUUwLRQEP1NLn
EQ6iFdi17andvtJBay3/pxtMsRNW5tW0Jw0LKx3h+Yh5fesz8u7K24puLzoG6ENdw+Dp7VI3ON7y
X7OlHdEG9ucjdT7E6I8I1T4UNuS9nYCnyeisnutWFRwfqkNywS+luF5Szpb1DA/MzKL40m8FbK3y
EwXEEH2DfMNIBw/iDlo7bl43IhjtD4dk5lRV7A2hu8RDlGjC1lxYPiLyM6Z69J5GHhxRsK1pvanu
jGEFAePR3e5rhFTkBsqhmI4OWv+xl1kb77cDSaJ7PXWPDTFGw3BSEKcw4JxBlzF4nXLesq37npjt
Wi14fEMlwP9BqMKZnEzQG2jvOHGqMXjgYC71msUBA7g2tlCLLFC/fbwf81tW/gid4t9DaEOK33zw
GL9Bplkt4L/JLHgWrsK0HDXrMXRthR2iysrpLYQk9uL4/7InmIDCVixMc+MyUiNvbDCOAU9K90Rr
lFYUr03p56M5YYoNe0baf4q5rKoEsUO2sLGSvG8v8bxLhmAMz3wMqvQvqepJQdjKSV4fzbJrb1WN
eBBCPWHoRPLagW975mbgqq1KMBpFYqSG4IQMnV1pMPkBKQGrNQEj/+r1D0o7E1t6WDKouov5JQSs
GXIyfqNHRgV3JsG3OA0qr2mZAzcSrmhIj82Q9rBb6nsQMbK6XUgsJ8HN8gaweAf4nR9CHsdBCD/l
5y/PftXK6TKFKu87nwKe56JKbX9ejiwnM0Hi9I4qMnKbDuHCofH2PEAePCRePUc+q6iawO1+NtfN
POIp+NApeut03C4ZAMUOA0tuuHA6SisbQ0mGH6+DuJQeRz9qBZzdq5fDvztqNoHSaZDaKqlUHMBX
/SJ1/B1FjfDUvlmnF5N3J4w8fX+OGE6ppc1hD19JoeIgbbXWmy2eHsbeW3NnCEsnv5FwuWNydmXq
9mJNTdaVeSLE6AoTAINIUP7yY+yLhzDvh2vNFyg+bT0ThednSh33ozO2EXDgA+bCJdbagKSXBalC
O+eLF+hdQv7CXMIBKeNhF5auJk4KqhEtk3yrbQDGy3ZoYxBLuJ1/Aab/0W7zipSsj20+zQtXx4rT
fiWYp15VjV+hLxnYjWBUYx03/cN99ojbaNlVVvyXo/HGacc2RPpT/IKIfR9U/BgWiyUqXOb86dup
tdTQm3gRvlJCvl2F6eVy+bu6/09FgGQtRomVq2LFVGeYprwT/hb/RnY10uGhYFIoj8aidVLobpsV
oe5y+ATvk/VcnQ4hIKnUDQdmpXYwcc/nltQcvsfsefSI5oi85ddpyymEN2NG3loj5wzp8Js6GatY
ppKrcEHB8RdYIW5FLhFLxdDDk0Tua1ljygbZkCiUTHksm61M5EIsIKKZHhZY3kh6PJBk6xqQBpXj
tkRAI5uhT6kv/Nq32xqFDjBiufC7jalLRbHgJWLnX/csogx1oJ+5hj/cWJywIBoIax/MT0FUz5kN
ZR0hu7fqZKi27UENAgsoDiZAa6wF8dyFfww0V1M2aX/cyp0o2/Sd0+IW0D8EdoUpwhk12V2FQUHd
7Ug5cKB18zOFeUojM+mPifU+jVEr/hDJsXelqu+EMDHnWII/MlKGAiBMvHPBbj9gxHZS6AZ1dQDO
z638Gsk+RcKWxSiJj0p8R2JTxaxYSlSh8XaKVV6ACUO2QCPgoNGVJuYCm6KrtACsE8BYPhE8Tv/C
0acLaOJdo93It5i3n3MTdZgWl3gbiDLbvHJEBavzlPMD3zXZIDYZQYJ3PKvHa4bGQ38t9umeI5X3
1E4R2DzRJCUCizVGcndJHbQdj0DSbW79uYz+FNXCV8J0/pxFjjWKqEkPL+1WKkWYAd9iQMofGCi3
wBXEvF/PN7NqP5YrCClEqlISGTw/bL0Njp13YkZ3iHldKb1czM0r1oJtafo7UpsGw5vrEioFdV2X
UtSq48NUUinh0y+Xt4SK+98ozw+Ps8KAAylkGw6/WJxhFUtWSt3TMOWPG+0DWMSmKBVD2rcQfjlJ
aeOiaOK2aJh1WIOC/5S2Vy7AwwSGMwWcVwDxT5C0lcqA7kogYSyBeYbU3mrnO+V90rPttNq9W9vG
BTLmHp+t+yMvjvIr8e6JC241cg9aLnOP89nEWL5KOxSichADSbJHPT0hu8fAqfAR1u/5I01MJeIf
I93cMxCH+NbLtHRnW94ib9U/0igCWrlA9cVD9XSAgvsN8lnYO5CtveCgkheMzQp+4WIbcw8gh9iV
sZfL6SKgn0tOUdPWd7xHDqaG2s/lADeIdXHfcgsfgVFAXrLmqwWgb03MWlgxozwdHlWbk8G1r6M1
eM4TtKl5VoBl8gXHebVsQeBp+0jnKsoiy7ojH3anhUJT0pkAYaZBNlfAMiHEiCt7zGwWpn0AOER2
7ODDPut8tpc+jIJ7Fr5Ujf7d55rOA2DNIDt+NacbAbmru+UNEInb+ysI/MR3cA/q73CkQ4PpB+/w
ueoU0Op2PkPgyCMK0Dwp0xG5ldeKrXrnJcn26uT1Qj8/WXNFrCXBWc8FgSadt1tNbPHoHtCuuQxn
QhdETWDs+BRaM084ixK55o2+0RgLV73EofiFmJAngR51ew/CGU7GFh/tsz5ey8FDejncX540SEbF
j3iqZix4xeGPhECp1G4orHdg5xSt7nypVuyPRf4a8ykf55iyp+OD2Qp+E5iUaL8MTp85lUyoO4hC
y+ZrQn+uprL0GicyRVc/pPzavvYxoVntjPbpJqk9WsRUCtrn7DVwoLWqSzx8D1bxpjDfhxQIoxHC
vvoVqwNUfVS21r5oCq0XugZhsLojmNKP7vXxZ5t3b7kEry2Qanugjap8vVLNLOJczGNmMG6asR0o
RAceCjUUy+mNcP3JSA0Vz/dtEO/6eQYmU0QEYZWMAQzr9PEyHjGX8mH0I5JySkmFx0Jms/7N03Vv
C4ZEgSXRTLbMyOdRKyFR/3NyRi1D9UHf0bOwklLNRzmKzT6TznM+nT6j6lC/KXZIpwciANOPYL+C
QcjSOMrAG0OVmngIPJr8r/dT2mmVV515aSHgKxRZxuXRuzSg9tiL8aaaA6iwviSzEg5ZJuXfzHma
jnpPwYlQHSWVX1soTwxbGNOKuVhhFKlkFsRj9o753otK+lBaahomlYN5KbKTfBT0izuLi24tcJqg
UA/9rHioU7OMsFUmbZsP51k6fSeh5HGZ+Jw649m5os56vH9Lhef7jg5FH/SQrt7T0RDC/OSC2rmP
oQm/8SCxOZlY3n0LeDNw3p6pGUd7/Ev1Fg8E1xqWK/D5UhTobKheY00nDaKpT6GKOrhSpUhxFsSU
GWOBa7wUZEr0kFQhFDV3AZ8LyguHPOJzTY2sdcguOE2bv+FhjglINW3EjC/7PPPIXOAk9v9bo0ob
c7/YA0l75/rDpnduRJGRq6xvozMGzAwTeWdnnGp90AF2f9pK32IXk5OLR6gPUoWdKn7QyVTBWTqN
mBkaxVlLEKFIgcsfjo9CPuEOio0iPhVbYykAykxhPzeN2qjhQSiDW+KbVWLSblbYyr3OoWsK9A/U
MMlTYcEZuxUsthTMWMyscXUJRNR8dTZpfIY0Dcvm4agIdaq3QVozzU/MR1w+/wBfEOx+Mi+xVqkN
vkk/46e7i1h2ZBiXo+fEq/Pu5A5kf8LHoL7eNDCR1qegiVE1OFxi0/YvMsyoASf8E7gWWwy1SU2e
yDh7bj8SvzhLoNmOe9wamHX+yZH6EYKEL/pw3PGYVaOt2Af1Mg40mXOFZkkwUtHW0HA2EAGPm5Nv
7urEOdb8gTAkeec9cJbjqRE+nxi3Dwipz/l6fit55YpgNw7I+bGsrT0WMrzirl9lo+xmIouGBkyK
ehQT2/49bVES5ey64ANLlEKks0r7bo9/fGp1Yz7Y6NBBptgJfX8Pezxo5hzZ9tI/BlU1ssKcbTcd
WWTlyWE/StGTMe70b4Nim0QTWKzJTVdx/oKPJmDIDdoSpsd5w6n2DIqyfPi4w6mD+taz18LIhqzD
cjCeB0ZlBCofYLp5TxJBrPYiAHso6fl9LMYlfK2xP7sbnfS1b0rh52SYxzURP/aYl+HVhZia9lhS
jFU2V2NCUx94kjVPPbnAGsVjN3CaPCbNSukNcjxNjsInzDPSTO3ZnGp6SQjA9w/Jjj/4wHQ2FppL
+f81uO4TVZaB56u+qCvV2m8d3HvJlnG/gYJMCa1D+aP89G4eVOTfUijIhZDyfrYuXGsNybPaksOz
BbEDD6F83k5jWKKegqYbvTIo+DEQX9UVkaK8lX6mtrcKdA5PbljuizUt//ty39p4g09ek7mj+ukd
a5+EtKV3gPCRZlvnw1cG7T8D5VZ7BDci9ROOnCXXOIdDOt7bSAg+Azdh/8FsVuBFJnp42S1K5RAM
EO9g+Yt8rMS9404YM/RPxH77s/sKoEAJffnKXl9K0tVb0i+UJ5bXn42rQ/ZzzpJRVsvIpL6NoNKN
jsgjyjvdW0D7a7nhJCqxqjsou+PdsGm522AebtvJoV2wew2Eu1pJU6eBEKTP6Mx7HbzawcNVpR1J
IHJOZBA8SzxgBBVnR6F56FUrRA+xGPbvmn1vM/9LIFuDSZ0iDXV0ycaiz2HsLGRgCyCcjr5Q5igj
M+dbkUIs4A2Z1nuGixKQK+qf3s7FhoC2LPW39RDet8ZCZU/o0TeehXmUkX0cVXbb+0+Kg7al135J
kkAf/QNNGYnCJhz32hjMaJvC166pP8lgTAAKciNmHY0kKAcyEoU2hBwRlaDHTB/aw8lraxk1b7WQ
MpAA6NnHYgrYuwBXEEIDy2pZR35t+nxoV9BeQkBGYa9Nd9Z6v0quRcKNsMy+Vv35MegFn6LXT9Tm
p5NOs4AYH07tQSa9+5//jvIgoGBD5RmLQ/xw3sI68IRRusYX7y7YzXXkdYODwHjZKCGESbFyIcVC
8xIY8/Wdnwj/NN74kOR6YPgwFUEThBq556IBl+Sj7GJHuD4gZybQ9sbgFJh96ypCS3uMy4rhnVTl
06GKFy/OfAHNRka3v5a9hgh8OKA1R4V0yoysA9f68I1OVWEWI6/iyGP00XomDv5r3Szr5UffbMSA
aWPicchc8GkBsgNyyOWT9JC9UzwAPfnxMXzIYxjnUh3OTCh+uwJBmYfR4KivV6Ci92/JTeXX+6aF
5ItDzf2MQ+Wwq33DL322nQgr8RZhcl2wrgh55nVisN/EUlGsEWxjwlATr5tWSpmgAwSHGY521y58
9sKYOqdu4+5PbvFgxFJ6+bviqnYYbvpF2JVVur5V4NZ9HEsF0EyP+Ga0ydETJjBKbRq7/BWwfIhX
Au+q1lg5qL5xCfkLwY7+6v//3KrAGuuyAt60jovTlrwsGXe3pOE+LZG8t2vgbpLfne4pqj+1OJC2
vDvkYOqV/URoRVQX9blimPlVVh2qHjTuzYBc/y3nzZzDxneh+oX+dVpZg6Ige8cylF1Fr59aY4lV
hdxGCep8Ix2IfDexZSMgjncMgyJ9hNiVInWY17LNKVdYH2WGqSgc9gw9ChGMAPeLlRIjPiQ1rlKP
pU/NOMo2q8rhh+97VerhIM1Ejl/ocEoiY7UqLTwHr5Fnn9KXNxiu0sngUyQ393QpWo64pv2nDUiI
/+uBxb7yQmyPRXcqnSAgPDrjHOQejMk4g5WXSsGbgSvOhBT7nSADwEZX3DcA/v9uaTwtx/wy6bJs
HTRhQQKhdo5LaIA2aF2n/FBOLFxPqG2EK7F5kwhZC4R1M49LZtijRwcD+3iMYlinqsT25mLldrU8
pqoQRijii17b9cTw59d+WTELm8W4MPUksISrk5KLtraYa+3pekHH7hN1u/lAnBToHEUwjwVHUXjT
d5g9C42umhHJQtdUJbMHqx2bWk/Tl3Hq0+HlASw7ozKnT44qPMnTyxHT+3fUg14WsK8lQIRvOTtL
3+zZjaeOM5DTdxuw0YE5UFq9m2HGO2GNNI1qmGgdhPWb2hOliFdRGW4B42RNPionW2Ad/TUEBWUH
isS0rr+7EE54xdcOOj+tFIJOuiVM1GDaoASmLmXOuPWDQ3XNWa/WfjLPSTOvlK/tN73yt7+x64Dr
rbOMMmkUUQ/pFLZqQYiHndTx3A/uzDiY7WIT0EQ3sPqKtc7e0CC0FPTFmOh6hrpKk1A/kJzTC/qP
gOnDzvtGZCjhQDgRpvRIECbaChthCDy/XtspeNmOqWqYDtTiAh5gpQn2EttX/8uao5pgxf5KYS1y
gjDdazM+dPwM0ZDKnvvDB2r3QkiMVQXqrdehnU8uOd2u8/ZT9xj4X99B64mjOd5gfGuTqgueZWjA
2MiPoZGEb3E4tIAsVh1WvmAwoBv3B51uBiBer4sLlZAvzwyWngJ/UJG9LoswFC/Db1YnNOFwyp3D
k7jHh0zKWnXfYNpnoUDLg1U23vVD+a2lvUNZVkF5o9Cid2vVK3Q4FRdE0YUxtvP3cxor3T7tlNhi
JGu0zwGgVNZ5PgqsLTlhSbl2DWnE1181MOq/YDVcGUXINoePw9SbnsqP57zTCmpoH7hce/CEvymZ
NN4GzeO0WiK40eIZ92XRtdZIjpjpg2332U9LwvMdDYIttV5pFzXHk+h6W8/tutGBGP67baNgNHAo
G5D80PzBW7Sx2sJk7W9NtqSk/PTPaacVEiyZ/3n1RrFMr4HlMlze3lIDIb7U3xQC1oKYPv0v35Y6
P41LCyomuff3nIHl6cHs69Igslq3azDYQd5vm8guI+2YycSC3I5St2HvJ/Oeb4th7olWHKf0HCvW
kiX/h0LS5DBuvaj/6si2+xAJ96OAbPzoOeueEq949P/EKpOV5ResYyiJSaWwIMof8+lvk8ix2Q54
f0QSIu8ISSR9nhdww+lNB6VpUFNsVS/N1p924ZhMD1VItqK5rkKAiEnrus1aN/P9h/1rayDW/YRO
mrabnxPq7PvB7rfC9M20wpisumrqUPuhPPv1V2F4YO0PN8tvppJrdWz5NlEO0eFqZZw7dqBpZioD
Trbbp0Lc1fb9ar310e0cHTD1bKWuVMIY9mv6w09OGIBR8IZRf6zBsgT6ZDBOSeFtE5c7HGhN6fSH
AvRzcFYXZZyMVxmBYdyX4nqByOlXhCuRiW10eSYFB2s8oT9z1JJiBbUTaAow3Js2mQY6UP+QMKmh
SgepWXQd7LS+uf2RXITjtzp+mW2O7lzpdsXRFwTrrnTgg5CBBUIvVu8MYj4zu9Zxf3EwTXME6OoN
dfykEMtvMNtfMGiE479qGl+O/lYv1RVJqZhqIK9SecgiqG7Z/sBmlEzORKfJDWJ810rs65JhZ5Tu
0peFChMHpouMkx+mpM/nFsduiCFyvmsZ4tjiZn1349hryiNNa38GWJsUOJNI8W52tLdplyg7aepM
7FqJt/RN/Vrkf4uf2Unr3LO4BWCBjQwkt4BCn/RQiYrFf3ZUHftOlWfuicZF+mglWDiZmS+hRoP0
MsFLs+sXnXF0wNS9wLV+e4lVuHTZmObzyVA/0Ufbuzqpi+040Ie4LuM4GzdotNlVu0N+HIZDooEa
QC+ZN7zPuOJa4Ke63n9Y+xNWtt3+SPgIbdFDOgHkHguxsgg/OxVxkfmJZFNOK7fmbz4CQugR7JgG
VOEo1OPtQRx4moaaATHyD54OklQbIR4RPtNoNrSW7/hWeMhrmLd3TYs7E7lj3DOprU4hmRKv6kzi
635VXWZ+1HQSPP7EYfsPTIt9oSY3E74GdNh+3qAN/8vEg81bEu65TkUojloP62OP55SlobYk+lTC
IJigdnF5abUbAWe/OdEZyJqS+bKkFpxxzmQ/hJwRyn+cO8N0AGTKjEVgXgoxC3yBzeqmhqcLbbeN
N1+rWRFo9HTASobJXdm50KLAVUlSmm54ZdgsZjZM+e8lXcCE1Q4qcD90YnC1Pkr1MKcEKEvjK+km
JayrXf5JdOo1QZJMkfu9EgX2Z+pRWS11hkZTOnUWkmfpZMIChW8NK0hgtVwJcR7f0LaH1ECliiIF
wWxmv/KEAGuGEJ93JXi6PKaWHQPxOiqSPjoJhWspYUq9lw214kvTwH4G0QtMc1pyvFGVh/6wMIX3
Kwhm7/NqONl0y8SwQ8+8mGNVlHfi2DGs58K/i56uD9cIO6izyxkFPVSboDKaR0UgHq0Mh3cL2G9N
La87xTIhMnA4D7s0VUnFbwO15pPh2zMNNKUlzeGbar4qT96yxayg7P8W6aRpLWNL3P3SFdMpxJC8
l4JGFY2NfumLRJWuRkVPFAwiLI47g/iP5zZnkNEnmZrr/uqj2QS1K9a92S7eoq0FsHvqReddwLWm
0bWW/L9WFndkjVVV/S0HVqG5t2a5Wddl7Zh7lSddPcp0C93G7sfyQlJnZChCZC9ZLA7u8aK5ljmK
6a4GPlzkBzP2RmNc7kJ4UcyBM58N8jfFiF0VB2Yc+f0RuxsMDkaQ32eUJr2T1yVA/3cHdRqp7Ynj
M1WXErO3yitwqo/r9G+VLu32AomU9w1cnkkbLMZiqEKJ8HJFJMM9OVD+5h4QIChzeXU9zQuGV1/C
YR5dowefjElDxuhrsQM5RB6a2Ykx4gjj9kVSqipT4xslwo0TdcH0yTU6oro98jKQBDcDnbTIEIMq
pK3KdTEchPIJ5q5bhlJrOxX+EJKuhT++kn8e7kn4I9xVvip6qxMs6dOYdH97xLOuz7+ywUGcKxSb
TsxZoAvwCNXO0XPKMbE1LD9GHU58pk8uWi06U3Z9t7G2BFvVuTKR3NEZ3r9xkYOsAW4mmvUkvdSs
V2OZ/71RLW7/vxjrI+FEfxv26AqPmZJFx9q7wJdnPU3NiKMFkLAO+BCEAYQvZ4bTvk9D4aENb9xL
CZ87K449RiOa1kBUWGAfLzeDwoWO3o7QeAKKq9AvvsOnTKKqJrQ/oEcaGzXhu61Rrp8tXdLyrwRM
SjpiW3W7SI8ySR8oraxPyVkQWzmNtoWPm+GKixeCw0cIXKYII41P+xw0582K/v/jfXbUEKV1xu3R
jdAhv6rNUMKN1ht+qXkuWkLSxe93Mb1AwvcUkYNgPsBh94k77ulvd7v8MqKVuAwKzdcO8/Y/UAiH
/zCETpsjbpN+AJpg34Ps61EmAcKwV4IPhuMvAumeLzXPMNLa8wURwuIjUjF/Ho2tcXeqzzu3Tq38
8gQ/bxgRw4pMNwSBCFs+z0N/azcjLJ1sKDgUtiKPyHy9b9VqqQ95ealS+u28sZ05HDTXa5rE4lqy
dolq089sGNSjz23ZsPkkVcb7WTgxkFE9Oaf8Tximk6dNkR6Zs1sMSK3OjdUuNnqi98Zm9VzMhyaw
5EjJ33jEmiS4x0oExRX+odiCbobx/mwV1rvZRfIkZGv9pmwq324zIDOnTNxu6jq5CaoorOdJpXmj
7l/chLOfwOew726/l/IB0za6x7yGssipE1F9WSbrvfqRmIzFUBsCbKMbgBXneT//Ztnm+YbDm2Ma
wz3y5hnWjARxSi63bvmnEgbVxlbZ/JWejNSWbR+So/qSRylbs1SUU/u8W8Moz0tAqP01e2gggqQS
IJZ+UmnYDNIxIo62HcGff06Uff5o4a8Q+FVgCAF7Mv11CdtdxwApCQvQmo5MaAwSDe7sFYkb4BjV
vgPzJsaUcLNFlwVoi+s3BmR88muuTUb8gbvIoS/l2Ev7ILexZX5DgUeTiqxRiEWZ0j/DP14/xSH2
+La+UbBoMN3xT1yz+bFehwzqUSuiWmVG+LtthDAVOZHHUUcRu3zW+iMXsc7d43BUKujyVzU6EWIz
LIRtVdUsuta9mUNppAZSPdQPVAMo+i7N4YItdT1lK6LdEMysQVADk7XWznClFt6u91KYzOAimJBN
bn4uubrYiu8sBSszs8Nluxa+NZ/+omp90NZhEWDo30Yb8pAhmgAfaDNottpx+E3xcuOjjSc6CRvR
a36xDtLnI3V4fDKsTg4XI7ed9dwoQ42VUXM3AR/bly5geBNlzS84JbCX6w66ArY/nX7t21DVvqH9
1q0ezICFkuaGg/ZFO4nWjU84pOBSDfcQDEsFOT5I1W1UfQKgOETiST8AxaAT5SIK4w7/kKT8qrJr
abWcgV5l6pAJSybBDTNrfzaIK3XiC0LiKg6FeM+3p98rSgS8FZz5lxh0l4bxMc9mBvMnTli8HWEF
CHgGMslHCt+dQNrNMWvLWhbPDrGONPG6NKRDNmVEfMrCqyO8Soqj5hUTDLO/42TAenGceZEnW/J1
HlolH5ragknk1CCOB1kFMRPXPAMQCj9GkZ4Y0Xiu3IQ9Id9Y9FDs1Qsji5w4DjMgTsPgEM5J373b
sYX4vh+vytVk+cm4Sm907QFhbYOarpJ0FLPEpNeXTCYbe+WxbmtZko0VSTiHu9mpqcmsAF1rWf5+
qlsU1JQxLKYvNoRENcJpXiKrwicOX0qgPhGskOoVjsEhJNjJqj53I8kG/xnSiJKNZtPYGRLhoUyy
OtH1uzrDO6mU9eEsO0TDIu1Mq4nfewQBZ3oONo8p9c8jX3vKbzX8axtXGzSRVfvqq9KL3sHeE1Pl
cK4N5lkjwCMsOO1zHbEjM5MgzAoLezZAcVj2R5qTUbDXXnrQ0q55tKTXEBTxw3r+TBJtT5MwCyUK
vCQHj9Y5+ul/znJK1RwUNTzICkAD7aCyzcpJ2fAyu7wf9nalp4q84EenMeiq08TSjLesAobYg889
GUO6nrYHqXfMWt6zqHXW59ZIn8AkwMLxLL1Y3LMe+YI86YMxH3gqW+cGBAXS5V1xA1tRypNvxlOP
HwsOx0wOBXHF2WxkfSQtyZQD0sTkThQPxaM0z/jVjckgFoIiUJBXTKvyrAcIzwTx3zd/P1Cb1IRi
HpKsPgZWiN0X8+lcnKN53wHr88rRFv5Bo1hR0OYty+9r/Xy+TfPqcKezfnaAgGxFMw1XkEvAbIZq
DuScXXRA87wNtOOUv9VPC8Do/fClIXNHzedrl5zF3Sdaj31Oy8E407YziecywmNf3PY3r3anqh3n
3iLxklpcaAcGXC4HNHaQb4iIJUZiXYVMiaIh3ke328q1gqe9hsvKwx1QhVmoXmfbXKdS6HP7hhUG
nuIbbpF8+lZUWUf+hhALPfI2+siHLf2g7lbAYG7h1dHehA7uAVxAxxKdsvqsI6PSar0odchVLOWS
s8JPk0rPLKwOLk3mU14dOV09ite9Se5d9d24V7asm7J8mFzeFnWKt7aSnxCw7L6mHFWf2JPWGAyi
8myGRssSvSBzYFm5XpWpAeY1pThq+snImdcrbwRK0ky9TDt3oe3OoQ6FqqxJo/qi0fwM599nI3HN
L03Kevc15+dn1aENuc/HaKpHVn4g5jGT4xc1EWyVP7RByd/z1uyDnL0X/j+Kpl+Ap4E1Lw1R0wPn
/n+MHfsENzssYt7MkDEAVwo/ktQro9FtYAAaRzzGLsoqLS20Z9pE588OXRMPn155CNleXNW/Rtb5
IGAjjeGnVlqXYeGuvMOxlElPzA0vsRMtWAUQRbaTAbRV2lhhQU3g+oRj/UoDr/wZjDMmSSdpubhC
GT2504HImiSoru1fBm8nOZRgEDb0+woOOob0P5bb9fiFqJXwwqp+pTeX05W+gAh4jZqQV2KPAOP9
y3/5OL2vwWwx/FOeK/xb2oTAyI0GA63O5vXcC6BX8hfYlDfq1TRUBxX8OSBBFD+PwQKed8mEN8UQ
1/0/nBpqKdEcIqIYBAHj9omp4oqURXI5+fd0IvjWRqD179n2BXcZx5CmoEr09lLHj2A3+jkmHs08
BHx40SOuqLaMXJ+mhE2sH+Xmyjt4oI6WQ7hlR5+RedEbGjX88Lab41EHa32NAhEQ5QRhxm1u7TNY
YQJQfOTlRUZjPcbhuPic8xCGCVvRxhlvxPa4hVpv3Ik0fQJVQqd0kOQV2fSUJC8CHLl5eKdWhhdE
4Mx6aOh9hscY0qhh6X+lmbIMaOo3zUxjNfGrQ2/nZH7Tisfo48QLTUZv0EEa7sUAmhKDXv4NL7TR
TIP406U7yKsk3/ueIzANLaq5fr/hRIP5KORnIW+YcO1ilSI1WXNmoOmvH6cfvmVwDM9Fm4pK4jiz
EDrMj51JpsrpkWpSpgV2fExjnfLIZWmLx1tbJMy3ydEfbf/k/BNygrrgV/pZhfvQgcpEp2PBFGiu
D7C1iOOPk62t0D61FMh1k+vq10aFXKLclDJzbxqV4Rfg6wdnbdCCfdVw7r1EZGAMZIVJuq7wz1Kk
+kLrwF/XVtxtH+Cf9GyGj5E0YtaYMplpQMrm9eEUBMSRtj6T83txiV27/YD9lidOROoeEZ5UXIjT
3rLqHZ8Spw2aofUKrSqLsAAGE1ZVTnxvZ6lfxVqz+QxTtjPKbMX+W0YxQ/L7EKKdtcYmXt5S8X5B
ChsQvWC7cehT1EQMRAmJq3/JrbGuex834xJosyvBgOD5OzRy5acszYNAxSNgGHSRVCQmr92X1yP5
O/tv9dxMhXtiIVAeazsdR0XBxxkNGjU+Yf6UqaXbgZqTB8NbYgvPjn8siNiYjoLG7X7LYyDEeOKG
rjvKq+6ou0ApxOrs0mBSj9dDmFEP75JA4FTSvyxMH2VagUwA4cs6LCR0tJhDLxtz7Q0Oe3xAsnhj
3GQgxx6WWoHwg+k2bU+cTh27olrovXs5acTIVsvbJjFVzxRq+CmVhyJD026WvEzRGMuW7wQPv8Ii
XpSyMW8mreA7+6N1qeyd0yu0/+npEVQlPGkOZVoCQxj9FGpqbHD2McUQnRkoMRlW8Ja3kKdNI3jT
Z3X8tVwSRozvfr8b4vmrPJnCTRqdu4WF4P1m1NJjxNL2evb6Z8azh0oPQUPkP2kcKGPxMMqEkjOt
f6dIO8jD/YtSB8JhBfopnCm9OTG6zWVujsIBV+rkHGRop3trRrnyHLVRPbMwpX6r+8wxOsjOYGWA
MZARfSK2U57GwEIuZCqFtXqCC2tORdE+eFv60UtRAvbYiKjZpjDiSo+WjM8LituFVYzBrrVnGF/B
xHZOxVy/qj5bJ5M+xzYzgJMBdFeM/tQ+15cXfehNuiotijGQWtwsX5Ttpo7be3eac44o73U5O1QO
a+Dn0IrAwCT0o9Efo2oPMM7U8vjJ6V4CbMTJfPKX8tbXEk82WRyR3um7s8/6kNg6Oz/O9MEClneS
o4wqAxprZVz8dcS4dZ3Q/nZbfg1/z+61+stUSnsm7itggWtznMYrJQe2SC417cq+ly8AFkAMfdA9
iKnbS2fiYnijiiWSQYYNK48NpWlWFfqi19aU3pRULBMOOFxIBJqvsvkjmyHUcqgd4BDANztG5ejM
Anl8ADTmj/hOu+F8bzun7m7X2TVcAnmYJMLs9oWSUxKvyWp+D0QnzCzwM+vPMOaSu0uWB2Qsifus
fL+7T23iMbC6j1N1r8hK2Nhjr6TYWIKB/JXTWgXyQFRj6O0XrfrNz5RSR4RAv2PvkM0S6S6dcw/s
+2gq7jZoNoLan+QI+vZy0cpy+2DEmDF7yPIgFnre/UEVf1R418OVU7KuM20rt+yIONTxjsTqxGPB
ckdyNM3HjDHvMdepe4ooGibZxL4PkyT1uz3GGuFzbgyIgV2kKrx3msb/kRR0xXW/ZxO9cjIV593D
FK9q2/8/47hMJtgyrWlto5QaP6Yj2FLAglYP1+lEihRvFgH4QlgnQf8+fxCh1c+aITh9fkebIyOI
3HMRi4PEm0iWTGH3ET1L+nD86oAwNFlbBjy3ffGKW83mVCdIQWBWMuztGDWzc6qdwhaHZ5XzuzVe
LubVdLlJcniDgAkKxoyl1OinzIGbUPNoJGUbXO9iJQZozJrU5vyd4dT3LcbJbN+rbEjbjpxh4Pst
4F/u7D/QNy6H0f1DAGj4TRn0t6nh1RihlDooPgV4CcaMsxo2DSHP8jVQ+5BbMLrmEg2erag3QWuS
8tBo+cMDsW2HQz1VwRNu/VwlVCRFJLown1PClsY2TCWd3B6EInQCiZQ7Yi6z3f86nPj3UvWi6n+9
F6qXOwX+2IlayKed4xNTvFYXG/bS7qLglFmHSJ4CWR3AtUr1lD9HxyhTLVFMZvf7jAawP5alZVIK
P8d27Q36JNq+RnRjkvUYtoe84e0mg/3id694/8UdFM+Ebu5X+u1q2ZdbLIa4Stecd3H7r4IcxGC1
1aeQssbmOTw8uc9kYm7GPnLt6CwQ16xfqtdMxXvuKEIzU7NQqBVaW5WEXG88AMeFjYJAnygPxyXH
G+3ed3jhzK9bRcw2ihdYcbQYmcdY7likqPkGncHngtx4cAqJNwuuYwm5T+CSIXOAkBQWo9lgjuoV
yAeRjOx08n3N/Y9WcDK3WXC1vE7qFZWge1RTAUzn0OHlnm7p7mtKyykmLJDAunt52cA5DZf7oIO5
61NiW4v/HfGNVHbDRV8P2i6/7A9POBhKOcWuohSlD6Cfr+fUh5VDWmhD+WE+uSI8dW67gKhCuTxb
mA/4K8gSRtICataA/3IOWxUvV4E9vElKcsa0DDFxYCSaou3mVWU7EXtJ+vrlySNOe6aaQgcxiyOy
0Vzm8r6WAAEHuZ/9fab8fnYkACnlrBN6za7i3UWkSYOdHhKPAhau3ClWipmjnAplVK8woatNNPwm
jCayuXtl6KH9lua12L8irjoWyrXE2HAC/EpqyFVykR2bj8o2S7fcUqU0cu7XZgPgjzFj5GxZe16C
K6CggpLJ93vLbkGbUS8iLcggXevOh1AnuFBjwdUlJ9uAn1Sn3gSem0/Un+1sdA4uflXuRrNd4Ee6
ad0PNLTjjCWPhFtOAcrK8bZC9s7tNsnZLH1x4uJ5KUIPPK0h+9tMz5eUVYVKOs3oEyCGvLXU86Aq
zg/n+MagA7XCQtZH+ITPE8AKuf3Pz5TLQFZS0B52wECo/nEBSBl8Mwt9A5Id6xuvspNa3CXpxMY9
nnv8trMcIT08cLsnP7zMbrB5lAtuN+2zwImFm8ksMwp6oYxujmJ7JWBeNvFOa8m0CQ+jGaeSwqn2
W9Yy+QbZlqfVnv74joNMpvAZFXaQDh4PfKqUXgtyKyWXrpxEnWSpX2zgakheKr/JMRlghW7JZVBp
Kzlb/mM1A6XUVfY8NbFdYu93hG7NXjmWEYsgXE0I5hlJYl3U9JUsTbfO4Zsptgv2Tapm5KfaHQEJ
fiY3wVJ4dRo8lXMKcGhkT4HJ7LI1s29aUZDLcOiBBHOZsNyACLWKavZpu6YdBtDSIGdbHe8MAz5L
9rQHq0109xZRC7uBEvvxxnFuN/+r8BzpaOpnboUnRefs29iUj+ocdLl99FdjuhEfIVVzyB4iinmD
Fr49/jkVN6xSwu+RUP1DgD1+TZ3aKvt2IMuNU1gk4QovbAgd9/d5uslZDUJl0mPZdjn7en3ni3y9
oyJfNgoTFiXMZZnfKOTceOds8pHuPMviU+kwbweUsFhMJ4y4ggike01Ii5CR7/VmKjdtgvCS0twB
YStb62YvDTu8oodAD1FZ+vbaF5Ol4XGf8S50CjpeIFgMuFREF1mFDI0iefrj5aerv4s8vb8dAy+5
0K98QqjEpIYXOMUTS+DsYChZgvQatFPWwB94aenljif8B5Rm95uEBnxsdWSiSU+qvw2if6WcGUx8
WAonpkxZo3HyMTQnw6MsqT8vCxm+XXk1LpnhKhonC7wuiYkq/2c+Wy4qyKud4cRSrJ5zQZ8dRFcl
bbF801DuvRBfu4G0ec0bKnFlP2fG+UD7oOklJYiFUni6ulbeTBVwBcuN6nONUpM8KAvpcCNSdn2c
9wBzN3F4RVXCTGfrvJYyqV6wHJc9Fu73kkkVEIxgtRF85I3IyjL8Q9zhVuo/mU9xHoQZlCJWGoRx
jIAayZEHizlPoxHzvLg2nazAYQ5UACT+tM9fWB4PD1IgT04uX9ZMi5ogvs9+jQQaPU+/NMUO7KYd
vLFGuGJJmbBi1GiNznDUBuhcOhFMo5FhVo3b+F7PYeiRU4rnZ+O7mAKhiq0xqYUls1zO1LwM1zqo
KR53zfimRAzDWNDbZQkTCQCuOutwvDPEB3Q6M/2OLBMNmexyTlHtxX16dPukKJux9/S2rASBlEbl
FBqzhoJneAqEJYtQw0Css4C0L05q0m6JPntLWL6YJOIlFzheDmXbNJ1CEsPTuO8bYhS7iiUn5oUw
bRWLasJ/imKLocGPKg5s7PFu+WsjEzKqIhyo/d8aofM72Zrd08zeHGWrlva7nU2efFc43Pxk+Hz6
DmUCvRo4dbLqykqSjyjIuJQyWkj3tJmDWlOyvzr9zaux++/jXGbb9N62N2U1yOfjoJ45TCprQylh
lTvjzDSS94aRolMSDxyCNSlg9iOKmLS7gt7WQwDG4KeJMMGeXpH5KQnKRYjZPMsG1V8rAIVbUpjn
E4N3x3vl+5GNFhgQwKQQ3z2XZvBUgaWqLFTY5um0fBqHddBTFN2FBPHaCvdum5dGXgr26uYqJyXu
LHHo6krS3s4dentDdnQOSNl8gRBy834GzwJQTwa2eHM7Iw6i7Yy8bGvb060A53tGNCGi2FOo47Lh
AaBfI7Ls9WBsegvSCtRTQpLuWggohsfTcWQz2VN4hzMtCaaoajr1R6Cf54L8/V8uLLXJxeMAiH9v
Df+XOTJeugiU08QWt890tyIuUZ/s6JHqer/+bD5+c/TSLnjECkgD0BaVRd9ki+7Vg3jJRlTupSbR
jokPbi71G59bCHYXKcWlIloLCXOZN/ykPqvvHj13Hb3ZdjjA1j2EfeE3Yb9p4r0Sv0+Ww3ywyalM
7HXNfoPjKggdl+jNgFYK83LH19/8n/lG4d1D1onug7Y+R/zFkfderCmj0l5SbmEi8w83cp/ZMT+9
RhQL96wBJyaHyQI459GYG+6Ol8JbOUTyymH9bSs5a0lKDdbjwpEym/ogvDmz/S+3UzD7KZh1mSH+
L/bTQd+YzDPQlMVlnP2UzqQahceSabtWfsswRoL2onqnaZ3oGkJBEomKljY75uRvoc0/dZO4tbrU
6WGgUmE9wAtkVF5ae4cOJ4uXdyXzyN9h4lXGLU5KlOpFDo37RaH7ZvbtADYsAVFwSUfWaeAdyJ9m
DAP0/rb9Wis6Ek3Y/7U5d3OfuC81mKTEWdqoAjeMqyX0Me9rF6d+mab5qvFXLGrjC7wrVhldC5M7
02fHmS6igUVuoeDxITGdnF2QY+WcDiMyBw9jCpVp16FJWSnhJFGSxU3Q7Oum2tptm5pCU2+QURoF
DoFWwwYtpH4MqGX9GtwO375YblQijFas6AxKN+VaHdn2eHqYf0+Uxuz39pf/RdyGuxQzyAwtMdfL
G5tY9KNhRX7TTc4g7FxaNMQaSEhfd2tmrqBqkhfCE2SvTUWEIwRrLcwrj7pdhv+A1WSk29I8luPI
7Qx35Ie3cs3zoDAPNLgTRP9c1O9aQ1ouxPBHhEyDhHyxleVCexe14iKVcOmQhB7d9iPJM8jIwWTd
2kiegN0lvUE62cvPmLq3WFSTtdeYF5wOjf24hqaHh0ZIHWBZIx39oh/QaOxwVcEtJTxL1AhNMCk6
BDX8oAeEoS0/xA2OoPAC9uzvEy0VOmAbn29jTX658KM3NWHjzeMfCvqiYi86ls//gJY3lw+IRmea
Okh6wMc9M3vwaWPhUMhwlV82Sz1AolNkNx1bob0iesD8LCeR5igDI3oSN5Ey4KD0jcgWnqSpLZgg
2AdjoxcGlTpneve/MSHqzIb23n9b0PBcdbIzMNExh9/a84BOtkmKMZSZ6WxQ1ucDlD10rTr5EZTu
3cvN8GM6OCAjs2fZVsyLBcheqL3LY2IVHmJJm4vaflfBO4GBMs2dXWxG9pcRMQGEVJQGd2EgnHRp
rTmnhyFB47wZKrDEJmY74yBtRRyVG49LaMTr+fc+jiH4F4x5neSEhjQQZ2ABp9igGKsrpQ4d/4PJ
QXENKdYPNzxCGCNt1KAifTk9rx9AWTlFwQ5vTQ76xUwNkp0MIhAOcr0frMo2k6bIhrnJsgJmk9Ej
+Y0wgc7j4YZy2cYEckmuu87M43PkvZsuF4AdrFs5sRwIJJc2CjayQa5C0aFcAK9mQ0O/IHu61YpE
r/vyTlHOFTgIADvOxrvZZbG6WQauH9qY36hZAKioPnAhAqfj5GQBjTXhoO4KSGROHKt7Egqyblum
nTJrhoTF2r3a2Wy9JZ1d20GQbqn+tUfCYhwQYiroO0SbQEZNdSfbYMsuKa51bCcrD3wZoSi0IJXS
qpgP7x1qKf3D2g1Ft2A3p9lM5dE3G21DOdugndqvVUl9ygmUxWsDq4bugH9BNZpD3InkM8gm3nP9
lgMa+PizwPwv6Ghk/TSxWIawVe2Mx5ms1QFLpU56pmQpHwtVc35ytQAaEbZhGHC3b6siiAVN7sNT
4pmj1U/V97uQBzurIuhsQlGcmkr749rPpVgv0Qf/WEnNUWrZMqORoIfefmWxwYNAe/Q66p05LnHZ
N0Sv9PGx1CdF9ZZlm4Y3bydD9dFZ3FRHSBa6WbFTPrAVsqDhaSHiUfNjrpvDMvqXK7tY9EaLneUh
VYaJKq+RtKUB1GhL25jJoI05zzJKy0AonneOx5cA1zvMF2KXdnifb9BHVwAFHiwDlvX+px8RNJU6
uYA6ub8D/2fMKYkSMlnIXksFwhPLDhanUOMWMJQpkY0VKjrQX/RRSTxOMX1b5MnZ5j44Eg7zkLdB
f+DYXGvtH3eLDW7XCgTDgd8iPJAasCwRLCqL586MEDuKwg==
`protect end_protected
