-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Ag1nJdHvqpcZ5m7fdDbYoD41RTSOV71bNKn2pDcMbGR0OFRvs14jKA5UY7OZ/XFP50yUUmWRcamR
YKsAhBDYZqRUEJDRv0mYMO3TfHONTf75eyssGuWs7GLbHaXqM8q+gm5vxGPLVB43KXFjxmD26kbN
TIuyHYoDuW7uHw5896CIPP2vHte1YFLUFWxh0iM3JnZBQWIthmaUA6tdvi2CQw7W0BdKdKq1WMu9
X+pg6ubJmosUW+CchMg+mthTl0JHo0RUxCQ9PWD/3+Xft1O6ViJc0AEqWFZHqKCVyLa4dtfAzC5W
6uFKZRTPGrUxpPe41j63mMcc4/rirFR5WoJO2Q==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6784)
`protect data_block
k8OKyUoagvPXEzS9iYLQOZo8k9Sr2+ZgMAL166f9+EGFAe2L/8eTJc096eiH1j7f8o4c2Aj/eUoT
zmCRezhD8K19g3XofFd4Mu2FvrbjenNRI9OBpZ1hIDlKY0urdiGh7IXFVpjOPm0FHj/EntkzgNjr
1UvXtd0BU2AxzaRk3ESNpf7ijS+Eq0Ll+CHwqmUGHNxGjolmBsXVL8y4HVa3LJ4fux9yxx9tFeCD
hHpUsDYpwU+ldV1WPsAiDclMeRGymA9xlYpTk7RJurfPzgOeEfOkVCZ7C8/sVkiR8S8e+WNbekPO
8y8it3ZAhCSDQuiLCzf3qDs+LMrqJp7U/fIwyORkgoZeRKmK/EBwWJue6zvZQqVx/vcuCuTgBKqb
DuzMBsEzUijpY7TsrOClAHjWAaojAm65AxgJyExlYBAWaDIkop+GcHy1oVY4Cgh+rsT7bfx/2H2Z
Iq+D7mJDsGIKg8tgp2D2IMibeE2oy9Nm32s4cwN+DR6GsvY9QhwIJ1I2/7m6bBrNvBq73C0EUPtZ
O2XyHbYrP0851P/7YVsNERVFbGrHVNRYgiDj2f2McJc1dnXMbJxgs9GsF4//XNmy/8dP3V9zvFmt
zM63ZRyR3e/+flc4TwELsCHOR9PzQcxiwFwo9m3cNRPwKn+28L/0owtlnEAmxSIKoOhW8SOWcnzF
ClSqeJycnK5E1tOpnvu+YaKXt31V5KSAC786wTF1TjkIyiPOngaDtDu7fUEVOEsA03G96jJcqbsO
6gbr+7dfaoFW+MwYpzv6jF7ma6g36j3KvfK25hTbvYJMW0ekSYuocj+XG4PbtWNBmup4ynONC1+g
apgUQmz6me2pBRm3gO8BAwBT4J7J23eV9GkVFv2OAJb8jOWCCDovPXPBTJIIei1Xd1kQicvaGGOG
iwqjOYsIgs5damGpeWLbNViV+LbdD/oQFi71RHLMHpgvU/1JsG/+zXmVBZJL1Drp3ZH1gjcPwYG4
pAgAWV90r7BsHFVJtRnAr1eRvk7ZClWBLTDT3SN2bIe8AJ8jkSJuS/4zkNjpoXU5lATs58fmPmjV
l8mrGAkJblnglNHvnb0Ji2fCSCn76ikZtHfTkj0+W9eYii8ej0OlT7xOkhL6QQ8h7KfOePv1WbJH
pFaqzhaQPjSjQn9yUmVGrtKlp/UsgxKbC47sztT4BOORJJ9MxKTmR1qvuKtdbRN4XWsiZaHt/ndc
3avI8gxUUeTTTMtV9wDTFwJ0ilBDYz4C2cqxemTFJOA/eERADTVjkarfLtMkOsyFsnvnKnZOzi2a
i+Bq3IFHhZnOhRdUUp11lAnt7GFYUsg4BwvOuQYZkz6wtz2/fQSgruA9RC3aBzHzHyCxAyKzNq6m
cS0CjyYq9zH/Wv1xHEjz9WL0WIwHTA3oihB0ymj2R4DzaCHEWy59b9x2kUM7VnBQ4OdkKMICWPgK
2ZgXBTl2xYACQusbjJuXJz8mgelyxAp4vBGcwHmZC0q864eFMvgWBnfmshhnrSmZjG7//cBp2s3h
fvtma2X/0ijg+RXsKq265Eyes/iib3K2ctDLWFA9xhgVd/JnZ5tSAObm3QgabbtNet4gr/8p2fUT
jUoKv9TmOKiJb3rdpjkBP4fgZ4g1y5ZNbFm+pNuwHDJ6q1b1fnMRUDFr95fqs2tOKx34NROpI1fQ
t7OReDTj7t84yVmb8EWrSxNsb4uoupu9WN5uQcjQNO+5t8dSwKH6qPw4T5BnjmkXMEyoRxuCB7dh
m/FBDM2Z3bPJvZyyA7IcUEohw+x9l7JM5ZD1iR+WSV2VUI4YGy4CtUlUJhrWuUHNxsGdXZ4l+IHy
B5aR17LjmHQatj/Ey8giRB62QYdt9KhoBNKRl1JuQfX5B+WoJCIDxjNf2QJ9gXPKoNLTvWDddPGs
UrYwilkSBEEqVDh0xVfAhqLuuRb4p8o0EhHFAmMgZDD+PnJ8eym47mTi1h7f7IpzXMF9XqxE430g
oZpcpOP9fE2r07ywaK1Kd3+rdvwCUfPjwLZhgS2AaM1YqtLcoqCR2xef9XfEbhHYy1apipxr+0W6
He0JSHKYzQoDm+R7F+4xnrdbLqRM+vXUj8p/ThfcpTBOOqpoYeKNyJgN/o0Wodvsr3vp8w3ytwF7
7wEppajNco80hTqLui6v4DIhqwnrcjXHaCl7S8aRjX73vxszy46k1hhBJQZ08KE9lFmDaOQCow4q
i1QYzKiLd1vdkYnb7s4aDqZR7SWnyDmp4Nk3qb68NWnYAgf0fG1gO6+F0agFG4tl1dDZ3o+MaETL
5YPUyaE7Bgvkr/aNXum5Yzu4gKWrgNEGHaPUc83pU5kdGUdopP1Ep29wDM6xsyR3TEHFHz6ldY0G
5RH6ziZqf4bL77DHxdLR/C1TFIPUdPDU0rNikdhNVCjT5n/smNLL/2AVk04axzqehKt0qQ0vA/GQ
aeLEXiR4GmmnQzeMeVizNb67DPlj2sgd83kb6gXtoHIbWSFZLL3+uHdbjsyNePuN6BTH4opVXPiU
Ye39pC1hJwnrdiDCtKEH+CZzmSbxBTiEP5EWJv9qdnPrQSQkrGEBeFG/duSzM6u3LYHoqFimg1EE
5uw9jDEzy6XL4VxwI4k5jRCw4ClhKygZFb93VW5RgXsdPCXSwX5YFglK1sbGfqlnFxDvHkUqC+kc
+1oLuskIYIZs+n9ucY69a9JaokaEYxnwbnTzmkwlefnvTYHZ2XxSX9wOPzhySPpUWWcR9X4EZoXB
kUbh0zO0KU1A4By9Duopd5S4L8EHqyGMn5fi17BGyrJx1UQptknNNTea99DmbTH9Cu3TPT89sKxd
0R6jzsRreYskH0jMT7DDCDz/alCWq+kMH1IIGaHwyxdKWIUrCef0DqGT6pJm/f0wDkobj1jl5m4E
RAd0L0G0bza87FBu3BaZOJnLV9efDWh2Y9k8u/zEbw6ZjeyTC5cxRCV8KkakXBFlAgqrLAw8ziE6
szlcXbwTFHnHTcoGhxk3d8PZlrO7Ejg1o6Q/HfTqUA9F28K4Zbmt2bOBNMhq1W4JCvKPSgfkVEe3
zDXUn9f3y/a+gfDbMmq03l6mb6j7FC9asmyUm9SF1yvUmTLPUSzYbYlqk3Uur8kGKVvKum3UuVtN
9Ca447ug3e3gY0qURbdh+B/Gzo9934IjItHelt6MNGHdZWa4/ah0bsp8OoH7BHKYHGslhkkw3/Ef
fPV1bLTT1vnYOBW9wF2KHtVI5FvaSX3WOF4LTyw3yLhluOE1cgTKbjfwW03VDcXHWFCz6NKIuZXY
d7zTiHVQXD5iW+NAt7TY2H7MMeW+kL5qI+NisWHXVN+/1akL2S8lW7whSoUZIVNqxwpYju4X/NwL
xy8L1Fgho2T1L4eOYvZGVcmPh5MnUrS6hu/G7CeYhlEWRI9NHq5GKQ7IV9UcuUcDJdwo28eGdKdk
zWPQ7SJkZFfoy/k29hetbi6/TRswZjaokJT5ZrUpm8q3JCt+bNjUKcYehWpD80tm0kdyL2HRzMzp
rBIyayOpuBo75Lu+ZrpEIHWygOKLW63BIW0lfINIaKT+jQEY1hSZMakNA4wi/HKgIXQwGVvkidmx
udgJzUqs+LR9u5IB1ZMBx3eZe8ObM7JIATdYeX9AJ+YGn18ORIzYXZpgr1oW6J90P+jn3GigwzLW
dzQVE3yOsrVupZmcXRGJFHJHgSiqltpRAp1FXECwqiGacxLhSqaRBMQOgV1P9QcN6Ir5DOWtx2Po
8+kY+UbuCcCd6JmMiVPzb6BuzyaBmwZ85PA2oel9F/+K20E/IVmd9h/mLOBIKeQzqOrIihWWqjr7
DnyGlkfw04UY6oailMyjH/tay6Fq7Yl2gS5CPTsNWG6d9h8ezpjIYyMzqdDl1dKukZOziOu4U6bL
pbHBk8fIiZxmvSYUzFqytrx5ZMUIxLMup5zzKmhRntk5vbwvofJEqDNu1Qdq5Th2SRBBvb6etVjo
l4v0xnQ5DDi6sxCboHjYqBxaprwLFSq+wM464AwPN0KMAjUHNK3OOwRwzk+UCV6b6UIB3gBWE+74
r+ld0ohuKcejI2vwzB3XOh+NlAcuf88hfqWmNNePcyo5ZGU+Io8im/U32KsuObomEeyzls6yCXmj
nJ+jjJX5odreEpXjQRrDnK71nSrlWtBpWAY7kb4R49Zzjjef+i1mn5UkND8h81HHCcXMkRCysy83
c9H5pHrsVjFJKlV0nByxhPZncFR9l1MzqQs0LjPRdCxeAC2/AkyAESstHMZnXb/7i7A3AvQnWxw/
NbZ6Tvjfmc/1krjHJoujS4NYgeuTWduLX4i3UQnU0oauDGFHKUrwoxtWmULd7mZCPqmskmkscrnN
8Cuq+96zsJUuLAG0/pVEWtkloD2DH3zWuHigHowO2HSpdAAikPc+1NsVTmAd3RdPC6zAqaRhxeiw
/7SNcxd/nnRb3qYbMG7fZ2csLPnm3ues2BOquF3x6+Bar0zRxhCxmnl7aD55bTqxsckWaMj5mfTz
QlWpY57o1tnrkEvJXfPPpOJjkLIZjppiat/RbcAfdK2LDCmPzHatCJs8hxEAGSxGzNCoAGZfhUVQ
CB0PesU+51oC3ohNNpHfuDHpWKtBOuEC8RSSgDaLFK247atNj4DGfIJcbT5tOikMPKcpwtQWMxNA
vPXkst7C+qkPbQ7ZSQVsbm7OVP1xVU5FaJbVf15ija+3aEPcS0YUcccJvb7L8DZEIuriFPopBcsf
o9OuRF2Jjv5YRxe9/9Tar1hJPoIAOjEog9mvyFNIRHzzov/q8OmJQeflYzewcRlLNACyffSueRlR
DP3YrKJsvVz4wwrDvcrJgwCY3r0eeqXtprtTS/Ox1xu6LGgFyLAXhz8zZvlk3CmQHbxKyp8aI4MQ
5eMXiV2vXz5boc1GlOIDeSeBbSI7TtwLjjtaK0Tng+0LBsZSAC9zfBM+uTqW1nSnabnnQOScMTT6
dtfqfhyeOIuLNXLsgH3TEo0+MG8ezrGZxE6CyERBNRgMEvmlPL8R+UsYJ7ItyoqeJooJE3Mq6TMX
vtRnlScrvP0lOqxTBAiPvaOktEcogruOLu+Bo/k1icNFB7LlM9x+9YwA5KF07IsOTtvjO1suZWS+
Y8l3d1KpuiD91uU99zOGlJZKayx8PjQpkVSU+vqgA6WeqLmGgatFsvofjXToetwd3unE2PW/PTuE
0cs0CIUhq2ja/PIFAQI+j21mLE4WZGR2QDo01xDvL1HmO+gwkMdxyLYJtxK0yFl9SopUTHe8BBa4
HpoA7kbR2TiQYlGxU8Jg6Q4fOdT/5MBOnuckuK6EVYkYFHU4nVgRapLcdu2POz/hzm309Is9hHxq
1V791xAQJJrcpml/H9yupIpxKE6WEu7OXRJzOcYd8taNWVaZGzSjHhJCR3x75jcPruuFbzPB247R
es6FhzaBGnf5F8n/DTt2tL3SDPZwtZNAqz92Y2GaoMkXlKQA1ULtCOE6rFXkpO1gqBILO9RcKION
w/Zc5kj3hyWdibP2m9rEIFYT2Q+e8UIML5UEc2EC/kqSLmzPfMesFueasbIuZMkeRi5UFP54rXbI
8wsR+ZGUWl3QGCfDd0G9JjBo+2+ljCd2h3PdPfFMGPh4O9x0mSGxf6Y5/HpdpiL8VDFq9Jg8NKl0
eoBXS6ljP+vW8zgjtQUhsUYFHQe5LbFPbjLWxVQiGFZk19WTxmYmjJSQrbPusUDgU7gycRI48UmO
Ig7rGNAQtUeu8mY1AIY+IvLCYWK8aIY3FtwL5hcgKzUJihLHlTPcPC9uKPVi/9wyHb6AtPBogfYe
ybDtgt9CUJ8V0tnwQcGTF6mVXRcDGjsXcDIdIfncZovBr+8AIutEtp2NjRktFDOM+K4kMiBtn0QQ
6ZQK+gn9nFzmozUkHUeQsBmcTp2tbrq6bUHNR6CUXdkWYby531O42UmEE0diJ1VQBMDqoks8K6Fs
n7AaXVAEftlqvxCs/Dk2e8SrI9L0mU3hh6+e2LvGjHOwQpNKxAuXIrRK8/3k3wHaretDBczRsY9Y
Tb5Bgi10y37298ppuRCOOW3MpKIS0xMGPaPpKkwskDdiRrhVubx6/Xm138l0XT1DCvh4WNoMA3/H
aA7YBf80ZnvtEUhtNOa7Czmfbx9noxTf+aYYH4tfGvZ/PWv20hiIWpCUaT1gmedMWBRatAI076NL
bu2vgSqBfJr1W/3UjpbEN2//dxHDSZ/v18NTAISk2LUtybEKVett0+Qg+8Qx+gtzcf9kptU38WS1
S6EYt+IKjl4GFOFbzhxbvkwdH2cFMjNuFWuUHcgaASgWnkxJCb1JgS5qN0gLHYwELrsgXdU4KkOP
2g92kWffJnXFYyC3ZLQzxjdkU1x3Cmg6VAM/3IZyXJ8ReQc6BZzPmhCDXKCfLA3crVWArL93Le0K
goh7Y0i4KXVNbdIBjGaVnhRDXUNk+TArmFcibAXxNrxX3rIadNcsi+nM1vST1Zy9YJg1+45dc7Sd
VDCaASTsr1fIQUYxTC701ALofzMX3i1D+b0qVwh+xCzF/3nLTCp0SrvAZm3PyazVAQA+hj1/GYwL
9LWniWTbfGOqHleLF4157Jjus9Sz1bHOBNk7RbZ34WeyrUxDW61UVf8ZnaU6H+yl2nYeWJfG4Dnl
h1HAdqFZD0gNHczO2YHmy+EPe1GWFKHimlEayD7Y5cLFdPouP7FKIHR3+ptQBvcxTN5Va2HIKg1H
BFdhkxRdy0HRTp59FH+MvwwOT1Vc9esDAxG/gGvh6wksVwceso91OrUQd90K+Zrsi2BXlxIXJoQJ
6mVROjVnm2CeNbLTcjNb1IXBuhcUFFoUcufe/PFIO0yvECuJR/nGXU6BPb0nkzvdP3SkpOhTaV2X
LaBK++Oz5NiJpqr4TZ81eRmwso6w/G/Ggb8VcuYJlEuY643ISwcrbY/j68H1z0NUt/kgu56cav9o
qmOPbiT2whBNcO7Upi8s4XFDfvPhR3mpU13I792wKwQLlu/KzktituKUl4nDP6sPClx1cLRfLQCT
7xirChyjsOqJPD95p+ZjUR1mqhy94eC+DsAV0jEN7AXIRuOcNLexZX70sLGzwECafI4PmKuZPxu8
Tb1wUHX8CQsSnMT/iHwkkqsgS/mG3fM9a3wLfTzeTcPPma8bFXllm7sNByji0C/0cG5m8R7BvZf9
JK5GHcVXQZb/IU/ajL/gVMKpH/uFs9EpbGs6f3vUMFBxgoNODakb4McJqfJyEtU23FmmtlvEoZPZ
BP3ZDTm21syaERXt30L8AbPGF5QhzWkp5/e5xuPhn0zS2yeS0NkeH+727Q4jHr+2+Kv+S5ESMZQ5
u95v2UZ2n6eIRsBz3L9bHa43n6JAqlqoMLb7w2+0GeiK+we9E1a1rvp+mSzTk1kKPh0EicigNH4o
IbmvByhdRYnk5UjmBqsY0o1E+FjCi48eIzOuFPdMwny+VbbDWUn6skePZpfbwP2DAHwNrBedONai
71HpC8LYgNXIaODxBXyi5w266/T7GBbj/pLZtOnLUrlCgx+uEAijMjjwnri5dcKIMfPnfebJYy4L
/1HJWYtRjnJUv4yIXQ+njc8+uNLe0uYZLkXDUl5xUPQSkrhBLD/6lsBO2m6vjA/Q9f6Ag8z3VW4I
MF8w4SmR0Fw4LPyWqRAPkEx5ohYdu0wULcrWaacjgt5OwDLw9XReb46lOgm5Bsfjw3m/7gxWrDB4
tmlOtwfgR8ioqxzKNYiKuGI7Jwxe4NFW5eojzpP1JrNdgpJMrzZyr8OxQk+yQU6ZamaSQB/iErEn
SbC0DzqPwQLM82f+VUtUeclYnoqNObB9kIeuRRgYRtj9h7ln8W0g9c+Y1/UaXBrr9B0IjyHd0EQF
ko5ax54grSSYa+2l6Ic6U9UWfYBDoUzp5X7qb2lrCAikJkOx3B1RvaNUCRXBiAcDXvZEqMZlMQoa
gN1XysteKYuUltOfLSgErHOyTzWCfPoe12Q0z4vFhhYu+pLZxj6rC4QL5TrjC7nQofxa6KRBkJ3o
Zs7zcpn83E0Jg2gE9bbodAhZp2Q9QAA4jLZ64rPWWABpqq7IsjvVIfkt2c5bgKvYoafKvhLQHgIy
S1B6yACeTeU3nqZVQH8Y4xvIN56GrVdBMwKZfp/hlbAaILHgUJU9+RXx05YfWJ76d+M8u+o3yFO4
qNSQBzw1ReZMukuSCl0GBVCMgp/R8JsA845RBSRAlWTX+TYgEQSse/Tc5t9gvinzYe02JyoRb8KS
D6e7iYTrsb9WpZfdo1WRvW4gFtdyRO2Bijy+dHESgabzMrdQgYwV1RHAWbaHimjEG/qCWjrVjZo0
dS5JsyvLETm9ahoGbX2xJoO/9arhYjjjyORpVIq82riIVbHtV8QZtkM7+ikctVATUpvPLAf5mJUT
ME5v1MuHR1DIeMaAKd41l0dL+ZaMqCBbRYVweFdRz/aevsmiXJBqVc4sIwODkMRSbjHX7lxJVh6k
bH058JjUDO57j7IUW9zmbdb97k3+dcJ0zLS/eYXmOGBgJhaTAioQehv6Jg5QJfj/vI0nX5reYHv/
NwfN8yTka9rP8nc4m6R1gOM8IlNfQFEMc8R6bi4vjEOdsC+nkxzZY6dv9lyHG4f0vSOqEXdXlMKW
JB9NvXlVmu5uUEo5z5ZDaMCeqiqLOZQifTRsL+OG19oJlD2xmVLIhbHKDxYXUN39mD22dCOmUb1R
KwZVmbQdH+0DCK60lNdTiWifoYYejhNxGM81v3cJp9JYVtLyN1Z5WDPJlpwrHKog8ZUbfYu8aM5C
Ebq66fHS0om8a5N6XaWdEqDW2F7dgEGL7HuX9U9/2pXHeuzmbTYAXS5zv4N1xsVjwP8v8v4AZte0
JYo/M4iX0dbBqtVio3ev3LoyRZwhr+dfd+e2aNZI+KZsgblb9eeii5vwZSi938kzX/tjbh72DOn9
a6AcQ3GGTPAYsYqse4J6+sD17Ks4Ts+w41Lc/5wicoUsn9+5N/I2lbxJl4DP/lbFio/naSofjAMw
QANhaDbaRrqH6YPTQ1tfM5OKYkK3PhJeUe2sBXbIUjBXPBRf41e5emq9ElYH2AfkrCb4FBOGftvG
sg==
`protect end_protected
