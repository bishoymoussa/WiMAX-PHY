-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
xMMp0iztSVf/gn1quN8wGfGsrYgiDs57QVPwH9W6H1uGWYYzNTw403gdsOl98sBbjCXttYVX3CrW
8e+WFvs1Jgy5uzz4PKPRPMofOg1VHljlKNRxOzuMaMEJnDm04QImRGeh+v81C9ByLxKk00FXXHkG
V0SySrIeFLv7JUEWgogtxYQ8MmGsUX0S3HvS6LwdpVrTfcmZ1qP5vTVoaIZ/O1kEcb2HfLEDnb/S
w90HETLcMC6S+jVAU3DttCuuzI+RavyyYkMXJn3kRARTvI/sEk7rODiGzN3O2XM+IRsVuibmn6xa
KHjId56h7sS2H8VJkxdDMNp5/KmGXRcziQkt2g==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 13440)
`protect data_block
RZMxY7LRyml4ORkU6iX6+nT6izE3sYkkOxo4SRw/PQMLOYje545minUnKVnVRuj3YfUtJY51TMmi
qCxegL+8SLARuWxTUNUPX7OyIDKxlJY6CySXLh2BG2mXDkCZkzvhX5euQfS6UdYq8BTQGbExjW2m
2My0TKrWJiEsOH3Ol5fYT763dkg6zXpE1LI0UJxen9SKks7CFplH6Y9ow2iZmXRCbkz9Wy3hCOVj
yrk5myy9BAIYiCzlT2XSccdmnBTI2pPWE6qOsqXHcpW0zHCapsHk4RV+obt5lCInb32Q0EkCtwAh
VbGZb+Jke0i1NL/Tos0GJhQx55sEsL4EIFYO3lR4OX5WVt1E1hIormBqtHBwPNlBavPuM94VBqCZ
Dim6nV3l1MuYvaqGSS2AxY/FPQs7kNoHGBjLFN2VwcXfdPMJ+WGBmes82trOXDaK3g8/n+RA3Upn
hgkEVd1CaQw+b6Bw2epmvA3+qsjcIZBrBwcuqVWfEpnH4i5yBar9bVnc7+MqSRn3JIfhCPeIXNNl
i9eQ3OwuNdK/HAkTHfCgP/Fb9x7JedRnA2OW1TsB2ue429IthUs19lKaQ1/FN3Du341hgpdgm2/O
CXmVQo4JUz9kH8SJ/vyKf46LHBRU7J6WHqnUjuzNV03nqkSE8IbultpOMq6SX0ApQpwX2B5AlE++
m78o7yzBlnUvMbyHKRTTyifkjBLKr140tJy6A5KwNVaSIZW2aU16TzdQ5tfOhyii8wfCWO3dqJpl
y+YTJGHtnKm+PJHVFrLlfrZ+IvOwx2+B+gfjwhTeMOGlWgwwrUtREzSBI9aD8+BPMqal9abWuNh7
EoxSL8kQ2orwi7Bvbh6dyESeRWUd5sQntZzCIDS9r4cu/5dbK8hXZ5Jxy2nIhRLzz8cJPI87c5KK
sR+jGb/+fb88djST8zyC+szCLrvfRAIeakW5VxshXcfd9m0J1l5FTZB4g02XBqz8Eeo+h/+V30Gy
C/gV75uX8NJ100u2VMkW+WdykDZwdy9Wh0/3OoyUPKZRjMNTozGgmkYn3vDVHUpkStmpov1kdT+3
ao1n9pQcbNAjT137aW66hBSZlsUHWTPgMr9eF1S8/aCmXj24AskJMAycr0Sq8WijfhtMXJ9LL94R
ZTXl7rc2rTE0O4mFFi7rXVjKZpPVxPM+vLnxunEVoZ3oa5xAGMGder1Hk6+EJg8KM239i27gye9i
uqCVENfmwOTqheMD14/e/SVXJr1OsSMWn6BPh1FiZvyizIvep7Ij7nr1tqH3jcZUzOL1M/oYfF1j
uzAEavaxTUwyVVeZ/jKKkc79Z2wVSrZhqNB7N/01ubwzKJLdPzK9r5wK2dSwAHob75ll/u447ayw
W+ewvYyfUICruYlIndW2xd5xTxHaLCwOSjb506yjZBP7ffzbFvPHFRGybCYP5MGaNROf2AnnXbk0
/hCfrJ5HxW4Bxq4Wk7eF9yYyEtWXD9FO1it4zy4BDDIMP0qMEE/LvzDORFko8UMN8nGkoYEUmvnR
fYtxIM686zxzweSussVYI4DrGtrktSj8tM/atoqSX6pvfRVeDcCGyQZ6BgRwEaRR0wjvvNfmGQQ4
pFSzF5L4IdvguaUS5AUs9npZGyY08AyqXGRBPwZJbhNgH7xxebjmbhNzfY7dqKSvRl7140h+b9o4
JqwdvCPI8MAw7ShbbK7uawYASULbE3VJ/l6eDSVhMCGQlZXs8Xxg7MnIcjYGpFChmJVkV6dRhzYb
xe/NOfGp0erkM9yUKzJIW/1YeT9mxXfb80I5tKOk4iX7tfSlYEJ5BkwJkS7xYwwrSp4k0iyNRuwP
rW2MxVUWEdlQNz1ieepoAOIl6ujfVNfuLXLLbqtHP4DZafoUh1VovGttspKvLDOZOoYTrhyB5GCE
mVt98/9L5PXBTzv1bHmwoJ4skRjJESUGQIYrRnmQs6iXcY0vexj47dA8gq3pvqhFhRJPsoS6yd1e
Aoz/ow3CRYitqkRFHtruRutJDra6inWXUOKJxPA4OFbGHC0MSMxwSCxAVyvDPUgBYYWCn98CJ3kh
K3m8bkjEpBZpPtXKEwCScZhq8SipXQ0m7eM/urXbhLKpFCmFGd3bGU3uzl90KDhkJUrJ5BMcVTte
2kwKLt0hEkv3a53plUTH2mo8XtXI19HuiY6BWyrEI5m05bGBR6mXIePnmpElKDzY3pkUoyGaCWbM
tNesOQ4UHnp/L09ErOpR1tysvT9S56I5nopInafItt2mquD60S2Xl8C1/ZX9XfHasPcuBk3dag6N
3donO2yNqA9B+GrumA6cNxkdkjLBU5v/yOjtRKRgALK3EDz7LotgYO9TwgkrRieSar8F2M2nHzki
huDJ6F/scuqQE0sJ3C+qhWFyykN4o0MCr6yiruxN0W/CUkESUydAJkmgWVKWS2B647jTq4cdnXOE
3QxTystYUP+JRTFNXxhmuACeSpSdjLGiw6m5WOG5FPqEUbfZvSMbyHQy0je0q7gtqEOYwQwasO8b
F71mkm+qQxtuje0DS1CNPB9ewKXatjpHjgAN2KVFZW1WyuNbvOqOzYtNx7YS5gGhRdzxa3NPvMaJ
5b2jRLtvn+RnbJuUEKnZA1lR8uqk27+gDlKCO2DeXPz9SxVg9Qf9gUMu5x4xqV8v2M49ZTNQ8DRW
jaJahYvkhiOPWr+XlLTXpElFPfjk32ZxgDO24wZ+yVCZhukmZyPWoGMKybyzdIoALcM4Otkr4lpF
Yft2CUcOfABhhtns6ukpCmjAqw59aJ4wrFK3thrOGBwf5KXP690A5G0JEzidXWcyLo3pObJ4Ub86
j3a3XamSu7HmUr1/5VhNfP13h4BYCYrtyZDOrjKphJfvDEj8VmfgNQSoFmqYVpzXMpe0gaHX7Mw0
LqL2arXRngrl8N23TAfF3aOAvx/neP750JiOvvHPik5FekKBAT5Tw+bmndadReRKZBYXFNOyTr6y
OVzQ0rtbvll70aHudvWcwBOa6tB5ge3m5PGBrv107ebSveCQeCjrPbT7CNvEhn/0wEGIxJTe0btN
u2OUkygIZe6jBW574jFbpaH1KFFyTbHeMVETi66R3F/ntWYsRsbK4iMMsaZ7EEGvOThmKQtaEoqP
NNgkZgRMFKWR5m54rKXT0if9mNoaTrFApLlZQytFBoHec7ltVfiYzydK7r5CvoKu35OFMgvNeJpr
tF4IJwBcRFDQYmLl5lkqUwXCwha7sVOKzq3K9pbptBoNRIcmqjFDZTkg6jefBX/hecu3xuIrlUN0
Y52mGPp8fXNwqvAA1W/8BzITkxG2ZuQgNfjAGssDZ6e3kL8iX1SG7R7b8waFfpSq1v09NYZ8PXFS
oo6Tg/dkvHxILOpPZHQxvCdZgZgnvHthe9jcJFyt8lx4qLxiWkWELIN6USCuzXlMJdltyyP20MOR
rcKoDdl70dVGpbxYlL7I9EUfgqe4RpQapqDPAQwZje+p5/FcyieFuBE7E0DoWVrsC/FYQxMYFAnN
O21ILwK12qXfmHlrUpfLSTMuEfPje6yA3s/gOSYxMA9BR5G6rn69OXujBJjSIr492sZvSSnUvHdw
aYXlRD8LyCVsBmjaxwbPL5b/fIBfRFEsF7JnCNXvUSFkr8wppi8Mt8TrKFMBRauTlvG1durkUMXM
1LJOLNkw6f6sQvIrKQCqFxU8gIEBt09NPWNisAMmAYeVxpMpoV17ZnQfY2ti+fIU1YfvybSifuMt
AlYolgDtaYyWUJamCQCTH/E+CJNVr3oLTwKPzqv4CjrNcAv2Y2PRK6XYQdUh378KImMLO47ApMbz
x32bcQoR9Bfxu0zV5ciJZe1SzAxPteFBFu/+RNUamHV44zUAdN4rOe9YOGaxNTtsDURccXDIUzGC
cY36DlXgy/HhuI9SX8Acg2BUhiQ8fk+YRiU3YZxWeAJ4zvtyQm4EMxMPfY43W+7wXYUkhNDDvJ6d
TwET4qhqiCK0OPIX87klqqvy64TjDNfvpSU0qalxFRX+iaZZ9KjLRRQM7ICuUT2NJ0HY9HE1GUU1
JedSTcPdYbEb+9hDqlpMgNiOZy5MI/zu0BMezAdx6wvfncw46mL5r3IId1XTQvX7hKE2YtI2oUwt
hD4KfyeUMabmCZuczv7bhZXjnPx0n83F8WasowJP5ov82Nqw1QtbTa760/ClGRG8G1JBtL7Oidfs
VlQNe/YF5kK+cnkg0rnJ/EaETf3UMv4cU8uZA98wBC7xPZyRodQkfQBzh9qfwOCj5CqMymyahW0x
5uL/noa+DRkzpRg/Fwyh3imDbCb6xWGw8qxGy6HDDilB7vxiHZbnJPPwmVgNnmb0o+S4gJ9idyTb
DikVwNlEyc9y3HLCTJ3+iAOelAjh9u4MTQOw8nDoiEDywqJN2/nKZkh2h3rtkK9EN4CJODhjT7un
G5Ve591Lpl0+FnDuZ+puxeg0TSo39I1iI5g1myoh5cp+Y2wb7halT1HjfzvoECGGe2n/6m5F51S9
g2hVDFjMCFe5pwZOwW2ktoPqKYjhLtBjGrYkJ68PlZJ3MHaio/mG0C/kF/7OW+tp4e5wW4JygyYv
CEXP+9hfSC1NWi3qQuRJKiW+C3OhUtQ/1DSkNYy5qOjkfabrB1DDod+E+/FBpuBGI9YezkO/u6Sb
H6GIl44/wuPBvp65sQMSKwz91F6F3DkPGNZ025vZDEXgmjjBdGZyWpxNh3wer7cBN+sqq5MOZA5k
M/W0YvrIghAMN4kSNHhyIO8digWkX9x+9JD5K/FkbMZkbTa7f09L6RXGfpDEZHOZiyRSMln7BPPV
d7fqT+Dup7SUnav210ENJULwwkOFyMnGDUQBbcfgLC0Azd34MGIhVRSSsGvfhx4+giEtqrFHmz3Q
6QJOv3QC2qiKolQ1uQHmWfnce5Qn/2GtFyaMOBj94pSKVuU4G4FF2gz5Ro3Ij2fAWCnJYTO7IfIR
mAn4lSoNSAnvVpDZeyCUbkYXiTxI/IUYu41qrovowyhWvIDFdoKxQdVGCAmp7rh+fqCOLUfeemp5
+oj4xtSE07v2+ZhCw+aZVqMaxeep2sAdKLa7yG54LYHmxY1vfBJ3mEFyc/gxUpPsU98u+rvJFeh9
zc5QtOM1icAWH75wz4MoQqTB+8qZgvJSujeuzEncYtsX73r9v3KDzHOV01wkqxcubgXXaUMCBjIP
Pw9gFh9CCMEPkIWNy3nfuHbaDWjGKp1WQQPGX6yNEK8zxhgiLGufOQLBwPC9Wg0ght/D85qYNF7C
orYyehS1gAlL152UPP8QCluUELuH7xW5eHYBn8NbaOTKkGC7OZ/J8rpq97D8Ec1Gy4QxAqv95bHl
cLcRpQACX6ZhOv03ojnItCUvJsOvbw4cFWBLgG1gFJHKmUWJKWzO8tBzcsZupbyMXdA6NGYoPxXl
Yqed6V0Tvl6JbPskGGsX71Kqe1Pd5C52IJjGpnnsI+CttKH+akPwJV36Sl83/Vdsaj62JDIsXJR2
PU4YDc31oaZYLWrdJpNTFrEWThkRlWgN2A+UeTYsC7OnKWjlrzUbA3BW9GXtqqWo9SpukF3HjUn/
hW1M16Tmk6ev9rXXtM27intJIJWUKX8hOVqJ0hHp6MlhN2MirXXvPuzMTNNDm9DDqQ117hZi4CjY
ytUa73CKT+AwCbew1e/xN6xrRzKVYf2+5+3IgYOVGtcSWDeqzsYtI5/7fSaL/030dMmMNaIkZZuC
koeWQubsKwLRVjun3Pb+qzgegETrPQC/JIa9Q9rKEvjl0Wr1t0PW052VAZ3fMhLl/t43uw2Ia+LA
wwCpbrYY/1vnUeINmopiAR0KRhasHacVePnLBzMeyDTgGIVescwkRzl9AArqIWcyh70XTOhFHaiy
Sx3CS1xjlB8EC9RwwcP0Ey/RuR7hcwsJSgYv+2FfgSnagDQW66kygxT5FLUJlob23tnLgUKBDQpO
BJMgSAlCsYxLfyQI6KP42x1pnFWbo+l4X6n3eXC3u+DJMHIZFDbyOnxaE2pqu5YREj+2lW1EzKW0
XskLcOC4PgYhS/d805SXxgELbz6yjTAy/iar9HOgceNU0hEn2XN1IIo0CIKUni+Vlr4tOFMMEgkl
NrCJzlQyIh/eju1RlkD4Mh4W8seAONWH+IRwAyD4otIYtrRlvu/5L4xSDxeaQ6gh61J8peO+zT9A
8rfrNfddzDu3lbzG6W3hP2DYtXmssux/Ousn81DUyMt7+TUWRVzhPUS62mgfyABRihF/0HnUkcRa
GyGUXZhKf98ctRmo1ptl1g2/FKuS5LYA+5LO+AEcRZBUHLhSR4WoggEwwln28u+EJJ4XID14VZBf
lf2mK/CXAC/rwHQR61BFgGQl4iD3GhW8vNwQVJqI6UDoCWCBWTASnbwkC03WIoViw2ZPESJbYSd3
HA3XkefiX41FNneTI405MSs4mKBftUIWYLMb0aptyj4PmWstZveK0pK7rB494PjHLEsYvRigKUVf
awdfZz9Nz++HCcHiDrz6UGx/tgLNqWpMeBDwZLskPXFUEHWwikS783RmkrR/omCTaqm0zMuHaX4d
zWtEeMH596kxhjwjOPz+8SU54iU1fhb0SprmCEY1HMPAuMUA9DwMOQ0J3zvwVbNNOTrG4/sBNTHl
KxoO9amYUE6VaGuG+8MN/YJTJIktQYPt+kA9gpCzxeJExx1IfX310sWLaXLQ44e4Z//I5MD/pYBw
rx5yLEbsmtYOmugNvLj1T408F7/uL5/W0bxk3+Y0O7MlHmIAnVRLeDZSMPerVs/p9fEKFca9ZICJ
wLwOJAGv7npl8D7wRRZ0qNaWeqXz34fhOMBDf+VUsbzgbVSQVsd+t56lnUDQQio1SUAix8ohgzVu
gUDen9Oek47t3XMXH9xzKHDLvHgAMZB0SOEgEBBy7A4LLRm5j30WgsfN0mMgXyNxdJ38iKcnRCD2
Y4NRrYijNsKNRvBHBCSbVfO7Xvsw0n1Sa/lAvAMx3E1fuTSAw2cKOI7uj2WjcX6lEnOaXYNus+wS
vNg3XWNcSYFCDIkRY2RgPzdnS4QyR8o4BNGEyVIvHHzE+iSLypQm8j4V4Lc7eXJCeRg7bgw1Rmr8
7LRfOpymnVL1tG6IjT9k5A6HZAoGj5/YzIRDYkECx5+CRkHY8yIt8u8Xd0aNulbEYJI8Cc8uZAKw
CwdFDeZAcUFvkHwJd0N8E76cJvtlyJ2WO9zGQeEd4kVzVA1Y0kGgOenGHIsoSh+gvv3nbIk4glf8
LYbOC9C671CONVLWfKRFpx++l2uX3pIsa7dDQeXsfeBtBJTX9bt4yd+J7TXIKd7iaBMRH4vegEgW
I0hwR/8OemdybK9qX5O4hPgfm3/2FS/jgs7hw4q9+08Vbe6Dilit/nPy+KELm6YpYSa1NO6hhF7v
VkOjtAhe1fcXvh7aMDmG2w/CebfsoFHPCozXUnDTm4e0LsnvoOj5Rk3wHnke36e+Gyp9IrZMqjsM
RMnYoMuv2Y0ocmVeR3OXoaEOg2uy04zXz+mZYPs/bb22QZDZ2xs4yMouuIJgy7qsvvrNbhP49Xfw
SQmB/kngjVDJ/VaUkwr21gfRvw03dHm0yNS7uBghqMic+GEtn5mDAxrhyzmPV16HgQKopwSFlAi1
ReS6Re1VQC3NPHeHOXuM9CVXCvF9LuSG1UE+Z+R2yirNBc1mnFN8cUS8o6YoKYYH6qMOarW1HU6s
23PaRnKvjxuiYMk4iP/XgyY1gw0oKM/t2tdDcDAFkIkYNLrXUVNBq4KHrAgKid/CN+ra2H3Ha9qP
VwvdRII/yBIhHufLCI7DrhDK9/N1xfEPGGtQEqyZ6c0CE5+SS/090ZrZlUjnAmSyAiAxCu+/odiH
4aWwWSI+fRZKMkmAgZT8k9ioywLfLmPORZRD6vwbTx60/3+K+D9hz9rfQNbVsKv2Oh/d9Drusuze
HtxOepIZ/91Vt37Cp3rYE5HBlJgZvREJ4UGVRyfz4M0N5n2ALbKxLPySTtqxQiAYot88p4zpdngT
f3RIsrX2bTyIRxhFXamdICxZ75ybCex2bufaaumhjJWo6bWNyHvfBopG+L/hHemvl3hSgcT6hrMY
IkGSaY8uTINW61ie7QN1C/XEusSQRss1eF7E8FEj8/ttMSOcboIGCKCnbOgRwP8qVZ1XqOJdA/Aq
1OsiymoILiy4s+dMHuZRAVIAciInjE/yixvsx0SCXWtwq0h2kmjSWT33vDZsowPZA/Cdy7sstASN
ECri3KAw9N8Je47SKwI5i+mlJwv8Va8IRmKcepV8vByLUsWbYqtZyaCqJsrnCAdD5RiG/gE4ujEx
nf4fjZ/5HEBJVt+5NK4DpllncYEkx7nKUOfzjeQc5DcX8tl2A7hKGezQ7H7s3OisE9hSWBG+Kku8
KqR6CJXpM1iAYt1Bg1oYmWBqe6mEjlbfspTs1Smg3vcJHNvc10Le+X9XUUJTkiiAeWLoytQeZg6p
4OnWEg1UTFDbKsR8IDYXcUAUCPzL1JzEIli+rDb75/w7S0wti48I2kL5Hpq9vziozkdMuFIiDlLH
bwSVF38vA84r1fHJESBXjfNrtbIq+o7xrzhPW0S7qJ33bfh56ZHjVrKiRjjrPdfJHDOmO3/qBIJE
m3f/f84mdrQ7zDp5QTBViu34C5H5NuFSBJP/Uyop6dDjojxGWG21kQuvAnNAUCQE3eeAoD70JD3q
KBlvJl7qZ5Qigq2k2NUs3p8YK3m6Z/ItdsApQXZPULmMk2wN9omkCuEVADCwJvuqEx1/KubuXN4f
1usflTWhFjSo8Mg1YiUH3n5xeVLN1NGh+MyA91RQi8PT9JeslKnxWUMSJtjJrnf4cqRxX39xqNIa
W0XISjR20+9sQowD7IQw2CoPuoV/Ed+O+PM6soNbousTJn8fSPg3cULrFg4m5Zm+AYlXcANT1ZTN
M0FQMM/MOM+5IkcwDM3+kXiPweuRcUKMsoXpWQtfHjC2DkXAorp6ZqSdL94TMiEbP4E2BdXBrMS4
S1OojTS/HAQPB+Wk/iMLVtShz6ia2AhSwWeCPlH1vwBZmIoIXxTGr857BXZxW+ciXAiKTjwzWSRd
Tcu9mPxKzVYVKGhkzK/LkjQ2/9+mh9aypFjImrGuGqPR9DnTKB+HQ7YTo4idP27WwoEZeVaERK/z
yYn1Ryh7kNk/hfenUd5h6uVg8mmbYyg/d5nmB9HNth20ykWf1BU1x8lqmPfeNYQQzW92PmYHqh7I
OGJ7W8oxnpZnjQw59mavdvy+n4BJsAEa2vw3SZjtOQyvrA0BRI9+fb/7SMMHdHfKt5ZIIN+XkXYi
bdfC2gogdBSS1fI0vu+RfCowU2P37w4xnbR0b9l9diizpSvpB9z4Tq9Cl9mDmkmUib0An5mt9H2i
3RffsPnHuT/SgEuR0/WrvWlF0ziRGNtAgRZzCegi6G/fQAWc1eqIOndCQysI1TNQ5w5u6/Tz0DHt
nJrwxjX3HXS9o63HUsodIKQ6IblJL1IF4PhpdCjKoOgjqsBJPoPiZFrpte7aJoYxtMCDMzTUo1Vm
LGTw5MxrkooY0yn8J6cmDTzjZx1knrCqSlTNxLmRLbByPpmB9EhRvkDCKCW4t/1BawSu8jpCG5pe
6g4iZbjbhZqLIZDHiRPuGCKf5sJ2a1Q/FrXg5EwscwpD00MmJyBC66C/M0GZQiRwY4Z46LiOn6DL
DeglsYOS2UkUkwYkeZs9qOKt3PV43GLfZ9wrcS7ECULBcKaA/ISvF+ECCv3V9QWl+t0eQxY4hGeF
XaD6qHfaJ8m7patVjwQ3hIysyXrGTOR2jfuThqFpGeHxRq25L+09VaRE6JEBTpMiy8+bYrKkfMVD
OQauAJg59Qx7XGtrHuP0i2sko9Q+Lb/8eKIFypmaR+z2VAvmWAyBd6a6fQdqjOmpS47xN06iS/Qb
uLxEb/bkJ3rWoltQrvb24kZVAGxKNN+K88oKtMxSFkf5ZexPdNLS4easjevbt0NMHTVNJLEH/wmH
nEmqwZCiKbPnLN9kH0fDK1f2/xF3IM1D3vi/krXSFuNtOUREzK0HvXlhkSq/kwsGXu0SoaF0kLUe
hZSIoveAZ2BtomhB3l3A6XmJ1VdrFcKtosGxbYeb/PnkzW5PQZGYRt+3uU3g8fnS4mXekmKrS2cT
d0797YLtZzrYCrFmNa1x2Jy7dhrCufeERGx4z7AmBpxsDTDBD/kIVmt/pV5p/MDJo/mTfylYvceN
YIcwQWuMbQp3pYxqYLZL08BWsD1NJSd/iOfF2N0ONg8Uy8Lvmm82cyBU9zGO8itLR4n7ofWVKkPO
YbUf+aQMELiYUZ+ostIvBOxvxd4ZJW/yWnAMZFkbqrDf4jpGgIgwvTYqnkZ1c9uNHL7RwEIw+KxP
4qqgX9mN7ZNDjWe1Nte2U6honrpLMciDKAdd4vzYIARFzmELkPTGCoRVJnOdaP6jYJ/e2ZTwdLpA
UGq3VnZIRy5TP/mmjHUXCWTr756I3F+N4IqXjoAhstSSNIw9Xc9YiDAjdMf0aANn9Lijdc2Eyw5H
P3WThu35fEk7ABbyXDqFVXJ60l7LzBfr4ZfJsBd42Nm51bbpmTEu+pbzYM3kr5PoNUJk1BeiUdtQ
xu/Syk0hLAcKFynnrUp0XNHx8BQY4TILUMbH+BtpxcbrYA2zKaBuXnGH29cyO6UMJas5xjLQkUe1
d7P5/acM5U9y+X09XWsFV6mIWIxBfnZa52usUrE3ePgfLFZ4uNw5cowdtcr8tFuwJboDlT2vaOXW
aEf1l1+QwgWcDcSn9vqL/DBW4j4syoaCFxch2dxV3rzbzWQjGBfZX34E8HAEQG3WN31UWPZ9idHa
oI4429WEGSOGog01yU7g+AfXCmFZGx1348LmyG+9SZi/JMGMiIhZPugIYkf10lzwLZcZghnIyTRA
AmBztf/K0ZJNivEdD6Eh6buHRc6M8UvSg1Pw6DiiwJq6gWunyLl9kDVq9kGQVIFKnJQmhsqUsPm3
5Ml0sIcMHTY8t8WR7ldRGSXoF8OhIxH/FOFYqKEcS1f15H8OoqjfAz4jYAhu/t/WU95R26FdcV6U
KmKkLQwTup1Mmmp08edQmozrM8IO1MLXU0rhP0zCOVl+vRANSysOo4nLTeL/qJF5kbZUQZW/0wt3
MU39gzGiEarHAhfkDg7GN+HEX21XPYFg+i1QGCPNoY/1YRms0nQ5ZcK3h3orjLYsat+rUpZ5fb60
oL/arImGEhiPJ9GSOgNkrpURf1unzxN4suHQXmGFXUpoek4RSfCbOqj/BTWSs/bNrmyycp1h5aWl
DbrYMbQbaOs2HKiYfj0nYnCSuLK0qe2XIfVjOZPESNh9HaJ2DXCoMVSuvgSl3Kd98NjvazKwDlNt
P2EZ5uBPuTzbquQKH6vWZ918PLkkZcIOiDC01+OO6vwIBd+VZYquKKTqaulFwZJ1CiWo5iF+rdBf
xzQmPiTDVHHvVB/6mwOYk7GEOGeElzz3CpK0QJD1r1Ry7/C0PuhUqfUKmB0/Urfr55q5XXoxtS7N
RjrfCWG1U2udxzzyg4OR5kOfO58Bmp3PTIqKRO5lo10b2fo+sUBNsJjcLoR73QQFpxiz8aXpsDat
YAHvz7TDtvr0JaELpxTodQFQI+SQJ4x4S9t9/0jzWSjFp1f+8Z1CwPJR+DY9OBVmzHfJ1SgPC+kk
HKKpoUIbbzFSvDjSWgfTyr/y9/tFkeP0AsehRCrGLFGmmJxJ/W/37bn+g4aSFroNo4uXEHNaoU+s
wwdZWqLydxyHk7IyBX94FczTncRCc0NCPGyUZfSc7JLigv0bH8ODntk+cHEjxtg7zrllP5bucEqS
xZGc1jfR47ZsRKIRaUdZ/mpDCo+Yag6G/LrKOu5HymgcHDSZjiT+YLTXUyBNdCUXlKZaT6VP5Qzd
RgSh/0yFq5nBYQ4CQh0v7jBcMHTx7suUKYzORj7ktKOHByM0MMQMCdMPLE6wF6zf/DZHXWFIIiSN
eMgewSB85c3CLBT4s+PCrqyh0QA7yCVIEO2HMULE8zuI5DBxEWcmcYKZh+fEVV481zxHR4Hwq91d
Lk6U4IVhH7eoBs5389EPZ/QYyI5ARZzjD1iX/2a40Lug1SiQD0/IE+QsIJmPoddUeccxgpDPk5T+
ZpJRXp92brFdu3+SGeNG/lXS2RQIxdBwNgekeTJNbtEmW0Kj15Nh/XWOceLFitWGSZiWHtp8LMkF
urtXRFliY+Wf+WsSSDULVYx4qM2vsXzLB2ncffrx3FAhsBZYJnzCnlXGn13LBUbaKyog8gpqUajI
MIotG2JI8b1ZC5cEoaPeDn+eaYErOCFou3Qhtck5G6nhzZ+rHHjOXHoq3dOPqlKar8dWnGpbJvu4
EcDoPV47Hmjglagc1L+w4WDD/zgO1qk0j4dUiEYorAkbzDKWmN2FWA9FWt1NNKThcWV3vJubIfN4
U7pdKVJxZ/55r02cPyby5lhr/fWY8buVV8dv7rapU17NAatfNl/kVfj7pc5TA4BdouaurAEbN+Py
eT8ouMg3iuLT6lseadsbBnavqAgPaTQtaPXI+ed1fzpGu88rBdluCy18ISCAC0xd+fefvf8hTDuV
55ztrhi+CnInGxYdvYZEDIxClrUEaFWo9L35+hFn2e+HdDYYA6/FuCm78Wq+mnnqUD7WiEuECF/o
cG+61g5AXG729jmI1NwGadaYIq0mWIlz76JJ/j3t6or3sLwvj4gwBzA6Q9uadWNlTvGyuPbvkBfc
uEaVmd8ijJSZix4xSfUAeLc6czd8yIoCyWSduogPqKgOR1G/BMreaT+NpzrPwH2UfQUsqVj7YYPY
3Hntz0RyFIkMy3UomfSZTJl7+gDDA1MpQNstcL/PVbJQq45EEYzwYGoW4OWSoRxyPaK7yEaDer7O
B/UmQhxE/OUmstAzxxwlR9jHkQ813qbngLZ+1vvwdLCR3zxZ+scEFHdWtiGZrnuU/qrAuhmAyW+B
muHslKNBvReFiuFY/1Jv2tmP0ky9VjTWcnHOR0U4IzN8v6CFon/JsHnw5Mm1eQ2mCm+uZFCYMlVX
lbTpu+t6HCbYFtTRcvrcyz2PAVzJYfDfrBKrNoegno5QiD8nJcSJUxEodEY4JjH9BkIuSypodqpW
VGUlKF9YUqN2oyCkLGBoIHM8PSrz6McNEpJTWpNzvTgNFYwAYhFZL1BGlnK1gQAGiXPTefxPscP+
WMAHSNROpgtTMs6FGQ2UBWp0qEOpgmpWMOgpa34mxm3SZzZwKl7RCGQUK9jVi9Be/Ppd+q0KDYMO
1XitmrwaMK+e6nc7hp6AGaEG57gi9ex1Us+G77DsTZTLQuNjfBgQztBywwSayYWaiQIaFPogGvSe
CY7lVlz1ga1ZzYQ03v6rhOgiMuxFRXgxsizG7E37WVMPsOOeCBU1aRM5MkKrROay6lG/dPzaSHdG
U4YGAhf529qFkPkFTJu4bjA624iMrZy+zaw2AYdNNDuLDy7+0dnCwUpMPzsPS9j39ir6WyqIP4Ia
mKVpgCJCT2yEM2ndi6m1CCVV4ZyIDs2b5dPYEt4m6SwiIjPjoktMpENY1whlyNvF7yo6O2kSzaNv
HrujI2CbxeYOYwUsAZ/BQFbO7rGlJczjXE8mQstJl8BYmstzwn+NY5I11Oja+OmtKecE+oFadjgH
NWBPWi5MPAvyB6ivStknBmAKIHqYDFikW3XQER4HQNGBUDgO2vkgfa0Ssjgx4udLpoHJEB4NI+qZ
GEflw8fcRstNq4qfEOsQK4Hznpm6eJpwh6TI3C9HuP3umoayldUnEVYqvcWg7nP8HLB93b0M9RbB
8rH5WHlhFL4BjgYA5xRPOTP4zdtfcVu9/PqO4kXayj/Li0WqIxO0NcpHtiypTUAov2ShWCQZ557h
Plq/biPCjyTMM9JlJf0abphENzER8GYopfKAd0mNRchEkXvz8VgVbitBNc4OFE+SRRW3BHYLT3tt
KMMeXrPCm8F33XtC3tBWZNXom2DPlOAO7jDiaS6J3sqzY3FDumU2zRlcbB34p/lF2eRuXC6dOLG+
E2N3JFVyEP2pol0ytnXSB7iNIKMzVQnV9882AzCdDE42xKIoz1uQyT8O1WLdCMU+WD8BzLXNdtGa
OMsjOpcivO9pUAQjvyoD0VetS923OrcrznjHUQBq9v4vhAXsW9wBs29i/iYfHkiiz295YDvn1zzj
ysk+nCmk5tFMfRoY2lDtmkECtKTquGMLVNTFKD/i126h47lnjmJfxpyompmF99l0wBfiQCRIV7Ir
KssR+tKrNsSh/vsI3cu7PKe7Irp7s2QnjTY1KfZnvszDW45WMPckHv3Cvz3oJ41RFmeZyyAvvtIZ
6rmqerz7SwI0nBW2tKgttgZ2Az9DrTq+bhy0CpHjaUlFPUU7D6pj5lsqw7aivAqHE9Jj3rqTMNE3
Novae5XDQIybIBdCp3FVdje+a6dq09VSIMa1scBY2VG+mGF4FoVHyMW75alX7tkxkp83D8XKPNFx
z7yymRVhO0LxDm20F73ma3VB2DU4rs5Fk/dcTrSVyGdHWeW0JhQpOoqxe2fSjSO6hbwDmh+6sADa
5Rgjnd7dnHwcSCLKvdoJOzuzqHnfYFWC4ab5EzXg5bZxP7JNnSob5Mxoe2w9pAlFog4VS86FwBei
5AZAL51VDFGS9t6h9+Ob9Fdl0KQYx2HotERo5KncZbr7sENr0yZOAkwSOlrss+wojuzbAqC20fNH
n9g+ApJqAHbqZVMxogzcApgM82rwzP0zz59YGS1yQ5DgO9yUcfGkZedk/rJaVn+umLCdvZPLW/wM
qSqAfqnDWrP1/6fV9cZD4N4AcIADo8jhyuwb/70FqlQFseu+ps+c5Bnf40xEmYVN909wFvN3W9nO
pe5gRghYSoj4s+H/uJx9dL2X2mn5WUOdX6tFGIPbtASQ3ETmzjazBXvRD4mKhAgCzu35So/rS1vA
6d+58V7LuYGOlC9aw3niGmN18iHQIkdd/1p4TYvHWI98CuXBwfkrL3+d8ZlidJb5KVOdQFm48QB4
1YOFkvvO6Z/BXRxQHsSKvOGPOYe7mtA9koYAh5BFO9xYFZrDcna2aStbsPT/AO7QIlNTgTVWpFbL
jVGTcZNlb1HPa6J6ZkLyM75A6aM2yhco0ZyupiIxRR/VKcAd9A2VuyzLsJEFS1HiUhF2oe9JlPG5
qmKHHXR6vslCTym5+kCRWgiyoTF0JGqzE2cSeXhOzHapds3QyLizLZgTcohyIFpxZ3fW0pRcf8C9
dYsT4Afft+xlB9/OgWT3CTJI/D/9zfjXBae9k5C2frh3OaNFsvb2QdOvrIJ2J5QNbPNBRAXA3v1n
SpF790hbFwN76iBSnK4fWWkTQJKbgEiuDAw9lV5dg8Hz6ddGSPSQCbGiiuL5qfPREroy7yMUbrvS
23c5/0QmyZZjfGC0gzm3TjKrmprszVfaGnYCpyg2pNkmfhpY3CQBdMcHB2WWXrDjp2kOi+qSFPXr
iiuyBJRhMnFDZ3qiR2zLT1BjIe4CWS507we2hvh7uAPd0Y6NnaQKU6zB7KAQI8WDaGMi17bXkIcp
EkDludlW7nRr+KDPX6wn/NOb+rhhbgl/8sozFR6KQ5F62K48avfEC+yZM5P0yiy9IH9sPbonA9R8
ZK0VjWiLKcMnZWC8ks7na8O2nAOCdfJQRo+4tpKCEuQ6BYrVDsPWHlcT+Sr3pkelvv5xiyM+sbVO
S/cSl5fdSUz9MmmxDeCN30G2Q/R9c4jF1/wlbLX9XqHktejKNHWcIgkcAZdcIQEO5hSzwaTI2RHL
L+OgNu4OCnLBdEGUtyZuLBGGxRWJOVKfbm0Tu2aQ47mUmVz2IO1r15ViGvpnpRf+Dxk/XtvsYkHR
GB8p/oohqTmjvGdrKzqL0z3L0UrO/WDy4IIy996nAzP71lu043xp+Ie4Y8D7hroCI9m3v41pQn/p
VC4l9NfITh8tqGbKvgIiEmJ7pw/7j7HTT6/8APhV9xJ+TqC911aGt1NFyJO02a4OOjB0lUP4YWrd
z52MAlHEC7fKrYTo7T/58NqndOgsr0CTKvfmbPTBLTsoEKwRpc4s1MIBdS0VhnRKQVPI1IcQ0fbb
F88Vnio3E9Z/IFSgjFDAKpwjgXH1TM9M4lstSlPAc5zVkygNzvTXMV9Kc82gv7lS3Sqb7PjpI0g/
vMCEfE6HTGbAzRPxwj8mXKJZJxOYiBKE54VrsEWpttjrK0AqKXANW4tRs2GgNsSr/yWI332AcEyj
t1cFXVw9K+V+FLWG/cqY6rpiVnEhFOTtElq/94XfQvBsBjtT2XyKQ+GLMqtOa4jzcS0Y5oWYztsz
48Ll8MceEQzUKH8M67+LL80I67WcJh8GuD98Hy10dI8oTLte6N0YAATsZptId9y+MZPh7e30GHi0
SRE9HBCWRdXjcMMTbVr7og1/dUHpqy0QzZqKTT8BLhog3do/SOslLe9zmx7Tb0e2zDY1vgtBgYGl
7QGAOrYLTw9dd9Yu1fefT344KPDFnnTwkrCyf/DqzpCRVzDO5+RfFPKr+j/aBv4+FYFmfE0AOYci
35Lz+gngU2CBG0jn4lTu6llPkoV10PEIDbSfAjLknuaK1GAnAgJI8sh7Rx/KOsPPGHFZ66Cv4lgV
AUWHLNRHxSpvImZJ8E0zqGSG/hz+J6g0m44mGjbb36/OqKxIh6PZeAwvctts83wPvSzzX2oDrKT7
ccdgTU2BsgsH466JiuZRm0vGA0U1WoSP5UNi6QzmMfWFSRUSJx0vKcR683W2SEu3RTRa74OOfzBk
tDSdRMpieWAjvrC6nwnnsjiWkFMAJPjXF3lbPyM8yQmvlFqfRmZRGQ90Xv0MCzbibjaFhpYzEjAh
D4zbwSxtiDkmFma8l8np2DJffC+UAmHYPsQUADOM5zgfvCy5L8UYocy5ZDkl+3jl+vWwqXOyhjSZ
LRflYsiQ/d8JLm6dmZTDUj0hkS96RJ8vqrYTKcyD9dXEyfq3zTlQbS5+YOPiyQW44ga6y6S42x2A
JXUFinmNht1KJWwqcAMC9/2Jz3i1TYy86QWUfBiI+WaL1yNXywRKh0eRm0wFEj35kij5hqWPiZ8B
vQXJVWXviDD0MXC33cxgWE/68xjKsBlbrUy5AZSnUOrvoFW+GB3Ik8Vs2sM03q3gksumfq/0WYAz
9+f/S6BVe7nACNQBB7/E1bqU8ztysD8a3Evtbjqiata0Ygt221zA57aytW0eUOH3uVYKD3QZwMxh
hGTV3qXj0NR1ZKiiRLq13VpvnEBz0IMl/Mycgmg6N3zGki8RXogbc/2+4nJ5VKTDJ8ez70yz5trM
XH0ZOQ3SAoAXQbK6D5w6TZByf9g4X/VygSpLHNyyr4d466KB7I3PziG4zGOvkXoxz60JpsHy4tMI
S906dJbpgU+mUX3MtAuvgHGvc3U8haOr8UQF7jgW/Iy3pHN03kTiswqSm/hEo98nsWNLkNdlxuOi
ZzR/Mj7IuhsvLXJVfNlwMLgCxVvcD9mxXsXMDgvQ0GgA353nuiGmE1dYRBb0NSJuzOxd7Q1FjFWx
927MwShC8rk7gvZH1eCnOy0nsEsWY4gQsW4tyNRGz2xmjlMrDgTPVvG+j2QmHokdH7XhxTYU0WKi
lGoYZsnlY/Yv5040JsEeMldQfTRhqI9CSxjaldECMPjuq8Hw6rRFgy0mRYgcqPywGqMoYX6NqeeU
XuERNxlbHARBTgnZ06GhuXwTtQYp+x3fTZjErm6KVC7QZc+VVasJKXqK+m2y11RJNxaxoFuLu9gh
mvKwgNfeYfvZuGa4nPUdshjudl8Pm9HoSAUxxk5ZwOmt3zQ33uLDsSFoIkxm1QWe5bwMHdwW2SCO
Q6MrMTu+sqthcMjCA0IanBMli+tPh1XvcPVSyNGajf+ILqysopCwX0g/oIcdKMdBJIy3LInnRyPy
tgGeBVv2TFakQLDOSkOiktlPgVLX8gIWV3uezHa4Qw4XPbk/VHlBXRkeFeON
`protect end_protected
