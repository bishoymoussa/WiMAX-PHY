-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
yOtEyHo3ra4j/E65kBKbbeKfUuSoMmifjhbLg3IhntHsXJtTKnWTx/6XSMRbQlqVnz16hPLed9zm
KMDybJAXyHUUSY+mSf2T201TcMyMfs9fTkB4V8jz9V4spvG5DS099Xi4iOTDZbg4seAo03Mj0LH/
SCRgRX3mviQf0BPMaAHdxz0HHFK4zt/9DsLL+64InWb0VCrogpFK5tBge5TMnbF575dx3OXLdMPq
+h7JMFZgpjGa/H7AtXFYkjdDRfkgekIDLMeqWOKPEKkUWNqL2ZvOe7X7zu6IYkmhQxfpIDDRk8ZZ
zWFvrLkU6YTpsV3rjmeAjkRhHWt2CtiAenRQDw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5280)
`protect data_block
4U5rvI4bGDqNqfYzSLopenELpyaOyGXda5LMzogtUpuu5b+Upuz5vlfPV7W8QnLLM21ROgbTGgOf
yvg165is3Ndcaw4kpePijZL9t6KrwBE4YRZKusoLqWB7+xGyrAmTy8PhFpyuTaJcEOvb5fEwZaSi
vfIYogj59Svh/MI7cTEv8TpWGVx8PCSbwFpqaGq5ftwiDSmU3jycE2l05xFxXDSBPHnDAq/nWfH0
dW5+VvIW1/TCwjWjYD11wv2zIt8aXpXfeNgQwYJSUNLvRieMJCBqqLw4P3qxSsJNvp4pjUWNndT5
zbbE2Y1N8VsYzpaXYy7MMOPaD4uC8W33h9vk2eKIxP4UAvUYYNrL3D8Pp7Y9Z2NeZRZlvfg93ymc
8Z5bGpmo/2lpZEctktrMyVX0ydbHqTejNM+NnY9AJwVSdZo6oG9sfvdEyDwM4PAyp0tENOWd2Mz0
hK7ralk2THwev76WD7pAnNpiekhw+7g3KyYoKdDn7IOy0qpMBxEZrbO9I21gT2bdlkiK44rI7dsO
fJhZCeKt4OxYAo5Va4MBykrDSiKFarpNMrN53KVw+1Rp+Y3yDF+fDb4A6EVis92XuXyJMzCiN3Ex
rU92JuI1OxPEDr7gn1AZqNiXoQ+ONo3TczEKztWmKMzaWPZmQkMiuspTedGXnQgmXEhAl18mMDqA
/WIoEI9qoUdPnOEx6iLDJ8rqi39rHsAGkOY12RsWDWtJ67WAgdmds3eZ2XeVPcjbcO2ODXymTmap
qsviUmmt30nwXXvlaEw/LOu7/M2Y7Y2iG/piKuQ+2OXmEBw6nrQ/nDU1RCSuOq9wWjBujL18fw77
wrKL+XkZx+vsXtjWBWMlIrm/E/uWZeGghRe8Cop+J8PB2nE6K4Z/pCu8wABi8e+z2H5SZTmBbrp9
ZAnsseI0e2m7aPEfXOBzgAf7dhlWaGLXOl6QZMM2sg6gofOQAcQW/YC/Tp/BFZk+uVZbK1DYkTLN
e4fwm7GbcBT+knV/kQWTXaTdxNjegxOBXWsO4p+JnA3IWSke6upMwx1wqq92fw9Vcg0W7GxDP0kh
7v5cRvW74+y+DNly1d6ZvkyQrehl6lvhAIAOyt+ETrjlSv4UH7XaPjrmXNStfZ0EVxmjdjcugl1n
xz8itMiBTx5Xti8JuRSdW/FXxlFZnDy5ZgiyiD5DLehgdvaht60ov9Idqs33rpAnFhNyNVgxJSak
+5ZtRE6Wq/JePn1SE1Q1DKpxrxtRSIQ3yNjkIHtKCxxM4nRcHl7wiwGFO5wa9BYuVIVMQ0fCMqgH
9SdaznPqd/4KCtuqWFZh3f3BKAy3/93fK6Bdn6pSztUamp3E2btG5j830RlWiuSvhYGg/wEgMM6N
UnsfncqKHpl9s4Yrq4+qUtvv2FXrFNhKKN/kz5ZHfwskGqYefQkuk+OmvX20qB2Oy5n/yPlfdBg4
rDo8cxPABvYqHh7PBowJiZB5I5C/FKr8suQdLCRRbCHjw5PUD/iiGepygO1HhPI2yl5L/3Ktbhto
uFDB2d83IJ+dO9jAqrmjwBjGH2cmU24V7v0H+g6rEdzbO+jAHNgsMGn6qmA97kcWYsN6/KYgBhQe
EYFCLql6jnvMdlVfeem3XSGwP1Lq132lp5PAnbyW0yGR2agwZHvn7R18i2aboIHDAZA0kU+Lv3ab
l3XtUEru14RupO5A1dXvNhlb0dnhTbKowO9fzRNDCzKd934C9XBXbp3PIMtjMXe3ghj8UZ3msj0H
/ie83+ZDOMOct8yMkn9Dt0YViFPhTLa51apD7vh7XkGWlgSuB+sitviVIn3JoM0VakoQRP6tC653
cuUdnqH1jLywN3/1JL/PQU1WnDE3utEuRo9nJailB/Z5IElOqsOcLEYLiHd3hIDlxNEQ4JYPVAjZ
JqdgTpJgq4HEjA21yYETGAGh9SaQjLhjO5144koJy45fK/UXkHnzFom2sAY/BZ2pYprFlsRaeQ0j
+RZ+NAHt6ot4MIhsfTl/ha49ALPZhX/mMYfV9ds8xc/OpiQqWtftAIM4U74HthVNEdSg0FhEQ4kb
v9x15T9/x9n2aBQkbzVWIHrisrxfWVHPyQnfC0b73IqLjmo2I8A4tKi91wBNNCM/rxamtWCA/YIK
nysWeOVTrBfnUi0CPk4g1HYOX5njeFfaUkizH7vC52htJkIsHFOlbBNq7sQZ5Hgui6dWyRYfg/Ux
DCzHxV4z0bJwXGO2SwMVDV5dfhjoZ/yPH+onHodN9FbMEhHBXXkUnNHsxUBug+9XszHB+pNFzosP
EZM8b6oy3tbLNs5aMLxvPJebF5bOgC+72xeA3SlOZ63FqBHOCYvbNmTC9G2rPnYc40q8fQ0IV3IX
WWNju7cssn2J1bsrMQGndNXUhLMq1m3NwEfPWoF+aR/cXZjnIEyFgJx5j6EeuSRMgipaTWSyM3gl
TWaGPm8xAqfYvuprJYpR884l7X4+c1rL+iNO4Fo5LW5JNQXOV92dFP5BePkAI04DX5Rn55Btck3L
+QrZVwoX9IMJbKWxuHH+hU24xDe27lF3Oq0AqPFPW7UggeOslNvN/DrLSZKXhKgiaLcfGi96x3NC
yxS6yatoNvgaxFrTwFf+FX4/khyMzLUWohgZr4QGIKMgGihA7fvKVROfnAuc7SX8S7gWwlDAURqN
pCLxnVnu8HzoW6fF6qVMCD6+80airfzoBaefjAI0ZJhUjm0wghU1Gt9Wjfcc3RernkCHdWzPkZ6n
ZhPPF4Ie7ZhUyRdShjHBbYURs5rUTCkDFdSZR7wF3YxXxPTdwha37D2ihxc1IELL0kZKtMiwpkFT
LluRZOwtCj+OO07SPDbW0CP3MFFyC8zuZNh29vZy4NW/jwhsqMHTgOUHCqblLFMdw7vaG3QzncFe
3+ZQ6WXkUYRdp48qRsW/a1YGC3ufW/BUFT+Qgojjmdn1Nmp2++9rHAZROU80w1JNxxfXBYMxRleU
nZjScbZyHzdeBVpBM/z3q+BqbP1BfyRfQOujvWEkbZfx+WXhw5IjugwQ2sYN6SaHKmlqbdcmiffa
3TuWCoGzwERWO56COs8V825eT9V6Hu03cYy8gtLf6/0Eb706+gbJaM3AXfUy7CsUSEDj0DZ1n/fU
e74Yk4kMBPEgG9G1g/I5Gf47vZBOwxxyJXvJy+RMxYSMBbfNTuzXhT+uXJXhXUmeKTQgj/3yfON7
5Q1H6/RI2meGqhF9wVfAY8w8DTbVaJNg5obg5NTsJMhnvmJdCSgi2hUNrAgw2rEFTdHE4qYCERxX
XcN3rBnKoycgNH8R2dZXvdYZ4Wg7Hk2MJ8ULZOtNGRbzSkgiE66FZ7C5ilfuHVeh5ubO9con8eNk
To0mnqVpGAYNmP0mVm/GDw2z/xoXyKgy+55zB8fAwL759ercG5dZBnWhkh1tZU5hogh9Y/SjSvC9
u0b6MtPH+Fl+2Pv8kY6C4KQUiY9uighpw0qEtN2eeyw/d/YPfK7vowvPZ1zxw1lsZgwBRSDY6esV
E/NykOMZhwZyvCZM++y5avwwWNfP3+u0GTVT7J3USXfVDPVto736CezZbaKFSLNYZhguXJIxG7hf
lP4TeoosDUD5B20P3186rymK+ago4I/EbLfqC9OgTcbwWTtaGRMvg4NewWndPY2oAgaGdSGelbOY
6Fh+k9N3UBSL5F4VQiTVA4X06r+DUSz7xkKHfkWwS2p67upaw29hzeZQw8VPWWSEYfN2run7NOXE
oCTipbDqgZFWGAbvY6OyPlrZ4Btm14DqlFmVURz+WMe9+15FPBVGnxf4SdmkwRT1Jw+VMK0BVi9f
V3kyDCKGy4SBwJ2PoqrmJXho8lDj+NyLdwF72dcsR/XvZFrQ+9jEc9JoPhI1Ng+HCNFknpmQtt3N
/3P7qn4RlZsADkd7d4L/vvd0UkDzHaAIxwxLWlqkolP+OrA/kllcfl/+sFVmN2oNvnIgpC7NE2K+
K3khe7qgwz6uM/RP8O58KSplzTzwwoiNImjGJMiUxgHQjKSjdKlhbgChoCljQRKUWh730RpCnhCV
XAvqzDvbZif5D8Yu7xZFgb0bNJqQWDPUFsX0nTvt3rkyp20JUo+mpKOZQ0zRzj2mAmgplDREsWe/
+/ioZMFF+P/hE6kSaP+SrVZzKKDh0MfjR8QDIZ1VteAm51onKRjg/9oWiCMqTjSFfX1QWnRyDnJL
1kDa7NQZXD+Q4oR+6j9ZCC0rPfAETM7dKxO7K+n9pCg7sc6KJoOl/mHnT/1jLBrzoNY5fAqGeB21
Vc+FsIOmCydsd6ZVNvxoJrsrlhQSjYupZP3doX+dB32zK0AS39LnaGFMgg0VKr1cn8NbddcqnbAo
H8qNKx6ZUfzV0Av2Y4B1zjZXvV7ycBgG2XZagqWGHqd5gqfEfxE5IbIB7+F/DF3076jEOpzRzZth
hnmUt9HQseX0zZf0p96Du8/VWFN8fwDHW7LT15X6BgO2GPNl2vZ7NqaHPrW4zvSDzrsHBeJYj23A
IKaAmPb9SpHW9g14JKxqq6r92hk1Y+9KromSHrd4tmy6ESxikqcd72ttSLDlTl82uynL+Rrjgi2m
ovJkmpN3Dl2BEtGQcRgwgZ7KqsD30P03jEOIzxoRkpdme9AtiO7R4H9KEW3TijndhKmuSjFwBt23
42HPS36446wNBUd58snLkpqOukKqDX+M+pyO/5OhKoC0BANPWTGfvZ5oYfREv32tCifm0+DOoQ0K
L311oDt5im8FVUaeYYkTZKgTMv0WUNFQYPpKa7WMdS4fue3ebMlP7KakxGY3Q2NPBsfrSqOYMaOO
XftGmH5N3LzXsje0ly/iIQv52flx3ToV9RspkNXD/+GstSeFiaDd50bzjtKq/u11wr0+jJJz0m/5
WnpmlfD5dflP4gfKdGRzaSEgQYa+0wRywXVS09ERJNNw1bMAMih99v1HkOxfhTi+gHCge3VwBvfz
2IUl+br90MVuX0qvYQujZKtYHJsHXLBa2Lhz1aQSSwMEeYcXA7FFOPPN+B7fEJ4a8n+8zYaRsm/7
BLh7R6zmpk6WwT2+9eAufXJauVenoQAEBRphggqHQTKFK3kS3yAVn8xpa3POIxpMoyb7ff29ymuI
sAT22OSeA5xQE0BfhakbYCNIrLWrOfhNPJBhQwowzVZM+3bQP89qJdzJEkAsxy3oRHiXsi1oaeX2
dRQJP7BVlg6F8MVpdTu5GrcXU544tf5C8OhqB8RWwqTRd2PuxXJtdVdUvPfy+ypuuRUmlvkIJbXh
/0eTSD4NFs8oQX/oVrR694VLtnmoRVuBXwigvb8ChPDdA1Uy/0mc6Roigv4S1eE7csTr7Q9obSZF
A6bbrLutU4r/nI+Hm2xxBFAWXWrwI8MT1rT42DZo2n7+spGWvZYH2YsZrCVYN8Nbij0l/56ZRpYV
Ae5MMK6Kk7S3MPtS4mC+IuHUhS/qeVpqapp3dLO7cFKRlftz94pcnDj3Vyku8/SQ4qjEKCTKs/oY
JDp3KkfV5x5VGe1g8Om+aAPzA+hvHsKNh8RvYTLDy2IAvIthqsrmCvUFFJxPtFuvrn1NQyHSbm6o
935tupydhoAq/L+SngVFIg5+ZMaoXJvn89naoAgmL7kj+JtbF9/eudbJCyGpFb4YiMtR59N+z7aU
2/sobqrOkUlFXjPp9/WOtUmS2K4isHQan7ellBrewQPykZErQ6Efdo+JTraQ6ZNvznWbB6mB1f/n
c4ZGQt8rHeKrDueNOPNJ3CmVZOyllSayYQOJsGUVDV3dlv5XuHNWLaatuoF/nLBmE0GqJSVClL7h
v97BJhIruv+raXWq6E0NZQ+Ff0Y6rxN80QMpsVYJ3m8VqRSJDOpwQwEbvPLSJeJFBjDs4GrCNGQE
o0vTe6kzO5rmGu1Qt8kPm1Sz/Tbs0JFQqibSIbmpQwwWd4NRqzPAY3ws7340Voflej5clrsXM8Ww
5ZNZzosW1FvG1avO1DLSoymEj/EpSqIoKrsCCmxIPtA6rGT6dZVO4UOYvLCKt5lRPbsc7VRT2F1u
vlVkEh71hgyW7k2qp6Fu12FQE6RT/pfM/GQwpcj+P+KF9kwyG/3TWTPPXWdWxaCqrNP9BcbIZRFY
8WMZmPHZ/tASza593E++Bl6f6NK0U1Y8+8/1VAYsbWVu3lybUbHCiCUUYpm8PVoGZzCmj6PWpiNL
UF0X5yBI/8sb4C4Ji0Jf7IAEtME2+Ku+BTz7fzdEVT4QJO7k/Y8PSY313qoBDNVdBz14tgLKQeqc
U6BorjZJ56xvJ9lCBWQ8Qz7mqqesRw/gAzcXRLtoEZ1gXkM8LGkTTTEuMEoPikvAalJJ62C0bZpk
A6RH+9YzoNHC0RBloFY3zAQytSWrTF9EQBhLfXzczbfhCAJXSYzZivbQApTfLPviplr+t4vNvtWq
bB63gjdoDgMqVRHCMC95HxeXuh1kXnj7U70uAkdbLpnWCa+DipeMSv2QUGDvqt/rwqo4Zxmpv2VL
ECC8kOjciw40SU/0H3J35l9iNJ3yfm1t3E91AsdUKwFwUlsc78ARHKgivoy/qIPl8XarbyGcGAPC
CWki2wjFSIBejzDCMA/Ni0tR+iI2Y8v3Z4h4KpHvnScah/Fej5oHBSPyu6xjkAkuU2nFpmPPQh4M
dKJsD/lFq+jBxmtq90QAZUmmB2ZebnWkzzbJOmozIGZfJuSzWpjSJKSgwhQNHPwoAzZrmPqEdFF0
aomLuRvit86jouQopNWkrueRHo0LOEpYzrpMh74PvEDHQbeMj20uTdLLhC7JQW0OR6MQ1zmiOo+P
n6G4WF9X02DRUWuQkqV+9qb4ZsWJnYCax8t0XA+X9Dkw6bwxsl0zmcEvs/axKTyXcnWHxwTNBxIe
k/ZG69KVt768CKsaLtLSEah9gKdMFcw2s8kUaes1U1ALquYXndU4kUvT+pikfQ+LMCdAtHX1ox4X
6i1BMAFZ//4iIPVXX/ejGW3/XNBbnLkvpQbNjtNk+6Fx91ScHrZJNnfBjgprP8+8/r1h3nbW0bdn
832l5PYoBQqktchMjoqMJ7cQ575huvw+NDx2Emo2mi5uSpMy
`protect end_protected
