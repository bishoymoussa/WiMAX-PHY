-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Cs+OM4zl1MOAkHNWF+Mh3Zr6dYh79EVpGAXobiipPDNEFT7tGySfVuxsjhR0tZ6AN1gouDbEQUQQ
pHNvm8aVwjWu4PpFjeY6pfBV/GBINrIlM219rD0xoRu/JgODuGVTVh3sCxn9fSHUCrMLwAvnSVVJ
R89mrhlcs/in96QiZNezgqQ4EYDPv/AuXiHnJ3a3TICtByC/YB2jrSapTeTXkGttQAz2DW0DcaQL
rGW6dDhyoCAloKbZQtOmVDyxRGcnP1N6UQM38w05smvnItctQK0vL/RoIHlqLLj/C5GkFi7v1Cq5
QitJ0UoNPRx8rtSHUrh7vzw5LLdzu0VmqIX10g==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4672)
`protect data_block
/vMTFgT2U6LLODuSei+Jv9aND8afYHQL/y2q1EN7gPB795WKlZP1cwBoGF7pmeKJT1TQUCwcUrOt
aw7O2OB/fXv/m7FCVmrovVm2mmphEDs/I2fv9HbjyqXUtRFM9Aa/B96M/j/sypn2F6p7PzanoemT
1LF6RUgLRMGT8Yau+alySQHaa75TvtRG1ot43rs0daNtWY1GsET/gGozMK4CO1kl14YdktGK+w06
L4vLsNvcQdNV1jLzhBOBvdbPMRGTcUMGmK37gj3RDKuJU0Th45KFsO2hiHFS09xR1xAyXfR0HAG1
Yyn+mLVXSz1TVPyHpLKYsRpBMmhxO9UXEO03NvpHbY0eUmf+vJtixt5av7wfolud05y8uphr1Q89
ZchJpOncFbaRI0FH+LwLthnGrIMJWOGTs+mdKl89x5wFM4vTBXA9SOFgwAvXjjWoUDgqS/fmjXZc
bvfYE6KB93IyrfufFO2lLjkExPKq7ArwBg12lTEd4LhP/3rax3amD6lscPXzoZMnhiaFJPNgtruB
R2w/wdyZB1GUZMRTEQfqCbksjahdUKmevB5Q4X7xrrFTTChyc8U94+DLKfYFr66kpY/Yd0BGGj99
zqOjrtJUdnwM9vGc8NaNsXWMh77E84UvYg1qbx85cB7nT0NJE96oH9KtzJ8iuAWxCNPb3t/jCj+R
PrV5U9n+seqYDBTsWaWpPwO0WVU5lGNNn7UYcVTLo3jQUtQDMcAD0V8VahJD2d1eQxwFi/bVow2f
jnCKKzGD+7CMDdONCCKPx/mnh+yUUAw9V3tQyW41vWsQV3LVbCY/5ujWlY4wtaaIMqRfIjbof2lq
lgky7SDrxecN+vWfO7TAgpOltkCj2YVky5YGN0MAX2RblLIbRS8t7ZEbAc/PHkU5IqBrPwe8LnH5
PpMeceuIlXUBvlKntuFPcaVr3hgf8Fkjv+RhZbiHEjv3qeNetKriDT9+PKp3AyMEh6HJ+AQxQKck
R8xL7A3Z/wncC6T3MoDDVyOPmEHYnE3vi3MJD4jUzw8xICuAxyosvwAFjVfPj6sc4F0U9jswVAsU
tbQXkc6D9l1fuy20rDPFA1gzdYUGEQwZzI5vvTboFL1Q271M/j3RrOK8q7KgDemaV6EZkmXnpoS1
ObpNuNvsEtvD7HFWg/BJeDDlwsn5DVK2MzRpR6X+nKLoSIy6Wn5zVrliPCqNoo1TkpmB/9RdoNS1
DaAHeJUlrcvFjANvY6iWP17Eosgz0DPP4iqfzxHm82JCifTVg7fGYoIxQaAHWuXJ304sGJlBRO3A
agK1Lxn/vzi8eFXWjAuheGKuhm10ArJF937ZMoEoTMIxQtUC0kCsIKtlOyy0mSdkOE6nEdsHdVo1
uGpGL2E0yGSO6NHs4qzrT33kvRrRWcSyJWxvUEbS3EV96O9Vp5/5mKTukrNN0E+M6TmMvE6Y1Gf0
fzOcorh6K8ZK/OxrCSYUSG35AomOtmWkX7JkRPHp9/Jev4bPm4g+q6XchlTwq6qO5zh0v0aB5Qqr
t3Dy7mF/X8WXWh8c3FXXQ9cx+PEjMENRnqCbo7Cc7to3ke1t7k0vjZ6efg+0zPovWvlzAWADAIEE
g8+7CFexDulIK1a06DIP1Yzv8d1CrSvVmvc/aX8+fRL/1XvdH/sEMA8KV4BEKgdRqxu7Exsd7dIf
PD5w/QLEEQUuDEa2PQmr9wJCP8p85IwBTgqkA3kxnmse6jkzV8ZJhrRy2QBmK6oditdMIZC49bmr
GaXJGzDOFrIxNpYE3Kl9KuyMBIBEz0N5tRC4rs3/buhVpvy3dRGiFFe4stcWwztu0NXxH8QxcBEn
jIdVT2ApX6XyB06fSYAIfulRx0OdFeJpCQXadFxqNzs/3oOQQGx9aKCptOzZFrnX84QhTUe2unIl
kGrBxfIjUVDqk6Ubbw6/jydLSIPDFdybrjG11pPkqB7QZK3FHKPjiHUw9wsmFU/WETqdxivB7O+z
0mdknJLH/H9zIgh6BmHGcwPeJSvxYOjCAvCz0FWdwKJQdh6qf8tQZFfEtOvLrrN+syPQzEoYchoG
DUirF4KYOcqcaXwwYYfbZXU0Db/uU5vvXlGac5gOwKdLsUXm2sxyKKXwtF4QqIKwLlDYyawSp5Sk
OS8BO5RrdQCiZvhFevFebRbB32dYaIBYnPjsjyYfQBF4of7GUtMQyiibgfWQWH0EMrFoL+sfgOvT
um7HI83Tun9T8ir74uD3gxyti+IEyf/BkZzejLcF/zJsSiDI5cQsDC+YzMi54AAvx+XnqV5sxH2H
jqsiHSGXNV353Z6ZRMhyq/vNwJbIiC7PKAWxcYZDOQYdU9bUJYHML+Fe73aQrFUsHUNNto2I7MgS
AbtKRuPPBLv8tzpKSMc+Cu+O6q7R+H4Vqtc0Td+tKCI4ob+AwF5tV+1vYaxEleibDrp+WTtQmK/C
zZvD3I9A4HMa8+H/fv50Oqs0axQhAXnD4tv9yw+L32jXLH0EF8GMmwJvlH5K5y+YrNy0GPiv34SZ
hESb/RAik6y2VQT7bbV/7f549/HC1PRVhkInjMLcIPeqFrXKwxmmz3vnFm9xHMTX6ENkwwIHH0EU
MgQe0PtkFTIBHb29LLbIwb6M/EzHfRJX77tSfPbs74w3Ln2z8sMojHdNdsxp5BoRFfckfLKaf3Iv
TTTAVMYFclKIL59/U+dsRBVdeUI72Gm3GHFQxG9Mhl5iqUytRE0HAoXKRVLAAdPhHlqiaObS2xxD
oIj9miu+Sva4hAV7NUytuJgJ6nPicahcYSfCfnRVuqkcPOB74TaqTwkUR66ARNSZcqq0ZWmaF4eE
VLWbkWgxPD2SWsQBGaacjKtF7pMyT6QGd/e7jkr0uGXO/1uzUc18vGg8nrRwAsUR7KSfqekA7n9j
mEZQ/6pcO24bi4hYwhtDrjEotmJKMIa/TL3EAAjkwNDiI2aQWZm29pZkkPKQ3bTfYdZjHZz1oSHC
xeiakJijtIZIxxhvtK0DFeCACqljYSJIqHVfnHcg2pqsqFUY1vD/Ctw8NtLxC8wjpvu3T7ddVn1w
qnTZIOfqzR6VM7w0LDVT6K/M6Giecd/QooXm4gfx3LJTpzymQHUHH9SsUusp3HD0Gfvw54CTcGy0
VmmRPN81WtEPxi1Kum1NvxyImBcZNa2v7MVN+kHv08M7zR1lESh/Xoupg/o9/uAiFDiMeDwfj4NN
uEK0cjKWWVB8DKIH4eITqNSs7w6WeU13SgG3aCayqp/r6xJm1Fx/KrW7o0yBysLJIqZe7FRfF1Lh
5yyUAyX+vZDzqt0BXYnMKYbB03bQDpn13BR7dYZgWbcdW7PKBnmmgRC4BDhFf/preVQmKPKcHkTI
L7jINfgc+mGLJ3ONhf7LuAvpJ1PhT93/wJqncu7aYMYHh+//Fui9vB7GliNjIscDmv5HDFbyr1t2
lsAkn20F9FNoPlUMu8kM03rX/8dVWYhIULgW9z17rdgbH+O/U92aI90dGode5pacRuDwWcilMDT3
GhgE3UnZCi+dBg9ZieU2UyBxCtJN+Ci63sgWwApFvkpbwh1SapagQfDd1nAl6l5cq0S2PevXS1Yb
5h8VduNiu9mN+zcFy0FKUNibr0BXCnO4GVa0d6R/H+fb4kmMydByNswDGepwaDgbO1P8JUtOiInv
UPstgsTVItpCq8JjV/NNYGVsT6JBRcr+ZiNu2g8SduFqDktmo3F3R7UMs2ZbiT+rjKNfMTimFJ+w
nWxKwOAaVShckvs7C0eMQv+mQapegF3PbVwKvxydAcXQIBR1I/62apaG0c7+oe2IlFmv38w6aZXV
xS6u+r7gaOfgcZeqZRF8SsvcBOs44L/eP1tcN2xKYk3gWGHQt6NWLpc4qnzZaN4r3Rg+Dc04hP7E
+g32JhxySgBfXUBUvvV7K25qhmT/JEeXZcDpC3tKbtk9ZhNLXdizWjjkHJWMBlbK54r63D75jtZS
fhwl6NVs2SkRN/HPZujLujq3t81YbVSpv8QgcdKTqDUfc3YIkaCxsemyXpGw7oQagSzCqr5YWhqi
6NvZ0kAE4OzSPvbUGRj8mi7VVbzpxpIzL34y+4uE7+W1ENhRMJounXDsu+ce47MMyCIa62FuFCt8
oyuOhTnYJnscTS2sxKkk/Yqe1Apj7HTETOT+6Ayh8aT10+zxoOVyUCeaDUUh7BPSoxrPSUuCNxlt
xPO6DNvX5s9H/8/icsw9bj2A1qkGWoB65JsSiRd7Js0dtg+6sS2/Io7CgW32zGKB97kMTq247hxP
5g1P4Ul0nEHi/Bkr6Rw34BW7frgLj9KKTP/SziSgEnY2gaWfdSpAhuNKqCDJjlRvaP3J5I9a+JhO
OF9UpPGy8GKqYFNKdfCzeL0KroKdq3+fjA25AhnP+IPqj0LKF+8vKPkuX2eZmCui1OQSKUQhSqMA
+Sv6mbkKspG8ENf74h4f+lzCkfGLPjimQ5q6Yqv1GGe5mWzZUZ2fk9Qz6ciLu6mJZK/fNJH6zwni
Lxvse0nP2uNc7IQOuVm1nsJqlezVxbL3yweuPTRJ0gg9ZEWurabxT7rvO2XZU92ev81WKyser4La
7howb63ctTwQRGi9gxSrCGM3v4jaXndh/FupqxHOCO1DLMZgVhHOxMDIM1pl1365x4Kp6VMbbKbL
3ab0TaQMO9XjTjNyVwmEvSnJBMGSkDJwhuP2/Y+FWgiPSPb3Z4FcHKiF+cFwlvA9Dy7npiY4ZwKM
j9rqyKn26rZxWSJqyfHIMZA9r4uS7nKVjezSlnOG8zDsz6cAzKb7873x2bEJeFSZlLUCZLu+YHwH
3hPVsfXFWoOtZe6E9F0KWmgkWexK4a0L6LrW1ZkGdHoKTKUekQeB7U2F8Vx6UN1It6T18TbER7am
XLcRBKOvFZYs5LFeGA/hTupUUXqP28jHgBQvNETBheSCmLoSgdme9L7iWwTicw45uV/DxPSAlQ8w
0wy7yKjHuEFDyTd2y7aLrOW4UcnAybl2PT40j4o9rBg4F+TDnMcSSG5zZl5DwqggY5YowBuuSuaJ
YbrhxAvqkEK86udeqfFgTXAUJUsQsJ4EfjkvG3HORdUIdm0nGeod3+T0owPHLbAANTVRhkWoT04A
5QxArkea0K9vZxBidMhB8NpT76ppo1uBz7fu/SZHpRwhUBsUhN2uXvGxYMNbDP+l0jArwh6RqSBt
wNf84ReuNG5yEnSx9h4V2MEneTj1jgUBUEwm4+unBzj2e9o2HFvO8GiM8rYziBaoyrwSY99E+uOO
QbT2YLPmfjjZ2BneOLQDO3bfa1re0V1A6W4CDVm7vNm6B9dX2ssRLW1baASpmAOl9TXw4IfHa8E+
QBQPUcoaiU5T3yZiZMaPqgDIarLKmzkfeprheoGSgWVaqBAvDO+R/pLVVzJ+5m0rA6Ld32829kji
ygw+9UHFL4r8kqtzktjZK+KmdIvuJJXqe7rQLGDszRKA6I7RjE+tJOVW96rTKPc+igys8Of/mqZA
z99qgDorL4S5lLTnzR8m1mTy5r4B2s7lJCae3Fa+X9g/h0XvKNhGUkkwRKmcAdc91/uXfmBtlJvS
MATK/NUSGrwW2APOeEIqs4/n8NqgYEvnIfuksYmAaSb7qkVHbHWn8/OjbtDtIZEtpBJ791zbp4GV
cNx6uH+AR1avwVsi4OdfsUHl4YJ3L5gO49omS0OZIwuwb2Aw40gQeIrifg3YTKNTNF1mWokJfe4q
OudIvC++kawgxi9fvbtEk65jdovkwa4wU9D+EPvjpOso2kBpHfg3PdL9aPxuJy7vZn49zrs1ivZ2
6zPFj7L7y1LHwGI6tvsAkUb4t1AL6LS6mfSONcLicJ9NPheVHjzZ6omdfFvFn9WSffl65KSxKggW
PXhPSP9ckOlYbS9c8UABKYe/HkXbBJcBOlInQUkrPc4MdhjSNwEKtVx3Wf81LtUxHtWbf6o/UK/Z
TmZFgv59F0pxAGpCk7GKOrA50EanHaVekV4ZGonScwVMR7QY0ik4Htitga3WPqfM7ev1XoqE6WYx
D5V6tZdzIVaNrXPOdqEJhp25PRVSC4bX8u5u3tVOVXdB1QenlvRXow3hoxOd9PFbzMAApH7YI5Ul
xBEgAM4brAcIhmNCNT6DI/G2RefMsSv9w4FNhfMazkIxxlPFbcr9D62G9WOI8+o1Mkb+KO1jcfhq
u+a+qcTwb3dXaxlN+ASjjxp+EnvpJCULEafdvQ/gbnFUo9oJN+RitrrMAw3HnwL4SclaVKtLyg==
`protect end_protected
