-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
QSBdksr+8hAtAmqXcAgK8BplVq8GbbPKaJNSul+db7I+68zjsQJNnINOqhsN5V13eG6tCir9NI5j
0fumv4NMeYbMsRKlg/7YyezGFVcGBBX/o3bD7G6gtAE6U2ylfcodPxb0Tm17rGK+UY+PB3XoxWwH
XVdV0QUdH1L9otYE2+/Uwnh3ss6ICwvWLIdziAszmT95CkVgCsrxysnRlMf5nS6meym3u7a7hzW/
lxIoKVcfgu5Wg/T/IXapWNSPn69rOVpKxugTQS7xkxb75c9s4b7kE5BNikacmKIV71pcNDTT2Wzg
beeTr0sxBTj9/u9pHQUTYBESBPpWi+AyUVjnfg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 30288)
`protect data_block
S/pfHxO0IlrtceIrfXSyeKa6ThAGc4sWgjxqJCXQreMFybOUkxt2qildbOMsVvzCq75EWUZsFrEO
tNVtA5nYkg7+x4zUGcg4tvWTBBdNV8MVkgDM0eRAMKhKKj8UVH4dRJ8mAxEIkLUoejdPInQeOEnQ
JeJrMDCelrGsY+77QMFPImutGAqvcdIEWH5hAXapI4y8nDq/UWUvro4wI8BsA1QniZ8VLP/tvLOx
FqOpCcTiaEkhaHJZb5GUh/Twu9JMCZavc2BqC0i8uypUT4x45QYYBZzzcdz0fbNhEHp4GOMqRzk7
OtoKwvK6WBG2/OSVE4nGFNjGZeEVO8su9Ku/w529n8XFl++KnaXDi6nebGbUU+QjGdynnV+38+6H
wni4PMCW9C7XE1BdL65rFGMQ0gk7wf4nUnFMwRePcfttltvItlJxbvA3ynzoxN33mIuCXnfaC6Bs
hYXf3aYf+H9R6I1mzZBoqZtsqXNhmdloxFFymk5oaZcLKlNfWL2H+gumeaNBdny0hifLXkAF1Dvh
XJargIUYB5/dLLSWKCMq2jnl8rFYjK2/3yruxgoYsazWkgWdeTtlBeZdRXkkkQ8Xn5ZSlUixnmDl
slB9mojb+sV1MbNLpDs0P199nM0i9mForpwS4CXXzxjoaGq6gM827g5p/HzI+urEP0S6JOL5RRxg
QZNER24kfc7iv8EHoVfE99C/YfLsb1lWPnCWcdI05OU+dkWIeCAAUK5KNxv3WQDBa9WgbNv/NjNd
h4txclttYIYyEMESynLMW7ir1Laq0HVkp09TcH5TMLx3anPO5Hg0hILH29TfGBdU1E1DbioCPoyZ
AKg4y4E8NoZMjTUmEQCiym+ScuaTIJlby7cWyzcBzS/aO+YfAn0sHevUmSezO/g6lMMfbVlknUMz
PduP6F5497nCQpAsinRMjx5+LfqkVsXR9THFASHin1N0rH81uZshjwP9k/ivv3v/1tNAZnorhbVM
1l5QiVdL3wNKHYNcng6HtBeplaWKiySJf3giBhgH82YxZYoU/Fw8htJVHT0UNJNe0eEP9dAiuvuW
D4Kweas+f59zN6NSVZbLoaYjpVNXqP0oA1e6GEQLesvmvwiUcV53Hf+SWKzkgffmXGNghI8YADsz
FSfrxV9HK2Sl/szhg5nUFXIebcbKPWny8lyOYlUwb8nMoDxOss/3MGL6qexrm3che1m+gTcfid+N
+0guIS/1JHb8zwH1zxblMh94NvThCSfmMf4/dQS9t4gTIjYtBrjFOzI3aR8irTCQtpGK/hhqvbAB
/oZliAzDTenE7D/yACnUMdXFFH8mSV+PGqeHoedoLbWfJ5pF4jA0WXCFRUt4WH1aEXzg0fQ/wQnt
Vg359z0w/expmiicXeXIqVxENU64zl+I3hZHJ9kR3bc6N6OAavytZ9Ry1IQmrFJ4rDpeWimRbyd3
1z6oPVD01YrQzRIl+C6mCpVi7pFfz1K0QnQUHMqybw5kicYVSQ40D4y4nZUz3xXLuaHx7uBwF9JE
svTGq1piHJB16B1pvy47kZzjojkFZtBN0uSIDCOUGqsToB+YWjYfsybxEuzUSbcTsZ65XSUZrtDU
XlODP42wX+wAEIcUS4XIYsaFVY0KQ1b3MW01MUirCzBhYfW6/OWFoRgjzhnn0VJo6gGoEbDX2Iqk
b41sT8cMZIOIUUkZVY+NWGJznnlu3mogHFDubAZ+vO2AkzUOQAm7077ScpJezw9QqRfto0EuDf6X
IqhQPAaMOfBjY/Wp1m/ltYTWT2Uh+GBxhR0fLy9PgPRN+6qTDLmAMOC0WTYhrxNw2v1DjACCf+Md
9DElOQC4H0CFmlAQKHOuT9y0GOAwkUxQCZYnjrv4i8V7zy+zpLlI9uwDxd5ArtXL5C3emcdXVnJG
WcO+1CKO07btnjVsWDEjAnmD9HrUQ0nPeRfGr58YiPn821io6qg7sY/mVue6612jhptvaurzpi4H
HpyZdvGldP/uoZTx4RhBT7COIKHtkzatZqd34KBp1vVJ/opMqy7Ol6awMlK1EH0YFp15h23AmNGy
opU8NyBjzig8jxSWJiWhOgsXiedabg17Ih73v9j0cMsaQODfxXtoSdmSzS+cXR51RYo335Ov8uNp
STUb6I0OSWWDKC0BfcgmMZiHRkjIXlPHgzNbiBh/Q+uMH+mj4QCM+UE6/4iV6rNYXC4qYcGJWpv/
ktelZj2CpvqFu06CuX/LcpiWtp6uE3GH+K6L/4YT8U8JdcPyx+ySRmi/uPD2WNxJqRw0/yZBK2DZ
Y0qOewFgs5lQZApykzrUho+zj8dAXvLcQoXBLFtxkLkVSWTYzC4o/5XHntvshn2xLNCkRqotmpgZ
ivMJgcDWjbtCrG8nOjh8w9yGC9K44RVPT/bRa38ugg9lKuj9cobhP8H5wuzqsDoFOEK79JoVkRfs
+kHgwwWJoku0nPbC2Lq+Zos+/ET3xf7gt4rOuaSUOq3U01+R25GGz9sEbPx+JT51vJcNqbzMiWhu
4dY+4AUV5Uo8FmOBdLj/udNRIWSA4WuPqk1OMsrZdv8WV38nVZSMww3kzQRMndej2LRcXBZrvCFO
jgDnNux+6LEWGsGn20CTV6MBxkYI0ld84WJ2ajBltefMOxfiKcn10AoNhaEID7A1aLj2NogEAb1d
HwBBK+2e1xlqK2EKW6Ml8jTA+JpF738UPuUJBsfbCI03bIzwKU9t8yRef1YduP5lhq4BT6Phmt+Z
R5i1n8TJL04c6y2DWKqSFx5zJVtXU3QXOV3vgLwifR9w1p9tqJfFvkwdaXVVUcQXNcAm4rxQP/V8
04E0YLgJlmC+qfECBfjdcIPSR+Tywf+pF34PPoM5OcdyIiLbbnH7XA9xt8MQJX615JEQt+OvJhrq
Y03NWt1zI6fl+SQMN4YRd1myGxywoIWz1+w3Ps4e82KXJGmfzjG+JrEV0krfPvuo4TbYhcjs7mrY
Iu6eRwVGIhRDfphAhaim0wypswSaZxDDYS2jSl7z1ycM0N70p3SHvdlDRbJm3kpD8c9JO7l//M2g
RY3yVaMEgVjneEIJUa6oji0Mch07XPABbTvMZXwKgeuobe4N+MMbfMKzyR4SJ/tohvAMD7DcxFA6
3VcAXNr4S4ATFNREIOJukOZ+Wz/nijYZt/SHMr+FP7gEGaSSjrK1CqAOKfoCepDasdcTNmhNWEtt
MCxxIcY8cjYNn66jMMljqmgq1jZ5af+HoUlHYefwUmS6IOYTn1BMkylqLi7+1GgZTRMjw0PNq2zI
NYMPe7oCUsbECsgVjQo9MDf/ebzy4KtGYa4DVune7bnekhsSNixc+po9GI77wewNYdMHFVAqFfqb
pKMkpES0MbF149vc84VUOu75JGrzyEqjmZN3rcptbbPaegDigTGD6GHeElumqnz9QPxAw+OyaoI2
lpwKpQjtZ/Gs6mDYt+/iYVMSx1L0Z+PylmOFqhj+3QheR2UFkjNHXz1Ylp+AvrAbRl4q6z0OBnaj
u0VRzn4RmqAvxfbMyLWfi/xteBmZS/azAPNtLpjMuPW9uv7dhKDbjM9ldxVfGVvbg2auEjUmaTPm
Uv55pyEUEc6+1KbtQkxXmxx0Wye/ZnLGFsHVwVGnD/EkRFWbldzsMqw4OhPQSX1lcAzkEz+hQNkH
OZEWreJt+dZl3+inTE8JYOaRcCsVVX9BaA38ZYuv0dwt0UdfBD2MGXWoZIauWEL5StS5R/KshZ/c
cIg33skncoIyzgwo0Ez3ZJ1wQZb3xfJAxdK1ttaWTWVYupmRtpN/Rz5dqIyS/9xJsORaWaVnOk/W
RL4lQCZwnOd5i0xjVj6yYoBXTAA6ShF/ObdU/H0X5OREN1uWHYYaxGlOSr0KcADW/OeMhhGPIk+P
FQ4ovYmcGPuK5i9Om1JzpFIpmLEeUl1rpDY+VkTw0qWVudXNz7wr3l1KDOGdMJwi+9Cvcj3Gojqh
dm+oIcmIuojowF68o/K/kxXSueSLjbImVKFC6f4Li72GPAGolOVIThxM54yBY74cO4GLyjewMAcW
ZnJzPXDKWHf6eVpRGr/I4Dqy8p2gANEh1SNoVtDqaIq6j6duuS/HHey5C48vovfJ23CTVEB796NL
ovMdnMSNggV8HdDZKUH9mjtUlr3sGq2re14ANC+VSSHk9RcnA6vvrkPXz40LI3rVz1XScnsSxs/N
0CQn96WxFagdcAfEDlI/9BXfwYYWi3Q/7wddB4Wi3xkeqgnbZ7BrhsbG+WNP0bxVW0YMIKq3nuRO
TvcyzbK9QwUZCGdmiwdj1LC6Q66NS81PJIPgBpYulo/0/XG+YhqwdDxJR6HQuySFw//klKGttlhB
tq5JUjdoAB7XkhpSlySxUB1FEsdzd8sV/xYGSXEtuIueenFrhQQK/lCgFsG3d4xyhlz9Gl6WIT3D
q4OhcR/ygRYLolfT2xmLQ+F/brMDTLn3sZk9ktwMRpzk1DZ8CfTsX/TZm9SjtOZ1Ri+N6npOzgBs
QU0LBXNy3nJpuL0sPKkyuq/AMpxVMkoG39B6RzKXqyArlXvRykZX+3EcHeRaHpX5Ml0F+5SEbg7d
Jt6ba1pzuxZIl7bDWDc7x9oOOfHCiKC2YeTsOCFo1PzZfpFqdu1KJEJAXvJAMRsf20LdK4qsi4y3
NdKT5gfQ3RfEjBwN+CtIlRbib5IzgrL6aEMgKt4Prp52IVl2CjX2OxKCXcPOeWEVypm3toM/sqsi
BK8sWw6tLKjub+6/I1n6ClNofl3gpqVhFOuj30LHvmLVmLTTUuSPEvCp96sAWq3Kscc8J+3S7Uum
re4XoijrFHqywycdsUT5yRuE0aDQoq4/j7/q/3tglJBX6O41+G4q7DbKYJ/dHfqGVzg59mpvmCg+
P1hTSDCs1wO4mF6qwm+cF3R07pzkbTqS4dYkgjdO902tj0w2eoEwbyB2TBCA3cIu/xvfHClUspIA
4DdC4I2L37TAtYcCPzXtiarZywOtzDrTMuj2mtGgNDfKew+batVpEUdkJDvxrEQ1T73YXxIQor8h
yvrTKEmTOiMSZY6WvRnHzNTh4uwxW7F7SSM48/PBSIWSJm61ptHtaMKnGPz4mkEg3eRp+//QeVb+
SwXcpAnVpqjTxwN8efjKTN0atlicQ5gtLG9Qy1HfAeo/Ox5T+SrIKmVmBXrfi5PW+5iEqjc93kIu
vlq6/TAlogrwCFcsB9JNzuSAdFV4wNX9e8ns+ZffjhIkgUVl0eu4ZerWQLTY2JTgpPAR3Vfnayf+
d4b7YEr1kZ6vwJJMu8VojB3fGz5PpnM4+ZCKpL9qYVXEjPlawlS6CAREUjFNvrn0KyG6iz2g4g/H
z6hKbwYnUNWUykRYVFsa7kA4OvFxRjSOqp1Lu9cPFKxTkN4Qe8E1D1ibGSq0DjDteXI81Zfmqr37
wrmi7XUlzJ8LTEuOC3nLlkPHT3EKQA0clgkHer790CBAnGD3AOhAKj2DUF0AucCPH7qhi5atR0Bt
1R6OxrT+SUEBfDKXWqkec/3BsZBlpvpTD8cPsS7D1l8cIHNrhUzwqwsEDQGfWQaxfP18iEmt+xUL
rGVi5DDlMfp+74enOxURH7B3TTTEtq2nOqA25eAQfSGvN4fb4ir3yGzKfLFedMlnNP5hVgkQpN/u
+Zixli8Gk5x3/tbF/JutZcBd1Fpas3zuMgnc21nrL8oC9dr6WM1eJdnP/R+/k+knMXqBgBnns6nQ
gLaFzdC3nIqKXQmpiHIU1YH7iDIH/UchxpAyOX/MOX5wWqlpUI+WBMVdbBnNY/7s2SL50bllPEPZ
JtLkv8gXrVGDylS0XuXpCxS+0Uqzqtlsr40yFbUgwzwIPPHXNA1HftMWJt6hwhnGZCxtM9u9Qk/f
COx3yTMCeD4MoGFkKEgzSlPI89Z/4GsNGC0Ua7sAmJ0jMef60IPIlKmx1H2qkAgKIqNBbVA/lxyx
FHbqU3K9OgsrrEE1kQeDZYWSaPwG1K7E6I+aB8WNNYut0sXnk4tEI8PBswPamlFLbSUPbE4vFJSO
J7ygXF29faTCPXQq8h6sXBZlK89n4otG/w7rkBpmwQpZAQVs5oUuvkPvgseBoumrRQ3WKw6q+M3J
jhdb8TlLcC60sb571YKyKw+bI0gqYPGBE//NNYqvQFgk+aPcWyF3XipySRUU3/RgCk5V/ghfPQCW
o6RlTcnQWYmgDsGaT5FZ3oraeVq9jSSm2a2exQHGYGsY+jI/xCNnGGxH9pzMc6Nlnjbp58T9+WAl
WIvlXl62vh9jfgZ4ibIg9DnXRthKt/xpxKwBWX8P2MERulik4alHgNZWy/owNu6y2GbP3CfaHK3S
C12Ixz8fEwHFejES44yK1lUZzzO0fvefSoI0c+P3l2ngVj92Twk68VQF7vOyP8rEOOaCpuQUTeBc
jVjXO1ijEt+AWzFNEkVLwD+m9dbnw/l1BBfQMto8UkpZrfa5yJvU8wF45cWmgI0Cga+5/8Jv9nvD
yaKFJ8HnVheTykXNr7xzRFi1G0qZTWRMCmtPAoMJ+Ny4/Y5ydivAmgDYXNhEbjxU/kGBweHysPWU
ThALKgwvyKAItoed9l2b4niU/yRoLHGBI0uSeCio0ZN74dkAAdg7zqxPFgm5VFAfNz9b7/0hbIn3
Rrqvtqeod3Wg/1Oj26gW/FZEh2jLEshuNwLCwcjy0BwRC5b+ZL42P0U7r78QcTIxsG22DTW//0Gx
1NXLtynlKqimijN2x81L/q5Pgh8KIcz4EpKO8m3IB3s+hBgIjZ+MjwuGKWHaCgI4Pd9WUEaHXU+Y
7CJ/0WQVNg+y7h/X3qX2fN9BalQlbZ0RAKyE727GPre8wzyd0Fq5FRXI9SM3KVTO30Yq8iUFGTeu
MTcxMrFNNJZzr592FzhtRVGgG9apAgPpd1fZIQ9BrkpMpbXf1SWABcQNltsL8Nk/BKXNsB6ygTVI
fCZkApN02QklXVy3fHA40j8etN+5k6hBUy5A4sPlr4qsoZbAxLHvWlNer3I5lvzSMTASRuR9OgbV
A2kxQLyxB+lbquRy59L9JoV8SNmvXNd/QNU/wnz7VmnPeu2y2qk2OJvdfpGmkH5RNf0tepMxphW9
F4rdcVClcqBBjFQrKy+ceiUSMjdTaEnPJrJs+f7+SKbWGhEsq6371GzY1UKw/lYyYqOV0FzIznlZ
53qrkKZfx5/tAse70jLnNYWF/BGC1FDAabCFvi4Yo9jbOblzUoJZDKmTJKDYL1Hn7rxNll0lValR
0Xtd2aBd3SEGsk+qupKS1SrHMuxTy/wosur+l4epIuGmk6Z3eJCDtbAScXunjgqZm99/34Y2DC3A
rM95wA05ZL14Mt8CgOowId5eFfJBzbmg9EJFfQ1bC3xnD+/JKoSGWGKTCsi9urUykzMycaeKoTKk
MZnXBKiNKo6vbKQRHTVSJpHPatTIQwk4dOTyeGHciI0QBX8nmZGtDVT0tglByxEYRXVnBm1s0YsP
AoSZmgPoj2ZxGbkkpUBeqAZsEXYfzeOZXcsz7sf2cwhNBZL4ONKOeXplFIEdyUret91547qmJu8e
0U+XFaiV7Ecptwv/gmSGnUWlsRnYBl7PhsBpChscT+AggTA+GyaEyzE3HnIcSFfUMrdg4OWgfvbb
zUuhaty+3Y1LGCnWITws+dX4LGMDN1lCMebpAMIiKlYi2PfPb/5ogU8e8n2SvJ8mcPD2kjeQZ5al
3bwiV3jkrgvzexyzT/7ig2XP8KZOldfzcieWX3Dd2s2IkEHkDXBXwabSVYmtqhdDrEZ9XbpL/mX6
984FigipqahiK7z3D8zfe/G53OKJJoDE9Z7czgYr20DYsCxPpGwNOAz1zufIDJj+708IPUwFFJrm
aDljCDsHE3usz4uYGfSzdcQpa4+qmu2QMYTzyeOrqtMBypN7dScu9mISCSyMSSPR8neT0T6xfAmz
gU7RWSCVBYxCqK5KUGImrWAgB6YQLk1OU8xsh+Da7MGdfs5QAfiAtgXD1aIUfTsBMS4ATVlH9ULw
WUDhzlLMq1kM0PEP3xrFTazWifNqI1QQjXBL591Bo/pqCO5mtY0blyoqRNjNV23zr1zbp3le6HV6
e2Kgj+rCI9u0aHwVAmh5PV4UIjUJQyXJfgqUMDgHtzkccSElBHKBothFkNAJatS0uAMiFDgT/6gm
ickwSwJLB19HklSCVGehHkGoB56ytmCs4X1/74hOm3B0/pfxTb8WgC3vGgWfQo1ZXcN+a6yhZ0SM
N+QjX/TGs4HIlVv/BmCqGwmtXaW0jDSvWfSfrkZLF7hD6xtNpXJh8B4xC5c61DdeD7OyWnzWBvE+
tKvOn9yRxbXfBsrqK0kZdlcYCkTqbeZR4e5dYNEiIY7Rs0rNJLpQ5Vg02cxS6Zym4gwYNZil7w95
YJNhg8Tg2Rwvvypaj0C3Ad+2IbcRfMkaesEf6DA7mUzo/elRY0ux0fNWAmYs7yEq9rSdHnCwiiLS
WRQQts0j04l8obhFLt+uTagqdyVT4eX958fmQe1qmUghHV0ws/aXRPMrot+YV5eqGwDjf/6sGH2B
nZ9o8yD72NbHUskJsZ5etaoXXsnKj+Oc9YRAAt91cGNdd3zWYdmCTwCUJigiJQrPew1h9oxR1/JG
iykzKeLH8it+TsCwg6loTiC/JKTyDehjSBfkGuVxWIifK52NNjH+3unmHdpwk6NvQ3g6g2jd5/UE
ZvvMpuzKUFg/XM62ehFOfntT9/1yFumq35C0qdmMuNeKHw9PbfJEjjn0pGQLG0ecnuhIZvNPTiHd
c1o85qHxHUoM8NJ+GodgbgtAgUJ2TfYGc1KMou8fK0TBU47iutXxHMW9xjuqWE5ikvIwsQgBqb7+
VKxbtstgJqW7qpqjUTtZvcxv+kWFJnsRByooGBiZcJE+reIk4sVtm3KkAFZCSRuIO/IYLmdUwSwY
9MfXSejxMbi2PiL+CQViKiG/x347j2lwbagPOlKt7f2eUyD+BJSof8NhN2VO6oHGEF8uxznku+SG
17kt/+ZAuwv1j7DTbRL1iKl89257Lf4EEraY1Iww4kYZ0q32d2fke+z03KVYnvSlXQwfqRgEYFz4
taMH5qNUxoKqCRmPVyMksIvf23223Zw630mciW/YdQejJO0L+IvVFEgeMesUGPGIcXJLBOIW2Cwy
3IDa7x86+qj3Y77wvfOwMlvA/i1EZIu4YnE3grzvGzunOn4x8HgS8YlUZdEb97nONuYKFo0OkxR6
XKznleTpADBMHZrwNjWkF1aV8I9itYWquGyE6sdwQfIIdW0x2X9Q43Y1vCjzAPui/rpFFsLK7CL1
xxWLK1I6fs/xp4BMvnb1tR3zj5jLLVZDbKRa4UW+YA18EShZ6SNqDUg9+e+XyKkFjpn8EEjwfcbD
UjADh25XRUW8RDoQ2J0BRGFzXgJsYq4vTu9FC+y+vWJTx7aQ/xPfE41d0bxvIYQiHGH0Xne6Hacy
aLX7N88RXxmlHXsxi+TnWhfKOSyxO87qO2Cj710Fh/DknLU3kR0WM2KmHeCN+5iSl5bxfxI1r0cl
hgougDBjy39kaa3SPyAwmapgHsqSTw/8H5smZ34E/6nJmXMMcbd5/ArdRxQQh0vSRZNsAkyTm+33
0oBXxM1rbwRFf1JVkng0/LRTuc1rpgz2uZyKBuOzupp1qd1wNRZIGZqKPr1IEnDh6MKdDIV/sJUN
q3HuNbuVGuR2IYrXMFtV4Z7IjSOlSycc9otd88mmqOdbhblW3az/axGeDHE0BYduc4+gOoOTcKIq
BgkPbPxSYfxnbITKgl3G8+mc+oaRASWHCJNw48AeGXbFObF3Qby3Deq6NDarP1sNTzUx8JFaQJqL
An97kdQpLySl6Cg5hLRctCXJN6bgPT9Hi4j6dfns7l0WJ3y1rNAIUMXDnJCgE35cUyAZiCagGXFH
7J5xpW9vlr4QeRRa1fEpsjiByH3xpOlKa2F7U4/acM1+e5vXqX4b1BaYkiDPthmrm2n4c3Q/aEnt
gkiFopY+l9WbCI+JyCcgw448Bw3pAAVbOb+Cuka+2u4fzhUNfXIKJgMKyvRNphKCWB+bmGA+E+zb
/Re8l1cMBLwFFQ+c7UDhttRNm5PsrcPhcE315zQKE1ut+lG3meZMcthxtEfMPS496VhKIvF9lgYR
36myE20lQmwIQvzRK4sWnvn8Pcus4bINzwsnsUFL2nn+Lts1p0oWbUquPsrKpoBB7EmAhbXbKr2K
31Dk0ywT2UzDQdNYkXwQBMaY74B5Pewd8xQIrsi5WAfzuuPTkx8OtRo1Z/kjAjs2y1bMDGzVj63b
FEEK+BfVVTMTk7AiKPYBiXoTOexg7VefBPv3SsrgInRft4UnOSTdn/Xq+rDuQBa9PCHtiyCIVP1y
0rTRYk7Pccw5RRhS6FPWXJBeeioN2Do3URmorgWs92V992Z0gWxZIrr9JUd6NalIsCsbwFJQ+bdb
y+nEjEjMLg648G9ha6FNvfA/T/N4FWy9TNM2/J7MIt/Z2wlNjoS9xOQ9SZ5RQKc6uWT3lZjK1MRz
R/UeOSZZsI71rhZDBfkXJksnzSW+HgpBTSHzjxdyPbbtyx9tm7+K896HiKnpaJkS4j6bZg7d3Qfs
w4Mfz+0fl7gC1BTFOm+jPFwvgXVJPaG/LJ4lULHIE1qV8sefZkYp8fYO6tCQcASowDfmkj7iSgkw
Cwr2EJAC/6AfLEscJhZE1TDhHxhezcEp5SFxoXtS1M/E5Ix8D0F1h7lBSMfu/hDN7yj5nwgAccva
vFRs3NVAMLSrzRSXWrippMeNVkk9TXItkgxkSQ497m3ktmRGPgNLhGq8L8qEO+r9cbhRT7OI1umk
dzTTdDGQn4P8sixZZVPD9zKsM7hYwRhPu+zdoY/aoTI/v7uJ5dHtZWvJD/7Q8Dkv0A/7Bdc6AqRU
AE72GPtYMhgkXqCMajsyFOrpnqs4mgmqL0XK8KsL7008xdaXk4c5kduO7xCGajmWHh2FyEUTJe6g
EzE45qnsKSf9smus6jEYWYve1eNeGVWvA+YM4GM+TCcjRzCVaOu1DhZhbbpn8tcCAZScdIXpC2t7
oYv5tEWl4xUeNZOB6aexpzoPmuFyWCoh7sYE2ihaoJNfoIWcrgYG/rZmqkZ0kFaEKtcizdDNmwu7
JtJfzmDjxB+mVATUT0VPNp0Swlmt6h+Ynl1PwrvGe67lB2pJnCGZkpon0iWFynO6ryEXVtIQIqfH
+AfRR8q4ecX9bMANBoA6XlEEfFc97e8kWaUd3JqcPZSywfnD64FKq2jfqOQvlBhxUcy6JZ4v7Jm0
KZ0+sgAkcPPlxXVVnts0DZxL4sXxGJheneyTo3IgRYSdnQv4qCoCwbGCpUUM6LkzUSoDWfXnh73b
uE5syRkdZxn0lgbdmJYtUm0M01UYJPuDTGuZouk7V8mZ/2KghR4hCs9GUTePZtgDcTtmYKhlSgCI
T1N61Bp5gaw4r6LFG/vMKZz7Y/J7zd/ZgVOPLyvHgqGJ1u3OQioG44NiHpRoGY+zaD3SQgRJVCl8
GdEiHLpWRAKLxX0sJ5HUeObuuinLz3RPCyYYNcrbO63YJhOHVFxAQLO+nY91PlsravFGLnRvDg26
8Ud5lSEpMCP9u5j7XCa5HxPYAnnn1mZW/acX9aCaBmJfdFSyuocFczJi/6yhrnD04dLhxUJzwbEU
3qVplTpKdoAlXxR+wqsijGgY2k1HqsH06RedIxNwF/X//v/65+KrMsWw3qXhgauOHeX0g3jjSDw7
2TPmF8sU7US9gV9AXh2JbXmkh3MHJT9zHUdmed4WiWnCNTSAl8kwbBxKBZ8qsRZm4btvJWEWw6zt
t9FoZ9T9GPnqI6OA6cbjq8CmlqMWJ2i/BlSgUGfrlJq6JsyKKPB7oWB0zRZPekTL8pyC4/0vdvao
+zCvVeTcqdKyoZTcFp9FFExAkgShRqpHtIiq3NOBLaCWnK2PDtuXX6earM0TuzgQo4FpAmPIZtFL
ka/Q7uxcoAL4Rdubt8M0L4lVpwppD/txhK0lbTyjOf2i02se71et4l9mltmdbVkfexE27jH0qfHR
faqo5riRd7BkmJCit64Qnrgi5UiAXBAeDH1qtxN+yjLTSHuV54AQCiFZuM4zPd52xDy1Fuso9zDw
Qtj34tzt2STC08BCNMEYUAShIohfjZgsbFaTsOunMi9kmjEyzt+3W/GdMA+7ZrjV4a6UmdCzrhzE
fCgs0WC/sPPr5He7T0D65kYZYUeWqj20bbuz0K5HtaAHd3N5QmujGsrAoiR2GaOOcDyZdwtEsrOJ
jqSRi/SM2ongDW1hvIENaGyO7kaFJeHuJ8iQO9FevYvpXRUgTYSXwgM+QPsDasLW3/FMPGGEyQg0
eko+WA4Udp4hVIYKqXQ3jjoK/NFqI9DIKra3Ff6+MJsXV9tqyD0jkwRDDXXjR3Y+PUTkKH6XLFNj
WjtvgP1yK/w75BamAOZ2VctWiYQ3ZF1m1wTSwWaxPDlfoxGqnELlejBAlUuiCneiBlKya/9HqupF
g3Siq7OHvBj5JH2ladXTmUG+YBhbmFQZ+a2zRYt0szBR68JLxkZZ5elMZE+/4STCFikkytmWxbDl
XNqBqdzt0AYWV3aS132ApZwogmpBCtLn91Q1VnhbAHt58e2dJxi7qqZzdwRxw5YDEg4I09hf0yZz
flyqgfwHSexSF+YruNs/OXuoYf0a6zN7ToZc+hJq7gL4WAW/ta0Q7afuGkaZCi+K8t+X1wPNm2+E
gEwc7SnSpQx1dpCvRsjvZY6CVuuDka/0l6+5MH28ulB14avlz2spumZKlbtT5MnZEjJLweMjk5F2
FA5lzzPPjZTrmByZNMaAH7DFNRbyQlPa7TPKcuxgyB2CUd4Tj6w6SqfI7K0GB0JGfAz028D7aXsi
GXq3bLoPBE2KO9LcTURs3xduM1zTqi/OvuD4Dtgk2zOxB1kdghX3lWihDAcGDmMT9W3lBZju2Trj
ReffcGqkcD73NPo8P4MFivg6eFyaADjDn86biwZb7wOXB83sJIBNq98GiCEOLRl9OHec0Boalb51
v8STNzzW1PVQS6fAHyHtBiZXZw5xfCrvqrnLa70Uv4cWHmhe3DLSZnSHPontKP96uVv1fjw4BQsN
zl5S1lLSzc0/ILu+nyRlp4Pg6ECejcItIcfmt0tN+Qv4j6tYEU/ANp+uz3LWe1IBPG2nzH3eBZju
UjfwjUJGvJRhheeXto453z73nx9hxHKaAPSKOrY2k7+ilfZwpzTLw7mmdAZpF2kVg7LRLGEJ3nEa
EVy2zsU+erOXP2KzJQQJbMYUqVCRv9Sv4NlZMqqZju5mbekcLhTrVDABbuXfogVJymh4tSkt35Ys
QXncg+DGue+r8dwEe0qixrm6GE6u2wSYoBGCA/Akhm2armYWcqYMfcILn4R/3X0G9VukJjB8+Ghe
98j/MDXhCIQUcJaMslsoj0nyBiHju13z5ERmPBvPVNvcTBFBC8bXtVMg5ylGRoT7IsppJjNWNykV
46Q16DcIjRGayIFPJH//isbwRQxZUs241/R2sziSTebETwp4Iy9BM66ZuaNVgFXvoG68+Usa+Z3O
+T24wCcApvuERF7ppKyrTsJe8Y13x7Q3ltlm76P5B+UPk7d9Saej7U/hVW2sOsgcsrnua5hMPu9J
OE5y6kl6VelDO53LE1Tx+vPwHyNGPS8+wUqXsfZ65R1cH/yR1e7v1XwTp/NoDEoNaLNZ6lAzBuwf
bnt+gsBdlzY25BqkPRODiVg1KbGMB1+2pJ6Z+lwLvZd/H+4pd6W0TiyJ8bAey393JOcMvZYwPSJl
zKwHg/1teb09k7/b+V4l7DxNyT7UEUVHrXcPhjiFt3oWC5sab+NXNeqMQ9lEI6QLu7OC3TS1qErB
AFLmaRlfCSy3kalbf/zgUjBf0asLph2ISHGWhhHGjkQ+m2Rt3LDc6Xc7lmD1lpE2ZX4U+1fYpScl
Xg3i64tc/ydlBNO98noenaYJyJB6rHjsDlPjbZVRLEuIYlmWRpHj2W6BNKbjtw1LvdqpRuM+IVfT
o8dL4x/46NDqEc0HW3slhXtftM/0p841fZlg9XOfEbqYbm3X0tkSCc2j5se+og+TIX+lRJFInF1/
Zds3HXTDzNvzq4VQFNfxJoU/j8p6AxhcAQD8rrJnnx24hBPYdDcocNMG22cT59i81w/Fj1Gb+wR9
PwYAiTHh7NgKO04otTAOS7sIBsy0fm64OV2ccQ5BJF6Wv4b+MpwdQgKsYXlo8+r4xfUcXsfv/hEr
gq90R2i550q17pVxzEdNujHQ4iUhMdcP0OVjKOUyehYEdHHgutEORZVES3jrh212+tJl9CgGdPkh
3ZbYc+mZtlz3sbvKAI3f5PC2FxsOMO0Q4s5VdWWBJ8JqutVOOqH/ou5lq7NNup3M1ebjoDXHnPQh
Qc0g3PP+NQgMJfurZPHZiZfTtipCmuuZh5c9I8lPQYSjghMgt3PToIsiUXrTU82dKk40eXDzmsAT
OoTXyK1o2cEM6KmCplKZDpQSSE17epWeOZKSgkaPiRtTYvpVMHzKuNIXNpuYAiHHtqgfOrQ5eRJ5
liezJW1LlXWbAhGOmVMYvNDpITbD8guEJN/SQMqSWHaNCgWwU0lCqtpqZ1ueq2vjXXQto06AVUST
P+KGLoAQLsaOFQBqpk9tlcNlIYEn5d1nlCPI59GePXoZsj++5v2JAI6VnKNM/egLD8jKNFKBRLSU
DXuOCg07UKnbVq5jzU7q14zwud3gKP99UJMslq9Af2eLG3lg62+36B86I+6zRuVuwj28/ZKmhE6f
AGtVnIyBv+HpuzLlJsljPXw2kS5S0WmGOPCBugVy7pirXLzfWKUKtQtdzukH+eXFXvmaFdT2WAVL
saiYEIckX92V5y/GbVeqZ4s1NP5e6dXce/xY+GBa8fqEaEWVW78/jdpuNG7TCvD+yuhWdCFEgJ5C
WmGw4biIEO8dCKeb28ZufzOd32Q2tsuKC2nFMoJyRy7/lZnWcyLABvgeqC786vULulrSu+Zrm97e
esBSanwVA9UxtgTe+z+xW9wvQuFEVuP7D+SVmjRjKMu1jawHfTHlf+CaUx0iZDz+aNwkJIRHwn8z
y3srt3Cs2ZW2oBZsBYx93LaOkxNu+Xa0vnX0v/eZ7LnbwVvJmsa7MsREFwjbvbiuDLB79dcDsQZi
WSOnntWmRH0lvU2bRUciOvrEi5YCEzbyzxeMip9jWF4BOjvGqCuqgjR7A6BTJ8mmCwfRuukraUDo
CPTMjAWQQ9x02ZU86b+GkO+wvp6veBuuz4S6cuvtXusSZ3LKSc1G8zOnJbvwxiq7raM98jufBblK
0AOs78G8jfyqq+AEZbadBCdX+WZLh5+c/SiedhcVKY0K7AiCKOJ6COsX5hpB2wCxzEBkhbRiZvdn
hZTFiY0z+S7ORYr/J1GDGpZj0RYVd+VJTtIEey1ViwmMcBkhnDWaFKnB37TkTm4GbPy2yk0n3zmB
Ruofque/G5NDs/vjIIlFbfo5p3FrqXtfMLtNDjcOny3tsV9rEnmQQwv6jqj+p04niiIAGBg45NiN
+dz6tAQ0oVTnAXY7gQPV+pleiu/lV32uoThQ071abaeCDFtK6jwFfl97ZbpDbYvAym3XOWi2/ZQC
OY+YFyW7HqKz17CG4jxFhK2Xx75Fe6lXX3rU6751PxiYw9CVI9aVSLgwSET9C4Y4r3b5FfP6/Rdb
LL0Pe6n7jx4QgbH+Eu2bPAW8TfneVAWFkb1e5whAXThNo/Z2H1vSyy8CboyaIGJh2VfTG6hkwgtM
fGyo8k7OMwPp9cCG0ZW9f1BGUh7i2MnFhJLd0zIXiIvvYwzudsfGOK9mbLrq66y8uNUOv6Yfa6Hg
6DbsEyHEColQgv74oswCsLXNtl8NGZKee16SMQKJYzwepo9G0fKjZTD51Ad2p8KyTXtmCcWpEvZT
jlMvbyhgiyjJgAkxqDXfUz/G058HD16TCccbn+gc3LAteiXPnmWvk0vuG71DlTWBNG2XW3+gjvcy
x1cVM5uYTyK1vU/OWNWE5QohWEHImpDPlnpOhi4xE9r+1MctDVuUSt7bbkq1v+hcwUsiRlqfJsUH
le+nNt5xSRSK6R0+Tow+xZF7W2NFVAZxg2Ci6YL/1+FeTC35wnowVPx540diVtJMU/8LjHuKKyVx
QKCukWP1/rjoZvr8dGZayA+4ee8mnX1fd5uNWkk2FK3VR2ibADvpopqhxdyzdffNdEs6zCBqeqbB
V0b7a18UXysIQUxwuuTU2iX4gu7lPxvexzCeJ0o7IFDFPoGiiA1sAB3Jjoo8njHHA+gADd8k29H6
+wvGeTD4jdVIhDYkah33hUNj7RdPmfKDa4J1UlO2GM465U5/KfexVGouHGRj2sSeEu9HMh1Jrk5e
iKwLG0f/79+ttKEDlL/2MpAS213gRX4oFUzgGDbJKSUmvFBAResQ5ZNvXoKp7VCOCIcJYfwYsFlC
oWvX0kVKmzIPXPKS1aELwKJsvL29WFaMY9WmUjU/l5SgX0mBeLw6ncTOc+IOWpF1M134ILkQVK28
gQIyxX7oHgpGbcUMGylHym1n7+D6BUrpJLvOlbB2mGnucDit8LkRPWF3C/2VzYQZLofeM6iVfoZY
OIY5m3O5aQhp/uZVrlAzDRirzIvByEpUWB69/Evzh3VIFZMVcKTVugICINbUWCEEqqgByDb2WEbv
1bZaZtHsAx/UkiWqzy9lP484ur1H+zZklPcPq9PUzesAjK7qXcguWm6r51uVgkTDcr94NpDFiP0r
9t4fK3TxPbgT8+yqmlvKJyTKCV74lk7ctKH8VFqeuAVlBgU/Xwfcamy0g/f6bwFOZpNbp5wzwMGI
+SupHL5D0HBzMKGELWopvz4FExjD+vLI3ZNcx+ijIvhlvEYV8BfW6FfdkpwJ2Y+AeoJMhTjORYEP
3GH9ZENYHyITXKejwa0slag/zluT+zZMj89rxIrPw8Pxyv3W6ZuE5YJm3P8ZReDe7K3NIYfFCbv1
Nsp2y8GFzgktkhV1YkHLBfiUJ5Ven1xR5YLoRBX98dTEmlHIiuoViloG5udCd1B4z7DRg5XhUlCI
3oFYQxPMb7VZpkT0d+c+STDjTtw3e1zZ4jGMscM/tgLI8vRl/JVGBQpH9Z0WtMWJAOgGAgyHxdzH
0O9+KveJJg9IrrfHVgT90Qlm78xDJJ7Rd7YO1JR8JPpBLwZ+WB+JXM67seHTKCnAfJcOohajDpHq
Vb5eE5F8G3JxtuITu2EnogBHaKqXPBBmdyQKQy9JFochnR/ydQU0XNynrHv9WQXE7l2S7dzUjry3
5A8I2bfI98UJKpzdS9CeEsNhY054N0nZSrstNZ+mH4IQS9Wy1wGk74cSbzdZ2f5iRkAjlRzF4rPU
50kUFlXcBdb1tM9M5XV4oYciBr12+HzEDWm4nr+C8BR+IJ+Ezf8pQ/BG/2dBM1wME0YIBNHVzw8U
bU0/xjriT7c11mIiyFGQY1bXcrFnyzwMmOJpo/dmWz1Rul+miOKc+rUP2nWwQG7K/S5YX9C4ddw1
n/+VD63qUKgWsZ/FxpEMU4N7Db4t4yCW3vbe4InetzXsmrs1xVdR0mxY9ayJvbbzOg1Qm3f9n8ax
7lq+kaxKUCfxQNImk1fDMcM84M6WYa+JDv2aUupllwO6eVEajza3oJnbjVykUKY9Wga0XIxYW+h/
LVRK544d3EI1jzhVidGJrk1ElVmRZGQmwnX/5q3LEziZg9OuKjt8tjDxi7vIFtRwZl7UkzrdoGHl
Sp7Xy46KqAKiZfli+l4Bu9uzHEnoizo4kdq1WqelecLB2HrXw1TEp6rUMuhZJ2JyCxBifG9gSeS1
qExlm2qJ5krH+RCZz88cY+7PvLgIeR8MmfruyCSS/8X3kAdY69RvlwQNjVk6QIlgTPeTSdpy0JYm
27oFjRCELYnvuAZtJtuWRt1z36mYgGF20Vwvn4yc3FWezIaqzyiLVXUBcdR0OYgW0E6S/R2cdpvE
m4ElAjq1AL+CR8Tad9AoCUokxx3T1KuxEzkzTphM+sGAX8OFrST3yyyvO1iYCrptQK2Pe5HdQhPJ
/LR9NaDG20p3qjr+RBmMtZPsOllNIGGg/sPzjWrHkxTn7IEFsauDTC6ikKqH6L4Wgv/eqDArg6/b
72QSe3zj10eH91kQXMZzO5tTJWNj8+xTr6cAAjmzC3aqLQJwEyNPzgV/Ba4FRK6bJs/UhvWZYELc
exMNx895ii4mAv6osGF9wN3VRz/8+o64Y58QxdMJtrE2CQvdhd7wH2r+GUdsXH6WhZP5dv43lRKj
wk97rnFV/6HweNQjMLWW758sqCZQtJ47HLwiD87jFQfgrAjFKEwurDghXuxFo2Gyq4eCMQw0Bb46
9h5bFwmHNGDQaKGKJWsi2PdvEleIAfdgaMfDv+F4xxcQQGTcJEKObCaJ6q4XMN7N2Q04Qa4lJHEr
YDia/e6biZcsY8f2NKVdUi0jKimYvfCf2TJ6lKZhUCgiy9hE9PO1EyFNE5WVQs+3HHKcPgi8zNfh
vYu4ecvnX6g+OO0EEUTxC3+cgRrMI5pdPc+ysLOt6XzozobJTnqn6VP4qn+oMlvHRWkk6kw0hEiZ
7OpIKBHam8NLAIwOSMYg6aX+la357Oj67B2YtCvwtntIsG3uTf6vy40nbiKs3eKyhodLrvRXsGcx
IerGBc8Pzx6iRGOf0W878rAEdz9uc3CGLvGMtyc/4o/Bxk7U9F4xlyRKfnOF/bEcZhIAuaRhPzOt
PvhHEZ07neRr/R3k4kVN8NR3pnnbAWSxJSmgNUpuuQrJuqYIQXiosnzYeeCAuFHlCJ2RF8wYgsPL
C8g0t6xXQxs9RZ6Y/m9VgL1KNmdYGsnT6ppVYUdeqoygXwLljYUPEsibIx/9apgxsZo+TBw16xWe
QWlg4SFSkhCmvx9FXzYkkAbMpo+XYNIfHaF5Y3ABvGL1zyNhI32B68dj7iiL2DkcvL0pewZ104Av
KNu42aYkvBHAdxq5ln3h1zPyqvy4lqyZRWAymlOOTTPgxBmOHdH0tPBDmm+ifQRZUBqOZzRTyW8S
P88gai13hm4k3uRq8qqoZszztRlt6a+zz4/8poU7sDBKZMXVX4VJnl8e0coqb2BBDVTTp068Zfo0
GvcBcqWjikzxmIvEqEXe+eeyr1gWnINlC1ywpbecFTzrZfAt93ceR5Bgs3luetk8Ir/E7Z9lMvcH
W1aneR8hDKHCq9yWC5daXOVmbTxMXfXFuICKf0NQlssFm7ryA69vVp/uU04TF0RnS3ykwaEwFqPc
FaHpVBRnkcpNjdK1XHBvDi2l6sJVLz93N99qpFyfuqK2GS7YtZuGiSbHN6K94oaz5Y+2Mj2E70V+
c6Dg0iLQRAxzF01/ADExIBglBvra9O4SJhuvNvxUex4k23oHiGBDPBEtpSdIC5FQbFR62T80HYuH
F6MjTHsNBSBkGWtQJxqw1iHZol/ypjwpj8xoEd6mU8QbO/3SaRC77rzS97mXBQCAsJgQ91zmYRp8
4SL2IjlHxDlh+wTZNNJTMv8w8GcaGkY56MzGj0+xZMb9S3YNpFyg4xrfCXO85VzT83io5Ejj6v5n
n8p/4OLb+R0MfGHlEhwRcllPpKvosJqBsg8kZVlZAv9CoPIXdoqXu6iINSrnivuevuERsb1PWYEW
2DZY1Xh7V2HEk2cMBdmzjs8Sj/H9HmRyS2edZIKC9X0Eb86sLjfGo0RbI0CNLG7U9Obar6A+XzeL
CKMByV1+6t1shfRlzuPnoHD8IfJ6aLYEXsdPfSCWorXG/HBKx1+D3m7xcq807tJjFDbnwNwSNq3L
AYIrdxNJFajayz7ZcqEpv5/JakBkNWIYQx6NLMk7GfHtnSrcSgUgdfXYjhw3YN6XlyYp5B0AS82h
uWOX/ujKfMk+JAmePIhMPPAWWkJZOXmAcLc6vrs9HIzEJaNBG5g/YDqzVSnXkKlao/zHvRjU7Qo/
jMYl9+KMQYZxo229HPpNLj3b/I4Nie7P1Br3C23nC4byR8PpJf43MTdzKQPz0qVCnINrfVAUEF/U
SLim27zRmT86NiNSlrLpwisZeF+MifNB3GeSkZV/DT1QIGNwR1qXBqkug1Ve9d9IWV7ymKGji9Za
Ne0Cf137+AQt7sZio7EaUb+0/C2cl/bPd3J/lIBuUoa3p6u/agGGyqDVgjWTC2K1Dt3RWiM4adzz
CqXBEBBtSfDwBcqHjqXHWghtVJP9APD1Rwjz+A81PUsXkGpztEc98lcVORRBVqYl1mEiLIQasoR4
PXhV+BfDMi9BltS2sAmEWl2Ht0SNvzQZGfCaGqYdWnJiPi1+kiLkfWxTOEGDzFhZoRjgldYxA+g0
Ex485UUq6U6gkXfMJ5uAgwV0CQHcahdvUctXSNgSYnBBGiHXEzQbk4jZv6dSMHgNKTOxMSGnheq1
DnKlm+yYO5tYp4/DEVcBlG0r+/Oidd96WDlSQZuSsPRZqIfSikAPaRKoTP6hU5pBgsLMR+1x47oK
95Iy/PTgDGoAwET3RU++WzvIZb2L/ccrJxwemnMda/gLEOJ7IATjE9Q3TmcIsCBpM+zewH1q2OQG
U1bmfDms92sTfkai2QwXoJ1pczxdEaLTuyB19YhVl9BQLh+Rx3mRM5JCiAjl5EpXCaYAPuNBNzWl
njJm5Jj58ywwguUfWnj0pSj1NFwxEx1PTbrB2M+RmaLTtaHGXbZfjw4cuHLyi78JCgMRgz5qjZXO
P5MGLqtbJrDW4jFzXPLW/1UVyElY0lguAxj5KWmv+ikZaTc36IqcggKVddtRvyv6gv/DKZ9yT8nO
hoZEY40DrWjkn6KYBBJW0jRVpdIvgNS437bkVg3VR7RgUFvykb7++CF9SvOmG4ulo0rhuS8ALV9w
1GL91Ev0G8BjSLf+9mbuv5jboiyM7P69/mJNu4zGfuqZMqsmCCn4DIZVvpm+Y0zI5By6ru4UNgSm
rlXkvwyQW+A9e2E46oZH/IteL/uBgSzXi9jM3he66vradWrUXv5AL6qs2u4qG5LQMo9p5v48RRgf
BmY4EU02o8JXq9vxkuozeD88v5eUx902PqGCWgbXvKzukv0jIGqDul3AQDq2+UoTjbYT7/QWgcrw
joS4i5KN6x8y7frzVgInwn/AyvJ5dPdU/GmJA+VZSjo7RWite7f4V2H2aveK/Ec4ipYYylOu+lEy
OhdviVP27YIHH0dUlyLdiYy/VysfadaY2prPvSlNO5IKqWVWmGCEcRKPCK2+6nDpZnKyElUKEKc+
lMlCXuPpRYQ9yYM66cAy1DDwaJZ7QAIBxVM9wzJ47BPuq61cEcCJgYSMhg5FT4YMGGekLOL+UKHO
JdvQTgjF5E1ap5UyOfbPgt5i0hZSsaEFxVbN/vKotmC0fB3dpuqISIjQLMdit3nCy97EnCKl5+Y+
GqVWzMMhSDSjx9QV+g6bJVEt9etBHp04TZiQnqnYZnhDhJ0cMVCQFNV1S3Pz40HqgheX1zPg0OKV
4sxwpVyjk7k6U3ROgl9+cBXfTjmwol5xXm7QBtG+3RsR6kz467GJfGK8L8sSgD1/esuMNl5p7/PR
7YnKUEEIa+0YpsCcxSbQXsxVJJALpJC3U81wFwRvCUK8NFLjWElOeRrYbDjWU49Qq8C5HIIdKgpo
8hBNwiVDG5tal6+M6ANuszdVLNlnBskvfvCBHC9CDzerwkNlb64KptUT5BO0tslt7tD/ll8mZSKQ
cAXip+DMbkEQjYmKxXwhaYFeY9TE2J1VNMBHsVUmY+Wqjdt7KnlZlgoyRfXIqakPdfBJaEK8iuOc
6TjYNxplNLY8836eFNYOgRodnag2OmlbQGfLs8POc5kte4laDZ+AukREK63i/OwYMVMuJ8U56GJd
dVvYwRPl0Cl7ptcw8R44knhzTE3oFpw70cNEP4u08hEq+46WfnRsyZlf5R0+H0z1ccpGOx02AdGV
GyA7FfvvHWS59/QKo/vRfSd1GhlYdJ5seWl65z19EUrTrYqgGNRMrjYAftLxAZO8itgvNdTNaBzi
MrDWoTXVVZUo6ISVq2zj2wUjeQ54g1/boHNexhfHHpLHgHfkUDLiuEx6hROnnNxn5ie/cZWTunml
2cvSWmT8jfulMdNXb6ByGWSPnP4XtR/m/izGdF4plIGoLO9DsKrNtQVIMdo7igH+XXQW1XKUGLKV
tOyi0um4a3wgW9rCR3WR+3sZm1DTqGeBfpxeUPjJoIh9203k4aMAbazdc2tCC4yBOAt9xcnFbHft
r6k0N/m2075PWVhE8koGPpc4QCYgBfoATxCzft/OQ4B9pm3A30VyuKgt9j1QiIxyIVcGUzR3OyU/
BgBQqqJP+8OjIXpotDNJy49cdknIS7fv9tXX7jQ0BZYnL9gL11A2QPP6rgGiECHCO0C0LHaJ1C1X
eMKtJNKy6fC5PZxY3SlBE74vRGHKQUTSjUoHADg+f4B7wsw/OJFTVHiEl9DoQ43nbDRlK2w3t8QO
S1vO1OiILMCq08/GRja5G+Y56a1VwBMWv9T4/qTJldSkwDR7mz7BdCikoaWU5PemboHcT6r5QPjV
AIdo/lNfMzbpX/+B21oVjpbOMAX5u6fx9leWyVt7zRALwEP114sNXRsR4f3aYt1RLP/65pXv7LF4
NStmiNN6eA/7gx4F2BK5TAMs2v5lEqeavkXzHOwMjO0qhm4pVQNyM6QtVDpmv1ncL43y72pUSrqO
Jgyd5pMTZKhmnLZ+9yJ3t39pLuF1rgKLj1KWIIU82tOUOLifihGe9WXCEVIvd2MsI1FjeoLsTZZq
F3hHcBEpq+d4IPV4esC7axy451LCxM9F1PXOIGybxL5huv9eNoZ3vsds47yt9LVh7Ot73GDrH6v1
aqd62l8zffXjM7pz9PQSFCXLXa1aVRn+QpJYMwYhY7BJsH2b7S0sOXd5roXbGXGT9fOVT0gjfQNl
uOedzP8h51W1+KIVcChreeViVrptrWVufjjbrML2adnSgUs3vpDRzi8ArzD7y7DS4NdGF6vVpBp2
mWTYb7qgAUSJWTa5HWTLCVD/0b1//D1o0PHEiLJZ5D/rHjU8qhmRGOW1mwIWmm509ixLI5XGb6ld
SQWkB3VgYg9BYH1BQonbdgTLqhJzonfGD+ttcAxVNN5lKclleZXWaigRwgoGGFahBPkQxGKdXfdN
An/6kblRwpWGBxYRFHKHpW+7iR2GYW8nMWtNepLk9u78tGPDoxJhW1qCzH1I61VLZ8y83nDFfoiG
6ebMqCL52Jsq/KhKyaNAPJxv/SPF38iGKFsnw99VJYz/rf++YPY1n+npMjnVVoc8NlgCCHWIbjZj
eHI6gv3pQ4MrFC77O7yGC80ta6qr4z0DfIukXa+TTrwnEcsuPap9ssM6/pYgrYNSB1ly/Uh0BbMH
AYNXvrIcGwB3aZ6AHrqFV+ygFdA48SekLK/C50he+ky+Ay6ZyRd/JTuVVeZuaQVk1ajF16U4wGit
2zehrtoIU/2eF4bKxISpf7SUPJEzf1xhoJUKQrSMHal9nzb1lENc/h8QFjgZCAwJizklvXgTuluh
i+oOpB/imkenFIuMPqMfxvm/UQ8buY3/BIfCrfw26IchV5HwuAg9WwvokpbOBnqz6ymKPyK27eE0
NmaBo8Vl1U6f8SvxeSrsCD+IAL1pdkjAZKjCJKIMyyf21udC8AuGxmeAKFUAWfA6jQshhmc5XCyV
vcHYZtrUBJUmAxyh+PM3M+v1ltMPTDCgRc3WdmsR6TR3nMG+7uOf92qq/7jffyGuaRpTwhkW+EF3
TcvIeaH9XeVRe7+Y41tEMfqSaZfPnsz9H+SVUYhpmVCvhrSYRkRgadg3+WqjQ1WHLKVNrfmmaeYP
vzlt8qSzreqak4LIIPkEvKDZXXi+fD9Yx4r7CePJQsYzG9bwNFC6b/cColid6PItn6suH6wiX2zI
U8QXFHYkiiNJTRKe7TxVgUpL0V5eKC2O4KLszIGoS5Zvxp34BuLCvJCi2C2AFYHSNcdM7cFrtrCZ
6SFGPXk7kwUPfOTC1ZGcjTbLxkdOkF+z8hkmHwJ+ASmPaBDSPP7ljtISJKyTheAeR3ysagbRjmAO
ko2vnWGqgKrFoz4FNyu+PT6yEJIg/8RVPDaANw7ab+BFnMyR9aXFHh8R+jOQpH/S7GQ3ObwIhm6e
Vxi72YvvR3QJKD94J1QjekPQaLCHP+ju0TmGXBfVWcIJaKaQePfSAbr5dLF9OfzEmxkP4u31vqHM
n2l4dPp7vKQ54TZD1KrFgUeg7tvQET4e/fv9qd+YkCppsl37ZCKUFwvzrJcZCvbSJ2OJsl20v5TP
/miAv26PP8Zsd5GA4GpluySviciaMuuBzVjlv5DKtdOQEEiIDvg1Cosp2OdwPOf6k+r5tfIau37B
3vkCle0S8LSBCjbJMVEkiNlNFT4XQTzzdgt4/c29/dWa+8hQQlINGxZKFh7mCOqGNKchInwrj8M6
QP2Ng3EFjbjNcuEAv70mR0grtesTcewdocoiOdtPG9eius3/evxyICTQ32173RnVYOG1hEtA/O8m
+yeEROPH+Xusuyzd/6I51AFH6wsZTcqT01C+EKdULNTP2efNuMa/6qWwgDfHPO9d6YqQOvXRH0Ej
QcZnt7g25dwUMO4btgHQ8ZvIrM8MvWmAxrhGVVOOKteeObHVzPGFpXKoLtcNdLjA3V8rbw6h7SgB
X+PyGWD673ne7N8DZmff75EGRph0vkPR88G7i+vx3+kqBUaO01ZxRBYpOTDUC+rS80XbBzcI3uUC
POIzl57wzAwU1Shi5idqnfcJAZq1aRc+rIE9wSrHYkrZCqeTR07ghyyGuKTi9QoAWf55/oXF9fYG
h7hddwlBrmOxb2GAjxCGwoXCshVgcJGPQmxVtekeRGD3c22YoPz8vz5Q01Ue+4EBWva2kREM0ViF
XWpg36xsEeziVAJ/KAF7ioHv4sl/wqrFH+/xCwXc3fR+1bH1gucZ4b3u6Gk6Pp2pjYEe4KSqVO19
In0xhZT4xOCdMIeLuwmh3Vgq3Zx9D/5rneXODREi1eIP+BaJk/wsmhyFSYQZH0Wtb/qSoJt2hg6t
WEkBP222z+D9OejOntQa3xbYWCmA9ADsoSsKW/jPtVJ+IQHhhg2OBhRmICtYkcjLLhgLrmcamd3u
Bkp+6lfqFINk7lyRqKxRmYCY2wG84D/LqUvE/NhviZemaAdRyL11ShDnO5b0xJ3Jn8q+uvb1jEdA
O6equc/un7hcolmGvJ3OzHkxA/cVJMDIWM04K5CQ9tYA9szGRu1YDt0BE/H85JsuSfGkMC+PF+NH
bNGKl+yo4unxe4cycXpsRdIOth64Qb1rr1dh4V8Za9hLt2RYjWTHg5Y57X2tmOZIBWR1Laor322b
cMoy8pG8HvHpSKaU/qM37HouW5+UvbI9gWrKLDpmBprQKpavzSuEVburCGa+qyQDAYbHQf7ohif8
t6kiyIEB0KmFaAuzW84ziIcEGtlq2NuwixxtP4MJ+R+mjY89BURJ5WQc5r+EqkatbqW8U748vT30
UKPduTgb7DZFaoMoeJ+nOtBlpN1XqQzMIFJyxjwPVaWE+PqV7HYLWlTVtxf0kVJ6Potjp+7KaTSS
8ZdkKQhDQSU+P2uHQwjie1H5ttpxw5kBjQOr/c2+LQhPqYTxkiFvIVilxjKe+FCDTn75Wf448hdl
EPzAGM6uxv3uE1XVVFaobNPnTgIV7coOklAN6m4396v3yfFT58Dt1DkfNFwT2kje/Pqz73vOlDfW
71w6fY6FWWi8bnYaPc+LLbKUmxAht/U3R/8d7R4m+I/ERPUnLZSdeq8JkG25d02im7cUnfC5yr3x
QGz7+O1HgH3CoGEAiJVC5XCANdoCkdne97lgv5mMBRWJthuoN/YaVe844t/hJasYg0F10lgo+EsF
V/aMFaR16PWcG6u7JTcaOhWfnHsXLvY5tQknOCRdV88lN/YMw0EcpmwuOCqx93Fnt0S2yC5i4PQ6
EZP4Bo+fyYhq+v6qXzlzOZQCIrm+ZpSVlp6N7vpTdzorJ/U8yswPEwBiwovILWCtDKz5gKGJMjds
vHR4DRj1J6LqNOWm+Q1i9QoN6TA1XgowleMsZBZcm1AiP+I4UsCxIBZ/olgClLqbYqa+YFoeGW7G
aFl06fQFs4KGyxrnVWZPUE1QgK+5Mwx5b6/H186+/ay14BMTCAcLvJGzcngQcr5jbTGEousk6RTx
cQJCeK6uaTuHFrxP/xaq/nD8jeA3qI0S6ml8lWgpnjLHSziE/oMsuOSFvof2LUje0zS9UUORSW4v
ix1wb9QECR1k9zOPoOFoYU9ta925L0a9mYCEztiFLy7mPl9VX3Vc45WE2+zYNjmUkNe8vjnZOlui
XR208p7LgdUvqUSgN59AhTUGyuzmQwjlB4ER7qepMH1Q3C09oxNVYfWulNdS5+b8MG1tS6PgNgm1
vPiCFUPpDTbjw4vBuYfWMFVQkq1rpD9wcQXvcFV3kmS0FRI+Kuhejn8JcTsvk5/6J3cy4AhXupI1
1gxwWyzUC5upmH96OtYmD8Qa9/GHUp5IOmAlxPUKKYk+Hq9MBk7Ii7dv/vHEi2RvOK0+5cCkHr2m
jBxJq9TUCIiLyRv66Uqb9zPSS66k40vifBrhWoOfZf+GfZ9L41hMPPS2MUaxEJOhMlqJm7aa+e54
i30uWgNp/Ob/O+BRKs3nsYnTQWE236cXiCUvgA63EpECMlIotNMgrGg7y5U+sP5tguS1Ydf1es4c
kgGuys7mSBe6y4RGf/2Rhwl/1sdqpxBUu9Dz3Bs09gSrnx6JuzZ9y6f/MTJ/xySIT1u7VzDYMCv4
wyszOrgKmqgjum5RI13lDKVdnl+VfyWsWOg38Pi/lNOz61krj3KPhGwJbN55/lWENOVRN45mi1Jb
vn4NixJLVrmlQdQidtlxGwnhwjP0HU+BubaA9jglYP6MO3kKD4YkdqYhNoo/jrqWtzIzEcwO+OUV
rjkisUA2BrEELNslkRvoHeooyfpjI6jzFHdE7sFEKdwM6rD8GLzmHp8auli/7INI6N49ps9zZ2lX
Dd3yQBkPllho8E1e2SeS456pjvO1x1onH6bkDaiLjmob/+sfT/Towf+1QrHN8Vnw2LyGWjMCDdoq
aEMpEYWKxYdy8gyQIuNZ6bIJYsq2WLKeRIoAXqpOYiQ68pJUcuoWiKB6jFmo0pr5MbK0lxsKrVF4
FMBb+oMZLiFZyXdKFAe/7F03ZvetSY8QVCKi7M6OkvP8A0UQ8uUd7zBN9nw1H/Qb1hb8Lt0ypohL
K/jfR8Nre1mYPMFgYQpQ80czVpPWE31SkEdtYuJiDTx98zCvcKdIPD+vjDufHbaP4AgWoLtIVUAR
5Ze8dEXxTc2AeapCMw7PqW0v2DniewzTKKBtUW50vD+BCkKT7KQEQDkOpK2m75uXbB7FxsmCmzC8
z5SgPHm8f7sJMDSOuSvP7Zr6T0ofk/HoIMvrUhcAG6Vw42kyDIKk7/k/HCyuG/Wl5+TmJABgB7DV
89PytSyJRZYN0sXruZijV2LrYwEpBX8CkY8//YfmgauaVykhIFuY6JJuSNbQtmGcDP/c6sp7aDUR
WL+bkKj76z+je7qiOLr7dwHnAK6MdnrRGxOprDMjsnFpQGR0P5fFPDSzDAv4y0QwrGseao8iByRn
RXJK1rS0+LzHZH4gn0qSVzIwzcl/S2DRjBcQSySYedAd98AFYo/GdLVrSCRs5QFWg3ZWRz/+/47L
yR7ZfMrzW12jrka99KLRnzQeOYd1NHP4Zjn0D8mgSvEKhk4IQ63hQ52fHMdJvjZE2Us4aXyMmx2D
s1TxkY8vCVdTOUou8+GQvPaHqWu7jTySwP+6Ycu5egDue6D3d7/MsbcBiagCNLF1ptABOdrtYANw
J3vvA3Jih3ZftH2jpoXDq5wNy1mI8VNBa6JorNTtmYTy1vOwn9KRzeNWIL4fpmAiTbV/j4hXKrlD
7H8yjc3sB1vyjIzsCoSGpSEKlBaA5qoEKn1N88QufrV3W1whBiyfX7Fjs9tRiV6wtxWrw+4ZCRIk
hjFhFiYObTfON2omfaRi/iwNBu4hkT/2DoPSYHH4pDwhXzEEb7pErVfLItXrAmncNsW4U0RgrvtX
BXoDspmNyiwkyPTPMwS6Yyvt0mSZ7Y39bsPO47veGrdUOUz2FTZedJFHkFo9rTC2RbzItwK9Wuwe
Wng8QGlnWP126+Ltpr1CUOPqXgNwjANQVp9himbR6PUE7Dl9YnE27sjPwl+w0csSG3HtJCJcDlH4
MX9K+lgD50MAdFurvFQw/mx8ozWFT3OJgQAhpv7g3hhwAzzKyTwODsJY3KsdUTwAA1GBXsaYAj36
SgyhzhngvRx03eIRiWVM/3l8xT2U/qWPasXbjGu1k/3xHauZw7SQeUOjWMUT6GXLP0LFAbzvb4Sr
br7ky9fRRstaSq1Z6D0VOOyt2eq9ijCq++iO3bSnB+whOQ7IZgl4Q8bt7idel/YItExjnShVKHHD
xWMdhmvUc1dae7Sq1KR7kG9XdyzunTsvBVuzz8+U9XYP6jQM4ZKicFNsJkfqJBus0uG6jHFNNSem
cZl2fhdJ3RKIt2qmtMQFacyCVtxJ9m43EbSQ6xUQyo2oWAliuPou0pO1l8ADXbWvFBomy9UK7WZO
C9gZF3x/889xVVEYhC3WAwCWpLNVNDjUnH09YZNBo9DCnkx0C1tz6vTIq5bZRaPFdli7mzspb+4n
mxU7RuwPl505d73cZFz0Bh/OLABRI9c/PQY0gYivPsgK6Rky9s4EyhQIMFym/x2UZnjLKJlkdOKE
gdekC09uz1qNwarxh7KnKu9tqngS/x0X6YP14qPc6jKy7meQd3oSyCgtuwssK/lERDBI5zUd0oH7
HoJY7oBA3VQcuV5CvAjZ+ndf8Uy6BX2YDqESxrBDSNz2Bnqk/SZo21JWArE2rFTUQfSXYCreAjoV
A1Z+Jilti2DwKa70o4ClM1tGna3uaQJHPqw/9VTK3aP2CCLLBsXiq0iemo+cHQ7c3lmr3g/mflbM
xF6G+MfYWss3IYjJNRM3SRT/3JeRNQ4gZfddV4dDNc+KBAkHIp2B0ZPmeWT4rHF1GnqZOVOhBHfI
QefiFvsz/ilLz46wHaTmwrhYLSq/GmRaG6Dv9i+kNQGtkNCQjLW2b//ypmcPatR9EyU4XuxVoVl1
SEQ9F8dOGBVDTVh2u0Vs1FqqQhVQqiGSmi0eGUwJ2xLrgkdArZNPm2J33F1JQaksYF9Vn1NhKApW
Lfvl83prn53x+iR34nVI7E8auZ4d6YNJJySAcCUHGqgY8tA9bx6ctIJLYgb8nRYiLnsyyykfXglP
bk1mEc2sRHoxCiG/zFMcjePfbWsXCm19L6g5H4cmXXaNfOkw48Zpv70Jtv7LXKbpz0f96oFOIj3+
/jfW7fM0GLPj6popS5Hmq6RsYRIgfdfxAFdRlxOzF+Hu5Yu6TJl8XsJfXVGSPHyCXtrW5MGfHlz9
gL5IbQZ4BG7otigFvLQQDy1u0bgAVUxYKoZNYR33gEIGFSDjtkHAFYIwOVpDbxA0DFMLg8UJH12u
8ZF2H8q2akPPnmZGWUR0Lw0PL+QHwKrDHK+VRtKo57En7JtD7KFWhuhP/b1OsI2ptd76A8CkY5s2
0jVGV+BhPMTxt5xkYK16ownffvEX2vtHW7JXPFzW35YdrOtuOvuvZpqeCm43fwQIBN2/Cn+uKyNP
LeuZhJW08N7GNK80hJqbiPI6Z43JMWcyiNQUbzaGuNQoy2tGn9I59N8bz8Y0cRN4awTqzZV25Se0
bcpJT552GPSwZm6zb4qzkmRSGVpm8j6HL+62fu8xos5oEOYI2hgDhH3OtYxuJTpngwrhIFWTDaSX
rI0bq8QRJiZuWjnLWWLCBTuI7Cr5mL3Ry/JtqC8YjnDzhrcwn/bgHsZgRv5zxxI4aPYiMKnCoGhT
mULJWxAyxnuD7hHflGsSV9i2WDodvkPdhfWDYWXGWX7BGVeHzzftxQrSF5uzqL9S/KISDqyyC9fw
ow4ptY+RRIHobPggohF1vUR2BzrpcPR/H8bilU1ubFHOWljwuBrPkd7vQS87/oiMA9mxbPAt4xS7
kkBTIaoUmoXliKv67xyEGQrUqahAw22a3H6lmjcaA2dl5LlbmGBAcL0woDFJqmhQbzriGJTs9Tfl
y+JVnmixt7q6f83NdM+aW0eyvLyFxEmYVa2OS1oPAReI0tlhaLxhGS9XxMJKaO2RV+Uz9yjt8Wfm
GWu+O0JQC1PTmaLUoAaEU6UaQUh1cY2+mLI1ma87lIvACzLiGeUFlf8al0v4V4tkXQdiEq4mBblS
FL4ZpJ/J2O4xAUbx5lc7RTOvjUZeMoRSDMJIHhCgKTUOw4pNc7K+Q8+UzXtiXExMvkuhbyRgSbzI
azDV2w+8DTJHi08GIGUQx4/5ciGhvppr/tqlUrHtbrgNSsWyI+JY21ThEUa1zUCUV5ToeMah92Lb
tABJSeTcxNW/F8bWwtNodgcXc4H7R0iPzkX2KA9quTMS/jVmYeWe9STyZY2svIFnVYFPcG+MPPqB
PT0XAv2P5z6fAtL5KCb/EyP1CSAqEm7uEQa6Ou2y5JrEJEdyv7qT62Ga4KVGwEtXs3jyOnV2Toxl
k57WH97kWpW4EiBQFYtXhOezCJuubSELdAvnoz0ggiySC+8u9z9p79Ber4D97x0ldXrXH+4z7hOR
vCufL2B11b2ndhMhd7Swki7hSYJEUAHd+0AwyZs2ajiFs8LwUslk70XLYZULOXR7E2kCXAied1d1
hE+t/e5ULcqibs03V1Td3l+/knh4Rv2g8eTfo0PLV8AHdCUd30987B/BXTWVPpXV+nz5SOYCr590
UCpTFhqkzfx5Epi3/IVGQz8CmrX7xxI4Ea/aRYcqq4FM4myfIVfcIg7pTY3SvV9Fb3XXUFgTwItE
2e5bftl6uaeakyur4ImGAXSYXWIWKZXVuSRmncKbLzyVheBnP98iMNtyUwR/9Zr+EPbHBLISGJvj
m8fGgtl7sryjqkMbn4ILNC4AvaGUzhx3otqjFmnjv0TRKvHYeFd8JN7f3ix6s9yOrCDIJVhBfN6/
d3RKQE28IadM+Y89uDF7eEA+YPApuPt8NmWUhMjom6Nlc8PvkTy5kOAUrCDT0CNZZY4b77umtFbh
5S4OTPbb4r5vRtqxMIas0jP+ToPo/qUu7CgA/6aBR9uZn3cwvUcS6ErB1bsaZphUm2ZxdB4lSZMn
2kxXE8pR2AYhi2Z/V4z5+xpsXOiRHO/qoQpphOK09+Ih1I+Pc29TgVUGt3JglgNMwqgf20roSfdy
FjS7xrL/mpM3hLSxaWzm+xotIbqJr3k16/vawJmzZIzDf81UqQJvzjHv91MB5Hwi+HIutK9/CPPT
kduRaCsz8XhTyBBta86EJ6KcWAlelU3JE9ciS5Q+PT96nFupG/67e8xjpLoD6pMvWA8Jtq7PiNcD
FZaZctq/XPLDiEYpB2zMdyMoioaMID1Nu9dEAPocLBHaTm89dXS4oK4Uemi+88ratxfP2kA+XAmD
79jbKBSrqFophBP8SN2nluX63NGqyTIUqrjC4/4P9VFVxK9KfPHJAt0WHKYagCahR6LwMxHPqOzY
+9M7/BIgSnLMdeebg3vUmSDePYi2wOao7ni934qiz32uOIfJnUUvqprjFrSYu1gK2V8nU2kDQ9+y
5wjwkSPg88P35SqIAwI6eIsaTfbqmQ2hzt0B66vmar+9ksD/HtDjN2ho9J+yKTOSfQEPLgGeBMtB
Vm+9/66UEFta0NQLCFVNTtLDJBgBV2fsYyeZ2/ZAPkBB+HaWKfIxyyLVhFPi74y3XwBt/36ngYe9
8Qg1P2cOlJ7fqRD7wYqjBryrrwokSOPusDJIiN85u9/TRhwc2eSvz7rzU0Qe+m3LjMdAdUoZmojZ
OXB3DvsRLr7DNgMjE2j9/1S0CiWqY9+BraTf24NWma6Nd1iyc8PvggFBDUpiiF4nLXp3j5laQlIz
1+c+59Zm38XKhHJoBxqRLzVaksytVsh1M1Z/9A1ZcO7TZ8+FhY61bNRBnpPNnHYaec2ixQJPwImt
ibgzpev7mPvf2LoeC13YPBw66QBB4bAV+Tbp+RqKHlRcUfzTd9hrlGl8DowVl82Xn63cMR1Rfgtv
rRimqFIQaSV6DsNBgsHdcqckiG2ANMF/KfQnk68GoCWzqDxPT4B0rN6o/fnnOoDSIsnqyfOYBoFY
DFmGcapjq7oVvpvYFr+nvG3qiCFDq+Y5FZ+eFm32aE2/ftbGzibuEafOhzi0J0gUsMknaV/v/C4c
pIMJXPQP5kxCIwu2sbfYsh7e7iZz9m+3I1tbQj6Qt8Z0C5UC8cihayHBSvp3/RD00H0BEZYcedcv
XoeWJ+fkr+7Ipo1FHqvvR46s8b/METVgpanCGt5Nl5z42xAdB0NfDpKVwXoGsRHxLQaLO9dz3FAM
kskAXY7tESYsHmEPWPQAsPkpvjmEHWa0aVwe/bE/5VXs9skYdDVZKTNIO+A04QnPEmd9odkPOZya
X79a30A8Nn3GugqfTORsoIN5FBArOQ7sYr9PYnyDHvsxQgXSmfHg7YwyKkn3KoLJOc9OiQZ2CXHs
pzrk4vgS2OPva8Gn1n4+KT1W63t2O14jS3XBBCtLs5FN9igBgbhnJl9r3y+xFnSahKpfcKpF1Reg
utKY1X6JLZUS36Jbdt82bObs4YVVLUCukFzCo6uK5mWxrIlFA3lKbNsjghLkTYqLTeARBccniH5g
RNh7d8CCiQjKVQvsuBf7M52thL+0FALlasqr+tF5Uzp4QsA6pJvZMIO02hSS6AfjFylOjDwwdq4f
gg8LSHTxPtrYnSjEAKyrgR+y7Sw1VQ3nyPNFKzTVsdvS0m+OOI8suGgtZ/btSTYld/EKVkZsJB9k
1jAH7cbR83jAJuSeHvyk6Vyf8aAHIvbBXeUpZTA14HRxEqShKN+39O19pKhPnrGZVY1WDn8CPk69
7R9p4Zha2V2LW9r2D6sqdFCnKNHXKAgNPLRd2oIPJ025vkccGxQRulSe0FiQ/kfiLuVpFQOBE2Ex
nH3VKK4YUOOA4ZTMvRLYjW+cUQv1jlUByvfyo0rEH0HScm0BIIlgoEV4Mdg3H766Esgl158gqLcy
Jri/Di5d8kWiqaBbI+LwvRsG92YlIKerGseKo3Dith1KY3rWufCBo4nEGgZNhBuCVJYG51DeaEG1
Y30VF7tpI0VB2iM1fvS/d93gboBrKAbZff1jQsQYwkHixSakD2mRO4WZp0NgWVwfuCmy4O1or5Fc
c3awGEyPzeNJjEQEVtD0JK4KBXj78eCEmHnOCDYXlYHbO1IUvtiomfgWGc/UdWdFCSerJuUJwwlT
sssN1uMlmalA21MNvL63Sdl2FmoPA7tvyF6tiWBEgkqOerorL+JfGDKTBiFN/A44FeDAkl9CnaSL
rOthclx+Oh1NRIL8odMDIH3ZulrD5GkxwYEEWoXJIl+lXTCLI3sKmqZ85dyhkyBdYvahxk/pZxg/
FZeQIV//KS59H4FAoUR+cwcHnv2aUmb0iZ27XIO9KvVutbdIpJeo7PNuBNrivZ2SEi8xTy5t5udi
ISM6EGQHPC0h/KH/cr9cRWe7rQeGHgNHL+F80DOpmpA6qnMpJy+yPitn/Rqsb9WbuxkuAsPqmLeJ
Tug/Yb5DmXVgi77kOnkTdNfE033j5dOdXGGXoZirf3+m+fhAJOf9O7M+3Z3+KvrIRDu50vSHG6QY
42aD4YhaHbXLElvoPxcgEghyxEgL3L0UDvC4NofWmIS19OXkFP6ifoe9hlhz47fJRRNXHuhSdrOB
k2p6pg8ctP8WngUfYMD8kwBQaDJJeiu0XybKMHYnKT/FTvZ6Wtw+6LlZ/nPY7+/n1l3ErF/kO/nR
XdvBNvSIhg5MFmbbTZ0/85hf78PpnoeATX2y0hjsUON+FHPz7+pBdb0/FtqqWvRDDu1wSpzTIgRI
nTKgrR7HvpskGeULaEQ6tVZ9eceJPYChng9vhcqntMNm47ZtUleVxjKgGsiZcgendxMfUERoQ8D/
LTOXGxT35ETYYOmg88Mx6/Bn/mTZKnocgVR4j9JizjsL9ipGOfCP7Ql5HskhZ1nIdzh4F/I/dRI7
RRKpV1n361tiBs77jWLJIAtoF1pduDSw2Fj39lSS55SKF+ANPRJbtD3MsoUCaiPm0ZgCL74pucwx
T/M6ufuuBDwi1kPirLktennVBEaSoAU59WmpwRgZZyzKNS/iVemAYx64Sb8c+xrNNg+SgFWm48R1
XGhGinb49as8jC+YeUOxurwG2+aWTJU2vX1BPfhxwJB85Z3Ao4oGgxnvVYQZWFHtHZBIOUlSS9TZ
lVjrD+VEO/m6p345KI79tvBHTL6TK2r7b7plQFloGVAWggsLkw65HhG3jfdfhe22zTtLpdNE1pyR
yko9LyMDOSCLMP0hlTob59j/IY2txfN9CIV36VHKkKaE3MVQnFK2C9KOFjgHTRSOCVqqnoi5k/Vj
QE6PvQ3cM3P3u0hsv7W/zOWnHYMDWdnqCe74nDrJElJEo9EfgE1ACH4VCbRa6x1PQW00x71fdfxG
awTI6cNKfW4C6GNa0JwKBRXhMYTzV+gAR1KoMTo9AhEqzWaL3CiXTXMu7iD7chY2+KIl9tdxJ+Dv
ZwHW0bsl0zmmRBy1PHXYGGerDov8mEarJcTcOwga59JBRAOgNfQKm5ppa6feliclL7MFXjsAbOLn
0fQLFegv1JavSd1ia3s2O1m/fJGVq4uGEjJc8xZlUPEYtb2BPdRRwMDon+AolU2ty8rV+g054p8v
Dd4qEb+M4rtUumiZ/Ldy4uKER14XWWdLFCgqTMmVYbZ4D0/qvboY00oftFZc14NwkD7TpNCZKno0
AQGNj2SNtC/7y8/A6x3XAycDq/thJyhzKBjzHM6mjkn6rahSS7PJzZLW5YMLhKJ952dphq0TlXM6
ndsVFJc1z4Z8m9Ib5Pqwx5CycAgfnwThhQ+9b75SirNdKmhjojphFbNvXjd9wOlBwTFN+xCrPs+S
qUcg2lqWhfKCU2J5H4OhniwRDrvE0AXncgfMS9ts/JfwWEC9HHxhE9TU/CETMK+/BGwODv7qzMQC
YJTQAu18xdTs8q6NOkMlnwnxXOyzzIVJqZFSzt8E91qs76tCHe0LnkA4dnT7/8A8towMruLxnvIb
5VYjjkO6BisEMU/uyAC1ag3/RsE2iWMsZihnjtHd/g/yxY1ryvRwOwEwrGJ9Xjc6gLv+dIlrZiGs
EsB9Jw2U/LT1XDYBB/kqlIcxHiSzHYMwGf6cvjV9UQwiFfqG1ynizEFGUq+FL8Am3bDI/VmoNoOB
Tr6mQvoqhOYDp6+Vqrc+jblVPDqE43q6amH3j7FrnFGctGOFA3ON4jJS6WQ5B3Y9C0rH2d38519h
3IQ5YDqFYWCBFEqIoHN8Zwd7Qh2Oyr0ThrHg4uofv8oPDi+HZBtdkhKf/4VqIy1f0Sk4qEGG0pa8
y9/rrnX23jhLdO00cyJ37bqOwS6kTGMthu3AouHqTK4Raq2dErMCY0TVHXG4bT4+kMZBrD3YI1fy
xQETTLVwgFkorBNHu1jbVgGvdhFcVhRze10qz2OunSVWQWPaBU4HKQCQjYr6z27Vb3OtqOKBuIBT
ddi+MmqmNoxZ/szlabwwmWxGizwiKBr9TZEJALQaSsMuUHx8SutbQj4+ND+oN9tm7kicR+rwfV2t
1fDcfCf58EAuxqP8ml0LVXEPc7zU6HapzSj6E872OJDLa+U3WEtQ+K3TkkhjONYnK+7Sc48kwEej
9hC4JLDCUS4W2BJgUku9EAkrTioyGCZfdtf3clinsbP9ea05KYBC1hz27+Ivbig9glo3KUaRR5et
8TEdHP8SqZugdYkE6lqMgZdGNAV/N+ooipKInzN9GkaHJJLO4BGoCd+i5GXF799m0L78qy/BSDpV
+DokasZqtpuLLLUP6LjadtiOamanuCvRCAiig+WrUcAUGnjaVg1jBSafl3o7fxZvdvw/Y7sD56MP
9MpDWN8yn2+WqPnkEnSrZNOMg2kM8wY6rPVVUkEXQ+ZVLFLPxFSLGdKZwYPnXZyjeUch6ENIve/X
l6LKiBvC4IjsolcEybonUvcSIO9nPzubxIVBEq+NPwZlEzMS2EUZaa078ckRlg8e888m79dmQIjZ
by3hrz5nRlJUoQhOl8sRlX6SvuHysvIUj0CdPZvs0w8poMRn5r+cznuW9OpT/DVc3oj14NDsgtxD
ylfNeYbtg+/CmwjV7rLVg2cgUyyphZ33uJZm8aKVMYB6Rmnsythac4Vga+WFKJJO1/99XJ3HFYur
E33e0hGkKllhLwOh6WhIcvo6b5a5GxUjSJKB8fNx0BZzF+64mh5dZZ0lXvW8qmJPHMQwG5J/+N8a
ZZp2KKPxmVUfibGEsQc6J5MLeR+95G1PgwD2J/PmwzjkdcwEJu2+TCsNFSi0NB1LxVlTlD2hV1A4
rYVdkBZGrNqLwDDjScUMQhkdB4/uu1GRdeLCj8H0DeYCVfrNl0l1iCU3m1EpqlcapjQ7bMd6soGf
F9RXPT4HoDG0R2S8Cg8Li6U0S0+jdy2BptbGR0tcesEV/JaqmmWycMoo1avqpRmhQNixZCfP2BMj
tv+xtF4EG9PRGsaoCWi5J4Efna2jTlUEE39QuDNHBYXUvgBLnw3TUuque6XT/fiRSIIZYMKqKG50
FMO+ZnSY4TsaiJgGAZME9WvtZ2lYAbQpVyEf2Mc2O0XrV/tIz5vceuMKGsCtBkSCepNvlipLWrHq
AZuV6zTiYPtOHvv6PSZsIKX7h+E2x3pNlqN1MfoCSnl+zHO4YK85lSPFnA1HGSD9AXih+ID70q5F
Ii+Vu9uq1xHo7EfDk4iWRHoQEkgSsxORJmTUgpiNn77vAYTHc/R3zkXz23m7QnwpIwT4H26XMbul
kNel8DdtosRl9yagz63XeAJSe6Qh3SbbDCBG+EZ1oeCFx+mvYWuLgwvywKtymokQr40YQPsKWhtK
L4YnZ/w8XwtP70wS3bY3j4c5lD3JNYvULS6Yzq3OhL6pN6ooe2GvseCTS48wuoTo9aOb1CsGpKu4
UeTvglDGvi0HJ5ZaIIdLQ6Ub6rmI2k0zbSNbuvbIuEN9xnotSznMsG0sdahUDNpjK85eShq6y3i6
99V2qd8tn1wIsZ2T3Ik5Gs+gKcJ0LsoZUqq7lDLLOZdEM0qDupnI54G5Nz2dij/qsuVFymeVbFCa
cn7Ou76bLgKd2SofdVMR+Y1zw715ysKYWn85jVWaIUKki+Y5Vf6/wngBwUkvYeUqgIMYNULCh61t
iLa0wTM407+ipIkm0o4CD5t4y4J49+k1NaWU5YyHmxK4WijM2e/rHptsCWLwwnxSawEIqAA61j4I
aoxX1xw1eEkgV5ZZbB27WJJZ/9TceKxTLnI1fUnspeJ1Y3AGuemnH3Qvuij44FmC/rqLoAjmTYCJ
aoPwR5TFVwvXKKJ3v1jAG6Gi6c999SFE3v+eYlL8+PkgTjdUETYqnUPyZ02m7xrdNSf6l8xNDuCV
0prlVa7ubaGoKl0LkFMSjyaDw7lkpbXvFKGkcIQrZAgck1wg3O1HZ7MBcriXKDNkJR42mMLVMCCh
DutyT0oOuZsUjaQ/1O+g7bcZ7BC8trGj7xNK0o1TA/C40fOuDs9QfDmMkcekou+TgmQuOBQbyIMU
C04KaOrnQvp2rVUgtw5iCAg0r6k/SvghEUCk9RQorQyztA21zPFjUf3Z4YX1akLJCVuTqpsXsCXj
QhgYq4k5YsR+Sjf5f+qT39atbblC4Tc1+dp7lF5dpWzA15kbukofujh9bB5ejNJWhOTKRizuUWCn
us0BdE+ZFByEo+EwSFznIwIu5+79DVzp70l92Ko1/J8rIsJaKI2BjVR7NjYzMJPIxKN+qD4z1qbM
CVrdXgQOc/+kScHjWxHNbULBNQkdyekMWjwd+LZCXcis75cbwDbcL85CQSSHTKmvIEZl8PybgsQr
86OTI+kR5VpswjvsWXXefX0Vdg9dh8oTUMebVKI3m3YZ4+PkrxZicV0M+iyL1HoVSWFagREcfD6r
M26YJR8r7geJVbosrG3+6OHTyB0tum8R3nnFuUhZ+ZcmzH41A/Ch96xPsAc3D7hfA5ACmgBTgSHE
wb+PS5F67SkiMXYBukGBfqZQF2XyZgENRIT12AAhmHJeY4mwnyZ5fblbFT+60coyM8n7WaNt33nA
HxHQoAG5XGOT1h37zjig0jx9hI30+edueRuyS9ZO+lkpU8mVuh5ccE8vx3eX81tZpmwvLwyV5tem
AguQkD6F+YGa6H1XOT/FvN4EipVP6fkFwXUVwdFpV/VNa64DHdace2OI5WhzE5T9fJPLcwXHcNWW
urtzlXcL0VuetNgfT+GhDzlTYctz7pX6+JDg9qHMDa0PYY9x4c1OlNUG4T0gwYr3G/SX1f0tF0OI
U8ULq0+DU7McyidxQqIO2YaGLFh6zzze3b4wVZ1zZr9vpvnT0NHJ1J/nM5g+Aq9ojULQak5/eGtN
fNBrNzkbnSYZPQjuWsuERWpuRcWwcSn5jseSKPV7mKZotSb5NK+mLg96y6ibjArknCGR3TpwpqC1
4a5c5GSBJBMxBOo7yCqfl8HfxGWj3Ik50A22Wk/tkVtYuDINFC34CH9Hb4Ws14DbIKSARjrxusR7
O3yLggkU+hF9tRnIjQv4KbFr3Q0jG+4fIZe6I2p7az6ZSS704c1wiPfdhyd9JadncaW3EbjwTcTu
Pz+8lqm/ityy+X8NdjAU3Z5POaiCkNyzejy6NJnaLMoM0Co6EJNaXtYL1iRXTzMn2lHaKXREplDs
PetgU1SljQSy5CFXwOtbv0BH5an0BPyN+hYnRL342yaSfO6GNJgYzoU64A0+Ih4jZBbiCLx6s+lN
rCL4tdxp9/fyWyYUPD1Z1YjOo4xqOfL+QtnE+E+SfVp5LG0na4xmRVq1DRA2rU5nLGkf6sPoxLO4
gE8E5s4Rl9wIDlZI97g7YC9yPSCsb64k1cp+du1dX47YJcBD9J/wd08fuDovwPC53sxMcpqLI/pj
pHW85ZtkLcTxVVTeqoD4anaxJlOLcNV411sVN3pHf58TDZhwH7iJV6tfDDXIt8UvopCuTx58cMWp
s8BzMhf+P8oCnE1Ra2cSCZgs37A4WUYHVmfHV5tUf+nKBLJuTs6Dn1Ex/6z165Pr4T2LhpEZij1I
DXzsGcTbEFh03GyxdBmL0M9FLQX1WjqJkRaN12b+l4oKTe+qf+sbMfUW8Z3bWgAYYxDhCoWeOPz3
LL1lJrqVEF/vmclFBjC7k1zcuY70aJ6LMR8dCvX52IgxfwtpGGssBXGioQlzOYA9SWwhFgPTOhWf
bBX74ZBvmrO8BJaTx5/cOurq+6B6zgihxCNxjRGIRtJODQEgJwkS1ZSW8kAgnmkDZAW4sdadP3TK
pSPeR89TiymfnfJ+oJi83niEjOrAwdS6rlAz8km5fcZ3aXQI40m55QpF5KKfm1mVFgzG9SBbK7uU
JoGk2aYYYGTDk4QDWC/0repa7wWqaYvqCgHAdrKBtjFHz6WqrkcUNOrQSj29wYKQkxxwkcoK3AfS
N5ehQKVhBveY1EDGIQ2irmOKHpM1dxXvTTKLrhY+rpvDE3QqT29ffBijjw4OPbia6XB6PoG9Dm5N
YrVMbGg1zCN3PHueO0XhsSMeVdy7i+skgWJQBpvgSfv4DtNdm2HMua68GL5jlB2JXll/otk9hqOn
+Mcv6g2yVjn/iqmP38+qd8WQL5hypqNESxU/7IS9LeroAk9S7lenHOnoVeiq95rJHPQ2NuCOwBLL
4djCCGTne0UA5eGrKpvKOqakweMSgkkY0T25cozL2khLjcPIe6JuLoQBrbDm1bubxEPM2hELj1hV
UEDqUOtNRROsH5VDzQ+stNIwffwoBrVWvsx8jxAukycywDbD+mrbPmzaXmdDpNIHbSy5Bv6zzC+d
eEX0+drhRJyhrvwD13icTV5qBy/0sLccnCjZKgNQSlycFNU29EHGz0yX2UEx496KZmWN445zMF1z
QPxb0vo76WXqdCiID8Nfsjv2PiN7ls9LBQSrOLfLLMhOQj3QVUyJis/xDObo12MB3aEPfdTQ5XXY
xBu3sdUXyNIPULeoC5FAlQf3/ef+IleiDTxpTOousUktacPgDq0Pe3Z8VXIvvPmh+ZL5t8qYA1Hl
S/ZilIujHhfpOQoZ+CfCf5CokwIDgQshgtmosKUuTWta8jJIQwArQRTNGZJyh/mI8GMeypzHGNU6
rTn5TK0wwc7bAFouQkBSGAG/b44szT6E1zKpct3IjEu4UVdfVhkFJE0gzhBLc1SMY8aUPyE6hVuY
ybeMYqIfHgxA+Rl0TznpoWe/yz4BuypXlseuDKxxUlH9TGHXXGZs/WPSpc1s51zSaI2oWdLKfO37
9fc68qlib4TuMGxC5Si8/ok6tGCt
`protect end_protected
