-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
qXuCEqM7I8BjNVVMJvqFEvbCWDqCJzcBI5oSAPftPmuRT+CQSfCvetAq8zpS1yPcLb7PmwgyqRQx
XneODOOGGA77SQFMrN9qoVktGCriBHDti+bYvVgZk+piPw6RkJZ2cSAauW6xmYBBcT7GvDVbWGBS
reFaD+aOoniloWqLPNOXE59qBXlu8eb3iJ0l20Zmk38DG2ahy4yEWzZY5JMTstcAs86NJjij57Pm
jh8Jq9fo7DZoRVOfsgfRmIS6/cjN6f9LDXJuEil65fm8OQHq7LtbtKPvGMfZqaTPighEdY3nJAg0
lBZHJL2eJzxqd1f4W1Fk7rWqJNAsdgt5ATfM5g==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 10752)
`protect data_block
TJJYidykpndB67eliIZMBSbeMJRLlztIPBT6faAkUAC3Md4bvHqnGlxIuqZeo7BbfvUnCRXTyEV+
YjYIQljdmIYFNjRgjKP7aPPTtQQVpVCYSGSgCm0Dbb3kaI3S/krnDtgjAjWVQTS6lcyqqS/6YUqj
KIDwaP5kIFyQVVk7OAwXnx8H8fgR8up3+25ClkLDkI8jZwrMd1ZCc5LmlN6xz1uGv5rgYmJCXgqy
5+Z1wpe6gKhxnC/XkO6TEk+aFc4CD1OFssqtjDci6F2eDZ1YPV0AmXW8c0xcZyyaV1j2+QSVsNOW
NC9Tj9/fPa1ADGPxvIl6ftGyScoP8Hd4Y/tbHJ7/a08o3PPb8kaIXsC9icNhs8xg0Wlg40ggZtXi
k2z+4fqg9GpYa8VSYSnzj1DZi75oDqJYAbnemIbwJCxQTt9wlksUsNXfuI8f8ZvWkYIAXWBHUxMS
vXstoVbOohdctlv7+rl1LTikAGD2OONL95MFAwg+o6ZCo2pGHK32Zs9AG8W/7AIoJXeRPCKkzHx/
eoK9bDIGt0TNvj323+HJaONLXbUyqYiElWnIeEaTn9PAwORMguoQnxzDEc4gYjEfkVFtgL2gZW6y
eOuNNFkAbWKAjhRRcRn6eaCIgTlIYyAN0HSJR4HVRFKv90lH5+hBHkuRLQFViMedqKFfWZ6QowwR
ZXg376vBMrT91quzP7k5ERHKF2Smd6Ct78D8sF3ZpxJWXtCZmYjyaDnfFW/RpEENuV47ppinBIcx
T8cBH96qBW9mYW8L9im2TkEgpUhK/SYN/akHDzX8kkRCpAW5zz+sgo2gk2KeThmSatx7A/4MTbKy
PMKArGu7GmjyHJl24R/x56fJPG2iDLFQyFG1G6t51gfufFPfd8RbIDSqW0dEYz6xOwSitkwZhaj6
XlyAvAiAWCc9Jt/QvcYIb9K3RQ2DdAzlxdZo3S7nJzZs1Vo5XqXtL4t10Ross2dJw/g6cshxT/L7
tFW6xEh8YqMWkHhc97rn3AeyclXKTKgmCpW6CArvbGpL3f2dBL3qztkAFh5MRwFd4NFVopIpoWCf
4mr9kyaRmHMo+1Bj+3lhU6ZoOlMRCEAzc1RGCyAEDusf1GBK8BtDck/THSxjvKtc7wC1Gwj4jyyX
xjt+BxZYJDT73xqg04W5gCVhry/569jl2UyquShza06CdBs2TQ+7JGMJi+refQ/gGfZvpTX0W1n5
/cKyrg3UmD+vIA92PDKbiGHUMuWFr8v983dZoGabsgcIl/Rre8sko/Du1hNuXeNIGJhPlqPKFeX0
h1cFLBQh/RRA7wxgmktFDTOxaOYbGgwpTvn/8Ct6yWqrfGV658MPffnvCkqbuWW4N6zen83Hy8Ny
zmz1ZeW74NPMp7Elz7hWH0Gz4m2IwhjJXd4nZBjtWMlzEYDO4tNRkEOkVCeYeP4ZsGMBae5wfRaW
4EWy/ZJ+WK5So69m6cAIi+ff4ozCQOpot14rcl7acu4UNZo6nzXgzV8uLs+ynkgj29xvRnvf4KxV
/URS5srsQRLOOR/U3c/T1lUA+5FRvdCc/wDBLN5wyH47Q3TGDQLHWkUOscggo+ZEp4OE7kbrcsMq
o8RtyK5Y8X6OX1CLwMiHhHM0+vl7xYHVxUz5AB0MZITAcFNobiMAGzdqycRbEhNfGRChfs5FZ515
R6dUlz35KYJNy5Yr66a1H6udDmEUJUXYkVkQNvt7FbPZa2AQqPt2cbPc6sIpL/g7Mp1Gyx8g8/o1
70jhqJeZOodD4UOAdOa+sQtehS8r0NTuMCVf/AWSZJkEi0fVovnvkQuKgqbOCd7+7YGtG8oO+Fgt
+1+zTd8oWPpI7UzoUALtr/23P2hR72nJ+XYoCzEDlHVbHjRoq9qsVuMjlWRjHZPb2bD/+GPuyqZQ
NLbjH6z5o0fY+OhZb3Ij8CJvS3SSn+Yjfo53auG92B4wjwx2RWbOrqhF/6gDjDohlaGBFQiFdexb
Xk5IUdwS+wVYO5zIVdjdZIepPfmCWU8r1/DRSOK5VcvudajUV24VOOD+mBJCwak0oAJPtYuEFO7k
1FW+YzZMtb+JzodQWPabfdB1GeDyJpv2rfyWa+zTwNHiu/tAlX5AQrk97TJY8fp+zaw63ENK8LDF
LatQmZyJDcM0A4P5j/xRocw1x9vQllBenyH8xsAeCmQaTh1yYfdQ3kW37FGBNz7bcchLuuPv+rSz
hnO/4lLcFpFBJ5n7EW1LaQWPxNvO8nN0DpYDoIaM5yU5i2Pqw0uwXu9o9pDzS5/5UdMsknIcx27h
hbcKont0RdFqPjWP1QzJLM4hSU6vrubVZ9RD3HbteP+17o3Z6aGmJZuilAXd4jp2kV839V+ZPvcn
qUxbG7qxg/fRWSdWzhoCi+ejlgB6GpUaA+IHhBIBgJqSHjpVipUwy7SSbNTEwSnsAVjzd2MeFYdQ
LeStWMLIxUFlwlRGt2CcHMheqxPwAarzEuKHx0/JyDL6la9JKmPRUD6DwLlAx+MT9W9SGNxm3Mlt
2xZ9/c6JbCLsN1u6xs/hHivBl6VVlBvlTofMIvB5AUxD9pvFZY9W8AY0lkxGXhPK/OdPkg4LNU+b
4Q7ZChMbaBumtzXuo0wSCvNmYB+kTagFGsaqLsgntYSGzaPE74sDZkw8ZLa2NL3WiPvjvdKbWzOA
2KvPnRL1XhkAm5SCVCSg/ExIE2yrLaWuu0w6ep962hTh5bu9E6ZvxZ7dNB+CoWUKKcAbWsmo/ocd
+XPSM8Wzs2SJQpbQRegfBFNWZ36p0d9BwCCcT8t12nQvscaXhDq8b6RxVU6fQablExZkwUIOI6tj
xXqAfHMnfMOTyzZ2PytT7HKEs/qlZgx3DgM09F6sy61+7W8ksrgK1CuYRGRWdAJj54hJtAGAmou5
6qufR09KOrHwLFzeHkXYM5bWGMmAEctcQFsaAkCIyNCyZTcmWFGiPbItuBNCeCbgFzRpGbjqiCaT
Ziq6aYOZEeR59hIYd7OigdffOT+69uGiT2IJsdTX9alMkNf3BQekVhyQpjS9e1UVbpDXzLokDfsW
SEBLWQ6WjJAglsI2c+v6x/OzpfSNNWOiPcxbJGXYPjs6whVHca/kJF8TGPtaNCfa7CwziZttoqjV
zPl70sbyb6UiL0D8xKSqzhPOw9F5nSOz7Ch5IzPoHClcq3MLbQTUijrizw7nE8s0d/wiRFD4+aiR
WZlz4miLrpEPF6RyDUH2E+iT4cXQCVLmvHbhWeJhGVHKI2yeyROa3sl21FunPYEoM/v4L4hbTzaz
zd3BhTNFvSrijRoA04VLOmeGhIyrhm1zwWCJGxnPwj1vzRaAZI7OyGl+U6GCeVDvPPywpqODVjaj
Giqip635YlMMXEgMUvw2CtcLYk3ACaw5Onn39O5dUfPHp7YgZp4oqCPlYoq82W7AlnD2YHs+7J0R
PUcCOkxS6Z3/765hvNcSDB2oyc+bZpLzMnk4N1cx2uKgBuwXXzBXUfYv5b/D6G12QZVlrphUzxYW
u7ANB38ifj5H7nOWntmKULu15vCO8M2YNeot1dsl6ZXYoSSG4gh+ptEyY68ssGi9Hoz9TkcSCYA1
flDM9HH6rSAsJq7k9SoZqdHQrFXpJoNbT82DSzK858mxlZPy1P9yun++i64Jh4B+lvt0+BAXMXVz
CDRGQded1/KspycVAVV8LgreMdun+7GV40O3aW8MaKaS0s7q0k/SB4Csur4ZaYTP9AMFFfx8wRSt
g5Y4cLv18PoXyQmZk9P1KtCspiEOc4tJ+oZcgsGpZbyh9JkZAZotMdLlbp6JryLHOT1DDxxL++6e
5uJqDqecE91cFsq5mJ8VqEVvFf8GjU12aK0tn7fNRj4o3fGGlm5wpb6PZ4RYdWoJeLZp6Bab0TtW
NctcSO/+UvfJWi2xtOE6uw8hraPdkstNnAa4H5IFZUPY6OHUXvS1bB6EjAtPSct3twJL3QKxwpa4
1dLl9n4hClNiTcgCR9Ykidwz1S1uktonlYGYNFaNd1G1uDeGDnn8o+TEDCxRmpnrNy0YtDsUSHRd
O8FeCzVBQow8WoCw/ehkLQoarElUfSDuoiWt8FlkuAgCKJoLLvh1wUHpRxqhcgswkSi+sufD5+DR
BtD7TZgzc4rqjYqMhDJEauX0hPFaui32zLX6XGSqDaUZTqr84tlCFENguF8qf0wKz1CrRkk6Qrix
3aWEdJW/+5NL6Pf4039NTjsgMR06CyDZsVBifRgbbV4seV4SAvuyDgCozUJ4e56fPQix1B+qa+da
0tb3sMxcsy86sJ9pdwkmEkygOcnQ5rAmFC9EzoLiXyNP7ERDIDEYSCnq9Mocet1ohw2x0SGnACBu
xA0BiHMqzs5A8NneXrTJ0OoKLAUHaNDGF5h0qt7pY33NOhaI1/M+DfCJ5L6t39RIbNw2R5nTGbnw
9zz4lGuZMY2kStdbMTjTuhLsE5GvDZav170XYnKBMMiKKxCkXPwkZVrSycNrbuJXHGl/brKEFCKL
YkwaS3Qxvv77WoUXPTbAhaFdrRCiHKvAG/bEwmmMjpPQKhRXy7ppab1+3HbvquhXfragPkJouQAF
ORSENx/jWVYOgbRkJV99pot3gtliLKIP0/iON8juLpyoz/C8qH6lIi2Z5zFMoBCRJRXV/RlQ+Rul
3pj7dbww23W+ae9Y1FjxQ6wUZM0PcIX5V8V/A/wx9uVZH4lvzvynIkB1jOMKMG9sp6Rw4QIdn0AW
H/ZMGsQheldoi1BIiQeJyZk5rdOHIApwOo9IHTtaRDGFJ7WlzPU9l7HepUmWG7/iKMhx9H9aU5xw
XmDBuOohulBgG1x6x3JJHI6ivlo84WkIIaHlcorpAqWOWMlNeYcV5fgaFIagzZnTkAvV24eDmj2t
sU/USCZ17/GG5TalV9rtKmF3vMYB1rKnWzz1JksKvxqubNJwRCaa6Ee/efPv6fCtv1Ed9aBxRbeO
By4o/ExsIdc4rYR1KlWt9/YN92F6qdIbFpRDhoNRXSZ8Mz+YAZgV6X2pTnloqCqFE8Rnpc/L1eUo
vQ34uCA43dzccuqWWTQbYLzrDcHD8b8zMAfifOiCha5fvXjjuB6XkdA0iOwYNdQ188GuV8qoj8EH
tNx5CdVeuJyCjpvec4xUR7CFPj1R8spE44uV4VIiGw38ydUjQ0SP5xDzVlqW5nAMju1JH8FULfFU
z2D9QeFp76GgEytgE84NBbCGPks2kvbxBJkcgWBdejirw3rT8eEiiYO2+d2edZ6dyv86JJWrJ5h6
/WzkwTr98ryPj0ZktqWNxH3g0BEkWmupMQbW7nOJ2xKEHCSApn1b9ahlYwgonl5dtH0YLs1BfqHE
aQS4wE47EDy9I0xzg1/8nfSfzgcjb4wggrKFJeccHmndM9iojMvafTGfUpRE51YBMirOIsq4/fNd
LeVC6lcd6vRGXSmxEcMc+Fn5GZbarliveFFzjILc497CEMEn1fiVcwSYwDIBKFVIDmZvXAWv/Sit
X30HfNY/MeCFhbnFbQB4PfktEIaWXtRcnRIyJHNTCVN2G0vPt0a0gibWetEJNHRw3adt6CyIy7SX
JLVx/YW5enmdspkItBeOPNrCCx0cO0y3SlEAZ3ptAsVNXockhn603Z7u6kiu59Ysc2b63qeqJxMu
dvy6dQaTw+qXnl9vJeb8iYq5THcYg+s4BTr3Lz9fgPX0MccnwjOMIuv41yv8t/zGk2/xTPpNmy/q
vh7XpOXNB/aqtY03pcgtsySO30BHvZqEYK0aV8ywDULEoe3lOenZ2ZkRA/Mv/PG7xh3NLpdgkpVR
/xDvGB6cZECf2SKrTbA7PI84B9QIV/ettoDk1QiuqxlfEbDAI2+Ovfh/LyEUT+m6Whj7DuxtibzV
GECi/sMLXBr6AD8iAt0b7UQX3n+59Cc0dt4fNl6OhkbYE9/IgHlUdMpJndUvHvV9BA5a1qpD4Wwo
chJxRgH2wxtzug1m3bkAi8elWpBkeAt3mFCAkkbZeuqIP/sIB3JOadkaZJ9HtylE2576fF9FMTxH
EsI+s4htwMNMQf3D9dav0xpxIVGPa6tHi4d5DEgPvcej94velPt/DfSoodUgjFOX0jmbYuahKJzF
x063yqnRi6DC76v2owdSt3jVrm7zUD6kZ9JYc5oUMCCoYSgkEhh90lrZInv86+1OxIKChka8r07b
83WJn+9AVhZ8u3Z8UrASA62BLG1dfnQVuh3WezWN9OZuJtOW0TYUgsQtIbtoFvMu376BJqYeBorz
iS5SH7rR7yywx3feYyz22yEdkQ1K8hO7bP/A2VZyt3TpGWbvyBswYDaavvgWnwB3QHaPgR0M1+XE
oqNmT2Iz6P+gwv0vFv8iYd5yXE0YtUJ6U59izMqFbqmzQdrhxljl15RYgYgIOj9kPDXqSVvfKvZm
suMs+5xUSMuYQdd3zLYohmRbCRPWj9NH5zVYNJZrZZBwHrL0H4Ac/i3QAN+gATPo1KG64H8RMzEL
M2GguGI+axvxIUAAzkyeJ2ueSaLPz9/4e02mdEOVvi1f/Hoelp1nFzXzctantSqum2y0z8H/KNvM
sDooKH0+oyD6LmwoMc5S2XN7kE3zix5X5u8feolOmI2E5vHOLK5QZSkYyg8uBpxHiEV6HJlz3yjZ
/JXlfLgfYHVRLEkren8a1kPYKm1JspGyct9sCADG73Ko1Qaq2hJUfPLE/cqcjNC+wj0vBkxlE3Ed
FiK3cJ1Q7en2FpM5OhotrI1EfFTwy5tR1TpSys1/q6FsGJ2eQnSPT5j7SgNuS0Ed/fYSqlC4CNPJ
cQ8qkT5wo40OZoDAk/rAFxvQw9m4Mv4zxSCVMsr0P2APmB/aNTzO/hOhY/SdgC1AfsTzgOhcDFSU
HlgTKAMctxFnUZ/1qAfs5V8uKTNV2Jxwx4QrEMmk99jQPIVDte5Xx1n0JzyzEkEaLVPfuYm3tPKx
yfPhjP43iMIC5+7+it6cO7C4V4xkWlNy0FamxqjQRkx5Sc0dD/NyvgkVlhSx9ZlcbLAkn8iRjMTb
UAwcqPpxUnlDd5Lu2qZUg64oMeMXtNb0R507R3AFRYr6sf1bPULfXNCZ5tmS+PV4hHipsvhZn9cP
s9lR+Bfd5XIxsb/Rn1yT/Hxy2X2dmv4tiHqNeuVImFmcFBt+NWn34LUkKRGntPmYHyNnvWuOJ4Nu
oFZxvQ6rTtPcwLH9Hps59jUitIgfW6+jO/S+FNB+ZsPQBa1KNgDm8ogUrGUChDLB8z7uD+8JGblf
4DoRi4yjF5nzopEnUJlfRJVIbUWugxWMrTLkyZrlReZS8pcb6WHrL4vfGMWpm7Kx/b7GbqZdRgnf
Wlja81CM3OvV7W1Elp8epvTr6UdNUOMHZYnuVk/vP8g6v/eYjv962dmtvSXO6SdSSBJLQxGrmDc7
xhEK8M1EKv8kpp/zDT7IcMYg75tYFU2fKtyg0Sozq4RKuwKTSMgEoc3/O95fc/rfpPSdjrILhE24
ss1S2rA7ZPRG64pTlCyLf/mJUQrPiei6A1FWCzBd9Azd8QFwQyEn3CSUDsehDNUskGxfPHXJHdQt
11eed+v6i6BRgZ70nEtK5+lVBW/vt+wUlpy7Twz6IM9YtDaofVSUiosa4TgwFGXT4wr6D5RPz2sD
LOOVu4736hYZNCXLqFxgYWQMm6PmSTiGLH5+CCTxRUg+vXNG9CtZ4GL1WT6iHYZJRG+tFErd3Cla
bwEiK4t6H7vAwGjXLpHbDFCyThBK7OPCkXmYy/JATnnEVhncQ4htf7iH8FAVK0cj0Izz+lgx2IgG
Q6XZHwz7lSus92/7nq3X38+j5J/fThR5fC6/Eh8XopelX9AD1MuSOjAjr783OUWGFHJkjChFaM/P
GJeiFpzaglwXthlLWAIlIeD8XlKwBxBk0pqtADLNqOYN3XpWW3ZqNPH/IMU8O0lc8zOpIHwEcc1d
Z7W8t297NRqfFJiuAPCQldDoSXBgLK18Qm5aTaitnnk7O2iFshUJclyL1S2lTnXAvbtpXNSNdI38
kEHuMNxTp4SIVGGBII51/VM4MUJ6Y6Gmr0Dh695hN0boq2hu7Q2mrndPGTjO+XkYpQn2ow+4VAlg
dbquatNiZxUTWo9nUHmN88/KQ9gavtXx8vsgsGO8Zkc0TEVg3/06qs9IqIQjr3BzWJuNbUU5ybhn
RPlRNUD5Ll5f2K0XWZngEPnSGIyP3w4mVm/KQogPneZB9OCZ20cthmmGTdJmig7bkL1brpZWBWoY
KJSABkC5SIQ+5bj0Wzwl1ZC+VI9Aja7wHKHw+3Ty9gvIekv2YKB/Gnco7gl3kAQZKh6X2s/wnB4Y
5nJNhXHP1jPVDVVNl+aYATKqe1ypKMLkNUv4uBXtTaKTppCsEW1ehGiEuTVahkf57jAFlMUdu0gX
vXq0golapU+aXSbgtDEZuTidPyzKqUY/h5P4K7ZsSKIvR6Sl3ishHPA/b5VUBaaDM/UEL7RUKU5p
qBngOiZbyLCKnsfocGKs0rSboc4+STG4JPDdBQUrnYk2zpjWLtaNY4g3xKAInsqSeAuLGt0s5EiR
0RphPlau4p35Gq20z4s0CDLrIJY+rijnZ/nRFbCDB8yBJ/3BpmgFEucgEMe2xdU62jqumNVXcvCP
60SmuvwavCo8FqZTdDER4TUytdlpM0Bnpz+K3iHcLB1WHu+YjOyPJEwmvz/7YL918e1f5p0X1RAb
xF0inIe1LqzVQhJAGzaMT5fWoucin62fKaE+Nh/s0bv4SrNpcyqpGGI/meglt/yJnwcmr0lliDXR
vmEqkfftKLBotC8Pv2xfGkCQKLB/fCi76L23osVqmFXWGSX9k00akqcCqBxTavV1IV5nmeGU5XIx
eWJhzP+xpQ+jrl0BeuQIQmXLvhcR3IZo0M0FR50DHEYT0bONdCtEcq1+IM1rX/FP6vZ7AhRRLTIg
Lny3OjFkHfnHd+z8y6OTX710XT/syVQvF/RVSc00+kidVrW04pEk24f0p/WmatOYEQPNavRV7Ebw
UMVWZOqTw9Fz82tu6LnAwC8t4j1ZZuRkZdgkVhiA6sS5SwoyJAjGH8tTtlf7vhJ+tSe+LS6MVagL
lWfNvy6uQyb45vNTpBJhPj9AtXJeY6nYhWZ5UIl6QEUR66U/vvjLXavyIvJghn6d1iUNl4OaSiDv
xHnSjW8a0ZPVW8fpJfsNdcstyogrAmRtZJjwbcpT613wKD54eDzkl+5/ztXVYDxMLPhULuyZdH8P
RrGnV4ZwSToj8l4S8v5Iwe2P6xHd+C6u0LDt3kMnZQnxX401aqHLYL+ViMoN290PZGtv9XgvXPvB
xGElgRJ9W+t2qn8Y06aCsfwEt+WaL0Hh5C120iPBITYDi677Mo85Za1tMZmcNChvtMbubeLMcf4S
a/s/uHDyfNy/ZQBYW6H2Fqp6n1eo/QDq7lMw+ejbOq7PZn6ZS4//YFnzYN1rgXpeuIel66f2GN94
rJ7Ta3AoWldOS+kyzX935qHUq1/RvBApTrSu7txmZjkKZC28MNqs+SWxLVJoWpxU05J2YAixMPhM
xB9m6oDRSdL6OI5Lkdkfy7/hchsdRFFqubGrwBu4vWsmR0q1Wj13iMW8WMVf/e4BlTea5Yj4VIv3
0ZhvnbFR5m+kLODzFNycv/aQQTX9/jQ4j1SSxW54ghtoNfhcti5o86/VvZhJYCSqkEZsWk3nP6k1
Y4YEpdEfznOl7DS9jRnAVCHdKg+lWpJU6kOPdkSqfrSpRYanrb875dzZIfLsdQUTiCYTp3rdkMob
6uwVVIk2tGW8zxsp5EFS1pOCD115Kvvx0wqhXi00IKWXpndEMDx95YBMJYjFYFFDcnn6rM5ozz2v
q5QYfFciMfZ/Hb8ZlCRgsIQTzum6Cq3kdy+iVqShD/opNo8nD82iL2O9B836KCDKQJ8UBQ5tOqOC
TI/t2ebyhS7pOGMiep+vEVHCgIXUSWlgxpkQTVEjkpOgt/JUJyns8j/LUP/Mmv7Fe5SvzEyKJkO9
2Y6yf6arZqdGUmHF8wCZbFwYxp03dNqA77QCUSD4Xj33VC8WusDj38WeiYYFmmXLCLWU8PKoquTP
bG52KB73J3Q1NkQK1ZShv7mxyZWAdxtZF2Iv8IGeK/X6s/ZU6eLxkUYH8UiHDJpqWXjvgZe2D3y/
vxbPsRfF8JoGsWLl6meAA6LgNp3mdh3EEngjbqLXyiMaUqAUDJeW6qIK1WZghmWxy9d3NMVsjXCD
tW4dRq6SPZ5GHgKj8uRA6oTBWJoQxYgUTBGjWP1i2LVoFA8GjDSK//ZFP/Rku33PyD2hoHPJCe9Y
HuODqOGKy6LmCvLPUP7tqbz8OKZZe/I4yZVO53OMFI7L/Qq3aXNx1OCl0HcTDkkaJCSMcCusSF6u
ZyQGDzrBUTgnf/mN6GSFwP9+VRdpPlHhlTKYzuTvAg1/9E92NNnN07VHBCWqHTz3ndyrSLyAfTp3
nS2kNLN2xbgQNefeoweZunU0GhkzDHD/2xrvpLshDoNSSq1XgqVxM2eioYF3u2DB3pUxe9+Hf+oc
SM5aCiBKuKAXZiSlmlLCSRGF0vMiD2p8QAxj7jtqpsOGcvoA5fVCSrdUtYMnu209UBsKrwj8CX3V
GDio30B7G5BDBdQLkXsm4teYGqMFCUpXhiiTuTvBtrTjSxhqi3OInuRvbTsYyB4txHGeiu7UPJbb
5Uy8Wewrhz8LH9O38BuZLuqrrhZEAtJjCKHyaVK46+N7irfdP89Ssyy6cyg9JFAvPDCovhZjQZa4
whwwlxKpI9ra6GccdUyIrmxf7aTkTJYethXNOkY77qb3+kxtF2t4XE+dI3YMwUxcEpuMcR41CI4/
+pubG9gt/n3WIg0zQkCZXNLbkRsjh2yRqmT82OSGqe6uluRphUMNMnj3CYGkDLJnsWukJdQeX/rV
nm620sVf4kg5PeveSBf+DzTy6xoxoE9plyCWMCqoD4BSJEl2dlE+myu4rtTzFBd9grbdWA250kI7
EoUQ/m0kl6uudWwtS4SP39HgjTegKquypbE+LBrAjrbxlIFR5R8cne6yFqzfXy0B1w39W/pyu9q2
u1qjbM2mnMrigiYH6KefpJZUb/If0R/aGQpN09NXe6bbwH9AGy0s2ycXPhOwYF3g1LuU4bZgW/LT
CA/Cgd1IRH/enbeVP+IbR0SX6q9eOqOVmxDBvkg5DTdNVbC1D8wveo8rL8LSWDdP53ZSjIo+F/X9
u4Bk+30sJTCCpAVmTyIZZOFf8tjs8DvOnKyCqyj1da30fE5YBmYYEQrXlKwvGj9Qwt9kNk7u+Rti
qJB3M12/57xZ/HHatYzhdo6VrR2FIovXc8qKbnsygty4foy6ruVbxJ6qxbrIXxOWJfiJfeWpDVI5
8IMKNaQwrz32CfklqXUHnFKDtR46hjQF578Pj5mfSoC5vhGcdaPrFsjRqe9TRLDHaMPR39tDgvjx
RC/CecYRQ7fFtBTlBFb8llVcAcimvyi6dOhRgvIBg8osdhfKnclqy5mkFwdklVYQaemF5U1ftvqf
n2xqTqgZOyHOUbAT2QBeXdCi8fVmq6iFtdww8/BlR0UtXh0uZ4GrF1aYKsFTIS6vBcTvr+e4RyIf
Hgr5it8EKeYi95Ej6i0gGDsBdcE4m7DQ9IFxCKo3ofeucOhu5alWE4wVA/lrFa7YD2LT9sn0kTEX
JNgvH/mBj9zAPJ4ddiZbvM/RkWE0BDRAdmdbl1sVyrs58RS0DAyU3PQgE/uqBi9JRlCL4PnWtg7U
b5shIoHLf479/M7VzZGwFTnC/T8lAQEYp8Axnb5Mv+4g19GlR+kSV+FzkXK1CZsZqHIZZP9MpwYl
gKN47wGpIUu67h6Zg8Ja0HiHV5YaLeuMOtKbvY0Si5ZT4DOEJjiyDewIo0MuvEuWdAsloEgffVT7
/QAQcS554TcaeQKeqmrcrOcDmo9WE78oDvf41LRKCjQtpPbdhlrdn5LHi0tZLOYB+cOy+nffy501
xqbzQ7MWL9xzCmVDlbC2v4+OIZpLgXQfBlnuBWYgvjJ+WCsyQwTav3Qqj5xTUKEz3h57Zzw1P53S
jStPmsR64mnvsHYcUS+hIVsa/dJTEH3qCsF2B3i/sxVwQ9obZSb+4r3Ezdt5Kko18t/DIa2p5Fif
Dqnh+PjQaGOTeqXqtYrHhDsu8hwV5jWnX6EOJXYI/ysOhqaeWsZQiZmkdvp16w8c0MpI8uU034yf
zH88ifXdRqtX0/WcURdYwLs0c/5/WCFl94dPJwZ8wjEKF2kUSaho0cQatJqauK3+gdl40m13Dhlj
vnnROnTKMBfMj/+/8d8hqaG2luW67ae4qEmY3do5SavGshV3E9RBTJssnhXyRyYPhVPq4QufyW8k
XxO0pProg7k4ll2gSMMg1S0R3KT6yGlVCcyZWv+3POcRz8xtfO5MOpbytvO3Rh0MuK5h+tWI2YCB
d/YJZXg67v2yxugFB72DZe145O8sp2kmWLXme1UkMm1PD01YDhp5I5XKnfq1MbAIU9NopE4VihTK
3movkLl8NinM4MqYJKG7n535+S+bIci5Z+bjA+eFcs2hYPH2BwmbSngp/s03je66qZuP8oTu6cPc
CfkwePHXvgQoBc2pi1ysKvucv4tifYWuou/Dv4/shl8G1h91oMA1A5iKk8hfTNzx6FvfnvdsdNP2
4DHi3ki3J3vJ0QEyd/7fpU4SFxwVbGdtV1n/F/pPESlteD1tYze8zeNsMemhHVFigWr82eSMZkTJ
FNQJB1eEXNSjq09lFbQTk731VzlDq5PRbA3RZWBTXYDCwYMLpvu0qpzmk2JhfXJlHKOOBoxJNLtd
axuBebJITRg2WTC0pnjGs8fJWkd5dKd6V7e+hCLUQ+RTEUysae0Yx6/UgAgaHQKUNJHHwzs+mpV+
W4X1D7DvFJ0+61l145BpJLRISN4Sgrob4FxfCCDzmIJTcGix7bKnWi1SOMD+M92RxrS5kJHru+6N
U4CRmmHtB93rPy67JyvPEixbToYoIYSpU3UORPquMUQmmGOg2vcSOT2IXStvZkUnsfpnEmv7k7Vc
oSywO07H/ysRUTi3r3tRdazwMwy0361px1VaFiLp4rU2BvOV/AmkS5w+lcMuWWf4c+tnFAK6lRor
bZ8aIyq30K008sdOjJJFTRiU6bxkyCboKi37vM9GQTzc71z0m69+C0nf8at24Z1/1b5u33Ty3xQr
50/PqOIM9SXWEipaY1Pz9OXtUgyFnU6+518tbkkdzEPlyhIo4GDz3NEZGCgJgg5iQY1/LCZjmrk2
Lnch4+nHq5GF1ZO60fEynj8EqUbiuOo/lIPlGaXYZS99xQcYUM82WRJr60XxWDgDK1nFeLL4JLbL
ScaJVFOTSgi0ZPl9nNks5C+Sd3Xq2CkVqrtktrsfGmwSOB2nTNpioVEnTNpy2j3ZYXhmwO0FBPB1
k6T5Xy06ql0tcJFXc0qepMzBkciNcREOOwtqGYSmxdtqBd87I+drJ+2D5Ir5g86Ka5a0oVfrjwEs
W50qDJ8ZSqkMrpR/nr3QHLDi/SWqkXDjR4xeuAGkQX5L3dgJvfbfJ0QIeDHnJ3HpEk/lK+dG+TeK
iJIS+zCFNuDFooJ8Uc0PdKdyF1VRe4pFRxh4h5RRTZnfacR4Bh8K2LGYxfdD274/Kqd/6QL6sUez
X34/AtCUE7COiyfiyUEC3JvOCswjRmAYQUohJT6dpJ/xgky1eCVtNMhToPmZ+K3juiXmpChY2rK2
rUQMutYyH/pZkZ5ZeSwlZKlnXHU8ByDWE/ZWcArO1lkHxPI0XIRt9bbuToxCBn19CzKUIJNquI41
0+Y3FI5wzlPYTL/Cqtr/TIQMGYikEfcatIorLmVxv0u2U2MoYFP+1K8qaWMG0D7YTQQ6WY7wGKVc
BiaRmY4+s23Td7MuyFNSpSE6Fzbkcjn21VYbU+gl+2TOZFS/Od1+NIH0dvgBTYp+cZeoYYHwqUi9
jJZLbNNbTe+0fiyipuDU8LxuLSv+C9Rg5BIN/fYVvrXqdZjdu+bCK0/k9VtORKwyxLq2xQhJJZfT
J6fwmOxD6araVwq+uuuVu3gJP3nFASURqA13O3xASFewqTtd6W0w7X30+r9Zn4h9XBqzQpDmf036
KEfn1nQU84qhszO6dZGTVRnH4GK0yZ9Z0RSS7N0aaqZhbaAidfWbQ5YFfcatrokYD60JBSBZVdiz
1Bv2LyVD1hp+lX7Km5KNEgRoATUZwzXqz3cjAppBFjjAl0u1MB31UoB9QJp8tPRWCwlJQi+qqu9r
wZ6OQx5svSF2cUOKVWMbn9HdqPIXyDtVIjgCGNeLvnN4Euj5E7iw0QnXpavWFrxF9qJFkliC4vdI
whTNk1nMVfsKWWMSqqa72YBHRmJUtDZvgchBJBLd4nZ7t/ti
`protect end_protected
