��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$Rx�y�<��wA�*;�x���@�̦�W�X�fa�M-$u����n~�%���P�$��W��kYَ���P7�?UMfT��q�6�U��k�>����~�\N�(�����X�e���/6U|)�X2pF�]$h���d.���9E��WG��L�X"]�Ad����ľS���8od����e�GT?y	7�������ݵ�^��R�q^]�鍦�����s�ae���h��L��P_���ާ��YЭF���'\��68�b�[����w8�[X��V�F�0͘3����q諵�uW� �h�u\V�?@��_6G�_�*�G���B�絉�f������[�G��U&�����~�F��AׯK1�`c��[<��FY���4I� �#�G��x[X�=�Q1��`��R>(�w����R�O�?����7�,(�H\�#h(W�EH=�������yq��Ѿ��aF����:�U~m<|��.��0=�P/���4ǆ���T(���(֯��D��ф�.�SuF�O~�a�=�e��ȿ1���#��h���?��k�Z����]q��yRt���鼿:i���+K�H�eO��
L���؄����ˀ�4Zm˜\D�;�/�^��A�,)M�(�Q!b��s��	�#à��P�Ԃ��V���zs�9�QVq�7�o'�����1<Y,�rL1E�[�ڬ��c�&�ܺ��X�B��$Ł"<��׀Y�/�t�����oyt+�I��&��tt,�dp�(QR��R�>�����2��Q�`������30�q&:i�"^��?[�Ci� ^,>@Rl5dR��������h�O7%�O-G�avb�o)� ���7�]�?�u����Ų�hDAH�f$�W�����zS��j^P����A���v{>O��<��$�u�N˗�������ܓ�����:Wc��pql4�J���>�n�w��
,,��_���KՋ�"u����"M^��G�)S���/�B7�y$�&�jG/�E�p��5ϭU!a�-Fq{O�%p��n�>kP�m�f�J���(�������Â�6u����5i�F6������HK>�?��=��(��^��(�NNM\��q��>Bm+u���FG�xo##W�r'���KiM�����I�]'�۶MY)́��4*
��W�]M�^p��*96�"�{��lq�XX��z�E6$3ur謼�E����*u�K�	�sF�
!D��V5�m�b�ڂ��J__�vg�A� ������#�w����@U桜>���2�Gc{�]2%&�u�����/�}�y�	n�v?�T?��؜��SK��ҹxm��J�h����gV�~cN�j�Ļ���~��������B2Πen7S#f����3�8��ņk�!X�;�i���fLw�$��Z��Z��^Z�8�QaM8w�<���\e�3.T�xv �z!ʦB�c���t"����J�稵c��N\�l�[�t��܇�������&��qE�wIswE�{[�E����6�CC���=������~)!P�ʸ)p�����[d-��Q�P��-���l�hMP����!��#[��t���8>�>�w���_|di�I_Κ�lz*;�6C!&.��𴐚-.dQ.M��|)?2T�`���H���w��c]r.�*T�g4>�vD;Kfi���|X�=��r��?Gv]�43̃oN4�5=}t��|Sy�@d�r�Hys�T�(��w�"�6��(����{K՞�l��t���2�&��?��?L;��&�V��O�hnԎs*�:�	.�0�s�#�����@Dv���|d��a�
VdXy7� Z���k��=�J����.�~kF�q���#�J�\�/��Ƣ`��g���%��$if�+��g��of4�ʹ�k�aB�W�	&P��taZ�Ȍ"�@���CO��	"M̒p YÖt<�mN��Fu�D(.~D��x��aa�W�m�7��B���l�B
a�z�~�����".�C̑Ɏ�2�9`�+�'5(�du�z��f� h�T��0�F� ;7�\�HS�rt�J�Y��kU�M����	� �TÅ�헸1�(��.����p{w o�{�����x�Fk6����#O�=5g2�;��h���=�9�a��U�_������_'���'���������l@��~t��\�ֈj��8�숺LW1FTR-�Iʤ�,��2Ĩ�:V>�+��2���l%���L	��\8���6��Q��ߥ����Z��v&2��w�����g��U������i��ĽA��&Q��-�M��n��C�l� IF��Eقcȡ~%��p?��A֘�Jgح�R-��1�-Ua�KB�d�lUH\-No�:Nb
����	MءW�U��D���f�ӗ�j<�&�������<Ũ�3��=Z0�J���?������w�7_�����^y�^{�-�q�ɱK⚛�+��nZsA|h[p��i�*�.�J�G��_+(+�J��\�O{�_e�@�fϖ� �g��}��-�j躓�]��&B���~L����r��qrz�&��mG�ڊ��0�w�P�R��f�.��;Xe��|2��p����c�s�+�b8	Ә��ԫ ��a!��r~���6��o�h���]����$�[��7�[�@A������;;Be�L�$�ٙit3�
�5�������[j=�uK�zR�����c��'<��nK-��^XG�d�Nrg�4K��&
+\�Q�Z�)7��K1�	�4/#�9Ǵ ���*�QJ9\=�%��Ǎ'H9u�������eNy�����9�l�	���z U��1%�:��s@�Tݠ��z:�����~N<�NQ���[�o���8��Y�B(�<Q����u�2^L6i�'U�B��Zy�ޢ��i�a�a_��)Be��6~�gQ���&B�Zg_��E�T��I6XǬ&޶�!����f��(��+3\2�2ߏբ#I�� ��4خC�Y:�?�C����=��.8nu��0D���o�Z�C=��$��r���O�T��	�b����:�RL0?u��H�<����Ȱ{~(����{�`:M�G9e$7=���H���|%R�Avp&��Y��et�f��!�\���@��!�~}��l_W�
u�u��C�ߔ�E��v��r��9jA�r�uq߽PP���fm���2.,z��:��=㕮�ZPA.�V��K����A���K���h�?p�[]L��������J��*���jr>
#-�����xj�(^z6%Zb���B�)�<6}���QoS���-�(��=K�?���;�R8`LV�"{����Ve&ִ�P�_�;�oxd�>��C(w������!�b���#�u��D�t-gv_�jH	c���,3f����G�Wю�_/�O�yD�T����Э�ě�q�Drj��6�/1�'�N\AgA��%���s1�y�J���c�
���x�h�q��͉C'�;>���^��{�ɟ'�I���c��s�����> �G��S�Z͉��P�����BG��'�=6Tγ=#���'��p��=���,�c��2:�����[�x)�Po����ƺ���|�obJ�J����D[��S��{\��,#�9F�hC�fP:BD1	�c����Xl�~���o�&��"nԃ5+$��ֹ�:@�5SMMڊ�@"Ji�BK�'����Rk�މ/-�#��5P埝}��ޡi������{�Ë�T/~K_�Q������6Q�����k�^7JfSb��<)M>oS���|W�ߧpe2�N(����߇���Z�v�`Gh�:8u�^/����ϛ�o�*���n�$+�����j6q����}�+n��j�5w�?�^�%_��yݦ�>��c0;(��pD^�e��6?�����!�؋�GЄ�`!>�00���%�W?@�r���\���mO�.�U��7��*�Y�)W�`�O�D���4������)J��l.*�jBh��^�q� i�*5ʗ�Q��8"�׃� ���Nٖ��-P�Aōl(��d*��ɩ��p:�B�����3�ܕ���'�i��([�m��i��u׈�a����j]���>��,N��:�T���}M�Et��"r"_!��Sm{�쥈򥏜yJ�in,�qdy�,�p����S\M$�||c%��>������¬ǵ!�a��?�L ��J���xV��À��<�M���ihNch	-T���L���CT�H��D{�~[�3����!�\��5ȁ��Ecw�1��&J�[�hS3b8����5\])I)�k�g��I����5WFMU�'J܅`�߇���0��S_jgw��?�[�#'���'|���?7� m��DZ̢�b捔I,MYnL�5�؛c�������u<��U�w��SK��x����8�E\k����Z��t�{��@�6���lu�)�Ʈ������%�f]��b�7�ɘ��F���C�Y3w��3�]}j�)��(�y2gB?��	��O^��H�$��W����e2A.��Z�0`�1+{����=�1�V#<�V8���l}z��+> Rm�O͗��ǆ�}�9�b��0T�g��?�����S#�n�l�8��f>�8�0��l����+@6�.���2���I_s�Z���	�>sVA��OwH��Zbê��3�Q�F�SA46,�e@�#�.���g�tlU���h[T3Ӝ=W����%��;_�	�-�\7�����p��s�Œ�]�Y��;b|/���R?M���ړ�	 �J`�'YF�����^�/�\�)ft�[iZ4t�������k;g�/b��4x�E
����ށ�n�>��	A���>���'�N�?�-�L�:Ќ'���nH
�zʆ�����c���ʕItb���#sd��{4�U�!Z�H�2�=!�jr�Ch+�d*p�24�l���E0��B��;絗����f���a��\e.i�e�ݽ�=ɇ�+��_%PV+)��)|��:���|pK!'���m���pzB��O�S��߫]���Y����o�%ȗ�\{��IDfHz�J��4�"I��H��]��T�������Q�:Y�-�����a?W���z.L�y,؟~T&S������5
�@#�@s�'�*�m����ʹ<{�R�7Nu�v�珌����&�%���t�@ܾ��d���_�%����`Z��)��D��`����dEgT�F�u�p���O�;���9�&Q2��6u?��W��p�Ώ��+M|��q�4����(g&���c{�.^`;�1Y��[$�$�}��[�"���	�]S˷�0���r�^��gֱ����l��7^�[YQ��.4�jil�����<Q�A�g��g��Nb�Aن�:2I���A��y���u�E�p�-?X�Z�-�D��1��<b�o�~I�@��EB6�gж�Ub��Y�e�$O��t;2��!�R�"F �V�_�ґ�{�W�%�S������P����-�J�S�c~�����.?�<癚�+���0b�I�c������!���M��Z���
FW���J$���.�+o8���X�m!u�D��@Q|�c	�[�%����vd#3k�\�Y ���6���z����9+��6��'��Z��2}5���|�dS�_0+��ao�lْhm��zpBy��I{�	��^�������n����i��l�笘�A~e�I��_*9���d��l<9/r��
��������ݢ�Z�͸]��wچ�4R]�b+��je �Ux�+��-�L�e�WfJ&Òy�'=&Qaqti�<}Q	�C3��H�<�5Q�� v��;�@��&����uл�`%T�z{��D���q, �d�J��L}�Hc(�yY{���;8^gÿH��i_HGv�ߥ\Lpas�Ȱ[��0��f?ȋ���������?�.����#R�c�e~[7G�ibur�
%��+w�,j҆o![N!�9dъ{�i��b$�ڇ�"9��@�䇭+A���j��}I���9g��]iro �͠� j�nA��zI�&�#8�8�k���ʂ�j���ө+7�r��r����T��+�����/Ul�vK=�͐kW�	���G���Bl���Ȑef"����5ٲAR$�FV��S�*�2�j]�j7o̙"�c�\�L�S���!�.�/�Ǎ��"Ġ�k?fT��{�ɋ�!�T-�a�Ꮟ\-Drd�P�����_���0�4a���:`��0H$���::g�j�]�/�*����
��և�9�@�b�;�=��ě���᝜!_4.�p������1��FyM�thHBu���ܗv�F�+n�)�cF	F���y��|��K�̿�Km�����g�*��F	�|B�J��VGt���BD�+���W���d�I�W�&��k���;��6(Vo5s��4ѧ�n�S-��Zn��ܘ{M/da�P���ʖ#/ �x�Ͷ8��?�B�]�����z��؈����T�	T������>]'Z�<����3c��^N�ݑ���;�v+�>4G��~�Ϡxg/ ��+X���qE�Oh��W!�Zk�mr �>��O-�Eɸ�8�@[�+d�ձ;m���m���-~o� �X��4��)0�h��!	陏W��tp�H�OQ�tC�zJ�B��'1�v5��__B�yY�YkG�.L�Njː'_�l0C�A�{q�_��	"��D'�?u�E�����ʍ���f����1�����1����Pa�&E�Ϣz�W4`��	D�� ��`Q�����oSA�b��_ݧ��D�:����ڍrP.s~�՛q�2;��	3�$�j�6%����}�*��6�"�_��?MJ�3��Ec�x!����~��԰,{ז�v|(�*ӋD�U����]�)�)O�~�s܅��t�7/��I܆#���k;��Qx��n��J�a��в�m3�l#��S��~{sS�ף�k��|-�L*Ɛ�$�ù����X��`� +Fhja.]B���[i�)�Yo���n��9��(�~�*AbV����"��jp����C�؈m��1�eQ�$e�Yף�#\����/��ϩ�ʣ��a`��Y���1u9���~��ۃ���Q�#�^�1ZN�"������>e+�:.wg���|�:�> {�4p�W���	���a�}�j�^S��#̒�X��s��z��qJܹž<l���9�K�����M�����~z��
�,���o(̴ֺ".J���O�G��^͘!��q������M��G��^�������8h��Zd3��"_�3*@��%8�w�ԭ��=h~x{��B�@~G�bp�ݜ��Հ�'y�� �E^��mH~=��F�Cn,��D3� �2��;��E��FѪA@ֻ�Vhe�OK?^{�%Gﻸ�-��|*��exReԽ`�����l��>u��v��2�w3�.>܎K���j(8��,���E�i�1�� �I��>�B���<X �Q)e�j�=�Z����fl2ʩ�.�S������X=Nz��*��z��=��JKT���+�l�@h���*��7z��45�~'����[��&��Z���ˉ��~���Y��x$��m\�u)%�0-�ɕ�pwh�I�Zʹ��4HҔ}�{�f�s��g;���и�j͇�baO��9�6�h�t��a>,�1|�����"�W��Y�wi�7~�����;A�ͤ�4���2����e�s89�Cڌ���L�MpD���h������X)�G�Mw�߽�b�s���ԅ� M�@�q���S�^��v��'O�w���Χ�Xk\�]M�4��xSV��OfW<Ϊ��X�2\�1����G$�����G��|�v���j~�.��ڟv�P���'6
d.3�N!:s����v��p*��ă�!	<ߖ�F\�2��@�����	�>�0����}�z�(`����L�J��̳��֙6�*@��F��ʊ��	����k >��0��K< ��5������=�a(�Q1F#�k�1n�;��v�W`(��qZ"8T�F���q�D�o�ǥ{�}�{�G?���3&���tu�����!Sdr5���y��g����ȕ(սp�2U���1i��Q�Rb�ļ�A�i�Q�v�������9��Gj��|�@ț?V��ź�4Rۂ�Pc�Y/e/#�e@D��溤�l��.+!���G���'�������+" �XP�I��]R�%k����+�*t�ǡ�iM�&�t�ġ�	!��W6�����9x�;��w�8Ϋ�5�-r����MJ;����HX�}D_���@<��ʭ���*���6�>�����V�]���Z��h�Ml��|k�c�P��
�M��r�#�B;���H$T�&I��?̮�§��P���С�J�848���j��g�IդK��O�8B���:_]�F���2�w���]�E+�l�+Ь𺧬�ch�����98��tr^D�qǈ6:�?�g:]����_�'#���7E�̹�2�j�:@H��[D�;��c�G :��;�̏SxV��s:����Z�ݵ�� k
��.	�N]Rl����w�����QVbC�c�Es(�����V�N{�|�Wk���:g�	*,�$5�=P�X���v���Jvj,=�{g[d�:��a�'`����4Dpy��G~n�?՛i���dp��%dwd��>���{����K�݆h������cI�6񲕒y�����Gr���Θ��bT�
�/��A����M(�sA\���XA��,z�F�i\2�{��J 4,�X�"05Ya�o�ͳ��Qk,�  ����N��բ��a:�Y*9�w8Ƅe��	�j���7Q����R38��E�����(#�r��2�ߐiq�7�LL��Q����.�Mh摍�U��3�BO�����K<'oMT�v�j��_AS��đEc�b��*�l��^�e��8���u�'�E� )#���w�֣�$�d��P�ڇU�@��.�n҈�dj��)��VBlAwD���y�e�s����R�20G��4^FV�����+^�%?�Zp��)� C�� ���X�k�5}�N�Zxߗ��.����;����a��"I2qE�㲿�� ��iuO���%u�Q��h��9���)��]wƽoe 6��F�S!V������*�]��l"TEf�>͢�|v����"�
��"�%����F`� �}=B?��9���%���pM�IB.��9�{r�S����j��
�j����*�H��%鑤9�������0����i�E����&{h�$�x"i�$270���H���8� ��,pji�6|"��b��l�����QZ��ũ�9 59E��H-E�+5 ����u��YQ��~���鰬F�u|��� 8Tf�Q�S4'Tl�4�t���d�⹏�"�E���$LF臿"�D��}e��&,'��:�(�~��t�y��"q2u]���˓�W��h�����i�ÉYZp�ֻ�h4��&G-Z�Uޙύu݂?�qp���$�6��+���Х[���j��k/�v�4lS۴{fh4NXzbD|*G]%�2�3xn�%�z��&���?1�̠z����k��h�* ��z�o�j�*��0��.�������&�T��]����T���f|U�q=}N��Ѭi^z�D�QM��z�_��b�"�W�ݫ��S�u��n{���ZQ�Z���h�L�h&��.K����,.9){�|�Q;��ۅ��ʉ�D�,����P�7x�A��tXs	��fp���e��)���#	������?���k�u���c�6���2��#���� >���/����|Sq�殍�N�o+]?�G���g�zӱ�*V��O�+9)՝��X�R���db�Lv�G�*�7����ʊ����2s~�Yf6Y�6���4�7R+�8�t��X#��d��G>�od}#�p�5���+�n{��~"컑A��;z@K7}�9������I�_tT=X�*�|��ile:�a��?��`y����0R�%�p�p1t�Ĵ��R~K�d��t���	[�G���ɺ��j���ՖX�T|N�����(h2H��u���=�k��#�k�l�H3��sI����>���임?��f?x,�1��e�n/ �ܷ�?�a����!�r�@��rVF�GU�|�t~��le��m@�q�)yZ��/��1ie� 	e������BD�3��#���C� WfD�2h5 ����E<C�%�+�dPljw��y�~>��ot4����r��:d(���JګI���~�4Mu��\ ���ĳ_h�5G}�Z����b)�\`L�����x)~�4��C�[���"�x��`N�.:㕚A_Π���"�C����
ř�|6�)�������u�Mܻ���#(��Pu��Q�H̠�Z�߃�]��
�4���+(n�4�^N{庮��_��9N�#���ugv*>�7k&6��|3�¢��I�BV�;5��ʌ���<�xC>2��v�jo��P8r����]�?����a�!E'�M�6��[��E &~)���y�A�EH�a���tj�!>,
�@/a�x��jrʀ j~=�k��nk�D��eR�jYZaĆ�]��u�*�ˮ��cKߔ0}�m��$�I��o�)$P?9��v	X�dG�Yv>|�	�!/U<pɠ\��䪣�Y�nϤK)�ɽ���ƺƀd�cW-�b�������t��k[4��4�7$ZG.����8!���Z �dc�Xׯ����H����Cݜs�� �/g*�yZ�T��ՇJ�FĚ}��"k��8�[]�M�DO�Ҡ���I�ֹ9߿�d����"랺�	 O�ɞy$�(��[^�V-�x��˘
v���XWU�\qov؃��i\{�J�z5�O��ST{�\�'�#G�J\�ףj�oA��<	-w�1?��{$�Xܧ���C���	���f~��} ]�E.{�-�355�0�{���8�
�� �~��C���#6���<ǹ���JeW��ϏU��&b&��|�b�n{�P�(<h�zv��D\A+�r�	D�س$�jװ� x������ 6� +޹��o<yP��<�$�Lu5t�g7�����%V���J;LX�&�#FkZ`S+�-�ߥ �o�غ��[���Z�`\?�VJ�K�pR�<y\O�+��?5��cUw��b}�W�d\��N��:>,fɗ�M��Y?|@�[�	�o���Xq:��Ԍ��0#��m����fk��Y-�5�9d9ӎ�h�.��n[g���A�!����4򼩯~ �bE,3v�d��_}Z�RjQ�O�nN��j>R_4�D�#��-w�2�x�%5@���K�'�=����իBX:'Drn��;�����[Z����7`̦�e��4��^�	ΫqnZ������$�|�d�C�K�P{\�2���3��Ʌ�C�C�&�=�*I��~��6�~�'��5�����lFO�����+�[�rw�`bi�Θ����`�XU&�/
;'e��2�|Im��,	D'
�1�2q*�6e+�� ���/8@�rd�ֳ���B��Ě�A�+�5g�w-���q.a�{x��k��U�_,������۹W7��E�<*(�6��'C�E5mv�3Շ}�!�5V��J��k}�3�[�� >�m��i_2��T�MG���x��B��m_{��M�P��.cuӪ�fS&qs]_|����]9��z������u�CS��2��u����`�����<?�,�(=��7�Q!����cHk/�i�p.xm�{(�t�3���P��yHŖG����& � �4ڥ˼x�N�M����N��4���(�(f�(��L% 1p��_\�y-����J�8�Z���bi��C}{~Q��MK�ܿ6�$2�1*�C�f�7M�BQ~%�L�ʍQS�@��?���]���9!���P�g��*k�<�ym�P;1��k)Q�lÅ�� ]�b�!{���O�����,9��\��K�j��ZB�c57|te��~j�7m�LwȾ���|�۶��]/��<��cS#2�[2������x�;�[D�|G���<B>�g��h��/R��j'і�inT&�(���A�{ �� 	�a-t{��$�*��0�>U��s�F������ s��N����Ga6��/�氢^���'�K_@̸`H��̸UC,�㉈4��}g�K]�����u�JJs��VZFo&]%�|��mK����P�x\7J�6�Y�[�I����ӥ|��W�K�ex)����|�E�8��__����\��
��e���C��̠b)�d�VVR�Qj#�!�����+�*IIL��pN�B�~�cއ��l�"-���a��c��Bv�	#�9�j�fZn�:�j��U�����h�n7[<���G�6�u��Lp���a;���n)޲�6(����Bc;��XU������G������c^t4]���n3	�E/}o���1׿���֋�rG@EL&����&�R�����ḙD�n�:����%������åB�������[Ȏ���(z	>FB�=D���\�&����C���x�{@	7e�Gi=�[�G�E.�'*�S�r�tk��� �E������e`���T�H�H��2�J�/����S\#ҷOF���(c+�p����/f1#������m��U�R�u����0��W��=�^G�䜿f�7���8�;��'�{�n��+�UwJ�i��>s�ϰ��)��N֮+����C;v�T+��;�%�$D��5V=�~��~6��SZ1�4�! n*̌�vf_�	��__X���:M�sc�nP�v�쀚<�Sj�٢���R������7�G���9�^�������K���|�wcΠf:�gh6lE�N��]N�9��vsK�rB�{�	�є�r��ݿ�!L��͋��we�h�1G�Y�y�c�)�CHQ��z�Iﻦ���A��^<��%���ː�Yu�L�@��:��v�.b�b���J�s߁�@��_�ū�+����j��e!�{��-��(g�ʫ��U���|)2����&�]���5:$���vGt�n)��|'d�i!U�}JdM-�mH�Ɲ\Q �	�Y���ˣ37�܂[�K��'��*L�XiO B3M��r�f��Sz9���k�ĳ�~_k�>�8�7�ԏx�*�\���Hs�[,��[�
(rQc�s�ى�\Nf����Y��M�
��#���%���\	�ˤ��������C*^?éҨh�_$d�u7s�A�N]W.e�h>�ׂ~�c�cj^u:�?J]R�)Z�NՋ���l-���mg�2��
q�w����a�	�-#���ҁ��Ɨ�q1 �ىq�1L����qr��A�a=r���X���ґ͍h�Օ�I�-�=_���ʤ�,��c�N�{�@��1�y2��VEl4 ������Pӂ�Ǧ�2Cf9$�U>�a�D�;�W�7�O�?8P�FAR���D���1���H�����I����&H���w�V쎺N�`��ؙd����'!:<�H�$%�B�'���^vB#`ʔ���3��TD���w�s�6m��0�%��Ř%�uM�Lj>��'��a���>zi��U�"��j�v�?�6%����4>�O�����;:�n9Te��0{agjh�9\S�_,�up>�;�4o�ɏʁy�$������VЪE�䴡Q���"##L��0�?����L��ZR��ֳ}a��ܾ0ۡ����R��� Y1}��}�E$\m8���T��i�ۑ���0��-X�,���x��1���n���P���u���2p���^�;�w���'�72xc ���M�0ǩ�����?��xm[��)巂�����%r�����p�YS�,Nz��,ӻKtF˾�ζ,���S"���gN.e���D]�hZ��1�N�B�6�+z�8���bӁ�ª,;��[�'��dj~��V�:����#����C����\�M��ڗ��ؑ굒䉠] ��L��0�n.�:���ki��pil^J�D��NY�ϡ�l���W�����.���{��P�Ҧ���r_NP�����w(�pg~�9� D]]YS����(�e���d�
���.��M��m��1�dZB#����Q��b-Ǎ�_=OrZ��e(���q���ch�\`�x��KJ�R��9l��M��h>	�`���'�0��"x���P>�w2`�@��?N��H�^��	[���^�ց2�O�*B�����o[μ�}đ��z��%�Z�'Ie{�ސ>� �}��Ь�h}��b�X�0�k��84/<�!nK3H�<��)#_�Yj�v;�4��e�8�"%R/����W��ZB�7�Ǽ�y� h��ꙜXn}�&�Ù.�����fKIP�Ar��l�_��{	�r�<�տ�����˦V��&u�E���l3Bc����g�rChN�l �X�mo؍)���Kg��ֵ5꼄ԥr�/�B0~���*㱶��[��g����g�\S�%�P7�c�}�����(�+<Ǩ�-��z�@��!��h��.E���0*͋?���]�6�ᬷQ2��D!�*���rdX�MJ��,J�+�ڳ�i���ƶX����,N�����ȝ�H���T˫]5�hU�hl=�ؗ��4zU�Åi*4>��']b�W��(�F��G�yX�<S���ږ�>\$�������1�Ǿ�Ŭ�j�5$�ҕ����V�$1�#~�*��V�K�//�?�FA���	�)r�lP����5pT��������f�7���G�KL���ز��Y�Tߞ���z&=f�CZH[|���O���?�`-�f��ǣ�E �3�2Jޮ��DV4�DL�'0��Ǫ������� ��c͓��n�u��Hd������Uvؗ!�@��?Pc	n�]f-˕��s<^_���̳��"��������5�S�>������?Bt��|J�*G����!RZ��i{*��"?� ������D\:_(خ;��h��a���{��Z��.�����~�#A�읻��N�qm���%�)�q�b�B���(V�v�~��̚�ن��1�"c~��ƻ��1E���F�")�L\>���k�(���*�`qs�Ia�W>�5]�"�N�c��piq* �/��P�:n�5˛��7��<k�j�l�u3�QͭD�P:�^�d�9�d��]��!�3���G�?��A��u�d�
H%}݅�7�q�M[��/Kx^�ƍϋ3�
^mL��Q��{�v�Q�_�q�d�[Z+��s���D��~f��:�:[]��eą�T��y���p2�K2����ٶ~�B�_!�7:E�"0��A�<⥖WQK(�R#!J��#G������(�fTM'�L�f���t��QϿ�7����4��"��1`���a�,M�Z9�J��J��űN�N���{�O�6<��Г
���m[�N��l
�ŻgS�ƻ���C�u��ިV	�R˓K��r{ ���'��� �G�W��f5sC�C�����_|�@4h�t�/XG�LZ� ;���Ŋ��!ӧY?f;�:�Ļ��Ѻ�0��O�+���Kl���-� �hEh��܄}J焹�߸'OQl/�E;�jI��?��@?3�m��'�gP.X�R�+����9c?I������gx*����&P���+�t���>�2�^'��(�y��;��mhu�X��/^A�������*8�g�4J��<(5� ��gW�Ɔ 9�Ȯ:
?fO�ʗH�o��a�˹-�)���A�����d��}Q&����R�a')3�k�XO���	�W�ș0)K��Ӂ�p���5AĊ���߽@�y֝����n\��>$��~�FA�'�'Ղ��C��N�`�_�h�>����H�C�ly�%��T��3���Я��2�k4� Ĕ3pY�n�5>��@Us��eOP,�5�एx!p�K�io���~�2HK��͋�g>\�@�+/��rIZ/����J�3��7�ڃ��z�{f�Eq�AW@)x�n��U�K�j���W��w��4����[Rp�^>�'޸Śx��xe�7<�r��s���S[8M��09�~��w�i�[�P��1]��c��n�=A_V	�F=	�|ax�P����Pb�rШ�Z �����6H._┝��~R�#�W�� ����7�h	�XABo�V�F0��-�J�p�)��Cw�=)�6O`p����s.׾=�� s��m�Ĵ���eE�ٰ�p�ЛP���KfcV���D���He[�s(X͸sH��pJ�R=�*�@��+���\w���p�פ��4û�T������J�'�~����K�̓��M��F����m��Ĩ�5	��1��c��C��j5Ķ�Y�m��̳Q�wȲΨ�IxҼ�+�f��8/��/-���pbЈ5Z+�=���ow�0��S�:F"����W6?�ܸeh+�"�+G��C�A�f�h�_������k�7�$��7�ΡX 
&%2]��Y$�Z/;��	ۭ�,%-��'A&�*
���IPD~�t��՗z���}�CS�i!JY�'�9���X����6�֙����莰3�*4�H���
*C�U`�$MM�S��j��%K�pkޏ1O��ڑ���@35r{e����t�N��Z�A��IGM�����z���?��F������;�LG��4y+�򆎇���OWG��/�1�������!�Ѐa7���6�(���L�hO��[��� 8�����q��bp9V��TA[x�R� ��9��}�)D��+�%�� ���ʮ�#͇���h�kd*�=A#g��VTo�m��\�� <��}�!;[�w���BD7-�lzR?�	�)n�|�p��||�bw��>�Cs�R�@�J��Փ��	R�;�1;Y�y�s^�3���EX=4掄Ғ�0�2y�-9���޸��׋K*NP����*���,�gC"�mxF���J�ȍ�)��q�5��m�zfbպIg0��3Z�3+��&�����fE4rXz��x�
��@u6����9���M�(��y������"�2B�=H�|�	��wO�D]�B(�U�
'EO��x����g=��%�%
j�C��UHs`vӱ�0_��0�0�F��sr�0��
�D"}��(W$Yrm�vϽ�X,R�[�?���O&�I�v^s@+6/�_`Cxfh��"�ƚ�vJ]�lI9�[��2�Mͬ��\�M~D8p���AYɶ��;��\B mm8����d�\yj�YRBzӖܕ����2���kG��V�{m������#��9����; �T������%�C0���<VV��e��S"96ywi�;͘�xҵ|�L�Q��yhDI�~�OP���B[[l��Uo�ܯ>�c�	H��*t)�Kq��0�������g6�a8Tw�<�����e/�H�_�zt/�,d��]�� �5vvMY[�[R�*�\@�����#��ha �Vp$ G܋����iG�YE]�ī,u���6ܻ}�^A��l��V�zu&���[Ag�Ǵ�9�#�}v�S����v��,&�G��~\�����5�m�.��y��N�T���;!�d�w����������^婶��Fc�3��n%:��E�=A4��/J�i|��ץ��Y5~��b��/�@�܄U���Yř֞%��d�ZW�"��x�̛y^:�Re鴵�C�����U�T��$��7]��G��f�R�,����ၶt/���|���C�
����3��I&q��A]�;+}q�4"#���b�&�}�N�U�i�A&���)>�9]�e�9Fa^g�"r��7b)�*p��4�{P^J*T�{D�\���62ѐm�:jm�3�7Q�|T����\���a�R>Q�w��jhtYI�۫*�& ^��ШZ��Zv]��z����P�p�GN1��L2��Z�jr��v�R�������+iB�ܸ���0�vwt�"�Iңx��H Jt�D�/�c����/'B9MR��<�!�N�(|�p͊��k�Ex��z�+��37�.��m��>p���e2���-��>����������E�W�A��u��i[��$���n-c{),��}�P���ep�o��20s��ӭ�)�AD���D۳�GZ�>}�v-7��L7�N!7D����I����b�T1;)ȕ�o�j�u���⯕�Iζ��jw�Wy7�QN��JCl��Aѥ�}y4�C �N�ѫ�"bn�Y�@Q���� pJב:��&)�27v��c�]|Q� �_z����3Ի�����i��y~?,e SO�Y}����!��[~�"����T�bn�-�<��d�8�w�C?k`�sͯ�����!���	aժxp<�'�� �7g5I�R�|Ɵ�#$m�m�ޓl+�)��exCv`����'��w_g p��&>���nJ�&�g��̶5m�������*�*�M��\�pF�tS�kC�퇏����g�ԚG+0�M׬]�2�N5�
�.��;b	ʤ�ZGb5�Y��M����i��D��W6N�������0q��uu!�]I{��

��NF����-�"D�x@)s7´;�3�'� ��l�2��ښ �_(�q�p5�^:����:해���p;���.ݏf��`�YP�y<�#���o���<h)�G�/��4���t�Q���5�|�f�؎(�n�v�t�?����p|K�Пm�-6����AΓ����߸�&��'_�.&�W$�_f���rj��f 4���b\��Bo��L�ZߥU�R*=<L��+W�g��`Z2�>$.�I�gr�N7�<��ey��>d��������9Ҹ\hKe7�E���u�����j�q��*f�2y�O��:-���H�ə��N�pe�/�m>)r0���&�6���͙�G�m�g%hDvT�@��#j��]w���K�]��n��ݣ>���4�m�$v��I:$-s>Q�Q9[�8��^��m���"��:�su��xJ�W�g��ke� J�x�2��2us�棴�J�M��fI�2�00*%�b�3�0kT]�-�˽8z��/���#s7c�un���a�����?k���:�p ���Ć�d�a�̻w�ƌ���rg��cHiӯ�%�X8�^�����e�ެ4�]���Em��8Ğ�#��C����#��<#�~��(����S'm�{���ٵ]K�B��͎U��;GT]%~I�1�x� \��]�Fv��G�`M�*���>�[@���')q�	�� ��u��������ipHSz�(��
�W4���C=�V��ݭ��x�e�v���x�u����x��|[� :�~}��vm�2?�����]�#�q���v^��;ĩ��)���]��V�N�j�+��GA~�)�C/\%3���rI�����Ƚ$�]�^�`K�C&+�~�����~��y�%�,�ĵ�5��"/�9È���W��q��<G*���X��c6+I���F�=[���p�Dc[Qaϡե��]c6@6je�C�z�]�U�#��Zw�4&R�y��Ɖ�.[B�/6��Qei]B�E�OA�h�����^���o�tB���皮�f����w#"Mk6H����-�K,a3��t��|0%�>���)@o/�E�����s�B�?�D�L��`�ɽ���W�\*�9�p��Ήfu�x�i1��)7�P�|Ġz*H�xuy�6�������oо�$Ka����{�Z�f�_��k���pk�g?]����
�gl}{� 	Z���h���X�vM�]�< H�MX��G�6xu7�]<]������ևNY�.�cd5^[��O$��	� ��R���9��K�<�О�P��*� ;����7��` ^��ZaR�뀐���8�3*��L7 PΥ�Q�s��g�8D��s'z�n�˿g�꟟�7����b��>�+WC������BU�G�{�kcS��{<�a9o9��tZ��g�دG&d7ì�*õ+�V��l/.�K������X#Ŭe�<�J�f+U�x��S�H�C���0֫ ��9���Nź�9s��[�bEh�_�����N¸��l���Cy Zҷ|us�G�y��B��A{�qB�3��r�!<�J>�}���K�5�K#uz�y,E�0�qf�b���g�8�>�8g�p��s�	�ˣJ� ��ֿ�H�����-�-5���"���a&�a���{��������<;j�����-�K%��Yj��f�H��O�~۫i&V&	q�a�!Ԙ6z��ua�yf\�N���:����h��`6�0w������&���aP(� )�/��D�ei�)v�vQF�~���9��Z�u�Ö�������Hv턆%G����c���`Vi���5a�p����>�eXH׀p��2Bi-E3�̌o�]/'�#_�OmP�Y���Ǆ:t ��?4��4�;tEh����?ʽ-0�W�_�9����%"#/��M��η�{��Q��k5�����Ҭ8N��l�ooϣ��ʝo��`�@����A�
��Q���z���j�4J!`����@;���B�mtW1̀��F�ɞ۠*]���'�!f�x]<Z��~U	N���TG�Y��gt��I������$Չ���R&�������h����"h͏B^ �ȥRX�4�V[������V���Q����,6������T<�26�ƀi�IJJ&��v3��F�x���9�5ݺ�z���4�N��*��V(��2֣Zc!vJH��9fR4 �%�oV]V _�D��޹��X�
�i�v�DLۣ����""�cm�r�a��=�$��_�^�V�+���@��L����2� @h�hO &i��Tb!:���O��X�w�^��x�~W���\V�!"�ۋ"�3xd8�3K�тJ1vxN����!?d����H�8׏���X;[J��� ���-G<�-����ԯK�b�ݯ{X�|��s�61Gu(�-nXָ�Ycҕk3{��t&l.��/�.ZYz��\�n��?���ltX_�_�P�<�n�$#�+�}	��f�]�5�+�L��h<��[�=(~a�Ck0����D��O�@���L[��Bv���τ�=haa�����Jf,t���	W���=��h'���Rǿ,Re�TS5���Mƌ�7�R>$�NJ�m�J��m=�`>c��D3W����'v���ffW��[}���z 
�B6]�뎸�F#��q_�2�tRdɿ�+_]C܃�ɝ��R�0�&���<���:�N��	�)a)���t����ݜ�.�}F�4$�k?&�R�o�^��w.*E��8(`�S	b�����ӻ;�1����GB��2��u�f��wX� ;仛ܽ=��[��r0��L͍�θ����Nf&G��dԸ�g�1$���u����� ��H�i�fm���Qڊ��a��͹�a�|�'&�_9�P�kTK	W��a���[g�� Yp�	
��4�:��Z��(�5���r�����O�=��ۅK�<@A�:c�1����P�>@�������bC	)ɸ�z��4�됋Z���9��V��	���!�~J��NZ��z
��]d焉k��o �����:��4١� (�L�ܸ�߷��IzWc|�ͩ�Vs6������&�����`0��585�rr��9���ϑ��� �
�� �wE,Fzk��o53*C��-g�O	I���?���{���a�i>�)\�D��p���o�n��W^��U9`u�����9�N�0�bXP��E$�׊��j���gS�m4$a.����U
��&��vd�&hܭDݔ��h��*���	ՏH���4fন}?�Zb4��j�hJ�g>�,{���ӽ��(QD���/� ��y��:F|������0���j�Z/��2�|��l��rF���5��
�𼹯wb�y� ����4������r�o0Ha�Q1kc�o�2B�S�e0�]�VU�zDQ���J{��]�X�!�)	��-{m#+���q�j���}k�N]F��PG��A����Q�*Y9#����{�D���+�+�ޟ���Wn࿤7'\^_������XZ�] h���,�IH���D��yIdG����g�f��_+(H�[%�x�W'?�kT��˻Z�:�/�-�c	'
)���ֶG�G�p2=��.<d���B�#��*������y�Xa���|c/"S��o�ߩ�o������0��~�/�礱���� ���2ǋYWɈHQ>��Ȣ1�� %[\��P�h�|>m�[_.�A���F����G7v�A�6Q V���/-�T�,ɚ��7s�έi�R�`쀜��ga�����MPl.�rh�E���y�X�ǘ5�����c��x�p9/sR"��K�`���"�Qq?�������}�j̞� ��(�A5�p裁���d%���ƫ\p�^�e�B7��Wa�:��̿������L~���7{�)��
����n� ��uC^x�jy#n�^J��=�G�di�g�Z{��]v�>���v�E1�����`僸&V�D����l}6!uc(��|0�@O*n�7i$,��R<��/bF��� �<=��%X����#����H%���l�� �0�]����Unȑ/����t�ZN�x
��E�{���HQt(h-j���ؙf�k��T�x��S�੉��%��X5Y�2���B^�،���Q��͜�pϦIs����V��;q��.(
��ζ�+�Zxat�8Ϙe�CF�M���*l��9[�+ �	�_���Tgp��Z@l[����.{w'#뾽Ŷ����}�����~I����.��nm�φ%E�.�Y����TT��>��Ut<?�7�X~*4���O;�Җ��\i�P��E,N�;�O�"1n
�N�~�朮DB~oC�G*�>�h��+MӉ~�m�ā76��ngF-��Y�/��e� �3����/=\��A�b�}S�l�4@�����l;�Ͽf��z��Z�p�<��&���4���(s�B�7�-7��	�J���_Z�
]=�,~�\���H�CZG�=��ȃ�b_J8��	b ZHw�|�5|��<�����҉J�o~l=�T�%Ke�0�W�w�����>R�̴<#�<;i�R�X�
E�6w�g Oe~�!�㔀��2���]��=#�wH��m��P�Q��d��S�d{C���~q����Pj���Y> ǤN�Կ�L���w�G�{��*�0��.* �ϵ�
�8�a��.�Te0�Y����/f�4����B4�=ߟ�{��*��t�	�>��_�`�S��y���!.�L;;�:���ҢMI���A�w;4C�[�I��;mqX�l�|l�෎{Vd�x^fw��e�j��ũ�lux֎qz�y�(�r��2�gO� lc���ߐQzW�X���A��"n8�N� 2�,�|�4�-��������N�P\k衧�]�i�7n�S@` :�����m�}v���:���?6 �W�')�BFVA}rW����T0���bv�9� ����ƿ1*�6�1Tڵmj���"��ԍ(�X�	:X׊��%].Y'��<�\�8�d�!~�?�����;*�B�L���ÿMp�>�|� qN��������\���7�;����!���h�ͧ��(���3���l��Y,�Y��/L<S��~5���7��6����
H:/L�H!]�?;��D"S�����̃�2HP��D���N�@k�q�O���^Ӫ�\$ӳ�E�<C���&_���f��"�CS�w��(@��̾�l�:����@��@JR٩2vS�s��=�w_�IT�˚W�E[����H_���]�&,�x�3@������ĵ�{�9��x��ud�-��R�E
::���U9 uԺ{꘵Op�����S-�S��s}����1"�Cl��a#��+X�Ν���4�-{�R�r��k/e'w�UI��O/��7j�����O�଻��k�ךx�U��������MW�sr�R�M��B����r#"c��4��9�78��|�s;����R���J���z����`!5ަ_�6X�n��r��X d��)�F6Z��OiK�3ix~M܎Ǥ��@c㵙V$��1O*�
uߴ�FH<�H�q�$�����{۪P�D���0��1�7F�l��+.�-,��K�?���[CIC���I�Z��=��v��F��6��I�e��g/Jiɂ?��_��?��QȖ�>#��'�G��]Mx�� 憘���Q�dF�����<�C苄��_%=a�N����F�����4gmI�0Y��Y#���ml�H53,*��\��N���ɼS�Pr��������2��r��sa>���H�x�Zσ/'��3r���Z�}�C�=L+��.�=߁>Cp�qY� �Cְ]P���t�����=�_�p���مH��S�h11c�I
�{u�+�г.�9�{�z��*#z�-(��9ƺ=?���sb#&Z�
M�;6iQ7�&(����#�	�fDxW��������W�{C
�7�[b�X1�ɞ��}��om�~��v���kqhh"��'��Y��o3��9K;�d3�v�F}��u쨸6��ܕ�'�N?\�c��)�L�{�06�4��T�<��-1~���n	�6��!������^�k�x�o�	��p�(�ɢT�i ��Z�_�x^%b�Л�.X��D�1<�ĲQv���4$��2�ΰx��|`�%E�3�7���<D�5q˼�Gm"<�5�^H�@8��uw`,�̠�HpO�q���_%��o	�[�>B�`p����>�
}�74���`�%��'���U l>�+�\�)K=_��(�$�����h`� �ٺqV��o�x[%2]�(�{�ζ� ���^��6O�~��C|y�;�y�²WP�htѧ�d������JMC&�SO��FF�s����|��,�.�]��XhE�,�W}��sl���<�;�Ūg���dMh!I�:t���MW? ��VImԬ�'����G-b���/c�z�'[t���~�<�����)��ڃi�3=��G�T�GŇ�$�͎�s\Wy$�ԕ4>b{� #{�"��9`�W˫s�����|38aS�C��-�w�t�5��g��6A D