��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$Rx�y�<��wA�*;�x���@�̦�W�X�fa�M-$u����n~�%���P�$��W��kYَ���P7�?UMfT��q�6�U��k�>����~�\N�(�����X�e���/6U|)�X2pF�]$h���d.���9E��WG��L�X"]�Ad����ľS���8od����e�GT?y	7�������ݵ�^��R�q^]�鍦�����s�ae���h��L��P_���ާ��YЭF���'\��68�b�[����w8�[X��V�F�0͘3����q諵�uW� �h�u\V�?@��_6G�_�*�G���B�絉�f������[�G��U&�����~�F��AׯK1�`c��[<��FY���4I� �#�G��x[X�=�Q1��`��R>(�w����R�O�?����7�,(�H\�#h(W�EH=�������yq��Ѿ��aF����:�U~m<|��.��0=�P/���4ǆ���T(���۪�!q24��G?|\PoIMT�ֶ�1����NEG��z�,F���=�wN�Ԓn�Aچ��#�J�}�(H����*7�(��Ղ��ޔ���P[�.f;��dI�Y��^�#�;r�������<9��m���	B�Iד��@5q�W�M��n��إ�S,���5l��#��K!�)01?�ڎ���������N��R\Č�B,C��Xf��A���z����
"�L3���i �9��j���3�e�Ȁ,WR=޼a⡆��Rorg�?t�)3�(x�-(ؿ��C��g������%\�����d��t�!>,R������| KZ�H���ߺ��rqk��z_�q��~����gioq�}�~&V��tS��t���9?�8N�xw�vߊ�a�����#L~�/���>����ڈ�^�R �%�W�����cU@Gk3�׹jbs����"D��γ���Eu��;N��*��N96��is�;���ǒ�沟�o�J���z3}�x�!��!o�Ev��{S���l��8U(�va���P7�����(x�)DP��S`|�ฏ�7�Y��q�~ i�d�D��[�
�>�\�K��/����f�7�!"��Ȧ|����+��%�'|�g�I���ewc���|�V�,�����;��T��J0x����w��:�����|V���w��p�@����Z���ɝ�K���_[V�z������@0�̋�.f�!�&��Q��#K}ǲ�NFl�I'���MR=%�){�C��K�V�V\G�+�7���Wt�f̽��U�O/!��6.�9��/)�w�%!b
rA��-����m$$@� ��8�!E蔩zC���;
g�A�"�9�7<�pH 1�k-�#�A�@�#K�`|���T�(B:="DVq�V,��?����|S6+��.��p%����	V3���7���/9c��.0xuy��|QrKށ`04�'(0���p��4#����4��ٞ�ɯ{��'����SB����|x!.8��vG�#`��o��9�V��-�Z�ǖ������"솮�f/�>�p��mglz-���<	��&t6���X�|�Q���8�H��)���H4ڝ�#�'���U���X`�a1sߔ����l	�@����e4SvBk"��"&]ބX��式�Ӝ=�n���`e[���V�S���6q�xZw���e�	{�R�øS\����B�I�g{ �e�	q.��jx�~9Xr��4���-Z?I�����JZ�<����v���/�I��:��[]�{7�߀����"����Ey��Ny�X�:)q38r�8@�āҎ&b�]j��^�q��(t�_#��ř�˒I�f��$CojcP8dO��N-.���!��̍�yh�+ͶpVj������1�9�$��+��W#Mvc��S������9�(a��Y-���Gl�_�t1��U�L�Z@��
�� ��E�-Q�v.��o��_Qܪa�̐p~%��o�3^*�Jt�vI����B�ǹ�X|�Y��f*jI����<M�~�e�Z���mą#
�K�h0
�����0<LuzC��
 �����q���A�@�>����l<����n�QDz�s�;���g �U��~��&�i�u�w�)�&2���2aĶB�R �3,!v�x�_Ђ�O[=���;�q�x����jJ���h�$��Q�so�j��iI��9���jU��ɤ*���ITl��ou�sEJR��6_����܏y�LZ��3��'h(���`����8�ESe*<+�ܻ�Of��ζ�#�5��V^�Z;�����T�;qȕ=t���c(��:�Ԅ��WonK~�iд*9�nD.׮�7nM�9�=��c�h�j�4r��],�0+�3�y`���]�Z�/ed�\߃w%�<��;��&ǉT�������&�Q�u�~����icK�:8���0$��Ϸ@�� _���D�r=��%�<S\���xC6?|P�3?ਐ)��:��*�:}�Ǻ(,��@@63��.g��U���0��ZKi�o�����zNKV"�dn�h�}�L��ʯ�bI���>O8M�N}�0�LWZ�'w]�#Z�/SĲ�J�����T�[�~��Cg�cvf�R�u�a��p�kN�ƣ��	E� ے���&����YPi��M��jo�P)X��>�}ET��T�K�6	����H�P�q������4�Gvd�6Q�b<�'4��_YV���<?[s����;*���Ǹ�Z������\�$�U����;*�BFIK	��,H.�T
S�	bF�N{'Y<MS"���M�ET�|��u:���^V��?��	� ��y����e6R��ay�=tb&Ҹ?U�v�C��^�u&`[���7�mI���&�C����~dyvRPX���nMU�X��f]����Ugژ�$	�y��$0�L.-��>��8��(<����R܎Zo���*RWp:oRA��_4j�!�(���r/	��1(T�+�cJx,؂��(�:GE�Z�߰�8�hQ��%ڄ�:d5}���6c��|ԣ
�3ᅘ�7�W<���Xoǅ��&_%`���a*�y���b�2���ԭx;���۱{W���?�"�g���V��/sNL���	V[����c�ݲ
�kݲ�MB�E��f��P(�[�n��6�j�c�l�R8�`Qx J�D�<G��/{G����7t�p�*�`�]�k9��k�M��2놟%2��ދ�5.9k��������A�K#�!��E4�A�����7�ҡ{Z�.я|^)ہ�)(�˅}~�����V�S���IN��
��룰u/5�6��K!H��ɌKV���_.bI�Lk������𕉋���ݰ�Ǜ@J���乎BG�ڕ��^�#/ �.Q�(�����e]�:^Zy4ק�,_��L1�?����.(y�����m㷾��C����<�؁�dw��M�� G��s����� dg��i�j0��* ���m�}L[�\�1�Co���Zm1�,O�f8�#P�)<���_Lɡ�j�d�My�y՚� �o�b�����̞��z����aX�;ٕ��N��)	Xz0�G���a-��$���ܹ�b�Q��Q"�a)�H��	�*�0H�C$QMޝ-�`^�� �����Q{���,��~�Ջ	��`_oJ�0}gPnЀU/�(�]��z�7��I��؍�����#��2	ï�̍$��k��ݽ�����L��b���AB	r���4,|Gg-�ԒN��=	3�9C%?�HJgB�,�����0��a��K޵~������4������_�4��tkF�, �!Ц�A�Q^L�����Dcq(�
,�c��98fVá�{2����8�~X�`/�_9�����U�s.������I��#S��'���܍U�M�X�
7"���ii�N��wCt�?��CQ��58g���	hI��Y��$�GY~�>�A�c��,��P��*&ٻK:&����B���6\࡬ciӺ2��L��뀟��&}]��dro���5^NY��Bژ�c;v+���g�PO�iS�s�̳a�t�YH���:��v�������
�G�U�a�x��1������� W��I�1�w�����.XM����Ȩ�|[���Ӹ=�:} ��<芛x���N�(�oM��&��N��$��@)JM�}�1P�9���H�"���b`=�XE�2�?�k���=M�}SLd6��0��w�>k �z���}��6F%"����/���)�ƇG,d�0����������,�ĐJ�P
���0�?��5���)g �+��ֹ���P���� ��d�vZ1�'BN�n�m������_=P�ϖ�E���T�� ����n=��%HT���������)��**�}��^��c@�����+�<��`0�}���!��J#w\� :��wT�IE�$����tM!H�m�\�O�䊺5�/U'�J��	Vs.�~��?��06ԣ��)��tJE��a���mc���k�vF�O�hQ��`c؃�=�u;�&w8PNJ	2�b�'ў��ɉ�1uYG����7Y5����@W�(#q�[ T+M�}�x����EEi)��QB��e��P�H�aN~߅rL���W,�?By�pZv=)��QΚ9�H;�NR��q��*i���F3�%����B��{���[�r��
�<�6��Рb�yԢX�gh�ǡ�Q=g�'?�M0����%��\z�9�)��su�����4���{fL_N�45��D����1ԑ,����&x恐�r��bo�����/7Ϳ8�&���)i��V� ��^	^z�D'
0L:(�k�y�R/Zt�0��� ��I� ^�g��=�����zv�8��pK�m�`�q�:d�a�0�@v���9xX�m`�tUW��7~��p�ލ{�(��1���\_Im� �e8Pa�����w���y#���U=&��m�����q��8�׸E��4Kz�� �?o��7M{����ZWR��h�ݹj*=�+�z�E�����k)�ݵ���;N�}��+)7DlJWD���C��|�c&f�Ii��T�`�\�~�h7�����<=jd�,]�H�����W}�[K�̉�#���S���}NJ~�*E&���u�I'�M�2�.x�I3of�e�od�������Q�g�-���kW	�䯗��[�G>��$�y��3�Cߢ�pΡ[�^��f�ޝ|�Ӹ?iH!dw׸����'Q�[Zd����xk%���$�����ü>LQ���
�!��8q��q
T����J���-/3�V!h,�4��t09{���/� w��<^v4DH7�G#$��U���� F�w�=%1!����w��5Nk)�c����Q4�Fe6h5�_��y�5��s��[���!�O W *;��Y�����J����$f��7��ވ�8�v=�	�F�99'.2��#�!