-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Ia62bQ+8POq/d//z/VLYofhUrNMgGThixTAC6Z/DhfrtDWIzzwIt1mj9HTqeRYCPQDU3Kk53YtZd
VHs0mxRxUOrt3KZN/NEad1f81w+in6bt4+qii+edUvEhgzssQJhFENzlHBJkjLTQG/4EGCvASFhK
M2vogLZBMTlr7w3cPKuIJ31yG7vLqqq90pkI/O2yecqM5+mBwXCv+n/wH+CqSjDPGy4ia4yNYmSb
2QX3P0dxpr+gkF6dM9ZVs6YMWAn1htzeBkdxVX4azfDOvdDOiUUPEfmM2K70QIaGjVPRK7IAif+U
b6OdWBW6/Pmt3NhErFncS7qQVVSHw1IauiSr9A==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 20544)
`protect data_block
CaF8sI3eQ75DTqPz2Q2NiwXUx2jqkSafbI5ah8jRe4w92Zviab3Lc4VccN6rHeOYd362lZcFbXEg
NJicAyy9/DRtiioYJVi3dCui70WmHJ0K2PrgIuDKKuPLSfnZohVPGg6vhmiPqvdFh0kF9kQvv+fE
HFYCSKnQXLQmOfbIebn9XBTaZZ6cj8thzDBnhYAPW/To4bUpsG1Mj2AfrvaG1cpQhW2piYB++txk
aabxpRfQFD3ync6TTpvuEP3M6kpSmKQdnFq+pZQJdG7WiPOX5GQVdeiHMYsecGFp3S49gO/APc+d
bRvVWnQwBjNXv3VFcUekPJWjJuX6TmD8uFnxQmKjHhdYsyl8SG5bYYlJCBOP1xMwzeap1AkADSfh
rKXt+5UwvQTytZI+vmdZa7jbuWWXgTFIYTwyeplFFFEHa5t/aKZgZzaq3PQi/cq5wGDGjxg0JLqk
o9T6TG3xtgHPDjzM7+7VgiJqVky2+9qL7MbUmKO9sfNH3KHyRxCBNxsRYMxDgAHxsqQh9hzvOHpE
NZieTEGBrvpluoG5GjWDBvDHoDuL9z0FdiP0E/H6uB917bmVGP27E5hn/7gw0ZhgxiCZNLYma/n1
Sv84DOqsflvY1XwHBRZnkAOzHyn5RyrDh+idfiBppY2+MxlOKVK+q/kidxOpEkLBZHkOAwKC2uV1
rlhBjs7FRSxw4S5TMuH13QpRDseS3UYxInfvFgVL10Y0cULR7qVYae/bhQzTB1wWNHLY/ioS+RHF
ZhEXSlcmFD9yPjj1fQw7X8V5AqirxI2lGEam7VADyeiylizsqHbtOdzxxRnTqxfyWDXV3+GVuwVK
Qgzp1DZBC4NEU9C8Fnh+gGPFFPhpnpxb6JZ74X2fLh4h+bt7YjN73++oEUH1rPE7J01mUeoDd5pv
077HOB4qucSnANw0u9xfyWcf1puAAGdw5TGPsVHTAmzdfvetijjiSp3M+mb6KyBjWUtBjgMYmJgb
k3MYjqu//+f98dW903W2GG7oIw6IHLs2XndRoNCcfO2eXw5/y3asUWlgxMIj9+r0ezj+eUUfqcnn
THAyE01+hjaVnbOJRGgU67LAGo3OKkEMZooPPBM0JpFWwYLpnCWvLAY9mmU6DaNcrFHhbgHtzP4u
VlIJ9LWBNqEMhLVP9BIqtxGqLvww00yVu5gA2Knvb0aWZBCoT/ZzNXctPuW48r4CmfwzbQtbP4oU
ihEV7p03UybvgOvdI0jr3SaDHs2pvU2qISNj4gX/9aVGTvp2y29cmgCJ3QirIC+lzpDIpotBs64W
CfqJPky9fyrfQJT2IosRioU8XCf3NipVt7BmkkX/FtL2vU19gt1kGXgRlmvoK6smX9hv3hpNt8oA
WP3cpm/WpUWah15VSIic8XtKSd7J7QAI1hiKAGZc3MALNzlXb+ZjdxQVjSvW4KX0pyOJCA9EBvRe
BzJoDvUV/4xJblIYy+HC7a0IvulgD1gYdJDfEM2D8sNhcBsM7YRRx7MnBcUvKeIOOgvkHK9g5KbF
YgSlecPOxH7E0gtW1nnolzLxh6sRV8hufWH0dLd+Bne5BpvFHzDevTT+azjmnyg/u6b+SVxDzQEe
+I8AG5MqnVHUJp9dpCbIY+o0GGIPqJmxZuu435qUm7AANrekhUrLiT3vCl1tcxwUykxoA7NLBnym
MxxVqpUwDo5DBTw7ev9yDaGaas1vEO6AUooOXfyOq5aVQm5xJ6sLNqZPZM5K9e84n/DwSXckYGhL
y/WIvErulrfyibrmDTnEW5fh2MAyuh6YW6h0zXxjYboJcJlty6xFz0D7z0eY8BWrLKw/h24NH6RG
dCCtHmaGUDx1ihePmrA8+lX/bJYHnCNzATFHIXPtMkAe4lDIJrONzw4pQ8Zx24HW2GvtpeYL/CgC
6TB64b53iR4pPlV0W9j6j6K3v9mIpIC8WarYTNJt9VpmKWJIg43qeAPhBTK7hFKY5qWiCzJdTAKE
kkmsRCDrMT3TQG+XJ7mbQ1b5AqnV1h+2V1uw3s0fywb5AorE1bnjV/erVhKmlJilI0O4ywbuJM6z
oV5aYLGshV42YoeUfqes/uxErHyBE3jz0bau/pKw2tZcJq8eqhtUaeK6K0iTrMeDHdET/aL5mel2
sCzJZhCH60wyUyDJT3Audwwv3UybHqpqMDihc+oflSWXXGqc+LV9wQ7fnmhtHtOBos/sysWjnRpi
gvdAjzm7GK29u/KYjyjt6suvqoQn0+YiTn5R9NTSxzJoux33b007z9FFuAyq25ImrewTKmaOrxLv
xfby/PGtqPWLxm3ToQjUB8+nZmdd2QccM7ABjBcEYgnFmySf53IY1SglMyK/26Q3HtyF+qxz+XTV
QYaONGtheiIx/i0m7h9PS6mhgCRMeYOPvDk3wUcpqGhW7RbCe4DO+dvgGsfiiPZeftDMopPILWTa
US+gkIMsTE+93ZPlngJtFvmA10MraJ6tkUb9U6JJx/6OtozrNkqs6H0dpKdrThjd8sQ3xNCDYGPZ
xPBjZx1gYOs/nTnD+xKO5vEb0oM3v8KD3ywiDH4XA6D3SwfIxWKsvGCXZuXZ56XaNbLQjS0aIxC4
vhRVCYJq1w1xjHl/jOTx0Y8i1FjJ1uO8Zs3ro16WqujaIKyFDSnKnH0p4kwsDz0AVgbiYLK4q+nC
h8PS7hL/BPsKT+wWiSUQgQ81tZfVq5Sdt1gN2HzXXBo0IMV4SZZwTnQTOwHGIej+87b3oT9SiM0g
0NBTC0gOmAgEqWBUP/BpOmZCwQTMY7LYCnEc/QgGi/jP4kpywp2UYu6OdSitbpf9IDsM24vqASqh
r8bNQ5qmHoRZ7PSSkv7Bgk0bC4PaQtUmK0LY0iCSHkIfy4/IoRKcxo+iR9fBOGSxH7BUH6q6abXA
XrvNnO06CnsqcxBAgdWfb/4F+iBgrvDIjRK90uaxNk7rNsh8Ka4xN2/+a0ynLZX6oj6TesG83BGc
qdpM7ygc27x+6upifLMxueZT5/o71A/2MPLDMDcZGONrq1Fo8q66SuutEgHAYaXFEKj1y5X54sCB
39tWznmQzsmF5OzibBI9Ojm/uPgkNDfFb+t+hu9UAWBG1vPPE+VhPGZQJxwxTm4gChjXQWhkwWSN
XTIAKY43hUoZyJRHMJacImjBQhOk6vY6mvF46DTmTDtknvTeuX1DOWlLc/lnH8N15tXMxvUpMpza
CLz7qXDHda/tLgei5s/9OmD1pzGHHZb9jUIJf3MQjohWtJzxHy53M+6yi+QTL81Q6NinKq8ARrwf
2uU5i8FgsS7++rE9uYMI7flFr8vXu468xrw/wy4Q2csbUS1Ao4xC+330epyTb3LFqN7JbKVt4i0z
JhzFVj4YCkr7eNOtzXcYQxSHCGyTFF4u19gaChrFPmu7Ss4WuuAF5mu5GrXKr0oNtkAV/p+ASiMD
IqDhWyt5uQjBRBGt8afPV6Y1fO2+bpAs7566nNS4Kje8ogm5Sajdn/vgc7lfHZkQVKXSbkwsa1tR
BiPv3q1MDxVZakRyEWHaT+QwPP9GzChjIQOkZJmowTKc2x2+sBM3FL4R7XH0HRN7bZlQk1Y0QsHJ
/BDPqGsCcFYS0EgoyhxVhMMMp2Na+jeGAVJ6Gm79FjGBWWaGf6EBP/tZZ9cN1gtOVIA5qv+hcepQ
sH5mbk7+g3th8j3Xi7KdUY9R60c/m34LaW2cvZU37QeycmviQfRPlauxE/8IGe6EcmjnJL97AOnS
UqgWNuGKj2LWbMg1G4P6jWy8YSiZ7PIDbz8RTnneGOMCjzKkMuCnDS672oAia/6HIVTH1/vHCm9h
ZedzcefVO82SOoneDMVN/jO3Y2EnBOXD1ifXDf252u/enhPvcXYpP1yXBRpZhCstDL8/v54C0xcv
OW6kyYgx0nI6XNyma7Ay9EPjY9//KzQ1JB46PwfzCK2EvUqxebPJqx9HD/cD+vo0AfRSslXy5EWp
U9L9dd8i2v+X4/WG2A1RGOawauWWh0T+4yTPSSlIzM8cb5h7HkpcYgUxb7ZFWwyFmAr45UYtupAU
56L3aUM1HGtOb6aqCKHbpJXa5b41oRvEQAuhZm6O9bRD8kD6QJPAzXxGxKgX4VODKaVD/fTthD1N
urSrCD7fzXeRMa0UMoMuU3ZdCkQwkcV04jEUNXayem9W2YM9qkmjsIRLOOHAJ+jgLYaVygmUj48i
ovt7JS7xdH7LSiKan86qB6P5H5MxjDcIHD5rW138uKGaz4MEHNJtlrySr+uZFpDAylUUW5JjZSBS
N4i+wqMvxN1WAHe9zopNeu5A/oXbycnOOXgIrWKe66Ha72DCjTgYMPiQn99ZO/i9/tP4oEkW5TBm
4OoYOnjPekhlN65nTmtjXvgJPV/h8rYbHTEB88K3C55OdW2H05pBJTCKcQ4N4tND7DXVkazUOvCz
X55s1OgxR1ztbVGx5aNyLrrI9kJfofzKK031Yen1mwL0Aa0bG/woiCpqk17MNd9/1Tbm5SP8xh1Q
WDXxfLnbS0jKsHy28GMLUlB2Nv9ENGaaVsbEnBiH5w1LEFYJYMzCgRZgWD1eoAKfYkegaQw4LCAt
0E5uwaSJOFB/1jYGq0wlWnFONaueKABADbeZ9lUHJjRRLFsSn7/51O5Ec1Wq2XbbqMrdB0dz/19/
B+9pC7F+DstH7jlIMevqfrCZtxsXJgEE8ZzH7002H3PfbtWZQSxqLwszEc1vYzox/L0WsizdNP79
HxnzNB9P0QjiEHd6kpUveNnQ3FyII59yeWd+E50as2SGRXPO0Vp1rCh7arb4/4+HY//4b87K9BlC
AYK3Hsaqzg+UG3Md30q/2pv8zgV4E/IOnfE7zw/LuNlVovNIFI+NZXwDdk26oiG4Nm+AUcpZhyxA
r83b0uGVJTEipu0VFW6YHU6DK/E9qM5mQzJdm9cmQowd+19v/G+l28f6KPPpRxHqXo0dKducEE+6
2WZCisA63zzEOF4NpaJnSZt0X0hbiOXezEStBzKKrOk9lB5aNgqfxJwkB5oTLE1I4+ZgVl6uBPer
c78p1zjEiheGHLHH+RLGf1T/Oaog3D2da1OUJ/XhJ+8/6rmmsiY4KLTzfuJLgkH8EHLjPS4zpG/w
D+bXy0Fj1o2CM2B0Tu9jcsdhxAZbi+nR1cCFQO1MdkQawO7qUxOdIQWw9NhQ0aKsQhPP0BYQgavE
nlc523IK8tUJaA96KPRfZAc4PSf11ZFdaD1LrsZp92ZhNGz5ub+aI1RSHW9Rl/0z5KlsGPeB3jDg
w/hYmOel1XLMyc87RJ5CZj7a2ViWDAP0ui48ldOhC3Iz3y4tEtE+5+WVtQE5AH122YcCDdERFaTI
ZCB4jcgm3vDUeZOmp+1BSp/5YlAthrA64b4dpxFVLDtHQw2aetYSWDdTZs654OCt04B2eOsx2Z0r
B/T2W36u6AXv8kDNDEa+/6lJqe87ljdF8DiDoElYeKgatvtkbOnzJxQSQvXY5KR7pz+khFdCDHJ7
lEHUgQDrbkVcZBRl5HwcK8WX/G7PC+ryT+j7/xCmljlwmSKwV9MO5nkI1m+KKE3Zet09Pp1/a9i2
UpdLF2E1NLqCe1ax/Y92l4KQGtuFRS/JkjF26ypwpw5wHtRVgRZBxiDDC+vWObnUC1x+BgB2EE6W
sLo/5U9UJd5ctBxdPtAGKGUHZYdzOAOxrk4FcAAA3a3Gy9ncuCTloyTuubWHbYHOHinsohIcskZs
Le3kS+vWCCsWPJbK8Keim5A3nH6ZYPXUXFVVena1uMVjhbkGhxgOjxEW9F5EL8pbzWUjCMdFW/nN
u1Rhh5BH6Fpc5gGZ43Paq2xBRpFTlN2EnTthbr8ne2NXqWWl3ohPZCEziQvAlM+KwaIuh0YSEyGa
blSZH5DX4fRrD37iUSpsKrzcgc1jDryLiuW34PmV2+qqoWdmRq9sE7suwMotgEUIteqwk9es0tMY
GiSNzpkjhaBg8TuX0p7q29XaVzJftCXnblQvH/H2rXhS4LK5QICkao8MF5uqvKiBLLPdBmNCj7Dd
ILJMQ4TPjTrHN89LIxVkUA/8LR4Le/cnKsqCv7C4qNd8kl+OTgHgjzCrZU3aGiDhr5vjPuveo2+v
8bKkMRBniOD9RQ17zdwrH7KEQUecwfVyOrOGeXhfjf2Wjz4mHzyEqIB5tiRi2DrtVTkf0QT5RT6u
dK816LjbE1lBny0ExZ0v2bi/7f8T1G70TxS417HpssSMK4tZ2SvCCUj4VkhMV79Cl8E67nl2PNki
RMyWCDnw8/erXSIEvwu9L2DoDvaIa17rMCFyL37fV7HyA03S9hF8tKpOY4v5akbjdLjv/DCP2MLW
DcUMb64DzdKPBLSx0lwZYJl7Rx54YiH6Oi+4nQ652so80oQ3cdl2iX8g8Uyq8Dwh+64NBXuruHzs
9N4QzAOKWDmqeUrMFHoCDvQWUdfY07U0nxO9Yfp2sW7cRGjKNQoQW0BWMPtFCon3groLa3XI6OZV
q8KAvgl8fvUo/yVADtAKwqYd7Y1wHBgIM0cfqemcooJS3U33Ekoa+1ShF7nfc7CBMKYvAz2Tt2ot
WiPylnrFMHNgV/wNzr9ZOhBtG08vNmXqlmbLlZWl5Shedjck7RQoZCx0i999waYuNMeHPQIJPfdh
0tHYuxHMA5e563EVIdzCocaQGflD9nJ0zFb3WvRdV3fDWkyHx5ymSvis2QpSfaIy5GQLfd4nZOhV
Vb6l9487tuF7d0H8mBEX4GjO/qzfJm3/ah1js2qx2rqr+keWuhJXWdNaVJcoPVz0eX/eFdZLso0B
zb5kW5W77V5epjgsinDnCLRd2+Mm5B0Kxzb+FL34qGKCmVAD2Hs5fpKURm+US6BKKudepl9JPWzo
1Tnt37KWuPyesekNUFB+YcgjWAaewz3Z0+lmhzcSbg64MPqIJSvdf6arRz9ZX3YqDWPLdhb0LGWd
6XKgPLRZIv6ZtOkq4UgUDWsUA41Zn4AKsJl4eMU2XUXlIOAnlCHZfgzrTloH0I/qskTypem6H0vm
4dV+gyQJ+VE8a6sIZ4L9OW8D3alx3738pDiBXTmR0+Qqq/q8aSKiHtqAF2upPGdqIg75AQyWQ0nI
blO9ppJJWBhK3gPbEPPNtdp5/y2ha/raO3Tjyk/PdPJ407AUt0BM0E34hqz+NdtotV0cnAixJTE9
LQXZDzeDkAMLzKu1VxVtt09yEt7HfECKgYa2ivcOv4ZzRwjtE1EI2yEI1570fPOkIPKfUssAprjQ
fnOMVVA5Z0pJT4JsNASXbtaJjWDIUXN+PPYNptEfVi178x9S/EEuDMi3i88U3VkZJkW483h1TNOV
dYWn+jZ9FboNZxv1GC5Xe7gvfHL4zmh23j6PNF2lDrfLNJwIutZqbHVbywqtfUxWABQ8F3HtuQzT
vYzv2Qg5003ZB7AxnWmZKu5n1eBxgsiv/0jSSFtEzRiOi2pL9mCF0mBb9CMRIIibR3RUHZdPj0aN
8xgyFHxZ70jTr6Er2f97m5qpMYeLHNq56/Kjb2f2kH7RLhUzllUz2INkP4mhLC4vkbucY7xtCLGm
RZ+3oeOB0DUKBzVANr4TgK7dqFt+SBjUI0fYhTEE6egXoPP0MzcictU2lb7KAIcllCpBTAKSZ1fq
O/BuzR1Nk7RE71/oHYajGKFNUeCq0GmNZ5kOvpZzs3N61KJyWHwnkWEWlPUCZnzFpuUnknf6Pdv6
XCkbYXsHUaZSHuWO8kj1TFiMwpo5DnGLZRfFBVDXAjNnSQ9PeWjpVm2KkCNe2zwDOS0jnUsyO2pg
I4M+H6K4iNqV9u6ApeYd62gsCbFJfhe2YtiLrDnNNj8KGb5LX2YH+GmwjlCKpTCEfkFnbjBS3ATC
2zJoVUTaqhk6ObY4xcDu5KHqoveFkJVeaBfBQ+mdfjZ9lGHyRHPLsQuwHEcHMO1qwx5kUInSdJ0v
F3p51pKlPMt3dwq/gFb0PDlhr4oM4vSSmzMr1RkkBo+ElwpEsS+rpB8QVC0hA6cHHsX6MiLULhX0
rBhbQLHpGTv+XPY+iC14XZK49d48o371TZxVWZv1dT14c/Ukbnwoa75eptF/JQYlhvExa7dUxuhA
5x+Aa5xh8UPig62NFgxSCxf84SDQkQ061oyXQ6HtqQ59r7eiRAxxR09YL6atqJZKyo/iVT/NDgyr
BVNwbqcp8uSIzabPEZto71UGyUzBJ0mNZRZtttDnyEAPmhbtzWgvVwEDG5xZMxFw46hfD4W67CWA
8WLWZ782T8YlX8yQcbP4mqHmD1dLMlPRxn0pCGBYKU9WidxaAGV5cjsQMTTUuAoAxPxfFjASLIid
n1HAUb1ERNqWDqFnr/AKAdgKv1J1YeDnOh8Gv0Y5xtgBQbQa6v+ogUxj2Lq+LP+dr99ecdhuQxT/
JkVI2W5Jc8pgU5wNg+Lb2OR17+GfmvtVhK03RH7GEmkEqxAXtHL6qFLrXiAjnmJaYT2r3i2sCgbu
5mndgfsBhwuEBhsToOwkfj1Ip5bdp0zVvwhy24DlVUqc3uiRZSJ7Xb0w69OB7XVJueEwbxi5bFYY
WsGqGFj7EDJYGD2bvZC0Lg9FM815IzOTxvewvWlAiUcyJD5bpwJWMS6iCK+fBLQQXN2CkL4K4RVF
1yuFN8s3fD64hBVsVj3DSTp56qHRHOutcjMYEPSf8kfnFai3dfktoBnVsCy1Baokd8PgpGwGNj7y
VMxttLUem1mUrWJRuP/hRd4rlw/DUO7LRrb8MG3Fnj+kNyN+jmUGNBk+H9U10yskfgHg463t/dxT
Ml71WLDum7K0Pq5LJIT/gBGjPhjviZXt/C3x1YB/J70BK5Jqv8HDcPSTXY3QjENSy9vFDbHFhvbb
1eyyzEA0kLadFUFMXWZ/5VfVXd6cSNtR/jDAPcoxZ+NEN1x+QMAHLvC3rlbBOpxc/FrkXET+tiFc
9pKTJi1Hx82qUY3vKnNPl46qscwngj8UeRD7LiDQ4b2f2QtDJ152qF8fFHjuJLjgMBoRlAjRMGUg
ZQnmKttNgVj160QqGqtopI0UzHrkQSfV1B3h879DxrYt5l8pSP7rlZwiPLknhgHzndfzNiia0iud
rd1iU/hfFx9axVna3nYjsiGow2+oJeIZ237LVQjR1+UL/La14bP8uGVwbYtQFQpiKu2QEW0Xw8O/
rdCzdCD11r8sKrqEZr4forb/6UmuMhX3UqYFL7Ge7MY+wJ26DsvVb47M05fCIszKGZ3cBtfymbeY
r5fj/hrPQfEtJ2S6YTPkjOiN7qV5sv1NuiHaaFF/Tm3TCuI8WjtVsRiK+46p9T5gn0cuOsdecK+4
jU3E6xsZyNxhf1mfOCBlhMJ0I2laojjz8V7NALNF9W8YrpeyPcn+EM9GamrwaCWANK+mGLxRtJgz
Tv1iKnSsD8cTLEKTU053qiqDEjAktAd/pUj5H8rWlXiOsT70jQKcA6D9uEwrxofmm0Z5+nC7Dyi4
+xiESmE1cYcBHUF4imd8yKq11TG39IK3Dwr/ULXjPkFY4I14zP2x62FIo7G/Se+8hDcPIX/K4Pkq
nhqa79vwCuD4WGUSrjqCQMwnkvgmwjUckaoFisxdkYGQbUDCUT9isYghZv9E8MP3eGv21g3X6toc
akIggJMRaoSxdpElFODjW8Wi7ogWJmM6Ut908jFjPsaHmxBcNtMMLrIaT8tb/x8LU2s3bR5w2Ndj
649Y19ggitTw/msxQHX6jjHQbpPjNV3UDCNh39yTUxCGVt0lK0fviyJxSdCCzNuMdFnxotVLV+3u
QE8m3HlAzJWztcA2aTJAYkCxSyfu0qMCi2HYARHDPuj8+94r2ymXtQ+cX/3FM1vVb7wT2EcIn7CX
T8KcRa7wMA1Xe8v8b13PRiBTsZr52FgxIFJnEyImfiWqjE110D7x8nzoXoXnA5QYD6EsuI0BDDJ5
oTfZI7JOIekivk301qV5Ec9XMBUCj1q6XczTKEvzXpGWBsGkgO01MSaLTMha1Abr8kaIkqVD0x6y
Wj60+ujxsYXUoXOtxvakzUMiN334Y74FBxqdNtndkg3Ahlm2N6I1mZbYKOGSt/kmeeHx9ls2oXUz
lXQr3ecrdgWalyy6muYgNZhTXPEAQORp3nlVltkbUN2VomKFXy+YbD7Czmr9pGfCKDp6nRxaOU4A
jdpNGhF5P/mkF+qBTha3g0FUiushIeKvhSzrZX9OzDm16hAvUK4WpYUFVwfpd0CgCSf6YYBNEX6E
oqPVW3F9UQAeSWVQOrr1PLDAHNOZy7CRxglbG38NNvdMlmkEyTqXGABCRytiFAwdoxNS3Fn6itVi
YwkJ9WeBOzjn0JWAstdCDMGOqnIUwwWxcsy3E1p9dof9Qjd+ux5TrLu/2Zn7ql+yRq3hxcmc4V6i
Pi9mu62DJH95yBDjQCCobVfFrcldPzpOZFu5z/60ZWPCSNiRT2pkGvsZwKTi3CJ4kyuiAqHwjxX1
+SUBunHBFx/nJaPhJCVSJk3MbsPiQjyhibL1Gv7Ezr36yljoCIwRQRGGnFfm/JC7E9l8ui2epHMI
RWRApbHzzxEQf4u0BB5+iIhdayC/V8wwBVMp+88YzjkB/bWe1B0JK/0a6hCSSXBOs2MnfAR69ln7
cgCAGv4uVTwebFjX7WGwCoUzQXTQzw32Dh3RyrQFtOkx+jp+vJ55FCXD2w8+LGubUbTeaahWPAaH
BHG2eWtfxiXH0T7FxX0nAALYWBlrTEpGylEcE9pngLPqt+wPKcpBinENjP3SxfyyznjQEaZz81P4
z/GSXLrOcj1LeQzAviaRzt86CBw3MsQPHYqbZm+gwcs1hzTLBHQqIIvCgbudOW5vkI+Nq8IqNnOx
mGhGLriypth3a2HqajzHeJaz3xbTLdl597D4Pkw4UzNQdJGT9eCQeBWREcm/zV/NaZlVd4fooLuA
qJ8GD+5kb5VEYIPRu3YekCwc6FAJM/KjhJqUyH8QlBUJ1mj6HFL0QZ8mbUY3R5egVDMAj/wJ4P2u
LkMcMuccTikW9QcLaZhG+zlnep9Kly9JDaTrdyY9WXPunIvELRYdKsA/d2LHqERr6YJeunR7A/GX
fUUuf9aZKoojOBPG6m8tG9ttYqH5MLKYd6hD4uheCA7vCVFW/P8tI9XKIWz4JAcEzWhqmdmtl0wQ
wVga05bf+DO5zeP83Cw+cxSD0UR8W4lSpr3znZdtJ4e9ylUZnOYkNElEBQDk+TqviK6g6RP5GMEu
ehQGmR8ApCgxreL4YZVt/YBBvRwtYkxOYFRF661/MlWX+KqIWyMK7QTTaoYbqC5jI+UlxficY32T
QnjUacATKR+KHcUw+rJsuumQfYvHpky29zoxqapL189t9MVVBVQ+dxaCv3+uEnjXxs4Z2sNeYvZo
Ugr6yrebeCSY8xdWls6/9BoDpYYUoKJzKsLcBfjGvrwFRE4JtTUgTVmT/vAJsMCse1w6wepQe9fz
WLa9dd6r/E9LLi9oeLZ3ezyZemxlyJDHV7bt86ZfqLVOEdF7hhbqvmINtGFW7V0ON/33upXuti2g
D6tJ+V1cq8uj+Aay5ThDPf0xWUlrqh91gBufPZfmRxBc3WLiMv+A70RPbzQNFyYmndJ6fhDO+vW5
tgBiZr+rb2Y/YoOegLlMjYJl5pHZO0NqQsccYpADUVpzGwU02OoVd4isMnBWeZsLx45Dm23P+wBj
AMfkMTMszmaffwcAFzIcuXwVyHa3FVJHEBsEOxdenpMdDVF1BxFCYmAETL2Mlx7+S8lsu01GPc29
c/GA8rZyveufu8obIqSbYhnwZeW7cOd6GE346+79pjVaLkojHR0cxVHfT5JpVibnC+MbFXNwRHg3
FkIlZ8wIqbBW6LS3198RNN6B+000IHaP+nJuaM6Bn/OhX26E3x7tUOQF1gY1gCk3RHkB4tPwiVe/
ADkQYJGjYJjiGhp5SlfT5+KyxwboN4ft3mPiOakykUz59Xt12Y2TGNAnuiHk2nHkSpYzkK0AQoNY
Jap2gkM7Hc6tPDGENwpGlFSnfywP0b+TX3jAVd15OU1HTpNrxU6SJqhe/+esuO78n5NNsjwbNnfF
pzSO3xKoiuQGe0H+7ToUo5Ic2ntqk0vt8ngNxLxkEkUh1YwKLAL0LjIpVPNPetlxVztvf6v8ECpZ
rsCsdKX8tZtGDwD87jH25OBcXyX31ot7nXDyTr3+HzOLSzqBRc78A0n2QKB3VlUGpamip7NQwXO9
A7GvzuzKEFtzfIQKt2kwilEkDXHyXE8Mr5E0dllyFMKOle5Ly7amsw47P37bLzWtB+u9ykQF3FnD
SbL7rO/QTBNlQAOjX4Zzp9I3oNv1vmFJLbiI91MlI0n55WJcwdVrms3taq0XY2ATD85QbcciyUQi
fKerNtirNtbcWhqBB2/mmo36+4COwVl2lxjB5ejXp2X3bjgfmi4byKtCLt6dXkOCVRQvmBJVC2yX
ShFmENdRmWIhTPxtyV01IjdWArdqC9kxr+ftzMfA9IA8DVyq/OJrazOFMk36gEPKW4FeAelDUJ0y
/1VZrOxARNOEbqo0LNjeXwcwubbtd6Rj6028VhDPoc1x1AKpvIW4avKvCh+DtwHGSjChprIZ7RuT
fRzC8nysGwqcYwdvOByCj+3W4CLlraxD3KVETr/obWHCRn1zMJ+pPrAS1mjEfDDVZ0zsr6M4xQMw
N0+uOd0gcjl06/TBK8EmWXkPEFKJAif33gquX8+PjI7752wYgSaEkcbIMrcmGuIj+Qovq7aTLK7b
6j1rAhtmz89RfW2AMuVd6jZ4tZiXzeBs9qpyMQ+lldA7keWIerRytX3slYEBsPF+cGYVYnzTNY4G
2M5mO8eqck6YNIPH26h3JfkqmPlejxvR8hhJRQrkfLso7UC5nOHqaPYMHuDEzY5lAxa1h4rQT3r5
QRypDzKgmtHtk5rMa9lnaE+eNmQCDLHOANj/WfcbxqyJ1nOXYcYW7xsu7CrkPOD6mfCPQ22sGb6d
xX0Akp1ek+aEltq+GVO6MaZde/2t4sjYwJx3WChqpx9O7lw7/x+TXVSksfQfnBT0oacOYcf6JgRN
wvivgGtTTUX7g9NVzOVDX9zRqJwxVHBnLJ6yuWVOu4zloXuVMUQTLpdKDEvhQ6d2hW+PIyZj9j+/
64Kdobp91GcHgcELeTwUr5fnfKg4qODwzf42ZIOQOkUlCVYlQXrlzfzgn6RlISYNMvrIYjCftDNc
Sm/rq+axph8AdkF29sFcb9nISWO/yV5ceR6QhFUO6CtCaKh/J7UVbs1KzYe4cYPvbJmkXwaz4gRl
SSyd21ALT/PTeb2hs10hc0pl8qV8Lo1bmVs2QA4zvjZlDaSPHrlGRoHsmKvWd3HrVtb6VmB59sr9
i62rvmUrknj4IQ5Wf8l5y9kt9KVI1qFe+CS2aSR82IWHvR9+6Ria0J5QHPxILHuAKuTz/a+17abZ
JlkrlAlwPMkNYjEFNpJxiBVNBxYDD2+TbnZkEET7fQQ4nowDGDT0MLA66gR12lQvgfLEtjtrWXSl
8aBFu8UbemcPUvpN+IWpPsf9lYvKi2LRTtO+HW8WGaHzbWWdVPU/4nr26wdienzalwsiExu1b2vr
Qg9Avz1+urLnsVtQLpP0CaxRocDuKR/qgKvAd6ZepEP7KN77H9LzJ38vr4p+PWDHsm8l/BvU/XQM
ezeyHZ16M/QAKG2StMYZLoAwwQeyaiA9bYVubLlhoPN2cOUBPXkpQ5LHcRt26HYyWKjWFEOK636f
gAOlal+Y5pkczW/0M5E74vr2zgiRJ4aGFzF+9opRvlkpW6HA/b2Wr4jzL+ewV3BYmxjsk7YgrSzP
Znvn5tcaflNphncbTadHfN8Dl6kmaU9LkLbKF6LEM9dKU2JMnHOlzdC7KBQl/6Nn2LmVGINyfBn3
mKe3DnzwWtoCEt7L/EkeHH+hKDAHZ5j/rHW899p9b5pFAVvsUL9yOiGbIGlOGw56UIrGZ/QuHi9j
ApJfjKd5WQ9YjPKGQ+dD5BcSiPrOfYgBtq+J0M4TmFzoN/F/gQNfzzWqXMrjqwS8UC2oHMBfnl+Z
/OIb1IcQ0e5LJN//O6ety3sbCxixsGQpRx6YytTuDUH2nkNOPEFRuyVASoNHuKLbCpmh22UsIDwP
CvmSSBT/tuHD/1Jv8n52/92xE/453c6nDk0kbC+HGISwRgCfYZko5NFfoxGyJ2rx4SF1vPeXIao5
LfpmKXEJvQLP9QenA9lbn+0fqQKqBbKkd4Xoj4Okf+6KGyFywUi3XGpYFazIZ53XjyAsEEdlR7/c
npWkO14skhp3tZqDo+4lLUPJ0ITZeCXR4SzQvBU7P4F4nO1ervXkzJANyk8hUvspfvqRTeDdUIJT
V3w0IVEjbkTEHXL/D3MLi2BHKbSbEAcTcKPNKUjYM0hpQ2iWoWqd0/WxSG6JGlWMuGr2rw7HdTHA
FbzHmCEIGbrOTHg5Bi7ot0hUtUAocZuv0wWA5Q4mOY2FLK9MN6HuyWQ+Fj8wdDjZ4kzNNQ/zp2ZG
JtGk0nm83UtuExGztOn/YjNrKHmHjuWfd8TfjBe+ob0jqZuA9NTJMHwUY3BvFtfDq7L1gScwg5QR
v8T7EwBc0n+TroWpvDQd8nlaf1df80ME3vwpTURedDiPfhXalVF/nhYI5sMuN+p5w2g5vTsHmxpc
PeX3S9eRPVlofPLGphGMlEAeZcFkNaW/uAW0Wo0CuKwND7YCZ+PwZbXk5Dk/RNb/CxgYpbRruOE1
EgWgIiKkGtQwyAHavbNb5332N38sxfi01G7a+ywgfzehNTZEOQc/myKx+MCkcX2gpdTv5pIlk28D
479XAYOjBTkn8KDjVnUzimd8DJuA/EI9VasVWBW9mYoEi9pBha/tpQK1lSHX0QyROShDmZOmfd4J
qsUcdksHmidL6s5orATP7cMpJNhfQfWwXkUOa43epRbp5SHRBCDPI4Mza7DNR6bQSqi4PyoBTOH7
RyyOlpqPSzM9gktuxVsrkJCI/xAvUsgVIZ0HChikmA5YkZOhEjlPthMcbAK5AaFKlsS3VF4Eqe7t
cLqrkS2l6Vq0UT2dfxB2BDpHw/BH4Jh0szWiIKIc76NlSvNO3h5e1Jl7IBkwSIV5cZ/4s9tjb/rp
hvGtPPUQincpAkL0QkahMof6TqByHqceNKO1qOh6lSto6+c4ijlC0nBtp45j04oMr6u2gnEgM0Uk
c7xCN/YN6JpJdLmedMGleN0LTpZqim8miU3hh8exT2tsvF59ao6OwJAiQ45mKrgsSgYO6iIdTA9S
7ZRyeOVKAdKbZte6ygC+5aJUcT5cBB7Xbf1HBjsXEVXYk8jSsbxkb0Tcmovn+3gP5JJ6+LXIHFrp
ZKr77N65Yx4J23UfZ9znll+7UIZihwfK/5vTPBvIlNn/iVga6bD3bubpu7mrCYZduCoOetmNOzf0
LvnzMh4dQevsrQPqSQoG8OLDh27S0Fm0ZzO44upIYiIK6/aMcsbSvjh+gJuMITvBCR9ZZU9vzC/W
ez3Vxx3WgOBbJ6blYpN0J71C6A4UKpih6gotUXDjN9cw2YoUqOMIGkQlKtT0YbG6CVAJTcfVUy8G
F40cnZ7sRLWJUuMUwLT0UlyIaS79xrO9i7Dw3X/L9ROt0YQIZJAy+s44XyNaSHwqHOzBR+mw2eH6
V3np284eUuops45RN0e79OdHCqEqTRovlFNiml1GtUuLDameDB18xB5VptE/IjvvnLLoEzGoa4YD
VrckA6ylbMdaa90axoGj8cypalMqP2gZG3Q7Nz0ttGdUIdfrUCJ/mQKRAZ+N7Ted6pMLoP7EvZui
inftMR6EkMTlxB/eS3wolOqpoeq8AX3KaHi8VVrnGn5gnt1eoPo/59FoOY3RdyGY2bTY6a2CH4Ll
/0cRbgSbXhcjEJjdJnREJNuhVuHdWmFF7zc/WxEpcsPbhAxjjlizC8ybBSBlp87OHAdUQ15luEFj
0tGNc7uYtygQPik3aGgDrwswizwUMlIIbXfvps4qBsrvDvMK4GEuFonP0YRlc0dM6RfixnHFq0Fb
wcX5Uxu1y4fQQVuUWalRdX0BKNYosvuhEWKvqqW67Da7pEDhuzYq6bJUFbKHFP5KakuO6PPSTsu3
hBUAx7djRoxCSnbKRd0iM9YtI3wNNY5Wt0HXiew6a4Z4kA0ZmOTYq83C9thHGfpmT+CNzX4mLiZT
D6X4y1Kl7gfB6BcJ9NqoCiSyN/m5GOzQZrjWGLgUa+PL1Qwz5pNckS0yUKrvni3/n3NOTGZbzk7w
NfVbJ5FRTfJsBtVWddvXRm08HMqvObFU+y9zj9V2i3dWzz/kU9WEaNMmOXd6NcN3drh7QBbopzPt
NCYDOjNAEz1hcjANXYNJ7ZiEs3Ph419jg0W7FTxO4bwmpLs9kVLf5ufPTzi/hITSfbkcG68Ymur+
A6Y18+MzBSRmfmRyQSHbKJ3X8Ig6h/64xo95ho2g5cTmnoo387HcWWG75zw7PKzx3W82lagcMy7v
ejKELF6RpnBuSqMoydhvVGlZBWSU3sWyav0XU3Yx2jIG3XcrPjQDoosFrs8gq+uek2mx1UaR0SdQ
zFmkhQd5yNIOJLHRQCIGU25TtZ7K32DSVfH7G69/5gk03+8d2JxRJVHBVlD1CBESRuM9mByw30N5
NFpXUNBkpXFqQjAMVg7MQCpBBMTAYmmfDTbogOa+dJH/Pkii/wZQvjII1GEHxNpijXL9RZP3+BDq
weh6qbKfUdqjUjo/fOa2E5t2CE0y0EXIrwtknYeYa8AyABbsRRRltkfOUqwgwSboayznyWFDNXaF
brn9dQf40nERIDosS1+KCoBa2Ke5cQWkPG76obvANuX7Hx0+uXry2v4XbAjvh3SpbL76TZ1XvN5/
jmziFd59CxwZv/0W9v5eSR9L99eFSx3lOzeCYxVkyFE19HmJogndB5WmCEwFKUi9HjCFJeE5vT2Z
C3ajO6zOFPbG1tJgG2v8rUekyukZg8E4DXf07b6h9cEj2hofrVK/fwGHw9TvLg21i7YAi8io4yxC
GI/RndFBN+MHrvpEMFtmLxGXKFzZKCDvxHu79V0UJ7YMPCbcHFWcjwYfhiFxHhxIRO2v0vv20pen
x3qHE7zf0a1Nsjh0U9U0C68iLjodxwqsldk3uJwM4YmB3De8xqKcwMhg/+EccKqg71FEZHbonS7m
GSPfDh455eLsJ9IChuE62lPFSJpDcbV/ZV9PCwSgIqy/ahspralVAZlDDwAwsi4vIZEzdWKaeKoF
1xnYHGkrkdVaYJ7J9Fr8vx0jeEzHlEdF1K0yj9ms/IV7Fju8eX8S9Yi+fe5tcEHKLdUDnJ7p4gZj
VIGPAZf9oll+WWH608OBYI0EzztNFGBLIrgVx2jrVX7Od3W4coLuAAXLTwJhMVEIoPtVMFA7frCh
dkWPprbL6wtcT5PfBQZoJJtwVtMRFjEFKPO3GdR3alReus23c9KGadRgSq12pXKDqWVDYbpYUrzV
WuW54oLz3Jqh42MN23n7rqnMl1ckDcCJD3Km2Pwwf8Hc1FEcxF0wNj8igEJu656bmqlRn/Mww636
a6B9NRVcCtl/EfVm01Mx0yLSH1g7EQ4xps9JbuanjXOzXWd6xyeWFn59+7n0o5mImVlTf0879hiR
U5TZuo5nz/+TXtND+cy98oQ319SgAcnhGNRPHP58uSHcfDWHgNGbfyz7EltrwyXB/AWQISSbTHQ8
lAmC+FN6crOyTekVaUCaOYtp39f9BSBWohqIAruWITM1+UQzCqkb0vGfuZ0AZ9PP1nz55BP+Gwzs
z9ku3DkHqPWwE6gdWv5p5jLVRAlMX33VfHaN3avSubOoDcaOWtqjRaG8c1PIWWrBfIYHPRZOpLKL
fug+4kCOxY6A/R9m0yWOtDBE2l7pEXZALQnfpPytp2JGjxRdYSUp2KhjRJwPu6Scc1ngFy90/8XF
yTF/fFCk6BfsWtK5DDRQugrMQdv6L1xz37O6C8yzCSkt6VHjsOd6cDBFMl6DBjwgpehkGh2sQD17
1gjWZGqsL/YBNDKcerVJ8oR8dVhoL4RCQKK1y/jh61T3cSKirAJsIGnQMZ69eWtGBAIYIpZDdFu+
V+n+m2rZr/WvHlTUnxN7pCeeQ0DaIqyYiWrasFW3ng4W6K+Vp+ifZnoPt4sbKGWQYzTvbEHArs6u
hOGcCn7dTJh1gbNy//irjCSxDttUl9tUzOHDUXRXjyAyWGL/NWSaKCiWDy4LnfZEfkZ4cEFy1jA1
xsrwS8eZ+PJr1Uu0777PbHvhSFucUTSlSPbAJ3G/KnS92SIudq11pjikfXfpA6Q0+hBmT8Ue2zqP
P1mHuBiZ0guLjXuviSwstBDEiHploRsvS42xxO0J65qGvdxR6Dm0zV2hvvu1Hp0UDrAKnH+1jYSI
3i/M0A8jJMpKLIlKtf6zBEZmCBaRbKhHOvUTPFG4AS0+GEs+aFtDxxhW9pTcxhXmPNRBqW6PB5iR
K7mSm96FVPIUom1KP+jfxvb5Kt5qpSI1FHd0mRhAlLzE9JxRKV2VZZgSa7y8dmiigcPglEVtInd7
wLqrGOqiGkHU5JaUyOak+BaHC/KhpfwizclyHaLvVMyDz+Enlu5PYw2QocBOW6ElZoL6TJ2UCcLi
D8w291CpoTzP3X/opEPVICPv7xn/5h04RzT2l8SkufwEamUlJ/SrzuAK8YxJLKAG6rbUdzcbm6W9
5gyELwXUu6WR1rdfsgp9hH75MAdpotVZRq93O8ZeAdWCM+r6OtFBZzRtcwZ3nAggYa6rhVMNSCBP
B+B90tMqlMLN4OGjMqtD+BMiIimfRidiPb6T1WrOQJU5MJEnPTFn5XCkegqE1zpoDFgdc+Jfohvn
z6UQvsC9T8EsfVUkKkh7WiRZaEBizupWpiS/Ib62jPrH9FR+d7huF3iN1MYeDGElKaXrF2+puyQa
4Qyu6WjVELvCjir2sqxqZ55x9KjFc/3sSuKo8WrcXKEmGMlnlqm8kRNAsW20OlYjHY5Q2MF/ngZ+
I8a7QmIEDBEfXluJ2w1Yq1pCdiOrQJzENQnSmOrYw0Nwzm0xIHb7Fak/PVwYxGr5wbs3gS4CnDHi
U7wENq0w8crFtV1jfEZWR8uyRW1XSxBPMgq/qMSscgDmzT55HpD2YDl5ijTubM8ok61+dqsMEBBo
BLzb2Qb5oru+PIGmFe1FCQYhezCypNm+luLOuinWRl7y1gDQloRWaiWKKu34NkmT+LKfRKzNJ2Kb
Xj7TyrGCmINVWiXQzTjfmn4wKWNy28Oyr3qUd8B4j9S8b/yUF/AB5mAMdyE5C6cK52/RZiS9Urfc
iYU7Crtln9vBu8/JDREPaYRuELzHw5sgaBkBV3hnGQEE6pVBFGf3XdaHbFvti3gRDGk8zjiiptfM
wsbUNlNWHaj9JDxd+QSFcxmmHpTp7b9Jmjc0JvRAFlVJYzES4H7tRVByhqbc3SJlJZLtwBKvClJx
dEUmXnQGFz1oar5k58iHDgCB/6B0+pP9FVFgW/ZCtx2Q6PAlqovcU64jxEDNRxCHfeuiBn1/VqP+
Q7erau/z1HAptlUky8dY+FePtwimmtPec6qpWKedPT6X+X+tN1eVSNnxqB0PlFcCPM0E2bBCrn/j
4ui+TnRYDK4ZEu8nx1wcdqoF0x4BqMhfE7OxJEJYdQ8n7Ku6QDqsFkpCskNa5dDlTdWBQqNtXurx
dG5TaDFUEtoONj1eWwdn7G76VYp6iJU7c08crKMx9RuuEQlOClGWRuD398HaY4fdszribbc9vwkW
tNWf75VIliLKc7O+NkHZ8Xcc4FAwREFrxjphO9YL86z68Pkni6yzVaBL+OUyXUUCz0CxxmM0/xZQ
duXrc9km6VuWnsvcH5mW1By/l8zIv3iSedF4vs4xnPkKDy+KGTYaWG9GtmNIssTULvDKC0ILjJeW
0dAhZ8+nD6RtEZfy+N+XzYv2GXCZjTGX4KsWt4h+LKwt48CzKfUZ1ucPVEukWgZghHnMUQWLsfKm
rv7PlMlH2133Z3xLUkrvnBQA7AxMrvcF1HzfdVG522qawFYLFVJjEVJYwyUA/1Sm5M2Jh4IK+rgY
qLPVwyaNCYa5bXJIeai/ttkMTpEJWcasA80nQoas455xepXnGnqd9H6X5zdKP7VtENDKLC84NjG8
BglhkK0OH4dJBiOBslxYN6/jzElWEmc/duELPyvwRbqgyL7oFrizxeztASn2f3V/Xn2AMTpuHpB9
462b6VjiKoDLcmemAG7y7sCxo+FUfvkkPk4gFMp0FlNeXamOS0SiBv1+mxG8Mv3Lg3HfS2uWQL2J
CG+jY6LjJ9LVon8VVXKbER/tjAGAwGtAzUVOasTQYt0pndA2J7Sls+bZ7JNy3Y5tXIK+KdV6kFSq
8SCbXvZDy2wxYT1WempKjQObzn1QowRKtuoHYXTPtt8i0cPB8JTS2mdloZERL7uj29ExGXbMQ+Vw
UKozGd8uEfTpDjDeTZWK8qaA9+rUSNDTW9sUmbDmfbYwp01wIXzsrJQO1DHA3qON2Nlze/tlUzHU
HX/+FsrcsewDZIJ8CKtGtdUg397tB4L0MRluud7L8nGuczlWWvfKPtkgNnQJZEgK1CFtlgennm/3
01w7Sg8g2X7ekvfAp6gxOUbt7IaMJ84vvFdkdK7jSvrFyPo7wjpXVzBxHjoLS14C9E4r+bPP2Czn
TXAl2QBS3dr26hQTaDbz6hlSfmIJQV16bGRjOQQg1PJnEpWhsyt1XAwbheMD8LCKVWts0ROpV9Wo
GVhLQu16EMaujBKBXPlxXTrW5ciZxhx67jklphTV4ZEAxIXpMsg6xk7uAXr+SjlF7X3xeg2mQQCp
90w/1KiTlr09fPpdY9u2610Wo1wSOK4GAgDh8phl+HJpaIjLpXgtylc1WFpV0AHUTP1bz+3HDUk4
ll6ywXOmxXIM+72z2uIZN/J3EwHkFJ3yGilzOGBF/S8yjGIe2FqdSsG21VUdSBpo/jle9KyQa6hj
j6medKgHe3N/wbVoA8ykscue4B8jdzlsSTppxRXopc8tQKWCgMuXRq6nZKko1zCJvgA3E28PWT2H
kmUwMFBmM6mvP7dVJrc7vLUXBPDw638wIjNos21p8sHm6oJhe0p0hzK8HmMXy7h7VF23P1YSvroT
gyAixfXBP07JMv8vGf0DKfUNXxKgFHhgb5vGXx6CpWqECKjQh79V1TrGTA2rS1dksceIADLu9Dzw
gO++wMBnuZzXUY+TLi48lzjMYrQMmBTsjz4Fho91VyrRs5JSLByIXx58wQ/YH9dxP8qJDZ6Jm8vc
Qs9lTJz9NjCDXUeBzmBVTblSgPDNAZczvOdTy9nulCt7wteAAaaCmrnXqkPQ3UcEL4dgB2R/NcG4
VF7RY56pmjnwJuFro7htATKdyMitUnyCeuHDyXMGPT3Il8DmLxeZx+L3NCIGJqsrLcoPUSwQV/L0
AK6l59Y0/I4EP2VWdLfxY2aYHtkRPm5193wJEa7QrgyvGFdPxgUZj3WoRJ5g2zWRy3TJfnYtisB7
UOHSIcrgc9uF0GXnGnETA4eJjSm0K//geo15aDVn+OO+2JI71PyJqaLPFGl+XivgaiKxImX/s5XK
wSVl2TpvIT6XFh/G0gleXtPGQ5K8aYOMSbpXKn2/o6D0Yc/A+fvoaImWzT218qgefrjztn2IhzeX
eqEXrecgzk42Uy2Ck0MbZRIBCnPTU94TT197UXdytKg7HL6iBYXKzDqD7U4bvkwp1e1XB5XUh5I3
aNYJV1KC9gBq3mmaR1K3XvtxdPV1DkrdcMSED/RcSc7SLb0wGdNI1uIN/tJxFLM9XfRxRvnR2qTJ
AomPM9Tg+wgztFsAa5XP7pE61WlV7Un/KJlmljd3LBy5EEalxqmrOcF0OcXMcD6SPWVGMP/Eidli
+aO0W/Z/+LzC2rEZsiazoTwF2TsJgcBzhFJjG2G2WpNLc69DHUUUI5ZndUK9tQzCjteB5oXqblEk
xb7O73uC03bc7b29TaJsLmZaT6Wy+uV3OwKZT3dWJWCMwApfD47TJB3303dvgXJsQTSMIKjExcDk
pdwnCSqV9OFjh4jqujpvgfb3Bw1QojB2b7U5KU61Fc+yCmwkGlaw42hrr2JGYaPvyWe+4ZYiMS22
73CM6c+xZQLGdkKg/SwzOlG12K+cJ0VUc1ph2aff50OcAplZXJWwVW9ZmLfhW15B1zQtXsDo6hnL
OIBpeeXzrjuf9Gi/X8gLvSeyjy716nkJD+mNA8o9tjyxnKMyfU3gq3W9KdVm6o6DOb5Qim080cEf
sCy13uYxMchs1qiw5/X6nAU9bQOETaO4fj0wBKsf6ZxVwo8cIR+ZaUpWCVzFwfkqyeL2q8IZ/Iwk
1SttLmCfpf2TCD7+fFvCEC0E2o2K0Y4l/Y3DZVo1d+Cx5gHqVV0XyGSPS8n5x1Uiy0oE+QZ9dBlk
QOxPzyPlQ+ge2jcaBzNo7SkWeDsQmphIljVFG32+hNr3jbZu9fJ8oCOnYZQ6oGkX/6YyZCgMv44h
VHBlJWJmlqFwtEH16hGznY/nTBDh+as6ZtnOLoGEZ2pcv2+Vf20x0UYAr0FpJSk04uRMVxOTm8z0
SAXpRNnQN3275QeIS8oj+5evYWi5smSl+PAdzlcCD7N0bTxVl4rzQSdLnWEObWgKYrdW+nqqrP0v
KPM27nzVCSouLwq36tTIjPRchnfv/5OwHYMDsVIzBa4I62HKx/7lJRYvyrUzOV3jY4IIW/yw+1ro
HCKhzT1T47D+8D9UbMLT0tYzYdf+M1PUY0fNWN8gVMGYz+E4+QwdawSZojFYTCE0FWGlsTc7NPtJ
OAbZzPtvONrlmZ7jrVT0feGh8o3Jm/2I22TmnooKj2oA/vqQ7CxYjb8YaWkn744ph4HcHygqjApI
yqLE+Yp/xo66rdsvIKckWgXVYhRo+8USzSRIKBW046DBQLgdlvXFG91211Et2MuCcpvtXILznQeM
AnSWTYMjv921TBc3JkwWjpAxFMhcah26mXyn3ye2F8QeYYHuui9ru+51MFRNPGnLEGazBbGGPjUx
TP+J7PdcZKzf1BNVhHyq0h5ax/1n/Qdn2IU6sQP5EibgQta7CKRD8lgQ29Hes+62v4u64BY+PLqC
cXOslPc+MZCYgbZ+t5MKe18qBndVpSEJGXI+E2jeW7W6icSTaHmPMPmMQjsqSSBcla4vMJJ0qak7
Zy6W1PCT3pA7tKMzx/mrP6G6LOMl+UyzXvBc4cXmE9y2aU0cVSXUkafwm/UIH4TNQVu5lSAxL1th
TYkFD7CpDq+c9h+GQblNS0ueCIa6trEkXahN9/a+vjT7VWhk8xRVXXLqWffH+OQs03oe9rkao4a+
NLyzxf8x+y/AuXJh+GO7tr5rVkhfIjqoQUyuB/jeI687a0HVrGT7v+s65lRdFn4ZSMev6gorjG9/
r8QP4/o0Qle2CiFAwkcMRIwVBIljPlmhkkFxaD12X3/s4Giwg9SSiZdkmMzcC4q8spE52Z9B2rTU
shp0Isl3adBSFREBn/EE6rHJBKcSkjTACTs9wWRsgWhB35TIU59UdHuF3SoiZL+5rHF/+0POUa0B
kJF0tYabw9kvkVapBEAUSM1KcsLfjLN1sV1WFpTxpz6+/8wu8nhZFsFAGK5ACM/FB+bGs3TU4RT+
s3f1Otsq1LWcgRpbBZZM/eUcGU0r3ff/vFuvfpSqfqBzHyX/L3ATnUUOIg+YJ13/lc27n9GCb2Lu
SIMIeOIB4N0el2vUFe3+PwkmhX1DzrERciKKrLIVNKWvXX9OAeXquxlr9MC3Hlea8lBkcaeQpgzS
srWxyQhhEFuHcr3QRX4UYWqO85MhegdFNS83VOiASjfzhybvaWm07rhLGdzZ2vMU0j6M9ilYbGRn
a9pjLFQJ57tu2yolwowzZcogoirO/ePuJifLsbhNbwwz1RcX1ZR1AxH8+91IoTm94lkiV+r5W4k9
qELiwMgzDZFB443Ch4gFdwQhue/FpDFm8Gtyb7G/rMYuYLScpBNi/gAynU+Q/YzjGlRCXhOxTMjS
yT7w2pifULwBRmd8P4y6RnSZKSwizRqH41+6Zoc3+8uS13Tp52A7YeBeXo6l0juQW2k6b8/B6CHA
ED5tYbaP2wgS86TsJzEhfZG39CVr2BRyb/HcWy19O5YgL88XtymNMHDJy5QlvPpmV0PcNZmjV9cb
tQA5jww88L9RC8Pczbo+r0SNr8mYSdY1n5dxLDcVnhxB+sRDQ+MuMWK/Nn1bJL+09LhmVHiaeD6R
OiWLXusYui6uo5Uc0gQxxwjzBGDrewMNwwOGefq+4Zs6LuthD5K/j1lfdZ1Q8wtR/3oX971wlEZ6
QZrIS396pBbvwaKzTG7QOEfl8n1SMaxE8d6md6er+jun3kVm7z2Q7X54FAY0PXVwWMGQlkWXKfXp
GvZG82QrOvGMZC5cMNKyCajCOyuwWLLcenlK/J14TgRhFp0YAtE36q51jJKNiaFU+tN8jzH/iDCq
B7w5zU9OUml7aTtvqhW6wNafmq36k3gSoTrd3n6pg26cfzHYPIPaQHJNMia4XMSA8YtCMbPW2g4r
e6psLH/hV4vPMd5lhYnSTR8QqWcoCPAfRqbf62j3qrIjM+tsHR42xOzDDDG9D/qPx9eRo52krZCb
b+ZNWmjcm+v6KEfGVU8RHqG0+e0tvydVY6AR2nfqYCsEoo0G+5Dpn1CIAd722B1X2hP4h1q3Xp8b
eeT3ia9uWUgLqYEP3Md+RHiQXwGQxFWl3OQTjNOTwS1/HBIamkKeIYvtTrrhi2f9czBQm89daggB
6vujLUD0Opeagi9U+MCs7gixxFDqT+x0XWvwMu8jOyYpz92HUERuQeD0dEiwDmqAWHKkbB5iHhfn
ZoNeH8Uo36cHJPzCeFmNvtHXz/7KQSDbxKM6+ELc2koU9pUD1lpOIoOLR1u5S8KzqXRhLjlcNjbY
MxyDTraDU6bEk8AjUyzCToy/P10k4ml8zLLPUJW6zKt0bUqzwknYyX5WvpgydVERc++CGOJO5aK/
ju2BDOndD43Y5GOTZbf2MFYLUtezm5JQ3ZWyyBciXTSpm+BFTanG7LAA1ovfdlfam6yKH/rfh75+
YG01n3ZRkCpGM5PgGykpfGg0W8gSUPsXurvUN+Gb8AL9u5BiX/GxdGZTstiTbGzUEMrEf/kaB32+
oP/h74meaEBE7sEllAeKJWmOXdir5sO+TX12mvF+Yz0srUmuCHSORFxqQ8pS3ikEme4q9MveBDzU
yizzDUkzkO9CtQp1E0Q85lccAlwWMSA6I3RHXpKwUApumeSjQq0DN2gR61rUUlkV7xd2l7tJw0Vh
3E91+S0HoqD6yeCBmms/fU1/miAnzX91rxqeqHqlALaFrlgE9Lu+u54Lm6N7xaiRH8CK4u5gCYra
hEfwq26r3Q83O2mddPeG027cDa1KF50Ev6ZEURxWUbd+VEiIy9eUBCeH6PQNJy9+KkeZlhoIgFg9
vefD1957Kqz19FwYTgbY+it3fgr3l5criC5mWDjzRKXt6uJm9ZFRFA9flIwEUcYY+X7cx56V2vLz
p61BoYet5fwJBuuQIfdhmBU9iMCM4Fgvcft05GyCOYhUUAgUuHg/Ehfu8BLslFxu5dHP2p9cV3rE
xZQP7fcGcVEAFfIFmzyGyFgXiIskNe0SjGBi39eTB7AIz7isNK+KNic4duLb+TL0Y2Icpxt37aea
IFAnSj6XBatTPV+8Uk6dU0gWidM1UeqUAhpMUqpKcQTs9YH0sNiPA+Hm9g8/bFgec+zPmB74R1my
07HeT6E0KxZWOrPYrQ9YWJYIzNXjxpPoR23xVCPfVAGHiAjJSYJkZ5Id1Bqj7ayIzNi7cUES53Ec
vcNR7CM+rubKNwi0zoGmONHEW9CSacNgfMsptDGYk0VICLfTNEPjqHGq+mF00NdNAD2cQ/8Jy6Vv
ErWOonWylshmlEbbQYh3hOoBGasx2nTNx/tbCePFmuORHcbP7K4YLMPkQNhxf8sLXqwPwsRvaVR0
4rEQiRzW422ZKRj815CdKbpmmU+vwL6ja8wqN40hzJl1q8SLRmbBvkQwPlJE/iURjWxDEC9GD1O4
BdAxluMUii0nBUpq6Hq+IQcQ0dk253j3GawAsOOnE/TW6GcCR8lvd3wv04AhPryol3b9ee1sDvy7
Q6KpgPQ6kewu47LHeY3fsbg/M+LjZCKlv7MkPKgsQjmMvh8nJsCpOiyDnHRBAp+7BwZU7Z1wzv0M
GWoBhL23O8DYjV8kH2UvLZ4YuVBUVI7QFqftG55kUZSIehQiG2zhLLettmKSC2dVC976ZOkXo5Q5
qXfMamPfPSJ1j4sNYxINlxaXEUG8oFEyXrLrlMARrjo2RGPHndsxbN0xtfUOXAnCExk34GjBUIX1
8toch/IQBBD6nK/LL5Y6rsGz35laiZF74U96WFx+6CfZbAx9QzJDbBx7Fhr3KSuL0PfGnRDqHjLl
TsVlWzJ3FQjfWujse553Brq/k4XbAef/3OOYKpfPCe7KrbgWa/i2Mhe8nqbIevpBxDXeQlrlhekt
wLhDATrqIziZ8hVr+LFJR6gDDCosxEoKEYA6dWcReVQ9ujMLVpzI7HG2E0FoHfOM0CzzpmBjd5I/
nObgpmmSQ/ctQhWUgOotiFguGizHf71GJLiJblNvUIdLEJjTJigqNgBYvoq0Naf1EZPlUZUtNDsz
ZX3EeZjkP4t950zWJn3NNQHiIudiecRBYVd1tr12EqA8G+yYNkG1MUTEsyjUlqPnwlglJYvCutdo
qdV32fiwpXIzGRwphdHE0yjtuSjY0V81BbBjsvnLO8BCSRBt0G+lPjCGKbUccpYAGdovUFVR8oH9
/mm9VYocQDBxTlXY7r5gxVPRrFQEAUdha/qoB7esggXCuOwHXSF+ms7fiEn6UFI2hVjkoCOYJsMF
OY0nqOcJh4Ig9qxwAjIYP05k25V0pZqSX6lB/8nMNH/IG2w3B1Z7UH1WJvkDk7CnzOvMidhSd/Yj
mzJNXY8ytenxcXsmTeTrWfKBhv/EmMOMCyYLy8/NnyZ80YoEHhhRthLODyLW4J9JxAwpR+z4CAOn
FkkVXaJaGMPVJiQs5zMxy1/E3DV0CdBHi3za6F/wGybO4n97XHBR9sv1zuuyMyE/1ebphFLPTwTe
/7BD7hJIxtXSQJSWuplvI8NHSnodfBwXJFdQNAqgUkEwdOanshakGAf/sV92OjiCLqtyens7l+HK
weUA9Ce57ewd5dgLy+417p/ay5dHC//EfA78KnFuuVYYDBAU+JyiOBpBJRWuQ0yjn8M7rZ2C7FpG
ClRHKqspzXqs4dn6rHdW0mpXYp2gbUQerok5lnTTui6KQ1gUu5h31OaIrmE8vStk3QQCQNMb4bLi
MihBe58Miy17T50h6EPSJjIpn8IWKjXHSZzJ5RlschdYQVqltI7ox/oJ8tVQYJjaL9H9wjJPFETJ
dQicpkxYCpydyuGpBrtdtrxWhDl8L9xx
`protect end_protected
