-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
SVbJcIyh43Xd4yLEe9FQupQhPrs0VDCaHhCC/W2JZzpvI23mjYRXwHv5dqchR2m1ZTdP3Dwxpeax
G5hk8V46qyxNVJO33I0mO93aZwgjiLqeGjLnoJVFZ3nZEdaMR2sQdZ+Hp0XuEJ1zEWOp+XBPfSOO
y40CwgqeV6xIF93vQdNfVkZvPSImRUfd7X38hlrtjU8BU1S6oUf1XH2oMdxtc+b8XOWpMwKRF1bq
m9o2Gx02KQ6lvmh5/jt8fEYrlxT5+0G4a6WSkKrzVmQXBcdkmqsp8VhZToZzxX9xV40UsFb7UKRD
9qgTXMQ4jmZcLGlnnR7QxIDD4DThlKc3AvUbCg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5312)
`protect data_block
e52078SfLMZX1iLGNUGC38auzCnJ20jGDjTYm16I30VekG3zKzdEqLUXAuRpb9SrFNtMlhV2ZUDi
FHoa0me9ttQbQpqUdthFqGgR5VHKY5gNfCZxvMaIeFyYsUiHog1anW2iKUBJlVj8bZxxVSGKKeLF
C8kfAQZYkXC5Yj4olsSXURgYGRv2hQH0oXUmeQzecNwGR3dVgt56hEyVblsBat9nThiUMYVSgM6s
UOoLqaKcajaeBTHTMVyaPZHMQstIMAEbQj94Q9CKrIhBZvh5EkesvFPulzTthRqydn9rzsQR8kFj
EE8ymrGht1kljPu1QWq+spOd7sbD9G1rvON9le9hrLQUwH0ndyLpLIHyo7e3XcxOJCGZ6E0nmfWM
1HPsr/mDFX7eakZeWgdHgKPoU4UMohs88d7j+JdaKVJuYTAyjfIKObHEyi10yxP6Rk6uENIhq/8H
UENObpGpciVsCYoAiBDhmazvdn7mVUoMRdnBeE6UZLXG1Qiy4+fVvpi+2d4BeWkV3Yh72UEycsNe
G19BXGM0ve5ENV7aGBxtVlhOJ39GFXh8Pllym/45irB+RvcsXZTVoJCh7/n2LrxPunonKxiUkvk7
w4sXc73L1PmoXglOjXBzcWS+0aacuYxwPtKDs777IatLhMl1NlpMyXc3BbhMMQo+bMeR6FcYiL8G
+I5r3Ssk8LJRN/e044tnoNY7zbh0vMaXj9obl8js5H5mCfDlPtRxLCz2zZ6tMzd7JqybSBSab2cM
Op8yT3PDN6q7NPRZmiuyfrZgTCAUmtqgUwLHb2hoTAg0wIx8JyO9BXfqw6+ssIlv9DqT2MIyW5vV
jrPfA4A/SyJIx9skq0nyqio0qw+XkAfcRrM4EXWcB860zpLJgnYFHTzSqR2tfCl6lC66YSZC8oJ4
yAsYwsE5YV9GuJYSQsnGkwsDhxow8bB5CR9ouuhwQcIdjeFtSCcgqEt9LOLp7nKEXFOncfseFdJu
CTIiL53HUsl2E3jAtk3+Jl2uSLVLN+86QAN37iCP4xfb/EIoQDATTuEbvmZQnrWygY+FyJvP+zei
uhX+8PKwO4QXZcmCXOz2CsaBshB0hrmLWZr72PzebPNsXORFrjzlfpBRyGK/BKjy5LxtK3IGRqb7
USHm8nL4pfEweaDs24c62ileRqAcWQ5ws9O8VO72+nq27LE+XLHZ72rXr9kottvW3VkimHtj6BOo
jsln0R4wCO9Y6U9Z8Ow9Ew08CFEUfNYt6+e80RD72ihYxTP6Ln4hEn5WJJcoAZ6N6LUiLYsB28TS
ltOIJTt6cMQJToJ5tM4geYmZSopdzu27odYby8q+r6T8hNn8NyVIIDDz0jLLM1hAgFKr+rDliMjf
zuQhj6xlg0Uz0elPCmPjXFHlDl2Fb6FRe7HpET+8IfPzX6w+JCAWrkF2OKR/V9WRZy8RJB4+JzIq
+0ySh7fqpAVIbygT8EuAJ8NXG4AdFHTLKISVGnxLRCeOkXCl03U1QHqhC8OfF8vmmTnG0c0u8Oy0
R1IjqQmRkEwU7CkrGNxtiLjNiu8AJrl87OCq1RGHekfRejKVparewBBwNC9NOFyzGXv7RsdUl7bZ
FhH72wSpdRYGYwItHPRnBrXWFV/e0VJKC0ZZoC3iOPsUMFAYRtgyHauBuKJzFXVh9638v55mNrp6
G9Ut6Ec3YW7NcWiacXUcuBEPx6KbClDrv8LIGsAAyDO7oI1bh+zWZMQ6G2C9KTEXpEP6qZqarn0H
RMxqoHVhkmXE5Ey15Db4PWOh5OAH9i/XvdM0lcRm6qDmEBTvYq9BNkn5TZrrJF6We/otFBEePA5N
uKT+hMXCIihCkpRrEUSdB9z8pkfd3FO86QsPbg+pQJ4YCAJLPDwxPIKJlrsD4eLiqG9pFkKsW/fE
kCSJO8QHvdaVi3D3PXHeUPPrL9jMmwnbRnaw0sJ484IzbLZFduBr8givEkseFgd5ozV977f4QkTL
AC2J9dRuhxrRjEwIrOJlsdgnQnwbzPWt8SGPxT4Q6qvHx/RiGHcMyXqJCAk/OBD8hW1c+Ce6wplJ
WYCq6ibmlWwODAtNLe36pTN38MERyI3iT/BGgG63PNF2NYbPnxsfC5XCWxf88aavw9sVYq9N6Hwy
BYIglR+yVaVG36hUwj+5OipkbFNTy49QHXJOMojp81T8na+5VUvyHjjsFhgiVNng6Q7J5J3D2rwZ
c1vCyEuTAc3RlWLRNBFBZs19ajvY18jcddskA7dZNoiYCAW2/sr9PBzlqxm1pCJJeHTWEUVT1EL8
3eTYlteLw3F47yFv1w8NxQQsTksdgqH+enYMl8n87PzihKL/QMcvB7ojqqCvGaxkZDAtwg7292xL
kATsq7Y9E8fD7y/b6XQmO5APdP+d198PnRufNf3UEUaRG/Sb7Hl9XxHxOmgsGnWUrTJusloCqh1n
gabXVQum6UIqHcUzaCWesOJfNngw6OgUfJZ1rJrqvSowxaZUsSWhQdDMjY6tbwtaLI5MUnJlq7gZ
ny5e621mSzf6ng0jBzu12tpltOfJPI6dCfs+zaeHVISMzUC+QsLdvHhZm7//Bm+b7w/0ZxoqmI9L
gnOUXMjSVwwozhCb4GcGjbOyD3Xf5EtYprjM8lGeoKG/uX/Qo29ZrOwJVMLWRJaVaS7ygejnKvIV
NgvG+x12FUpUHWBJ8bw0RlDpZTY39V33WK3dVATrBW7l8xEDVLkYjUY/vDFTahBBmVEpwXiZTXtL
zDFIEJEwGV4aAvKEvyZoZvSVko6EQg+Dtd42mnYH3c3WEOEahf2DE49uygIguXl+stOqpkmdNTlp
h97MX2dXwRS0eW7bz3YaYg4pxpx498mqa16IJPPcruQuY2Zf9aEwEAO2FigcRQXI2G4n18Lm1Ns1
4X/LbNmjd9aQgfar8Hr1uQPkfAJNMXP3oiRBIQwVsmQ5sGmnvteh1GAyeHPbE80dpiC63NU0cJ52
W+dl0wDAnTI0SB35ntsjo+EfKEHI+KfxjoDZ3v3khV8pnJLXy2NBSgmtwKLdNit+WcE/vlH5hV+K
EUJuKMbplfNEIXKMydB8BKMbGlnl4jo0lZusPvJBN/TKnzW67OMuVOIg6fPr7qYH7YeI/2PARf/t
Zt/sU2Dh3j9Xg7vupmnTe8aS1rjr0SOxC3m0X06B1vZ4gX/XciLXn3H5HPXXh26cwCv6kXGFAG0W
goe0xsw6deRwnTFoV+v3G8RBXjEtIhDjeUZ+gNXxoUO90EHnhOcjwOrghgfBP+XGAolMmPiZrwmZ
NK+sVw35c1WYxotIcrX8S4SbzUq6yxnStlbUw4OqlkC3C7O+b8vJnL8J4+TxfB5toRtjOcB6oWoH
SR9l5wA6X6nLZgKwzVkjzy67bXjicVUB5er7a42UM2MSpYcV4wgFsFRxkSzaFB3g4nrBMucfgz4+
MK88Dpp1zHnwBhykPnBLaYQiMvPMhXrjBFHoo2tF1KEn2l6Id7Zhp1ILdCIgv1hjrFc7pD2S0CSl
2ZMQ4/2/lTxDM5nN6oqXLmXXTX3m0M+3ACmnqGoXvfVjI5/45NCHyMOzGtKl4VKFvXGRkISF3A+V
Bd5LKNum7jKNtyCfYxV4Ty8kYDxS5re1uboQI9lwYPbiQx5qhUK+RU3mm4mHYuOW7w95vcm5CedW
bVKPfoc385hAs3pmkxDMoMevT6nTWfpQ+UfYFeIat0hGM9tgLRzm4W3mLkG6csSC0wPpPc7pGRzh
N+reHh71adFGjkromiqwjasQo1rE01xih43qHk7NFIB159WsXJvRQ55HOEWPUQ85rorHLmTJ90qR
tNodpDri4FOAtvdESb6ob3liiVciz07meAh1rynts9BpNuJq0+kfYO6hbnWmzZxuSnv1Na2dHpQI
MTzE8/dKzlptjDcE/dphPjQGsOwXs+RFcQafnK+WUlbEl+HrmmxRh6evvHpeGE1lX3pX0VlPT+o/
YSrex+Kgqj+ugbT92SGiIlH7Pr84b+jDepMwexPVhzD/moP20Phlq3VKgROgh7hG0vP+GGyzE8pQ
E2u8fN09R+fLq0Tm++wc1I2O1qWPY00FS15qn+H1PNOcvN7YlWCWOFx34VhKWWcbp/4kV00QpUWD
yZMiZmAkE6uLmvjtePheyo1nyCoplZou4xEy9lqLzNw50sR4R6G12pAfujLR4kCK4wNZQLG1b7uh
UPZP1lMecxfLNL39r/E3FfxFzzdh1rqE1bIcA0Oqjs5YuHqfbe6pOtvE/n4foH4msSGHOq28UBv4
mXvUOqyT8ij9hxrRH8o8/Wt/ruwFpSGsTCBPuecMzFifCM8sTc0lLaJ1fBgn30s2GGRv2KDlHC1/
nLdmFNPu/UrYlaW0tHBxzEBXykYg3V5XPHzIZD8Huu4VcGVMMCIjIYkY9DYnxG10k9aK+nxAsUnT
z1DEM4zpUw9hBcAaBgrWeOsQ5XXylG3RgynowNFC83rbouhHH7BiGA0k6TrqN+lM02zps9viVfnq
aI7ceKraOUtBkBcf5eBeGmvQDuHLCrosU7/niTPDosQrXlL6CwUbMuNobIfszlwpGCjHbWFSdnXs
VAIeav2RaiWx6OZ2BcWPQrkCF5joF35q8h1wLbP0kx3QeTSDTtDsqFfL2fjxWF5inr3KjYuBO0co
ae23D8zDC3BihTsHgOKoXJUb3YrpAKjMaYw1/8v6GgLH8hVb8IwzSu8hzIYsgsSpw8wdw4vzwr/C
Ph6iyXBaLh1WP5sr7IF8eFPsBCeOu0Ra43bQZrS9bSDEERkcJYOr1Wj1CKEXbrUHvokbQi7Zd3H0
EXnxV1c18aWrrIC/loNjc60ZlVwOuJSd6UlyZoxuhEjaj/0XW/oUKjc8/ijqU+RQvGivLZMn3K0S
yxLzM1b4arbk1UG2VPK+iuo1AlCtD3bneB1DyybaSQSNQNbR0+RVHg5heu/MDipGKrSkEzUuK5dQ
dzWkamiA3MNdBcwJ4Brjr1H78e5Letj53OA7t0ASx+Pv2Lvon2JQb+n9HAVHVpo2MqvLC7z+6eZ6
OyVLykELV7sqVtNQsnoUv5IsuezXSbo8xEFKaAKBDpMIzzFsPIjhmBwsrXA+AS3HXjs120U8oVEQ
5QZTWn/gNNUnTauW7JGmQe6laYiV7SYLouYyH/mv2nN08BLvLN0NHSGfEuAgjDEXBKF7t523HWFE
zYIAuRgOqOFmR9Nwi8M2IFoSU9tPjK12s9pQVxIedLxmLMf/AXhPZ9H0BTZJfKN/MywbwxCl/SRe
sbXDYalIBI+O4hjiXY1poIoIdpMFPwy+OO60jqyXmXXFUbWnqK04WaHy0Fnbf8GCXOg3WCdSqA8Z
P5ZsodVOFCAyIBhfCCBqM2bNM9C1ECGGTqGxmpfVcublk0+BMwExmPatSRjB2kUYarYPhejO0e0k
5LJJmRDai+/a/Tv5Y/a31PmvEOvxyOSd0wsgS6kn94ZOhF+Nz8XEWG5+bwKLI2TOpE41BXXdQIdA
LGnEJBlZ+PEHk5bUdn82I6GIRryT0m9EFTbMToTsFNvpt7IKSIXkG0+MFkig9KxmCsoBJj+QhTCf
045DAU1rVfMcKQmeo0EMeGGs6jatyYOA7tNfcDhTKuglsJGn5Vg7P8bu6ZTx+WGV0f6DrYIEb42u
zG9KddsjokRLWBw6Me6m9AqI/lJRt2tDlcVoyEhm7T+8HhnlCDn5cV0NyO9HJtN+ougxh6iUsG7r
zsnXt10BqC6mKZxyxaxbv+P3M6w6Cle6lnPdKVPaIcc3gY8/tgzN5XtOvUodcDtJElU6WtmYio3L
d7AeoRL87Jrrp/TpkbrnxeBky68I1V6atGKeqASNa7M4ge9BVWL8NAJd/PuXFCQ9LTUzqfm1HtUb
O9+oNPs2hHchikK/offU0TnFuiDyODPob/YZAcBxbL7d9UfUIoRarlENvC4DGhAcNUe8gFUs07zF
Bq97fEao0W1Svs8L5Ir5uoPJfjqASaG3XVU+EttDkEz2FCkqB+Ec2h4bTjCOmjrS3tctF7sWN2vX
6meaNIqQiA8LWK86U0Qmho8owcQNkRZ1TOnmKsZCYbuGoc4V3vb49ZfP7RJPvHinZrn/4BrK2TZT
67+vRFIamTroEn/vpE7116ExhjMSynUQIBd6VsZjEESkD1IDakFk0z9FlnFFF/O4O6IvLX33QSw4
6rjNNnK43mgCIla59YVbhYrnMcR6wp4lr88zfOUinm2zzGGzDYTJXqoyWfG4TMl0TiibdiKjVqMD
4LULqbdtYUmsCVnvJ1bKax1b6TsM5zFYJnGSWz5ljKg11E5NOb6Wa3MCZw7KEvJ3xvSNUY/4czr4
wPvuQxHdqzmkO85Vb13KwwM6sz4AfN53J7lXc/+HAmL/sxSaaIThd0cHCiO3ajaIPjswmI6NilvW
PtmVK59879+8OiTvXBCWEcPgsnZ9CeDhLKUEY2T6gQwr8P+tUqQlEtaBVlWBvCf4q0JGtliH/4rB
Nu3P3EFuKejOLChWjsogv+50TJc18NSE/IeNH2UGJh8K6V9o8ZyshWop9k9aZHIZ8F9ATomlHPF+
iKMVwSNTv5H4CIw94JZG1Rl2hEAsTN2AzMMb113cy67LU22nqbFKePOTUIqiqKneJYlsyXLqxkLP
SlXxce6IJ5TBNmqNOKwurVwuqmD4REmnXIObHTdcfkhpQdSf50/blD3myQicZd2UCFiwgRgSurKS
hsT/RPWP86gxTGTq8PyAT9WzsCsiTVL+dyve3oMU/o3lOZYVmkIvk8R7NtckqsR3Tnm8QrCDDnyH
1FLpfDkBLg22+e0XdF4rHFfS6ub9CUY01PWJahpw72FaSIGFlkkoap6R7m4yvPy0uuPSxFZaSGel
kFwb5TljVxlbWf7SSS0jr6mk+oNJg94YBQjv/v7UJsQJSp6nu3XHjow0pfnOjA6EQyZA4dnuM1Wq
upce5kNCiJ1Kx4GxDOvrEQlndpu5ObKvSqXnHXFD99AUyDw+k13SRtsn8cHneyxs7kNR/QTEyPIV
UK6CVYnCx7+pl+CZ1fcWsA4sMOXRS1BGfZcJQNTB0X+nDERgp3ifh3nbr/7/FUb9oBF6h3cbAmRo
WZigZfXq+xu/o4k=
`protect end_protected
