-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
vTPnvHBHRcs5naerxHAtolxgnk6baNvQeLgUEqeyaG/uS3mEh5j0wlhYnZ+Q8rCTLvILOgVX1t5z
JTNw9l/+m+onM9DsJ1IQp4WfknnuiW5M/fcS4U4z6ojq4Rs3XJFZ1zKWuZda1sDveixYzRuLOydi
tgZXpid9BF2v0rET0UUiA/lMDO80Qql5kyq1sS1dy/RLZiH5+bG2wJj/9zNVTRWsSP9aONityL9O
u3ND+vE46YcjdeanMtRhLSxiFw0WhL8RSX5PVSBdSt5OnxWL35BC/TgobpnZsYFwY356gxxi/rpT
gedwdPQbglln30hxqCTnK7V1UlDTUaURhiq3Dg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 100896)
`protect data_block
Cnx2wSlq8n9WTl2cghOWjRjh7bDsnhjDI60XmkXViM1fmxeIMYQGuhgfwhp6tmI4BKfDHfg4DB4F
JW2ltivLDkPatTZASyjZrykW+pqvcXl3JQmG8LVX9IrUr9s4z1fFQEGoHEcg8huTFq67JDMuHQYe
vj54j1eu8I8YkndjLv4pTkM/XVuAwo4MXnPb3zhQDzm0ZaVcNq9D4klyCtcRSv9BBZPsUBYIGS3u
aKQXtWLqeMNZXhi1KfIxXmqmVrz44pLGr4SP1Afz9MA4k/FH4AsY4FTe/Y5mXZBVn+1y7m5xjaP1
RGYZKX9p2Gbxnua1aSbiB9x35tRuR0ji9//5OcCvn8DkGCThgrBmJO8WVEd1i2TBgChx0blilY+1
Z3/0Yqt6xdE/tkmBCn584B6kCPmsiIyHTsTyBUX0mlCMTgPOsIjJ2nJ3DrHpDm1LHjL6+RhFXPN+
MQCJ56tYYToMnU6TQBnQZlqiBRpC5dZR3CY/eEVBjvLmBXjxmLWz4x86gB0eANhUihq6YBtOWAXd
uU7w4WaN8dDxl4aLrDKILIz6w9ngOsY2jLAwWc3ChULWhSmQECiSKnJNzThviiziDF2k9EugZXBI
nRs5znsd6CK7vLZhfhZCCP+RgmynJZUFsxJt8aozS0lkKvXEQD+f9FXdwXI/eJUWYaV1AHwW3I5v
SXpyVfghVyj7HljNUipIsIcXTZcBTVeOuQBFbyzkPSZwsMt445oryX6XFm63RDl60LRP+UmxMbTZ
eP1slkuHTusA+kiAaf3snvRI2iWYnb1XKtc9T7oh9Y2uo3aeoytblf7WiDOCknA8nVtstvRL3T/Q
6tw/jZegjJWubYGxnc2e1BK6zGXp4phc6cdCcHZuKPc+DwPSq0aGVRg9AmXGsUK0zgbWh2VQ0imV
SuffyirO9BHGk6upY3sMq12DqBZgxTcR/T1X9IUahLdD32AKZO1H4GZy7g7yQ1wlRfjKoWEcyHWg
2B6zI6w+3Ac+a4JfITBaFJkL8YEXOEIuFXXtw+iZUWpRJacjpTJMp8PHpHRIJfGiRbULKP3vIuND
11jne3kgi7+3U4K4IN4bNQNwyhD4QMNM4oTr0eXTSBDCHclEa3Cve/S7UTmpl6W9GIk1Wclu1uiw
zI8mLXQR6YwdPRtcfwbSKXlxqpQVUxJVWOKGfKPh1EjgmDAl4O6zQgGUW9H5wdP0EdsCvpWy3bBw
lQBezljZ/7EYm9n1c4YP4MEqDAz7A5J2E7P0fN39R3MQvf9GvAooZoT03K+tcp7YNN5R8zfDjv6R
xz4kNWvlK75QS1WFbtbsxo/yv3RePQP9IL+PIvxcVY/Xt0DnYfM2A0qG3oargUqx6uEkt4LWMseM
P/+29816tIG9jN8dmjUgj0F1G2VaPqMojKPNb52eMvGUHr+fjIchZFJPmRhSHup0/R2XIs3ThNBw
OYJ6hqA1/6ryYQYfB170X5S8bZpoG8yCgc9DctGxVcrSjSSIu+/v92xtEIGKbRSopmK2M/9oHQ4A
DMnSSqrNSzWqFObe3TUoKCW8uA8MVlzrLroLf0mhiqKxqvhCIRR48CX+CCcUG0YpCD+L9mjkoa0w
Ks9njJAUWtTf6kuvrnoDuZQpbvI8+MuOO4JsivgmQJppKKwOUrzO3OpbpTTfUcy0dyUbm5Hv+g9G
rVEGSBuXkH4gaOQfjgPH69kyyYYJmlhi98uL/bYQ/zQh6yGWQFCY/IvCXEUkNNPCQYKJZE+p2TuK
W3WLSYuI0e6L8NMBV2TIwnpll0WP75mS73avJlxJJ5SOgqj+KrvZY0K8hWYNtQpcG6ShUdyfv4n+
BchCjBKyp2uvYeaUsUik+Wl73BnUqNADyuU0ak71NXQ7B9cnafPve9qcKFJIwOOuY4VYRsOa0wyN
yzjcreftIrMBt5gcQmVAT5h7ye/ovngxTFqqb6aDS6U28UvPLVZ+oY6KygEEE/b0hi1PGUIyj+Ho
OuL3/M/m5xQ6R7xA5GsM5ypnJ+FQqMRzBFjBMqlygc6YTDw0CQ0XkQlud6hWi7Ca9BDu9bvxa8kP
GCUJiDcmQEO6Edt2rZzBObVinAhQAB2FpL2i/Ey6265RAj+Mb4Osfi8y2eE6BZTV8j+2vbcVgJ25
yQVOsUU9DcuzIpFJIGsrbT12vkxYsNrj5HiI7Zt5vknbW5Al8692JVJfX6KMdGQfKfCCahAod5YT
uPq9nWivesyYoD55ZCTCa9ubqTyonbA5InXRMtyaRN+2q8gR6TezRZTdZLX3rzouPKc1leIHYF/y
7K63pXroVy8a6tQIlmlqBKWjxMi+GkNsuL9TyVZdn7HKcfVhBojQ4DDXbMBJyH/u6d2iADLFm8Nb
iEnc4N2Ojr65TiPp8vALV2E9yA9dyf0qXtAgSJxwfyybrffxzH0V9lMPliuHaoMewHR97P07qWSm
ZV6Lm0aCe5Ksskng88Nbw6518Z2gEWugURguIE2siwYHlFIjI8wERX4Jr61mKsf7biS3sz6kg0vr
CONQcsPf27kLuCak1A32t1cMRO2C9UMCpjd39ZC4ZkRiXjfj9CfZ0EvDFVke1/MiCoQnlVtLm1gf
KjwkA2izuV+GR3R+Lroq6HKr1PGFM/80lIaa4pvzqo4PnqXtNS8pVgHiz6agYF3QhV0uXYyrPj4i
Z4t2dclNKeEIsmkxcb+7u7zX6VlrpDfN8oDWRdO92zoGVZVUbCD4elZ7uZzRTDHjOmqb+nsC0CxO
OIRKfTY4P4bsejhou8Vmov0c658LR7afEfknfyeUCBrCITWKNwdow+2iSvjk5TOsN5Ccm1ARx/Mi
dfQTSh5k/LK2ZIbcKiVS+fMh7qL6zieFvNlsuHURxp+DuQ11tuhcd2TAPzDiMatYhLH7kxtnqSrc
Q1kHF2XEuB9llOEVDSvI193OO5PyyKDxBjQQWl24r+FfWETze8PrigmxlP6wB/JLCOLtKCjAvtAs
yXAlxDAknCFRGwnZcGYh4m/HrS1z+Qfdp+ESnfWU/grk7VBiTstrj96IVhsV2mdnETykEqqDW/o1
pdQ7yGDl4mISN5N/R7poQOKe5h7ZEwZKHHPJxuYDoNPW+36HO05xnu5D387vObCj3ZPWddjtOJ12
US4VSZp5IP0m13PBhAAzDLygnwFOdiJgFds/U3NrTjKn6Miv6HI+/O41gDjY7ObkxZzXWEMmkutb
V+RM16Ezw0yByvz8aWUMsIgfDNMGTsuGQKwWnJdNT6Y/Vo1ccztl11vDAZKvPrTpPw4hmwuRYg9y
iU2S48DErIwLQtAaSq/XH0o4r4+/YyLSmocqczaS7xXeYK49uI+ow+2n/8mMRUilv+0n4NKVs1Zx
ZMuZUCMrK8rX6Duo/fd1eaWIEbbuq9mIk50rzqJTU/koqs3WPfH1XlNH8GYlA2/RW31SI7VSiHpK
WqiYlHAfkYu6rzdvswLbC+q4OM1WXRLx9FaVg5ARh2W1opEJopeaW3f3tNNdKlZN4JE1UQSqB5II
VYvx6c9aVFHQDa87DSAdeLFyXx7SlrumIVajyAtk88KYTTV5yHw+zWx/LB3BxxP7HBzgrn8d+OaY
RJ9OB9FBHhi1j4Jdza2xuORubVPMKrLTT4UOuA/1Onqgz8BnB6m16ThVV/g4tP/jt9anU3QBs9SI
wwUuG8TFmosOFyfmcfj57XtgB2GK4s6EvWyQ5qt049nGMV2NaBblOYzXUlCyLIlPAXL/0g4mvWpe
ZeeBmodz+QjwWEowJ8PgjfLWuvnWa5kpELwUxmOWVFqTr7enjClxKALM0xo2ZbSH++zjN9lXkbCC
7S1sEWlRILB5MbAo1NTj5u92SX2+Iwk/OEJGJlIq+rY7Qpr1BJBX/ycKjkHlT6rdaW6mh1hRh8wY
kK7IiDmRNLAxr7d71wkYvU27BhIvZciDyjA8qrpU2b83XAcRJiRjWgE6O0y+KO4GF1/tATj+LJ5I
mRnmDvO+UG1MnewtQiieQGwEuv11Xd8ZoDXJ0O7K8tUweTuUOoquTpd91pbyDSSxB4Z9UJyMa/l+
pwrP5F5d1H+VoYLRzCZwA3oDIbJJp3z6NfGGC2S+t/bzpOc9rdKj8zN3CQVK1t+HE1s9gSOhwGaM
aqjLvZfjP3BGAEk02+mmN5IBVaVxDFw9kGohS8j/Cid12EL55wztX4MdJZEKZ8iPhqv0NgaM8vH4
LITh1p3N4kKfDARpW305plf2fnAtxvf4T3uxwEtUZRCvf1pqkiapGctmnJ1HDC2mCpkcbogBCaZr
HpZF0YiU840S4irW/cAOeeyx4AD9G1LwiapKFMIu1kLW9zgdsQAqlZFiD8uY/ykRxXoVsxvnkNY/
7sCodBSxL63HwzEYR575kYdwLAs/ZNtzxrDXYsj0/CMGKVfznjdR9Vrd56Z2yKACvP81V3B+cHjn
j04+Kf9LVql0LDYuf76XOQIUTPJRq3zf/ut9EFMFSpls1x13tlUep+P2jE6lsahVMutYUirWeT40
cgaBD0MXGpCIv0yGWlWqzTqvuomAbDwfiNzwXGAZjTsP74Qv89RCKKJa48SxfkZagOMD+yp79oIo
8v6rbqdxA3UQ0VTlK1AMXfof2h/e3ltEP8uA26AshnInc8RaERidmOW+0iPitywtwTpEDlNAciJE
2gTGKAIg1USZ+O+lLAnIPMlqArX8fw8qgM0jJy0W2URglIXWL2ytv85v7WSjPtHWsHSEEZW8j8dr
+lw47HgcxtIrjUDZzYSVK95CwL7Y+5Wo1XvrFfvhREcuF++wvBaxLTNmCcTI14WffFrQJWNG25Tf
cUlgWQ4TPkVPVK9SAnHjulEJo/K+PYfxP07XwtCLCQCukKs8cxrDyBTplsz2eenlMOB8dQ5zjkcf
Prt4MYJQsTmhdbotpaez1KpL8UhIGi5a2XSioh8bqHF2Odhe32UTsT09ftutprAG+b0MdsOUx1XK
h8r7s7bJ69zxUZXyk3+MCrhxTyZnZEPr4CFUGgwfkq+SCrcistT8EEcfBIzAjii4umkRPy2+OeOE
4CyrS5CjCeKlb3OQwMhSUjTcVDSJdlbtzTknvVhSoJ293odJYwJbnaThN8ykCYozPpB1boHcwtbG
1za2LOEi7c0DtyoejLc7J4HLxohLM/oRLxJ9dV4To2OCRrSM3h7qjyLwTw6YDWy9HjTP2L0aBgUz
UJkbw0jehQ7oRx4e+wq83MBmoO1MoQAZof+BOoXnWA14kdMYYUqymHevBekN4tI/7+cwP4/RJtP9
6cun5qn2yBJWwOLKAqHWdwB/aRCYHlkizLSDsafzHPOqXom/Mq+lhHdsjfftSxi/sfc6KGTT0s70
H4MyO3dL8wgQQgwyW81w+0kv44rZNTGsqpyVoEzI+fI8UKSPG+JMXhQLerGcYosZhdGx9LvK7slW
0cuzl9shUsqxnEBy2ztiNIhbLS04MmqG8EqBbsTpR3vuH7eKOmS0JbqnPLkHp+R/ZBHgwjARxE8w
k6Qh47vUC3EVYSct5W6dS33JdmEo1FUhxPx2BfO35Lh2cTsMf7L78pdSM1z2meIr+cIK36hNficB
A6UEX8EUmiqczXxW6aTvamWCnaPdETO+Dr97xjmA0EZQi9SnYkB+IFr1fBNdo1skkc8BVHoEamkJ
jtXjVv3/8bovtXbymNmnBwMeNy7hOY8BTbPW01QDMmQmEXp6ILI+9rJfkE7lBYqYgjR60Q7aiSRQ
ge+QQwPGVzmnd5se9BgsGrS7QZ2PeKdNflWc8tsUXvHeZSHIcQqYSY3BHgVaX+R3qsbiUN6Zrsbu
JXyEMvKHZBQsT9ORVbWhsxJfQKH1qF0RiBwTSX/wuPfTeNLpXhy7kuSk4lHZ+buRTAoiNK0rJCYn
M+N0AkomoIsuvDYU+d/3mC9pM8KD68ikdL8JvqcmHsWy+6B5OIbHW48tVA2VmcxyDCZQNtPF5ppY
cqhHNmxXb/x7EvjyHkbZgTpDdYPRBKKac3+791WXpu0gCN4OdVdOntBgGyNwZ2058awFLLmGq0GX
kyv39k3eRumgG5+Mi8DbFvm0Fz1Kt+QMj9Xna9e3cO/nokYRmnLKvC6907oJELHqOHM3XoLZeGfg
+htGMAjcVpCgYOJjUPGuUy+xqaz1y2vI8azrvnIcINVvhrSHy5qSeUe0afzv4iRj5LXWTNLkQ4lu
TILlwPO/qa8NWfseCaXVUaksuAIluO/zZJ7+LL8okK1Fj97WCgElZce5kSgxys7JInDBCUrTdN08
53x2nTABQuN2eGOYRX/9dSjUdcHhuRbdrEhabBMy+ZUmDV+xSjhdfcr6Kc1TqcP6MbMJV7MOcgSb
68rmmML5FlGqKO14Pu5X6YxVndtHJyBQVCt9G+XL5dQGtMlBJIuifUAgb0HyEg0rKOfj3ehkAUWP
pOjRHiJnwgCO7dyTgAyBQrP//WuOqepb9jrKOsseU2QNcUeaJJ9uC28ayaK5JqFk5uCjtf0oTLyk
gWg23yysILk7ex2p6nsNZjrzfRel7cezManeIBYgFUByorW09y/eEaoxGeuwj89A9P7bgNnkjggH
EzahA9StI7Ri2IVc7NUMWvUodpEKUMRF+qA2PH77lfBXeCecVXZohvJSkgF9iwZ2zLQaaO6HdAHy
p5xCjnwCEWcu2qsy4Hl3gueQo5jjcXAKfyCHAXCDVE8te1w2jExDw/vZnzuT4C4PuHggK3fVwwBY
bP6coE/tKLRgk/r/uiMMwnhCy467S6BSCA2btLQ5UM+RW7lWakLLMmvwo6551KQA7xqhkIFCG+Js
ZoBBZIFeycGPL+GRbCuA1Pgiv7+gkAQDE8xHwfMjSGJQ/iVfSdad8IfnFcowSHzbe/4RhVKGB8Fr
HX9ULeSvlt243J/KYPmBnqrIDS1VyolHmScrl/4AN+bkK6iW1HwOiVVQvzXC0dWGWWCwxYtXZ0UN
zReWJNEexgwtHuQ1Uwh0t/cRqXxUf4YZTCHgMDA+bgNp311OYLqXi3Ogu3c48xTrvakww/izMW9q
FZvtEFTByNn7MlUM5tSsZvoSjxLf4eQkQ1Fe3dIntGRwcvMn4SqjDv20nFY3mB+/GapvTsxUNU56
NGWKr1FQtMcaRtNORK6LES05UNS3fau6ICg0V8I6ZYohJWCDa5hqtJm0DMhOkrAzblc204ZPYPbF
1xTLV/et8ZybNThudwyqZZ9DLeenw4QJE2VNg3bJhePrHtiIFEef70LpY1R0LQtjtwrx+1SkTuvK
N7mPvqEsqIwpSloXm120UA8BO4LQ04xRCmV6OY0XvhqC8tR4s1s0FmbJSOR7QOJSJEqDVsgqv9uk
PnHI9xEAxBkmAbnKmEQl+qP8ixyH2Kgf6ImivGNoJLIRrxXDhVsR7QG8yWn2F9BSax2P1DXvMrYL
paq7mMxCaFt/uqFMA0w8wyR8lpKQ/oaQAgT72qvnJ6F1QD6488aqx4bKLWwx3QfU//Ugp9NkeCMb
ZQUPxzbdM75ovPUoytZLYjtu7QV+Su+jVS7zHeHf1qcPy8aZu8yoWg4WHz4W4HxFIl5pl9TFtR0r
sheD8LJk2qH5yMn4jBTq/vnC87urXkPwd2F6cWQGRXPImgVvSMgsfZEFe+t+zLHgeHAJSBXGp0xC
PDKFXY4wllRXsvSjF+cCaNWLMYQ7a8kxtLi6FTcLLkDkz/Ip1PjF15fkp3+gyrabWBWy4dgllx7W
eMRTegqPftTquI7aU2+UHmdgjBJ4mcM8ki88yoGCgwkPXUAyDUAjWjXtWoq2zoOuTCP5yuo2Q+Eh
xIb3/5lOTKewQdNPuqCSi/291Mgelx0hicKpZi4Qy87IK4WgA/PIVOpsfuWZvOhmjoZQ6dT+Vzbb
heBdwCQYARJYeXQaTqnB/ARS2kLrOwx7Pr3374wCOmgotPjzyW+qCJ/HZCxWn+XDnVeqhGBV6NO7
t8HH1o46sC/xswKAsdlmi2zirf54A0/8eVIWsUAJxC+MXUlcy0pnS5UFNce3B6NF/TZMRWsJEwuV
1NdbN15RDzJJWIcDZyRJVMX1Oh/2NF2QOhmhEU0WZBGuyGuAUMeO4Fp8WVKsVwCuug/15JDpiWva
dlNDg0YLJpMAAOQLdyQbPw0+ep9X9BBglZZVgxu/CHJIfJfHbJWntovXbZt/hValnZgryYD0S0bc
kBeySb+lx00GocgIjzGjOeOl2CWNZzKJl7EU58ftokh5rJFeXmb9pisgOIXjkLs41XiJng5DkCfN
62MjPz2tOOk8db4iutoRQOArQy8GEvAZSR9QMxGv+ZQmF+iNsgSL7tGWDFjrX4l7G3KHlCD38/tR
G4FTKJjEUFjX2pTR7SgRKdRVc5GlXL6TACEHBvwLUvDawDTK3qty8n5yoLvkF3mfWEinEcpnsag6
lHFmuZvhXjTL4wcacEFX2ekghPRGShYhWticdvLe8t2dXUeP6RVwHSm+Ywy44PDeFwTmmRxc0A1z
aHkfUhMbXEFuxjTd433P0yZnQtM/o74C9w9mgGZpcRlp/IiG2A0/HHwqnZli11CImnvA+Ud3Bf10
TQy7xX8NZNBBDhWEPeX2ehDcskeG5FuLzOnGbs8hePOUwygonHlY6TMoQYhvOrNEPkMzSq/HlVQ0
+KCsBwuTIaRcyH5VycJR1fxk8RfXp4qPanYeg/OIGqp2ex71pFVO324Lw9tzRKLpPwiNi6cwTgBn
cWxoAPzj61Tv7rQAAtVqTFbJAj18xAjJQSFu2boDR67gqbCbUxafG4gTs9BokbB82Fr0hNCrVNUT
MhpDXKkojTI4EFlGv+7i8pNIVnmsufFYNYOdPcLzeaNLhYC6QlFDauTw7WFGg/nnJle8S381saOz
FOoLeDBEBfTIg20njrcNtDD1lDQcOf37K6+yZT7Zg5x/6DlvY8LtIklKb+E6Dl8AJYYuA7AuDWv1
EDgRxrjr2C2q+ijzFsnunrIPV3gghxahrWI6QATzKDx2r6bUxVkiTVAC+3zNVyX8F6BjTjAyrfBX
mHtbKf1Rb9UH/slKDmtch8igSaaQMrWl7I6wQKeSzZiKElCPrZJSphbJpcCl+N7qi2ljv/rDSCAE
DMaDR/9Zp1kPj5MfFC13OuJkvlc7qG4hiYiyfyYV9jZgiekimI8a9kB99h41JmXuwJKg3F2btcbM
x70L3mW+c5NZ12PQ9Y1BVmC7NbrRnBjeLP1TRVnh0lNM9UJROh0zV7el9moS4iYAKZd++rUG+4Pv
/Mpe9fF9z82qOUqhWFEUT3SAYqs9dmN1RoPBx0+1BS+aw2je+BIhmLsI5cdD5RGKpOTpby5+gR/J
TZvWTePwKHWMfM4cdruYZL0NUmX4/jtVbsMVbUhgOE//3VfRRewlHjFIDlosGSb3pL+71vODTzAy
j8kvzZEsOOocf3M72ME59sGxzbC3XcM5QNEto1IMMzZxtCQh23Nu7UHNceJ9B2Su7M0Tn2VFBj6K
bsUZgbkAIHBtHhPGV9OnaPBUzXp0dfqj8hL11GWMW3I0AmLshOr+U13kRjREjI8dhDDrWtePQJtO
ecRnKfemJAQDL3+Hj3ZrR6WxUuormGCdy1HgtDXJ4+gJ6utsYncNIpLecyBR4xtxTkxvt1oRhvis
ffUUaeDasYypEBlwU/uVpbOvMmfIuv4JoO88RZBnzT28Y1wyxNSC5FH9tOItZXpAAXlPtXUExQDe
+f/DdGVtyWHHiiOyvHtZJRmZyMAl0f9RJ8WbWunJp2ufy1oyzI8p/mUlOf6akK1NNUnaq69iyQeT
iJlrn3LzlNX5RuhC05gFpIr2uVkn6eYqabLdaUwnx4ffXfc60ZbzvnFZ6PVvHG91ypS8FuRK2rcw
smPzXokFEYFmSA+Vv2CiFxGR4eNYqYTJWEbgAKVS07UcwjyCZOpBtd9URMSqYnq2Vn5oYtNDHlNf
w4h+pMMY4hiWg/7MOJ+5nby0wPBqqiCe1HywE6JY5DqKx5TNoloZJlU+vi7u7GwhwvEzUWyHtAbU
XezhGMptzf9fN/V95eqMzTIbFrAtfGZ2kdiuipuICjBQNW+SYZkK+s1Q0YVn4LaNCrC9W85XsUq5
LgTXSMVF+WV1NjIz8iVKd2PfmFpfeLeRIjLnfdTtFOT8u2H+XSkKMouKsBRq0ZCpimQmM3xy8K5n
XnsOd1cWAUy9ibjhFk2s/nGrjrL7oLo4TcJ/L0BsOHyfT+n4k567jh8EcsR0vi0Hi2RybrWSqpQy
YoVhq3YDdQh+wTlcKwfDijHuMeEAZv4EpHS9APqoIlDtzUNsVJ1C6GacAzSSdQfJh3SGblDaYi1i
cAgJdvyawTPGOS9tVeOpTziFdA5TMICBQf5pFGaG2vbCAnDXBb/pQw7GDhnrN/rxR4/ATzblQzlR
3iKmG5z+AurFGfrQRi1xRr+fJ+ZNRpNeWNp7ML53lEfGbwn9kzARDnEygDKnan/s+SBWYOBRB+v0
GdpF8ZXUdAWSBBxrD3kagcEJ4DPQ1QEu3eomEripO54RJYHQstZPSEzDfBtj3+i/686Ccouj9S4a
s7SQZX+f074Ciy1cj2aXE1UygaCe21QdCg4UGu9mqv1exb4MnYVW088S/M8zJw2VUA5j5nZx5Jbt
4hx1vlXTq3HahouvQ+Ux1yxi3ELxqcM3bPUTpbOWe3FOYIWfDjFHFYnre/Eg0Dhx9glTIBLkwC1H
Aby+Izh1Vk/nFsV4+gaWBL6Ujc6W83ZryusR/Krhn2jF7FGgXXaBCjzcMxu+KtesMweKSOO5MgeO
PXX4e6/KDqWN2Gg2jjHdi9R+380C2O3tShWUFGjB0EKFb54B6UB+ohyd1d2z3SBTLY5wYl5NEO0I
UpCan55qRHCt6WcBc4KP1/K7eUhHM8A9PLoOpHqbKDL8FMlrn+mdhYZOTnU2EfLqOzZE5YtOkn/X
Kpar2GFjwiM5PbGlqcP3i8hubDOh5h6C61ZJ13rN1f8jT/SK/dK7S2H8yh0rFFDBYFR1KRs9Dcgv
PfbCtBApCQI708hj7/y42/sW8FSUjOcnnYKjiQG52IpRN3PwTkF+XGaJ3zGqxrAsuh/bKqRn/ohr
FYQCqMnanhzx/l7rmEixwBxgzgdcRE2cfFiM+Vrgz0XqVLbDnaBJpP3Ns8f/cLfa1amVvYpGLrWm
RTp2xt02P7uPnW5lVVRJHBPz7vQgpDQFD+GVjp7E3Px2IulVGZCBdOMFgf+go1LTjY+/gHf12EGE
NQubDcj5TDClFavcODZsdE04+tSRQJOyXKEicjGSwjFc8u5SnTqWeum1mJA7ykn10eNBaqH0j7Y1
/pf5gIV8B6e9sO38VvZNonvhZQFtofeKK2ZHKxGa4OGP6SVcx/0zlsFrhb2JnPYWSnYBagx7vNbA
d0vAheipLe6pUDhMUY7UnmMLG1TWXs2+Hp0/xJ5hH4OeHwtUBMy0e+fUrYA6J7zNrfVzQH4YWfcE
AjZ1rdlJblHets0ioV4AQWriu0IG86grQE/a7Ccun9CPqvg8aehs8pIWUIDDyBszlXmELJHiHdrA
jHQlXtjtvqoDfECqqZ3+idIjNpscrotF5iyNH3QiI/XRofQzyIYP9y/dkH9v0cS3K2NNvybU+xF5
C8b3XkY0NmdRU0z3lD4Qrq3dzv6aipkCt0xTAs5H8ConacHvHGKgtMF73FUCU7xzsV6d6DAvX244
hD4llamXqOJ48brplUWTvrONtonnijDq4iHLygifacmbggcOtLg11hUFK1RMgpZjSRdwZR9uc4+9
CQuUTeYSM73k5U+fYmnzOVZb3f7iVGvwfdfue27Bofe023LU+d/xaPkmcDmsEuC/+FX+/437a0pR
ZTI0j9N+3cGnwxpg9kV1V14CX82dBuDEpBXKHYQYujLmcmICC+ParepvPiNrWTk30ckYnhNqpL9O
2uWuyae3pKIjiExP/JXca5SQOhucx0egF6Mgu2jQTY0NKIm7Ov8eXXjmUMBajIgQpZ4Ae8XG0vd0
czVHG71T+GY+vU5/Pn6RebeZjK4Nz6EFL2yiHKayuldh9+TXtioxiHz8yJplA1gJe3sug+jddCY5
ZiJOm64DUs28s9GDVjM+UrYyntlEpKfPDXRUR9BXCUiMoSkVNh4kcwCpchfsZ2Zf7z6pM5Q5ZpsA
JVq5PYh5aX1GdcZSYIbkY81KdQ3PsGm/euscqa4kBD+XTk+8ZJtq4JSSEV221jpE94pAe2PrZH+0
5FyfIxX8PZpyVrcMAk5PgPon4Z2n9D5jLoxvswGHvPlFo3cjlI0dtFM4e5oMeFMqFQf1zGxGJlMs
SMY0FC/r6HHkAmDxG105k7x9VeW4+khZNeXvoqHmrZxlJxLxw9s8tJNZt6NzZL4bDfc4mxPQ7P/1
LggNwa8hIvUtn46+7XeKuTGzU0OJeUi/H9Ce+0xhpt4BqQyRR6Jht1mWWh+wjAP1Q+n6j8OUP52Z
WzjqIoBwWV9XhnxinbeY8BlrpuafBgX9nWulQDs9BNCLJTyb9pY5CsU06KTAJSiG7t4L9jd+6YAT
uztJRPwZ4PKdxx5TQegYbdUMAIoODYiT9SJlnq5+graUCirL1PL4A/u9ob3UPipV9GBFagXIAKqA
zTDwskEHqpIelubKmqQmg5zMnNi60OJvIXVnBZr/CYdljAhh9dZiHmiJHSCkCi91DGN1mahfhngT
BLWP5NiMGqegXxY8MrIFnsuBeqjAYr/1uuwk/5nWAyN+jjBEGZzq2PnfM4FbiFpz+rF6/dXpQbmE
SXLJcIGN9JemIMLm8E4oH1tmLSiwDwcHgTTGnkl/xCVMZSnS4CUsDT7J9LlDw+6GBTUariZ/tIAf
Qr2054/S2ajatwMiOFXoX8Wq51sgHj4YqFE+q8fxWJvbODmUbpR9qbO5rWNUOGPdMV/yEs0ysYy5
DzbWK/PRbW2xXA8uSsDuQDDJB4qkyObatrNJVOoAHS847q3Wj71iD6bPQS0ZB9gRJN0Dp9zltTNM
YbwyTLosedGAnjur1ElWlyed3EJlBbHsbHAT1lxFgLDrXCHPmit1RbrUrtMIzDQL1IsWGeva3X12
r/C77v44IH8Fmh5fDsEbfkFu/SXxR4++uBiz0QoD8V3K5GCcmhWYZdcha6k6DlcrfVAFhPk055pV
W+3K01+e6NZwVX8z9rJQ53J6DgI32uDkIxFed4RPS0407UgvalnIROBqTuBnJryWKlb3pY956vin
zCR1f+GV/EVlp3Y7AwcPTf/mO2RPpXIXBGbDYYYN44+BPyJuHDl6VtA9OPAPzWA+0XIG4upmekWE
Ed0MA6Xp7W5hlO8WEdV601/+XTq3ZoTRvB8d3x+5jR303qbkMS2xszk5/AC0WKc6JsGKWQl+vB28
ggZs0wWQgz3NAPAdwd8KXlIZVneyy9Ssiz/zbQqVi6E7x4VKNuu0o5swug7gMPGgpULspZ3zSUX3
cq8rmIptfDPG9GeELxjiHUAfm8P5w1MK7QntApvkYbFpAyYNFY3cfNT8p8zUHi8JYAh9KzgPvk5C
9H955otdgNcRA1tdGy7Zz/WgA+/QOhym89ZBmuoaU9RiRtYLt1y3gzv2YcGw/ntZNQ3db5TUGBMP
b0lh0ygrQV/Xfud69q2s1dZwQrQbgn4cDw2dW2pm2o+iUjFDLC0bBHgWCpkqnDWV7rG5aq37gF95
tWZO3LQE2oNruinGUCjUh476FjCj7ZkJkUhLPX1welrK6t+RfoHPdfUnxd7xXLVeq8r6uR0oUOIV
MG4+ybL+xL7/mBZFJwGcHfR99o+dNDSVk8utPlC/7LWyInKv9e958MhiSQJCSG55gyZpujsfa5vH
V0TtXBrsPpnhRuphYbLp7ne5nb7x5BlgHkvFKvao9yhMHKJK8gIeSaz9MtYg2wjtzDOIpjhjo/bJ
iMRDMziEPuQI7NHzpuwD1Kz3SYOaJG1Wv1pTnGonuS2TyVKkvBW2atY43kH51/yacLTL2wel1rO5
Efwhs9HnrMAkIH1vbI8zVb2j6Wu+Ss1+2QGL8JhBWwBF2AzadGOol7nC75QaGAVRPQNLLy4rl2gf
G4oqlJHEOHt1BUTEALho/SiPjRSY1wlO4Gaahcsgkdf/YtuKt6X366n49u/zr4jTgbZ5jSp9DUah
rwbV/iHaT/KoYG6Ptt5LpYcyv+eTV1WqiJRKMoWQ26xm1KabKHsjC0/fvNojbwEr3ZGL6aslbOQK
YRBnj3XHX8de2cXmrMUwlGvZh0ivGWx8TgmAbNNA3A6SEdamut0GqkJd37nWcBWOg6rxd9E/DzA9
RxQf1FQJp4cHVrI1IiAJtvtD7ffd7oUUTwmsSbSfmxWP4rkA11Z5kzcliGfX2pVpEeK92sQ371Nx
LoFphtkYzSPSCgpivyp+ta6ciiuICnmb5bL29G5ah+f4xoco5W+89jt874hikVd91cSnHfZyql3o
blsiilMSYzOXlVEXVWE3vws0McIzKzz/tHXUnTWaHBFm+MCcI2BBD6T2fWqs20MdCKQQdEYHkb8L
LqBaqIAODH7sBzTRLW0SBIWDCUui012RZ6eEM0Xk5wLuLoyre+/CzdKMy/r8Mm+SeXe2q68DzSX4
qiJXRawlK3r1CrHU3jy6W9oFPOY0yfVKNj5nIzLZdz0XCNEdHyHn0MWua1kXbxkX6v6Fxh4st6SV
Er2PNJ46Zx245D7Zrf/dzv3xGs9pU+ouork2J30Tq2LnQ0W5CvWykZbRCh8dgF7IK1RJbTqfojTX
iAHgoM1ezmgLeTdkphCBxGzSathzoM+HdX7XpxKRLPwjvQhdAxdCPzRRJ51Zd77QLADJk4s22k3V
uQcrWpT8pAEq7EUlK+UbMuVaks+S4lRJeRLKpPJyJlwBob7tFAlkkyzaWLxZAy3pNqoyWWk2Wo9m
qhrrNKSX4Rcc00zcrXQiYRMT6H3S9k7leEEJl05ef6dg5AGnnyXumgP/4Y+5TFrlE1sB8Hqeoug4
8+jL+hCxst3lLXuhSNrCFkqYeizsHT34vBxeVnbKBegb1h46v+SgrfjJpOTxpQLEZoSJiomiOwQq
kTCHFPQA6AgLtjDJgksXwPd86l+gKdMDDj3CaiOYvK5X2awC/UPdnlXLOGcR8aUH3t5lvzZsj+rF
VtZD9oaF/wq0KbfO+68y6atXQegvw/sqwwLkyLzRFJL0q3T7etgaeO0mByFnXCsEzYHSCtB8sv6d
vNyBquUNdFkraxN+5eTKv1eJPGjpHMXb/DkA10YlqRG7TJEweDVs+n1KoyREU99wf/MrEd/mbivc
GyQjTUMByln+TNqHdWCn9Ts5VPehel6HbydykM60D6/ervzO5e27ykjbXYXWyvzyOGcIqsGn51uq
tmlmy7M5kF1vV4GU/Ed+T8Q6NQGeyHRFbVFmi2gqMS3XV03U2No+vW4owGsN6Dxi4RCDzvGHR/2H
QTAWsA/33OspBjVlFwlwezRkE2ub6EmNIsr4wf1DyGn+ROxTP4g17JeRgrdN7GErAwYv65bsEu41
w2OV0K6eq2EZDBbfiZinTfcsS/xZnOW5KAJPqkM7ctmA5GA4uBtANfJ7QwHmCfb2XD3+b0tCFgmK
e1eJLN6iSnZIrtQk2siBCi+nWhedvh5Obqs6PSFWYVCbNWABG9N4znVTU2YLF77SL7NzbRopq0gv
QqoNbj0eO5CwnyQ82kx+4NbzZ8Twf8/fzy4s9ve8pkAWAiqQWQQh9lne7vjy4pl3d7ohZ77VWeeF
TLYuh54uQ1lHU6jDCxgMJLf9pvnJbaHq/1aol0phdxo2STnVJaCFnShuxQQtIo9Ql9P72VHwyZuq
fsyTRA0S+sljtqzYjz74jALCBTMxiGUlu5AziUWcygA+ZlSzyGip/drm0VmFncYclyYUadfwIYiU
1/e4JuDRZ9yJQEyLLyXgGCTT2r8hPcTFxDwnMA1vuvazLLenqprWyasnMSR6n/j8xLws8H7mplmE
XWK/fopY1n8/taNo7PO5w0l+k6GJBpLDKmfuYM6znBpPtIc1rMAHDxLQl8dEwFpYOius+j7HXiNh
CEE3uhesrEiZ64IsbdYVoPSoILSWvfwAUovkBlGHm1wmLp5plweqBoe7ehl8/wnrIk+FKJcRm1jP
8ZWndentbT8/v5/ryxbpM8HTMP/GMrR6YJcv//gaGv5bzaMn1+NLNs1HCwYxyRXamilUiK38yqVP
Q0YNsBno6DbQiLKVVZZ0PAbePzm3OVKef/T8dCKTiEYJ9nXaPhvECX8Ed5ftp/3HzjkbIpF52ln0
1LWliWRl+mFS7abIfgyJR7cIvaI+3b1AUi5UOpBdoLtV6uGQojUEPPG4Nxandx3YjrosoSD1gbeB
3yporHGfCOhVt2eGqZFdoSUq9zDUXHaZ1JW7vCxprXU9a4oWppXy6GL/jVwDEtBPUg24il0Fhp/1
o7g0UgUCGaNzENlPO5KfbwXq6wDySfS7VqBSo92qgrRQcrsrO3YL1QpLFEA27gZDOmrFTCSKFo5Q
xavg4Bwk2BRbqKda2T7iIko7cm9SrId0nz6Y2j+ZDV3TWbzUcIm8XApBTxjFO6IaYWqj5/z/q6+y
PrRh0ZG5vL+p+jRA7KNh3J7S4YyhBMUWdbS3RW0tYI6GHCdb9fs2UaRYBZdoIOe/FUxu6RCk0ZhF
IqyUbhImMYPKJYuroLTBPW3hlLsHQfcmxK+me5VngHN0aMqh01woX8+un1tfxh0qFYCKItuKGDA7
JG9KvpGlGEXNSqYfb5/abSnv70Iw1Q0F92vhq9+3mExDz63OVurV1MLVp/wgCVcFBCZIHvr1rP1e
sQa3xnfClmFsD3oX07Okf/+bXhbqILXF7B4hQxMBwBLlqyIn94xltfC1wAeR/gEZOK78Anja9mLS
iMQVmOiPeT3oKNYkIkA5GO23Q6ol94fJ4/n809GKX3h8xOkuyWWG8sS87vrx2mk2me7F7/TGZjrz
OI2ZKP9807kNBiCZmT3cuqI3BgD3jjHKiYd95IAGU4xY2TI98P9xBcr6OmQ8xz3gdSc2mQqb1gNX
BIwJfuzXernsxZSI9RiEBaAFV7rLK9MyrHemxMv6VoGcowdjbCTsyVBITCzPHmfqEQQqrhHd1pnq
f2Ziqe/Uv+u6b6z7XD1IldzLBF9YfElMta/IMY+GzKBbUIIs5gn0C4MBs2ldH3iFuOamTTnh+QfU
9SrWYID8DzNP7HVXlYqYwEWZjvi3SAJ688vWWp1BEvpH14tsZm/jsNz7BHUeQ54a1x2l1sjdi8wl
X7V1SBGoS6ol4xIxeJKelJp5SOW5IJXCcjhzLy7jdXLd/NbVVxPXd5LBhJR4F8FegpE7RVIGB5BN
/olbJoptcomQlnXX5GroX83xqKMZNGJUu1yZHSivWyY7Q80MpnWpXFNKee6oNInWvXP7DnDQ0T+E
eo2tLbUnhaXSFEENjFAGWp7XCvQ4Ztd/ZmK4dQsBbuQ/WYzgwWwWX7LUj9pmT8Re9E5xkcmpPVLU
68qkPeuDpl8o2tYCF1PJNwEGPS2hORRqBJTsfZrai6/gSHDll9GrSuz0BTkKCIbcMquNbAhirIGJ
IMzm+b7iwzKmbDOxd6W9lpx0shM/+EyLIbmG88C7KGTDAa2edbBHRWuvs/02tJDeiGe4ahNWWmwL
UDg6civThitCtcJFfebuoaMRW2aVwtIpNG+sznIZsUj3n5uJvUJEQRQ0Up+NvyvL/UI/8UxZwfrS
LY7OKKHtWj0xGsUMKSURii8d3iGIV7+NHj++X6auy6arsnD4TTSlKvAWqjY8jU+JIlm8UquBPw/d
9+CxPKcwYh1SeLibfJCrszd8+vF/6e1FR/idCvmGqAXV4y9uMI1yJPEw3y8KGiOI8KlmpB4kwrKr
gUTWhbNT1t6PMc39WEaH+ZsMZMyLERdR3TjdvwTpqu4ut4JLkEnr6trQL4HzrI+keOmywOxMPw3G
MlJ1QJDVhZ/pM7cfa+ndLiyNveJsM1BSD8ElxNiwJWd5MIg0PGrvX66WNPN8cHQsYTB3V0peV21W
A+e39HDeXcW/ps9IpVF26Lwhbg4z/Fzo0FshclSIDVZNPlwU+C+hrybB8GONk73s+wCgBrv63Dw5
21pS2od9ZjrkK7o0Rz+dM6kwZ0mzy0dBZYi/RQfmCUDzVe8/Du4Fslu7Puf7ahILlNQo/um2Wef7
4EDtng2P8kmrIAAqHNrcDUg2ijSDs9tMu5mo/d+PnKmAvOUQkAu8rE/XiQsNuUjGvAAQQktk6rhL
XI8lw0OVgiWg5DCUTrlZLbCTGaGIgNdMn7M/uDL+HpRJxtoAguDwXPXRmmsNQYG3ALquTnmEO8Yz
9UbSRMm2+sszuZo3IBJbf120Nehw24lQQPW1bvO3h/1ITdWqTmbmTD4rtgmAR4T5KHYTpevpx9Zf
7nZbfAC9TTZWPFnSfKr9gqD9W7U+bUgEwTdd9GwrVR214cP9H0ZEr0l0csvAsJydC1NtPfXzyc0K
9YSdtq4xQ6pV4EEev3KxwbWtN+L9Sl8/rmQjzbJoyCjz/TmCVoAgmaK5aHDQMCDQz03cKv/rlny+
K6zzJaxbsgG6CcNOI2XGhoxRug09nBS6JHBgOnriYw2jKHR9/lv18d9N7cp/N/KZRyOch58Uuxm5
7anKAgWNCLy57Om77aQ0rlMu1Bf80NllfwTgHRGPG8E4zNt6xB4u+GSOXWxMW0trZDu3WiwuEjFw
mJSb/HwnI2nuc1epaNVmslnDupgzV5X3zy0q7Dlv0F7JPFOaJhqN5u54HhHaT6NtXn/VIcp/8H+H
csmlkuzdtAqN6OlKe4EeOEUD0q5/WwxRQJaI8XgTtTuxtl/+Defz+CX59nT1T74AanR4KHfba/35
NEA+CXz11PEfE0nGuEtnV6POEmvhuhanfP9MVpZbyYBjTAI+LLU/wyFt3C7tQ/53rE9W/pYaK7on
oWXEyAod4tcf0XPcfX3v2pr3p7n/o202IgWYhX86wh7KBLo7lqNMosJ1Dzv8ptJwa9E11N/6+OJI
4zhQxyyPgrcKk7b49kfKKRVT7MLD8+62cNwaLfmGmb1bPjY6Sw8wvrxPgTGNvAdxBzz+AJnsspTm
LZGVKwaFG+EMl9tKE+/3Q45YUZZU4jNPd9LssCjKWLsFHFPHtJDDHf7iVUMha+iPGWDKVLoHdZ0F
K/QZRV/1f2r8d40IL7oD1GkHqqVRjd9pcsDiGNCADnhIos/vGMUH9ZLwR0GSNxi3HYNFIcrYOQua
4n4erDG7FxzE1a7+biuZdMd+AylceCuYExzPsCG0aalb0egtQsTCvmyf2NkWYnPeB8RBwV7VZCJC
22BYyTsI0KR7nzpS6OXGWSRh1G0p9GG3Q5vZwrxeyBvs8syiqA7HO4kN9JyBoB2NniUYIzPfDeEj
rHPMisoKrJd5HPlCEGf7cMIRk1D+AnLmEywFiBCt/wvCjhH+e/UhtDUZz37N/ZM0o69GKsFVWaiq
XhCWMSfQqWAmae6ZcvCnLKUs9JYV0dwcn2a22nWXaoL4VaksaAnxXjeL9xsgS1dD+iLOOLKtDeYa
HzQwiBj+ifWZM/5biJgkjjo56RPXnxE+ytkh6D6jKpZfLyLSyZCbJnfQYTBoG/3DpW1k2T0BqS+q
SO2xr2j6E5WyecqdJUiQBPbFIssQr08lOfEZ9XoDF959sY7bybuEk2qwZPn6mxqcWEcCXar1BOST
AzvHTyAK8Z/qOvS9NZwiV/cE+Zjjbid1iKZRljCZn5QyuJLLXDgPxPgPz3o/amsoC/xc55obqnZ6
iln0XtMlJ5lsGJGRXQIZbk2u/ia2jJgYxWI3JbM9GBoEgcjg1jCt+4QBSMFoFutt7VoSFIKJklDL
z0OCE8rGFz+WpcmwYI0jsABOe9comA86y0/aFzeMaaQaXhS5DtBP6e28BS1CieDE7LQRZ8UvmOGw
4WoPrqCy9OczQGzZJsWfQyFGRIYNlU4CObWLfbuPKtUIQLCtiF6l9E9mnz+DZvIKfvIV+kn6LaU+
hhLUj+W+D40rXr6y2cNk3kThh29wxU08Q9iPqv7MeZU3uAboRbZHDCq1t3LPps5mXtfEoPie455d
sYDwcE6dHJJK8hbBkEl0hmAiKzBvnytYL/hV4+BliuG/FmV98Ee8/FXbvHGxzu1XZHFvil6B94Ch
WhmItkbFP3S04e8TFw/2T2OE85sic222sh4Gh0gVzkMsnqehZjz4CN3MnNAGJiGNU+SQL/5wOct8
jE8rAVR9SifNs5woTX7mwLMhS4GCn4UCAs9ZriDMC6DMkttTTOYyDZWCxzIyX/EAdcpNoFZ/X8JF
//yeMTrtxjpqe7PFhsiWecg43XvAxO0ALh1R5/p7Epaw2MJW1QmZ7UGxmbY/lVgrCCCRuT+soXFr
VWl7mqBXcuuAGoc7j/7QmhjfYZfBv2i0dxmZ7KjAv5w8PCpUHPj9ZEMwHGK8UIk16IMZ8sUOS7qi
FSbvPVj6i/rzNtakIuCmYLJKhtf7y2sFdwwY4TaIsA3uBeFKdi5CqVakDd6DHLR+LCXKZCUhc9+Q
WJtx7Ed71YPEzeHt6y92j6ao16BIXAzWUlNq/F9RN8VGOqicIp0MsXWKQob7/B8s8cgde1dbRHgi
+LohqJ5uaRbpJqvi8fSQPgPJmOPdNDW8RzZTxr3W++esmrvgN0RN7/hHKQn0ehVXx6bfvfLXzdBg
P9+xRDJzgNQthmLQZ3zMSofiMCHAYYzgl2/JXztJsf1FWsHgcQUPJwJlv9a6mK7w8FFAz6jQ/Ush
4mzYq0D/8/EyzSXFB/3hdZCV6etlZMlGDwnO5QSHysu525mLB5MQMX6esNx5FGF9D3AEi4AWeMF3
obgqU0PQb3YjfdDtNVgKP0RqQo8TVme2jKmNwOa3Qgccti/zAoaiX72YNj0xiAx9fPRvYWWHqthV
osunX7u3zzth5zc9PWb6ROkNVB9+lWXeaT0KmBJhNoEcZJYbD5lYJAGf84/sMg96VB4ZurVyhW+Z
9jc4tzhsKFH1JBlyalDelYOUFPDQ8r74edFE7QZGiVbmytcVkqA3Vyky1jUANYZsfRahBm9hO8zF
3uy7piaGT5Wc2ezf1vNzLoWDrEgwPnC8fn9AzJcNQQdpoHcoO84DSOmFsK5Bridl11y5/2P/rc5D
1+AkvDiVvSzBhmhVtigxafdCxYRzQvt12sNBBlxTB7aJWGBbUo88+/FgrhHhWtDRUEEwHkmlprWQ
k+lxiUAkqRkECNOFHLEf8EBz/B0oM11g3SYUFCAsMdBetzp3KP1A0sf427vIMPZzCB8NlDEWl64u
3DoCE/0oCIgMgWhU0WVFKNJjgNyFRR7i8ozQ556KbvdGu0qc2l4TFCftAtEqDUYKlNEgnjAvBHfs
e2G7KpACR+G+fj9qDKhKzMcasQAWcuEbnExgcQC+2vjISTZvf4gXCr7TB2GykHzSRv9SmsKqnqto
/dZfutBvvWmnPG1N0VAuSiezyQWJij4s37UabfJ1JOp//hEFoDd0TKmSdZRgY8PcLrQlhTVBfYB3
6NYq191GsAC2F7ZMvsuhRzjW04jL4/gPq09NQse7x3ONkN+BqAXVqawwpA1wZmnL/P9ZMcPcg3Ye
8pzz/mJyfF3KPWhM0Ce3flimIglyD+yIZQNxFMn9Dgpco5njFFozag+c+fW0qQ4uF9zzW6/gbGSi
xctHck4qxifZax7WGjuzsnUze1s9AoEu0JDkOA18HAiRIoof1TfOWXb87TsmHLjw7YVYcA7us1Qz
dl6wu7unRy2771a1zpji+VfGWAGtsKTmg33qpGPwEcr5epjyvaTw938gi8mH0T8OanzMoXPflVuM
w5zoKtbXI7f1W4BCnEoaI2hFZwTpEzVHxtVS0f2x0H7RWI9dWoJz7onzshawdC25gOhA33iLUdP6
KWb+Bwz5gScagcxVkVrQJ3ZeikjxFPs4iljely2PQbG9/KG1NT/nWcVYXQqle92ErASJMNHDTnaF
kcyjO/hp75/upd8vnCdYc19fyvqn99bwBSHdBGFJDrqTrZxH7+9a0JX3jk9qTXyGXFol+lYMXXFQ
j3I8KMl/bApD60ceQ8AVXRvQlRhueus/grbu/MJBttdGPz7cGtvV0LwoaQQmxKqThvWJYO3garSC
Kum3rOWRdK84f0Zoprk43LM1XOg4SzPDJt9rHQzVJ+9QHNTqk8sYe+eQMwafjBba3q7SC7F0stBQ
9e9ZEOWUEA4CDShC/ZbLVQY6R6EbKYopjbz/ZOXzVb6O8JK/1Ga2qcjHq3HbPJubBwEQqjbRrs/J
au4Snvrw4Amrua6p+E7VhcACyW6iy+bPK5T3xdt7zee1pk54+9R2MAdIrS4gCMlCmHlsAqsAR4Np
3X/3WAF0QwYPCvAl1Pir3dDLnb11VE8sPXeD8Vpr5Nj0NLrKaOiw65zAT0K7dvKwg5z+YpFD8sDL
snUs2dODgIRSYa6Qe/H9NuCFUfeuMA+5rL82W/I87+78++Ox8vhqlEHGuKarJC/U7MrGKak0jfgy
UquxgD8aEEOOsHuM6w+GRnW4I2gKs3JScFdGiwl+94u/vUMGY8wp9iLYIaQJO5xCBzpKL/f76VXK
Iv/uRkeHQCHBaaYZyN8r28b9xF/fs5oa2dZgfR9d+46ucr8GWuo3NnexEJwaOJON7aYiqv2R4JKX
Xob6wL6yr79zZC24wuC8ZNZziMp8JypEuKPbJo5rs/MG/gFpY292LcRO1NYzGhQvlSf9MMatlSs4
zCJPh7y9kKGr3QkKxtOxtttU2prwqFZifQ1dWmuB7zPHsEid1ZAkAqjrynAdPr8WDzLzSxpXgnIP
S2xP0CzRxZaHQIe3+wFlVFa4o/mdfnqKtIzG7y1qFkh3ZSAW8S/64xL7IYmMg/RiOUp2UC69ZJqR
oXzxL2mTpC1DVQnawQw4fjtkJThgPbsDvxdua+upEGum9QiLeWTp/6xLupS3gy1UFR0GQvkXwO97
Fp9ZhUqs1hczRl5QHlZXQwjw1evjtJ/LvRYw5OSBPk98+39i0VH9/KolJ6P5xXCgJbmGxIH2Y26b
5Hy6GqtT6jRGHMDqTByEI9e+VL8BC8Gk9QBEKhurudd/IF99MsXTbLt+t1SDV+fq6JjrRMPFm18h
VcYmi1XN2yGgKqDAOOO4s5cTW+DE3EjYdtVDVRbFHhHgPtgh2cNf98T15FUArgFD7hMGeHydK4C/
R3zgDe6bJ08ymiriHg0MKGVeORTjYcAjAIekgpyiE3v7ljeRz6gDJlVHJGjq6g7memDvQycSMUYb
fs+fbGXESFvGUxJ+ZCzxoKuCquPU6aPZl9lSWTaOmXA0+BJACVylccKXMvqrJxsJUqeBwDDNS3D2
5P5VMkexpUMHtNuc5a6X6z2vSoCGW6JyByXwd77OYo0fl4MkarQAIdj/uqoS14zfx2MusAG8HcpL
UrWWLKe5KKbARnnwY4kDaq2Bcjw+3a+CO6eBnVSYFLj6xEKaToscfaecWqsoAIB5HEE2RanyGJ+n
n4jdy+znQ9dHX6GB/pkXi1zXBtm5XM8Wbl7Y9oZ96rASOhkZDtTM4Vh7wPkz1JgxvCvsf1j78vCy
KABHUSe7l/HaQiYSC3kRPCC/gsKCh91cnnnI50pGZQTFXqzTFk7sHbR8od+/Y5VjS25SM1tXxUSq
iWH6596CcbeyPANq15kC3zzn5YAR8rLxzOUl718NAqpBuyWPe1qQCRDGgjG4/5YlbICtBhWmk0Ym
1o8A85vo8/e4thomUuKV+P6MzF8lEh01eLvONKLhIiI2Md09TQ25HgQpy2uhpjVTEx31NQ5fIW8X
l5mtGhteHgaRurdJOCG8j2ct6NIFSLoyRhzD7SwCYRwCVW17UKd10gK7y7cm1mlGEcGFBALX76rs
4FREnuNgatOPjKIKkloV7Swv2ttWnB1vqMckfX6jKDyrEEvAyZ6E58Ity7igkAhYtGbvfPaYivyQ
3wr14aIx/L3mq9En5VB2lWpLZniztHn85tolCiOTCSwAYSCIaogK/RNjn4qyQihi40oiMXKe3qTV
ZUFSi9mCbzWbcjcU2iOhBDMJACxauBG1kfiSbT6ZyitanQ2/w5rM/2VkSAlabBMCeiMJg3mzCg03
TlX20Zh2xMaMjHENpVu/1ufpxpfab9dawCKi6gK6fmX3FerCzOu9az/svKuiRw7PxXxO28j7QBCU
uHZRdUYf0zDWd75Xinqk2Dq8mhXcIIRtMCvNKDFWlALdahFU6zDXN1oKffJbUHo9IXLY4tj+Imlg
YN46ERIBTawC6kaghD/wHKQCmAoJ7rNWtt8WgtCugs3OeiW/6ShnYRtDjj2j8W9YZh8LuVBu05bD
TqQpUMEa8DOwo57mgv2pLvsmlN+PqPkq/PY/I0xmw135vg3g98QbSz1eJ39IBCaGkbK3ZfANZOG6
ImaTfP+A4y6M9hDN7U+0ysWZ6eWTFtzDkNHyj4jDk7D8o8/PnQAkw8PknouJqzyKamUfGMsnsTtw
DNCZsaAsAm7OJe4ku7xGDFkd53N7K8bi1b6O+zFCvW/7mmJ2Iq1wS4aaK3Anvu1gZ0T+JQTjZWq/
RjpRANbA2LpIbJbLVJ02aip8kgLcWCgj5s/ea9bSLJwhpre7JIjNLEsT4z5/h8ivaenowi9E4CWv
eIZP569tatcgIeaOlddE5jIkF+X6vuRMnk5b+dn0bwnJIOLufrd9ntrqrU3FGkmqWJOKyWTZAmx9
QDfvLxVEm2f/MzLiJhvrcbRMqeCMlxiO9FAM3p9RG2ZMX5rOphOeDJJVem0CflkqXuwpQxVafpBH
ripbjJ3cJgm5xkO0I1a2UB6a/xXbloau7lHFH3jENqk5Hd23HHeblpEa+IPnKc7ICGRTxCuKy5nw
gHDxq8jSIXuimq4Ag52OZQe27oeDZEOcXaC8u387HVL+rXcS4n3gvaNs+m87vVr8J+rsT8l8WV0e
HG2uh7qSWMQWTPaygG/ITn81eWpsWnIZaDNEBL6povElicEEdSWN2BN68o46Pw2qThCYhdcjHxED
/pXASe6ZRvStFxDUvk6kdtVGwbWpskVoOOhFChkKEW6KmBqWlh1kX5PgIWGLnG3DlC6MMvZUXVeS
2u6UQsGKA+2gf3Rp+5AKP5oSEMKZYQDsmt9VB2/QWoUFuDlBLUpncexVNXDJu4BM0kk5fdJTbQEu
KK+T8YRMYkr3Od8hb6W2qaCSrM1Ei4ufB/6VB73tgrqJ5rTKH+9jumF1owYyrfWfa6Ar97XK6ull
cS3ifXFygyrBRCbIo08lupvnnfrFGK+BorrdfcGLX6Y9+L3Wlv8ElPSVWQhHLk4fe+avUC0QMXwF
SZjG+jzlEfPg+f+VbMPGjDvCdwZ5qL6Od2bI2Vr3L7mutDTZcxkaUF6qq1Stm6RvCHqL1Di5nLUU
EyWJUP1XIB2G436zE8pNMyrECUGj2GTJvxY9KC0RzKxpeMBV80Hrb812Kxr0SP3E9uuLoziC3hLs
GzHqzF1GKRx0Q4vAMA09J4iNfV6KdWvFzyr5QGdJ8fH9zap7B0h/DLYN2azk9qUBR6J7kX6M8IOA
0vOyWgViDUWfCp96xFy6TaZ75ylzHkWXNhmrZDetz9qNJJl5ZQFVik2EUUKOjTFmV/A4X21L52SP
KR0eTH10lwKYmV82Js4uz5hCbPKydzwkDSA4FeTuMMy5AJnPRQAWWafgID3++FIe6yt4D9VlsYHk
DFTCrJVgY13IBpvG2D6MMxQxXydcpIyXaIppPFh/nRG0PXr5nJOyPurhByaT3+lg1fg+UdtzptMF
VWn2NnYcuRyBm160gAz2TpINGhzPCTUnbgsS0YnHNWbZ/5IH/ijL34L8XHdA1isMhm1r8IH4gFFk
VqCUOO1RppOqTKJIrWGME6/xPJDBtztLTVbxJW23BCOlL2auI7mnTNp7m8rHei7JzsawVgbX22MQ
cPmU/6rLCCEUut1kXnF6GhCPmpjJf0Brh0gZf2E37JgGVmPnlxYvHcS07N/TYbfV3o92hFIpljrh
NZquvLUJyzXX2ICT9ZuxUFIh74NG1PqWwqH/WD+NsdxTxN3k4P3ZpdvratS+m9ZFT4DpDgFzIM1l
WxNq9nT3ZEFNlXDorez6ct1oWxoDFDTJtXQFs3aBfWIeb59NUqZX9TUJoomF6NbgyqKOsuR7CRvv
fMinFcr/kMO8kT3oy51YliCW1rszRwUCEkw1PVU8FZ+vOzStNX/7tVJ+Mqx7e0PkWx78jSDk/1wD
hpGcH4QtK3Jwu6bJxO6yM++9jGoKJnfvUoEOdYcPwVbcoa/LDbdOc6jeRcOMb0rMAWa0calDtyyF
0N4wrh7XDyY+XJCL/0EFuW4zu/7wDHIuQoewrLs6fbwML4MN5bYsiOxdC6fBbomuq/9ma2UW3Hi0
kaeJhDRJ5yBc/l2a+FLSHnnSpKIuApJzAylejEUlizTX6BAioh2V3iSRkrC+g/sQz9gZeX4srqtc
XvxVlWiQUlQlfalvJ6HsmGkxySc2Oc/BR6Ee+QJN6dk2fPLjgdj8TwfgKq+aigArUDmwfZFd3QIo
JUpgDLg7yN2Sc0+Xb/YB394Ao0z2TKMbtz3QCLxUyMhLJcJ87H600cP0ug0CtdadqaYpWQFcArXt
HZQ+KRYxZ6Xv6o4r1WjZi3xTL0IoTVdcJmMuAaHqSke/56Ts1VE5pI93IANTFFjNi7y1kzHUVX5O
GqpzL8TBDnMuSoWXiEqyO3LVGiI7LCcmBQ7yY8fXxFaYR4rdxsB42v/rBVlHeb51kQfXOaWtRODC
dS5hfQvr/FJIk+nZKmT+Dl4bkJIqYcawvv4Xtp4LMnqwPPKE+iULLhyJDO+6tW9tJgSgEVzfp3/G
3PvZXkEPYqgmYvH6O2pvrT/YarQdA7o18nLW2ZpJl5U6eMlm/zDFne0pxah/UQuGZIrQbo5rgKRU
/A5Uyp8BR3n8s9HRDZCBINFFZPySSWSIaySCJSIgYrN3ZsKcTknQVyztSDiaqtxFSKsLHdTYxLhG
QDyhr7lTeYVOId9ntW01lCfue1zdB65H4YCsGoAYuCgoK5IiwBY8WP8DF3eRGgMrX7C+nAy9XZg3
gCcA2cEak7cLvhvWGE9DevHM3QRHD51UbCmUuNUiiHj3E7Ao2tqZ0mENrvwpHLmztcy4vEnDPKDv
MCyGykhmPkg+3ZMvJnnx4M9SF9Jj2KGFEXZC+DxuzcvwMPV2xOyBomirA0m469kax8YE4sbv3qQE
CzB4hD+0HpUDG9VNFBaQ687FeYA6lbjlYPikmFc5jTXMmGA/qt5MOvBKXacrYAoNvDj6HF1nQYo7
91KV1Sp3Ic4SXGvNCPcjeU/ApBB5kMlG42RztD9QGNmytOXlODektA41Aqph2QDqEU42ZCf7NxqG
FxIOHQiLwxF+8CgjnZ+LsMz73Q8JJj3ZiSbfzvZ3zBTYJQRkV8z7yBO9Vj9EK1w52VuZGO54cUx4
kpnBjSv+65Eu2Hh1tba/A9i752W68IUkKhid4qlBaDPiuEsibtr13BTSEkPoKFFpfPUFWPSdnqpc
GBBYkVvSYPpekFfZbZz25E+gh3VnLmeS3qvHA3X7lCmg4PheQ/jlhZOeEtRn3rbKK/qqn0o1A+6T
mFo4Tday3AsdultoEXTDRxNmlEzzAGJkUc8MqxZAE24/86HfDh7eqmNGzIfDVKsMvOmJdt5px8Ze
CeYyc/SxoEmAGbOE1nCkauVvMuHXKCc0/IB/Y6bg9uK/oxi7GZ1ngDPD9+/O8ftTZEqiQt0GqmQT
8cTEyCJTGIEzzVLHe9SjBmTVs9HFeNbAsz/IVlgTQBXvNKaS71Qr2c+qPBr5nx0gDpds5H+1ubW2
S9uzOXHTC5q26sQWAsi8L9C1QUjlZxw48iNdh0nNoZW7bR/+81XIF7nmC6hXKwYXSiyd9nRDEuAe
H8d8ZT+AwH1xmtIR3qS9qg5Y2TolA5LxS9WuRU4ST+vyeiZizhR3uZRkjMqdGVfos6NIbwr4aUCB
dd21OZQjjJq+pPuqyAgPrKoePaB/JcQFcZomaMGNnvC0wtsRTPuCiFWDEpKJ4d1fhlE0dg1vnuLi
lN20fYgHe8ny0nmwRAZh/HoW/UZJyMMfHaWDXHjBZ3gDxK3p3X8u4jTC6TM3syyYfx9lAwveMbG2
0Wuv5S+iNj9E7CBL/kmiXj6IXuIEruv97obv9/HbNNiRbMUbCv7Z/SbvS1+ATLUu5vvtqMKeiUZz
ymCoMrIFkxiIuk071g3o2uebEDY8DDMH/w1yQLPPDY7PlgsvOS/z/RFpEyYskfbQYH9pYaQQDafZ
I2w4I4FBDC7WyOPGSxJtPOxJJDt6y/oQ1ybL5Uu2xia4sQ42fQWvqCmUm5wxrjUoq6MJqOmSKj/f
43FqocRQy25nMEG9gdVuLfFCDkwTBkarnYYaYcYAp9KIGL7TCEzAe0Y9QfL0igs24sMVY++xZ1o2
GAFAogsau4KhH6iNm8Gdh9Vu7Voyrr41uw/nojZk7vVzeK1cRrd3/Zce4V9Y2o7wgTO69meNWzsZ
HcwYGVNOcEfGWwy7ZV2hJysGbop5RNY7QItgxuuoQBJ6pESHinUB/G+N0LcrVF9nDYjMug+8A3Jt
IAExjlGxZDMlVAAxLn8+5bI+whQhzQZ46EZxZTksOLlAvggTm7wQ6l3P2qlUsLwYxbrGpB6bSkAU
+k0KlMwVgn3ZQMD5cEe74uKLf1MqMf7ODPSUtHQhTk20Z1+sUYNDQK/tp6zCLWzxsxvGhB7f6Eyv
/Jk0uoQkxl/gDC4l+VfbuyJWTds7fq8KW+B1Dau2OZMKzYFzxrcHHMI3kKEhRU9rtCeC0c7vj05G
j5k3OLJOj4LO98AXHRjbRF6Zo6kE8YtqcC9S1b7rbzxVACrj9CKTnSk2W9qNMFF6TmIykAlsweak
qf1V+g1oZYfKkeHabzoE7v9bCOYDQbR6I09qMJGG5ExIGc8ZxaUBZjO0dt5RWa4ZW0C4pwo1AGqJ
/n+5qUQ+jA+YmGgBqdOoy5O/mlOr9Ikd71ovDm4c53o+oq5rvP0uFs9zpXrUKgiXXsi7Ld3DGxgS
uZezZhasay4NelWSExCsmsJWP9dgdYq/ODD+Qe29ySqAPrfcj/eSei3fN2Z0RGoD0ecD2APLBIbJ
PkFFW6ZeWxO/a/d2nr0tE05r4HAjogaKpHc5qSGaWYpzNdzyxcnWt+B7j9mV9I4m1m27t/XYtXnX
XmmkJoaYDwROfx72Po3oem7OryIvoHqetrUnldwCEz5JTkp55Je+A3WAJDpRpXedrRuLnpg3o0SZ
ud3XXUe+n/dCg9B2zyhe998jDfHOU2X0BKT12KLrx2fiVHARhuo6bDk07L5aMxGEiWoLOxHyF2dE
593p8XZl81Q+2zzDYpOkhBC5emIuoUzqKnjDkQfMw878E1w0b3khl7pw+5d7PQpAROvxKAphoyja
86J3b0tX0TD625+j/UDJbYUg4gfrccw+H9su2fJ720SO+QECE0lgiJqmMxg4VZaUvZ3T/LLxrBBi
mBHJ0qG5398dVH3MjWjQ+h6QaKXMJKm25z28arnpl4+mpuoM1af+HGV1/iqkL3F6AgKcRzkUI51P
qu/Kn3w/3UcL6altasxxvbxfDmilOAqtbN/rpfHp87MmHm92RWlqo7dvH+dd9/M+vPAd4F67sQ7r
QhaNEKDSGuF6m5S7Xh9p4MvRtOqh+i2p+boQ6IhNPuu3PMr8PEgwVo/5TG3s8AjPBqPfqfctkJGW
C6VI8m8SwphwhKdM1JVDlJkjJz8qt3BdQnmXKQl4XbvtoFSh947QG4AyJb8eUMHGzeZuqqxGrwXA
n2E9kD062kQ/xPLovdUqI8fUYGVtSrd6F08sPJmSWKVicx84bL6HrCfhQ21NU/lDFMF6pIZmh6pX
GRTNtPLaLRWVSH7H3xzerXtnSKgS53M8+qZ12BjALFHFGGmETZYiLLxYvIfvP3FKe2xR86tBwxp8
tyMYFGYlS1qBcFrfWfTBeY/Rx1Xko9zdKLLrFyTSQ1KlGXS8VohW7AbmSWLrG+6LbZZuOy78cwcZ
SZ0xcNFOIgBGP0wbDG/9V+Idc9KH2s6PngQmnD63frC/f2dzeOcQ89hRi3xYkl77OoQ5jnqFznMX
5yHKY7ktL67Yaew+gyK6fPt3U344SITwedjilV+wluQwkVlf3l6vbDaLnQGnGdeB3kZiRdaim0vX
h2uaeCY89TZFt/hM7TaFJ/MYie+TFOFL6zDNoHqkn4pk9yCs4A9ypf6JwdGwTlTO8Sf/GH3smV8s
D0RThdCHrsqfIxzdDScswi/s9TfqxR6xAUqTe5TuDSoAyAJGf2btxFoV19Yx1tbkyGV/8xFovo1i
rl0DJm++knMxCkvgB1wgf2eoo9txaq/1Rbim4od7UuhbaJflERywzH7qT8TGQYEcaz4lXp+DKCGN
5VrU6DILwAs8jkOHcF1PsQPQgqTUgpNHzDB/7OQPNnyPKofiC5uFdLlrJXEat+4nUjuqQjwQpGtA
5u7t+pZcda7TrzOCeMYk7Z43BV/ELIr4Xk2QzEfbt7aglbytTqVe3YdB2SlB/QHTIsDOxxChY7TM
sh37U5BQDWx/DBsFX+h+MAIM3+fSqCzL3wOBEmP7he+9cHwHtbECk8nreq2QfW6T8DQmFHTA57rA
rdQ3eB4KBGEBdmEPdnhHyfOoVXuLd162KWFlafXzhC0ZvzJqnnX/I3mzezZNupXDotxCU/RI9A4m
bkWVG9Y1SrW854QEJd28CJOBRUnLCJhzuf/5YADYmvWEEDFKz2klYt8emdOjlyXL+I+vipZ2NFaZ
yV57QVZc99ocONMXAFHjsRaQ/vfKw6xgF8FwUCoTt5HrWqs1Kk7gTgMlaDVfOUiXNCdRg7AhQBk3
ZZw9hxpTvAl4LhGL+DUJWXkDh5cBFa1f54ih50ARYAHh4+gOJRI3AfL1WcXW9OOLtDGrqOTyI7eX
Uo83TzNgPn7HYSHSlV6fk8Yo3be5C9xG1RMPXJEPsEHz9gKMdoKX8FzOCpcUOso6Cfb6dmtvod3O
RLYSJj4vDRjsIXpkDoxmXZOuytyvElLg5kx/l/QMGBa567SojyFO6/CraGIP7SPHDe5gMwwp5IBY
eljHMry9y+4lfolbVZlCTzmHhrLDACs/9uGuscNcsSe0AKNLS/p/vmBR40nS022b03yJPqSV6dZ2
t9GapaDWlUKcVZCLM3RKjLY7SonXupOXQ+dNYzaw4TNj3eu11sY5Oyh2nWEEHI6LoBwZ0njyFXK+
XqJd5KvQ/ONkz3dD1enXtzfqeS0foCocPWArrYR+DoRDv7gnfTTJMDxqqTanjlp1qw0u3WTX4kim
yCaUeqhxNyeQpDnt35X/U64g8q0uqghD6sWOUN3vceAC+wea7ySP4svzRxGOkiO8htQ+gdVrPSki
E+S2tVUaFs+vWjBsLLhCkGOuFEcyNh6Rp0Iy2352/jv2f/LDxrd3IFQKnvbffCpiw6h4xTGXQSS2
pugOmGQjlTNj6JUnfEvrz3Wnnl+9+EnzGMaI9+5AHD4wkf8CNTqro7/KG5fLVIM7xzUu3ZvdtPqr
c1EqsdzBJGA6ZtudkwMH4WSwQFhJP3r4bj1y0NFsfZFlon9TRZNsM4RlCCA4S601MhGDuB4jw/7P
98/XmybhdrCH24r6Hsi4FOgyBu+gOGG7xGwyTMuEESugBpspBFjdd2XmWDK5SkypAlUcp2bqKm36
Lm4l85XK/12DZvhDmDN488SnKKS2hzLGJEMeMmeGYgnG1qfMBQvzBQ6eCliLWEQY2O+mN9u8vKC9
AAGNUYWzGsHQRK15vJgP9dsR1WOdNb2zxEELBxo3vHXJl2JuhADcoV875D9XL9OCSiLRFtGhDh7d
D76cOr4fFrJ0EAbiTFGv+9M+/gZZtHr7XBpVwFU55TPRUt5cYfXDgE+DBU9PSE0tHFU22PajxE33
CIm1H1BMffzw/tMH19DobA9Z99YuSzamQ9LASNMMPGeBLR3i7JfCRHn3aNw1DTnLmyrloVD1cGw3
uqlqU25CnVYtVCJWCsrjaCHZlqVEBvV2WaPIn58sr83AYOUdZR3qFY7clYFMtfKtrcccZzbkdMsy
Vg4hQ/08r3t/uV/fF1lhYfFVObur4+ANqp/uVn75jBX8HLeEu17W7Xs5cXJINTJgoChjD0/XY8nP
6VZ7iHoF0uBGxOdqV9LPOHcbGca5nrG60cOBvpJAjC7iEKSIHGVHlAu8ONN/YIxKyDpErjfkEHVy
vUC0Lv/xIiOQozPAUw4X3/mF6eGMy4OzsUlIqE44JBd2JqPEtYsGEpNo/kBOMPpBqT7P3MJFIBIh
ZFlitnuITLxAoJYNXNft92+NmXtqZlF+CaEajyjGFLl7lesxtS4OVNk5tgauap4CAMW4GQkIEnLf
R7ZIHphoxDVdB90YQ7J/M7VVBbexiMOOKkk4EgUijA+BvRPw+REEc9jY9TTQT2oqU0CxIJZLPW0J
V+3jRNjKc823WXYVjr3VvZupAuOtnwqVDok5VYiVLjE4mBAW2+fMG4ETxN1CbQuotIyo5e5aquJn
QQLakxH0pK/CpJ3fzSyAdvTtzuiPxV0a3PZaTY+PsMWIwobmY1gBQNBlrqs/i+9v2r5ZucOpYjJf
eReP47y+ElV9oBTMZvS/iIDiG6xQNJ/HQpK7bzpS4/VXZld3fkrJI36IvGOogfnV5vzEqAoaxlsU
7tLaab8BjHB6EgsdXNEPBA5tgB4GfEHl5e1jWgQtiDdp+3HENliKsGIo2QzHh5Vnm2IDsflHnvhc
EUImf4IlRw6uwxwmTjOAQtzo/vO+UkzrIBwQwCQQyLFM3Typu1vGax2Kzj7NCs4H+/0culsu1GcM
BFWIIgeuGJXnuRMvX2OtMGsVCbi5zoDIBV7yPx5ZeNLg6N/eGJTgO5CXP0gYMsVNybrSjG5w6aMK
eLMM1Va3WbhE10lEIR8I9yOiYwGuHUfHWmkUf/8X33SylQlUb+nYbdNP4e3fSfHrtIqkcTTxVcA3
i/LsQv7ktjJw+iBATJw/RDZcUCEnMf3YdWHHUQRU7eunyI4mBb8okLtKOKXfeW7vp/AEDrbsh3e4
22wpR/xC8S/TPKFzGIvgMrOuN0XWH+6QOAUjn6ZKHezqzJTT+V7AS0upqaRt6wOLd+pKV4f6fHZz
gYj8vOwav9/WZEqQSMsKS7QpZZOyCcOfQ86+39eZWorSN8XwTpZkDqWhksLh8R2aAq1F/7UvGC3i
glzDLMtxFw04p9yGlXJqTI3EdTbSUc6PNuC0KU6tTy2GY1Hxsbwx64TM8AUwvvG0+UC3YmWm3h9a
pqJfxRtwWu0jtN/KZfV+7R3P6kiST8cI03+lhi85YznYhLL1kydKBHdk4kmlMQcR1D0G2SjdJ9NM
tAEkFi5uLcEp4lTFBBlUIKUTB9BOMVFBSqtPJcGtFgfaxT5hbNV8aJ9lDXoHW/yWzx4TxSt2pKm4
lxgqfB25i+g3ssxHxSJpJza2TBHh0+lSXkYVaTTobyenUeGTUhNbpYZB0t4Ooiuw7ojeznVo6Ibp
qvOoKeiOzG/t2uf0nN9XXsJCH9S6e5TfQOOMRQMyu+nSA4RRtU4vMSTiHL5si6OggIyFtBBJaApb
/dgLzr7XD/Omb0A8BU7MZbo1djbVTKN0zjcE5xDoCur+7mChtgNQwu3pQyxgoN/sc6mXIxyDS8Hd
MjTza8gpq+9xG5JTTP7ZtuzJ/EqHsEZsh9jJAEclmhqJs+vPjgEWVHbcco3jnJ3DS5bjnGEmmung
5dVfts4g9gO/geJ/Hd2qrQ5Rr0pD8N2XXcUHHOifNEq+krLiyL4qoA5JinSvUfGilS2+QfGMq/JN
PmgJy4QQJ6o9NrqeYZgOshesEsfHFU8GYK9RH8fuT4Fmt9HXKjxykq6S+AuD5KuaKwVx2SsX9NM2
1zs+SCCgmgjf7N+rR0sv6iIJAcJ6GRu4arj86QJHaXYwqnTEppNdyUd0F4boVsSToh8gwSA8UE6s
6/eJmt3a2AmRW/xLgK0kWLDiNfXIrqtSR5eyPCIixouh+eXSl3rpLAhemzK9h7euahC0tnQULupX
+V1OAzsO+gRm9l6vT3eaR/AU3An214DW9sq5FSyvs4vR7lV0Cq5aNxC6S7P8rRxpxqU/aQrpNfWe
Dl021xccDKn1arXCKljlLw7iVznTMt1WaTdBExacN94vqOr+NhhVrbEaK0z6AKq1uUAlFukCJ8lZ
qx5ZVX7n6mUFBaksXKvmHHFlUZob8sq1KgAlR4Me1U1N51WHn9Cu/xQRIO+J1cGS6i+A3ED1Cys1
BL2kQT8zKwbWmIc4LTrS4ysxsJZUm9Iv3QGe256MFoF+AX8/HzsN9DBqmo+M3zs/nkThUp6SqvfP
hcpZqph0377yccRlilF85luB5c/SsKztn0LXXwzejoiTLsi0uSglILvd1rsU9BN3ryRlq8Y1QMFC
eQBfXh7DWr+KoItvk7B4AyADGc1P5QBtNedwo4hlnRGqUJpBkAGJM3GDUNrQiZN9skfyPO5nf2Me
pfhLx2Cpfjl9stRasiwsNoEnrvXB5XjQH9KG4wVWSYYAWUNb6azWV5ZcEw1kV1Jg3+iozpz5l8N2
cJTl7nW3C2yZoiHUr2agBSaD4lXag54NvLgQvc4Wb//XPJrbvTY8vvaMVfy/0Y+gGC4MFSqxoCj1
B+hs5YoXbl9VRt1MZl2LgGtEh0yvd9YlrRRTi0DA8lBg3HULGRpO3wiPjSYi1pkDfU5/uhN40e5O
4XUgRtvfj9dgVAhJz6gc1y4+FMkbXU+bkPH2FTwOFDwKO86Tw1wZeEG8go2SQWO81feSJJK7mRDR
/tqvbukiaRNBJiw8qF95WjueUpBeyJ4Nr6bm1cR+aY78yP3N2ZchMlvejrGJ0YD38GONxLI0hqew
iIYQbqRAOh8BDpq3QvPd02dnQh68gyTBQ4riv2Su+n9DOG22v4piUZzo0g04bL5/kD9UKOZgrr4K
cmkGR3+B7eh4J/Fr38jYhu3PegxC3YssKPKhTlqVGYzy206XzXs2S5tpu7lPREWzSknL4/zHacYo
fPQh0vVoWU6rIsa6CXwUxRSIKwfDEtqbWVXDVKLvM1vjxHpknsls0bD/u77FJMJD+aWPhI/ahF54
SzD1HcN7EiDRkmv2qLh3pUWXX+yJpdfAi5eKkG+JW5DitPMpTFSFx1KMYh/ShXRlSNjvTvymc9F+
1BHcIrpQ7VBsUlmHYlqkPIMTMlzFyzj98gAdwsmaFrSeWYfZBggnzz4szDxdqppqSxta3AAa/2xk
8HHskWhNU/k7CJuOZ4k8N/+TLLsRpglqfnz5fLOBsZYJK0s5vs7ihl+M0oex+wooDWduwWFBg1C2
2Nh2HhCugkyUwseXksaGKbqYO6pIxe1AkPPycRUO6krqEBKPOvZwyhU+eDRWX3q7ZdDE1XK4N9Vi
i5nBLYz7YQNQCCAzw6dZDTvQ6U0pAQc5z+pfTtswLxQ2bUWQ5V8x5HB7K5KmSYFVUO4oiQxWzOdZ
iZf3NRqviKsduKSZjtkSHQ2guYZBhK+ywuc5rlChlvlznGvZ2wmlyGlM2FBY8SIY7q6QZoukT1zK
BXatG113SXu4UTHrdUoqdKKHPly88ibFFo0FQ5vP5RzUsplB02uAOTOuactV0Gv2hXUxGEoq/hTQ
fiFbDFEzdm37+Q/U6mdBxsTFcIO0/5gBVahyOiQhYdz+kTwaaKwZ10/lMPEiTcpA7NRAhP8NTUjv
IlFTMDyZ4ISiN7Z/cyKkObve7Y1qfAjFqxWkfKhS3d8+HIWlf79Jo3xQRs+oSByKdWBJ1KJHdNKR
5c7Yg6T2XCBSnwo2nQYEUViYutTudearbNF4vNYw3TdCX+zAu5ek7+IQuaBritPMT4QaUFOTPQwh
p/oMslc0ChF6N9PS4FzAcB0VKkLrFJzu5cq3I0D0PQWTbveaWUfS0jiDmaaK5H6592jKCWZ90pXE
HGt7enQX9A/rWJafjaKLptQhEfTWaCc8isNHf873MJUeSZ6dRo72KV1FH206ckpdNGpklTuEJHlM
V1RE5iSoGNxCH8RulfqQo/MtdmGcck9qHMRpMVMn7e6I+DT+2ALKb07s8TtpbWfB/XT0QRuoyPRC
+vtjnjqRy7bq9pNCQ7QmUOidYWk4ERCvOXAReGSgD96LiNS4ujQPW2aJrqGc4dGMFQk+O4rAlhT5
LEGfKwIFneJomvRWZMM1WnEgNGLT74nubddVp+4zHFPQmA5/8UnaJJA3FeWh7k6J9M4UYZe77rb+
utsl5oWVlfF2npgMqw16ytsQY/DpiOejw2FNu2ZxAT83s3/lCLnwQHxuXBrRIEWRbE816X27BGsc
mkP730l93HliwyHG5ZZiFsLGUKQ6WdZgYe1Z0TsFEgVrU+aowBCa1z54p48dMfHBmRNRBmes31ff
s+kaalrdF7mpedSTe2wxgWyxBrnMofKrpsck8p/GE+EbSADgmiEBQz7hU5UhBCIPtjGpiO18kz0l
4+50v1ropiKiB2DsNC0bO22pk2cZIdVtaD71j1GTy5ikZjaPJTokRIK9rMBhKVPhVatEhJ2i2eB0
bvBwwiUw4K/zQ9+foKgRIaoEwhDE7qIlDA1tZh/Lpl/xuzwGEZBFDLemkWBROLLOlCRkdonZtKZB
47HCIgqyAF9q4EJgT9lLP8vT3PcZ1h04UuS92EcznubTeFmKI0qDl2Pa3M7rYbGq4NZ1K4TItCkQ
7NSRloDjqB8p0PrVCTZgNPflbwt8mWzfojzzxJImdnyySO9B/gzgIkvajitDKWFPgdhTY/MxF9FZ
t+JMChPLydyVtHM4O8PrIRKwH6qX4wIuBYF+0eQzKWnkO2HcaO7I5CkypCOw0BpyEEs9IvzGjUBd
5nZnGYaU/HthuYRSoSsGYQ4mVNyJyW2wYr2A9kZ+LjVJ3riiieJOYm23rcINa+OBbTY8uywq1jiR
G76Vmdvy6i/RoDMly4q75Hf52dhOqjzvvxPiEAh/y8gWBpYi/TIXAG+ZU0BlWRdcUvnYl3amROse
II7YxVThPifCAvVvj5yfv3kE8BF5uToqxqUJ5zA+/b9vs4g91kvkLeVYx5jWEvYDXzGYnbFlQvZE
X5juF+JnFKd5nuFJEcDn2O6HpjFqkzhw6kbZ+GWBT58E0dk5QxPXZp0Fms2l0wz4nEQcBqwjUiYA
1FOe7gl2OWV5qVOjNaozDGLw3po5CyAl9EhUYdOMHereu2PxElflbleml3yilZ4QIqRRhkh6K0OZ
SJnrdqqQ75Dv/NjoBsF+/kR+Al+fulAFiXmgrioIjLJs5nVxRNfF6087+1nFZhg32HWOxUCh9VSe
ouAedL+tD61Zb6Ee7Tc7ZFFRSN71pXBkE9DCnF9qCi908e3yn5B1sDnnkPncAKaf0Ddz2rLoYwP6
6ePqKOp0XHdx7Y/wvRcBRMr3ApuNY5ENOSQ3oE+nSfEcL6KoYFsZCdxgUpSnVv1KpJBxj5vTkBFC
ZY0G0V/sjSypBTrE8yipPm/GE21cfA+NmBmWvuoljgw5te5qyYe0PhYmKdWYWDOg9Uvmlu54ivar
8fIMgAegvh5a5xcwFvm59tiVjW14X4mXaGApWobIKS/QQsEOWbJ20ftiLIVUpS15I9w1lL+pO4hm
TnYg/GH/9JWY4O7/xREwoZaol7w075Ye/W0Wx6DaFebDn0BL/4zqc5XYJo0yeQuFrNG3LBCLQF0S
V0xegKj4JvWoH6nMdQ9NF34pJk3DswEb2BTT/0eTI/ym+btLHx22CGAojce1dEzjG945H+nzCUJS
YLrxRfhN254cdlkuVm9rG1zCb1sQzXfaPDE/sv86M7k1NI8CEQcrg/UrzE2gxJzX0XTFnz8iMO9a
zvTgisa+LIz/kAICXn3e8rgtrk6cu3y0hMWkYWN8PDxXF5l3wCWDij3cOfVcYjUUhMBVJDvX1rR2
aAI3D/aUB6h3QjB500pWuRe0gQqTbv9ElZnh1DNwJg+Uy5vel93hNHId/K/3lYR/E0s6KnbR/ob8
2KbAZdaxxa/+3nSdw5rrj3ePDhkMElZJml2oK88pq5v3usLV51LNOb3UwniVRBheBT7lH8JtmBBQ
rcGO/6pAuPMWWbShWExNuqLp3NI4ytKyatRnhqI/8vwSsi8rtOwpS/ZI9uHqPoeqlCJjQ5YELSUH
bWJl+/8x1sMiclN7IgSugSQlMmbjsgzf0FRofVo0i6Fw78zb9Iw0d6wTIP/WiCSVEkHxhI0HVTzG
pL3y8ZaVJEUj8UvYlO6fv4gQLfE5iz0dUcPEQCwXFxIoWh3i7k4SmmVNONk9+HFLRuT+uf7S2fmH
VK9rjlK10Bb2vETG/pNq1wyY9s0cUB/3hZR4R0UodK8m0Udbavdi3jMhiMNwTCnpLvOO1J9ouTZN
UEWDhMzh2B3DHGnSAiR29ow3FbLJiaC+Q/5Bdc1e+jvClVBZ3sURrVjUnouJp89nz+2UtZN5DWpv
G/vV0FXc2TdCDzJGkSNgetwqciPTxvESwLVfIpEnQF89rvpgPF7vybpqiClabofJX3ysVGR8PtG9
Nij6yYvMkbR2+YtqsDFbO2/aB1ut4PcN+wtasL6YTf2apEOSYUPmcaFfyLB25w/89NxRp2xuWCHe
DYXu7JiiLzzhs5WDlR/lM21nZfQPcbzf97QIKkmjSEt5FNm1ajPCDG9XcYC8vUUATLk+cGE+JtQv
GxjY2uqeVLTRkmEhJDOnXHc+xI8u86jz0blvyuOn6r62VinD/w3jSNNroE/gTdR8/mhu9WH8inzQ
4JPSjafZipg4kR0fRbGGx9bAbBYHtIYuydjGgY8sfHHc3AcgB/eUbOFY7E9JLBFYA/2qdbuLOUgK
eh1DPGKEwSCXU7NRA0WeGCQc0rwupD278ke2VOshZOVYpkx63LiRQ0Ap/ZWCe7xEdPO0bkoEcoth
7GKJmvqBryfLT4sj9HuJDHjGN4AR19fr83iuYiHvo7+UmCwmSet3F0rTe0PnoCCqYc7e3y+8o6Ip
ALFFDWonyrLKNahNYLrRssAX01Y6QXHA0Fodf6EDHGl17cL4jtsJioKHHCMmYoZLOMkNiMSaWNJ9
BhFNlVbJTmTOJtVQg11hjSZseybcyiyMJPjmOILOWOdj2EM7VrcYdfYjrFw8O8eLfxQZdQYd9xvl
z7m68+llFUxL+1oEqqCiIH+KMIGlL6BEMIP5eZN1S3ebGWOG6TnlkOkInZCUV1P3MM9Mmzo0FsOH
q1tTF14NhVfp5i4IPJMaxT1N0ayARNo2pA26rwOK5XLvvLrGnkFhkNDcGEsAhTY4kaX3y9aiERe9
L2o5m1IuGCVACefFU2huANdm87fNKc9NdN8c8O8dWRs2/N5OS2/cMoiRvs4M4iPF3Mi1M5j8YlZd
Nh/n4bghlxZmPDZ6RLXpsGsNfJnSgikgcfsrXxZQPTqfiIGfYt1pmVp2V8o+Xt8WM+9VJSj7FVX+
Tsu3WdUaTxBSvmKlnPFFeDFda46AWm7gv9VA0zCVec4OPULbRyWngH7j3p+9XWoWTsyUXX60d7BI
juDAWnWBBEzc6caAG6isD0QZjgQxAmN/MHgmEHyXtCYKeHnxkDetr8tdlTnQ/mylhcp+Mz9BUskZ
0qiZJo5xfPZhn7jMWmIWFNxDxa3F62h7vaKcAbYrm63TVUCjcqkZKzVbl/A6nQkY/t2AeV6pN6OB
VZakpL7MSnlVqhPlc+MIfunY1X1/V0j9z4LZ6eSAOiMsBUFFppICAfcjrlJ4S3hPNi+qucVJmYNX
rh2rJSSA+wN29+KN7EMR+0ho5lvUPQaRQK1VgdODdvMMs8I+n5PR1alDA7M6gHJwUrTpsyyVEGAV
nMi2HBqZAwtj6jqbE3tb0XfBv0xRTYNWFtQQYHQZzKSXTZEnPvpCbgGaQ+LV6FwmvaCV0YCLipv/
BniL0jfwoKnVhuTsoRSbY9JoiPgAmrH5lWXuLsGmluow7MqHs3bZUveGbxKkT/r/36EcHQrHr+ZB
E13D03/CSxyz8Y1ubZVAEkM7qXJ6qhveisgZ14XSNqObDpLR0ZEzppEN3WITPxOoCEHbyLNQF6/l
/9VvzZI2JtgBQRAzo/Nvl7A76KUCDcVPB4xGqITyWx17OHZWLOSGciYNsIpmZTUi9e7Mjw14TzZB
+xXati9y+GRnkvAUKJSt/I2s0IwZshoeS/Pr8IKk59y8Vqn2yamCWWRG7PeBEcRYLHQAnN3LKCwa
9Vo27nNoHd54ZPg6dKR45jWbYGkaPF7zSjPfemEy8olGxP27dGEQSeuoWVQtuINna7WbawrmIOj8
Nw+HfAQULY49BVZtZwprfMjWc/eM1jk6nRKG97uIFokK1o94oi5EC7TqGxSA/2oRwNPVuksOuVyT
8IUDZXBwcI4GD8XX1jIGIk9IEEk4lsmEana8rQULWpsvSVz7V0a+jPGkd5ciCrz0CuqxZ6F2xxLB
nJCjTkPJ4d3o0yrH0WlhqHPBZAMo2/ul3sebDfPm5NVWfkrpGtsRjBQa6adqerJGhbA5encpa8FC
Gt26ybT7ibko0nVWpyK8Ygqfq3pss58NTHfNjRHmVUM82z3MWSxn5PaMkZWm0P6b+k6xktU957DC
2vKYclMMM3lbcQKsU8cRA0UtoqwDZxYUcAsTaJEe9z6FLetX3dZrx8TimPdU56G5HTb6/LH8saIY
+s3wdVMMP5ZDjGJSt68RVc8741+qQ8S2A/Vc8XQAb/EpFJL6wi3e/1sZGZUuJeel9ekE4dmMUOCV
68OcHbfg2/q8+wOrIoPt0OKd+ivtk+LZwAxbToMnHsDbOX41cG4Wm3+OHzkBfQ7QKgXvMK41dXv/
jfL3U5b5kBoyguLQDGOwmEjcQC3VmVtL5y2IPjCFhJiWn4q/Q+MwRRaatysX0YvanW7xAZWVOTnL
GXqvw+bhHxGl/YulET7k9z4D/IHiB70X2ploo979AByS+cc3U/MLC8VXJ1JRwmQSRfXn5O060M7M
9aXYvNPNvSBtAAtyuhRxOI/gTN5uwd46BJ5LLg5rfr/wobV8cfSVeG9eexeCufMpK7s6MOMku2hT
+sneQXlXT79u6ZA/Bsw7fC+DhwBKLdER5SyIYVVs1ufSUR1zPlNxIu3yDHFaCn2O9wOwH05PkGGm
Ed7Co02hXy8m2OiZzcKTh7+5rRfdrwfgQ8jba0pfGWiSKWfW7urJoMgJ3TE6hw3P5rj+3RJ2+a1n
Iix4PRP3SW54zR2I+GTac5RzNebeCt+IhkBBtwAjCYZLkPcUjQoi32FU1NWcfXD9Tlb2OXaLyBdf
xHvG+MQFKUverIRuCC8reOrrwVhEgbLTNPOPAHJFuw6t3fZ7QfpwF7zDUrNGQB7m7m5JPExxQint
/RrH0LBLrEPR/+6COWf1piaMiV8oXVM0XI/Zm0xk/rjWP/7/Z3Yqt+bE1WXO0R1T38aqCUc5C9Hz
6/V9jUifGcAwXMWPq4apuKHnaMDUoZ/3IVbEDj1LBHfkQ9vw4g9Key1DS4bsTGdUrE88gjaoBhiY
/jGik7EpZJymrmch6p9Wu0EoDDqYWreLWEdfIblWJvtEeMzZ9tbMq0/rrnTlVOpu8Sw+WgbQO9SZ
TkbOE+yWXZxzRQIVfGRA01XacVdrFqJqn+WolQydHQudx076gdv+N9mdjZqgSHko+BqBKNOrfIIJ
eIW7Bz4cqtHb19+qHNj0DG8RYVym97BadLFENLq9TmE8HjG4BP/244oYVwUUyJb9H7Nch/9Eltn9
FdXwZacQzpEo40wKLGfzef/74XAJE4gwTs2opGtyVFHrhBrgjHdKVYw0T0xWuFM9tAyNJ+bqRA3t
8cPGi6UAIv68tcQgS1IhFu7A63EYi1V6vIGEENw1p25q4k6h8WELWScjb2++9jbUkzl8NurQJRUc
0PZ5ydImSPBfz3Clr6CC/4Oc2513MaEQEKQwFyTHPnlGOfoPiDPh05WBM6P/ek3exRBFi3SVE2ud
ZXBjtcLdTk7Y2L6mu+I4L2XjqdW+HQIELXGoX2If71aeH0UJTKiHWHD1xnO3iSMsSKgbO1bkGhKl
yhl0Mkjyvm9B3r1rUTRWkLVvTRzt4xE8O5+rIHXV9qLnvi2RbEA1B1qm2SERQl9PQckz3+ZQUEUA
gnu3YIuYaKAtsqe6cJ9/0/T3kZXR+JaN645jPBq/cThy55WKjdAp5v4wdqyCbplFudFFlA5SLQC4
Tfy428weNvlF+Bha4A7YZYLebcUsAejnIEO4Xo1Waf7vMTiNx93rG1gC2wqFpsYybhBeLtdQYts9
u1K1hpgsjCI1WMthSt/ZIWkPl0r9XxUKFWxnzE6ariQ6rNgdU+cwGYfUCpqkggw8J53hrwj//JTr
67AluuutT8l8jBWbHaq6oVqTW2XgMhXoQ+6o0/8M5Dbi5Sg5sXWrEvWX5hIqkWzF6PXMGhUYa2n9
HsskK8yalohBpjH5bj/Zw4Xc8CFlAn8aJ6mEtqSbdHxq6oAgwBCEKxD9BGVBuS75AUL/+j7BYUyy
h4lCd485XHhYapoJ5Cz7SeMNgb+DqtDOqhTiaWSxQtpNhC7iCOCq3mEZm09E8JwS5/YSSWtn3XFp
HcNrmSZWmNGEexYWeScUw2NT+y1u1eT4s9Bsp9UMSf1WnrCpPqTHxKqUC0A5UDlb0HZ9lJCp7gDf
gf8p3cRt5oTPWXpxzLhI7hDLNOig0P9fDlZV6cV7ZwLlmYFj9EfY2ylX4wOtb4Yj0BSStfn6wvT3
Vb9ys6qPDLjcXhDhOjESDaK35Y/lqRuC4IyCxzk3liQ9YQmagrbKTdE3y/e2lcppu4DLr0LrRMf2
HyS5EJLC9/GL0h/meq6wIhGHDtFREv/t7B/QGcpIdaWY0+dBSIEvevhHwnZ/jNq8RjcdvF8tcrQa
IObBvHi5W5WIC0zBAV39LQ3oTrop8asU/PwK/AXuYUxGPYTqqdH+rUwPg0gr/8H0Wvcpj4S86fLo
z4TMbKkEAhnzHwZr9qPcDiS72rC6Z40dJnFx283K0GRm9PmnAUNVYSdYbBfImztdKwNet5CTq/ee
Fj4vmmu0h/w86H1OsaCRPODheQUhiomzahYFdwWpuy4TULUVhnCgxjtTD9ku/G/C54ekP+qGT46U
xeeXw7E/knl0oItk2bGg8JEGQBQZYD4dzORjt1MpedihlBmfDtFiqc7BZoRBX3IoimCHR/c+r6lg
4CBcTibQjI3d/m+e+DUAGjCS6fI5VZcvzu/Dl8F8QOwwS+QpO+NAEBnD7HxMvHBsFP/I29tQKF2+
oc3I+GzLWKHEmk40zTD2oggiwEEZfpMHiUQSVkRjZyj2hLpjQ7pjCgv3YkVV93EF2ISs8FRvLw43
mniix5bpqfmGVXRQqFW3FOH5OBG7/G6ySL5v86lD4HL8+02D66r5elQQp70AhTx3OLUaRetDfgZY
f6ptv33kzIAIPj0F6kLUVwpI2TA6oP4IdN31Hi5m9wRRSeqPDIZxWsUWdrC+A+tcpXxlUDjDyxi+
/P5cnyI1vk5PLT45zH0zQhlWjLGKMn1lrg0V3QKRIDMBmAceUavahZpznxWxvOJEPJl3EaZFh6Q3
0BOfsh99sN5uTCfTcch/agkppYtzW1Vo+Rr2LchEQRQHGQUpmwZ51ZqocGHKjPCDVGndLthD4jl7
4EyBKNWJG3YwXp204dlrZlAmRPY0iNIwMZlfhjRE4dTdzWL1aohzjCGLYEj1L08HWd57LgSwezR5
Zd+PAPx+2vfjNGJd2vTJMyz0+Q9x8/9QlJCUz7c62ZcnrN7/t99Ql8EM2kliZEE/CU8CFnCDdvaS
YmF2nZS9firg0D2xeo2sNlD03mNLYEVrfDY6c26IQ6qu6yiPdDkR14V80RSBarHFyJSUyCbrOK3r
IK1UQhH/VWfcUBeA/gquyrcJytyU99dBGBTeJlr1rdTr+L0TKLZ8UDqqMM5PTJhNLE0uMsEI4Ty9
KaQZ4H/EF4zwUFlFVooWD+yFGBK6crRUfAa3ywZXqDdlF3tMyS66AFAzjejK+FusAPGsJ1+M4LRP
BpPF0VdMnp29Hn8dsSBM7o2Xy8WmA34g4mBF+pir/XhCHgIqFzABi5Th6M7RYnolZ8i1CnQrQxrU
WTYVnD2ZCM3FEi2GtBf5tn2TfaZPN7y3rGb2L7Ac8QyAenpa3l2FOQSWdkaaZMC4OpOdTxUlD5gA
r+eCYtAFtgxnhIrM4wUGM7F3B3Bo+wl8+nuqUR3mP3A6YZAa9n1yVmSvGFYeubVGnf8jkm4SWB4B
KT6Net2Y6VQz/ms+JmXQNEaADaS0rrLjVJymHlRmh2Ov11QqW4Y2wjKrAGiJzTpwyL5etGnsCCv+
VlGQlx1Q/Rag28NG0/LQSJyUQlx0XRmVYA356c1V/joFt8yfEJcoQ1YELaPxvfEuJM5WoNFMFjjR
MDdPNiAF5iYXYak5vIurjsthXjtd6p7/dZad9goC7NJmvliGWYTmEV7lfHdnZgPAA5fblH2B0Y3p
fDb7lXtdk/xq1Katm9uDTkRXBc5m3scvZIAID9c7GOVCbTe8XtyYu7KsDBFg5c2Tcdle97IKPzVz
DGKnoswJm6BwncS+HwgoVuUjuwlqwxbByw+3Xd9BJzQdSswJ05kBCRMYNdSZnFBpcfnp8Z7JeRY1
E8aBQa1xFV7nH3mAyRAa5LKCOZb64J3pGfB9t1dAwLizdDlBLlWcBgTHiePq9H3qUjlTT4ZQNbKO
hZ/9A6p/FQKlU7fMFg38IUtucptso69Yhw35RAdlnjrFQITvZhzs0venHP/IzfKzQo1+Rtcktlo5
RB3fYz8gfuCqaaDgWbepBtMeF3sGx4KkXEBbjlAFBDwFk6d67omnLAC3ZjZgAbF7YjjnGrz4Ik78
SIo7C79Le0G47FanYMq+f9Aa7eyc1E0qylWd7xicaDBTNQtVzot9JoyI9BM5Scqs489w7LeOl/r2
GmExB/SjS+Oxb9q6lm2odAW5IuPAkCrBIpL5UZlbiCdlrpn//FNz48vQG5Yxp1V1b4QYU5v+XWb8
BTR3lPnhnfuILPfAD3GE+vgygBWcFUhslbItiZFKAIx4y/vgS0YnIs5rrTa5kLpHyqJMg3bFd8HO
6+rMbXFYCBSxPXfG6SimxE+RfXaWh0it5hFiFo7CrELWhm4NDhldlET25nrPCOeKlGgVwaKkqhou
2WRPamtPWs301ugr/mfPfiXj09h0OJXtMgPP3S02MEStX+HuarQakY85A/PPOTBPF+ckIZfDav+c
+JD8PAwT+7ayKgY6RvXC8Agyi358yo7C+qk1N3HwRDANGSz/qjfI67UJXII0lZRezXF2cUhFkB3L
mvnpsrTtk9QKQGZaNVFSVUL/Zaxq9K+lCvqs+7RryCMsP/aIljvQ8Am6xkPfW//ygskgcibl3Mao
p3Ao7CKTkgHRH96VQb2GBZzDtZdJnN9YY2dYOg+wTTUxjy3eOinaBQAzMiPUBNrqAHGrR8xNhG0X
4uW5VbGcHAElIe4gZY/78qOCi/R4n29EvBsKxK0eLbi52oam0lWlnGTrX9EzTpRei864hXHZA35c
LLdFa55xidT1Y+UAvZJYrpuUhOD6y0FhVmLH4Kl5y80xXxkCGM0FkYCElS8bTnsnJ8l8nyeiWQUW
FGG2oSzIE3/wkdEh0v7xtMgMXM7ppwmIAc1wpL1+W0xPbKERaCVAYNMbiHRu49xTz7gQmVfyLvEa
b1i1jSl4AgUuEAkC7MjZwVxSZdDx7EERkuQMrJbaNZp4olrmeKOTcDk2LPlJgaiWlju10/4Nfjnq
G8xbJFwPAXWXNbdlGtkje01sgj3Cx5n+sNzKk7NUkiXyeWUIEsshNUPmdGZd+Wtds+GDv3rk8zAD
yQ1PqfQj/sAZ0mZ8KvqBeJifStPNqIo+YfuOlo3yorjW9gfLYow5Dty8+dRBm/rbJIMm3pDemw1q
ULG/3ddZ8mfFs4T04KxLzswlKdGuOJaGZtcExLBrFs7caYNh/0MJFLrxTRBR80C1FdJ4hOvommSV
NryS38gP5nUjq0eEwzOk0adiY63AvPQmI5McTb4BvKLor4X1dCwB/5sj1DtGHQP4YXe/tmcSz0YW
u2YLcE4HMxcI5er/a39YZESnXbCBzOcklAYSnQTYhYkO3Iv2/bQ/2drmmfxTvkN2jSAgSTa+oMdW
MN6Dtvl9gH78NpeSeN3I44pgbHUeEgt473mq+aZX7jM8rjqB2eRQ2fY37FU8WxKQaqwJJtQBP/BK
fWO38vT2ZJ8SCICHvtxpChgxEV6heBip7ZxKHF4zgBJp567wc35TBmIc58twQ6FrCdfPPS3gvMHY
yiiPucp7GsZd5CHmU7VUHHzjsAEJwmN7mKk3romX/3PnFhQC1fGTMCsD0b/ABzZJssy83H54sguP
LBjuTsfoni3mcvCaBYytOfNKZohFEEtRcqjakV71urmWCMxk77+ONCkwhp4a7HbvfRX+i9v87YAn
CDqdSzAaPCxOf0/vBgzVAKruCnavL1Foudhf/6mTYLpebxRAs0Lbx+aq4QLLTkvlIm6YaXy4Cr3U
a6K2jJVZg2NtmZ1CWi/mlMriNPbGUjl5wpfd0AH3gBv1m46FUsM8UrecN/TFz2SIEJ/tqF4/YgLi
9s3UdPaOiQXEIRY2V9+WU8GzctFmTWoFLMnrSiMnZQFPu+wdcZGHmnGPfYAflBG7tgK3KW+ZQ0E4
ySFZ+TxhMILT4Ql7vMalo8DpjW0rjpokUITENin8/2VD7MxqbXnC7dVhhjdWPkO1IfFAHbuH1ADT
Y6QS3+J6btoj6WsezZteNn9Ke+cyuiKjA1FtKVjjnEAWaDdOQu4nWE59gCb7UhklIHtm7fMKDvjR
dwaGuQ4MaFmWNWgAa4nC1eFwiSkAI3RmchbuCwyDQVquLngKsPovjcycSabNerBvful5u1Gn3sdN
HckyLWpi0XIkjW22CqVvHobKND3K5sq8nLK7/Uq2oJKBVZretEEKB3wKMg2ixi7SGvuKhiKKshQ2
foP1RtpAan+IdwosxSAO4f5+cRX6yflPVLNwCQ3U+CIz9coW9/CMtVObhW+4aeeX/8U+XqPrxUY3
lAXM9aP3l0bhycgbs5dbzkwihqwenBO2KmCpmZ31IUD9gpCugUAwAkiisrTMv7SHPAVPbyUH6sFp
SyFgjKE4wdYh9K/4q4FKgx/xWFB3AZ1TACckH2PqGV9wWkj+cdObZmMstfx7eW5tE3PSPLUaWTwS
gX/fkfHNzoNMPSqFGQSXkqS3dZGyEhTnQQIn0J+lEs2srmFMnUK3LJZ6Mey2aon8GwkVQEvSD+dR
p5CoLpCFPEAIOTSwSasj8g9usSgIc7OhWg5YeSdk9h6ksMWKt5S9XQdC2qbjxGJj/NpKe0uKpQu7
ksTtB5CbyQpdvaHASDV6qtkOLftOA8Foki4n8Wx7FgrJHgbMQBGQBqGhrxFoQJZ16m640NLw7eCz
cA5O0cbB+ljtkcF9PdUcHgCsFVg7+SR3/nbqdvo6g7Fz6AUkBflp3edNqVYe6Y7d/jg/9Y8yy6WZ
9MCgXfBARzgLFGQArxMw6QOus0xl9HFZTAYbRtmIi+jVdXa+VUmaJ7846B5dq02U50dZsYgoOMlm
N07P6J9O+AprGABhgai+QaHvNZrWcoZKxUy+NMrmxuN8fuvSrGZk6B06Arw1G7+6BMsvv/ZpaGNw
Gyowjfxu+yA7NbxhynU/ufxzRdRlkYXweUI7NNkPAITy+2ozv8YEjy7QC6Lzmub669uG0qUBCT5P
nhO02A6a2Vqgr4NP3mZfabdrskkTpswvidFBxj9DHqmlO07z3FUIYILURz9G1xqkoXzSVmypRZgW
hPuVHVXvjx3tLNHwBJqMNiLPQpHE7QfGfY6wOcydN+pZEEaPCHTbgIA5pIYM56KNz4celDMBPdiY
gnx3YelRKA4QKtYGN8/S+D2ry6iW+F3bqCK/EmLCktlaNGbhknsrxY72kO/kuYJLdBpVofmhxnpB
lwDvgip0suEjaTV19x58A67OKRjTJis/Yxx5HxB3isUd8xMAcze2XEQjM3gj0ggQYURmffPNQrnX
bENGdVvl2N40tB4yxq1WZGRjmTY0+yphhvoCql4e80fuYipHl4NNf+DOpntWpnHvQwCX+lFhIzFi
6L9qSmoNnjF9cCszDaV/Ydrv7la0x4oct8V3h0BJVIlnnUF98+kTQGXqGLmWBRnGz62/68yFH3bH
4E3fejIPJXiwtNN1djLjkSMP3Eu0jzN89c/dU51U8c88xjO9lcq9y/clxtqQ/QwEv+X6LQXb/f0c
hGtCxKzbjZ59SS5zRY++rJzCnF+ZBPkp5wZvcMNZzcu4g5VAuVaFQcxF33ZeQ5MGt2i8ShwYakn/
VQ1VEWlTpsrH65DQPl1MGibCCg1dMQutlY1L9D+xrFS6Z1Xqr2C0j2IWh84hnOeg0TVjrTHTzyU5
qATjKPdqB8uEeQfq4T/VeuZqXQHxjM32WuLZ+XgCjVdmgiSns1YKYOZdwIH4klqsmn1b51SBxLmh
jEVxvj6ciEYFU2cke458mtJAI/PYkMUtzc0XbnzMNgvbImRJKFVP/agoDlg5M6XLnO0Tf+twfoyt
GGz8KSPwKIpvgNpLI0XVBMlUNY1yIhJUdvSquFOcbhUdZEt/98FNHSIeo+3HJEoRHb+KIE9nal8+
leikAOTM+XTUb8I9CjUimDkekK6vWX3034R+ClouDUiXuTWUJQMAIqRgyPD5Sh4N02RImvjHyiDN
XO+r/KZtQy6dHWwLeiyz8uRVbde+nL6BgDffrhf2s3JOlev6JpfppGaDmh6e0kw2tbr4OVWFYdsd
KSuWILzGCx1WymPjkTKwUUKoRQ5RVyEtud4aa1aRXYSoB7BoCnC+oK57dfJoJpWU8nRnSMrKcMW5
t5d1a4JSszAyxwmKSXZ/zqq8+oWl5gARjUnJgUC7jCCMY0VcoFNySjTVdLXCfQkdbqcUE8Euso58
SlVnD3AcaWF+TnjSghIYJ3Agji/xBm12902Is+Db9IUh8c5kAZTySqomWDUZWUQKPIiFOZSPy/22
yNPPnYokXGgvCGADrAQGzE50q0WFMTD0f49sJH7gSztOqUgt+JS3FIZulHXmXi1/R0MWrEZLphFt
Jssr+ItEgMlLL0SCsrafnH9mntIRTzYWQCLsvlzs+sKu8PS0ktmwNkrhOueKQqWLEUspNT6okfgw
NP54IDumShR8E25SNIzHUo1NBbnNmJygopx5xGMl1BwjzEPOAVWB5XWkA4StJODSfGN9o+EKInjX
AMC8dVnDikpCUGRaIJ9a2IXkY2TxKdPHAq0HTbikaWNXlZ5BSDSF3sPm+jJjVVplywshyNHEcaN9
kd/txAwLepvo/vX5ceA8H2T7Ch5r6LxjPD7TVQAkdbw5zhY5H0fwrsVy/NkM3UNbeo9uyZpn3ecO
kRZkb1yNDIJMU6B30Cp/y4rlstpVFfKUXwrhq1Eh7W/bnbxhfw7MTXaclcr7uR0Jp0ONNxdErcS+
zoyI58DPalW1BvqXH1+TNHHQYEx7xpLGJMwzVFuW3d7ZkEpcym7aGsURPFzO08TSWidKeAgAuDYL
JZfU4eV7rIstP3/eg/PMrEuoUkgxQgwk3GkzsqoOK1w1yZCwxMsUvc2P/7d1N1LMBorUEzd/lyWD
aVrm86EcWvdnFdhkWpDlWF5370+ktgQPgsa9L7IBTBRIyBJHStgQA/ihtFQSJzK27g+YTfRzEHS9
HMv7O/4DtLSQzNTsAxAylurhm0Er3vW/ObPhnS6hNtgDwLd7p5nBrGuDz3o33lXnJJ/sL3M9zBXf
st+zEWIKGQah16ozj6VIc8bzclhKvH2Xj2re+PtYfokIIZqePSGnFJWozTojunqI9pYX60e51bdR
mB5voi2gvJfCLlW6Gg7tKcbCi4Hhy6MrSA6PHgPHLQ87sSLGyFi+xlcnnyrEib51NwYMc0HWkMe2
fzmrd9IW77ZQWIlSGkU96TZhgSaRPPJFi0f9xiGGlTpQQsjbVrAxzh0aTMuTNqJX9ertiSitnnQd
K+1iIPGiWcWB47T2FfHtOLZqlZRRW2vxTg20PW9uc42zug+AFyf3y80Z6PrBV4vZhQZUQTHFIDh7
Ddy1UhW+vfwnqQC0D5ufQ2iltu5WxewV8S/piSdrzZW5MxvMZbVdRXD6v1D9rnCvwKt14z6Sagqv
1i9QYkAXc/AkZ/7kiyr9+4fHGpq7gdni4yisn2X6arckfQRgTakn18rQgb15EVQZk7z/XFbM1UAW
TnijJ15/vlpL3BwOpiqw8iuX6vsvZF3BIYrnvPmcnGlOjt/Pr3lwpHP+0CIC7GRqBdAgp372es7c
lpNWTqMCwE00Hhj/Mh8k3D+xBYkWE49Nb9lgwJCeDyE+bQRmwTe4PPRU4v5VkpHTTAkqcZkWbJg5
X6b5wRLh6D5sAczi8pEUpUfJKROdUhy32EXwxtLHdBR1G5D1jKtkXptiLqG5tC/xtic2sX9yXY2w
hcisjQ3CXRGNtkgE5Xe2F/6xEqi6lRks4KTR5s3clEQONbBOJl8kUA3HJI1Y+9dIOpldq+iMkOQJ
6FuGlCpAOmueQy9IFzvVR6upZugUxcwVGJSA9n4gzzRXgFgZl7al0nEHGLT79VfAPd/shma7kbuv
LdGdwzEjkzK7F6RJ9qj1dFJP+jsuZzBmetOiTuVb4e3DNDnEl3dIrbmoxXt2eS2AHhO9p+taK7+B
gq/FLILpEvwQ0H2xSXRU5N6RaVcg5pJX2IhKVjYLixCNDWKMFwkDuaFkuV9cnaiNjR/+3DkVWgmL
TW+UBlzfU58zwUPVwF89osHG+7QHWkJ5wDOEQcxU+nbyN3xcw5QEK70hkQFDS2e5wOitdJlQUVvZ
gLAJEMfNPestg5OQDqtOIkmi3GWkrLO2sWNCUFpNdSbEUWUbcMPYR3Rxd3jmKwAMJn3DhZyZvMiL
U4/nwwtOsbWzPrqkFg8tUJGAcjr5JGO8jmRXLKJbMM6HjhVijlDvfWM4dAQ9zvLVYVq0EidOTG4n
Hg3zsDeqVSQUnpzjtuZMdaDIIwFPfQHpwrQ7lCuDa+8UDFtNfAw0Y0sFKP7H1f66Ka8WlXn4eGrq
iZdc8Stt4IGgmvR8rN3rC0tL1PVui+NtLgmoxRsjUcgBhGmn/5iOYCmOhd6e10WauepBR+EkmDvQ
l1bFwAud4FAzQ7N3aXFyAX9cvoQqtdU+PU4jcg/LspKassenXRsoWtoy9pD2j4ekODDk3gFXxcvH
IWkCIXG4K8H3bUcr3mLf5DOtoxNMcnNGpitU25Dny1C79JyMsLkPn3BMSjGGvKdjB/TBwjKP2/L+
GaWqoNSI9fzrDZSx/f7KWm9riFqQ2MQpHueiix+O8L96pp7OcAjKjRE375o8lOoq+bCoMsIeIbMy
dutm6EkZvSeNwPuhVSP/+vESDOFnwCJ7cU3DpapL0+0tk3u/RfOddq77EDF7nDceEPqt6eyyCsVn
8T3ei0dsDMMVI7tjxLCpvs9YpoFnI0vSfNaxDHE8EkMpbDiZxBQ6/Vjp3o/1MTp8mDtrCfcuxxM/
+yz1oMQknMfRDcxJY3zW/PcxbkgMk8070Mo8+HVr+srHVRsGrZKue384i906OsYR/oPk4Xb9Ns7K
8Hzk6SgX4eCgOILSbT6NQHGTm9doOZzf0DdNyc3F4+nHHdKVZBt7KUFfU4GUERJelF+VePCe83w0
5GDUENa1nQtyLEBoGUJ8IxbjJUctctuxMuh06ie+Zg0C6rToZub1n8coDWKJjN7mfoIw6oPqBcZF
Oau7HS3zTeTbA/sF8NFiVpkxeWoMv3odcPwvbgs7KvBfG3Q061BILsst2jSZIq4eNwZhLzPx19ne
xrKNk0vTgapQIUj/5O4YRlBRfyK8qfnKY+JOuey726iIqBR9nkhYBGAa36xd6PXbm45a2Q6yAB15
DNaV15lG+aYxZrmmNmJcC79TgKJBxdDruSdfY9fd0cU7nvvNSvebelVEDkFYVzgQgi/GqDPo/oja
E13QrFbaWg31l2pwKQ/NU0kUAwDfi1RBUVRaCiuJ7H/zr6AIVIezw+D9CjcNQPQWFKbdq5YvkV85
qN39Kj2ZWZfHTBBfG0K9JV1O4vnMYLNw98jNL2uaEZzp9seAtGXQjiuhtQ63EcDAczeT2NM2NLqL
XMhnhVNqXsRx+pXhxKDmgnlM8BHQevtvPeoqYnY78IUgAOs9qKFFm1o2a74Of1wjDG2db71tKN3m
tSlqxGGDo9VldQhvnes02EPGhgK1CjgZHYeMEM8wnQQ685wt6Q0ibn/PuGzjHMFd8Xca6zuNcrkY
lj/lNcQuQ4hzTaju/bAxUDaJTD0SQcYb/mWZildHcpBD3EUv2SZuNgPgGnZzOcxz/V2VE/v/PZp3
oOx/XJ3ZK1AoGxOYeWHClQHDYXyZ9XCN06nO0PeLt7tLBQzB0cbstlOVYNyVCG2WyUFfvJ/pbUk/
dkFyJ2GRQcd2QeBDE5kOXp3hif61sLuRJLHiKvC9usz/2RZIs189BjLlAQJmeyUSSs/esa1PKOST
9QCR/0YS69NakcmVqLC0h0oM94vFkubll4aKHSwkMhGwGEBU4PsOGbte+eFv1SLnBPWVc2ph4GGy
JU7SKnOYUUebMsCfWRfGVMFAY6J+brAzNr+ToSzotrAIE73MwBtK389483b/Z3m4RbP9Cw1SnyJx
wdSFyMLEJHCjNRTtohz+9eHbBiwGwPKh5m9pkRlrcoBIdiVfnWO2Feyo54TpbbXIbC3lwGQSb43+
DV9lhaeUJhWve5W4ep/3E7CzCHorAEeHb/AmgmMfOm11sycfLrB57aTGqdgicttAvsVjCamApqSP
dSVR+ZX9RWVqTtRWTmgkeeupZ0FTalE82EWS33wjnsb6fBPl8aQTX3gxPsBbB9cMh+MKfJL1M0ch
akk63Tds68Kar/t47qNAI7xHKc08IT+vKmOFeilvNp8VrPQm4ej/0AQ9tAbI/YBhNHi7tzoYODUM
XPFrD1wMl//4ob2ALIJQrixTN4QB76Mh+Ihu46ZFrVBfGdvhUbM0c0lcFZYeqP1Yj/+mqixvNRJ4
OQMVXCl7vbbBqRW9dIt51sEerbGnFPH0mClIXCoMGCfmwYGvv1SIcCxm7Xh1ZgBrlKnzqSYQvLQY
CukE+6mCQeBNnHt110QTu5a9EyA4F0bNvfOk7FJwsdIVLwEPmy+1Zou7HkJf5W8JNtep9e0obWcE
8uOLLN8JBfnY5pSH2w7hMSBUD4lQZqeqoxIUm/+0MADxc4DEQsscOEBYcB+oGDOTYrZNANvh5Q0T
3ha6x1rHYXJjU5ubXhEyLga7XhObBQKfWANINUVHvzj0CKah+/ieSAxSPhy2nJ15PIrAB4oYvRke
8H99yaDpJ+k1INmaNiNZEKu43js9M5xE6KzvnT/Uo99ma8M6g4Zt9OsX7Q5rBl6z3yCJpsRfLF+3
QgXuB4Zie1IHxGnFX5nY9t64H5llz6KzGFpG4zeJlRhphHKRLvpiXNz5z4sUy0iSkigOVFJBzXy+
XAr6eprv4HoHFk68VG5bDJIxRLpfxUwErOCN2hsRZATRm46vhFcev1AO68u9B61p2jCH8lYWb+G4
oesQWOsKCN/9LEL8FjOXyPnAZmxa7jjaWiv88Nyk3YAlTcJpu4wwiNbEr9LuA5KateY+i3YNGGRA
OEM4m/YPaqjQax8fFnBsvfqGLN2181NnQ3oN+DDboMCW0EKSjIyt4L+slcm7fOTfssGctNM2gG81
b+pshopT6rcVqu0HovvG0IacY8a3E0GnBeCdVOWxWYO1z0x8Mr+PTgiz9/eMi6nOqWnlBP9TaThV
kRFuuwfvMQNFR57exRPYHd+GBNZKWyCapyD2nvdt0JPUynNDGKS2XwoF7Gt2nh2YeBjBGsYu71LN
qPmumWbFR3KK+sAeZsv/lKTo1Ty+eUDiGFyVvSJnJISQaiPz4YWVia/G+KPdHecOn8wW1lgr93od
oZ6HOlkOWvIUKrGV0F0sJWPk65dXz7DQ0Ane32hK2clpj3oGR/fTa63MyJt7mPIo8hQywRXRniRq
wJhUcUyfTKkATbBVjgMFSgYHH5lrzpyivIeqz2wXuan/SBhJFhKUUofwXeWuLEzCfyh1mEKntRCS
0CSjTi4GbFTl3bGVZt5QglI2AKN85PPisLJhiT7zNOHXFWmq5E6d4uILN2mg8ajNYIoO1KmL2rIO
0AVlEz2kFZHNl/2pUWux5wSjWFiROS8z5izCAfLID148aw6QXv7tbC2DwMJPVquuY1h5/pgLOtLa
Usrc890wUhOiQAyHRBm8To84WCXUdeOtX2s1xjsE02KMpUsR1yk2kaAShumVNJX4BkyX6uNqFomQ
kd67Lg7IQHU/OoX7Y+vVBMng2Oh4AZfeGkSBddnveV0UyvBf0lEwD0gNSHfVbUj0bULBdqNO2LvZ
zMd33c1l4DxAKPQyVuplewPAAQb5EHGh6iRPYxGTZa2minSVxcQ1MxS0SFBBOhn5pfa4qs+NiZV6
eOkkbC0dhr6e2TOs3TvdRFiobQD46A8ZsQUXEnFhM83YM9leJD80TmOgFAag6gvu7WPaqocGmunP
eeRTZley0bt/WDZiGu8xEvjBpb3kEY6+eBON96xCbhBC5/Oon1bJN42hG+nlk78Dv7utFL8xOFkH
grLfYPIik+cgtFt7YbvIq1h/N3KcU6mbORygXKt5M9NlYkHL9yDpINas8RGn1BZnap0suQYwJumT
7CEPgwEVw1+GrGO8a65909waofv+Q0DZAgxYtr2YGoj5G60N2HWjnIRR2fXdG+QNW7OQORsJ7g+Z
kxplo/c7YFqA3mdMpIymPLjVCjraeF7y+UEnneYBiWVEfS79q9P+FoLhrliLRlrGSM720e6plAKL
fS4HXI8jQATeJq6XUmgo+jDXlNkTORFRnxWmURIoCQTTxAXAbfGwp6lfOIuz+T1JNq2STm6FZtzY
d4IRcdatEmasMdRClTLZ9TN1IftTSEcjrXewtSUYMF7L6nJHQGydUAmRF0+Sxn7nU9rZuq/9rHlK
SXmXrta6jPxuNvt6w0L0J8qlkdDoV1dvU7KbdjgCYsEFWBO4yFi/VbsXFGK2HJ6QlOZjbrmI28pI
MIxrauzETMX4iucPq1Ltn3tPdLtznr6TwkWnFg0grkSMSJkZflPOKU3lSvuBDz8sUSudL37sQg2W
dysio5E3j3tkoM4FVBR5ZgB6tLIUo/bwANJKMgVNwTzkAXqon6jay0N965B8va2qRIGrzrHe3XFT
9WQoLeDVG6cN0zxEB4WFzwTPWIMTQT/RS8tVzDr7x9FLfvDGZ2tJzlyexkv2FIxzr6K16E+STXcO
xlUSJll68byj2fpM5GUqt64WwIF1RgbpyG1cfGajJ+M9A8CVWri/zBVlLghBMhhgI2Pmeu6/yG71
WleCbqR/NKuUwgdaTCC18eakyF2ER2ZJEXO8B2XIofko/XM6X2pWKhA8wC7NC7FClmzNIe9GW9aw
oagj5wkZka1soaRRzPG8fihcLWvS+4Z4S7ykxLGiwDY5g55H//ip8pTnnOmzllAPOh8UGB3YDu0P
GeCMTX5PUTgEe8cs06u8+VZzjUl9x1Sb5h4yoKZYq6AH1pWoHNVQic3hjVoRbW0TRLZkCY9eB+KO
Qjgf/+vHL0UwtEpxBe7qYvE5wxk366U12NX/JAFesUeC4MW8HoyBstFpXW1BDFwxdc0PnfxrdesT
ot5izC0sC9+0sVVYFwEDrteHE17pO8FVLA9rNfCK5JZOsmX6tJ4VOBMnHeB05CdiLJZMsIPk2iw7
jU9ujC5F6z+4ZQ7AWrho3mo3JKR4fisgF+I7OD8IriKFUH0OYd5DbsYTh8P0WJGnTx6St3y0u2uu
a8VNO8oaRhvRK6aN/U5ZHv3V94h5nBQ0ojSWGvRuxb/ybZAVX9eyD0Roi8ROEIheUnG36ae2+5bB
UAtj9jQLbfwVIGhy/v55Lc/jNTwSF6mI2/lgdpUGI3WQqwGPTSb7dJXm1cfntQ6IT77MGEj59Cf9
sTqBm0JV1DqQxylc6Iy+iy1tnVZt9RrTl7VUOnCI0fYG3DyAC9vbNbQ/3+Xbi++Q0JBJ71p9DE4i
Q++GKsW1cVlpA1EZI60b5+vdmjZu2wB8PXCyKNx18Qq7w9Zioc2vKqwiXQQcgYzRB0OTm1ojWLXe
dVtHkaHRJzEsQXM1xp8nAUObTjjsIpv4eZIb9Rl1xmkXA3aYVcj80NK0d61kRu8tIPjj9KEKNXX2
YXCqLvdFgk52iF78tJxaZBqr8LW4FwzHNuUB2cZTiNPezai4c6ECcWVE2iAYElHFrk4holHCYKZn
mJT3CdWvyPwFbG5cF/9wKIbzSMuwy2zNZAzQjawH7T47GqvpQ4aPeHXEad9VFWmEvJ8lmSpSvAY3
Sj6x60F2dP/2G/Ejatwxb2xQwDZWRm8i0zlXadpWPNGXFtlY0VH+gppSuPunbqK6pZXf5skawVBs
ET0kY3H+V7Qljav8ucgKWEVFTQsx/pMTqQD2/5cRkddkmZ/2MFQjJpS5VYG13c2fQgjcCFwvcEw7
KayHg0ruNMljxieuFO0Y40camSH++HNsgeEpYrluii2mbsQWLi6ShLjUn74NBEZdNeiC2327WkfJ
IaPkOGNuR+6H7GiNK4mK/9t4DVmoukMxk2sm+LwCbL0adYBUu20gf+7NaAv3y6wxn3qhlhFTpRhW
FVfE2XEfLqwH7iCzXjW93U4stYxiL4UwVX1u2tPXJJXh6lqk4Ncm/MGu6y9Nz14v/8Zu2aXRTDSR
LVKCXlK+wp2uQFCegs70SGY1XTivfcpU9B7ETJf3e/+M/s70nouJk0Hz7QdKdEOUtdfnJgKpTvOA
ar08SwXQQJAPhvmlC6OXAyRXgAJ6Z9V6iHgyeF6YfxkOGotmVLGeeW0p46a0+AMDqnxzYb4o89lB
5pGhQQfuXAhS3ubk0FqR4egOXvTGPU2xpnhpBvr5+/OqOvYNiv2MB8mZISi4bEyH75aLMcqfjxv/
ZVNfPhjy2bc7u9IljUaqkjPvAfHFUy4gjvLaFCasspIcgmGC28jHwqqRluf6OS7mvl3quSNwh/rP
cGhdkZToyGAXxa1NhSev2aQ0UNHLZXpGADy2CpRQug608t2m0pmvrUs+71PvcP9fEwvKlSHz/kso
dv/JkXj8pcYs262ADBJUp2fk53mdGjtqmrVD0zDC1QCMSdcO1SB2cylsBa8SjvFEmpoglQcIfzum
mWL4W10ipua4TCvVYKUmdDGTCutxqdN0xErj8Siv4YP0IYILOEbe2kQl0yh8O7Z3aEUt1aF56eX4
1ZvpZuWnNRI6ZVytGYiYXUMFCVZ8aDa3phBAxLvMc35yGYF8qJLJsFSe9VkDVcCa2CwXBRasz9Cm
Zw1tZhoP1IZEQmQegGQoJ1jkDULGIxWOCHYSuivPA1V6+pvRbgFCrrcUnZ8NJ68PUfUs3UgcZxMN
mKGY5KfTTUqMMb++jBH3iJwOGO3y0KCjl1i39wS4JbriRAHaNcW79DrcEUx7zY5jOiuWxuhJEQQy
DNzhj0QVzTXcCn3e57YkKWybb1iaLNbtAKyVBB3lL+0y0KRd9OnSBEKdp60yFvQD9xwIprSFDI0A
6n4q9rGy7JYRGg7H6fphZBK/Ug9ec7Z+jRqKjAIv8vDqCDF4QZ/wobsQPwYMPX8dOmyo1AK6Gojm
bl8YDFkC+MMcZ42r8mti5vZGiUbrzlwvs2B9ZE9AqKSp1hjP00E+ZAH07KDIaH59R7cQdChcR35M
vY/6GtNaFFKLpCwGlMg+y6seYcWMwVHlfeKTB5/MM2sk3nss0ik8+h1GTtKqAJlQAVyHct+54mkq
JvBm1afnHuEzKwvIwBdtTkr3NHw/z5EuIqxbT5r7YjmpvRxjbLs5fLcILzLBBcjYTwTBM5jo6ofK
ycY0ooV0v5khs82DFpWyGJHnYWgYo09atptHIEr8o4Xv/oAwVeVT6gkcdIvabRvHhHmfRvb5VgO3
nfvKbXiEF80whwx1bNHgpGt68H/D/L3xnJfdrzcqmMnxvSTPAlTSWIyu07pH+A4zWY+d34+Ab995
U8Om2Vwjknb06fvSDQJgy2MMRLXVYx7hrYc+tdlZct+N81TvvQ58v88B1Wgoe5jcqmcKe+VBGl9Q
VaCjU3NuF/mt+ZMc2JpuaAGjsniZYia/2vGOGmy+wc2jwJ8MoN2lXTIFm/JUq90kFmXqvt8WDjNl
Fsc5nBH/cbF6QpFjq0MzV4wjG57UEMC4oXGoSKZgGcxV1rH6sEJ0+kMZogjNhJeuSg9l+GxUKjJ9
hAuS9nH3x42X8QpNDiLHUR7yqmsOo9UhYacD2eVdSg8dJQYSRV4IwU1Y360GX5hO2BU42UFSrK5H
XXuJNwPavaD5oEKfcAMGtibIhv64y+TyiDowjzF/MUkdXVrgJybmNgswIJ518vQLbt8kJRU1pbch
XHt6JrGeeRNH02DXpJVRLnekzTYQvFmvcL9eRhUbHmLDLwX43JDd7pDDkNvmMVElgojjQfdVewM9
XAbtxNkHlj9kuop3+d8LO/ZUfW51QkAhkdyo03Pd5fiuSyxDZ/ru2Xr4Ns5V2oxz+40mCMPNK0E1
fMx0BRDnnIFqHN3lSshs8yEkqhalhdErh8vHUUqtZCqZ9lHicEo6UZx0SgoqvNvXKsRNOQQz5lO6
cAa7og5AD1p7D4fDeQxCm6LlJaPC2OKhx+rg6jZGarJm9CJ5qs9bLKaUuuXiGrzUQxPA+hqPx2Jl
L4Ff9wN/JK/2PvvA0aiTNBvj9P7jwFE6mM+7MIW+W9iMipwk3/0m3GVZQjE8YAzbs5k/gQ4aLuYB
K2b4bd5OlLWK00oI3PxTjQKQEVrOJ3DCsydNPkL9W6Ocu7fIbNgg7snqHngMEW6Mc+3eD4tZLork
FubIUA0XoLY2yCTayTDYAAzjke2odQsOagwAdB8ma5/Q/bf1dFtOD5wi8o4CQAVV4L7FnYxX09m3
n3WXnrUxxonGZVpRewDZEwAnmTGmkJ75tpRrstWPaE/YBUNyPm5c8aGbl/BTzHuUQ7nI9RFw9SvM
crNPKPIbdGBN5AH71wnbEoZ0HCmdpncF2f6j6c7ayMSyGGy8xDp5U4iM/SfFVUIP4wuNkHPsTgts
dhrTEP0S6ZnwzKEATwqc4W4JgugJFx2ijUffjW8jeV70qND+Qf57VytyssQXgzZ+UN4826nsmHbR
lsGmjcMKqw6Uzf9QPU35GD2E0yCMTi6HZfRdkuJAiRAr95ckzxwv5kS0+2Vm4nyV0CXosc6GE75D
lXxF/ZPcYLQqLnl9/HOeZ2YCl884H13OzkycCM4qomQvQN87nbSXFjYgbuD3GOO1cqDKUAGECaDu
LLZeDU0qnz3lTCnV5lKh5GaOp6g5Xb9UNUn3hEqMUblMaifVxfKbB1Z9ik23rfvrEfHSP6BhPUph
NZC5Su3QajXr5W2dSOfaWEcQ+d8Zc+6dxb65lRmks1ySbz5gDGDtCZIB2h6IX1lqVDT5OkyVeFZX
YVZR2An3rEjVrRKJ4d87YnOVoz+7yeRBT/JISs+pKXyAxRQJj0LSgEWkcqhCyCSXVEy6cLXdmv+U
Qj5QH9ujOiYeUCivhT/OTsU2W3KZjTDyxIyRzUSL+MnsOpPkuBASb/4KChQjeH6mTHMzNq0JITKf
poazi2+LQ8bTZoCrWKG4nVR/A1MrCKn5TGdOR6OsQoeeJ9JIKYmDLiXtpZf0KmF9RQh5qv79jezo
EQDXecEgaYtgOshvBbx7zvIqEA2CgBuNQyD558jSJKS88BhD62dfk3JGVG9JUbfckYSvKwgobJz8
e+3drJ80Y5aRkl/kFyLRsN0EDuHnkv8YcljXurudCnwV+mJaOal8yCW8A9BhxPnW1s/fvXFzMhsN
o7fW3zALSdtm9YfMfBVvfRzelEPcNYqUQgm29cti8SHkicBWMoP5Cnkqir/KCgllP2g0v0HQ0S4O
b3cjWjoZaYltTvpp/dQ08rTsDkVfLKkJ4NVyuXr33Coxt96hQur4KFwzOLclhqmOrYOEaZgsz21Z
DZyUkwkWmxFMfSqQIuCEkWICw9xMAv4SN5wU4jY8Oq4Ql2pIPekyaBJazVogyYUbtUSuHwE0DMP8
iokg5Cte7tKsfsWcaIIr3ptajNVnyJX+SZcvztnlLHjObRcEr8/XVXdCl7tRidJcJ0FCZaB65brF
afj4bL0tcodoevw7pn5rg8I3DKdBNtk+yAt1qHW5TAXOS8/fDQDb8RMzyDZkx3E2ihTABj9x75DR
6l8knrLQ1EIfY/i2gwl4G2MiCrKma+F+frsGdtEAQHaclsiYSY/B7TucNaJ+3J5SOZwMgc6dxZVV
fbvSAHmOcjA3G1AhRzHzWKw+V+cGxaufbQ7yGQJJ1Qb3gnFLFibBl0RldrIsHHw2Ef8ULsZ/6Aes
ZRhDrx6/gKFXz9KswReYNdH3ou27OXrE+KkDlFUm872keH7dvua6PCMdrjei3qK5efbCP8uWNAP1
qnBf/xOKMFe167LFmM1jKFJ9b9LRx1ofdn9GH1Ddrx3UHdbwbDMy6cgypfIfyyjD9QzSqpWjYysP
Jrt0a6Dn/R2vMQRcjB+aFZY0S+ehVY/5ngv2WC4R8Nkfqd4yeW2rQ/I1bTh4SoDxGrDSk9j0S55L
q8/fYl/R8FBVl4WoBT9RLefwdlqdhp0J5Oj3GI7G4sAdrDRiY2zud91LHQqMqvHWMpYvZeQPgF62
FdVMWh3LayGV2Y1U2IbGt8fTmUbXPk8KY6nCiHz55SXldy3KZmRg9j4UsCLtoVjF2bz83vKpgdAa
q6IfspOXMA02suO9UCL8Xi/of/xom/cU+mUygb/IKpcSkv4gdylijmiWWMFMIWcHUrQKGwDXnEnr
gFOy5nzO8YP/Qq4WTd7JgnYH3nSto3H7XZyRJCZF9kBh/uUV5HXogGafO/mDNYTyf+1zQ6wZ1SbO
Sr441uwL6oo7gfN7blqU44GeuxTOTLMePeLelB74H+HTO53742wjJZsFs/uoiBXnhae8bIgV7gof
LQdsnz+OaVqUxRblDdxd3GK0TH44wVjcNvxnM4Dts5sCGvGhA3QxJpvFCKKoWgsu9S4GQVGvEjGS
0WTs0O0/a6d7FI+2errK7fF9YxGJmudK1uV9/xuTfXqJpywd2NXBobZjQbkXNh3mcSzEU5p3dQxb
siCueaLcSa1WUgnlrb/q6ZJ8r4BFswtRtp8fI/OsNRWiwrY7CRgIAHbOoZKqkiBxGkxz4dinKC93
NY3oTcYDpD/BCu+cTLhqRNuCYHHMQuRKVNA+yYOnCrpfcNA0Pq3Lnfk8CLS2DNVi1Ot4Ie8tLazp
dQUXWuEDScuR+BEk5SO8cyEq2nAopZLK1hl9KGdSwFpu9IBCSVhE3A08v9GnMrlgdtb4W3jZk2iP
omfYkbm6eHmXiUMWeL9WJvFrPp5cRJDB7lwt1WjaetHlmGnD+9dBsBaui6Gh6ZwFX1lxA1Tzsqe4
0/KawRe+U4CUmi6jZZDMQi88K2Ued1R70Wzs+F1QB19TU0x4d2dYiyRQFtDAhDhZjQGXVL9pVzCe
4TwgLKaIupZoKaiu8puw3gKoGRbGe5M+rA3oWo/tm5KGMSmOr0g3SURljmmnzc0u/3WihkBFmSK5
lJwvpDNeeORg+BN8p7NZ7lVHmDDDbG+1v4+fW6STsdvkzwGe/sj2lKyCeC7aAmG1bQosOK0jDzRb
OKhsWBTpmVJ+CEsgyJTvloNMdI5hO38GuOCp6NPUmz8UH4CMdNJlbQCBcIF9+Vo9FJLQO0IEIwkB
fEY/W2m+b7tlpUilC9ljY9EEovI7KHdC4n0nSr6m4zh2zE2NGWMuHpaIkRkQG17AujgKGl0awbWj
UyP+MJezFshVAvb4ctwPYP5E1W9nqXxiiOHyDoAb4aKsNhKnqTzmAyGcZAv2xiV9TEL2376zMNuJ
MnzhJKSZPWDqOnpUpkTZ9hnhBVU8D59TkgwiDOq6iYqh3ThaplsSK/lORzkTVB8mb4xlgxymgebB
L+X2JACRWTbbG42kZkXp4MOLMVJ9/rCnltPwQE8o702dFaPI4/biGa+OkYCMDmXX9YXdQB8P7UFh
hvEtYz6UjCgl5Kxvle5qcS89A/lOuFVCYSPtmgKSbMRyp16oSh8xrwRRDNUrUqMjHE52J7tiXPQc
TudDtUJxrdMKOsHS2oEQmpEMZfCbq1l5Jj46KC4nPsdmhrXXEtMMLECoVcOn6UvvdFxJFRwvMg2r
aIc8PxD7+g03qyfhIKrV/RKcPPd0nOctRxD24Ce35cJnu7w0o/b1rJvRukO25EpZfwJIrMpkm9nf
IftGhrhrh9AaYKAGFOM9GUcKuAP64YnRzBjuUP8/jDDbHix7f5X3/g+R35V4AH9W0gP9fc4+BPka
CVdup0zm4X3J77D3IO4BltMJLW4ZSVAyDvKGsCPoOW65wNOXv6P3NCsrdZBxGxLmDUa36STIwMta
+P7Xaa8cRnyGkmJy/etHf5TUF5u9+q18Qz0eG2VM6nS/MarGEcT/cGGI5WCbYJHGE7tc3i52/phX
E9ur/Eue1OyopZ8Sotav4Qen7/LAvnZ/6o3nS7dnqljQkO4RUvHWhmughpAEc8aFh9H3tMvFk93l
t4KI5ClbUZJgKI6dvZ8QrbIYaRP7RSNVq4tvD5yyGPKDkg2/BDO0sZ/ogSMgOHhKM1in3BC6p/A5
CUeIFCqnuZj3e25XbscJGX21MRwI5OZgpXSaWV1fZN/lDdmO10bwVOsEDYPOYiZuucZBzXUZxTrO
9zkbadn/lv4Oa1B5rzngqa0NzG8L/M/g3YKDHBiSkGrSca2uqeR+AayXzR9S75pjaku/v74ew7wd
elKdl7LBVfTfsUi0tKOhp/o6B2E2XFZQl4bo7cu3tfnFn1T4F/xKvHqINs/CDE3WFjaujr1QZyBS
HO7hpSqvJyU3o/108gxr5uCrU5zYn7/p1GwtrKKqVs3N+nZ5IXVmUmWzCATt6d2IS9MZqS4Zenoc
4eK0zX1jvr0EH2KIQgx0eVyvI03he8JTuMHyt6InBEPBUacQMlRDTOLEdZjZUFiAl7ODqI5vas3S
xoc64kuOZWInRNxrTB1c264FwwX6r/3EkO4mjE0PrYEPd9MEDN5NJmtspNIb0fI7AjiGU6txgdOZ
wKKJzwSqW0D1xtaoivJP9jHDN75eUVlXU7aKVtLBHjeP8wl0c7euku8sxGBgXjVViJONJdRBAzrh
AvBqWzPlCNeToDivdOg7Q+L6NU9ewtSK7qCIqg7SEtkdixPiyIGbqA/6f8tcSzxoAcjOD2HW85OL
mKZtpMRI/CyMFg4xgD0NoNaoafaoAdX9HDjEWIXf7yuKi4jOY3L6GjkP/aohpEXJszWK+iDC6oLk
671AE0U+1SYbbL0FAPxFuhG/CJ1UArPnw1s5LJBUJJbIWXzIHCMzsBAi++4JFJFaXr3e0btEDeAy
rRi79B7AWk/aRRtL8BLU21fHmsDXxY1aLsgyHLQ8SsxnbJF4u6P1JJLuq+Q7AJDLCKH8Mk1wEtcM
k7JNJslenF/KUK3MUHzHeBrhI4Na5nurz14VG/RRk+lJwciALHKgvXKlDUGOFLSgolCfLDVdGgUC
nfhvmU6EMMOxOUXQWBYjVksS0bf6VnPdlWIFR0cJFJzwKeM1rFgy7OUaMAAbE6HbBT+oPuZUr8o6
qzzPHZE+6ivL+SlZ7o9iqL7elJGqvNAHLfA+jojMGLB76G8098vN0WYLoclCP/dWY4trzuPYvap8
9vfjmDXGTA9nH7X5MiJ57h4ySbiVYCWfzc40oT+FqxI84DED4iaVozJFXHVLSbQ8Am5Dh/rgc7Aa
qp2cGj4uULBljPP+MDKJgAvU+ErPkV3DtjiiihoDpoMcCgdN/NruMnqYk9UghmicEt6xi6tvl2tT
w6D0MT/txR4t+l0nX/xXqosc7XB1u+NWK20dp9DkOQnfag3Gg+NXXJ2jvWrFmRnPHB69Gmh6DNBe
TXtW0hAsq6GS1ipLLORA5dQ8Mf3cptNEin0ACEvbWkyvaNhWKRJzuXM0tOkztudlyLZ2PX/PHqZg
OiEmzrtlEIQbpAoRFgzREfAKBMUu9ME+jSOmfVbWQshRge3+kkE9O8my7bUNHslR3yFphoYIYlLR
+uIXljzprKRmkE1oCe7v+uFTNDy/WXM2wgRd3fr9r5/rY/qUc8IiftbIoQ8p6m66WOqSMCpoPdMv
MBEzFx1niKjKO9tGPMSPLb6PA5lqVVO2e3gq1Mutsh8/ZqLdDq0kYPUG8De4kQieHhI40z7wGsOa
8ZVyyBddkx4IuMJXBZw6jHdQAVjZbQjExOMonJWLNaIH+6ue3bZZKOPfF3/KdJxhGehLaYzVvm1e
97/eD03yO1W/rkFVl5+TI3CATpZvhqR5GdKLyqwwjYnBerIu46UNlR0R80WIfsH0jQK1UEKXUpQ7
ncoDWJF/4BNNeth7W00LfHcSROaI6qjKAtSG6NcyJVW/xWApVgWG3Wx/g+k46uPjE0AaEZyebx0d
aboj6oTEff5vAjMcmFS6abF+AxY+D8c7kB3XogXqse0Ltp3zZqp+/UpDPX+mV1SUPv2mVSGSs/X/
8YFmfOHHxRD9Ws7/RsaQpWdRdmn1ZWlvHP8SHfs60VBrVAyVVQA0Byp7a30Qd/5Gs1W4z4jwwYIJ
+kVghS070YXwA0IhhKQxhVmh/D1xDz607TNNwYA6KOogr/zt9jN6ohZ+e9EPzxKerjJNzzEdZcC5
Jkf2f+B9LeCJccsau4ij1uNwqgsmxjDd62EjxKcHuTvQm6KGI92Jncp3YKFs69PF24BPFe612wTo
tpCnqxTnsw13dxsNGKlRvLgIwWtuwcbHLMFiMg6Rj+xucg0+rUPiZCKt3fbNE+e3WQpq0eyiN44A
D3u0AY8Aq2SASuWRjFCYvYhqoiMpLqYPAM+TsTu5agDcPcFh6HneRLCvrrhgJFgTZk/4uVIS8VDS
WAjHpJZJxur+xfJtx/hscPZTwKSvx9GhxQZPcPjf7yXm+bRS0L7B6FzEyaxoC+WLo9iZx2xMsHH3
9Uo+8NVLLeGptK9ht4jIgGbAtKoXJ/ss16XyMWNFY9V7ZTTfVycZ63aG3ljiiEUKrmYYqskK3bbF
nNj8OaX13RxYyfFrt0+HOblY4NK+StsHENnBZg02BSkRfb2Whvu5VpvCmU0gN3LwCcl83wyW9D7b
hnXdpoiPBmZgRGwI37ILKEZDGxbo+H+LWXQxgTkvkfiQmOctka68KDG/JKje3CQa8Dw63hSyKc8p
a3zicIPixl98++76PYap0j2Gno60tMq0D3hs+b0AMIMW/GIEV4p7P82Y69IFI6jkvDK5TEEbkqoj
28LUam7Hw4/savTBvlQC2TdhRY/Osi+VWxz/50AdSy6wREXkb4kZSJhSsSltvBRwuUvdZR/UrW/5
46izThDVzh+MTtSN4M2CtjedeA+3H5vf3WdhWM6VzNaYDkzVRjTsaV1s5kB9SOAlOd3qHvFR3odk
v7JJmFmy93AlxLy6cGPqHrsiJYelh45Cj0c3Wc9M1uo12jIc+lMIiyKkPFoHOju65LaDrwb7ZX0d
1vexqIg58VgNoVUIeYdFXcjaO0/etnbLfOP1fUtSqXPWKzrOFljK7kYx3JpQmqUBM28dWu92gscD
b3E1iAf/vBNZp/qhHQCSScOuVBjy+JJeP/CuW+YH4cwTYIPVWTWmCgDrs49yKsiCa9OzJix5f2d1
uL2CcgPAjTqOgG5RpZ0oiDu9xT5wiqJiH8q64cYtwRZWZq/YPf6zttrMB2C1ExU+GUdEjHR5pfhj
tmyK90oTJGIWMh/+YFuREo/tpBHU3XGm5H3enDXF/qv+vbsxhbspyIky0R+StJUGaOLSz46qVQxX
9hMSVSoY6AiyVu2U6fVz3Tw4FUfBK1Rx9fkidJJ6QzhjBEJD+5LiLAu9rFrtZ/fsVSpI70mfkZe0
Cm/G0/n0NqUm9M/RqhvLY0Ogt244YQtz1bNPui6zw5nB7gKaLyFhkMmGefTwTDs2wQQ3URzAkF0z
sQtVNaawNqIaX5+K3FUS4l7BD7RDE0eqq0wAiJwLVMN6Litf1ZBb8Bt57jkWZpB3PIQlr51eXGUL
sE4W/9fjCB0OpNxQ8PLs3yDntTcFSQzFYM3MG0yfYi+GD+2yN8AyYaZSsZ2BWS5TvbVojaJzFZhG
VO8au40UhwyVImQr2IhGg1SNdcsCw03Mzrm4NhLpCv2lYdtMOkI3W0jOAplB4C1sM+nIZOyQny8g
wo18FOZXmymmft+H9JdOadOnKTYe+si/VDVAfps+2YYczz9A/re3148rI+mUjzEekYH0yCoMqQ7Y
Z2HqFSlNZiZA1hacXmcoQZDJfv7qh7DTALfEXh27bTOjNnhRT3wMINaEAffI+V6S4Jky5T1UKLCk
7zmla2XWQv3N+R1JCVI+dKWOkDyr3RSof5c/nydYFmnE4znAoddmHUx0Te3NyPmaASSZ8lxhtKE7
LHBwAPLckkUJ9NmY4MSJQ/VwoBYDDOCQtkwVNlJ+J09xo7XiYUwQd6Zqzpno6xKQ1IRDj9u5Qxcx
WQ4HNIQWGIRDwGSLTDoAABXF+YYnG4BRuWlK/C6a8ZzY93Ol5LbinjUtxqbbk3nfgR8Wpmworc7B
jb9Ai92LqQLGpE1LaQSXpkcETeaUh1zrF6KnUl0+4Wr4D0Ktzf9JnybjziY7qyBsMAEdl3zFKumG
W99lFchfR+2bNkPsHIUEURH5ho0JuaOYKWjfR2QEX/YSKZ9qCEOOqGvuGHUtJsHOLTQwZtiUOsIn
PdRhxbF/cXuDmGBLeUpqbvyQPkXJ1QE1D/TgS+46OO0qfWBIhwjbtan7/yzzKVhiN2tqWNX9hdnQ
UHlWkaY5dBCtTZaEpGDj+iyAeDzAolGJFZ+ay1ZpmnVdPbW/kZEHFSpaafi5Rec7GeAKJ2/Q0miZ
Gy7g9GXcP5NU4C1pwMkgNXQlkhH0bMOeNoE5YBpe9sNA9lZwUj9tHq2kX4zovaURgowy/9cfE04j
MkIq9tWyHTvU5KS9ynoxFC0LttQ3rzMfIqe64yDrLdsfiPLS63jDslXtXnmH9EXIvGu3dp8bAZ/X
raebY52VMZxlEMqL7YWtqYt+PzuLA+w1CrQpNfSNQza5tmqwCHo84I787rQSiawlRUfWji38IM5w
G8V5FkagoC10edHZQ6mpZBJUEffiu2mvrJEpW9z/imq2J9ORQGmiXZnGPq+oPxLP8t2C+RC9ebdo
rxc0wuJp3Yx6QeyyBHoKOsGoZxpOkjQ1iphp7WuDYfMOHt/Ufoo2mbsGHgFyUYEgYurebRQNJgXY
iYkenVXZDBcgZSrTNcFdbV5MEX+tLkB/w+kZjAOnyP9Hq/7oGvy1lEL3bOIElGZveLUKOgN8vGPq
i2bajjQbdTkb7nvlITuTF2ztxB6uFxswIqRL+iByRbKMPupsUHl9npjne5+R52Nh8B4DM8LKYXP7
TDS0AQi3/5FpYTqAas67O5G91d9h10eCoz5tt0dF0Q1QLyGb4htN5osPTQB8blrYW1PExyu50OMH
L/up67MYMNNb0RZBS02p/jvpyifOc9le+h8adTd0E8lvzxQ0Sp1lwwQwvbxvd5I+xWMdHQnhcd3e
aMmD+dgFQmOflIrQbwVc1mzsC5EiFTcN8i3iJed8ddyOorCrDSNNorFDs18sJuC/PZs8XHU9E+JE
1Wby4BaTI3V9/WDlH9msg4UqsJbhvOsGv5glLOdas7KLScGwdeg3Fio/g0XjDJMKPzknNOvu02N0
uE7GHjF2h44FGTaqbfJ4HdjAhfV/mI512eJk9u3dfro8AanLCpTrcTSFqkMWu3VDIQl/1W8YMdDB
uGODd0XnbfngGvbGacv1P/p3UiTbnB3R5LlzmxaNs2U25J7yA7ji9/Xd2Sp1YHOHhdOYyv7hFmG2
HFt6HmQxk7pfmK+a8eFqzm3Mn++uHrmbTcsHm1Rf5Ck9YxsipcDPTlmRpjz1yV/j4aV2zgtvhV+p
1HYe/pmEAYIj7EC7vigfdryJxWC32Bz0KRLFs45zyvDliHXHm5P90uaUjrH4xloY7lYGW/6dKcDN
UPQQ1/cJlGA3VRQFrNJw+xHP391aEWIZ7tcApom5heaNdPiXRI6fpFgh+tzfplhbU7PRR7XU7Msu
t+jgWlyD0WBpo+TRoErpzuj5VP3qBNh5VY0q9RHfzqXAXhAQpMLfNmozKX5TDszNk2pHxQMm63ue
yxOqO+EIzsd9fGWpseSATO0NhhOHc8jgXwspfgIOsbReCeAZ2O3ol2yj8f2EBQknESQNJ3lYzttK
9Uhd9JGPBWv2Ob4Pys6cZhG1Yr60PVaSYLabOirzfv1LsiVJrLk6cK2JLCsguyqQAeAewz83ZTL1
zmueGhIlhll6c9vzZ2lHEwFbM2I8Wtu7bIJL/Bjhu8JoXy88zednkjadCoDgAYo5CH5pOPQvhDBy
QTS8vky/zVE62KGH5nPACUtYb7BHfmtLz+iwRSJ648uGqVBndlSxXEPBUU/2HPVZtyXfnBIpEDgU
yf2Z1HNPaHRNjC6PN1QbovWvAeJBd+NELe03M97tXAcgMfj1vjAykOKms9YypuAcUmhy25gxMcZL
by7ioV9U+5ni1WXXi311jmdvVmdRMvMmmDk4vLE9HpmLvZvU8f/lvLtJvnvdEtKA1NSFe0ljb+L+
Z7rgtLMlHPqu8IlAiS7AR6N8KFYGRpN+2te2Cryte+rflXiE8ayvX+OTeedfHwjADVdYuppAmv4d
e1TADDqJbsuI8BF6s44Ng4vPCnkyDLAUD48cP0ljqczsi55Ic4MUqn5FeFYrDuMB0TsiiWlp1ar/
OO3POnc3Ktn6P6HsUuMXXnFJOCbryd1fsDbCGngCgAP+MwB2sydJccu1QnpfExXwkJu8ElboU1gV
2npxstQvqQLBObaxVy3jGGhWLg1SrAnr0aTMtIbhkRmmKi/5kXt5/QXS9XfxFDDUGjvdzg83ovOU
AFoH2T3xz6xJoArL0007+J/W5hOWcNWdq4ReeEOGda5WNuP1T2OuwN3GU/wZvdUJr8c7nNz4xv+r
Aua1ysC4zD7TcPfy5mGzp/XMeBhSRXEhhbLbtFlLPRzHQy+k8LwdVgxjshOwUTqfF06YVg5xF+l0
UxpXI73082JniDehY+BqATLHMhh9FK1SG3N8h+pcgtc3Bn6Pl03WGwXNBo20iGStaw0Dceq2WJsL
JjyZTP70yqYVjRlMYmFek5r+4HZNELJB0U1rvR72OTpe0X24N7IPSCtYlyq+1jiv7QBtu5ORapn3
PW88yyu6SJaw2cAPsQk6jlzpDtn90Jj8GpDNWeLcWdvr6z0N3gDJQzKfz34TYiRqOIKFtf7NYaqw
+3ewn1ldjaMUYiDvpnV2TBiubm/IdILYMtsLfCUwWl/0jnO8FFEP0Tjnkn2eMTE50o0vOrtY+I1J
dcXLKxtPW1WyoJzEfMwJWt/FCg/1e60fZaqevQ+WNTSG7fhqLaX2Sew459C/BxBxnIaHzGoB0gTq
CEBjiU1f+B1Zq4xIqb1O7i8wGleIGtlZbgxZCoY0cE6PthdN7maMBGX0j8SQO9UpfNbZbbweXafd
J1n3Y9So2ECGMy6FjLx/mYvBzbce3thWgArpdYEWhBk1gNbK6GNQZtbiU/BBpBsKyXjwYhYEhngB
zS6Qme7MTwnITK7Alxc/vAzJzE+BKdm7xioRhzuj2WHwQG28Z/3N05fdVX0wiJQc9yYnWx9G5g4Y
H4BEK1M4Sfso/snwBvojKxPDWin3qEZIfczUT/688vVzC+/7U1+uyEqgYf9gwiep+c0sdkzY1bFe
z6WmqjGi/9WbMJIb/VaV+kOYkee4YR4wXFA61n+EisNP1pAqK+7FPrx/Po+f3LYL0dcFwGV0cssz
4lorO0mj11KGH+faG2rjCcZ5hSGhAGjkNFFgdP0OVmtGDhUFxpUL+L2lGtV/kRUky6lKrY6ps8z4
Ys92Lqqa5FDcCHZ2NlCM8hU32FzOafgboINlK57kZKcfc2kEFeOc93yDKwLIh71JUcRZxyptoCl9
FoN3fePwoF9dOcaQItz/NnOH1b1S8GvHiiDljeaLVPE8FeLQ1zmZ8kH7cCNekYzMZwIKhlG4ONeu
AL+myIuxK5V1lmHMI61xRWGFfSfpE9rEnSIVa49DpZQTGM17vesr2ppSjMIIYNrgDaZ8dxqaCdCb
2eCYRgbPMVoMySiBBwpAWXJGEccrXM5S92i7BA0BFsPoxtlM91Dazv+U/Gy9xk5/3M6xgiwlPelQ
9sTnZoZmZ9enJirRtXG+zDNp4CKULqZmAXmp4RAG1Dh86G0joCqCo7MR7n1zJ/C3nwdzqdbMxWko
hIJQXzIigSnmJGqciE/zE+ztMuBm3omRaYXvrcKF1PGodpzN1xt/9AtiqPw+sE4whdtXPZGK+ing
Ln8/sz/K8vecwxGL/8PDxbhkskfPzTxOMbo8jgTob7ujQmVV4Vs8dTz1vJBPcAEz31yx4VNRZaMI
8bfAwQ5O0dpfyRKFSTZRNMQ0eTBskVEahvX5SWf6/yrE9DUJvcxMa5azvSWtJOdp3FITTAA2kB2Z
9VjfxPYlDf218AB2ef77ei4sSwHyDUUBZGWNAsP1hvLM3RmfIXJ7qnZvrutKkyrIquOwIwJTit2U
Y0Vk3puTj9CN94Mu0cQ2TRrfZc3/Nq31JI2JRQdWEDXYK5b0Xa7vgMuGsAj+wkwTLAdp/IsjkY3c
H5SiUCPfgfh7V2Zi8JkFsMDZk0Gomr1dAnSwFOAhrSCqadrWK69nyvi2S/ZvtnYz9pB9H5I3nyri
kPlwgzFUla/FV4Om9GLZUXBsiN4upl1XcbhHzR1cTUez4kgOHyVzGkLlQSdMp8MA1xI9aVMKuQ1x
mLJGEaYLC4Hv+Qp3PF9HWOiaZ8CKDHhqEJEeL3AJkil/eqEeCst96BoNHCRdUALgFtm0ueGLiC5F
UH/rmoQZTd49llcY0r0hZKoX45xHgUfHm4TQDvRXhbvTveJmdpIpQO3FO75rIqk9cnjqzZkVI+gm
ozypBan2IEqqy/5KB5WkToGmM8PJm7o1HFLK1J0kScHPsjSm+LfSpEg5P4Bl+L5ys3qsAToiQhx+
N7PM6IE6XNypEI56j2plxrTSnBuBtCHHd892Cil8yUwl1yeTXriRB799zRiGPo2dwleIOVXBGIFV
A9qsMS1I+TNxY616GAdEQVxgyF3nN3gsASLwveR1gGvIyQha0uQ/76ro/dRLuPugePm5ym3PwXfK
wASRBhAfUB0H0ulU2ER+GwM+O1+eXp5UX838rv8dcj2AXIxUG33YYlE3KTwPLRKyoJSG7oGeXh5W
44L0g2NtrgDwmy/7U51C4vZ5NBh74xl9j0p/1I/EBkIr9RyTNwzSSY/l/G77JxUSL5zsFbfCoY7T
Ar4vz4Q6P4nEWkCNVP87K8A5XksuFl91SpBxi3s85letW/iz6bGQ029DoJnCpkTGud4yCgMl7Pg0
z5wXluTiPhcZJxHqcMCh0vJKTgiF4Vdr+pVDnDH7il8Xb0x83gtvLKO44YE9KbgcEIRMixyMi8i8
ZuJMtdsDLcyrEpo9UQjkLN3zeM2ld21K75dBrk+8yZJU4v1Kat+IqVW4GbTrvAHenIltJcIVJrL5
aeFtZ9OpPk8xhXMhkJontoYNNw3OwtjgPrV40rnWFRk8SntCXAjpKMkWSXeL9TRDSTC9sjPYQ3QF
1bdGoWJdm3QIKCqkGvshx0i8XkzD5qeivNTMi5hgRmVwp7aBU9L1LIHFvHGf72lq6VN/d/vh7CJI
m2BRALvW57Dobb5B8SBCDagns27vfT+XUg2JzvwKl7ybc3LI28vJn5A2duf2tnYuAkWT1+thdBYp
1CpITGylcv6/E59O8oPp9iVv9sUGGK/f77VW/zhGaSl0LrFWiDUiCsbxvMTzg161ap/py791o4g4
TnGnypsxYgBbRxGLQQaW+cf12/UAUU5JBmV8I1yaICw8nK9bG68bfLE0ZH5Flw7ZfMbZmcYHmH67
FQsCF/h1rtIR4cSh5HL71IR/TAIfATOF3KejtQGD9V9BuTeIAbDoHw0pPKmwzcyV/XgGLddRnibi
/+8ub49GtLZ91zPuSDNpwInX4fvjST6lP6kFB3Hx3jlb6TdlDcP01+w/EVDo6pF2CyFJ2gwd3+Nb
aJkzHgUD97iuswamJxfd45G3YqjIvLbpuU3FefqrlgLi8SmOjLioTSyK0vkzQfQpOMLMHIr4dLLE
RXrpIeuLbvni1rTOtPfb0+egaiAr81BwlR3pZO7yPJSbbkp7Zu9IaSaG7CLRsV7Pi00H4CE+i4I7
3D9fYcgh3fqt23MSwqmWg0VdOTAWLEo4RDQZfWKmlM8WOi8osR1ikEYTZnV27r/jMdFEA7g6xSnz
g/iFxko0iOPR7hPcLnqTIyH1YT/q6QAA5o+amqEWKV7Qmu5dTOWzB8d5W2ZD4VMKNyh87zrTWm3z
dsmRnJm6BKuc59i/JNC1VtH4kxnpcg5VTFDwD0dCE96ZQjbiFMWNpdT4nWc2mLvP6BScoylrevu7
x4JvKzvZ3ODfQDZtwNloocX3W1lv0cVNalakEJ1suWmuiYMnKnIHQ85X4Ifl7VbhB5fuVOJ8d+7c
1Y/R7T36193aPTeBtmx5IdxCfiXKphqsZaEYw2zYOviRaNbVuzaFpDJNA+1+nwjutFlR5eyLl3vO
JPEoXGlRucTD8CtMW7C1ovqiff9ocrhrvpEpNNZiXYeBqNQjYhuHY2BPydtx2Cfo2o4edV1aNmWM
6jwl0obeQAYm28QQCwkOaTs47d7umm+oI8BdDw/R5ruk0H/i9zxO09Nl7XTNGHrTXLO2auyOdgyL
tFy9ofjyeP3x1mHABw0kiCYRUy5aYMfs2g8nbQf70BMgWLagjAtepUn64Nn+xAGdFiUZhvND6Qa3
5XuM9STFR4Mb0ipfXE9GMfODf6n9Xqq9mReI1qdivPNZcbDWcvsrX5aVpHlUQWtB5YPBjMZ99DZ6
7pF0xIByM3286RyQvh/S63/Vqk4Ze5cJr1fdaFL0dHK1frMH+GwrUEM6pLN5lq6YYlgeTEq31DWT
36Huc/VCdnmEgGc0Ngs3bBtHgNK6VPYXLkkw1HeahmButgpvc25kc69Rr0jWZk7qjlkoJ2u2+aAC
Y4Q5Qi0KXRHMoGFnG3te/FtomV+PFx9vkVwJuilwKa3VUSWL89eSPnb/R7jGynJaMTKP1J4iFFAd
Ahnalzck8KYB6fr/Xr1BAuZqw2sZ5ZC6b2uZq0vxnbZKecGCJ8S7IJEIlkJQlmDX21I3Tl1PzGKB
4BGW827K1EYtDC91CPjzAEM/9/scXGa8HeywVP7/Mtnpr0yOjJaBo/0vDabxEKzMEWRGOUAOnugB
oVne2WYBBsKUA63kHqci10Gp7SA1+tiLttUzt2WM3DzwAUUDPv7ZaM17n54+9uZ+aXk+2JHe8x2K
SVm9kcBlJiSyTzlxA7M/djDtkRL+a+g5k7vL2/1AQWRCZ7tNx2U/1hBOesw2lXee6yVqpMCcZMw1
STJESFDRIjjlh4vz86fXX1f9MaT7JnxbqtSwalbRcrVhtAcCYFv2b6Ev7juwZzPwTkFAEGA1nD4u
WqZ5sNjob7o7BBqG+Z/sGY8UFRcvUuScTRYvV0PZELxuvYLzyMxmC0VFons2qPMcWbxQK/Of7m9+
9Uhx8wa9CQrXuaKV5KKQslPW/MldnWrx4ZkHRnTwcoTJIa88d1KB2/ZvnwkVeU/Hk00WD6YPHggd
oAxakDXF7m28nmDJP9l0oXQopt+h5EqUjtpQvGcSoVZ5WJlhhs3RZeLpXqnWx8iHFzZmlv6v9kud
Pk2bqgOGIFql21eMHd1uhKGY4Y+BmwZ9H0pMgLt74t6LtYXUmuCiYR0jf64e9YH3jGxesu8Z5qAn
WJG/D7bBkoElhltXA/ILXAMu0Eh0neZg4piNZhf0+s+0PExfztIo/roxy+1uJrIanxZ/V8yRSWIb
Mkyjp3wiEFPsH6Z00g3aO4h+nbppEg4tvu5/iO9z8CZQTlz/Wk+95XSO2atbnnAwNxs8FbSESZPH
Gu/8c9vjvebqdL3L6DZgaVKqR1p8ME8sUkYgnRggqFLigwxMLLnbW19P9ffftxAT/nLyW8xbnhWM
faD6MBIJ4VSdxSJcVGLgfnkMqIAW6+mED7FNJ7eDsC7GDxsnMoRk3b91slnImhlk56khu0jM1pGP
kVD2FCnOUFS4XlxhPyA7EQngX5xaB3HAsB7mfg5t5Iu7pYqqNvBCLmR8/WB5pR7eJawstiDc4cbF
WvdydPo4y54Kba4aE5fwYpUKMhGvvHAQBykVp/sTyAtfsIyKFhRF7TT3Tq8eRqktz9YrjJ2hcqBc
ITeay9h3dYQ5Tx6HdVoMRBgEzRODeKWzRx6UvSSZPt3iFAikR2kHCJpam4GAzQjnWpGLmUa9V+/a
T77P/sSlyO9sZCI0qZ//CwlOMwlB2pU135njTokghjJwvmNdeGjEIwDl38ko/25iW7gCgaw7aPJa
ilj55He/qqOAZ1GOVRbGZ7Ln3jYB+ybizIycixOQRYv/5I2ohy6LGytatzoWJBjB1ArQOzXTHxyZ
PFd05LK1R209GZdIjYw/xxz8BYTxGL+KihpF1mhaamIGinl63kJmyZ+iqQit0f4mGFPsFdDQWaqF
STqHSGnRpvGORf51x8rCtFygbOOvGuL61wxT9z8ykDuuTXNIS3webwo5DgbqHFwGEMod4hlCdrRp
yFLN96fG7Ju9mldYo6qv7gVU0i7dGsHgVXzo+BEjlhB2cNC1Xi/EPBH55hBfYeUmTYqiDBvv746/
fHh5suxQAdYZvPk5idFqY01PVMjn7kkNdVPtTgfggEFnnDTP/AOfB2kaMFP8A3mj7wf0QN12EDmo
QXJ+T+GLeHv5CIviXnU94OcWFAzAsXAv4XGRWEdydI67nL61l8sPtDsVrJ07rDnzXENmAjcvjBgI
Fw2R00hruuhpd8QLSVy6yEXYVrOwMWAAVCVwZo83kiYXbKrhsbuKP+MOAbq4LzcJW1uudjqtrWcy
gsm2UlnXLjcUMsKS2kLa4KJALLCHHwPh5S+aawvaEmjus3WWMjcYdl3c4KPAC9BbX5eocSg25XeM
96AIvQz44xYi7+jHTYteBWQlMo+BWoDKtJaD7dcNCmwmZpm7O8/mOBoe7OLTjoLcxnqiJ82SiUNQ
1Oxiw09LUTmtQGAQ2e4hUM2XjPI/RvL4kIrkiJSQzJnEu0O+2ZCJHP0sxNuBr02jIKuY9sCDWcRz
eAIzhVciU0QIgkPUrs1OJBzYdVh86ZJCe71gpeA5UVIkz7Oqon1msK2IM0KSp0tD7lMTs09F/RYW
qGFlTOyLH/1XqEOYAV49wNbP0H6Bkp4e14fIpjrUquBXI269neYASLiXQ7HaCqOP0wuRm5OXUHIA
wxnkroIIHCKWf5yBk8IF/9mby/3xIyo7emxPUiJZOSBzb2UMVb1ltzPrr9cPK3Y6yclrSXD5k0eu
uYDKyUnG5LV7sLVjC9vZp4zXnZihst1/FlOVMdiEv5PaqVfkJQ5DdGxE+77ioMnk8gTOOMfZUceg
52gzBrKtzXLP6jdylrjhh6cbV5DlwlT62XQNbD1EiE7UBmkoJ15uu6hVtgwjg8VgTfaplwIbBec8
y52zxpsjb8wEmc9ztXSzGmr8ftpIMyt2augjUFHnLrHv9vaz5AFC6EksRqiAUZvQUNqQLnZ9mSog
mlwt9JslRzHABmdxX2bBN1Em2iR+bB8NPF5R91S0S0NjmJpxP1hQKlfr3cSsGMWmV8oqg4oryu9o
TSCSuBPCRC2Q1+jvcCs3aA0Y3C3Je+6L0568MXmXEP2ptAdni6coXMe5BO4lbspK8Ovfn0QTb3Mk
qcLGRkREwSczsHXDIUq8fPMRXc8+xgrX5PpqPCwjLlY3o2ducbvs59Ur8fIVurw2CeKsC2tWPGz7
RqSZn4PcUL7dYzlBI1AgJzZYv2aSNhbeNeqBRBPbMWX8fXOEILWXBYTExKftbuUDMEuNXbLkp/hj
lTQDwCH/+0idZjh8h8sHgECZwPnTpYO+cSTJ34ze0aQHCaeQfVvfQU0B/qUqvsdiSp3iBxhRdrZB
XsLkp2/23oX0tAAQ5kfhoQAsYE070lTHRTMsFra2v5GDQsdxbQGx30LiqABItiM3Jx+rorxWZVmG
9B4HPmzBa3BzJap5Y7iLxK30cotgQrNKapCi97RKvqjuSf/4UZ8PySR792d7+qxlRJVc0CZzTbCW
nzfxuA/sFFtEQEKHGKGfxmX8ys5KjYHRbiEmCYgi1CTmQKLAIEj6QCZC1qa0D1/SLZFY1kbBxZUw
jF2xIkfjiD8uSJE+y0c5IL8GvH12yYdWl55C3qlo4q9w7YiZ4zCZs8cuSJQ0mZpxNfVnx5uRcRzc
WMcksJLOaM7cdc/ToFN0MGeIN8U7CdBqzjP89sKErNYWECajz4yEQqpBJ93LQHb0D8BBW/o0Ep+S
OPfzjbpeteo8MxP455YuFWS5O8+7nkOkyiXlGUCX5JjBL2mbyISEZX4uyyCLufnYFyrRpBz8PM6b
Tf3vntPUpRDJP8Y+G9maOtpy1mKJ+UKX2JZBo0rpIDXG5EjiXzsNuOwlXBarEc1h49IFXd/Y+zkc
a5j0viwiYI25pMbsZky0TUBSQyEuZtTVvJWAlMVJuYSIqMnx8l+2XjCQIMGKsfQBwYLfhK31MVS2
I1xvbf/ppZjVoeKTrdQtHLrmJEp0w9NwH7BbVSl/O2OFqIO6S7WWGFUuxdeaiuMIlvE8qqWvzGBy
iirIrcC/sFoKUyX/nJuRpjKz339J18NMwZ9BcWvBtlXtZQ5KLcaHAEopoVJc/EoQ3PJzaPV3xoVH
UTp6+NVZYheNens2E7ASgBO4kQ6GoGBlY0fe1DjxHq4GCNuOYsywEiGKOEO2wIhAGyzXdaJRU5aY
1jO1ps2PZcU5x/FtgezujsSrv/qKvIhe9nCRHGk58fmTqO9bj/aZyQBfThVQeltZPN95dknk0y/M
HItVOMwJcgySiWHWCXUqQY2Fbgib+LRGFwfc9hKMP3k6kMJNs98Frcot7MtCzXXQvioDHZGcgyRh
j93HpNrTayVYWLl28fzWf2X6Yvk+Xhzh9MsFmDrO4jtTQ29ZyaXm1nSwhlDfqXksOfy6OygkN/OA
AH8oQGL5rFR/p7RLs86zBpf8JKcifdJKNRDFzlTEACzIQi5y4O+7eJYLko8tx1BUPHcZqnl7n3Yx
9Gby90SQRFcn0xgryUDGsdizZrpJES8dKITZHfLGMga/p0vrsKYVA6CjK/ejs4FjMJCQWnZPVKnj
g+RcNqvudILMv4pDvvEaK4Ys/7uOz1sRF8g4rW/luJtdGCIRffplmZbiOZBLzj0Qc7qBn2E3L3Px
s4OBlBw1BPq1m9ir1nlSKyqyGpYgCijRTGUsGuGPk8paDbbwFrIgzcOcWKtKCETKCtqsEHWj18kl
4X1OdWTz59Zutg7eChswnIkwk22+fcbhHR26sjyV0uqit0iQA52quG5CSoqVENuR50WqA5QfO7JD
JeulVWclWLTwbhY2yR4Hern8kR08w7dF1IWADVYzmgCdSQVuTEla1itEFEeZABWVb3d2d9EqbUmq
ZNjtLo8e+iIP4h2C+1VwtS9+DTz/M9cXwqDJiHev0JQ/tqW5ixiqOYFIYeshamMXleOGXxtMzRk7
5gpBNgtfQ94MydlE2oLeI2wRq5cHa4aaDgydPlZwopPZRK/LoBsoADUjLjTHGnnmOhmehmSX6Ps1
5qqj0jT/EGZViBW+YuIxSLsFb29Ujn42KF7o39WQx6FLGDzFDQq6O5qbnCeXGEe5udN5gB7hRJeH
4C6Y6g14A5rbIMbr6z3/fzNa/Tm+VRMi1ABlQouwhHtP4Z7o4WIa0+i9p8w5Ddx+GgOUgIlgGr0E
AUUIaZQVumtMVapcfE4bOlmSg9xXvYerYt9oc0pT4F944k1o1zkXVAzbjV5kr6wgPFRgSw32/Yf4
mVsp4Q8Qn7znGPe3BdAqV0mJepkwibEoRC0a+UcmgEHfs547DNIp5RPiE0zVL3CByZJB3oUhNzqj
zVfSqk3JMZ90liXPqAd+8teTLvu0BpnQgqkpzs7av+T/o2i/tOaKzRzH4irAvN/nGgRNpyvD8fpn
v+6lErUAEV+P1RUMm3BKqjyPqSIsF2D+u+t54l4d6nV4OCGvoI9YSxz7n+jasmlDoOCjeFRZxdJp
P08sDrk+5Q1lS9gDYOaYos054+qRvPdzso+xpPMWFe9YKSoHlnGs9UuUsuy44lwfV1Kcxkyv2wpp
/J9VLGVl9QFVjSewo8vzV4D3vQaBFWM88zokjyPongEiWUbXDcvJSWnb/cwgcaKR4BCFDkP5tYrp
wfGm5pTMIepEtGRqH2DlUUkbCaZXHyW0m7pWUZv+agsEawlkEV+/2nPy8eRSbX2niChCQbymE/12
B0AHyGszfywjj0giPqhHIie/FOmiEibpDkNrI62DyfkIlKneYd8+55FRSIQEEFuprciyhqXt+0b1
JEr1ZieKsAiz64kIcKfTVVNMhK6hFvC+QXsUX/5cYFJwhvIrC4RU+G3Fijazvy+/GR1XJtOw03mb
GVf3Fa4FlFIbtEAhnS8j+0sSbfyw9r7cJj4EnJ4xLVNGtT05cGZuUadYsqPUH+DOOrV4lVSIM6Mb
8NmqbnWxnuGI+RMRrHcJcojas7i1QBnGnD286xUUHxmw4fpMrcHGsc99YggRXe0L6DQKSqsM7t7M
9+PWqkoE4NO9Gzws5iZ/Ju+fRCPIz1WhxShH1pTfmZSKSERBOmyhcNZMLqObdyLbkl98wM4W4Jp1
zV7kilJf6uNNsN+m8ExgHuSTVFNikPkTF4LIJKu9mXi2SmXE8P4GBdlYme3rl1pnMcIHgHG41sb4
w7WVXJzG3FXRlO2LDLJH3myIyZvHZ5MLSEAnozISUcbsNr4BYCqsiR+cZHgOX8DwUN8BdgHmCzQB
qLyKQ50uCUEIPIEwuiVjpvqCKMzqMpskG+cTeAOkFxwbAYXmmr2bAF10V9q+37ad9XSOVqw4wddo
uVf7Sgrnyg7w/K/HPypyq0+RC68d5i2SVSQlfvszVT8XP0JWUYNsVWI3TQjyZ1dVq56LHFYwdM/x
I1AA8kSIzsmbDdBvYC4PGghPbX3kcfMOmZusDzl7cjx0tBELvkIcOMXWky5ccsirUGGMbDjXEoPF
nLJv6R5uZcpvblssqZrw/F+bklGtKutI81+P3G68PopKm5auBw/66DUHHzoIzaeEPcmYAkCmC0Vo
NNITeWImgDscboqrpoDYqOV9QOyqN4mUNK77XZXBx2KpsFWcnXivdG31yT804N2hrMNhaT9R6tJK
M0cFPmDhK9XC4Wz1xkitWRoXEShrGEgJ521IgX0vtyq/2Ms+EtwJf4QtOSkhWTYs1EFcpGhV4drz
xCO342t6AHNNKmJvRWVd0VER5+foXoFzaidhQodESyORzuK1+nxvfNsmUpNM0o+wcAnfm/zwESLm
50un3Hepn9xW+OtL82mAVdhYaV6dx0z9XNFKp0W26NaJclC4xWG8DkesZfX0PnMoq6RDkJtV4D+T
XBaEuEC6ptBxXLPUqFJaZNZCJJC+iZ42AFIwxueBAcICfEOG8Hgz8e4MBHC15ooCKWWlO4gMrNoS
wCraLC4YzFMmdS0k8/yVBk3dOa1YFbFrdXIXHHso8pGShsakEsXjh9QwNc/QMB3f2cBTYlIIR3e6
4zHluVfvn9n4aaJJjpt3yphBHQryRUJrVBtg2Q3ahwkwl25ofgD7oMcUYIaeQGs0ONy9omEw6SGT
r3Y1KkHMgv7wDx8zmkXIz4ESQRW6NQUBtFTWZgNfaFSClY0umd1g4e/AUIsa5uWdzLDBBLrTqEXj
63b9cqMssa1ATY2uZ9l0i7dy4s6EyjEKFs9pf+Wnuf/u7+HR3hs3vgyymTVNsSlkjUHO7XJSZXnD
OkrgkY5EoztX4Dym7zyCXbKw7O7pmBj0n6yql0qZW3bFiiMeot0PtlJ5+T6GX16fPBRuqA4iZ5fK
X5TY0Zb0TBG5ruL1wsfTHvBp2+BLvwsQoE1iaW8tzCiKQQRn/YV0lnvg/9c+kO4Fwekae6/Y1kcF
Y7HKsR1y7Ny2rgpaGr/+NtGUkwdbiXPFmZmVoysHEheyH1Hfg2Uy+dQkKdZ1hDnoOTsd4Jq0HwqO
GVyy5jUbtvUaTuN/A+cfABlltp8QMuu/R0L/g615EICXv2BkYZb7s3L0//a112E6IzLH03W5J/Z/
qMtNqvvlUI75aNj5IGUYQ5mFi8+sKyU6SWoKOfFGsp+r9hTcFUjKqQlbvn2N8Ch5wUriVVdGQe+r
kShPDGOIpz9meqPy9GvtLQhon9Ho728Ec/EAVgV9NFUzFhEZyuLRv/mTV75jldMQ+XzcvJYCFeX1
xE75vqFnapV4JgHwY6AjhdLQsofR5YJhd62MeMTW464zDb2M0FwsXt9/gIeqwDcQHhVTc+YMwyri
c6AiaTp93GbtEXojn1y4wy+sU5G293dcGkxrDRsXaYdVnAC2ahAp6MGmX65RaOZ3BhmT7FKw6o+A
/0mL2gzQ81ELJbTbQmu/tenkK3te3WGqo6kRqzZLhPYWY409ngnABrWz82SfQMd06jec0Q6O7Qo0
E1W0HbGwYTzVaz1CnhHGPyJ4zY/tO/SfkAyVVCn2idL1Xh2JAYTj9Ke+qVayCdqaliiGZAIRERsa
IdOYSund21skLbFsOHQ+5LYjb2QKvjuzI60GS4a5VaGe2QsVhPM8XVOh7yVTcge3vaqGPfWmzD1E
8Ock3LqyCEIASv9R00mmvtdXbTn9c8+A6Cmn1w8kaO/wYph8iEQDL00w9ZZFNeVXy9svmAljzSJ1
J0MtkATjhRtmU7DnboO1DCGQH/zMroPJ1M+0mOvstSmGa1jIM8+8CVJo3Pn5LG+iNNoUw78Rjys1
n/P9jI6pnXIiLN+SH1Wh28nQpKLDylyKWgRN2xVKQxtL9ZvYjQo0T8CBIOUkBZob2ReHt8VZa/I0
77kyQE8EVrf+Lb97buaP/zbLtf+eZb6tLAynZyzuWqqC8bM/aOYULYhbPhb/kCZHcnGYAjzHk9KP
K41EZB1aHqmuhOFYNjv6iO4TpYSJ0zDSjfVDg4dJLLU9Ru4ZPPYgwptguzE15um6F5wkKLU7xttY
jhu8nBcD1ARYTkP6lY5SOwqHceZvl3lpcT8Q7z/7aI/nmqNKvgMbo0bBprSX72NexRLNvBpFkWEq
1OB+oG6ZJSySVmOVK2/CEyWE0xIZJejTXzw8QK7aGbBSruC9+QY7xQj9ic7pFMGg7ggGjnO08pfA
vNcSmJhXp5e/ikM5f44bM/VRwXMQTf/BIMdfWH9Wf2cnxDL5is4lDNc0huDeNNQDNR+bYZgdEsVI
B9116HTnNgCNXKC3CzWxQC2wMQ4ZUpF452hzu3et9/rjUhz5qX9yusbLGayh61cIXwqgfQ+/c42Q
GFOCxF5EQwI96nPNoyqE7bReGduIGK2WB6xgz72pzJ0NMZMlLRq15FCth5PWjKCgi1gaVDt6yEc+
aPAXbE+q+LSCg+mWHl525W0+wUm9m2MK5p4balaS6C0DOpooCs1+XozpgVDe7nizIllMg08N0x5G
08hsSPAo0aEHE3IjKRbyKf3e1gfFUhLsGdAuvCjwB0Usu1THrZsIbM9m3UzBG6yUyqwhIaE2R2GL
bu7MRRV0AwlJhoyaF1R2pxjxFLlnQswjyOAvlsqIGcafHFd5pFWQOgZKi2MWCcFPKFWmr5IP6z19
n1IEVriUkwAvbC2z2YJbQFHO/btjXSFqMT/6YaX4z4Yp65pN46d1srAsBaJzBMV2Xq4ftcsBSA3B
TG+jR3XbQb+JBVwdY2zozHCweyt7/D/ibNa0sRoo/tFB7+WTjzYXN9oABmOtmgkL7nsrkqiMPxMg
9gl4Mf7boiNy71YF3g9ladjhN/ucPicA5QMtOEnMm5EOXP69fq29BlPojJIxBVrOadK3ZXV7n+s6
Veq9VZQ7bM/MJeKXKM2sjtlRXO4LvI8xBa1xk5LBGSkZxHnDVJQ8KEAknX1xXud4gMuiaFMRvLkg
kzK2G+wiBA3FXvolx42k1JadT9jTh3nK+8N0k3Yr4bZg6nLW99FAL3Pv6WKGG7nZVsW91dRxy/Wh
5vzf/TDjNK/Nwf7UA4rLfbeTuynBaj5c3TrSWhWksDrfLg5F3yxPXtKTHrZTYcx4WRI9+7TaaXge
GhYojY/j9VAwSYQlpB6FnW7bVN6ZWoSJHAVpyvNOix+nx/vd+Dyqh7QWa6OayQelaeXQgMZYmLRG
ngtMlJS4fGxw+CU/gbZC8B11Wi5RF6WkD5u8/65ZkIMZNuHRoX7HwHZ5yjgBYuuaYuMZSXGlvBVS
RsElbX//3w0vk+NALenAkqbaxxa+k1FvkthXDtDN7X4Qi/ne3QrAkxaYenwSAZddiORXkj9uWsFT
msErZ8qKH1hGV6vTbuuLjZ5DopRrTr51Vy4gxLk3Z5/Vyjzxy72xhbqFHwS1MNMrC1sfnEdoNXIC
05B/U0oSZpPX4t8NFsiAGZYY70lrH6d17/sMqlwqbkQVJx1If9Liz+I442HS440pe8/wzdzUZt6f
kd2B8X81Mk110IssHjucnGG08tGSHGpFcRGT4YYroBysIP37BFoKCbYRipsvZX2Ia4xDodmUD0rf
KUsqjls7bmWjCpceIH8/x4XE1mrIfRQGfcyCPIlLZCsbxnthFKblYDX2dQnAjO6N6aWYVrPePlkY
UAX53kj3pGEiW4+ZwXevMMLay8Hw4CQe1powPrViZ1LSkCWwmoR6aXyz4dZGFo3t7T9QiI4r9Sfp
Bp5GCmWldfD4sp4QHJ0TjZK3uY6vm6uGbGn5sD3J9N+1YA3o5SpfPEZ/vV7YlHD1BFmxuoVuOnkN
A5v/kM1YP1JoEvLRtbugwFK1Pu/LknDGaqq7/Vkq2A0KkM6k31zeePTtig/LwIgBZXv9SITJXNop
DUjAYTG4hczk3xzQa1gCXbgXqPNsHh5YDTvoMPAZCwcURgIdQQ986lmlvjdgjtmla3jUF1exD3zi
Gx23WnVOWyGoc8dh1t4225XP2bf9i179ji0KKKyOYvDAHbA6jGlybleNtsVByxQfYt7For2Y5S1J
cJWIM09i5yOdSTsmVcO1H6buPCyhMVOpgw1NHFOuTd/PiNVDNVbvyGYTWZqwMVsMocMbzKYBBUjh
QuC9E2ZTisVr/6+rXL7hzxxpo8P3blGgEL0p/CSVcqx05BXNDFExUTSVjLMT87Z+xuWwJabW3VIT
06pe07qVWl6bWjahKAShs9Ls5rdBBFk6NTJ/go1NvQNCpLBRFOrQ6cU0yVnaRWgKrYMgt+RxioZl
eck3hmIn2uUsMW/1lD3OaLLh4Lk0vagS4FTrUIEyBpegzAT8hIY4OQ1n3LhexVPT/wqH4uhiyrx1
f8+QLSun9QKV0vHvPWMZtJJ092h/5jq807et9sN4sJ3Dnqh7lygc5kn2/PdTSyGX2HCP92jzzWV7
UoMjzHMgcDkkHYelA9afMGcMnIVT1WOd0SkiZWCY/NSRiEfcPA8JVGMlygZ4K+uiZzz5TbL/iU2G
cPP6tEfA/XlHEg1NkXNvyiufPfWk+63sN81sSEswWyXvgvBjDLry4TF5UmNJmHxmV+Tro+Bns8Li
/29c2NH9Fyig9uZrc85KWPJVHf+lD7B8acWhId2AZ6eVnkQVMaLGcxR67+MBXjCMm8wYKlBUyHwB
bAc49K6Rz0AyMfZRNrhBAzGwnoYwRMH67QjuMQH7vCMW+hhQGZmHM1+jYqgVApkNNPExV1yMcRu0
/uqO5/VHfVG5WXwMikzGjPQQXigqcaAYC7765lYiec5ebHJBngu1iSBAX0iNCYsW00uWXpn4ks4Q
0F3nLXEw+zC3QIACG2NYz7ghRO80N5W2CNK8xyQP4EVgxTknGPBNDi/+/Uok/RjPJl+oPf60aIEi
yzdhX5pZ7A1WOKo6tXVFS/nd7MqLyaCht5LAuGpAnkNmOQmccrgOUV3t3w8DStoL3oksC7lF6Cam
fH3GLjzSg3XQ5repNwG02PwSmTMlFeL+R8rWyxmdvBe+q1Hi1RkA3SrhPEAp/ZEp7+rq5VvQqjrP
edNMcfNPDAYOLPjHiXKazCpW++SIvKstFex50eY40cvEhdZfc+fksp1lJVi7kWCmNYJSUKsWdNkL
cG02dpEIQ8OH2A4UJxXzDQCZyj7fPR3yTyqCo3gcD4eQoZlhHm9/wFgogylOeSCBUufDhh8Y1xEf
eKE0bbJ9P36vpN4cwtp2vY6KOiPDPuAZGV8r2RPtjh/OtxuVKTRWP2L3ejMAD0AgYcRxFYy00gpw
r+WhYMujKuO6PSBgK+1TGdg3CYRVCWKvVdiJo7zb6ro8j8m63klVGop+iCb6v29g3R1JNhWS5DFO
JTMf8vZT9RoWRJz3DWOXXXZBoRIq3kvGLtU+JO8297Mn2JEqW1l11cogVwmbhZ3CtZA4bE4TwicR
Ahce65wWuMfD7N2bYSyAZQ9b54H/8/b0fk051fFr0WScmm1cIKqET6TR+bpN4XlFS1yLcgGue7YC
rQ+iQah8Lg9Kp6/CZGEoKOts5psmMje88HV3+YbxZ2exx8ykFn4Ln9VOgvovUcGLhFjjvXRvowsQ
IHSzZvzkomO/wwWBOo6U+BaPby/CEmhPvBe2GIgy+hG+A2T3SDML4cLVgbwD9ruAqZ+lH234ih+0
JzbvIOc9o5GBw4GBJ3wSxLTRbITxmSvTo6uWh6QK+7jPRIdlB4yzf/8JdlhgdaUhJh7bGsi9Lobw
E6i1WVxyGdqNNSdW3Eko3L+mxlz9fsaoNTyio4M7Vzgp9LhFcT4pyqyPXtNVj/fkvIFwQL9EgXib
/Vixrj1EATdg0JaXEkjxUhdyk3/kmTAvasB50NgDEDcbdMNAVj37vZ4baWy5hUYTLJT3YZ3b26Q5
WPbBZk+PLlLq2SeVXw9rvTnbh8uxpCHDKxibTWImjM6MaPwNDBYm/K5ME7bXxKhPpnsae55Jk3Q+
IHaF0YcC28T4FQzQoMEtldFneb1NEvi1KGp++4yb3/jcDaMGYiAU4oEqCuwlRS6cXqg3V4vb7zlx
LtaST0rNDkYPOwBKc2I8MzvgH50j/km501N3A10fgfkEhpTyKy29D3oez7kB/Ky1hwuelEJlp3nS
+aM78s4uzvVFUD1kA+2jMfRpdipWiQ+//hULQfz8RQGCV+fBB6JKTGdumKVnmMCqSyOdk/QNNR9V
L5YO5iL5Wh6Bc5yjY9kGVP2+IjPfZ/mGtMmz71LLH7Dm7qzuvYU6zJNv1GUTFF0FP9NTo6mMOR9N
RGmdNGCC4YOiRwdQG/tX6e+/4uhm9EC5Qc5W06aSRouh8I7W7KpqG/kMcVSJ/V0Y+SwxxkFHAuTu
uPqwdeBg/voN77s92XPNym5ME9eFo2iEkCnhaQSTj9Ep2g4BgpcKlJnuiR7UvRc4IkUNkqH8S+dV
1p6eW+TkcE2BZelOkmCHKKkbO933MOJKfvb/t4XAkFXccDT+uOt8b2gv3uCN0nifqybYIsoVvy0q
WGF3iVrfEcI8JcBXKRsCNc6V4U719L+v7SCze41qv5BlzgE3ZjH4Z7AtMxTGD8ABMz9A5dWg3CXP
3Yplq9BK0Qzm7Bxo3lA4P1/yY9n6QrVAb+kX1znA6Qx/95072AbvCVa/Kgw4Dux+OicZI/ncNgpU
s8hxrtoIQNv2n/BvaFMxYmZwUnJTzPivGccvMz5gWpi5AtImOfdCH3v4B3IS1NmO2v2fU3G2a2yj
Nnd8dy3tuoN/w4m16OX58mrtnfbxgnsq4tiWYYObyVTIG89PgI5hTs4Vm/Z8teNo5oL0etzp+a9A
kV7UCK23T4CVyI4cff1KIu7qZOTa7zIk+Dcj6Gb6cjFc7S6bBOqtpeyRDuMdFkoFxCVtvJSeKIaP
xdFeXujLlUdA+A8u6dLcYMWG5UfAybhqwttopt0QjR89ZZfjeiF+llH9EcSHZEeNMyec+0dLHSak
Ebp28CgmaU0Jyn9jWRAoaXbUDNN0gT2WivVvtva2i3N3M9BPNAlDJ4fqHmCQ1GEuNkAV5HOG/Ej+
fL6FSDDICEPXsVcaYSd8eJrWJD4182uGEO5vInPA9najMUmWGzRruuWcqk0z9yWwNHUZqPgIX1BA
lShD5dN725O9b2tTiJx1p9Wqoem4833pmIXQazXHMuZma0U7hJg7myi105B2LNC+utWNdZnlu6mO
XATZMDst3gkY/gjEtf+pd2I0gmNoQA7/LBpjYendTiMaW3Vyl/M46i9gRUMNsJ5POvE9d50S97kL
OExyY0ClUNp/WQlacZy354FYvxAi8GM9vQCzR9+OVSDg1ZQueTjMNjXlFL2H/PpkolH40DdgXjM2
miMAKoDr7FQq10ABMQ7kh5jjxK+ifWAC5MnIOU35wda4pUMxAeRGzMTpo8+MQiBCZSMfqcDLRkVW
SOTGxm4EVhC/qn2FbRGlqixoiIA8OxOK5GCrlkQsd/3xRQbuJmqBLSO9b6CZs1xwh+c1JuIqz9kC
DbsNfPSvRBrwLjSgnUrLryOu9sXGHdbAOg6yPBBDE4UQyebv3M8uGejNXqfouWAKUx+rDR9rNAXx
5yqG5/io7YBaSSUlUMQAUjAY2XTnBDOIZNm1S+0YaaTK5SBOp+m4/NkrvDcnnl0m8Y5VCQh9Z0rz
7uxK67YcXxT1RaUDDymwuYa2LO2fdYJ/y7fUwYKy8nZ/QyplvGfKdMGRWjxuzu/Br3XqDYo83n1/
2Yqe/y/fNUxwouwkQwc2vVT1SI905US4xGbFoN5vbzVRjkG2BTul+ML1rIqS4ANWB2YJRJm2YvCM
4Xn+3IO3jf8B6MZdkfsRDVPKdgYY5aRqSLRPZFVNwMOlb66qaf6EA2VF+Roi2d6Tzmkx/wcVS3nG
8NNJFwOc6toZsd302CDWDORHFQfIp6zqatCAPkHA63b4sg/BFQBykz0j0vFK/6iYPVXMjVNC0JWJ
oN8SbR2QZopnOQP7cyqHZCrEpOzwLYtMfUIstw3Pt5IqATR732kfah8/ZhVHufP+9mbeQjXJ19q7
ptQQtFlHf1pF38gu2akpjI8tvSvfh4PvHrNnC1yhe/ZOwkFwRsZ6sKX0uBh+3RWS7+qUqrlHsXx4
owow9fucQgdtkfqB94RNrFP0iUgp0xCLD8i+2L8N05rah4h7ZZ/NtVKiip4QarseMKZRguux6qFd
PIw9xcbbzjVjrbNDqeDJlnjK4cdqakhWt42R7DfMXI09iVfMNtunoc+sT8fzDpwgsuhajNI+by/2
C1XjdjLUzHlrgWD73zj80xIunZj28/31vlLY43Y//wHf4Oh9vPVQSjt0T8AzNc64eVnL8wM+FB3J
8wASZhWS5iQ72Y7ny4KVv2Bszo8OUdnuC/H3xI2dnMTbuM0TSML1o17K/sFafEFm6tSRtideHNu6
sQNw4a0CXzG+hsGnmrmytZcFCPB77FhQZTH0R5VciaCpes87YTxxhcC82ine4PWKWZbtGfDJvd1u
fB6hkK71G7orGVhmIQudXvZLpcHikIbrWvlLKRg3lB46d2wsfjH8b0mpUBc0DqdQ82kzTVJ59A8h
ll1s8dK7V59ywS+wK8eyO12A/gJuW6ficfxfJlrabT5x0a7LuTJe51M4DGAXsyAP/Bu1NljDoQSW
q1E42no+k7H0KbNcxZSHuklkMqOzcEqHKwGE6cHWl3tflOyrpaEdhwR/A6AYCWMNK5uQi1EeN9tF
ieSGOklu3wBAAazKXdROvH9T2HZP5mYoSG7/RN1Ho56tsuKexTVtTO0WuBS61oOjuMLuNqbhl1vJ
2DOk80MvwI60nw+pUrYj90ETHSZAEatLuguh2UAT+LMXwR8RyQ6/OkqwF4UdxPKelx990tRH+UyY
FBXYAuOpwjs6gmXFVGoUudW/9i+7QieCwcuvzTPnFzyYOp08bAx2omlb0J/7Q53sE4aAPj/SeWLN
kPwaWnQ8JpzYIn7xy91uvRVtb/7zE5/FOpszVgUTQAD6Znkw/+4kIz46L6oLqcm2PdFxQOPigaAB
OGnmTzSm67vFliNgPxoESUGNqFMoyslMA7H7+G798UCNEeHUY6LoCr+9x+J4X+nJzwUjp/aseTQD
GBE8/A33eXGv2tE5BDfO8ExO9bP/IsnC9bj6u96Sa6LeDf87Pskd8EVvxKrexihTa4QIs6Auf2Mv
pScU9/lywjwI7uu3S9PT0+EBiH5Mxo55w+QWD3OwE1u88ev5uAGaCI1kUg0zJpO9vMC8a0IpNis8
e7D/qxpCzk1c8Bl1mKiej1ULCJprZ9vVPrdnqWziNtRw1+4S3tno1wQEhWBswHT4d0U+vFC1J7X2
1zMCZgt3MlhuQ2vYddi1X+QRpYee2SqHNUSErguWwXzaK8z3AKeBX8jd+qnXP2NLY41kQmLIg+uw
toBkEPH0rnLrxet/nAEbYvnW9LW5u6z+yqHmG9NvOQCRy4gPCz2FjbKbtWOQEVQO3OXN5eIjgvYM
5v8w2tTrh+sAGCMRGgOvV5GzIYA9BuLPoxGCspH7VW7zrSIb9W+3Wd3VCFfeOerutRlcrFpr9KxP
HNuHwvZ+uhXeJnVmU219DfO1AFzH8cPsdhbmVPbGizMxCKqwhtc7GxHBMxMnMe8r+pNOrBfRqDIz
VP3vUyXZso3s6HbedjEHdrD01i2yny51hWwIUoXEPpbp7mhWK7SGD1vFKeKTrMM4GVYQVuxs50Qd
AeI+bwD6RbYFfc24tIcm30EXx8NbLI4A9EqbLKu43lq/JCuF90ix2v+PD1yf6TwXsAkGGX8B8pXG
ANWjGp/ex50VCl/gmvW7Om9bVLjbAEQ1xY/Fh1T5QBfA2uPM+xnZ8RjfiGylr8e/s9OCZyWJMXo2
FInzxm/W3QEjg87fo8rgjN1RX7QqnUQtc7xcQD4X9YGzd0OFJFuM6eiptM6ZKTyTSlzs2vVxV4k8
y7PnU+O5Q0P8sxWLfBa/kn3HO7GR8Ilw4f9jFpYhCjG46Si5vY2VlT5Wj1WcNf9rJNmE9UCd4sTu
Qah5R+xl718zGgiqOYhQxRMMikj4WtL2QR01P0pebmPQKjD5R1Dkbytk3VRBxzeCdAi5P3QDKwbv
qiWrV0AHAYPnUTtQ+JFeAhl3Tyw3rMNXCTzt8E8WcQc1byxup1qPjDTBueELHDbpojt7jvSvU7ob
FAXJWfMQpGnsbXsb9x6SsZmiiOAEZnVmu3L+j2VtU7fVjsCEFJbAt0wmmUbQczXz9c4eRdcSkcM4
LSIGMpZBSkRTwAaWZHr1LGPBOfQCENkDDavHHQ1TcGtbNZ+vqsxlMGkDTsWs2wv9DfACcvyvFhBU
22A3kiKjNIH0s/22qFWAFRl/Mb3w5iRPSNC2CWiojJN3SNvigW6i/tiqKm4XqXxkNZ8qHCRPItPD
8uypWA9MDLLDk8Zv9gVKTKTY5Cb1/BodLpo+vCLut0n6OcfKdYSsJ/PNdGydw7tJe50BWZ7ArhIl
RCws+Ocj1bQGWlX2asCsda5gLHs7Lbe20IH2L08lzOLtrH/r1CJDh8NdPaRpTohfwr8D2HzfEvr1
j5CeU9KHe/IGdPXomkYBHfMyxCWwtg9fuPZB+bAraOS9LAij6wMJjBcx1PLNADbC8VI5pfa74eAX
C1q7CIsni0Pf2OnoLWGAVh6AUUsoxixGAKVAga5Zcjc7Wu7f6PVB1OW9rgR6ms6eCMZoD7GroI+u
3wzsLgvZlS7KuKHVfHFq1nroPF6yMAIEuer32uQzUf+vuVMKQbrwb9+fyVpJMIsgLU5HCcSNMXgM
l7Q8YDswNamnc90Q1cVUzAZH18aPV/fqlqTmAkjOO3wcJ5qjw+eRwzrmKjt4bWu4hw+8laZe+dad
m/lM3Omzm7BGjl5Aqcic0kXWFzyAT3RFXCzSmeLyTIkOcgUrpMvsPLs0PObqQi/qnHK2bLk/3s10
ItC6cXQmVkVaDDmQZ1TNTurFM0H3GBpCLbaPsIHuqyH1AoP/pPdNAGcLZx5goSDOjY4CxE4NnYdd
nRRBhsv4awIghkwNrS7VM3RGM7VOdU3qN9P6WULgyficlQHByDU3fUW4LANpxJVhlvVib+ViE3QY
ZTCsCi8wqaoX0FNcMoEPSZXnlP5CPy4AC+CpKR/Nbnn9t60JVoMD9PHmIAyXsXmTYpvf8epi1erP
tSEJAl2oFcnlJ+NwwIyDZu6OHW5LS7P9Q9BamV2zRlkeaxsubtlsYQuLZw2G9QZMcPKB8QgGAi08
IFgf5F3iNV9yotP5Fhj0Y4qAm31gSKPZTfr0GlNZ0nBz5f3Fm7Ofb6xo7q8hdy48myNNzQZlsmMO
OKZ4OTYNfqI0l65Y1zxAWGDg3mrB4BAvUwAdGFs2lmjdqcfQn/tG7LMPvOSwtjKozElYCJgQvtSh
XeLKlhyUM5qdgGbHHKVPgHBrRuA/Hbg70rq16iNIT3DsxivLYfsjUxCRBMfRLaNzr1/OuEtYJ8Ec
qGz23VgyY+S5P6wLEWvoFdkOcGWizZg8rFgdfQCwTBMg2FR4BesorAT6yfV3tXJaCiq+XzWBtYd6
7b6wIVFT/8ardEFQYFkbyAtBgqepvFy1KhSnf+Yd6GVeasGnxlOEGhPiCOOMKQSdOxi4PpOtAPja
naweK9uLpalgcr5RMJjJUDhLIAvzv3bri/Z6iqu56MN9USrdi7fGju3UFGVLtuTMdftbAMnqliR4
aIcJg329J3Gj3O1zI6p1A4xVm8Ge7g1ozh6HUQoYOl5ek3DNGn/VMGrAeXZqpadxmmofw/fOAaRe
2SnGix3uJ7JUPIQ6mF4vovrYIbrrRK2YBNwMVfPXOHywtdYwsPWTMMVuNUP0wK7MKXWgKakqn1ws
X3Ramyjo5NqeVQzThp2k7ioMEte9IOtI7wWwB8btqmjJdzhUHsfhY+emAqo9WcvaeUZMBmTRu5g1
2dh2VN39OMLGBTBidoaIQ2PJF6A5/Z4OWlTmVGbIZeCVKKLLtrRF6LidQ2qaU6C4TmyLchQA8oB7
14DeDhlTaJ9JW3Kdqt3lMe7AP/Kilvcu5GSQNJNGZv7n1fhzyeKLWpQIaeQ9K3THlsXdntmWOwhe
/UJDolM+H5zzF2N5QZuWt/zLEDnI2XCnJP5TuOX8Vx/1hESSgFUojVcSCXtrfRkHF5ySCanUqKml
7441I2UeagiaX2v1NKEYq1WVDwWwFuzmF4MMWY4UVK9yD+5GG1WKQGc7sDfkla+QbURi/U3uh31v
CI9qgO2gIw74p7Oe34EFoAfMJhN562jBZbax4tV2Z9ujlqIJYLzHZktOYnncJjO+R5JP9bSdF1Ew
Lcx8DT5912L2YqV5oBMKPwicMDEYXS8+8+RYHOlcLOtbCpgev+VwWNyzhWsVDXZ3K959/X01hqCs
aLeGeG18IVxxQhpkB3EUy4J2WSa5GFQyMcIUC6iu5QhTO2lB5RBFLUtZiILFMEFrhF0RiU0y6u7Y
YVa9HZDLGEKzIou67LsINFehF9cfEM+gsdM1Bxd7ErbUGvMtVng1vBxfgqTB1cOlEeGavWxPZMUw
V72oNha7bJMrS+hlzXSlacaBR2UpQYGm8kfYoJJrr8e5dNZIaNobm2xlBlqW3CU9N6iQCXgSCT7m
IkT9z4KXAJuA6JXb4kwMrA51ogQmi/WeOnPgbuaC45D/ON50sfRPSg53AccwxDIKb7PwwAIVs72a
tT4swvNhhcAZE4a5ZiJg/31mp3zNmIv8qC6JsU4BDq1UDOXCFn+XjzQiYjLxHkAJn6vNoxBCQFT8
1pE2GeolW2GZRi5JXvkA5WccXqcAAYXiBxGWQ5WetP4+NGc/5RJqq9/4vw4J7CneI2bR2em1Cavz
EVhFAyVZxDBzJj0FXrjYeWeJnVMm3zvZ+gOOGPpARvzZW7JrTgRD1hEMqtyXPU35Lq0qt/eQjy5w
Lyd6uUP2uFxdiGabig/Jsi0k82400/T992l62DbChm7gFE8T3Xplr6+bSzW1NwlfKatMsW/J8plY
4z9NVK56FJnF05PDTuFOxuoYLJswPlhQnr9eyJN4zL7hRiW5eOKHcxWZGIJ6OxrLy9zRhWRZdYZH
W/vmre7rCaUa52MwiejUXzxG13Ldabc84W1sDv6BeLxpHtdUp9PNcNAPSSTxCkqKx1N6iJbgIdvP
kRQpTDSUTDRA/GecWtpk0hMBv5xHkjBwaauXImvMw5E7E6rOhhc6SahmCNoqLL1aNTniZO3TUsWI
a3RR0rxoL/B8tMY8PcxaRhJ5Fxt7JXQlxWpgkNay/MfvToL8A/SyNRJ75Zd8jLLk7qbUkeMYkunz
tVI7RfVRUcsN85U8K8vdYfLgTu7PLf2H/p43NBKx2/6RnkNSxUhNjmf2RAeZepYzX171TZOFRNQE
0GmyWAXCwuXN8pDmeb6SUjHFCsxDxXp5O4OYPXwM9ULqWp8i1TRLPU9z9gmUQ13Y6lOOroE4yJbA
rI/FbvavwW1rE4aBRrCJF/hDhzj8kDjqSm1abiQJ/sNaNSzkJ9MXEzVVQo8z8ChMBkrAZCtNmVNR
dYAMLIK2gU3ErHO072j3FYWSsbKxG8jp9cBgT1RJUV92CcnzmXMWai7zMXNberM3etwp+bAM+l+8
QQB+kY/7xHqcbEBkGKyNBtleqjyznqY+uQ0uVG3cACX6jsMXa42QsZcIw00zix63C8VfTOW4rBbF
L/EodGdkFr4swg0s4SD5EbtRtPQSP8h4N3+pYPyzRiiSrqFrQxBHudZgysWw1wdH7Hd/ioYtGysY
px/kqwJ9K5+L8d9ubSIybEYnXxPpw01RtRiHlWdzXgdilgk6Tq778XLWPnC60lyyYC5MsOeYFSw+
eaYR+4br9RxvbhDFslQPkSdCVkXExDsetU7qTAI/RGJVT/BmskAo66OeE210vUU/q3DaYUZ3lFMP
lRdxIRv7K+FEb0poYJsHfV+/4mDXFbd1qwuo90PMjqBxw8wKDqB9d05SFZIHerx45ZWVfljuzOA+
4QV+Yrs0QiRtwk7JnaKTTBZ0P9pgjUehzgnYGXPXdvKUbaC6rjr3dE3SPePSduLnL+f6AWqWTAZW
a2BARNWp7iqIsgxLUSyJtUHjHcV1EcBTt9M+NHJynUiOKEnIeO6/nA6nu8yrvwgjbxrJoHSZQV1H
OkF64HtttLKwQbZn5OZnnKyQ8pJGr5RCuHiLFbO8c8cSm57HxZpFO1lRKQncu6RArCEMenJ3igDe
ujmeyXVzI9REZfXSy3MRBtI+L/wg+nwS1iN4FWg5tEGAmkaRf1qSbQUtHFoI6dARG29vMVkFRF48
E1cKtvqJBeNVS2m/RZgM4ye5Fv0IfYnMMzjqlE3p4aBXXSyDKd8bHeknq5sRAZT8rEdqU+vg8wli
KE6cOrajfHd6VAnkROurdaomDyV6IOzACgEEZAuC7X6/VYoPpo50V4Z7hSga5l3+/6l1Cjkvvc2K
IEA9yG2CZ7dIFcnAaU0RSXpv9W1NOLkNOlTyRRG8dWyMlUQ507XwXs+W/14DkcDgRl1kbw388+4q
zz11xgQ5uk7ikn8y/XXGxZTfaRyMVfYtsUZhKm4IH2gdhQ33Ts4PG+cCFgcZTuEcDr3CgwKYaDi+
f/QPhnswRItIuXKleL9P0pz3odMW8N3m5JpWMQMU0YaoeGy3xwnYhhzlcG6wndgU3MPA3Fu6JMDP
r+0mIMVo7MT0R+Rub801TIAs09n6t44ZI7bNs4bZNpITtH+4zdfwxtNOsHGNCNXHICZAPK5AkVx3
bsCoWAeh5XxMVRj4oxm3ron8ZPuSrIRXGLezROXI32se6gYInRO5szI5XxpxZxaevFfmNGv0zscA
8H4jKMt8Ow+3RFX3b7P+Hyj/H9nfeebzLcbUDNFjyT3jHso3AXt1BQPZyxQ2ajoeK8jSN9mu271I
eCAMynl73VrQySOrssHXXu5dCYtAq5VhsyWAyL0l88L9ed7v5mefgsFrSd2lZiEsPqZEQGUluiiI
uY1EmAM7zNtTE0nU4slKTyu2KOoGWylXXZ5iFlmAIuxhA5w7lZ5ReczrmaD+/iZGRctkwVTSQabT
7Os2ZMVrTDEAyPbZdZAwCWeuEIkPl5L0t1mF+67Y5bZJ1uMc1UzXGiHpipGebLv2OcDN98lVF/Fc
g9aSXBspqov/6NLB0Xp2T5ap0J0NxxZGGtoc7LeqHswX2N6isp66taY2tpIV8zN6VMOqUM++Z/Hp
Sf3JfakZEqA3QN9oFZMn9Qab/MMjnJwu7NaW161w0ij0xaPI6btTE6yClkI7FGtWV5zwXrAA6oRa
7eAM24SbG+NqXzqYdBzIAASXP/fVS7myGtIccDc4omJ/7z/e9qi9eHCE3oZcIMn2fToJ8Dil175T
u/XIUj54kR/1Lx3DI5v87WEuOZPXyj5Ui5dj6EepkJ3ZOOmedJYpcqWyVHV20ipYJlsd8sifkiM6
hNhwJkeRs6t3RF1AWrsvWSaWzFifUy4rZOv5GT2mIYHXtW7lUBVw+5jYMUwZvZ+MfqHVYnY+l4DM
XEnJtB1BTpZjDyU41J0noEBRSRrDeOUFC7rKClQupngHcEA3x/SvNrDZOG7mBKzH+L6o9/XTva72
VURfbZT7UhxE+1oTMqn5DRDE1+u5mR4mTQguzBpTOSnoWhwCh0BD/t1r1Ztc6e+jfgH1NV9u5yRI
8Xq7LWoKsn6g2PmnSuKZKcJqbLJvw4MVBS/5jDBo8T1ETfRw5W5X2R5NoUV2BUNTyaTbKwX153sF
z4pcI3m4st3vwDQXSLSfhJf8wMxNWMkEcv3WQLxW/5ivDkkVXAdB74x+cekitQWzdIeXsabcY1rt
gAgjXaSJk4/ZIHcw8AaURT43iT0enqEzZk0Zza9LcWPTgm4LqqqFWTnugGsSycwOkTrDFXMgMBtZ
EhpNtA5nQ3yCJf81qFXptasRZrwaWwTFupw/E+YkHgyZ9c0sc1By94ZyvnF6+5f0q3XryEAgPexl
TzR7O9I2IAgxEbIkDMTSt2Y/MJDEU7oShSvpiwhAIDk4uoH75TMZlPT0TUBPYEuXImDb/99HTnpd
OClg+TXe1Ja5xP4e9JbLtZA1jnvYwnPtx0CsosmAu2qmWAR5yLemk6ZBU5IUOOFdiJ9rbmoqOnHQ
TpjD0rJnasVjntdkYbIqoEAUrlAnfuS+669T3od0liGsmRUj3/WWKiXQjm0lKxaYIKS/gwMWMOdo
jXHNK3XKnXuKjPDA+LpzMmxz+sfyzpEz34wX0lcklNXTxcCDl1E68qZKXM6NGHcKueT9rEx4Ed1O
oGcvCYh3f4IbhZJf+NvlWRbiOofxZTnuxhnbmMa5tmGafzQE1EIXQpYkTmUZQgVYxdR8YtcgHr8v
UqdV1DuI0NfdMXvIzA8JEdusvHKWpco/ZvhLKIQUF4fq2/Lc8LAXMUcrLCTxok68k820QM0XU0sT
bIxIlWmIUlYc8C5qaHWpT5Mod+3NNiAgApplgNhgjCbO5QdJ9C+eOXL0E46oVRQDUONf/+hycHKr
8uxvy9i5z5QdFxqcoxW6hwPPVHDkfEyCc/RbkWL9XfMp52XSlh/wtYR70SC/WeWPlrdzisLk+gma
P8HmFnb8FA5LODfqcDiO5UkpDNFZx0LfIuiNPme1m5jxZZX28mhQy6g8xaFbdH183wtylj53dRo9
DDjfmiyOm3A4MoNbYFZ/A5qv0SJstuKMXz8DJL4SKGqOA0sH6iYf9gX0DuRJ+4rwJnM6OspLx5uU
IUqQkRPXsp7ZMHO89IA29zOVgtehll85HE81tq4bKhAh69Epx93KMcPjIMwRC83oAt7BGtaSQh9K
gjoJFlnf9SgR7t7IS9NOPFTHgOpTrBDSFosyA4sR3yTqp3CQ/Ywdu/HZZjROrnGbVoQrYvIYYe4P
S7hiqCbr9Z4jpImc6/kxxIERXlwrjCEhfe17aOxOM20GzXHXUnRsK8mus4R2d+6q1NnEbu2bZ8IT
CjKsfNnKKkpGbgUGyM9TPQLpegvCVaEdQs2JBbSlVPm2HexnuYGKrGv22hisl9huH8rD46jt7Mle
X8h6GYGYq1RQPCEL5IDf6exNeOkD2CuY95Gfxw+f29LhOdouNeUzzvTURcJ+g2J2D4aJW1KrHvvP
qSoVXAJDWmcTN8od3c6Ju7oZsdYpxww8qTA2hKrUWAXBQEyV4ql+jcwAe1/rPEu2h8pTUzbP4LOy
MBQPvemPAUamGAWyvcpUQ+zPTNmczbVVsEvZgcfPWuAoa24/GEFqg5os0f2Fu8Cu1dVGL/7WAAWg
/tTBhPu6tTC0c1NzBSnqSoG1b6h+vB9vYWlrKjiQ7/cp0goP3BTOC/S7ZDVVyNc0QBs8mmXjT+aw
cbdK8UsA6KQcZuUKSUhKXKVRjMDaLB9TyRQ3ZPaTTGl90ODfM5peQJCT//+/jDd9pGXngO50gd9C
zc+905coN9WAQ5RbxMx1w3D3NULd267V8hc+aJZLuftJ7DP7kqzHLhbagDcY3nDcsNdsKNtwoF1O
Mkmz7MP16yvYdB5nBGYHMdx7s9UbcY6goSOelOzoXaVin8tPoSlXv0BtaC6WWlQ9Uho7K2wAxzBn
17xrlgKK5FYBNKlDFRB4h8n8QqUVhaZ7ju1Ki9KaAXcXlHoL7QDZY/Nw2miBH3aoWahOtM6Zktya
XIjSuI3HoRl+gU2A974K50u53EwKEixj/B+F6N/XzvldFIg/T2fASli3l87BnzwZmcotHKh5OQeK
OLvxl9cxRFHZdVn6/g8n3GVF65h/LaH5henbjI58xP3L+FwXNH8ILZLXsizV4MQbPsz0gkMiu588
TkQ1i3hdy7mJ8TyDt37IP6f2X4WMggrxrwLLE/2CbvdBKB/fJM5+gCXhmCqYGFHIg0VIkKNE+gm6
AEVQ2P0Q3xDufmwB8TEg3NT+51nlpN+x8iYX/hbn9c10HsHQ67iG78b5zQcZCYSMOOGT5Zb+ZgFB
iMAnY68XWJXsaylDUTgNJoivmGd0TwCdyPCkoF8h7u8b352DdjDy+sgWRiVlmkHFPw2HWWg+BizQ
Cm/bWMQ0oJ5hVZGvueVOr1/PS011NGPTPxHLVX47ClHZdWCsr62ZacJmODnXfqDxCjaMUTKUdxJ/
MHMu5mBrbJ+AZwx+YUQrfM0iaEDGQo0CU9ijXw9VLJAr+H78PythUKX/+euaercYcnP2Qm9GZIZY
Mmm2LO6LHURdjM78/WaIyb8xGreZNsMFc1m0KtDj86a6z65bXTo+csoL7uS8IgFZ5RLGPmgnEUNJ
ejMQBq5+UJq7fOmBwwKURWOGA1WNfY7JMrnEDSknA+lXZBUPu2/F48MuVN0XHSbCGvN+au/7VxbQ
n8KOj5f9VvSIICT2/hMuFJpZJWw4xqCVnsY1n8TsARUow3PIn0UqisLQ+7HGiwmVx8x8mHxjwaSh
RL1REPQJYnGmJWPC0mEn2JoAPbz/UgooTLCOX/KQKPwzaS8KdkFNWfAi78GU8Q/XOJcbD9AdNtn3
z4JJWpUyq4FwvHbMuFc2d66gZ2fXzdJkz2RZRTahO0gl9ZlAEbt7SkyhcRxpTHj9OP5Q4+dhZxAO
g6frd+eczl01x5a+kFcaYrtT473nEXFkzzseZnAyBeaqOU9vNWDv7X1SON35LqV7hCGOZFKDQsDg
0/jueWS2H1eDn9Fr+v35yqMT+gYT95qnUEeci5SUhuuED1h+WPlyaLfpeahFEXsZJnVWni8iZ2LU
1vKyqCTsoBAocf979O+e8igMcBVRBQneFGfNC2pWyL1wUzAhkVtXpd0eJEoHRgvroDPCzqQ09Esm
O7pNVcl3eqtPafqEATDM3rT5J4eIKmB+k1y0ZqCTlaBfI+0xMugUW9SbacZ5yn/4CvwDD43UQrJw
yQBq6sW1nfDdWZOxqMN4LmDk8kJJHzUYBwORDdF+AhMylG43YTXjq3pLNLYYajH/6EBLKivA9XdU
cF7Nyg6qyfl3LQIxm3XJLygv/lfk5wuJelMvghByEklT+Y2vf6tywZSPugs7eL9RILh5FdmiOzPa
o5cN6Cemb/jUzHsr8mbuOsUljKQsEKGkB4DYMuuHcHUa2YaFaHgyZY1YAOjejsv7sjrCi+6AxJsg
nd5jHZ1l9WwTICHcJ1gBaQI/54+NSTsLilNrD/Z29PTu/73wG6HkzyiPXXy6SLP7sEJnBHBiqap7
HW4K8XOL7V7jVbdDKT3L3JZUcwK68Y8fzlCE6oRpSmoivDK0J3vv4zBOMTTzFu1XgWprXZJmDhmX
HEfP71ujOxotFMCcIKhEo27l/tNt0pPdGJGV4v/TLppKSoXytofsxhUipqBUZdzTUx6BcNTmmo+g
yM5kJjhpobIY0iufPn/7tcHgYajkRmF909CZE9aR99b3SR3Be83TcnhanN/n8uMaAzxXVtSTQyZd
0rpOJe+OV8ZNK/3JyG/wNxXLCJnvHFbSBmc/g8g0mrZM1QBXU0bCUzzoW8Z8AadJCPz2uYcxJmAW
elHsvcYDYiO2xs1YxbHKBo3VmTu/Aj8HUj6RDQHyF18M6mRfihJP4rlj7VbeFTaPRDYG53aR6PI2
9fER+x3PvviYdgNiXzRXS7pnKQYvHkWNj6mI2Iu5GIb+aQA1XMdxOEWQSvbEP3MyIX5q2JNHhnWP
gPWDmeeQ0iBVdls5CR7RDaxaLsZcO+2oVE2LGw4u30XxyaopWNB4YK9Y2BbI73RTB5FdfaENS3cJ
dRB5iSEHD5NXaBy+D0Hkz2Jeh8/ucQl2Bm2PDeON5Bo/uNXIRd/ovZefpsfb+DDDje7+jzcYAnJM
bUy2wE2haB9gRwijHuOIfPKIsXezBx9aWpi0UIzmhq1fjc69hJ+l9uOHNKHqvbOVxm1f+P5MkGD/
UzFOX+iFHSVxYw8JcbH3GcNCC9MRIUjKtCqPSPb0d25MLi1StTZpTaNynBKqLZ2jC2MwKMWA4XXR
Akqu2H54edTTsetzXg7QpfwydOBcq6uZ+doo8q/0H4sC5YT09c1fTjc/GHSnjCeiFZaOHFiTdFx/
TV6rPcm+ifdbDAyWkedtwkcnX0orv6p4LtPH9QLvtpJkhHMnYCjz55O2ilcZlNkjunaU/Bj84ODT
ygEPkuo45BBY6sfYMZ+tzsktr8+P457WokoaCx5pJO8pVgrudVSfV1O88Ryb0LmyFbo2bL2TDaqF
G5KcPQKy5AEuCpl9FO3cKlZ6nl8FNFcYWzjY2kF4DU8ERdTAdjUT18nEcdmnKF16Gz04lX+8eTFJ
412HRsrdyhIDHnVV5KXtznanaZ7Ob/c23VGzEzsK6EG+k/MUlFn3pL+VOufBy8HIyCylYf5lwxyT
ihgcWEbUPYwRzkSAf6esyc9bu4rcmNLW9wKnKs5m727od2n1Ri5AIi7SHV5LtojRpBFz/mQ3Z9Cb
mLLzHWP4qYakmBqvKsct4IaL0Z8Gwwckw6zobyJAm/6iPgRXNiwFDGX8EcAQgBlM/zDOJ8WrvYTC
V6TcL7iwSiQKqogbiWQ1FFucJMcBg+ZTzy7UjDgQw1mKhgwhTQnDOnRDcxx2LWLSqQ2w1+j1RO4y
OJkc0C0mz1r048ofwSWyqyhW+6FWCDmh1VjDP3oitYPGfbVud4KDTuJXm5eR0BiWlWaM3rv61zl/
OZzZk2uTQI0MvSiaOlxkpSiAiO2SvnKRfCObDbAPZ+4tjQBMqJIzPjSWw2EKr2ArLMdlkAUoTsOQ
BihpeuuHr+7SZZCvsqqLj2OS0WJsTrg4V6wVeno2nVWP9tKKDbGY3SEcMwPTj7MidPQuTHn90Krg
clJ/EzERZExtSeVTgEsqoC8NQKCBSVdzJ/HsY/sr2MXpTKuody9XR25eczX/IegvL0Oe5I3fpZz3
Bnh2le+cfHZ329c4wlwPzca3mmjDPaSgXD4+JPsE8+n1PHZ5scbeS9gNA0LM8HWZGiwGqel3LFBx
yooeOCGhA19Nk2rnEvUEnocWwfG24xNcoP0kqQzj857kWgCiEVOzIHRguz8N0+4Ol/mQogHILyz3
NbNmzTM/VPuJPUqrkGluG1kR8uro0IgOZnBV9H2/z3L+f7HxfwnqO4/eKFf3PxvlybsrAKpee3A3
4fJve3PPirbQ/+TYS8cJJGidI3J2X4TO3gz0mlRdi7Ry2D7hpUkYLsBVoxM/F/zHiBaLOQqNTUkQ
sUKAxyObnNq5D1AB3LGJujgQtrFDn1fDqW5IzIqN0GD7xsIfWDepTbZZJgWdIim1FdqCjSun6meA
RG81FOi+GHTan6RKPqKwPSz6GGWQAcm1X2SCOtef/zYbbRIEIaKM4npWL1aTHdRyJu+VqbKEQq4A
xV8fGvi0pl5o/0EMCmN0NVwz2XqRawwm9BOozwwHl33e/HueBY4yfok8opj9fF9mwrh3ATOnK2Zi
2/mfE6pp6hRtf6RHHk4sVQuvGPdZgv/Dq6Vc/uNt2uAgLIYj0vBTIZQEHpllmDZXl6nliNvkW3ul
GcQiCjGZIpnp3WRAsImiYNSQvFLoCFqjoAhCiKv8nwEswqMmZs6kT2ivAS2030HTVrzk4dWpxhG8
YXeRKEQtA85cLC5mENUkLpOW0VXwOrmPnPbuj1Cn4C/NHI9uUM3y2yvgyIglM/X90ZMwP36774bq
Z89qCvzZuOdHoB0CwbhXC0TPY6eiSW6YuD9VYdeLSsmNl39O6BFF0u93oHv5/EY9LNr0o2FIaGyg
xcMmL4TwUzEWbVl4+9XP/tf5i8LMB06pn1FV9dyzjWNPxZVIPm3ZBly2NT1BaXgLNAv8eU2ViAUY
tsNG6fCjJlps5sACchn6puLENcClFk9cD4Tw/GkZC5TptoPHPZ2dKJBNuuAhxGn1Q3BiZ53JfnXS
lY3BcOrMB4d6blD6WjAlPQur+IOEsP1CHxlbxxl/vfFRIC1iUA7X+/9GDrOHiBBBmODaBGtGkDKm
Aka6GR92fOoHsrGio8R9pAXW7W3UZOge7vhhpG+my6h21u7NfUWId7QK1u5UDYlK7Fxb+rxAYxys
ZuTf6OiRDG/0Q/BBXjEovlDgKqM3CSDL6EEOsJOuysqkw2D8FhQW06OpRlSwdOxNNroe04iSZcdE
OMTnccv/qnuNb6HEHZLiBwnITOEwdHBmVBJMH0WeNOMbbwlH7H8kz/wKR6TVxirGL9S9lOAOsNbo
6NGxJWsevhoIsHlB7EisPUaQVmbI1Rw9jQOmyN3yQ0aYDI2gWqvkXpxCirbYh1YLBJ8ls+TZ6ogO
P4k0l3jLKfNgovKH26e99m4r7jBag8MqXTQolS74God0/6b3hPITKS8RCXi7NFiUCoNF/ZiuVciX
qcO2Zwt3Ohk+E4N2gzNaij55gDK1BKz/47LE5Z+8/vGbwGu2O9OXIHmfGR8vZctcGwwQyEVTNpRy
OP1o/z/cbnEkA6oLuUd9gECINkb9CO8Ye8lljSrNQjCwOrMWy4Iv+c3DWHCQDs6llwJx8vtkNmQu
KPrFdM7j83UW2GWQLHSc2/EN39Fky2HqKjOXG9Au6v75VmfvqwNQ97SVGh42WoXLN/to4wQFlJbE
/pxkRuxXEp2b3zTJTNSKianiEhYEVC4rnW2ZJXc5yoBXrMthHdjz/I+ONCs4yh2jPcet+LV7Am1G
ZE1Fd6qf5fSgznM5ho2vXr2+LGy3zFCkqKdN/nHO/5DIWUUfhO4kcKg0vMl0P3u4MO7HS5JNevmU
x1WbL+vX+lK2T0mvvdHdnZjvb4pc4Grmv2Tz8lHtLab/P2x/W8OsfpCUhfhkd45jfs7xzdjQDvUQ
tte9562wkEXPI1ZnZOjO1wGaMIRSb1Rnhj8ZOiTQ+3iaNXljEJXyfNcrWw52j3mnZkeFIVR56Chp
MctQ5p0LrExv3dPl9kG3ftpKS5n4BKxgkbfKftxvjQHi5W+zrJ5kk45vTP+DTOdkq8Dh81EOOZ9P
+VpPjSzkuP7ighNuOuLEP/hOmYhgy/CbQ/P8z4lSMPiYC0skiwKZRYOc02QoDmeFuodLtP86rpET
o3B2WD7qfRlgaKS2fYfAJbt0GhphaKtSJ1ctlsDN6hhKOXDtFLhzlHSTfjnzamSLKZl/ML1P75id
IYV4MLvmhjwePzYHvjkNOlu4YK+lAarBieP7s4OsiExh13iYv/4kj5p9Rhfgsi6ffEh00AgeZ5mt
eYK6PcURMNR4b1VZJmurpZIcjEmHlqUZdNpvE1L/HpC540y7vJpjv/6eiQmkpRuzkE0iMBaTf3I5
ZAdRsyhXt6TMjXM62/f0456v9BW7Phj1TCazP3YaysyFX8S+ei1Sj6sMYQfkj6dDEiU9I5tsZfOi
jg1hxBMeTxkkV/GAJOErgT7AyZrtUcw78LTESSXA9EpS3BmApqAE7u8rcjWjKoI8j7awJmaybNwr
g36UQ3Na5AKIio6VGK7tt1mYmuD3GDyaPbAUB+XHHODkcFw04eUv7JtbQLHltCKE66zIMCuBBPt3
Dk76ZuUwasKqcgLX+3redIN1MuDuxIAjfEWoIPfuQ0fYUVFv9IGdgqPerOfFmUN7NQwK/jvjWCTz
d65rXsiCvmgUIXziIUdFX2/bmS8X2d+kXVpgvcdWoJC0BT/HYNBX0aA7w9vPDwdenyhVryWIGurq
3335IlUtqWTdiaVYp7PXUpUd30zeAqjkHZZTOWfLHv7ZivYugut+r7C12iJdqNSgkKMMOPhv2Vxc
u/EM3dKproITsWIVUnePSc0wWlcDXjBHOjHkl68TUv7TlaCo7BQZuFyCQ+uXLCzaCPbwTYH7ooDe
HM2/wox3rtn0Abx5b3g6LAgHPTUDFsGeGFZvHve1AwhqeWmHJaGYE57fmA+BeiAOtppe6F61iz04
bzlDNQtcRabMlSMnrIabEjfXBJ+xgGfX7insX0gru5mmwFdYZx2RTRLs6oGb8G5XkSEMatSICMEW
w23zjNGzEZ+8JMkwlhSc9j/raNEx/jk7hANWyfr3/nxkdM8mQUv/Lmkz1S1t0d0lNUlro9i4HYbU
ATii4LsH5Y+rfsFIhFoYpftZ/MzVj8/GRhtb8s8yLPilnsDrsvHW8ZkAbNWhkwbVIgT94RX8qVCd
U3WsSFxcKiYoHh3HTo/Jznf1+qiBFBaSueVK+YuuY4ZeUVd13LmU8J+BeAMZkcimdZHOfmW4UeKy
bg0Zaz/f9L4psIwUgJ8mAuwFVktPXO9k9Gjgut5uAZC6Rf5ldXveCsxKbHGGRV59cB+5CnyRbmCG
3308XFKeeLIxsRh3qW0wQLF/FeRNcyyl8iFRb1Pl3GJde0cMeKxIzlZf2fKlFsDE4IgVu6ioDaDz
QL2GH8D8Ck/S2mDJpWn2YN3ohDX9mnO81pAl8iMxjtVKIvqUSHtWlAzYuHWb49aPZ+qgvUcfH9yx
QRyqZIX9A0ATsYyUsElTuUFqyyRka8Q5VH+p2yxOTL5iklHgQ7ww2BXpzvLGzvZQ3yS/msZpqkpE
pP/dvMdCPZiVq36Vi8Z/bRGIZbZoceQG8nH4lOTPX5FGMTTKUJXiLczwEyzTDorcFcntsx6EUo13
71CPp8NJwBfkKgUd0DhBNO9iEpyUKsN7U3Vx4libPsZi9Sx/Aq2K9wpjlwx0ZdJlcCcTAEy/ecKg
rX6ZUHFvewl6JjtYU9lZOZjzdUQDl3bE587JrLX9LbcoNUDtxShyi+sXDab/c0akjlhlcVhWBPoC
LjOXkVqdToyZ51meqT3toOFGl+BchrZQjyTqLvOVKKuZOPU0EGg/Lkn+my06wDDd6Whcs2gPRjyN
EriYdB+J6Hr7dtyO8rpj3pdPjjaPtuyGJIeLCnMoPtC9U0MIQblfGHWyqbNpQNUfKZNF3N4jBM95
AVMZ/6cp6MEmAl0kFWvOZM1HFgziJzO+YmzU245YWbL3y+BEt7jGKDjcg0U8+805iOrWmsw5gRb6
zfTjCc9H/tkCYXfvPCX5puvwVEMV+FQ1nTqBy59MztjPim5tymrzaOmkL3VVDDEFoufRNhAALk9f
6yfP3W78cjPLkIORsr6rBaK2dq11rYlxhyKNPI/4FtnOL01arujOvd08+Fbn2Lxcrf8aSYrwvtny
o4/0DOQLXgTxKbphylfuRHc/ummiY63nl5Si2B1+ffk7EKfyPjNbl18ic97M9XiDrCke38Zu0ChC
uqX71t+I5Sn0mIQMT6pknAXw1eEDSE36lgSF50yStA5IMthGyVMjVoXoWNAcYHPykrghY5ZYy4f9
2/cW3vk92WsTMhjHBvcdxUtPCc1kO4DFXJLDp4qgaaqKt3aC/EDC0f+BTPVzomiQdnfqsOyvh8VB
QMFosXPi5sI8q7GpMOrrrqxfBtXOlNNwJlGp9wg+zp/FjKJrZDUBFel1AO4lucXaLCUW/0t2kJdV
Xx2lhYjQoGXMNRFsB/Z6he4XRLAY0PqDOsy8UBaUpTjq9ov3wiiDxPj228lpD9sSoSpGxAK+juhy
Ds429Pb/PpDg3jxdcRRDrajeVMOuu0NPSZLtDMV+noyBq3lJr15nUr36cTIiPzwJ8JD/xVzpmaf/
Dh6F4tlzUpMwumbBDzgiVtvVzf21dVi55QbwRJYjEOjldPqzFFlsjs4UFDPyZVUO6N+9BihzELDF
NHKYEftMiQ1yzX4GZ/uVqWPn04WsP3YzsNhXt1+/g27Srs1t2RpI8h1iHe1w0WwQn+3jXHjOULYI
/akvVM4BR+WwwQRM+jtYlFnsCGD7EtPLC7Wxuby+hBfxAZNk5+PEUMmRg15YCR0I4dpPvKuWgEJk
7x4xEq4pntBPaJNXfd7SykGmIylTy2yi/bniSRynrfzfBT6mmUZz03JLI++0zFX+T/AwZqvZG41E
w5NSp8yEjHVMPK9XrQ/dZ58yXT/D4gDJwuInZ8LV1xEu8H6HkmhV1TOQ9BW2n5BhrZtYgZEgYiy3
ku+yhT7Te5eHwdkHAEW7Os+DHABUQeZgTiKjbcTDqH7T+DctpwtEoruqBnS356itK70PbaTOJ6Ms
K9o8H9OrkxLSPF3/2/wpe6O5nGtpa1i6ldVNMT/jAQnX1VDbNnZqMG9dJyXlyCYqpimFqzqFe+Ml
3WmnKzfKYz64+K8xHlF51ywlHc+/O6pVb4Xzc6tozc7jyWphis0HNzgtvHUszQeHKs7uOxwITN3r
q7BJyDPYqPiiFmfkusu6l0TE2lzp67R9HdQTgbXD8w3NWoSutatTtMr2QiOiSf9ZjFVOu0NpdjfX
3sB+ZpyhltmQbTus0is+4g2DH23h5524dN51UmPxLdVGwYAZNxCGHVi21JZIC9L6SzkJxJvNuDFx
0WsTGLQD+YVVXT9OXAS6ww5ITQjrp0Nu4rMURgwIy+WUVolbliYipL20Yrm0Xsl3qvLZJKVU4Gdb
pNVjHomUwWs+PLoethMN5JgND/iq5LOpabTKHy42TMZ7HcZkzuFZxhTPqqUOmqa7xrcB7spEgrKh
m3lY9FNBVF9r3C0TKs5UOKXYeJKnpYRtnuAHVoFCNmjmC4WLK4mE9WqrDRbk6obTs4a/tYpIltJP
fpLaK+yDEhlKuj/2M6/bqffYWxRDz19tRlbtI2UZNlseCAzI/aeh63M6CPPcmy/CD8W6LKpTlYEU
v7hcg6N/9+X8NGNnut6lI+vCzF7zOuPoO/ZgOLCwBlH2upkHi9SBQbPbKnuZ70WEPbl5UfThZyvo
dkd+94eYoUfpq2XTMxwlnWuurUiW2TFrGdSzOuYXya7vh3zRi424f9uc8h83Zt8oaHZDHxz6WaYQ
RAfIykFfILz6hsIjZw82sEqHpEQ1zwmlWs8qdPBkOb2aZHyHT4ZlQOPV3hhg/kjWwRuhEjlUA8Bz
TsUt1l/h7n9/g9ahZQWqRShI5uF+Z9o/e5bZJITCCyHTQOHP/cZFqck04rhZoKfEs8SmSOZRTSDx
eEHF87SRMzvh3t5v3u7GdWWsnuiiM9jr/2vILpZKotvxdJDtO3NR8l33W6G0b6r7wcc/1Fa7WUL0
aic8j6L+91SAaMJlifq01SeRes+3SGCvBWxcpYfC/7pFIOpY/1HZ6BEUQr5+Wy6AJoeGgTch6g58
S+j86p2pni88LVe8gJP0x983d+NyQcaKjnL6gUUVXWEwP4U/5HtndDT+ideGBnXjUHJzYj9CBAK/
BPDUsvijaa4fbhzvlNlunspIP6cjQiLKy5FQZw/GgqTuSViPpKVibH9gLVkUiW+GpzAKZD+nh/Ul
2k2Z2quLRh5oNcfNcgJTp2tcgAzy5xlHAZa5HtlNkAHB8znxUugBwDgcNoVKPKWuZ3jQQVl82822
pEMeWJRK78o6kGPvsSi0usQg9ES6e2FJIqKFmPsgXFCr1vrb8NazY/qknH8ubEkBK3ETZ84vVjq/
6o5P7hsSQ365HfXANogvpS5t+V/BDCO8138JYFvD+/0aaWyXXQLfrMxka3LpeAawDWI6OP4RvZPf
41Lp6Rr+LIaF8k+hh5cz7ufxmZzmMK9yIa6oyb7gAOhdtDNGJg/cMo7kBIxISHXRtcFto9DszEIy
/QeSgi4CY+7cfLad5UeWqZvKfT2Yz+V0e/M2avSrk6NcjlxsJlScy6kAV1cx891NpkkwBcryN7R0
C9u2PazEDJWBMhox4tfhpmQZO+Ggtrobkhy6D93MwLDiaovXstvHyNIik4WXtvailK2vp7dUOcCz
bAMf2aY5STi3rkMfwopVGavtiXG6I4LjMgRyy+ymGISERhjCIugwaS0Vqov9TqadlKIBqSjXUbzo
87Smk+Za1q0xi2ZK8LbGLJVGEn6weWyukrKhR96oBxP8kQ/qBwJGP7xmu5l6gCvL0s8pkzE1k2bC
T7uYxfOh2FwOwsKNQopHvvQRSl6XFnLpBbFfWGg5SvNudHmlhnd7opTUJMDHZweJyn6vPNuMf02B
Mc7eK0Z0EMjJBOYqB5GWcO1aOart87lPi4Xt/Bsto7KtE+1SjSKjijiW1CpSp5V/exn2p3ehIqpQ
UN/U2eIxR5Cf8mV8ZehWOr0kIRBjhGrfLEuoodqhBRoKB/RyXzJSr2FUmt6uIvJtSwZ8ICNvAEhr
1Fz+k5Lf3HEjdXtOiBGhSV+QtFtmQ7xvwJ2r3O73kh255+xxkutAaqrdGvhEVSHEcqjHuHK5P24c
6jOB1Tn4+WVoomBdfrrDLvhUrPBBJNrPS5FiQNPqZGpxij9FR0hreiCqidxN4JC3vKJ0GwiLF3WY
hk7GeULWR5/kMhaAO++6zBMhOo1j79QXLWNkJIaOW8jltMNJkVvKIcUULDEZCdaSa6+pKKW2OnRU
HUwlZmOIlb9Qcc/h1K6M6YwjH66gnBOC5bqmp6GkElEWasEuCimrgw1FmCkE3shFQbMrg7CEQCDC
J6XQM7bi1yTHgO7FVRaJgQlr/5x/6w9GY8br3v/QYoQBA4LHiNgnvbjf9TWi5ZowW+kSSFXy0iF3
jjYjhRxl/28upjjvN8m4u3EM4I4A4cWacjHjRn+OcP6X/Ru879s+3Z6WABbOdXsDfQQzTDJTBnFq
+wt/+zGWxqaL6ExIZNrzbWJimTIse8tfpDll0BjVizt1hwx5kIyol8cH71OmzPwpiq+HQSwbWfM1
bPCtFvWvl9A7dEAw4MGQrFFKPPU3sfK6BYSO5BJc3m4EUrFJ2unKYXKLACS+wtj/l7eRhS0hoEXF
gndHPS+NWVs1vZ+xhGf5nc2qUkm53bD0o0XXVLG6xZDQENMA0EmB5AD1bgG+7KXSlgqo4TqYJlHG
5AMwTX1MWMBOMShnYqOu3xkAdsF0/2wVblPTVpzIQhZYpBxr8l9a987SfLm21D17lCvelZqNTFAZ
xIvifujg3rtjboj93sZGFWOzZ6CbY5n5z2ysJK/UlCIY71VOZq5WdU5I0E0nc5cYgiGafmHoJiye
5n2U659ffq5qK4JTNXN/XLMsKsyfTmMosQOxUrsZS+u+uqF0S3GnxmPAxAHkSfOEoVWpcFESvSQf
K1dqRl0GvptUJUTQZ0hNpNaa5Svn7l1hQPvGsWWyJQHWxEcl0SVVInHMe/7Pbw/iLW5h7Aekz2/N
hKOhjlQOpBMRT/qd6S29tK5AhFDYJUC4XOJJ/Wg0FlqALzoSy3Zblb9JcRdnmm3uH2kyihsZz3Ez
k5FTlV4uLES3vbmYKoviTby6mEjXp0wIsTuCLaW4tQW55aAGOemt6OJ1Yl4bRkuADlW+PahkKRlk
oTho/G5KQ2eRDpgQTUV67E2Yz0KVkqbUOMSXhU5VObw7ZoO6iyCcZjflH+iB3cu/sW4EoBtp0VA8
IpC8z2P+F6xLZhQZ28m01imGhvHa/bu7UPRHs+00ijCz4glgH5iZ6zp7TNyH13yrP9Hrx6QrCgqA
0LLjOmmW9HE6ytbcSHDoOBcmJahyvqffIwQzcwYksbu0KvAA7dBMBwH3IfHU4tEIKgA0WXBFbqAm
aIkaWrUBB3AsdQotoCMXm1GvO4zAps5hgPeoUqotIOa6OsZv1XUGbzIOMyWrvj+rwY3d0eIiUIi6
xNAie2StV2N2Wm9mHtRLjjdKBGQBtPiITSszTnt0RgyxkmZSbs8rw1wQGspwm8O976teh7fmOjrd
1IbldMKQ6KHfLbR4x6ZxGo+5DCoxhL275SXs7RLEqOLNA7QgIVh9Q+Qpe5lR+NZJJ6ujppkN2k4X
DZZq1C2uPsYCASrxEqPZXw9bh49t8ew3nUg0AgoHTOVZwmun7Hvm/GCbC9k4fZnup265uFnC8Fwf
CZla+kv21J3S6WDyWF7qIHeu0HDYtessjEqV6J0pVtLnK8KbyXWbQqy889x8kuXW8/q5joCmd09Z
akWGbmFzivHhmSq+GkoKFaUAc/NTxR3gq/m4oLblFAhqzYyT3tmkjqgoNvjYSa9SfoMhMOrobJV1
eLIJupFPO67atL5spFmhHwP43FiSBOb6mLE/eJb3INca5IX4/HKjyEJtsoUp9/ryWuFFH+UlM6qD
lIklxdXmoIAaSh9TsNYxBwtjf2N6ydtBsse6gGbOFVM6kJNRF+JcWnkz3nFlCxh98Ag4/gtKZ7Ah
a9AnZbSmPPUFauIsgJSqS4zelQpzB5UqDXMBIat/SqXzTuL9xhgECoxCoxDGxoSjH1WAtUtJOudT
9g8YnzcMRCU+LN28BoBBTwl7lhCuFfTP3jXUgs5+f2LTkzqj5VTWpVP/5ACAeil5gl8h+7Oj/jyC
ifCaqWnVi76ImJXgjtkh29EDeb/HcZ40bAgftm0/zj86gX3rAFwtPoU47pd/yzbYenvdeOb2jTPj
YFkcEguxYWKfTL9rSekvpgvt5DZQFLDlqSAyo5eWlSJrHFRCmmeUSfEb9INoDHWo4lv2rr+XbOMt
GMof7pUzXhLzSOYZQxubb/7+0guZRTzG+29oc6i8YC7+X75JE1wRajw2PHbMQO11UxTS79QAaDLA
9kxQVD0NclCCIlmxAbUvEiIdCZgpEDO1dn390UCk1yUc72RVcdVU1wGFPuChXz52+99SI6B4q5uN
v66BRAjDRWk0JXQJLSr8SZfN2C6HM/L6cuunRkbLtbBSkB6yGGXPqHfNK3PrLjiZf+kcNTJW9Jm1
Jc8izpolMOUmJkaKeE8t6eqat4QAbFvMppGvus3CMtYsQFgscGOCJZXOpM1Hs7SkAhzMHnj8ADki
lJH5FjRqu7pS61fdIX0JmnfJcChG9+pId/oQDUMlwPG5eb9jmgQjKfYuWvgRmppEWlNx5KxcPCEk
S3yreMCS9kqm5suuEPvi7JpptkncEbGcFTUd2zduLOntP0NaYs490GGqp5u9hH0X8MGwjUvHPKlQ
VspysunqcNzpVSV2R2T0X89Rlhayx9yachP+mjbAQYfUgrj5WO/aUSo77omYuFYOp4NF36bret1w
xkRj3VaX+dH/kmp3hLEU2OY2y7YXyYRrCpOK/9FzknzJhKMWwD0fGlbk0r7W0zTyMmY94s7qylIa
ApXMCefLhSZVHFaQe0Krb0udrs3Z5XiEKa16i/38VHPinXKLhNtGZ9R1JM58Va7kiC/MrWbhjm6h
3vfm9voOWP5mXsV5MNJgohCuMGlm044e29YhWM77+qhRwKjFBigBRZveiu/9JpdmNj8Q3GM3/vj3
X/DtORVhULDrS8dLhJqIoZ3NBoZBLg0RV5dwgXughkQXKVyk5iG0JVzuK8LZtCs8er/FYwtLTOt2
qbvwILg+SrrNecrzJjHmKJnfMQHpdLwJ1S4ja3T65KCGYRsuplx89FmAIeZM7YV9vBK5Be/ZmKfX
nQ3BTeHDHVIpyi9hSJoBKOd+LhgSlvf8dRlq9wMfkrHzarL1evycpR/WBmbwXkPnEYBPrIvJC2qk
KXPz9tksGcvYA/DRqQJpMShgUeLcTfxgcyWBy9GCLwZyyCYwKAAcOwhFb0kytMKOWs3eAY3WB3rN
H4PQyD5I7exOPsujX0guNWa2e1SJHYaJMUxjkEJ1b+Ij7hHDGNTGv6ehw7jrIPzTi3awpkn0Hvoy
H1MVH/kNoHaPl6zlXM6jtlatvCHDwW3szBuOCLjZo3Ve3i+gHbODyvAm6HWjWeeCvgNzNz0gB7vs
fLw41c3evgSaXhviwW0q2XKYlvQBKhbpXSkkDr52fEiGzvC3WFXDbbimmS3sJAgPGq+iP2MaVPbY
UpaQRQpNdQPE47brzEAPam4tZjL/HIR+X7Zyw+xfNw107urMCiDUhhrvNdo9x9j1xsS7onoyxVXe
9kJxJ7z9m5Lm1JH5AcdcadgDfIj5xEkDKPQ7Sy/UjmNgrVdibWjWRaE/hIc8xHqbm92uqrbyUuF3
J1MZSpvSR7vGGh5Z513MnjMb2jZHab6vF/OS+PIA2oYBd7xQZAeAPDb6xx1w3DatOywzkKPmEzab
VVEW2nv1bREFaN9jr6GDAFH/nysJtdfVvBT/lLXwREAj3rJYDhYb1Q4TeMRWExiPOi2+rHVAOQQK
Rzq0Y4FujBt2ANsi57C5X9yFNfnXfB7mUQDeSA7oP9kBKNmk/R2GTonPxnrvkxPHDlkJBB6VAmo0
fEoQNov0RHOCWG5xKeyWOxQBYyK1S/xlGe29NH25hPBI2xQodeJreJ1zLG2FL9U8yzyHWlZvOZa/
ZDkgKtiKJsFlq10Y2Tw1TzjY3ZtBOCTenun19l2wPDDBwTq6ugKFtYb+mVsiSNCVusS61DVh9J+i
eyjM6a9ViSC86xK1cQsBk/oLHXaNt6F/DqRaTgLi0JgPepCEhgXEBz1Ag1lKU3u0s2KBO8XoVfqC
QltVWblLjbDf+fRKf3tSPH/XYUGkpfjUoJp3RjAFP0wj3hclPQAxvS9Lp22QRWos4ecp+0/g/y2R
cnudBt5aJEhnZpB8cKoyy9Il0bCLUigp0TZqTYVswA/hjNG0iXVX0KbhxkuuyW0/zRWC82IVAaPk
tlySWKZb+v53fwrrKlN+fYBjl6JmshdNQx25oQuY3Dz45o7Zo2dSWBdWSnNBzZBguWbBeXKoTvVN
6yGC1q8xqWnywJA+Gr0OFjrrP8BWFOl6SDUTF+swh9lHLc2iXC1sw1BDFUYGeJY+CQJj3bi0tALg
5eHEBTYd3kDTskP5MujMJ2alV8wCvlgs6Aiv4BB14a2hGNcvnzdYlTTe13wmZuDBiUwKD27ysM1H
dMXsNcvew58iXJil9TGbHoyomPr+o/NvIxOGnHM9i42d7epOZXh2PlUo+O9VwY4vyTEmphMcIyVG
yiE3qGcILSLvx3L4YwYdxLBl2+ErSim1gWq0CpL3tIODLw6CIUOpAgrtk2jmbyXZTGBrNmaCc9dS
eKHi+dXqQ06OK0dKtTSRN84gF+OvCfpy0/jWgaoY1qP88pGiwoTtOPbBpoK9pvfw8S59cdSxpuAj
MVX/OGLtgoVzTaI2F1FRzqeWYAoZYym/zbze5nOM969KzPfBxkgukO+8m3LAUVCCKG6GVHVzmyQF
7qAx9rYyJIOvKDxX5v+Nt5V4F96CLk6At5qJL08jEvpoC3q12/fxipPMdIsTWnetaxmI5XHFq5zh
MuGIusbHJVuaLzvCjzDFSE5XUSTJH5/yiEOwPBFCnIf0llro19dy027FStLpycxrWZQ3lkhHbplT
uETo0jYH/iT7x1K1hlZ9UzPQhWXKAvqrNRQKDq0D84akzxkt167ximf+MnwTSoyZek6vdXrb8Jhq
bQ9KyStmAiw0Zi6OrbIh0SuwCDhUDu61JY7oliBGJzOuRiQb/PWy5dXKKv1ArXxD2T4ikXM2aVJ1
EXy8YnxICsTsNq3UPXJ4VFLl5EANp5P6uzW5bWF6RNJbBF60JS1KOe9LN9CGH/U3+2v1zE+8uMAU
xMh0+y5tQZ0fFvxhJqe0tQo99IJjbULx0vWO7j2hT8c7QMqbWjBanIdiCjBftvrd8jVihBieBkGJ
Defh7hLBxd+hgqAwpJu9Mv6lZdf9vBpJVIiYajkwh0xX44VM8Yz1e/i9yvYU2cYkuGxaTNb2KdRV
MBRH2O2C69FEAvRyIfAOlSLfIYkEgV9Q9VvxLkeoYC5JO+UwK9yjzakvWY+fR6N4QkXFcoKAuLpe
ZaYtP0PZbwkX91v+VPEelj0mN9q1frwoGb/wqw3RGOlnMExW0NAxbp1CddEJizDcbrJIcwXOCF9A
MDL5Nlmc/D6vQCY3amMyIyooR9Gc1i/B7Ry74ohAI5si8wvkeH05/LToB4N1uXBDGhb/JiUtQhk+
WWD0k6KNvzxolHllbd560E5Jxiq8H8uib4IWKt7+Zue5tpgpDUi7jdzlvpu3DFw3jlv02cgDMkLT
vsK4yMJMIquLPB5ZuEuLGzJYfM4fbhzSsHEQP4tnF7vHh6HawYA4sb3RnNYzNzPzd1FZFt8OMq2c
VXQ1wdlU1LW3NWAcCugAqCBsRDdZiCJWCZWVdUzIrZchmRPEp/SexfnEaPrRIXb3dn4qYGG6FrPn
Wul5nUZH/9nkYlL6Yv2ofGi3xwEVqwhVqyh8OIXNwrKayoqPZdrh7ohiX7WwM0FRAmFjQiJi109S
eEaWN7jqqIoYTVhjNhKTW1cLYqQ6jUVmwK96MLkdoeolXTXbDeSU1I2ii2g3DW/EYHokU/hyN/56
esAMwR3ERuo/EdqX+PMQF1erl/PUQS/JdlXM7E4bMiocbvjSCCey8ySEC2bzBOhRdpLTSC06Ttfn
k+1SQboKUoOq6I2KZ1L3fmy3R3oxYYXOl7wsnYuwKQvhZD7PtucoEPjLWQttBXO9HcscfTE1WRXB
gfNC6CZkujLEZytEX3xDFFoHs1uGG1IOq/PW+G8w7v7MI1Hr80w1eJKZg8sVDLoBjzc2jt56jxKA
fQN3qyuWMyMUUShP5q0nKUV+3j7E2x7LUU4zKeVsi5VqNAW3yAdXBGhhHp8uYL/lGFZFr5gfmOtL
5DgEIlU9Zu9UEACViA3+St9UTsr/tdCkO43+16UnIDz3L1s5x8F2X+eUHUyYfk2KvMYAgs9M4xot
vqdxODKKq1tiLPCiPBfgoBemQduZOOXJtg8yz77kF9VexBex6qJ9R9bFTLhwxi0rKnQmt1g9Tl8f
3QOkeMBciurM6nM1YIJ7fggNOqCiuAjS4xdOBr6hDNKs2pMBdUBG8XxhsVT9QUetyVgfW9I9jddy
40cjdnBJxPp9aEazo0Om7dNFeJ34c1hIpvk4RBxL1/f36VLxeP/EsXgG0CGg1ClpF9Ki4e1559wk
X2D6fFbQR+ZlIdZ4fpaB+FKmHWAOyjmbj/Wnav2Okqsq8/PEd9kjn07kILwxLpRjONCgCw+NEOs6
TdYwfzw8hFMgXGeEUiSUrfyUVfoeopnO02rywlmkmKC8NRRg/0d/MtorAi7w1EeUQyolQex4a+Jx
+PfPH+l/ItcwmwdUHwRGemKd83TOYK9hly6pF+eRvho2IJwY0Pr4cKzsEOrUPCxV7tG9znyPAhiY
NPpBiCsNhdjZLNLx9RS91QMqi7nADifq2l3ACERA1SqTp3KPdKApCMfa8jlrAUv1zYo+JbOrHprn
4Ke2qOlsjAu4jRu0EhtOLQax+nOv0mmrQzzR9WHk/v4Y6GbK+M5jqfSEIaixXuDe5GLcdRiNNFo7
SoEx5whO/kRBvJCsng/oZxVa5F4YncdqBIIWhdD/dn+KEme3N+de4EISwJpZblMxP0P2KWcOSFRL
Qmm2BdNwHLNSIUvRQeIUnTH8DZKzvZ0aWI/RWkrYKD5Mva8pIOJjkD2zALTJP3Jk6PYx4Xdo8cWr
g/l0UheBeJO6L13TYGtf9pVOxNQks9MqKehL/ogs/NwSbUuE+6BXccjWqhm7/IDkO00HfSZ0s0yA
wmfXUcf61hFEMS0p1h1qTA9xQdwbO7QYK3V54M+Skq3IIinZy7pj/jXR0G8T1/YXxJWJ0m0CNcTV
/JiVN7t7opSreQIiiX+jvK4Jlpy1NJXCVM4OyH4emWb4ZmPbsTXzT3kwMO9OeO3IH7zU3qfmiQgy
qJAwNTsAWGFL/SJy/u/u0dRzl+Lfa5P9RKCKRMNsz8gK7gv/O+8sraW7IYItEqeMSQO6JjxQHfiB
R1kUuvgVNfVSjeN4P3pF3X8Hvx3E9mtQEddC2LrwCgdAUWeUf589wwkwVv8hTSUnRA5ZTQni2nqe
0/KMYgZldc7abf+0vxyrHI2X1/ttn80Kvx2Ec4Xh//CFPhik5/7Vzee9W0RE1aa38lZqg/lSyY99
EkYEwKxNK0/QZgtlPDKdNYGbjXpOJaHcV+hWU9hGe4HO+k1M32K56sksPCUw3XN6VyEW2VCsy++U
/tNVYL/OVI8TXv2cn6icT5NYB8+/es9q1fl2IC0aaiwCt+XT5PquTym666S6WfEPXE6mOPLyxHcm
phb04og/BLCOKMIKfQNZ5xpH/PDs1GapPDnOLlTzFnfLcjiD0Zh8pJyqA05HNtdaDlmVL8Co/xOK
IUz42S5PdeWdGSxMuw43X/nnrigY46x52hMCHkJDCjlm4sKrR4PfK3HhUBpByD44HNDrgzTviiaT
9fdUgQqFnmkEj9blVPSAb8nBuqX8Hlnm8bnqaWfBnJBrT3ewQJPhjZHjSk7QgKhsoOnjzOuMq351
BltDXr8urtxF26ZnID+XZQlySSZns8PMFlMgMzGM6uaycg1XS3hWmJS2JdudpU/EBb/hBO3vXycy
HEQ7SXlho6IeuTyEdj0Rou6QMoQkhoWy26DUYh3d3SxlTfnbjeCM7LhmsiuCoUwSjAliITAF3YE1
Ate1KvmQ9tvTHXdPrrQrCelKIfvOnUGZ0im1qWeLStyAkh0KjEBRDrid2iUvVHmHBR2oQoQ3YQPU
JnRc0hSof04TDGeKGpWpGQ8FnelmMXRUiQWk9sCLHmcFUm+//HXurwRakIo4LBKbiFITBIVX4Kc3
kery593+8tMJWZXYGVWf6Khonbm/5ke6KWYGJC2qXtfJi/35hNcIrycCcBqLLGb0iUYeKMtPV8aj
hQtH6L/QL0sFY84egDrxYezeEXUQl0j8doaTE11AsecNLjvJgujZtCn+KrBLB7pw4l5divKz1S6D
4m0gSAh+wcbnvC4P5hkbOhDOZ9G00IEpqgYHlRN8IyeMBsP7Tgr/3Bhm/Sd2IgkYaTghVzfL7CE/
Q5SzyvulcluHk6rjNkxu+HPq8eO7K1vrepe18CK3ewqShMsHQ0ydOVUdjmumffMSJIiH3B+6pGiV
nKVBwwZWpUIeTUuV+EkCHm7rvZ+xMj6gC2KEaA0xnfAh9j0+ifOfVJ5JesrP8WpiBk8dv+ZqTWOk
3yWjFIC+4gXcmf3rwSi9tKifM0fQDUNkX00nVQawl+6yPPYgNIdM+vhsiY7kglf2h/7sTsj0+oNL
Ek7CDgiwUOUq2qFPw7uKR6bApaJbJCF3k9kA1l97BfZgUJ7wQ4rP/lLGwb7tfOVhIuwhlWdADp58
jKNl5i8fbnWbJpUzjRUbO4fFKyZesbW5iRDn7ALmy6Sq6IjYTyHoldp0Ln55MA+sP+KxgRz6pVpl
5jcy0yOzBVLW0l5oIoqD2kCXjFQ76ZI/KXEIfJYU/82pfyXWgtVChjEpJcNrZQdiYpcx6ZR9Ou0e
FIkCgQdCYq/1ytAWGaNxXFKIYVwcjhU+Db7RkwO+/yO+qfymJOLxUMyORVKCt1xz9m4m5dSnV9Dq
PEhq5BIWD05qnxffKi+YsGD7jgMmdObIbc6CKyS7Oeh+GZ2aB8LCIXO4bBUBapUC7oM0LOcv0MXZ
hD041El53WKAFOqx5YlCvCrvoP8GleSBs/N+Yv0GLfWJJMJ4327jbq5vOCBpaMxMHy+HTMx4aXiA
ZHC1dyw46ZoZ1uwY/wBl2dvvq14kbs9dlxjrqzswjl/ptGYo0J389FZwmZDz0Et9CM84HM9H7kZT
7g2aIPrSvDmEjn/s2yAv7W0a8ZnYkcRIrHCI3b8oZYyQ0HJpMybhJkN37nQp5hRHV0pOpWgewIoH
ANC0eyibuJ1h2VRfHEuhnuYrCuVk3OVxtb5FqmS0PP7+AJmbY1GEyuhbCdQcuhSG1SbXMadeMsb/
hLorwmCbkf+mv2Vs3kfKPhC4eeICZa3rT1Yu9UYuCHVfpxODW/lkg4cemLmEdoFFmoXgVWuBjCkF
pBETMPrxOmlCpANc8OUawxU0oWpcwnKH0/wWprkAqcHDmakXxi9FWpig306vU+jDVLBYS4PQ3dAZ
yUb+hNAWLlg1EC4R6EDhv5XlvIY8dknHZFeHsVDBlWzG8s95+A/4G4T/YR5P99+Z6XK+7dT0jfHv
kHmEmwdalAJwC85BkrbqWJdvh1ueyvLQTFBuguFcUFm7nDfveL5QEW++hQ8dBYabZmyK4W+ReYio
f9VzPzpwHD2fUAOYej1+iyaIr6+09Qv+B9kodDdaslTRy+ptfXpMY4BOJ24ZJEKRgwuikm19W58C
AGIZkaF0Y6oiKlzii/VOVi1zAO9jRdgLbHxvPZoomf86L8Gyf2vklEvpktQPdmKAIj9HrMpXUFDF
IJtQPHri9G+HTRMMy3aZyxurbpcNWjb8lgR3KyBz3mYGhK11uESu+KoTDOA1qzRc0SEGdi35qRSa
eBVOUyd4ZO1xK81RO8Qezf9spDA1FOGz+O7u6cJF3VV/IIiZWFgTfpImbjO1CVWKD3+30qrvQLni
AXVseympYmkSQ0ojts5sn4AyVg/aSAhkKWbwKzEyECRUtPNNzjE+h10/SJHxNiPNrZA2fwntTJOg
fXHSfssO4TK0/w0+RX+DAx/EGyi4rwM8PQS06NdtG520QJ5uv+IGD0ah0YAYmuTv+vjcJAW+o3YS
ZtSSFIBXjf8a+uVKM52cmL1xDwel6aAmbVIJ2Wb9xfeLKP1V+4jNtm1G7cQIV/FxIdm3h60ci7S2
MNoDKH6Hv2qTslm1GQR98s0CEyH2cjqFdlb9TJ0R5iFdHbtXwNt5AC9TpLEPGEkTaJAhPZA69XOo
5Qy6iUIkE2t58KD2y9luVGao4fHHcC8VcjdrghIdn3FmQgZJF4USSP++V4xEYJLmLizu024st23E
48y5N8/m8g8TZ6Kn7L66H5FFv0zKArvH/XjVSUI+p6ClDU3VQNJrx2cOfRXpx9jq+Scdt68jkh/r
GdOoSIZYvVL2pbR2lJ2kUgDBSWu9n7WVwh7fwb1VBqBqJNP4ACgVpDkDZ/dnLyIqySGbhP+zAO2r
YzGlOzOXORJ6xsi7TlSSAVqz5CV5ZB9f8cSrdBRWbOZfzqReopKoRpsAEk3Ni2YyPBeV8RbfA7jm
gAGb4bnVTemnRSJoiu6Sxonpyk7CRNgvWfyRa9QkWKg/D9QJORF3PZl8UIQemSBQTOLTuxbcDB2x
Nxkem8gLEzjZ+RFvBrpzW3VPCHsM8cE2W98fOV4bNDUg3G9YayHK6KZiq8OwW2SCP8Tl6a8bh+4t
Nl5LxuizKR+7qJ7nk+bP/Krb9fyJqEGUKzl7P3zduBMwxvNJasr5tBT8I5EfOCdXv9EOpSn/WJHO
tycPVNtIfT1BdYZTcxoMAgro7LJPoCK/+6v2EHiUyNWybzHA6Vos3W9zFa7Ve5d+DdVY6cCm4IIN
WlBwk1trRz9nA9tY+r177OnVJP8sZ/TScdLyPamIwJvwlBw3Hnq4Axi6nFHyBq/BEIDkLgFPKXR9
Bc1r4DErlOwL1wmm8jdTCcgdqyLfUi/km8WR6EH+Wq3QDGD10Hc24wgIwXUVvzq49gqyGT9n48IP
OhyPbEcBupE9z0PvBmCjfls/QrkTd282rDRk26SeLcrwgdXRhAFDo5k98s5LdrmTAS2acQ6wq0Ka
AwY68ZftVr3HwvlhL9uJr6Piyfh5orCschmJ/+I+jTQBmtrM99ir6I/0dghBW+s6B0UcVugj+yiK
+36BNApLpP0U5+ktDXuv/WeZEBZVfzoNOWA97ptUYvLyNWKZYtzEPoRw0KwiGuVDSp1X1Of8Yprh
ijsErdQKZJ3lg1uEDUC37XY9pv5sLSJZ29/nha9WbCBWpIGR68Gha43HUi49+TLbLgzYBeuhg69l
92QeX+28lOuFvXjAwQw3Ga2t44kXvPBTrr/liYiMJ7KPBBOHAtSZM/jBZR2gFNekeRhPhGs9TPJB
cydn99AA/CkpgTf0JPhVz0EobDBkq3zv6yyhFD1Xa0wd3h5EHf4bvfXXFFGC0Y1P8ypF8zNXDCTa
PJiQr6z0SWBkYu75t9uCcl8knj078iNXjjhANaUed0t9gMMsPKkcPTpXj8L5AKc1J8x83LGrX41m
JwWw5MSj3BEAMxalS24+iBYtApMqH/3bWE4wcmsKG6l8yZCI0aVKh8xmGk8K6QOl+MrQLB0e4QHP
lhDVZ4bxUFLbpYH7pnK9M4wonNFGmR2AgnoeO8WxlAaSTCFoMv9Z5l/CtGnfySMQRiN83Jam0o6y
M2iEYUzedZQM3M6U7ts8W46U64nzTvkzSbH5E4sMVmdC39nJUhO9OyPZChZJcE8PoaB7MJlTxvR0
wI79HJlRQ04gTQVf8Ylw+lZ/GUT2Tn8ZDDWLzqGEqtGWMVNFP3cEg4YkcCjbA/8BS0T3CsqmgKEq
N1t2nrVcqxGI+FzpiBoB/Ivt29ox7gUdmJ87giVGmhcqoYH9lIw1jZa6d0C6+M6M7uQD3bObcPha
C96WfB7g812MPrE8/vKhPHCKYSidoNgwBKA8QeEkkAw0elyQ6ZvD5M3eHFUwTGDHsYmjbHp6oBWu
7AHTzc3cFCHC5OPqVs69Ge/sdCp3ynfDwiMcZjKOrgQ99q/0AemHzaSmHsL9eVDf2aj5w3edKdtG
qBQ5vMpDCnw45+L8N2PJVleaFaVba86EFmtAdFTzhblEGWB8DdUtTpcBaVu+0nzGw+439EzU8rgS
1LLssNOcHN96TJNpkg5Lr40+8RFirS9MeJrS/f8K1bfUisU0IZ1MWbBj14KD9+0suKGdgsmRIeg1
vcigo4oapFEDVCtLQOocOosHnrJ8geRx1KRDGGPPqJlQ23La0WF8udYPsf+eRJnEy53ldvGKqY78
3Ggrq4NRETtUAjjGn1EiDzVAaHwqtHajWrB3ZSCZaB9yfty70wkIF0MLKN7WarXghfoLNdzC2mqJ
1YpG5EpaHDZ25w8DpQ5CwBKjRPa7Gb1rbZNHmsdlIJT2PzsZeFwIFo6TT09hmeU24xQmv/2M631k
KOP+Suf5a2Qcc39zN+B+vAmd6sZu7G+ig1nyDHJ0fZviImppo1MhWC/5igi3gDY5N0D1RRee1yMV
Q+GOpEPLLilxIWFLERUR2cQh9GXZ1/4pm+xPwMTTfj4NjGeTlm+YgLG05YjZBmx2itlWldKujELe
jESzxpnEC+2atxGnLR4PFryQa2u6RXMnCQMAEFWdkByflXSzEyESm/yvCJvn0hgA2AAGgg5caMLZ
2jtBwRXivrGuLGEqtvsT3WLAIbB08hJiWKYjwqtBl4fBERFBaoyWE/wvZcNlliIhTOI1pLvLflTN
ENf+zrWwP4xYshvJ+/5vEiY9JVLJVHwLd1UGy+rT6dPL0pVWFLAuCEf5BnxIk6rrP5qrSMDDhmFN
BwVQ5UoluBgrUtJp9pXBF3uNcV1xpzJo+W3UsChmL7FqAnZ50XHF9f24UPbGJ92JB80hhLybE7K+
5gbaRYqag5bQVoJHznvtS4YW12+5FcMKM9s7y0EjUPlWwfSHAZUS6sVGN3Re+bGVEv7i+asu8VPG
/2X2zHpRMLZVoOXEUe0cNgdI8uU0/TiuIM3xDyM9e6n/5p2M0w1KTkgdhZymBrgVG5i9H/0Wullj
qBQhG4hzXvuUUBzCBvU3LPbnxfejAK29F19TEmiPmQb3qLTE+RO5tiZzdEzVTuc/WijcA77YiY+V
WUdgmJALuCQz39PSDI4XKDZwFv4noNqadP5z7Ko2bWX1TCrsI5fSKU0mzbgtrBHTjxnmGK3pgb6c
DgyaZ2LtbYkRZcXFqArN0VACvsI9gDMrTx3LwdtSGJdunEWEhLKAfzua0+qmKnv7yNUEYhiaSxSK
Dif51L4EjJ+qXP3WcWwMX/4kILExY42qNq2t3k5Ae1PSHsBXg6fG3GNwSw32Ip+Ncw4SL3tIw5Z8
T7wDvDiczQUC70YX4XbZCAf7WNJh6UJeBy9/yuqlajNgbBwL/KFzkuiYDRiS7u3rZXXdond3cSm6
aU2Aj/AF0uJ2QYgwk4XOjn1kWNWa9pGlAvb5dEqVpxgVxhAZ9ZVOkujqgm0BabqwGLmr49HeYNdj
Wnn2qo5B+bEmA9UnPklJFRF4YoF2Diz4QG946um/auAaskF4CaGoaghmRe8owPna8yIXQBdI/RFo
45Vzp4X7gHSP+oN3nRGOl/owlcZC3GwKZsYEM+Hb1jfrx9dThaK71RgXCyHe6YxTsaMs7jbpr6Z3
KyN7HB+IC4aNirvPJQCRpmVwRAfzZc2sVkVqP/r+bAaQC38uVoYmK6KAPR3LQdGXa+wNH+qV/G9G
hgcRAyRyDT56LG1oH5+5lc1wrq/Psmg221p13W3sgIUOJ9ACcFTgUZIbi6YRznb58nF/Wn37fv+S
HkwbK0bgb+7UI9KDbohIBUuneuQHg7U89/IKyYGPh1bVhwodJXi9qZjxFOrkOVz4lGg8dzLFsN25
xxGRfchm2VQxfj1+HJY0GO6j/L3pVZAidJxjrf1ia7V/Pg5zE9w5TKzamINKygO6PLaNTgvrx3ZQ
sJMcZBNInSyECcc1NZYiWoi5s4Su5ckQWYIAvYCdxDkkR8aIm5RDY1aAB6q6J/Up+stR0YhH6jt/
M5znBElFJyrb6Y9o2nJKW/CwNnQANVEeRHfw9zwLRIeA9a3hNxQGhPtxQXEKmIEKZvpPqYhR6PuY
DGX9g4lee0SvF+fjv3hey3Gr+NcreBVPwXn7o2YATKuhUlrZVxD/u/1p9lTryXMO64Q4lq6LUAl3
fM3Y4rpKYf5xrVbpf/guVfg8uXDQh66GgFtdrEEwm15z3vseeXso/rG6vA4ZBja359oTQ4BwQ33t
JaG2FfutWY5uJJz3Ayf2X08oxQ8xOg1VMIQ8OYfszi17IVu5eVlmTyy2wjn1QMD4hlvp4ze/iED6
5PIoK5EUyZcbKDZGwUEztHvpIHaXwMrm9jeyxoGONly+e4AXDRyId1F13vWlO0ohxhXP+tSsuxZt
PghQbIOOF0l8pyoM5swn+DE5Rvf0vG/5eIVf0beNzqd5/kHggoKgxR/NUqLnuoKmyBaZHYHoTxvF
IxIm4TKpPd6yGNE3sf8TiPwzj1m6LrM2HeBEe2I6ZbciIp5KCqpaeeDr3wHn1T6TEpg00n8/qOmv
Fmh50ywnJaoy4ljBtBuIiB1loLMtzv44jJYH/v6ASiABUSHtjTTe3Hsgv8JszoVeQTsbWhR8lS6h
jiuoQ6wpEQ1M0zwik+ObUv6quMRbaiMAZy4Vd9+9bB3P0uAuv2UGyp4vb+ok9pwFJnHyshoc2kUC
CxXFxmlfMYf/95IGu5xhAlN2Pk+bUFhIYN4pQvaMN/hY8kxgVAcWbrbd3RjKYAOZLs4u9XChyft/
LdmdPN10JTXWPExpyODIhLSLYZ8czU89TCqhzNw9civ8LP5m5gIWTTM6IOqO7oV91hr0kHDuGAE7
d19Gs8tcuGh+uGr5sOrnuaAu+CTvTxdNT2Q0hj8vrZOhl7+HLfaimJfOECgpg37vDDRSgdLs9M9T
Y6RQ1pAicEF6E3mBMuTi36d7JDF+A5fck2WeEd7Xy8PaMGgkLxkeLGRY50ed09sGa5ONxk85s2wy
uhhy7QN++PVpedOcEU3a3f2UGheWeH0yuXSmXcCmB9GE1C0iea07dEtQRITEy3QBwMjdV4DSlQuk
mx9zzak74Em5kq7sQ1ejngQgXiDZiEoH5K5TeVriAFdw/D0ZpLs5oWmOUGTX+YkPHeilcFCl6u9x
D+gIhA8oN5EOHsLTbDavBcdGCFegPFGyc2TPDitqBxMBCNTR270ofUBcI9ttmLpQH+mPC/7+lH/v
lC2a0gzdI6MdoE9CtW6zZyq9N5wN+ZUDRtEZ2OOas7oQvoL7GoF+yn1SxVJps7/+OJ7JkhSVWWqS
EPEwEZ9w4dUk7op6bXOPX/+JhhVHTsrEgOkWONfX5XVb1jXvtz9QjCojQ6LmJ7PkJ9bwR/44hirr
/ZgLnbkiPpV2QBoBj+hzpLaR40CrIIZksBoA4cyDeUp8hCtt1CvnDZ0/2/8rx5Y1fRNWWu+vG/It
LohIeppfo0+eT7nlkQnC2gY4uFIy3M7oIQ2VSerzrvm6RzxHevRn4Hnoksaebp0Xb+jPd3BM09V9
MyrtYYOqBCrR+ybGP5iVRpOw+8GkuUsN9TQn+FyEWNOTpGcPsIeWxv4G6KIoFrQ4UuzOHVmyu/9O
cibs5TS4VFVJNWavpxt0z/ja0iRfG+A6qMluYVZki/RwbFhBrKGoB2JZtKmzS6FwFzg/dgSW+7Qj
IBRvbl9DIEulZWk+L5jaTeLoNaAqd3gNtRDbVwW+V0vgElbhQBL3BnYuQOP5THqv3IqoJf2CMOWI
mpcUNsJEJWaitgRmlc8zDn+LBOWSGq773qd4ff+tP5wCyGfJX21hYmhZiyDIN4QdCvD0rEwBcDOT
UcSM69dKXdiOxqtUwJ9Yw8UUeog9+ZV+i+f6lIXvwMIRqM554e1fdNF5lg7mRYh8Mp3es9zn1TeB
fiOmSqCD+SZndXiIGCL8vVCp7nai96Sk4wK1jC5f7oYOQALHoRlku48zvKWVdy9/jQr9euceC2/8
79XNzkVXyPbJXnCucu3BBatv8eDvWYFE22Soj0qiBbwk9rl2NqKZi8l05ZmwKlNP8iXQI0T9xtTi
QYReUmu7lBizytEWMu4TAB90JpowE+RPUP70qOuthFmvAyCqPrUnLUAtKIUNly3DrpB1tFCVKiRf
ZAA6DIq1vRPWgBUv79Bh6nEUtTDF5xWCvpG4kuZJtsQVf6tDkn42lRoYn82jAwLDtavpkpATo7gp
qy6w+xEfO07gh4GJImGg6U1cqtK90pSst33T28YMDHEXG9rBrCYKRbpuM3AAfjlIpGwReWB+GJYQ
MCJaf6qF5ICPDz9OnOLyx9XihdcaR0mgHeJYGTxuPudyZenXRuzDqSQICOb6iVmy0LObEEBjT5Ar
3bTWukgsdQfijq8rG91VfUibiO0PeR68FOJ1bmGhib6sk401w44YrmnRimCsTJ56+PAFi0y6leWH
paJh9lB16XVwVN+kHiOwmuhyRwWZ0LCV8siqYH/m7z152WxFJtQVB/c98euRGE3GHDm9MqEXnYTd
CRMwAW2k4HkDstY5OlhvGTZFZfPaUJ6Q/h+OzdaAEkUUEvtl3g1tpbq2Re+9MTgk2KRHEv6ESXqw
YlvoTHdhpp4kxRzIJpbMsIMjkZjScyx2zZM3zZvmn8hFmVWhjyFrtEuR/GnBYwo+XoiWZkpG6EQH
xpiYCOlVcrYI7xGyXChdkGW2RzKRNpPHmGmZ3Q/3Ov9GnZFHwrss9kKcRWTKzmeu7gzW1gdEEy/f
SmTZC6G03PoPdNx/BN3qheP3hRoCYmFdTRqqDh3QM9kS8k3Mb4o1k0dIGuJElAVhjbz+oqoJdnOK
Ffg4NkEWNVrgQfXGRBRsvvzGcVgSlEDtPeXbS4mZY9XOftSyoLDCglbrPhM5fiwdF/abFV2dYXeA
hd7a12ADcxz8QvcIm+WaELsdaZ675pCAVY/PJjKWP2hZDaUP+TJvZfUGrfMppwLyq4mO19JQQ6DJ
SNhJ19A1oNQURrSe7KJSuzbwFt79cwPdmmBDYfOTohIc4ojH5Jk29+dKgXL0R9hIyUShrtopGwQ9
r4rnLePMTi1+dasnF4AA0v53QGUHYoa1guMa/XPcNPp28cG5VsyrnOgX65/MnMkN1fkw+3zS/7FF
U5MVwy9m2w5ypmWVRB1iBFvRopsajbWQApGZG4bFnwqCiwRsGnU5zNttaijI0lwM9y2IE3BzWUwp
5gjjEWyKB+26iVngy+ZG8gpHzndAAFtf7qvpTa8ZwZG/YmI0CdLfb1ENSuG5nBwe04j3iAr4e0M/
6eisIL+OCu5cBsHBol3+r7UEBLmMugYtkQ7a8J0uTzY6tsKzaTTy+ONvT7qFlyraZ+Trs30Qqnij
FiDR+7IZahS8VNQ4W1qKVsqOJCQ47+ZcOH9e/izG4vEW/vjQS3TSYz1b383ImwLkfNso+MGb+8Ml
J9gdi7L197qjmgHiQsJtEi6TRmzrWiy68WUZEam9I+RhMhYKdX+kurHT/YhE6B1Rojc2A7UbDj/b
F2TeYDyPzeTy15OqWn+Fj1VOwYaIV16lyoC6f78H/R4zhAhuMI/37lNMpq0ufnq6KSIFUUmYKaAv
VdCjWEFrHAWR2uFbC1p8K2BzJLEzKVeTyWPEZ3mnC6txa/gv7U3w2Fiv0MbvgQ9NIvzcaN/O24Zb
2BJXf7xrDI9UqIsiaLGiJL2P0d9yL7BNLd82XU+inh4/xa5UP+ZBBsBRYqricO3qsohf+7eQ5cWl
BwTF8KD4TCQWNIO89wr+5Svv1jUvEJSfuRukqHj1dvpNDZxUn7dVp9wtGfO7LMvr6C7WjjQjHEU2
PZhJu6kPxI+eDh7uLmrBfJmvxLNSrhbB1r7lj3b2mi0Gz/NVUJgwYYRTrQQY5KXVLfBRJTtgL2wO
tFqFAhzUlO70TPTyF24AEGibaBWW518Azm8RZ3syVvlrPCqmPI4QkNSsGu4m1YNGFxYitoouBB0/
WaMNO1x0a/JuER4l+6T/CbTo62TT6IjlMT3LDcMbHiOcfCXJl88Pvn6Rb3KtPys+VYc2ie9SxHEl
GBGF1QrvuSniunVBG5kpugVfdGL+agxn8uyVDYIQ3t6mBxRifnvdTikzu8q3CsNgSQce5P6jRNDp
0hHEE4e0NGd1FOxvnLJl8a+MSLkt9b4PJJlAvhCZQ6hrV9492YAPWe93uMI9r0w2U6ri85YheoyR
SM7Vh5DlucQlmQsYIh4DJ0rPaOwi3DEmVePHg8uZ+oHrgdyvbpqdKjEopq2RKk0N9xmR0+6gJ4Sd
meMuq/2ESasfrt2BrbiCpBEkdy9CPjYMjmw0V/PaNxLZGVtFEGIEsdoAryPBJJyBcUofJOVdTArZ
OHWYI8iHouPwcVoXKsqxg/8S3G3rPok0j7SoWTcc3IiZlAbsootBGwfWJ/I308xUH3iy8Rqozujr
3PGh9yhaJVphwh4i63uo2ySKyjZqolT2CZrEcwnhmVXmAxMmUjpGVfI4l+UzzSGSbWBSEhaYGiU2
NB77NIqMZAlBKwzJkLybd3UPoYfWTgYq2eljy5NmbwX1oDSq9QxA4vIsLWs4OHylU4cZIfuDqQj7
k0CBMpUJkdxirqDqNEYz+018IvFKvuF7/eje25kTARlvAEIxiMPZGr0+yD5w1nwIhU5LBIvZcPXD
dYlmjOXpefRd5gffVqLRWo0Bs/QQCjml7FAffX94JYRUrxdu07Qkd+5UXhrFGGv1zVFyYDYkJfF7
4Y3mN9pX+gg++HF3Kw4xjNXJDCQoKcMcYg/Ibfr1+EQDhD58kPppRo9V6Ce4IdBebQjSVgdmQznj
zoqolLxxfrtCt1+avXUOshFvCjNaaCceewsIp3zaVk6l/ttXeqapocusenDsODvENvfdIgW4g18D
ZCl/aOB9epYjInEUMeznVwZwV8bPzYuxumzqAyAMbgWQsVhMDOfm3G/iIGrzc5zawo14iHC6Yw6w
TN/9zkHKUiO9ldz/oTFiIY4b2x37axl+ZPqLkXxi8IYf4f1wMC2Ip0HBlYh8Bj6fFjocptYLZQrS
G/eCgkNOKHdgdl4LxvSVX8VItzTVwudbWOoiS/nVf5dDU4rpen9kK5fyfo+JmLt0EH3c5kzjxaMZ
UwJgeKz9rfyDVbXBJVsy4eDOyM/E4s3QpNSbf93VCSpFBQFE2rdzaSAc9DulX9MggltiBbyDeNUQ
3+4XhC8XauH+PoSZbZxqESVYjvBLjaquPMr4n6LXPKPoKi6uLT+Y8DAD0NKYSIV2kZsVD/QVW8il
sh29H788I4vAlbxRdrVAr3jwHN4Xba+6QWGLTWouMG32f/beqzRDxqBbK7aSBdx+kHSOU+im7GPG
6oOkkpnYlzGQO3AWsSzSdfIg2EhO7QiFQ2Zi1j2+eN8QxOXIL1C+aLLXlQzkrNaC+b9GXoFmvjBU
hCM3UpgZFTqlWdULtSNXb0hFZk2oNZ6MoyIqx0U+afKEIKUVKE13TUlilPK4XNRCW0qf4Wo2j625
Pk5CM17XpQf0LTrS4q9g4fsgU4ydoisl+28+BdZWOG6s4jspG+MyLRIF0l2gaPVWIxYWKN1gMm8b
zwxllACPebOhT7rYagJYZIpuqjSPc4hBGxzCyLcqIYm9rsdnR4ehiIKbuVUguEFm69fPmYAkaxPz
7XPsw46/z+AF2Ab8kDGv6dgrm2W/Yo7q1IfKspIUmzowT8EZxDOzsI45WK1DYRv6+YusQ8sCX+Hd
SHrwS9rg+npc+BWujjziPm6otjeaiypxxA1u/cgo/v+sru0Obq6MK3Z2y5IcRh3QCu36GiplMH8A
lIKSmYWSXrBqF7B6smxsoQJfspxLgcG8WbkAruS1sNrFYfIY5kIKdVJbneMgmHRYQ6/7AblpLYEn
7thfr853w8DrUlVp6y5+eYPBqbfn+29NwpZrk4IXd7TUAhqNXH0qVh4mF7pOKOHIdyLkapdCILLt
jNh1MOyTAPZ+ncTyxszLN/4Dlpo7F4IQ+c9aEB5nNK7ZeuMtNeTTgXluUnQMY1tZgpU5O+NgWxAk
cRcXi8mJA59YGHYcIYUv1+caExvia1Ee64GcEW4qkaLRLJnc7FUm/w8dfwKF7iK+DbmOMwflRHLH
a/zfl571aLxp6qOlMrNzhhB97Kmefk2QvK/6nlMFfPeXsKor/j0Pf+ASaj3BAs5KfVV5OU7ktPsh
OMvy1UGNApLKqqUGU5FrCXOqP/R715Z354zu+lxDkKPo1ariu0jhABDAP1pJctgqxeEhlnuI9EoY
Verq6Yu44ATWf7sXCM/dFOTHrT1KPz9o2WKxDDSA5KFtgC1dqo8/xDi2P9NAAfVjtNMD2L0Z+Y+1
ZdISFSUTcvlxi/BNY7+W5k+6L8nx43kS/DL+eQP0OmGUyLgr3VILRftdJMkoejDMzEkeL9Fa3BdD
ieAG0KxmqIGdMMLxuuBSEclVBS/dB26DHjbJFuY2kIYHRuP5MAt3TWQkgXRxFFAyi/lkORlBkoBD
+l8qjuSSgCG/dhpJ0Vn193c8/qMNr80QkY2CNKzFR7bkKwBQ9/OV3KVKhlB/NgAM/nwDrHAHa6NX
UOA/taM7nM1ZonfXcWaV0XcpshUAtJQEYvEUspqR/Kk5zuEJJahzY6g32HYGxjjCvSr4xcLWK1zy
HQKfclmBxbEKttsw9NFHF7visp6wbULuSuiBHa+tvVcQ2xbpaFeVDN365K/Z9dslJtQkjvNFc+3l
GOPFYtnbZgM4yR159rTAFzrN6IuNvoMr1tj0+YF9Z2V5tvTjoIap6798hFGt18UTacFxqBMR7DRw
4TrF0Nu22CztzFKf2POfZ1XbNg2HpvQ+c3lrrCmFcBRPZyGrAveWRVqdMQxUCQTE/oEtPRTO9/ga
XED9JKfnGbqHgby60sYWPoGeuBkH6pesj4reHBs6C8Y1QDPkfb+K5r8QxEXUiCMOZwXbgOhA0aXl
TOwxgjEHY/p5DN1BQck+JaTvsyM4iRuSnboYu6heXkhasR/cJspM35q5/v8ytzifpki+8WuOuUAc
Dlz0KfT10WJLBzG+E7fidWHtVwxE2b5dbe/bYvwGhAMXnRVovobr/qMPtBR+HPeLyWBLKt39w+7g
BUIO4GZSeHIepQfH/QbtXsJl7A7FY37wn3t0TX64HDXMi89ui8pkB494yyE2hCH+lpGoouYMIuLY
0KNM6dm6ZpZiXafmbT+8aXDmAEYcQysUxf7fHYBlT7SjkELf87hRnoUQEWkVL8cKh7p8kbPOL32b
s1CdyWyrLpxY3Pu7VA4mcy+VnmUh8iqDTmM9F9oiPkyivgndDia2zh46elN7/pKokFOHxEtiBBRf
7m9U2UuBuSd9Pe4bCOfOu9PEGt6quTMSOiP0gT9e4BFF2cMVfBsgQfZOpENNZE4ajM5TYZddK1hp
OXIWa4yp94YjDaapJXkQJfgrui1IkHHXaR8muYZ6HpA1sO3za3Mofn/GqzL5vXqIEN0DoF2eZLOF
6YVIyG8Y5GOBIWnpc2hIt3yTofnd5SVJpE2xA+h7O/4T0aD33zG7D21QI9GRwQSKQJYfg4OtV6t2
qXZWwdcnu8QwUaRUMCfLq2ZBplljnftYrrqsTaWV/kaK6slW7kiSZWhLfHszbkViLAJ4j/BexQNT
rK5nMRxJLsnVIwpCIV1muQybk1JATHqNL8UuXFC+80KyPVZ9Le/wsai9Ewvk/rx9QUQ1FN+gHuSn
nE38pfrJ/Xr6Zjav5K3myuKwZfU+TkYVH+ytTAUIbU1TVfcpznhJIUHB0bPAsd6vSW5DwgAS4p3D
Lv6AP8ekdDeYE3vhz4LYoQYnaJ2dV62TTeTuOBFxxU0S+KwqGfiVNQDIiurIcRoBs3gOZ/JkQ9UX
XBdng/nqx6q0BH1HSXZkAr+VDUyJcS2aRf0o31J487YiXyGmZ89/xGaUCPsZUO6m/4TabwoCc+L6
UkwJYh8UfaXyyZ0w2IffQcknwWuSKg2oQozdUFhacmaOvpES0R0DC7MPyHSfuHsKCEb6Qa8nNrjK
FXDpXLHRrNPBdYHonumVpVtn0vQmu+z698bJIBFUc0acrFXgFCMI11JvuEc8RRuUc+IsPu4qhkys
RyB3I3g3WVR8HdqAHTeXcBdGVjGUhDwaFt68RkvJQStHMzd8RVOw1/lxzwAZ8IWGHsidr68NUPLu
cJUPvaW5dgr0Ed3ISMvxKat6/jN30+H39Y358RE3wzSS5gTOcqIonmfWn6rDgBY+wrR1xnS65ajb
9xayNGwYx0Qob62gozRb+FepocBMZgIkoJiHkKCj/QO9fE+4hEvGv+BaOiRNMhBJfU0A26JrXFd7
gk6QX2fDgTLkecVlPvkC5by6Lm6H2XczBnM84L0TmMN67R1I4/erLKLUePV4lYA6tv8rcxKQa13B
UxhzhI7Vl3EkIzPwaYWUELERRuR4HternDuL0uOv6cuabE09zZNoI4SlWcB5bHCK1ae7/0BfyrSI
dc45nGJRdvUGEJGQfLv27eWlMqo7ogRtQn48nnXCWq3IE4ooexq21lMyjITLmdqGtQeEYoOw882e
tI5Bb40A2jnSZ/teEboeMfdRi7g9VAoY7bZxVzFPgW3xr+U0HGd+sJplocWOzJcb3v/JXuchq8a8
DyzIobfLvmuyAW6jFIM+7U784fzlg3H29vZJ27htuO5AOpOBCWjfoJ78zpe4h0FclVSUsJL8t3K8
Qj/8y2mmDjmZdYE53omhsgbPoGm8tr7PRkpAtjTi/ICyj1nIO18PClArXddEY8zyUUOCO1PBoJbm
k621JVz51F8l8MGmuAmAkrR5GjbqYfwqdv/XI911Tn21UmjQpIJLK22vmZnwujRZiUo3XYx/VRVg
R5Si7uXJWHd1LnB0FdGr3r0L1RHzfBOvQqHDkxPZtvRGAW9Lp0MoMIPbygBYs4DaxYOIN/4S+Iri
H0pdpdjGk8QfwT+edW+/6csKdKiLV+OXz5Og+8SgoKjanxe/wNgj4Z+X6QwwVpH9g0gHYvnJnxt9
ZoMhm5Wk1uu6puSdwG6YOI4+UyAQby9UmJ50EStbF7uQsHo4IO16kN6a7uSu1TOfgjeZx7sAR40n
GvHDfMjMzmCTbahI11AyEBHMN8y0kq+MwVWE1h1ib1MV6mbSfdZrGUckGFgxtYN2zmUvazoOdI+t
XgqInTMRBIHsBw4MyjIt+eHkgwakIwypYyzsUI3oW7W2gNJRvBKyHrihPgVppOdh9AMyE2q1Xi22
e8ckdkv4mzXeSLIv25sRRkl2K8fQbxt1B7ns+8648ostUqjGSiDJ8PKJUmZSeOB8avwd7OtUey+A
QRBDR6tGqF6Z22b+us7/p3UXi1H4ieUG6RhD6+ZzRLu+Iml3wUkFt6O8FN/swcDk0jihI7agHy/Q
7IanfY0YweFSvq8TwRTPps+zNOpqqSmUmSTlQMWJFpRmJWvLQmGfNFrFE2yQyRpeLq5sWWehxfOW
svN2HiqhuMPStOek9vcYkv+4iqdH0qGK/vONdJSNMktaEu8ZioIZc7lJ4Zod+V9lcyZhSFcahx0X
sw2L+fEkRKGWiliczj6l2RwfQLXOInfu/+SLY4O411qZ1Vl5KyyyRnaTsRXK4X4PceeCPjUGVrKJ
7cdyiyFt8j2L70tbSlb+mnOu/oC349y5lY0d6sRFCPIy5xhCoD2j7DdHbsUJUW8K5hZZJvKBtmbD
ijL92qRgC8A938epx1DwPObT8iyCopbYHgUVj7RwnjrFpbbyoI/ip2chGkAeOragLeK+K3B/ndEr
MILzEaJ7wG12yJY+34Y5T4JALLks841+cWhE7l2W2WK97w1GnMTLGy3/cdr3MOom7pUzZC+4Jv6z
gJ7YeNpxcf2iqsYh6gcTGTJ5kmGnjU0S4NZzagPJodydcfFNI9e/Z+VGfDSJzP56EYKd1cLZvuCn
eyIMWYsO/h8nvjM9PBNE6dijZTeFGmUHlaS31S4tHoDHpOLjhekq54V8wZ+obnTok888VipyLynN
RVRQK1zuXCqodOBIZYVR188d+QK5Mjk7xD7uZDet8kJXQz8NvHuPmsg9V3XmdRF3SGv9USg8mmqj
YgpK7sb7VzQ4Lg9L8oKtFQPMF35NbDo36W/DdTeudXDa3CJ8zq6NY3YIwNwwKd+sIFyC0M02Ul3v
l8SHdvBcg+fgMxCcwEeavQCJNU48nE/aLbl7VhfFG/pq0ntn/smCunFvyIuYiDNbJlcFfknuUr7f
pgx4XG8T4hLstjaj0SVq7NHHdfetS3jJoaOIhDMlj8N4LO38ZSxgtJxwgzp33UXJSdOmnub0PqRc
xdlAmtJcpbV5nxnJOAOw3PASQMOaHw4dAmvT1OlxmFQz5OHYkBzpfQs0ZdNPPCbnH0v0TwWwKf1J
cg9dC+PSeFPYfrVna4FStvoks69H9coP7I2olPHi4Jvhc2sD9WLQNZwYmnuAWmpmoU65CoxDMWYa
eRUxw0OjT03/rXVHzLLzxGfEcF92BCrV8qOOL+iokQ140sJPQ8fLjPesWwsG4CeZLU4LZgeddjDH
bpdwLdJA699XxtLcd5NYdTgGaIqrik5XmfNNPETAnNwheI8gZJpfyl1BE6L0GZdd0nYcJq01zMZv
zFgKIkNGZ+HQp7qx5S9nAUbyyK5KJsYRbFfAu7e3f6g5FKY4uge9PpN+IzJ7Tw7wpz5zmcSiLOMu
URPUlTD4IgA2j2J0PSvLeuMmfVS5mFkJQDDE2ROlFJH1GGG4TRoLQvyyR9BXbU8+Qb9p0hNprjdv
dTvdVRd4cHOM4THf2P27DR21cM+BfJs/gF9znW/VUYIeUecKpuKJP+dX0iPkLmlb8XS/Bwu37sOW
NqtXGT2V4wVzf1SnzGvHNL9JJ4QhN2fxb/zLuRgea07s+JcnKWDOGG4kglFUhVTrWZB/V11Kx+ou
3sqSx4VvO5uivkrOS1w1DXavDTtxtPvLP9tH/aclaGB/WzqI+dW+6Ac/n1SgbOOH/W+onP7P9WxN
4/RDEyY5YOT459SKG9o+vGiIDRkd8CwZvteMlk5x/X0o+2H3pPUDgsZUw76Es/Gp6Xvo3RX8JROi
mzi8J1i5/djbuSKEb/u/OPQXR844MpLwXz4zHYw86H26e0L12RXqHJAdnyex0lAD5peGPozEAluX
111T0OY266E0XgGPi+sqPZQKulMaoUMNgYBkBblHgzJgC7FEeGzZqWrxkwz/lhGYndX+W+sJ3ZlU
e8VTa8SLBsdTQN6sXffYWBaC88cRtyiqq9xogXszHDdJSJNEcZ00ocfP6lwvfpg0WeKjo6ADrdDT
t0FWqJUsJoGQ+8yxSKA4nNSaLQ0PQu7IVhjBuEZYYg5yskXei4g3HJVdaXbvngBbMuba0Z3Ho5hJ
GqH4TnbdgyJ76iZ84VyN1EhiiM0vOp36SWNdhTgtYNI7TesnJ+SKacUWdmm1XHM5/XGPkza+YSf9
uLh1xBcHfSsc6E0NzYPbVshU5ayisV040lMGsirdpvEgBkFuKT2VommCHF9bvKxcoqOzmOrbJwB0
gSIycZ3/5Ql2GuTgN6vflxrWBtkNk48TECkOlXgE7z2vo/d+ih+vtkxpc8s/+9WLrOJc+78+0qU3
N2LLCDGbWqI+955TT2SL038Ig44eU3jOauUyzha4zDP1YmT5mWttDtdvGp4gr56Hk0z6erjUcZ+h
0Znr7+S81kr5nnFWYyfD1/1IYSr65q+B255CYRHG5Ptdo2if4baXUst4t4C5VdIYTkplTIOW55Qj
5mKgS5RL72S/7qIyrX7M0lTS4X+QS7h3xT5CjcotbaFjrwS+RE/OuzZ0TRiPITZi7fhl9MLiPFlX
JI4eUB4jt0LJuS3gAmC9Y31KFbnymRiNG+ladDwi6YzNJ3ROJwzmH2RAzTtv5nJBFwTC8Tjbya4U
pyf9kXLeSWZ6dwekoT2Wyvi5ci7NHd6aMBHLFJaOf/zdJ6Xvu/P2Sf/ex1TbcCP9gsg9eSn/TBsk
pH8pu3JPEblAaIEf3ySiTBTSJIm+3eFsGQDUCbuG2QOMAF5fr9x464ghvA8xJbhKkVPgC5dCj08O
FZ3GnPpyehPfCtTJvpm+t1P6YzqQqDri0eLti2TOYAlPFAj1EVPV/m7Rt7juwiLbqZv/fdzFiJS0
+c+REzA0mP9F6jqM+Ljjpvhj+vnzEbmDEudrwIncdRcHbmwBN6Nloe33fTU2reeZ1vfGEYbW5NAP
2Pshd9wHpeJFd/rMKQ4a5pfTfeQh/e4+eDQOM6MW1oqIYBUJxAFcEzOJ8gbycoLgglC2LXgTmyC0
Bto6TsgLch3DQq1qKHkvuRw1Zx6mzZFo0aY8Js6EUlMDw2TfmkaJrw/4qUJC7VJEpQV3yHajTrPM
L0Ez4lQmCR3nr8NBUfSo+IB45b8NYtkAutqre2/0PO7AJ3VsrZqOQhD1xpi9iyoEQcZDGirKM1fY
WgIJPH14W68AroNnkXLHlkPmG8K7y2ITEjqWsAyDtfuHHdzmhR6wbwbgFw0VsFFAIHQwF8+MfQJr
YxLID4iM/uUwPht22A1Qb0t2LQyCLsyBq1edaaJ4dlcD4DgXqhNUBMGDbqhSUHXsVxX3GZuh/oll
wcixYzfTu6w2eFWI7Tc+kviIfhOrdQCO+0tdhLjquY8qxvfnG6tdGrUugvQQSGhnckHAi80js6Ub
H+2EfccH558M3dlu8Dlda39cojyYtGpK3TKLjLt6iwehg0bvfF9Yvge2dPOzij8Ach0MP5rrEvAP
jyj9WJS2HF7VGsHsKA6TsmfqUpX8GQ681MvuAtBxHIClqdmhz1WMXys8Ej76aKWJKm2PsUWGS4XW
qv8pmBYCvN/URcqCYPUEAFsvr10//PO3sLFAHlkIHs6rNZJtgDMn9+LyjlIF22m8w+vP4mG9ia/7
x4rNWviOqQMbnbH9HaNBvxv46XU+0/VLtnkleAJ5gzTaDLYUwVF8R8TlaQOD4dem192ZyKIKZhFc
JBx0t6dZHtGbKU1osY+8Z5gqF3009ZFqTCSA8hIpS5rdRMyKwB8Yjz+zSGbgiqTCfdYjpV3t8UrM
f3w3gFrOjSqbJPT6Z5UY3meTvw7tIDZNjMImHLkJ/CZQlMJX+JUkR221cJXV2QI6OWdY2XvUIleq
JeVHbU/RXC07L8yI3nHY8mGSj/H9c4vt2RWeOzti8rQRp/dPAmUL7hGxIrrYOJxAaPGgJWgIS137
e1AKXU566at85NABya4V+4+nh8/t3SbnJVput5NYLnvH6z2d/7achQDRH64R/bGpP1OnRvQ7ufyU
c70nVcDna4sVgG4HCPT5/xvgxCoDoDR+g0BJbNIyQL9Stp/Xm3tjfjEYKW158fKwWCMQFfU2Vbyg
ekN8bXZsPLaPkb2OEJCRZWIG9R8v3WBQL2qPqmj/U1qERsQiYgBHZ1CEU7vKj2xHiDm5Zw9SCwql
jS9UyjAR
`protect end_protected
