-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
L8zgY7qOhN7Lmu45IqKJDW+IhVCBTOKJnxRKXefxOpvoeEsvj0ZmgvFqXv3OUeKYz1dj4dp7b8bN
vE8ISe145eOrRwRK6HGOV39hLEllfx74xH4QpvQGCXYwTsv+h9ExRHy2snk1aMN/6vwX59/fZcAc
wSOpBMloEJTxP3d7WuP7HQfJ1sbpG7XMminSd5X3lUFM/ejJPPUUfaJlr+o8LwveS5QOgZnozm2l
ubE55ruCyC8A9hvniujyGwRl/IvJo8ov3UxbQd9iz7QL9eWJNqNHLqIirINrxgY9fqTjnyRkPWnd
OLjxWcWiTJ/tj4JELSS3hbutZ5cjitgw2YgVPA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 86768)
`protect data_block
Q+Fw8wPB4gq34LBW7Lqbfcr0KsnmxezfZLrAN0p3T9awrJs+qqO2pEVEcib2PqgH8DUPZqYxpP72
kr458N2FxXKAIm9jsdKxBUpyNM60g5Iioj8PhU1FA7rEyKvFUReHGQO/9eiqqPFFvqVGGP0KyNQ0
NeHckmzsZ8f/DE4KeY5b1FaXQzgZpusVfqbXC1gIpYndsK1TCaQTl/hc9bEBpfHnySQp2my+HUVF
pNgZn6HjpNr+RCpFMTSzpROYTvxIj1dv0oZYDU5A4UwA5NAjnPMY4fpOOCFe4jAhtyeiXdDraQ01
KkV7RERczkcRJeLcFjouAJ6QzetnPDhUDZchVhp+UFSVEziLey3l2mgO3Wsh3Y+fvExnt/sCZw5X
MFg6+V9iE3f3sKKpx8Vq/alF4JoEVH5Si6NK0pGBd8C3qOuQWXx+qeIu06vqvJbi7HiWNqjJpTMl
U70x+Hspb8AKYAPXXbURrmf00udlF5/5WEDBMcDa3GjWzE0oslFheIh0oumrjDZ2OnHfA6VlIGI5
2MMsom9fFKvMid//M4qoJcwHhpNy/AYRwI4rs3IG5kZn86wFx6hBQk5JB176YXhY2VAOG4MJtEs2
dNHLV/SB6mkGjpXVJbX7fpVKcYtCsnAOz0MVQhbGohT1qasM6KYvjRnrgo0Vl5BEDQ19jZ+pgGp5
IE8ZFq5sd+6UGO/8fW1zTK14B4l6/4oxKD2p2NBYymksCTS+fbmiotzcSOpFTrpLggIAXXp6bdp2
kiQWTmucqiegNYDdkAI11mxVyJjANNh8uY55wTfkWiRtzwA7ehMXn3D593ewOMRE5IksYjaJsa+T
0RMT6ycZdk0yvaGYE0Ajvh1ZY7BVRHK2TnKJlUmK0VMy8XA5eHONibXSSk8FVW1tMKkJ91nF0wbB
WqK3ntSceDyavI4tpEBHd/l4RI6+y6ZOWe7fukWAS3mecxbifOQUXVB0VvfVrvI7Zr6KY32EYXrR
tbqReo9t/E9qJ2Twh9TyIfKqFQoqueQfN5RJGTXtPblkCZOvCvfT8oP5rwnL+zvG0GCyMaUZC5ng
V8IRF3+vh5AL10vrpUKGQ3qW+rgB3O0hT56h8y3HtqXEyv3/kDHjgWx5tbnQpmfveOcKFx22O4Ii
ksIHdOvbtEm/xpLdGZkRYCCsYnWdrNhSUfG3Ic45vap0nG9rayP8r5+Mve09n3aawmiaEYl+E6Op
C6b8+Hi44l/BTEsltgLuCrlZ2xYH1cQ2eVj8g79G7QoLIX+3sr1NwlOtvC8786WKMrPnb5YOARA/
o7tO/5eXrnfbG87LCq+CKYs28Sut3SkVTVhCyxe+9/fTnf7LgD/kiR7qg2MB+EdFH6OHo81bf3Ey
TplanNViCAlwMCZad4+URTjlmZqs+W5IkcTvgRHq+FhsFSOuqJp7AGFJuP8gtkouxBOd/G0XfSjI
Ww2XD56/irXlHUJ/SuYd7xxNB2NoJthbNrL/kM8wVgaUc07zc02Iu26S21trC+/4I0dbW4LE9Y9z
vq6cOEBrNwPgWQOVgejKUZYH90usaWhishF0TrJe1KMbk4kaVIVXu+7lmAP3F6pxAZn6oYqA92kZ
AC0FVkYMbC+6S2of41nGzMAwiWF+5VEF2vFhWnwfG7cWNWAi8P4KQsHd2x6r7nryAsnTx1nC/cg/
/GAA3ShvNwoosgi64OBThZLuswPc/4tXyBXH1BpGntWi0J0adOZ2z80y+WTond9LjSN6e4POVl+8
29WeUR6tQz8OvaXRvLig0dESG1Q5PGnr+LL+vhmROBmSoRzyStD58M6CY/XsWQk7DId6kxDHLihy
h/d6kRAuQ5kmRO+iOTXoWeKz6YC+4qrFeOt6BIp6Hh8/CigJomy5s8lcCN8xpoqJWBMbiXSRkbm8
Xf4zdh3hlhTxzyxh9lilYjksWxVhP+Lhuxos561dh3J1wcIkZ8wGPoBcDOWQmSrn8YfGlfdOpeV6
/KECLJHAxGMM9mOmZL0n+jo/WFRKkdxaH6+VpUjn+xDvzl3/EBqwOUCDFRqf+7gRtFm+HEAY/lz2
VIdPzJ7JPhPcX0EXRIp1G5yrpiAEouWzRZmw4kJii14lIVJf8o7czCt3plVFIEC/+egydRZ9iJQq
sZUGM+4ukf0F8FuM1XisgkOdFH5ZkiRChRGAOJhsxdu5z6y3Owa5IXsl3rSA7H+d6GPLAuXOpoMe
WWSDvoWk5LntswtUqLeNMGHVswg/4OIj/5Qtec/ORtmopGADwk64rXgAbXgk87uuOJXRLDu5QU13
is37Yusnx5YF/ZQpQVVRlmQUiKFxdGDTApCVakbyHIfTozJ0ps78Kk1NKbKuvkAVa3DYQfvikrwM
AJTLbFKTeJ1e8knm0eCOQonzmQV1P4a9Mln7eeilYjFAR2O1Oi3u38NZWdbEm/FcS5nOqlJIQnEB
yJ/QfmqY+9dDsb+cd/n3yFgImpnyUwaRcKb/KFbB5YyFP80W+mHvNGU86RvFKjbwf2Wqq5vPyb+N
/W5oFRQwjH0sMkUHYPRTLyRIBXbTDqx9ZT98WaxRv1Se6nEvJ9xBBIcLXORZEdZRCOKDYi1lBHbr
lt7KmzLDXdp3y67GRienPZffewBoNOAvH4kqlYe63pxo+oAjRVK9xsSrbbyT/bT0TLS7Ig8nKII5
Rgfh5M1YcIZ4hcOlKj9cegq+MlpAcLOio9aNUvg2hF1WxntIz4pSeyUuzJo3YWkn4UWRn8ava3dD
BtxPZpfmqheK7roKv1b3RnzsUozOOqwObaZn+YKNDMqK8zA200Jo0Kyc9G4ZWciq3kdAOS1k8u0v
fWsYgNda28QUbqMXaWgJBeejHqA76MC04IwWPc78Qdnmri3B6akUC6v4BhUeZeZNbXza7YS55joJ
MQVzxH+GHITiNZjykGC34lTxQT63ByRpk7Nc6JwsZqiuHK1WaN7aYL+n80YK1M/vAlgUOcDyDi21
+Lm3vt4X5tvFU+y9xuL+o7iLxhyM5gueI1zEnXrbHUrPIfkvVLWiUToI+BihkHqQZBsxwylY6e+H
p9g+fmJ0FBHFw/iB53Je7JknRvdR+yYqYWswOBsJPWlKPyFVuMNA5CzhJt1YGQcf6x0j7FdZSZSm
dc6bWgf/Vi5EJyU/ttrT8NQrHN0opwFfD+dy4oZOxHokNz3qc28SO4sncX9tn1K0+xza9ZuXzJwT
wXVF62yRsLN34weITAKqTINKaazIQY06TSXwA4n30MgDqDJxGTEzgI+q2vtTFfEa6zRPVgUrHxfA
HKxqfqOe3mc/UrQG+9MMBWEtXAEGbNlyMzFwZvfE0LrZ7f5WPGqtdkX1UgKoidtoc8KzLOF/GfYP
jgUVKto88L2aCwmRcNleyoGqv3mtGXdh78obChpJmGyZM6FNxoti+syEOSYMeGXwkRfV8ewrnHJm
xvIYrFL78/qASVJh6g0qr6czmFpdXxqmHRVZheVReH2zwUIlEwqLVsHSpATYerOviwjLUYvL+CP4
0gFvuKbuXjYRP9KCo/0xeZONypsI9A/NayxwTX6TAdAhaWxEBJXs/T3r5FbrtVkgKgaSRuFZVCoG
doQnjDKgx/kN7SVeuE1MnbsWxPr73ssPkdNeKTNLH5CiFW2MLu3KStdL9k3TyjyF3M9sJdHbD2eX
a8opEKIZL3EOoKbjTnaJVvlyICWVpFK2fYK+PhWmjJLnfZhmHbMz/UbIlUz1hlPJ8pajoI7b8j/8
mjTUtRenKMN3zEPJiSpPAW633hLJIjCPNONk0A502wjCCulJoPsW8h46LXRc8CHkpiji6A7GLkoF
DrM5+X0cP6342eL/11x4WtMJbzh9pPwS+wc6o/uRIuFNgSlvDGw5Kk0cXyJrSLH2Wi0UIRXc2nY8
GeVgiPfA/4+zrRswXDsicPEF16yaR+kipxCzrbdRAUvN48mzxPe0oWKk/0sbZ2S9XkLcVbASXqwE
V1+uBOmIru3mD/kesKfriU3ReQPmfverRbvNskpcTlcL0g+QhAPSG2793h3Gg0qJCWrLj1ytWS0I
9BQVj1AaH+6TMHO5ZJUpRwN5FBeesepLuxPIN16Wu96tVIO/RG8t6u0LzaFf2kzb2g73bM/JupB5
S5flECGJomr0qL84l9CUnBIThS+QrOHjZRTRhFIL9/hZ/G4ekVfL8CpIO9et43hIMPPxTdiCpIA8
9/gV2qu0iUQ0k6Amxb3nGqT8As/MkJ61MMRPqAnly5j9ttPN3J4CTcSiJKxIkwFxrxQ6GhcX4lST
LYEtN+AieoYq0mF8EP/wnqIVqoxL9p2vzax+bLfxx6T+ublCMiSwoeRdTQKZHqJspSioXKuRUPPI
fFw2+J48CwhhFW1EmM9ch0w4RVkn0FeVHGohZSbcUtiDKU15cGI0aD1HMM+vZgtDquw2rm3uIQSn
0mFadPj+A5ngI6x0HscE8XUthlXxSdv0bpcwI8rclN86HDRgk69IC3zFaiH06/Dw9qFD8BiMsXdz
AYp2+7vo2e2cN4tbAVGz2GUoorbaF7tMTOpt5UE8oA9qmuLu1iazjGJZQgy+i+5Rh6Dr6NH2jbMD
s8vFdI5O3QY8oaivlU8BOkiUvC5OvoCz7DkbsUIQLL6Qts3OgcZijnlGvQKW9eCAx0BblcwLm9wR
ZuvRzU9XD+y+Y0c6BWWjHdJLapCxKu0YeKB51rEGBgP96M80GpOt1AMTU11nAbT6kZAdh0kB8jSi
Gn6rVfewk2dsg63n3tG53kw/XUlTuKMBL6NEP8BsWfMefFEVEi00BgfYXeOPB5n9jcGqht7CxgcZ
sviHNyGcPcEUl9RFksQtdTKv7mlng4e0iMwQ0aZF0PqasjG7ZCEj2VGc6RrdJpVkvpyDex/ph/C+
kwk4dltk1kmQb36nlt3BcMiHSnuGPuhQbcRiwMWc1z/ZAyFyjtt80Ok3c6VUG/aILbYsK5r/UU+q
GvCqJXuBiblODXFP6azelCmJdCMj/q8k+NFDeqpYYCJIsfpPtHgwtKbYnhewSTe4P2EUBbW0iwTQ
2ZZpz/P/xdlLtW4MeqE9p1Sv85e38DD3U6XrFPZRoceQ1wT2uPVsmocsATRKflS4d/BO0kKk11lk
ohSaBguuJo/vvvg81yk6nQzXmC9kNXjRBF6dAJ7Ipzpi8JSEgXBNGofMhjXAVPSjzKMYAeMDEhu6
UKDKRZe6rCGFg5R8f0erpXrgcE62jqrC+lrgwql0ynw5CJkLI8arHcZIyjUuF55tBqckEcX8TQBr
2p4nVL/PM6vtG/M85HKaaR60+bppAfTLzFCAcWrhr9Vkbjr8H5zzxrHIS/fvjNLqdDRuZ+zf5puf
5kbKkZxGUOuVdQaeEnjv/8ELBF9UPM5FzKSiTVFvwqdfh3J5ZIrjWxOPhsNlzjGFk8H53kFU5q3c
n+NXz6ch3JuMcoaffoVEXtZ4N8t19+wIXhXejWhyuawGRcq9pcQYn5Bb+94SW4ttgfrD/F0MAYZS
vE2AiDpUm8sy93Gt1FZxroAO+fyOwegF9U6IwyuC7WdXdjWKvBcs96SdClItGs530qTSJB0FwCyV
2ilMVibYq1QFsv4rxcQsom4CpPQi4koacmyajWyHrL9pZxVALwgtoGhdGIEuRG1yTa9pfmUkS08O
U86rsVKhSjCw7W10ldTGRx80EAJ6dWBRB7nwzaDeDN7guVG8k+vIGLS2EiDFfVxbdKGE9zbEfk7l
65xYkF+Top8eo+PUtPN7GVH4lwWP4FFYDvIsP23DQ0Njg6jUQAU6pCIVCyBEHdOsTPG4xVfzuvbj
v2d/Ae+wGCRpoCd8sJJnbmBuQ9CpC15qF3wcG73CEuFcQZDtDj1eDsy4KjeqMoHxsoXfmKzCuzG+
W6CFkOcW7iX8Vr3X6en1ZhsEHi1nkljn/cqAjmwcvo2+I4uRRE9v9Q9QOiFlK59J3OWYNRO1PFua
GlCCd+LA297ID7QNB2tlPFREpTEzArGJy1cDzzHiBbAtTdd3/FlTDLLp39Ik8YniaVZgUr/YGFcA
GjPVfelvTO6ZetWhwDJXfDwC22prqLLnrkuj7Rk8LpEc/2BrZHy2ka6kkyC2KzVpJIgS5NxvV1KM
PhB5P9j33CSyxDIO+6RVHNr9StCPmFLnwdQ5fMTo2/Xr0gg9B21HNMmCfSYKBkOftfY4qPXU8isD
u6OWir5fKSQmKc5RNbhVTe2K1i/25ltb0n830rBffCkmjFfzPcjQJppdTUv2DRGbxfSMJjeWUzz1
27Jvwf/Q/tsUDA9PdJTeRNUEJyNTenPQ5t9LX7FPVehNz8ZJQSyWxzbUtKg9yfNdu6KmSLDgLxdJ
YOeayiPkfj89WCwiUct8z7AX4ZmjCXoJus3+gpC6zF1CzkNVL+4KOrN0NOkmNwCQLiZDg1W8vvfp
DbADp4R7GuutX/LEt5QcQqyNoFW0N3NZOgGYEXNBMw8AXr6+bY7YFJ1j+UqtZ3Hq/hs8KXO8ygi+
oG9TXgfe4Frsrc5UH/WLv/IoFOJbPgJPO9idnTEPtoouHRMMpyDPQLWwOiSd26nLns3PbWs0kSDX
46LwC254ImmUCtlebS64xSbcgLzbt86qEW+ARi4gL8VdzHc08RiJgNPaCRaUf3+I9C0J++T3maLg
6eCFEuq+RqaWksxJNWuVNyCEFY673ns1EAtRg/XySEQq4Y8L7I2OyjWVFo/S1wDu7klT79Wy36gW
zWtqOJM9SLRdamylpRSb+9ck/ZMsqJIjR37oBcb7+sdbCqn45RSJYghQYzUBvLN53zWQe1SwzAUD
VZN/H7RxrbzmKlodtzUev7xCCmlnmlhiduAaOBYO40lUllgl6umcu7/UZu7vC86Wsvt9QHMYBVZm
/q666Khxt6qbXbL8RRsXsg6c9XMYmRJCCzGFxnrdw7TBtPqJCs0fTbxj8nJrlhUj5y89exejbjQs
nuif56a7tIjw6xS5N7lpAhEOK8iv+j3Lf0R8KwGtlWloPiopYzVJfjtA64WuDz48B/s8/x1kWh2R
o6x8kf7nPL78ocE9BosSrJ5V6DNaxoGhpG2ag8IyX/iw1G6NaqkNYOW8v9N8PiWrIrESHu1I3UmX
Nh+eX8DZb1sRSluOP1qmcLIL15LFTsSBaB3dIxTlJBH/nG+eBgipfyCVbaYyLz8vr+92Ku/j1uGr
yXh/TMPBeW+CLB5qoZBawi9hjzuMLFyBHO9ZPjIqy90rakhJ+EE0TVwCl1/JJ4Zt7z6q/qSdWhMy
0Wex8N7zRo5ykjBYKcWssPO2WNv+m7QtLHuCBb7ocQSmnOB0r4DEbw2e51+ClRyGWZTAB91NOhv4
hOIa9TNGUmS9H16uRLOlBqg0O9GyvL4ITOZXp/HwR+/6dsHZY2kVFZJAQJ0ZMm1myQwX1wF9x9CT
dJljH0Z1Nv4zieRHADb937hz+Qpw1aYHIOeN/f3FRVDBL2FmSqB8TG/T25+VRa5Et+ru9vSFJbaS
jcgP2fSRu5FiIJJQhfHzxEf8+VnUk7FhE3XAdUoKxxTrDOnPi2wyfTh7DFhrbY8GTKubKuxVe1CL
7Y18/kMc47u7oW//bkW2TnMeEvaG5/Wc44AzY7r0Nmeqbtjkk5pRvRbtvu02QA2yq2HR+O7QcPzy
10z2LzPZU6s8D9jnK0Q0i9OXSfQPxqX/LcmVMkyLRfPLcoaO2tsVZVALZFtaD4yVSxq8q/3qlHfc
I68FRlIsFI6sOrjN4X13lrhR29tmQqj0xHoyA6R5lkXFZ9UF3wo4bnTSz6YxKVahNcwbDZFK0nwi
pb+v1Hjs2U2IQGUjlQ1nNuxyH0wBx9wZRf82Nxf25ApfCIJ5cQsUf+gpn8JcRKVgMVTYg1j6SSZL
21+WIj7tSp5tBb5HLKohjI6/m1u2AOOz3diuVPEJ6f3LhjKVa+6Qmyglfedwnzp/gvI51JKrEH0i
WlkOMWnmj6hZ9apnWdqEhkFkSau7vc18vtoXNcFKmUIcFxKY05mqpXfB2SB2eNrc3rUUn6YaYXii
PCjxY7OWPku+K/BcTT96uMyPE9Sz5paE8t53S67BpXtD/3IMnmYSjGmCodAnskaXfvAUdoY9xXfN
qqSRq6Aur1htweMqz3GUQD4alga8kggQUA4pW6cvBsAtThpDATi+d/81B0AhIRWqJeF4Jfbb2qJK
UhshbRW5ykJkpzaV3ilS2WDSh+ARU8SSzQ4nIY8K+3o40bLV9iVgnFYBYAT59MTi/LMql0+uiZd4
SpaRK/DKr1DNKDiVAnEJ0P6RZlvp5bSdpK+U7T5MBxYg+I+mlYRLQqet2VQYnrjUQtMp3m6MD7ft
AsAiGFs/IWyOSz9SIRr6w5tvh7GnGMZXGGrIkfvf2XZCPHroXOAe+SqyvithdPtse8iXLghqpyxS
ZCS5NmYN7o2yupldj258wKgsks4LbMJymW+bKXm7yzl0i68Xn4S9dxQa7Il+DqsFtbJa+xOFmQXQ
T2fDCJLkPg6vRlg2wjx65ILD5Z8OXaplUBsjvsIH3M1bueHVfiKiCgEHq357jGAA+TBVheJel/U4
NmXCg7g8eKr0AFGmOzgayRt4798q6IJxVB13zS2afxBzhTfNCF3dTl9t9rZ/CZLxPwtCGmb7Tbll
q/6FEIlGpKT/Kckn8uaUcmgL3qqCcAf+duzX0icoyN+YzDcAB8cNtglfpP8TB5KvmkcbFx0PmJvi
N+/QaMRyo807aJxrXgbXIyeaqarIEF5UkKd/WVhsVWuSWMFQLheJaK/Gj4VE1EmkwhU4geqF+sTC
qBk+11L37Tr6O2nyLRj40noPatBcRgslxPlPlppyee+/iyOyoLhzLMwchNrqL4e5W689Wo4/ctBG
rbLqJWhIQxPspBgbp9t4wEo02vRyTtKdsZus3ryKjtdUjcrrJmtOoXHVmFTGphlfwpNofLdi7WrE
LbAPakgwKIBZA1foCi6HerVeqXvrw4Un2uM243mZcfhReP0JxhqWMtl+pOdSun70PcL8AlsR8FIQ
j9q2uwW/L3RfGBw6YZsT9kBJeQKOfpN2hEIn/60r2xG7JmTwTiHDh/ZWU87pBdnW3u1awWyZcvRU
0hsES7q7RPkdOnOOqmPYych/AdJSTj99HDtMwOAZPUhbdVLiZajSZCqoDf04tQIyrMetXPAwf3p1
kWW11n9sYOK4UrCqXfvbUnNSg3n6dAvXaTLrTOKs7k1smhqZwa34qhAZiW/o2FmatYIPXlV2Ocul
ikEYsEFx0Dlhy9XVsy+zADz4rYwr8aEqsmbfrJvzffRYjb3LavcU+8M2GOfqfj2iZLN0kyKPd/TL
1G6NW7ZuqeCPTTlUCOu+vqj6Z6MuR/9QaCjXuRFSzKx7/6wBPAZU6eFIjoXsDGDtBRftYEYhjiha
dMgjeVeaGnY0idb5Ie+kXp2IhJx4cpYYQ1OBq0RS/8cQMmbVLEAE7YoTCyzYKIKXVSksZqirqRjn
UiGq54CcTD3j44EdW0rsaTmuPQOOo58oCpr2Ks81mgoaz/kkrAyR8zddVOw6jUjwY3pkKMOXB0YY
iQ+4KHfl6qqERTdxvg4uizmstnaYi6pmFrlbap8JfBMQ35eHqat5B+SYFIMDp9ExuaP9em/x/+vQ
6HPvWNb6ioTJZg0CHNC2BrCbIXWepQNSUpEAM2lpEhWNNTJnsU3wMKxf7G1GwaVA7oQ1gzcc3h+z
V7YX1/wlc5QEKIDEAxXSJCNZLX7ldoIWoujPS6RQNQOOGZrzsyQYPQAtYgMP6K3f54lRg6k6m2EN
Ku9YKmXz0jNq584/QtH2fXBNtPBRZfvyL75YvNJsYglum89EVaJ1BnyxNgsh4K925adWsjpi2HVT
1TBreXJSFjqT1YzgNc+2DycWj1+odbXYmsavsm59ELeQvfYEd/rj39uXe7OoH5knfklcTlFyK2Ri
+COYs+beGucU3cirNyVHhUppmVVyj9LDwab0g+UVdVexerBLF/q1nxa1JdAfPJFvOZmyows0UlTJ
uVBLUTrzj889erCI358/65H3pWUptxrm4iS498DN/x1/uGejtnrkLmyPif6p72ZVJBWaijKDUEnb
HPbdj15uIs6eIWkEUuflCt8msvuRBacrg0QAEQ8MMxIJy5plm62gIp/KfutZnHKPdvEW8sFqmemF
yG3lMglRd7OBZAZi/EyBeM2un+myr5PL9yodhZVWsJIEqtrszcmMb+TM0IJRBtTxgV+caDPA3LwY
wM21rQ7lFa1fvw14pn+FIlwWMfrLg0rrOs01Zz5OMoYoWvXcmHHdmdZVxvPmuVyxCUct+wNertoQ
Gabk2dakkZdzYmXQOlIHlrvuItQHumZ3DH5fkaw/njcq2osm5fHWdoC9PeS9nEeS8veqyeoE4NN/
NeAnSUkeeZIx4SWYTH5qeK8FWliVVMOhX5eyHhnX7ontn5SFbglGizniEHxqSiIZM7eQKtancUgR
HLN61wlEasmEUY6M0FFN2WKGpdhV4d2kr5X/Guys7YqRJyYgUbyMiLTMquA2QqNFxCzKTuaAIcEn
hf/I62gOKOrKhNH7aSIFKjpEwTIVpFG7Gn1v3PZ6wm9hnAP4IIHZbyks/WOexDF7XRTtLb1i8SvK
dZgym/HBdzB9XF6HBwyJBW5J3Qnn/+CjQaL4ZbBj+bJh5xDs2f2vb4PiwNrSHwef3TOTYqaxJgXt
mrA4Pzo5M2s5HhZ+hZGA64TTsTUXTXdIGB780FPZJ3YPBTOy83cg6JmBFKQccsx3PSsTHX2ky8Ic
Ewe8+KrcsxGyH7EvJ0CM0RA/pZ864KgrGTVnSGmPjZdFyd+8FV1/BOLGqvYK3wCIUzn07tZo14k6
jILo+LeFwkIgP9giBZtmgKqlG0hXeprn7tV5USgIvnVcY4ZuYSp5fYObP9mmk01Ier0jyikEEf1N
okPfAV4gcoRIKd6vVcnEcE4CWFkhf3XgD5Zle8TVre4OM4ie1wo7yTmNwLFDaUZb7Xi54hMCjI7p
meHzYWmerfkEwfOmM8bWxS+K2plxt+dP4R0bGWo1SMicDlqdr9/2QtrNgEMmd9HOHJNLDsHOOVWv
AaEXhYtf46zu/40fVNHbkL7fp567bpVaSRx5CG7R6JeI7D1GiWjd/k93BoNLRoVmvElBfdvRq9uG
t0mR7sN3J5D/8vwp1Ca8oX8pzzXuyo2J4Zyvv+WLAchCG8/PZFRrOvezLt/t25cpTm2m6nH5Iksd
T4Hx5DHULpkLul5qLfLOYSS3LfawUzLqrj5Zrk6euEVDniL6YPqwMDISQLxSXIMMXtgGcwnMtfpJ
DW+RhN5plLtyKzaOxeGSS542Sf6+U/I0Nn8him7cfZrnbmEnOgHQRejekVlqxfHQXaMWjnhZ/D99
7bSMaba1pD0FTSmnsoOb66Zc2XiSsVsF02VPV6ZZbSRWxkUjL7hGGFR0r+0DTS8klOuga2SLETja
MNzEbZjg0evw8PZCCdigQqUPmkrqWY1odvbfuGWDBoe+TGlGSoqY+YUIkfZZf/OIJgmmrzyjKkJc
r1wQAJ3FZOpxv7LUA/YCYbhGeo8cn0IQYK3LfLPCXnkmBL2ZS8tLix/uHcHyxFmdPn+HJgMIDlRo
v+L+XJUYM85+1pDK+n8IdwBOnA6MSvkDxly3cqqjWgmOh289pjzWNIk4aaNiZCnN8508Shiw2NIc
yzlClAX6sfHkqcKnYSyW2fWJIkLS3HO5XJyWhod8e54SK6UG4j54cRefb5T18YdFvUw++Y6/PM1M
2Qx91Y6UMw6ZI0WpffEWQV8TnNoQhgM53WATc4JHQvMxVc1PCGWD217v6X4Y+b9B6Z38uZIY+XTW
TOPgTAFAmgVUmNfaS2xOaBkd0WDuOrB7MnLcNIeXrEv3DpSZFjXNNhntNCtYKKQ/8gDSe8vS8w0E
pUf4ji5lo3R3ynKVBpIk+cwf+4AvggO5lDZu27UC+SgjIJ+sO0LKjv8+IAki5CQkLcH6GLFNILUt
1UvVX4CDbhRS3Xvlr5Qc7uK5q8XcPZUUZ2Qa6v5cWDmuSFqgcQOoPnaOpfGwGHXV2sBqxfWyKeaX
uMtUL6/1boYtRdW4K7PpIaAd5ZQcnjnVBXQDB/8Qf8ZLODN3bFKkI/nZMn3rEb8F6OcznQAYs5O8
Uf/9QVy7hFispctcVO3C/PvGKwhNWKoJfzLASY3NRimVUqPdPNbwBuzVrd6qDZVo//nvYY15Qr0Q
7UwkQYxi/idSUftmgxYu7LmKULw0Fh9MupwCiZcG8UIuFa/WdQiiDSd6af4r8viP2xd2D0wVYxX8
+5H6+4TE8qhZTEYt/m/SJrue7JvJdPLUKHtK86AXzUrLqHGGN5znoJEmsCdNdcevHoVH/5Kca72n
531pPXgw7bG9gYzmlsEfaDlv9x0+dqgtcE8A1uDXhNNq1sr7QLW1IHvHm96KhUEWOKuGW3G7A0LD
O3NwRZdbO4WvxIAUHmqfLQ2OUs0IXHcbdVJCam4WKB1y8Tvn3XH0+noDn7mI79U2T5dhOWgiqIVl
ko8VLD6pwnNHL7pH3698b7tf2LjS4hCIsWZExSSsdf8W2RINYnp0rCmf4zevU5jGYCiRRjBZ4ASO
4JKvz0iduQIm9N+bR8/zstkw8hRu7Lw554Pmfjj+d/EYbz9r4QiihoEn3/d6GDfpGghZxk53iipD
6CnLabw7td6P8pqv5QXSfv0E9xhZHuG6hxdeteE4Jr+FDPCsiERFQQmRmR+cMILMKiRAmdpsXkxU
Ad6OQnmSjHO+W/urMRbq1oqBpuAqRPB8gOIU01VUmQtj2Wy2fWTIWSINSNZHyMXt8ktOilTkNUMg
zRf+qdZxuQBdDb7VbQ0Hz4DJr20O1J7nC6eOpEOMKRG0yc0T/c9z/quJYPQKhb9r/TB9D5o/UBjQ
Y69LkNbCRndT+YQ674NFBO9yV9SOFtlEiMkrXKWtKMrWBlC6d91fbDPjRSzLc9aynR2rXWgGkzqB
KN3sPC2oseShmHuzRxeQ6JHTU4Edp8ueAoKrMhHPD1dvXTp/2IvL2SZ9rYnd6hMUS/vhWC2tFctx
5hIRruSAMf8ilYZu7rHuPoK9bXR/DyE7SECxME2M4T9r51ko2LK39OPcI9Mx1ThBCG1byeoFQsjq
vXMk8VjFJvsz2q0JHQ7JPqLGpyj11dKmFNuxj6S8HYvbFVR8XvHHNBGTpvIAiNePSZD97CPjmoC7
wtL3H3vd7SQhcWn7txg06DYCTg9l5iCyBa2N5d6rczbWNQHnQIVmLizk1a0fTtdBTz65k+xUGdu7
bMON8eYkMn4+FwPNHn+y8yx+57hNJiYq+nbLj0kE33Go4lrZO9ZDdSCiBA7ej2o8hV/jri+tWvgh
PRmII5AZI/L8MTuj+1FZSte/l3jQQc79Ehl33gy8gW8zQS83P1m37xJVaDXCJB5O4RuI5thlaLNJ
N3jR/PomamCrs/ue7NJUhO9moaooVPpqzj/6BTo9Nnn3ONy+CDO9fK/RUiOAGPe55V7Ig7SquBCm
jNh1FTbkDQN35rabAZRqvR1U9M8kAmUbA7kpszxtLb9q7CsLoiyzZx16naoZqHrsLoBHOy0Lmk+G
cRU4mdqdgtCGnOFpibVtcr+BB/3hDNatBMB5hLLGITdOxqNwevIhXYHiz/lfBRe6D4w64MbJAI0N
qolLlH9ntUtQKcMpxv0VE8sUXkWn99BpOlowA0T05H+Z9xEyf4MFZW5FdW2dGIgjVwuoCe1xtUNU
8IJ/SHG9imeAJQ6QUwONA2ny3el3M8y2OcbZA5kPXWHse4O4ee8Bv1Lf0odqHnyJ/d9dbXctgFzm
z/8pMJBLjyiuiibz8bvb4yg18ZaRO0+aMOp12A7uN+PpPU8x0rhZ/FBNu7c03VV8nJ63oFqxJbbS
HAv9Fvz7NpJwBpzlqikesZke4GS8QIkR03rlUfaHXF+tbElGN2xM2M2RA2waXmu3ZtkAmDeU86RJ
3G8g/AAcnZGbpmIWsS04KKtA9owcHCirV3d2Hx9jgpr1T9q8mD69Jdg5KGszVDS6zRGX1zYTzHUD
rj0qfUO3kUkOnijzwgT75Kru4yjiyt97mMA4n+aCrK2iDSpGzt6vx+Bg7Pkvf3rEL2fvga1pC2Cr
GLLbKPyYOim46tmGeirD4/9p+enQLpbSpTVVOcwnnfICqaNlJ3+0kNpfRaq+JtIcrEQ2N3mjj5Lx
YdwdELPDghGFkcM+Ni/8bPMYObrYee5nmIlrWGAXIVgURUu+K5I4ARovt0tUh7QpH7MlmiZC7rAT
6w7eqSdJtZop9xQu+nTUFlKurHig/1Sq0aUxn6yMYJvBV4w9w0tGMal+6ScyZa/e4LKo31kASuiZ
/XuNH9f7hFruSCo4L4sO3eMdNPGAMcCnPieaYZ+F/yZOqWqlBl3Xh151dp7PzozuOofHaO3YRp5A
90YWzDR9ceI+XZpC0DuFtmf+wzEVKtvRRWrbXLJhCtxCCsuNjzDnHi77RhihyZpkUtF5CMhXx5vZ
jDWl65LCjwmEWlDOQgTFJi+0ydmK0IAiWaXtDbcABBfdIpjp9yLLNnCjKXCzx3yzyTAmhoWk9eXF
TRlAYqqQRNGrSZ/PeKro7ffSdYNvprqB8Se3BKazNuTrcYh1BZZCTKEqK0VImsbDEjnjOha5HF9S
nBhTLSegrYQykJJbsTGM/7fsUk4Atimj/+TSiJBBJ7lrX4FnNATfmAjHwaLoRDiXPbecHZCf1qvl
UuBAaVvKBfWEBt6BkOupooMFU+YCrlTKWoKJkJ2gR3Dqaq/JeCVFMLzDAWsJIGMt+P1T+2H7elEF
Ib2/eucw4euM3fZVpm+XaurbJ0y4zRXypZlVpKOdI0+lbzem2EXC2MPoWfDsr57I2QCe2zgOfgHO
grfQTY4iX4DPRaAPbScRHCDqd+syBr+OYtSNcQqZ8fYzkPUgUy5zwQZdaLuhzLshNuQWQxkNZXC2
XS8MyBKDIbta/QiRqfGVMLbB3J++ZK+aNbiQFiQ4iBw8ah/EjFypEehGgjFWrZrK3kKOniwpQE9V
q+NwK26y2EdpqfhaHSyzntL0D+UkV1bU8MMd1AHh7pmKc++/r21TrJkhnOn8Fv/jhgxinu2RREP3
X8CCrKdnNiEXqqgzo0t4s77BkjW2bfoahHZLCvrTu3KnLVQq9v7wCG7CsswmYLTJNjuSQ7yw+R9Q
lgrVEZrsfSlZRosr9NGY1DvWxGOS+ShL2tLskGi4CVva2ajuII91aeYqDiMxcOAf4ni6JmY0IlXg
CDr2lSr3G6aTWp38c+79yavC/azz4EAJLHp/PUMT3mYFgvzsHNOkMig3cre72NIWK0W/4PIDBLXI
BNzhSy4V25sLpHFD3IH0BSj7tIls8P6CmW1vhGIBAR+fQ8ANmQzLfoL8fhOS7DcLEQ9hpO7HoGPi
VGZeko7KuU0WotsiCleWrIveZNXzjMxo7btVnV/naMvUYA+dPYauSQRsb4ecjyKFOaNthOzv6ARW
IN+6S0lESPVYgoY43FRgRNq6t1A0tM+WcJu72mpz4aR0JMJIG100ZxFXpD9x/EDn5gQXROOLJ2CK
cU96R9sTGLKZrJmu+jrOyFOfrloDq3+7vIWxG1vHbfkulHzFGpI53IVD6TqbzCx2+k9KcxnP+nMn
tOMTb6emKHv8uXGyzEsUK/cvuO2ht5kqkIM2alfPusW+lCgMw1epkCfcn2StOcFk6jV7/BnegPpi
bwYvn6f7bnbkIhfEXfzHlhcfbqEJ4f7852Hil2PYbbc3xgp25jz2/R7yVVOl97eFYm/kZBQAztR+
hZg/QB6TmOLy4gqHZbQQnlPkPh1N5OEXWtWfuWnyCDUNl8iYBtKlDMNZGycmhWPK3RY6EU46OAD0
l24T0csjWoy6soWnIvbdj5j7SKSOoTvtybOFM4umUY3bmJGGuuVZivIDSEbAgCrwzBfm6Nzmg/cT
6ODUknsR0Kw9S3DaFOdUP2IfDwCvrrc+5GzSqodikR9SeTchz+4Pr5dB3MTfpum96zuQTow2BBh3
In066BT0ncKaltcVCARl1RLKW6qpMPD+B463Y9NEmA1XwVhhu8teWIUUd+9LVFNPG3IwJcM/G0Xw
4XRi9gQNFxgMBpXn7rnmOl5aDOt8V1BnsSEOIHRdJ/ET+A14M3bs39u5tnrfUZdzO7u+dbdyN5EC
a9WyUpgTlg72MHNequwGUShhjAnsYEK5BIkhF+8LOsj3iZjh7e8+Q4Ux6ZWCzNcDp0M2zSafXNtC
ESTKDItk8Fw0GoRkguX70lGyszV0txvT3U56kUtBwG4Lkpxp5g+3UQ4EvT7TcWDEjvqAwPAOqjQt
fMPHjO+xri+3MAiFHcxz2Js2eHklUegzvTD9IIv1b8oyd8PkYUUDHPchNZtnOiiTYouVgtJcxV+A
9OIn3onKHnIa5m1RWZLAyxiCq2P7DWnGLkPYJKA5hjdNdhBmp4q/NkdRijAwhKT7wLO8wlIBvY9Y
ZoHUaGWRgo5ChmrdyWO1CMKDb0mHSjgOZlDVkJrGmAG0Lx+vm6BbfY0GN1i3aoKX3AKeZ5bd+ccn
VON01+Nak/gNjQhQqX3/FxBxN4FXmKp2Z8VPZEzKb40/v0U2jKjiF9mpzLd10/rFkr6XbuP8pgRx
3t08tl9fW7SdLkusxBrrS28ZjL55qh0Kk9FOtZnUSylx1QrE/QjDHcOsrYtTG50jKFsnsUGDUgqr
sypo5idjsHA1UT35gUvkA6wBe8k0bAm9FcUNC5Qrk/5w/SxS94ELM01KH17jkDmFjPEuaJGF47EI
Bk8m+5ISRySQqBGF1jnW5leiLZvskneGvLIOEvikIe8YQtkr+Pz026a52a6pJDNX/WVlomRcCMpg
voGGEPz/bbZ5leKMSxD2WDdWdFZJO7+jhciSQm6Uwh7I0Pg78Kfsqv5mIM5Zm0NdCcSqX6KAwzsm
50A5aSWVzS8y+4/lcN5e75RX4SU5sluS0M384SunZ+ZvF5qS4jTpwvEyFwkrg9sevXCL/lzx2V2M
f0W1T4CCvrQh2iReji6gH9qkoJrxR2SUwdlUhKpfW8uSRGjmPQopT7JoTM/J3o0KCm80fT0L0WKX
TxqAC9tJjbaTQdvwxGt0Pa0JDPgSRNkyCK85iY+74gfhhU8pP7uR6g78TClVoC47bFJK04MSA7Lr
aDvTLROjJNs84DeoAn8V9uykCy4ULWCzFUNEaly+13cdMHbWIO8EnR64CfXXku6WngLMqYQvgA9T
FlxhAAOuEDj3PiEL3xaLoALncCQOIyqYKGxvj3nYbTJAXJLph5pRnDgaWG1VIEcdag2cE+fqr18o
tL0hbrlZbOv3e2EEfa3yypd2JsrKZHcLvK0FUQNQph3zCiXyV2/zd74G16W5lnPNSCPu4OWU+BAy
FpnaghuccQumc+SzWWZfDaTb0kzyftXwEVvMks3tfJ6kuUQxQlqGsuRiviGO6f2QsyjhDlzOQO1N
BDxLEog1atArYFWu7IFseqDEZnYNHtR7M8h52BP021MkqeVoQwq3BtbyKJXwp31BCgNQZqWP7rFG
rFWBeiXsqllpcyiTzWr6tKxk6zttrKLmJRqzavK2QfJBoqbDyKjaT9VDY7tyV3DVoka5/zf3S+UK
DIusBGGkDcUmRfwkucoTESzN/ydlvP4hULceyngCpRxSvduTuF20ZFgqxSgtkX0Vdsmy6fiy+dac
HPMNIfrEF81o4/G/fTw+MhG4esHNE8kE8zzM6Vb47fIiXjINA0tSlBEJbOsy1HYOgxSdpeVQ9eQt
HPgA1PoukiRqu6r+gQXNT7QCS5wCCLWp64FY1kmSZxYsJ8m5y5HmdvzjnE5xyVf/UbTWfnAzbJY6
LJ3txL9ypenCwXzvEryMX/9X4zEPj9sGOiuSOjLD5iHDShlBoHEdZBvnsgibGSH+nv8kLYVAdUad
ERyDMIA3apZaLV2s6ftNREHrazWzY4ltYIOMxytXH8vmSd1pF+hP3FlijON3UfXfdtgMEkwk25G0
AWkIzfT9YH16sOBU8m9WP81whffLqm6U7+xkntvR/2Eijf5fT04mHTvSJKAHn/qIQH0zC+DfIRrm
M8x7dD2NZo9c9hVEurEaKETtvXrDwtyfkrt1nDzyzn98Bqwhpuc1Ge7r4M5IIe9JE0RhYyiy+WOU
7A0ErvpdQpOfObG8B1ROlS4A6SvORqH4lxSMDolWwCoMiWgkCSs06NyZLbT8Mghrr2xys5C74lX5
N7XDLTZpX0CrnzhW79uyCiLHYD3dRfZ3fig5N8EdIayBF/iZVjhmcuy3ncDdtP6jJIo/gilOBnBL
4FpgCV24fIM/u0vcmLMuBi5DI1nrs62V+6oiu2YwpocTTpnC9tmnthOul7/39VzBBs+jfoSZqYBp
aLB+sUGNZEG9JYSLR10wV9mQGCyrJEFCQT3m4RB/k5UUZV7HoDyoKtIyFe5En/mmUrE+Uz3NLn9J
MZDl/pVQKK6AnFYyZb9HcPLESDQZKD1N7euO8E4ali/+wDMVkNT9vKj++ZRARzdG4TCZQivWrDpM
n3mF+nmELttjlM0OnakY/VRXjUk6vaLEEk7Hcxs7c8E+H8582Ri+BoIHmbwfHdIHYHjjWPs5MJnE
pLdvFouRJETODk26ftc26gwM7g+d+YL6YactkkyNWLH6D8Ku/QN4OOLtgJsJ9qnHzRs4bCxvH1xH
0jB/CIwCBne42cTOEdC3gOLchJA4Idd/bsVLjABeyTJr5h4kfzTF7IV/MquBUWCoIFWpYv1+IYe1
Vwk6n1y4vmlqK10f+1kKy2N69fE+XtLfROTxgRLElIsCiuRsn5T4W8n0zjS8Gbi+NjNOp2gleplv
O5rFOlqMJnD7YNxhxlzghgDHUFkTcaoLPbsFbAh8xcnj3QEyUJoPWL3aD1A0EgvTLNwp4oX2eJEM
BU7DXf3qZrlczlEIqu4ZINASrnA08E28NvaWASzZVYriE/0wjuFlxTvZrU9oGyTg0r9Zq/q8IwHi
jTxd2u78fzoonAUVIszotu39o9zmn34pqhY1sBcZfc8hTLks1cm7EW3P5gzMbA5xIKarAJCJVxmj
jctuUE/2KjsrFTIs2WOrr5SvMmAw6GCk0IAqWcXwjBxzWDIWLpbgRVEAOuIeMEYoQyQmraJuG1tM
afDPxG1Evwh0H5vsOGmtwFol3D+z8F9CZ5/o8Yna15zdTvJs/ZwEuZuqzkh7Zfl/2ZzYlDKXkBup
5pEa5gMUAaBcQfUPK1GyuwiqWJrqgT4rQE2P8ghDz60uEHF+zZ+uRl0qxBKjVR4ksIO0oF9cK9JN
73DxncZBwY1W0qlLm/yFlkRanCqaLFJrBJL/CYRazLoE4sg8l7G3z2W1CIx1QrQA95zHOf/pYpJv
DKfDjB24gYQ7RsdWQBXncOXghRYW1NbkCOybri0aSnh2pKWYNYzOyLzl0rL2FnftrWE/R/3PLklQ
JTA8Y9HIa1wCYocPnnLPs9wre3+W9MWBRibTjIAllUB/CjkX9ly6lXU281GyOO1VvAJRAssR50jw
gbXSgtuHUuR85nvl3Dl0CSzt7aL3uTfo5yM56Zv3fglm/FqtGmpsvFBrg0+Ono2gbwknzni5m0dh
0inQdAnLQtSRj1bOXBmd4GAQN3RNG4HoxUqjN2YTL2UTowyiD5nWSLU3jPkEk4j2RYbLeCZmY4Yz
UFuNRQZ5w1j/axxc+svLFXq1XfcJ1m9dT1HrIC4mB0RzJBfCoshIGx0mUK+pw38uvpxY4jQWv3QX
07q2sa6XyfH4UdmbhwSIfPuxwcxrhtVUWMyr6ClWUy4P3YT5eqUmztb9n/ajqXjCKCXY1pb8TfPC
lS8RoJDyTQW2qREPGEZW2OQ74CObQILMgavJtEwsTEJxZACz4UXkBAz0RyN0BxViHE8AWylOMPJQ
4fJeuXuPZtMd0tfAdaDrlbD/BtloA48vMqIhL8fyPAVRDPK+VFaSLej/F/7eQ+4YHRG3bWayYZgG
VSB82ju47Jmpf6URn0UcaRc08f0dtT5tozlfP3z13GMzZYhbp65jvQJ834fCFWsI3EXUVfpX/qwc
jS5x3kGHHZGkGrZ9lf6bXty4qdfc0oGV4AYdSUKmgBtdtcuFdApcES0PGcX6+H66viSM+6I699HP
NhAAVfhBK9HRuuakssSVhpvuCgXjDsFgrXqBiOd6BJttsb812ygmitrj97BO8S4qfeWUs26rAIAE
Q2F+FazkcDDIE+u8lQLsW6zCD2LHC0ELjjhIjp7oo2EFXQRSKIPi8c3UmkaNkMOfyxsA2Akwzn5C
VbMObouwMyhpuPpHOqTKGMZElbj3KBVwSvaO5kVDpFC3DUlwlKRt2xw2NUk3FVGwybuJIf+QPYIE
dAXZs2Nf6YziqKzS3cJCG8yfZr2QB8Ytr8wj4v3gqd99lR6JWL2cuoKBseXPkEIltD3CjXJ0q0/P
iq/MN0WlsMFQaCbZ8JGb0BsDUaIezfbt3Ktyk48Dx/6XIr6BU1EpRc+y4n5xy10KCJSux4GlkZ6H
uOkLYqrIyfeToiaEImZdMyMblB0KGhywByMVkowZ/D7OuAIwUXF6fT+ST4hJUAiaRS+jdq1nX8b2
BH843q8E+zulNGQ46GHfM3S18D0L94PUKlnO+F3q8avW+6JV3WWQXQv7S/JmsY1bs0sLWnE2xR6f
3QyoJ8hqxhPCqTD+Ni4gRvRSBnCZd6MhScoZqs8f5MUzeFttGXcz4XCwupRhdQd2CgxTXx+aqDdl
2vF6kQ1iZ1qGXuzJZlZpzlRhd7iCNJMdt+mV8V2gCwcXQmmDDXGvFpsz5Hu7oOFObFae4HQY9QAL
pfvFOeqzTUu/zEna1+lJWtFdTghAkaSee3zguDFUIgBNpCAtgDjQioL7+6bTs+/ntq6/uX0AyqIE
wlaOALzcOiAHtzQvGWfS/nwMkjvd+d1izEfi0Pry0Kg25m3RG3cTM1KkVOpmvlQgnRUYD4dpZYLc
EbG0yxEIvtZgIMqMNw8cNBmLSEp8hdkI3AyHfZWiGPNmQqAYeRD3y1S5+D4kxtbfKNMFFY2XOj6l
5bnJPDXsAlELCq2mFX//7uRJGsMdA+/Trzi+OFYlZfVDJAJmXG60ntJq430Pm6Ui23wIojkeURJ1
192E/YKWU72H3q1MKRcUVDpMS/W1E7mMaA8L5IuZ6bUJs9bl7sDo6nZ93v/CxCi3CBZSp9MjG+Nw
QgGDMrtvnjKTDFTrP1t6wxjnHkxYgIr33djL7RyvGUAsQYhu2TCF4Wj0I8fcPkNIIdbvOI86TaY8
3PGuPRCRbsfWr2bufKxYSBLDOmJJCPVxViQQVC81+alN82Qtx7zwPNf/exEXyU15LvNm+LXsqHmW
qPvwLnolkLcOdaX8mPnBONI9RGZZQRnIRRMdLUB46X5cIVVTkcaIRwOmx4YdieULF/hDb0FlpGB6
kyIhd5x7fgIlRV5R8bVzEhl7QyiWGJUJXgeqdAW5ezmIoeXKgaa41gkLCTRy4XJxdZyhdd/Ta7jJ
c431avuQYZz7m3NLO4bDK52FkjNhQ7PM9cMbjz+R9E39ChEuIK0OUBfXdlIyjNeSD8xBQIxgUn5f
Gykw04SU4CRY9pI9KDdDp3cpQgmHOHUjmV5mTpmVN1npq11r0Hp0lELIksL6cxmaCbvz62Grir+G
kj3KSYARC0uh9bb9it3ksHljSMRzCn+INcY5qha3zKbF7aGMFinxjoqOCeEoWC5gN3k8RTzPJNZw
9q+swsSrPCyGFbndpUtXGJfmT+TBAT7U405AM9JpuvhWhatfyKgyEHL3mtFbPOnrsrm/fRnqgrl/
Btl9qaXjwP95z/6Tp77enQh6Btz+kyEvS0zFFNIClHYvUWuG6N0S+VwPQthD9Ne+R4FVg8k5TFHA
bHlxbA10IZp+6Cu6/IlLsJUyVz/KeUEMcOZLpHQWv0BmMG28WUUrxcWNBx4Dl72MIcTdfHjse+0p
LIGGREuTX71llwXF3oW82SZ+aL0nHV8TcQHFP5ihWYeGDjJFDPK+G0DB9TUSTLBFxDHKrBu1+4y3
OnsG+SEz/7LRxnN0QHeoRNoEbfrUp3PQleXHZgdIKg3qE2U3v/RNLhyfdVGujBiIR0XKRDIJ2Z8o
z/I6bx1cLXH4N3258+OYbCPIdwwKn6IPxuE5KoK+t092Ml8vEt6Bso7dw0/h0eZwCuV+yTMXHmRH
9dQXos15JWsuzTMTk6T0LZ/HnCTuOT7Ca+OR49EHM224jKHqpnjZxnq9bhWyJcnGL5eVEkrdGMV5
deg4st4TAjDNjZh9PD681g28TayY66cgwJ/txdfi336cDH2S2wVsPuBdBMOP/r1iVHonT9fOZDVG
Z8cfOy/9rm50qpsJ3+nEcTP+OTeTYWcMEpc/5ARTjQO2GIHtRKi57PWmk4sZFMOpeHRjHe9giB+3
KG3cLFLsRI1bAef8X0nhOA+VsRtC2i9Q7j8YWFEOq29UZgDoSWcanm9gPR5NNPLYnrjyVWavqfhN
TKW1CED/1HZiFGdFT2RHoBnO9WsjDuvJReitnNzZhjmpbpp0WMc+QAWaZCxjTdhYPmHNvfwpAleL
jkIXTD3bJI+S2fXJDnkzc5G+TFSYMBdi5hWYdN4q5BTb1yJenUuLh5r/Q5iF/nUbnsQTrnDFhC71
Kp//eNIDSN/TtIJXoKzrDUjP2VJa6QaKVQ6J9POW8M2rYpW2PLSwCK2U4ssCu9J85gjeJFSi333Z
zbZJbyZIELzN8JbnJCkj2ZdT44MFzcu+e/QzYq+Xw0/exaflvdCJDlD1ulBPlcuEpwiE+sulK2OT
athOFp/yasCLsoOv/DHSZjVECSwiUhAob8lB1WJJoBXvaN6JH3nvwC0jhjF9Pp5Cve4F7r9Y+d0I
kqoi1OB1LOTWzz3ln2YnxQUP+/M76/DRaQBZS14odh+2a/2mJVcRzvNtHlaK/8/7sy3cffNOl/iH
SRen4NaxnqpgJVGjuciKD4Z4H+nA9y5I0fxanlyzrgkW74hCsN2P5q/lUcDkWppz6g/wKdUm/E4r
gaRTuYfFD2vtfUSxs2mzsoGDn6eFbKxXvc9sXzlUdJnHQ3BeJLdfjGB6qGITz8LZzdsvV860B5Uv
HL2njA2bQbS6AKnOBQuRVgLoMCpfC7VYS/Kq3Ltc3xLz3BvKDcgyb0vJWivagJC58pxv3r7lOArY
axTfXSjrp8ExgtK8mI7veVYnNpouOhWEkXwmTP5je9jiJ7UOYlocmNX/Qya0rkIGX45u04Xd82th
zR5aJ4FQeR0PDpiWCjtww7BzmxzqcHvnbXzpY7lruhtpQbTEY54YStobn4iuZZHP2xhSUvLU9yLl
hjpbfI1EZSM/LFJiJW+B3jRM0D1cBZ26DG+SCkj+6nYT/ql05hg+Z6rD86/L6FkwG/DQUFXUuH7k
yIYmikUQebP6Tdb7FXFkdKjybfpR6lhBK2OzYZYkDL64bf0OQr3+IMcaaAONgfeUNv6AS/AEx/ek
MuMiPysLPAoUAa33v6lacr7JrCs4KNBQVvKgC9mmgxLEOFNpL8mlZMJhDuPmv5XDsjourifASEJD
tl4oe7x6Bq6j/hkDYjT7eKvFb6dkQ3/ltK8ljK2l5dvoCwFdB9hFv9MRLTjmV56EulRA8ZBFNP1r
aV9SXptGsPqoFfAWqnN0qiT3yaI0CBfXTzPqLO4NMNqP1C44WlAZCoIiJd30/SRQqbA4fy8mxM7q
wGjujV9ttYcmrsgXCa+vRJnpRnF+YhticKF2XXD6w6EfKxbH9lsKLs780ottF6zfAMeDGOzFCQSU
s9FipPdMmedGacUU8Z06IMbq4o+I2rv3YuhadmNe8SQtrCkkJcag6MNEa4c513dh8D41nmk4J7le
AyBBh+fhbxjTlS2X2tw7k6teEij3sJ2TRpPxAq5MMFgT8lMFEktDUdRySZbV1v8lgRNOi8TsnlWA
GM31FZMUc1YJ+YILQ909tsFtdXwQDVl2RCHbUnFC6ug1j2HWXeQSyTSh2fRcxMGPpc3iMHtgGPI1
v43jmB/SCP0UcBxQQyWKHogHbmS4yUcc3uiwC7vsmakpxvrYkX7pc+BRnTF0pB39FD349HVUFvmE
wXmdS+qT243pMsFGJ86Y5VyJj+NHPVJhC+niropmnaus9WokJTPL+628JY0/9CGvSTwqKm/g8SgY
v4d6b29BjfgEMP7cM4NIYqdxoiVIvMMg0FACpt+TZntqoGa+Hyzd5BftkPvSXNM/R71QaPb/RrV9
EOvfxU7KBu1gvZvxisWWLKVvLUBNPECSez3Du91e+DkbJ+de948VKV55UGJrdKpmwflerFxlWsvU
49vDgoXgfHjNndCmUqQa2DLFqG08ea+8zxCaBQdCwcOWnk1VW2wxNz273JbcWFeGjkgTYAsDtk2R
igfunu7sZNAFZdQRlKV38df13loc2D4x2yCtKthDuk2F3TLCnOthL8J/lqoUIlB0+oodRuCG/0vF
AyTHsVWceJq8OlS4X+O4hb8coJfTX2U+lgBiMbSFhHruvwlec0sKTfOXuWXMaUDz6yt2jz1+GKFU
yezlFKDZO638J3GWfB+7jhLK0hk+u4nioezrJEdJEa10EoUESx80anflr2niXLXWc8nrzECacVoF
xrbNcDZZwz+/gI6IWkTm2190QqMfWCydVymA2lMbRlAgCD9rwSFbqJPchjcOCgoTuZfx9Wwd7rjU
bKqzF1W+NE1CMqm3P+rYB7MbmJjGIJxuDoXUvU9RXW2ipMFi6WRo6bR8qSNk8477D+Swaxe9oLRs
F/kPsq4IyRolGpZsdYvTW3S4NsVTekLarmgmiP58OjNI1MygBxxbL2cAjLdcwC8G1MmZg1VUJo3p
6sA9n+Ez4Zy1h1HVQ+z3PIxM1bZIS+DrTiYn5i68MtgZ86RvKHSp88xIsh6l5orziS+AEvksp52j
GVrfQ/NSnZmRbTCSezgYMeU3+m0F5f5jqmkquJyiN4ZbBkJ8t0KnEKoZRGJGcfsucxWy36zixEyN
pLal+NYZ4IM4UCIU2k0D87Yx909Lf25fV2vzWkjGY4/4ig1TVMVeYQVflQmaNzwfhRcRfJqdggW/
txw+M/HIDK2HrSNgJ6s0LetP16g5JQUF6mrrBetVrzjZtAxk238MkwhbMGbsgC28gE+Wv59Pih+B
BF8y60zWANtOwtzI7gfLVhSWU+gWvI4tp6Dlc3nP4jgqXciB1HruR3uDLVIo/q/WiFl9GXvET5Be
bV/zvWhaaOJ1eEsDme3O08w1u9aNosCDBRIre3glrByKOJtfk53C8xl2izYajP6mnfh0W9MpRvhq
vJZ+XkS31z8c0RPAQMa+/TqhWL5Jl7RCoytfv/avR2zmIeiRYF9Pyn5nEVYKnoPoOSYXkIe0eEd/
Xs5p5HGL6Jua+bbGr4zQp9HxgaPgPiP34LO0Sd7XJufU0XyVa4mRIRnu2Pp1FBrFTNyGXHcqGo16
PCzvQfGSrKWCzRE97WzSyfWYufvYDD4OsgLLWwmo+7fIyN4odgeNad0o7s8BXy+nd0On9krwuis6
XQFBClZ0exf9zR8y9nBtktz9XK6EPKyuzwqVjeO62FTizDzPLEYyNvvMi41ctFuDpYADKXwNZcnW
VdHsWXgKNeUvBMYjjTqVmCQ2UruJJs/P2V+KqtZtfG5QK4W4m4PKsGy2RjL6n/UqkIeRurTJOP2q
ekk867V+KkTft38spKGvQLkqCkEOgWRSEkzRTMNwzEcxaFHUBnFqBcG8OCxY/lWq5R4gNs1OiN7g
Q2SU605xpPe+e/85PdcB0vTT/NkfTAhuEEWy25kTACGlQFOiM0vS94yR8xJ323JCqK7W5ZVP5OIX
hJw+9qZZ+kY3rSNlZeDLMNPPdhfNN71OkJp1WNY+4glpY73tcQTLp8BsjSXE129adZMclkNtUkdG
uzaMxh6INi9dERImudZcJ0tzehr9zTHM8omKwFh4VrpqDe9KzkpZthFTHJCqeLRQ5IPob9Xer/KP
mfcwfFcJR6OyP8eYtsoe2ybo3qlUB3uXSFIFqaTDuahMtoWB/cVZIb60LwSlyOSHlxPzeB9ZuWaW
Yl1z/+8viOb7csjn2BfJbXMpEN6lMRv7vY9ABW523EY2qkePGwoVkjXeFzvSwUygSWi83JLrq969
+nsYukJ5OiaOMUFi3V8doVdCVMC2Y0mb7kIHZ30Y+kBSPXYg2dttIky1sgMrqDZ4mGI+QULTMrlu
8srBW5fjC2zddbq4u0tQ6OmRb2pYVAYAQw8DxhMT424AbCjnNLOER//gElzQ2ra0Ppuh4aeRol8e
q6aqpKjgKPabXNQZ/fg1SE/DpNrCLMtS0yBCzKgjLnLYFPrUYLTc7TYyS/XrO/OYC1m8kJNMuvgq
u5nSgQB7Q+/P5z7NvP4fD2buJbFKpKMxh91bOTWkHrlB9EGNuFq3pcK+8v59bXcliy1EGm4wgDs/
TZREB8Tx11UE+3fPoz53ahdFNfepfMCccnj2Fmt5R6W4b6YjKZav/55/NRtkcPBda8GOOk+xFYe/
dLHyF6iS9t9FBj/F35dC1rzc6aoOIpu3P/fYw2u3UKbdDSdURC3np2w3BS7+RKsM4LfyebgeuY8A
2AfxOit4nEgOiA3JdhZ0itipvwBEggrxPA0+nI/QgFJTgmrSMjOfLOfPCbx03Ig/j/uTzp7UUGjK
O//4wRWKaDMEGmTF7ITIQYmAnct7otQpMf+azccrJ1Xtkt1I1jnisdEsdU+46Bz6Dx8yDYQQ9MzZ
qbftHxXSQt5jdLKKx1r4Xl3NiDRVEDC8SvNZf7P1dVRU7h2nwWCeEA7V1FrifuIckowVxTVunSuQ
87tn1UqlJHaSeH+U233Ynlgh7X8MejcicJoi7i6ajlHaxmCJ/itJlnpde42y9lbysZW4PFDTfSWB
pR7CQgluscrQ2I+yMH+4UyA/4rc+V4YZb8U2Ege63aErf+Bc+JF/jh/TbM9BKQ9IaEh5hhRLfcrX
mgASKn495BefVITxJxq+A6gTLTvvwyMHnwwdk7LCzU8GirRe7lLQHLEXEAGjhUEmIs3a9nhTwulE
RCiFfrZVxTTbayvRLZrFerPj/ZH3k8h2NW3bHziMAdSt5mzhHgMLHHzRFzPqkwjfUnEOjYR+PorC
wboKEC4GOmudFgqFWLcQiv49HlWOmJXSmQe1tTwZqdeEw+Y66PG+OH+gqwMLDkdJP4CY8UrKMDy1
OkADWKNvLI7R5CXLtcdswGFn2e+XNagF5TRas/yPf+BaUS3s/AfMyAdmj4QkC+ZS4S74MtWNEV4f
l3iOyUrgJjH+o4KGjf7N7r02yyEH+KspJUyVnubVTUEza148g+81+9GZrTNk/e1V6HBTF33o4rir
yHRsBVhfx81bXi4QjvozpsM4nmfbzHxEzXhVN+SQhn0L28vKxARufGcxSwDBsTs+/QA2nlqaLu2c
L1gody6t3psqKMmku2J2YvAdBg/xBiVcX8dt9qDmAZ4VQeAj2fdAF3t74Qsb9J8hWu4DocJTr0as
WUhD6m1AYWZ837S3zpY/lCAvpPNUbwQHlYVTpDQDEyQ1yFw8oqbG8tXzXU/ITvC/KfSyWCdh49dj
XsqqIwf7o3kK8d9jjNWBi6KzJNx7xgfoiepuQrAhH9samsEsz9BJhJCxkkYWXhrOVJKUSNmqRAnL
9zMrZFgBh7YYJybJXMkTejYeLYNRKrlj+mlknEhksqC+tgtba8OM/MqcQZug5PUNOzm1OiR68ztQ
R+ZmokFS4w7byVKFUkOSpm25DfjxX77JDcB76mRYqFGw3JpjKI+KFz1IWWQUnmwrqlTs+dxOQ5LT
mvk7mt1rhdGc664vQntAUhaV56LKYYGuedmfhgp7ppUXNPaezQfqecskLoJCLSjFQqyadZ0oVVG3
kDH5tMUBfnqfdGIwdauAwrvswB1e4BJVnAogjoSWQgDbnObKjx0yLgDYrtHUYLjWNhakIdN7+xjr
ya/HbPxx3XS4DsNKHHwfnbN0MVz6kVRJjKmY9RsiOj7YN1Z4RHsofyl5Ncu2CTLYWMGMwiUJLlUV
4kNZTys01O7cAd8ZTcf2+AXJY67RUrtCBNg4wfHhFhRSHgXcsKvD/MhuyUMMOzbvlQEXzz77/1se
pa9JTwGilbFe8Zrag54Z2sCSw3ToTTrcm4MZQSWQCmtKANsKjVmKvXxQZVQVH9NQKENc/VaptrL5
DWrdz6t1xcbbnSwRQInzOyIaXbEBrqJyPCkvjvMGnkGCCvneLGZ51VNTCKhibA57P7rtpZ4Z5i/j
qzNfYZ8tnmADI3Glm0Q7AXzHJHHHMJshXG8alxRksY6jKIREiJtnwpXuSqqe0pgcOoigdXXnnnE9
7Oiz42JD9xthm+PQhn8TN0ie+k7N7fMlerr83lwZVSXlTDx3Yo/zCJ5UfLz4ZTJlqjWSywjKvyVh
bAgwnKFFJiR5kU5rsGFpJ/IJ9cObT2U32W9XgxYA7lYYYCdj2ob20OwVyuPiXrytPr8DBg4jlQZC
k04OHlq0ozitKIgPZA6P3MwHM5AlZeE4xAInmhiQnI2xdiYQRoXJmf3siUiP8NW3J4mI1CyxE5md
IS90hxpg5pFQHByJvLjb+fYFaaZjV4oGKf/cSHd0pYKuate3xP84N9ll3lT8yTTS2pO0fJ7LZSLY
LARnkhHe4uDa2oKv3V10zkujw4t9/9w5AF0tMykM2N+EhkpxbkWqW9hVuXf7sRUY2mlxK+n1+YE4
J79gOmixpMubUSDqDXtz3ki46xUFwiT5ugf6zioCfa3iB1cOzBRhCrqlvm5wbMiBKgl4Rzs9j62U
ONwgHu2ZkYuyuhLCU6SYf5JrUEv4gshwFhMBSaa1WL1H+bOCvFT7ooRFjf3lFFYU6WBb8z6wRtL7
lIxfoc4XJi1d3/TW8oGH0Qgq30Zus+E7S+bAM+TUf55A0F4NPZbCvFamsHwBFwotbHtu9Bvc5MYt
2nYoL0bHy5xFsQNedBQzSNkRb77LQZGolcsdfM35beRXCc6i4xGjmTQ57+wdPgJUcMpVl5hR026b
A2xAlNGCOX0VM8/MEYQ/rc7y/91aOsu5fhyir5tIiPYkzFVNeMao00oZwetU06QxBi+Bxd9fD6J5
L/1e+JYFfB4JrY6b4Z675yl4Ybg+YOJLS2yrMyCFkpI864IN9CRvWX2cKwdTH8PtB2e2Eh9Bszwn
5T2tloJCXWEm3vfhRxVMgPNk//wszxRFqUb6qBtGScx5Okb1zReEox7ZGavAuT8A/iEzwihjvnGc
GgEav+vQ3N4Jsr0WSW26unLdmg0Pm94xMCgj45rDEpqHHnZ4kt+K29p7XMRJvHKvOsSdP+JRgCa3
aBXVRqenHqh7p0gQLqbsFxaCU4bAnKQ+hLhnlWctFCAz+A0/IdjgIiq5GBMN2lOygKzDgsU/ntcm
L/biBHfZbxFRQbVt89+AYx++j/WlhaIEJ9bE/3rdiy6gs56ENE+f8BYuTVXYvJ4odiERu66Ik46u
l25wWjfyyyzijfMsjHDtdc++/9+RjTo74l3HNA30LUy18mOkVsGCXP6TS0zFucChljPkYip8RlEZ
+5uk8ldR7FUQAk4Y/4UxW33RCdLs12Nmyh3TlksV90OquxV0/YzZfMjjtG0UTsDBJgHnXOjgR0lK
CGlVRV2rhhC9Vq5f12PDq7kj6RALExLTjkwLKEY23irY1xP9V4jIuF3OlBzPBcA2cOMdkFbYO7Y1
Uz8jiAX4OMrgUOiZXQJ0E+YWpov7oCyDDU8zxwZfPK/+tbPRgpahF53GCiPPmmQvH9WEcI2es99J
lud5e55Tnqj3X8qeJT3IBsR4E4+da/+92Kbw7+qfH6MG/Ob/Kn28MgFr7W/wWOqdJUfx5OlLv8TD
L6CqymO4D0MI6W8uPCZxOBDMUjs5EwmX1iBhcAsncV88A49cPXxWcB9wqexd6NtE6POres5zGzmw
cLYbZA7Dm8aivOXio8sBwuwWskEMADilQbfR71Hgb0CTVrScq18mZ9MTGUYYGDxHblfQwArU8Uxr
L9ER0c+u/CAJ5JCcqik9EZfiRHpZDr0KE0dVtEOTUOIw6dCcUS3RZ9OIIjUf6mtSWoublgUb0bdW
IQtE4F1FcACHMK+LBCWmHF0irdaFLuTyhjmPXBM8pd5CAAoepQHloMkBHpy7bhiR/9enwMS/dRAu
eH66EVBFh3uX0PPybOw4DcX3HFjZpXR18mWdV99j6TNw1D5Y/YlQxN4EFjtb75Su0KtXbxoWHMqr
ddxO2CecyAgzk4XYgDzOKZcxgtbo3a4t0XoUyU8K737UUySH+1IJuMHaeWGFTPJ+Qu2SouC4bgca
4KwfYmyiUohuYViwPDUPsV0GfqIuTWIch2w8vQr890ievh15g77TdAulAcx92DuBuBWu5RX+yCjA
a4+L72ewLNDftkkZg+53ABqwtzZ8wWD8vJj0Nups2Wv1OQ2pKoXsP3AOsI40DoOIarTxyex/8y52
lSRhZa+zXM3wxbHuWdINZ9uCvXJWrWNzYArGw0yyHbl52I8MLP+QIl3ylvu670DjD8eHvKEJMN6e
NkWhdseHze0/mG+XgJdQHkhta3zw2CBTsI2d7K8Ds84YhSjm1NFwPv6SkTlRblhLqbURLnjHSZn+
jXP94ZRgReR+B6oRewORjtSewwr7WqQHzkjCuO8F0OG6wfBHexcwd9mjA1XY/HgNvDiSQIUapvnO
H+JRxbB7+0jNiM2YHWph35iYa9EV1nIhqLSFplfx3UyfDb6JiTMwlwnOT3X7a8rRqO4jTzHkprpR
UYBXdOFDeWsglobSwjsp3s8rUs+o8laSCQQT0YSNWUm0yJzaM/ONXq99FBSgS5FpfS89qJKTCIw6
nIwUaam0omCqvmq8Jz+kr1l2duUS1gXOaLo0q206kevMjU3k499ox0Nlw/So6a0uHOj4rw5LMFzu
n5ZsjgqWs08wTn1Kwc0Db3T0lPXn0ajix4G01ihwDyXgeO/4qZSfFl9UDl5ZQth/AoEKunu5y5uH
AaiEx1wNkMEbTsrghmi8KdHOthcZkYNBE0PKzpVykwNuTLfUM5hDSV5jItr7b1JfWl610KXNEdFz
4/0rEcFvtW33XMEZgCGpdaC2HycL2oI/dLyj8AWjzrBJt6DW22FHtGgfUcTVVclTHSLYFLgzA1XW
jvnn7bVGxvEKyJRAmP7XFz69/ITKpih7Jx7HKoXp9szf+AGykAbOWj48Wo5h8ffuUhpa8XMqfGEY
yYZUsaGElV3uI1LbFONZNvFeGRC7ERxQyWP2uqHx8vS4L3UfZ1g8Z1NTjL6QntxF+4LCt5S7Yhnf
AwsR3EG+kyegumnRsgXWj1GJP6VG1GHoiOaa3zDNvphpGeSC2/29EDtkD+PrnqHTJXh7i8rDR5Km
jb/hqZ0OvUCqz8aMJk+VH0g/RPr8swOtgf+lH8nB4m8ghv0OXuMBCCyEFpuuFtcHRnpFvwglKS22
f+SH22lqykIBJG7FulWykdakNTS/vODm7kQZyrRJMcCsUG6LZT/IETx1gV0+/Ez/GlThuilB33kb
i9AkejZF/3w90osqXpT/VKvkUD6dlqvem4GpK4rQwLQ1n9bwLhltEohlkOvC/aRtF9x06dKOOabf
nbUDlGFrdOcGzkFEbLxdE5NKbYrsOFscilKlF8JVi1qp0k7QQdS/cJRmYFZaiAh0Cok71DSV38CB
esQwhwZHYodrZUniO2UneKxTQ4FjOXQJmx9dyukfTV7cdmWZa1MzewmahIEPNMho56SvrTpMPQSB
kVyZ0C8UGTRDXqWwhuIlhiJhiH+RIERDWj96UwZu/FzboJs1hUB2LWQ+rQOusERwUk5mCokXkSlK
aLSE5hkBNVxmauHdeDqMIj7Sr8RUzsmMthZiPbNtL+MgeBqywkh4UseRxDWnw31OoiPoilEIx/WO
ysfzhZLawFRRjusJX9iVJt8I4hIqn9X3+J8Ug0xETIWGo6E6SAESnoNfntvLau0TGiM0psNw9GAk
sjpX+sv9rmpPXgrv4DQdYG4vHRqyAxVovlRhJQPGMW5nAgPM14KJ1HqaRpHQOIov1e/Qz9JJBF1o
EsF3lwxXARhfPXL5kJSN63BmYFhydDZgYCUUILigM2zis8TiTdQmSlVSo9bhMll7TCiRjRmxiDQS
zA6AKqC3LUHVvKyC003jXbyxunFTeTxdPaLC1VSvBF7Q7/U0ZOCeL/lied7io/IC+osa9WezFsuk
E5WgM5z8QS+BeW15xXy9OJlKsTViwNS5ZMkzOwTUgUwudnrLLhSoCOzn/gXWNA9lQAvJx/4J8euc
cSJdNzAr4OV0QpkFFR8V+3kvPt6sqUfYj+r4CmTHOYQuD8Uwjs6Hlk2JxC9+z43ZRKSKXuR0zZzV
orUhX711bN2tmxUeGFg+oCSsmdqU99oS446sKkJjrWu8GZS41NvsUiq7lzbNYnpKRK5ifD4jZU6S
9PcqJNPb1b0noUVJWY4Dt0hSlmUr7+iUh/XKyZkSbR8w7Yq7tqgZQxAWiRy1yns9vKmJyIlaB3G/
0+Ua/PAdwJnqxYwLXZGXrxv2Hv4+wmEKGXvoWcc9NapuwHIJ714M3/kDeLOfx3NicFOchNsrhOBy
P/QsKMk1iKp5yAPYJlDKNXV1fdo0YgG4nXmnOWzqLmcbmaUxBjyg2S3+tgdhOBkGIAxUaiV/XvNT
Py8rpRKTmJsJqaKJRGzkaDz1g2wXqC3GabJLr7T/F1n55/6wvcshYXFul00tVnWB2iRA4iUCBQe+
sOSMax8LBZsSgCGszHgVjSAaD+SRHeXEKQ+/1to5zlro98PIRQIvkMhAjubu8EGdAr6sTDO8Pdmo
Dt2raaVM/cGelAiA06fv+WxWT47qoIPM5nutWzy0VDJRszwLkKq5QlwSvhjaPDWoEGuqXLihSumF
egEtbWIAVtZdyn5CYu9bcMZAjysP7VBKlUEBxVfcb1wYIzwjtgiBZJH6KZDoYLEHk4xYrtDLHodz
Nb/8OHzUvd4DexQ7QRKfnMsKXygZh/gyWwRoGJFsZZaciYCTyIZQ7HCOtAZddqrZMblb8K6znq0D
TwJgsddf9WwckHCcova5zQZ9F8ekH3oiY30x9fjudTfJEX6UCMUKhWB89U2T1SLWPQ02p2fwN8qz
h0UjVYsNn8a6hA54LyvmGeiwikeWy3mdTCZu8fQuGCz2UjEwRA2VbZs2WY0HUtWDGRWL9+MQjuOe
cLnaxyxeZOnOwBE+SSJDURvPMcUwCWMuoV45rDPGHiuIQa3/JF4nvDrA3qXDdSMmWp68NS0JazTs
o2Xk/Imn98eek+vbT/Kd8TEOYkPcYoTXHpBKym2O4jeNuvjUjSFrCMROAnQ4lyAe0En0vzaufeN8
sK8yfE7xX/HiapNf2vNOWnAUXsJKLyJD3YW0zsd2hNAMunBFIkndLIQNGdp2stZ4hb901/TuPbTm
qaSF1fGRaYIv42J+Mv7cTrG5djS5u5lChu00u7YM/fVEjOe3TeR5q6PB6sLCdEKuMO9nKv0wHkwD
+e+CXggwCvIHnmB2791BYsmz0RmT0xJrHwM42Tjt2eqFLDTZsVBU50jkaFv1GQyNrGLt8cUVVJYS
WbxHADB0KBv6rfWH1t5f920RAD0+8M3IC7fMmu5r1y4GC84v4EC6ZQ4TE0HpaVJlrkCVWxlgtVuB
5o3465aIhuJTgdoBH6NZH2OzCEKpg/Io80VzPq7gLZ+eoKLglw74z3s6GSg5+qlsBpnp36NOv83k
AY+QiVRTHTmIqoFZ7w9eF/CaAjfIjVlX/7AwUa8eNX/13OMre5m2a0+simwOr17X0sf/PcYQ13w5
0oQKiSAiSFgLKaKiJzBDj0fu8wYdnYLLqh0Gc2PG7UeyHjcAJpXXAKYNchkwgLe84RsFEFMG8sWE
RIdHs4rxMqDfOzi0faS2zi4li4KSekUT9XBkbhWNC6kTPsSnYplDVUNfY26xcER9Mg4FiRbBdM/3
9vdV+3FiE8/zNp/fXrn3g9RHO/JDzOdavuF+xxMBLKsSBIGRYDFcIQFeF/3v/2BgOKPJBx5M9GSA
BvNQCRgWWwEzhl6Y6pG3o1fJKmkiYwb89sBWZWCSErKeB8lW7nURsPaYONdouTXd7tYTcUspzcZN
2DrXwbRBsFx486fWukYf1cOaNldidWEG/wrJlIE+S/VULB58HRx2aJvaZkeSZCS7CKxQ72TqgClI
Tosi236pJ5TEhhfCtTFlAHZuQYCXKHInhdMeMTha+z9YsoyB/FWypaOJB8s5/akZVr1PUPHmJRng
88wxSCEMgtdEfgvqpUtCvJh7D+BO2//qXGrbt3C2enxt+Q7TQ467J799fpTX83Wo/qXXtuk894lT
lQsda2h0ZhxU0CSaw2z9ZZHhdo8obnvgmepoXovfPeoCjUM8D8vZQ8cBg8gAbinfcF6mAWdJkEKC
Vkfi1T0CWi0pCVGOZjj5j9+Jp6l0h5mXT/LPIUoEzJ/KNtw+rHS2PayeXxNcfhuhNX1Sx3gXMemm
HeNORhlBdws/LjcK7oip9qLYi8VQxPmnGALjUG2BHAVPQIbe3JaJb3wXsO4KTL+3HDvccVRPYhtS
yMaAECyw6znWyvwUPCoIcX8YuZ6v7+jCVn9UZNnr6er/Oa2HVBJ5KQwlghUkRxNvNCziiGs37uKL
ss5KAm6/v+M1I5rqvGQrUabNOzUyjixTIFtsAzpagQWp2+fe3xI6MKfyqne2ltGaVDu/jUC4XgP7
gjK3mnVhgId2sprG1XHAvjMFWilFm1LHwC/hgmLmL6fbWvUGe6dmvf6lNVdqm1wo7QDxD0AR815q
XhU6Q38dkmSHzdVnMAK7s5hjch4GACxZU4Jf0m6/qEBeDTXMnqpRUHCS8Bc+urH6om8rOzkTW0fP
OjRpqKwBgFxYWjgfuCSwpU1bMqRZcE20X1ywORq28Qva5J4itf56uRkVt/VuRMr21WGIfJxQRxqL
GPgfzuuqEhI+S8WXFXeJc0Lah+YwWwleL2IoJEWyRFcnzvV64kpNDXgZ7QRcXJlzD809C52F1O3Q
QQjiKJc8onQwECYiHRD2e304hSr+YqV2vTf2Ec3mMsBzOzk1VP1488qk1EaG4hEFMW5E5KXgMRZ6
ILNEtmfY0lGEolgiyocxAyKmmT5R+tZaPN85Y0Zapqt+/ZADLHW5JjbALgnZqkNJAYD4Wd2ziC1s
cYV+2wfi+CpPh6IvzjTyGpQ6ihSdlaN0/5v0gPZOYUqkA5CTAgwNWRNNbtCv0RjWy+z0DxY8JnN2
0Lvv7In+/fZMdRgTVhATZ+Mp3oPQC5vewA9xyOZ0lDSJ7PRNfmimXyUNfjvApRLaJZPCov9rr/iF
ul0DMFf/XACzaMiPdcE6oCRQGvifVXIwXzsEeO8OwyUMhQTLG0uASpF55A6jQz+8sYdIY4xVyezY
ZNu4WaFpCH19zN0uzn4PjxabbIqMX6wtBDPWKRTffcyJJMgiluVIjXYZcSzUIUmI3+GVeHxSV/S0
BNjxTyxchwlWBq+qAmlsJiszXN/nvhNtPAyYVCtUYZLHcoi9lO0tln33RjvEN14aYbgSK48toBep
xssg8Eq/r8od0bZr7PKFhfFQtSpcNIfeD+6VF+kAEjmdSRSRvSgjEK0El8SDJYQRZDTlMBl4kcHL
H04TTOdsvzpNP7761eVmE/6tIhIPIaidEHtSCzMIoCYg+8lYQ/aXVPDMQD8AjwXrgQiOJYz2pUWD
fMt77KyOj07ylEmG4+bXER2sWolMiOAwTX1ADiX+alxRRDuL8OFNQ4yVRkLWN8/0xCjeY72FakJq
CT0PKZ+qMxGu/4d82LDo923KzXAUOs8C1qH6eOltz+EjPi1BGU1onaC0+M6GtjrEQgD9r/66DLgO
J+/6dEY0jtJSYIgmpk1vt1e0G5ilZZo2vOmdbNSG9S8GO2cAVPp0mQrXLG3Y7l04lrpXg2TaJTYu
bDT0iLDwCliO3pv+0C3LXTl9aDgRs+Pz1ubmeCgcLM6dh9+XvEXWRcLSs+cB7xlBB/jhTYnY9NbH
qdIZQx0zIRZqZ/EIG7cWLAxEviB71+R7mdZsercB7k5bMUgtIWw4XHBp9yGWCP1xBUManzVhueLj
eyfn0sHlMX9ZtvAJ7T7jyyd0KRqKK/my6ciSg6pwHmqhRNE3y6bHE9bScE2D9aWbi4v5ftx3Z6n+
LHEhufK0Dk39gSNm2VgCUKCBRKNnpXCNn968Rw2C5iL6pvkmNPOJ7+HGvE6kvWzInY2lN2y4rPqy
mUIc7XzYy8/Um4GvHHOc/gTEy/2KCesoxyk5LMLOXqnNr5tJnCHXqMLTC72yI4KmvTM7MSSUEHzw
R+VbiT519UYWfNOT/YWmOlHBARz0KmIuw04fsLnlSSFe0S1x0YYF0fE5vJCPpH/d4D3UVUpmZOBn
PWfngWwflCjM3k6roBcmoMvoxZjpl+AfBgDbfDVlBtBVOHjQ3QKqxD1Z1GKpnGBbXHfw2KriWmEU
yE3nTTNBeL/HN1aApWy0ICpaaqwTqR51XTpFbRmhc4artURbQMa3DVqxdGUr67QuSobqlbVV8o/v
E7NcPGM0+JSMzJrTs46dZx02Zv/EDqb+sdV+Veqdl3biXabRs3/HNS9aS9v3xdC7/+RRmBzrcc4R
s/9iU14WENOkvQjPLhGgYP6Ob3MHPJUa5D1GY9Ro8uF8jJabbM8wi6LBBAca51m+hKASLzPbEHO0
Y3Zm/RPtw0+cy4nWZ1Q1MvFgm672w/YMPMZLwmpvOqrPoXlTvLh9GconmRSMVyywuEQsHS+iurBK
NgOTyiTvJVHkjJhWgwLHGo+3M7E9tGVC+MSXkijUB+H1nN0gZ2RenCa8wu3iWjLXaLSLsbTMCuPB
LsG57P0QDWkemiFyNc8ZludeA7jEnWRaxMyPZbuBldg4/tynXtDhCqsua+4xHYDGyhP+zQgFPcEs
vbipVS8ylb59DKRSV4c3aj/Ubm7huGCw8A9rfcKdxLGkTrynor88VGwZr5rdYyGooRNEfjo3B3Y/
O1andhiXzG8szG86XLplPOrJ7noqgC4IIs23xeo8gfIGNpW7b0lMDMlLxjAV1eTahFDFmwDwLMsf
gFb1q2p3xpIsEayyQxElw1u/qiMUAmDiPK6vQfZd/BrAt7fGPXwWrREFK7QTDk8nPk+Gw95wbuR2
0hV7K1QvGc5LkQyjnPUaBWcedNRyT1EDV2dEI9mNAvj4FA2FpnzebXGwnkEQtGaa2aegnqeMP4e/
XOQAP8uz0pTbEFGzvdYuAvvp75TJvm/19Tz0uj/L5GRzSXQYdNMvwLc3ZGvSFkLblktc/W2SBy6i
Z5wO/bSA57ct8JX5HFW1Z6Lo8q41pW18gWYZAZ/Moj1sp6D+XMLexWwRES8Sm7oPbzGgzxc8rxyI
OVWlTpkLYNVxuaId9v/uxQk5rX5htuGf9InwfrOBTIsRWOXZIXtaB554WjguHuuSc5sxBS2SmoJZ
wNj595UDIkAjJoaWA1+mUu8Mu7mPNwOeJH/EbWcC6IHuVppQBv18VaRKbE66xxSs7nLaxlyuaQcv
+xX4Ciju363475gCpm3reo8wvUZzCPwBjYktpy4EcIlD9dwaERLcczbUnuLX/hlEPQGERf2XO5DA
HsJkSwFT3UrQaUUPF0IoYvpR55BP/f49N85JIdkG+yrv9B/CntoPYT7PXcLE0JrEnaAYw5jP/9m8
VyOYwVYIKI4tbbxRf2XPzSy3iNA6anBGjZQF0VJCxm6gkai6s50dkWKEW04P6njl9c3z/Vi3lGpk
Hmi4vDfGsLovvBS3WEkO73n0D5guAPMT28YdJYsGE7MptTtVeBfCcKjA6hz0wRbBcnB8tLlM9O6s
BFY7bY0muH6TCp8wLrpsFLDPCoi/F/E1CmEYodS51ruEQ7VXZAarISpdY09zni7G1MQ6vfqmcDvX
E5zrbGlhpCl8xMva5pj49pjNqD7tIeog9eF2dXfnDWPiSledd1JhDdP0sLVN+dPtY/vCL8j0QZ96
TladerRAVSBp57EK/PLkU8Bb8SCY8jpvcSAc43VUWyQqO0DskSWzsFwqegxJcQ5xv3kKoNgsrTKO
U5wto+Nx1mzGVbRLZgs9ghYzvJa9eiVyfQGsSIdklZt4kCD8+agQYaUx6gWcQ6bC6WnxBTpWKNBX
30xV9U1gw5F82wMgoo4TfUqOB/japeCLhWTCkyrv+fL2ENdLT5KybHvnnoX3IGBPgr4kidY3GGCe
1ITHiwn7FINCIZVYicDOFvk9Mz6UZWpR8njF9LfzkLqDsX9VRqkTG9Pa3s+GBq/SokKsHzHnm+pl
Xn/qwvtq3iAfyBmigaKKqho6EC3C+YfW0jYCBAs3ztlNpG1RgIoqTsQS1enfzL0LMikKOTyECeKE
vOKbllXeJUsqlOTwKqMOS7Qtj9Dv0EgXGEOOtlUb8n6mJtOjalUw1+XTqu1viLOYWpy+8N/OZ1V7
4uJeAIUKWz3Uy6xEjr25iX/6Bnbw3sOfF39pVTFpUaXDPTfY/luVVh6BmyB4dIZzVT5ay58uHsFA
hqyMcwT+OINrCmKxCj+SZC6hfBeQy2itPVTOLBaSdOEzJmDuxe0ADKFDDz9DZd5RXD6jye+aY5va
N9DysneiggQepqbPI1az5OZHnwEoP2khpVNyrngFkE5VVRyPPLgAmniCYRQuCQNjpmRndDFngKJy
o7oMttvP07yukgpFalPpMlNlE9nS1qLw6gn70lbM4LZ5lYKCyMgFTWMXdMmMl3sttS9hbKG1KoAD
e6NBY/TDHwedjLarMBKFdzU/fmTFCnzPW8FPk+vuswDF/hztfmq/0+d6NpwZrWziSMVrCzWn7r9o
szU9QfQEfjOgB4EKptdevM9TMfo/JvGZz5ax/OHLOJ3vte5KYfCUNIHZvuGnb6My0PhciLhQwNZp
9/Xfm/OEoExgsgo+bSVnFdUWcX4TkuqYNceT8ugCCL1x9Ko4pCINTFAKNxVPTm1mkKuvwVv6+8bM
Q7EU22of+dudBXHSdWdUnRAdhUJe9lopW/7mmp+sH7XFSzmMWkA8CEl5JCz33ze9VGpEfX21k93H
7gxWO6+BzwHv11891AeO0GVAsCRjVbRURM2sLc1NPwExexdJGzTSoD/XLTNkW6MmmlGu0PDYKPmu
eSzEQzWri64z1DMgkpYKpofoRyQI0q/D40zuiylTvNSvIlgwVeuhSAuk123JRnjexhydIvS+UTK1
+i8o3S2YScYmwl5U32sqqPCclEb3M/Va3dxf/gqzr1eqBjRLLPk81V+L8MNW5cu/uaQrPWU3tcEe
s/9LLOCOhWTf27NbqbhRK/eKCUsSRuKMd4chlNV7nWOabHku+a6m9tsdLC1YZzxWaDnQHlWYAjvU
rRcb7TQ+Vm8NCdau0RZd+y0l5/ae01ntbwDobMVXx0gO0XPOnIhRi6EN/A5ZpUmJUnMwHmmJj+xJ
PedA4sDu1Ok2ZrR4WPOFKvuVJE4VAyBL0XcMExTNoNXeb+f5jZWN8ADvfWUZIIjJJcywinvcwGna
DrFb16MUiF7ZoKDe3YWMCKUqjluXO70ipBWvxS1x68ANZ+0dOMKuvrmvi+CvUEUskQ2D6SZDtNI5
2QxeJLXLgb7yBcnMJkkrY4cHvuHe50mFBDmpgbsTXSOVEBB0uFkELHp40kvOAWRQkYGY0N7EyXTp
htRZ3qNmW7qgueg/5FTOlPd8eBmUeiHszA4SGftX0xur0TiSJcpfB2ZML2x9Z4D/507orTRxDBn+
V6IMQLNvSEL9jmnQk7nVrFDp9MCWjLgZENNHsyzE430lHNixJmoHjY0slIT8m0z/DW7cON4/p1Nx
8LvH6YBq+fjLEeTHNfj7orATuz3nanmqoPM4Xc3OJgOEES6YjAl5RPf+KAFbF85xjJA17AWVCVU+
AgvsDKCCX4Zhs2XQQtGYV0yeeP9GPRI6o3bUY59iUbA+6k4S9dSMNy+NJaFZk9R/F2nt/GY9Nswk
D0c6UjyPPPUZhBXxxFoVoywoQHfCc+uauCxMiGTZlDgNql8A0pEZ3SOaILl1i3rObrcAW0DUnh7Y
EJo1mGLGGWvRIfNTa23hSJUpTHCKpUZw02IDZx6v4TsEhg6om6vhcAosLvpp4ZXOFeoOI4m9nf95
BrQHR0pS14uhdVTUqvt0NFxM4baCJmmzlVIl+lcSPdOHumPFQDtcZ/vhgRSr/ebwfFFpGuTERMSj
yD4TL8W8A86DYOaYLCA973sHhL3EW//cVNktZg82pqP8AyJfdSJPDhWISs+LV9ilt5GKGobY58EV
Zbd22gw+d3X6gUJubjaDLCKhMBcW5owI4zQgkgz49qS/hBdwlyLiBbjWFhv/nzlOmu2nZmTDDBPa
KcwYGxq/0qWpIO8j0dpo+wXzJ6K9P+DVhSIecSY3/YqWhRjGzvxuSsB+1WCMGL3MDoxKrlkm7q1d
yHlmdDq9Oy89EOWY701KrdHKSjpS1yN6dFNlKhJXYGr9070mzxu++ImpeM5RrWRxOLXmXjAL3XEy
kp1p+8DuOWeYYimzNryLKR62oSQsNNHf7SA8RqH47HLHg+NYKZNeUOogke+XJPr7ybTGgprjZ4L6
+ERGzRkHQMf2fX/Zm3zBlwcFY47xVdsDY9F5P2Gu555pe8/kdYZk96bYDEW+vpEfyKa21er7qk2n
KmIH3kRlbj+sULtQswKNWd5ZjYdkwlFea9rxLfLmCRhwdhA8QsYMw+X+zorLDrOZlawDuh1hp9HP
WjN/b4/kDfOf4HoodkHANhyE8o4sflJ6aICCV+y+rjOBJ0bTbG+xLkTOcQVcpKNlFDtHJ6JK1Xi2
XVLaHYvliqLiELIIdNO9+QEf5JO9sRAs1MupZJWIuv8dy0yexiN/YWJq/G0d26I0L8P7433cOfz5
OJAN3wC7FG+P2Pz4F4s+PwrxIa7RZxxF9on3Ijz20VV/nwmQnDq3diD9XmDca7vOgOKzJh3337W4
sbjBHITTkbkkPzkS8N6roA35+HIsqgyeJnS7yuRTdWXXHb+W1Gdm4BmqxXCq2qxrWi5US99ADBQp
0udpA+/71/vNineCVRjPh5LdF1MNYk/pZMs7ozzk5BtkUCgHkKyAI9BoJGrbz96nfASAfPrLOQ+0
TgJBq21m7kbp46Ck8lIN+QvrhE6OLqNRhyUd2qJDKXK8eN6WVcSUj0ZWR9jhOCEW9P+fxkuAv0qH
kuknewdaCZKBUMuxA2bSsyAizGjQdbbRcxhHMyR5yC1wk4O9U7znetK+E5Tc3wf2y8Efqy6X3Rbc
CqU5zp/PEqA4Tc84XN7tebKf4I1PtKY7gPvyHhDBrv3cwsGI6kzgU9P64vKYR9O3Dj1M8rR+Wug7
kDQ/i42jSOa/iIQp9sLEZ9uYUKXFbin8f+nMRFEjchHd1y5xY7CGPEfOTAZJ7Wq5fR0+HLcUsAao
XDGAoCnzcOb2KiLv8tyLnEKHy38jtRBx28EM9kwi6i8RRn0e83+MKOhvV3fCoyz9AimQapNLSr0K
HTFvqRLlrMyy5fsn2xMTFYcvfxjkRItpQFVXxnG+IvUBaRdhG1BRwidP8U/0Rx51bzUeXHYK2ioi
rMFE5e6rfB4N25DVxvEbuAmWSPZdSrtmOt4FlslVreLsf9rP9tc67cp5YvASRblSCM5ZIozCHzS0
WVAOLizhaTzZObJkHQpoNJ2y/lrh4rAaIqsdOSVzjcdPG4Y5vlqIwvoL5vVYjWdQ8qT/8QRvNTV1
oZvdYxHyk+GaBEHE4CxkepGkjEfluOw5JbJeVjvPgH3JLvyyxNzg27jIF/20EdvnsW5X142fOOcV
pHIPrTk5/R6XWc6xE+EKmylfz2pHSRGBfSLNPFxpoSRPSHioQ8CoW/PWBhxEV/+cVOO/ZHWRk569
cR+Bieumhc5I9UKO0mHhIzHMTV6iu4V7PV7/zsc43r0EFwlmNkyxBQTYX2J/cEGl8/fbMQeefGbF
wyUIX352G1aBQn5RUp/QQG9S8wLV/O6pOHGAamcClaCJydjpLpiMSrkoHc/x1d6Capd/cMEM2+gq
AbqRKZWenUvxKFj2y3C+PxQjLpACLURCtjf56tElh17HnMcKpOpg+oK9mHgpOmcy8ysDzFUZ2uun
djtJxgiBNRdvIFVupSWKkFDdFwm2GYeAa+oHtyP59Gej9ExzImvAhBlMuBZ823laTHKjPnhiFwxz
Um6ClZMgRm+wzI78FmfNkrRl6U9ozq65pPIfXmdE58OgGO349Tdza73IwNP+FNucQbzGtVBbruCx
/Ov5ea5Xln6bCMdwDJKruqQsw77RnXpevcEDZukk6cZxJYlqxzMkLrByizN7ghO5wtw6YrortNI5
lWjp3NYoXW0zQbhy8fqMN8+8zqnnLFb2CwLaFK++ev1EhRxWaLy5gMHmon+bHjVcNAE8Nx3emL8L
4MqypKFfHfyY856GDKBO4q8tk6i/gpzX0j5rBvRI/RAhD3cP4UG8YfFdBmk8GVGUmzUGd+SrDi4t
izPcLZViShZro04VI5vVlWv9y3kwVDimlczYFpG4HnmA3/oDauFn4DW5yLlp0BfeGHlFHjv9+2tc
6JVoar4sEqv+s+Wg2/2YyyvZtsYx906kFOEF6d34ZfJJSPugqwqqi7KtD9FqS1UJwPKL61gJ0G4r
IqBs+Fe2z0Z2mTYXkNA9sDkQU0USftS9gKEejMF6osV2yuby6FI6K9mwbbjF0LOjYGA4z+4Y6//m
SB48lAEEfpIwQZCJn5ZlFFJj9dbOXZMvBhdXIKQxrmXc3Yj3jOb08r4vCFSjrp85okcuPt1JWqCk
ImiRjFM2F5Lneos7cysiofZ+yTJpldfTFm04KvmfwKNfNyBkcyhEPvZ6kKXvqPCmACdOfAUVo5B3
tno8tScKmvQIrGGdBTTF5XzTXmFIG9FGyhTwWe1JXu81riEsCs6KLN3WB/IBKuu4ef+0/0dVMzl0
4Em+R8zboaW8iC9sOnhwZLPrGknEaG16xGBsVEfkK8hWyG2mFQQnBE7sLfH1vhagt0sMqsAZMkLw
Z8SSCNPYiSFK2F6lh5885e8LVC38Q+YucstYkA9XsEFY/2CB+e878pkMcN3/KvNXZEqM2JtA3XRs
LO0LX+InmAyQqKx23p3L8hvxS2pdG9yyJXkTfIS4WQaXwGvTb7qEbaTSDJ1WVb0y7GNgzc+8I9qC
cs8VkIautDph+ym6pFL0Ucc7uHliihQOv+gIGtfud5Q7HMetu2kWrZaUjU8IKjT2IwMt5C0SSJer
TZThAWOIKeqAHG++tGN5dh1Bp25KlH306Xtx/d/GXm9nyQauX70CrE6kdPnNgIHjac5tONWAYxk+
ihO+Vs2EvGyXs4W0O5jiN6haWHxVB7mT7jDeHRnUFQJz4/DET4WZ10RtBUC9pEPBgP0PWZNv0NpI
4BdS1ClXZjaqXT0lkd5pp5wJy2+JdZzX6ifvS5GcgT81m3711b7w8Pw1qEGtgwaMxYhM5azg9Elr
PHze8qztnjMZ57Qhcf2AVzKw9ubSk5UccH8D9jjHRHOUuurJqn9HRoxzi5d2ur6mGL/bye4qyjDX
FhtYtzT/6s1WjXhgbSG5hQahw8VE8d6YZ/crxkPECj/jFfs6Uv4npnVX1Wk4zVFMPK0gy7/V0wlR
N/Zi4IEEpnOmSZ9BcyNFInhSPvsPV5uFYZQynP4c0QC+C14XK2FOaayvqoT3J8Nc1cq9gyUedWuD
/Bd+OzYHAdP/oPxxAN1rYlDMhVWp1XejXuDaWHvH4Ns1KRT9A+OPICHZWuu11k2J/LLMn8p1rqKQ
KfStZdmvNb5I1Gj6xZ7WvijHxunnOlSBMv8+8YpSm7mtPx4TWfnkmENQ/eRKrEwecUaYuJijfEyI
/RthTtEO1xVZxbdXPXBeQmHxV+NvhbPgwDypH+Jah1KotekcDAayeEh9VL1YDVgi/Xb6RdcCjvM5
+P+hlp9xAtQ3GARDfI9otouBHvdxc0xUTEfmeUD8iA0H/eR9KuQDwSqoIjde07dLNq0xYL91zNw1
jRQQjoUecIWv8alNZM3GxvcOR5ljOv3uTjd6pqR/rht4x2EjxJKStatkMyHxfBaKpEUhdK1abKAa
RhGp04An0UgJCDafRTG0EIcw2KY0ckK4EK5fqNmT5LEmGIpYjWSdBB2Zel6+fBvyqUlNjBXRmu45
ykDahJDn4qnLy7QOTvW4bIrGQlynQrB4+BaxiL3dJCj1zflqukH+yPGq0pV5V81RAiqrxIsMBKvM
ZR68R5foWQMfKVD1oUsJF2b4mC+HitFZ9YXsGbmnLrpvH7hO5xUPrOwG6tJYAjOBhf1+uwxUa3VH
tAGJ9hlcuC0JCuhqfeFWkj+gTLzoNge1Y86U8ImaSdeHY6wnHE7hGhmkzJgRORi3/lbqws29q2W1
vJ+G+6bsqAoztis+v6wE2kZyO44aFC+WghkjTTvx0p9ZUC4EM/2702WVIvtzRhci9Tz4lAhBqC8Q
wXMvj4ssN7PFET+28Q+BfIrUpWPrWu7SOehUuDW6HbLJorD490Ku0mCpxGatahTGy7C+ROCYf58F
mZF5RmNVvBCdKYJMV9+eG4yYavBIJ1v73ebashNGosHlWEKx483sDUbG/TRavf4YI4EMmON8FMI9
/1ufLHVPGHmZKf/zKyeDb1WxvYBHABYnLzVRCpaElcEDENe11A4CsZvdTDRB4BknBMuFPYcyNzMa
OJc5DFcLgD6i7g72HKnbNuWnG7B2Ubg/hVrKjonLnFx6uvZOLXq2aGhooSveaRUneDhEM39mNL9E
dhdEikKW/EjlFB35G1EGf8m5SE6cb/D+1wVNJPFdMBAWHq8s1nFkk9J+04eFIPdpwAcYEN0A2bG2
tmdhF5iSDyisP6alSkqx1ULV4u0NrQWF1rHpbNE79XQiLp7pqSOtbbmB984gqz0d1/e9PmkGaNyp
GE5+YQ0yeZgwT+S7nVq2925/9u3M5ekunKzKdRCn4+TGTWupNjyL5wmXWLja3RwRat1zUk8tmtpU
DifHFvrQoYTV7XehfZwZbEdSBJ7/RlhQnXba9ZXQM43Ym2CJ8rYpO0mJxgtfuM4CBlv1aThMnxai
ldpU0E10lRRQK05SbJuzKzZtktt3xiiP7orCcgHq7BqgmPqWrt/YCNgwt5dBAXKezLWYHsJynPv9
i9xiuTHxb1naTKMejRN8SXheNPhC4Eldwu5bYiL9J2GZRRVvrqIUWLk4qiFVG9eW1pwfrl+VDob9
uEL1YHXRgwxxVlqJCngAclmOKhZcDzrBsL0LzgmCIZLXDKvQbiSLgdnwdzY7EPfjEUnlrgyZ66HO
vXgeR9JYYrHGNIJqrf2DzV2Jtnf+sz2HqQPQO7PkBKX6XbEoJBghUKHryBK3dBsAl0Jg7FFEnBw+
vUz1wQb+XDfiAuWK0ZgUDnm7N4p+fK33RVNIuXPj/DT00EE4l2jG0XKTdpFKQoyAGEStzx6PKbnO
iOvrLVaI0nfW1WNAwMM5A075dCc8ji+bbLM8pLkF4blnpOpExXYzJ643N95aWVjlqZLl71jxmc4J
cp7CODtk8aEOxq9kcJE8yyfsgYC1wyEc3cWRUTwGSbY8q0o49YIzsPjdUpNvk6TBHe7qP4x1ir1F
u/XefffiLA6RZP1amlTOxKbSv7lxKXt8NFe4ZCt1mc7j8r8m6CWWfPDjQ0fRlMOuKX/x6wuuSFdV
/2yAVqM4GYm95JznxZlDuNQ03d7onKsEqD9tCRwHYGwb40qPK+mZdgEzqPzOm9UcD6tenEPCyamD
jw8i9cgXx5QhKR74HX/eFlJ0ahUVWYnLpyCGMnRQhnf5sD3rLaLVs0is5MPyo1MC4fdDM10cmKt1
ihPYbCL4YCCz8Y4jl+WN0CJY0FgxRZU1Ja3iKRqXHQYSYpEzP5QXiqur7IAB0zI7LoerJQu/hO/x
u9MW/oimJ4kIktb+iScpwvOmj7j5duiG77RFUBzxoXHcmZ+2i0Pw6g7monqvL3rgtsjdld2nlPzl
+hw1vYVAQ25nau/RfpLJQHqF7BK8T0S1Htbrz96IAhI3uURtBNMjlftCqPy016A+mrlAGZQTar1R
rseHNKZtKJOxSkRU9NYF5Sl3WXvBZro+ebmPZRaT9ftNGrYhSmsUy9enAdaI82mTvV1llsHYSmUf
UsW633T123/geErfB8Qrb+cBkrPeWaHX+DMHf2Un1XLMKlJaQj+pPw1ZYQ7C+jWu8X4hrlbuEkGl
Yc/6TVGbwPjdzEqyaMXZkUpZSFuD7n63RxeraHE/sc0aRdY0MBB2TQzP7YGadryGlrHee7EhmBvi
c2FzonMaHFvhJ02V21p7G4chFLwx76BbF1+8yDbRnkr09QRjj7u5GhSASaIusQz19s9k4wJ9SwAj
RtRBLQSnoGREwSHTg7GXmJvOtvXUVFUSYnie/4k+QNIq88fuYejmgopRd2LuMaJTTRZ/c6EvKQRj
Dc/ZdfAo86nh0OVmSclmwzlF/wFGjLc6+Rcd25zHfHDMwOu45iLfqmNc5QKGevrvLRWRnFtC+Yty
C0y9uct3bBBjxcdcxk7Jj34RLEthl8q4eJk0bkp9RXFm4fENCArqVff7bm6qsXXrQBuSCKtcuPaX
380GQoHnSJeMobDX28faxbD0l8rkqFi6Jkwi+mAggL8HcpueUGpCdhrBxnhTAqWRr3NTsuyBFimb
84SdN2J9/27p5K8hMZb7eB10XvWZv3Lrq31cqX7XgrmLbme2q6unnVIC5UsB22U8mRlNxQaXDDQs
57ND/xeCjSIsdud/JaaZ/B+Ac9KzmlgZYG6GoD0gtkL+tj8uIW2VpbNMT6HbGHsY7s0TGsITBe7e
jKr/GS2x1oFRamCSRduKmhbadf+XiQmIFJ3/mHLaI0C0NGHxdEzavRCAFV/bdDXjlr5BNP+PeRr1
80Hz7G4u1bBdDQfrahZuTq5257V/RYWngLMkWi1uc7jNYzVrhXSntRzRpXjL/atQu6XPUzLuN62c
h1UGUgUWRctukjJ5eymLSdJpG4b3xiBY0P+2lxJ4ldBSR/jZEmZNshVyFX/xLMVprbRNNt5lphZG
Q6Elr2L6kpJf8a0ZsKbsrPSv0C65AbX84kH+THGwTKRR/oKgdvf5f+ZOqh/Awg8WtKa6qfYmoMUF
qRUInTNc+td9CnqlBepCBd1KeeTmS31HThkldUNRaCnBO75HCR0x/FU8x4YQQzREsO2CjYtejFdx
oPRaAIwU61Bse6bi7p2prh9yfoscD4d3uDNXHBXzffRSkJ0NsPBYfd9+YpI/4lsml77PnUGlHovu
FEu7MrQjHNMPgd1POycmTkrIm8QCok60FiofXwCliBV0PA+2LalMO9f1vQWtYG28uKE136YNx3q8
G4EqxgX2kDk8unfNi5eGJcmCtONERSUquVidGh4IjPy1Xbf+ExiR66JgRDbfP/PamDXTFtxzIjXI
Zjbi6Qu2o8BZJKEKxEb5cMr88FmQtiDHhCQPciQtgCM1hLIMuD9A09Lb4J9tGuLO2XsJt6EQXnmV
NiKHger5LH5tuQ9P7jRX5Og6yQosxIxMTaC0NN57u/j/YC7DVrY0NHFOpxz75XkDfQfochUe6tlC
8fQhlMVqs1On0hyFK3vvfMWNNED1KzhZKolaqHfSrw1MjRo3D0UFEKmNofD05YXmN43LhjhkkYF5
Mc5a4LGym2Y/qbA99KEXvmWUNf4r4AtK0iI2T1HZdHcwGwjQ03/cA18UpiDQWDttCBy5mlnpdOV4
U/knfzwv4dY2UtlldgCBMpXvSD/7HnuQZhfgZAaCC6he9bE6AUn907bAWdahkZewLSquy8OVFH1M
IMFmgDHHwGJtVf4rGF0zf2HULEBQ0CojgMbQRvTy8LK671GPF/iGAs8JtQPk+HQDe1ht/I1IlaSi
DDXNlFIh2PjfCMsCb2q0YAkawWm3u6yJlc7EWipBg59ZOfef/mmNIYXmMlnIviDjvKov9uWgnL5V
O6o8Oe5kWPiACZje7807SYv0oePd/Y37qikmesacv/gVZxs7skCJPrFO6G3W1YJZ5VeG8O6ezoBR
hu/L3aYZuk9mAAGmLRXOPrURo4YlMFY+LUosmdGaUkPRBoApGvs+FNpzXA9KGxOZKZa6Qpc10gSF
Rh2CanBIxOa16d5b+JwspOkLAqOm+c9DKOVKjDn7sECfgGTCYnis10oaLTZU+mgu7YS4BmogUyPV
Rvmx/AwpLeQkUol+RBzHaVtGO3c1f7mEh14Pk+x5qJTlPeqEI3oJQGbMxWiXjXyB/CQpJi6DcjMT
DQwU0875uNdPUOW1ToqXfH7ShuCL2pGCU93CjJdF8sb8hn4DtJqxI0uxnVYfn2chAujem1o8597m
aasa4oANyclk5f/cKmNy5MznQ08/v63d2gB3FBU8hyMo3ZHmrv6CikLkarfjetmYgaiU3Iqj5WEr
LXRwlFasbBYFVj8btgJSM/JfZgtWfMIgcZH7goKcH0SkSqg/obVlJkxk5V55tObNaMvZQFb5+cXf
wTPiuSYqSmsk9bdnvSH0TadPF1RXRbNxXF0iZNTMD1+DHiT3/x+8HnjhlNWFoZ64kx+GoDyzfJIx
j+7mEgFJcq5BusjvX0U0DLVtmQODiT14C5L9xWPRGGsrosd8t7U+OJqWHLppVMC26FbbbpK9XP/5
CobucDiWH7uGY+/0I6xljUJFJkok/P/HmUYk413OqUna+6FITM1yRR66ilFKNUS9ad8yvn8DGGtX
EoKdpNS4Wf2tEOZD8Clty/QyXssxd4h8C4G0Razfi+D9U9xlxq/98ik+jb+QGWJfMaKfOlkEEDIa
LfCaEvqdFM1+XsDXsp0NeJ+1GS+kcsWOTOdPkMEB2gxt1s0UrT/hjHGokpg7M/mTsTAsy5SFKn/p
JqxnuutqxeNbP1gfF2ZCYJoD0nfb60n+anZoodQOzgcVf/cnJkPfJ71JM/+4UR+euZUam6HUCNdz
ISaE/W0g1ZhjQe7jB2ceoMZRxHPRxVuOPXGndYZNQnjDwOhpw0TchnSV20/YQhTvOPHQ7ZF+OCIN
jrE9ovS4gI4/kEDUH3kje8Zq1vZE3W8A4JMcPRFF1/VNYzWRfeIFX3jrANv/nso+z7BdTO8ed9Sq
WP2Kr0t63CjkpSyOX7csecwuU6GfepFPKYpujroKaNOuD68JQnMEoPhSao3gdb4soQj2ke+GqrKn
l2Mz3sL5rnijj8QpG/4uZJPEpe0owf1tUGnxYMyYvTiSoC3GAyLyrxLmgcz4Nv5bHXnMzXqvTfp3
h79tISk16pCkaMZ6B1JmPOUvxyJdsJFeUfAhiVwEPc5d4/RfZ2jENSuCch6zZ8vqp7ir1E+pMX67
CPZUiuxGioiH48EiLHdnHGo9ozCRMHhsn6pFmMkw1aRaC1unjaLRdiZFZ3YloZfvEb8zvGWACwns
4Q+tArvwkbc0YyuIHwxhr27rhky+ULfHldr+97ProBS216paC5npBpxQfNmhKshfAGxGy05VW83F
4I7y6td8lL93Y55dxLMEUDgttqymzJsc/8glqsJVux5gC2vY+uxQi4KeHnqNq+UzauIc///N31hW
sD/qWitd3I34s1P+t3/egXaCbxHBr+KeBahc/wyUS7bfNz7FB0CQlpR4rO7pS+/sh2PaImeihWLo
bX/pQQUEAPVsFhrn+J3kqzIZZ4DEPY25g5JmhRVnJstFnFpz5SwtZ2dy0TTUgjxU4EKJuoyJhW1j
xv9soJvZQ3ZcZFmaKUnK40DA1bPxA0EYkTNoOj7dQQKWAc5JGNMoPmZJEJS1YDf+TZ+2HOCwOiZ9
MJB6fnh9E6WoU1K1KYkFy22WvIe2Xh6ricsTPxWGWURv0euubJ/pVIYCpNFTYsNYX5IXL2fqR9Pr
zra9/W25VY5KM1sijNMeGwGrdDuiq4e9C8ucCzgYBCJ5nSCkrB9l50mJRuJb8RFZ/vaTeGSYeLDC
+fCW99FdwjL3OhFYaCOQQPevySA36O3wvN7c14ijlHkWzm4a8OEAbTrzIg3oUDtKzq2edduN5/5P
lXj1B0jCcGP0B460wRv0JmPXTg1Vb2hoEw46SK24s/prKmrCDctxiH2vlgiRkIKE6rvwO3LFqep9
qqnN9INWS5EG2qhbR18F2YP59tuhPQBJsATRpF8vpGRk3fMWHAQQFeTdELTa+72vRDoRN1Q+dCTw
r69aYXm9fx83rGpSQfoU2lvqaImqneF6X+LV6Px1kPS0w9oC4W9Way9RdTfPAD1mEfCFckfjxciv
yu6b1Ia9g6ew0kqUeb+IiVUy1EbstSP1Hu8qBE2WmqL6/plhsB/9VOI5azBwIaMCgw37slr7bvAg
l0Ts+kVUNQxu9XIkZRRRtblKQM//0TIIL4LlJNxaouz1iibz1qjW68rNIUzqK3stLLmXZzIakXaP
zy/dpgICnFfdslS5Ug5tFatWVSajkIiErM9xW7lc5bZdKyPBh+bPCtegwx5l9eZQnH4B0TtBmB/I
VCy8DPUq/+CKO+9znZL8DI8jO2HzUKq+eBL/x0xNu4Zy8LAlGgWZu+6t1ysEqsInas3aIx+bU26Y
9s96t+na0votjR9IYFe3N7DgcuIfZXIw6WDPHZtikeuogeJrToFH+GWCMdQjyRh2lnOO/Us1yFYr
HiAWrklIDQT16saKcmlfwsooAcSN04TvoDr0kP6lP3zfIqCldN/V4C0F+yix3bDbhD1NKHht1QSa
1PRCSnV59JfgEsQv/pR3GQzJ2dOzGQIG0erGJebyBca4z6wD+FytOtifzk412mkGA8tOVvAFby4p
lzf+qgUwFogHpj21air5ZDu2KNipPljTmf/6SjhtHICZz9onXJHBOANVHAXJZ+xdRG/fCSsdGXJl
9lQTfBMfklAiqFNbkMZKgJ2lJGj8m6zE4tvbY4ZU9p9kEyhKymVc2fi+yA9N2htZf3S2Piiq43FP
1VKpsjaFLoqrT/N0nJbZsHreQrz2vqe3DYWRFu5W4dmvx8LatGQPzHR26zNIvcoF3AyHauLsQFaQ
TEN04alYdEHQo32txL/pCYsbF9jiwL/wupYRqxu8zl+XG3cOuCIYn3QZg0TlL8YMNZclDjRFLuxu
65k0/gJvwQaPTdrm+owh609C88f7urF8gIo6iJNimfNeQJPGEqRA21wANHKJCVQX0/gOcEBBtwBm
wjQNvJVP8quV7seAKwAhLF71idyk9SfnlaaEt+TPwTn7MUMCaHlNxSXofx6Zr1hYq2nbOXuPpIu0
wDq/aUkAocHdhnJ/kRXNvewmy/IfFyDsV+EisKOW9VEwGr87z8vfbahYGlC8ahl4oqy6UX0/pDVn
aUS1BCUtuqYNhnQ4Mv4nxWXnaGW1d511at3zie6190ZFxpTkEakyE2WDSF3W/ifddbSZaFTIcftf
/tHE0vmhAlT2bmxqINTlylg6TmK+//HfL7b1PPQLRoBdYQOV6JONl6xxm7z6XpzxoF0kQPgVPslS
WQKckW5KP0OU+gMBaFBounHq55fezVxG3+aJP+giMkpAgrGRGne+mWDOmaIkuOzdEf7iJBhqU+2I
tpgZN55cMJxBKJ4c0k7QDzeCGVTu66CNbLZjg+q73lqFEwgSC5LQsWVvTRFoqBmrXn3ElpWSVzzx
lhSrDK1LLdrPX/19YH81tpM5xpLf3KsNAOZaP9geAlye62KoiWU0q2IkyVEiIgKshGtB1Lji2fSy
K+6ksk1Hb1xT3FzH63xjD+vCE3s5JsscMeH7Dg96zUEnNRBCRWCkDkw8aLwLktVE9KLY6gkDd7Xx
BGLKtFDO2dEjnPtMEwNUabjMwug5SmrYERo0pxtMrcqlbENYcw9swWD2N1emomIKaojEtkndAevx
v0st8PsLg2dXRj0H1cb1kcOvoe9kJGi04Kl5cUQFko0aQ9H7qMPvR4UWkeQ/Ii4WXITZkpnHTcNx
VIXvmZheGdUl4Mj8e1YCjNf4D6f/hJQEnOF9o3BvlaASS9agWN9kZFVxH/5y3poF0q91MUA/igX+
asruk8ZK0ezn0J7DzS3mgREzQwrIz3Yr9b4pP/VhczAieF43LQd85zCKtCIBFTcWkz0kYAFoa0s+
q9JApLAPr8hFgNCPvBWhwIDGfNTi2ma+E9h7b6lkhvGk3zvHV79Uvlx3rvfv5CzzBBmPHhiF6gLa
XUB1yfjMiPC4iCNCwvC7i7PfWTs0bu9vRhlsbJqUIEn+BMijGdq6Y7zvVv/943Q5h8TBpK3dvScl
QtG4TJ3a9eUALUonRaKFuRl/qBooFyS1ZCjb1MZ2MWu6lMEi0ublW5JqDdHB+YC1Ysxis7yiFGwf
S/ZQ65OqskF40XVCyiW4oy8ziBR/s4EH/7Gj0soCKak5RJJTHWOJ4gZJkEk7FFdCZdBOQLsnqNAK
g/3MKYVQmWmabdD6Bp5T+yWLTWOj2OP4zfD8eLGWH/s1+BBlZNBUEd1oq+CnAhokxXHxLkqbEAU2
SBXRvmBi4tfHu6H7MZVvTBzX/5d58Q/FuaK1KeGw8fxsopQDswQ8ANe9C1LUY+a0bO931ByzcdmK
q2J9vKS4R0ovK1QPeUQ3zGrd8JVCUPHL5d3VzOl2E5YX8/6Nc/qXk1HrJZcTpArR/lvce9SDuXYR
/9mkU4fb8u5/6udVVO6RXOaz/qr0Ccz/t4b6GLtHLjgEeCJ/yPjx6ZoThGA26nGqsFq0MMZTvPwG
tcta8g3QZUTGulp9y4vnUZuaXaqEZKN36v2gEt9fQH27A/zaN5UwA0EymfQZgyNz5c6NK9ZDZhYq
3Z9FqU4qY089T82HZxbXSWm/5l1gFTGLEzVOlEGNoSNuX6BmG9HNuMBANNVXurk1OibhJ9yUSAdL
a+mZ4J8aXbSI2hBS4C87qczxuYzMrirTsLg0bJAD2bVhfuNgaQjaZ/9ZYrW+XwFcWai726CFM0Za
qMGXe28wHEJTnhP/P2MO75llfRAsGDysUYmSRhqZTMvNtsHlzVNP57ZV/0b1e+aFUsZNDtIZAKuN
VOtG+26Nolh8GvKkRTEf3p4AFxmX7lz9Oqd3ZOLklIolGvCrEdnrDunQU7z+h6RkiDAbwl3/J0gj
ncrx4MnoPocVJlDBx+qlrlr28gphdkDGMmNkSngmXYXsuyLqnAfvzCkFClOWd6mxAu4LsEAjErIh
3yR0paWjXA26zK7nZR5ObbcIbZ3mf7HqLVZtysqdl1q9DAmsR0mzDjrrXpU0u7jMViTbdIipY9ZE
pXxnp6JKlNfE96pUYVS6bGMReIRtluopEkfVncWMccPA1IKEX+aWv37MRkadavvWCEZ6gXx+CV23
e6vnLjefV1Od2bEqYuKm7/KRKpGPnhrjD/qol1umDyPGASSXrh5jtzU6qFuTw7EfviyBLX2nWyZ0
E/n+0rP8GC/IZjnH+2TIYw0oQuOAil0Yzr19QHKn6AcU/datYpzM/UhjQDE6tzhfZuydO6di9/FZ
1T8X5VoRGMpDQuhjh+3ws6jvkYdK5iZuqnvhD4ucTplp27+qRFMlHTBEdN+ys2P4Q9LRUCtRFVpS
wNPM78nXYM+yJTVLj1fouOxfl52NSPYHnvT4RU8N9eqZhR35bu1gsqy93XdR+M/WpyDWgY7HL9tl
H9JkI+5NFdgAdalsPsQQuDD144lRoht8e5T4NMLBzQlv7biGdZoddezZxXq7DgNmwpCmbplQcJuW
GL/hnio7Lp5ICAPbZEEBw26jwpSs/fYg201uUrFHML8pbH0iQdbL4QjRSl813sWw4CKwdexsndUF
tyuqzkO5f7pxw/WSvF0yWy5E+XyzqlIyP48SSCGg3NU+9pnnARtJubbR4/MCX4H7X5AszQzSqX5A
s29HumCkZ68U4hTQAzE/7NW0//KZuwCA8s8+oukbDxbwFB1SRPpX4781JwhH6YZlWXx4DBzczk9W
wbNlvyBA2b4yBNpSX+IVjmDA7CsY2dGtCIAyF4pznXIlu00FoS5neeeVoBR56imBeHtcuHkGq0X8
sDTsHxIzeyQQv7l43qWoAgaieMxlEoYmXbZCthTCMvrmckqr5+RzZ8VzaxGGB86wGstD0MAIFWWa
D1hBn9OANwGKMHufdGRCcZ/GO1+uVXlFSDspdy2JHpTS7edWINKwogvkjOARtioOd05EH6FDf8wD
M62eXOwRiWdGZo5c9xbjUCcrfgOgUKF+NUDeV1jW0RrYzVpu9U056hh7dmIg+6ekH3/MAkIA/gjC
hsoVl9rjkxQI5/S+B2c1h3oU8L4VHzGrmOl4QMKGp/QiIqgl4GKDLm9IvgEyp2IGf5vBOBK4amjV
7h2wKQX5VpGyvOeu9XeJwxG5KeYNviRsAepu3bQd2014gDI09KEHuxFsv72UtbtRmylyj7Szl67q
ZtXBwCL0em8UOxzz/zGV3OXfLg1k3NVC6Xh9BHeEi8Fd2Mo3xaEWPCGcghnFgq1+kOLTks7Wg9ob
g9nl4R3JvyMZo6on5Mh6AZI2Ad/IZPbBFVK+autuj528NKzy5BogyCMEMWDyL/CTPbT3iprYwVXq
RDXrF4Z5D3Uj3FJJRtRhT0uQ8WdQomuwllyWDqs5w/F/BIHb/X2YT0nfUAoK1/47xFhCqVrV+7tn
vX/UazvyybqeXNT9Yz49X3GYyB03m7N92q0Munc006VcdmhYbbdfum6T8+z7CA53jXo8orOqqlhB
eZ609jpM2P06uNDW3Qfqy4OW2IWpEfkrsTwnfUSVv033XTIW3CvnvesdRSpwU7W3DYcXpKvpU2jD
BAHoZOICy7zr9Zx6WS6R55uvwC1nmOmccb7vOgPuz1dxkfti0ZuqwRhjS9dWDsET+IO/e6bDrNU0
s2ydR6FbVZwFtvk4PAXd8KxNEnMse8bz/ERIk8n5jf4+H58k8hQQ1mUMwNMCYGV1/Cd+0zKZlSbQ
BB6+wPM/lOnGVIhiehlwM3ocFbWjhlCWoZ+1jb4MQlZie+95N2wLkLRCp9HwZY8YS6/ctAdIO+qX
tzfxpCk/K7pIPWDL0Sirej/kzDT+wwQoqH+m7dzKXz+TTGvFkUjwvYJSU2d6KCodIKJoQ7DXcfkL
V60NXqGk5cW/lNZJhH2ne/9aj/YF5FxYuXsg0Yit71cXeGYzdREWJ3KXEQSxeHk0APH1d7mV56bS
D486/XEhwL0hsnL+w+b5elicUYrxtnXH7+BPBv8w4es09zqLgmKj73v3lE29C/C8UVRp3FnXWvVa
BMk8W2bFvYL1+ubt9rFu37+T35hVQAAsSNVDhAfCNNBUJieqMNm10lObTMp5WtjdNNLwo+wGJAeK
O2tmVRDldTRfdnJXHr8cJhdCAMIP71BQy+g1qIFUgz09E60AJHWDkawAMllKsLm720djcAdRy/rt
hSX2yCjvamrcwCuLcYtv+iM7Q5AT+iAQqHP1DFj3BM0+mYWg05kQEtDv9I6UfpcVAJfVIxZ2D7nd
pL5SKwLmlF6BKEUCCxeaLh5LjsAx3usqsziBIS8R1g8Xb44erhqgKPohl+wUALcjK2yNQPOhvC92
BQ8dEeOL/+WaOxQbIsU+sUqsvzZnPotNxQDjk0sfLU4S21njYwFouiDHZ8+P4M96PqyC3F21wR1C
726g8zQv9dXUBb+IXjKTj/tdzRK2fjG5HaFuIFDh9gKIz/TQf37ykgXF5hre6kzuQNcdF/pvDD+z
m1LI/cqysMGjqexTIo6jHyNvPikpppAowoKjkFaKDNYvj93PMt92uJhzJV8aOJvmWsdbkAvJslaE
RQJayvnkUbyaeIprpuB/760jG4400MBQN3KChU1vJ9sEpzljAYV+bO8pyMw6QXyOQw8Uvqqw/IvT
2TT4QTeriTf9Pi8LwH+L3AkkGofnuZ4rlpyXAo1lgd9tZ620AbupWrzqjdr5WyP7JhWxFhZKlWaD
YeizP8VTHOEjkAY8TEdfbB+wg1OrMAszpL0KPaDm26mp0ECwQ13nCJtoWsB6FhZTLqz+AE+SEIjf
kSkW26xTNuQZDoY2swwM+c2PIvXHA79L5Bq7eKLZcvBtbOwIn2Vt1l8kV/3l2hVjAxd2r2q9Sp14
pEc//O/IHPMW/uEDMiBpfKiOSlDaM5qmdWuIq7inqIoiC14Vyj8l/o6MRQOI8AWGjyvOmHaF5uft
WJxDgbiqnoDL6hkbYE65jiQsFFtAdDNqRXxO/aL/poYcNbFuWtfKJsEc8dF+aMhJzL+WwH4sMkD1
F+5z2d7QQ+EvrvWpVyJa8rUrSWy+HNkL7BtrMZGiH8PjunfNGmtFw22YDLlo5pLehHoIpFB+zIgi
ayNrdrHxRUVM4dhGZhqEHkAgC0fXTydILQ3T+OM7VQMrAEi7Q0tSPfkiFCtDswwR4bLtTS5rseoX
DqsuAhLhkBa7y3Ef5gcpX5PEB2rhp/t60FOTmTeb6iiqHtu1S54Nzz/ZweoBojnXq1yIkDgj1wSw
UuPkUW0DqFTZr2MMMQy9PlCJiAI9BEHM1U7FERp7p2nuhPOJKt/w0Fet8tyi/bQhpAE/imCBj+hW
nwTD9tNPPqcvtQpw6hVOPebnnUrx//6CMngoPorkIObO40tbM8/pr2YCFmv7OvAAa0PKAuvBhs/f
VhUIaslxSXH2aeAin70v9AU8HC7GD3SqAJXdKf/A9HZdsBCps9atkO/6ZsXlfdtAO1xNcDWk9tVQ
vWhYaGdY1e3DbTnk8oR5UftFdfiiVh9z2C3keTFHSBtFfDU2P07UO9x1kfOpBSgHwfvvYltayHo8
fGr5jsTMnJ1/jqXQ/v8dNnK+b6kz+UXQ1MiwyFLC3KzkcQrnGYuajIuf+lTVTkgsrRuqZHI4OiKo
7OA4cJmeOsxqIN4FPHfcyGZd6TRYDqAcLaGtSRn7udkVmLDctudlT0dZ6TG0+Cr9jVCF5xmoSouX
chvQduLMEeBWeDc1FKhMWX0LxDuM4suNSrW5iUrv4PmuFsdrpuM2N5j/OP0aZB8ZrmjZvtJFvAgO
2lJyDZzCkWFrf2Id7ExR2Uqm3GuZeCZv5UhL41mS6iFC/UuIhiul+9oaZVzlUiFEWrfgiVALryBe
v5U07nlrESZCARCQ3bCiCmm7B1gDlwHwc+gbmGDRVZe1EFoi3zRC/aq69y3EXvP4NQTC00+38QGj
ifPFt5epG/8aVWhaGVLGk/XEXSm/H+Fv4+uhh3B5FfjjRReCz5GPooGI3SwHf2QRcNzN+BWyvIrc
kf0wE1PSDlauspibWTR9lmB5eE9rrirczWva4Pzz0UZ1FIEsfsf/6Hk7PSxNrcZWps76XHeegQUK
3pSdKJEqmcagTHesMXpSG0sdvYC4zUNCRLpT1NUAopWyn3tzPCeSW70Z6VHBwT72OJ6iUmhgDNp8
4oVE46A/rPm23lkBO4dypqQplKqwNF+eKPQR/jGE+SNDWvkJGr0wYsqvYly5yUpHHg5XCsuXmNS/
eT//zQK6Fa+cBo/kVVVUMpMP9lWYV8174QsQuazeV6nEgRkO46bEAKp5rpygTDnL2SYAwUr6Xyrw
q26SUS8BiE06xNwilkVsDL7MXOklI3Rvi0ddWSF7wGl/iWhudJjpnNyw8WnBixMKPT9PtTeggbgF
p++/UyYUiAOgXrlT3aPjKEtbCXWKsvphCDA6sXu5tF4BbN35eEPcqH+5NnlxfK9o5MIVegN3lkV0
+3t6vcEjWF5X7NEg0JR7v84xU5qNBSZyXApQP+znvaOW2VbEOfEEABJE48tTYxYM3bELQ5AKB06M
1vy3OWSsL9mVLG42at5ayevPh5GBcqpURg+AAFnfWN+E4+A/+s72RnVc80a3VfLMIX5JwLSSfiHK
w4W+gqHUz/2us0Fmi0YXX3LI4R8Y5NLLXGbweyO0ktAiltZzDiq/yaAMYi8lkDwUdfK7RCfKsvJN
nAv+OnQ/VoEKnkeOnbfI1mJFmDwKvVChIYytxjtPlDWVzIwoBMbZbiWoDV5Lq4mhRFulaca7VN6/
8FwfDPVWtqH7ZLstIaQbswCdvS1xpVRREjUYLuVkPY2fmnfQu1fwZ2i5r/8cbCAeYRqBJh5IWj08
OEe52E1zalpshOkP7TJNfMo017V6654ik++MxEwxEQkTYdk2fXw3l7eogy6n0EDUZ5lzpwWOWyja
eq5ekLV/lvSSZ6N7W9VJrfFNxl1E2o6RuhJ7istcmyc4ATX1eLQfyFnPO5TqKepanYM2OKmNczLq
ItFC0atH2CZkdl/+qLaTM0gpFE3VHK2mk5e2VX/IeDt9pAhFs0ct5YTSilNL8zSTLALgPR9Clo0a
ZC7kY2q0JSCnJCo0h9glt7An8otHrziPV/6KEVfvavGlnCc6PVcaFL3+EwAm3Bo57SpT+yl6i4vu
0dBFh7y56KHL0GRAVKkjY6W+EyaMkbyxOlOhdkqHWYBnhM5kqOi4Gn/pqF+zfz3tCVq5p6UzVlu5
caZS7kzRVFCay4JqdyFkb7wk8hF/3TZkaRpzgGHATD5qdasQ3+Ca5vZevLJ8r+Nwukq8SR8AP3za
W7mtzdr6NKDTiv+CAawx5/mSRrTlLwNBu45+xFiPPBKZFb4iVEPPMId0wiRpHxfyt1cQ3FpzPRHe
jifKAqkvRNFPNgbh34NdPf1PO0dep8ShqHwRzs1vpfR+lqm1TZQiLxLknkFGNDr/CI12KCNXWLyV
LeohtJfQ1gX5t7/K5wCpms4b+1mYAF5X3y50gmrtrp2zgpS6o42CvtB1R3dcgrdnDA2JrltdDdRU
IFKxQ+NDZmW8KsGFXee/ty1xbYZX8tVUrj5KfCbqIPasv0KMbZxhlrPEqpczF08qVBedvrIm07s2
mT0ePQFwp5G2A+UDXIFGJdD9vKhZ3Z5xpNSUoWxZlcit7CL6Wduv4ld7aiw0zHWnwqb/qHyWz4nc
jhuPmjBsGM/TlU1ZeB3lLJ11ctJlBlal0FiHDWT3dvhPUjgafR5qXAgwBL9tXw4P8idNtyYy4+6C
4PV6SbdovqIF2QQuvGM1IzpyRgVwzXWsMmRFWHnXqao4l5EBRV1qbRX3KDDLyvjrbKgyuXdNa0uj
B0YwRWegN58av+kEBbyOnKWwhO+tDYiATgOgyguInNJdwkiPzEIWP5kF910HpnfWvZLx1xgiEKQP
6hR0u4Ue3t0QQCal1l9GRv98wnCw19P3p+mrA/qSE0ysLW7jKZFsmfC9N2hNNdrY5MDbYJcoLvlz
3rigRZ2n6BQ4BeFIzXrUNH3tFQpdic/Ds4YTiIMUhCF4Bh8Xcj5KP9nAueYvTV8hr0jnzfEDsiQ0
1h6jqlo8xbY9RxFtr4hGUtrZ43goZ0d6qqwUx/fcagJw64RGiNTcdYFaRtjzo0fNsAhFKGjLTGJo
OYD+nk21uEC78Lio5J7DOvb3J0aI6hwcwKMAJDFeGnUrjXPZOLTWcewhp4bUStM6dCOPM3zp5oKR
4qpB9OiDCkiWvFuuz3+8dnCvui3eYKqZP7XXtoe0CT+fYzw00i5El6+2UyWfhiz0MrxUoa+ie4Jo
LDs6zCd/1F/cXH9lr+PFt/DOp0PAb30HaqL8/2wTjCw3KuBW+QmDA/XJfwQ5eDw5T8ty+Flnr28I
QKPni+WmtlWgvAYtkI2IweA2AytCLPDEUCjG+xsepycwhuWazgXjaEtGW6h87fabP/O0QtFN/2Gu
6GVn2z9B+O2ce9EtnuZL0leJIIC9YWYiaYh5cykaLwIISik6Nkuyip+XArlwPirBJcxt/z1qO7Qq
KoXjTFCl7CniwrP0MxLygCH7mlaSIlVNTQif/oR7bdp+/jcT0GTRTcf4wPTgwWsV3JH9n9ZIzt7C
prGY7r/rbWqErpXQ3utPMA8pbpiqvXg5AglmpCIF0Sy7ywcZA4jybXgwDlNGqp2Ykbv2FZ+X0mRy
U6UCbMZLlM+vSbNuK24sKJvU5ysfY/eXBiPt4jptp3s317UHyB5+CcuLcZmPZGm9fJa6u4HW+/4C
FHJwPZeZBF5+cE0guWYTQbPCF2WYOEayZwswSrwhesM70UQDvCrnsd0NIEGUfORE+84kbfxMClzq
dvNYFs6qqH9bGa8LZPGCfHQhFfqbTwMkgVjjCMLr7Z0CwXnfffBwcepy8lziNzLIy/MnovXuqZfb
5NF3NGrkhminI/rnmL9h7WuRa7qFq7lrfqxCn5E1edUoHbqLe+RpzgxHLOMCRn6Ta8lfM6wqKH9W
nqL57VGsvkduVpsmLc0feq0KiYGaPhYyREBzMd32vuvoP/MafrpSMpCq8/Ealptm7c1DUdxddzyA
PNx3UWXrJD2ACmNz+rMuOCMTMjugmqNsh8b2ef9ZPsxWMMHvY5ldRbAT7+b51opEKSII4HpNR3id
plI/cFHE7ZhvqEUvZSbSt8z2RmAp/cg87LkJc3FySBDCpkeznuQ/Adb+tpLEWPw1IasFSV8IeMx2
eadDNXn4XzUSJmMpGvpkN4ZdXx7WRdzy+bnWRrdCAYCVAATpLKyC5ZFV6KkExWlPh1RDs/d2zteW
0jdkXNd/yjJuSmMMZPNDeT979qOUl4APtj7UCNrXV+nnpE+PicqMgx6w9qzELE4dehu0EXRoELif
3KxqJdJEUhR/Ku+VT7Q9vRTs2rp2e9lqY5AXJyg2pui8kAxOfbEdMmM4B5MvVvcsTxLfRioS8iui
i//Yp5YGQT7gCu6JGF82jTvxIltjyDAbmC8PllBfEIKEyCUpvLF/Q93XtOV04XYjHVchguEr8DYa
PK0xLnC+8pTs/YBaHzXHC0EpDHNoMgQ/mQ6VFZEaZYQFZKmII23nqEI5E8DT3otGpv9wfBy73Yy7
CGwDF70KEMn2b90QiA1qytl3rzre9VR8cclH6nW08ZhqygtPzvD1NTl8fR7h+/n467NNn4PT9oWc
VcIik8iiNvDLulo7ISTGF2l/eTkFmpgPmfJZmfEeK4+LYdIQC82bPilfOVEHgg8I7XDxin2cH6fS
MQhfc0n6rmoDYzHuJb3OI85Kyv3xadMXNuwkl5rCQ2zZWv1Rqiw9X1dxfBcL7C6YrC74fnnpBuaj
wiDTiQ9+lyiXwZbxUPJOav5q6sgPTH+B2oDxRXr0rsFpfoaOPgb84X+QZY/q+8gFq5LACtE2zeke
TH0/Zc39kefM8rOGpUb3ADH0HCDja2ooa92HeKVCRG2qtCVU3a09MlUO8lomAJGHqteKRO+wh+lo
ehfchToC4+azhZOjHi/BQ1vQ6n2eHYk/HYSq7GnjkvysKG1/Wt/3M69SQoKDe+Yk9AesD22+RHJV
9uDwcssODcVo+OBOU8TsM5K9lHwt3qBm9iXExancXiGW5mh0plO/dmkWJCEEaRsAmwWX7O+cJ5xR
WzJbxARUh/Ril4qYf/3zl+SgQAx4W7sEXYiiroBp5MQrjGiyWKNpmQzp4jTN/cy+L1mVukjNrcSP
lUQdm3pHwMFFJyYeir9tTO85y/Valbth/BOoc+oQ31AVYxIPSrFTJ05w1o4KdtI9ajOwcgGOJoXO
Rdlmt4q/1lRyIW4PdelN0qme8TjmfA7Vcj0pDvBIw4XS8hALmrNECnazkeep1pZnrfRJhZyhRA47
KEkrGkUt2N+8l4ia3sj4ha3FSRFM3AhHvVjQcsqDseTtvJoCXqKacD6ZFXILgf44xqMEaar3Fh9C
9ieeIveZ1O3V3neQdttRCayDIvyEqgCXGNnuCEUHEADbXGw+RNLwc7gJfnK6xiqOU7l/OfqU0ft7
BhuzkJ5kJ+GyyaSpuB2w0kqJAdsL+mcd0I1nCw3jD8Zs1j2RIxBi2JKLGkR+B+5rRi4E1mqKRTu8
IJ1F6t8K8dsY1OWTI/UoC5T3s25hAnPwXSO1syzyj6Fp8RWgFDmreIwtgufNRVXJMwjWIx9Uk9ce
Cf3wO3jfbCHTGh2IAdp11jWaO2e2TBoDAOf2v8oTu9M/t23Pg+/pqpJFy/pUl1t1BjT7XBM3Y4vy
t0JRymzAdGLoF3l3j7SqdLvaiL+T5by0KCawNBP8nczfh4E+NbIqe467jd3JLK/AT7TlXoERmHRB
nS1rBZYSoVtAzOJKbf9KHns8srNqWX+7I/xkboipxnEyPWnrbAO8owNyvvQ0pZotoprZ/nBhu9mj
sv8sjii0TtuwIyPqjHwPLMZCNR6L9Ljnlpk4Y1eowQ7lmPhKfqvYRGbBYfCc5NJ5lrQS8YcWww7h
V1Nts/oUYtRwtxGzXTnVSfzDPLVxL0ZQAknLV0GTLcl3uDlR1Il7noSXWrWDZvKW6DBlD62BXoCW
/ZfhQuzgzsTvqeMNxJumOtz0rWIkR1pamF75P2n0PY60G0lvkun4tPry3dqyKJcGmwYwnl06JMwo
IuNoqEThgjrwIYK6L0dQebkFd08X2FHpzHR7fibAk6kfr+T+2NruXqkfLpqUmlUbMpEx5LG3TIjm
A6TiJ9VzWWEcPLeZ3JqCDiUXS9tPSO6RstnYRPTpZph/Gj55DUiHUZUkMDGvWzLrB8V0fXsu4ghU
udccMviPRkXMoVTZFOs7QO7iKcjlxWxcLv6UVp9maE3vZHp8VVyYiv0qGjQRSE/lQSJWHXBQN1A3
WiiI63dpPHbosctJWDZwb0dsTcCaMewWSOCP81z6lZVFL5jx6n0GaSV0wpaIricRCEZk4MNXL28w
U837U4YTWzBAKhVjbqSafB7eKCgUpo08XmiAM1LlC3THr9k2l9pYAr8+FraV6H/127ls/od/xrjS
aah+cLiPqcC6pI1lypPaaYObTTyJQAf79fFrS4EMCc/MfQ5HOj/azAgKZO2OY/Fp1tG8oOwEw5sG
tsLdu1esYxt/oawYr0V0RKE+MKslNlMl83h5QYvc4PJ7o9sXkKxTmnA8Ahg82qYMpNNR/NXGaLH2
8jEZ8JZN3uyHSIck4eUAL9nC07HbGjSB4gjrgp2MshvGctH+gaT8oNnnNn5sslXVN8BJFxRBAMEQ
L8gviS/xkVY8n3Q5yKf6xPNxCsNd0/cRLzwjRDHN1Qy1XSczt8SE9jWh50fFKgaGari7cthK5fIs
ma7fxPOgEs+B+yecrGB6xgl7LgVnSMCvqWt8qf/15UqJSdeskjf6vGTzhQd1JmKJ/FObeaIczeSJ
fNgab+022iiYBHKj0CwiwaVfQnl6KNY/wKDcgTid9dTGbdgRhJSvjzV/eTd+W8ODyh5uFRKXNy8T
d4uxXPOf1WXVD9+bM4NmvYnsJIKDO2qXIymbW003Blt8aTEykpZx7EaOhUVzLk/Yc6sF6F88nkXc
N36Azp0bn/qMVTzTXhN6016LdsK7qn4SfPqjlTayDM3TUtonA2I1SsF6QgZeLV677F7oaF4/SHC0
HesqDMZ4VK1a4GZesUnCm1Q4OoA4qPYORvjm6ZfwM2tz424r8pQatfI5EHkIEmk3AuBZCsPH6tCf
P9kNHHNeULRANCu4Xu8ly/q6rVCi9bXxAtekzw5VblPkb5b4tpBtzf0LlF2eaeG4/Hh9P1modg2u
/uoXtTyVUujmF6YlLRJmZMUmpd/ciGnorqk0UydqrndLm94QxGeUI9aTnpNvn0DWL4/Ktqdhq+Ui
j9+9C122yU7odnk5ELBCJny7N70Z2txANawzcr8tsyBUGX5TSrFcYSzGRGIma+RckxFdg+Iw7fqS
kBBqcapxcjG2QO3aZZ4zB5VmB96PZ9C1/dKL6nRILyMsj3Y0uVlcwFbdEbyLSB9qdQlLycEi82eW
n1yT/1oRoBQkKf1Nb5KKZMbyv6G5G6TYtoPHvSWDkmKz4XPFIYWZdyPTE7I/DCbmTVhcuFJAlGbz
v93wPXe2SkxDPxQCc+96X0psnPE9ryd4JfMEBBmTUJPlxwnKvO0+9TSwRQKuBEQC9qfVLe9GNqvT
CpN39LzKRL7UIHWJ3cBdkahofbl+0lGZYpp/S426DJtfKDJBqqQbqky0+Dl0M7NaBtmMBGuFNEMC
z0qGjpOZyC28gxTl14w/rbe88IcPTW4YCMHIO/2ce98yFlz6WyYrWVr9RGkgaDno0unwghuLbJG3
2QZQS4axAPRa84MK07ZVhzfnacvnwp0YEdO9HakCHcq74usqC0uL2WKVP101xCjLa3wfvIuqFwbm
JfbkmU+l9XKDoUGT9QAjdEPte9ITbl6gNfgv7/6sC6mOG5iHTKLGsZvDWu+Gfl+1dttc//7oe9Ut
SMT4Vb3gv0XCZjXAo46J1i7NVNsGvRCsOgBS/YJ4HS9ZO/leMaueSKxmRfTwPYO0TvhGvc/dQcre
VCeSk03S8Y9twV3siK2IXKU7ROpDXmFiUDnr9sRypapFNiT3+3U//LpPRjjKvo+jEUjHfFJMhwgD
tLIfCYyPWgceRegtCMXKXwkJAC/vjYMWCVzQWzm+K55+Mopb0CKvFwaazijlt+WXE0GUG2DQ/xlf
a2vGKHgsCOMB6NhP6FgoX6aI4TpjSq0RyoCypocTCzU6FmIEyyWAGNsXLcpIbebKT0NMPzhJ/VrX
z+7G8J7ci9IMnP+6uZzIzRpuYhfUrRFFz7fiibx0NIMhhp7NeGAVt+xgGEd1khXrXtTWpDFiV0nS
3XryeZT0c8Hqex40a9BL6VsgV66KZocSbAEWkg5KJv0zhAxFsM0pDesBjjLIykLUZZiqMh2JKkwZ
pLgaOn45XETx1m1A4xziVTYd/6ObJFuG0WaYlQcOUVL/+kUHhDtJpsSD5+4qjw4Lma0GRnJP0Pc/
TXSBH6CLPB/UtGFJ9JB/rsdT+6MCh77hUfq32Cc9Zp/EbCDF2Xrb6ffTCbNC3SAbrw1z42xiV9g6
h0Ujojg7Ywm3aU/3McYYdue8rM/iPj+iJtwh3pjLwmOfW94i3hbZGdsxO1igg36u7ybT4zVo/alJ
2lFSMLqvFwqHC7PyS+HNWDJqieLGY8jeymzTYZp3cKPcdW+EOHGwymzv2zW982YIxdXksRzDsUuK
5mekrZFgZlBQa+0Ytpl0CGL2jQNSIqL3smjM803CCr3LhXMFIw8VyJ/PtccpPFXW4hZ8gh5wlz2Q
PxKsReE5qKHWa6gNdOOMLOo4E1ACFJpwhUXaSF3gIRPc/LBmeokpu9AqljbdSaF7B588IEcaxabW
6lWmvkp7mR2ydeUeB6vzkYmtdqhKTU5fejeNF2Un9v4eZVwCnXZ92UNvtYACX0cUUGlVmnPFyLCJ
77VqgszDg8EtDytfUBMD/TcgT+pHflF3L7P4kIUcHXy2Bbxn0MJhUzFwtW5NaDC7YqMzH7gWsf3x
xzI2yOQcViNpZxa0WbsGAZUQD+UaPNwh3sNWDZYsq8LPkgYJi9hvesmnsinqrDB4tc9g7fqrGccw
DFWU4y4EJC43UxPMvLSFCOOvqiI5fqk+gP0tkL8TopN/wfueDtWVohkDHPPFerSu7sH33XvfugWM
wk7vxV3zmGD4iJm0eK51yRMRnkm4IGl2PdmfvRKduqUNVxhIBfaynPWRVlSbb07nu1TAHGQCUi4V
m4Royy6YJClHZ9LjE5+E0r8kTEDiLQeHWhyvAoBuD26eahXgjMvPzCX5ZsBZwGkUCcXUMqQnPr63
EArq7uNOgWMEn+yAQjK9+15OFInfcq/fo1Ix7GqyG4UvCAQI6lRc+k6RODvgkQYJqsdvwKEdLJEl
GGOFVkrDNwuj61OjT7YTKZjOUnq+/qrkPkyuirrmxZsdLoKUgL5AHQtJLFgP3w2ixXuMKtDIVJAm
L2m0b96rXIG0FDiucx2KXppZ84EVzYfKjt2Xf4fCMJGiLzlrHe1F77qmoQ4vmFNAvB7CI5k8QQNV
jeJ+WDuRgUMDWK9zFub+ZVKxdw/hTk/WTSE5YDrdAn/eWdh9zPhAowTJCPllbBxMK5C9yE/+GzVG
0amtRTINyGuzAxHjpO4yPQ32vlRmdS4z54Bxt/cFXF4AlVok7ublMSzSUpNbv2ZXZSNq1DACzUGC
ePzhnAIICiEE5XXix1qcUcFWXrDHafUzNqF9HHlP9l03cyHJPZLeejEDFQK8/MyawDvfs4y2Jdze
TEykj2WmQ8/KBPfx/tDd91hcx7xTWrBeXfGK6P0y7tP61Z1KnSSOSmPRnDnmQgnn1ug074RymmSU
1i3N0vzuLk4XOJmmfJUuLkjeEFS4NogskX9IA7MdcP5vligQ6QlJfn0QDZ1mHOnDpn2TBWr9lisz
n+oN+aZbFvmKl8ToVMKQCKYMmOqeeKUqwIqSZAB9mIWZrjPd73S6YaPJFa6mfWy6t09NGHBm2a/4
b/gCWol7jpi0x4/LFVHRSd+h89++AEDBjUfjzZBh9XXvWGxlY/JCc4erXXESSC0F74Rmi/YxvkJP
e55wfNDcsgOUcByLoLOjviFyWVX1z/tHPpCxG8DE+3uysf5SOfTSv+u1ltxL9umkp2SU2yFdRAoP
tS5cLdaZv7qF2SuwQoK84HGiTe0Wt63nV5N1zucphdIMhY4xG1jmryplMfOUpcSklQ5pJkkdzH9K
e3uyZEXsf914P0yFEgO3KZRfrlv19OCaS17SHXejew0e9L5jUBVUCK8ioNXyhVUNElgW77XM6a9l
/Tiic6bYuH4Pbt9fTz6DP58MAJj3O2UsY1lo8bgrz1Spb/LGb//Yxsh/05ElMp/rV74YbO8CSmr4
epPMxRwiwiwWoW2TwsU0OzNTm4k6UCwtOFP5RtcIJcsu+6hBUoGLgNxxiSSkcWj2T7Ijc21xFsIu
7HqfQW3WgFw0r3N/U5jo+AbqfW8eIvXwAN2EUc0bcxhoW+f2Q+bVOvksJI6MpIHX9YJbRJXsDThB
VIURCJHv/YEk0QQ0cMANmEb4hbPOPQeqxzb9SF0Z95X5zZvHrNYeGf+ZYinYYbRvXRIuBsg6nUQz
7MFvb875zzMaVwmlXeCJgEQV/22/poshL98PSUhQ7OqxgBfkq1yi4YOimXvCk5Ybm4BoADxrEXag
M4CXyJMU/DdtD4zU+NKTDCJcYdNUs04yPZ9a6iqFkNHsKGefFqBW3dUq40vBhQiQUaiYabqOAjpx
OfuVh1IYyBZNsEBhLP5Nh5bUOHdEEpTPXx+oMZrvgmMMxYgNzrRc9Gely4YmxrZ+2Q/MsR7Y2Al2
Ez4mO7L19iLwUH9U9AMaXajZ/S0qNa6lbmMmIDTv72fws4YYDCybJjOkAajcN9CHb9+FYG/S1iuC
XFC0M6DR0yBR87pvQyvFgeZ5hssiPcGk6SmwUVMSsySbGeTKieVj7u6OFW2sy6JZBwq7pFp7w2gy
jhPYERLJxHOTQ3Eg4IQ0rjVdkyhMfSptRYhXg/S6Ztsde6mWcNPk1XmB2rjghis/UzYzM6abf/7s
sXrUkxsCalhn9hNjOSGmsEXx8cZ86XhOZOZsuLdwTw58WVKfR05zsKLG9aC7CucoQyPkbeVed7WQ
6+kVjq0Sn25o8ucNn2GrfYTYoB/y8g1js3/5GteRyZA8WJr93tvgJz+m94KwFs55VnylgTjVUoxP
SpeYk5XXHJmhNn3wcSYWLWwZJWcM3oZxts8yvqOxzxmFtQUn83v25BjTKzASifOIx+er1EZaJeEq
PJnoRWGOlv4HD5E1fA7sjNhZQpIvAfcuOwGF7EcCx+hKOaH/BBV8yijPW5dpkgD/4jsCe3qt0UFU
MGaX6T1RLPIrEpPHY/YfelWvzao9db/5WULUri24M4BIkSGFy4taX/xSTSPjyPoNOFgeaWf5myz0
d1Mcjciqe5WFeF6i+d5scuY9DHlEdCwtnUhNkgXpe4/ogNpH/NTe73Etyn6ZnoUvB97oNWl8r+Bs
ha/Lnhg4qU5MyApN1mOM5WqmKVD1X20JEuS9r6AbMxpFAs5Dx3DI/O/bDhETix3f1F5PLlDUsAcH
maLggGb30/6L+P+RiOko7Q0zhcqK9Rs3rVWMiCihg61nyvkblv1xEvy+gziUumw2pLyHML6NIlSb
eM/0d+HxzQgqTJiEu7uahdh2O7KOPijUTBojPqT97Xh3rJShXFTGsW85fmON3WJQ+Je+gYP2OKF/
yXep0B2gtfMEGluj11FmQNAQLF5ZUneF9NhWOU3NGnAqmw6XKSZSNUC2jvoEt71ty6Rgi/EO7+to
P0z2wunc0RnmdeO7HycksN8eLu+ZHf2qP5D7CQReZ+0fgqxWLv2RyGrbTbUXDXR3TSP+keIvZE0u
T9kZC9rdAbssRTTC4wNr5CL1/CwUY3WH+OYH1FTLgZZts00D/izWepwnL5PFE7j0vH+OIAN+Ttlr
8GqOK1RccYlFs9WoXsHtzpRw9T/SFfJLkToGVyE3i8w1wT5z/z3KeS425oPqjR3bmSQksJrQD1hF
oPZeZOKO18Vp0ZVCYfBMlZtdoUKOQqrTVAG0OFU3bD2Va0pW0y4kQ2f49ljUESJ2iV9XBkB7x9WP
DhN5K4Dp5I6UaAcI+jxdLtFImVEchaN13C2FQCwbBL8XUgDUrbEFAiCdF0BOhk8A11NR8V+SfeP3
z7AeALQ2He9BI0a/oS8Ayoz4JFIxxYImANjNJO2clg7RRZ02pTxzRdgrj6ZS2QZ5z5996DPRPrxa
e9GOUXpUbyiXWgIeOOe6AOmZll14DndndcJ65vcHKH/V8QDTs3KqXgu7LpAg9PrTGAhRRXlAiMNr
yp9lxnF3TQtsrcw1gDq0YvI5XqUYfT/CrdI/UnNxXzlSofdmF97MfGRSiDyUI+REgKbxLie0LSIk
YxeAShOPD1VJAlBVYaP0jGfN9o770ct7/wWqZXb+cGEY4YBch+UPNEnR56w8ZgyhaopFizc5XuVQ
EIJYF18zfv6ki1TZ2PdR83d61MDt5Rg5xZnZcG76+ZiOcDXjXDVREwjuAg8Z4nW40idvcnljrwVY
bJI4CwxruKx+y4upBStEteouim2KSmQb/zmWHBtZkMlGUNTz12zTJ8ZR8Gh9n9iD5KSHwaK+6PXA
r7Wt7EZHyPo8uyATQSM5KyKnbBrMtQ4lprJ7kzMS0URjA1upV73Y1fTC+cN0VQlEnsMX9BlElof8
7zGyF8Lu+of6/vmIpdb6SnopvgSZdDq/ZJecID91Dun35RmgBu4HyQbXuzh277kyR239mQu5zGmX
nJDnGqFQZMVtEHjPsrIFVGlWOz4Llxgyy9yWqA4tH03qnszrPgzWp4SaW2G6zQeKSOef1ebAVFxJ
4NzMiRS2vpy8e+CnKmP9Ol//5qgTUKxeRo/DrxUquQimK4XCaPtN0K0Rdop53zyIlEoGd5vuoN2S
C8d6I4XYAopNK8njVHQOdyO8kUxufoSrpUi8OG1lj6mqOPSXR29Bz8tD8yGe/cV5GC/i/UntbaVa
tMJn7qOjZW3MXIXlIHjnytz6k7+LO8oY6BdcW8IiiMyy+RdLSB+QcMhV6N3PxMiQQxDfNFZXiIzt
NwBrod+o1deZtEClurbfPRhLUwzbmJB7y1K0sMXe5yWwtIgYabrQTJbkTT6+a+CEEyVBbbhuFpdU
MX8kGB+v0c4kLhHIKuPVIuxozY9ukUG8hAFo6AzK20gP+uoAZOJ7CI0G/UZdfwkRbnOHknHQ41vc
Ah3uT8lMvr6X3F7bQ3QRo9b3ppdhODoJFaGFCLElqmDTcJhaZBt2Oet4pDBkQOObhtFxDENt5kUu
1INtwrzJXtvzjuutUwct3fsPmMGJGoUXVOrfDZ7K71EvpeN5ahjNlTrlNCGzNPtC5HdiawRMUlt3
gtu9CREYRDGVrQSUZGx+yy4uFVx+WrdkivnKQA09YgrFkg4CTFxwBbyhAqQ3sCHgGqWygP1D3NAZ
5ZoEiGde9IAv+KHhqqEhcxgSFrhvl/ZTREDm/RLLSM7V0kcqZb4tLs8VGhv6Chskn3A0jAU164lU
r1umkW0j7SB2TqvrvKlvIqPQ9/JBS4FPfHYq8cNp993KcL6fzbcV8UM6oeQWecDI21ooKipu92cX
IBhp0GzvFGuHp1oBamN6lQtrMUTo3o4RgDThyOylDtVTCC0jbE1oR8jw/vfWTAUcdtFeSSMMnxBZ
TxBC7cyr60RoolSbs7Tlvd/HDYwVQ518auOCQsET8QiLGaEOcklcIYUAc1uymSodt+IjsjzbbBE2
Ey/2cwSATIADvYJWaGZXI7fCvdhGl+J3DYw2bQP/zHPuBkp/RUy+4afqqyBN28c9ZmeW9jLyCIcM
Qp/4h4QaPZ0KtfAj0UnBxS8yPga1WVwbMZVkyAMOsuaUG3zM1+/2dKtbXOewQ6K5jARtC6HJKhjy
TpL+NfLsfcg6vONr7haR6jB92R3RzBVCzMU59nHRh8GRivZ70i43DH0gTmvfEdVDJYZBOdgn/xAt
63n6iNJaoOy4Zx0kjuFs26WypN3vyyKkBYbLAHJEQoXXYyBrM2THWnkjECSqCOEVWFu/fEwEfQIJ
i/pBbITn1g2xDoAfabTc4B3Y15eshkLO1xNsSzU6AMBpZUryu4V0xTcagzBBO82tpSwUOzs5GpMa
EIqNURSzvv5zZOygZ3NioQ/1Rozivl4KHmp70E2YoC3iTsFCx3OCMeTQEqwzNGWVZi/vntwLhWdF
Vp2KXepo1Vf0WgSwxL/8i5rA77w/FyP8/BqNF3DjNDjU3RVQggdQcSFm5bjtD7rNjmLPPR+FJLEq
Zkx+/sSyRUq5HTKzWkgRgXPjfXd+tQp6g91oU1EKIcrPLU8lfMjRfdL4tSCcq5E1mvmRA0L9MZWl
IeAdQa0t7nAAHFYTlV77Bb7/u2tU5raJZKnrDOCxbMLtgR6pnnN/V0WJi3qCiP7OJOXe5GaHrt15
zH2RFKc1wa1bF4S1Aj7IuMVeq6R+v5WbXoUNRHSn0cZajdbp5aApAGyPYCxK8sy8fHg1CYstTBpc
vQV8WVSdGkSl0s/3LPCGHwKsuehGzQK+v0cU55rehDqi2zJ1PCpT1GqWgzHr+4CNejQFva/lDj6l
UHmN3ntceAKOMY1KJmJCfxDV5kbzwpYdlC1pqGk3w+D8EOTpkF20qts4wVAZr7/wbJO+ForQkyCt
Hxrmu8ciu3P2KgQXnmfxQV0OlmlPmIeRi+aZTPQ8UZHJmX9lvd3yIJdnaA0oYt/+HAq6LvzOb+rW
o95Ej438+SkpsrnaDeWVuGTLtGMbm2REFIs2V4XBhFvWQahWvAqMMYfTIgwQKcqLC/rgZ799AQI3
vHgLKgGkRTb26R/45uSoLVqACLhj2BfWoSw0J8ig0FrzpIafyCw81xW25Sgpw2nP/A7t10vhT17T
GAzYLEcMVh/LtTL4lWMlTvrGyXwD43unHrRzgsjr80yf9BnhQWNVyWswurHoDghRlDeAuEGWb2Yr
RfHP/3DAG5VNMRPDbKOFEudXFRgpUJXEVKDv+2eIXORV8udIJ0pkl1CPzUOqufUOjLzYXtEjaMyq
PKIXrjmSSAQZbJwE98wopuM25Bu/kkONiE8CQ/9rwhT3Avet2aw/ODVSiFd06QHmq8ldRSVP8FOf
ezLDc9Rm395BZXcybTQXIcescp3IFHslaJFkTVQtDX19+Aa0wyidLM16RLoed7Pp5E8q3I5uRGzl
sNlZUGHi4p+t/bYd4FBe9OTSV8+Hljxic15gFmJq6MsxieOT6XlOpOwm9gOn9jRpHOxNNZO/G42k
jph+l6FG9giLdKcpOCITKFBZMDfGTZMy97QMLiSkqo4q1OhVElrjN2S9b4roES/mX04Xk7vuiLCz
oO+8mChlTeWRdVKgzHKm36AXR3QCs/y8wvXzzm4+L19uyWqVVIQ31fM6rfsJzSIgDIPpzz/QRot5
kr2VBckrEumEDpuiZW4B2WVwUC4UBkWu7RBgp/jwvddBnsiRNeUGr2O3G9eX/gKlvxgEluVKVXKK
zBkD6VFyUfUB4ueeyyeDqbrmUhNgS1+Bj/MZXkGjmL1QEaLidfh/d4k/Xoi6VYkxtwP+pNPdpaqm
LRpA3gwJjgU+Sgj6t+0EZEbpdU+yJoElDOx1j1kYqvNdJ6x8kc4i/+jj1JDyIn2vseDcA5U3V0fv
8YJYMTgANcPRW3s0KRpmupOlL8oZAkadVU1yQcWyaPw0KAkgFRuqR1980P7ytjqc1ktq+1rJN/7u
oRpaSW1OWaWRPOZDA4ecY/OG325/sk+mV07ub9Vp5QJZ+3aXRDDdeCicpyQyU4QV/iBLYoVZOJ0S
gxNrFJ9lHUuYmZDt83fnX2b4X3rKHH/7NXZop4Pwi4b+sGa+52TANJCeFuwzA7yJDjy8qOz+yKA7
7vHRMT5bW9osKjYdpQniNL6Q7IzSep0ZQfpuvjeEkOpygM8/NqmWklcXPBclGsQQkk6sSA7SzqjH
aWTWQ7DQpIPvvcuflQBjY8NQ7ep4Cokvfhc2DHA4OBl/YovwElWNo48RLL69WN4bVMqpWY+O4+j9
g1iLdMX1zin400FV0IkqcV9tXohmsA7ASEsvnR1D83TeKvgMbEEHVpXXWYnghuL3ZIwu3Sgn7uE5
mxHIhm+HqtOMY9/ZiP7iR4UJrfirZ9OnkpFULEOKJVMZ8mvDElavQmhQOnHpJ6A17Wujjh0zGSyZ
Xlj2y5dGsGf3Q0gA332oBqIL571YCGK8Q6axxN3/h8CZeeLFsCQJCaWqia+VuJP9y/zrDyuMYQn7
wW03vssMd8nnQnDLY0+PwobyqS7lnIAy3Th4GRehuuaswgMqwVZqwNlpTixGWfMwz3sCwY87y0sA
2Loy9VOnVJDYBuJA5TsaysYzb7j+IniEHYRqNDz/4U1pxP8+cEiy7NXpal2q9Mg53Zp4bRB0CCuX
y77zGuC6oDQSq5fOcy3jgEaVYSTpJcSYMngVwMq2nSCySvB6EQ76iCgi6Qqnh/2WHpneTt+Dr45n
Orteymu9+STZFwTbYYt520p80ZPk9t2nmLvnuYZA8oGfmnrYrqdaqEsAsiVZbNvGlke1PFej1d17
dBpZnkto5rxwKECv79WdGGucHgRcTVseUi1x0WdMa99f1Gsoen+ooj+XpMRkA+O4xzubiOEhGUmY
UyRrfuBZDWlfcMkUv6SosXh6SjCegxw6zEpJGd/B5dd+goOeaG50u7eF+DG/vYF7l/KLECnDyhLy
BkZ6PJ+fScir4svM0UoymK7KdC/CamqT+Kv3Hja2/ux/9U4Bg3+JOE9wGVdQGNipHom2YqANbjuc
sosqEJLShzsRGX3QS3icTGko4V2RMvq7FCUKoZQogJlQRkTX3P5rZZV9KFmvSoLzmyTzGRlq+baz
+7Td8aiSOuXZsTzX7S/Ioh+zb6GNYWB+JUQWBuEpCcEii9aHrLnMzg5f0wTFAsF+Dnup0/d6xs05
Ta+QyWOSo/wkkbCAX/mL/RTj14DmLCssyqveQ/s7SSYxvk+AWpbhFwYKDmY8j+9gTD4i6I5k2jGI
PudnZV1s2UYoepsc7sqFe+D64cW18IHEufxIfyy89crhJYunz2pxAoVOyTD/d3E1vGjShzwHMOSx
hXs8q7lli99DFovDHd43NJfY/9oytDzItGvzx1UvcARu1oQEP+5YhUpIl2SEX/fTX/UdzXMGmVcC
PaBCi9wauYvdChrraKCEjuBNWP1IO2ds87P+Ka4+9CWHONGxOBtnohVKnaH4i3fvY5XqR3rI/Kz8
X4bM3mU243e9oKBuM8efP4Z74DCnlLrCaCe0Fne7gtVxpgMk2EFHwdIMxNedXJeH27EwpgFoufc0
BQdwPmNHU1AGmWnGrg0cPkM7gihm/qIyW77raHyTPdgVGbbZoZZFXifaWh8OuRSh/a21AWSdWrle
tmf7r6JE204UGwNDAD1l2YgzjYKfb/XVgTtmFpV/06jLHdfU5+LEXzcgiQfAFOHs7rgSKJpwncEI
TSMLy6VXjrmpHloGxGgtRtedMKukCHZE3b/r8wSVQ/JLLdhZegyDq0uFu/EcO7dK+uwzMxMi3Tjq
yzTMff/4X/g4i220p10tHvt7lPJ0r2BicpnTbLb6GzPCGYa1X9kY6Lw0Jq1szev0E9sJzYWnpZgy
5CGhNuCltdvR3wDV5HMz36qzKvOu2V66Ticfu2ay0YgtzviNGkZuyj+yNGSYRrZzHXBjDPva2wlc
mvuH6O4gCMANeN8RSuO/lpuNGsn5/t5ZNv0Sz89amTEg9pv1jO3r9Wj+zyBPeI+aDsQ8+PJIvjEl
JKf8bR1u1irfizHMfJrHB5AEb6IjF+f9GndE5d3GW5ym/aV4rJXF/l8EBuzLOEALFGvqp6gGMpfB
/KwFbq7Cd2VY57xvLqt9EPiyinfhHEAK6f+pBgUo3yo/NKwKae4xcZ+gNKYWNAX3y8bMapnTlxa3
koib5DraVp3rthLH1jjxIr7FBaC9l+Q4gRS57SX5fMNAzmm1hovqF/RinsQlLLPB+m+G+dmvsERT
UeDKfwKmOiODtbwg3Wk1paJbQeP9opU+tlfk5wp5hBowO4rswu9IXBPb+43mjDqjkzhHRBLPHQiL
omJy/JfXxLp2hU26+gFszVBYPBX6LNyx8nGR3cpQGnnSsaz2uOlsDJkzUvprHt6T2s7OD1byBqhN
SQdHp/ytYeac8my6USadO4qa7FR0JMBqixGnmqXTtevFIRfsudlDwHVWxYv5Vwu98WHy818Wnh86
a2e8Bwb8GUnSlLn6vLHMuXopRFJ9rGoe73A0+G2UsUtB13ONPJfHssMgLWdNQWjH+ca10vRLJnRo
hTG1J3JQQoGoQLyYHFUIuui+atl7cP1zb324T6YaOmVV98ovtKDAJfkYGO48HTGkaOb1sGlqO4z5
aGMHuHiV/YzBnLmkhKt8kI74YmjVd2Xqt98jLZwUkxvnG1xAnzLPVuahWJM0gluEW8cLWr0GKfLY
9uhP0R/wGiOAL9MW55L6mtOzwm2HTMdICn81e/mjc5bfkZjLeb1HlDmYr5pkFA7NRTggPiC8HoKj
weuUMsfSAbTC+UFpzAaWzz/uzI6o+h2G7TTWBTwA0Ui/NeC5xNkWnTmM+cWtr85dgcWIQKhbhNTt
OL56JLlyrcGlmpTwZHNNDjqz3YZplIXAPyaGAjcA2F8ZIrk5rCTiXZqt8N41/aVAZ5je+G/UxWVa
jlm7blnabOlUqQ7A79Iou5y/CxcYn54/q793dGNvVfViSICu8A4qytiX66mEUmB/jTpv04zJGsuM
S5pMENjPeev1vQPLp2rivR/Kf9yT/2QRa5z6zbngo77C+uVLy23sNRwUowgiwZZvc40NSTXIMx5b
eoEXBi1JenZbkQo6H0lmPtCsRSwmbjBUcS0wPtmq2fgan2GsXPWiz9Vu/Er4sMDwefzfx6JT9q2M
nDN5uCqXSWOZbdU+MO3TbW1/pcgslsmCnZtWMoqreBVwMbd4LNua0cUoaNd8DLDGJFAJ/+nX8m1I
MdbW3UJvI4yfE++qX9IZ4CzBjsgwT2Pz5jAi4ZMcX9MLd38pHhi1z8zM5lR2Ru01Sy/snoELoKMJ
Ro1pgpf8IlKRQl48ggxUt3pBGFOMoTx7xNE9B52qzSfWA6D6AsRTo3C045W4BpFnRDgTNOkAummi
Og6RfF2hFw1ofYMWR/j8k0udbSs/Yw0TpdOrlAxjXFQd6OZAv7nMh+XiA9bnaFXYCtTK6zu7YFd5
qB7aDSucgLMxIEo9hB4TTKdbJ8mHPIDX71yH1hORJHnbDeHcx6ULMFAwWOe4a+0DbVTBigIlVdxC
YfGkUAgLAWsCWgOavd8zcjgjehFLtHLXIacMzYhZgIQvn1foAgAmyCIC23NeFqDf/mDWSGFOFilS
QUE9gweOZtVg1TkTByJ0JjLiup9TG0C11hj/GxMyZ16NQixpXRnD0zIjVqo8IR3QAgs63XHrFX5K
4eppEFPCaDW9GtV+Xfydcdsw4MN2jsdbgTbutR2C02PFCP0KdW56Oh9H2tMTHiJDOnBW3X+9O5K0
8olYjEO+B4hVqocwxI655gl2eLK8nKdtnEXi27c/MiHrxkmLnmp3cLiADauz/WeVCiv1Xwbs7Zq3
fLeZ7HoauSxzt5YVxxbCAY9wkt29QJ+ZmATY+ZGjyWyOhb5pceNpBhNwOWLdJbtkpGUIMfN/VNfV
/VnO2ntOoR5YDVw2zpOcNML8+XocnbRJ79kHHeAnVmH9Izu62BHDOYrT5LLIUbDGbJSArbT1UfEM
u12wM1Sc9OZt72X5B7gCXX2YyIrY4bWaAkR8T1H2xfT4BshXIfSULPkZwG5mNLKjpsQmwTvZruzL
NU1TcvbSkuOWDEF96Njl0cuB8zFK2EYaJT/NYQhzJRgp7Ct2RCMiGjWQrEXn3ltevQQ+QXu0JHPz
KIC4L/KtvaVH0m7/XI61dMm492PXyCfItoeQm/9KvfTk5SE47nFd1zbRCipAffY+DGkmbtxDJd5s
E/UT6A/i63IZp/u4qdEVMMdijE+C+tJpTbtcwI1rQ2+VGO7sHBkTsliiTx+fL2HxyYtUXKelsB3d
yJ0PtiaKVqVc3sdmNEAdKdXiytUxeYuPd/6gl+MuF+A/bcK4CXi1+654tzqqgs7OzGnR5hbgltOg
NIdNFGNIUNcJK7ybp/DxcQDv0IV/Hg9jDu+VMuBCQCOAnud1n9QKnaDi1GUJveBN1fPHrzfbfLpG
aEg+Eq5fUGrkJmmNo0r/EAcgj1GynUI9TOdBmbL/cc6p19tRcKkpy2U9f2oYit+WCTQzxhYppYd5
mKBOwB+bDAULcXZHpMMS/80XrD93VhjvjSACIjdXAQtj2Ki1tmig/r8u8qtqnCFZ8PreeEp2YQJw
8+Kiq6zHAuQq2KdWDOSFrLqw3SFhqLpDSWqHI1rxtvB5Zi4I7gNnYAIbXzYVmb5++aUMtUZ3M1RC
OGpzeXotaD6izm46B733wKMLMYaQ9rtKCiWLjThOV6GX8u09+tKj5kFbLNH5yYhuxx3KwBmucXyy
4chX6ijClita1mR2dJh2xcB6Nc/iFE8XUTaPDRK8lcl54u0q3KGaXqpDFccFf40lIKTrEPxSs9mb
2HnfaWv+X8maMukZDf/0qO6xpAwdxCehB8kQ9i07r3bCMfWYUMeCZlqhh1irF4JqivmglDiarxmO
8F7TvmDLWUHuvOFBYK8r7Z/mTVWnRA2ldDuDUGZdhIdOfV4wYET3mfXltZAtZrgDWlgRbuCWWhhy
vFSeGDsu+A2DJ80NCQfiqJA7Zcbs/5gEubfenbjkhsz+8WvmdWaGJhKsDb62jcGomvudF/ejCdKm
h3woFoGL6YXIU3oH7Wgh/6KmvR6lR8BNedfHJ25x2c0KyIwu0bcOvOzCiON7Y2KVdZfshfHQGEIN
nhEc/H1PSgDMaR6tGXKNR5F01AZIwAtkrPlUmKHHkkWvvPwTZSXlC0CUl1ZyfrgslgMFdLQSCHec
xEq4p4X8wIGz8FuGHeVdKew8bHQRpiKW2fYok25CXEJ0+SUXzGUsrFipqzSSnkD665mwD77lQtNU
t19jIxBg9D9RxQa3uvI9g3ItwFh37iseyoi69wuLzPd2lg8mDEDLwEJRC45cD6y5xp91UXI+17sX
FKQFTWxY9tBsc2X2ozfy7TvVKvZvTtKZFRqhnZdIcARYKwf8dQfIST7coLbElP1osS73S+UQ1wY3
y9txy8VXR6Cl57M+4irDf4QYQjksqrzRv9mEf/ZK+0JQsSXKGEiD2DqykseJKkFm3tM5hxRWk0h+
wd8B9ByCm+KUxOSu008lsa6gCf9hhxUuklbWg+/sYjLcnqRS/Mote0rylIOdFW4+KytWGagfUaz7
s8ob3hFH3MeZ3GZCEeSEfmwJPIUInX+ZbvCzFJwmu9jlu1qDMZqGLFchZU84qIuVHIrtHEmfp+Mv
z1g9BS8PK2ZzLzUAazaELREcjrwYyQdwEJ3VXv/5c79ICxvR9Mg6Gcw2jull5MaCJjapWYpMdX68
VJ8qHGO05d6o8y9ZHzAXMuSydrWXTMHH73KrgOcNKXGxT72K1rBGw6AbOhuZTR3rd10QJQUQqLBn
50FBlAXP8sgUKj32UwOmt7NMcb+PiXzDTVtF0hayAYVN+wORPdxbgbkNjee2YyzLO9l8KK2H73ZY
4RT1K3inAbXDayfxES5x5nh895HQp+ZD4UjZ8iuwm8vJ+qSbyd/dPYAwpvPLANsKspBhDyfu4jlf
Gf63XXnsTVxcya+xX2hdN69S9e8hHxLSpOoVr4cNI+6qZayZbMZP4J8Syfnq8LD5Zw9dkt1NB5Ai
wRAvOobAxJuxTInvBr3xZOJF8CNU6FZAjjlevLQkzfIBGiuC27JsIMH47FDsabVq0t3d2Fl1mH4C
nxdF020kmTyXv2FDNI2Xy6Zktj6Dce+oOVBI7tSCWq01PWoWuJgQG8pNpV4DpRS268fVnHKkMOdi
JP7Okp+hMu4fHlGKW889Nn+dQIIWil5M+jzpFu8N2SFa/nKW4Y+WhtPkVFSpOodOWS1UuzUDX4ls
eCJzwlrFYRt4nKb7+tBCPnxZkkrsl+iAjm7UMBNzJ9It8a41STAiB26oOmzHNY7JPiFh4aBv5tpm
ndHWZiRTgyHJHSrwQF/O3oX1oTvCogqg77jFyDIsYvCUocekUL6i1yP+cj1potaYRs1SilluwHAX
6R05Rz/MyxIqt/tROOZDqctl1EBuCuMYcq3nhf8XK2EKeUHSu0zbuaWy/5bIupkrb6HpzBOTRzfk
FbcSN4Ed14vtMhfdFRo0xVRAfY5vC87/LhU2pyPTgy0aJw0m6DCj5x6SeTVQI1mVpIbm3W3vlTcE
LPNEsSqIJR5NE2lgCff+DAACVVMSuNbYP8CYUxgBRzehxRb6P1FCY7EcI+mi45dtoYsyHhSR/joi
1udFM64MPRU6D6GzxIRNFeCQdy1gHDgPKBhbTGBu2xdf3IVa1WGxUOmNFxyUR8A3Zten0ShCyPFi
T/CjihmXwnSpFDG18KZizbWGE5dvp6nEw+20Aewb9fu0wWIUgAIbU0SVWBTVXsVZWoTpjSqWXuF2
N1ViFjX9YkvgNAU3zmXP7o7TGx0FHqOSGsPys9oYcgMFbn75IqFcuFPrfNd7ZTghNJlAN7/ZSZGz
vc+8EOeQ3E0BhMSVFUmDxDiMOg5movVWGkYvsmh/tF4YsJzaa9GDadKrvRFW8FoOX2HQWOudEMYO
25e9E9Ps+hXWIvZIqdFearqujS3u8dce3rbzBcPE5D+1qVAg5BAl/MjdvFM6GG9Xu2LxRFx0xnz2
u0GEEhTObSW3NBQWI8hIUIduiBXXpw4/wxFNN52ArvDaUJX6ySWrGfn+aSlkLR8aOmbCety5DUxn
yeedxEj5kEUikw2H80q1qwcla/6NVXkz1j7tBY8j+4vNNiJxmc8sbATxBPxWQWvY0jKfb5vNwu4E
2CM0g74kyJ174ctkpC1pcyHrXPJFfzztsTl/QQ0sUu4sp2QcPDUEXiVNXBjySjt7K7WsgYcogEEV
Zb9iSfqFYIW93ZNiJlof43hwdKenr9DL6sqOYE7W05klHFnAOA8Ow1pJ3OQhN4+BelEpOFupm1Aj
XnriPXWVHFpM+gInSWcRSEZWZrMElI2dQlN7zytgP7+HLvXrvTWW3dJv10hcjRwKn0jF9FsfJBzK
vAJRQ5PAYawC0O7yX8bXMrdBuWLMnTsKjRIfVfbKCV2Gs2Jkn2cvaTWcSxrJLUWMznuY47UBecqj
y3lu6aEwyY5H+qbOCO2zUnqlobZ/uufT4YFrx0K2/jqE6tWEeC9yW2auBloXWyB+RVovKjjhSs6U
NjsaBhZ17uBx/DiWMmXG+CcmeesMpLTtT5UrfapZMLge2EFVU9JOrseKGCC6fWY5jVU4tsaFtf9f
NGU5/OyklB1nfIbdFfYnsFDSzNed+Ioby/OnsSdBt5k2tD068EZHQYeJJ9NXrV6qK6z9j4v2DJO8
uDQbuz8bf7BD0D70mNTaYHyPHNP90KmkSoXAiXLU8WZ0IxSWzJQNCaRnaEQl8CchkKN2mblYwnUR
uZUj6mkYVAVhhucBteGjCCtZ6IBCQBZAA1g5yW0XxelFHfjKS1IiM+mI392WjR0gz6/GE2Z97mu3
e0x3Zy5DTPop1J/C2IvIK4BO1U4uXuxiuQnN47MlkErITfcSKHrY9eaSXupppOPjK3uz8J1AOEOO
WVi/jSoNGVXebYDyw0Rk3duAYPjNjV+2i3/ygksWbelg76BD102sVCUnqIORcM3bllzmhV/hihgo
0BrJTocoDI7FDI6tp1RhCGgUouFUID9JJMkNKfCRAOrjJwzc996xv34AcLdFyDiuyWQ6xnKwwCTK
jwyZ+tUbJOnuaLLDKDMDgZsAgGsekeCuRMr9vumm7ZrruxZLiYVqdJoHF781QYowow1NgX6by/gt
1eTPxTGF+ef0Si5kKKCynZe76QKXr2WndSnC9jn2U7v+SOxSLPe8MR81Uj+GOQbPUdBvkW91qTTQ
u5MEHyFk7Df2A+OIlSv8e/am39me596xjl1r5UHsTMqkTiPxh0JGGhkFCHbnxoVzEtMuWMF7/h4k
0kEOPDpPb0AbTg7+SFx9QBuXU86a9N7FzbUOymzg4Pbqt2PXK1ms7esJblzCJxtlDIxUVUcjpR5l
40yRgpcAzYKELFEy2DK/E7MitQQX0COvsOkMsuhQI3gUialIZvBStzN/FP2WFf14DGeed+YyLYF8
L2uNPyByXbhU9NfA5ZQfA3Q6V50zC1H+vgv5KUm718BrI5EVQXghCBtIaxDuaZNCh3bw4l6SRnlz
ne/ZFw5UR4O/08JOgF+Mp0LUtTOnQYjTKX4MlpUks8014oR4iHz/JV8R1nrZfx4v462N/Yaq5ytR
WlTQ90VcFyDJFqbTLAsbNl8AYnx0HEe38RW52l2hpZ3WZiTtmn2i6tahbvJf62V6ziV5neRcPp9Y
/jp9+STFw68fNvD91R1mgP5Uh0zftWh3wIabR61BtVYOhY0I2doKwlhoSdgiu9T5+26CYUOXkhoH
wxxklkxpdpwzZ4M/SlNBuh8ixCKX2cuT6X3pUquMR5xoWJJd8ZwJZr/qWM4MNMJBgZVjG2v0JCTE
6U5kNYLSjF+K9wFh3OLyER8Vjvf/nQU4S6FpPZSe0+2UdXEgE7/qG6c5ENNWnrBCaql90oc3lnyb
M1PpAjvFR4jnaVgCfjAbbLcMmdFq9ByAZepWsCPBYO3fedVP3uJr425QfZ4rO0RUgcljzLjS6caP
s/t2DU1icydn1X21yumwcrZ5bLG0dvw81uEqUJf6LAVeODkyMX4vbKpEsGGt12PwW+tPGIOuwjpa
NT+JjLbJa7TJebvApEenbCu9BJtRr5UME1vfRLNtD4BehNxn2CsoBmuDWxDs/vyYIMpwNDVxAATJ
qnNUPwICkOSMtoxyIShhIoXGuhFw51AyDioY90uVH7UyYeffvfj9yBDE/H0JuADZSjCXlsm1Mfzh
JNf+5wl5I7fiRO0HXft8GIK3KBg9aUD8NNz33xAk/1NNEzsK/To4NRkcFbXDxFU1gso37wqzKta4
xsyUODmjs/Mh8A63RjQoKo4aHkzZRpCUg+IR1CAu3f7V5Vtk30izMiEQbWLa4545kgq62yZStZmA
C8M1bILNsjzf0mb0G2yhqKvNvj6OdApd/LXJ0z2EOWPDZ5AZ1PpG+3scNipldBovECObzz+CUxWk
dy7JCAtvDNcVXDo6Xt0ZRW6MReAkVgJJZkHbHV96YzSTYI9DRuRq5VLgj3yQy4zEgvYPwwG8v7MH
9ARH4Yqemgs9Kz7P3SUvjg13cBcQxDH4uprwyeMSAJ+Cy8ZNgIhtdxDTg4hoU19d6MHI27Snm7lD
/9C8X6QogZwcqk2B5xohUcaBu6iYJSfsxcmq0kJ5skzeHTmRdlLldZ6xNAK54WUkwCfTSfLGNbXy
4BH1c64n7yvpeVSlfEzrulaGHiPlsco/x6KbleYEeKogJEPfWKtYRVLA1T2TRvFxlgf/9XWJm1ko
Uw+QeZnyUwTEL5mxRDenyKDmPZNUv/CWkIyV5EWMxD4rVigIGVcjlpV0eu4k/vJW2oXpYjq0MpJu
1dgCPkpiK2QQiVuZ3MLOqKNbm9zMhiwg9iw7V/Y33HG/CI9/bSaUpBE8rIZaHqKfLQ5p0dD93Sy3
lIX8SCrVGI5AzflTyCYcRvjobXO8L10layV4A3J8OSsDAnd2SRaeezB2lITRQeUwrX/emX/eDTTj
0o4DiL9q1W6gb1UBgDg70qY8M1xKD6cKtDHHtBmIwA3rq1ds2D7kiSur31OzPETHoGprl4qhfPV4
EhgTJx/wusx109RSdxdKTIy1dPn71ldGq5n/HpbcCg8dQhByfCpe5ufPpnJYfDyY/3U84YdWPJOo
mBEm+udNNb2DF8mSGCUg4HJZGEm/CCGL7zhOUrPUpNEbxXBqeIW+/NS+uAT+vTgeRaSxT59CbNTt
Ao6HTwfgWYekQrxWTAQFtRATuRngxR9NmURf7dfpP0mw9/RNhj64b1j93N1UdLvhNQGN0wXbfZKm
4AmGhE96S0PjjraNOOHPVcMJ9THjZavFE0jFOoschSNS6cjD3QOZvuTsrZ6WibV8kM2SN1bYTMDJ
AGXWpKEcsN4ew00mDY0e4rcpPIiMCW9DrhxzRNaJ+oi2Sq6TmoVxMZ2WI6hp87Sa5x0HtzuSzeA+
7EHhP1CIUMTB5x+7xW391xYsrHzcCOtces8Pii8icE2JEJ3acOhUGuxg0wcPelisb5gwtDBiU66m
kqas6fbppqt5AKtM2GLW2ZQ45O+YPzgRXCUZ+pgqUKFp6qC0c4o33B5QV39nw00ZcyMAO8JtgKlR
+bVBy6aFzs6KLLQjx5/fv+EiswVV91zPvAeTaeuRY5F+Mz0Rd30tbZfe9QfkdJJpAI75H++uTpon
//N26joaoTN/3ECCLeMtbXx6257/jvjqeCf1M5CGQyDpoh/e1hBPxnSfUm2d0LOErX93e8Gf/1Mj
4IK9DwGX6/EInyWwaTRBd6f01ZMgdnAEytlkBOr/WCg3LbOJrw6AO8v5ZjMtNMlJEC3TKndnbQAE
5xvd6zpMIazytrEnUAVNqS004mwR503raFy+MVSHknWbAbbLLKQN+jbEwO60LB6D+6fXLyyzXk/t
nBcJ5VlU+CqCRSA/jd1jofgk43tk+lTlM5zy5PUAOMjZBxqD5X00ow1UTNCXYcjV20aQ4bWHoAmA
w3dekm8BChPgIStrLO7yV9E4h7ODeA33r41i9TcjEUbg1M6pRBH90FglCjVAzbyzXmEp9CAloBJr
vGvWCH7khkD2e3hikgWwKKFzBLvrLaNnUQXXk8m9PdZrx6iBHUYNDR9KfhnuqqWmLJR86lTHfqIR
AMLVPG9Ij4MVOsmJvZ2VtfrEuWLEhC2YY3k1JzhefxqlyZvHPnaq5Gz0jQWPU3HEmrYQbpAVH31e
miMxgBOGbwG9QmYIhrRYYlRob4ciPLAp2KrbVWDbBCoqEaQKc9zMh0kuHvQNre0QUviXutD5qQKV
kXDWU+qCAXr1jj/vGQEvSLirXWeUDV/xjYhlzZneNcC528i06nLD6rRakIei3gpCjQKp0UGA1Pn+
WICVxwdhQCZhcqg65sRZtirPWkgMlmPXlhMzu1549Z5mWGARX9CruobcojSGP29Tpxmzh1xnWQEm
VWBt+IR0T7FfjOvXkg1jOmqHL1edBjeiYq7Cirw+UJklZEzzceCGNRSD+bi4Qf+QKUrawWiQRSqT
4rBFn7itJd6A+JOl/0BmrbGTtKSeatpI4jVzZTkPEhaXv16oTkS9kOVLD/+i7aBu1Vu/t98KoTQe
KAIv2pWI80INjbBtnWgPZJJHaRjMACNQrqfQMiy7eprFLhu3SPgYnMoYmEht8gC+aLp8kuDMoz2R
v1ze2Qitil3FaouDcJctM1CL0x+I47o7tMn3ZoXzMhbtkcQEHZYEFYLYixTkxBt+Ml/bNPGh8PGU
pPXptLCLn6GLiKo2Dyq1YVmsJ3pXtj/so3LwmOx1onqmwp1dt9C/USUylvN85MmFcwPjleUcHQFn
wwZnijWfYeohLOWH47yMa3xbpHvdM3iIjnMd7J9abRl9+kFr4077fv20o0krRXTNoSPX0bp9+15o
sdkyyzmuUN0jPye5RfLSWTy5C9fsy4V0Od02/aBDacWveg3EcOD7zJruCMkR+TGj9vhvaESIe7UP
ps6PmsgvC8pjci1iwaIBhgduyZ7yJAhn0RtqFAaasmb/IjTesjzwWCMEznMo/vAHc622O92NX6K/
Q+DLYNgtnokK3HkHZTblqhxdW6oVaQC8/rUeSxOZWOE/tya5nbJYMlFpT7wJYqOf9Jdtkxl/+lvq
99VOaM38fdfD+2epWQKPZF3Fnm1+AgqODIHb5Xxc+yNgqFF5gvab6oQRcb91O9ZuMSVYLRKLamNY
dOAyhdbCCo0vKR7d5exng+1Yn2fRLY2WOmBf2wjE5bJHIbaLQRIMuxHkIapjjtLoK+eAM/1l1MFr
r6PJcwzs5R+X0TQQmaJsBooBZobQU8NCB12viYN7XHW4emPjwlvifGXBEkJ2zHgP8jq1UG3l0KXc
fNZoGP3VU7nQO+iV99D1zmkmit+hewNEJBfJ9/iFWFsrcf5RJ7zf+oQbaQlp0psyhwFpj6Kvzj76
4dLCZaBIvKie4bXga6NQuy6Jhp5nr8MPUJlDLGQA7i/53o8oE3cE6nTXB/In1KNRxqu6zyqAfeOB
68RBaov3CtpusVhXOHXjisl1InYtu3rec2CGU22wB/Ltf1zL5OvPxq9270HZXiM8P2buBif1bF4k
TGosKugkAdwucLiVoMG4sf9YiRYWfyv7nXifqiQrZOa3RLTL4e2c0yippre+eQ2N5hP61ftN9pzk
szoyTv/xW0MLR6DRN9PB0KdaWsDhjSNXl7hdREe24RnmVZdYu3+SWuYD8JpgjgXrsmVJ8RaJ2geq
480VPWUFMsA+vMU///h7G/BxVOmZAzKMQg7TRF9kVyuuPEC8JXOY1NX/aaXqRHI0p9R6+oVDTXe+
axo/U4XsnNsf20db4PzMa8kvFUJ9sB7GrJuLN6Tz49xmsQPwXWpKdVZuRmPurKSssGDWzDbSzbtI
YclcjuKFJkEcBxturZTNOqOo8n4RXMUFcnX58l/5U+vUasSltuGjljWvfK8Hwd8tu8wRiVHqbYCo
4tKrZjtuO29Apcj8v49Pshnr4DL82NQctpcOjIONZNkb1c2aBhnX8rD50Zk85RTpyZ8UhzWjutXa
qtdZlj8t7NxIYE6PYJLvLPvYR2AWLnJw1T/49iTaQt/Qqi94l8z1uG2cTG73RJqVkbqN3FayoJZX
bVv3DF7ebjWekdha76aLp7qYS0M5Lq8qNYWX0YYkMg6rSON4dCpV7UEQCC2xskSp+aZuX4Pfu+H2
vTo2b8nWJjIEvIXl0ok8v1WbpdnpmWNn97rf95Ucc7WosSRJQ+HPhnquDzvBVKq2FjlSCKXEne+R
rRVI8qSRpxHA+eM1n47GJqnmt8v8UuemmePw6WvB2wtEkrkHnJFJVlse+zLytQuCOHDfsrnWWz1C
j4DGwdg/eLeQ7Bv1IYg/op4IUWwnZlsJ7eu48f11C+Og3kTcJ44BD3bhsDJITSK2D9RY5XB9JQ8a
3uet+qJcrkDEpFk39I9SgfXi7j0SExt2z3VucBWZQswdgRM3U58uuNGpSrAoshLoSinVGFh+2sCA
9F7YrwPFrUwMzgSS+xBjuLhjuwEp4PsXQ61EndZmL4bvDECG+xxnNPjHpGNmRHhoHn0SakqDpNaP
uVw80TzfJT2JripJ7kZYBv+xEBV8UpFNMAJ2g7V+ecsLPeek2w4rHPdkIyGFV0oNLsXN4TxYtULX
kIP9Vjd1VGmOrghOuqTr5DuH24RSDdP0RL544I5k34z85lb7aan46H/lr2bypTpd9Cw7dOfNTR49
ywpTxiUk/gvW0Hdb4hIRxK2Je38LYAVLJknPSOWHU4Uqa+gfFslTHL5x0DQTKK2qXEe6yYWWT89l
qQmu2OGCJdaL0lGOVRphCpUZb6Yh+ou7/RGHLdHtbgDzy6Snj4XnL8cdRtGJY/TKVww3ABavGtOp
WopHsWbcf6c3lWyxReXWg6wNQuF/exVwPI4B03MyPDTg3U5+hoAHZhxGl25nM3Nwd+vdQDRqZReQ
J5yBY3bT5hOfF3B/+mXFKJYeAFsD2bB/QF3yNqQhh1CuapwrKkY5yFCHzP2DGA037bsx6S+D9ArC
T+7BSV7vOFt2lYPunHiZiRY18wFGkbgluLvuBSCcUmKudIxNFCGCcWKcLGONZy3QZIpVgxYYX3UO
jZuYdIJBLoudnaFPXkbFr/zYBrg0td9Kk6wP392aBMz1g4KrseMGaTWhEDTzELG4zwoL1zoCmwg7
d9WUcHb0jbAT2dMzW7mous36/cNRxgsTnaJeYujJdVUV2MyuTMwPzV9Ploh65N3qqA2Qki2xWNLG
pxb4ifBkx4UXAdemC6TbIu7oTTOHOlpoP56TNDw9aTdmRqC9Re4mIlBercsPdGyF0etnXD37XBge
jGQien9pxWY9Y9Y4Voz7GJwqvc5R63x2ID1kbm5A1RExNq9ELz74gAUw3XFxPw1RNsNzZl+AJV7I
b8XUP8O+xp4oO6Y3BPmU8F02sSPOnth4JSF39HyoPA1AUgK2rTyxEHiL0buDdfaqAZcaz00uLDOs
5z92FClwP/Jwyx/iLniwaHN/BbFI6j7N89HF2pN8duV8bvngExnhNq+Vrl4F8aTedtazsu/jjjUc
+DTPojXBq4+q4BfYwIWStEi5lc+2HyU36DNj2S+B74I/dZdGxZVsl2fFrouzdYQVcLOpxzgsoCPj
FbsqYpP4q1HiK1XEiR3WeTVwfj3qll0D85y+H4UeVuFkrpn19yb4cDDjNz3fuLdTv0W849SVoz/5
MbNXI2cDvjjZHttCZH/t+z3ImIsTqFsuDHyqbENTdwbZSmq87+KIj4wBzHS8D08bsisKlqPldGwr
WK18t2xqn6FmwpaBXON+p6bVwFHOTZ7+DewkJxYVeTaUhz9qj8m716C/uuAcbiyOafqN5EoWXx1E
CvALMAwfdaYOpBsO8xW4k5PiBlDuL9At1/igjcpP0N1HvcmntGyYA+EMpCGWN82jCrLdI0muQCJz
GGAo+5ksU2aUCrvTDkf9bcW6KzwsYASu4Jg5moPlgXUtYocT6vVpTTrokVAP6tKc+hmLOYw29mbv
YdTDPN1SeiI95FtVLweuOIk1NehRnG7HfaH0Mc/s6mzs7wxeJekz9i9LjA+8w2PNqYUCiZaCRp7o
u4yyEElYrs6I/avxkKDotkycrscvd3mc3yO8XoW6roWEbXe014vCl0sEzfx8n+kJCFGdKjKJlEkH
xdmv9w1zCRchkUlvaDfzwbgz5C4eBtmOBmQDdWljJeIGA6PDthAm6kFaFcyqxcfb+zNUeMX//1Al
mK9hhA+d2G7c2GjcDpZ4rNq3VkoDn4Z74ZYamVS5XWUOQyjHeg5YyIkeE9buHwXYbYRz51NAISvq
uvBgBCLYBQTA9+Zy4d0fZycbNywaNfd7zFhjvlJZRXFSQNt++5f7fuS42Y/hillnG/uk706zEsF/
ZPCbE+CYXLPHBLDtrr7rf+b1TZj3wxJ+ZZPnOC6DOZerrE+LSuiRnRO0ddINuTox/Jrc950Gltwq
mxi2dNpFyz354bfA09ykt/SeqEq2f0NaHNf/memd+T8ON8UqR2kpjdWtk1pgMKGbukWoLR7tYOPr
wwgLOqwVdWJbWe1GcJZmYW+RC3LkYaaGazlMy2Mz2kenOpCAgOflDR18eDSNnWOLtZJxogNOSvJ1
fTWrthYYKTttVsJ7M6w19oMOjiWmM9loT0n+u4jNm6TXgy0qpt9zNhE4UOsKMrOAU8iCdULZ4r4Y
onqGWZ6AXOoI4ANmCPcixqjxFGWEfBLnTxXGysCQVfdJ2bdZ5tpBtNyVX+VqoryP3r5dx7U+v7tq
3COefl3ZFLeRN+Bd6ftgCdcSEfbKxCxhlVDEth2NRc1EALm1gx1hqZQrJJ3rw9QNf6T2TI4FWapz
V0jl4m/6B2zUYmYhr6oMgxA6ftGN1cq7fpAjNCfyF0xv+7zrGi074BeRXMsN5mlMFlYvV8OkpDVn
VVH/44lPlxGqX2cE7k9f3NT5HjVHFt+7waw5cObQYGpFzPWnEE2dN7CGNEbGVAmkKgZ5vwNE13bU
gUyW2aOwahIuN8XUbg1l20e1KGY3dqMLRtgCFM3vHDUxZcxCzSt89R10LRfeT+jaXyfODO/Lg5Jq
DLRv7A7HpmwhgkaQmE9KxeTX9384VKpo8HjcWE8PHxiIkz2ZDMfaMTiQCCM6HXtHuiIfcxHS73zG
MqaZW/WGOBh/kbt9Czr/42sOXqAC2RfHqb562wFB0hrD0POpHTO116uLCTw7+r0/KpDG1ifK0EnU
Tv+ltR5hAv2KiCaWoPlnfbVguP+GGY5p7HW8BJJKSIVRFnOfBp8QIoVIiUV1RhNKZDIgZnMglLze
FvCfPURnVO9HeIBVec+y/uyf6oYueDGF8DNzU+qnbmy8dSDHa3ZptQEBjVmRXTzPFQVk8iT5qkmH
hpOUYV2UnEIgq6mZCkPLy5twIxMmOlJxVWs3RLirACO1KXY69Yvfoe+VBysZqtaTAkUxelRELIAH
DStwrNy8Rk+jXPIxyW8FNYZRqJa6J6o6td2gjTM7kGTTZq4zIPvn/IwHsHiDypZucsF587BdA6Uq
kGGTqfv2KQ/52Fqmwd5Lt1cvcsQL/MQnJgRFx5N1uyvHztHH4rAp+uZbOtGfvBw+qgDJfXkxDQe2
Nd0qe1UY8Usy0NbkWfTDs1EesFxDOT7751jGXuhBJRCwxlwagiVAORScpWdvi4UBgwvER6oTIxUH
Or/jHTnslaq2bXWiBav0g/9X3b6RkdskB3w7XUK5UR3zdW4GWw/kJjCq3yF7yOCAwTKjHFDFimDf
kYhsPQqHW58hdfdjFpEa1EsplKzjCGRQgoqwAotjBsc8B5m2AlUi87DgAl9QTT9UZqziBA2kVq3q
hHFmn3i6G8G22VHDvaoULPLSIYOXhjBag5N3CxxbBLgndx3W7rUIi+zD/NtcpJzDgJp+bAeZIgJd
52H8iUS/xej7KpGd0kUE7scl9dEoiM2+ezggKtIPeqV2RskcK4M23n+MhZadycYoxv2resQRS+WL
9ZzXpWEu3zFQPWr7ASi4WvuQfw9Ks5Kiz34jKXpvLR+vdcWL/CNFL9oOxYV2Pa6GRS38rKTG/8AL
LRC2YgsDj51+5fSDq4BjsJ83C12djywsI3Q2kZR6ghoRIB98WOj0VQBq/FreAu2gtnYzoFsCDZfc
Ha2b7ae8B3JJuhxHb3p7mIftp9wPSBKXjVsaG88dQSR1xASJ0uljLUMYy8lOZynvwUOGW6mgT/TW
cs2rH1zVYAWf/urglZ3djuG/Jgz7s+hQqip/VqYNXgVR0j3Amp78CXQK7EHUMRgn60eQaF+cBgjl
6FfU2grV2y9qJgfO4onqBsjKtT5I1i+87Hc1ynBQhw0gFZFBlnHvoITT8QtQRt31dyAPo/bkAtNW
q2MCs21/kjwo6NbL5iFQjnyE3uKwlASqJ/RB4rR0dF2zS51LLM+Yeqtm8UEcB3lWADJSNbhQMgeT
R8UUoWprZfxPSan3BoQaqvoomHZznAFEoRdFtCVGASWrMmxUzFW8QW0qvnipimoyklSvNE61rSoA
lprGtA1P1Pg6AFpW/L8lL8doeIrrQZbDQ535vY8Z5D2dSG+o20aV5Chh9wxsnliTpqTUevOtB1yy
hmth7ElfE4ZAAiA8eXrac7WXy8i48qeIPcQTSgfKxg7bMWDPL1BKCwnkBDTySfl8G4fA9WATazDZ
Sh4eqWnj7LqcDyW46dYMXeTwbtlsSwuErFJfDZhknffi+JBZeltXwaPKkeggFrI3QC2BOX4m8lWX
jAWldDneVfUQ8D0gWJSbyfoP1CwGLnOhu+6RKwoL7bSvxFPZy92J6JzsLZP3n6PWbJbRkv03Cy8L
P3uk1O9/yOHF+yC0ZuD1N6nkSIyukYBJEyfk78kb1XWjmElW8H8+BUzcFBN7qSecGS0H5Ce4DYDY
XsoMMu65fBlP0kqoKB+x7WTdBalOHJ699EfoeeWAAzWiT949q1c/CgO3uxa0gIhGTeyFqVMoT/J/
+Y3W4xtZTloXaQ8i/KEg28NZRPwVcjnoD/4mf8oVltVQK3Ub6x5O2tXFI75CDDYMzhP3iWZ9Say3
pkSsc5e7chii6UDPGoRxY2tZwbFZeb93lVNeqg7d4ZUb/vfo3Q0QyjQo1Xua0LpLmDtV8V6GVfeE
g+UzHzdfXeRFVxDzCwXrvr+ko2OpF7T3CztUV3k5GDqkGWh7gbr3XUdMuexbqnBE3iQ/MDuc9XyR
noUbvS9XxJEiZvZd0Tz07BSoQMvsF+9ZAiZICRPRMZltw+bNTOyaMF7E5G+mv9DQIHIokp6Y9lwV
WH+1267bhUObilA6+6MX6TQkp5Eh5T2dXuoXgV/G22Lrt9bjP7oANXrA9FDhoaYyepIvgxD3+C+P
TMp0pW8orOWhndQqWJdFdnmbxEX244O/cOOcbG5XhrhKp3keH1OVExnOjCX1DJ4ze5BoeMa2dsuy
HY0QHm1OnkgMVKlE3/U7M5radKRHqZgxOZUcP2dWA9KvRx95mC+1/Ou17HE4VPV2wLzvSgiTZJ0x
BKb7GX48K/Yw2TvdNfnHX2mhPCXs03cPE/OaMAecK9paZidSlkj0RYMRJVJpRXlMB8lZSKRhXTK+
vs1ckumF8QjeXkqxJGpeeCUxVIdiVoglq5BD+teNap7sXDI/2S3vGXrWpOo/weXCOjtFojq+Y0wz
wrTpm1D0gAW5wT8yROwdrUfz8LeAKQLjyChatjXmxDp3tNXG+mE+tHpv1HdlFfNhBM+hkvslBYPb
cZWXVXXtNGK9NEjG+3DhA+AoQLd2QuMYr9Xr3ZChpN2H1atfeR5Pq3FyD6y4Ou7X63HVdp/d6mWI
4vPodPiNReHKRbkddEEPgjXN4osGAjJm/LUJpCwDsT1zNJRSqKNlLF5EIMjkj2QDHc48/G4gQD0/
EYBxFybe7uAjeyQu3c2kGn4ECEkqjhIo3O//MuQJ6s+zRpu5kcjeZ1VK2FKFBRheSqshmdkYcVJ9
vlxIyxq5AnbD5mDc9WdnHFF3+d10xgwak59r7DDyqmmnC7SjTaTas2FnbtvCcth3pP0oVHuKpPHy
Z9lXgpCzRVeybNIR/bzX7tFxQ3FTWZxObi07D3347Gs7KcBXwArrTn3WZbiM2hsOXPJ+srhJ0CZM
o6kBSHR4LZuOuEWFIq7N3uj1jQEkPE38aUp7p3pgjvSL4J76hOwpV1IGbLrEN4Yi1Fk5Uyy308Rp
291I5hkVtJx93E+e8Klfem42U6fabyWau7PCRMSaaBJquMliA4l/Ri2Wm4qyJRi79rV2FS9owL5s
XvdHz53ufeBRoO1JcaU5eIWNs1wdq6BI3UGOHh55dGJHeG39rNvnS/uSqzEPhX+K6QUVqB9MQSw5
TFT7SFjFSiIynLhElRO7IxbYcJkvENlUzfmRsaoeJqZ4mlxx91B2BlWPd7JJsTHyFlXPgH+V0qHB
tojoyGr68OgxFinVPkUibOl2QmhtrVZ4bb2bB0T9oU5iyEH9YTD2Z7J0r8r3g1Bno0ty0mTK0pWH
wQ+QPwlsuK6sO0PcpdxWl2DTOPyeXBE0i/eKjdctp5T79T49i0w2NY1b+Af6rMVpgEQRYfa+UuEH
PNmeH/eUW8H+mhD8YZax7NDh5biwwYpumX3WVH63Lx+G5hlqRiDygHKxH0sgQpixmdQY9eJlxwLp
gzuQzXgi1jCJjAmpPpT2cqrXiWS7ERd2WKI0mjKkTqGlU1Bnnbyw9zGcV+Pi6ygZ2G+nZ/uAFQTS
E4WTEfUZ0PVJRAVBxZ3xe2x2XTNUVwD9DBioXy7p8sIKoCRVza3+lNJ2krgPHySL+XYMACxOz6gV
elEUs2nFjiRkMU34m4II+t67fL26AudKqkosYt50wx++zs7IPD+KY23vf+cDnLRndVzluMIaMgb5
TRgzk/yf7voED7oSW5pl4G6Pt/eok/kcWm8QIEhF++7FiDQHcvHSmVvX+72ueew9IrJXOSgL/A1u
LTnDgiTPCDXWBXTmZxMmGLoJiPWwMZb8nbl+9SjWz5C3N+2FGqnnJVcWJ7BrzimzoDZnYbryBAHN
xrSB7Ti+WGgvRm8tG5oWeg0BUPgh8+3nBlN374Kk+L/i6qtmLVvE8+cv/zDKW3VyCy0pxKPgweet
qsVzaYE1nAzAMdqRuJbjbMZ/Ju0Gc3eGV/XGEGPoaabYUkN8wG1/FA4ebVE/1YM9xAUH5M+YYA4f
eexKF2A3pEt7FD6TEu8n5QoNtShFLLxQS/Rn9jHH+Txq8IyWIPjFcIB+v1s93x4zBWDMAx/Bb8xE
uN7cpv/5KUI5Us3c0vlK3c1PNF6QFSoZDshLw2D6hnaUoj6G479snyl8Dt+QFKrxz/7XLX71CHxv
SYjYsDjHL+k88M02uSQ/DGmwd+rDH3nZGvaylI7eYBLlt+EBVVX06YdYiQpHMtsgP4NrImr4ckmz
hmcRnzO6tZN/t51UkScEuxMFrCd4UeNW3IrfAU3HTbg5NUqN873ZYZAe3VcrKsTRqAG1OMg0dP06
k1p8szZa1SOik+sllxDMwJMYwgUOZ+Fx6tarOv0JGTdHh3WiKJj810TGwE9jehRVTB/gzyyw42S/
9MWZwXE8vFZj0qqIP0y5/WVLHENRFKhYqNlA+LPGiwuUxiqIiRS6kLXfYXZAT10/9tRhT1J0WLR/
u5spkNcORsWKBIi6Mjjm8CmiUJ4uWX6Chpd2Y1zPel/sntNJJAyTB0oLnqXKbwHuR1h/xi6o7brH
AaIpoeDfi3cvP7jx9dtTpObVZSYGu2yL+2pv0PF5NV6KOEsG4dBVIT9BX3USjCoO0oeSNrkhQf3f
Q9BlfTUOlYMezUgOkXf2lv6rLxSRlD+n904gSXBhA+sTzGc+JCNRozehqLqykEtlWCJRxx+Yzx+P
WHUvLcX+9zxMQ6/VPhBxk21AMH2LSFY/wWSW/QaGqppw7R3We3yyv2uaPe7FQhgdwe4zJkg3d8UB
2hcqCRtjo8VNOLXTSb67YK3sSaOQLRzboo6p/CRZdVon+kpTFYJ1YPMi+/6xLEj26TZRxvWY3qVS
AXnay32G/S5SFAfHIQ9bq9OX38RnlY8a8nX7hxtX202ka2r/gDH8pyX/QbbS/Y6YvEASgDxihDFr
TieWVxVMOEDwHjmKa1sexQiLmW3nEWvGXNK18cdJPjIxfehb5l8FUnKDDU0Ba9zUzIfVUo2T28Ul
FqUYPM7hi+Nifa7EX/8wciRiBtI4CerAKKUXdY/fPhztR2woY1VfOgI6JQQJZQ8D1pwSGxjRkUXO
3ZRTjsQog7L3O26+ZZemiOVGIw/nnGokeLtYBDUggJIIHq+UexR8WSwk0trdsCdcap74TIDe2BLC
Oheef/QbrEwn2+KJjipmO4bry9xfB7XlMe199br2CNZ08oWlmSZc057ndaaYsYPa2qLfC7Vtc8cK
y2Jo02TJykTq23ev6c3P+fZRMSP7agZVeN4hzckNhZHK7Bwu4aYRsuFMLsXwMU4zHi588ELTP0pp
9zb+UvM1VtlhlRTgL/4ATsCOD0sRp8xhVSYlJAw7wGqrRskoWsqxcrpOw59KIwekgScabZQWoBgV
/89COIvujH+K3Sd/K4IjeeO5WTi9ERhPhsGWlIceWPGGghzYUOk9joJvhFpdRNmAFX6NCQHx2pga
RX/mC1SZq+TYjhI6jRf/8lK4C5lFr0S2WafP2lVK8lXvidhCmnfxsKUtf33nmRSGDLjvftft7KnE
a/rfneyEi8RrtsOC/hBEStvTl82FEL1zge2AAVxTnefV0HX79e/If+HhC5/1JoPJHdzW5/gyG5nz
NVj/S2VxHTInK9VmslS4v9NmghQ3azDo/C7DkeniG/GmSLzN3pXyIy4TdnL28vUnPZEnss3RjOGq
/LD8O3EWhRb4YJGCskXQKI9cugafUsIJBpNLPDhbftpkx9jcxMFRMb5ADLbhs1BG0OPZ71GFatW3
pYmmOoa3k3q2XLpo0oMtmV2fe6Gz0coW1Si4osZjZ1H6HZKp+EuC6qKuHiD0yErT+KC1PX8xgfRl
cips0isCLNKWFCalA5QU0qecIWhj3pQk1jVCkrvWivUnJoVCKih2R+W393xzDsQgEHUzytG3ZlhX
syJTAeDXDeL7xq8H6uCf/oaMocaSU+b9RKrFv/IuvBV5UfrQq/Zcj4AtwOxev3wm4TLx4k18du/u
zeVdcd4y1w3D1a5rmA4YAnL2zuY9S5I6zXuc2nJZccvNBeVUpnkspmAz879HFvtcR0bddFWGgDs+
0HEPPYrcYSVSnS/79notqNTjS1kBkzYYfQijLLgV7cYVLVsNnaRRHBetEivHKKLMnyOGS+AbUUtx
SfmElJdf3+Wjenc/jmv1CY3LZyrWO39IG4QpHZsyapDzsvflrlBJPhTI1qPm/CvSc8TAz2z731ry
vAx75akRsgseMqNS0/FtKbSt1O20xd5+RF59N6DKmvgQTI4e4Ym21d3+1B8bah/ImvWohD/Oxz9l
v6+IDpM8KCck2xNQy1byO4upw7Uqzmxn+3wj/b3DO1wQQ6nWahgtV5x/sG8vFgjNQsYWeQJMBwmx
4Vi8Rrzot8EH0QU+akFq8E8uEZfUwNXaPj/rP2N4kWwx7cn5DI1o+0MuSk5JPllXKu4hMntL1mpt
HXZ05xwcMUA6AdvZCGRoNRdes3T+BSFueNhw6s6ZcDBKB4txDPG1sRiO0zX7q3OQqreFnPj0DnUZ
TUNH4EAsCqCYmypBYWXA4V0Ip1onvGh9JuBkQG4XK0E4fQ/OZV1iT2qtSkAdTBmwI6D4t+93gSp2
oufpeZM/rKWF0emTcZcDPL2WNGEoYifmBMD6JUqSbXlQFEq8B3GG1FnGQ4mWNesR4uyQ+Kbs5mZ6
kkZsenvrGCJxBkONSCXYPaOqJM7WL+yse4BmqeGJE/PC/UMCbway0EBtVKWMzFWtj8MGdXrYU0Tr
B1PXc3GBugvSWVUAIrQOuQeuXsFobJ17TjqAB8pBDMThBtojpOcRr2gYrRhebAAUmNb+NX0EYQqv
L6V/TtaR7+KZXELiplzw8w6kgVddj9qmctHIIExiSUDPAF2rDMD/U3vmRhKnk/PwO/+oDvJEKhlJ
CAivCQ8wAMhafTuDUQbrivOm8CCp86D9qYKDi1oi/+a45YrIQNUKQNlOYClnT0qxPdmnaZeOxgR0
zKaLOcDlb2VnMriCont74OvVFi/VF2ybP+5O8lwb7WwatHjdO1z1y53B06WGUe5cfWEQAjQaiSxF
s+F8fvGVlOSo2pggX4dpHUVKtiAbcDLU2k7z2ss/SNUiR32kIs5PypGHHqC68scAlVBCH/pstR9J
uA30vw71maBBluuFfikr7O7OZ6trvAyEqVx2q1otw9ccnssC3Ak3f32PVagq0N1/UNsaetJ6geGC
cnld6NAwDgz/LtfpA3RG/N7WORJuQLPAcKtcU5SrcgQecHhOjXyJFUP7KHLVPDdfPYesRgvrI2Gt
gv38Ew2A5ts2RGSqqSnUI6jtp7+tgZCKZGk1kcmil29AQMr6gYlIo2jAEzykajVtG/eOY5HFyl4e
Ib0VxuRrpO3s4+khYDj3NeoAf9J2IcYNV6v6QaBVYpZGH5Ce78yIt0p1QIRPgo63KT+8tz4WHGEK
xPRmnpPXhBVtzf7LncCdj8dpDrn1H9Ik4pfKQYDCEkW8XoQg8UvKr5+HaDCL2r8Af5yUbIVyKbUd
UoIyU0972ISGORNFMIYNoFqKwEdWLligPgkkn29Pgf6jZ731+xfGLZn7YOCHZnd4NH7nU/yJG9KI
6dflvMSIeB/qt7k7m+GEj4JXY96t4XPRf9WEeWcSxw7rZatDTsOhwU8W6vNtEIgVohrcfN/0g3AG
Eb1x0jj0FUEnMbQq3KseW0v+SnTpZUjOi275k9Tpn3O3Me8NYMBZXSMVwwuZqIoN7Npdp38emCCO
KYQ0IXYZZczAu1GOjeyYGv1yJkf2Yb600yYzElDhF8gDd2dAPIWjkQ4GM9pYkuZwS7sxLautm4Rz
k9BazevBXFJnSkTmYS4wsrHIkat8HrPFsTKqixNwwCTOlK9Ak4waAvhwEveoQ+I6CMKMfEnM53Oz
On61W7e2jXWHxqq39lZssSBMf9WF/7dNIWRm5c7QmA5SEbb5T59LNA5+7/Bs23hL3xcqhVZsggaW
XXjk5AcjrXnHGMf5doUk/RYy6CgQ+glSIZCAGJTPFtp+TgL61ewLH0/p0I2cMBn11ZVKMYmfy42l
lLfSPbSy6RWPKNfwl91wSOflncAWK1s1ML+6GgGGCC3rnPWIPlP2d/wa9aSiOpHRVJgkMnP7Zpxb
mVX84Cp8fqsMVr3DknQvXA1Zlso2avkqL5drl17JfHqhq4XWXzGxWvRPLCb2DIkanSLgwH4mMSlq
KSSrffBcQ+O5ODFvgETDczWEVYHh8bvNkv3bP4RtcFwdY4LphCZfclCs6h64P6hwLRfVEp+L89Jo
rSmG1TH90l06bAbosciPw+6HJE4HjXmOgwmDz/QCuQz6rzRjTy8n0dgg6mrHhHzepPG3/odxq55L
aM7w5jCmKYG2xU71PYmmsrGpNf5tQf1x5BhfWh3dZ/3llJXbbe3YKKG83zrIp8LLYk8IKOB7GvHk
CUhYX3mTcbkHCoxlKXfoi3k3ylFo3HvlSUJYfeNztZeUpIfI4hFRdyeDRnHpk6fS57y95f5KT/77
SDKSw86mCamVbct1Zzsnzv5yDkPxEdiYyyLTkc2YfNSQCcZj9LHUHCpwI4nrR8Sg81rDN3QIRUB6
7vZkjKWkB2pHj+6rctSQuoRq23Br7PWoaKz//QXqTZZpE1nWQeNA3QFSmY0r9he45DPR+Q1ibRpR
0/VVw5aM86Za7RdYSjAmQZZmGa9Ifrs294eRRRpRpF7M+NXPJQ4rVx5/pWM1ssQ4/rcf34Wn55hA
VxMinzlkAarYrkVS5uJNFoYkh75FH0o7CSkiA+9OY1Elk9isH6S3bAAWl9xM43hGnTfFNO937egv
8SSHPYjBn/0fuvHFBTNJLu39tDF5QegvLeT6kDPvk/YAq23MSgAC3SuCpTxt44maJTdN5z0QZykP
gAO9yxe0SS9W5m/6Tfcjuw2RKvquhX9uUeqyiEf/qWYAEO1qq6nPrvyrMX0GeQwX/L6B8j/LQGAD
wV2lzH4TriJMi74erwDQgL/47zLJT4Co5X7ZBBDbBb9GLQyvgfp7MZTZT3i8B/MA3PhFGRsHG/Fk
dYT4TqR6jaV4YIr3LCzLKTojAsJDXhzpzLyd8l+CLP8mPvm4FH6ZqLp+7AFpuxlaJYMYYz1lmLvW
pnbeWrJqBTJ3Ml4c0eoCgmqDfXmcEMqFV+XqGQhZXkk3JTGzQbpwO5r/bcEh5hqD6FeTHQ/DPZB3
sAKc+CdF3wYV/dU3DaZhjk7+J2mlHZlq/Yzw498kUJ2o2mcrUoltzJvBZ1AfVp7d2xIZH0sXTX+U
FV0DKnw81XsYQqflcyntQ8s66Mb9G33OWfwhEO7e5CwyGX1Tl+OdpJ68e3CnJo0EdeXpF4VioKGt
gBvO/fpxC/Syj+0QFjkwWhjew0P7NuqAE5BrnXJ6LfSBKV7n+aToH4LW8umNi6NHJRQc+8Rtt6sa
m7rZoh7gFGn2cpa2dEkX3EWqW36dJuAU8QYhotOPgS5hiOJWflhemnJUQMDh5bQAOuJnlRbmXC/T
Pq45TKOkJuq+zJVNVJ8xKp83rTBtN6fvMtKDUUWAD+uLIyOAKlvoWjPxUFiBlE2zK9+EqrZs0GGw
naPrpn4AoGH0r5m4q1G6k17OlLKT8leS09Urc9e+koFPhR664ngFErB6OGQpLUDWXsLHVjDQHU/s
3NFj4TLWeFuDU5iTFUd6FrJIBKEXODnFdi6fweKewQgl5oX2KYUUNUC1XZg1i20sUU5tuQdRDdls
2uaPBoeeaLbBzOHBe4wSRTdHaNIOZKT6mqBNxZv+C4TAmQWeCKrFWX/PXSL4TDhdAygKd2MQdFho
LkknTJjtQh9JdFiqHsmCIesc7QrZiTX+kjDHmzyNtukU8uZsjbhBDQu7A95hkVyY+5UUl2lzBTtl
FMCsYb7iFWMPf3UDeybWzvGF06AC4Y70EHonSVYLQY9oT/LoElIJ8jULwvLdRGs0MK30vvxy8nLg
T6B1ybINyJLZaZInTR4kwYAukWLeMigM8b8zml0O86Oj+lPKYpyJ2PAdbyGfbb9WYCtI2NB5wpsl
D3PKHyrLAnbyJXP4DvWJORhF3osqJgwgkLP5kLhMuI/3OtkXb61eHUzjxeKpjH+tAB3xrrlSqdqn
f4Vdkn+wLEQc8WCrGEbSgLo9TadjTNLDiW/q/8spmSt8BwyanCfEQ2ZQIaSh+4YgWCahLYzCmzJQ
yb0HAVMKhNKx8g5+G4sq0doOulvGCJINBpFexY6wiPp/m8tFyTN+6tqGHBR8/jp+z18EspryMzUt
x5I6jp/BXmNvzUwaFiWvpVboud/w0aIwemjEdId3YxVYVHNk3t+018U6CSRZSWNe1Slyr7qUsoiY
QJmeEZz4CqWaD56MigNg8f6+qbTDLL50Cn12y4N4NEds+Oz1aCqgznBOBnrgBbwVvRLzMB5WSSkV
LZi4nY7vUm9ylryIKnwAhya+UUK6y8CNrJu8qu7yMuaCm6r8JulkkOtq1JWDD+W4SIwYHZCNO3EJ
ymHKQZ41dH+jpZSem/8t1Vy2eegIXhgApunbQkVGX2WzWF84NBS6w+whJXWgyge6/7ufMIxa2+Uc
eXRFZXJ7jKg7HQNSRoHL/KtUj9ifTREuzyx1UX68ingkWfrT/knrKad8+Sd5MUC4jMGK6VxInyly
FvNakAOHMj//dKEwwrlxo0YcOBk9iWsLtxdises/UwiI+EsbMCPMuKHPEJEgmL+46Sg/BMwaBG2Y
ItC1YHsRXgq6i+pYFRoAJSwM7yNu7yu4DufdLGiKzxspMK68gx+CkwZz56cfC0u4nM3gGZyaWga/
CzzEJfU6AGK4F3v4l35eGyMJtNCocvBW/OaNjapQQ/v5woryEINgSZKhcST6MeOjddT1UmRqpHGQ
I99nAFylgdKFFCHf7sjH5slR67s91o0CVdlh7WO5wVseZCAJ2bdwPobIAVqf4foqUIn3m+JOCckj
g5HN81imh58kJcySss8/3Cp+F5hlFi7BFiAYYpEI/tKpQ5i+pGDzcagD/AswxqokqrsTZyLZeiKE
+l8oy+KBc0Vq71eqOOxD78GrynPv44kFkSa+dsgFr1ZB1EP866i3hkGuJwEQjkQNnonaUhQuLPU+
IYWHDdGP4spgNQSRidK1o49MhVY+s0eZZcs3ApSOdGZ5/sxq7QjB5Dr6RifAna2jgliVvDxDjb3z
jwLI/WU2NtuqjpOOJ3BWfdEKZYupwZvUno1HsabUgj30n3EjGq5q0tP9IDry8Jlhc7RqKCwfce25
qMEXPtSCvO3bL633tRf7boB5/DdyW33YydfIA1M+4ZM64+gTvBZeNoMOWZzNKrWjBDiim1uxvo5H
wBFFGncwdnFQoh0YLEblpTdOfW5AoyiD8qNRK0S/TkOFgZHuNu4yiYt7dvw7z1N+aDB0EXJCwHzZ
aFKWNSh4kpoyf640QIERK/2zrcsEVwTj4pxNb85KuODgK56SkGqTCON5JLO8DgREb3lyiHzSxRX/
qGIEMPPf0kSh+bfk420mo65x6sRwwLt/+itrnmcY0UYlrulf4MYJSzjNNAg4IMxF7sVXXdCv6MW2
/MEjC8XRMNfkNjF1BGlSMDmbeppvas2o0GJ9Pmgkpdr/TRmq+9IJAAcGnyNjc2xWUZJTZeTbJO6S
aE+QuQiQAOFJqeD5tRyHw02AxWCs8tDUog2v08dJh29mlIFzqsNyk5M9LC5L7lLeqjiCer+WGeJO
bJkmFh/Wvu6kmM/ppUHe/znSMpVgxKqWIvzfYVKbvYewNilrXJVjVM/X11zeNAfjdiVBAnj6bYQ+
gslRMBd6EFDKnMLoaEUos5/DchakIujXuU3AwiStp5qeoSKhuaeWzDpdt9Z4klimK/XRw46ha9zS
RykRljvevxpX0MI6g0To9AWpL8LanB/mDlqvY+UopPcFhWbQY85msgdqNAt24XdJyMzw97RjIePI
X6CgIvGdJzDlEuaSzfEfo5AYoUzY/rxXH1kv6RQ9iFhYYzZnebH9E0bscMgoTdj0OuZFFkG2Uylr
nxNKT9B5sms0gdKQ+gIS/6ciUo9TG35fb1hts8JSxJf7qzvejWUx+B3oDnO3aqgwkSyUW8zM9T1z
12EQ2wHP2/BCVej9uBp6KvrovrbxVg2i6nfobp8/uE16ZkrJrYyj3f0rJFskCQW/hVyaplKLVBkn
rrr7MuzmWbi4/rykZZQwaNtlVQ0ljpqWbkDXQSim4rJkaZqdZ8ipjaG5NqBqXlWXn3M4rE5atEfx
N5R5z9Fb+wTlPfGA1jdRTuM7rOM383hJkt42trrZxvSCq6Vtal+284kJfW3jMPXP/+8sVKznihNX
dQlRehIzqsiBk2OK3ZDLMibpIBTo+WZ3c4YulWSu3mcr5PJ8m2i/3rPSJeuBZnOGJooxyKBy9BKG
lSr0CJU4hIjzs7x0JBy1SFll6O4Z30xjbNOFJFi8TQyTQooLr7xrh5Pxzv5INiRTHd9QHQeG7Zcq
P3gVfqUauL/zwwddp2v0VpaHatsYRs9pZFjK1XBcN4NjbA6O9sTN0XblTvDU2Qz3Xj4ftqWNkUSQ
qZHLiV5tEP+k7nGefZKHhI5Z8hDLOYrTolgJgmwgTkX0coEMNDnG25vweLI1OthiugjM4LxE4GcD
XxwuAjtHMZSZQvtrnGR/Rc5Kby68CNmyTZ1w12xODLvrof3/8z8QHXY1LeUVY7TTYe/aIPMn21/w
7faWL4M66f1PU97hGhPHDJ/r9UI6HBuVoHiFMBo5g/FxarWHlr1Ko6Z0kj+n29OHwqq4uVaB4ih+
zEwmCK8zPycednQrOTsz/4YGMTBR4LgxzWNvgRIsqpKjCto8PcKFMYGic9K35giiInbhNbNCTf23
dr1L2GM1Up51jDtGLozfMtjHAmcyigQURbK5pW8VUU8GHs+a+hPhNmGpOVwIj3Wb7nWG3YIyuwPX
+xmStsAx2j202IGjEfbbIDKjZWIjiqDe82jJtCZ63X9kZYO8Nrk1b1v42N8ADwpZkt4frTloar+2
3ZD1XOFyy0AxaWKjRyGNR7q793mcTy8xsFU//Af2wlMVLWfgFYXnSmm01PiuADWsl/pWf9k2nc4b
2nhuCzWLyl2vtCl8V1GpyrGVg60Lre1XAJg7iVBv1iFi93bYpfH9AZFyIFKncxEyHi1M5GJkunKh
uKjFakE0Yo5JaCuD2SPx/XCBsdYYo32KrWmzxFGHb3P65+yDwi4s/a6SE1PTOG5VoVBJrKqQllF1
QvqDKFpla1UaOyWtEvHkjd9sbJ+gSADeqTDCQFi9Qwa9EA6EcWsmcg1gSrQoCxOcmKe290Oj6PMY
BXig6ogREYv30rFyIW2oDd0pyFORukmJsY/2jbiIgYucQ4z0d4YiJh/nHkvb2ytttyVrjgiSKA/X
Lr7O/D8UTAtY/fpJmVq6JDRJ8XaqxtkJppiTYSJNFQIas5XKmHDblIxo7SgCxPCbSDsoqQdKXhfc
y5AtLL/MHiCFRPW6q6qd0AoS1TRN/h+7T3IqqdrJ5M4Z+gEreE4q0S+0ADCsTjtYAXSR9+2UcFur
o3n5BSKOK4mHbzIXBSv1hHjCUnJynPu2WJ+86aKPP78RaX99a5VMGrXVzDad2ZlE/lgDUYU3B2/f
KGVW52P5NyPNv7TTPLfi9f9Eip48aM1BvE5dfrkbJueCgwEjHnyB3LnEEIdsM5n0qH0oIdLbcCfO
yUGCqjTSoZHX7X7GHo7CtDInui7go7wlHwzuDn5vkrcvGK5zIyqUvv5Sm0axzQ6v6DMJpAI2g8k0
8KzjrtJcmZu8zNSupcxbBpWtjU8Lbt9dar946GelxeDe7EXJ/f2r6IuLF3e/2w162RdKvhTrSwQN
EjtG3bhv9hZRPcwO/p9rRfwYfcDFD4IRIYhJkS54x5UlxOQf864bZItOxituU4oMoHPENTqrtyg1
nrowL/oFKzf4bi37Y8UvkLrOFmD/bjz7P1jfSUXZXumPWZWTUa8pCXQbElJp7xYPTLYK9J3C/aBe
1KNlKXiyAxzWcMPpSTjf/QzXTHjwoPtZqPaMF4SHe/LHs46XrQTzp0QVCUdbWyAy4JPQ36rolVFS
ylSFPz2MIXWMTT0cN5xQeSyl9oO9Z8But3uKleA5YPwB3v47I+KYkpT0srHvtEXoabnMQbxXhOlx
BgAvWpMngS2nIxxd9ctG2/e/V8ZCFDJL25wKb4otGwdCBu72tFQpYd/o7ovEIM5lEB2g94eX0Ye5
BkJOs3Vc4HPpVe/NJ73pyajEmKSp5eL9HAivIjT62sZtvQYdtNtZinQJ8ILEvRaswja575gBdZyp
dqlwwjM4zD1Zf6xD9KgJ6KJW4SP/EBSL7OP+9e9twrYRV99no9BS9ps9qHwcet8fcTJU6DpL8/1e
8dvC4/YSsVKw3KkcMgWZp4kw86YWBJS7NlANf4tZmvnHYiJ82xZDgMqFQ9msJjfp72PzULWqf7iz
HKSb5PSY+mVjp0c+GxMl1wKDIXlPV5bjZO3HxHIloKESpjGbdPG+Lc+kwojVVe155eTn9+EhkDJe
wBTOLjXMxUdMoUfsKmNptevaoA86elsuAOUR9eUSuUhl1zrri1SQmceqJzbE2wBnYEBpnIi8LcTC
wTAYbjpmbQuB4ZdmLsOJmUgIEVdwkbi4SFMA/5pUZv5fssiyw/CN6G+WmS7Tk+Xgfjy2FOooCWLA
R/FYrMyIq1DaaB3KnZNMftVb2BYvZHJZurgGPgftTHaQ4l7D7EfqVZXe+3xM/sAW8t1FAziqh7s+
wc8XVJ/swaQWrrGKZNdxQaBV/vuk1LINo8io9hDUJ6tsQVE5KWPk6utfJ6HQfr23MtMXsyIaHRkW
y8VjUYrWKzmaqZlZST86OhBbpwBeh2kpeHm9TnIumo1bEJx7bz2AF4o7B4aT+gXjWohmdbaqvlIv
37PR2yiHLhRtDCks4NAY+7/TzFqebc+TfSeY8e11gCgemVLOBij3DTlB7//HF0eXVVVMTEh7RloC
JnCAh5tf3j0SQKi2CcFZc+PWpR5fNmJruYvxJzxPpirf5qtnG258iDaCb00btxXGXkLhY/643daJ
8qvgetpBNNpPdxHYTT/iU5CpUe+hSPFJTDWS0ynHxUVFCJwjzarmhuD9n+CgfRR3cpBc7Qqn2SOL
nx/+x1Hw+tWQWSh7vLDL3/nF+XGb3ewjPKGQSeeNqmIeRDvjTSCDsgHJqRaSqsuN09mB4cM1C4Ig
gqEqpj0aju3v3KJvRilv1GeoYR89TmF/j6yFhBhLP9SP6B9c5hgyrKDojb4RTvMG779awrqB/GLZ
Ykmt8C3cVoXPBMTK4RpoofGN1U8aRHWkrvBhh7bc2AlQ9gndQ8ZKg3JNOmnUavKtTDJDXAr5M1Pf
u+7HQVGUV1yOWbcgDyzZiLjne0pn5HprLU6JJrVV/FMSHFd6zQkw2L3rpQTKnWaHcWr5ud3+t+pc
ivZLImeeWX1prdpJ17bgeV5gxUiykTeA2y+XGRRjBrEzjUFbbqjHk539yjUsVyQGj0o+wFsw05IJ
oQIiVjHeW+SzZD2p8Mn8j983qxne2yYehnS8fzCCLRyc3pJYK8jORPifd+HeFVFRAX8Eqr8/ry0g
kD1RTTRRUBoxxedXFSWEb9q5fJRB1K6ShZ4HztyuU+Ar6b9qNdtzBou5/6CWpheOp7ujDsAP+Gcd
f1/8FtefMDbeXMVko3UMDrlNnLgIr3n6pJL/69lGew6zxA82ssN+ISbecFqfYQaeAujhxH2XZGnG
OgYH0Sp9jcQihfhMDYvZ+DEJcCW/zCMtj1UaIpbrBaFcjohkzH0ouHGsawn8sx9J+v9bb5t0xcxw
296grRuloTB7eFtr9bZ7Npd4cJXnDamCjV2/zwSDLw1PpCmvRzvoDjZ8hE3mRvp/2tlmFxc4D26g
ZBAznNHdxEAxnWVIgISmYUPa8rWFM+LgdHQ3/fQEHlo18exk5s1C6si71EGinibrz68Ix71Cumx+
WZpUJJpwJ9CS/j0uJN+GKPW+Gv5WXlBiAKriyrRLbN1cTRsBiWxBuS6t8W+Lej/LEtvjSO02HRTB
j3lEBQQFx3BMivIIO6JnaleoE2Pu9uoCR+kMjAyXxYMx5nZX2D2RAT67fT0vYxXR1L+YRxdW2wkK
V2yFOp+HlPjz0fcy3H2Saaozg6/96F2bDz3uvaFZ/FeIchETEMHMKfnmYXwZJnAM2diqF0apgR+T
pTBwfqDf1EOCR368pA+rLERhmzEApxzTGDYSRSMYGkLUCLvR441PARggOunksyyS0hCSN9yBe2Px
NJSlJXiBnDQHlXkzZ8HIKhiFE8h0CoUTVOXPevlVCWzaDe8EobpSa92t+gQkZFptjjNR6Mec11CK
ctvRghGnElLgAsn7iaMB6N8aE6zrcbOoM2D/oDJTReewPA4uKjOeW+ayOQQE2+UEcbckG81HaY6E
9rrh4+SntYoHbBAs7djcpWKUD63Mr1W56IplbIBqZ87/eeFZRU/zSaFn9aC6fC22ibORyPownc1l
bhBPMgJ56E0D6u8FKprSSnOsTs9FP+x0FU3lJNEF9NQDW4ohKOs0fE6Gi6oBCURWSTUZnaPmIJbT
7PXuJOABtMF5lfkbWkrMCp/edBsaiXmPDxyey6QcQSB/Aftuh7oxsYRQAIlKnPaz8+ykMLT0mpQa
Wz4qVj7Vc/VjvvatO1Xqqn/tmCUjbndV9m9uot0jbAl+sCMppLoHi2Tl9YQ0KM6SSb6s8KQprZD+
qic94JMBrDiINLAFjiMNdL7jtR4R0F2F/1u0UQ18x3Yett16FcjluLtPhV3m8JMRGrx9eXXVsHXD
Khuuc5R79h1ZgqJK5VVGqmIuLzCsBL4fZY9slN98tNvYFuN3dEFwc2DU//6eF8yixSZKaoNpuve9
to1DQJ+nUEik1MvS1jZQdaPBnh7VbxipY/cHhoNovN2D8rVHr7oDnW3ie6iNlr5XNy23ohSsDUsn
P/I8nksknKsUuWj3iRRXGBGeXUGfENp4Y519jYaniOoDLqT9gXfIwNTCpGNwiXhqCKYNTTQ3r6+1
+pM+VXSgehEzNmr85YP8NpJaehn0XnE2jeIF8e7ftTjbgX0M3RfAnC6ZzcNg4+9r9IF/+iQ6HWPp
ldDGbFomuykwBYl0ZPRx0fYpeZ28iT3mir6VuTpyYVUJytTZUneNquw0/Tnyu7LaoWQZH/8Dge0Z
Tn0hQ16W70BdtLnLLuf0Ved21mjz7ekMqYcoTlWE/f0QorfQxl9tnx1EsuWVp9ul9AMIkjmdqT/8
1fy/2aplrLj5b2VnCjXThcmZjaxpq7W1ajxC0NYyWGV5FIlRjl6N8MF2O7JxV4kXHX7L21n5rgmM
Yj9oc+8N5I3nz4AjrD+dRvdgHJJFkFlZObY6bLXs8XlZjnFgT8b2aDophSF8AkbiLIu1cq8vwzQC
mzyXIpCQAzHcy3TpbbsCgdK+vez5gAeIc9DMtiIT13Q6HdRI6tCutgL3LNagsI98Ph7CIVGjg0BN
U51Axzcj2XNlwg1LNoz+FOCC54aPHIX+gHxrjgp2rajmVlZbIY/cQ/MSddMLjyGcaEI1yL1KNrfO
iJtwy9OgS7hfbsm2iIuv24FYlu0iWr5h6oIGJSx/Z1w420sT7EIhCOL/4GL52/x0Xl7nHkovR+sY
lkJ7OvOo4HI9zO+PBth6z5p21qCTfV2Jcv7qX+QNEZ4CmCOG6j6F+lCEJ2Q4sHLxlh+eELf1MVyN
TN7hJKSKJNwbsI8bqq9cwCqaH+Mjl37IbIqULtytg8DGM3wvLjbST71aKNQ6r49jP/1Obvx/hISY
3ZFR6pIHl+4m6VgCNLcBgJbr7p/P8nEtMtRLl+LqLuaVAEvk7/TMtQWABT7Q4ZDZA4lUhvgZEcnD
UknUbxfQqmXfL4Y417K7pmERRG/tKRoxSuoswFuWcDagp8X2kb5bebF8OC7jiz2eEHSHjiUqPIId
vqQFf9yiLd+F0w1tCfFqmgU1t1m7uKNgi7i4BddmfNENMO2Skq4RN0TQ0siFL5fe6LMxLmOAtekY
5XefdTjkmx0EI+xxO1COubaRSl3yRjIafwU4e+/sNkF5o0P10XH2VRhFjwUQD6G4HaljQS8u1deU
qvf/92eI8yvaYjVlyqUteHAKYUvFNCkwGRvb4Ec9FabIPbdVOKCaRQBOCfBmB8Xe8zbBqjYBYzkK
34Yu8zaQeOT9aR1djRB7zo/WBwpZWSf5JalWwryZ6Vn+U3xNe7iW6D4kgwN4xAYquU2Tz9agxx06
V9pAw7L17+imu0cOqtqAEWPrFmpVT5YcYP6/FtUV15vXqZygV0KvW3S/+892og+H3GxbHJxLKFuD
Vse/J4nZi/+hfAaZURW5U1DC8w0qBI5prS/dRbt6DHJu+XFxKtPSgK0+1CA7EufwV7/FO6XwKVjl
mv9OJZUwjmX2TMr4j+9btu8H7HpBiOB4+ZQDEL1O1vVDTtcU9tBYQxEoWsYgEWjWIqysHzhirbzt
OosGpXEhZHabhRZ0HqYL0XnE6XsqOUSDH0AIE3S+y//NszsOf/kgkXZkyv8C+amEhJ9zjADHgPUW
ccDdvZYURfM7XZKccCOqSjxBARIlCkp2as3j9grRMJCI9UmqTFpMy5knx0eTFlzuyzK1/4bRpE09
+zR7RVEBcXVCoL+Q7O4pEjTKcw0Q0XbWimurFFbkcPm+D+ADBQ/0aGalSPl0dHPjXILCIM3G0bC3
QjC/AU1RLhmfzfbXXZ74iWrncXo/8/3CiXZOFuhve6m9IWYE0YObVtfv0gvQBUufK05N6hjgEbft
foyZ+jlgOWS0FuCV/BBLlJ8Mw+mwpgIXi82aKEUqaG1HEtMdwKu0HrcbGO8geee2PyH2/lZ1W+Bp
00j8rcLdv3dXUBygkuKR5LXCefICyo5hBZfoPCgGLyHyq55B4f0lTuexNLChYOKoPJvnhN2Jc/Vx
1xnTofpqXm97R+n0lFrXlVUc57pCNqxMvnVSrwApCbVprj1qdNUCgY304PPM6ow8Fum4cgla8IB1
yyx+3d0SDv6T1LZygtNtYVSV4pNthfYjQtFX8kb8NmidZ712pBf0QE6gtX87OrKHSPA9eI3++s7p
wPXZGra1iYm6fOQx3BImHrT4hYe/Ci2WTScrF27SaPCSNGI+RtOLhu+MCYqsiuTE3MpnuT/YU/H1
aIi44KTF/xh44k4zxD/1Tw2sYYSUM5UVI23XzWzhbq3iLpNwQpqJk25mCd0j775psBidj/lulc0l
vdYinxEegjQnp7Nnfv3HT2YCu3E7Uh3cIRJKX2sWsn+I4dPd7ZeCRktEsQWlaxWr8NxHC/lIYmon
2/wVinhxlBGj2bXWdmdYVtcexmbtJA4WLSzc1YGJl9v2nDqQSdvhyJP+BbYZFoochsGGlrkhE6Cq
qggDTSqHwd/i2gjx7id3ac3wjG/BoXwFP2eZ92CJ/eBs0pAaYEsRynDc8bYcZc/1PiFBC3q2F+fj
AUaGKc3lXt9gxXhyoYnqMhmi8KTDf0jiCXUo0xL40FIqi9UkjathmE0LbJ0qtpR1n53nuF7qEXEL
r/zyfGZYmOQLZi7WqWF6zobYxpmVGO8Z+nJdVliOYC7F5FvTE6djjC5cMzaq0zMdf7V1Qgn2cI+H
lPQsmQfp8wAktDTRO2z9R5edTL23rVuU/YdDtqN3qepP/6RogBSEnjGrtymqOLnBKNzKPFNZsOS2
YMosiGh7Kq52GRvMLFglqMwAzjZEw13k+Zl1q0IvwePcq84JKME1BKUbcWz9ecnfu1tYGt1S0rVw
YeD1rObglV0wyrFWl/EL4SyStaEtmOhvMJRX9pOKL6b8nhKeop98jwBOj2pcWNZOE7Dt+xagtKmm
+mXUrMNkDRvJRwibsMS/mDTpxcSIcwhT8d4GumGwi3uz1Gs1RODeShQUKYWjXi9bEb6p50RFjHuE
GdDGvU+25XoMvDwhJexXabBJgo48F4+Cw6dOSOGjT+zMsF2qM8URGJwbhdz2RaZJy4UC7SAcHYbY
bvHPalWkMhQEYUP2NVdM922/AfhlLX2RV7dkBDRAC2WANS7tKDpZ/0wW9IRg2r1AJupGt8kPwHoM
yPS+gEnD2J919VOiBdMtepMysg7qcfbb9jCtEWJri7RUmd5KUx7oOwrNQb2TkcL8cBFmZU/wYpa7
vW4yynxgJYueigzQKBjo6izIJF+4UBRvpXnbnvB4+XDuwezm9B/uWfZsS3PewR0KxVDpv6tDZNzU
l315qlCeIR7w6o4iC1YOLk1pIpkxdPRSGq+/E8dIRSEkVTr55lLnxlcDzpFnavh6QjajExVMsrNv
uYQiwYVLIVjE975w5+ZgpnqhsZdiHLyAeVprNTGNkKubgRosLy6tEShdW1Wuff3owhFoBKcMvlV/
nzGg6QEGwk2nJsC4Pdpc2mpsATA7IplIOCzRsTBwp7I9+1GJdZlE17g/f7L+XcEnTNkiEYCrpdR1
DFMbbI+juQu8jU0b7xzXDyMhKIv2cVF253797A2y4TaONfDlGqWe7glStCrRwt17f1pljdsrVLmY
x5OvSkSn4Fmfrg9gVsbbXGnyUs2Jple0rMKZddnVF0rTcQyke1tGd4DYhgTZNgc0glOluMAhTiYh
JgVMLUsmDRrKcQAQuYEmRBFTb35r2M5NlwlXZpFmJiOCa+TF8kBYWm540GHWv/Dw2nZxYj1VqIas
RrwB8Vx2O996n7mmlbZ9RcA/bhan1wR49nmJbtrePcSBlrjyiTp2vjkaGhIyQERGv6EE0rdfHHC2
h39j1BwDKyFVHd+bSXrBC1rZvDNVLjuZALRs9Q5Pd8xw5ABQFNYZ2FuSB0LiwWM3c4cerEILZnzc
2bCMgmbZz8QbEb0jLM/tvqI2Ij086Xymwf4qMgtj2lDTBTdGzaxQpciFoi5GPMlwo0mgk4XCoxYY
mwS8rLRXV1S2m5fGRJU3gg6i9H5Af1R84CaD7tpQRr8kSMRiUib2X0Q5Wf6oEX5s/KdVSUbLomUO
akK9CF8y1FI88EBhf9Dq6dq2cf7qaFKkK3T9BqOb8di76GRQn4d6b8tuM4VsRbPdBZs5J92sRrxJ
werY48imvTZpSfaTJrjctVERSl5WG0o5IWjm4OAwO745OlwEw3ZaSfjcfHjdxFupSMhKsvS7tsOX
UXD69dV4RKicOMXDvAjtZDqicGKOSaIK/rWh9B+a+t5Qqkv5hZELaV5cstp629+zJrAk/RYq0bk1
DVnTDWROTS3r02q3a/OmMW75l0h70BSpRn39yc7nQuoBF0mdCmNsWrXiyuQtAHT6uY7382u3zXNH
8eYpl5ub9b3uLogwrjBZHyFPQauaeAXIWW5Pn8Q1mOba/2nc8s0aIt9PUOLGCW1hx4BivquyfNIN
KkEeQzPLcM+FUVXrRjrnvakaxJmrO/Xql+LPLiWH4TMuO3Rygx8P1pq7yWkOHeeiuDl/qiTnBICs
K1EA0H8VMV2+SL2FCLyTubV6U/fUqy2Sn7SZIms6CbnzJo9F6oL2VgqrepLYtMJCkGkZ+a4b/i8Z
cIXne8UyXW4NAfzSFB6heQGZqNqjqbo0ZRoCaOI074bgJ8+T1E52K+8KHLcmsMDt5u+OH45vaCgX
ItRToWAwuU8l32ufjyWRInLA96M7M1kbvGmuDjSiSUoffF+U6LMxWEWtW4Ym2jwyuQd+UC6FPBsW
t/1hjJvZ798H5Tz7XIa8sZc7IL3d0aJRkGr823PUfuDmm+oT09fU1PHUKcJwww2Vp4vj5NxwOHV8
hbYOFte2lQrlU5UtOAYbWlTdxtZw/Qubqwhsgqr17Twq7bqX+VEuc/qpKTD90NuyNmKtOEtNBqem
hUXZjTFv22bBH11LVya7vDACSUlPMY14WugKGLIEEfccWafvm3i3shDGrjSKD8VRYxush+jgFn99
DEHUMp7b6QVbrRHprZmOvQU9EpvQQIMdtxN+lFBNKn0/bjFDO7DrMySIBcOzA3dMgYcnYvt9hJk1
dVCaOFSQnsaGL8pMRG3bpOV2LqJlLkKQRJNJHKlTqNIuH3rjlpiisSyneUrVqzbiS43OiB2J7vQA
QOk/uc79eS16H7P1M4L328C6ariwQUB2qATDMfLPDLiU7sVRHympfoK3oOMJkA3BZiMVsF3+Og2p
TXme3g8oPx3A2sC/DnT6MU4yd8QgpVLRX9mwQQx8+fuWnYW+Ka1nW8PCzGfh3Rh8YEIzQTzEySK3
xKC6IfryLNWlDEUCw3THcyyCN3pEaDAFbilbbGcS7BmcmFZD7VAfQNhIpLlTHzB14+BAEi/HCQAX
OkZhbQibeWS6OHXA76Q8De5hPjWNMlFQkQigdttI7N8G5DSFzLiixHZxe7qcs4gDdDMnSxLNRULK
ovwHcZqD7e0OxOKvQYzqpqFsY8s1dZRpAq74ddJhx8td7C1bdhHIpnnBbyrmdw9ZaFT8+S3hQjH1
8WOPlY2OmgzYlQ8x44U0Mrh1+YBq4r4VxQQyYxb00LPPS/Lp7YSoVFBMCYCFhkHhy4/Z9ioHYyrK
oNLRe4Ly0SrzlceJl+0kiEPJob6TJvY5gpZWSEZ2SMFZYIZgXCzd5NsNmIGX60f6TG3+m3Fi/rjK
6oSA/6FSeyT1Br6Q7KGwTjmvEWiPRu/XNlUYZ4dVlm3OiZ+cldeJu/JPfMe6NleITfcLDBkrnEbu
QL3yiseQ+l4y/moP/yT8+JnzZUlcidaVUB7e4EORqaUgxtUh6ocsdqpfcMcuOaRXuHMEYTFfO6SY
7YZwmU/eCv55RcYC2edZpPJxWxBrUUGxs0H5G+owJteCYw4dRi0ggg9qfU7PD50TQ2sJx0deKBAy
Ir7YeeAK6qYRPuEw/lf9OJIg0WvHwCOLSlUh867J6FDANIYCn6jDLLzRB4pxLdlzifphcO0+ycNs
7na2CZMD5UO8OtjP/KAMNX3cp2cBats5MfTUW7hJ1Qt1qG92/ZeINXfvpab7k0u9Mt3uufN1d3Yz
46EW7u9tWxhe2NXmbrmjiu883j0rihS832umPC9Le+NQwkHsQrCIvIOZQrgs7WyV+DPkqwbVyEms
yNYdi3BM03H1rn/TN1ypeBET3hKwvTp1q5xNRsdWwZi9et9DakELFHWeMwi9W4qpWWB+J0ePQwEF
uz6rjm9F7lUqNlsW/xfzG5qEFiYGcmD8XFgqtPgLYd5PKpkEyeU3I/nKR0aq8HHEDL3r/VLDkwTj
dWO8wrRIJ7kxuOisStfAJSWh+kEBEFEAGOgDEZXX9Tv2odRNUOZGswmJEeDp0lHmsIGNDNyP9rxz
QFOED8jW9kQL3hHbU8jE5LeQ5AXw0zda0FdzbRCjFIQrw5QZ9tzoOUUHC2iEjM93mSsSJxzxrvBy
E/amdyIqcipnmmlx3pa2jW8zWjFn5ibWcjCpp2ae5RnyXhD5JxF3S+Wz0Y1zy74lLXhJ0ok1GCf+
ElLHx07Gd5a/PfNNOZJRDYMmlfQZl9/OKIV26P3UyM2qnpDj2ILVT3yOIEPCoJRq8pe3sSKh9sYD
aIZrn35kxGH8eUtwAWA6nmCtW8DPnvOMmvSCW3IBjLAQq355jwx0fgTlz+VDALpTUNSTHbz51cWQ
zhxcwKTOTbt7KMwJWBPu7LSERHaouyIqVSXQqCpnBzUoRN1B1PrdFAkEDGyuvQ5OFjFmqWUPTCyX
JgWG4a7mfbOaqhtlM8gWw2Mz4fona6fx4kp/PcJ7PQ+vb9j7Wv80bWWgSDSVXp36PHEp5uZWwcM6
imNls6JPBNSigx0q1nAtbrVU+NtbHOPGkGaaTv3jMzldLc8RRyYZSmeexx6v/TjKjD9mNfLg/nk5
R3oK6GiGbdNd6rrMwcnqOeBB9q6gwBI5eANzZHE6KQMaFuZ+u4cqRuGlorlmpD9bvppR9Cyfvi/K
arhY5HYUBYFVI2Trzd96B04WuIodu3NAv7/aevyo8VTxe3Laa9ZETYgBAUpY2yMrxW+rbQuOBPxD
ezVBn+w6ZKxUR98yWu7zelhLof5kGD/76PutZSx6DgfHm+zeMx75whlxIyIIw8vj9N2DBLcjkNuH
NHJ7z0ywFjqLGfteufPBGrNS0ftNo/3NeXNAEporocIt3uDeBYuyMcvF2xwkhee0MxmHQMOhlVCy
QTEg8FlxtAn2sP3NUBC1o1stF6MwZOSp4yi4NUPuGfPb3t7CTXl0B7r2QToGVl0A42hiFxo4inky
P6sPizi2CZjehoTuLaP5JffWj47No3Ra4gY/qu59mQIRoHJwiv/SwYbr54XEAja1F4Wgo5Or33yL
WPrKpEdaH9/JZEvq+i/w8bwJmxrbyMGdDRkSZPWBg7T0wa5yn0Y80KwpBxZjZAmC9Z5Ezeb6f2Hc
BZsAmb4o9bG1E0KFuViR2onfkXPcK2sUiOoa5Br3n1ii4BVdSsYJnmLL94o4DajHpddSIzABeCqc
ZOXyBAWodewiSIvs+slRRIA7DqVZwzP5TnWyvruRCd94qzi2N+oLNvpjqHLbJWtCBnkgiSLnWr8Y
v1ekhp/baVgGyx18tuHNGkl0VSC1/rlB7mHN13GjUe+QPh4UlcZ/sItf5cn6jzW6RDaEjJdfUocO
ZPAJxGxO/KKEcxM3JE18nvemuXk2OS/04X3iGypgKstKtuwofjily+06xXVG20CGHNIEQC4aJhMz
JydVr7KectW3YvyAl5iUitkwjHtOwMkWU6nvliQ56Saot1Cm80XHh6GEv1u7u2vALbm/fUvhcKrb
v9vWFCABevWmqZMN8HILTHwmoTRpC7rgK6/27KNAyrNzbByBFqKlDCpTzM47cBd8VdRpEvpuaa9X
kU4yqypKWKTd1Yu5FjR3mloJrWWetJdmbK4ORvBQrV2CQV/GpeZtEo878NqkS3CUu35CvUT0WACH
TsqVxtvy/mr2PMhL25uX+fbYhhrRV22zRd/KyObsraYSuUQaVmptOsWmJC6nBZqW0+RdWNdY1urk
/SCOtleAdQRIjWEFmltsj9MbRjQkURMwguySnrZQsyqox7rVYj81vXIfwY/jtTD0kx6uHQtJT9PG
edWK7nt2cm1xOad1QdMR5RYvBUZaOBRZnwpq4KXGMs34mzYHPI9pOE6dwqIcX+XIB4vBrCM6pFFS
ieqTwxNE4cksffPb8S2XoUVF07FgYdR81U9ktGFzEx3VH158eY4t4jeY6u0ODJQTs6ewxivvh4N0
uvBl5mu7x5pppJRgsSgN8hAKoaXoTlVTS/CsemMFFyeiLHNKhKivLvTF6l2sHGfrYVBSw+o+baGs
46BBGRrcfpP1WMsj70sKnKqbV0fQH+rf+1F6uQDAOsDlTuVFhjXJiepSz/CCq6JY6BgrqNTaJoTg
gP603TBTxXvTgdv4EtOiDrEN2eiZzXajsYk6qluxnLota8R5ObgjhQqFf3M+gfkN2r8SAqhfykLj
USRL9uxwMhgW8oPR1nHyIDiiaa8Y4lsrayrVnJ/6WFPz/9whZau5XRRUzRGCCTlupKhuXAs3vutX
0Xd7U9ZhLe9krnS6u3yEdTvMSUxzlC7d/lzpv0Bi376HoN/VcdF4igB88mYOIDUL5JTYIYSXrJ0p
p/xzqwAdR9voO3g7CMPlf8EuNPIPNxeWHX80J558BN6jMtPq4Xl2hDYNIq5WWTA20w+Y35Iz01qz
NZwYhLRPeXS4+u1xPGcXjYn/7+zv346qSLMrY0/TiVvC6WUvm0Jek6srLIRsJcy5y2RKVzRS1jvX
Pjnay1p+3KKlwQatwRcbFblDrEKUz6fkMMTZtIS8sRc11BigcuPWniSb4745uZm5sArNMetVPOUe
nXU1GZfU+tWYd8kL2y9hqL2HrzI0rTOgj1VIeQMu4Zq3al0a1E18kTUtOpe17MahFSOeP+8q1tsv
/z5GjZMBYWs09DNRRjkxdMRFKp+XCVTUgrSBrtC5ImNtbPvgYdc7tcqNnBqaksz9ATMQ+/qKmkCY
v9GuqaWwd5hEYEc59zY6TAdFuF9SGZyyMVPP63dBXAa4j22u7u84MqQK/NJY+F2GpZCoZ3MTal27
sqC875ujpcMw029QEOOIuc6IdLtRDU67iNTrixbgOT9BkkomwXHcfdgICh+LLOSKkhEgsDkZnT/2
mHDYI9BPJaTmZlu4W5+po5WfeIbbXm8xo953nRokFRi2z9vYZiTQhUrt+cJg8rbKAee4f7XawmK5
mBLphnKiPaBJoGemyC6z4BlQdTOiNISdMblVdMiaY1Rp9TnuBiB6u2jMOLLLyKhYm/fi1xff+MJB
za4/MRqh6H1iv8CEQezrlJ6YanIKJhzDZveZ3dzU+GSnYLMZbtDVL8oH2xUHVn9aUaa7C9/UxXuB
WCroQ4VrpwE/3HrGgyWIhwanjMxz8gdDvEYJo3h/yZxT1YzOnf9BjVqHCE1+cqRDKaJswffd8h+3
5KL+xfPIhD6yaWDJ8tcgwzzos8lRikH/u7l6+Rc+NPJj2oU0LtTFBwOTYHoleBZgDp4r9FuDp5ju
WHHpzJ0lFyvFt4iLulLeLCtxXLLQqx0YV0wH4YVbCLE9HQTQeRWOi/5FOjBXeI0+TyoyWwEU1K2z
aAxPqUILuHEZvl+C7AEN0aQ82GH5Yv6NUxCIsn098jpktKrHknl029H0MT8flDFIRM2QpQc6lNdU
CGMpAJ3uBP9rbpr8trcJDxdUmCXLKAlw1vjythIPMeAB+kl18ANWYpQVCC96o18JK0ri/ryCX2E3
2ZB4+LEc08Q2Fl9KeUAxdKd6QTNdvX10DL8WpGHRE8DR2xUvkMs2QKGXNfGZgyJAaNqCzduFps2C
xscF/RLnEmfMQSMxNWttW+jZ0sRvhe6xriIox0u49Hzu12yhLQI8qcw4MzMJJYyuCUTVAIwQH41W
4s7S4vYUlBTAwDcZaf8QjJBsvJury4NGvvIT88FEb9nKfVh8ubcLQFdWFpeXcqZlg8SCWdx0elpK
jPBwhQM1mCX8ijNbb2ZIHvbI1s9vnMUVi8B3jG43uCSWbZfCaSBiHWJRUY3yqb1W4Pp6QXkNKr2e
t2rT36KM9ZdAS9gcMKDKpzUtW3FVEn5Owrqj+gzm2uGUaym1N6wgA17/oz6mQYuG4mZZ9v7G77P6
d7TQ2RVzIPiVeg3hsErch8zeIjdTm7L+2mw6pCpK6k2mlFZFbSs4ZR5Glwjw3cxXIvqGo+VKaLJG
pCcl1SHyFXJfWgea4AFd/xbvTV+sqg/wW+Kq3Rws/E0YwOtswwt52OavaJ19BJPxYh7NxkyjEEMu
TrtUvRJAqezxh2FGytrQqo39V3u47YYpDLUy6JBS99kSO3HLTcuX11b48wOi17oaXAlnT5ztbcKp
VxCehQOgQH+XKXrMPz0SkRCmKvvj0bBi3BsFfDOaCUYTE9DtA2o8i3N2Xjbsahj8HeAtafGMd7bd
BAbZyuZHy2sxCGvJKdaH1Y0vILeU2zrtGHUdj6laq5nk/QxjSJwmRUiJ2ZR9ti0Jq5VRKGXa0/9j
bJkvq1E8PatCFb9U13Msh1pue31rBT8DoUBDjdDZgrmAYDAiIxXQ/vpv04Sl0z1W9EVy8g4QgWVA
44xS85a8xb200yPJgFgtEXvGDTkilZ5OxDggcrQD/Bq7oSFDaZ9IwoBqshpjgiwhnWRDkJZMK8pQ
2dLXTm/UgG3RLiRXOvM8xrOffNcgUGr2N1Vqf+dR/M8RJrIdBuMEC52x2Xv9oYz7sDlekRgOdPuC
smnxVZGiHpEhRyQLNoA=
`protect end_protected
