-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
ZLvS0jA3lpidFWPRpB+2Yrqm8tt/6nluXw0QiAnMUnkIYa4+MlAM74RzenKLwLmfllqEefs9Ytuc
7xURblrXsIK5NSamxlEbMkqXcSFQlVTPlP7+3esU8cuWakd9xiLPjgTjBOqE8tZCW3B7DGzBp3oW
attVGdAGaYaIYCIAOYC6YMXnwJ/oWQOcX1hXeETKhtipDxJ6jJKA5dE/mmVAXUBldg3iKsqBWjgn
ywP57r288GWHKp/lO/hcgJV2h40lkXS2ulvoQwfmdoq9bdDnTJXeWhODmJarpxRw592f/9/wTy9s
TSVgua7O4R+zji9TqBDRCHnBx3XFgrrSAUP91A==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6800)
`protect data_block
x+cML2uQaOLwZxVKqRStAEGCyNRA9dshnzOvNY63IZSEt7fWWW4wnPGJppuE+qkyjIoU/JNrD6wZ
oadCNnZ8/T+MnRnKf5sF4YG4fpmDISJFGE3VDYKetMHdOY+pYDPvjZVLTRogewFOLH4o1PiH3zoN
DzCLmQsjt7ICRF3LT9Mpy2DGCUyV4vZiieNgHjlYTv3zsQUH/2mUd+98Wn0W/2+/S3HigR/kTdYk
1WCYKXAekwMUpXODIW9uCiRmMHpg8RDG+bp5CmBFZu7qQqvmCEy6nl8W2EqfKqnZjQcuIw2aIRjp
xVsX+JcajQ2gr/xbIu5vHQyCDrCpfAhWjInPXPWy6vWhyeOir6RmZcXePjo8Rof5jPmVQVUg2ogX
4C41OSLZ+ovNg22g74tg4vhkM5iP2huiHfHTDpOqZoFdJSRNVCz6a9PFx11vi9zJLzifqatBqyNu
dUit4VSxjEwM2GvC5X/apgka/uzf3G8p/kC27dn+viRK7fBXtHSIGfrEs485RJDVl58ArLb4NF0j
xk12SM65RXSYoc+PDyx6oQblppSyF8edLr1UKy4pdoRkf0OQmuGWLb+MMvEhdvV/XOtb5oMg6eS9
kH2OpIjgfH0WqMlY6D3IBA5L2bvQTgC3Ei3gp2zMPntq8pRWaDOlrxbYcSuElmIiuZWs40uSseQu
CwVU7tkdrwwsO+5pfBf8Qf2ZzL78QBkxrSi8KvAjv7+fppLiAsnDlA7DS/opmo+u2Pv0yXyXpq8m
6ELskMun81JFvXJWd+TLNXo2hOpby5wX4/sC9wN3FWeHJSDwmdYZUv4TI3B36qK3C6VX25eVLhL3
seXP5yXLxBusHKJ+StmQGDr7Go5VpHJoZGaNREc/36BhEO53jRq7mvjGtrLiDWfhLtyRrfMHfNYQ
TGnavLvJHCkRWRO++hK/6nl0/8VkEzeF2WwhHHbEtCNuclewdBB+kNhLPOds4jNFWAK+N5L4v9ku
EIqaC8Lx3SlC7sZQs6Kby2MEJd8BonotjRyq9OZpAdSvPkQRNMdOpV8vcpH3OYc4V8XrKzMq4Lmm
lzwhO9HFCH6UpIDeie87ynPndRnmRxSPtzX1VVfHz5/aU8xmfYl2BTtfH8iVJ4astAdZgqZFHesb
U7yG96XEGqOnC7ODPXe1OzB28LKX8WtM99wyiBNJmWpJHN18reJQ8D7JLVesv1OU9Tkh8oxMR4bQ
2m9PLzfEX4uY5V63SZ9Ytyg5C/OCLmRcaBzH+QX3cjF+Ez8sQMidFTNUl5KAdXBqZCY2ZLggG+83
392xTRrtcvsl6+aXnf58G36tz9fxLrAKX56j7G4424NOvk9cOUVv5zoaBszz1zRvSQhjq7/2zfTE
QpojYSV6D5CBxkp9sIFBmBEEi5ZZH14u0akq0ClfYgeohYf1wCCIjKdTw+2pe4NB0Mc45DM0DA27
zqCAU4J9XqDqrIfOkthM1gmvPksMaYPLLbcD0+zyYDJY6Nug5J5881twJC07Nq/9ysWbiDfbOj7Q
O6cEQo+ApCCY9yfy7UsYK4MZ1TtdWbn5Zw2MS1H4MLhTKyoora+rUfp1xbPhm6jZsMgaoRYPlUEC
b14u4X0gt18cvmS7yoCjTKGcHu6UA2+At2p4vXnF5NJspO6T3HILpzRp6s8zqCZwc8xB4U1srfrs
W7Zg7fTzolsHfhXJIIr59gAXFS+Pfe7fGVOqGEAF3FPYayc2Qa7KwAmG9NOzrwJmjMlgsDZx5gS2
1p3AyPD4wJEc/eTVfhHUA7fb+Yyz4bKZFlXLb1E+RyEDA3mpVcVt7IARJW913RMhiJrDR68zzdVp
oaMDLuV5dwstJGuxXw365H2Q0H54U90+pJ3BusoeQ7GYiYjd4iZFE3KkKR36U4vltP5BOXzxWPPs
bKj/UAVhTdvrmKucRj5ewM90RWNmOggw5+FiaW1WkFb3Ar2JOX0ova6NLkL0SxX69F3eM1Opg74p
1qAKC3CwzkIKmqdrsCVaAr01foHqv1+VhJKFObX4lL73UXV+3tXYvfOMdhXA+ySOmqx3c1GTg6Vo
TqYVw6v06+Ql+GhpCJyi57fd6FTDesCg6gm07mkK6Q/Y61uHpzh/iwpkG69u+4hFwoHq4NAzQuED
LdVmPJmiZ/ISl3g9ut4qIEgZM1K8TpwGjFzhsk6dl0uOAvwVKadq4Cuoiy4Lxwn5zSAounNNyuwK
v1xtset+nXuPu5OZq0pFTmglrS2dcbozJDXgM4BP8EnEDj1GGsc0NTVpjvrZfnh6LjQGUOPtzJFR
dpv7i3ETrwGtWtlFlKwHMmVtkXFSUIX7GxqLV57BgwYeSONO+MDpOeDff3a3JZKYHg1ebey1gdEb
T/vJ2okYmed85IVZHjG1a/D2P6W/4W0IRNJewCeKTinHpo+BifAvJwTvUSs1iYAkkY84j3G0TLi0
6Iufk/13/U1Li7sJ423S8nzfAnTZg1OabnAuNx0dSOfeLuwuGrhqOrePVVo1UsIV3Hbku5F+9BpD
c0vr/ogWWC4NDUs302AgGszXkrGqWWwMj1ez7bAsZHIp1waAFX7aPkNJt1/AQ57TP23iHCYugvsq
xNrqSiOcX5jUaE5OKQOmlHrRtBMfC+Zqja1tBEv3QmtA1epOx9pYNhRiHT6dfHQmeRmHP0JMd592
fikL5aPXV81btf8quHRF80FzCxEyFP7oWouvSAauaQWN6sRbCMYsZffwm1Xlm6FNrKBsA6VKtUbi
D71J/zem+QysC47dS/o5XU1G3Q5CCPdvp/79CfU5kehHsKJj2Ku7og/wTt6YGnLy8vHv1t5dnwd4
2xf+f5oAZ5SIYSbxi4aPu5mMHgmpeO7WwaYEXhvl23C1KL1nB5Kg9KoGdcJLqkC6SHMWKOMS1mda
8765FF9CujDuHz97wuwdpEWj2t3UG83Pyz5zCb+DA7YzxiKvTu6Bi8m6sW+C8gMwXyEtCJekFXc1
nUTthMPI+UOeIcihADbi2zJB6VaSgFuYD/4Ve+rWbl7XNPXd+Nd67ym5eRqy3Bv4DX4pn3Uwipm+
ZDVVZm+6Muha3sYVbB2IlsAiLDCqTBUWAfu1S7s+SSZnlK+p92CYxdLr9I6C+VGJt+Ot1ZdhyIK8
gaHIU/Rdb+yEntVYIADammQDN6xwWkK57otlDMx1zeLQe533QgWRH15J8IvF6FZNjEgLPjUYPtm8
1vWw2TL33X+g6iVjoHOP8+rPYGOol9L01JhAGMy84zh1nYuLs46X4DXtEisKch/aCKXFDB2ln02M
LscTHHGFlMiyVAy0f/NrfIYiJV7SffAlX25BGh6E3Xe+pXsccqEIC3mD8uMwQf0nLijfGMLnhSMe
v7HJXA8ZY56a8maWxl+GPLn6TRC0tDfAGKG3B6W7mcZ7V7lVx40A5GYjDsrZqslx8UF6A91GrAnh
SW0umtlcGn30e5w9vw6o0qJbEWDQBlYky/lrdbeo5rUwQ5le4HB1x01LrAh/+h2tzdYrXHf5JWH+
4KixYVoUJhVe8Ns9H1m444LtUhhhOlCOncGtZZ7JkkLI1jeaXFM6soC+d5EvOotNPZYgxyIgJeSY
QrNq8luqzmINQ+PJtWDQ3r/diSTomcZpPLi2uR2GlnYIFi9h0E/2MT1J/XTfJ55WlZUYiou+jI2m
YHJjn78AMJS5lJnmrzRumu1nlGpiouV81kXVLrIlksb+mlFOj0lMGv1r6GpC3kLt0PaHKxcS8xmR
3Y4aHnFFNxtmKIvLQRrvszTNRpwbAN1d6zEvM8kgHMz/aID3I+vln2WeqdkJ2ZUiecf+riYZEVux
OX+kjge6SBok64jwLjrFHHmA65gNmupNWPJsBELSPXveqkTxa5re5tvlcVJhd04ZZb1/R30HUM1b
87cFgBObQOrEWHx042LZgHhIJJOJ1eE3kbGhV8NMH1e4JgUeh792nAir3+0YSgeTQMZAjQJkA55J
38Wnj+SAUo3+TUfx19PnJaM+IjW10Phb5fj7iE0+u6v9Zhrx8YLuYH+xvAo395Br4Mvoskx/NuDw
/sh7iRQTr3zC2Y318bW5iCA6gIfDza9VV0qoVGlBrG1pEM6W/DoxEKRVUAYJzrOLKz+CNIT+GVh5
06HZUqb69WJKGilwxOTbYiA8gfhd3ddzv53S70wMtKYXw8nc4NKNf2Z7CNdHMcedVx/SrfuDzEWq
Q5uhHJJ56M64061Cd8XISaUKAhspivzijlt9mvnwWQmGvE4rX3I3apVquPT1AU3SuoI92JEySev6
Wk80/nMXQViRTvqLdSUnWD+AOZ2aHHQRKgBbYNva0mcUCaQdfTnzBdzrNhEporYFNWcABGwhI2Sn
9M1i0obv/gw5DKv5tiJ9Ln/cs7rJJl3NcYjWSloh5VpYPYcJV/QWUuj17TkxPvYpltaJ8l5ds/Kj
7Js24beYcypANf2du6eKwCwV5D85YXhSthRw76RDO1FnoVq/BQ9jw4v8Rr+dcSjWxiCD/8PbJ84i
6DAWuAbTUWnI4vLUhnd8GUnnzwSlkeOoQcmXCSgzoWXVsyRmt07o8nHebLDZYuPIUqsPSLNDe1xO
tiFEPYhAdHVS/yf20of/pv4ybl+N85XuXonljRHa4xzXahyc3ZfmoZuCzTR5bMvJ9N9YKh3xfCGs
tP+NgA7NlkyStvYmGgEwQwNCjP3JNqJCZZ1iNoxNgvbrlZdvm/sOEVfZhj+pqMMeKd0M2R+OAh8E
b3wdVFNQvHiLo/NZ/jkKOVjvlPdFmS+1QQ0uLo1aMzdWbz+5QwRPcWqLyUvnatmV7+mmUcs3a1/f
z/bp4YCJfzlhfv2wJiYd+BMQ+d3YQ/QK6CPgkWFLSns0yDNLdoGJIibRKtTFdXvI06c1+dH5W7q7
V7QiLlgbM49i2Uowne68F2QUVXnulzHD68CFVXGrwk+3lA1iXZ827qxCnkMLJ1go4km5Ok8yfUmJ
dvWbZsyoYqwNub5PSMVlygDbNvc+xuMlp2bgHiFpOB+ESKOVT5dAxs30WgJVkwQOY08/hjfIAqsc
oU1IVSjAfP5rjDVwSDeemkh9E0nNUs12epTzz7Tklo2U6MBiVWlqKFvlUpUPetkNkPW5Z/N0DTGD
T2O8s0uaDY3eBVqbWAvEtFCzNEvIm6fVwawdh0u9NdGn30DfUQjh0gH4+woDkbP0w3JpE8Hb8s0S
24OWrRKHCRSaXqsQ26+M1UUXjiYXOfIZjIUlUt5e592DGUsHoo4aBo369lWWrZT9R0DFDb/UA2nM
f3JZ9J9Tu2k2aQzxtRei/zYwty6yc/LgvSBb5BgC3SOUIfLmiA5mg805i4Q7ALPzN7QWgiIPsGOu
RsC2mzxMH7/PXEJKd2TiWqZDPbHshpmupfTq/Lx1K+j7AbMCXQgjYFB3l7+/Tw72dLvv8IXG7oSy
W3bLmg/OEzBCwG3UdnkavYEQ9jgaqy/Vo7v5dvVkLfMMPhavy6i8TGnmL3Gqy62acnzQ8r5rLx8F
UAMlWp7z4ShC8/U3LVFSPjLxvYCkYusD3DU1BsNC2bqCKYwhMmWZmTxkjk7su+OPJ8K422G9g7DP
m1rTdeSQQTKzv8QSgNpQofP2sH709IRRo2CKJVr/NXLrmL486mUjx9IVgmI+TTw+rJONiIfJNVEf
/haqWH3F9B6WC6n1ifp5ds+ZIjcvAwGc5dp8fLgCasigeehI35R3R3c5YnknH/NMjMfebCuY+9ic
6X/nrGDAFjSVqOI62a5gry/SUrUBRv5qPH+ULSVmJTSZXWP1a22N+nFAXqMC+gUqd1dPxsTEfYej
HxAnYTvOvum4u2wcqi2/Ka6VZDN76CIqZcvA0jGSl/2DfzL3hoZtQgTqf4YUnRSRO32NAfP1eVyb
+A0cbxR2srFqefzLHOiulR9ytgHFsni5LB9V0iYnUeUhxNUbNzdTkoY5xtxxuGAP3mSbE5ah/75D
vpe3D4znPkUXWHHuzM/GMQ6NIE3r3YXrdZ9yARsdvJCtYTGeHSsr5YpU4kUft5VlbruCZv957BqG
Bdh/2KjsW4Hh6kauXPRV2gpeJXnJ5yKvVqgXiOGEz6ud/yqPwNdS/8kswP+A7vEhZMtfcebZUtm2
Tn0l19l+O2F6ROn/6G+lj32IjZfvUxojVwZayaGkxJfUTD0u0yrhtfD0UkM08562nCKcTQda+g4l
9YNuuZ64LdALkEreGn9pb6xSKsWnsF24NqQ0TtXObv2ZuVV2cYk+LeKwqvMfqO/NBYsmmfXoCsGP
aMNb8AQNsxu3Q47Mmu/Qq2d0lH9qrStalgNZsCJnys8s4nA32/wMKurPsEVEwU2C8f+FYktDj1HR
SeCTy90T49o2NkcFI5ltWQPLp3pb2LxYLt2eIcJ0HZPqVJX2j+nZ5l8+b4/bpSnuyILY1VqAxiY1
7Zfz883Mf5vQdyAZ5VGfq25P1zXCg/m65OptUhw/emg3CHkkF6BIrkh8nNwFJUSHIATV9B1K0yrX
s/2vNoN36gLaF5spl5+n+uD6sOn3fooxx37OqQsa44cI9EWDbSaFwLd4OElvZ7v4ZF9DWSIKyT26
rJ6D+9rFe7f2RyoVMH8cCnhVXJ2Q4rqAYdbZEmh/rus6qwWIsmol2lPR5Q1InM6X8LP+ZUvRFMof
RVt/kfockDcBy3YuxHkUHownMoQSGo9QBTcQPqjvjvbMaSz35kDKjCuLYyO6Vg+94zH6YjHhV+0k
LFWuX4r6pk0sN4+f/GfZUtAPKLufZw+nK1QqBtWGd7qjwR2/5499HVk6wYZU66BhBeG+nyHjTQPT
tx5SpU9zQ/OmooazOl6CggiObgw5SxhT8JpIUeosAMefWIYk9lx//B1MMdC6iQjOrlpjHBgbaznw
rIrL6l3OiTvG0qMBEC4xT0pvNaHz3KzsO3M8sR4NJXlhaazhyP+prtKVxk2Rk0BK15OdAIBXlrn9
ko6OQCZTDU6aBSQiEyznUzUaRxK4bIDQ0iBjSCqiN3iFB0TiPXqLltMHhN0KmNMVvJU32SuaL3jv
5zbgaWGImruSpJPsYEXc1uPWWsyS/9oHo7gq6enTZwVvI47sqLm3/f6sfpk4/ATKhm+6e1544hWP
Bgc7r7FsFcvdAAG6zVIJB7l3J57nAEIIXjpiMjb4amrPWqFhcKhUi+g+Z78n5KJb6Fx1Sm6Czaa1
befLc1/xlPjMLRcNNpK42rbgtdk/MopRU9b9Uzxge4CVU6JN+LpbL/YfOEUIQidpPWlpvVwLyrwY
eu6HSoZNFj0yvLMB0Z0NOyHRghIY9jWTvn1lQYHbFhEqo+izzn0anN5MIsdwp6PTr7rclushdNrJ
ZESd1fVBWPZ+JDabQcsaPoKufkZVMHPzMrmBod2Bv4UYzOZCOHEFKTUPcsmZWeVMlc9yrFXvnfgV
8Hj/d2XCf1pO82EVbmMNIL1gMCgPAmaZtSm63dDxFW/1OyJxZE1clk3hITEOHgriTl8ZKvpH9VBu
Lt2OkqXrMaGwoAJVS3o2gm5h3WXSldVvnAlTE5gdAkMkuKz2keiFB1Gb1mLzThhCn7FQmAtiYOaC
RDc3cpA3Pgdqgdgb9OZ4eFbhADX2d5tir0akGJBBYSMDA/BLI69QIp5GdCA+xw3H+3kQvNsoUMLR
MDKOsIXbSkhAFoYjyxVQPtD8YHtiI37UtqERBCLlFsBfqAKOGGoje50LSeRqsRP+nQnyUZ24ydhM
/TyoN02FZyHmjiyIK1Une5fzd19vj5FCH6UdS4L14OVEL3KXty0YOf+tXQZEtvlfbuIhbB8RLT3T
xtCDgneJ0UEaG+hLLASP/QD9dfWoNyCG9e147kE/cQnaTVSnejjxnjyvo9LbIoTti3u5p9p1ePxd
pIN3xiSz8ofA2clLjLqpTjiNc2XUnaeLYcQrcC8qffOV8I6+XntVF9u4MkupnyCrUQyypKAuxDB/
NBVFQt406lle4Bb3iWqzvByAgN5to6DolZehUkeBTsykutraRTaUIA4TKZR4raYpypIbK38XTapb
0xJ5H7A0yhVk0r60x9HZjqYY+SeViQG9EiUIB9SProYV5Qp7AeDo9W3njnTcFrLZnMbD8Ea/6lVi
4VVB+bpGONUXjJfddVNsNBsKdh7UbPoV1kJMGxJbhQxNPPVy/xv0PzW9tSMw9qHt1V5qOk0K9N3E
rrT+2fmVgmxVLP+5SE6T2dXph28vuWiOxLIg3daUkKqN1Sylke6dvcfciDehWETAJqjdSoW9epQN
KYZ8xl8JUHm7cKubzDxEJUZgLiR5fUXirPRay1Cfj+BBVyKObeON07frNwmUK32e/F/CbLQVv6ty
0KgEiUjgXo5BQXMOOpHo29zyWgnUFmQeH/ZmFhN1O4tjqn+Hrv4+s5TqL+6/xHWCjXa1LHMTKRz0
C1rnzdvKHWrdlLoSeNfQ+GXlDJXecr6s4oSroL46RRr0DnVehrWLqFD7P83RSWXcrg0kHLjbObvH
ZcwsqzRidDTq4ErJaZwMYJr3HqQ7UjmVBA4cO7QewpI0xj/TkFJqR8UdyegDFdgyQfatTzLcE8LL
D8w+4aB+HLo6Dg7qSVfSsvpQbhDcp+VomDMhS6gWAhBZhZt1SCrQdZzv3/8PFErgDiwq6LNOHOlC
L388MESWhl/6Uq0hy+wsORnxGzmdmt1JMgj+wWIitOy8FQA1zSi6iPJuu4AffrW/KBncuu8206er
1ubQRlM6yWp8mRfrmVy52qRTEQmtUm3WACbzMjibxqCNKn09HB6VoFhgvWA6Ys6NwH+Q8QMJ5+8t
gR9nltOwfU1DFR3iUPgqYBWSBM6gWv6peCqF7ONXtTVbNWQHQvNJZbyOjrbSziSVW9l6F8jSp0hy
JMem0JNrXSNwVtrdrr0/sKPRp2QJoSZZop5xSlgmLeFcHI6MVa0amZ/RbIcDjOLs4jZVPhkN2O14
BTsbRynJ2zXf198nqxkttKhGjmWskTX8Q0U3sQhw8TOBwrONegM53/sHxhOQRqLLQIX1W/cBMJIh
yCMDuMRe2DZ5TuhrqtSrEikcZGX0ak1TpimhCXqgbgUahT1SzAoNvcCGAsxhxxtnWXksqighqO3+
7F+TiJWq/NxHznt7UyBVBMg=
`protect end_protected
