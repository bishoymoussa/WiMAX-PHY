-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
zWkElFg1VCUH0TzoQUwsnial6jzdaLpO/cQ3q6rpZWgg/6zpCnpWlz3KoPbSMSXHU8men8V+Bn+O
Yjaf8Eta7EcmIz5oHUIwzo1ncoPe8883tKkTrE1GYbbdWizGmhf0m2hRIoVPu+CHyjx6KyPJvwYU
RjiSsl1pl7bRwpm1vOBV8YMy4+mAtUSwE0l+1vfKsZryZ3Y1s5laFLNQy2HCD0YWVNmkX2UuFGjR
X/W+fS3vckTvlySUtPCt2B7zMLc934hIZ9GnPmdMJ4V4xBnYdoxaHXqe/XbjJFy1FcUcP7BrQQkC
mb3Edh6VkrqmTN9HHxKehJeg0+8YcC7SehMBlg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 9616)
`protect data_block
02wmvpMFj0jx+OI6wO8iQkHQ4qD3oZpGdsO/ScIJn7zEFUAZ91IwooDXZNuT2/a1sJGt5GlEbp+p
XMeLWsO61vKyFasvY7nT/LGOqbGrkcZZ86XbZ5E8/ZFJO+G2XUqxXvGazKCMCTu60NT276rSz38u
xWy72q9xByn7kOgkNpSXPKlRHKNldl+WbmVnuI2SN07OXPbDWxm0Q9sNgtN31Bl7e86zqKKHbPOU
QOUGV4hzTIohWJusPWwzs8ttt52+WEk/EbSA09laQE/IavtSPSXAhazZL5V65WD6Sc4gb/2ib0iP
+AiXgvOwp7WSMpRkn6+kKY/ysB/lqdBdjsJwh1RNwYqPNAlNxjxYrtmu9CFuTVO1M9jv3WKUy7Wu
xB8Lg9kVgNto4HEsfy42VZz33D7p9jq4JBAtnFEg3Z64y3FlVse+WueF3A/laQsuB7mHwo6o0U/c
8LWdn3MZwZsBbMIIIK9Nrkm3IvdTLyc3KEDex18BeqsEIn6HEC4VSCSQZhmEcErNK2PKzmXmRuCJ
3DkMf5VNMx/DDw/WEZtWzJnYZh1FI2zzu69XNyUTHW2DGwM6V1+G+5yENOMkCzShHChr3oScxH7l
fhsst3JmimUMKSKI+d/6fos+bgk6XXf+uXoUZmI3+Us1txim2uH7psC7lHaMS+cUnepFgGOL/o1c
MtOYwupXAiu0zag6QTmROTZN7Nhv+tEQbCBRbfmz8/xCqwbw1+xBH5OJFULIYJW6Af4JXABfcRE/
6tfzRwPIodcBpwWysBDry6i02yMO3itZu6qzKlhKRegnF58oxQOBD92RhwVBU+BgU8FeuYvjVC1h
u9rS6Qt7gEDC7C5slPiElbRnEwTrfC9AMckiG/f2OTusmqNjOZbIWD4EEfTx6xTshZwBVKNmMq7t
CR7sMBEaHmk3aqf8epcSgq3h5rKdOaGE5FKLxfyTFS89y1W6ypNDuY9aohDG85qwvKqDm2RUg4tH
Vkz1QvlWH7qnVC/8Op+ZODZyhkGyx6Mq5x6Pd/aZiQLWLzkuaLh2ZkVxS8NK88cn+G8oybfAc14Z
oe5P4aAq+5fELn3WzCYFGyb5wH+nSqWEfT648lP2NA355LQslAdAEPPbLc1Mh1d/CEeNTXaQWAtj
VG/VWs3x4WlY51iuZ2Ep1rMH1KnaVf7ouMJ24dokOGCSso8lkEezE7+OKhWQ661FeYmmBP9nQDjs
63nPtwyUbC+6slgZRUPwwb9Wg9/OoRhYmQBlMDIYnN0WcikWPnH74SK14cVE3dsBAc5FjVLTk4G2
Dk4HcbgheRrir9kMwEaJMU095y4muqsh1qM8dvdKK3wj1uD/hR33wqzLazB580woomNDHWmlMV51
H1ZGlGHl0pYiz0m+Ydkn0rvbiJXTDSYA+z5aTIL+KZpG5N8pKZd7qJghCsAgKoJghEW9TRk9IlsB
htHHqqJnVgMC8fXnX0ZSLWdY4gjH15H2PzAkziOIFap+vMLFx2zHmqBNHnAiokfhbalY0FHXsCVL
xGDvGChqItPvwgaPZZL8ii6awXfzRtJVp+5B0H8DVZWVgs5F8ncU9u0h3TKMHi2R7oWPyIlOrzPn
SNRZHFORcYs+ptr7ofRMg4BocWpnv46atjO2HPkSi0WhVhM045FCopBk/mrdRuwiF2mBmgQ+rrDp
dDIHgWMc/ONm17O2062sJ02uVE2hGApofjxv0qrr3m6b9E6fF8BaS5GQvMRU28yC1r7sFtMIKFga
kZpyaOhHTT2jqlAIewY35Xl6DWRZ8R112Cn9ka2xZaMhaR4Ge5AXQajHmF39nleFD8zv/uOHobnN
EqWJ6Qiz0+FqJXcUG0oJehjhEplU6GVyKmpsLOrmfwyjR6dSwuzwKMpm/oMYtyjcM0SnOW6Q4fjw
TOPxpVEYr0ZYNjTLKGLn+WZuwDxIOydPDNjh/kRg3UkFhCg4hxHCLsZjy+Px/VsKS9hadtD66di9
c4HEP3Cy48XQQ6KRRSoIEkehH2yP0aOuGaJuWyHJa7eQbsziDiFh20mNk9NrnKDbtQOax+1TbGhT
vaFqbvdW1fvjzDNN2xHtUORQs18mtDyQKfaeSKzO0QcFVhm1YaYqgY9nLqRd/FgEmNsm4w3lgrfg
KLv2OO6G4P3ZIhJAQq/CcUJSkvlWDezu0GwLbUorSJ2EHGHikv3N59X8/OBsO+eJgVT3DlPjOp8x
4N2/O9e42ZEo2qHR1jF0B+9RyQCML3gQQCB+hadKajYw49hhugkmW81JFdgdZsem/uB5eytemtPX
F0B+8cvMiXNGjMRNF09HLoBMyNveiNOVTym/Eqn0u4vFP2c/3RK2Z0TavVQmh753b5aL9Xz+S9Hl
l+Du0Pi0+k7NljHzmHSADaIuxk/o9nrH1x2pMn/vtpqOaN83wGvaQACgLIgK8z7u3EB0vv7jGbY3
amrgcCWtC2uP4aIXc88w1ks1NiNH3oJIjwZQfFn1x27L2qRT0qwe9TKdtDCefFLjnR1daWyJfQ/D
rF+EERuQYB7seRZK8RL7BDYB5xNNlDeGz18dSWU5mwGNRYjBE255p7F/JV7TPq0XGaAvb9gc4b89
45K0GhJZhuPERVzPfK/z3OmaJmivR6vKePSoUthqi7B3T0xIyo4NAHXxi5KagSgAT2miju87ihqS
2wJjRDitjxlRjhsQo+tOPTB6+GhYdTAZu29/HzV6jw613Ss8rR/AtC3W7HoVkdWROHAzoeeZa59N
9RmUcHfuN8VZ/uvJVFF8IC39AbYck6Kg1YYWrI+3g67eEsPzFWAHM9nMR0hIknSh7A0Pp0M6YFJ6
wVQ4x/F2z7+gkm0W3383YPRpGeczmKBbTsuuiQSgPA8B5N3/9NR68eg+6pY2WyyRiGx7BbgXPGRv
NkEbDgtL4h4v06oL2bokqNCAP1HbdhQR8RzZPe3ZuaXLDgI2ENbzAUV6Nj2Vy++NGkv6UGfKytDZ
St0qY7PeZeM93lpvO06HzxNQo6AC0FLjyn4Y7u0wsCUof3xVUuhyVcJz8z1q7nMKbqMWJmt4pwak
aNme/jGrdxvPEDMngp8Kq2HFWEmZh0w98eA3DgJntbLXEcLaiRxtcUQHQb6S+I+h9Jgvhew+fqnw
n0tiRQOX7oI/IXQTe9qJ+PDdkUz/MdLo5RlIIJPO2oe2QSbe1+AeV/+6c+9adIXMJFpotGLCHfS2
6YHaGHxOpHLqHTBANlYIbWONgfGIO/04VWVnQKGKVbfQ+rTCSliij0vCHmbu/a+CpjovX7mU9air
rwneetajAQhmjI3o3mjBcqU995YiI/4JExGRhEfxbE1sqPUSzmnH2hdI841meLGiytlasv8lOXU9
3V0sg8SkKx0hsvZ8GM6fsyQLdrxM6aFjkp0kWNY6WDVTTLRlFCmh9LNrfErfdofU6Gno+ND2R/pU
UNbov7CDUUw5iV8u4mE9D5s2ku4F5xEqR5gV7bidARZmzcON6nBbnk+oQkEQQrvc+ALKMNGLRGzm
+HRduLIGIiQDj7fN6cGd9mAtExMwZ+esYcjgIm6c5N/C+FLWgNEHpG/FJjUHWWv8dQDrWwme18vL
UYYbyDrgl/zsg61qSKiF1MqBt7ptrxk2YezmBwBrM9m5iYRC6+c1YeMnHWMx7c60yeC9Lrxe7nyf
ZwpDjOjDI/PoxCdabrDWb2f8g94SxApxsKp7tZnd1Z8RcavXiRixfs2mtZo4NmVfcmhClPb8fakD
ry3QsPs0dd/12dBeA+OEb4ALB3m7UjO/f/DiPui6jD58W61NHDCD0uKI8ACK9YA5Q+vkhuIzMwB/
BQlNharmkmOAktJH5zgZC2EdEQm61AxpaKrVv7Af9tFS1mMk+VvUsTYh2Cet6IyAhE+wtFaJzDhI
GJ95Ys47eJ6ugqqiP/7WmIW8y04LWUnvuWcky3yZsKH/bORyfaYhQnjWA6cObM3XRKQtonWb1yQ7
Y2Q5NRDL0alWzmw7mZpp8arQYWRYh5g25NA9jc6k1RrRZjYsP/tbPDMkeGekRJ6paHeVXk3P80wJ
pWeS17W+RBZ96fsmB8EkfkL+uyH0R/NaZMnl50oDDOVO3gybxHBIR29dn4NEzcZiSEigHVkpYAQG
a1VtG1ltKteGKCvmSHedsjP7/cpqVfF6ZQZ/Bp77MkKhMO97B86cTtOtyByt4Unqp4lhS8PqXIGP
KC5S4RnEkaFGaixz5v21EEcaTihMRaVRsCc88Wmb9cnTcqf8Idm66ESS2eNaTeJsxzyGmSNWL5mI
w7d51+UTREpEr1cPsZ/KYiWp4QLG9Joyyiy3GZqMFyppHLb4Uh+KIYmh74lSihMvRcl6VfXDHUuO
gEA0FbCy/bvnnyGEZLuxiz9ih3mbP4vy4R+HDU0Tm1LVEGIXeRG49Xhk3J8tOH3MEw24CT5nfyrw
PsP09CHqreF4Xj+7iaAgt1eOGAImDB8/x49VWJXUkbQv7qP/pB1o8tSnMlyajrVEBzzgMspeS7TA
xeSUyXaEUPJUYh/Y+EDrD4U5tz0i7BKB8zso5BGPhgueO6nRR3ret4unjLtfcWGCQ3AdgCx0sNn5
eLh1Hfx+RNXAdwD4QBV49GiQ6NGh7sz2UFJgdvU7i0rCWbbSVUX/sEsuucwiN1CcdOncUM6Mrl4X
5UaB3m8kunpxVJ9gS3AdeT6t0SJ4Exd3dHT8abTE1NeVEG90wjK/8T5vzUvo1OzBt0LWu5pdd1Zq
Jwtlfmu32h+Iftss3IKMidGqSdKS5YKBlMZy6trhqcvhZ6hcPe8glwuA/zD1WOdrThQFc3mWFBQx
QV+b/H8nF/8WkcUQqttqo8+x1tOng9HzdnBA/8bBhowaDVwltx+KgUJm3Ndz7WhkR85or3dut/Yn
AlWg0m9MZYTV2m/IC9M4ciaXbLVWXXICmBTdEMRmdSzJZdYBlcPwstvy5egpxWxoCQXvPBEKTmwY
PSJBzS/l4e3njfUuynLYxGnXyaW/MyUsG4XDI+M232MNeirJxI6KfSq/Dhcq3r/ax4cdRx/H1IzI
wyp0oObsEuNmq5h0e8VmeLRt0rXrr2FpihY+nWyUlyyHu0VCGdqEnFhQWOPpAybvaCEWRZ/TJYEN
5MvoqBMqCM5Qe0xPS3NAAoSA6uNQFOS0HrfMb2r4JR35IPGR/4C2Q8g6N4EV4AlqQuZEyePeZoGd
EnEzLm95btae5/NL1iY/ybMe35MMdKuhMXgG3mCOKlus2rSm8qiJKrt6AkrNUPiksZmINdM1zT+e
0wmjdI5W9v6pPWThcA1AYvMqO4U1ixMIJFZTPN2h1cq16MaL7oxpnuU+Rx0wZk/ZXjw1z7B1EbxU
0UMMQBNKzmctP/C9xW202fCrnYhFBl3lwgHYLHfDckaIGTMPiApMOjY64ai9E1oojOr0X0wY3uY3
NumwTb4DmPiWo9RjAxTzv8ALmOtDWyDZV9EjjzDu00vKu4nJtt0q9Z2fO8JzuKUFMbBqrqzgMqwm
40vX2C5+kPjrL2xKEkPNpQnuAOWg2HRRxjXAnIglmljtFRo6zIoyQh77/5TiJ/Fq69bzdjduoOSM
S043u79hcMfjcNVhRbQmXOWFHGfFP5TnVKSkFC3lROMeLEa1NPplUMwPJOXdjZbojct/tilJn+it
GtcJ5mzNUD46f2J8Bw7fZzFAHomz4vTc4YvTwlqhh6rdb8ThkWFdpCL2nuLEjvWdZuEm1fJd7Wa/
a9IBFXvAPZQuCQ0tRd+QT+wal+c7hW9N8wUi3p0cR7CCy+w92uRNPzc51+xaSLEEr56qoy2bjrg6
zl0Zc37ex9GNnc8mgNUVEf8LXEIpsNGRIUyREaBqKiol/7/Pt9JN0xh8bO97ZhR+MVl2TRBlUTyD
hIJ6GKRLT3dgkey/PlLRRHL0zBnmHErb3+hGfO3+P2AqzYdaKDMPlIihSjbK15db/TYb0LG1XHBj
8rIK/kVWnL9uO/3QAf+gOJxnzkrbO0Vo3LjWOI6w1pMeZNQQPHieZxYrQydrYba+CowzHIP+SI/M
ymtxrUQgUohWGbXvankoJ+jNj1xSWI4ry8KUez4g/rRDImnn1niS+/BXiwpPoBdNkGpn4pndkBhj
GSjvP2GUGe6mvfh6ex1TpCUbUzgKZZ4RwGlxYzCfr9zW+fYi/eo4akp1aq90usqnclrtnwMBY3ER
aKCJpiH9j8pU4+BDbSneBcs74bPte4NVFBqK8SOPtfLs42hc+Hxdx1m+SCjrh+ayUhzLMsF9U07h
JG/ikgVPYKNpV1hcMRsHKcR/FWKF3jgjFxgNpK18sH/wBFJjjLKXN3WobCyUBPnw2Th4t5qzM3j3
7Eo2O7enZEUPKKdQBw2oeR68ScfPMdUecYB9110Q0Xqzr86jZicjf2D1ybAoPMwQyhJ8nNRPfcwM
JKQrzAfmVAbPulSX7cmPvhns0WOSRSXgRgd9VW2xrKJ2TpSj+tMphuiubsGFhK99vB2bkeHNnWHe
ONCZWdz9P5aDTHE1gmIea0cSRx+53Z7lF+N4e6ZyCIVQ5iEljlzur3UL4tX1GHhYmPVTKNPDL3b1
V36QkNXgM8U1iOPI41qUztLU/WulU/cUBGcUVJ8JsRU6nxwheZlDS4a12q43BsYa7hEVTjvALjcl
MBGsbcQLUomEb2O4NOqoYTHSYiY9+P17hYopJsLgzxXL6+wCbyLHlA3XM/O09i6VqJYKqNQj9ms4
LnOy1FdJJ8brqTWd4/MJzDMiwlCN+L2+nDKHwUsoXCJ78gWcGdULJZTBc448ENYKmlab6VqBEjT4
cI0ZvSm671tc54Wtv4auqNHJP5FSTzO/5Tlp8WR8+e5h3zI6aI4vyoFcrE+9HyyhSVBu7vxhSxjR
Y1uQtAPRD8pFwfytTrEgutZ+eCtOQGU/R4HWO3TJG4f05u+weEDxIjpntMXQpO+G6KAa8AIEvWeV
L8WPUKD9+WKZGIZ/5dser6sRV2ZqtJi5+dzQtlJoFTBxuZMn5QgdQf5O4lCMqHzQ+wZroujqsBWp
Vs9tRLJURSn5SqTT/qo3YAwy7Ts3lnrN8mNWEZKZDC96xHpbJG4VwQzRsP5vXruI/Ni4BBvePa/n
joxpMAX7wkbldCHAElEnIa3KW9gQGLPT4X1Rq06rfooPM+KtGMePFH2NUTdf5LwPONTrVbCzSB00
JItyHIuA5MX6MEdmzrUcerqiApbxlxmC27A76K0aM5i69o2cLfO3jzkXXQUhU+fhGdo4MQiSADyR
I3BlPhgsv6YgAX+yyDqbij3AWDoYs10aK0YUdXI4n+KjLE4SOa6tf0fBlqVoPsQsfl0Y+j9LYL+Y
UtEFcPOsnBlTAzEOCh5RMHGoveagFOrfzTI/sAv5gBA9uSLXdDDR3qo2jSBHMUAhHREeVVC0RXr4
GQ0hI0J4HeG7FETm7/ALJtiZwHcQPGIGNVkNhb79FS7Oj0XYbBnIy+7BP2PfI7CAT2JXG+li5/Zo
kXra4meV3aIhEXSL+O+cWCE8Zefk+c3yaL+lWKyFXgFgmiJm6HivJ5I0d/0OWuBEHZoitaPQ/0D7
OCiBFYzcz+xkWb0MOm1xWwiKeHd5V5B6aN2d1xKSUg6sNSrerdlGSU36yw5zKH8EJEG8enHUn/a7
MjnKdKqmAUC86/fKhwpBxemntjtMcQy7SSCAiKym3RxRAa6qk9ST0SbR+K81ObRVfvynN2fEDR4S
w4BnMSu/AkP6DHbocwpngGqEvrfqoDRz3jRT+TeKplaa6DTMqdzqJWsGJRYHiNsStQyqL3xtCljY
4jRGH/o4K+vd6n6Vx58FGWTRjmAAUgdfFCrdB97xoaRnN1hWam4c4Nx70nnvnBx+dtzz6x1pbUzO
0cG8eHWUUvir4oNMWbhiG0KROkvJRCvLYHIisenI7uqxqRtnziYnU0+WxQSpReMZ/8kL0RgHeC9+
GmvSpcNVYLyHxHbbTdgSMrRTgx1UJRTYDF5BSZML16OxheeO5fs/Djfqy+nPWOgO9b79Ocz8Hi+z
NxkCm/1MdauNNPyAPFp9NOBPdH8Ztp+gtYTZKgdp7IY7l2NjFdnxM03eHFD53XE4MCjsTPOsLbH9
iutRbCsyTXyvj/NpzAYz4nuJDlIY0lGzr2QYKAZAbo7PIz6Wl/I9Byy9AQ9PIhHPbcXqNJK5DNv8
hVUpPMxTKx05M4e7khCAVHD5JXrVcOpODwIeq05Ty8AIKXAgm4q9EqDkXDNizK4k7lq5xe6MHsK2
siBLYKib39aCFFJ9DO7G5ypbYN8tK8DtOpl5cNzapVStJdL3M1YGKUZFZWINr7IwXp67r4ETsUSb
PHAtKhh1sDQVMbjGA+Wvb4W4xyg6t0PLkL6oOihoaS/lWkCEcdbGsPZv8uNikjgUkeUnB4zN9Nj7
Ud0yvRS4z4vQP3c/x5yE50gUA3Pfs0k7o7oOxbQtWCRMxt7GbKUchFuM0H0XGeWsHefsSb1NEVCy
IifHz1bUpWXIIt5Swdf87kHqi9RlNLITBQoVS70OMkmD5FQrgTxTbqdBWinULzivIKAAI+QhY1RV
L5BUT+pTfDk1vkebfq6yyzMPdXOukW2719IblbLbTDoF6Abci9FtTgEuw0l1WalQEFj4TB9jq1H0
I1JDNcNq/uE0vnwhIZEzEldH77e/z62K1UJxhM0S7H+vFG9japWID3TgUSFNYO0hF/yxCQ6ua+Px
Znh20TnGsp2x0Tm3+Bac8SA6HJYeHE7SjgVDU8tRnXZW2IdC7rM8lMnMD0ZLH9HaWs99JMAh8H6X
OL9J9RuVSvFTqvDDkj/lbSe1LThgA7BOOTJTa0GmArVKLsUHLXaxVzVvgXPb15BTyVqtIGGy+V4b
sF32o3HEstNgfOSSmxnP1qplP/0eYNgwd4UPLmQzv4LCuLRlIIjlP3kvOUX4tdb+CSsqNp5TxBS2
ujS77RKNL5g7hMuy493y/W7DpRffwsvUiuO1bhvV+/OeR2RJCcxmTzb1gte3yj+Z5ix9macNzvxC
YRo80hPSYfYOs4bFB6DfFHz/sY0rF6g379klpKzUrxqgLPldzAU6XGhsUKzum4FJh55evL7FND4v
qxZuqOoY8WRy1n3Bhtu/GOsCPKjxf8vgkEzUJGPIMWxX9bPu7T1OtdtHXaopj9g4u9bUOnq1JYmP
XoT+vlpICgCnNz0IRoa82Y2ruoyVXVDF7yYOfP9ykVidn3vdWbydGCYLcoth/y1DY+QahukeF7u1
0DJsnyv3MYJ+kc7gzygnp+jUFv7FKlKunWfHKbRPIahJ7x6z75zrHtCG0e0PCJQeauuh0XN1IbUb
TG/NF/Gvux4SjPyA6OTybrNFB28NCglev7o/2fjd+Ubd4iy24lo8J2YM69JaYRo1xcpVu6tQ6xby
Sn7eukGRKG7/+dKtBCWtHU6gS/FWmNQMTu6KCj9eztf752aXOeh+J4IoENUj5N326E/7GjKa13LM
RwJa6CClzq05v0McNCA1B6xf5bztgafapKVDjgDsRkooCl8lcW3d0GoJDIgpTK57BJAyc5RPkcXj
leNMpzS6r66+OUxj4A1IOYo81sSCXFwAWVIfp/7kPSY5qrmcag/NItysaPLWa46oz2QUwo/b4G7C
+mRMnmwOkQBdOSUZyKxuVjQ3lOMilyLDFGFqqoLy85NkmFyfTJRx4YNsLtebRvhgjOQhkHdX8adP
oKkErBaRUYH6qaXXxDo0rXxCRu1YzqQ+PS2TIbU7zrhspRZUui9CKN1ZqZ+e9iZzBJbv/XTHywyO
V8rOa8nDK/l7Tefw7V4L5o9V4DT8kkkMn7KLQSsE4QGHk16iHZVEWSlH3FX6xzYVPwsEJvzTVkwf
MEAuETTeCZDKEbn3DhEB5fsY6369PWB+HWVGEsT3ngRFj/PMWn+gKOtJJ+DzmY/ZkvCBc7V543/6
qgKEIeBe8Yi7Zm/4S8JeGxqHs0JX1vjc/RAHf31jUJu/2WUiuAxExKu/kGqzr0p6FGJFiLFU9klP
DScpqF35HK6xalIR44LJIzBi9soDjZXBnWcYXGB1EXMwNLYbJWMeVy6mUruvnScB2eyHp51dq7pv
b39sJ8HGBbSndhTbq4Tv5RJDnhViZ8234iqDMGpZfh3UlMglQAWZBtArdYVxDQsbFeAfegHZa2kS
wpTWXl1ao29Ij3knbAwPfPt4U+3jK2HU7ZZHTFlXnEBMUqXGKOmFaQU6i4SNxYfR/kFSCjKgd35o
z95zZBdj1TiApgfpYghRgFJAStfcNaxDFNE8z2DmrCqDPkxUY4baIZ7xLm1C/YqS/gEhK1qjPn7t
mXYL/kkQjTG16xTteQtPQFCNzeJQqSLqhmAZ8srg8aMtATg2Sko1IMerD6am2A9lAjEZsqmFP+Nu
9PYYh3AI8XSIsloPo+65i+ujBcWmQSmFyRba8VmgIpZOB2GvZkwdgXndFgr6rHC/e38YEPAm7F5X
kB5WEwXj/0lg8YOAJ64cxYTVdKtXPQba+rMXcbcQRCKSJlfGaZ4OAzL80aBQemwqOXU4GXbzJetn
JOsAHvChAMnxappnVt2VeuuCjBgkXD30iaLMbjnZfTEanejPqI6n7vibwKy4v/TRlZ0wsUkt/5NJ
XdR2bMwv1WgrQs1UPyUQnNoIcvZvyoXZwCaH+hXidUnjdJIFysUtHdprG2Qx39OxgZaUkCgEC2FJ
QDetGzYGR45zTWJv/oGCkxkkuFblFZQ1gXY8teDtirEEbKK647aNqWw37/HewzVz4E79O787Uq8L
COJvwxPHspQI5Re162CE+yUdpRenqolWhPBNM29As8H7LPIJXugF4OTAF3O1+0br9duAiLPDMBkV
K3u2lZto2tEeBK+DWfriknwKuypplL7FJ7LuYFHE2ZYn2KfhkUuREhF1+16CW3i6vz9Hsm35AULH
lHdEWpTbyZE4XdjZ/UI+crKBTZVJ44+94iuLRoxBPbEtHtwX14iCQkON4akUEixTn7z8Lch/wX2d
ReTxNLzmSyLTcoaw3+YL8OoWczWTKcbVAq3Oe2kjy5gpnVrswIyIWJEeuzRRl2ys2Aq1ZgQ0iL1C
LTPKVS6HA/D1/UYJUJAewWVBlvoa5pvogwvh3dqSQl3o52x4NFo+gG/EZ+OmZ+hIqzdjNXUZvYor
Cu51HDXgF+/cOvHcmoFLk5CtABShKPfMei3Q2tPPOqL/MvkoGLbVEdftE+exFuelMV3rXhU7TBBV
sx8KFvc6P1j4/vBBxTiQJSxSbJZBE/szeqR1o/svWR/ti5xURzPWEseCrS2H/7eFCLYj38h82gAJ
TlYq2Oqo4CAh69huIghlLQCNZoRuyffiC6Y9JR4Iw52jQoNUUsaleOp8YVTBOUNw597BjB3nOHr6
ONV3b75113NsgKVhD8vMtfYwlj9GqQ0dRSiIWGX8GsjDaGqih6qlQFw3XbkiVklVwSi+4haRmJuB
+9Owujy9RyIjDTN/XIPh92pjGAThMc68MZjoxleV01ZMujU2INDpaCuYoNUB5aZymYPXVv2Vzd9Z
lttDAcWKnXRHixL+RfgbM+4O2uno/Y1ZelD9LatOqwbgn7J+F2XWC+pmPVHi38qBHEm2qbAsL6uq
VLyKxFuzRy5IP62ykKMxSBuD2o6t12u0MbPRBe5A280Ak3e8maqMtwqG+uE0DZ77umcrPvJma6Tq
JtXyznpxVB5pwluFtVCWO5SzZMfPRkqye30DZAEb0faqoWjAZW4CGXCkSVRfpdRgRdjAbYxLubWV
dtYvDQQR8RsTvfPIBtdENFFqHF2PtdT061wDLTCW7h20rSl4udjzKB4z710tt5nqnu5IsAax65vr
Z5+paMtS+MBuPE+Zn+xeLMyp/pW0jgHx6mDQIipurL4QZxgoShvT5ML6VrWpuTd9n65UE6LgxVwj
S33xPEXFd1/2e3rkU/KCL/lOr14+qgx1r35kQm5t0lpFTQgNbMoxUMesxT7dDDpy6/8pDB6Up+S3
S/lw0NtcaroaPXkfwzpfwhWyLTaWgGTZ0yKzU9QEu7Yi/GoDd6otmrzKwQX1ediVYvKSPblrjQ/N
ma5TelXwfzClJL3urrjhVtysw22E7zew+GE1AoNqZv68b0nBHZhoWaFnES204VX4PlJn6hJcQ2mP
FKPt8+RpFXez8WuSywNLyFHp30oJ4vbcEMfxWaI+gqlTwMtG8GbuWS2n1uO5iVZ3T725z6stRRfi
fF8a/xRUcglo+hFFw4Dx2RZlaLOyURLTiVn9V+1qjl0rww7pE5nQK5guURtMCvYetcYEsYZxG7L7
aOwI+2TNmeaEoMm5yyO9JtpQVIxMe990JJ5hjL2Z2vx1qALyy1EsHMfRPaqv8QeRiBxyp77tz1dN
DI0Gan42p82noInhbdFY39iw6y2Y1VzEOpvdMyVVPG/HpT4J5OOoOAgx2WiHriT9LAzSFz4mUAvx
kdHA+W2m4+uooMZmomsejti8Zc5yqmcu6xChX6aDDAcnzsLz46cszxhQ0jUd0tA9F7ZCtCegLELd
UKqq+Tpo6whShYg7ZSV0MLa/p+iHEJMghSzxYld/zJevaGF/M8nOkmO3Y0YQnjkUYM4XZ81tUhGO
Q1Wq6VHuInkw/H1QJgmAYqh4TJVxXqiCDuTE0Gvd6YOkbAS4pgB1qlUt+OMryFMYMgM3ms0slDH/
hFm0y60rkMFR6BvBDs0rYCvQ4S2xT0kiiiFWDNwm8QTPFGm5h77ZiaL8NkkbkJeMsHJHKeEYJKAt
w4mAsBwXYe7ZVpgyQVLoaC16jiB6cCtE8/pX8b/PlWATIruA78KCV6U9Z3HsPg9HKr2xjmBh3zK1
M/PMxCHvtFxAUmYi/L0puZC9icSbOe/Pw+93GKXWO/xSemblH4M0+A==
`protect end_protected
