��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$Rx�y�<��wA�*;�x���@�̦�W�X�fa�M-$u����n~�%���P�$��W��kYَ���P7�?UMfT��q�6�U��k�>����~�\N�(�����X�e���/6U|)�X2pF�]$h���d.���9E��WG��L�X"]�Ad����ľS���8od����e�GT?y	7�������ݵ�^��R�q^]�鍦�����s�ae���h��L��P_���ާ��YЭF���'\��68�b�[����w8�[X��V�F�0͘3����q諵�uW� �h�u\V�?@��_6G�_�*�G���B�絉�f������[�G��U&�����~�F��AׯK1�`c��[<��FY���4I� �#�G��x[X�=�Q1��`��R>(�w����R�O�?����7�,(�H\�#h(W�EH=�������yq��Ѿ��aF����:�U~m<|��.��0=�P/���4ǆ���T(���IjS~���2F�k��t�"�����x��GI���MA$QK�_ҥϾ@0���m�q~`�]�N���,��6�YC�VoC�V=4C�h��2{7j��lj�+���I�k�x/m�BX�nH��>�R�;�|�]�o�[��j5.�gZ�~<��a+��I�P����"8�K/K�����<2�K₲i�lg�*�۞��A�څe.�)j��QЃ�;���T;>��U�p�+��rj�H\j�I2��[�\�Qc��=�j��v��˗�-�0�{W�ÿ�ɴ��[����B�3���JP���
z��1��M��!�͟>yt^ه��1Ά�~wTdHE�f��ڐ���f���=b�ZzF��~���@ūU�$�u܂�y���o���xL�*5��g*N$��0��Ab�qy����39c��:�?l�+RD�w�����+1��l�H��Z]���ɇrs�A�O{��t�~����xf}�X���/h��3� _}	��Y�mC0�=n�J�Ȋ�F��^ɑ�:�*s�=��| ��q�ꆜY�ܲ�b��(+�;ۼ3�Վ(xB6G:���U0��&�1������;	C�|Ih5�J�w�tK������0iKk-�i��(��d��bz�cE�0��V*��#(��nۍZ��y�������:��z�l�8hk�/�������۹E��=�\
��0 �$8�ܜ�嫭ۃ���d�EMۂ���l
J(QK�*�6gB��ڍ<!����	i"�e��H��ڌ߃t*����X�q��8S�OW�_�4�D���#>H���|s����ۇ4nG:�9�hN�	��^@�js	���n���*����bo,<E!WFĔdI	��*
ݹ:.�o�]�1�E�P�m��Eg�ؖ]}0��^�P�Э,�lxË��^rB��~��)zwY�9')>����U����t������;y���C%Ks;z�t>�R��t�����F/J���z��C
i���#�.r���J�^���[�Raܬ�+h�(8ڏy�3Av�|5��D���<b�Z�<��3ȝ�j�㢜�	v;��7oQ2�T[�6^�ƉY%"��5&=*�9"tr��de��'dg+���[����녑>\� ��r���8����ZVo]��9ϻ�S'|�B���Cna:˦�(���A�~�ݖKX�?�jȧ�����T�B�tZ��ӌ�\ݜ��Y
�\��t)"ڐu�b5/�P���r@��pqR.��vȳ�%zF��xRNLq�T�� �%`v<�3�O�gN>����&&0���K��Χ��i�C���nc�$&�a�^m�Gy���'5z��y��Xuا��Tz��^]$��goZ^��F���U�.�����[qvF��h��m�/~�󜕌������w����i���I���o���Bf�K%&}6�_{�Dq*`H�@A�no�*���	9��`�^�^�p��5e���+ÏL�L�0�Z�޹���}���'���=��?|6�;R��RGM-��H^ө�Eo��I�F}f�>re� �ޏ &%���,�Q����Nh,`-Z���;�Q�һ� ���c�Υ&�m9��
P�����<��gP�<Pw�{�ͱs�D�cӌP���+��H�'��w����5ov�c�|�hEZI�s*��-���b���M��/����X)�����	)�WصX*�b$�Ȱ�]��\�x�l�C�*A�2:�r!$�E�321�>c�@��ԩe�l���M��iQ!�1jm� �A�<-Q�+E4� �{~��AS���⢷�|��,��n涉)�xj{��� @�8%ե�<m��3��8D�:�v�a��}��Y$iSi��;�[�� o�/l ���_��(*%�ߖ�A:#�P[}�J����=X����!qgG��J���Jl��,��Q��e��e�D�լ�:�_Ɖ��A�)Z���R���\	P\��DwbGDP�J�f.4��yM��zA����E�\�8"��&�BY�+q��Z<�a_s+�H�`�utW�&N��Z�x�P�au\�!!p�Ϡ�R�ZaM9�G,�q&�L:r�z�����ڐ��P@���_�3���y� �W}�-��J���L����H�FP�>Ϊ��6�S��x�([���`�/=?��=^����H�ip�����[�L���릱�U��c��r�;E'�:���	���ّ����-Q�(��Ŭ���\� +�/RZ��B�%w�_����2z�M-מOazj�Yb4��&=�O=�n��=T-�?�n�i�^�?�3 V��R��7ܺ�,�r^�@���Ω�S}t5SQvN�,�ZID���#&���8">����?�	�v9ů�B�"�֦�d�N��y�s�=�t��z�!�H͚�4�d�#�-h�	��L�s6�w����Q�_�l�L�a���n��.��R
���:��4��\��OV(�-v�z@a":j��F?�>l�v�X���/Ÿř;�T����^1B�fe��j��8���-������U�����O&�/4���Ybz�HѤ����%�k��#�!��K2\�-���吐ZLHc6��͌�̙{nt�̉��ŰP�a�_|�S@��ئ��������d�3�I������mӱ�B{m>*V��-l�[��}�D1+���9�wx1�}�h#��ӆE�8�Y|����Ա�5��$2��g�9t�%=oh楾�� .+Y�����9�g�b@�w�C,h6Cg�Y�� �2À+Ŭ���Ǆ#)��|--7����c�����<���
��R��a��/�B���6�_���T��)���*�O.pӎ��&!x�V��dF	���+��ǂI�����\���?�������(K��G,D<(��z?6��`)��|�֜��M��~�!`͋>Ue�RY�6�mN�/�_�Ӗ�4���b�@]�n�_�B�&��v�����va�;��\izt�|-��RƂ�7""�������~U�~�YOҍ'(\A�R��^�W�ˡ�۸�b�f_*�"�Y��᧠b��Kx�[ ��@��_ߦj�8*���1N�d?�V��2�o�쀼pD�"���QƓ�zȪkh7h*ɼ��:;������{��H�˞��,Pd|P��}�k���"��X��qڋd�֮#|����kU<���qP޷�����+��¶���1u���8��X��W8��ї-|�����5mp�F=�a��h�É�D\d�a�cͳ-�j>��?gZ:_Z��������?� �*�iw��b\�L�۷�X�#Z��J���ZOc�`A\F �$�����8�-r'D���v}��VPUQhq:�3��H��H]N�_I������	fY~/����3���/�R��:�ݲ�*{ ���O�����5��_��dV�Q�ͨ��\7<ц� ������K�]1��?�D���¡��r��{1d�k#�1����2��ƃPn��@SW�#�Ƭ_��r����E��k������e��Ӣ2"���#ɋ�͹�|ߝ��b61ąe�_t�Z#�9��>�G�hB�G����z�զ !/ M3�j_@2~:���;߽�[<��ƵR�Lڡ�gW}�<u$o�E;]�%�>3�r|���*��z᷐��h�`���SoĤ�k������}?u=� ��eC9�����U�����}t�2��\���;��1�)�g���&}G���՞���n�N�Q����b"� f唎&˿����i^u���U��C3-���� @��N g�e�]AU�A_�Te�1�x�y�ڵ���\��/�S�e.قdF#l)��Q��x5�g����.���3(�`�{��?�5�;�yJ3eh�,@Ջ��q<�)�C��bm�BqQ����ÑY��i�2�u	��%��E�(�����u:��4g����i�K���AP�N)d�(���@��MS��Y㾎A@?�ѐ�u�G���Z��Y��w�^�ȹ�|ٵ��``�d��{;f�)���6"����'?0�B@�����ϳ�1�*B��_��Q�+�:�\�����:�'^��a�(�X�y>�$u����c��q��3�����b��y5&{�6���#'�ꢲ~�>I�/�re��X뽞�r����.��>a^��V�& H�cB9*D4}j�cyQ�.v�1��t@����vۑ��؈(c�y��N�⛿ ��.9��2;_���]>�N)̰��=�(���ػ˽�����T�l�ows����-g�q��x=|�xНeb�ּ	v�4�{�+5������C���I��p��pf$4��ý�x�����q&8�.Px%����QU��+�n�&�8Evz�IzN�j��߉>��$�v��/A��i��/��k�fbe��@���d�7e��S�I�H������:Mf��>���a|��&�,�A�4{�L�G�+�����b�0d�B�lSq���W�d>�|�@0��0�s��׃�-�qn����<��\���� �
H^�j%
��[^����d;5��,��=I�J��ƃCb��J�p	%(�`��-�Y9u���P�ܬ�3�;��}�����1҂;��?b[��e)���<�*N�8�3��Q[$u����n6��b{ ��a���n�H�HN��\�Lb�>�g��W���g�<��C�!?�:,��P�U\L�%���\S�K/jwm�Vy���M�^ܢE�v����p�+������=�8>�<C� Ք0�q5�\�ꪕa1ٗ {��Jo������L	W
�"�)�]Y`�M3 ���t
̾���P�8��s��v���U���S��&���(�����h�?�Qy.��"��/6�6���"��{O��"�9-a���v�" kҹd�Gk��U��䟈P[7&��Tg3��/֏�yp�O�<��#9���	=Bp[ ��{�p���I��+���ȃV�%����ӥ03U@��C�-�>�ܣg����H���/��RfjD�Un�ֶ��� lBF?�#��4$La�)�+�u&*l����Qn��T톍�w�gON��HίQ(��~��=�Z_.�Dј+�n-�N#����eK��]�>����Z\���(Y���Y�i��zb�\�B�@qH�����{q�V, U���YIw�^{�z��!fh�s��\s�_��4]���Kc\;�3���Py!k�bd�;+@$���,���#V��g᷃�0^:�G۰�ZfmSѷb�VL%z_S��2���~t��ٌ
A���Y�-��sq4�8A���[�60q�ŶE�SY���m2�/o����"�6�1�dԪSh
�a�,�I�?͜�  w��FQM�fkr�Tz^8ss��/�qc�\@�n�t�5�|��2����z�����+�=FU	�Ƒ�D�2��	&����)=p��|����s�_�%��h`�f��W����#~��!�v��V$YU�ef¦����*�S-���z�H�B>i ���5��$��o,я�<X����m��ZD8���5�t����� �S����xjL~�6V�H�d��\���|��/w�V�9B��C�AK̎��➣�Y���oOK���
i�@DahȚ,:�',yF0��>��{��i;�]q�aBf�k�$�(�o�����j��)��Qˣ��x"�tɈy�[
�0n�Ȍ���2W��yØ���j�"Y����1bIQ���������9�`ڽ�sg�RomG�
d�C�=�~��Wg��3���Sٷ�|�<L+��J ��b�%��<�?�dS�wn{,{sSчb��?7���g�J�7����t:Zə�m���Pn,��ϰ��}K�G+v3�
E���������B>����\�o!��T�I;����u��U,�����Gx�
K{�L�B�r])�1�&�W43yx�K��1|�a���P)��D�tO��<��A0��dfZ-$©��ײFs��`����5$���+��/��l�nœ�=�d��Xn�`5!�,N��@>���� ���s7mJAjF[��w]g���l+��zn,w[(@j���7Dd��g<���[Vx0X�w�[C���+JJ�e	����g���Y���~=��p*յ�5l���C����؟�>K �1O�z��c���T�b�����{��
At3?m��aB�&:g��bug��z@�L�~�X�\�\ϧ@-GwѴZ�@���q���G&�Y�'E���H��3"����(�r!J!��{�*��V�l6!*s�
�����;;���Kʧ}��{kf����x�˗�~��(����Vx����{C���w��Xn��t�Qo�]2�^o�t��Xn����t��\��$1����K{ZzR������?=��:��b��
�-̤'�w�6(��|�\f�@[O��pe<C�I�k�qb��5	���8���m�K�,�1w&��LC����@�\}�� q5l�
3�]��P��LZb#�˸�Ħ�nθY"�/rYd����=}�t^��W�u������6Ť��F���W���ў~F2	��H��)�����.Q�q���D����m[���(�/�㳯3�8s��@��l����2F������HF;����
S�,]�s���3J�ÜI��l*�R�R�T�M���s�uϭv�͠l�����H?��yE;��0���6"{�:����~�`��F�>I�96�J�D ���{eJ�Hr,=�/t�����nX��5\�@�j�RɃ�Q&@��"�p~}��1�J9~S���9ڐ�͋ȵ��G�k�f��g|l
�����R:]��\��x�Ϯ��BgxK�!��D=�G�����qֶ�#�d��iI�p�$�Q���>�Ȱ �"��>3��r؊X�D�sQ��g��4��v����4m�QE�5�(S�/[�$Pen����1���ä��OW�ۚ��Y�%m���`����	�F���z�(�ʻ�Vt�S�vk�iI�Tq�>��FhP3�Z���O�]/d6�գ�� ];Ɋ$�`q?xKie���֕<���57D�K���Z�D�l�Tf[)�C��(�vO�:%
�r�rW|���qt�q�����	}��i.rs_�a['�w�Qa��3j���[q ��v�/ɛ+��n��%�쵣��l���oj�Q����A�q��;'����kF������NS$�۞�ժ��i���xPQ1YC[�����;-���l�*��'��7�K^��]��h�vL�Њ�wG����y,C�Q9=�U�fG�Z3V�tH��K������̖��U�۽��(6���~���70��^Tjq=Gl�aA�p�!������l��>Tl4H�ޙ+qZ��0"�����}X��,��k�a��~\��g� �#�僚`��D��ER�Ι��*$�:��o���t�"Z���F�q�x�R��XH��b�y����UAЅ`�M.��%�2Q5v���$�N�ZGˡ�����B�S�E:o����%N)�.-�z�T��g�Y����3��0���Ea�A�%;z�׭y3������koc�"����y4�^�R�^W���S�=�미��9�~`aG���d�,�;EQ�iX��*����n�|zF�f�.,` !�
CԷ\üMl��}�;��j�/�~V��)V�N�JT_qWg�R��ǿP�\�N�1S���/b�
C�.ק�MYKA¢T!`��
�� ��_�e؊m�S}>a��6l��Cլs-�b��������'f�N��j�t
Z0��0�ާy�t���jق|��O���F� ����e��E��-VA�y�e�8QX�89~ȓ2M��gI�A���+��|���q$4z���i���%ޅ��t{h�=���?���h0Y��C������y�"zA����x�JE�۟�} %��~;ڨ�4�0�I]yk_4{�"H%U'�sp-����������ׄ����%x��C��C֘ޭ?@�O������LC�G�__L�.[�ZH��$��/�!ż�ak!%�������Z���eb�ߟ�iT}�K����ս}
 l&�\��x�����c��SB`g�T�eE1��f�z�_Ͼ�)u-Qa�|��5����G�1��j,3�Ф��T|Q�ݝA��Qę�#U��y1�����D��
�����B�C�q�HЮQY��F�\-�pf�Wy���u4nc�t��L�P��@q3%�@ܰq�JU��:�/��W����уD~jS9�.Gp�?�5#���2�:i:��uc4���#����K��<���QX���i�{�ӼY��� P@	��)���5���񙾆�V�EJ�F�2��Lv���-E�k%����mʂ��m�<�ʖ4�-I������2���B���5okm�X��ɫP��o�,�q�9� kH�n��5�z�%d�Y�^�Ys��r$�>�/���5,n�?�����m��gv�a�1��=,��'�_$��Dg� 11���T�M �=H����?J�ǻF썾��rx��G�O��|�ݝI̶.�7����vJM˱
}�V�}C��1�L�^%̲����v�͇Խ ��y<��|���a�CĜ~��#x�D��瑍c��х��)������ʚ���p<�<�� ��fV�V�w���9�X�-yU���Al#�T�LʏOB��p@p��?����on�W	0H��U⯜�
���SB��"�,i�-�1���J�Y���T1z~�����:�j,SI��@������2C��taH��_+�!��b���fbT���+�/��g[1�)�҃]7#j-�j=�?�!�TwK���A$pl�Rw�J�-f�B[�k� �M����;���d�AU�eU1Q������?�x
F�P�F9�b�חb��`����ݹ2.υ �Х�����	{��u�ͬ{lT��$�CZQ�*��6p�1V*)�*�!({0��uk�a��0���1�Ǣ	9~�W��m=������j�U�y��Um�f�x���!g��)}(�;0h:�	a@�����P*�kD�=�[��_R��R/��� ���v=�x��x��e8���Vq�(4�����)GXɱp��4�V�d��Z����������5�}]`j�����R�,�$�U�@'?����z�܏ �Uīz�/)���	�x�~��O��)�	�1��܂��Z� ���D*��+/m�ѕ�z�A�D�<�$>A+�9�u�	��]�;q�K/XW&e���&/� �<�'4^̧�H}ó;�����S�6�z�.v$  wq4��c@��@��,+��o+��*��i�z1i�T�e5ߤ���?���7���u���|�$	E6�x�E����a��m�>c�q(��nv�%�c��޶�N��t<uu␙�ʚگ��%YR�����MX٦�ė'_���e���@� �8��I�C�+�������P6�����@��)��?��_��eJ�T-�@�
>L���z�'S0���$�8�8�+���!�&;sD�.S0Yԧi �//2`��?^2�#0��}h
�m�X1{��b�lD��Z���|{Y��B�QP�H����5�NWz��/!Q��{= _��$��<��@�ak�95�Ģ�MI��]�Y$>�g=x��Yf6�Sg�M}hn���@�|�o	�����Q]�Ŋ�tiC/���'j5
4�ʉ�H�;&�DOL�p��^�~a�g&�*+y��u�i�M�V��-[Di����V����M��DL/bQ^T�t�hQ���hG贇 f�Z���VZZ)"Į�7�A�ÉW����.�^�_3<�� (c�V�f�ݳ�*�c�O�Eo�n-��+��K��P:�ٛ�,��H�$5��O�4������l� <F�3]!�8��j���_%���8�4]�D�up{I&��Z#{�H�o�Vޕ�_%�Y6�Zk�R�|��m!V��"�.TL��4����={/q�v3�K�[{1��5ض�0�<kVߋ�o��ȵDwH�����Nq� 8�w)PR��w^�����O�U�[��=(;�]W8����
m���6�I}�b���K#O��R�7A�������Ʈ���3�,q��c��v4D�*�-���fs�w-3���MG�*\�h�s��J�Ei������j��9�@��]s91�A3�
�e,�\[$J��=�
To�L�_������HRz_7D�o��wԆkr��r�H�q�D��p�-地��q��v��H��4{T2"���d����S�ݦ�lB�xM�=��L�*���[�-����y��}���1ڊ�!F��]���-�x��DN��A�J?+��r���D���/W���y�u�8KM�ZU���jv[;D���k��R�**�(aV�CY����Km�g�?uW��w&T��c��bMڨ��|�Ѕ��Nҩo/�S±��������j�v�q�ɀЍ��v�����릀�.T[�ޮ��%{�:�V�v�ɍvEj��#���j7�$,�*�,��}�W�ݒdJ7U�x����R�n~׿�u[����Y	�wl�M��g�X��z`�N�<��%L!D��聚�J�y�柴k�$�t��|!T��������Mak=�q��)O�w| }�M�6���D����v�E���X���<ɣ�_ ���~����d������Mj�/TJ�e�i�8�����<R�#m!]�q+���6v_�Ve�Ql/n�N��P���0�5<mA��ݟ�wT�Ċ'�g%��W\��x��%��P̳sʴXN)TFK	�s9YH�A��w��>�4��-�ׂ�j�L�Y�b>$�����oR����IPa�����k��K$�{�vk��s��������w��r�Ea�P�Ѐ؀5|���#Z��S�$wa����-+�UD�!e�Ԁ�/m�Q�`M�T����>=��@��~[U�⮚��(�I�'�� �� �I&BХL�݊��X4���ZDц昆��