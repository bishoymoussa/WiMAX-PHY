-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
zX6Bwovcb0QMnI71D/3i7PX9k15weC28oqL08uDrIELScarxs6D0PFslztDfONikgmFck8DgjH67
X9huSLCHKOlkk63SwCBw+eBjkOGIxm1yN48AHGQHeF+AV3fFL6Emj71wubkcV3A0dlq/HMmFqBBu
CGmielUeY8iO9HuT+4uYzF/8ERJrAHubxIIHGmxP9NrnVzUllqWWgKFlL9xbvsDQpEbyf11vWVT0
kZHnZ0QGRYjPr45/i5dQsclnOPegocgmfCrLGUb8WntMWWy5NURcOZtlsY70rum06AaUdJdCkiuu
kibv28NfRVcaVJnC0UW2eIHPFRj/05u7sLcrTw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 47136)
`protect data_block
czZ+6EnBraCGg8A7ZFozE2r8qjspL8N0oPLCIrEm6wz+E0fH2hW98mJPAVsqjsLWqcuI1X3j4roE
DzZn8vmEKhJP5s3YC1U2ayShvLJYVTxY77+2tieTUpX9tTvZj6VTOj3kUj7gNnDoboKgewqhzQSm
5iTQPH5Im68z3rSWMhn5NW2Z1mARp0POiK2C0SQ4QJ81/yo2AohwpLYDmlGp24Zcl5E14z/gCxgM
2hfdbwnEkMpn4PZLulr01/0Dk07Y4GJzHfbMrztWWU/yWIGIoT4G0cZConb2BRNaI1jcARkVvTGA
PDFmw7mQ7zN8ppLe5CoYDND/RNicaIZbDKOgL3PZ5kJsmJU7JT3N+lYrixQ9s19qtRCI3xqAK09m
W03Bt29WbRKNqcI7S0hzQQAK1JPO/bBl9/3XztsyTsMEQoTuE5aen3+bjQtldw9Y+7vbBTbxHjX2
X5wS42OIFjDhEo+aj/sPqRKkQaxwO5/JdiSYTjgdCZzr3AJBU1h/6m9HutmfQg8YKfM08xhTav1w
31pT9BMu7SOFePKvwv0xCWK9ePYy/I+dwIYixJFqHnAVn408lVk84lIqupIGcF1gs7Q0VvPL+rS1
XgXu+SWJV7dMHWlcJ8/QIwgXafusXUQFEgyBbLyBhbdxy71bJRYTrglrq0BEVjvc0ItXj9emHDNJ
mb252RuHECcOJcHIq/2FPGJH4IjN+WJKUUQ5Jvynr7jcyZ6rxHILG6dJtVFIe1spj7FnUkm+3uDt
5MwfcRg9CFitgVSg0hdxVPdI2W1T/RLzQcDRKCndTxgQ/GnZTkavcyYI0j3PCLhuIHO1j0hlFlbu
itLz9DfuQ/OvbxHfxHS4pixq59FrIhgcrsNIB5+yTcrTwhrB3N3Ka2VtsVpfWjUK7ZeBjiUuD6OF
01Aqycd+yhDorIxHXgWGYSGpR58fkMjp3IWyNN6XKegklMi6tKZ838SUv1uhZems8BENHLlLiaqN
Jus3+O5DiUSc/7D7oiPQ0pLGF/NmCO7EFWe9JPuc5nb+nBO52f3O97KG/4k6tOmpZVaiP06qSi6B
d+JYpSQaw/N5z+Ar7IAM8DTRsr/ZyxeNp5iweFQK3qscHkd+K1QT/mulasGYivgCcBe9ywM9123S
QXKgn/VJikolW8omISF4sm6ZX1iZLXAPcrNEM0pvls5aZNKDjCPDhgZlLyIpKuurc1OJ0JC8/RVZ
DaEEP4Dezv49fDPvrs/O2WgbL7VU3M4vIbhbQ9MRxwJOEiwdn2U46W++IQsU6Uy32UFzRs0oQDds
KcNPvCKP0Kl1D+b6UxyOfo8Ow6sF7NjkzJf7qph2Lbk/RxsthkTHTAxph/MO2RISYXrs3+mXYacu
q/aENOyvlb6vkg6qrsH5r171QictGGU0oOlH44lMf0+2wrZ8MVSq9hWd8FTDyeK3Xy/qi1Ivvbky
4H8372tndO3wMNT/m1FGcMIOwcmADcs0lZETBs2Vw1UFcaGu7+PB253CApX33cHxZXuSKA/j/jRY
U1i6LqOg7/phOqR0IpA49/gPVGqEONfoqITCSvodZrCD+CrGnVAQfVz+XdxP1Iib0287GHGDKhIr
+JWcyIMlgv5IiflzD525XDY0EQ1uyS3sl/K5rp4XD/qZbWC7KkjtRvHXIRl1jMDaDXVmHZxiK+bn
TGVwsAYOJolWVykebOId+Ad+ZsVuf/TT4hFPBfaukCsKVgblxG7WhjzExaAn7RVZmTCDAIJMvufJ
7XvBRELlicnWJcYPvh7oKNmpfKBW9/93A4NjpuxQX6mRDOH6Pkr6zxgUAcawQaAkBjeEyaDIisvF
Dlr4x2ec3Sn8Cdu/zKnflypYZxqKNvZg6lCEoB8kc/eeMF7FAZKTeA1ZMczkoe9oSd//rju8u/2M
HsxVcynvdTwYb9qEb7q8FxzBfVPelfYhfgUfI4s/sDg/SZAOJO1QzQlO/TKZrjDOc/HpTujcU9AI
rxElSJ6M8pvKP+wdTPo4LS9pUn9K3rSi0D9YYYOsLBGORG1pe8WmZxMMkb19147xuaMOZm4+z1kr
3Uaxro+AVuA5rt47jmwbaaQ9pHl6ckv9u+7OUDXECaMEAfrpignyCLS5NZr6CRx2SElJAOBQQtwO
uQ78oC/TfsR8I1qXLJ6xIISvrnT6V6d0qjQ5BnW8Bu4vRagUQTCdvC1+jVsVFgziDNM7uHmeowJL
7IhQIwnFonFKrqPxDkfWxvOAXJSc3BhJtRnK1G1NcU+a30DXDf2iKrL5bZg6oyEcQ2i5sTnFWm3e
0agsBuKXxkYArw6WL9f1loPx55Rmpayb3sSwRuGW3jR2HWYPA9pZhcYM8i+ChkBFL4N/XIhLq+Gr
yqcZiOkS1Sx7n62jnvcmyt+rx2jN84uY5D+nD++xpPcdrK/ymr7gSP5BRkAGLK+j4C4H3aPX+06J
IyRDyt2iXG+UEspIRd2NbdTlyYM6FlMlL6g6DqivVoaiDyQc0tcT4WleBM5Y6XsSKaVg31XTEMd6
oCbNPdj6X4PeWWcs8ciIwcpJzhVF+d0AZJ9U01EOEglgy2RMuJcmFpQkJfAiAUhFCeKFVjc1gVF/
6L84Hn6xBFwlieAXJr2a8QRqMtamSmK4GB1vSYE56Sxi8NvcKvDUfsGELxVWJ3gylBqwETmRCQot
1jzHyKoJSlmi9A7BqeadA17CKaKb6TqwZafI06H7fjGyBu4jsWmvRQM6MY92HXiBjr9jQHDGdzKt
9EiK8d6iUwzpC3c+Ys56t8A2KguXvceYdS5tDe1gKmaHg66UtG7N4SD9RfXmZ7MF9e8648Yej4B7
iGe1lP09uG3DAHSSj2z0xfk7nN5u8gkrn4J8PIP4nH4pfG9M7Ybg8CE8T30SV+iAGc1RYNnUMt/v
MUZf2Q8fw0kltpX7hzsfcOyiD60zRE6o+HiooS6eIl6supDjpwa1ernbSnwW3WsK1mhGj2Pk7fEv
gBtDD1vBu+OV0QGcDXBbyTNnhSU/Ny0Suxoz0WIa6ETOeW57gj/Xo/AVKlEmap/UAs5eyaCpeyBQ
hDbtqhE3n1DlcymgIkQADKF6ISMsb3lWKJHb/BAURSN8FxdBsOFoNhaCcjeyuFi76HcxArZbySTQ
46nq0mK//yzIyg8ukQPYqA0g0fiGNoro9hemP9maeGxhrtBNYbPLhYHd5YmeY45Iiww7q3ZX9PkF
J7XGqbnWlFe9h0cDlxSDVgs8QU+06VfxLi5oAJTdqFXs1o99DvhySf9gFxPsKLtaXjpZmPFLuO4D
ur4PAtOsY5w64u37scm0EmxKLeAf339sCkyGR/8XjdaXOPGFNW/UfXUpbsIUo8qMWdxZU5cqzkUR
YMFDGwLQVlyrRjhuCg3F8ManL23hjXLgunAruvvK4kUfymZxjbFW8iiXiH2x764jpX7MBzq7lpW/
UlmT7E7taqr96QWhwI4aYw71qQ7lCor8aybMcZcFN0iXUDiX1OgdI2xnJfIl+4uKsP1P9nfnhWew
+dDUjc70+OXQf7CU1AZBVBH/WKmf0xZwrg2GJczTTx4Wi4wRkRC3DX/fh9RsKBk5NZXxlH1m2H1+
0jkDWkOO0oCt3QaqfbBVGI8AVFc4j+PFo6udku7uIlCvEBUp2+LPHFY7JS2dtGJ+eMPfF+BiOaA5
3YB4RoOhkXiDOnr0S5eTRgqNRsrNYfqZBd/tyVD2+xlwrvHQjQYWKcjg1I7sfGCoY6W8pXJSGW0r
7MuPH1BaluKFSmN7Al+mg2im2emvD6gJ5V5h4Vc6qtO5XqVqSa23Glnrk9DuaRhT8yV556pq/gAn
NmIPy0+chSgIlzPtZO9z+EICy9+C7JfVSmLApz+hzMWMGgI0XyvQe/RJzYDGKj6ZiQuXbOtQwJPn
94BHkSZ4f+RZ1J4mM5KbQwdI30VifhgZYZVM3B9EdHNYXreiwLng68uQVn+JZSxvGVteQS+bz0Z4
x8y9zhI04SM4b//0S6zt6vOE0q0YKApQI2MHJ8yeNHD4Cyd06qutChAyOsYqhX7utIYmEAm0tUkm
hyFCLBlVJfIf0jAxW2QaygCa0YTE4999+H/B3LeuFFGPzshkDfcdAx1h9Iqm7H5e61AjoraUnAdh
GrGYHd/9LNtQwIVcmj5+xLP+adf30R1EG8Qrg7FFsl463YfQYxaRBSQx1zgI1g2KkMVvJjUTJPSl
moSO4REIc4T4tfSYLyNhb1079oAPJOwpKpPVDrxKKrjBCCLWkh5FEXCpyIF5zqMt1mWXP6LPHDQ5
GhcPC1fIVP9kuZ6hYINv5UOgqImLyxYkxn/gCLhVm52A5riQDKAJtSMrXcplsjaItAX2QMjM2ds/
iItqsV0Ncn2QvarY9+d4O0Kquhu95kxHqE7umBaNjgZRfyipSe9Z6FiNK6ViT54/EQ6l/5321XCU
DrWhTjvHa/cBtV5KWquKNM7QqwXwxA+aII/ai6iBgjduzM2Zm/wD9QPwbouSTbEJDtnVqQit+E9I
zpFfQaD9uk05Exm6EwtdjV2ryAUrcuxxaU4mUbtE32XJ8hsHALYOQRVtFf1LNdogYuZPeq7S/CvM
SWBqItbtXRZF/FnjIvcgOB0stqZNV8tq0PBmt6FWIcyD3Nhra789ZRcK8P8KO1UqRBbVNtLvfB3R
tR0kzFdfHPdA83kJhof0IBlXUx9b7ubNHEYq11XwiitfgIDlvfK3SiAFmJbFurpAZck4IuC8oSSK
ZvVAz1xdo6QHomLqRpVuJXW43QzVEtylPnKJYr1S6NOCMIZFTLWmQxaBrBK7sqbvGC+afeBOY3YX
+vRIOU9632dJ289n1s7drSu6nNuneyqjS17MHFV0HXdLWxMUoJcYiA+VbTDaCz72hDzptGFwIwDQ
gSxGtW1qF65t6YxkV/KVjykqhrqS7RnyzNyDtYzSs+VtvoKSSlEfRtkQen1EPDxLl2Yri36gh6xA
NqGc2frqDgcMRBhj4p2awYysRwebQfsKJRvlT6H5s4yfngPc9WFi+kXqOtXCPgmhtDvRggfHfMZg
kBIO9mhvUpxcJBu5+b2VC8xTyJ4gVjGLcZdfyQ5yvwS68h3FsHfsOLHWGijw7znzeZB3RVl8X978
YEEl1ncokKSMSqAUTMFchgnAWh39wyWv0fM46FfUpVUht9F6FJ/KrwRvnFnMxAFcfde5yxxQkeuC
MvK5nSRZLpKmfnnuXapc/Q8R1jX1wLq/71YTksPFSoi5IuJKrV+wfUB+GRh/iiaSoM9/BXcm9pQH
yy7ELiXuzyhI0r+uO7MuOHI3rnI3y943IGSOQ7odVdRSMFBo6ubXqBWJ1F/Halu4WJtIo6jWocWr
iMJ460XSZgJ2j3arvEGtIqJpBsH3J6A3p76WCqbvDJ7KvrYf1pNHw8bAeMDrRjDOw/Vs8X5Buaog
d432wnhKn0GGB4jpnwgpsFxHfSoqVkucUlFP+T4IJAEUgn7Xwu102QA0DeVotp1zFbitDh+skkY8
qTkOqEbxBj50/QymtqZ0104veyNVpGO+7GFI4lxuZe265Kj40UBFAYTcvyLg5s/iolnNLenAGZOm
jIL+LtLWmdvp1h7horcgZMhLdAGDkECVEpbEPquWCiC5gngRkniylKCtCiyz1JLVl1NNtDfgqV17
UFXLGoBXxbrWW6VL5h0gW8oLuUzM1QvlJY+tVBABbitdiUirrNnFSbbjaOioaG2bW2VDb636oy0+
gV/GjdMx1u2MimwXAGndPi004e4qFPX52w15qwZcaeGggHDb9/ei/0Azbudj3viX9L+yS88Omd2Z
Vct+XdGXSZ8DlRQsFk/GXFjA5J4PHvp9N0u19KSpQe9BoRbKVJkMmSn4pq/AdIqyb+RBUrvmly6M
IWoaBtMy5IUFYzbVOmzGrmPjr3iNC4D6QHnRYDeru11O/b79VOa/CYVaqdpYAmqI2A5AEAPookUK
JPWpMSH4ZL6IdtXN9Hyyb3pgQvt/eMW2Zia/gtoAJcAKbpYSzozapocfoe43POYrdJoiFRD19QuM
/+tre7g+UIKbk9qYiwxH6gYk4yyuyTjKIiRqT0UEB2WEH+T27dxkiqdBZ3ceBLbYZ1Gfn54p7d7d
o0mXxcsxIeXeER4p2kIq4EVdrL0966wjByM8xFfswOtgn3gPEkGipdRhG18H4QUkLhAlD7P7hBqc
iqrtUVZLZdOvmfAbJffXneD+Jc+JMdj8qm++DIuonkRGdtdYAOQIr46TkG45TaJdQOHDkuvJx5Ir
vkTzWQwMH/uOogxT7z56T9qMFB1njgkMpKNWL3od4H7Ik90LDqu9tjR+6obhcHTtFf3scEusHlSh
VfRn96fwHZP6LYrBw4Ge68RsVIHh/t399n8Sr8R045J//7dl4aVWoE++QLkrx7384/AEUDjO34jY
vTBueAHX9PU0lYjV2N84F3Z8HTnqnU+Vs9/L3yPgFsiofFHAS+8Ktu7WqRk9GaiwZDdxMJDfaYdY
eK9FsGBPSnlIfKY4qaSDlpdmEqf8TooZISQzyAEM3hB5fCyHJgsT+6rONG5SOBW+IoOm2LMEs7Nt
H5oMAEEM9zzCOc1yKzvtT4roNNzbWoa5QV3IHO9+FPXa6VbzfzywxQ9cTVaml+RpLVDKmpdo4r6V
C3ciPnT36TT3Ehkw4C38pOeWZFQnU4BYCM18HXOWwyJzZoPCy4gkRpcqTRoGcR5B/3t5RWTzO3oP
eVTLsSkpdHetWwks5AlW9M2iNACz5J8dhbgTFQSfUVNmpzp/c0d+4pVeKadh5azHEssPkBjydzph
TIPPq49vC36LuQjNzYM8N9ZBymLSGBytTXCcmD6bn2H/fDaYzk2FYuBb9Y2IiSxBF5saJdDmVVMz
NN3/BA6JAGzG6jDVF4MI98meRH1uacnD0ohelWR4/Cui9f0/BntRm9Zdr8CNmMTwi3mpCv74Sz0B
fUshLCzHvIfnw0VW/GS4ZIvEAEt/WXRxQ7xQ9EwMN9lXzeQabMNICfG7YJKYY3HQsBqsLOZgbzeN
3cAcPelV73UR0DpTlZLODiCEzIaHev5u1gTY4clJJW1+Pw0qwPyO2epX/u3HN8h4eJtIXpkMRpM6
Ipa11Xt0Jqho4JQs1DySN0ev7WFTWYMgjgzXhpli//dmtRkRA2UmmmABPupqN3MNoBX5cPHOAcLF
u2x2GGxqysurVXIL/YNeQU8bBYpkvgB7OYUaJIaWkjf+63fJGwGZ9mBFrBnZleSnmkFD/txFn9Uh
Zk2/I5dTvdgTlqpQ4R74PZgtwl1sPgMMSPNaUL8cEOZNLwul5yZ3UunuG7LcgG0F6KBiuRVkfJA4
BN6HR1TFuXDrsZIYVCo0j8LIGHKiF8fGEb9AakJONHPaAEReEHnA4giEI9SoikebSa3RrQTXgn5n
uOdhGQtCHk7sx2G1vOjnZUQdsAWQwEi497H2k229DlXTnIigu5H2Swjp7Imjoayd/tdBTx7A1Tn7
eu8rg6Asjwor4K8SnPD0wrTRILdYt2T+WE8Fr1IEg7KXyyxTNLfJQDxHCh9CcuRPjBQUnfF6d/Gl
Ln/FkDldQJRVW819l+/H79ZhsHIMnq+wD41uKt9heKvQeu0bmyk8MaRrbateXzbUyLbvVGE9SlEx
3+w3qnBBngqkpmzI27plsuyDLKwJaHAXPSKRXoIyFD5zdC9B4mw6/QU2w/U1EX0NC9XWErAQvb6L
ahOsHfAdruqKlNP1YBPqwDCFI79bmvssLYsYPVaiQV79Q7x0XBFKLW/pj6TOLjyjQY+CA1sTBFCg
hrFbsauRuhNGzUDhVezVi0po1OuijkNIOZ4BzbdCA/qVYsxHSG6QFNv3J1SFEGAFANOejhA786wm
LWcRCMc/+D1H7s7jIF8M43Ch6YMiwuthDqGCL+muMNoYaP8zqf/YIHZ0oeZcvCu+AGiFnlOnr4hk
Zp1r8GzAs5rYsDjaEmNke9mt471Evbd8K+LFFyMSN/9IuuXRzQHplP+irWUDgn4DqTL+A8OSERvZ
vrT96KpKGNqDyF0VjjNO499ySrXnB0arl/5by5pKW+xx00OLeYlNODse9xX9uLG8off/170Fm56F
dcgVtBpWkZHtbIIdDlXjgoBudazXKD0Ilvsgm0thcMiCXVd0/lKqT6WPKyqa1lmOkC2Saj1sg6yw
zYZVFd93L3g8L+LXVIKsufDfyn2HJChKSUW3Vh12mQyHYDSdRw76BGBUY3oAIGNYN+e/NMmyYFfo
VDVyib1YXnTXG3+Ve5JWCFmSwkDa4LhHbHAhKXBGmhxUf9Fca35wolCuVZHe6YF1o2ARbbq1t8mY
69Y53Blm+gN09ItZmUJuR9I/352A4sR2hKpQfLRZF3AH5vunSzdxb0hbrxSB0ngiW5ZWcxh1XqJ9
5o1MVTr9JU9pNmBnEaopReOBO3d6tfDB8xHGtiwoD/0Liyl7uu6uyLCgworabcAX68x4pMC7KovV
4fYGoO3FSF7fVXIF6UKe4EpvXwTRpSfaTK/IpwCkBpmbWIRKpu2R3HEbdG/tNvlwMkl2/e0AuuiA
MtTjZ5S6dPJRKvltMJu3XWnZbwq94XUxMRX5jb7CUzwxl8Kx21+iTD2ENrr2VLc7kTczksaUfARD
5LcfD4j82FEISO9bF2arVjIRwwYaiYIDUuvKD/GzLbTed7m0qEYgpjwTWjGP+M/QRwHT5ibPkDhD
Ms91RiRqsOrmad8ceu8hQr/Xv50WJCHPSWyQBqHTFuLEi4Uo/UuMjIdkWBwNxTHOxXuNGjFDd5k/
iIJ+bWd1R6tUD3p7GCuCg5ew4ljlv0EikQ3vyT5ElqdFVBikspl9ZuRQDj91GBKJj8i4GfNmG/xq
JPPztcDRQkSEAoY6soRbjyBZqHU/tda/HLzjZAtamch4UwG48UFtgAAfUxjByMwRYS1KAUj+coy8
qdL/G6crYAMMnNk295cIvMdjtw50LTMMj7qLBszN9ofCWSMFO6hlpAPym069/ALjCUfL5MKlJCJi
5WynANCLtXty/X6FMMZQfUfwlJz+1HwEx9ciiaYrOdahE6TnzMVCdVvI1SUdkytOsAtoCJaQGU8s
oKFgM6uYCv5mYnyjPZ6BxljwQPQO5AjLxj8UQ7JNtW9CwJdlCNd9Tg3kGuBZMkQisfxUPdotFbWb
bUxJg6d4PH/xdr1pSs+bwXEsDhgKM3IEaX3x/sPBhQtPJwRvB/i2qDUCbL8T0bUEiTjOToua2Jyu
4I0grepBAQ+Pyb276z+4jfIDQhLLKZCnYmOFbIZA6EZxwYU31QKhV0cuXlm13ODuc6QaGaWnpT9s
TnqHwiV0kH1g57/pXTl9H5Ou9xUJZjuxUmNo7ak8TeSwXB7jE6ifh5zjm99LwcoNK15pNTLFH4sO
g4HCeQYJ820ui7vkL/2Og1c0Z2feeaQUDPVy+/Ag1GAV09DBm4p+AKPvdHzRUpVRgFTTaRHxCpNw
0Cn+O2g3ZdNPeQq8sbdzhyIFSFElqIIDUrbKsxNy5XfAAjw+Wsm5T2QiISYCgGzDvaKiBFaLcQkB
NvgEaxDB/Op37IqCTld0FuOO1y9dGhl1SmjQWFDVH+Y+k7EN+iXST9eM3aJmRIC3Szg9w2uiwLAo
8CJv+en13HUetxTryiNsqi6HchOBlgrtfFsyqNFsHn5QTbrZjua/Tp9jmu8dDybH30nseVHYIk3N
gFYBIDRfCfihgWcP7hm8swiwlgjNa/mB39TtsUPa0kahQhYzrq7qdeXdbZYoS5vytgO/OAj6OXOl
8YfOlZDKIe8puPEhHAKz75R9mLuu10uFfyJWDYh/f0xq3+n5qWbbGihswgx1zzntrW9XUGXKfM73
H8uH6++Hoq7Pi03d9i2S99U0XzgKjvAg3DGrBRgAjfd/HVgsNnTAGSapszquhZhze1YmkEi9efUy
01l5g0U/oK7r9pLqHnAxp8jO8xNChCp4U0/J5rSn9/hz1766PrTTUCzm5ARAXGPCDCR5ZCsaYnGl
U3w0T9o8hDb2MhAmkwBg+g/HNNb56lADxkhHJX5EmhaZ3sMXucTHOpQfYy5QojaqfJ+FkDJjsfOf
AYhzgiB2eOCbXXvrvEqGohTIseQ65EocOE8wojW3lA3cpEJEEW1Nqz6iNyBvVHVeZBRhTK0uyyoI
kLZukXoTZYNhpjEw8Fkwm0UT+gNhxlXwSJU3JjNCUGVms50ZKDbUvr2GOdmCRRW02+H8ZzCDyBOF
djQ9nQQSvfJjwGwbJFwIJtFOCXfEPLgsxIcwjDllk2wXnH+MIabqsod+r+W2GwybekHhcLNut+6g
c94Rg2Wdv/4/3LJw1y+YSRPbO1ITNscoYuYO+p6LEagXpVdkU20D1O7hB2nP5e4mkHQsoALxhkp5
PD3oHGbx6UPK/xmOEn79ZBPlS86z7j1NLT5Cq2kxsqhH7tBmdkFW/0NVQXv9BURL4hpkaEYczUu/
Cn0v4V2y4pcav/168WSQhFT5h6PtU6oGIgBICRDQk9D4LxeDoVR0K/YQCRxQ43O55jU7IJKhPw5s
74qDqtdc9BxWuPu5hdUcAeUsgCat9+ZsdYgNWlePWJq7l0+Ikkf6NQ9UEFyiodzAHS/t1eIJGlo4
43o7yCi2b5GFxrtlmdJNvpqVVSeQytiTnld5D4suCPOTPvm1ylaQtpwzTtDao9ImBLqs1NhZWsUM
twTwHz+6pUvdzLdyx1swZBBx3Ihvq2KyRfNer4zxAlb3DzZYuqDMYjYTBFy26n9neV73igLDtWsy
Ylok9gW3QJXdnfkPOAHWP8fZ6bwzx0nUFWjUV+sjK5XldtLhr0VlChmJbKb+yoZXYWepH4fHVcqC
NrNAmBJU4GUKPpKvQXPKy1nVfE6I1sk4iV591VoS9GXFBPxL/h6g/tMXLj+a7C5MWKyoR0IrM9By
+SgdUSjK6IEVHV28N3bT/2N0KOAzp/bj7bCUSvMBBmdhLBqekCqWQjh0I+WJzyM0aVAyKm3dw3Nf
SKxmHYn9CgSwXPX/sJWMo2IQUAbI1mWfirSkm6Y3GeTOL3OtmmkgBakL9HONt8LXeQe3p3HUrrxO
ADR07zQEnGX66GlHl+hbsGQqm1mBOmo8pAZm5TbmYJ3NlTR10Bhr1qQlX2yf4LpRegOjukp4uBQa
JYKgjFdzkQtM/yMGo6OkdXx5b4HPY734BNhq7pzAF+4yDs3WFNLRoDdvYZWfWV97PX6kf6VpeU9S
iSx8PLSaVcBfpiOAlwqVKyaMw6EWe4SlP8a+p5+Co0/kGuHM1cwe9sx4XlSjtQmuv+HYpjURayB0
mWhCNhbuSACCg2nP53o4dEOIAaYqjLbu4DBBmpUW5C0MoCQz1cz0Olz+/81AuwBSFGli9DXOs912
AeqSYtZM4RYSOKOoQddLlRwooE9osCM3bJ5TMf/zW66ajMg7ny7vjcteGyv+0tT/p/dMtjNhXtEk
nXMkIfVivxXj892mngmSHvgJ+gigwhP+O6D58zrv8Oa/GyOqrGxTKK/cKDOkpIsUyifY8R6ikF/L
GjN1TqwTbJTreF+HUmZmCUdFv8aJOP1JVzg4aRauxkCZ3xMZcD5O/bxRaYPyujgOkRITSoqoTbiR
8rgA/ihIaxg1rk23HbvwmmeZeqDVyu2vLHbKMqS8GhjOtYNb+CpCb+RHrAmaGEAXqt1xAWxKZrLj
vlgRlnV5jSJ2bXsuth5rmVNOwieYEwN0bwYlZATHikh1Ys3t5ZCjPDvPNai3Ol/moKTOUuKmYe/s
2IFbX3m5ZDrWcG/qSl6VqIcMaoFM/OYyCGtePT2updL4iX1MRbn84iaEyfgP8HiuNoJSTOSycApF
/zipLEDI4GVNyVDUv+6uz/RbBuRWzUlOYCq9LajlC+e3/iwuvXHJkBsPwRl+30z2EIYV32XHOsVx
/zBW5idYrJrgt3MQrVlIRrNZHFwN3rHBcjIgGi7KQxbinNLyHCPaUoRbIWqnVH+oRLqKzRl5edQM
ZgUahAoOQTb6ARHm26wYeHh+02TdhRxKjPIWS4Kjdyspi0XMzzmzXAnCYWcAcWxfQCtUypZTKDb9
jS3uTuGzKK+ricKUvReaiywqNFy/oKSpDTDutM/KNor9W2WMhnBDdu3NWL/GklYrSlKjyzewSM0u
s7CJ78rF58s850VomYj6rsfeWtdXPxaTQwZruBvUUwXLA9SGl+5BR+Z493NXY/U99cP3Rskykz4v
57frM/FnbrV2WTIshPuHV+fa8yxDFqsLWhzu6BPuyBNlWzyX1QW3V439S2DwFb/EQqN6HO3VkOZE
cxRpbK60m3ilehD0HDxqDWm8nYDL5CBcNNvJbF3RO5fNKOZ+ADHp0fLDErr2GSiEFSzl6GWVNjc1
wptsd9jPAjemXFdmRWyEPQg6VxgmEbmt310JWMv2K/JGn2yEj49CZ60puTxVUS836Uq2Djcpj9NY
cZjzdDGFO2/dX48oyo6UftZung6X6vTm51T6uttDbaRARIj5PFE2k3NHdzM8DYWXMp6wHU1Rykd6
LueEUcNrxcd3gke/7gmU8qSaaQcvz/iYEnwnG3txeiR5og42lz30EsmuOv8IeZ3sMlxOXaOyIqC4
9KQrZsR7kLJTMG2Escb0Ed8L9x0imLt08jQ6guS8+M9y4VlEcyUX9fZBj8WJ8yNkMe53KtnmOGSj
RdRziMpXMrysfEjzDfOn6NWTS+bnr4gXCMzOmWteH9IbyhGgPXwEAkAFDIxhDw6aNOJpDf+OnYHc
l1bR3l8mRnHEYOfKrerzWrj3H1ldelNydqjLRg1CSttIvNTpcZ63A8SayIgkZrRW/TmUjx5MCX2i
Dss1V/W4rfkl2TLBzif0yxSno/2GRpzT8EdcAyhOMm/M3GwPmt4XK7l3sTQ9qqyjk3QFrAxz+bNe
Wfv2cFuMF+w1+LL3rJ2KXnmLGaLWdJ0q6Vh+kaoAvEBvRnWcjUGHgN2/2Z5RTh2kkBA9Ps0cwPIR
jRGnhGneccog34tgm2rmEeoJ+Caa2lFTColykkRPfdjU40w6rNtRIGScz2cHxLIPMyfbPSudU4Eq
6+JPX/j0lf5ewxxRJn+QAVlPA2wJr5QaSAH2GTRbOEPDusio49oOcoh1Zp4fgz44RuCwZMAOaPwy
kicdoll/zrtBHHtTejQFPJmkXh3m5rtG6SC4KjJ7ankjb0EJDDjW8C1Ji8sbIG0EHA9WQQiRu7xZ
l1xE/cC4uwn+G2H7p0LGb+iCiehcDWuehRIXSKRsVncl4hEKxlNV1C/6fVyqRRNaaLHOaE+Ya/Cr
KrorLqcjFNkM0EIPSozXh4C1RAHhj3wfBNWYQsM3wppTtdkVXQAhrdohMUMYKpr5tBAqLxxjaVDM
cIXaAhPQdGMwGVDnCPi82rXIV1SOztU2gPTCDAF8AZxx9npt3Z4KO4i06Z8r0NMoi6GjUSSBAgIG
3dlPXXMOTuzdNU6X216f1pvOdY1h7WWrOF2g9JQ2D9p77q7mtDSZ8TYLoTu1ug9T7W6wgqAM19gz
qKgLDBY4q+HQgQ6XiburbdSB771ujlHpBtOKXLwXGjtc+Wjh5nnGrOO+5ZzRwpQZKZzATHhySRR2
+oyzJtt80+ahijzQtYshLJoHFNixOXqXfzAJxTSEE4BgDpU3AqvpF0SOZ9LVBZCjiCvFUGnzF6Pc
Z2n6vEoOh/guxvnoX5pAHp9IeCBOOtbgKc0gvMHuvefGxT8cNCqoTiaSQz59RFIKVFaLYm/7CtP0
Ofrk3KC2ZTmFYOxD5hk8c2iIqrofPqfxPpKc/YB156gEU7PKqJrDqnnsx4FasdjzJA5xYVJ1eFRR
I9DH73U+dDOb/WnhOXmHHkXYuZZD2RKP1NkS78U1W1aYFitqO64ziVGLRjCjv0cd9bqquET+10sI
mbLJIkrbDqiiEfUpIK7lp1ZVrNn7clmBbZQHBBEyYLQlS6aPY9cZ2PeHWykry9VWgMiWh03VenoV
IMN0/U2ED2aAaWzv1PZnLoJsaMOdBdjx7qvTT9nUbfJIqz5XPC8J//RXgvwtdlGyc+8GQOViLx5b
FbYA3YefDzLab0OT6AODgKOEjIFSIHRy8geo92rQvKbmxP9ynadbxYS8F6JPyY5k91gocgrw6MLC
+mpMk7prqu5DLlDh9KP749Cu9vvq+1m/la7CzGFUi37FyjlFZfEmusu46g7Wc/gB2qnsHZWiuf/a
oMxDk055yhJf4CA0g+qGGpOeBoEnEU1cpanwu4a/XS7JZ8vAj5ErqzCjEGGPPvh0KtIkWziKdUzT
t5PCWxj7/P3cOeRGrfp9YbCwh5rSIWTDqNZriX5EZhwo1oymTovr3mZ+F3WTLft5JgHJ7e1Lxac4
8rcv/VXSOMJRc38fc8RXzTrBR1MoWfS8ZvB9yZIKjXXww82dWmGT5UjFxMtTG46YjGoKwIi1tijT
ETYMoLZ2sNBDjN1KZfKTNmbWgtI8fTqjVQBAuoMGS1MgscBZUPNhpYiCOwK788oruv1nQ2BR1rrt
3ayZWfhzyGRNSwP+Ggq/GJGEwbn6duAw62Sc42EGcfhGhMGZ6b5BXSwIPBAeh2+xDjC4A+lOq2oP
sQ5WMKmXV+xx8khda+iZFlke0M3mApBXo/pL+Y2EfY5M2DGQldriFUFDrScVB0ch4i4SaBy9dBms
7al7UmA3Htw6HWf7RjBSZ8WcdRfNvz7beikxeqpCh3uK0CWIM3jtjKvhLlrtzRQve8OtAxJajwT2
jcwjq3xmzDSjtSbL5Ry7Kbg424aCExsDLudwKW54n3lylsXmJQ0aZ0/ped9BCAtuJzVTU0sEIcj9
dqNn0ARKqzMmdYQ30erAv+vO6TMlzgGl0zyv5AzrJ6GjJUhw9H3B8Z8QLi6fTNl6PpwpyXe96T8H
HaBWgJuvP1MMChbPrJxzO/cPwcL6lQQfbkmNQPFtRXA5WnIJp9nb9txP6hGdO5fCylYyFRT3aPmi
RQtD1SZC1opYrL/Tx8m8l6+6hqUxe/Q7A5unxkY/dzTCgUZghexl6cE6WmGKULK9DWlYeHtuhXhw
fdU1XRIcSk8dK2t4qTmIA/fyn9UVjQLZcGLKmo59eACxLQS0QfQD9c5hnnnARHR5Y1v+XBZ6pRg7
KeC7+QWwxi5xsaqJ2WPvV34H3LJ8px0dw5CRVdDpuJNeTMZsqKdcbvsvXJuVmpd+7vNvJu/E7zVL
LzDKl1lNdI0Jq9uzU96Dxfm0x/gSt09TFhLeMvOS9SzwRHyd5ujtS5wKvcYWB0bckKroY2ZSjOvF
fgcF9mJ2LtFtTNSMjIS6ELJwwPfCJpW+sOaah3YDgrZCY3uBm9DSxflJVFLv9ANw74kLWoKLlMKk
4vkLLxoqyppsI9/PLcJtPWclQoUvxzCQMj6iPby9PAIKju3MD4adsDbKDBH5gT394y80p0cTDgnZ
W9ewu+XaLZkFb+2j/B/sH/WmVSi0WyNG7HQVHKRq/J0R9jORgb0eKMvcUEFwnvuoOXMNvcAYzweA
9AKnx3vMcuZH3vkYcwVXA/K0ToGeFXE/9uM7xGeay5sld68SEKU1a4CLDQyNpatWyvMDrZQJTGLw
o3F2DGz4HRvA1SpQs7zVIf20xwGGK6fTBC56xxHF6+nyLidwDiMqQ898J0mYVIHxFjDDojxj8XbF
e/skLmADK+wKhjvHCEyzTO4/opfnxVrszKfVbtglvHe05M1gvr3ZnTQ+mTdgOMToxNQaZ36Tegl1
u13bCPZpFL5aJB8IxTLY1w5SenSW/5FKRjxdlLrV/effZaj/Fzf++Dm2qw12b+eq1VkP2z/mUoqA
mP/b7p4GbZbcjhQ3uItiaYYCDUKIpMbWsbYH6lhUGVjhGMDwGxQ+nsLpnTMvMcA7azdykkPmeBP2
skSvgqeOK90jkCB6tdov8H5PLoAROtkEe5Wg107w3/Zo+vdsSL1MeSLNjQLVhSzF8LJ4ypD2lzuH
+si6ZlSLAOTAFioD2gp5XwdXgjA34x3l16pKGPIfMTzigm4sB3wkOKp9eggW59uTpvfScs50Mu/n
iR6Z8mroTejpndYMVl1h9DNDUS9sV+LsBBaE1C5WZYNFbdta4Kb/HSOFADpa/6TgK58VqW3WtZp7
M1eh1ljzvcYZBdF4cKsNhEfI8w6VjBZLxSzNZXMh4qW7fW48UFp0/swYtOc32pNpUXd3BO9I7SW2
E/6mSx0s3upGh2A3ZXJDzldne9cbT1J2Ncys4eWMpp7Zz5ReEC6k2izmGuoejQHM9A7YoY+ROm4w
Bu+MuE9YmpTzGE9TNQcDGMoZ8uX5i9KT+0ym9MNjOLjEjFJXyS5IyGSMRUtbRoNieQ6Odww+GFAJ
sUdr2K8RIuEbLlKn5qQ7bO3VW1Kq5koFf9RefK1nJKNmjIKAPZzD/GP7JS8Kwqg/IN/tv76gfQr7
3ah3EWi9bxOwKOTk97OzEaxqT/JqeBQdaWA6op07LcchFjN3hsPNPQ6kynhgoBKjluSOH+nAEwyk
EMEoxg9H9KUw35rSbBLMjLfpnjaEUXJqg0NVH5Sn7ZNv8hlzwi7KwMSDdctNI5liV+Ds9ZO/xORZ
GnUWJD+ooGnAzPd0WmPlyx9+ehn0mnFQsOeJ7ezkifHJWVAlfyLpFe+LHMXjonpHjrOTU0Qdg8Np
NkUcv2OtQk0+dbxY1eDWB6dneb09WZ9M7qfz3Wf4vmDxR/iYaOWO1Z2a5HTFEOFgh3Oyh+IKiYBG
c+vReK2N435rd7NzCeredMAEEgVJsmMzu8QUCmJDV/HKrOhhV4ncLFkKhq/VCXdUiuGAbFcMdY/z
MSy0mMa/Kk+yMGASXjnILM2HO1SL9dA/isqreMalVjmdWxwVBQAt+sYPi3EJ6LLR61rvPiE+Rygp
iAkF4hktgc4sMFR7RnX1SBg3sy2wWsIcM5u+/5xjYkKih7CKByW0oOcpxFVslEAAGt+sKgwAecGn
CJZkz58yChR0/Go1w4ATzyDop+trIHvZIU7vMyZAfDq17q4yGLAnEhDS1AWywfaTpuly8iOuC6ut
33/hL144RU5bEhN8J8351jIyN7Nq5qU77Jo4IeXxakvkQRQZQkZNV0CrJyc7mzdADijh2H7gcMEd
zyjZNxyoRTwrHVKt1PItwBTmioVSoUmc4k+26M3VRR76ztzyoAw+MEK9BG+BJYK/cpC8CPCetSKG
C3S5resemuLFnsRpNPIv2ouydRaLAKG1ZDfbY9qtY0FmqTvQJDH4taWA7g5yelkXZQvzy6pQCWcX
ZqmB5gB/eYvUplEdcU+sfhqzNf2KS4Taf4jcqK4CDabNTqllr03uuHwj/OEJ2fi6cId/LFApvSxT
d4kzOreL+IHDNgXLWhCM++7DVD8aZ+Ft/JY7elcW0LoaNbkdgokZe8a2p7Mnx4Nqi5dxAaMqMngv
H2tm/teu4tPuCyPpGAMw+dFzTkzAS4hZo+KEVxl5VDRmqecC8dKHRFuSyMxJy9hDDkiglneMde7S
m8eSUAZJy28L/x5R/R5x7S9Q+bqFdOmpnyLJUK9wJxzEDu9MWO+cNUXjw9yRM4fn/ddcSo6GELP/
5+CS7Jje6vw8bWt+0UA7CTcReLEPJfCvVKOt8UABqTVtGXUxvfBt0mW2yu8FKOs1z+BdTcKLx2x9
e+gU23BTvOyCQNzsw4zBZpuJVTRHtTjvgWCS6ZDv3h3ZtchixAP4aWHgMNRwyuWHugz/VZgWiGAW
36zBNrCrjor4slu5O0X5NUBG57wuujr6lXK/8Y1GsD7YKkTWyYn4CJ8xkTA5hVu2O5v269201dor
dJaIi4V6ANcYHF1GzTWzLEmY7w6D0qUhm2t0weh+lliWMGJL0JeuLJj/TdEmNqA4gv8V05Oi3CXG
VuaJNpvsAh4k5Hf85chUsXRpzbpI2GYD9VCei6jbMhGDUENZQ1Q7QQWcp9aNjMMAuaRC/1fgGoHm
Z4NFMW3l5YuRZa9VuKoosrfe9WdZUEYmAWx6pd+ff7067XKzKnvSo2hFh443RsyLBf7AexFvgwov
Z47lwV+Nu8fu89rw3p4HwbupW/h/hbjwqlo/jKcBQ8esGDRC3KKUTwGJdSOFPFS3y5mQ9FdhgaYr
Xcg/75LPUhygodE6ed1u+PeNSo7HZ4W+Lxgema4IL6Fqs77LvpxgCHd2fhw4bw9u0ja5YfFb1WA7
dg0GfQQCX3HgYjnwARVRBC8vLcrFgBQ6t/t186Ux9HxSBtGkOzm9PsooG8g68WwbOQbE/Ig3tJZk
bXT11Sz5dV6VMzfj8XMy0vNilWfbYVBfzX6ni11b1tn5C3UqDks6UjtLUCC+t8RFj9wPsVg3CDU1
bP9Sjp1O88b5HeOY98hcY31LqELqZ8dHE/Kc7JX6hxkobUuQde9/rgNUrrPqudDwImAR7yopT82t
q0fZrP7LB969Mfh5tedO7OlP9WJIXK6/UVuEQ/RL0u+zXeb+xQSF7rJ8liSrWxVotuisrtA7IKRj
aiF87SUQGtigllt+G+MxIrZw0DXsIZIrCKSZQtRNju8yupsv9KRRM1O2yn0vQadN8Lin2yAycqgU
/sKA01kR2xkOdJonv63QhTM5+EHV6byFgaefhOIGt7M7e1CBjLmiOBtGX5Q1juKB5/LndxqC+Y7M
sSnNsAFt8/WvIRWp5lsPz6+t96sbyxS8shaod775Xb1MhApKH+/RqfVwYmon/smqn6Gyc7l/KJRV
UqkK7fmnUciMGunhHAZjic25YL3GssvjqfdAHE0U5MEqT2/D7wyF84Cxr8V/uOYc9fPbZYoErcT8
9VtvNzq+toJrHcSikY632wIjbezZ/D27hlwu5pyLFgCsPD2sIECWQGPl2urrg23aR2b+6I3s6I1C
3u5Ze2p9PCqkXLk8N1LSTJ8C9xf2LfCxYyQicDVR/EMsuUDz1fJrO3YW1RdEepSPFd0wA/qqZ1C9
oh43s8p6RTnqmsPDZAT8fjeJaDvpIeJBmOiRrZeEY+WXlC9rO6llrH9MPG7l/cs6PyJ4EexPYwGj
CIKdbzBTkjrcDiIWyHU5iZyjBNVbxkbia0lSnhphqFNHoK/qxDF3rMhgTlN7l0jzDAsomXE36ysb
wsnBcEcnYYlkXaG3+V2Nwo2HbRktXiZ3Joq8RXp45RLfdHvigd4qqTCV4pN0wg4BIvsn9CTcTbSU
EknbXLufaodaThu+rJmJr2nD8AU9LEYmmYLGCJd6g2ifXD4o+q+zimw+tOdVmkODT81e2mI9ZR19
WqyGCEagQauO+e/LpBC8Xs24sBNysOeYvj5Jum9X2KbTwZcgGihofAGXIslcjOnilYF8zN3YkIOh
t8EkUsSrNngS8S4x1pnuLFhyAgUXlj+Gnb/kxGE3GytiR3nkPe0OWp9PiaiJXf3B8lGv1jr+EQny
baNVvHlSQSUcj//Xq1VyVerNOkTXyQ4qTkNImopXfAj9Fp40LzZER/enQB4b7b9bPM5zoxmy/Rrc
TATGDiBvwyvkOlGV66JzD9uHmEnUtDq+OpqsKnTF/2++tqlBkw81lFR2Cg6LCL6bsrEpO6ce+g8a
04bacg0uY5rrmYiVYJJzQoaP11qZbCsqtHYVsEXqcyg9gLMWr+to8PnrZAgwMVLANjjbJ0UMtYwX
KHSKTlP9Njk1BGwZ9cFbtB6mgyCbswsN9ekBM/vKO6GUosQOQcELhOz2QkeNRnQoD5cXP5hJtsgi
JSbIHgAFocmw0wNFsayz4vq8Wg4Ga/hjmuAgn64Bmg1cUd+bhLkw94XM4YlLGR2btSJkQ9ctMito
gBO3sdssHEVzkRjDDOV6R8L2C1srg7lVb9fNibXoZPa/3Z2JQbMYYtpz/glz+mt78x84s4HZJ8+g
Prx5QgLjLBKA8OEObos2FL4HA5CtO2kDKp3gAywXr0mq3Wq3jBenFdhdhhS0bZemmBm7HwUnMXD/
gAQtGstCF7Uf1h0Ts3JgZIrpFC2iOXFuI0dK633zSYH2IK6uIBVjKn0VfHudOtXF7gVREvZrcWr6
FG1yX0F/WNathS9qs2DuzR2PL4cTu/2zxfs+Vhfz8R9F0xhoo34Ma8kLQm0jy3MpOq0V2RQ5tnJH
kDkT+uHS6aNkdFgnMYfZmIZvSqC/q6MBdTOtSJ4oAMRhR0YQmMb8TgKkNAAoUMZaUUU/jEwVnvyi
iOqfvz0E/IQZt1plyjTiqHa5vho8UwcunnRXbt51xQMxjKpj/sr5Bt1SLE4DWF808zpWPJFAJ0e3
zz1Zr7qqSqBUgnCw+SIRwB0mgyMs1BP8Le5JSGwlP/U+h9AYsFXDDFltzK4s4gy4ELrruvniTJ4p
pku3YD7FQ6oZk2xVwrnhPVBbq5UKgqXE3mOUumsaOKpQ5hq8x0ZzM+GgqxB/t6l/ZrxeTDiKt98e
nfvqs8BwBnwM2xmDYkg5O8Xn5IQscZqiiJAlxjHO/lG5qbiAvFllpBw7SmSwM4kyseNbJFCSJOTP
HlrXUnRnOFxlJ+3IYZj+28s4qXbA2/UbUC9QfYu6tXGCOvVP+GdQNZ3TaiLNWEvVAVdqBH0v/Nse
h4DYxyOd1Xr69lszp48Aff7MrYPPKf/eD6zFojmCIysD+4b0IX0tls2XtYTRecQiREfpMsCKbz68
FH8eQt8kx+P55UHWfMdt+zokw6aOencEgIeMZPs+atJ7Wq7BmCewDp7c7dqDwOhH9IJfsiI8IBq2
9KN8brStKSsx1TOF5qAHcDJXmUa4X5TMuQUD5SaYs/wiy+uXg2Gth0zTfMZOYqHDSo70iKZxQbTz
DwBF5l9u8ljOIqKIR7NlzidhJi5nkEzky3pv6Y5inACUuSQAbTBsvGEZ4d/KiKMcpOZBiouhiJFk
oYYaF8WJqCaV+wqjZMIpzRsJreW5WT17i1NdhGXMDaQnUw2VimP1sLhvAjtSODVcRtxUs2GEO5VI
P8dvfJoi1qaPoyElslUTNvwDasOgTVW62mr9bZCjqEbgK5K6VWXNJLBctZlA0JsVvdWyKrKY2dq5
7MMNbqHPZpaCLd795aSVXhJC3ioqE28QFODIUsAzs2z+umw1qQcSQntbSgli9UqWvc6wW2B4Onyg
QKWk4sSEaTb/lUV0sDTzo5Ev6ttiIHk8kVEE2LFLVK6+avGKM+l7s5FzuLh/CJ98Zi6dBP+k5hgE
8BEg9ts9NcpnbC1oHrbs8qUahOJuYTWLpOGXKUwPy5RUrG9Cbi63lAPnalqzSdiwuaJN37sYKRmS
B++I5KxghZY4TkjO0zSyU4rcPyK5Lv51kwi9YU++YnZ6rZyCdXipO7D6r80fhHtVBbO0TfrV6y9N
DBLPtdvJuo4ESBSF+PNRdMyouj4PDUZr61NBDYOm8FgxLoUdt2w+rSV59CMwr7VmWFEYuTdIx/qb
nFLHiSxHEFFakr9zxNBeB6bGtBMSUlC4dbLSmLCtzxVzGAN3sX6t2mRgQMJRCoqvKwrToAhs1RbA
7FQzYCIxt4+JCs65RX6w6hOb4MpBAAK18okzfy1mYXbuw4PPXlYiy5rq1voy5ZRWjH3hzWbf+Rjk
BTgQ0KL6IyZamdRIjCCKKTgUcA3g7+nKzBhHZIODdIAwN8ZMKKC2BxX/r5CUix1jPuzJ8KkyHnYh
wUVY2jiyE3SVNXhM10Bu8wqsih0EMot/+FO9SWc//XEFfjwRSlAbqGyoWhmyGYKiplHlR2ZftmNs
ZfxW20P6yd/ChcOBfVC4iC+Dqo0UbMXbQArumQhBuhmggwIlazMTGzSvUp39B+97k9cna02QA2Mc
dcn9++7eflt/zYDj1/AFrTMTkrcFFK8P/wimO+IWNgHqcrrw4c2hU5tRb5M6fCSBBhPUWHNidzVb
t8qlDQ1t79YNEn5yeTrt3+LlQ/ARLDWjILfe/aQe5enNh0ISzshatfByO1/MmQBNLAQjGdACJtR1
RuTMiG7/MQm6xMRxAqERmVdYwkCAG3TRU+QsAjDuZbpXRU0xw83fFRs+X9GmtG7bC9ZG4hYCQg3X
pFNoqaYELByD0evXv0HGGM78VgVEMnu4XBhH3RKRIjk0XuaRxPcyTczw74up1KL9C+lKnnV0QUin
FnqnO8ZSAoAwHj/SoxmLjA5zfjoNWSNliI1rjFe9Jl519qgEep0m/2qMMjIM8xspW4RWCZ5ZE5I3
eMHbEe7NpWjoRsbB/TuC7V7Zf8343LCmjbLbKrZ59cf7B1vomrYED1m7jmAjeOAGs92HP6/cMi7T
BclAJEO2U5XAs1gUomEUNKC6GiH9nXWTPiWJOfy9kxxPYC6SyQtyKGmlxHRxFSnGBs1+BXr/upAl
62Rhd+ZFctnUS2IS8HI3flQhAxNcfqPsEf32YQT1vcilbEpgwyn+iL2ETM9RuaYOOX8xp+nEjZXp
TOeOqBDiq46CGht9ufT5FejDYqHiZsN5j0zWiwW2AucZ5sI7gkaghsZ6L4CXFYmFYuqU4/JoTrRq
3qg6EHI8XNO3dOUH+z9hIdwLivT+psBmaw/n/3UNuGEoeFsV+VmJvsNdyWo3FdgPtkomUFxP/iAq
foo6OsPRqeIS4MTCgYKLPHv4WHfZxm3zvgNZMvyDpAyiZRmHiarLMtkfYV7Zn0GvxantwBsmpFIc
2KNfHxW9wabA2C3SPn2TfuwPw/uzONUm9yaJGMV/ZpCziQKjXCyTyvYDsQLpjkvBhkMhQhophHYl
1GDi2GpIrJVpq7mFqFdHcDyGkHx6N+em51p6rBDzkmqeHeXKqySgi81Zglph4K1pSIiwcPiWtQtM
MfihdfBBrXxA+lzlIdfgF4DOHpF2ajds9mPnUsMvs/TUuH7RRu27totGJsXD6uhCqHvHblDGw2sV
NC0mm/ZuHBencCrdcEapjQPFvm0fw0Fp7DMkPSzfmaqEQa1/MaES5ylsDzoxx4LieuI7C66vhMsa
81T2Mlt9B0yxnJSVDjlfi2942ytZseaFak7DxIQpNpXmfYT1Q6QqJod1EURuj0PVp49l9nLDZxXd
6np7e6pEKEMRTHwdxZkV7Wnfe/YD1VxHjS+uOx+tIukTIvHrfKS6cf4KMcAM5Z58S4wsHzrpb1zy
B9JxZxwGOUdIGxkU1BecoeZC3jSNtKYvFBF88DvTbSy82cVM8a2vtdSV1nGHE97CZPtLPMQpQ4BX
BI9ZDcrErS1HFEp+lTxKGgjUgNPWXM4p+Zj02CqpN5tq8k6NeGNR3GFgIM+FJ6f/UCL0yHqU4D3y
Gl5o7+cvfVmeahXGn5ZBCIf0/0JwWGY2mUTcN6PoRo0tJG/HwMD0d5BM3MQMfP01/EAX8L8hKMp5
7kEGOX82XEjLy4aA1lOUwGJW8p9V1GAG3ezGTqgXS4B4+/nxB/Q6iXN9m8nj2G8y6xdr383jM+dP
hHIc41x9InVzm3azdnk5vH8FgX8zEJUus72SDWXbhgN8ku8IhtTuvQY23fE2BMf6FNuThVajitXK
MSgmf5b3/nbWCH2681DQyeUtFLfZpM5cSd6WAP6CuyEzeUdGGt0bwv4aK043x/tnrjhaeOxNMcpK
dgfv4XFjRZ7yxTiRNbjDn11ac/LI86aBILyGjedgtAW5pt9/gChiomR3mJW5oV3F65gkzAqHTjMW
qAUJgBLV2+w7MdnVqGEyORLMXo/NtNhZBB7o0aO080JjM9/0RvxDZXr9ySo/hlsvhSnFfoP/PO0j
yHHa44+anXkQDuXtrM9goizIG9mIVng6MURgZQkbcfJWUfntjHaoNABwn6kv1qng7sQYx39a43a0
vSaJU6iywc252kxZrPFTKB/FruYvtk+k/p5LtQJhzzVpamrG4UIHhbhxnGHAQGlqTkg8VOgqtbFR
yeV7AQ4QXJKxR2QB5BGeS1wfHiZj3+vTLHG78oXO+MG7dB1VlHQ++ko1Jddw+ELSGhC53ql+2Ncc
lQamgIRGu0+KXpJxY4rbf6pSSoKAK1WngEsYBY+enSfMv9NamFhWb9+5zHIqbpiuHx8HM6Aa0DIW
os0bEUkPXGrxLUui0/oskVxa0rDElIyXdirlqxgBzXf+RwpA9VYHHBZsLy05qDHrrGfaJuZEwiVH
+tcpYoq2tP9JMCeNW2BBsWMrpinPutwM+AXnXOaync642+uauXvmhGxtc5aU+sSkmpmEVsclQj7F
Vcjs48QHQQS1QfyqL25gnDDALF3htpoBgdvVWyoQv1QzOipIFFQ/FpFziWKJUD679BUaO9ACZikz
j4fgpmcN0yl8BC8UrsZybNsG+zmVM+a6k/yRaT6AZIejC3rw00iVI1nMKBi6cIUiVdqy/roOfTvB
C0io7y5ENYbOh32TzikblZMGt0GpyAit2yjCBe6wagVVFRFUFjk3Av2rXYZgOM7IRRtFY94Y55fL
L4VwuokPVAKbHSfwjUt10M8wt33FIXQJdHGCX9r379ud9RVLJy9w1Z++i3utObRMLdVh9UVaKjjT
TsKVUNDu3WuMUuyb4cV7lgx1LtAYu7kOTiWm8JCFv4ZrYbgbLDUWg48vGeDYIIrkW5bQRK2/kaIh
jVQfUzAcSSIwhvDTZMV8OLc93VCN62nx1Upopk2dkLLYlyK3x8rXNkUpvfH914KAewCM+bSZKJNB
4gv7FYWIEFIBRrrZon88bI5nfGuyJjqWhr1G4mNO943CwT/pKAbj9pv9RHQLjHtZhhTXRPdDMQTR
tS8PE/86E7Og9dbAcc1EY8yzv2ifznUfhmG7dTkjG8edBS5w9Oo2kBllDdtA8pC61YjF1BUC6jbJ
7e3gVNT73b0bJllp/1WN7+OZiKM9VjM6rSAqSUA/Ybonh/dBl63o7+Z1hb7OjX9LS8iiX6v+Jy9e
o0KvfCTH/0IrGrO+SpMn2kxXjVCIeRJetxDIUTZW6zI8Zt8b/ci+255v0oXKdH2U7yKNqGRUlfME
VOT83Tjj548mHFIqY7sEYcxFYC0gAKQ0PTwi500NNsP7L/DZgLdSyzUu6FtXjkWZslfAjRdDa33+
mFrI2V4al3WI9Egq3JnYHu652WPO75ksT8SctS6zhZIQZCx4fw7kZHFEl57Hnx8+i5Af1OjnuCHz
dHldMO8MUcVRWx9AQlQUkfVjDbX/0k0YNstdRI18ZnOfN6quBZH1CVaqDPPx1HD5VgqUDZ3bqnYB
EbyqshUTJK84VlQ41/957Padv95ipdo+Nf88CULm2LonclpsTd/KTbSrMI9S1ROT5xGxtAMUibRn
bDqh/eb/ScYDfVTlkxbtUxK9FRf9mHdrtSVxJxO/xSPcw7XN2uzPIFUw75iVHtVdrYUjYHsRlahm
SUsnwYVrJq63CPOnqan1ixlGH4DtYmTF6aD+ac0jnM80txthCHNUk2DBZ3461q2bhKfbYdoPKyXJ
+S8nnl0dLEI2DYOQXbJ8r4voUZEt4jpB2SQPRkIi2KzOtO4p/7YI1Ogcg9TMFycMXP5+uiCrHddL
b6rXQvzw+vMAAzlCFr5cn31YY9Rcu49Gankt8HzDGfE9DZLWE9BrtTnP4BEnfdj63Eks25gJKlA6
ySzlCYUVmpefJWBBQyKXzfRqA7bnXi+Xs3nLeMI+IYN2MIYEHbxAEFf4PU6Do45zJ/icmMJm8mn1
iTz/u5WOCTzYw1yEFe/VClLox3c9mNeju4/HiyjNzHjEKEJQijHfPANS+AL6Ec42R18VwwTAW8HU
Oar7O2iNceP1a7xJ4zqmHKv6Sk6vcKnwAVCa9+x8kbD/utP9tbMjB6G5thRjBVi31bhLRTM+Vl82
QaIcDDefxQNvAZV6L7PyfjTl2/ylsbf4zewhTXlajxmv/BimCXyai44m/bbYDYoM/wdN216S7S3D
F1pgyA8YJ/+nzKT4tOrxv23J5alvN8AGNL87YbO8/PxY7c055PqsJ21c37Ff7lIfC0nbVZsm0Bq9
6y7WQPfo9qt92f8UCmCHui1H3clT5JSnroX77qq+5eIzUlfv2o+SiJrrysdS/Zx3hQcrgmYhGatA
Fdr+8fqth2CAaP41rPDwN6skIHLQF9/XalegwnanwFzVilo+qZGCONXIKKLxEw2AOqDpCHS4eJgD
6SpZpbHbInerqMkF3t1QeS6r8SzRX3SQoJWBPJz+/tlfKFw8nWau6KKscoyvd5FOIplkHGFS1JX/
fsoajQn0SZ2mcJL5D00+oI20n3wtQ01drJ4VR3jpPjEkudv262XmnA4Uw1nEqsW8B8JRXm6917Tm
mpcaxepvdkj49Y1Ycm6opW3i2zmYyZSSg1c1C6ypDWNN1aEd9BdEhaQZp8n5sigX9BtsGBvXE8cJ
2D975+UNeBGVECDE5oVfNYAGvx15klN9gpwelVHLDzbXNalrzgZEgEzQlLujgDzuMkaOiB46fB0b
4/WaSNRfv7hjSKxblLn80gwXsnFlh3FEHp7NIUaJC3FHTacWx4SXYNNUU30/NIqVPKiwp4HLGuGY
79tAhEGxi6tHE5Z6Nt56dEo1R5QqMH9C0p1HtBNpniDtz6Cjc6Ro4aeZe35Q+Uy0jTx+CbSQPUDK
i+6jxojMxXZi8Imu2KDwRT/INlSq//vKFZ8dp4JNAzCKxbE9Qh4vl5Ym/aZgLDhGNmOqIY3QtE8J
2qlPprAQ/otUVqOPqzMNzFCSvQY5DyPrZjsjn6q7XSwpdupxQfTrwhBfZN/rLijSqnPcap/Cms+F
bNCc5YuSu77eV6SLDTqCss80lSmVa8WYTb6FPnL1n/vK8ShAPBCxy5+3zFqra7nlh8+GmyCrF71y
9cgb0+sMmtV5GNb6pHax6alVV72zPdr7zSrEvYJMqC+00OAONfRRMcFK3w3ztJPqIKCUhWwiNwuE
H6llwBEHnhTDxFJPqogvqGOZUSCaCEiMDfD4SCU9piby3tq5cD7e0lMGk69Fi1izD1SMSK7xk1aT
bq/GTxXhnDIXXJTSofuYFGFIdZqE5hjuTHJGbswXh5xE5wtJnLg6rRAOBnVRORpqc+wf6vD0OPbG
7jW8lTuM8yyO4fNjL7cJh2Bgut9p7Q5HY58fkmzK6MG9c+jjUppqF5l6yCnGnSpXqIKhyC4SiqC/
rR4K8RKNBthZy8zz1mNy4fRs9U1zPgL/2BwMd+MGK2bEx5jPqWPnp/jXJA6iPzayv7S1gDw9DNF8
S9WBmVmanOcv4NprS651nVUP1Yg759fhsGHH5tW71RubUcg29aatCarCNt34l0JqbMgKAjFYx6Us
wuiUcJSvC227v/a9ZNpYi0C1pLcjyRK2RuEFji0lwq7zn0VHqBoHzW/KActOdB7XNkf32is8pVe+
6coTI4rVAetDX5Mhz6u7a0ThyrCnEzSYbGR6wtvN8uhrnjkoY4ALotytj6QCZbxReu60YQD1GAf1
POddStfZhee0zhinMvOLhgV/HaxJAth0TJ/pD1AjhRe+RdmMCIVTQI20EOIoadhKKEF4McEQq1EO
5gyJwttpA8dqGqsue1VmFgGt9eOmaSp367ftm1gw7U3AzIc/3nYWzMsDh8xMZWePvojM+hVd+Dg+
QVT8DBaPH0PkiQdWImm9xA5jujWSP5b8h9r1lTyg0j6TfoKdrEooxjkxeFZX4GLa81zYCJDaGXkQ
UYe31b+ooq3gckZrmRoExpk5dNGcc+yJSdgP/dAA7hbRK0IUcdHlFSVLiL/hRc+HZ1opqnC6GYgz
4C4kx4YY4kAVXNBi+HNXhIftoGetqe9r+NjeDBAki7cIzF0chBKDQVGrkKV0Q7V7VSDwg7br2nGp
wROgh11cmF6mU79nwNvlnEdJ+RGV0nNiTUKgzV4wEw0XJ2gzYp+2ZZZyJzTd4jd7AZ2Sko2teyQP
HUsd6lCbcckicrNlFwhdeJph83AZ/2z9Qr27fO9pYgxuJ4tBaEYdswfunEw5znQV7K8+8CQVhHSv
6fLhukYaK+BAFTfzDB8gvXEx6dOdg4SlbPHaLgG28HsIPEcWVeeaqIceEDGHyaVec+vfQbo/ZXMU
MukL3NB5lRj95sQJu1uPRCv/EN/beUx8ALvaegmWaCMo1HeTeuaD48zVonT/CR641Uati+rTbJOs
VMA7W2H9rWi2huMVbG1jhykAqBTZlPR9d5P+Wv3nZi2tfn+AoQons6LA9NQ90EW1xcP9phCwxf85
HxY9PkHzGSH5oUO6GkSmPlsjtPV4WCVBX5XKZZ7P1EmbnjEfzKOnmbmpkLr49kOE4F2y9OV3L9bX
IkFmd3Ul5a0H5asBU8Uoe4+pHPg/FQevyg9c+ktcbKUgEzGQSodWtDdRxezH6GPWIJ+86x7mFrsR
LgvJQ/2RE3SLfihPFtoZjHZ5JFNcApZfSqFpWbLc3Sk6nygXiE0ZmsBznBCk6d8ig40QxFFLYvS3
rTqY3fRvUoxdnNhDK+K6NinWV7/+iQ7lwu7I70FseBw1nXfGjDRrFrrGJ6ReG3AjWe/CXOH9InTy
hS2NQAT7lRq2HYhDKmWLOoKxFypQsYImwd0+PEhMWFO7M9y3NvdUGz5dDvQESaIsCtKRRH14Btt1
AnkUS0q+CSv+9e/+FaqgZa0yKDSEDfpmnoWqY9WYbGX98mqr+YOfaPRlupvRjWiugq5slN13AvBY
JDR3+AObJQjyW2W5erJEjSkiZrutvZ2B4iS/Wu4HhYT0akGjjcIGqJgxZyLtdfg7nhht3oJCc8eV
fkCb1CMs27NS0Vv9ivOJD4nZU0aZ8WdZVhgD8b6NWwKmURmFoNjU6jKpmlEdtwT7IzPaOgyHkBcY
0XvaQmKdL/khW01avXWic4PlB2w+xx2t/jj3cL8Krz6GZiBoNgMr2C60YujDpWZnM9PhLYPDTLzc
K0y2VOUM5ep5cDCCRXEBAu41BUVG7fzBrAGkvPb8UoRymp0G3o69iJKuXlchNEC7tHuwxLREcvqm
Ifs3rQuq/d//Ftxvv0+yA3tM7ADpf7LTQoTnJtV0KWyqJ3QUezHT55nOrayjnHDjBGUec193kTNq
heVgAgQPEYFcsLGr8qMBxC/oF1giR4tUSxSa4rayolEwa5g0yP1JgguLmRLTHopCf40yfCh4JJaL
OLut65QZxAsPIHcTvFCGFUYK+M7iimaopotGLR6hz7OK424p5O+VjPCPBlV98bs9DqUVnbr/bXlJ
iqnoIo3n2auh9zX3xv2k/3Vj4s5vaiRDKvE4bEPROlu3v1v/LrqQhcp1YVlCh37T9nyM6S+xfuvK
pPTWNU0Wpnmfq8yGDeUqnOD7FZhn4ExkrVv/g0ZkjKB4VZYGEwk77VjPJsCDVo126b9Kzed9HDLo
dvKX9/FzNoqpwF9WWUuYQq0XezOm72S/mZ8u4K6DciAmWGA/nMrv5soaQSDbO6eW87xoTQtVUj47
0qBdERpwbRlvMGrYEU7rWumc2UJiWc5IqtJDVsPgmt1yJCt1b1dQ3RyB6hTaYqJAuR5g5gBYK4nZ
KxJm08VfRlddbGVzxmycOumH1NnYFMg0tE/Ho8GM+uSOaHoJNQRvfjXz6dnZyA0CUWodJsAYO1ZF
MpCJC/vepojEhSRrun6iEuxG3KcEtfmuCt09Givjc5RvHz3yTYDyInMawUE0UmvD24RSo4zWGxTa
27dH28snlBlu+wWgi5umzNq6p2S7zZD6uH6+q7h2OOewTXlnpZGOj1+Araq+CpRsbZ6jHqhYIlj9
jYt6mUuQUgpxwbuJpb3BmaJe+JklGPz3tfYSn0PpHuCS7eCvHNumhY6ZETQtXI1PCjTURUioJOVA
5GAd5iHAEC5NSJo/9MRpGZpfQORAN+ifOPaTjyxfILXegxoBeFCePO1QPS9EXcy3aCW0xrxsDlh2
G7aO40GBkg5/yN56VdIf7+F5K4b5iNMNhDOKwi+txTfQFnrUBJj5w2ysStZgHfU56Bc72DJvnDWf
awGvbByXOLb1zv3uuBpdGhq21go+P5iTkCoil3DFnekbTG9L0POrpTead9pu1Ovng/a3GjQ/A1mu
YsabK6vP7GNPeoybI81gQrFMEjyxITIARf2LukBgtbIOSXux2LEKrfrlAPX0EbEIznDa8XY9LaIt
yNzNER2nk4ZlR0Iy1OAGZVSZrFSf2jlF0IdCQt81kuEWn8TRETrFn/RNPQsoUdl8eDt0yTCIW8Sf
2TY35gftYO7czbHTd9KevYnNV19hG3yGjD1wknLeHQ5Qex+LcVHgbiJ1q3DvXIqTm8jPqgoNAKt5
JM8/OoKQzGL8tfhfXKhn2QD35CWe5RizBZ3cKVAr/YmUrJeExCiviUbJqzsGihdX/VpSnB4KDObI
JJMf1cFCOozJNJeCjFVNapBPDm7oT8gECz127PQcJhb0+mzmStEvBL615fYyDYyKVKXVY6SDYMho
vhLdgBvIjxt6196oszl5CS/RtMUczI2qPj8y4McASp6ex/HKCrXelAQIzuNsEcYpp5lrybwKTh1x
1nBUYrc/vBxWSRkdAtUklx4mHTLjkdEx+aekHWHgrRQD5I6lt7DL+DPeBorsPsnFcfmA4q6kFcj4
+4vqsrVB04CeY8tBFJn7BTDFZTeWhfcj2H7/fSGNQRWljBGhuIMz/lAWadCycfeK35YHejWoNWWy
6Yo3ONnfL57WI+CR2xqlV09MwM9T7PJ1uU+zuwrTpmbg5Z3QGT2/YSn1vp8JcBb2/gyBLJpFycCA
XDHLi8cTzPDhOytySe31BOhO9wlHA4/GtVo3VrQTwmFtO3ZCHLrZ/UxEUHLXb4nrJ941U7ZLrrZN
26qEwhuJB4TimTUIKbZ0uggOsb9BcZvtZytbpNSar73RNCGzXGWKrrQXRPqr1TDv4U7qN4Ddy/05
2kbrv8KoCT4Ljb/kUyG3qa+FFT5W9aeRxvmsSvZUJV6O/A7bfaGVYMSfPJDstDFEHV0mvhdUVBHI
5vIgpeP/Nzl1uoDUl4jweoviEY/umMQ0GWW62/IL5wdH/uyQwlovP5otPCogDpfQOjrkuhJHZbJA
zbUYDw1lshN7ozP5XDohCNXTEKPxpOodw8bzBjYA2NcZ7w5D+BTGxhXJnwz/73bGr/OeZr17hBLe
EVOtM/nlBoHyVYNkF4PT3d09jjYrxs/o/M9EVb1EA9UCLM5cwM6o6yEMMRoC1+CnmxeDl20a3t4n
BPsB7qiNIA4tVifiaw2WV9HVk9uwcW1RQe38PjYDDsVbg+stJnXAQNKPtcUPz2kOIvNrwfJNd8Dc
ttHQRxSXjV5mPxDUrtoO5qG19rZRKun/JK4APhSgnRHRvPW1q/8wD3OXekoPlEtnlyRnTw7l//A1
iBnguo2D90rb4qCBNjgUuLICfaL8chvMv6TaPxDpy4RrvSjKUY8/ZqgW2N0+pP+lC0Up5b5lIUy7
P4l5YhAdaira3KHhe6fc68NcBpX7YHSeshjZ9lefq0Pu2Qoje6vC8H7XLcSV0JqCn/H8fS615RgZ
8GrSjy0KPoiFihbVBbD0yxYDtSjqM5WINN8sfQCj8VoE2MaB8rc4w1G+PqczHKs5eQDn1wHrvy4g
Rl0QVugacWM5TkHKFw7zlIRubwN8CyJtNFbDaDOnvbQdWIRFX4I9yy49hmApFqZvilg2KdJi4sZn
ShhipPqp43gRdDxe1XGs79PISWHCwOSy8zI0E/klHJUomvymrZSZK3lqhLLQEanc8YKN8RXD2k3m
ini/b4Sho92zSCTF9G/6BpBjzNArnorRZj1S1cvPR7M10Bmeon3OVEumHVdBTsmfetF8jN9K4GiO
xUAN8Qh+kJy7A5IPg5bLElMcivaeLKwsMIpZoVAC6r82dZ4f1QXRmOfnWtVl3lfl3MQSx/uaSnif
TkY9cC8aiRORxi18NGBLwUnq1WhD4jSihT2CTQHWKPnwhZabQAUb9sHPjsTITyuHdPb2DWIjcmfB
mcDRARsSSWp0mTuGkzOFZfqcJSZ4sMyF7zcG6oORA1bzR5A79fBMeyTyhZu+RneeNJgUEVxUqAMh
5IiCQDLXJVFj6gDAJfFfcoJYm/c3LAkrKbVG+1H4RlYKGR5p5Zw3Akz+M9ZkksOEymEqliyS/5Jp
637xXvpO3LgWI3gBu4JUr12mfCGsJbMkK39uibfLpsCYAEdSQSapFhHX5TcEmYQ2vkp2CxHdUvdz
TH7sDq71IRUa/H26X0pCdQjerNjjzvt3BjirD3879VbFMZ1KU9j66v3gtXtPEzI5Cnyr2ikLPHs9
fHpx0SJySEEz0Zh2vF57fnrdu9hhatTyiaW4nc7mFDLuZaqn3i6fUT5g1GqOdbMvLQWDyBPLDCea
5o5T2D4sTNqKH5Wvkm68JM3DVLqGZ2UwfLzuIR1MlXGmEsXmENNve7PtOzLRGe1V6h+LC7BY/0Gq
PupQ+gq2VeU/j4J8E8gCXCshRrXvaMPcaNwS0a3OxKNkDRLWk1pPLMBfgMGrPOfUpOcHEO2iiuZP
4a6F+tL3xGivrs7FQFZMU8HfZwsgAaU/il7eUO6x1S70U7VGyR/QMFWu6xF9hBlh+NA6m0RwR5cY
t3rh6njqXx4QNaYMQfo1rhRbg60ncW1QoQK7dIDLCdKO9hVhCz92cogNsZA/iCAy03qpR4HgL/c6
CMwkpDCjbTnwFUVEXiKrjLyoWvJ9RiEKw+e/ngokTNZ8Wj+6PKQVhvdB9ss4PkYVPHSFx6X7guCW
dcBdADccWZzayr5gZZSfXnHwW0TksQCk3OHljE36SRnl+FsL7qxpWqvDMXFfhVjac5RG1rVq17kt
u7i5+MfoiTriE2ciAdXnPXIw6aH2goZJw73hlMAYYxsdJGBCEd9KhCbTtX76XuGmj7a2LTfPK6Yg
oNxUeientMhpWWYhMo3VLSmpNxZJoKpvMMNvQSqwraYhJ0dwd4hOUCdzpocYqT66x4lu9SJ/4glm
aQjgUKbvJvJL1BzaBSIxFakja6A4ImQd8VdoIIAHaJxEFQkp+yWPFiUvpx/resnygl+9ao7WhCoI
u2qXWoMVeVCjp3cTeuxGhGODKozqzyoWWiK+PmwKpAiazjEMBH2slAjOMSsXR8SoBjQMPyz94Hdf
dIv7V60g+ht7kJhQ4v1/YrQL536cpzm1gCNCUl8CKTRsKQh7bCToGwk+G7422QXDCgKzmLlyyuxc
oipyXUeP7izvT+vd8imVmlEadD/qfcXgkKurvsJ8KVN/ht3gNAbg9CPmI8IM1tjE8qv3+wJljubT
PICq+Lh+/LYn3z6tOy7kdJl1KTUIYeEb8D1AMHOc3waWMOtU0qEbjixeJAKi2gNrPJo+R0wWMCKb
nHKdvxsBmfDzZq5vA8LoiA45h3Vm2E1cf6pNpBwlXdnhWUyOm8vuuUhVMZGLLcO1b7wvojCzux5F
V5O2RxtbSaHg22Iwox5yc4VnQxSs9R/sY70GCMPG17kz63pET5alwzRFL+V61rZ/CgedUGiaIdqD
0xfQLLKjPLOSddj5p18WtMJTYlZx57l27vEmNfEQgEv/RlMUM3qvM2juemnBudZLIpykw8i5jGzZ
m1oGkHXo1T9avlOO/VX4Y38rf5C9vdfBQXYph8woeZupAjcY06QguyN1W0yn5JrQa2z6v/j9novl
UpMXrbR0joJ4Dq1yPnvDW25/utAIPG6dU4ghoFWKARLsmkY3zYv14IlFlg4zSpEjreyxn6hD8ESa
0soWuO1by9Z/9CG6htCy7bXNrXJMotEsvuHR8d9+chyo8K3kWW4fiSAZWSpvw9ByfjjnBWb7/zth
2xLI+O7LAUCyPOu2IOVo7j+XQg62RF/LBkwfeaoadZMT3UJRCVEL2LmNLR73DXxAEPDdPlHDVMEf
hr97sZK3I6ZVZqVfuG86H7lTE8hi+xCHpWbF+VPqNjkvkjDUq5UdYx/yW8Pg8Tvq/qOrbiYNZw81
7IIcPZyqz19pM3UEwXDeY8iWRkVBJSaBhKara3FLlgLv2G22FY4sI5JBlJS17zPKyX8B+LHG4FMx
G6Pl8AGw9eiGXY0TczliZulq9Si8RMR0hvCB8DsTGdtk5SAndoeXpaSbZfE1LVxLRPFo2ytqx/Oo
Qx0PMQMOykT6IXLqp39KozlL/ZCwurWASjJjOiyYY/jgRo5a9gZVy/N70S2sLUFz7bzGmAg4Wr8P
Uqlq5jwCQuhu3H6o7/s4LCXaF7/w5LlMC8W0z+hELmZm8ewn8Z+6ixDZSKE9r/nGgve4q8VN6HHo
tZ23l8Le7qCngJMFVsjH9134rC7iinXqfOA7KuyxZNlMly0BfFt8jYX7hGCsAifhgAHXf6WqVbyC
3COulXAZd29j1yOeZZpx/QqUgJKQimZE0a7SENjsLcBylPFqNbTY4R/ktGKgiyGTyYeh9fke+isl
Cix0FgosDsL5yXB2EE1AInWAWLJnD3wBxDwP+c0QZ+8o/Gyx3Ny46RH7nbxN5rUneeA/acUj+Jrl
dSYKOtJnT+Sp7Np1Q3RcWM7xy6k4qYq87xX2+QVclw6zzry4E2meaEU+3qWISryhtMPS7CfTOGxd
ZTbH86iZsCbliMUkqOssT0HVqlrgCgFxGxW4f2IFkq7Ayomj0gEkQc+AqjMSFngrfxVJKQlpFpxG
cMVdbHDQ/RXrG07waYx2T/ILn1APCO+D60GeZ77GvJ4ewM3MucBvTJQrFVOspWz9RAhHIoItqZOd
OcsMJcp9CLpkOzbZWyInJgQY6T7HpnDThXXpQ4B6SmGdPvcwp9Y2/o234N0UNCoyvadFvhyG0hgn
O1GfLeNg9D7r0JHXbx8A3FEvCIYBsa3qS9gMQjianyUuOmqrBNFbdcfvmo1Fh7vQr7Hlddu62xMc
HpNcmEnONf+MjRVkYEH5QZu9Bh1TIv9dpf+KlKU28jYoKRs1o5KTQoKbAcsLa0SjnPRJSS0s6oqz
GsO3gL+YrZ4422UDGK67zbQ3Af3fwi/s3/wPbufUBiXnHkvbE17NEWzWWNZLaKtRlwfocqJbcZ0c
ebVqCmuvnuuAN6kibMuSmEl22rzgQZ9YgzblSMJlya0I+tTCvrAagD6xO7HMsFN8jos2x7z6bw/1
iZR0FiOPvLuy3TNVh9c+tFzkwHf/uxmTQQE4NfTm3KW6BPXMs2nSNohBiBMajhFfYdbTnwm2kgVc
V32PuP1oIjB0+3eh+bDVvvVMFYmzvTWIJ87j4BUEt0OOZuPtD35+g4OS5WW87znJ/AO5TK2daHIt
XQCW/mfHlw/gHkATPzJerexbxV38+7DbB6L+fjpO4SWGkc848TeLaG9GYREvBIsDhWdXO6UKIles
IDZrOqYBYJ581/6w5F+iPWEYKRmL9HIA9HJ3MC1SjG6EAwB1bVo7smOuU1NNvsaDXAqyVmiaBc6O
vvtQVDhgt6b3m6vWTXp/gJ1T6BcWU06EJy36Kh1S5hOOZkFjzsuBsFYQOefAfQagkO0pivwD4+Ry
lsfpqYiVGWcvI6Fz+yAGYyKIicp/uIu+EXdfWifILxfX3tfHQvNua5bcIkTSjKKr1VkfEUnNxLop
EyL1EvPw/O7609vtVxrJAcWOGUcTaU05jCty+6j3rqEikOrgxocdAQ02qvNGlFE3zwcjGsRjGabQ
v9qdkH1rbTGlh8xJxs6qGZikpsk1DzgFJ2DCsGRncauOBuUWCyHoxfLVPgOxb918AcElWzOPPdQA
A1Z8dEV2M+B7SY1qFLdB6o3oShtpRnSA8G2g5fTdRhOSjq5QXIp7aaE99KEf5xVN49dljilbIzJc
+Z9nuZQ75qlbYkN9YrpZL9QICtbCPR9BHtm3N65MYYczXycWzerTR6SbEshmUBrkVpLRN6smW5VW
zeOW2TgvrKVGSLILC6D7Veh+y1fa1oXmdKnDenT3ihY1mZbSlpYg71+tfJwWEa18tCUTWTq6/nS6
dPUtabNJ/FHmSzI/JyAWnn+RcP0NQ3IlbBzNYpfVtD6RMh6ebtkGLKIXkd2zEZhoTkIfHlb5irOP
uQSfYcdcEO27bqngVasXSScc9+hpAw9132/mW6wAaPBdt5itiGrKT7oFxvDliDjPtmqjOqOIZ8Aj
snM4rjD3ZSBovYZTUGAme/1dtD8dEZBIw/ZknfI+rJixFftZWwCygzAn0vv3BB9Y6f7RafMx+Gte
PUPTWwY7AsV+Kmb1SVlEGAuaIriyEdHhF2JY6a97XOhAc8IZAiFaEaOP6H9Zl1Hp03d107L/ZL8I
/r6PcglEufC8x0HUNF8Yi0GT3nyjfwEiimLqSz/WWtOT4h4UtmKjfXsR6teyo3Q/qoTH3zUxDJIK
fgixIYC7mKyW7wZqvWg01aZz65adwim6JRYb/MbICoyflagc5uOn4g+uhYoH8vROimfxSTsk+zyW
DrCyb00wg2tXhKpIDa+nAgK4TOBfPnCyKnTPsGOi8rLQVK+Pl0TdnY/5RpXBY9l9i2fMxM1cSpig
hQBApGQyW+ROczhtgRcm95cFQgGsPkurxSxdhNq9vpw/bTigPfat9dIt9znc05dQa2ctQdgkRZLy
BTDE+oD1THx+gM2YMOGI0esYqfhSxtCOG7fg2IdxRBUJns9avfqTooCkroTcmA4RXFcx2Ri/Nu3P
2utFPSCm5KfqJl8/5uIU2AuPg/0+9vLUWPZ2wmb9UVHA8yrqAxFBh8xTAWFs7aPFib9L6kEDqzNk
ZFRELnZaMdKDjFQn9cw4LgEBo6sR5pzhgvLeq9/6fNElktNJPs0n8B6YsyQCyjhSgrhAwe6b17Ai
jWX8Mk4rulHOVzP66XaLx6XUSf1OZHITxYYOdGz4e01TJS4qRD63R0O957JiX4DUG0nYC70q5QKL
wth6ELv7kOLCVf3PkqoQR0GXYFJRiaqf/pZ3Vs+20f0TqQf5Cj8OfMNHZ2nlunL6Gl3Nkz8fGK/C
zJRRnfi8sdTsDQZCaouTLD7OJrVTJ29OvocpPQWxN+GxWhb8wkZ09VVrvVdFp2+cAxgfPQUizU3g
7Vk9f++YdDZOCrUJ7er4ecQksLsOjFBs9bgc7DVx+tV1ig6TNpg+Ab+t9bp6fH+CVwGx02X3U7/p
8hOg9fG+pC/qJxAVG8SwJgskeyfw7e0icxG32kCS/u/UKkJgKh9+DWRDVMa7V25OxJx1ySWrcpjx
kJG4hhSfJKqQpjAQ7EVMjCJvVMqCwUC7lXJFM5hrVq28PRCoGmvWLBEU8D/RG+NdRigAHqOVh9N0
GhUtemXJ6XfkZ4ghGNBe95VuUYFrp02IOgmyPdol26UfvlfaBVE+DdIqkkwRbX3KHV6hqmcr/2dt
OfA8cQf3g3YtiGssjNPZCmxKB98K1J7N0lb6PrmbYVOYfa4SiwuwTLu18G9Q5sJ3oG2TU5dYgJsX
gJPyHy3dDki04/fo2njMtSadebbFa79p0TIzbLsoVsm51o441LSRCbutNC2rwxjsDTxYwfKGhxab
m/U7Bjcnx84smk7vEb+p0LpXB/iLKMe+dSPti33zG5d0+7EK/E+cOmEMwidDYiOV/dSHzxXTNnt/
owCkkN7XvgySDXKOo+wYOpw9SrMgq7RETNWOYk0Io76G/PK3wYMLnrNZSSCyYTjMHsKdzwBJZSTl
iLMTV5aOQwBPMeWOAv21vMrM6WbcQTnuywIUZsCpyyFs+NfFaSd/m1flHBlSi33Gg70KLn6oNMkp
NXVhu5hcnzDeDeeaGqWLehrygALdifOJTatqjs8YF+aMeAYPCv8gDAsvh2GWE2doFewG/ognvhpM
TA8pTaQM3/fZbiLI4uc5ucGVWMNV921dNPRwRsXH4ucHOK7178SW+1QjJsknUZdbqBdBgCh9QkMy
w5HSddWSNp5MvGXmePmBkQf4aLGvk/ZYxDyZsB790dlZIcYrP3fOQUwvggufSDhCCQs8lUvUVPKK
gbkBk9So/gE3i9Z9NJNQkKEz7pqvx+qCpSOoRv1D/Ap/o5KHhW83Jsn39AdSoRd3RPZUDp5pvDbX
YiVuAL9jwDAuZbCY8p7rLMQQIrZpLPsUi6ACQOfErG6ocmatv7fcViM1zlRoamzkmB+Am9WacJkK
Ke/SfxyE2D2D8CHbuvzPSNJ30/uL9FgwErOGfQ4RkSxLCk9BRTxhVBhC/5WsZ/CubkuyXqE1VIOr
NgV9WQ0chI/y5W1f67+wEwN+Rr0XV3sOq7j/b9y9nopmuGj4i/nWzsml3XZWbQKX6kbH78x1kkEi
iaIHl/pcbrrmz7xRM/PjG/XL0j2gqwfNiGiJPKE7Jr3gzc70n+U/Cd5ECiM6LLpCxIyGu93MEzmp
tatcCWwFKUHPO3WA8mdpHffIrNznEVagJ6JV+Jmq3YqHJ9ONPrCy+LRf0ZTZAPKs9lTtrSttrv9W
sA+SBhCZeaBTR4LKURLirpyTarcAeEVrD4nVLmHru6vbHGbMe0GpAZFEcpMmExMTAJZfkuQEWG0c
z8LmZyP7la5cQuaFtoZr9Y444COyEXZB0wtT9Jbcdz6HiW1DXBOOBJbub2spHHLNPmMMpoybmsiD
Av5aYOQdtysIXEJpnGlK9dOqgwbtrT7p03dNYEuNYYqiVdBPO6mSR017J0Ie15diE9qwPMk81LnK
2qa7qe5yrstNSfjVhd4MfT/5hNQUtCvLCWkpLKelQO5ZeEHsNKmuQkElOQNvx5nEylNbaE3cSVQP
SzjJ7G8VU2pByMjULL3ztiGX4aEHQMhxSc8t1VLi7D3yw0h0XWX10gbqQjM8iylyENahPfdBTt9D
wbkIYKIJ+knHTDo+GPXSNcfKrn37T90vi4ez3eu+UaolaEUxdpF/9+LLnBXudGYD4Pm4wuw5Z2d8
ySWANT08NfLGCvHgmIHlEyleiPVdMUfb8k4cq/accl6DzAK3AYy+Q8IQ4ZEp3EVpARUjrmAKEe/1
I0gm7eqj3qmDlkWlvDZjG1fPLfz8AkNSbIvFBbDTUT4zJlqY+mDYUUykmZKoR1WtxodjUj2Dmadp
L+oosPiknXywneWLMA66BJwr1xOM9jMdvzX4rx4fBK9sJRvDmmufcKPKdV6oLe9ugVJIhJoprRPa
n+k/hyRsNj536KHaFb1oLrDP6ArFvf/CSm2iYjiVUR9jXdOlPMe43XQNd66Yw77GQ2RqvoRKMp5t
+j0oAyX+lXAqITaQAgz3UsHmNbnmDbgawmSX0iBAWBtwyYHyW8o5buEw67lII9Xy/B5pdPGVAPJP
4oj/+PeuwTKImQLf7bCix8dTDK6kik8Jo/s/ytbuAWJMWus7hdEfueL6Cjfd5gESKn2rD1u/2A3M
BPUqWXhOGj3nTIuF3Xib6+RObhoPeVGpj74DS7o+VRsaP32W45CZYLpM9orOcOgtLAs0vUZ/oPXz
A4/f68shdoQDOy9S1vshsFCvP04RDP8cl7oiIOhD1akp5STly7n26OS1yJd9SscUSh4ccdkvsA0Q
j+3nQGiD7DbxgGt+1UP56vkV1n1I0vGmG6mr+Omfuqr1dfFJRvOt66Z3+BODqN4RIOvzdwvgwtdC
mrF/8zzlKqnYRLLnhaTIzoSWLDBZoKxdu/Jtf164SeP3xmRRSHZXlrNDg+UvgAm1076cfGYtkBi9
8/pWi3m6ZiRNJ78S82pbLQxQqjSnNIj0tf/vq6Hpj/NuaJa2fDxSSY/UQhSXN7EB47U7kSGCNdnd
17UaFaTLgwoDoPGmdHjn/JPV92DfOsde43xsz7J3HUPyZoDBITA9qUhCu5q6dJ8Iu10VkzYF0Rx4
SxUBm40iKXYAE8QSW/hvlBwE5iRTESD4zK9DWcPSV0XWHZa7auS7AF0mejjAIdnHlT9PABgQiGX7
gZD80gIAO0ID9hX+rTZ0cc46T6fc+QB2vBoKYjxLqpByOiyZMYjmxWX05FtNfHGzcDLOqXeHBghL
U3akrSfCTnnNHP277wni3W45t95pn2eMDILUdyJEwstIYmu7NI3wTDil/dvxv9TsxAtJMpo9AiLr
ApuWJkZoGgwsSxUyR/CLTsmL6H0glW2sEoc5SeG6kwlZeJiSoXSLqK4MskLs7vNtrIv6gilI86AR
rCpzQoy6mzckCSKKIMFePSP9QzeJZSNeE8AkBal0UJ8SqD/I07KpyTke1E+hrFfpqNVcydS0oDtp
bkBrurpO1GHC9ShmbNuGqvL8vo0IJFrYDKLIUtFDf35VkjZlUBFdUMyRezdJB3B8vBDqx9y0+gOw
ag9Zk0ZI0Yjf+gPmHgfWKZu9QTcY9bQEYVrt2X5/QBf314+ZeR4xCCOs9RhjiJkCCIA5gmXv6klb
U+tYgnavNPmAxFlKf7kKuMnSODMG7gPD7Lttz08+VUKY0TFhFInjBdpbIebyRWRFT48zxnjZMexx
mxzklG0Pe8BaUrn2Zrzhfw8IIllpJxkJ+BSW6wBCE+KmeSnxGJvKaqvjFLsqwwntqAWqmXjvHEJU
54uJOM5XZ1IaHlRcaYYOa7b+7QmJjrqaWb43d0YI7w1rq3/Nd7DrBDS7T1LlaPUPakJAWUiWKIOc
CoRhwSRJ9bQ/aehdmN9DhLZ2EPfhOmJDBXv5KGmNBxmpCkfxlvEhJL3diFUXGP9V3rx/pOmfrUcN
ZCvlUHumsuGQz1jk2PgTbg5d+7ks9wJcWDQGtrH8grNvltsbmWp3r+7Q2YSbvZQwVYPNo1kj5+wX
JsQpUHdtasObIPKkV3atjZKK5hbv86/Qnn34zXJok1VSjezmiOFEvtUBbVI4iybsEQ5ZsCg5UunQ
tqRSLSvHdhjT6oUFezKSfD6q3yJvlGHf8EGzASBFRvMRvdnLnRkhUPyL9n33faKs79jVPt4V0ZDv
uECYmTbnxEaqChxadimKmEunVC9BL9R+VEA5/1FQ4MausGEZ4c1FzYmPj2Ts+RPITOacIzdOWcM9
st37gR8HxhFnjmKy5wMk9MCGk2aaWhf35UQA/wpugspq16VyFw7iUYT39xosL7Q/C5s3zOQlbZAK
XlF4h4jHCFtwDA7QLXLoFvZGdp2w3YzNzhzVf1ah40+avuC2cvBeAyWTz4mCCaMMcXRpO9FMtCQX
8/vYUORzGqWEZxw3FdHc1TPbkyhJjbB3RAfvaDkePLHz962P3XzTgPdHgBVvbq1R97JODxc6RqtH
Xg3sn1XSxbXJ6exUxB5sDmHQT0Uur7RA4VIk4rYToLX5QvCc4fmw+Ok9cIse5OlE25ohQVn1/DAs
VsBVDyr61Q4ysRLx2zIfuXKu901Xl53IqsW9sPH8yrB4N3g4avlmNERiLBU0TqLqhp8G47+gnOZP
ijGHdOsYbtzKFuHiMnJoyIls6IQVyWzot6mydR4Y+FK4GfLVGlFvr/EKpytZ7RVFv6/v3FuEMmlc
+sXGW8yCE4nZP+D07LnTtEpSJAvtX3P0m/ZBAQ/HVsuZBvZAY3DnD7nyW6aMqMEwWLuf45C6jRnR
P025oJ7ODUJOeeFHerpA+CFzOmEiLumQ7eoJ6fUCiVq41b7rd299kzzK8mvl4YmmlPXRVKjnI7Iv
0RhUAyPWxxsFeqOdwO0tIYlLUTO2cGfbEabIopVfY3r29I4YzQE71KbAn/Qivg08ey6XUDswjKJv
hFOcLc3AEoktJjZ44Ei2p24lD/GJd6bgOVSDUgbjgAnTV5A1FzcW2UgK6L+uD42HtizjNLLaNxfX
F8RkTvF3Udogyy5ac+pNHiFTAgqJ+TbaiOjWPzAQoTJuMSOm2B3kbliFQTSFvnm0SDRF3KREPv+y
5YiPXbsHtzPZ8keMbSeK1jU9ewpDH7axiM7z6r7I7cDDlM/bAVUAOnjwI3pwzyrBPy1XGf2TmUG1
Yl7JIEgE88bxXzXBCtmdtykr0XP9In4z2ClIQHvJPuLe4Ski+h9ks3/OTf+6SIhNH3y5uC17dsqY
Nh3VJk8FF3posK4fudkganeI7FA9BW8HZQzdwRgCf2Ks8AE7/IHK+q5ZavoEcFTsZa4otchN3+sf
Cv3dmuMrKDZ5YOJTfE/hrWgEb//CKgLu9OrCcFRbRYKgnEfhoK2Rw3WfQxbCT8ZUWGGAK4x4hSef
9EiZY/rOPlOydw6QE9T7K4/hz2SbrOvU4P+OVPdkeYGuWh/FRMiE2iY1GlKSyGjMKifeeRQMN15h
qX7epRsDmgMuskB3sukpZsCIqRMIx7LUZBV03Capu6KVcf3sWr2KKG52c/i5Enzdy6SQp0UB7Hqf
Rkr1kT0oqqMb0d43hsIYE01/wkFxa8Ml9Jn0Apvb56tfAGFskca1OP70e3gR7nciCDYiiFzBYz0S
fxLY6HApxka9AVNApBs305nJtfBc9KQGwI+Im/sgpbZdQNQVmARj5SEx1x7DHKs9zx0RFXxZS1s8
rA8Zxwu/MkOp3q9oHRS5nx98X+9rbgPsv2AoHUHZmjFT6jlOBkkAQX3UgN3cF2ZblrrjVHpm1ZZj
FFAPWWjB4eWYEBA2/WsaJphlbDWOghbgLr5xSl50Ps/2NY34Zu4ZCxgQ8N/jZ1df1DzZzAzic/r6
6uwLowRHJ/HDfnz8ufWmV1kIT6/IHkyMyjhFEtJk2Nxfo6nYl2s8hD+P3ticgOn8S7oMzl79FuAV
tIRrIWKIsAJwp9XqpYrd3ZFbtZ7QZj+ub1XPJvmsrpRs5LQN80dxL902lOetLt8AYqAMbwZM5gUl
hiwSKUbSFI6Se7G9x+kaj4KxwxCS9tU0ZP0ex1hHWPuiiTTmPeue8OKG3Qq7XvZUlf2Twln0yWLv
aQMLfcf0HiawnhkTpGF0RN/eU8Vy3Uc/nim/p1QavlaMyXPEu8tuCLyly2d/oSdpxkp33K8qw/DS
OGHDq9vC4YQqLM4rq4wa7nwaxnFILysB/MS0gndieOv7uelN6F83he3DlUia5t/w34EDhP16w0x9
PoxnIUu9RgLoUVPMVMuYnlsKym94GjdzyZm4O9gBYE7yE30vCh5f+m0rM9OrggkwftA389y15Sv2
IzGywszo/OzQKGh4eITWSAxRz45y0O3A7s4DrDPUwau34d1PwXl90dxIhi1t0aYCZZuDX3PvHzPQ
B/E6VDVdDu1p3MYVg5oDcgO4h4wTJSUAs3sBYEqMMgjXJORuMVQvdi6o+9aAb8xy7qjm9LjubWfs
19l40fSrb7cN6QcEBg6bJQS/qeDPJ7WkK9CsqDtSuWKg4Bqr/b8iliJ7Gpmt+uykAHoON1WZWTB9
yaFJvzklDWWjtZxfRFQVXMDoSV21cbmM2qsyx1CeBkG04Db3af94izcfgnuptPzFFbRF+Gwgi1XZ
ysJJBsPSUqkuHSi/cBPXS22hJAuDzQSwbUSCi9Nx665fskTihcz2ICBTFVwdmUAJAx/CNDW3uvDY
qcNrbfzD3K/KV4srWRj8kxL4R2Z2u/myxVTV7QpYL36qI0NnvHro38EV3FDjPcyHYylDv6XukEVt
kz8qA322OF8g4tpv5dbx0M3hfEwCNys/tdwtn4LPFdjaFT3kxq7y+ryU8/rzz8xe1GCJNPpcuvVY
gOlCV+EvMFoRHJfmOXADpN8GPJupJshQHTQbmPkgtyhHCA+sksbcQSeSHJ4fGWZwe3AEbK3Yv7aY
BxIUa/s4Vwq7dRYlZNg5dhTeYVhnMfqo0kSXSQP/D0cNQfnnF5vcKPV58Q9CzA/M9PQN4IDXo5zi
gwrehDpEb0FwhiNBf6ZJTB8prG3aNUj17k5nzq627VyCZfeEuXZXl00wkr9eKicFy/ndVLYBVGRv
mRW/mVeuWTjZTF64Su7XbZ7Vp16j4fSL8Si4tIqQLnUYJfDzK5mB4CrrlCrwmuwY+F1RmZBqBI0R
wUkCuOuQ/arHrNkIMe5wT1ko7Nf71Vto1jRPK0kb/G2hYE4TFPRMKeNUJsvuoVVmRA+MRFsCY6XF
WUjHa5w8dS5oWJ6nsbLf9J1VpsD19v8UNRwU1/WyEZNjlDMy7cmqUV8dQjsYAPd8ujPIuHIrPuO7
litDo4Q2A9oMlQgL8lZJEeOVTe+Mn9fTFgxBhFdP99yDKPiJvb3XF+ww6/ToA1hGQZuNpI/KZ9Jb
QXUvV8fBJrmWLgBqyl7JiMhyzkslbJ29UCt7GR7VO57dbKsKRkI/ZvsA+wmrkikLKhFlTbME7iY3
AfUXay/sprlfwbFXXaBRv91uKixqBXAZaOr9Jpwr9xF9ygVJ4z4U57dHLr97OgyAJRxwQ6jPih9x
PLD9dmt1qqdqB0OOSMlzMCOsDajxRPbX+CnjAmBH85DA7747GSoLWa++g2lIATZObN9Ip2q1QF6Y
Zlb54kzm/VOVi94TZy/qOXwyeAeYGWPZ8ZMX190ZwdEYTvJOXkZ99kBiu2G/H8tZXj/BGRUL0aC9
KI8m4B0NOfoSLefQmNPQ8SVaJzMZyIIgY/oi0lgkr5Ypu9UZIqSqTVQ7PfrtPnIE1kiXfKiiHxv0
N7GKG0WIP0TdVAUYZqlizcTzNF2u5cVsfSdeJLT6C5qryRdUPYhQr61Vvq9oTj/Ekg2L3QOd6/w4
Moulo7jiiGTvYd9jJF7eobwYfB7CvlsZgSjrxUxc8wnbl+dU7MlQg8TRriiqP8oksYBFHUcgRzyK
BTGMO7AZD4rjgOvLp2h2EP5XdzyFbUgNlTPNPcI6jaqzSqqztgRsuPxC5x9xz8xUDHDZlG0C14HS
CDes3milwRjPSv9zoQhHA5CUwEXFGFgug56p/tsRNeFJCvH6Bu+cSD/c5YqSGymMbO/P72lEBSft
snsD9IUS254mOmthvCB8Zi83bTCBf4zGxc/eWVNVqgptL6FnlODFTdBHTbmMzl/uqURiQyfQNhSY
BUKJ5CMmGP0UY2MRdcmhvOMTf1Amk8uxNd9FzQjHoXOMHKx+Pdngi70bBPOQOO53UPPtQNYeElo5
HVp32uO8ZJtUI29Jpade/mbHbNFZcWnFwEE0NtB0jT0JyDm/R0cBSIVl4spY0jtszx75qmelrnnh
DMKMcg8xkKfK+G8zWNgCwq4bPuhxxF/YEZSlX6BGFCpF/ReEQSvMsbyP4GOqfjkUfV9QYXhQup15
VbOUMWJoJ2HsK/2Y8Bm2m4IzHvShZVCAeQ+31o8g6aLxqY/3e1O118udYdM5aiyF1J7rwIJ9Ox8/
oj+IpRHLYbEWrhzrl4W7832NEGZEjhtFopzXg+//LP23Pw/OHcx9d7ipmeN82tnLTFccEnQc8KhK
N47mfbJfPAwaRI26TuO6wdcrDc3yTNldtxapBZid/VHfjbwAPPZS2/DNGXFLC+OPiEKoV2eEpK3d
WN8bT3vlxbq9PM2w3VXU3BWzUBE3uqxHJwwo4qpS0IclFQkYR44j/5Y3qfCQoaXf4VSvOkyMqdRY
R02RlfRA9WOuPN/4Lac7+WiFlVCb53oHKyaP7uGKt1wP29E2vmXhPUokyBdjtt1mODMx95Ju8ZSH
W3kJ/dvkkjffSb1BQDo3Sk60ceOEmFYMd93e9+twNCsi0k2Ga+NHSfH3a1OHIBGPKiNG4oMlMUQi
qtjAopuT21pi9CUAwOtrU093m4aZxoJ9AGWnTPrh9Ly1c7EcmX/QORdXKwKd5U/C5wB3HDPJdg1m
1crBnl7+osgjLDQRCG3JpWaOQD5Dn9Da2mgx8tJMznaT07eiXI99ofkBw0SqstsPy+X1wJi69Oki
Ne185SlwfsZdByaGddGramkxf8ZDViNo9C1PEOjg3PQN+jhfpg+JJlO7xBsVdZl2S97PwvEPb4lY
ayFnHRUcBeSDCH2v5Dixklv3UzkLUSZ3RGbTTkkt0ncB/bF0oHw3na1I0ihC9lmsiEOrkm3otvdF
l1mEAlr1hhzcu0WkjRG74vyvN+8RWlPVBxY33i4fGpLYVa9s5IvngrOXbsbK0rO6TTrZmoSk9rbY
oBIMIIJvSighblccFxDl0uCCeTvhQ1ZFWYJtkT82xfyDyLR0WSVboqp4sQhwRXM1BTNDdE4P/4hg
Da+YI/DwP3era62/eRHvFWSC/QLdWJTjuJjRPucjtQss64ezb48dIImsFCZ6TkJzP3naFcqMkltM
YhzpYOW6GOsfoh7YRujnDeIcM7rGeQo4K186nlB7wL6PkKzWDEaRXsmni7Yq+Tp3GHtaR9LxRwPO
4YKDnoePnx8l8vxL9ViCntpDs5KE7+Cb0m+wMYDm5DrIY2dKLKBoptT6G0LO9wTAg2mLnom2JlrS
V3gD/nsr2pF+Zd3UZ5wwNGOWwoH9slzGJmq6W0vMvD8MBm8F7LtJjLaerif78GFe6YBKFPsDwWV2
B+k2+dTO1ONFJPmZAGrJPGUWY+31Q2FIHIoy/Pt7CaSEw9/HMDCyzAGXgnI0qmiXHOKLP2rGVQhR
zF5TVwO7itxrZIyUv9V00L8jjkY2wZrWizEzb5/yyrF33lnfAplZsLL5L8Y8ZDy6UwXBrmxNGxrM
BODrkygA5TyAKo1pixzya31Z4S8G6hSbvrq+NwNX5NAxNOsk/gkWK6ibMByWiQNT+82YrncEtcAm
/LE4J5zft+gb27xNoT+yVI8IMHANXyr969nmAfqaGA2Kfm56RnDyLHwVM3Jk+rC8fesoQoga790J
ngPogSIh//xdSFNLh4lIoT6yHpdDTAqIcf2R83qscnBXpIdlf24j12+M6hOL599gkrJ6KqyQraYG
1o8xaW7HrIjbJUaasU9oPO3mUYec4MA3L6wstWQV2QbGmnDqxyEVXltg3Hh6EKfteOhJGcNlzz1F
Gy41VQx2hE06uSoVXBg630GzsfzR1TctXp0LiR3pwqyXh/HaNYpJ7ONzAcxBQqzOfReUP824wDl8
ftA4MHXc/0U34D/xldWk+xNoQMRA0cWRhGAgJRVlRP6bMtPdgRa82ZC7RxDns2GT/zkkJboTIlMn
s9heP0qE1+35N38cRc/gkx/xlzHeAWeqie0WCEBhcDonJz79znWDPJFsNqsWU7TP6IDO9VAVixTD
BLmoBlJCM8BDKkZgtVCQL0+pdtEWhbzqdKKMQmLz+KXatdOGij7I+lB2qp5eUmOi30gjBj/uuyku
Zaq5VnQzgBmErqaEtDxJvJ319TMRu6DPtym+mZD/T7aLX1mBI0NJW0O232HJPNqmQ1bpZaJvC2tD
+2LYEU4PmcsW6Ap7iLwohpOSI7n3UTp2umGNV3rklwWWAjdnFLK4j7gV8OXpYkQbKHlfSzbOw79L
TCiROWdu0lqFl1+wyDQMXgcCR4TJX3aYvorAMpCHVtvBP3fcaGRE+NiRdZ+Mfb2zRMpFkDElUUO2
YQhafM/ygCLs/Hal7keHTiMm6Y0c/DLw/6SRiQEfsCjsGlbyy+d3kZLLauqRetqX/IfIlENt3eUV
v8W4aM0fzsNvt5PIi2MSiNo+l174Iibk553QI3Erjnmwme78I5/UyrpkONnNmPsjJbPmfU26w371
KWcfZbrvY+26Vv4Sw6t/69QUX/uAGUINW1U7v2acfJTV84PnFJNYbwOrfJ3d/DL/qrub54AuVk+m
fJbHh4zLaf2m4OOG+5GiaTg96d5pKdZZBlbRfaCVc97wZqb12Yo+DDLp7FbZqYXBgDEidCQI8nfh
Lw+kpJJ+pFAAFJUtoEKwOCa2u4Pf/yv1Lnb37tiSFCDPhuhpK3K1Mq0TulWmM0y+VVb3jvmOqbaq
YfRol/AwudDXHvfM0qODqiMBm2C6wDd/+ilGCQo0bdRKhgC66tW6hNPNkOyQw3HvHmUkwhptzQ0g
ABil1c2BMB/6+cJm1u1BMMiQZTo2/ZEPLSsEecFKRLmnvV3e4QTMX8ki7CNXSgW1NOy56W/GTRnO
fyLGdI5ToAn3MRNCDkBaWbBo20ZMassUVnZPfvvSnLNCCKMbEBa9wnuEfkwbpYCH3Fq2osPqIjbS
7ubH2bbWoXdS3/M0l4iGJoJEIa2hzE2VmTIh+CN/8Y/6tNg7iVeL5+M8PSH5c9a2wt+AAm+w0Qq9
oGLh1LJFId2F77uVAJZECVqtP995SPOGhwZqaC+YnmYLL7DqOqZfZF/WpxKi/uRBqji2UQ8Ucgkr
dDgRMgchwQeDTwVN/fd39qLyCFaIju/d1lJBOfQZ6Grvx6cBFnVdgg9vY/91FFSlK9Sd8T2Krw4E
W5r/RHOfxCHndR9ZS4+bAIkw/zPMFPscW4PgryZRPqFs1fT3t2yFwTBIWU/yVAKJ/vziN7CQd4go
Aa/1osINClZBt+Vqf4QQKoHFfYHjsghimblYxDs25WG1jhaKKCuExQFVCRk8Bi8CajWiv+ZFjvlL
8a8o+feLKlPJfFWT0P5I2GvlXaeqGnMs2MTQYkpTpQb9ifp+8XmHuNb58WoZn9eG5y0YFAgVD+Wz
xAz8+wqjHp2GfxWcijnIrhinBFIjtfLFPThK2R5ZqdzPLMOppUREPhTTZaN9jWdEw1vAVjIzJQj7
zxZsMLOeuaTimxO7HGfgORhsPIipc5gJ/KkTuluYKCaoqxWFAf4XB/cs953bS1A6ApqJ9m2qeCua
ASyfCnPEtKHwLefu8ZjaURJsLa+SmL07tt4Zpd0z4WIkz7zfFXiuedNBz0mf+wfwPr71vxVKZXgS
5TsG/ZOKwecS0lBaCp+557pfnIFRauXEFlGg8AAyHPJ4biQSeM+uVxFtLM+/O9wPdI+9le10Wk/y
A9BchEpzn07deztKt2GtLWKzEZI50wxa6cXI5rhi0vPPGVzRIvCtU6/Lv9XeBXX22RSxnY5z+rcx
D/gfIcGYX9p32/VWT79Q+3ooqBrR6fG+SLz4rp9tKZH82lDp9Lwll1I33/z9BYzs6HZAHIy74AiL
vtgcL39SUW5NbPjx0Rm9+F9D9AZ43aZn/gmzlk3JWJiJ4HzcVWXnMu3VQzRLsbgU2YnkhPJ3Xtdm
WdYCfXe1f5oBbmmymB949JIgoNm7d3BO9iV4s+RzaImTwvIgchujuCY2DkpPz61pIocDJFkzZg0u
wNv7sxMsEn31V3d+JWfexT18be01H98md7AtrYgCmamBHr3tl4D68QdoKf+HAFurz8eS7IDR0gHA
Jw5hofyBEW0C6BgpmTNoikbvDo/Mk+eCqrpYnovCUlJoDyFZkk9SL+g24/WQ20KadOTDlJLPTRRn
SjrIQ+8P00xcdNkJcKwa6N8+vH4d04IFI59mvgiDMQ0T/3T4p6izThXemKUbq1yxcH7nnF6n/doz
DtF4+wDKnT4vNqMFRWnDuiwEOyP4q7HUwdmCEXf/gpeCpfCDZRIjTiiFp6YcSbFy7hBc2/dek2jV
dqNoF+axJem3V/iQOEdIWqUcZgD42AolrgUHHRwLWwF5y19+9UlWuPuHtiuSSQefZ38z7gRgBPRt
+eLE9ZFXfbwHqtvL/p4ALPAn8Uc4gxyrX+FlPf/jCdMdwBn7qtexNEa3/pC67SOvVrdSWhebljfN
D7fQv0ezjM7Ng0EhoJVXgQmjcbYxpbCn+EIqIEe4DFWcq+pWGeee0yqJOfx5s0/xmzkity4vDOkE
byPKKDZU2UQb+eosTLBqDZT62t+1yOVutLhj5OASYhMJCAmovqqpJXUcaFaAd6pM2I40F2ojhmtb
1YUMpDzOidxdngKPK63nL+eKvcu7jGDeYqDdj3zjzbYnuqEzDBHCgS3L0OnC5qZMcD9tqq66yxzd
2MmheDOGedcUPBcxR8/e8uUrhdITdZvV/X0yY+vuU+i5WXli9+DWUCW5f/uhIiwBK1ucDo1wd3lV
PpfCYKmHfXKkmgoHF2+sTMkeoSs/zSfZ8GsOxZ+209yBuP5X+d0BNN24dZFUZj+1ho1Yje4oGrmX
xHWfAHCpj3ckiRaDWglOqO8FQZhiP0LSFPD+9408G/Jbv8Nc+8NDLeVyUh9J0rTpeZ2e3Bl5UlHD
mCNtIlphyUBRWH48aHgvFxQIJZsrVLXGd4DmtdhpRcBrllb6qqfJzGBqEtzKOT4WEJQ0vpV7u5OJ
nvpRCV4t/BiOazwE6GM8e3Li9Yb57m2plMU7tRHRd2fqV7ACqJ4Mq0PckhrxzqyUquIZVRpWT0xG
l0EKlkSuTsuqPfAzSsjEhCjjI4C+JuGxkLKkpEPnA2bhofmFrUn+Jp/IYZp8TT5wTUwPwpzaQjNd
jDW8nsxN/VbQlqHro+ANrdjI7eFZeHuJL3pd8oKCtgarLbIvV5gOqlMnMTUW2nmmp2np6M8u0Zjk
F6n1lWtvvQoEwhi+ZjeCb9pzyHCiVVsHilkDOdqwvdzheXMuzQxcq7Uyfx40NnzRPcAh3IZ/2NiZ
0KaAvsRrC4516PogcG9U0Fdp2POUPNWkoU7CBJlwejhOXcbuR50siszjCSXgSp5dn1Sgr70Zx+3T
LpFQZcK846DLiCX1OqLE3c15LvdhqxpZOtV+TRYlkAqXJLPuPxxcb7ouTfKqmbzkrgpOHZXJa7xX
OAw/PR7D99aW8u+JhZjkAMvY/nbQ1hED9Hwk9D8lVYTp+BHjPtNbXCymClBJfZtm3oc/Xaea8L2j
/UD2h1aYiAmKgcO/63Vjh6GeHYNy5IAO48wbxyPZyJQXU0mwrI2UHMXCNf/lNhmLCMHlUbbqr8Tk
ONJoKMjhqJ0e9VYu3GVdoojvSKKb4jBdWeJoInFRMBV/TjDrHFyewGPZT5uAWUObfkxPyWtAaRgK
JUI5YuFQHk6443+rgVsf7IMHDBTZJ5mVYKOlD0oT7/+lseI03w6TkaZsjJzPvFDklkgRusF0HGek
mlQt2NjTHnZtcR7JEvVWXSTNpd9GGcNDRi0JF2rzmrtMV+ZndhEV5F71pP5nlFxX1BEJhees3x/v
OTEkto6fs3ru/LNi/ASteDBcBssKBIs+wGyKKGJcQfu+fEQ5rxnbVZ8t9trz/DijBIHuoE0xyvbX
FwlCXgen81AQqHkSIeJ1wZiNToYDlsQQ2K3DxvPHzec0ApaDglMwju9zzgfOA2egEUyv6h5HB+3/
tF7gSFqh9T1dqdMSaT6vqfFtCta8hsPXAgDuIqO3MjzI9UFfqRCJ7rJH5upUJ5uNPQadgcElCP+9
YUx6rujtq4MHq6Oq9bU2LxkUxhtF6ewBvO88QhMIWAyT9YL/0DrqKtALKqGtC7zgHVWevqBvNdVN
/c6LNH9WPSfIHQ0kCXbWsJvK7xRTHQax/tVLRHAAiRLkZhpdrmZ8N1K3WDj/AZTPyibx7qAxvpDr
fbeNARJ+RD+tfIxQGnVChwXNT0mpf8vVnlwCYrPPX7HmzyVsKgEHW9X013fXm50XXAXaAEpmObnC
7903srvvwdrn43edshQ4v6LdvpuwyXOtD8K8Fo8EnIjWd2inRwLtfA+CmnCzACEoerSDU0K+2msS
NKxR7dUVBxSsOn+iugjy1B3GoyElG/lnBGrMkXbPP6RDM7QhNJW1SLmoIXCn4r+KAy1WLvYnmnUp
0gI0wy0GhGCTm8jJaG/eDWEoFNcQFejQm7Oa6A//RB9lrUKAxQUOVgUdV0xbc3FefaLfDpUNh1uw
VyeASFSsgtA8OTB2Im1HEzsy7FEz29Nl+CFujNBzrAcrcrriyxP5R1DiAjXjqaCUzvGzlY54e2HQ
GyOetv5VxrkZBWfqvcPJoG0tDhrZxKDCe4vcSfZmjAErMsX1gh7ByQOGiJ5rRWmew8F7meRmXYBo
xlXAcL7Ry2c3V+yUFe/kFqXqpmzlWdSNcwWvBVthv801+4Ri91QZlcJAhH0azl67AtZU5MH3pI9N
6GsFbfRzxEQUIVheYGhVL5aPoRUYr/EiMMUPV4J2q2g8ACT55vsIGeU3+voLTmiNY4pGcj8g04n4
bRvDWZmvi28rgI7pThShjdwc6/K+jo7FlUoWq74pwcf3wH9nQiQdGVbdZJGkAtbXAmL1C1mVc3KG
kCbjpTu1H9eY1DsjKxMD8YuaYO7L8SzgcRp6Azy0taTHwpJAWNtf30wTTWeoxpOw2pFRIddnMAA1
5LfggWrUtHxiHtsPcj7mCncvKDWCIMUCCCIbK/03perG6WQZ64wov53ONhSNKxsDcTHG8A6YjFS/
gD8UV+lce6MEKOV1I4mMDdVMYYztNS6aBWtjCwQ0INBpmCBxTti+62tR4r6vlbI8lY8qxNX4eq1L
MTgwrhxasd7A31x4Uw2EEhNWWQWuXrBOOmCplhhKlSLdxW0YDnWueQlwY5tnqZpaMb+3A4pROf++
8Y+Kd+LM07tzEcbObxOATSKygRbP/kJ9BJaDUHwrqpofsn3RU0Fe0kKrzcPM6AlekfMLfsYmMU/+
Ep9UaFAtNN+v2Sm8NXwVakG19cc/7Xk1qDkiEHrwqOp91ITtg0DPcBirzJ7qJavaR9o1uLHs04lv
IUDaSx8mmS6NkahgfBaeG2kJmAjcMSHJQyKZQI5r4LEg43KZzZXIKV1Y6o8k22A+CsCPyKBUygEX
P/JJchRrxuS40wfiANMs0NvUo1IjWzx33dpoyo/NRYFkJndxD8t99EM+VjT3tUgmXvCbAwnN6Vip
hPVRkW+PzSRupmOB96fRad+0AI6cwNDkYieQNESYQLu0OYxlH+igeUjwahMLhid8HOO2sJHraphB
+jfahRX2GZ5Al+aZ/B+hZeuMCeLWyYH/j3HtSbFvdU/OMZXt8M5b95W7q42z5BVUFpl03yw+MBQm
RDnHIQx9UjWvf9XA24vdl2kwatbqJt2ctNn5CnwoWYoZt3GzjKDejuJ/e+RCk+5oHrl8mjuZrt1g
L8YOBMGh5h4MSA18FSqq1+rEIUzicDxiHYQ517WCqyxYqG9hQFHt0NrhGj2PbSqiGJ48Y+df4KJ7
0wGlCSJ/NyKf1hPb2LPJq4z//+5nVFxL1I0MXohYIFC70XpRAgzX7gmgVc8X39fynjbAjKEcXtDk
gt+YME80fvqXOC3lKyatOJ6N/InJnDKybUYo8eYYN0VWmOt9e5pXpjet7JBTyh4npIqb4JxInBQq
PLDQg5IiotwFpQYn0x/JM3HWnSfwlvpfNysts1oIttQNwCdW2q777tp6wS9CxenHSgO+YTyWhKH+
otcM7DBf0bPeZPfn8Ts41p4wCWQ/LR9UQvLksBMNnRA/cLIZMqrr0u+H1rw+svyA2GLIuy9F70CP
v42QuEzoOKfE1ITRo3VSdrwrKo+hBZRFvvfidc/pi5uc9hnNJx/DQ7WEw3hpH05Q5QlEKgYwFu0M
hJ9EjT7jEeJ4ml8piPr1XlOM9ePsPjfJGAmoniBuoCsKS7Fmx/AESsIjHNFlQiZtjIzZE+1mm1mP
2gt40Et8YF01aRE/rD6E895EcGNOp8mWWlzc7jLLcgGWCfDmipshaxjimiIcpGc1qZ+cUXomb7NL
CWh9DCxkERpGP8GNPpefisyfbbdNsmH56tdAFjAIpbUh0j0HaBTglkFIE0T0eBBJ191vv8yKRFrm
kASiiz6zLwrzY2tjtAbuZAdSf/Gfm2DnUFDhAJ+rKLB7TfPqtNsVyQLsHcXgTK6p1FNkrWqaFcQm
Xl3eCSuK67cTm7mfnnS32XPgMBqvk1bf5pZGTVrQE8Ee7UBU6kkrNcjLgQQwlSZ/VPRUTpJpgNnS
SagEO/9wxsARB18CuuEy4dn2231FNzWzpj40Nmkoh1SfVT43CfPL9r+j29VRT2esiUjdLIO1G84Z
Qpid/TiX+4YZVnUoLKVifd3RgnAq2gDMuk1GMWDmcQz+T4qx+vHB4JwtsEOerpua6HvTOGKh3xSv
0DApCY5rkWNVg8gxJGWS8A8w9uaj4wdxx3Q+R8EJuRhZqWjg3S1wwSQu091qLWg7KOq4a6mFRWVq
WaviHMI+BX14c5TxgXGySnje6synbd8j3NKZlosROr/NLW4dCcuL1c/iZtPWpWvfE4ti8+QGouQz
jDMzWMiHLPJx423QjdhezK0LEI1PjpVddD2EYXEf7A/S50GIIG2FlJcxrz8qtoMixMEJ1j3HFTW8
oMbk/40PjB7QXm9TPJ6J/V2289sZXdErYuu3Ljv9Gejpahlw7kGJxX49ATlTRfwY1w8IMfHqVZFv
7LbRDuBEvlCO06ZLw/0pxphEpDQhMhwOLVfjxBgmFD7poQPzWI/nPs+51//ko4QBa/TFvEUTzkhh
AY037omzN1GYJxpqyCkBqf5i/NoyzdAUTFuRDSB/1vlAX8GVAdhawF0e8bm/aBZeyXhq3H/docri
1Wr4iz+QL+QtdMPT8YsoqJ7lDNDyOYn5J6Kn7mL9627iJ7dDpRKaZofnGW/af+a5MMkbz7SoD9cN
0DuKtnFWkn5Jk83feVcdvrtjp9c4TyXkGrvS0FI9CxpTB+cTeyjZGB4XhNn+9286UovmfkRlXqay
D/7guFE/Hf0khLmpPCHnnkh9gpU5BFDv91CTUXYzn7KzNqipF83odq48XHl/e7qPDcWHsnWG5z8z
Ry07RzsIBBWIgJChKyobcPOdSIfKS6ldgcvDhUis4KEypqp+nC7Rhj0XNWoOI8Go2aDQq5wdj9C5
xz24Llgzn59b2nWEDh7aUnfEL9HG4VVnQZJaAx2VAfUnIIZe3ZS8VKUJ9hQE/OskS+9A5Ogrk8Lh
wtdRKWPtQxL6S2KOHe4G2P0A4FCAbYzdf9nBaVRE3CpFcRaFNyiGF1BLPZrPqFEE9dgm8pRmVeUU
9N3obHwVM87DLS4wBP/ZTERNqau+cmtVqk4AMUUuzsGGJI9SlHh6lprXhkzI6yHZvip9bEh7DIOo
IWlNhtCiormzwjvNuayC95JxA1cdVP2qInegNXx2EG1c93DzcBMQFdvmpoh6BHA5zLsTwx06y6mf
TZdPkPjY8HEtBmeUeSrgcm8PQuJzw4Cga5pHYDtae84Vph1Yeehv4ryeh9q1b3k3F/4LY50gMN4o
0XrS2EeGLEs8TBdmruMRoG1OHfHp0NoW22ia/BHHYW62ovZPZdolM3pJMUgOcclkyRFWAuHRRTw3
4B6vZ9qjUnIiqYrMTrJ/Z/0bUlTMlofE8C/Yy3/QsIm4SgDt6MHpYzORC464yQOKnVicb8V9iY2x
s8dP4w2G/Z/mVeaqSBxBGsVQNE1mG6qrkS4bwdudtIk3uyatoH3STrXYBowLBGBtYDgQ6DnbzFax
M0Z7LUqS6RLzWXZdmEFy1jQIPBvFhk+BDzfa5+O2QebIH1CorVLyAPzfe31Hce5M5DIq+ndbk3ac
gHISCcWUpRSiJ2aeAiuH4H7n16Jo8lMvAnU1NXCKb994d0hEt/K6RSzhixX887/RKsG5IL8N/qFg
7okyCmTsFhuUIFAbu+jmTk+pGgFlQ74CRiQVQRG2Mx8TpI1xqeJ1JKlwCmBLbtEdZ4OE/0IQ5Yco
V2itaCnSwAWA1VMp5e2O+LYKw1njCctJm7eWhdkH0qhyYKImD6qKMIa99lo4j9ySlA5kuzeamma0
tSecVKBfsTR6T8vuW0x6m6lGO9QSP3npNGNnGQDKwb/XAl5j33fFvbRtV30Jpo9DF4oaI24za/c9
WcFhoD4nmMz5UDm5vL0jpuBNrvrmfZkOPvAerfH2UK94QXeP+ChvwPHekbKZVTwkY+bb9J7YK636
4rXmgKfR7f+sC8PlwrCWz3L2tB9Yon8Onca19cEL3DMD87bINKga82TnC9nJf04qFcdbN+LbGoRZ
GcQIoP81IXrDl2yfnZltSYPZgY8YBuZbvDJijCbkByrjLltYG7jsRdzWzZy6GRfFnQtebsYyvNvF
r2hpT63wfd8QtnMIS/lS+dWur+B7jMb2/L9PrsqsXLlUl1Sz6a8LS7nGrutKeZrdtF3G0WcbBifW
yYZeGweEKKHh+lFCWRkxRK7JCgLDURf7et3pkTu/gKIVJrj43MfzGuwYZeIzVCxUs+j1awzYio/p
LaEGgmfjK93T6qoI0FQnZdcoSGq2AZUTiE1ha1baafJy+ELv4A3zFa/r9q8sgMl2LZ2DoHn207Hk
rsSiT3gsz+HP3f/1BcmbroLRx3cNJsHmPwM0QDlpI/wRkl3zfmgPuV7leTK90KHpU4Ln7lSnMRfa
AfKkqLIpZdUiE0Mhd3bv7RrURM7EJpAe9j3pO29uIl6v6l7zjAHOWAgmLsP/HTEdsdzuauo4Z8Ll
x+YES/lWv0Am9dsQtXcjX9P259zgN/ni4V3Cp31ZFvr27y+U9cg8YNgt9naI73Nvsu+wlS+eGoMK
t2g6lQHJNqIe4mUTQK5cHx36IRxl2gj2t/IAx3g5apisL+1vQp9zMZxrsDmgWDkwSiet/n+ykpfz
4p2tx36N5d49y58T9eBlnr6CHsiwCk6GLDzB4IYoSgwQnQ0Rj/Y5+/93e9GknDfVyz1PIxVxrsnd
PbJ882ZfaVNTUi59irQS81CvijIIDKtUyIALbVVRQXN9vehQ+bFU2Sl0KjNc8cht0dWzHdjkgG4D
KyBMl4JF3QevB2uGIEWW3utBUp7VG9IKznKtIHwaoSF9IGZgB3tOUdM/x+lrNOSOEZF2YVyZKiRs
7MclcrRCXjl/yWjd2PedEqwl+VqAgx7jv+pA0JRtYpvVWRboKCyjRVsszFUmEqKJviACz6Dl+9sU
jfjwezrbeU3GC3xjpYZ45xGB390eiZxkbUB+VbSuJy4HbDgc/7SvUpEbmEDARwsI9Z+KCdnw2nBz
lwHXZd5BzkmPqvk4zCbV3KCTLIkRIsqWRgsLU0djcxe/tj9n6+nCnnReR32POwvjNnXddhcuuaam
zJk+ZXXIfEdZnHLLLaaoPVGJYvss3HSj9E2ykhIGtjHYxTEVgf9T40noh4O9cuN0QSkkTVtKStqn
wK2aRHqQIAHp7px2vzPlhjKdBROYR8TxwHxgA5uwxHHjDoCQkUGfDiLOn+YsxUGQ9bVBzygle8I7
tRtRTrtmjv7m9rg3Qsz/aejfs7H/VGd4/1ReuStJRklRAxp1ynqfV2cl3Sk+Y83rtyAAcT5kaL8q
/BJDD0l6CzbNKc7Ef3RIXGfa7vTehJWwBB7nrK1r4ylYiypibeQ1JVdGfxgfF1w9EK9KDXGCvZ6y
/7T12USGFccRsZvKKS4vv0ArSZD3NhZk0LC3Uv542v3RC8RUzdlEvL3joMiFZCJs4PTV2pM6xuUm
rkalcK8r6I2ZH10qFsZzS5aCxk1lM+loGoqiq3VTQsSFlAI0IW1tlDLItmUP/MVVYpEZ3BjLKfMF
p+yOjksJONHWgTKFpeXl2La9tJLdn8/kJsBaoDo3BZ5PGVg7UuTToANqjKuSS5IZXOYyloR/I3UX
Oqs1lpSHu0sFcbZq2AZK+NhkcVyR0UeQnmR53S98jFSsXvk6L5s8WGiRaDqmnU1wvG/4UfYTRR9y
0Jxg9gbIpMxAvdaylHhILgZI18iRAh6GwEpmNnX+TkakgQGWYX8Jm2dI3KyuQYbqtVjwYEm0i5G6
EaC23q3W7Tnu4i+Rfn+x0/1r/V0fyFJ58+j/XE5ve1rTJKWnx/VfWrfkJbeCUggUwsGPdXk4psrE
lRosFpflj/ufOWHQuyGJU67khgG2XN6TaTB/hSgBM+cWx/VVZNDBS0/YQc6Do+c9H5YCgSClfF33
t4L78aVNtBStGLqvqtu5SyG3HiGrVl3WFnjlBAErefE+eySLLuBEWG95Merzpt/s3Ih15hk8jCRu
ugDHu4D0aH6iSgH4ac6n0k6YQ7WaLIcRCmh7M2D7UDVsrMGO5AmKHgYlxc1TKiyowZZ7b4qT6PT6
PtLBp3DRAGDTs/e86YSqWs4IPDuSMmeq8xZH9sYW2C7GEUCgkeJyM1YnCTXgAfW/euwS/iaLaT9z
wdlnT3wIrBwcS0iWpIf/1FeNFw4tqmi+JczX2mq46Hjv4lxrH0ZkM1QCjM+kE5PubxIW5OLsNRyJ
VXHRR/1bMJnNXtr3SckS8sHF4lp65ePgev3NrfR49z4HH1VqHZWAtroYEigyAOL2qX7+VEZFSumY
eFvcWDBp60e5vYS5UHKiUBfvn+gNWunaAwMcy8cWZVsdreYToL57W+6MWGmO7wZ5R1vVG7s3Wcly
y+X2zEjBmKs6XhCTcz1pppEXTi4B6HnEoDin1BM1Fle3w0yawr05qHosBmNPbDlAulNoE+JaTa4A
8gA2EWzDDojentBKf9Wj2JD/eJIxQ4DSCHdagqGcGHpjprl97mux/wT6IPZ4peLjOjIyP5vndrKh
E8l/4MwLGM4+0YXSAT6jfw5edvQYHylcrjeuwTtmlsfCEG0BmLgcTjOKd1JVtgEBEs5IsuHMK9++
2jnIwFF+Td1EkxsTMjKqb2hkMlfcavWVYq/C5Uq545eqt9h2TL+sCUIQ5bjO/OT466B/N2t0izrv
EaCqyVho6foPpVPQ81KeYDvgk1U4v/Rv5SkdQcVry9H2hT6usWc832qzTP3VlSe9vXBA2u5MPyDt
spGSCqoRNtezwsUMFD+ukZm5HDW1QtRHX/kJwBIqK+/3c7VQbWLQfALzVlcpyUTaEQni+FMN6V1A
Nqt3CYVPeYD2QDFDisfF6Ug3K5GsqhnLXNg5HvmPcruEedJ7ZWCnDRaie3rBfrT0ccuDQeeAz2IX
O0XNrM9NOqWtHgyvsnQLWwt5rUG+R1bS98JXpbrSOI0QbQ44CSysqTSSzf+IjEgPO1vBrmaBoGL1
ScMn4JU923BWM5E5P/D6OWuwCGFiPQsgr+uEvEK196Nb+zr09nSB6HrQNbwwPmK9orq8cdoRVQyj
rRTF5Ylr9IWn8I+Y6NPAlT2C579iZjcRC5IRPQ9vyD3MZ9wcHh3RdBYhek2DW82MMCxbWHmz2lBD
iMuDUl+ICyu+nDKIUuS3Xh7pHMEZjmnDDOaUj+x00Frhv45bTaw4FiLRzgo3eYy/jOineuUVUJzd
kRYAT7kUEGZzwE5Br9AZJwjU4vqrH6gyJq4/G/E5Y5B8vqOjgGnj9o7vIIHcscx5bqrnfnMpBtG0
fE1UCpdAhCcrl60fBoXkRY2i8CWriA/tlVCWWYPkHkPHFnXvvR9rGCqzQ8NMIg1UULx9GcB1QvFc
RMIT9l+yvg6i2V3zuhbZYEq2fCR/dqwVCzUU/UYJb7RU6ZzBllfr8MwmXkpqwpgMT3Z6AuyMOnR8
G3ydztrFXlcK4wPSm9nf0TvsQZC4PjDMxdxw95q2QwcqDrRkjQT6DZGAC52IbzVq6+5DL+O7ODEK
Bl82st1bbDA5grCrMaxC1jDv4YVugdfenHIvcVcNhrtqQpsdDMU8XbVeFaTy/p8XRSDFuExIDp7S
LLwWtTsCaBT4QslheSFbuz38WliXczyQn+pBJxGikft2owCgIew48HGKiU9WO3O6TkvxZkX71HgV
LleKOAI9TbfHGw1TwKaLI5BWSBhkS+EjRdNTve7tY3SobDju75UrClJmPE1jvgV+/EPx4UokL8g8
Q34+LZN0wOKZtcsQW3Y35puUHdAqtYo7bynkMAACZ5um6qlMv7MTIRrknyY71h2xBfZMxFgWUX8U
b61Xi8kvRZ5fNC1ngbe8LgS/o7kwaDFpDm0D2q6Qu0Qe8BVxzTt1OeTDX9OPqxRMUZ8i1PqImf95
zFJx5wb4cxRG/zPMwVGH52UMQkLj3rm8JRRog3D/HysKNX6L0+w4QzyVm4Prjvwx0zlG7fmzOntK
XBOXJpUoH0dO2LIgCokC506hvaeE+oRY1JwZ90QMbGy98ImsYR1XvRZwd85RLSstvw9sN5LKzPff
M4NJC7IYgzDgLZmPTKWQi4518Oa2iSbyF86KyjKKnPnwclhpP/WQ+A5PBkW+9z0zWB2NIUrQMZcL
OCGcq0rN7PU6Hoi3ynQ3fBVLbz7MeEAMOgTuZSBp7qTZ5mAlubEM01qeIY26kyRAaEs5Zt80in8I
5jpbTaV6g6DW3I7HjTNDfoq6oCm9AkL+7Qh5+evQxi6ENRy+kllJ37HqFr3pfjrgX351cFLEfyEJ
dUfmgxU6NS3BZzZXsH0e8ptWQXVqfllV60y3Ls0nXcjgMiOJZCobwNkcE+3t94uksAbPe0jpKSAQ
M3WayqYHxpNgQdz6qSqAiPa7rH5tc97s/cm0kipAUgP2v6aFyhcieA/Y4I3IZGg6lqBaKo9nP1A1
dx8LMe5KGtqfqDQ3WDfZP8otVqwXD1i/zKLS4AhAJ6Pt5ClXf07osldFmXr4HzpbDyWTywsuR3dx
zLxo8sSL5yZZVSd3hLCagO8OrVKJycwUB++40Sreskq5ItLGIGR1l6uN/yD9k0YElwMhfJU4Tal3
Viw2WXJ1Mj6KwCZ9GxmdK/tofJu/X5v4gJVTkTca/A51efrytTPmWyV25FwjWseT1B53zSlRp+c5
PKnIoTBw3hVd7YnxXuQrraK3nf46HyXFgS8F1lIHb3U+lR6AzSw31pLq7hjsPQPTuLfzripDhMsz
PhSz1yXJULTTKN2Th7Oa7oCq031CFDivdyzfYg7t0KtFrK5l+DmvEDzhevjX5DGWPm+MPUQ0Lx9M
azSHrthA+tl6d2Er+Esi8oRvXLE9wS6SNCcoLNP3HNiAk9c+TUzKkhiMiapP4RUyI7QUgXiPOWXg
FJYBZ/NcDGPgmR7Hbz9R6/lD0p61w6dEdbiAerD2ZBYFwF0af/mwcGOvw4Aax10q6cUCz0sc9WqA
+Nusyw3Ok7OsYhRJUVg8gc+uSg42Q9+LftNL38MlQEC6S32nbQQ19a5qfo8FeNo5pXMyArJN+xEB
waRmdaYrL4+nF6Bry4hDTxeJPHqLTT55kUBLm9at42k0Z+ljAGFNMW3ayM+1Xum44/GPHaPINygT
i/Zzf7AZXDY+XMS5e7X1bVtYQYBEQT+3Y5gFJcgTWfVa+YSqgBC9Ei+ervLoqFgMDwRLT5/6XmRb
OWFNVH5euHyM5g1tMpV8VjHW5l5nr6KmYHOfyYaWkn/xY5tOhEco5Lum6eZ55wFYXfZ+GWDuH9oK
aWzbBgDtjc9gHsab1UJyoe3cpslAz1O64hVzuiV5DQ6t7aAMx0+L/8gwbgFSnEgTSHkXQ8jIX8QU
yxiNDNGU7LqZIx/xv8IEJECXWSKyvQ9DDHWlJuEp2gbhfQUfUxKIGn/+/1PrAl89yogG78wH3feR
UwNRh7E/EqbS+hXeGDDJZB0G6CCesytaKiNceFR8N0MO4ANwk5PDgooHYwMY4vOdO4yFdhWeYw8Q
0ld54vcM7Xnyy6nsh/JNT1z1NoWFwaX7dwmk9KKFM93Nanz13WUnCA5D4jbRK4X1dJSdxTcx4Yet
4H1s40owlRwXttVyhW8zFKWcXPJFeV6xa0wM6nWV6+TwzeY3GmLaGanF9mmG2ZBfu+d4sskOAwNe
81l2+J2K0nfn5rVaj+Y6G5Oq1bMaV3P8Jv3kXkx+/sQt7IkZdY9ZvSDG8cWTCwPxcj9NFwM2pWHQ
3wKortPY5wstbSeVDGInRq78uEzRs33ojfAT26bWcJf7ieaD/BFNXwfrdD9dmLPRmxjfgKt+aav5
YSThlsDfrmLIOqatxuaoxmHcqvFBFNh3grDvZ+mGqQC13qjx2Ye0/yuUkYIxqOo7Jko8uP6gZwx6
FAIIemfaN94F+WfUpSvNmMpOIdCMMHFKA0S1baND0b1FDCxkNx1g175Fc36CBdS5YxGnSMUW1DDO
GFh2ulSmGw3+DNX95bYUVcxUUuLJ/TZwGlB13EyydPEBc+fa+JX4/GH/Z61hCAygdP73GWcpH53g
goY+f55y56wlsturHgd4JMZVNP9bE3Yq+lwirQqGT6SGK+KgDgYyzCtDxgk9m3iKpb2HbnXY0odM
JXDFbZnejjBWHfOI8gelcQvBzlc5evrNVWNhF0oNUmHfolGeR+iwSRvIJZ+sAeXqf1YVPls+IpPk
pk74QGt7xmEt+izyezh4sBiY0Di0LxujzlGw/CDEKRLLunYOIZpVtIAuZ+wbH3KEXJh0c8uaS0wD
EyqXpn2/rZLmEapbfPYpSy86gXAy31DJRAiiSvW9urYQZGrPiGRD27ahEahSt7+amECYS5+UnNII
dkHBc27h8Ih/xJ0SaviQenbPOwvIbPTmtcvk7KodrdwSqGaZ+tM0RW1DxrbU0/nzGurqPr7UQ0+L
O1XVoQ//eZCl9Rsg6/SGyIF/xK04cm3WMjED2jpoICi8mRgbpDRdLrQho8aD9BLBgTQFrwJxej29
fMZjHVmg7sBZKzEoASFakAurfdCV2XqUNBmeJFsTMirtXlRaHzmPa3cffPN7BYoElhY5evRP+UFL
veUl+jI0EJ6wlnTxuwpwacHAmf6v6LdnpqWlYMptuva+AY37xmt66L0IhNd5ZzHutZZuyp4ncRJ4
ONteLUSLi20wmn4yMlzRc7/42dJRZDOowS8yU8IYFKt4ihxRyHqcee6eMsqHPZ0kJEw8KtJZoSW2
6BrLh5ozvhUyPN7glMVYPb+zyLsv7d2o5jtz+BcSb2CwCPWCKdOgFfWZ/CdsK8S+yyqD5+9ZbdaB
HsswVFbsWqlAgdWqWaCUbeFoWKD8nnJtlfrG3t35nUC6sIyHLSXdU7gHPcRDtNeNgFYtqhTAkxn9
tIzwwwYoW57eWOm/okvsnQ3GET+nJuClvU/vODhmo5PJpPVmYTkPa6qhg0wWA2RIvRvKrGjDzH6Y
ITwNpsAmSiHv1X8b4YFMxXsiBEECbp8ZakHhhackWBCsj/HxcAr+OOthJ2I/l6K0l+JK3Fk2KXIw
iEUN8zy2w8o5J1yGBYn/PTqPOJ0jeELVuIJHSbdFJOeftu3b+LY74Q6QajUBeJytrdauhK43ZH4S
qF4WrRgkyiY2KIjp0RvlUcCVhvCcoUTsNEWEim2C5cCm0F2onOiHppq0U8iSwoZ/Zwio2eAZAZ5k
a5oeogXoKYHn0Tnk1PDobGYHyrIUxhlwdUVMiqBsQ9VdFwnpOBEgM0/vwkm57nHdxT+c1pKeFfdI
wx848Oa3SwI/UDi/9JFrfc8nmfIlbr7/JDWS6xNkzgdl9jEa8c5bBrJHCRy6Tj/cAbsJfpyplOy8
BUvgNBC8NX2fC9LiGoxb5fMp7huBIHubXw3gX9JKhkAWydhF3XIiZApwfzZpr85cBFiZE0O1je19
VA9qXooz2PkXok9tZcW6u70Ew7aS9FAf65TVmui/FMKyk4sTz9eu8zbzQmMK2WWHyQIG9IaX60Tt
tSO9bvp2HnV/BRuQCoa9dex80/g4y5RIhnC9zaAlw8RTPAx76anliaGukMy8lRTZVAZNAFoUxY06
xJ1A82BTkjzaJE2D/qKU/EDwHz1hPQNRTnAoeZhRmOML0gA1rLTmQq+PxcWUzlTSmBaRmMr62s4Y
hR14fsc5muiNli/KRVjrPhsca77ubsqw7OlXpi+x7l5z3QhVI1EIo1+zOjYVW7uB2XlYevIu
`protect end_protected
