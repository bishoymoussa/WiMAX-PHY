-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
U5ImhBvsFQ6Qj8iUhD2Kx8vmAZs1lE2zSI0nX7IRT8WqYaBAPk+zdWwbGjR0fFufu4qBxgp4ldKR
TpjCe2eX4B1XpRj5b4A8ZBQdndZoDx9G0VyE4N+5rStaTYijD6y+s+uEW8QBT6YHrzttFBm1h70C
NzK/1MVKc9kDjgGbajpaUIAH/S6ccs5Wzu3CibC3sRZGTfr3LuGW7z+HRczRqdanaLxDtC88YhVh
hq4pcSIZT0s1UoufqQ90CJP8CtomruwfvZyGkWTfe3Lj9+Kf29iCJE+Eg17O5KheEeySgu2MuyHh
3pYD2xYBkmKDOmui0flWao3Hdxmjt8W13ZC6WA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5824)
`protect data_block
WmfpC5BL240i2I3DwyC233sATvafPNLWqdiH49MkrZq+W97VeEuVOVRP8BZ6zyGcEneck3nPdJY8
xpgASm0GoNx4nIpHCL0xt2d+TRNYNUvGMStCSR0e611BIdw0OyCPqzCwoOUebS51ecDv9I5/2Vlu
gipcP++iCt8LV7boKr5m9qA5z05JjGQzJgxBT+OYpjjbBrt8M2qeF1kNjBH6I2FzPqUMMXlfoy0f
IHzf693i8Yomw6JcqNrSA+jWAmVRtjaLELzoAlwmlYQkEJuQYXl+yeVxYwOORgaMYUpxJMnXt+ze
RAOT7OX5M/aIlg2kgSOB0gxFaCJqxmAgBh5zh/kbm606U77jS8Q+G9AextZslyP7wlT8+YTYubIl
0QlbivmntYJ92l4ejjxLL5irHmiZzsCAuQkz1gqjVhJH+eIEZtroU0YIjzkFgPotcXVcBFUF32m+
vnqkCHK5zzqwhk3J/qf+7VghebRs9NuF4rLb9lAsB6pKWwgaIwMqn6npkdRZt/hNK2UxVkaguRgo
E0cd546/doWhv49PfwGQzdWRbJo+5hxzhedofxPbFdjFpnnfj5vIoFpgghTTmsqD5+rw5bkPCRLD
L+2+RR7/ftTMFiE0n3TrVAFAAkqJQuqhAzezPwtPBgmurlmC+gKkVJh6ROrwpyWQ0+xPVpbQAl3Z
gGN0PiosjjmJ0jOGHmQhuDMTeVypxv4NJej29xUo3D/d5wJQKEA0BpySTh3sF4ipSguoQtr1D/Sk
i0NnVnjS37pyeVb8WgJh1CTHh3whNIAoEKrwo7kR4/nYDZWMqIrbrYUwEKAraU0RyW9gkYDTZT5S
Ju3tJi4sWW3QCAeShnq4SYANMyfjvhjlwWFtg5PCm4+8xk4ieT088cItRe2vxkNxG4JKq9fHt5TS
ckkAlLAXdzZj0iPAOjyzM45IWRtkVuvTIbHdCraNygPPMdP3ibBErI/Q8aPK9sMmln10f8azo+Xx
XzJIiCrEapELx39O0muS8J4WnuMsEU7DRw/Kez0uClInjqOuMPhCO/8OF4UD6fwwezX5/w5/Wunb
mKnJSbU8Okx9qGNxZ/hTBI1MkaWAsPHWdt8K+ZywGxR+fcTL4PdJJKDCQgYynhJENrQLEU+eCGtc
XPp1s+81OPqCxwv+nZA1k/7Tck77mM1kgY0Lb9UXqAyRlr96Pxq1kkcwspw7TVy+pfJZfBW4AJ50
URsDmQ2lXoDsPv0k1hRKKJDpHEsZyywfC26W9OV6BjU6HR6Cw6PMuqCBNvhzWl3iWyXEWa2Mhmxt
RP1+q4NaVv2392IKNZ91j9VWuFrtnhkVOAHz429hJJvsdvlTZyuLefJdoj5qmYFWYyWTgq6iz8GZ
INXxj1EUteVsAqi1GfYsESY1AiHM3Utr6x1vnJb2Cj3cMZlA9qbj6LSgN4xrjvMOgp8ssDlbhP8h
2+st3qtCAGHtYXb4x6nxUzBfbgCXLFM6Ac1rkfV3nAgfsBp1faA1LQsrUhsYHiFASIXJkfGXW9Zu
n1Llru2PxWbeDFS3GW/NKbijzT54c+ZhoPJYKU0adUGFaEirLSeS/eVbPJW3n+3zuSDE9A4o7PRI
/FwqHNk7jzoS7FgKMNInf3WY1uj4OTuWckdYCzsk3iQ+/mY9CqPSOxanOHpgknrNkX6KsdSBBGhK
f5YAkBCs334KTxDabTuu+NWDTesVL0skaxLUGkrzlPW7CLUeFXfY80RQR4PU+gWSNDYZvhQ5x550
VV5aP71JG6DZ3Yk3/ka7GJ4Y4WlkCGqTVsbFfBWQ4OKlXsdTC0+/oN57JTHHi6/mOE6qwFiRWHas
w+rdAF9z6Guc5oPgo4DP/dVJQzDKWf9AJ4Xfd0ZJ9Zzvr98FsUQfjMiM2dSLFDr9ZV5OHWQgNiAY
8YwjrMk/wgemH2O4CIVsr/vySeXL27gD15LLSS0ESdtdapTo0DRSDthgUmz6k0GFjYojXH2EHdP1
OwZMW0e+ORG3cqirlvkDwi6UBIxcFVI68udOndixmFBGkXkNBWAu5d3FAq/4ozRM6ABmD106adb4
MPwI/G7JoN7AGLtrsbvUjgb/rhpr4JCJ9hwnzMpPKMx4mIbhr9vKxxUXGW4yp1WP9z+GjaQO7HK0
+z1YqXEhvJc9S/nPjIW54DCu84LE59VbQAcapmiP+Cqp+Pn3aXtTyMbboAhH+zrxnX94ry540dM2
iQ48TqdXZBglUGfSS08VthtCteEck1DjlSFgccjTxC8Fot7LWtBA8T7c/RGZVR9nmmgZ0wdpa1Aa
GnBHlDwvr5hvfUjlfC6GT1TWcNFwj/jJSa2W6H1b+WbGfePXa/xAXo4HNlL/Q3hhvYytVOxVEx3I
yq91hK/ig+q7JLuI2nAKRqGWYQbqZytSE4o+lcGmKuig2kAPlWMmmQ96D9W/f/tyWneLKirly4Yc
TmbqjB25A4G1Jp5feRqgSksw77G4rXOf/V+ORE87/NxeirfR0PCe3ng3qTfd+aduzyi/cp8Fnovk
fdEu7zxBSR+R4ehkbAjsOOmvsOUVOZwztDuYwPIdwz+eIxTb8J+gncCiiOv4AL8jBTvriToTNO8i
VPn1WEuPkTrG636M0bdpyk8p9nme+K3VqcTZPvUjEBiWVFawOBLpdkFD9/W8nAijjAuaOJiI6yhZ
tE7DnqAXjM4BtE8PAZUFDapzj5ncJ1GcHkAx+1MdbXidS/Jfwm/lPUMxGj/flESYzDBxat6l/3Ag
CpjFNlowQjX9EVdrPcP2DLflNPlBsb4Im/qGTE1eZz6oDcv/l3Mc2bMG7l5JbvvKFUzociA0Ooh5
ny9x/AVwP+xxOOq7SCnMRKkgES6Vn6AA5RNrjAp204W4R1sHQXRnEBVgpDEPMaPQMZYJcTyHokTs
SHPYqh0MfF9wIS5X9LPnoqaLUBBB9L9W8R3jZ8prgsi311LYOGtns61NJOZUuD3sjSPP/BlDlmwr
ULWcdJgWJCmh2wIxXNCvqypbDhjEzyJUy+yB4W1W2gsX/xuuY69Z1VOlJEK6P2jkW/bgdQYRuhBz
qszFhUzbshU5Pju/8S6Mj3Y/rLIzHEVGp0+Gra0SCHdTz+xGr2s6MOcxy2GYLCdMXCpZgXZU20cZ
F97FhRszzdRKzlADFB9ZgwE17BzsmZ57xefBgu8JUzNIsQgfePR6bgsdyNPCzoiDsKhTVqWCXs+i
KWqBBgypApR3xxmpD2WfOPaGy5DUK11fe1FTT1iUKRP1ogCUAiMp2N1Ur5wgLezcoBq+8dZ31Utx
cITVIxwgtvFmSqBuIHYjV9bUnoFj813W6Dxrl6dP2iUZ0OLnR0JtG/BkxYmH+kvVig7wc7N+c4dH
TZtQw57zNncxZhUL2nGSFWwVf9ORRd9wA+5ZV+80YjPsoPfeUfikUDOrWGjnknAcxrnUtV8TuGkf
ZZS4g5IXfyNp9+NSTnrWfKxTr3ub75LMgpGqAZtIciieEPwdl0lnKhC3gjWmZyny7im4BL5Cz7BB
iAAdefHFnNN2xU3Y0iNBXmAneeL35CV2xTn4AOxJPhk3Ld8llrPNm2htWQFZa9TzHLPyxa6PhM+P
UWM3BnMzuzGUkaN3twnJhX0C/I9430b4dupTbMhMAB1Hm/N0hn/y25oF/4odvuctZJNDcjvUJO/b
VJ4e4DrNP2Xz8UztulC1wAI2infUSGOpWr5aM17lr6AHFZFHeYulKhKE5I3IduCyuYcWipoIqWzb
OgQbEKT2rzYwjoqx0J5/t26Vpbdd2CuGb7yCi3jfWo8fpNJxbWRfEqmqf0Gl4Fg8BJKupWRdTPll
ZvYDb4QjCtBQYmQ+Cuooq3YEYi5ugASKIDEOwksX7TXhdPfseM/bJAnLMijbBfNtKuJ5P9WUhonI
qyfHHoWiSEa5y+H153V7tW7vHK6jo5rmKcADKhvhkn7Xj2I92HRZc1k4F/y9kKEdmNNWp89OwRit
RA5JTUuyYTR7aZSPp3caGnNvNaKGOHjnUxWhVWAaAYbOMzTQFpBRRDXdZpTl5DF7oRp4/K/paCTI
MharQ5GtWxh9u+sSGcCeAekW1WE8PyFR6wYKWt64zxfpH7wa1eATTrLYAwLVlxilvDi2aOASg1JO
u2G0xXBv+QJUGzQoPxuX5fN8YEFPynqZKCvMRtALTCwRfLcc4baZds/mK8YNQlzMe1H1rbBgRyBR
j+Ge3IXNYsM0JFZcGrb24IFAAMo6eGUy7IFzo8NGacV4C6uSngszQxLvre5aLlaoxORCkOo5kPam
M1q3OjO5vxRve+98QyZlLhQC+BJuFANwNPJmrogVS5a7sRCW9+DxHlT10R296QWaRtFK4asthQQ2
dFtvT89P3YUh2ILYIT6jhHFvOdFW/sbhOFyRQRifBL3eG5KxF2U1zAF0JEoac7haVuyumTXoC8aO
hB+zALl29KdON7FnJs726IPc66tYAUR5I5KDN0B/a2A3r5pU1m+ReKXo0e22cocCJsyKe6L5IMrN
V1iJCkTjWtStpyFu1AXXJcaNjBjplZTdHJimRT9cOygppTYCeCS1/NJeGm0p5+YbODMRWxwUgMaf
gL+nhh72iVqLZmF4Xg7yAws6V3fHXTU0TQSahGzztXhcQOGOC089CIpT2LIpTJixMurzqQoMNXHx
npGIetyfL73CHIBWPk7SPdniuURtsPSUVbo/mM110xUG91NsdDP9FLVJDVILa8iTkVRoEm87pfDx
segUahK2Go+w/JEtgLTd/2ZkgGEzHmazq7IpSUGjUdnkjW7O4oiHtPcmlj98vTC517KVYqyJaqOQ
vBbrvGPeu81JAPeGobIv8WFDSOarWihs2cJH3Q61I9U6mm+tcvg3+fnNLmI2YmCEQLXF2VXgSsDd
XPmpTY5ERjdDbMtuLd0/IVFM3JSLrKQGNLYwMhH2LNnaqDpIVWx+reSwRRWISTD4eTKNspIt1rj9
gxvo1CiiTgC17dIW6wtkOHgfZMyyLMtjsfZbDyy7cAa6et9Maxfh2YMY/nwiYWYGOL9fIUD8CSny
VpPxwHno7Fc/OWD9u/xpws8+UTOxwfwdMgD1mkn7M9DQantwTXUlwBa5iX+QKA817XnCXTLsVGtx
bLcLaX+/SUDYbjuG5NnhiFcg1u9syqv8F8k6xLiL8klinWt0nW/UYA/iBvXU1k50VeCzvuWvE/gO
OsWPKWo5jZACL1qcdIpcW3sRE+rF2I25Dfo/UxRSlN88ziHIM/jYcPOwfs1oQYypQf/q4gDonVSI
lvlB5/X19IaFjZeNAAXrfAIz188xJ9onYxNDI7RihCzJci0vcfi5bmXp+Vh0eLhocKBQ15at75H2
csrvJKvjFOhv+ouVj92kUK3iZoixdcK4xr+/Xu/Cj4+nVzgDPLmuouyeDUfLOhlUhjzmo10aCJCJ
VfsuRJCoRQTLxHiQA3WwGXIxdq9jq49QbMMQPJknvOPM7Nxkbz10nKUfi/aQ7muVDctDOGfXHBt5
9nzvJx6VApEOj1THSDOMnsFwUs0XXJjDNuClklz8CUvkvMyrOBMyAE2HpPY2bTCjoGHgqVXTp4HB
4ZWJDHAZNWd1wzrYualsgfs08SUiy/Drgoym2deAe4Ny6wYkeDImzSMK9Zl6y0SmJ0dJ5ea7fq0d
s/OI8Uuo9LN+bQjzYZ83g+AfLXZpHvZjX7l6hme89yfx3HRN2BsdzDNXuZHJ7mUtTLanOZY9rfWF
v+DqLQtuMuiZYmEW51puIcNaecWUu0Z8srCuuVpV9j2HBRkM7j9Bb2kpU8V8nO+oY1rYVJsThayH
EVag/Lbf4vCOvVOkgZrRYOw+hGcwPJ3CMxpfaDfjXPQYYgybYA0yVj7ck14DOyDIJIlOGsxFqEV1
GP9O8E11bKM9zOx80jj8CRgIxTQCsyAmaLnt0vdUWHRfr1kC+j9X8roCxTiDGL2cjwUSCM4ZOYCz
ucRxx5xzWCtHYAVPjG4VXAsyyUoERjEYkdH6fh6mx4V18tdWVv86lZUbN0TNn8f2bmnmNaG7nsEt
zD0+suOvkBeaybA9nh3QecqytheUYoFce1Lk/h+765OgAxBHB1vphSw6Tuj2ZKfN7M9EaMuE9eYh
JWS38IxEns1JI7Sag8lnBoqSqW05Gx++pKGTWv6wHqu5e3xbBOtIxOI4eFn2NEY+scqvGdQuW4Wg
67s9sqnuwsoJjjm8wX+iPOrtzkq5QOBWuVHZM/BAS8B/6vtm+oGGBVE2ndfNSPgZ3OSWByQyCYLu
0HRqGtQ4CIUJnxT7eKWlZrAKgQkzn0V1S3tFYQhYG3m6SIVIe+a9nBTSrn7I2ivz86xeTUme8Owy
qIUc1MfOkQCOsn5m/Iiog3zAFALZu6KDbIjH5+UobA4tF2Bf3PXQOFMAQCltK2YEnWFqaWBu2+Jn
+jxKdz1VUyyHjd2AehViZXfqvZCljY39PChr6EFSKWh1vvo6K/dw/V57L4lUK2nC04m9e83Ygd9w
UtMLHE/0w9J8gxJvKcRP187WPDMcoIF/MeO2vPS+w5zL+g3dlOQ9P7xKv8mWR1PAGy7CwIcm7zqi
WKwFfA5rHTARBvarf1kXwcja9p4M8c0NnVJjGkK4zDaLzetJ4EO1SXAi7nKl95vE13W3lvsB7Qbh
BszyKhDlx7y7DcgXI8T74UOP7b+lh/giVyvq0QuvdOEhkHOKm2WobIwe9XAtcHJMvNAInuEr7Nt1
V+KvWX5WJWPXej5fMhozy2oE4SkXJFu6wGr3NdKwgeE+lRvY23Q47shKH7L60CkhZPiMhC8qgWl+
mRgNKKmMAo9ZMRfFHNMdJ7Mq8lxiSBsU+yMHntHIOcQDxsenMBUHC7GQMhGWi9DNRzZkCOD2+g+J
Vgv4m/zzDrdE26RMRSK6kFVNwPGfyj6uQvkiHcLuMbY2qHzmXaN0/gF0FgLsGBUt8+6464/vb/OI
sdxe0A6OyQAqD9JhtDPiFqapnceg5Xx/Y4wK8kLYGKaOgPr/QIoV/VQYBW7aH2QPAG0FrsGOq3EA
WvsT/1HhZTCl4zYr7p2isvdwR5iTq9UuSj8yBi+FZAAGh+Xgp4H8TG3nEHi3KT4PC51vZF+EK8UK
ngvBG4oMQp5P4owaxhSeg+o1dS1j0W/NFh+swkSpXsOJj61/ckmuiSah4f8CoQ5rJFhsqxFcyEeu
H+XaM721ZDpMpo5K9uak+WvaGA9GQFJZHCNfRB3UyrgRb9uJ6I/8WixFrgYrcpQrSxzbuKK+yBAc
vTt1PvRb6bnEiTGnj11X3D1QkD0i1uOSz9vDCTuQSO1QLIqUFSQUX4NPmu/x/EEa5RMAhcxFus7b
pQt9Ot6ONvZmkMmerxWoQaAvPf/G4VY7iRu9bAzrfttTB3i6W1vgnGw78PuUKpuy2q/vD1+MIy/Q
S/O6i58FADXDWyWuk+avhtqHleaunZyg0JEs7oH/WsGJLZuSENk2RrFakmIRBQmRzoLGH78bap63
U69UVi600D4e4TN3BFrzbpgHHQ7okVpHvrFfA2EL31LeHZwc768UFJpfPb521X/69OQaXPY4wjsA
upS0YqLT3mesBhSMo4xpU2UPxk4JourT9VRTU03xw48ucyV2FS2+lMyXJWCmRxcG+sh6homXnEjQ
7ydcf1N5721usuJZgJ5Nq7smqZ6ZEpBwhyoDNC2IEyGTf2wiYY2nqxyaMzo9AfTlsSdYUvlb3GrJ
N3CFAbasL6C1S5phBvSl8gsSntxzHHvhe6glca47XoBUH9Kwt2hWuN2xhSRMNFcfuukd/aLnQjyx
XVJmfXPOybpMwQ==
`protect end_protected
