-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
S0eqrapkOkMAfa4r5XtQao2HL9U3tsws0oYAI4GcZjrdaO2AUW8y67SYQ2f8s+jFJy/bDWNmLL6E
5WH3df4NJ3RhV6iFcx6vhIV1gTuRre2pqH4mJdNSsDgO5eeADCa0xcwaUuo/lpBWFLwcctPmcMCY
F3CmVv7FTcPnLNOIUlHYfh2CJFpsY39gz5JIoiXPIq3mn0WMepcBhCwSrZxWT2JR5eztNB7Ichl2
wwHWXrogYIfQPQKs07waC5vr7lmNb/LIZoTrfCUPaWeH33Yaq3gUDmEYu82KEj7LFJwIPspIrjrz
ftnVBBSVF6ZgnwYHsdaQDFBdI4n/E8oochG1Ug==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 7936)
`protect data_block
7l/eS+wCu4Ha9zUhjo2o826Yb4pkHjFt2K44tLq+JIx9TcSLZTQSoW4OjzuQsoBvXt8ffFp0AA3x
9JZ6wkbcOSZx9Tw7osBoDMpoY1rGTbnSAcKjPuQsc7M0ewM4Pi0K6Pz7SFijPSgLenfJDfp7U/3F
qYKxg53d2hRLTI96i7InJ+QDXeftefCFdtutsGH9rxM5qrKyEaLzIpi1dL0wLFgIvHPPDI997aGH
WN3T3IrZ0WuoUcGRhTLInKJnvsDiVFENTpetGiiQiz/VwBHFwmHPkk8Fa9FsGzat8IvWQg9BGvll
ep7RO0Ms/0PI3/mjfeN8f2oGM6yPkIiih/C1504+59rO3f+0slDGVBff+X4wHSOU6F3HGeRAv8zH
+Gy78jOr0TD7UjKgEDc48D0obX9XGxBSXakBSfjovR12SWzjRsXic8O33Kp2RuchQK/UVEaoe1gj
WjyRL3dtjTMEeyGpKUwjRrnzm0rp0tMgdafLqHklDsjxHevDqg/UUSW6aCkYtqinaKl1NGqYHa9+
ftDP3oIzjTC/TyBaKZN4inlP3ZDntM7tNp/j0QclqR0gRSKXwwceUy4rDkesTJXPMDjmgqGXoa9/
u2Z+AUmcxM4HhQrBBKjuTJI+5SK7IHtSUk88QXsKJ4QfAg/9NQeptsLVV71+6ACtfTwbSJPN/GdW
eeuLiCmEa+H3HJFzC7heVpiipUsiW5Ah23LwVXa0klSVjF44oQwJ+wRGLidbNqiE9cr4gTjl4e2B
OJKGPx9PgUF8W8MjK+3MPVGhxKaCZbrw/HRCDtFROHUaPv8mVAie3v6uUqyzHhHLqeuMx8Qi0QPn
tSiSreZImjyImWLeXmwDiW6Cy1qhhv5Xuw6J1xnAJp3kOmSHcZVobwCfjA06fKOSitnCXHfEw8jh
Yhv3Z/scA9/Jnkka8eBOrH17SJ0zeC0U546VGR6MX8nWIW81K1eHBVqZHX9Uzj4qW7FOkZfn6ad8
or3ZHZ0dKDWQzNNgkl9AiWy1R7pMa4jNC40vXxdJT9K14FaFWThGmOP7rmIdxH5vVw16J4Yz3258
4Z7DhZ968NXDC6Vpdy/yMAkpa+S0kiJjP62+XU/4CUNDNtdic4hxXd/5yLqqhleaGAtO+MsiKA83
iyyQT/JUKr2P/qjDHBE6CnMgd2MF2sYsyhQQhcOtG09UOnA2h44DSlyLSnNobsGO9kFdLOxiP7ac
fAVjcf0751Q5vKadbThZnxn5JDWEhHCVJD6dt+RyimOpxUgOLN2GdxWMWbMqJc9pkGZWDjsNYzOs
R8Jw+NF14tBG2cfJoRxM5L72EPS+CtxfMyCsNE15MIaK7F54lxRZDfbiDw9EbMOz7ClCtKi6r2PK
RfWLamA+n/I+Kd6hfMlIdPsX2ybAmLpKDz/admLAaivtJ7pWkR5EGr+jxnHx2iMZDccrpdaVa6X6
EPffONqImU8jmgM22LnaagfppJlqp5HQdE1LCCiw+Bt6Ssm8XMeHSbfPLQQgB1ODDYzawUYahAmi
tiqIZuU7PXd3RLvrXNWWxlkZ8NvDfmFP6lyiF8kMCA4usJH/YB4A5mnWshUdVkTrpzqOckdAv+9r
EK4ORs0YwdohbYFgykZEEWiuf0mJXaS+j8TW+cs1HoDBTEHbzqzDvE585vPfDux7zxylAh6OpPTT
5AER9MoqERrvr0EzU7E2kTwhC0pO8ukUbA4gzJn6JKfs8WEbnKvXc/9V/99JYfaRrOHRE/9t6sW0
RPvAHTRqAHQ0dYvxhxqF/fzHjnkLML5bEeX2JpV62St+JHUlWQo70gFtXA7yjsRjfuahfYu27LPI
ATllP7pUqbKGf7exR08/0PqrvJQV31GeCgyN6ZeoAti5r46aYT6a4OghfxNELkIbWyFeEpGlbxDW
h2axM9lAiAO0NxSEjNdZc+k+qaWaiZPh8uiR2oED7zQ/383dXBs9cO3+vK1jUaHuhuYWi/f0iF61
spAsNwupohH/fWKfgOkSxC0r4ptJjWCsLgO+b6oEa77g6fW784BBxQS/vBEMGNubFfpsBoqRTf8n
ZoJ6tr2nL8kUhaKOjwkT1yAKE2BLxvx9505DgV8WjEhtO77DDlIkHkWqslXg+coLuJWyrLCqMV2x
rLi74oz4hstHkGmjiusIVh6Yplym6Tfz3roJs7rIRljKjII4WVgZX9rWsf/ziwJEVszGD0a+pjTb
H5/w/xZFjt1sXqW0fpOzzBNfWDtOKMxzjtUYtMYDeLUIO3GT2cqJhwy+rRe3a1VzK9PgcqysvvYP
U0uORyrppMYlB3x56vOyKybXf9nFGaV4IdSKqQ3W00AhQ5K8SItz8V3dPmgFj0Bp/asMDcJKfxaF
ENekH17YbyT0Mg/gWQ38tp5TDkzmUVp53Fpx02yhj3QS2AKZ1Ctiy83joWNQZexQuJt0kKmF5Q6a
84lSM0r6XNWK7eIe/P1kuwLZTHn63g0xtKtxmZxWZyKrwb96e3IfNc8XBUf1DGJUouSvtYc/AZZL
Dmm/u0brNW8boJHGd+gyu8KD/wC214LmTXceXb1zFnkiy31mAmS4foNQUjiIXUvu/nSnulWGdJDY
ff1S8ED8EPd4xTNqZVM6asGRfjlEOQQlXGTJRERzZH6ERt1xHJJ8S5Mc6jW3xzr/NI3nHUSw8F9N
mMaQty+/goPvk8Z+9u8sElJI3gbL+t7spgQloHOWo0OT6X0rnnh2x5mJrL9EwQiuTT5EB8ZmWzIb
yXQQSI1Sr84Oj3Z+72Lpj2u3TCVSwEwd2P52djuOuFE/FFMigiJuhVOhzm0+zqfgbtociIMQDsnQ
rz+WvqckQRv9k0SBBkKZvd6KQb9XBF1dzOB3K4cGl1+4XY3aWJ1bxCq1Y1H3r0UBaDPSuVBuehZV
UdwcrbwhNhtt3Qt+xlraxcZ65A8Pz06QiXvH3Gi3M3+1kVyB/yptB85iFYORWaqx0UjL+OWdkXGP
hyca5+ZhGlNoUZfWUWxNrsmSFkPtnPNoWvUu2WdDf1rE+5mcHK+SQ5v3wIu6MQCs8L9YnLbg0qrO
v7CH8swPNb1Yt9XZtgEIP4uS6ZVu9O511w/hOQJxkfOdXz6GtSDR4nmI7LmzNM5kX/y7gy7RfVkQ
udHMQjXPMioaA18tfrF7qJ/QozmSKKQjNbErE5qt/hWf35ICshqsrDCpCvVdRXn5r79WPWjSqY5s
1s3j7NLadcZMcyQc2BAULb3woG4+XlVm1PPhPg2H8h9p6ZLVssRmSzmSf6H0QeVDx6IgP+fua7s3
lcXUNv/1E9YumwgomRyrLYqpM+zBNHObhYQHKiN4tX4SrojmUoEmceFU7LUbx5lnfGZ6T2bozOvR
O9b6miy8YJRLlBFCRwPaSaKiH5nAhrtAW5r4MprM2SYiFgA8zYHQjxIxhagbze4ACMmsKFfSUze2
8nm9qp2/+OeT+xQk+DJmsKk0cV5tye5cHvkyz/N8B0Xbu+DhwxS7PYw1LZQNPDJ9nW8SvBG10Bbh
GRCBzTcdsNLuQNY14GwDlJqnyy1eG8MyxOEUo4zyaE/aLC1mMMs2CDkLB4pdfDfNRws/e2ei/Gh1
hfkMPSaoSxztGQqQWjKrN/sSTi4a1LsPPn6XqWHVKeSKrQ3HlYyCAX8HL7HFEqCz0lyotxbTI9j7
119NfV7scBSanwyI3/OyhWeVe13FgaJqJJbD9dvaKUdQ5FgoKbtkXAejuiZJ5YZr8R4SVtOBBCEE
RwwN7+G0fHATcRkgDoTvwVFtYsoiP9cWYvJqcAewXiLkFYa4U6WJ2yrMG19KQXqaROKtnfdDjEgs
/l9wndJoc2zzB55nbiaV4IbfU7b8KdTqQSkhr6SitcfuSZqaMnutp6lSfRRP0PZefUEA7sT6UDtV
mvuMueeVt9l+FzK8fJTQ1OegrkaVT6w7b/1ytKCKMSPNutFpAzoFvpcjWdyGqxFQ/Yqsyj062PZS
2apeHZQv3p/8K66o2K9jpgDusW7+wEK3j38E9fMH9f8ESGjP3MnTH5UXDJYDLdNixoLNpcqUcAXm
qInF3dvwAkrJ8fC3JbyTcJG75YG+/yjFmkydiGw2+i6fMll0IyGTYxOogJd+Z7rSgtYcapSK4mCK
cnt/uDTJfYmBZLM3AB5yyQZQAPGFQ+PRSE4e9n9pmXkMhQQU79wTyFkirOWulW6Tjzh55mw7DtGc
opoHqaHwHJo7w1o45QC/egkElkBr2AG3dwfKYaXTYvKbY5kcs7yhjaoZbhYew4dq7wAV0W1gPqBD
CIVng5VKwAY5tTu+six5oybBf3b0AlM/fFwwVj2joZTfBe82dV7gG5keqdwkZ8dwYpU+da9Zp9Gq
amxXdzt5bJrbqLiBjMk0cPx1PqtGZWg0rC0gXJ/SzznoXIn6GrMJlSOCyuIFEEqR1GZYUaeV77Bs
ZIc7FehisBqme10J+kL/l+0RR6qBGKwOZ7jmmBTOeMGbZu/Zr+0Nkgp22ErJVHWphZBeftotZm8q
iy7zLnhFHLzr9SPLcLRzfFC7cKpzQWjLgx0GePiMoODZSlCmpdBtT/jYM4yn/RDO7OFXskBPVV2R
18rYPmyqyFxoS/eLUy4lvOixXpto11YEpTcvs/mHGFaO4bNgJTgxlwIbdIkOJC/YUwM3I0t3BbP3
qHNPZJ+2waK+6eVc6XK8Jm3jPTD4EsJt1Lkjmr6KyitA2SixHaV1Kenp953sB+3Ij0vkfzoIWq9l
MRZqb5ChLfXo32tmY/Z5PXrrHEjMeFYCsZfTXMpl1HeAv5GREn46LMBZCijSD6dteE88RdswmRwP
Dj7WfLZltomlM7y/Rmbxhlkh3mVdN8tE8PiNQzEbf5+xTH+hPcVdDrOyNKWgBMLKEZ2OEyCxE8Oc
NuOEp5cte8G0ugDemc1dhh7Rv7HDV4efsx5n7ILSkGm/0kOwv1fCbE2VlvSCwyEl78Pzk057XIkh
QCgVMWAy+2Y1Eu76jPbp9Hbk5sYGsBLaKKazvbRi58fh8J9p7D1eHxsXm+vlVrsTNS+WkInWxtnS
6YEt/0iJ0PRJYbfTxsDc+LKfwYWyRdyReKZF7WfHZ4k+A9+QROIFKYgRCkqh88O4gMat9cjvigNd
TSiqpYCKs4I9SPohuvflzkm7790noiCSu7mV98erVMOEjc9TzOvvurJIzUWZ9gguyQ5q6glTlvAg
7ns3wkL4eNAO/zyj6l2TzOnlaIGYBl4UbUAbWSmCWvJAXB0fKY5k5QOZ9qJA+7JetSmvDLEv0v/x
dIaYCY5FB2ijRs4295M9eJ8nIYGz5nCgAEuetEvcPt5K3zyhwUK/tAeM5K00o7D214O/Vz39oObE
aRRkTxvaMWgjq+Mia+VgFFekLAkKTwX0SpPJxXQCyrt9mecII+LrjllCpmff5wnqwVszHjygpKV5
ecQ9ToU2Gx4n3EokZL8v+UbxfqTRrM3Ya92gSJ+EwoKSZbI6GhgZpeWh7o76iJBxtYHYL2kzBATG
AbXOeC9uyHvoKaTRFECIqF46owosGdTCDxCeX6+S89bpcpVi0U5UVoVdjYoB0QoYMxtCKEZJ3tTz
n6jB20Z/UUjdYSpEVopjOYxKVDJpjepHG8zqMl+Wckx3ckS5S0ypkla3pwMA4D0Co7Oy5jREUJvF
3Gkov7M5PtXPlO7tFMc62Ecc1g+ys0Aa+vqtOWzC+fei828s2rv8pWcz25XhXvXHuzdacLb5oXLl
fDlkBp96/t80xwO+tnc5iG+kKbNKH8I1sxAPj8MGWrRUGyoYrSN/i9docJFEmZYbxnesLJnjSCtF
TPkYcFBPthQXm4ayzt5O+seJlH/edvfWgCoVl1sQDlEhUW37YcQ9RP2kaT//DmomhESXgedCvYsg
Omkf0YjHLSFiC6Z3SFqPBtR09k2AKlTcFbrdPvQo1Xd1mT/elFIQsg2sdQekSsAxQpkDMbETkDPt
92dTmwewv/wiQsogwQ0kEiorzABEizgTlG1YNxnlNX87oADpazYAPQmKjAansGjBMRK6Fjoe26K6
YphKw8Y74Bkqd/DG5Yu3u9FIbcuMXKGVAtR6tMVqgPMmwrroc83+pVeCAGI2pzHeQirU9psgVbPO
j+K7dst89SbFwY1mXUuL0mbG32I9jNZV0u57DiSlmYRPSXc86Blnk23ZEVEkbxLhklvXCBjHHTcD
aas+fwDNz7sdv/7o1k71g+ODkD5NbcSNoDU/EtBTNCVnlUNRZny9FbAr3OSwByNukUV3pQPpqL0t
vCO2pdzNWd9CL7W11ZIUMI7xO5grcTu8ibGtfCvMMxUq5vCEShBwS2scmvLjTNxl4O6QIbYhk2D8
nMgouGANWtRv3CnM20O8+7LbVx4R+ca8mRAQR/9Fo5cLOoMB6vBBvOjGQ7bT0wTtk9WVrAmgf0aQ
cyMhnp/88PEufmn9awVpEjxTM7jw4siMsZt5bxNZ34P3eeWi5K0jfOL9I4Eb6TNNkAE6NK0U/RE+
PaegI0xWPqF1PXwfKmtHUI3kKcPyf01KB0M8O+EGH1weshxtAIAdpTqYMjv18mTYPbk1o4r6oygs
BGTSVfA7V1AWk2ezA21FlPzMLjAXiyyitwlBq0YbVJUIUaEz1BWnVjtq1At6UbZHvetYfakVshw3
LNkqaKW+lvY4sJCMruIDv/WGLVoreQ27UfhqG31/3tv4pZvA3m9PiVjs9mPcVBA3Uxc7ueRc4hlT
fvxABcZa/G5MEPlokVSptL7klHMtDOcWibe2rt1DEgo68M9/pMneiVV6JMhuSQidnIlKudZeAVKm
x0EXTjZvTS/KvmhUv0HQxunnwUUy/Hw5QxlAcUqbIdzJGZXolb9TuqfjAAfA+q1mCLcNmWR+Og5b
OQvLD7BA5naG9mwoOAcGDO+1I3DO65FsoIUZwAUGrBcCDRSkWOGqsC159IZz8HVKFyMIbnVQaYOC
F9n99CMguGUJ215vnh7HxkVVPAwZIpfSwCFVL7r2GUBjKlASwfaK7dWnYNof+ZU2YcfWi3mtIbIe
3JupqrgDZqKnVRIzzMvDqvkB08+Xa27VVaJZOaWLve3mbgQgaQEDMeHtahn0fX4US+rLJ0xlMcLC
+QyhgOjUeDEbJ8tmeRd/HETYwNCq2SAR+v/3VtTBfVB+50cvrL+BzhDwI8knviLOKOTuS3jwT7HK
dO40iOIOVCvWBR6ikYvRGBBFB+vLzdmbni64uA2XY3EgNi1N+3uZgEBHC2tKtog+ZceAyL0YXloQ
HzTL+iKTVi8mpP6VKYhxkVbCIkZjQyZ7ggal5GQnxvMA4KUNuqZ3GuX6+D47BRkg1J3V550leYz9
SyCXm9107O1NOjfT83+aztKeD4ThYSoP40ciofdupJMmlZK8rPdHvTFcLs6Vttic7jROfw4GBjJd
+27gQrrTeAc0N2NwRTWk67Y8jcs6q8CDVDkhhKkcjM/okFEBDRbCwCyY/CugJ8SKSGxdTzHYa7sO
tGdjOpnnRmpDOwhX3atvcTDQjEw5D0QDTkSIRWXAQRQsrcEf2oHyCQ9/Lmitu/XFJmIxcXEDryEX
4VShMLT/K8AF+dZ8l5ywXIAvvlwv8GjCQdM97Giqyqx52xMUMIz1rZP308UHKQMUe5oFtOLVSOtX
tVn7SvuZi0PZyVg6t5sRJzj2QhSxrCveYw+ve9PYsCD3BBMV3j9W5+p8k8R9E7X83Vy8PYaln9+I
hJZh1VjzpHRXWoXlcBukB0JBfxTRprGtMC2Hgere1EUNJKa3LJ404gNTr1SFwKkiPEnsxu3acQT7
oYMqv2rgr9Jj6jN8UFe3083enYKZBDBotKS9Gjwar0fvcSZcvE+zrxilfH4QP+ImHTmKPIeEzTz1
s+TR+U3VEM2AHvKLYwHVoFTYwsuKla0FsDxuOMljn4VngKi3HjLA3pHLl1WdOXnU3reAg1/X64Bh
gHUfw5bA5S13m2ta5RHOOf4fR4O/mb3fPtLOthz/mYOyuZd0hcsB9FT0mquf7hURCAVXHfpw8/ya
s1GF9vzosyBKQaMR325YftjVTebNxCGpVSLwYpGG9+gz2Q57i0rGaV2fF8TQ294IxN+fzC/wFduo
w0UIsc2S9m5Imb+F0gq7EMFl97IYteaoof6UW4ewtxzNSQLhfI8ZKAtq1t3k29DKmhfHYiAjIxwn
lsVbpaPo60UWLzbpCyOke08v12w+RbGSqE1eCWazxuOhcVFVQS7Tc350n/ZNxPfDJOy07tuBRKnN
TMAXlvolgpNCuLK7XX/r1d2BSpdmF3W6j6r4G3Dfi5EvQs7jxgsA1hyWTJNZaXeKyzJoC+ckOpdn
4YuCyIxWENdGGGMJb0xz7NNGEFqY2p2uGLf2i2PTajOT+R/iRcZSsNDavZ9UXRLkS1h6mv3Iua9X
ASslDWIXGBOs7ZJKiTa9G7YCTKUHkSdtY3wtCJ9zBaROzekBFkchz75TRcgHsf5y/H5bywokcg+I
VBrdXjhL/O1XR8MPVfKt2JaB2C+bAmxbarHWzaVgmuPjYxt/QU5FPQkofVLGjd6t/MJm01wrPJpV
UoAAoEyf1Gpalh9yecVhpFv+ajqrYl5bP5fAg+f8ojUH//KsBZzaXqXqsn/YRxxuwvTDqmLfhECm
GzI8ycAN/cM668X/C3RpBQ2AtJ1CJWmYp0XZxp942uHD2Qg7dA0OrMoKiATSF9DxAlQip1jVNzZH
WkIdDT42iLEQd//Gpgwd7XIMs5ZkKbj7WzkPbrnWUZrG/N2nuav0pKmCtoDAN7sK6494v9WAYTbh
vsSQjfmJnGE7WDAMFOVmR4tMJajTh602zpR5XNsZnv64FcE/FRnzm1jlXAtsjuOQXFJGC3xsgoMD
73vrxEeQVaYRcaTTKHtBeYu6jSjkOmkyRh3dsXxIPA9nC3opvRxWyYsg0zF2B/u64ke0NZv4Cqbh
b4BUl9Jszvv7LQDbIHS/at2RvOZLTEgLx3fdtovHJyjaex3Bl+6O4iMLmaGVaDtBTDlZmEvr9jse
OSzhIikrM6fT+m2MoyTRUTSEARqFwfwRL2y7p0IDMJJyWBsdPD5iIG94MTOi1dWFfNtZWHAH/Pyu
d7owG4jY/y6t3fM78xDwyJdgeh3zqcIh3R9gWIjrVQq/v/kZPTTRuVv8VuML2KR70aB8N/4pQg83
wktVK2mtjsjnUgx182UhzL6pzGnhe6hyvX3A64tDC25LYWYOnyOYCvjXaFlBXi7+E5owjUKw5heW
Z63e6xQVafiA9DUkdHJbNHgqp+m4iSl1TJk1mE7N7h+OAKEUSRvTggSLd48QE5Rz449da0PQPF4m
OeJLMau7Aoxm9Q03yS6BbkeEwwgYoijwdHLxZLh88JyHB9VqNXkjXc3C3Hq7z6eC7F4IcSNKWlb6
3vnBCjIRzfHKFNoKA5m8N4VnODzyjb0eVx4o5n8w6eDUxs1JcBdD6jab83nOzoVydGIElDMyMxwt
MA4CKq2a8gJYTQhQJjd/TtbV4HFKrMipijlZbNzfu1TB/tFRKBlLOIU0BA0lvQ+pIVm7CvY5itRg
w6zTcUYzBaCesK0z3OVmxkCr15LlmzgtrGEBysdjkK72XYqSGNE3grVRtHZEGCZhVIQAXkRrYRoJ
n5BSzhqvaFDNhowWFWG2ISoVXjKUJE4UzTRNlKBvi1C0ag4hFslsF5Aa6ZlB/+GLqG/M9G2Xs9KJ
BIIrX8wyQaGHDusf305vD/XYlk5xYNwC+Un0OuhYSsBPhWcv3YXeQZ3Yy+LK2oj2p7bOLA7uJNtV
Qz/pRvFLFzJ609hJBPyDXYNQQvXjq6waLzcKKD3XxfTongwyZUhFFoxEF+yJYY63J7biwIy/imMX
ui2UBHlBzTQQQNU4tsPtE8pbOP9djHnlewj/iAGBk8Pt2k0xeuF/+xgEd51MRTKRvKWjM6E5FXlD
/FwlobJ8bUIAuTj5DJl75VZvoBupOINdbkDXfdPGIyMa5zNsmvMfw/HHqXV3FufqNXs0HNFP8+Za
8dhRMR4lMZ313y5U2Y+kMSucsMOBZGHdZqdzKiXW3QC0Gtq+HD+3FwyhA8EdLmcuidIIhrtBtn9u
pk64eMh+V89d4fkT1NAu184ZbtUh2vCBehghS+JjzvDzk6g5AFjEDlC4nPi+4OWPiCgC0WNvmP9Y
Llmwa+coLu3sX2uHaVNKNbcpmdXeZlsKcNzNPDVxwmMSJLn7Xo1gYLte56Plxfb8Tkd5V9IckcRd
F4dD0WUcx0shrr4gAi3U3HVYLXrSGmHMmMXf7p/IMlaBcM2PNF/YdDSfUMDVO+8Ei6BW8M8gDzix
ZDzKbVm5lEvah3BJEGYjGMs8mnfLBmGQ+OEQf4TTXFSFCrB6fTCqcA7wZKt1OKhd9Rz8YBovXnuF
XifYgT+ov2xe+lSxmwgWYUbVtBCFXGUDASGxRE+quR/8Mn+omugC+HD8G4yRALl1Tl4yGzojWeUV
/J77dkWi9q/3zp41xvzw9bESvv/W3piQ0XS/7oU0uEGT3sRdpIo2eZzxTyU/XTPQ7ElogKg/GZFi
MYNwNl1/fxqWKDSNn5NrZVtKbvXTBvCE76gqftw4T9aIFJNNV90+y3pYylaWrHx8ixYlztwwENEe
LmS9zKjbXhJIBmUYwA==
`protect end_protected
