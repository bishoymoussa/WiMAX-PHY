-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
vy77UkWT/EzRN3Egctc6Ff+NqjrNcw5CyY2kmdugf6MjC+eutrZVS/RbuR5suIhbOOsen8qnCrCG
eeVxAhdY91sRmK6vZkp+QLwcYD9etBF/p7zVG32MjTakG4ztBTsPNDWscV1v6Zr4U+gvVa/LGrMb
AVKEdVqMxUnxife13V5FEHEcaSfUqI+DcgU9J7H5E8tt8KDpnUvSmTOX/t7WX+ffdZAJdA51aslO
fNuf4P0I++uLuQNgRN9pJgtG1lnTZATtN8CQd86EAlLtH+dzFXqYdnF6jTrqSjb/0J6RvFTjsWoI
HP0gEtb+ygVXeUZYeVVYAkMZrBPQ/GOVWCUY/A==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 13296)
`protect data_block
ONzCy6IvuzAZKbEltvv43vseUX4ttgJqT19vJqFwc+BUCmpwOhW8FLK8hmlmERrngpwtxlPpbceS
/2i/Wxeh808pPIqh2kIYZk0QMdfwjvxsHkl/PzxPhBMmBKpqDUIXCdRvpJPs+WcltJjZYn0Ze+8x
BtQ3zU9ohFbkUH6XRNbb0E3Ftr4Zh7bwVMHwA/h1Y7zSw6z//0RB3DJVG8u79jb2cC6Do/amP+8z
gzwnwb793g2H/UyfbyrVCRXrvUvWmIhsHmcBGU6jeZIHoXWkdd4CPM4VeCcYCtuhDnrZ1ncSPzY5
OpJt3AQfMOpKFdOS57i/5/TynQ8fXgTrEZqu7oTavXWlhcsy82vURF4LSMxbhstQWCT4KZUF/nmB
rIOJyU/QYC5c5SZCfrngYmzl+bAjz+URUpQVaN8PfHFZuaCOhn8MTgFmsDIjkUtghd0cZToZ8aYO
iqkJkiOjhFiIpDJZx3tCfnzvltFll367mmxb5UXbx+SMnQr6Wh578bPvUY2LbcanTS20cC4MnVyu
Z0mwLOC3Lr8nrQ3Zm6Zew5+WkCN0nf5O+6nhkPvB7RvW+MmxYgeHgDuZyY++FRY4HmaESvbyNS7P
cND7sU6BLb66GffiQ/UlzjN8NajP5F68k6G2IB1HJaJ2/RYSnzhfjFejKgLzQF91BE2KTwwWg4qj
0Cft6g3FcaieAJ8xHep58HOYBHdMQ0AwmbXiNxVOlzy7LzmLwFcyxMc2v4grNjTH3fqj1M6z/yQg
b5ymYjRkoH1NEkNBdQqxmmHhyY2FJ/x2JttDiqfajEQbtD40Z0XsGFlh54jKTGuW2H5MZ9T2ezAR
OiPcFbiykBF1GAo4NfghPq0nhhQbwJCDvgdhCnqZzKwDePaHZ+SODe5RjBEEGb9cJMJ8b1tXmu1H
jRX22iwnAfXDhMrVgX4+w+0ERZ9lQ1IP/wkKtjscU+Z5S53KHs+eVzPAB/gRonkObyOvbpq+FkEs
sZTdTmKD5DPADTNmvy/72Qp9gcCddx4j6s1czoq7E4+8folSZtzeaQ8dPuIJQXBnUztiR8tCESf0
oNzLsGqjp6F3rSO371eemb7j99JqLed7A1PTwx9BuCjEGwrJaK3qQlKQMSe2OAFQKPiQa8HYFHc9
DP7QBAAKAycgfj3GCt4ANdGp07IncpZ9+CNxJXC0S+PE5JWgbRW/4xPyJD1ux5jEGD4OM4s/lgwI
0Az+19H3tI5HKGATJRBHeTgJVZSG400ivbVC+9Y5T/t/S3gyOeRqirLr4jlohNE3+bYX11qiG/5E
TTahDRVn6Y0T+TIDqWc08vdMLrmd8Ra/3Bz9yMCci1hOB1bOIlgmZZnG/qBrInSP4P0C/hbwGFQz
eCsL80iLmAer7UeOzmyOew3xcijrvuJ4cwRucTc/39d9hNPzrccJGmA5VUkEUpGNhrTlpC30GBcj
x9VAiF3XvB/gusXw3yWmcMuPUeUHamMAw2mRjDsbn6ikITymGEKOdhA/i35IJXgRCHjJQfKndXcz
4iYms9qYZbuU8lH6AZFNCS8e+4xoyrpvtRUntPBj2XatDhLSMkbjHOk3kdLqcWiJLBHozkHVH7un
dsN7Xti7bPi78FFix+6gcSmHALSGXjwA6SCkD5DHy18F2N33iX1kSM8PEFoUZw0ilukd8vCQ5JKv
0yaYd9NEYsoHEY4IesXwBRTK11jkF20T8V7sw+vtLSswUzL1R2HN+iKvDHKksO9Yj65xWv3+1M23
TpKRsvFkCKxx5bVIJbCNh6WuYRjOz6gt3rfUHnfQ6eQIxn40aOCmIw7U8N/bktp2I1ik57oQ840e
Ke0fDUJAUoogJ5aq1gogRxTQ6rYYjsq2pdjbz01kvZN6an/eTKc99uzyBEVPYd+i+1PE6N7yDjlh
RG95mfYkccqhwEf0753ihBP12btuY2Ss0QP1atx6YxrcQg1+BnZu1PnF1fVzjXx3p9Lx7I70Hxsi
u5MU7w5/L52hvzbhOaJAZVqxRmWd/Y0/wvy3uGzL17dO3hOAE7yFWkOl+Xf04LJMaf16tEn2HB8i
tzqt6wZJD6sP8NkjoMyNQrhIrfLnK+66PYLVm7IxJsMNS2y0ISTAdHEnnPcqOj0o5gbMP+UhyngO
NF5bB0LBJmydOJ6+xGCtfcow0/WNisRLFU6OOOGGImsk5JTd7jnHxU6fNvqeyMaWvRyxEFV/D8L3
CJGSWcHbDdkZ3fjEq2fs3AnZsW7mzOyHq9kRjrU9f7J8zxamk+91qI0F2vRcdC5+0kjS0p5Ax1Q8
euleFcKRDc2yMBRP6sJcJD/Hdw2fFfoWeg6Udv401tXDo+CXveM2SRpY8fsiefHj+nlG3+cjAedb
XyCEBmFL0dI4UVmBwWIEvAA4sv6zVWxY8b37nzybWj5MnRix8HAa6BRrUG9LYYyWWFB8wGpgJ9wD
72LE7NEAszfO78B5Tg81vkEofXlO9aWxHjAAMbOnjdbvtcNSdhFKqPipcDhtr35lUtsBTw+19JxS
+zAM79w0T+e9Oj8BTa7/hsStPrpnAZ5FPoeO8hptagwKs4dPESgoc2CvvHKL8yD88od1KEwBID6o
ItK40Fri/ihzX78cGcaDRns+4k8mSf92HDrf7Zme51lBUoN3jf44+bV+jFzE54Ir4p86Ux1UEagI
QpnXc9DGji/R8xwKGMa67QMSsbAA5ey1Y+QNLTqvThNMZHWS3oTxi+PSBCnWdrhits11unG/MT24
Fo94s4FMH3QFof+NvjaHCemt8pnYav+xkJUiD5a6CsaKMPVJdY3X0ixT8IDWG/CIukYJPDSfB3+T
RdRNb3hBWQRaDIYbVIj9dq4unweNyYuSegype0IZ3scKl8ygstP4PzyxsVKX1nuzU0i3cEHkz/Ef
R4Dui9fVuQBXGwZuvkUEyRHKu/3HY6VGgzvnBOpPTU55+QyQ06buRRqI2gawI7A/NwuLG0emM9HG
jHnDvYYfsCegxBRV6gE5HcG3G0SFO4p9Ksj+5BX/Txzp/qxaElYfojYBhFZ2imPai2on/Akw1CdD
Z4ApRuM+aB2Ivn19gnOuwiKBT/I5f8YAgdV5jVUo8ZYqJYZOZQNPTFbmHVHptooD++oKQKSDjQwJ
VstKTsAdEe55wIcnpqEeuLt3dkbCBT6WvHomd0w53RjipkZeweUP2sG0tIOeBMppvdjLTS7JjSk1
m0mZKaYqP/quELVSVoT6LGvKxIcqfdzZEM0K7j1W7D4n+Rdh5d0an/Mu3sAsrMm/9eNwGmMUIj8o
2a5cz1x6mFzMtuRCVi/Y8o/0j7LYstA2vzgpwqcL90fGbX78dVgMERmWMK8uur/uuCGlkRQdx/ic
7DvYWRAeW0ypemHrDRMzeg7yB5f2PZL/ighSkoKHsyjSR6PNQ1+CN1FjpTSGJagzdAuyEV0+VRea
qbfqZDEgZjS/oLivesVhZ28vq6/vFYWwKVbbtxJqX7l04Z4MPGips0Wg5kgKUAP1xXET4o7PKF+R
VdcpXXdMmsD5G6veRsnMf1tZs+AVzbsDjjRxDfTm0OHinJu0RUQRgxpL8w2IjWmnKibPnVg0HEhu
GFIcZlREuKTlvGHe87gQ3w3HfSgJtyTXwbGJ+ecTUFFL+xuiK/PNp0ZoaqXwzp+y+rUFZ5Ba7VVq
MRYtkQFj0DIYT9rp4/0UHTcXtxNKNFmZhuDJzFseviriM51ycGJ2Oa0JFqqsoobMylX1YfmMHd2V
q1tjx+cI+1DR/kgPKxuZ27wrHmAWc3MpuJEbLvfCUCCM0amH7ptJNpvq0ja93+CRI4hUzF+yG0gN
jSUiKgFGTscnL71mZ6XHAFbOGxe/2bW/faxHyqzdZFEpwVYT9h1sWaVYNikesI0EdeBQ7fvALjkM
IaNW2xSeLgrecxrhmt1Q8tFFVL7BqwaZbqtURHsu07lKlv07Mo5Y8btpeUCgKgkCd3VtFrskVji/
uu1/pdY50aetxMOthfuADzItFUgTUQwhaifhd4WBjXZ39qxw6DQ6z6tf5jMh9p27WTDzdleI+vFe
vTQbeD6iek/kp5rtoktZc5PFXAsIFRFLBseNTU/gV9fUw6Wh1r+o3d0luUwxGvNEQfJw+rwH3L+E
6uJUJsRCQq+g3VlRsF2RuZyHOutwTmzyZcyez2B1gNIMPOhI2QMferofHgmFgYKbJ/f3GT/0UBmA
AWNQwlOTxz/JZuvKx0Kdwn6AYhJ9eKEkHjQcuGXRrqrHPjvYCyVQF18MdWC1P5FFC/wOkn+UnbeD
kn9VfeN0T5cxFjHaCJMol0EVARkg6hJle87DyZkpWrO05BSgPnLGVAbLkOFL4c1yZGxRN3sesCj2
1amg+BGIfGAB5Ho3QB6JHS8V8Ure+q7KG4IVm95cEHU2/mgM9ZSB7TIAMM5EqD/841+/hqc4yzCx
gCeU1b4E1WDiTCJuumpIA+/ixBPHYI0RyCHV2brH4ySG8AAgwftCE90MQOSWqQgZbEabEbp4zPXu
U/FmbJzQxJky2CwAAoYJbrP7745IQ8ZeGXNbXZm+C4MSZ5USesU10rs3N51D9br7YA7ir9P6T8P6
lymhP3NKi8KwiqfpvBEKH3WDKhnZSxpKAGxkcvlhS4bz16mAH7p2HLRoZcDeb2XvKgefYHUPxtFL
yCPvyfqEyZtAsoNvVafVvk2MP+a06Zp6sL31dtTKMNJ0dwfoUiuTYaEgbvT38FBPQyYwGnU19S20
cHNVlkkw7p9bzF6F8Gxkev0IEZ9a/Y3B51EL09Tc1OXV+OHzheoGTvQLCp7wkQNHUU1HBCsPQOjV
8CGx7nbEH40mvwcO+uJrVXdoXyTDjWSfyse61GuQdLbyS7dBSv0wQGrrnRW7md9LqCseyu3Vkhvn
rR12olba/jY7yiDLe4myuHRLTv01i+YBypqG+oOw4LUWwRji0orNF6Wnswm+72nk9sMrxyR8PcVe
V/DfH4ZMQ5mofS5z5rY3rc3/NcYeLOXfAOw1pr7WKnc2utmGv+IXuvQagw7Yamy7zyLElCewUWnS
+ODBm86HvXR1AFG2w0nFYloBn3qzoXmPPEREASgLM+PNY24xH8inDCWlpLdUSm2C1GcuDhER9SYN
Lho+WEhDV+PaJ6fZGbvZl76nXDujkoWD69z1AExbH9eXlSH/qMfXDTukKXjM9YwelsYEVTCe6uq+
F02/dRr+TQUYRmlU9x892I0nxLc8hczJK/IQhCAijn40EmEA7SJ8hFn1wVKruS7WdRbLI12ofGns
HQ7QGhgIW2i704TxoiFgVVodIziW2ClXRNfvQYq/gZoDwxoqd/cYNhnViQSnxOg7YLyfcsy+DUYU
y1Ch9tzvDlyVostkivgaR0VvRPhmdpKYTXu2ELNl2NgkG7De5N7unA7se4epKHr5RNdiwwdufIwv
Zs8Gq8VqjRqKrcJjcx6Hi3hakKVrvn1iqLjwzhVjV6D9pVYjupmeMOh/L/mp8/amU9hNnM2D7fIc
mDzN7cQfm5HAYN/7iGo3cbGn3Mx8o26MD9vM46Tc7zxvr9wS5hcKPIatVPU4cXgnutx6x3jpHNYW
lbaXZLhnYDI6xmi+e0ouyz0JMDkwXk6Pb3Ros+vzI78ONWAqoy6CM3zKKMEnupvPFgoYrx5imBBv
lloasyjQph/FIrgBeKDXLtSn387RLHGRZwEOZnnNW6wNoD4BjcBrtA27DP8cT0B5RO4uh8XAEEsw
zmIfURDCoaE0iJLV1XxqPJIcxcHrWmDNliVICD/+7jsLriXJN5lLM6MzcG9ucdi4xw/irxSvRX7N
lCERlCX7X1r943uOLfwCaujKZB9JWoi12V4pVTpBv4jxZKO5hp6COM0VP5S1fDeuo3zOoHzkcZ6+
EKhpuPVM0aZqjs6WefJjqZ94+uNCELHJZIy8D5oJeu2jXYaZyVeQsbgZkGpIAjK5Rp/R6MboFrwY
TPHSFVUyF7y5RQxgmugHfd5TvTZWwSK43tUAZeYIaDDL+YtxGC6jaoUqQqrTlchAd+0qaVHW8mrw
ZTG4qNinC9Jh38zqnnuAZNS0fu4pgiSDfEbhGDZjdSB/A+SnoNh6s4P+w1Ez9z1xjhyUyEqxMB2G
CBrOqaetSeKQR2MxZWNnJdRkb5jI+1Al5zkrkDDCxa4gtdJ8IbGMseFzuid4fMdJxpFJd2bn31/h
G1PWLF2XPZ2sxrxB01nB/rfON8IkarSwCDh/g6orN2g3lwLTtmp7B1ZeV1tP6eEvOxhtkq0bWsfu
bIh4uhT64JKFK4szUslveWvncaHiJBU+EA/DuiEx93jcjTazOvYjE0m023P2wWlI9JdbAvXeVTW6
alw21wNUbcjY1qKK83vtrt4sRJoTItY0wvKrLG+RuFrsidHpJd18YnTOr4EA7Fq5Z5dqxd17zU21
Vwu/LbmaZZGW9w4BTz3Ku0FS6PUUUg3mFehgWA+orit7xip0CKsnpnKw63mLJUw9alJSobSEBTm6
IkKqkuIM0gleemq3mQyeaf7xpflJcmAnDMFvwqaY5mcduV52SGshRM1y+qLfkKLAOXmUroqapOaJ
lQHVY+HfvympWP0N2Ble3KLKu5NCphs9cCTdNvLzQULasN4pv1qYO7GStvCNGRq/NNnIqJxOFhEf
dR9Ki0NETsK5Yb56R2yBYOWDIXjt2hI5zP8QlrVBLrJ0Ph4jVi33eFGwZOPVJTV4+4q96f2UpTQq
iEQdhtxxzZeADlJxc11VhymLyOej+Wrk2irmmmxt1zR8LhbY0Ic5WKiOFswOMlHJNh2ImSdc6zun
PqkkcnH7MAptrhx2spK/ImwiB3kVS3amX0ZgLAkauwkOU9rZwctr6Us8XUPb3C4uA8wVIYZSllvK
197ZTo2KeWN9T2Wsh7dYhPRKo71FVL4oKMBTyiZmPM56skDJ2SqAGpANHonid27PW7sIiIpdzxQj
KIKHPcEgYblIQP1Pw6ojb5zL2jdt3eaObfQdT86QFhEmLU8MQS2ZBoPCA9L9UhqJ+WKYwL58dSfI
9LAC4AAYAbGwg26mtGJCW8RRbXdii9EaGrYcKYeSc7Fv7L08LcaJdXPHs9EHht7FHj9+poIhvxbL
eDddAdYZ3TYbXYVdRhNtLqMLeD+nUihenrL6YuhfymF9WChPvtXlvs9jUgnJ4TYBzqMMXTrIiA9B
vg8SXcwxe+W0zQIoOBxPtKcG2ro6+cZuXRl3fJHi7PZ45Dwz4+L4RhNV9Q6RlBqAiF0bNQVLLyvQ
mbuphQG71EUBfU2uzJkRjbuB4vCsZDlttdKTb5Qy2eJMa2G0MO6Kt4josr3bn4aoPtLA2mI8ZB2V
/YJU3FHawZkU7gV3iL7AYR4DhaILR/DQEqsva0+MV89iBAwgmRijezYLyuxuzucCfBN0PNQK/JXN
Aj6zRgaIQR0wX8Td6rXOo62VlB5xU4qtQUAZ1xBQbUBPFBl2pUM0zT6pyiVUioITULl5U46q17yt
7FxzTLe2RN2RBaux3y0oFp9VChMprvcl0LnLVwx4zAHbbgokcY1xmKlYcKi+hOaYopSbLmC/lCek
97zYxlYQM/BrG/4FFJW/Js/sDjS3xyTBnDL+tkB9Z6LOwgLXB8WidJ60xHEnLJpHtPbngRD0YTjQ
FzgBQ2HFd+/N5Ti3Rdz2UPi9jD/VeCVUwbInI0y+3664cDNJzb3ZDx3vcbGFJ4qSo8cIq+j2IAqU
UuPC2LcErNx5UrgHnkfblVfP6Ww34GEPYrnuLN58yOpWq2OwzQUIcp1WjS/dLFQA/oFUhzqvGFN9
O87peiowVshQOHX8k3Cb+ZZdph6LzYvU2u813g2e9EHwSL3qeZf9FOgxwvwe8O6rXwfSZzWhgOnW
KYxa1e0YTNSjN2nhHw+Wl1b97sLZg+hLfFoHOP3Yo1D4jGYr4wKU7DFqlbeNlFEd2wH0MtSCfU2D
dlKYPPPr5VGqCYva2Bx1ni4Lj/xuOE/6KzXiiGy1s+UlIHsTakHUKS3k68a7mZ7HRmuv09c9Y7gi
aGXphh7/OdXIjg/nwMTdaT+1bQnR6gvVU+DVQnnGODQJHIM07mIqA6AjE9XY2qasWhR70bZhkZ7b
G13f3K2wJRNLeIlsa7JBu57yHI3U+rnbsjUMinMhIVkRzzCbpZ7JWNKG2EGAk5hHvB0nHkaY9i3i
5mGM4/WK1jIi1gfT9k8Ek+gnKztU/ebMhr4MJo1P0+yX5bzSJdL70L+fEfonxKxxTjhBhNDCoU5q
1/rS4orJhzQsr4nd7RbcV0jaROw8ea+t40i3apRLsLbZnUb+ObjLLX+4rwHnVChEB4BqKpI37tJ4
GmQkCZwUEDivYvCRA6HWllBMVD58p6V9iAs1hnl3KfeYYVaYu0Rfq1w1x6ufE4ujtBXMp2irmwZY
J3f79j5QfePSinupaWOL8Vce3TDw7fxpUOdWSBn0Uw6SNEZwaai+PC2K5A1mRKaLURTtQD39JZ2g
UD3AOq+QtfHp+1bnfcsPmzLNEvcZAJLvE4tgLqYObbOja0SQ0CnbzZeYh+e13qXlb2ysbAMEPFHu
u/ZCnOxRGvUnzYGqJDlMbpFF9LGXuD+fpSdog1klI9sdoYj21w2ge2ufFCM19wVsLcn2QvKb8qNG
6YtgvRY697nE3w4qC+vZ9AEkYrqC40Tnng65H3f5KRQC5Evxeq0Y7SwXWcOgEFtC7GlAlgbTNR0B
Wikk/zDGtV0qPd9L4gEC9eeWgnUxF4MkH4Ai/vgK4102xWgwpMCThjDujSPUtSxq/CzuUnA3hNOE
eSf5ZHWRGTRa+g66ep7X0VmTgkBkWfQ34Rxft6p//Oz+zDe4g4xI6l1HubxJ6dZKR17MqkQOVIQm
Rtj8K0pRHwRqFpDxT9SWNr5ghRnzr6aFchxyS7acGd6Vs8AMeE93+PJ34N7iIFUdk7J7Fxwgp+Vh
tzvu0OmApLAFQBy1m1HUqNeHkjXY6KoMRT8C8AYNmWvQAibB/gGmEIQFHr8xBWG9rKyLBsRoENpo
1xLGERNVgy8wMq54eUKFtxL8VsdU7MIOGLytK+bK+jZPx5QWexhw3h6saMEZ07huvGf1HfWciOgw
o8Od6w0E/LLyFFkgEBnAt1rd3q9TLU8rPoFmn8MDCafbsFGqKC9SxNNAawhRw8KH686Nh9jwZD3I
Wvcmxgt+ICCzVnHiWGqzM4izstcKEbP8LeTTO4IzqCSJSdGxZzqqCLpLB84e8O4rqUSy6dxDrX3H
RzVgcZPY2cQX6rUSTxWFWSr14TwW/unslFpzOLm4AUBfybatUqTMvZhL4w6P8FHeyPpQibruf5+c
iKAiMCXlQxNl2FBUbvzCHnooKFw/8YaLUe6ZV1ZbrQJosLE92uQ8iRxgkXASD4ROSJfwHR4EsH2x
Jx/vKZmpW5QMOKMcxW7fv/2dkPPW4x0f5M2sNPy1VX9kcxZ2XVyim0O09qPcyXns+k/gPWPiRpQ8
KKf0qOeXcvbiY9wtilDx1UFG2D2igmTLMII9uZFcBftUxt65Lgd7+m06RwW9FYcFmRwL2R74CwtU
Qvf6Xoq+BTDZeyoIJ1YRXg2tpGwWa+WxvTvVwuXDVu2XKSnjg3qCcQ5Caqzwh4XkvIb3iGXoPRab
2PJg2lVi6ebw29Cdjdc7KOIN7qimd5m+ivgKnojskFUAlpyYYnzjUzNNQADsXB+k8g0xQEabX8io
LLzam1izTa899zUhqCAmgT1A/u4+kpfJcqpVY+mI5v21wcoLrHGvL+NagicDwt+9Ia59aDrsZsPi
Yl9yfXxAThjWXIdDzngSfCYUGsMqf5DgovKspoNhdcRJHJMuAsEzNPOHvGOlqoXvMrRxgwi75l4y
uu8kmOBKT42vnEdgE90kI4nWX7jx/Q2rJTqiF/6R4X733nW1VkoLL5va/JMSI45J+wy76eaWf8MK
7Gz1hLACyNjrrHbntL1se+GI2IuenPlIRuz+qy1N5E/sCyQB+j3X0L911tnQ1nDCr2lCYf5Wna0X
tko50pBowUYHSbZ/0tZzt8V5P3Q2NKxM7E5Ent6zThINvA6mxobr+6yjhYTJunVLG+w27qHipbvm
1DbodkVrx+jHwNVS2gpCn8QhZN7RrSShf8835//s9tgn/SGadjMnGCICg9z+x1G4H4aZ2up8X1RH
/h/nniBldjOWwJ+YRyVFiRUCV8rmQf0JkM4+W7wyJ6NA+qI0tfo2yat+70BqS3vcm8X6NdYt3BS9
6fRtDaVzVnAsLC+WLDcF9WwfCj/GkTN5yUuvSc7Tro+5pBOeZwGqMXUx5CAnphsn1rE0TZljF11r
e5uuTc04kiONtXa3iHgqgTI5CJJ5V95Tc12oX73D/JYEN6lDXtjvCY8ht0dfOxw4zdVVPTREi2Wr
ph1cWTYSt6YCFKVzsZ0X4e1eJK3rWGtNaujxcIQFQp3lwZmvlxcKxUjtjSQDEkjvA2E/x582eFnd
+c3GbAdlY6nNEGqQBJq5uaJ1FaefqAHLLeaBt/O+ggmHToiR7l4+SMkSpWMr4nsDw0jiB+rz9BER
+LtwwjH7icanF0BYVtJfp2Ww5NUfrNVgO7ggdXXxFldJMwegX1Dftvzz75+e8EBtl8h6jXQi7y/H
vwd8vOnaOhrEpd97LgFEog4S4syEfEtKMcmhge8MoMAy1THyd7ojrybinSqnC0gmyaLalVmxQ27o
ocBGtePCLnyXC61d9iQrxMfyn+hPyfcx2Gl3ZL4Tqd+cKcAJqOZsXreJ+wOunXCjN0Vt6x3e4Ngy
e46Vme+Oycqc97WjF6cCi2pALktsMLbE8ii9FXIxgKxg7boQFi9SMEk8UZPHbnWH9f2k4ZQgws35
qCJiHgcY6cUp+OPrEaeQwbdVrjemRkLPOfk6I896pS9ESMwUSPyNOmctikcOnZwPGBoYmInuDo5b
R5yJ6wsbMyhncqbAuj1AQBIU/FrpdSapAD4RseGsPQezP6+D0cyF6exL6AfFefKoHSK8URLxF9ta
hrQoQsQX2WqwoW3kZxuTqGeoOY7V3U8YLDOgxIuB5P5y9tyaQTLxtkGTJlcWH6Ofs8e3hhar0YEQ
R1MTHeCTz8U+7GXFGVjxvyHq0x2TYEF28TLbVxq0qFwfn49bfxttumFF2Z9vr/PdGUbNcBjAZaLh
xSH2Czfdc2zU/3Xsn4Z6rlWLGOawzxH/h3gYjFTcClHEML54++5XDQn170VG7Z6AKfITOwD8Wi6l
DvvZiuJcIDMhTBdpvsDd2dQ9Wwok349szUVJF8EwYjsRZZL1gIZlnQ4+ief25IzBKrlimOVCPbs7
wo3yLwnrKSIat30XSWRuXQM6HI7PyK4vlYEuLJMM1gUqQdTghcd/EwaXgyDkK1j8xqfO8QmLIV5B
3yIwnQusMHGpFSkBtilEvMVUlQe6WJjCmRoMwkV9tp3aYA03xNzRMsDA20JOI/K7F/nntoj+zTg0
3O8qJIjqNqsU/ugPcjNl5M8gu6lf7HXIGnE6prk0RwHFCmz3nOAL9WMv+yt/WpuLkbgs1KSMxpx2
ECDaUFPDEPQE+4/WaBLebJh5yAKgvOGs+AjzuRZIKZ4d5MttxssYMLljrTo4Y255gKz8xRQO5kST
Mq/rJtel3VK/UcJd9rlw8ZSXyIDRTBJELOWE0F1HlRm+nLpf3mkNImgP/AyJHYZcUCjsoq9XXTN6
VzZOmcQCLqKQIgR9lQKxF63X8RP1kgjQG6T/6k07FREmof0lpZvbwILF4s7n5sYz6G4fNqQrrVE6
736k3cIDIUpkjrcyRUyNOIkYA1q/GtzQLf10sz6281g9UhnrbxLZpweJ3DS9/JIoEcqib4HeUagj
VnfL7WWzxFXMniY3jEL/LvE7eWz8vw01tkHgehfyUic1jGeFnKQlnx7GzbZFyX+YLYqIIHr+hdYS
szC1OX0SaUJMrVMrpu9KqgyQl1uo0olHWuXH+OZohQjpWdONN1QFbXKekbwmg0B3lNJaYj8nobz3
Vxy0/FfRT+MM0Sf+oh+l1KPkM37tcI954F7/tQyNnR0l4dVZ5EIKFGhuJMLDbnoyYWr2sU5rDRDP
TatEE9T4rDlCuL0YqWCgJg9nDRhwO65G/gYsmPwJ3WNOcNDwQoJvjWlL5b8ZYHTsgKTjSIiQgEHx
MW0xArQZto/cmXtyB8xng3TyrwqzoMmv5a+/rlDJTKp90KFrZn7tUyG1UXxizG9lOp06wRcKQBjE
7H7c8724xd5+sLLaORNBmprBStekUg8eYVl1885s1tOiM3m7CvvSvJO7/PwJqPxnBVLMEZnDGC4G
1gmQhqRKcE9+vV5m1mt1eyn+1c0leJ4i1tsbRXs6AoHPn+SiPSZGVSiPElTawJm0Lu1Wya54nDms
WsTuQDwQrgv5a3ya0i4VSrAVSYZTJTojkVdUC0ZaUef3dKOCdxWzzNEGHuE7CNe+U0RjNWPWJRw1
P2Zim9qb8WsPiCyFYLDOsRyQJVdZkgtyS9CMteQs01SfxTfinV74YIjONFB4g1kzJ5Zv2idLTnWq
x1MNgrETGKLNbEjy7JdwDUIP6+Zje86VDBmvrOxXyl304HZXiRD9tqnezNpHvVQTePJqJfSH4Q7c
1g9Rw77QgxlmUTVLE3WLwf/AYgUyqLheJl03/6NKDn8tC+O3P4oi1jOzxGZ1aUGQ0B7SKmL+PGPA
DDzld8Zrn4RcEr0w3973iuLYYXpPQMMepETtzhj9hTrX9dyCz5yU15xv4vKmCa9Z1Mb6DbDj5IMN
W2VeBTikfAf+2sYW3XA+u/hS8HCyVCbCO0Ok6WNjS+DkUQoHw+h5xKZZxUgWTDRkESsElC4X6j5n
kpR/pNlAPTkCRV+TD+uY5dSSGzbb2shBScWSRErefQNi90OY5R0tbDMmmpdlHHtE7JytgsK5CobB
t0BfHzLSBuoWYRJNr4H1hnHs1w3nWZaEsWdxDirtKXUJlr2UyEzRHmmh0q1UdDQIIVGrZsxVCKGR
ty9U8e1aDy9ZByRLQDURp8Ew8xp6gDkfc56YR8QQNYuBpiX6lMzfKjYOdS4EqUESdVemia7xaDCS
QWqDnzmLcMtGhW9AY2DgkQ4NXiYUu/M+dA4V7EGJ/sOY6KM+NxdnbkDbBuFGhg/fqLQ43lmUMrOo
qI4vj23mEvbUnjEZqTU9mwgPumWDgKCn76Tm161VDNgkPYTQTdj/3G/jdZXkT3I5gCNFBqGL3ykV
8JWO4dTKRyg5DoKcNJ5dqWiZ1RtEFwzyb36DQzx3ihvXO5+4umZxrdhu0dSoevRtAltPFZrQJC10
RN78rV/BM90oObs4U9biC+9Rj8nCBrwXr3IqhsrEukHx+gavtx7PH/w/6ExihczHORKakFmfB4nO
efQO7LZxkYW5HQgrV3LL9NnSsTusxthyFSoeeapRGzR1WzOaJd9bppbpSlR3EqFe8kHOHIGB+3dU
XJb3MRW2elHdDrWLo30zLjVsLU8QsHwgKDurfwR+10pcaZ6ie6VRjKUeQtP+7ZJqJU2j64PEqpVh
ZRxOlBLjVAyL2oA34NxhLcH/GDmvjS6IY5fi164R8beeF2VlL7/kOprwZtmIprBdRnb5eKJpJkNs
7dX2eGtuBA/Wfig3EBtEFfdEuVVJ67kEVOWTW9G6NZI32Jpf7Wag528BmiqZCCbPzRwEdQOtU8EX
aBgcRFcSarQpm09W/y1ydCJYcx8j7sy07WR+pK1mAeiHWTVdDqgJhBiuF/cWO92INVmxmydS8J6J
WgH6k1pknBnX/3w8vQMNcnA7vIWYRvYag8SKxPZO3QVDvhnx7Kcgvv7tOuwwMwZDnPqPAjrIUocN
PzCrXTEnOj+rG8+8wzGPWrbj/ki0h/2bOxzwHyP63PyCUUdpEsAxYi5JfbgegSu00QneQ+s/MBCh
N8lDA72bDf07KDz0p7hj5NsezJowkV0jXAcFjYRRI6IIGFh1g+XrTgVnJ2OFvmSc+HrGcXw1rW3k
/6awGxAa6D2CUPFgnlcyhRuOPe8zzVuGA5HgxAxfSYSC/T0YexPpAeXyj/dFDbB5JAgRgIuwOR9r
8pvXCpEvv/3w/7Rmkgtpw6px+LMNnkvSFglAQ7FwmCb1Dz9O44w8PTt9bqJTDIvd0A7fAXnf8fUH
Q/4Izu2y73777JcQ94/wVSfKnXA7weMDMGmoRM7MnjYndCVRJZcBDvJwwCmTWHUe5sq7U541gKMt
QL9z1cFdz1Y0tQ5DRi9Q5xQJ/HuqE4t1b8g09uRiDfhaSJxIjFK8c5C5+urpS34hZVjEkd4mEd92
bHinmdmFkJb2EqOgWPvRYEK4sOEKSVXGnlTQkQg3+Yp5EX3gWLsdMIuS2/H/8CZ55CZbk72qX6Cq
zKUNHq7mQqSmczvdjt4yfobL2dkHAPXVO1IKHbX0/mEpIEW64FW1ZLVG0neD4sGXowioFLE5HNS6
3a19o9WjibP1bKfFDHaGl52tpM0JcZ42+j9nSBSLKIz26vVXkjpFjVtHp5++6EM/sY4zrEPyxK2B
O+fp/u5ONa1Sy7H9f/MCS9LslaC/9sysdOOs+Z8gOMpgzdcIlsaLCQr3K0qW1uvroEscsxJ1wvK6
79XYro4rkKRcZgRO0IgsCT144gpkMRF0mlFr+PL0YB/dHRkXixxsaDanzNzNbTTON5wHm3QSJ+CK
XHALFHxsjakiRzzN/nG2ASSQzn5zTabnyPsl8HjH4aZqKlGvhIrQrx/jHbOlTl2GqY/dMlEXk3d8
FrceTEJVvZq95Wv67Wb8yIW99COUiAgcXfsx3hH5kcQGhV6bwrbmlprvqSst924cT4XJ7pNORM92
Bjc1U6M+d8FS/z5atQJ1NJwzBnAz+3uysWwEoAOxIc/Beircjds8aeUUW5/6yIQEZxFvTAOZHjZj
//ppb7AZRMTDp427HE2x9tkHEeNhktNVZJoxJgAMn7FkuA8iCYUvpwsw2S9/nKtFIo+vrv+ygD8T
spALm8NjzoacnqMRP5nGu5BvT95RtfdP2mgvt4csRrLsIO9H0VzjfPe+7ZwF9LmNRHHERatDxeEJ
h4mZ9C+N7WyCqSa8LFXY6Ug0MJO1SWcpJ5D7MVBOVPmkQlfAy4gzj3PAzL6vwbKTpnEChIr8hBXU
/VGnHtNKOvdVg8b7Aig8zXAOJs4zLyi5Ppbcg3pxib4DXH75FxjLZYoQAmK9xGf0CsOtFqhwQ1FM
2f6l8x1vSWONamdCnTVzH0Wc485FajJEh2bdlhewx73p0lTExaTfN8hDNSrnTvBVAZ5+1Thdlv2z
CYvM3QgyktOdfSInlxtwKtGqNsbzM6GUnl9JpHzp5MzTJluMAhNhC8XeXyVD3aN+4XUkllU3mZ+Z
pSOr4WsD5kJV1LcaP8/xpPfhSSNRCjb8dTx9YXyTQTs+/ckV7pn3Akt4qEcT+ofN5kLuNgcH/yLj
81e9qGwvbQ/sWSoHLkdUzQSH/E7A1HuLZssMRKBpF51EryfNeUxeR2Z3qtge7dP2VDCJ2t48ubS5
mhMok3rwclGxwLXjNusFYLBIE95AJBQswQ8xqTn2VRHHxJ6+RBmCTNxCvNSmj7hvdKBMuLDi6fLQ
clSjHu6kIMXy/Qcqoq5cwOEgqG7AFKSEHwAPW4+ASPqkhUS5DdIKy1DKWErfQDs+6PO7GWVbm3WV
fvPqqNgvRGE+8E4pCrmflFh5R6hOhzWOvnd/ceThgBL/mc0/pyeLdRVL2uqIpfgao3E1mVGfHfsc
j3vEnCXy5KAynwwxe2JxEIsyWPiz5Qx/GrIZ4u6lO8RA7ZGRv3iwytb2lG3QX/r/34LZzcNTeMg1
RNgVI4/UUNJdofSp3iJ8lokFuNW3VL84UkbvbczpAT4pmgsMbtMbBSQ61RtdL15U17Ci/CbaMaQG
/Fzaj1+uRUTuOHZamnyC04CWAo4ifGhNUPqRPS6SBMmuL9NDoyOa+Wnf1kCtck5ZGcBAWBxkZs1N
PUs/JcqKyfGhrUq+Au0hotfJkL6LYDsM4w6ioAdyQ+iJa17rZt6rcp/JgHcHjR8D0vW9ViwZWPS5
ncFu7i4eqYLv+jFRlxpyA9UUrYofKfCfDeIlR9ItIL8HzcmlGaLuWG3v2ZB4KazWe57xajwPc1ek
j8WsR+nbRKD+K8GUST0GHMB14Bt+7LuYXW+QuPVZLq2z7h1bEBNUpZMQF86uFFR2DlajnzzVTQYJ
1oj5Kvf/DL1T5qFU5v4kYnZer1hBHsUM0hBLNKpHCVMVK9vaKzbiWoGCTLkbZmkrgD7fnKnvZx2K
r95bfSG9ADuMEdNz16tyjspX/sdsew/ecWinfZKV+qWt3UBgXTIW/YcsDRQmsCGo57NIaqNkNl8/
lnnkhgOR9JTRzqlKJj8JxJEt1NBxT4SOngClTtcf2tXeezlfYmxKl2FdcdSicesSsifytT53kUEG
zrTYnoQQQRlKXwdGLY7ND5+UnIv4tdof+YUVXRvTkL2Sdn58Qi2/08iBKYTpZdbteIeLVtB/H4ih
62zojT98st+WzXyZ7FKUtjqdQ01V2svxJoVF7yhzcksiU7GbVjjBHeTBGmzdX0o0Ue8r2k4JyOQf
1rpAOaoyMa2eRgUWcRXgdL6LupHiudruhmTDgSom3SGL9JWDoVE2fOKRwBDP1I0dnNFbj+gkTKOc
T5msnCO4Mkldv7O7BFFlNF4GmGyd5F58NkcTd4TnX9G0jTnjmJWL1q5JC+VvhP+8W7q/VGpFYrbN
7jkyksJoJZn69n/h7dzyNHyIugW8Wy3ekb6OPJpg30yASDbR8aiWz3ATkmYj01pBKhkjbh3O5VIa
8GfxvQJZNg0CbOnRwftZXijAmsB2LVkzJ22LZYJbOWHNC2pBhdmb+cjIsndluVTq1KtzmY1oRflg
/LTGRw4pJyr1JOSHmhRRCtKEdWzQJcGifCTPhUjfEPcN8Hk06pOO5cWBMlFEcdC3w6ppN5GXtz70
pEU9ITM2rS3DVG1fY1tVnu4bfLtYj7B4CU4FUwzIPSO8LC+CvxRbyGCrTNLYDZbFg7yD2bYdgq/y
VM3CrwFKVTHbMuuY/gm96lzwQX4UceCxCHEENjJG6D8mnRBrCnNocz9nwh0hQOLljQZspHSHmeVa
Apf79W6YyVJTTWWyRMn0Mc8MZTmxHMTaAeLEfz4+mAr1hBU8HFPqOmOgjs9aUuAiHlMphM9H8GHw
2SBeKGxaphL2ENZ7fDcvzSTZthL02KL4MRkcAHwrmX64A/I9AYiqipOBtQFDkRC8gH+T7vBAx4FE
iaSPsTDlBCmgZ3mcvbkWWUfU8dqm0zAaI9Wix1xmvlQSnDaoS09HEBNUFgOoKoZ/XAZvEmQgGtY9
wdQ6pChI/Gry8FnU/6hdibadntYKeOLtjLlFgDkzX1Di+HjkIU8FLve77aFtChMiUGVu1e/+0gUM
V2qEPNjmdCqslXYZ308Ncv2p76yfPHTk4CVVvkunsRYAEevVZEOXOyVkil/hJj9IKAFHTA/5NB4h
6+5otg9wjhRixUQ7s2B1SYxHX4C7lmvQSKbGPDk0s508Z0M0v5SXibuk3StLJYYiCFUVoCrgcSAj
HN6cSjTR/ujgeanbRfXeQ351gU9o8/2+a7uX2SttmIPm4RXqqPWCnRORrL2IbkvMNyZY0i4KA/ih
IULz8xUOvKmZ7R+G2w52qhR8aDyfuN+rVudvsIlW53BCHy2haLQlwYPnsIgQ/AAfnU7wllR2VTdQ
YQj9YxTCB6vN8G2+Aj/bmx1iGeuDhaUHZPfH8gcYsnXEsxwi0C4mKfR7Sm90deJHo2xQu/XBCiJZ
QsBJBw9ejp++QZEpFlEI
`protect end_protected
