��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$Rx�y�<��wA�*;�x���@�̦�W�X�fa�M-$u����n~�%���P�$��W��kYَ���P7�?UMfT��q�6�U��k�>����~�\N�(�����X�e���/6U|)�X2pF�]$h���d.���9E��WG��L�X"]�Ad����ľS���8od����e�GT?y	7�������ݵ�^��R�q^]�鍦�����s�ae���h��L��P_���ާ��YЭF���'\��68�b�[����w8�[X��V�F�0͘3����q諵�uW� �h�u\V�?@��_6G�_�*�G���B�絉�f������[�G��U&�����~�F��AׯK1�`c��[<��FY���4I� �#�G��x[X�=�Q1��`��R>(�w����R�O�?����7�,(�H\�#h(W�EH=�������yq��Ѿ��aF����:�U~m<|��.��0=�P/���4ǆ���T(���G�nze�C}L�Ȟ�-yV����Q9Sɛ~�V!6�6̐ҫA�K#s[�x3K��¨�삽.�[����I�����Fb�5l$�G{v��39``���)0 �#F��}���ognB�����%��_'�f��0�;����25|�f��߲��h3���>���<0w�1���<#�ܥYy����Z*������=���(U�~!�":�c�eۓjJ��2wW,̷m�wZ��ϓ!{ud/"�S輀YV�x�%�cՓ[N�H'*�hg=֖`xJ:�\a�	�-ȷ}�%��Lj&�K x�!	�p��5*o%S�I�������yz\|3�ہ������J5�KG��/���U�dn��*E ����d�$Sf$ӂ���8C��{=�,�-rwP�2����]���xl�,�\�_nLN��]�~+ga��U�s:�Wh�%������������h]������,7�d���<�&��Y%�F�����1��M�Rw�Y�bh�FsJ�R0�A2��'�����B�_��*=2uU�y�$�)(������;X���vt��iIg<0Xb�d�� Ԓ��zm�
��6�sG�8(Џҹ�S��5$\�2<������0T�c�x�(����"�;4,1�z֮��t�bP��.-�G����şI[�W�D���hF��9lT;k�r�K\�ۘ��P��`���֘f\6�iZ�(��Qz���7N�I�G�t��+^��f%:�qs�,z7��7��^>Jmӧ��`��쾼g'�V����Sۉ�	���M�w�+ٿ���(p�ܫ�J�p'�����Z�R�7�+���1Nrga���KI�o�����Ӂ�]���_�H$��6�����C�mk�C�:\k-����Lu��ܹ�P`\tť���'Y�#�I�����(Ֆ3�A�M���+����4�n�}��F��o�߉����i�����
83k�D��`�[F���|�5�W�'.���դ��V�]�6�$�a�d��t׊D�3����J�O	�m���a���q��#����1�b�~�8�W��-����w�0�C5�SEe�"����){ts�0�{_��^�-��טl*�F���ċ�X�	P�De���?���W�]�����$v��æ^���L���<>Q��;�O<Tn~' �Z	��?�==	���و@u9)��_}�jm����w 0��.S/�ă���ߟp���ψ#?���\А�j-���A{��F�S疍1��kI[כǃl�ND����-v)lFzo�؊�X��H����WK$~)�W��#���"E%���Ü'���F�(A]Z�������bl������0%I�j[H-K�	P:#���R��3Q�P7�ǲ�ȪM�3W4o�/��`�X�]6$W�&�OVw�7�k82O��� �H�R��Q*G~X�HD��jӳ��� Dī7����Q����1_m�d��a�m}dﰃN���a��CQ�o��*)����Z���\����������G5Qڐh�������o/��<���J!ob�� �#�{����CN ��3�>��<&@N�IzX��{���Y!�q&�H�����HJ2n��$�����CCk�k����M_��MլH����V�����u�~�3��[��w�{2]��xz}@Y
E��c"�t��9���m��lAS49�>0dg��*�7êQ��}ru3�It��1��� ���ߵ2�s�g����H~83x*txX�9��֎Ɗѹ�yt�6��e;8%��3'�U^�/���;��CK�K&����Y���zFf(n{���U��B��W����1�z��`��X�U�İ�Q���i"�]cy;�L�R�HKdrSq����e$K��I�o�I�buO�D7r��OI� (��x���X�e�\N4��68��7oң�L��ꆳ��
	%/$�����P~G�	��0��n>P&�\6뛬N�	��q�Wk@��M���>t���1ܞ����H�� |�H)���Y{yD�/�!q���^��Xi!QY���������ѻ�r��`G�b�^<5�V�(x��~~�5�[��9�R�F� RD���O`Q�Ӽ#����މ�m�"D&��[k):e�+7��>���wE���s����0�a��*鎽�N��e)�9��3hʭx���������� �m��A�v��A�ی�z�mJAE�1#�-�*3.�~���^j���䂲���#��l��Glx����x,����vk���M�!6$Bž
�݋9e�L����B�#3�#vcI!�?��5��	���PȯC��A
<���n�V��[��(r�{@*i�*Pe܍����D^�`\��Z����p���v?g���Ω���Q^ӓ��JP��g��U���vD�m����$�R�Q�10n�NXGdO������A���>�$��Ϫ���(�bn�,Ƨܒ1��v;���3E�'��,J5���-`�sd/#=�MXHBc�Q�t�'�l���=ܛ#P�NM���g��LHSn{���LGB�)��'\A>�e�#5�//f\�^� k��d�w��+첋�O7Z���^u���sAK[X��m129S�4�����K@��{ F��n��{P�WJ����%�7���a'�":2�x��.SA��垶�ٌ�xve��!�t�1w�[JP�z�P_�(FV��4P[D���a�b���C����aH���VIl:�x,�l�o�Ñ*j�Pz�������y2~�h������($�%Uc�t�m�OB)���N�m��&�ɰYi�Żv䚊TN�Wh��%ۃ���7|^
�3�ڑ����v�YhI����q�6 J3mm���bQ�q\�R�n6��J���.t>/����E�Y^�N��P�c���5�Pq��Ry�L����Z;�`NreO&<RP��|���U�3V�[����Y?e�?1�=K�t�����P�\�ٮ�X|Q�b9؝�Ⱥ[5� ɞV='S|Ql9��O��|mE0"���E����uv�f�V'�L������;��ZԼ����LQA����eќ���q����x~{���������gS�E��G�.����=E�ER�E��HPm͎o��5G槄�g�"��I�p�Q���([_Z�N7��&��'���Lq����.��%c|uw��ζs��@�+��Ϯ�6�;�NrEY�]fR
C��{�ьA�P���2�{:��*�����8~��.YEiх�Vx����l� &�`�����%g��.֘W����8�/.���������Ⱥ3� ������SH�dM�6N}s���Cφ��Fxg�]!�ȯ�����yS�R�вg�:0��p�%╮���)f<_Wc� �q��_�q��7w��1��v�Nq_pꑙW-e-�D������|8�Gv��CҢV��_O}�W��?���=W��eٝx���T�Ytm�5%�U9��C�V�on�⦓���W�Y'"UX��--\yNde�y�jL��mt8r)!�I��![�%�Y N5t	$�q�cc��%F�9���M/`u�+�)��х�/z9֭I�x�|ߤ�������Lt���� 	t��"�`A�����d��]��gJ�n}B4�=򸛏�Dx�%s�j�Є�۳5�Kχ���[�B���}�9|����o���ɀT<;�ci��M��v�6�yCC�ek�4y�L/g��K`��ݛ�>�w���`��թh�Z2_Oow��D�ka c�d;Ɵ�K����/.�Y�E,�D֤��ё�/��r���!K��G���E��2�]���п��&���r�4��$H`��Zw���r�M`rл�Y��T��:���Bm����𷔘"���>�N����`���w�R�����(�&�i�@��,�k���uNR\�H3h���_o|�ND�`m�S��� ����&So�j�Ƶ����������5�d��~��թP��xqe���x�/'@w���xޖ&�0����ތۆlb.�	yP�i7�}�N'��	Q����.���E�Ԝ�ò�z
�v��]i�!�\������7G�?�m��U�u\��x,"�R�W\���9���R��
�k�5�~�w]��t�P�