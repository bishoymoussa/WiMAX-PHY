��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$Rx�y�<��wA�*;�x���@�̦�W�X�fa�M-$u����n~�%�ArR�b���#�j��ң$��r8d
��K5�<���5����Ǐ ?��H�����e��6�j�F�K�B�e����Km�^�;R"n[����/D�}��q��eQ�J�>�5|�>�;ĺe��.a�-(�g��+Y�gO<���E��6!i�S)i���Q��2���l��K�^�%ӄ-�E�=�Z�X�t%�J��*m���X�f���)d�IEz-U�Kȵ?�I� AQ!LL@�t�S����xHq2.�L��Q����d�8��A�zmv��ƹn���eW�8佂!�y����2ڧ�
��Ҩ�O{<JǈM���%���Vɶ 틜q��a�6OZ��2	�AQ��:6��3�X��2~gztF�l��v!B��?|���<�\�᫜��Q����c.��t� �)qg�b�TT�0e�aN������9���ip�-2�^�We'T&���Dg#��r
5���]T�����:�Ô>\.֗���{�S(�H�-�,�Q��"fj}�6��N��+:�Q�V?��(����_}�O����H7�T�"�T�B�d�Z���	3�ײМ��k�uf��?r�N��;b<�9�,$+7-<V���Ci��H�����ɔ��k�:�%���`��&2�Nw���,Y��G�?�C��������a����[?�zJ�S��w8t��n�;� �Z��Hd1���0x9Н�X�7��4;!�m	�hHZv,o4J�� M���C�#�kei����QŹ�R}p�.D[\�(�>����$S�{Yàa��i[��w6�EJ�oj��&K�Pk�O��B�X�4{�%w�J.��;u��!^�:;�	1n�3��+�X,(Kn�$/���+w믦w�P5�@4T��	�&���]Y�Ѓq�`���ۤpH�卤�k�ٱDnw�n������C�(��29���t^��)vk�~�t�E]Iם��ym�EmSb����rSI��K���@��TW����(e�k	�`y|�+��]������s8k����c����;���ݦe>���9���s��ǂ-�/�xV����� ۗ�zxm6L�},��C��"I�kj7�V�2�Ξ���OLd[o���D���?��[B[�����}��\�A���{��Jɧ�~k)1)6��fۿ��I�0��s{���ǇH`�����Rl������fL,�qN�ځ`1F���/\V�%[���w9���j�W��Xe�,�=߮g�j
.O�&�Q�3S+��En�CtJ�4K�+�����E�1x?-8��%��,nThz|�=	z���kM����c�)�|4�c)RRc��!D4c���KƼ�8Uv��$��Vk��c�n��¦�L�����g�A&qNQy\��43rZ������F����e�-�~�DOeV�>j�z�w��l�:y��n@cr�-�� dg[�CW�Q	� �F�sE���D:&���aZa���|A�d��	�":�S�1�L��m��N��.��»tر�G� A�~�v@9��{q��&���5�����B��j���1��>��⍾�ޙ�z@G�^�F"�^VFX�P������E� q�o�X�h�~�6c��j��$��\9�O��ZP�����,a$�$`L��s��	�j#G-��;k(}�S~��`�8Nu*�� $f��eg�rs�k��b0�t ��аc�d�6��,�i�@�P��:\���ʱ�Y�;�D�#�owGFo���Y۱�c-��Ĝa�b�͑u���d��`�O��2!ݾ�݌ ��	��@�3;�u�%�Z��C;M�>t	�ٱu�$��;g"�����V{�㚿)���eHU�q5-� �"�H6���Q:�܇6�JZ١7۪±��|��֔���`�FH�:����u��2,0�+7=�j3|R�*v�g�nӋ�d���	�������;�;�_8�[m��fI���mQ��`m����l�$��>ң�`-fuE�`��[��v*Y='�Mc�K��}�t:"ټ+z37#d ��^�G87ِC�n��_z;���}��J7$B���)N�-@Jc�m��>����7O���Ǝ���ީ�ʴ`�"�흷z�d�˶�N`]fz�V(��)�쇅�@	0��N�ln&��vՐe+oXÏ�C�)	��2�Z�ã��O��������5�t��PNģ*�(+�}VZ1��P5u���I/�]=L�����d'px�P��&�����n�ݯ�$�%�j�ݰ������X*�^cUi4�!"`�t����It1��=&�=��2����|�{��G�ni�b��'C]iG�����!�xK~u����O��5�WPb�kh1.�5>�FY"��	l���A;��G�nzg���>=���5�t�+U$f)���}���%�r���3�dmM
JL�kSV8���U˥ a�ד�е����,��}Y_p-��O��B��S����LI�i*�gj�ϭ��68T]m��Uj^�q�b��e���Z,9	��t�H�+��M�0tH���+�u2��z+�;�7�n��\Hl��1��T���E��e����������H��*��@�@mw7l�/�Һ��7��>��aoL����8e��+l�,D��-�8=:�rn|,8"6d"��!���]/���e��n�;L�K�\�Ơ��p��}#�3G�@��̻,Rڳ ��@�Խ^��I��\�.cP��d3�{$�2�N%�$�<�3��Iʁ%Zl�^�}0�XThe�5�x��r�=���CCAC���s�j\�"K��쁚�(�|㚽d�g6+7������wct���7��E#�գ���� 6���{F��\�v�n��P��G5s���>��"��moü<��j�S�6F��^��|ì�]ٲS� Sː�� wo�� �'B䷸4j�x�,�&����൤?Ԣ��`��6���pT4NQ�Y>�yVfd��X�GUoQ*K����\nN�C:��[kݐ�GX�!�lrv�-������t����VX�Z`��4��A���t���Y���hq$D��9t(fK�4����H4���\���ԍ���G���-8�/R~�ʯk\��Q�yf�%]���e�`x+J�� �i��A��-*�����u$ش�����(xG���.�Ӿ��7K�B�O���t�e��b+Ɯ���9��2&xR�I�S+u�L�O%��B�<�F�kQ	��A�h��v.9����2y?la�|Z�lb��z&J�$[��}i���?n��ꗡ�(ԯ�+���������F��z`��{�,�Ӣ�(<_kQ��D-d?�U���<�C(���I2�!�0"nt� &|����<��'~f��d$5p��[q&^�cf�^�%�0w������	�����$�(�ِ�ʹ�Ek�Z۫�b�!�����t7�r��X���O��g+�dތ���Fpp�����3)�mM�FJ:	���
	\���f�Y"�v2�f��a0o�P����n^jv�ѿF����������q���þ�ˉS	g���׭��G�߽;_���:�pق�.�R�{!no�c/�y��#+זU��5�k��hL��	D��){��*\����{N=&_��V;�Ã_,0�Jou����^�yg^��f�FI�b���;x`du!�|�ս���A~�O�T�t��	ڛƥI�wI�?��ޣ��L�,^6��U=��������%��b.�T'pp�'׌��<��+��e�}3��i��[y��W��P�si󄧿]�o5ݹ~W"��)�by&�O!��\���5�],j5=��-+	s`mS�����m���L޲���w�^+[y�	D���f��i�+Ef�}	聤d.Kbn ��/8�:?(^ i�i�Km��!��8(GoUr�1:�����h#k�r�]��:{݌�7;�9�YG�Z��5u��tZ��V��(F���g����ο��8���%*�ߜ V����A��W=$��-Tu(�!/��q9B��Jw�f�E���]>�ͺ@�-�"�����A�n��Siش��fs�����-�}~YI�ˤ=������W�n�I��c�
Gb0�xJ���Tvzb*c��X2(����`�vU��ԑۖ<��Е����!����b_b	x��zCi�/�Q�Aoz�&�O��$�:T�t����J���v{`�jw�;58���t9]��7gaV��J��*�"�i"t&������L�>H����@��{�Vg��C;�@���Ak>*V%�p*�0���K%0����o����r�D���#��e����
G�W��z�%e!�R������z��Q�ś�4���	�^�t�hY&�NAd���`�(	`2�{z�-ȧ�����'��� �ӄ��Ӫ�ر���˔"A}K	��zb����K���8��s� Nˣ#�������U��ֶe�4X����l���2�K�vWOE��3�E��ȂX+�{R3hw�;�'*�1�@n�s�I׹F �#���Q5�ƺ�f�yGrd���ۧE@�cx��i�*����-�C�l�uUv)2%N��Fn�]c���Zj�J�c�U�j��<�id�mV��("�x�ɱȅ�#�}0�FO>�T��[@pbI%W�	'�ފ� x�#��U�n�d���`����_�xugFA�% ���t:ŀX��`p`�$A/J��]��Gª���qw_+�j��w���^Q./��w4;�C�$�H�[�z����D�]�¶"%-���&tm��U��Q�V���H
݃��������uA[�T����׳?�7sZU5���W�1�Ք�ײ��ȾJK���YE#���I�]�\���O�c}�U"�_t�z�ZH�y���rm v�n��s�R��e�����q66X_�V75�U?f�ͤ@�%�#����!�����=��%9�	���eO�������ڷE���+��pF�$�h��p�2'�h+`����|:Ȟ��xq��$��PB -��7�Q�o�#_�C�A)Ahs�d26NPX�_��Y���F^��v�ƺE_�ù���8襛���[�5��M�T�h����=$u��x��z�~
�\�j��	d��-ɣ�p��F3�+f����3��M�����	餖�a�����;�	`���24�8�4̭	<�}�4'Vdp �|�Yi*˘�>~����|�K�6`�I�48��e5�Ø&�׎!#F�+GsI<9'{��v��%Tߓ���8'�ǭ��g{|�"^<f�=4��� e���<�D��S���|�3�v�@�U}u����Rd�yd� Y�|��C�])>f������p?}�B�f
��ѿ%�Mˎ����*xU�%Q��k�h޿xİAb�@A�f���N)��Ό�󩳝�{a��}fQe��@D�>�k�ĥ�]�l���7?��S�	�w\�%��V4�*�W1`��#i�X$7֢���|5^$�_���5�+OBZrk>���f�������n���Rl�9��XlW��x�Y6��@A�����v���It�j"�PJkሆ�4zCm�{�u>�������|��v�)�a\�e��C'T0UAsm���Ծ�E��-N��%Ҡ�f�N{��ViuE�T����jY�{�4<�OMFHϛָQ��"�6D��IH����8/]�ڝ�C�IJO����B�;�5��Ĉ%a��h P��[�<���~Ÿ�%M?H8QW"nQ�8D�,->A�g�����9��əߋ����4ۤ���4(-Yч��T�0a�;��>�����,�6pI�T�d0;]���]�ҽ��_לi�}!@�m��-T�}���nCFΏ��]��.`t�I�HO�7�v��5�Co�����ܳ�~�����jL�����[yQ"6�2��3�#R�Ĳ�S��`Zī����)�>70-�LK�!z�_���Ja���u�"���e�b�I���s����t���uH��}�Q���f�\N��9�~l�4r���w \���?�Ŕ ya�r0�O6��k˧����0ޢ :/�	��A�%�B�3��iC�YB��8.l�u1��'��Uǫ�!��c�'W~�/uU��Z=���]qj��-i�>�uմ��y���_2N4����#�dW��b�ճ������-�*�#Q��ݕ���ÔiU>�c?P�ցx;��U�_�ݑ��#b��շ�X$5Kg�I�]�\rt��	u�toQ��
�`d�K���92g:���2f��
�4����N�W���%Vas����I�S,l>�nC*��}�J��t)��Je�v�Y�z���ǃ2~\���O��p7�ǁ%eAL��!�Dz-O�<5�YX�0k%�q����-�F�b�a�T���o��d�"����"�!��}inK ���^�����xF�Ig������^sU}��*B���z)�;��9:]������>neɀ�wsZC��G�S�d�Z`��\`з�?g�> �@�Uٿ�P�SP�u ܣG,J�-d��6A�S��x �!�3�ġ��'k���XA[�}�G�g,Y��W���>���IC�8��*X���ŵ&mw<�R��%�����(�y�)�~)\�;���@��)�&�U2�D������"��d}�X�B�I)uGO��09���)C�J.��Q=c��:Ս��\�=5E"�|fĐ^���Y�f�]ą��Y'g(�� 8{�TC���k�4�,�+��H�Y�s�B3��)��d9EX�����] �H��0B�<��֪�4�W�D���fő�t���w�NmJ�5BX��h�A����5��:�;�֞T��d��.���$�g3g�0���^�2��&�8�6�ў�-����8<��h�����d'�)����&��P7��L�\���d��P��P��D�������i�l)��O(a�������
�5�-������0���E�LC�!�'+0�6Dڧ�FŖ��*�,>a���[��5Qx*&��ɷ��`h ��0�s������7�x�0�R����K�D(��^;a�ɺ;�s��X*���lϕ�	��O�R��b'Z8��m���WJlP����L��/fB�����Ś��_�1�����lU��x �5&#�q���eF^�$�MQ����F��j`��%g�FB���XԤ�G�3�R��"=��zS��,&�}8���B;Ⱦ���0�#W���t`��ccۑ��Ȏ���F3�<:��%M3O�q½�+KR4�e��ߧ)?��U��[Ȗ�_�!^���YIS�Nv�hf"��z�(
���`�&���6��s�cI�v�ҶV��q� D�����]l�������!`�q��g%t��Z����E�Ѩi�i,?�� '�Q>>�(��H�z�)*u���m����M�x�������0��5���h�`�{�ԇ;�r���@Xn���p�륈S�NY�$(J���(5�X����_�v�>Nn��Z��uA�hd�~����ފ`�j�5%{19�q-=���sX���y9�~����d����֚��}S{��}rhz�Xj�!�Z�V���;���O>���$]�Ê���B5��X�J�|�	v�V�=j��Y����^#���.�gZ��
9C;��_�����`�'���|���%��#A/p:7���̢�EJ�b� �����UHz$��H��/[��I�m�#@#�CN���H����yص�v��Ck�:V9���ߣ�`�b�c��o�J�v�^�M<oVs]���B�'w=�Z���>Y�}�#���(y�vDh�X�����I����BCA:i�܋��nY�<��;p�,Fp|�j�H`U�͹�b'Q*�?WJ��>p�����`� 8���P�,�I�)�!�kk�B�(6Ksv��^o�X\����մ ���j]Doz�ȍ)֝��x�v0����ra�G,_`m4��>��2�e����.o7�P;�86�kYG9�Eۤ�72�Z ڼ�s�wK�?���'=ª�rC�ϙ���p��O��Twh�=��ڹ�B�IN��.#�E�R���w(_��<<a�Vf_��
}re�;<��h�F6$gM��h����?����}�;�����jS	�9H�L!O� LG+�;0@�YQ��}g��C���|n��������>�J�d�����_GhR�5d��a��L�F�i����^�����J��h�v2� �2�A���r�dq�$��K�C~��P�� ��Y�s#�B�$+�܉��d+̦S'�5�$ג���Q������{�4]UkL��o����Px2z��/�}x���r0|�|��.�׻c4k�n�ؠa�֪6�M���*�G5�%
� hvХ��X�aY� D-L��z�0�7��^L������P��{ ��R��4U���9%g����L^� �~-4�1da��4ή���@��p�
vJ����B���Zk[��=jNNڧ!����������/�8�s���K�{�(!N;�P�f�ށ��YR_f�M��Jyj��]@��8g
���p��������d3��s*$~�5��K�r��L�Z/�`8���r�;�%�\r������C���c�|�c���<ܸ=���`�Ԫ(�\t��S
Y�N�-��'21�2�0��d�w!� 5�C�}������#'"$t�[�䒦����=����� +�J1cɜ񍧜r�D&��Z:~�Gs��{�m0�w�I���Pp{�Q[c?���%!�ۙ~6i��.(q�n5B����;��o�����z���o.��zOvM�w�:I����
^>A.�|k�+!�l������u -�Da��r\�ن�'.9�L	�����r\K!��C�뼺TE�S�x�^�k\lڽ��q��E,(y�m�3�G}z�����x{G8�JJ0��,���,�Ȃ@�Bݿ����$҄���wҪ�#��-R�J7�@_�D���;9�����7��T����B���@X����h�f-Xa�f=�����7�?�yUF���LZ��g��KF�R��P���;�
 ��SԄozW��`����yAV��B$�l��;�(u�K����L��Œ�_#�x���ȷ�����o��%Ι�@�(0�� �v&�n6���ą�he���tDdY.��|���;�4�i-�Aڈ����ny
����XzL��EȇD~F����kZ�)QZ�XK�~'���^�̗��ɋ0�`�1����<y��6�c�mH%܌��(�'�5�e[�1׮%��c��ّ�ĕՙ(�����B�C�����e�!vz��VF\RQ�����x��࿑(�c���<����0c%"�񁒥��ˤ��?}�a���_ڑT��\/$:�^�=]�&^�e�����,�t��"1)�	�s�اv�ݞt*�ڞ�le��mr���y�C25����-�O�0���M'1g�>�1�6�̰B�4&�y��n{]R`u�E��ϛ�B�At�,O��}����Sq4���5JH; ތ�G�d&��~��a���=�Пhc��r�Īq
- ����M��'@ָ?�����le�ز;P�5ۜI%za!�l���0?��	�MaG�̝;��-4�\�57t�_��Ә֬���؎^X�!�N�g���� v����;�(?86�ȸ'Ŀ#��J��-��B�q4�$��)����2�տZ@��r;a�Yvi�կT7��]z�|٦���X�H�[6�t�/5���#���`sչ�ca_�x��:!l�(˙�]
x6ha��c�Q?^FM�z�G`�*w@�9� ^?���`�(l!���6���F�X�s��3^���|���w��Gf��1�� �ۋo�3 ����I�A?�g5�`��Ԡ�h��ƅa�P[;���c�PG�����Du��p��X�`6n��1���|s��Oǟ�8���T�Id�==��6N%P��Z��*^2I�g`�1"���M���T���^z�$fZѹ"ޗ�4��1)�,�*.$J��j?^�6k>\�r��Z����g,t���˭
��"t=M�(Fs�>�����iw_���$��C�9}�6B�|��!� e�����
U�eX(�E�ߞ�����]�y_7���e̤&�P�w˕9�_\�}�L;�����4mU������6
٤w5��pI��@�)a{O�O���0��ѱr$�ҋ�'�N�!�<�߮��~����L��ѽ~֡q5f�G@hfS��*�"'���0��s�y� �Ǖm箒����WI����P)�)t�_�-q�����Ms<gn���ZC�"�Z��$V��1��X�kb��V5���y�EӅ�[�-����v`N᭷����pt�q�A.�3������^x���1�)� �'�
+ٶ
�J�6�U
�l�5�lv0{J��B�Kv,;l=�|J|)��,[�>])�0?���͵���e�(��g��*τn73$��~^V���x~S!=H7q�@:�)+"��m� ��[Q$C�b�g�~%Xў���Ɖ�i)̠��@��Z�A�&s� �E�vС*~B�H@���*˼[$k��\�f���?�9�P�A���yQ+�}��e=~&C��]l�I��G)�y-�L���FE�����:�#T o-���i)Q�c> �K��h;��+�ڐ���u?��1rc�u4#TŎ�\3�]���T�f���V�[+��205�z�no��7������������׏o��%�Å�[N$^���W�m�f3mY�K�k@s�l�ӄ[mo�4	�UΥZ��]��-�k�w ��7>��ӟ��,�?7����z�\�����#*��z��L�v��w��$ex}p>� }�?��I֢����6چ��D�A-�����m�]s*�\��X9��Ů���p7�&=Hh�͈ô�<I���d��qj�k!{[w�~sD��Q/�L1�ư���u����jmOm���ޅs��ƴ�;6�Ď�x�R>wU��5�c	� gúʞ7��G�%"ΆA�7H�� Esj��<��#E�6KU��� H���{J���a����$��b�����3���,?�dU������,��r�05�;�c�B�����a�v�_o�N��7��J��#ļT9� �C3�o���ztof���� da��ʹ�����		�kO�(VY�S�%U�-��v"	��k�D5���4x��lĊ��$�]��DB˷^���zx:W�1@���Y�
��	 �t�	�W�����c��T4^[�}���f�E��89�1@c�yc�����6����ڽ����~��⎬lĦcP���X.�;#����Qf�%�1妁I�Q䅅�ME'�������yy�J]�8J���w&��;#h�"����Gg��C�~����[��1�;�X���8=�?>�j��� B��t��=<Y�FZ�����N�e��0i ��t��3���캶�L�zS�R���Z��YF�W1s����F�ͥjW�_�H�/��j��|��������c�@eN�F���o]'�\���	,1�W�օt$:�!*���h�(�e�z�|y
��#[k��a���3��Y�FHT\=L�O�mv�z������4X)մ�J�t(>��.� F>i��R�8p1�K����4��,@r/@c o���K�����h�G�вU����1I�+&Q�����ƤwD�e"�Ju�n�$a�`�~E8r*w
��^L?b#2I^����D/4��k<�����:I�Q%�@��� �|v|�����DqOzŊa�㯵wUG��3�T���n���[�t87���	ͺ�����/�-����Ya�!���!�'�{��.�ဲ�^����\\i�	g��'�u6(�b���n��`%�W-$���x�=h���s�^�mQ�Ba���s��D�K,ˤp=��Q�*�
P+B���b=�h�a+�b�Hd�Q�hN�=�p�	��k��;v�׻��ot�Y�؎�0����d\ə�(Kn�#ܷZ`&i܌_N��u�s{�%�2�;����Q�.�<�bRA�d�ߢ=u��fJhNSL-U���d�i��egD~x=�ƪ���B�%F����@��e��0�t����pj���0��L�]Z8.��BS����R��=Z!�WI֣	|�M\�x~[jF������x���W��jU�������)uc�J�h<���0	���*"d��\ Y�N�v�k�w��+�Vl�R���u߷R�7`bp��I�U{��t>���g�*i�~���2񹊌�q�GƽfID���5�}Q� sw���{��#�A��e�Y4f�u�
�$���%e�
`���p�ĘnD##���@�T۰��1�N̟ro3)�.̭�3v�N��=�*�o�v����~�]�U�@�fQ�-�j��B:+����Cti�<T󁜰D�(;W��K�[���7���l�Ȇh1�G.AЖN�>ie@k���&�fB �j%6�?��e�(�X�&�.�Jy�G���������c?z���o���^j�l�3�<��s�Ϸ��#�O;!��I-;{@��_�rf���0�`�;w�|㒑ET��s��JbI�-�;�b�f~|l�X�@�	,��.B�}�s������C�O��j��NC�Fċ�G�4��+�wX�%�����P�Z:�M5UӚ� ������%[������v�|��e�i.�t�r�gw�C�D�Y ���ڠ�iyk�������Vr�6\o�VlcׄG�Y���Qv�Rڲ�5����O_+�쀟�tro+鉍�Tri�i��?Ǉ&��Mwn�~{6�F�ZD��~�GD!�o�	�����۠��Gv�M�0i񽿫�W���o<��-�IU�g���%�:�T�-/�<�� 0��G��[a���"y��	|�}J1ʽ��M�:��p�R~��_���:��]��U���ѭ׎#3�3��+�C�#W�U�蠙��p��o��Ŗ���:⍔w��ᠼ�8��1r�L��f��*�m0p�ۡ�!�5��c�I�� 55��� FV���^]?�7AI� ɶKCj}n]�T���0�
m�f�
����4�-�ڧ�gM�Ux8i+]����W��OU�x'�E�ch�Mi"����/�Σ@˳���pz	�5Y̸^GO��(���Ȑ�,Vc^9�l�R��J��y�O��d�'��!�&��dO5�!���'+���>������٩_]�!�	��LH<�SțO�Mo��R��ŐL�A�u\D��"T^h�7/^hT�A�B�Y�`Q��&͊p�lrϬv�bu��hb`��)�\ѿ2���R�d�v�/��4��YvL|ҽ2
n%흙|Z�ܛ;����UP%��D%�=z��m&�L��p�bAHBu�}��n��0��20�A���}�"��s�t/�a�j��%�Je.9E/�g�@
����p툪��> �5�7�������S+�9����uc� ��J�!�<�c��(m�f�ۧE*��<v� E��n�C��Z�Q��-:������g�/1I!u�K��#B[P�d|%I����1DL�����k=����&fVr����*���D�f//�����۬��+}��As��%ŗ}1j�;��K�M�&���qV�f8K��[Ւpj���SF��r��0�%7�����nJ�-���ˬ�C�xC��1z�\N�f-3L;lq�	�\\2���Ip���Y�־�ݳ�/��&X��I� 7����a\0�g��!� ��O?���[�NQIz=-��EIمj,g�1�B�����~5?}���s��������o0���W���[�J���~�~��ݦ�"�`;1�&?K{�ž�J_���"�˃�ޑ�vu���K�c���LJ�6�����vz��BP���͟�S{�i�֭q\Y��� �Ԑ���v� Z�F���_���(.t��}��B�jy"x�ݴ��k1,t'.����Rz�ʯ�q,k+�">���.y�Zˉ��3����HX�ݘ2���:4�V���A�p�0{zy��լ3;��\+�Q�v���?���M\NB<�
��2��9	F*�hܕ6�|�)�'�X-��y�s�;}-;s�<��k��{j<]�84��v�����Lbg��G�m��X���3��՚�Ke�D�핀0���S�J�o��1u#`jn�L,f�?���]���Ʌ%|}A�lA�ɏ>mt�R������*��3�$$�{������d6
1>��f���|T�p�V0r=��{�p�Q�������p!n�r��J%��w��K���(����R�O��� �-b�=�tR�c
}��k�F-"m��>Y�(	����^����AC��������,��6�%kᆃ���9�@>#�"8�A�h����z;�a���R
x�XWv�aP��=�]��n�Y˴�ŋ7j2����,���蟥��?N��H��@'Ic3iN_�^����
tEp.p�Z��'At��Z���)ĬHN��^��P��:#�M�i���n+����9,uz���tt����FHө��B�#�;����ґ��x*��.�*x_ ��6�z�y����]�[����1����B!�r�#�*��	;:�nS;�a�ސ	X_1b�3�
QI���|�#�+�=�HU�$�^���fr�$	7x�cN���s�<Mh��_n���@u��C��!^��Q�$���~F*hcț��w%z�v�]����	r�
���y
��K�5�M�޽KyR�#Lv�T_�X�@b��b���ڼ���ν����C ޮ��s?�\ԑ����6n�$-!"Ƃ{m�f�B�I��6FjQS���U��_��(� ��Tz����_�>n��ݚ�M�)c�һ��e�g�ÊK�S-�t����|b#�i�����	��jV!t���oa�F;s<�J��J~��2��U5��<�t��%�����.��@�PI����Yk,��P��@����,�k����\(R��/:�3�?z!���H��Q���7�֓z�x[�t
�w#2��'(�/C����r̗��B%�%߆/�(��N��#U*9W��[2"I�2-���s �\��A��z>kˠe�」��X������ �,o���ts^^�N�?�zf�Y�M"»G�Y{r��U^� Z��^ ���J.I���-�N��\<a���6@>�CL���أ� #�ƭ��c�,����mж��0�)��YX��r�	!��]�� �DJ�Jo��22�IB�#�t��e֥`6�}pm}dkA����A0L|-~E�N�K\�Z���hN<�g�����bܠ[�=��Qa�{B��/�y#݄�q؅��F�&ԅ��)oB��ϖ�9��.�� v�C�ԑ���,�N�h:�F] 9F*�7kT-��i}O�c�߂@��^B���AU��$������/L*���)A}�Ll��*����HHtB�m���f`��3�6��1+��H����K���.�Y�����_%��~~�iM�NX�dŶ�Nn�q-c�s�c7�U=���}5�w԰ᖍ���t��Xp�=c]�ތ�C�-)qeHRQ������X�=% }Or[E��}���ȡ�L��y߈�;�̂3&k��op#CT ��N�gL���i@��{�I�ǹh$X��*��
��V+���}7�`ŀ1�Wg2��[��Ρ{�bTetP� ��h�sS�J�v��ΫF֚���+�(���K��E݄�l���N��X0>�@���#��+}�Nق���P�Y;�v�����p3	-N~�e�qvI2E����6�x���9^�0�ݢ��p��H��ΟUh�e����E�Y��Լ̅��k�O��y���A^�v	����f�l��&�\'X��NK�((���(<��ކ�L2O�l�tX�K�8�d��v����}rq/��y�􅔚��˟�F�� �a�n�BA��B��?	����_�Aq�� ԶY�9����H���6�|�+��0��D$!�z�KP��L�v���Ad5����F�� �*A�P�_���P���s�o2��8�^�-�I�u�cy�G�h��b�w��Hmz��8�s7wT �$�ܚlm;B)8(YM���H���1����~��b(/%��&�d0Ɯ��1���&���JG�Z�ի�������~�ԃ;]�v���3=�)Lc.��%G��h{�X�c�B�!E��"i)��'���w�Q�m���V���_�D�Nnx�؉���g����-��k,7�!���h��x,��QǾ����=��&{$�L���}�����*��m~ Z�=�!��ӺH�[l�JǺ���z���Z��pX@ ��� �X��� ^���ɤ��q��s�Z�x�Eγ�~x��������eD�M� ���B7m�`�Ë=,�,&H�N�E��0����sf���s"3qr=��ߙ���jb�����S8���UN�&%�����7[mC|UI��$+�F	�;��E�+���(�*}ISP�[4֩����H-�	)r��k�k����J�<�<�<1bHG�a�֣Fy�"4��2L2&E�6���߹𦲱��Q���Ę���<p�]�햝�Q�/�A�7�	29�4��9�F�ʬ	��q������~�x��s��[c7x1��0̟��Ar;�`��P�����s	A�U���11+�'^�:��U���U9E�N PCA��6҂퀌���L�uY�G��~ *��\�+�4��aI�(��CWx�{�-�[�2>ˮ�&�<5<�fb{'C�l�9G�ΚВPkOV|@���؟~/2� }p7R?����`��3����\[w3s����U�]�wJ������Q\K4���oz� ��l�enP�!>���OV��f�&UG`�.�������q��f�wy�T���2���W~dEO�v�B*� ����js"0(��E�w*� �f1��� U�ό�Ĩ�vu���`ā`��:���܄��E��AL4���*�D��W%>�hq������d�D����:�E���=d���	S���H(s�&�5��E�Vn���������X�y�6�fv��T֨����]s2��U����I&8ݙ����������R�q�h`�`̯����Un�;�ǈ#q�A�ˈ�� �5#Ҹ�,�����LUԍ����«q2�r=`TFˠ�u��. �%e�#��VVcOD �'H��%���1!:�ƀC�g��n�;2�$���0z���ܯ 4���g�c�u�B?��C�!��i�':oo��ܟ,�֛fOl��=�"]�A�%�[wiA�>ځ/�X 鿝8Jg"�cްԾ��y��q�}�����l��)m 5~C�}q�.��XZ�l�P���Y�wL���`7�@(I��y����(�\�l�?�&=.T3���䐑���"�3p����L1��IkF)����h� '�](�r?g<=���vg̩�J|����-�$zd֖����F0�".��`;��k,
(�8F�[ZX.�XS���Θ�28T��w6?)�vy'xV�/ed�W�����Y����]��0�*���{�G��ƴ��~6O�zb�H�/���xp��8�,ˆ�r���U��d7�Ĭ"���y�����)5�kY�-����L�6�9�ι�����^��G#I�%�ѩUUZ�n٦<��iH�8	Wutyu���A��-��4 �)�['-���1��1<\W*��gf�Y�I����oc��قt��/�ݘP�E�;�5�w�ԏ��c�3%����M@�
-�ozlc�4�==�bp=(ke�3'�:�J�D��t_�5c"�N�y�,��c�̕�L�U]x|�MЩ�t�Z�r��'�sS��
�����͔H���D�z�튣���������e�-}^���Cz���9�@5��%�9E��R��'�_B,ǐ�4w�3������e������J�ѽj�
�h`i%Vb[�$r������v����"hA�e�Y�h�L-�5;��IY�Ɲ�bo��R|R́��N*�e�)�8����g?L�tz�����l��K�H)��������0��5��@��$�/諲�6�f��,+����iR���uX~F�3���KW8R3'V��Wh�۟����&�"��U�kg�ƩLG?���p�"��E"D��$LTn�Io�[>%���yF���ⶑ:7�13�o��)�d" �\��T���Z1�V� �P6J ^s}��W���Q��0��m�W���.X"����)b��I��JK�4�TX��,�veQau�(��
��'v��X�p\�h��X�#��D���Z�X���L3���v�a��kFsD�-dE#���|4�s7�^o(����������wG(�0�c�m�fL�2^��-�w�mS܆V�At��7�M�h���'t1�����P����Ttm9��t<��	�'�BQJ'<��Z&[��7(��l����I�#$+��ɀW?���(��C�� �:\JNL�Ւ�:_�;�^��9�U��D	����PK��z��1���L�BK�y^�y$yK>��4� y��eOH�&L���2�o֞ڭ�:,ĵU�6�l�aimDmx���,��x}��L��>���c�F�b0+ �TþГ�2Qj���k��OЖ���Veˎ�t��l��	&�`V7�ؼ=��}��v�k�p�؏�"
�9>qsr4C��󠙒sn�I��=2s�*F�Q��~�:�c�J��CR.�\��=:V����(�_��n��<�H��rJ�X���}�n�i� 5�/�<fy�C�9JB�"F9����	�q�Y�P��q}�avKI�C�mn�D��CR��sU䭹"W���i�'%K4>�H!�	*�.^[6�dF@9��a�T��ck	����2��v������G�o�- R!�>��Qb���}c��l�f��L���1�!f�<b�B���;���9�IzDX|�1�.��OIs��wN�\9o��3�(]iA��z"h��.��2h˼������L�LB��ܬ�:�B��[D�	o'�a��Y`O�	o��Tİ}ly^�ŋdh�7��C#:�����Ӟ*��]��8��>����j�zt�-�\B�@���w����OX�%�O(y�H*&7|複v09�}�Y�ne�F�$�{�S���&����?��^ȭ�(�rL�k9@h��-b�t?�X�"���3�˵����@i��$)�,`�q�`.�'U0r�?0)92k���o[Ck�ys�/��)�OTv�n��x���y�_�l-ڙ��[�=
a�S��d�o��$
�2����Rߚ��U��J^f}[o*wKoSR)\�=������~���L}��0��#lp$8O��)�||��Zhv������A�j���8���:��?t�m_w�&� *2��N��0@Ē����a�Mm&��^f+��*�^�J-����s�X/Og�3���bAP��u*'���/$U�۽u����E�v�@w������u�kZ�s�x�'`EZH��m��V�!.>RR�jIG*4"��R��E{4&������.�p)��ҹ�h�B�t�w��֏<����̀'��<���� BH>�Z�zYWv5��$��׋Lf>nv��r�?�@����&V,Kh ���\l�-�$>�M��gz�a��Vzn@ؑ��X]L�� ӚhR���۩�a|�f��r�uF���ٶ���|����9�E�i��OD��X�yT(&�b�QOA6:>�C��_ڏ�;m]�h�����1��A�s���6�D��^�Cv>E��4xƶ���^�k�i�ISp�k�`����4���^�S��
�SxS�����w�1E��+��$tC��=0� SD�tj�`sDR�?8�G4�\��@h�8孉Xrb��r�?R�xܹ�jL�<dAN?'����c�}^)k�q8�����K��N������լ�_x59!T`���Sa��������݁�b��2�-���rז,tY� +*#�Ю�zW��놬�/�a�[�U�r��Q ��U�Ԣ��b3��d~�����ך��U{�p]��ʶ{s	sb�ۻ2l���<&��p�lV�V����L�C��L�������K��fǑ�%S� ��[@(��gpRY�Z���Dx�9��Cd�F�\�H#�(��kN*l���C���)y����4
m�4G�|#<Ti������o��a�u��(�Xs�h�g�)4��yq\�I���sV
f�rHP�)Q�ϵcU-x�`!��4�M��q�ؖ�����a) �8��_�M�Lci�7���rm7z8�������}p���ɕf�9t}~x���=�P�i�A�(_����	�v�1v�n��띺�d�R��j�/ig�t�#�������H� 41=��J�㲕[��C��0d�cX��Oe����-�!�5����� �*o�+���F���7�G�����fҎ�8��;.�%�(^D~\x��
��Έ�M&���q����8��� ���S���b��@0�	c�J���J5g+E����	�Zs�#�	�ڶ��f���6m;S����i���\a-2TrZá���|Ԟ�I����R����n9�[��;u���k��E�;x�����8��¦hʋ-{�e����y(�{/�ׇ8�`����TD��?+�Z�m������Q���tT��-�"fd���<L=]hd(����k0l!�P�ME��4<a��@jW��k�xFr�УM'�[�U�Ui����_I�������'�|�H��!�}b�rQp�U�FXoط(�hֱ�+�=����1�
I�4�S��۟�m�>���'n��۪�\y�?���G��L�x��=7{�-F:<C�M�њƻ�X���B5���.��&��)����2X�=���y�,ׯj$.�!�0�����Z57�V7r���\�g��XS�Vl.$�P�`C6�47�w*�'ɫ(�(�~6�2$\��lQNv�i[K��r������"-�b�Y�I��	=t����wp��p%�D�Z�����Z����5���"��.f⍊�[��b��2��\�~�㪫v��[K�G�Ţ����Ń)U����x+f����,��wͪvϦl8�0g��:���rĒN!�ܵ&���t-���*y&ӀÕ�H�`Y��rT�8śX����!S����8F������[��A�w8x��A��*
&�՞16�5H�UK� y.�7-��U���$��Ў2���Ɵ� 
i��sT2=���v�T�eaW|ka4/�L%�2���P/�FDR�Q�?�p���[��0�n��Jf��3a	:��,��Fb�F���cp�������$��Kԕ_u݊�"b��i
�^1l�W� �:�|D�[/=SDN[B��c����a�x)��c0��z�P�f�Nlb���\���6-�5b��� c��Ay��k�-��d�|��*$�6��Z��x�ܢ�"�a�_ P���:�}Y���x�f�.8��L�D����7��֢~,��ך���t��ߣ�xyD���;6����<�OLE{��k��D>�-\��)2������CN+L��/��֔��yI�ؔi��,�G�1.wK�(:R�"���|�ۀ�� ����WX*7>�j��:4��'�n`�_�4J���]X�֥yBz��j���~ yAZ�,���&����4��a���H'v�o� �̛gm��qx_���Ʀ��c�%�p3P+f�	Q�7���6���<Ղ����)Ѹ*{��"��s[��x�8��\���+e�:=z�
:ȢJ,\�C$ݡ�J�r��\�fF�� ��^�w�$�������=�N����^�&��+�
)H�#do/�uy�6z���.F�; CaQ�D9㪨��G �B^�c�>����Gt�]���q2�t�Yg9�;�5F'u��ǅ�[�G�2G�dA�qW&��/����1�̛�!��R��S�8+��S�)͓-i���H���C���w������r��Z|�w�K��G��n�ϻ�A���;�y����2�����7�,I��w��7��R،J[
�CVC�0@�p���ss��"f���=���NC�tdB\¿'Ƿ*������=�s��«�/����ށ�4^Vy�����|LK;zHGH��M���|)��{)��4)�ܒ	,I������
ٔY&uB�Z�t����B
N��B.u'�z%Y˼�
�o�s����D{R,��m^�(CI~��
 �wa;���|6\��ec�Sx���a�wM���~/e�SF�ᛇ��5,��5���0�%iu#[O�-����cI�@F弐�nD֮����B���A��nBo5�*x�Q�[���5��>|?L��@h��!����N%0|�־�����d��-�z@��
y�a.�hU8���w�p0}�sچz𪫁�R��|a\�Yl.�݌5󒯇�>����i���M��U�ݔ�d���9�Yu^2��h����Sw���cd+��=8���� ��vʂpT����Ѭ��0�f�B��:���1��䫞����S	�y��Yp��q��h�k�����p��ΕC텟��C�4[$O/֘��w+�Ѱ�{
��G5l�챀�gba�YeDfR�H��uj��Kdb�|�,6��Kѱ��
5:�=`�=\�ff��8����H��>Za�;0��f�Q!�[��Sx�$y���]���< ��9�S��j��7^h��c���$L1����ܱ����de���a���gi�x��	���>~SϺ�O��jq��p�y���G��M���!lSy��k
�J��� 5V�~�"]G�p¡��<�IO���!�(Ll2����cqS,�Q�,;�	��7%n�ʶ�P�+��%��������)t���k�q�y��F��H�U��Y�/Sz.���-w_�V"���X��!d�2�q���̎,��r���^J�����Ŏ��'Xs8}A�_u�.E�u#$��[��/�D�������z���l�P9��pL�����v�(�`7�څ���@�X���$5U�Ț#i�ZK)�O�Q7����5U5�*��<��U6�D��.�'*3��g��n�?SQ���:�p�X0 ��g�c��3���E�4u]Y
�M'y8����`"�B�O0'
��_��1*�уF��R	����x��s>5��)�Q�>n.�8*��sj������E��e ��Api�1�}&h�,+�ݝK���2��mD�a��-���Kh4r��K����#(�+��q�~�v�<y����;5�;;��aھ� �w����L�s�Q3�f�!WeΘb���F�h[����^O�z%T�v�NI�:�CP�2(Ɂ�RU�x��n��%ӹ޶�.�����l�D��ұf�]��.|�ɣ��� .��	�p���e�O�i�9o�l��}D\��7����	���w�¸ e��(�B�C`�G{����&�+��adT��w�uAG���U��ʠ[���?��cv`ܳ ���Y�o�� 1n���wM�%.��հ|{j��vv��������ٟlpb��'P�`9}M��=�P�	.�wt��Fi:8_Ct�۽WZ��u�sUxM�wU��+���	�D26"�#�S�lģ��xԍ����@���p�X���_Ū[#d����CU�㖉8oI1��,�v��$K�H�HD��Bl�0>-��:5�Gx�f�	.ꜚ3�Mxv<��lюO��2���[�� W�f0���[(ꙟ� ��j��ehwKXT��㆒���a�b�~.�X����G_s`O3z��=��*�8ΚT~v�X�#�1/���t<!z���n̚*���\�Rf�&F	�I�v�X>`.����aH����5)��ǤX? ���p�RJX�ݾbG��}rN�����f3�+1���P��x�Q������C.8fsW�i�"�m�"�<���$p�����F���-���@ͭ��@j<JR����I�m��Hw�P)b!�af��(�'�~�y̳g޹��7=�����4��c-������
լ�ft�gOof� jo�޼%M��ƣX�X���l��J�u��9��˰ ��F�O	���Ad�D��P�P��X4QbU�<ܫ>l�t�t5�E����]m�Q����gE>�NP�Ej�A?�]�KZTh����UT4�MK�q}������D@�L�װ�sǭ;����ۦe��G�����{L���`y���Ƈ\?Zo.��MT��Q��TK��E����nGʉ� 9\�X{oC������Qs�]i��3���E �#.��(�'ʽ�e8E���U|S���3~�pz8U)0VN�8�|��l�2��k]>�5�L��H��4��?��2;�G�M�|5D͘��ඡ۾'�>�aW��U"��+߮�}.Ŭ5�>�-��=�/�~�[��FX"��KNT�4�M��cH�L&T�e��W'W����A��K��ti�\K]�O#��2���r�v>|��ewN��5�U��m�`V�o�st;��R;,���O�DƎ��I��:RnT(�G�T�T�sI�:�v���bddt���� 6���$�����B�9�+#1��B��H�"�W�ٞ�������f�PM~�{z��ڍw���X�!�����vH� %MG�׫Y�	]��yCf=H@��{��2��.�*��d�\��s'�x��Lx|�����x��q�Wf��KU��u�JTG�$'����R�t�f�d !���SL��c�ս z �%!.hF9�Z.�Q�N*E"�96p�I�Q����-���amd���Y���¡Q�n�W��š���r`�^3���:���S=�����.;w���CiFil+c���*m�;�(�w<7���� 8�}��SWJ9�ɻT��X�=����1�c�{��|0�ɬՍϣX�7�ީ,�R!������<Sr�6��������y��0}�)8�(;q�`��nтO�x�vE�롳d -I��6����;�#�"��~��V�W
Bbߊ%���D�t+%�{$d�7Jb	�zk(y R1OqК�;�@Φ�H �V�@Z�;n&���u��.�rw��Z���5������m^��p9J�p�լ��u�Oo�;��@Na���"��,n]��0��=��W���N�<�'V�����b׾�qQ��D2�t�����&R�qE�P���k��]JwJ"��RM��$�V�9_����*��SOtнq�\�{���ۦ� %~V�(D����4LMΝypVũ����A)��� z���|2�x�beұr��?z����8txU|w�6�JgY僾$���_D��m\G�5۳|�A���J�´ͺu��TƢ��H�]�����`�tw����������a����O1ـ'Aou�N��W�Rp�3�Eք��/�]���C���)���u�fx�8�D�i{�yxY>�H�m�.��l���__���0�;��*="�*��J3�ˏ���Cg�`���f���;ڔ���6��A1�Fd
��s�a�S�
���Z^�MX�d�.>
.���%۟��<[-T!m�5�Y�.q7�'��o��s��OS]CN���<"��{�d$���K��N����	v����J�����[�Dx=vɿ*�����4f �Q�U�m�����.�T����
6<9��uy@���(���9{�����S���h���#Y�%������
�L�i�ݱv6�����2���K�4�*VWk9��)	�&�Q�&l�6����4I������cz�B)!_FӔ��>~��V�EM>ˏ�P�O�!�U�N2J^��܈/���H!��@:�L��2P��Y������CH����nd�Uz�O�[���2$y�-�!��Y>�>��A��K�v!�J���:���?c�gū�1]e�8�¢xHe� :�2..�3s�5�i����%
�Y+QjJv���(�l+U2�aH 1V׾ԅA��+OQ��x+��ӷ��5�<�kNn���r�����֣�	�+ �h�8�3z��eY��f^��>Θ7�OUz�Z0��=z��3���Ĥ�ma�B�O�Ռ4oL���Y/e�
�C���ŉ�
�c��/���/Kc� -_��y�4�}�C,	y�pơ�;����X��v+�y�1� �*?	&h�
͞BeT��X�Tlc��g*��Z���Y��Iz�}�DmH��2�`�!����ڶ���9r��.H�O>7tf�SǕ�l�g��>1SH�0�H�z|J�HEP�mds��� �%�W�x=���b��@�����j�Hj��͊�[:�%ؕ���HAdyd��Vo�?��'����	�GqT�kS��~Кj:�֚t�SL���28�䢒��:�[�DY0w��,:t��a�ZI���H|g�ި�>����XCtŋfF䩤�;�F��
:��fOl����3����>�{��s�-��V֢�å�nuk�wM-ZZ���dc�S�-S�t9���~W|�:�k�b�R��;wί��X�z)��oL>�q;��Y�aQDpO=\��;��kP|Z�P�QBn��� !�@����c�R��&?����0�b�#oMG\Y /8�M�K9�|&�堻L�_֦������k��;p�b�3�mCRC]�R:�j�Vt�/�?~�ν��+�2�Ӂ�N!ݳ�I�>$�L��s�L���j"��׭B�������pF���/�p6B,	��'m��J��Я�r�tf"�0�lS8f����GB�n�E�����F�����%؞$,�$���n����;q���*�����`"
�A��4�*��b���^�<o����F��H��L��?����2�@Ť�½��l
���� ��ѕ1�1�w��n-��۔��(9�$tryTFm2M�b��Z�o},�<v��������|�@�c�Vv-�O���2���+TZ����;�W�o�!�6!q�!��ؖ�I}�Lӊ�G@Es{#��(V�G�ˀZA�{�X�
���\}4��5��5"��$G {?eM<{׺~�_�Ha�?�Mp�WA���R�H.�V̛��+�}f��L$����
u�>V�o:C� K�,l�*��Q���Y<a=*��}Ӿ����VV�عP�u�-:����װd��j/�F�nZ#th����ۜi�ܣ�Q����o���UY�q�D򀵂�b��b����sl8�Ma��U�r,��{�4^A4(T]`O��׼3��-�)i����Q���0�v�>�l{�w��Z�mNj��"��g!�m����[hYC� �oW�Ӗl���l����w�����28��XZ�"/wb�Q^]�c�(��ِcӈg���9^v�CTk�%�'��	R�Y����".� �<2	���'xO�L���E�L���șg��ė�h��c|ʊh������ۛ��p���$�:��)��ލ�]ͬ]�5$�rj0�N�o��� 8V�nC�ؓ�ce�|a��bx�}ul:��O�om�'=4w4�mO��Xh	Ф5CY�)�^�E����	 
����ż�S��]��\S�LGR|�ȶY�UYf�_�k��� ͥ�*M�8��|+Ns�\��{n͜��Ŷ��r����6%�#^V}�g��Rl����H;B4�b'�ȦC���DSz%y���Xk�ߨ����f؍��Q�����3�Hf��uJ���Z�0
چ/4� Ց���PW�2��}�^�&�DMM�r�V��子�� &�xO4���5�x05V+�&iZ�� 4�
(
�� ��~Ov�O
,%^| 3�ř��uO�甞�e�$[E��l\��=�:��^0�g�r:���ENAIֵ��CD����k߃{�p;�� �~t�Ru!�@{11���L!R�>u%�oj���vY36��>�@ô�F�qe��壙o�4(4����m�Bx��7��_��ʊZ*{	=0��_:ꉕ*V��,o��Ŀuy�>I.��+��k�ܼ7��>�IϻiX�8
�~���ɡX�'K�pG����CrV=��bg��u'��u�`fA�Y��B)S�z�U�.��5�����G�	��G��:��,��P-�\����~�I����