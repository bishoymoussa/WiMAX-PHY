��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$Rx�y�<��wA�*;�x���@�̦�W�X�fa�M-$u����n~�%���P�$��W��kYَ���P7�?UMfT��q�6�U��k�>����~�\N�(�����X�e���/6U|)�X2pF�]6x�793�w.�'J���wP������;��y���k*��u��D�ED��8�|߹�G,B
�<]&C�~H�~��4J�*E��N�$)�Nq��J-�l�$vgZ]��X����B�1���0�m�ܡ3��T�00�S��(deR�r�Y�C�6%Q)z6�i҈4O�ם���*�j#9�C�L���a�[�0�P3���7��s�X�~%Q"gd�.k�W���G�Ԙ�t�����e;�S�x����A����9����H,*��U�>D���������l���nT3�g�&�17w�&T���~�#���P��O�B|&��Φ4��V�_3� ��p�ͼD��� �c�[�;8�
�Lu��\_�_?�G.l[�����1�w�=�"��B.�J]s�|FaR.RR��e��	�q�QD�8	��|�q���e�f��$�|A���8j�3�{&�{<xI��L��b�f�%��``��y�B|� ���6�D�h���Q��E%��I�����u#�� �	5{y�dX�H��[C�Z	N��dCE�nZ�'am��*��*�.IٮG����!�_��~%�3����W3���}�����ú{p/��W|c�SB|��E�gI�y�z6@��ُ�f�
�߭(w���|��W`�/��K��<��?�Jg�`v-�f^M�*\s֍����y/Tg:�ԅ�ij�S�������=���*�{&�\}u��<]�es���������ڮ���PXZ�\��A�����;R��aF���va�ڣ����bzl��#�F:�=D���<������������o�l^Gީ!��?׌�2£r0ʩEZ*u�X�0�a!�M�į�<YxU��YF�2��{)��
F��<�7�,��D�r�zis9�z|Q �bO�X�40���H���j9�Dn��0؋5�p�P�ݫ<�$��5�)YG�?q2�+��'�W��r*w8�"
�=�b��2�jM"Ϛf:�!%D�������sy- ��(����$�cah���퉢��pk��B�x2c�Z�3�Q���B�L?�6��$��ǿ r��r	������)����r�zE����YM��n�v�z��U��і?i'`�6���"lش�^^0j�0:ł�5yt�hi�,�wX �4��C&������>��E��W���Q���^�g�91Ǝ��)�vk�jk߉�i�OL�W0����3[�p�/;��߄��F��[�2.��% \��X�0�=�[��<-��Q!��������8�$��;9�|���z�i�B�5�o����:ݰ��������g[�(�Z��ޓ0��Z�M�p_���i�S������	_<{�:'qBq����&�v.C9�WlB���,�n ��q�,j�E_޲�7���k�g>����K��{1��0cuq�7!F�1�V�NWp0G}��y&��+�Tb�����a)�@�5l!$�c�;��\�t��K9��2]'{��Ң|��Bpa/!��r~�l$欓�+����`<h3Ig��K���Ѽ�z�36q�����x��1��pR#�E�˨�@��n�_���OE��Q^@���DAۜFCap�� �*��Wb�o��ƨ�Y�e�'��ILBz���"�^�PU}���L�uց��gb��<wX��s��+��Diz��C,�KT�x����<�$u[�J�y����JRz�c��g��S�$�ھX�Ž�[�u�2��daMp�"Mڲ�1��Os9v��T�-n�6�R�{��9���m��b��cBv��^Jx��t ��`໊=~��\v��u"�"�y�������?wj�A=ݗq�W��Ht�b�ǿ
<
x��տ?��m�r4������?�Ɩ�x�톁@9	� +H�S�Hu���m�*����;�ۤn�Vav�e5���-f�SW�̍,����'�]��+���������	�W�q�"����8<d���ՠ�+L'�����L��gKr�R���P��DE$G���`9�b{����S6��w| �)���t��6�ts���G�#?>���"���� >*s&�����(Zc�w��{` �2�%=BDJ}������+~�@�[�΀T�6=$�c�z0m�J��=Y�G�ӡs/�U����FaN
�=j?�$G2!"�o�~�YH���n�M�n�`�T��q�����;��<��2:�9���襑6���
�� 8j��w|�2zp_G�/#]�!�vMq-޺�i ���t�l��&�q���p#��QNn�
�ʄU�t�~"K�	���"B}�	a\����y%sB���d�����"�9N���D��]  ��*�W��JUd�_\7�4^އ�Ƥu����z�vY����``��vKz�F���o؂��NVp"!`�a�3���C�Q!u��_[X:�A6b�v�����g�.�L�Ru��XN���� ������!iM$�i#�;�`'��w8S餯p��c�b��<�����4�����BX�*+�a}�71NS�؝Q��۬��c��$�9˂��E����?��j��ٕNڀM���F����r��
�1?`�Yv���K�љ��dd��˔V�������
�!	0�x�#h����V`�=OZ�W2L�ۛI�+� ���B��O;G@EhS;҉ݽ'�t�"���pI^f&���~X�_��r�d��I�@b<A�}P��#6�f���/�-p�,�y���ی���?[��}'T�D�η4hQg;W�����4�zQ��7�4
rQ9��!ws-��9+��S�wxf�&��݃�n�r+�0���a������9����pRW��\O�����<u�,��%�tH�M�D�A��+���VV��ޞ%�PÒ����R��HѦ<+J#m�s����ȿ���˺�vv��u@�X�-]�'P4��3P$�!5��/4��0N����q,-��c	����Q�`D�x�n5��������n#X�����5�4 ط��&[�N�K�gN�N�\&;��0��x&����2|䴦_����C�<Es�-9k��+w���l�5{���0j�n^ƍ����[#����&H�0�Q̣��埘2�E���4L&_1���o�~Vl���eي�E{����Aa!ԍCÙ��1��`�c>]ixe-�}�(^���=�o�$�Fi3�O�{��=���j@��ܰ�a��VA�%{�p�bQ���2��P,r���S5��u���] C�.��������w9kF��z���-�ͦ�W����fjk]��H!pA��%��Qҁ.��*b��!�|�y�34�<�(¥k`d��Nqx��S{��V�Jd"Z2��1��3&R�"���qG$��Fw���o��RQ�Å�<�����e�7�v����r)u�j���^^�l�"��u�[7������M��*WI�?&����V���1usP7E-uǚZd��t�gD�Cw���rh�=��*�d�HL�����5���F�����k��%>��	NlS�b�����O��[D��1�	,7����������{Z������ȼ�+��ȼ,�E���kw®�C�f�(��K9��ƅ`v������a�χ0�Q`��LY��#��;�
�p����8{�yU3�y�J3�	~k�a���֜�pd�u��e���X��(��/���#�� L�Ӿ%����N�r-ľV ��WD Ú
9�@8�i�W�S�F�k�B?o��<��sB�Dż�4b����0�� ��G�"�?-��l9 ��n�˗I�9�G����\�{��,��x�7���MK�N��+*�yj�ӧV�p��X/XX�!o+��F��|6�m^�3a��~�����	�x�h�#�QF��.s=��
�6P�?z�f)��@�FO@�M]*L@Y�KP?����e�-��k/����U����;�>�糫4�;'��՝x$����B὆J��`]q~�".B�������(q~��X�����L!�Fٙ>�Љ@��}8�L�FL��Ķi�MZ��H�-�Q���������O���j�f�*���z3�S�SOv2�U|t��xߩ�]k'pZ����t=�{<�-�� M���M&=UB���̋'B,[�L�l��+Ocݸ���-ހ�FD����׽�<�Z�����$h�HY��
��p�\H_U��h��R*3�C-o����17̝�$��)Mj,n#O3~�3X[��_�#n��U���#����1;�WA�T�Ľ�|	��5����hP�����3�w~'����HTA��^܍��͇MW�A��Q1��o�.0��|��F4�P6f��b�s^T���ض�3�ÏC��2ї�)��F��~�~�����S�"�s�x�w��J��(3�����Ġ��L%�Vh���s�.G��G�e@ߣ�� l/����^gIΙc�n��%�g�W���S-<˽���\o������0�*�
&uJ�$�u�a�F�!i�j���j2ֳe(y�'��y���tz�qj��x�ih�R�+мlzI����-��n����t�X��&�M�,t�Xu�r�}�m=V[�|ۈ����g�K���Ty�y�l�1��9c�$O�O6}���H�~��kY����>d4�~k��Y��f�[Q���<<�]!�I@]m�Z��33y.���揲���b��չ�y���7r������>���qg��lC��^<^o�'�ƕ�p͐,3զ}��� y��kWH��q� ����`���z'{{&=��J�E��GuC���?�N�~�Һ���>��H���%M[)��ey8�:ٝ����#Z+��: uC)�м��W#,��_rH��I�+���e*U�k��e���G��#��]�03�)�)X�d�7/�/��&���BĽ}w���-�ֶ�ݔ�|��+"{�8+��e��۾n������N@��?���g��pA�W�#]��CPWN������𹴯eG-��8��ɇ��N��βe�Õ���I��`vs��g.�B.�,1�F��0}��6��4��j������`�a���C�G"�?�z�?4Ӽ�ːcu���1.��L���e���q�ok�����ǂ������k�$f��U�_?%[��w?jL��	)�4 �T���Y�@�suI(^�d'\�7�!�g�9�����؄P�H3HZ&�?;̒�#���G�Nf��!ᔚ�%1Djl�dH
٭Z]�[�5T+a+�;����2�[��Z��DB��I%���|3�����Zn����i??J�pw��|�hMFJ�>�
"R^~��p�k���,��j�Z$-ֱ�����4��{�!���Tp��o({���z*l5�R�hF���D�H��)��G�t2X�Y)�!�b��f��hN��_ �5vW��>�ۍ���O��b�u��ܔ�X�_ޤDb�6��e������Å\�͵��P�	
R\��X]&�	���FԠ���<~�� ˀi���4i5I.�O��J��}�z��	,���� F�4".�w��u��n3_�b�E5���>;�����&� M}�MV���q���A�����+ɥ8)5�)�H�![�dȢ(j���{/��Ʀn����D�b���Ss xEI�ч�Q;�f;_��
�4�F��3#ƙ�9?�Vd�|���Ə�N���	��V^��5�t���<x�������#��b�ֆ߀��CV�y�W�J 0�v�����?�=I!�K�]�m�E���%^�-�f�@���]��ȉ#��BS!�P����d9w���#��-F��r��`�i�%�M].RO�c�h�S�K<�G|a�D�+z��+ε-[(S����Fh���T�B�ഌ���iNePg��Ϊ Ttf�βlFi�@3L�"�N陨�����1:d9���F�c�xWx�o4��ɲW�g�&9Y�!��6&��rb�(.1�Ϳ�[��@�]�n!���t��W,���o9����&5r}BUp��5�;���{%a���2Th=�!0yq��c�5@�?�Y&q�e�����$��K#��#ٴ�:��s��g�S|�d�ɇ�!>����w�Y���K��A���f(�+�+_K�&5�� yA�7q�w�oP��CTEDubCF��H���=�I�&d����!��Xh�h��B��y���d�[�2_#��딾Ȑ��+B/��03Ľ����ě��갬H�6AY	���/\�-�Ȃ��&����u�E>#���w�K7�m��ۈ��g�,!����S��e�*���N*m~���t��0������?4cAa�,q����]w��9���P���(��������=0�~5��
�+��u�{�	6����&�cr��|�d��/�7?]�I���1>dK?�2R�Fm�����X͖�f��.�Y]�k���ht����y�!�r��5����������`=\Kؤ (�l�ڦ?+{U[�����	�d���n�? Td�w�}��F�({��q㙏V�7�?P���1�L�&�v��\�&�&��O�m@R�~�ģ�
�X�C����;��U��R����F&We�����I�1���^4��%�d��F���I,��s�{)�ଛ��������u߀N�	"n��Ez5|�l�ת+M
����@�Ζ&M�{���o>,E��~���@A�rL�{"#f��i�8́�z����j�ҵ��W����7������)��Yϟ*s
���]/ڃ\���:>����!3,=�(0�|�O\Р�d��~��隯��\�uYq���/;\1�FS�*2���U'�`�+ˉ���M�����.Pě����r�Kc7AB&���'��^'�� v��U*{EQJN��Fi0��`�;� U�)0�]��/��%q�{6/��S��!�y���#
��g��@��l�f�n�79�~���M|G�f �<�M���-��]��'j&m/�˸W��r�O��P.]js-�z����BCz�Y�<\�ڟ�1u��u[˦����̕��)���h���8�D�{z��*c���\U�l8�6)�F9D;3����<ͺFy/��b>�1���I���Q�k	����L֙�w��GZ���,�q�ws+(�����o��ܺD���K�g�%,��h~Ψ=w΃4�\��-�}���bz���|o�}�����Qh�#_棥ZU~���g�mw~���.������>���Zd���}��wjQ]`��� ��dK��dvLsE[E���3@� ���'.;���/3O�1�r�p���xte�:�vH �z���6g�$�<���D�E��o�$`�s�"��E���i��).�+rj�u<�}�h-�b-Ny6>	T"X�Sa�I�*\Hز��e4�'#'�=�$�{R.g2)vQ�c���J��y-�gZG��������6����̼l������/���]��:�W�v,Şp��u˟e��7�/p�Y�,-�3��uEI�f�J�<TpL�v�db�z^����qr #���w�bԱԲz�_{���f���о��q%ͤ��6��ز�c�Ŏ��m�R;�2�,}���zD��U��)||��(-�F���:+V��Y��e��V�i��Mq��\�L�m�a�ד��
Z��c��;9~_��S[�N�O��µ�
�K��쥚��T?�@��m�gH:�V���Z9jA1o=��(#�60���ﻰ�]�&�1�O��S�-�`�Kaj�U�y�f��CW�_L��#���@��z�����F���2J�H��!�|`j+��KД��fu��8HRJ�G�nK5�E/M�(v8_����0�S^CC��Nv��:?�G�k�9�y�a¼���/��J��c�ߑ���"^��;����1�?���xV����0$��]�(":��M��Vu�#\z8�O~��>��P0C�?x��w�|c:��0�I�ӰB���3t�k�-�e�8|̱o�c�.l�֎�:8��\la8d��&J�Zk�J{��͏�5� k�zMj�ۍ�Ҕ�O�U���{en�& �D|d$	���U[1d󔛻<��V1�iĿHݮ��\�F�[&;s��������&��_�ᶓ�kw+��,�[A�;aYG�uX�xa�0>]�{�(���ݴd�(�а��E��r�>��~9,��=wӪN��ybGw�@���V�~;���f<ɍhu�p1��:\]}T^ofV��Ã;G���Ca��	`��O�9F��\^}m4�$��A6��Pԩz��G;��ơ�4�0����l�˥U����-:�e�v6��w�����N�-5�e��GBAqx��	Q�ԟc�4��gJ�ҝL��L{b��-��|�0!~��B�Jj ��o���l]�D�y�E�����?+Qa���/�ONp�1�q���t�F�H��}��348��H��� �cm��yE�@��H��!i�O?Q��u8���F�`����u^�Żv�:�)��f��B�I�,�ސH�e\���\��X�ـ	��a\�>^���5,"
R���k���ksq��3�M��9V�g�r�����s��ۢ�!��2)����5A������?U�ͩ��>�1�@d�b��=v��]�&.�'���Oόf�D0V��sh�(�2ZR}ʀzZG�Z,b�����2�� �����:��w*� Jl.Pf��b�c=f7`2�(3�.������j�Z��*��L����A�i$��a'��+��m[�Cp�[9��p���:{�# ������e�����͇�v8GT�S����:�8痶��7i�)v��µ�a\����N�C���m]�lm΀¹@��3���l3� �;b�>R�$�U�b̨�I��W'� �<�^Ѡ%�k����C��a�g��ʄwc�������;�	R��=���/9��]Q�ͥ���ک��3�ꞹ᥆HA�E��M��`p��&�:Q���$d���.wGŪ5���O?T�|��Z!8��#��a�fלq)Zu�BODL寚��R;XP�	��(�,������_��oT|���#�ּK"��1�4��1�m\NWJ3��&��t!�1	�����  �*o�K�uG�����_�oĥ����;7�H�Hђ��1!� xێ%<��D��3��At/e58U����.pdg��'c��S�0>4��q�P�*-<����_��n���xb�K��5*ſ�f�Y�-����lq#������W�f�U�W�V�3+6�vj��Xv���׷0O��ݴô`�Vh
�C��s�|�21�^���E��]EL#�u�xj=����D����/��?JD)�	 �h�,a�n���Y� VX�n�����m�����t1�ui��x\�.#�fS�%!�	Om��.'��#�]�+�bA�i�{&����fF��d����?~�����s�b�!��F���C�Өz�X�k=두a%�y'f)�j���,E�>�8���f�W��^���e%��#>���e9$tQ�{kq�1y �~K/��6_EF��P�l��wÝ��ے?�
�W��RbJ�
���}�+����c:r17������#ɗk�]�M��q����@�a��W*������̵:� �����jfwL�vn���m�/�1����%F1�šB/�+	�r{��Wo�){KW�@������4�o��u�I��d`�q�����}�3(ʿ�`�V��1Zz�	만��V���k����v�K���RC :0�j7�
�y,�����;K���s�_O-��?,��^���'�,i`V��h'$C2�A�~�[�T2�h�,�R�M��u�	���C��,Gzm�O���K���&��l�W�]6�r-l��wI��S^�P��A�5;c��
���g�W���Pt����S��Ƀ��O�����x����s����P���ւpck-]!mΘ�@�������|�4�|����N�n���^�T��p�&[�|I����%�F�YK���-���$���tl�׫���U��9z�ρk�󀰕�E�������/7�U&��s
�^�9��ފ�⮱l��DQ@���z�k�ۢ��R����Nv�Q%���3Ƙ�N�ǃF�����y�SC�ֺk�-�3i��,P]��1fmf�2�ǖ)`oV.��$hj���5�;�U|�o/2������\�Ƽ_�(�7�FM������c�+�ᬃ�`���?�As�ű�E�"(^�屵���հ�X��F ���f>��_C\]d�݅���%�����at$�?FB�Ө�,,�9�na�!_�	P o�Gv6�-��W`��'_����h��#ݯ���1.���+g������?���K��M�$V��Z]x�tJ�~��t�ə���{����˩�CB����p��x���$��>��O�W�zsb/u�{b���!�B(g�����kO5dC�I.(�IX��e�<�Q�rX���@s0n�Ƒ�E�a�)����B�|P\�b��0�9�
7�i�"*6�Y�@���I�:a�G�1��m���֏�KF��7�i< �d���� �Ϋ��gM�t����O����X J�NP�y6�uM �r:��xĻ��f��C�\�j�A�xS��eSqĠ^�=!9LXﴶ�h�]��e�A���g��m�iګ4�G���zyk�z���r0bC��0��b#=*V�BNK�fx[n����Rσ�~��`\�-<���B�Z^A�V��_�Z��P�F:�t�v�Z��s��yFf��Gkc8��f�.Y�:E�4`��+X��wk���%�C�I�}��F��2���q�k	T��%b@y"*��`�#�9dp��72{�Z��]�X��ﮓ�i]�|�Ħ�#DQ"����x���-��ꐘ���#�!��'��+|at�x��!���|�^k6�C�To9��qft��[�0!��-F�a(	�6\p� Cq@0[`Oޖ����ͣ�����b�`RLs��G���F��}�t@���c�L�e�A��S�v���1�R�waՈ˯O!�	Y�.��W���Xz
PŇ4�9���[땉�����-�j�˨Y%
/OL�#����F�B�)=����no �҅�Es�ϐ5����oyNDq��/�T�֠9����x�����'��h���Pp�Wz|����7~�Mh�m+F��J�"c�/Y�g���Ů�V����&�5�]x�c�tT�U\�퉁 q�؉��3����APS"-'���0Y����f�_�/�k4L��V��-��ۊݪ�n���+��i~��f@��q�8�ԋ?O*<�L�����Z��OI1�:��'��\}O��Kt�� �MA3��%��xRV}�2N���}�I��v6�D����8�V�e���K^�M���i��ڛ���B�%���t�������D��}��b�>U�NA��w�e_���Nn������H���p4�tWR��a&�ܝ̳��z+�&I +�N��lZ���SԱ�o�L����k*���{��R?��ă:R�I��c+ &`��;т�����V:m�MN�q�8�Vx�h��	���CQ�ʾ³��!�9k/�r��}���|�5��ƄHXQR��������;	)�~�5s#Vf+)�����7'$�tyL���6D���E�K'�
��b������id/�Q�����Yo�	���nN4S?#���OH�՘r�;�ѿ������\v����"���ډ�!�^�"�p�&���ģ�9 ֳ��0����ݸ������qzO���>�+<X ��t�(H�Ā,f�0�r�Db!��&� ���?�I��P*^���V���԰�Xc+Y�ĩ�c�[�R=�-FS���2��6� �'	����}<b���/��G��M6�Y]��n��w͊�Ȭ�T���aK��L��.���l+�6��+C�ؾV�~��Ꜽ�ºQ��z�$4��i��F
P�Ӳ�K�.*�S�Ț��R�M���o�f�@�9d���`ї2����쨪�#�Ψ��<}�Ԃz��~�Z�8Ik��{ͪ�A��I� U�!و��c a����X�q}�IZ�:BA�I�o	r��^������(Vi�܂k�!�J1gx��u�C+.��K��Bon�|U���=�bS.�Ǟp����6zf�0�����%9ۛ��;���,Ê�t	���0�u�俨��&�O�Fc4a.�So��޶��w�g�jֆFC���zyЈ\�U
��r	1/7�3ʄ�4������P���4`�!6��d0SȦ�������+��j7{7� �t�]������*n��j�y2؏Mb��3��#;q���{���0kq��QDb�E����k,DB�KW�zE؄cH��"2��g��dM��hf����h�CU$/���v!��k��p�k�V}�Y�a9����Vk5`�fx.�*:�A�#1���+�/��8����C�j��m�d��eږ�7.[�/J��i����X�N)�����R,w,�J8����]fl�;��g�X	R?v���D'kH��oDZ�jg�r_����$K�o�3��/��1U+o���:�:n[��	��/rd|�-����� ������*V����޽=���hgR#�57�p�&\ܰ�6���t��v=�D��d��*g� fo�w�d%�+ͷJæ�+�a��#�[��PT>!Cly
�]"�/�R�i�7����c����t�+��[�j�:"T�KGIN�W7'G��)�>���Eű�۶��?��$µ)�|3-n9���G��e�Wvq>y{��:q֓s}@��ܴ���KT���lFvW(�,ӣ����!�����1x(���)#k���w�p\\�t�Y�I�9⦣@>K)M���S��.��jI�A��Q�	u|����}�tI��U;�O���A��-�Xp�`r^��O�n���ͩ�m�&��BX�`����S��?�ϐe�¸[�-n^�?�Dh`KǑ��v��~W!{Ch�R/����eLB7Q���M�M8�X�N�g9=桑9�@W2���D��Q�󥕅��[<Y(���qO?6�� ����?�.��Dߞ��okD�9�fc[ʇz����ר�X#�X�{���ϸ '5!���m�!�$�4.�Y�W��� %C��>��?��:`��c���U��o�'!�lV'h��2�m٘`�XG4�ҽ�vXMkU?i�!�4�#����&X�2N<ZQuk���B�sܕH�֫֘�j;�(H��2�8{��ł-����3���ɞZ�ӝ1Yc��4��N9�!J����N��bW�������B�gز�8�>$���RR(Z'!|`F�&�1Ɇ�1����Ò}���o��L%�_�Xe�߿�텄������2��?�Wf�P�\ ��9%��ų. ���0��.���k���|)c�R�2��;yч}���� ��%&�[ʙ����y���qR�X���^��g��Ekʮ���\L4wͶ�p�ZK
`?'�>o�(�v���yA�����|B!z�� ���1���w�n9j�m�,S�l� �L`N�}̊�<�t�5ӗ���t.�ڋ0n\��8=�s�t�}c�K�h��g҉#�N�����(U��9MÝ���8(V`�r_^cW��o�#�r��^�qʟ�,�����Hf�`<����>�L��=	��	$���a@GT�`+kv�m+�r_Bti��I ��'m[i���řP(�;��,t�mM�z�+���R^���qPjn�'(��6b�_��:�i�;~��@��+KJ��'�I�EI\���t<&���c�2މ�-Zp�n�F�@���>IS>�� E�[�~����3Ɣ��u 2�`e񠦓L�3�UA�W S�9`V~11'�;���{����!���.�	"w9�)L6ʄ���H2���'�f <�l>=@>'���x\ �R�S��x�-Ǐ߻����vM��uAb�z�x���'̍#�%e�l�&F��co�U�D�� ����	�<L�'�^&�`Pzew3�VD&p��=?>|��!�:;�)�7%�V	�5�������7}Ü�m��qo����e(�n���n����p[���ɨ�ctg;|( ���3�:��>��|*��kQ�m�S׻]�r����x�s�kG�ǉ��\���X��k<D-st/�����W	1���!W
<J�毊��A�z;��I�x�D��o�O���$�	�>�/�`�dޡU.r��;�� TL{}I��ۋ�z���[��� �a�̨6$T�Y{����:ז-��	���sRb�MQ*���d��b�3��.��A�e��9�7�;�D)�GN[���#�s-g~��D����.�1�WK������yJ�W�ҕRS�s���	i`�C!w�"Ն��M�(��A�5�F�nj��_�� ��s�oSm~uT�V����DmM����!�,��B�
=��:��Ȅ���́�Ê\f��W_"џz`�H\j���:W�\L�����T�\fѥ����C�"�P9�[v�_
TK�ɥ���@(��&�:��S��>0�`%{/M�18|9�e/K�/xw�!^bvSm�h*,.���(ޮ0���C�ɶ�Oh���౴&.���-��|�lħZ#2:�56�z����H�ຠ1��1�FH��Ʉ:v�F~��?��B�?��~��]�o!��6 �>G�8�u<WA��^J��Հ�J�� ˨aUY�=+�l1=>����*a�����{#V���@LRǆqN��'�He�{�<Y�S��}0_�0����%U좏(��Z��`B�����vo�VY��v���s1hyH�=�b^CZ���o� �r&F9����e��$��؝��Ã��2,��b��>�>�My���.(����,��q�P��/�H�%Y�А�nE�2��Z��#�(���S�%�L`O�k�/$������z�MS�*[O�N�5&��ũ[#4' "�K�a\S��ιޖn<���T���zd��ac�A˴1?:�!��z�k1���s�3��r4�f1�p8U��a:-�J|��Ǽ\�"_���\��s:�S�e��SNa�q�q�+T7N��h�y��&�Pf�%�"���52��76;8�lad�F�*j=
,&	���Q��jo`{�L1�g�l��Y	a�/738�[�IB����]*����)We!xw�!�X1���='�ѷM9���L�T?M2���`����g�k���G藬(1֑�m��A�3�TN��{ mEu���D�Ahj�Q��n 1�=.y�]fS�6I��	%Q�Q�GS��>kx��B�}�?����pC9�+��52�;m��=0o��݇Vd�x^I����0��ڼ�ij�����gZ�GMx�fj�؆qY�rc~s��P��J�7���L�Z�f�.]����ľk�#y, �����t	9�W�em�@i}`�{��g�����g��]�zz�O��(�l��h��SXBN̹�%Hs�A�X��cR�LD�ĆA�m ����9:{,���v�_/� PkK�ɬ���h9��R������h_�Ov��G[�A��D}zJm��hK����/�q�ek�(��gg0���D��C�����m,
����s�4�-�aNUs����2ZQd��9U�ށMd�1����$GF]1�=Tz�ʚ�)�x��
G�~]K�N`�>h)��j�I�T9��PD.h�DO&s6���E 
O��6���!0�����!�=�lI�N�|��d�ؼq|#��@jŋW��h�gk�@�f2�:�����A�qB��U��S���k�/�C��B���
��Vbz��B����Wʷ�ғK�P�r\
��%�
\���P���ո�ע[��1~x�ҠU)J���fVB�^t�}0��ηvb�{P���.GN��lb,�RZ��LǄA���{���+��7��R����d�eyU
�y�+KrP�i�5�0Xo�"`�|&�C�1��ĩ��Rs�:���1��͉�g��61}ZԆ7>h�q����!u�h"5�u$_SR����#�V)�<E�U�ஃ\�6���.T������l°,��'��B�S 1Sr҉'!'�v��:�����W�}��Iw��	� ���/-"�������[�Ă:==��(#1&{���V�`��N����qG:NF���ܩ���e��.W�?.+������
��81�m]d���cZ�/{���ѐә0s�jM
�B�O0�#Y�JI�L�%���1��x9uR�%�S��ڍ��8Q�ք��}���X9d9Ebe'�ʆ�����/[萪d@/��)c���ҍ�.Q��q�L�He��c���������Lh7oG����JY��k�k�-C|^�FcE<�L����{l�w2��� ����k�Ia��_&��%�X� 8�>[��`f�xq-��.�G׎(�ZB,��wsC~����mu��1a��=q��j;}��������ď14�$
A3`-V��PP�A�c?�Z&��_U������Fa��1)k(���v?q=w$R7�ʋnYW`�����\��5ϐ2�`�Ѷ��Eߴ)��U�j<g�Gɯ�w�p�ٝ�B����Di��x3W������]�w�ja�A��Il[�Ud=�ğ=F�E�@��2�6� �Q��"j�R\�3�s'5���I$�*b{���$	)�Id��ȯXK�nr·)U}�Bw�j0�a�*������@h=z|�׌W��n���s@�|$��38i�M���<!6��t:kҲ��S*��m�%dI�����;�g��~�t��5�L{	X�5C�HN�e��g�O�\�"h��x-2(��l&���SWw�`]PRV�$�=�E)�J��M�;f���q�[^!�h�ПR��2�!%�7�d�T��@Y��+ٕjs��I��{��ћ]�a[d\���M�)�;ؠ$�A��	���^n��#�R|T�h^O�OU6�7bã`e����-���'C7�?!׽L[|���!g�C;.R���z=��b�;S��y����S,��=�#��^S~�x��R��Hhp��0SKt�ҭq�����}�[��}���i�| ����iZo�< ��S|��)�93����^��qw�>��,�[^YY��ؓեU�_"�a��ٛtHp�@5�U��ۇ���M-�V�L���:�J�e��-z�E�vQ�d�*X������W��7�|y���'p���Eɹ���;�ejVN
�7 T� �bP3�y��"?���Ϫ�I�"��5;U�ɾ�� ��@�1qjet�)'ק�0��"���0�"Ƨ�,��]�K�;���ԝ�����x�s��{�M�}��hZQ�j��u�3=�l?V<�����F�/|����m��(�c3XI�gIT6ṧ{�t�k�F�۹�H{2���B.ʽ�ǹ����8�Gf'�,��Oz=�i�^�U<"�!v5��>܅���$&��,F�>V��9%J��S�qKL��_+��K��دk�VƠj ���Yl�ЯJ�� (��4���oBz��_��u"TӇv�'D^����#�ˉ�䁴��=C�:J��B	��+m���:�*}���^H���a���,��7_�)�m�����ќf:^a�b=�O��W����� N6��6����e|S�Ta��񄣆y$�
�ɀ� �g���G��M�6K;�q�Ti����i`+�yY̎���֖*VRZ��_��y�տ��B�E��+ʤ��T���m�'�%�`�-I��0�~ w��<x�06��O�5�Ӟ ���j���٦}D0J�V�[�Ӕ��W��:�za#��C�#�.�w���zp��t�}})Е����!MUM�Ner��3=���`Y|4v��#ʏ]�Օ&�jU,�:K:3#�%թr�ݳ�N�c�j)eya�[�uD_
�;s��32H��mix�#V%>�p�
 )���u:�A��:��v;	OJ�ͬ�DD�fnNO:�@m`iZ3��m����5Kj`p�L��-���K��t%����x��Yw1��G˒H�c{lV-<�wʓ��a9m(tP�D�u�����h-��&��5Yƨ/Fץ�"���sE2��뙞I�3
�o<'L�^" @{x�]���b6�x^�f��`�R���R�+)$�~A�D��|xl�����~aJ��λ����Q�~�rT��P4�S�H-`O�6_6=ĩ�\�;O�ev���kt7�j��%��/=��B�m�D���\o3�ͩ��y���h4w|�c�nq�N�(g۰J�|���hy�.�o�b��A�'Gm\+8>�Օ�k�t�	�������۩��-�2��I���Dϖ��Ѱ����������q�'��`=�<��=k��M�s�k�rvg֘b�V����Z_�!-�c�H�:@���"�OPj�p�K���[5�T@�{�͢ϭ�K�(eV�N|ީ��C�9;����ф��8�ٺ�7�T�r�V���Z#�t������.X��\�{����}�{GJ1z��N�&rL����/AP��9��c��0��W�΅-v��8h�wB@��	�w�	h�Ҕ�@f������r�%qe"x����,%�x��C-|���((��u.>f��{��a�ͻ1T�X^u,qB����[�<uB�_,Mc�0N�&��u�
���T[�?O�[ؒ0�F Y;|�8�=�bí��fD�#�jH��G�l����V�X�k?ٿ�7�{�j�W���O��P�ur��m�}xH���-��o�Ou� ���SO��H	B���>5���FxJ���0���(n�y���Jm�W��y����:����-R�x�#�u
k�>B���W(R�&����f;���]���m�9t_-_b��:m�@]��=�n������~�"���Y w�8�Ķ2;#��j���1rD�c�0��m}=�D�[�PW�ߜ22Ԫ�8?�>2"[�+�.}2���b+@r�u��GMU�!�e/��y��dӵk�?��C׫Epv�T�/�����e�DF�i>WN�2g9U�����j��������~Yr�!��1�Қ�L5�򩄂[����J�.p�1�j 4�.(&fNxI����Ľ�r�1-q����s�nN��Ix6����U�pY�����$ZNpDi�5P�Y�q̇Z
yߔ�ܒq�ݜ�?*��S�M
�"`�2���dD�U���*A�����{':�Z����B]�jt_��*��F��b
@:�6'����Jk#5ɸ���D�� %�N��f�x�lژ��u,�]d�2]���Ï��^�S_�	��G7d�C(� ��l�z�[`<�z�F�`���s�ҿ��v���֤5؆�%Ë_M��U�]��hW�BU.�;n��qA �\�#�9[[jA'(����r���䠲�( ��V)`�v�Il�G�o�X�h$"��6�oj)�xhC��T��2,�Mz�(i�s r)�Z����ۋIb|�����^���O�ZzȎ�}��1��(�K�W���XǱz�H�5���1o�~hU:��Ӹ����%L��IgG��˲��Q�o�^){6��*y��^KV�ۈ6���0<Up-q)��u�&Z�x�ԝ���}Cx�Z�Z���(7J=��g!L�����Ra�Gl����D�7�iL�� �捾~@p�ԾvI�i� ��K�x͏<)#u�>q�"^R�����)�
jG�����p�TT�'��Eu,��i�. B`Š�y3DF�V��U�$�7���D�����R��u��g@�H����o��5�q���h9��n�}�Ybc�&�z&#!S�o��q҉v��v���c���(�E���a_x��1>��TE W��dP��(!�A`�)GC��k�R�%���l�_MXs$g�I�|n2r��ȳ�(ܫC�ڧ����S�jpm�L��Mh�\�-����.��tl����}�׏�N�c����>H��ߏ��ڨiC:�AY]2����hz,n����5��.� �F&B�D��(����`
-�DqA�?l��Y���C�뤲F�ك4�9�B�zk��P��i�k���7-���)���8���+ofh��izM$�����9�#�rҷ�\��-�gǅz ��v=a��Zɐ��d��#}o�w����|[d3��^�-R%�yf��q�{N `3�_@+h�z��q����O�,�G'�K��9��B�-V�$���&jqeC���22ܦ�Dn�S�/��q7R��?z���ä\G��B5X�Y`�P�p]B��-��P��M۵?J�0����ڸ�d�<>�?��]�{<����C"m!�H�EW���+lv�V��_��nǊD U���=�ʠu`�:���)?壟{U�ģ��W��#`�w�qV>�$�k�c�S^.W$0�c��t?��O�+x>؄�8�<��b���R���;{g��&��(�AG�A����A)4�q!�wrе��O��9�×�VBZ+MY��F�V�yZecԌ��Lc;�{�wT�-JP�+��_l�L�I�}��p�<G�z�q�y�]�~�����$� S��T�un(̱�ܿ��B7����Y7�d���
�F@zM��sm'/t ���8i'����I�y��^
�]��Ք��WLiECu]fNXb�.޾V^���i6����V�>�.9@"�zx���2F1@�q��1�[�Id�A�����f�뽴 ����7ɻ��d�K�+5� �_Ǜ��c�f��gl%�'s��b?IOē�t�W�\ׂ!K^�� ��r�Lm�|3�G��7��SP��'�@tcy�;��}���59{Ƶ��{��x�aF�c�$;0�GA��`�7^���2��I1���j,���n�����°�^��C4�lۃ� ��M �-�&�o1��F��Ĺ�vk�uoجx�n�͝�&�.j`�Si��Zӌ�������s�X��}���@{�<Y���aX��cx[}^��ե4v��P���"�)Jm�����Ϊ
����MhN�>��ь�����B�dw�k|q�#�7��yNԞf�X�<���u_S� x��RO�"�b����34*!���C��-��US��+;���1�~W�B��pC��1�ߢ/��#���AB_���&I��6���p�$Yλ�!�2ŀrnK��*�ҩ���0<S�;ͣkp���c��p���`�7rs �f��FW��L&1��m����(N�VuB��&g+��Na���LJ>R����T��Sn�8�)L���.fy�J�Dw1�z%I�R�	:���>!I�QG��Q)�ؕ0��x��	V���4|Sӕ��\�j��R�a��>�A$_����F�����K1g{n�!o�VWI�̅W��P��a��<ZtȆb.�%�+'�*,�nTJ�^��6ms���`6U�e�$��D+K�3��I��2��ݮ��e0�T��]��`�R�O��6�ց\5Ǌ���-�,���Hn��ۓd����.���.,��A���ݠ����T0a�#�c���5ք]��ӲٷBT����d��D��\��fq;t�L}2x��c7
����WuHzJ�$P�<g�[�;[qӯ�`�Q�xx��I����`�Of�f�/h]�<Q�]a�F��m�Vӟ�4�e>A��.=�݂���y���@���%z X�B�$)�$���彨Nu����$$��tϙw����Hl����c;��ڜyI�I6�����y]�=�E`�\�ϐ��:}kp8����va��k��U���v���)�y��$W[Ӯ�8��M���%�P�Ha��g^��,x�"�Wz��G_��@ŋZĈd�v�^��1�5���5��F����!s��O]�ǣ)e�p�V����5}�����{�d,E;{HY�F���%RI	�e@H*|	�1Q'}~R�ǿ��x��a&��M</d?-��b]�(:���c.XXr�H�[��P�?��"u}hX��,�%�s��]�^Gy̈́	b�F�U�!{��t�xtXíb�Zq���V<�m]h���|q�$��pw��t����)M���3�ڰ�~|��8�( ����n�g�@Y��~��5zI$q�<[�{���)�'�(�"��8A?6�__/7j��׎�"�)�?�S��:� ���[�4m��kڍ�'�<T��߬V��7����'���.{�������s�:T�%X�XO�&��[mc���@���e}�#�I�դ5�oYѴg�y�PZD)W��:�R���{���B��ލ�O?�m2�$�So���Bz^Jj���j�gIvF�p��2���_kz�܅GV����G�~�j���� ނn��zT��X��L��_V�t�?rlF��na��Ztb߮i��ͯ���HE����[���9j'F#˟��Ru����A�a��o��1��p�9p+�P�a�c��e�i����Ք�BS�߼�
�ß؈����zh�(����ބ]����(ě�?)�����f|�]�3.5�5Ձ��"���tϸ�f/zk�T���&zg��0	s���&`q�AaA?�(s��Y66w�h���{=��hF,����+-�Q�� �1=\(h���f�/�0f<U��sK%V:,���pd@t+RO��l�׶͓��р��������,�.Ӟ�����H�h�ʎ�����U	���mط�5����\u�s�53�b����V�Z݇R���̻��s��^���v-�]���j�������G��x��1��g$�Y���H�� S�V61�X.Pӛ���6V�:S»�~�h��Z)Ό�� ���1gT����)o�M�ǣ2ͫ�0�3P�2��~�-#��)3����<tS��/1>�J۩��迈`��5H�r��
@|
�(ζR��.KQT%�5l��Uo.u�Ν��x1��N�6I�w��@,v���XN_�ng�t �*`�U�P���@��?5\=j��(����Sn5��o�Qs\�[�[z��3̷��'�J�6�����==��뢯i��P�Q�4��K�u�G+��~�H�O��`�׳DrB#��N5CV�%G1L�v&�(��O5n�-qb妀���V�&#��Z4��)@g	2�)���}KM�2s���ߎ�P��a�m� �t�r0�|��N�C�;��k:Q���G	�j�Qΐ=��� ��M����j|~�47������O�$��LOn[��H������T¾V@�n�d���]�5�]l>M�Z[����SK�	��+`
"��&Қp��Ӿ���ɫe���Hh�G|��T4�Z�����Zdd�]����[��������G$�0�ڣ�o$nx��cΰزp�b��h�_�mn��5���7li���,�yNE���x�#�К�{?U�Mvطg��ݘ�b�M��<��j�V���eAa�Ό��5~�;f���Y/����
^��/α�
���M�g�D��ا��bn�D+v�=PO��M�i
�jf?�,|YW�#�=0�(��I�'I;�˨+Q�b�.�B쯦.��	 �=���r0�6��X�{��8طl�g[�S�K�i��k�o�O(w�N2{f���h�5���߱;��q�t�|��i���~3�0�,>�8��+��,'�l��PF�P��d}�5nV�lrf��O��H��uZNǡ��qSs�����*�&��c��3>��Ш�ѝ���+���MR�6��.����s�1mn�r����û�7C!D� pj2=Ṋ������=G"���=D�Nܬ�U��K��RKs�M�=� �i���_O�����i�kԒ���`gda�\���(��$\�5�d��{R	\f�����]�,���w�+f0R[˶�R�."b��zS�9%�e���L"���=vtK<�(�6�'@�;���+�Θ����������`��#vƵ;k�O���\[0S�e~�(��|����������@g�J�2��Y�L�"z��qG�t��D�^�G���2���&(��߿6D*�u�A�6���ʜ���ۡ���2�$��t�,|�û4��54P�T����X��5}�r���-&tE����W���T���:EϢ����Le�1��,EFk�9��Fj^�.����c�z�P����'�?���|^�z|r������ �'�(��Ǿ����'M��
�'�ʚ�<�3M�៎H�mO3�'��P;�\��?�V����G7��~5����F�OZH{_���'7A|4N�P
�Q�)�K��e_2��4ͧ$Z%���q����.���:l0���9y0`,��@H��#'2�=xUC��zjv]GH�+5ˀ���fi�"W�3����3�쿽�kS|hr�Z�zΑ��!�����rx���Dǰ������:s�w�}�,����/����6����`��"���v���H�C^�<8E�m����2�忟N̼f�a����}<5!,e�htP�8a��	���d�S�fyz�c��8<��l"T<�������Y^O�uf�}��� ���޺�n�j��qg��QaH#��_�۞z2D/�z�oa�`�rC���Ĺ���E4�U�t�E���9�̚�
��؋	5�ÚB�2I �t��E��������4nK���b{�$}	W7���>��mTr������9���
RS��A�B�K�O�H�����;�x�<�̑�������S$ZC�^���s�,4���������d��abs��6z�RK��X��B�Uѹk�ȡ���΅�;f�,�%�������ٌ7����I/s��4�ȕ�_I�و�	��ͫ>O�"���V���kЩ��������g^��C�#��C���ʒ��XhEa���+�Z����ǫ�u�_�k� �\A��A���`" ����POM�������\�XD
]��z�&>/ ��h��V<x����d�*e�>(Y7X���p@~�{&c���߮�D7�c|�f'�IfcK�PNý# <��^����%=܃�7p�^׮�]$=�3ȂуY�rb*���4 ����m�;�{A:�W��Ϯ�'/@#?�����qݒ@��Rw�z�����:�o2�xQ9	�J~�a�,���4����Bv�:��#xj����B�"B~]�҅�I.	vW}���%�]HHp��I�F�@�-�����NrC��T��ql�t���d��T	a�!�]�Xe��o��
�mT�:�JN�X�k1Һ@��Aa}�꟯�ޠ��A�nQ��#X��81VMG���/i<����<\6�����깇�������9���'G��+R�ঐ���u�ÔoQ��G�M.�؂���:�!6�W\��V£�y�m�r����
0�憼vҒ��W-��~�A���_@D���HY{8�8c�����*�����@y0�c�8� @�x��.�������/)oWu�#_�-s}]����;����ק�����[d_��ڶ[�>R�؇p
�$�G[
�suS06w�Z��{��CL��p�F �+U�����G�1���'����	G�g�;��C
�ҥ�����y�d[�c�3���pj�L	��,R�\�dO�cv٢���4���#��]ҫ׭��\u$T�5&C�;�>I Md��"I:�>ȽoAWQv=Ց�,>xo�e�6�~���'���b=���}X<I���--�MV�5�m}��fi.#�eD�;�%�c_ݒ�%����zATr�{�^h������,��bX��#��\�
�>-Pd����|���,SӋ8S9*�oS��F�K��?�JR����!��k�D;�!�i��AU� Ü�}l�됭L�ۅ*�Sn�qO!w�W�]g���
�oV�+(G�a�.�g�v���D��FXI�dg���n��L�W���,�;T6rجԯ�l��?�m�I�����6�0iD�/C�zt|���J��Nйȸa�B"��Шϰo�� w_vfz�y��0����4u6+&�HK�jL`	�6x���&>��Sw! �6��G��I����2�}Lj��0��mb^��%� ����g��D�p^����f:�IƝ��Sy@�$�c[b�f��U٧v5X>mL�V��ߴ��]<�G�>�XYfP�q�y��Uj\�����!u*�`W@4t�>&8����5�t�=�o���|��|gq#����N��-����e9��A��B��	^�p ?f��k�.x��控t�u�U���{�>6�J�:�
�W8c?I(������x�\�3�$9��_w`Y1-�<����Î� .�r&�:M��-��:�?w�ѺQ��X��Q+&��A�5�1ɮvf������k�����nu��Nt)�"o%	���K�xR2�e�1(�b�v���������=�Gn�G�v��=ME~��\jn�{�g��ʈ<�;A�3D`d3&t���~�c&�jGi��ۓ��,��uU����{DԧԎ�^�\��Bv-�����O3G.�#W��L�ʙ�4�$:1c��8s3pW�9q��pM�,-G�ns�N>����w)-<A�7'�C�V��6pkziz�2-�/7�i�X��>�#���.��F���f�Ј�׷�%���ɽ���d !�&f>��q�ґ����.�S�{��jaH
2W��P)��y���/%0R�Km�ʇ���5q��Zk9�'��g�[�e�('���Y}��N�-^9߰<Rr�ӟ`H��ǢG.bdg��Np�%����Am���;��� �E")h��l?�]�d����� ����_:�[��K�5&�ͻ�E�LN�K�J��o֏5;	����2�M��bCs���^�u뙑M����R;�^4���cOWv戂��hq~uX<N��d|&=:U��e���H=���9l7z5�fvF)�q\^��3$�v��.\H�z�rb�u7�$`�c[R��.'@��16cKe�S�J�X��9j��ݽ�Ӏd[F���A����5��8Fj������ss�	��-}�����?�+��
)@_�3;��=�NGg	V8B�oQ�^�O�\��3k��}��MSF1�r��"k����ɫ�%C�I��=1����o�l0D�)a�,�f�n;D����ƦP�1�*]����]�8��a9��|�Άc�-���I�u�z �R�G��u)��4���*pC��$�ꅌw� �
���	aB<�{�sTS�Yk�(�˦*�-5�y`��������2�_�����P�,|Q��D'Z���������G?��0�
���-$j<Ǒ������[n��f�F�,u�^�&��ss�!p����Ɵ�'����B�F؁*���(�P|���u����8i���Q8I�Ȓ*��j���:ۋE��6�#�.�e��q76�3�V�Mzg���x7V��ȵ�|E����P�!{X �$���%l������cJ?��
G��;���%j�b�����#��ڙ^�;�ف�q��1��M�˔֛Z Q��d� 8٨1��=��剭�$b�2H�I�W&�G�)�„M�j(�˸��<�ºu�CX��%�d��+��(�G�V�@�l��^ی�f�rn�'�퀞��|42��V���{������x�1q�t��3{2d�[#ǂ�z��1D<%����z�1�����f�ﻔ"33F�#x�5���R&���KZ�p��
	:R��;�!�B���N����EtЇ��geѨ!�j����r�|����3`S'�N�W������m�д�\b���@FN_��Q��I�D�T��G�S���"x��<l�`��:Hh ,���K!�@���F`��tyJYgS�]s������e����[x��9�\#��
�
՘���m�"\U>P��w�m��(]��>S�pA��3��T9���#�P#:�&!
����@=Z������_~��"9�<6��a��0J��9� ��}i�<!0,r9�7߾|`k�k{���̋�5st�L:��A@�#ٽ~c2�!�a,Ū�]V�z�獁�t��ÝR�[3�ǌy�2�$�We�)�.��I��kGX"��Z��`�7׻A�:�?;c����j����v�b�r~8�{(����$ �B
.!���L�(zed��%�^-��F�&8�[ӈ�O�JX��{H�>��	g|�[�`��G���@<;\{����݃�YѠ������;
�1��/����lB^��B��Jo_$w#�٧H��[O��.��c±l�q�T�g����J�'7Y[qlsT$���p��!�=Rm�G ��Ñq�]�?�F�i�g���>��b�.�����g6�9�zf���K'�Ҭm����֙�y]��/6��<����x8�.//�O�pD�2�6�=<f1�F�E��)m\�o�y���n%�쒢�B,i�����QͿ3G(*t����"�i�Q`�)��CU��qe�2�
��*�����9#
FdEh x���d�ꛝ0�`��:V�0«����f�p��j�O���w������V5e���fh'^��l��Ye[�A��[�/B�k��}�.�4�l��[4>�Q���˒0�Jķ�v�|	I��$��l<J~(:"%H �h�y�2�)$�p��n2-�̣�nᘴ�,nn���$�A����cװ����P(�����0���@�x����A�g�`��w��R-��
�\*�����%l���$��D*��������e����n���
�!��Z�'���S�I3���'Bf���2K�����~�|ɪ0�aZD�`�F w�C>�b���p�r?6��ҁ��Ƭ7���8��ȿ��������7����~�����ձ��x�E�8��m�aGo����=�,�3�,]m�#2ᑓzj�v����16�@�9ke�U�D��:g1���P�3�L�c�������Ё��rVc�s]"�����J��؀8+� �K��Ӡó�6����$�/��K,����d�2�0�}�m���)*hK��6�"�ǃO68=�1O&��1>ml�M���>�}���o)M{(��yk��.z�y߱��Sˡ�w\H�1w~V���2�4��)2����wc��p�Cw�q7Ӻ�-=�T�@I�I��,+��cO�&h*��.c����{�}b?�߽��s����L�d�♩K�1i�,l��e$y'�OC��Jش؂qV/��SH�E!�����\��A+Y��a�b7<�n����*��Yr�&��C�sF��#�1�s� [�Jn�h���ᧇ;V��މT��E�Z�A�hpr@r�ׯ�[��%9�O{.�����_i1*el���}\d�阔�8$�|_���᫈�����쩚�ÆsU�� %���t�Ǖ8��g^�u�GV�����B��<�</�c�]�*�-w�s����X�kڪ-�-]��Ǆ�-�ˌt�1�X£A^h�I�	�U��Õ+���9�,U�G��n� p�g^ζC*L��|É}��]¼��o�R2%�Y�N��1��i��S�"����j���xx��vp��n�K�s�3>nă7ڬ�CL�-�>N.�G��o��e1�[IU���A�u����w1���H�4��s衝N�{��us)vܷ�pH�.y���AF���R�w�i��cX�f��p��IL�:qMl}��c�C&��śx�����sr�~6 ��e�6&�q�TZ_�N��aEy�"Gn�1:k�nz�B��T��ML�?i��J� �-��۬��ς�-c{�u��R�o�ÿGR	�7��2��f�.���2�@@ln���:��$u3?����.�Q��r\<�s��DU7>����k:��g��	2�?�EG����!a��6̊��^�D�Ђ�^�ȭc�	���P벓�)������H<�s��T�>�D@i�׾!���#�����!/`�"���(��r.=�*���{[���vȍB��{��dՅ�~g�.w �aN��|����0��
��y���J�Mh�,������Y�Pu]�A9�Gl7�5pͷr�_J��
]c7j��ܿ������li�\����0C��SZQ\-lY&
��tO��B[-ݜڹ���ȻH�L#��{ݮ�3��<`"�}���o}���_�\n�F3t�P�B ��&b�K���m$o�Q_q�2gW�&����S�&��u��g�fL�[qm�:bj?��}����H�U���z�`��4�j9��&DV�?q���Ax�@2)���OGLC��_�Y�*mfBuuNz#�6��|�s%�X��);H�Ltpq�mB؂M�s�2�m&�(К�N!䶳��l�_sު�7*l
~�E��{������J����U�,:x�WRs	����o��nA������3]�5ӝ�TG��
i>�Cqط�C8O��|�}ҫ��6G�=��Em|=ً��j!�<Y%w>`:�hNo>�ɕ�~s� +3�D�P�|�vjĉ@e�D�Zm'�`�.�B5ZWNbi���DO�E<B��t��(s5��n�[73��u��Q"Ԏa)jJ O�6��3�n��R�^A�;Xo�z��l��G��xo��)���l/���	��'&�����N���p�g��gq�z��o/i���	HF��,%4P�k�# �P@����!�����Z�V���*�d�\Q�=F�Z���4*#��K�7՚DQ���jӀ��������*B��Ơ��B�g���rA��J�G���4k?���[���	g� �Sȁ�'��z�Ϸr��bѯ��`��8�l�T�=�`0��IK��˜=h�Bwێ9"g��i7�)��Y�;�(�|>)�&���g��t��]��,cI��R�z�.��|����D�E��U����y����`�4=��1������Nt�e�s^�v����� y^�������-�e�[π�?3dH�͇����U&h������g�`(��LcN�aF�[���7[�;T�)Υ�~O�lW���mp���h�;�Z���;�C�M��R՝4֡�:���F�2��q����
7��t�p�E�5+'�x-�)鍖�]�G	��y���N�:i��,Z˦�^��Uo��겔�	�����}�a��
v�`=��{Q�C��Hi�;������ �l/��ܣ���A\��qh������7�.3�?�Ս��X�m�is�y�N+��$2K�X�x���D c���N�T�u_����"8r�L�8��iJ��H��7�.@�u��N^Lc'��픅v�x�E�R�t�)���/,hi,ϔyR���%<�y8�ۛ�&V�|ߔ.Ӣ�K��<
����g�v��f*?�@�|��~ޫh~�wD��b�����R?nJI�J�F�(��rҚ���oD�1�2G��[�|�⩰�R��+�nDuZr��?8���� Y�(�M�h%<�G��6h8�DAt���*�
J�`"�-��'��<uK��x��!?,����(�Z�$�q����P�����M��PR�e�z*#yj�4q7�dI���b��K���Y�xG\p}8�PUfå�R8ё���	�n
�4���T,�s��	S<�@�s�P�:��4e>P0F�}O����%fK�ȥ�G3�Ds0���RY��"y)�m���T��f�����c�}"�O|E6���}2�-츖e�:�x!�S$J�B�?��m��\�A�H���=4�7E��C�6�w�6,�Tu����d:Q�C�n��$)3������0��\�vdT|7y�`�|�^>"L��F�00�up�1й�_''�L�o�Ñ�s9 xWY���|Vr�h�oYǆr���0����F_�d������������m�;�H�b_��a�h�K���E/���/O_8�M~��d���-"Z�_���F�/����� �ɿi4����J�z��!.˥~#s�S:��s<�s�l�O��~�+Đ�"�ع�b:1�SMS�م��Hu�eG��dfP�-���!��B�:H!~w���8E�890�g�z9�j��ǯ빝�
��(13���N��{\�ޣ'v8����ޢ�S��jX;}3I�;M�V���(w�C(n�?<A�K�E� �D�6��^b�P�H0��Y%�~67����|(n]J�/��Ⱥ6 N����b�wa�uÙ�=mW�2:�W�B�7�g��9�ej��ɲ[�9�E	g
�����iek,�<_E%����/.��5rM~:MZ������_4&�������;yN���y��1,�M��K��W~Lb��.z7`N�����eǶ=5�������z��	���*�\��8��t@昢���<�cs�cBc���R-�g�� l��`}��X�>�e"	O ��m��=�>	�ݞ�͙#��%Tx3B�H�@���z�N�[g��K��=�{���"U*&��k��;�t��9��I��ze FM pd�?'0K*+��x�j@� O,��:n<����%'y�����b�)ė�ZH.�����5�e���ڶ^�S<�u�4��K���!��;�;��9*(R���!å1�"whm��7�qz�D]1C���En\�dv��^�jJ_,T�2��=�+޸���\x���޷:߮��@�V�5s��s��*��Yc����ނ�M���Aq�����"��|�\�����i SdI~mB��"j�R֌߲���(�s��Ap$!����4�V��R-'�����ٴ#�<?�a��D��C.�R�-�HHk/�o����O�M��n%��G�t�KL܆Չ����S;�vne&ة���̙���D��/�c���+���E�UD�d�2�Zt.۔�pI�W�PT���EK9��o ڦ��H�^�K����O#w`s�.綬��m�o��e��9��R�U� �ce�&�����_k�p^����O�U�h͘����x��!���t�L%��<0�ۚ[�זM^�����Hu1�;#��	{/�it�����
11�&���x)"��Y/`^g�-#��^�/��9y=_�����ܮ2�T]�5Z6;:q3#�K/��<�گ� � �4�'T�����U�йpP,�Ul�]RK�[e͐�����N=:4v�=�^��.��wg��W����8�1=B���Yj�nj��w��^���ˎ�U[)bnI$�!�f��'E�q�9bLm�1�����(Y�鈒�����o�!��Ȳֻ�g#�N�z_�6�GrC)pS�}���"�u��HH�f��5!���ʬk|'H�7,�t�� ��a�?=�ԯ�YN�<��=`�"^�o v$�D��Hi�"��<8*�^?��)�WKp��ߥ/�
5���GR6kQ�����_��hxCR:f� E�"�>�J@ ��.9�}���A- ���c��X�������]v�Fp�����()HhE�rJ�F&��s�n��*لQ�b���H��ϔ�Y��r8�+�Fc#�C:��є�R8W[;��۾�"�i3'`�x�������bE��P�eJ�w:���$��G�i�����:���V��A�P�P�S>7��i�5�p�s��6����I|)U��bЧ`DYb�&*�@[*�)�6��Vm���̀&#�ޓ���t����p�⬆�hȹ7{'ZMr���z�W�LZ��^mӾ�sP�x��શ4m���H0�C��*�R(�6#Ϙ��	��h�����2�Q�-��D��7�F9�I�9M��^�0������k�T���s
�א����. �����f	�	�g���^��O�')6���(��_7��Br�:{N����_�>�a�X�2<�hY[��ݺ9�}$
V
��zĿ`ۇ%���U2gO&_�rX �$Oۻz��|�7LŶCE��M��4�s_� 9e���� �3z�t*ҍ�#ږ���o��ְx�9��S�W*���gYs_�i�,B��l#]}Ȳ ]��b���'�?� ���{�f�oPBP5��ɇ��,�#)J�5���6�#�QD�
:6
�H�L��l~ڒB*'�;�|�x�3���	��O��Ԇ٘����Ss�z@��u��__�)�Ak�HC��[M.�c}o�u;_Ɽ�y֯�+N���"kp�ĕB�`%���˓�u�D��d�	�*{���I��3P(NUG��-Q.Q�)�;��:Y%]GP=�D���e��&�ݞ��d�ς��V5�F���%v=\��SG%fIN�	=�����a�W%� �R�!���PPX�֖�F';�b��)5g��,�e��;ӥeD�/��b��A��5[��C��(0>W"�Y:{#��R^���1���U<&�S~!S�C��&���B�9�nX�ƶ�ℱ����e��}������������x� `�(my(�ԹIJ��� L���:����"��JKL�~D�c��sS<�Uv��A��!Y*JQQ����x`��ʖ�ZY���	rX�����4��Z�Vt�s�~�Y��tf
�_>YM�#���A')�g@n&/�<��KO�� �Q��4�k�(�iP�T��z�@Z��׃Ki*�rY�¹�����q^�hv�cGRk��Ю1hO���S~@���x|�p��9����W7g{)��M��Bjr��]�ٱ�D��b�IYB-2��bv��H�f8�p�/���,�\���@ex�rtNzX����;�8g�g�����8(9}$��z����E�8�Q]���������CRrf�֧v?�^��]�GY��=!zJ�Y�Ǌ��s�3�y���I����}C�����`���i��橸"�u<�&�<�ɝۻ�!�fx�/���.!H�>�lO�ȹV��]���&e�8�s����R#�h_�7��VP\ٶx�w��(�ϧ��Ѕ̻�k���>a�ƪ�,�F<��$��	�]?�^AQ��>gJ�G�8oe<L��Y������2;�à��Ju�N�d\���y� �����!���,�tni�L�O�0g#���*�b��d��{;>�z, ìAx� 3�B�� '���AwE��Q�j�귱���-�W<Ր�p��+�n�U1�>m��SlsN���ը�n���)�b�ʋ��.d�{�X�)�a��%����6���0S�
��jC����yw$�&`�|���AIWc��m������D ���e���Աw�u�ߒ?�����"�d�$��q\#�W�9�ﵛC�lBk��!��OHBF*��
�������f�&V���66��A�&K���_�������W7��/FZ�d!|�9��Vcw�.B=RzӨ˥��&f8�n8S �#��o����W���[�W!d�XB�k.���1��m[A΂��3�W�0l��7�j�,�i��
%M#@!\�s����s�<I��64=$��BRT'Q���|��U�̀ᤳG�P.e����mgt佋BFk�#��_�O����Q��z�%3_�����3�E��2(��<�鉏Dy� ���T�_��(��h�t����觰��=�p�U��|�������Г��W�25_�RC
-w�4�TZ$�C���Q��T4dt�wS��1��AMO����(|��^�
녔� Y��"�NG+�����SDUz6,���|�$�Ss��w������l���#�S#��l:��4�$��7��g�-t��/X�2�U2����a����^A����_��e��ex.�
�i���]�OS�;BR�+sӞ���l�)��`��$�:�THMJ?D��x1v�Z��0T2(�D�5A���R|/WC��BJʵ�:�TĒZ1��*�P��pZ�Z��}�>"�u?�f�-rNl���=��I����!���yp�ɠ�H�s�XV��_��E�9�6	��r'�%�Q/
R/�=�uel�	zM���c�s�+ 55�L
��`�c�s/ ^rﾥ���8q�@����W�Q�hħ��h�cMo�)ڳ�����Ԁ'�ȝv��:�Cn�iis���ΣF��S��BPf�l����7�?�f;�����b�E�7�/zdkػ�	�OĪ��}�Hbw�V�1�Ǯ�Li��G�"��� �"C�� =��<ov�[�HZUp�7���"||b5��-G=а-���fd7��Y�w� ��a�om&���ꖟ�T��D�<�3g�r֤����^���W�榧�
�.�>�D3����E�\�W��e��n��������]��B,�/���RA��8������バS���NO32퟇y�GǦ����)��;Vѽ���I��0X
4+6L!J��7%s�m�=��,s�����J|j]��b�0R{\r���3�>C7��x�KT��w"�5�Q�yX���ꨂb&Z0�#�o�|���X�
�*g��!~�t��.ˬeT�m8�����8�k�g�� V��c	�n-uzx���Z*�'�*��c�=��zK�	�.�d�ĸ�����>W�J\1V�h�\:��p���ͧqfcK=����pc�Sf�ZO��2������S
�h�4��>�d��Q�k�&��o^[�w��^H�o�3ތ����^���#L���[�~�RS�b���}e���(_��mh�[�Rkm��A�!{��)��!{�!T���ۚ�\{.o�9��aͳ�Fh|lx���\����ܢɭ�y�����5�MT������[r.GL�F� ܢ�%L��o�����f�C�����N��I<T�iw5�:� �����3t��T�Ʒz�y��}���� ��x�E���i�t��R����d��N7P'�'�QHdo�p��[D��xq8[�RSb�w�����	�ۚ�T��H�M�9���DB�τ��2�4����|h]��r!={<4�?hQ+�>�,�Y5X��p&G�xbvE��Е	FQZ�=��>8�o�Z�����;t�-!L�}>c ag����m�p�P�� �^�D��u�����ˉ��ﲤC�w�)#�_�ˊnQ�R��nպ�BQk��/��5
��B�f�1H2��sM��_���vX���𘰘���F���߀�u�%�*�o��Z$����׼���D�+���Z�H��pl'����i������YK>��֕;]�v��!d���G����Y�>j�RP�1�}TD�V���"-�/��I��kkl��˞��RM}]$��:�ބhB���q�0O<���B��6����pV�vu�j̹k��#8Y ?틴~잏���%C�^�QMR���@����t���Ȉ�_�p6k6}��������2��0�P�"�"��-�Z{rG	#⣞�.�y�! �tH4�@�VEI�g�%�6�
;K���L��zY��:­^�� ~�����G1&�v[֦S����3�B��X��ޖ-r�%$a��B�zԀ��#M�Fve=uw-Ą"U�:�se	 ��7:�j��ڲ��Ij��.�W~���O";	���*h������W6rр�IH�oT����6�e*��k�ϖ�����y��U_�kl�_EK��E�MK`�M��y���%��w�M(��|���֜�α'8 ƚ4t���6~�4+�'j��9���h��<��kE����n�ױ�9��#�lCU7E�xn�n��P��>x
���m�Ո��֧�X���貖�� +��U�HÉ$�y��hUs�,y*YGG�Ȭ͗9� Me4�O�s�����> �O�wt:�����.�~p.5����ĵ"�EA>:�����N�J~1�8�;�R�nV�J��我G񋛈�O��DO?b�MCJ��L>a@�ji�|�x�=�Z���-��
���?V�p���0����~Ӹ��c�]��H�g_�s���\����WV�����ey��o`����6��A	���=��,��'D��BMRgI�W213:oV!�,���3�-�����I
��Y`���TX�ӑ�����\�hɤ8[&;��Dd��$�Z�ř�E�60�K����9�j���lt,��탕>1cbD�>��`���ԼR��I��a��5ȥ���Ƅ�]r߶�Q�u�����uSl��b������Aao�L�E�<�v�f�ZЎ]�h��(�?���v
t�"|�K�>nn��1%k���E ������-��7\��G��!8��-ג���t������|&*��2٨��'�uz/5�q�y�"� ���O�%�43�~�4�ZI��1�'�_E����3ie	 ��3!`A�IX5� ��E��?�P�!&���6RV=ωy�2�g�E�Έ�½���}�S矾���6-N`�� ���&
�'�CB)@_I
�\=,G�73�z.w�ej�U��c{��(CA�����M1BF_U���5=�gM���+L��~FH�J���b���8C�i+&Er�ᴧ/��g�.]��m*�d�կ����mb# v�F�<0,�Lĥ,��q��o����ਹ��Ͳ��B����B�x�&�y:�\�.K��9.�B��]�}�-�m��(��X�S09Ч�l�(v���;[�=��KDt+�9�ej�������S�)f�#�W��2�]|:������L
$���������h]�,���.a�|(��3{wS� �����8t�RN�հ	�) ��(�o�_�-�:mҁ_���mF�������ZhԴ��>����4�Qd��f�j�HƑ�\��z��
go�ȑa��PN���eǋKr�?��%��C(y�e�7���F�0��l���krbO�^.����v�U}O�q�0�L@ D�b� �S�������xx,�[A�}����r`��x�Ҧ�G��i�fC��wk�l�ڄ�7ra��3��9Q^��"�4�žH�e�At��5c�saU`���9�LI6�Bwɿ!��R�|ft_ۊ+�,p)l7�l% ����ȇ#�gY�(п���V1�/ [�K�NY��K}�����E~lB�:��yאWa�,��E��d��$g��M�k�6���^�.�@�ɇ��Ȗ�v���iڝ5���lf�H<o��ٗ�����_�.v��6��(�ȕ��F~�#
 ���C���g�O��ɢ��Y���l�T}�L/�2�A� �3.>�ꡝ�`�&��LWn�9Ó,ସM��n�)�D� �n��.�������XؔȞ4�qe� WW���Kf�"����3apmu�9�陪�1��g��b� ����-X��v���5��p����#�գ�@���Zq%�kߐ���Q����EG�����]eX��1�1��j�$��S������?7���<��
39/�и�Z�t��!X:߂?a�5�,f��2��L����=a���n$�L1$Y.�o<0���Y�E<�q��T3�XZ�7��XԤf�8�K�*�5/�&�`uN5�� �$�lr��@�bdc?�y�{�c���׾�p7�z3��+��~�m���J��h��9�?Fpr��bJ!6'�R2#.�l�K������m�4=f�
o@8~�X�����\��W&>iE�a�˘�v��|u�Y�t]
��~壇��T7'ao��þ5��͗�Jxb/���¸�1feWӉ��Y�f�;��]BEx"Ҹ8*䗈�O�hC��Q�]+��D��>�P�(~��d�Nu�¾�I-���_�.Sz��Yė�Íګ=��hK3���=\x�U��Y��0�+a��o�A?�M�%�$�!��|B�.���WG��6ר�$>��B��fFr�ôFϟ�$!>�M��ӃO�K|@D2f�/��9~��kG}��k2�A�?J��%�b���tL�H��_�1��^��+[@>f��Zؚg��7/OP�XP������ �J�����څ;h���¼�s�IVN��OT��׾�2�5�kބ5#"�ǡ�&��ސ>d�:e�$�_RP��o��o����vMZ7�֮)�<�B/�eI�¶~���@���	�q0�pN��c��L��@Ӎ��TR�=@�1%J� �[X�d��h�؃H�$k�D
���t1K�u^*���q���ze0;��2N�[&��q�Gѫ�G��B�]`���%b���Ȥ�sdH�wقs���lm��D6��NP#{{�UI�|� ��*�!78D�yJ^s�Mh&�Țc�`Yc�$�	ږZ�����qsM)���u�duO�2�8K4���/�^f�u*��a�Cy���8�#>\�{����
0�;��m#QSl��@��}��W�vVS���!�K	�r�0�ϊ���m�~���7�����"r=��Y�\��(&jd���h���ssW1��u�kl4ԭ�10I�����$�ϴ��P���.Yk?-|<Z�@Fs8���G��\���=�+!$��YP7��t&(���w0�<��X�%H��4���$0cy;{�w�ܵ��OV��<}�я>���$Ȯn�|Px��η�5�8MG�d��T�Ծ�����0u�-'�E�*�����!�*0��km�)�L�����7���Qt�Q�:J(���B;Qñ{���%���5�1�C\'W�9����F�d�Ȍ����lL��_�.�x�p'ĐP��=8�Q��o�fj�R��	���iݕ�.`��CX���Fσ��ܠdT.x��JMa�䞗�[-���Q��W�!�2�ˤ�f�7r��O���l��^���R�ip#�
��k`kG�b\��CS�pf���Z�ņ4"�\�H�$��u?��Y}Z���^�|$]E� �V��J$��gz�e5뿄��Gぱ�⇄U������<�R�Ws5 ��4��䖛�~}�Mt�W)X0Q,�.ŋ��e�i�IJ�&�f\C!�W�M��գvW�ق��Ѯ D`&� �WP"[�`=��Т���1/˵�̗���	����N�9Լ�� ��Fy����%�I.��s@)E����K^)KFZ-ߘ�_��i��� ͹���tz�/�_} ��p��W\��f|�T8M�B��F>���_��Ή�o���~m�5��c�$�l��&\��\�?0�yO���s\96�K~?�	H�[�@��}�A9:���u�.M漎C}��j[�;�tBw0KL1-��Y���ê��XA�y�N�&�X2���Qi	�qd�<��r���J�V���G��?W�q/%��'��R�S�Y�9Y5�f�����;��(��ǎ�&�7y�-Cʦb���R�cΎ'�Ei��~'�-d~��M��N��wuI�0r�:���>:���x��K�4�����^�79�$z�!\j6�<]V���MJ.<��ZV�CN\��&o
 C萎�	�mt�f-e�m�����	�8���b�PM�\"��i�W��v�����V��� Oӈ9j�f��0;c�����ƨ��-.�rM���C^���z|�.�H@7�{P� �\T�.�`Ǡ5��pF,�oQ#����8�� �,w�̈���{�K����qfЉ�\��y���}"vx?����kf9�!�ާ�����E�1P|�\�4�{��.�7������v=N:Dy�C�H�j/e���7�����i�*��Ӕ�4�钜���J���G!s�\�X�8�R�K�ކ���#���%ٺ�D�H���W�=�%c��H}+����X̏�[=`i�I��jh���p���#-�VB�65�yq(c�U�G�7�6�2 e��o�eHjd�闕a�^�u�\��Y^�XX���Z�t��?#�Ȑ�J(���{]E�h2c:u-���ͩ�6��R�\ad>���]���feWX'�g���F�+���VϏ�L�_ �[����*���@C�4���O�ɯ��b�wA	V��.'��ud�K}"��:$f�؉��մW<�I5nG���{9���s�X�v�/��2��Mζ���	��ʔ�\�O|A�jQ�"��΍t������#�5�H1S!�6D"���c�s� �FY�Lw���>�/�|e)Apjk�Qǋ�UBm����o���Eӊ ��~n�Ө�-��#�=u�Fhr&�w��}�QZEq) �!�à�hߴ�A�u����N� T}{tE�X��8a�g�F�� О	/�F%+5�#�|��}������.��#YO%�d��Xn49%�'㽥���Lm��[�<�`v>p��[X�{n���T玃¿ֹ��w�<0�&��zʷ�_�)���A�T�����[N�~G�'t��h���(��^Զ1N��Ӻ/�;�������Hrp�O�ыYo'��]�Q�"`AÛm�`]ai�t��v���L�6 �κ%�����(��r�D�Ɣ͔Cx��=�G������G(��./�{�W��7����v���uK�bO���/U#���X�KZ���p9�Ov��l0��d��+v�E ��/�Z��2ŗ��e�,��?T�R�j7N}yyi˿�c���S�[��*;O:h�+$�Qޭ��V�	��@h���+j�[��uW�o5*�����-����ۢ�"�ب�ɖX�t���֓��wcI��o8��`C���n�6��S�=�K�v��X�o�E:�0Q�ά�:9ύ5�!�E�F�`����L0�K�9�j�sa�+��#MY��Rs�^�S�ߢ0�㤷'd�dߌP���I�;�U�Y������v�Y`o������s(�7��`#1���bV�ޫ�7��_�F����AU��=e�"�ɧ;sI\I/�=�w)�U�ܨ-�lYk�N1�/�k���v/x�� x��h��s��pxr������k�\p�x.\�*��9X۝�(K�y���^�س	�b��o'=\S�nl�KΣ<Y���L*u��F�4�u���m]\a��<�ډ����}����2@R<֚3��{g�6;����x�ͅ�|L���#�ϋ���g+��o3?)7���jI������	�R
9�
���Y�������)JU�7kUl��PC����r�bH�3K�U��۬d늍���95�^i�o�[�ޑ܀�ke�#��"{���� �u裩T�C'�i}����xS�_ީ���ij��mؐ6cR���v�(H����DSW�'cg����MU���˶ꨄ�Ř�32���v�,_X%����#[�!Tꅍ�0������\Sƒn��G�W��h��u��OT�R"��w��- j�<Dt�W0�m�c�iA�;5��K���ǯX����rI\s�M�'	����C��)ԁ	���t�Q�>��-�کV�mPc���5Y��p| �%$���F�^ʴe��?˰�t�P�5�u����u���J��v�o߮鐽�0Z0p�����8��N~�ٗ�ܚN�)|�G��C���3� Əs���PSF�]z�>W�����1�)O��?�r�v��:�
p�����f�މ8��<X���+�~��$/[���¹�_�,<[s���X+����x+}�"���ۅ�]�@]���0�' ���P�	�e��4�(:��w�V�ܥ� ��M0!��z�81\��T�~��$��	+K���m]F��`1p'��#���l�J/@l�J֞+�MU/M��=�_���X�$@��<������B=�!�H�����pRB�m���b�CDGh�@8��=���V���}#M�h=��V�����_^�܂���Z:�r6�(ߨ��;�`�K����_���X�����-��8k˪ܛ�۵a�u���|?��a�\w�; �i��G������m�\+N���8Y4o�� `���V��Y�� �7nW.�|���c\��9�Uw�j�^���O�W�l�ϵ����x���8!C�J���>ZY'�D���~¸C����'������4�O����!yw�U�x��Y������O&	�X���멸��+���?�!�=D�Ia±���P]�v�&g�;��O���`A���٪qdiʙ;�G�p�����⃟�7��x���a�)c�`k������\�G�.^e�g��'!�뒡6�����0����$\m� ����a[>}����e�/H�5y%{bH`'\<�N"y�c��q^"8)F����p�bE}��k�_��u���տA�M{(\m!�w�eu��ʐJݦ:Oo���gk=8�Bޙ7a��;^�Y��������S�@O!c�n��۬�<��r2)Al��j�I�s��-g�����#܋�,v����Z���sx����-Q�lE�%ƉP�d���^�x|8�OiB�iV��Y�n=�i�<�:X\��?�v�r�����J)���[�29���G��i�&"OZ���j�!��-�J���J�U1w���6����D��|�.�����vW�P�n���R�%I�x���KmBw�Y��S������,�'M��mQ|}#���î�1j��8?m�,l'�� �u��5�U�`KX��*]S����:�=\����͓��8����$2��1��J�ۦQR��)Ĥ� + `���]O��s�e4���$��� �K%��|�ՄG�=��s���&���;����!zDHݷ7O@1��;z��)-l�}`͐��#0p?ճ1:��i�ˤiH>�s��<�Y�C�,'��r�a�y%�~�Ҏ����HE�tNg,Қa��qd}P�@ϕq�|��Y�A�\VLB��*qi�%���"d_�V�T/��bĝȸ�t����Vj��R?F�AN�w���k�9�W ����{=F���}u��C}�@~zC71���G-�٣�py>�!�-t{�dۇԏ���'�^ky=e��o�N@����
�L�?/�"�6X)Ȯ�tA���t��w�q1��*u-4cP���Ta}P�q;�������O��Tp~�r�<Yv7��i�ߍ�p���QoXyc���a����Ks��AC����Q�V�i[E��j��&H�nu�Z�⪴DYV��N����s����d��5Ǐ���Q�4�����H̩
�tF���?����E ����wt]�·���s�i;~V ��oI�Uw����JNTl2OIl|*η�@�9�MK(�I/xoc�^�e}z��� ]�5�X�W�J����+�~�h�e4����D��8���`�>�T=V���3)���CI8��{m6���S��@y��Nڟe�2ԧ���.xF;:�"��(`�k��K\��'j��}�A[�8��ȉ*cd���>0!����� �4��o!I�^z�	e�G�v1�C6�
��#���GY6�+E� �dd5
 �֍���6p��?A�z����P�9�s�v����d`Fyd�۳C��RG��-V�b5�� �/��b��i���Qy1-Z�1̆���߷M  ��,[�6)��1�F-v����C�:�9�}������j��h=dm�W�&?fEՏbj0_��/��Cy<�I��U�K�;����z�a�U.8Dq��ʻL����t�9�����ܰ�:���-wr��s	A?��\��sjE�)��������,�L�4��c��2�(�����0��(��S=�eJ�3x��{��<�3�	����w6�o�ٽ̄r��z�B_�.̡�G�ÛGt�`�w�%��>f��	k�2=Fs�uL��H�j%5Qj��B���>r���Nf��9��^�������Bc��4(�l�6�dr*�T[@~Z�8���b*�[�@�.'��SU�4T�>�Y	5�m��{�py��*���vå�f`E*兛OHF���f�0�k��cF��~co�s���g/C~�+�c8���2 7�eAcς�API `��I�D�e6��	����N������Y��`���Q��8��yǈ�M�W�z2�~�7w^�����I�0��9��cL���������ͷ `S���u���i�r��ln���J6wE��i����z���2�y��tO��Ê��Q�P���M�c?�Z�=п��߈)-����Y���&"�d��.Cn��vtF�cĵ��Yj�Rݣ����0���/v�%u`$���Ş>ă�Ko]3�������֍�hPG��'���J��t���03��R��K,�N���4i��+���gZz\�l4a�$��,	���T9�y��b�}r��E��L�10Vy�q؃�=#48�Y�VHG���k[k�TsI��a�,C�7o�4e���8��X٠�>���l2{�@D��L��di77��lT�ٓ��C�K�y!�a}P���58f[�j$9��z��A;.OWŠ��"��͸k����j.��
b��ܜB���Ŏ�� �i�y�פ�.���@������ۮ���z *��n����()h+��^s&1��] ��W�5\�\;I7e&0F�mWZq�K��佑�u4O��\6��-�VYئE񟗤���:�5�j��H?<�ʴ^6s��'���ٚ�������m$N%��f�i���}dȖ�Z�Џ0#�Ũ�x#�=���>� H�J���	JsW��Ih�'Łݨ0М���p�쭾����r� �{3=&|#���H���gM~{X��d6>�	�?QX�9�C�=}dF<;=T^�BjǡEA�A�R�u��Z�������+a�j(�=�l�4e�Q�`�$��iQZ�ȱ�� �[���Z���������� P��f/EMn2�N-�kS�x7� ��HE��^���TH@���(�w�Z�g얎��e�6\&�VV�0h�V�'#_6:�\�	z�����d�ex��=4*�&Q�7��IH?���$t��E�L�p�Y2$/�CuT�)��se(��0��<� ����.O��vST����m��5�F[��7rH�H�ͯ�PQ�*]IfmW���0�H�Ytg��YOʵռp�K���śo�E9}8
cW��=�o�RJ%�$H.g��=t�vG�E�W�3A�ף��������3����D��~8u���X�XL���p���+*�� T����*���2����b��
���!1Pl���+��'��-U�1=���ͧ[?�YA����{�R����-"�I�ٔd�'�fΕ�M�rSTʥ�V	���b��tDo�M��N}�4geg�x��(ՍryO���і�?��׺�C�t�pu�/�,^qDl��8�y~������+����xE2�5I<���9����Q`Řw������)B��1b8�/6�&�M]�����g�h[z�������-��5���@_��c��z�D�Tevp�j��|$?�[d�F�z$!��8����'q����$��V^,��]Ê�����C�_����9ғ|j�I�R�1�7���^�7����z�<�#s�~���~�����Ϡ��ÒrӘ3�xj�� M5$�	XB$�~��	Jaw�A�S��j]��Z��?�Cٱـ?O����ڼ��*���i�Q/�Ys�b���l�r�U��������ا�?����2�7cH=-�C�)�c&�q����l���?b����%Zj)���B�8��H����ZO�Y5 �a,o�4���(��a7�ؼ�Ody�0Fy�L%+б���1�SʧK �u)�|���7�6q��R��ؾh�hdA�6ׯ/���nid��C���垳�(F?��`՚X�\�9�
;��꾄B��̩z�3���b�l���5%���Z�¹C!���MŘ*Ԋ1�:�z�|�i_�il� ���[d5�Sua��W�Q�n�=�Ϩ,k�g�^�U�����x��1�Ǔ�����y-�4߃B� ��V�1Ȁ6e��H��@)��Xw�cVD�BM���19Fw�W�d�i?�l��^��7��5�=B7�Q�fyG>��|^r��ܧ_pm�^mޱ 3sP�!5t^�:~/G}�arP�b��"��et��#����Y(��1�����!h�{c�����O͜��d��u^F��.���޶�ٴ/��۽]��`I� ��X�6�ن�
����H(uP��PF����`O�_'���qF勀м��0d�~rj�]+��̃Z^�s��$�ƈ.�5)����],I��V,g-5�Z�rvqw�ݴk�SEc�}78������$�I���5�������p��uxљ��׍�(�y����2��ņ��A�;��k�s��������}�ĭg�%^�kn�u����͙�2�I�^�Ÿ�o��`E��g��2�[^�e���]&q���U�Ĕ.�SL�Kq�~@�ͬ���ݔ*���F��1D�!KQ�15?�b��
��Ȇ�{J�/�I�'6	�l@)��F��(��� q#�A�Q�(�J�S�K2����A��Dx4��I�Q�yU�>s��a<�>+�WA�5�EOrvW��&�(gbϋE�u�L�UP�*�4��\�H��wy�Oǯ�u��m��ø��K*�=Y�A�x�7����aш�M�|
�t�y����7h/]���A�3|����˖�Ēy*:��NZ��/��Eڻ ~�����&�/\���3�Ȅo�����&���Y���� ڶ���RDa���~õ��06T[I���;"��Z��n���� _�8�ӆ��S�۠�0���*��֨S�d���qV1����r#�Ĝ���آ�'�`��c�
7eo��Tĭw�6R��@&� I#e���WLak�T�PfMH�\����X�HzT���ǥ�p�ʤ��㼄�~94���P �a�X��ay>���!f���&��"p�bk��)��NP��v*��t��:���ݍ�F���s�mpu.�5��͚o�?� 0�c��D�~�ۂ�k`|h�	�9z��J��^���t@"�J�Lx�����ݏޠ{�m� [��#mlɊ,<B�Q��F�P�u����	u�ߴʾ��o4D{Q���(����rsz�hcxDe�}>��:y.�ܛ���j�0=�D� �+��R�0��o[�XN/�tO�lHڧW�ȉ��ʅ����{�#��&��7���jR+���9���������OC1%10k��;���7��.�f
=��\��{��X��b͖�3<�z`$ƀ�ص�m�1�F����i1������A�4񡸹��R�w{5�Tͤ&�̤d3M;����@�8��?�0��l����ZrQ��1f:
UeL��q�'Q��#޴&�I/����椛8ܬ8�y�eL92�,4ǜݜP�M����-g�D,/�F�П�U�_��a�IǼ�i:�+2��r�VMM.f�W/�(�>v*s�	S����0�������T��
f��&MJ]�$�B�����;Ū	x��:M��WѤ��Y�Ȧq�7���9���P������*�n̲,����1��g�� P���?�a���}��6e��˨-�`H]s�4n�u����%wr�K�.R=3���D����ۊ`��W��p��+ a��	�!Ë0�����o�����j?�Ti��Q������,����u܁���wL�0��'{�G�+�Ty�ޢ{x��		&�����:����\��m\��������������][nFqg:y'�i,k�����Jo%��&��p��aXg����&(�^	��x<dq	}&�,K�=�O���#S��D1���7q/q!�FI��qN�fbW&P�y�v�_\���V���V$pd��)e�<�?�dDh�؏&ޙt_�t�h`�]��4��b��L��q��.�K����^`Ey�Г%�Sr�)�g�^����Y�RE�F�a!:B�)��jE��7���8�$��<��R��ė�բh|�#�;-����iXz�%�ڶ�#��D�c]�m�i�#�6�� $�F(��¼wH=������ ��Sm?���h�gUq� _�������t~�
�g1��
�kaCv�+~@��.?Z�A����L�>5��7���Q��B"�4a7�JGXB+��DۂfA�CH�b��	�<ŝz�g8�,��w6������g�R�9�P#l��M���ȵN���G��z��:��X�NL��_��y�����Kusv'�f�s"J��e�b��X^�>�8uB� �a<�3�ɰ�o�F�*q�J�7~^�\�v��ʠ4�����|.xݟS�����7%�,��O��I�H��x��~zd^��t��A8�:؃�E��]��E(�wj����r�����ڦ_+���=XC��o�����\�0h6�;�T8��r�2Cՠ�&�)�x��֙����b�=gh���a���q��:�w��x���٬`�>ͷ��}��m����p=j�M�FZ����SM�p�p'#T��j���h�5����v�_N#��;�s����Ә�*�������2ę�^r����@�.�s3��,��F*�>C���2�2eNU}k�k�:� 8 _�?f��s�P^aPA3t����Z�x�>�k{H�s�sK?��� !`�z�)�ɓ�8��Omj���Ɩ>��i<[S9+..=�\� �ύ�R+.H� J�n(�{t�8T�{�bk��F��<��"��@1� �ƻ_ޗ?���ʔm�'�C��=Oµs^�