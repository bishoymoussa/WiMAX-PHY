-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
xZs+415v5lLSXTBo71NHiRbtXbWMj/THFp9ZHrlce3Zed3cVoA36r74P3xvTniAzZN172oXHT2C6
WYMOXC6SjR3qSEMilzUuMreJC9ICQh8WY923KHvbfMqDsf2e3kGRbtePkFu0m2goNmOVPy8cJjUP
IaKWs2K04Bjqt43QFNl9WzxN0agXL+sWfpkCN9K9AqgAkKmxF4uokQYvwyAI0qdR15u22G+iNCGa
D2ro2jP71rFmjPvJubVk4eMX5/GBsXB5LDFh9RSVFb28aUbmMjP2hYN3aaoF7kGR31Lx3BvGWuPg
m04ZF1DkMSxK8N4YBVbogloZtGbqSkpIVVZ+CQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6208)
`protect data_block
FbUU8eQhkH2cNr91c4qLTJ7y1TftJWTHX/t0bRaeClIlPIMOhmVxxHBlmmlBzNLjDhkVViJZ7uHc
JEpu+OM2WyOqa+E9S5XkKZoDFz18oMW05S08mbOJ9YB+zd9TEiKQW7L+Vswsl7eBrcsm2KxOrrEm
FajRECbdN3UEiSuye5GuT6SMs1fkvcAbOaE12NAKgNzGGHy+VFJpq/rfUgP7pKexKU1vUKZblYO7
Qbc0BNrm+6UmHh47I+P6+Oc4Qz+ODTXYwSKGUjMqi1FT+yaDStaCvrltFipnQy12oI4cdSSHh5PG
qSkZU+tkILR+H5CQT6fNjptd72OJNLv7Va7s5hE4qmgUtv3FRNXAVBdDuVQU799xuJTxXMUJApYD
XOZzHK3qbYsq2Qsg4oezJCV8cmXG0BMAJJMZHH/hF+6rF+ooS2S+/3a7ANRlBtvKIGT/PH8TkBMu
wNZLCeWqKsTDTTHWuS+KIlgA7q0PWIsEWm8SWJ8cBh/KCVYxRPNXlxcw0qFAEciTHoFIiX7vtPcA
I+2QzfDz1N78Jh2oyUKsJ5bYQM/LLjuRWFNNxvUXXORzHn2NyL1v5NnP+eCiv6KM75JPj17CH+QU
x2tkTzVFsnYp2J/Eo9TYjofUWW1WeaDQgNFyDAOjvuB7SqUnDoqjIZhqZAKgd13VuwEXPKc3Pf67
fhS4kPVhyn0Tl0HhP7bUzkhFq37CjzMNP0QdJIdZ6jbX/6lLQBCto55yXisC4Q5tp0xVF/r6cmir
ihpWj67EPmDo3qwsz9cSJJnwYxidatukf3G4lqQEwES/0TXpT1OBlcCsrEcPkpERT3lkmhlRktze
D8Cb2XODfYlcHEtonmZK4vIHXoYLXuylBLXVGc4s1zJPhxcY7bN4npe6B/Q8ur5OaTv7ApVQx7gB
9Fqb0jAOfLzoGWClUzBOkt1Z3DMYPLj2edVoJ7hsmIUr50dYP1vb4F3Orda4wCnfb4HGnBx6aNUE
ABtYe49Z7J+oKUEGL5oJ4RFoCxm+2jbKJ+707ET8y4CMkPk4G8OPROefGk+Ehq0ui1JX2a08dal7
nwko4zdCpf0HADv+jZjdSQCmtUy59bz5X1Bd74YocQ08C7ZpM0LWXpQ9BylN2+L4ZwKqEsoxYlwt
HloEFiHKFgqf/n/dTLIB9+BcyxsT6EdNOoNZtxQmLqQBoj9+8FeFIDkieUXSuIH3EZVSLMYtOAjF
EMGKTic2Og4zCVTo4t+ThVXftSbfg3oaJjxsk8gNkZfsAREq5yTjCOqRLec//SZkylNtL1ZghgqW
L/lKDOPSqpPvO4ZyR6aM8YvO2YyYNUVT/05vn9xw5hcf8ftu4Xov8FsjDDy6swWLAwAkiQc8vkmE
7K1tyDMSWl8MmHrEQ97IqGHVFhDqaZ26xz2h3nQgm576z0JD+mvapdv7KezR6PRcqpf+9Z2/h1Lu
poxc+eFERPiFYcqQclthYqUIm016LVvz0OKBIuf5TE/LOQwMwKuaqxnvhgJe3zQp/yBpsu0Tdqui
nnfr7Zfa5QpPRkCfC57bCLPLe33JFouhJJhii2ODLdg8Q827gcnMcNScuwcSw9DLMB9t3wfb4fSX
GW54xeuogGzMSZMkSCzf7AkRmYILP871mEp5P+bn/ZcAyyw3O6xoRLiL9FvSmyYEOOwfjoMLOuY4
VVXbHV1HQhY4wZl22akk41ON+hOHPJvsAHjkXwhehw6jy0bNfT9KiLGHclwF4WjES0ap/UMmnG53
Jxppg6JwPHIrMkKMwwCHby4PY9vkmkXExRH3+pnUZ/ivDTwGn2lXAM/9Lagqv1D7/RK1tk/h1yEl
FQHzCFj0PpuJe+qlVzQDMu5VpVb9w7jG9B68fDSic5uX19NiTADkfCv8Z4mJ9/18Ti+1XCbRA0Gk
+QXwviiv4HVv61bZiaXl2VRtTXrzvE1pY6OLGw55NYVwPteCcl8Fik/HF2Wc9DwxRvj/R2IuzxCL
hyrm01U5NxR9SqXr34b2Mtzf3/Gy+LbvZeQUP8kIqXuZFWQaYA+hbTwwfwkSbiTHfkAN99x2kv3W
+UxCYtvPipXsPCALZazDzxao19pwu62hXHj18zVWRA3pniSKbQIKuitlekMvZNTg18N9alQn+YC6
M2jgLO4XSguxl/BhGj9m/gyJf2IzlMQISOjmUE73Rn9D3Jr0gdbc6gE0TXE0Ky7Og4W9FiYEtMQ2
EM2Cfzmx1Li9mLYdUOiviJ2egTNWCnN9oYF83eGXuIIZkdvDAw5mDlhaQCjHXi+CUdmT4cgK6Q68
fxBPAORhXhUgBPJttuUgsG4SNd1U4t/aKmWigvsCC2GJ4FXflxus/2br1B6MY2rfJPjbZKB3lyVg
WY1I98oiDSe6CDUiDvs9auf+Cm/44DWVKl3Pb4w5LdPHQDeKK1t2ETj/sSL2hZVpotpwO2cLhD0u
Oym3B5t7cuwwEctAWS3SkmCk6B6WalM3acBWliAWFr/XyF+8DpTY4xULQkanK6Hk4dxwCWgTYev0
cqh0rk7qGBgY90+TPToN4fLcD29X+pT3zB+LejkiAWF5dOh/pnpCuO4yerhlUYW9H1YUGeq/zRO0
glVTrxGqE7gV+v3ac06PLbc2T167qHIdq/R6r9AzOECLklkD0xN6UcBj3I7O6OpWAI9qjO6IKYCU
DBJw/GPQIahs08N/5e+d+fDRpXo+sQEODCASlVGW7XUp7Gci9GeXpSvNk0jkvij38EcyCF1i8U9/
7rDzv6ykW9DdQuFz1CADjqfpa5+gRY9T1eCq0khX4Kyg0+EyfXU4h/IjOpfDotTWK/y5TlGxO877
hT+Z+HUgrtWFUc0Gl6ZpW2L+SJLJ46aMwigEmoEkd+qQxaXXKqSbh/Wk2ciaHDrvmcVyEd4XIfWV
6ZXRXXX5AhUYydkzdy/1cyqnKx0dEEybgLIVnFIYKsJq75Pt9JB7VK/TiQS900Ym86Y8Shoju9s8
HZ68P+RGRY293F5sFXSLCkV1BsLcrD8CXbsIJXk5kLyvQltAlj14aAi7BylJaC2AKjr9UIKD4G6O
klc1v0Y4bJalTKn2gPI8zQwpmEbX3+Kwc0dKqNlYh2PzK5CKSonYcdE6jrgIwXMsrPLPL/RbTyl0
jbA3XkaYHfEFKyx/ptD6ww+Ti8igp0g+vZxux5Lql5LpgsqVg25mxYWikHMy5lKEigJ7lj18x4Li
5kgZkd+yy1pw5jHejbV7wQIDjib0DvsxNgWuuBRx14QK7B9q1PODGBK2RcZPLYydnbLSxfeFOk3R
AYvZ6ANqvwqzEubBdzYuNWs8C6asd7NMJZ7T3jgtQmn3BpGCvnNHM03xJDeEEewFCju2mePKFXsn
WQTZ9xLZyo4Gqds/JKx3ucb2xaQBsXBP28FY7dZH9hkOySXJcrG4Lga3T5nKLp7wKJktG9Ffh95o
5NCeIUv2EJVEkkqq/xk91/4z7WGR7wi3oEZlN5hWnhaXCcZqYFb+YkKSUaLPK2r1AMFUjmSUce6q
oh20yfOcxa7+iMX27qL0BZTpdm2oAYvT2/pRY+v0jzAKhNlcH3slrF/AuccWPWqAge41cKOcAWpc
fyl44b4tJoUIxyoasO+TsYIb1yfT07j5hMK3Nz+NQ/l+aLZE84o1m5vfSC4Q+PHfnd3Kb9ULtC87
Oned39+Lhv9BZBUNkHedRO0ORQZzj6tv0/EiWysfzmsedmyGc97n/NU2fSvya/NJnrguM2m0xLc7
zDqBkWqDYYncN6kDZY6vKP6AdRNbovFtY3JxKqgd5P2bN7d82ikaMU6qQI8UTk+Aqp9tsuR/TpZk
liGdN4Gxh6u5TNhcR6XX1SYVGSI2Zx+4GGMlsWS6FNnk8OcLadQk6K6BmEC8QJuzx2M62Emoqx4O
EpyMddXD4T9suwVxcxTPpG//g3uGVRZgwypLoombsW84kAg7DBCkDGOIEBMMj6mOb5obHk+r1h8d
LPTytNQa7879+KKWqMSD+boFVTDqNQ8kNBL6mRsOuwsURey9LH1NK6cCaqasOq4YSC5MT0omE7LE
IvmKk8xCqbArSG51lsohX0z+v8ZM2TuWjq7EmhHFfhEMR59H/A/UqqeaLFpBaov/GARy2BEoNGwZ
pOESRAaSoJbbkvN7Jwrvl1oAiwHYOcM2+xCzI8ETQYOfrTQRltH5Izo4GOZCW+gxtg/ggPYwliId
0vAWziCn5AcSvVXOiwoQkcC+AhZUpbePmx1lto6txrDZmLwQgjIzLO1AYazhRD6tZNpD2cRiTr9z
FtheTeV9Fcv9s99cyLEpY/M5xTU9nmEI+JpBhgf3e3GvCwwgSOTIT1mPU20YcmZq4qBY5Ko4TvIn
PPzlIlE5/kGCTw0AGoZr9wg3L6i3/nld6bkx634bKbtM+HBPUY+M4o57/T/1q80M1LDG5YZD1/Q7
SxlOXnLbK6Png3Wro4+SfUKZV/OTmuPZcpsRDobjLyQrFxSetjH4aGTvYE6QwksNjAAODmE7pnt0
5JvrnM7pubPo/unV3R8G+Ieju8m14yRzHObqgoWjuEne9r7LNTliZxhI1boos679UsvXxKuH/u7G
0A8/5HZ9SeIGUewZ8CPHWRvqpaix7tw9D2EnGDitzRXU0mfftPLtCw8svFJ60q73J32XPS6Ldl75
KpqNt8a4jv+lV2/stJbNWhw4pv2dNVXFVbtlTXClB/A6ficti7XPiXsmA33DVCM87F41Lf2PGffn
yWfBpV1905cRFnlZupFLr/1iajRaBqhyP0UesQaWZlWuh0arXolyfOBwdGHstI3btb7xrx3D1R1N
5NR54wWI55grnt2c7VhGATY8T4ztlVIb2THqJLJUb6jLCjHZLIWxO5WeGoWKmZ+cjzF3rgnXeWua
3DPEbsn9HLhTPDnPaLK+2hqJd/+/y5JR7MGiy5K6VGl677HlTqkYLx1i7DTU+hGPA4syZ9eE0sAP
c3qylIoJ6bM8DoyFJo3cRbW0gh4RMRDvFj/L9lH8j5nJNo0YCTOI/HJB+j+S74xigNSYDn57QNES
hBlgIlxLFW5GWhbwyy72XSRa2iIfnA6jNaJx+0wbViqENQQwq+dtCwsz0MsQ2X6+9m0Z7EIvVY+O
eJYpb7T7+9J8l0NA1TJk/kgPRho6ZCJd4Rx0iBOtAqx95S8VQ/tmXmayedIoFlSHGX6ARAUbFM2L
ZL/ew1qphKGTlxvHbL/j4TpS9heSVl9vsz/U4Ob2lAV3rwdcnvM3I5tZAj221//NKOCkD2CJnJjk
5Eg5u13d+RLABDjhm2uQjbtUoXD6X2IGc3ioelPeghJnLf738FL7JIi/1FwpTWcswvJhA1zPrtS9
eEu1huLxIi9/wfTS6VHuzx4MbsA3o8WwQNrfIxQ2VCQrodHd47c9JRsXge8DbAs/777ZFakHdX9n
nJ0Wo3Scqvd/QTrs8OXlvA5nEdlPYEjTGlwftK/pvTc0jyHzNB9G6LnYaqktLW/pMzn3h1he5/LT
PzupXroK/rv9xE3aqt6x7RfyCjEI+IH2ZfaKWSQlMh4cJMESRiibIMSG5hww2IVjlSoILBQ7W7xJ
zj4gx6gkbmRmVaOfiNinFJSMD+EULYB6uBD/FHiYCxHJuymD9R8JPc1Cavcax9fLv9WLQ3ZN7LV2
Q8Jqo7APpXy8Fbfn9+bez/av1N0d3y91vrlrL9rypfQ4KpD4SVREVYMBfuOYvxPMKRJIuYRJpPLJ
+/IjFfgt4w8c2ueu6ywLzTJyQjxuDkhb+wTfT9F05zaTRDtPMLr69TIn5yUMPjhj71cx5yBFqk0y
3BQowp6Ax/4MYq+wvH6w5I5A1xL3Dd8ZrCehrfaJZcudhGY0xoKLJMAP6UXCWATWJLruTitsRRSO
1HzJuz2BG/tynQsk70pM/q7lWFLjuFlz9IM6OBe9x/se79pinkgg4rhZJeZew6X8oX+TRXXY6r/s
TNSggCV3ukk0N/58+DOTBqyXk12tBJpbWF/N50pFhj1v6fDY5rL3J4YYyiVYlNTec2rF7/9AzQ1b
gC0crc93IBehamnGtmX6B5dI12DuDGHNt5qg/7e05YQYXuxtEkzPzp2CBkuRv47s5eGEn0FWGqAb
DV6iw+9sNDGINnyIXnYPrPHV6FVWhHeG45lXHLoreucmVoTVmgHvY4dRi6UWt0wighBGUubs4dTo
GU2QbWD5ApFDVy5Z6oZCi3IaTq5ACZdu/aktlpkzla04yIhR+UHRNMXKo4jMBszhpP4fAwIt6kGp
AWW3mqHA0qrKerx3QVzgltitxxn2sjWKdUvWpn1moz/Sa4+pPTSx9ZEBZkzQV7sT+SH23dQqrzYC
bWGeOG2u8mm8/DDF6W1WZRxRApKxAZFwUTP7DxJYgNw29J1UeveI7fzpPXQ+0qMU0yliq5wBUm5J
Yu34SAHzSpLRlXhpOz0zM5yfiX3nskqt/y548SIvMkLUFS2M78yRQLyhpGvnZmb3PwLmIOzItMoi
TSLPrLuBBh7w5EXTm0DN+TLUvCTn+E0WaQwyO5vltlA2Iq/l+MPQpqvqSDkhdZrnSiXNoKkCpCi0
v1f0p5LHajnDuxrHIwY0WSeBGnZa9ARX4YWUTgrUWCk2H8jWdg0tSnjbna3uxq/Bs/jusSzq8N2k
ooTGjvLpavDIkVzjsesAV4PMXn12TjWjv6GFxn/UzgKjHt6g8jpOubolxZBbWTaqR4Qjy1CTkvI1
eiRA3Vk/l1X7nDxYzf/OoHB5qoNd0465EKv8m/sfgKhhK3csoyt9Oy+AhMV9NLDBD79G7CvjpO6e
HJUTvzuLSJ8VxIgPsYpnBBaPRHNNB7DuhB7OG2O78M4WICaASLQ6aGRC7UXufx9O7lA0m4CtmUck
IYty1GPoH10bprf4hWA7MsSqAzUqjxomi4/mDAc/ps0aV85nvAucrv/OA2Q5MZXXeuo4LT0Dqx46
52taczCPLcy9aNV4L9a9PuTQL8PLkvNL2tqq8Bv916SUSnyxnCGGcFTFELqzBAasmw3GZyCmhYPM
aolAJqk0BhGtncx5iZMxLs2Edmm4aefu6f63VV/c1KhZ083BVIBtO+a91cM13/97ZcGqLll+PufV
TVQwhofWNTL13l+gd7JTeLD64jv5SgesBF2wzoF+hgnmp+N6Bm3LDrrATtbk8ZLDBJMqX9ZAJQ97
k/kimgZXEVdrZsWocD/w1tiWy2ngfL/xIF37/WMFVV/2SjbbgT4gu7y7dXIZINHvibX6ujP94KAo
lnHqLvzbde7NdL3s/BzBdoHeWCnpwbTl01cyn0O2r7g+E5wcqmR9TchF6V24G36TGXJ9JiC3hbic
YtOg8aLLlRAzeFhejOGap1wevZjTveIGO7AvbfARmowQpnwUVEiskhX+K5btv3DZGMnZWh7FyiH1
QZ6wuGcopeWHcXDoexGtbudMnwrJhNuwuDXbj4n7SecJzNRBQc2HLLOzCyuhpuQ+tFBMx0moqp5n
1DnMsADf4vXtcx2DdFE3ZmzYFktpAALz1XbMpkMDOxo6dQYt32M62u5wtF8Ly8WBsGDtoTrX6VdT
mIbRTDocWMQW2EuVM2V88VZhe6D/JC7gbVIn3xlVFnybOgApf+4cLqJjt0btypswoy64bdaGMylz
jPc/ZPIEltyz71uSrHME/0QOO2XMdX4kuh4WTXtDtxDjksM/VQ61f/awIVse4745Lzwsx+a0ltKz
q8Bn+n7srlaz4GGcXt9FAsVgI1tohTPgz8WZXJf3WeoSclRe4PYg2nbqXqZzQ91qKdErFWt9UMqO
iSrF7kMrzvOCIErjvZWZooNdQ6TL19WqRRBDCTxkscvdatxRnPSajXpdvPMDdlS9AkUrjwaocZPg
SJEy0Uaih+mjXSw01OSTJGVXwK6wcLH/W3CrKzDNbMuOQzuqcZylJA/Q9nEKVqVXyoeQy/MIE7iQ
8uaz73ZXwdArx4fYWOLmfjhLtah2PMxcne3Gn8ivAH5W18VtEGOuzLNsHjmJ6CQhDoXA2eYujVzF
78x2mOPeZja+v+zPZBqgNpY1GAnQ6A7syb6FZSaXf+AdsStMORIo0CPOnjdiY4mZtCFLMFTqayrE
RvVJduOxywdDBQkfA9JhEbeVO+7sDPAIqiQfTU1JEC8jXJCRpamkYFW8+ChkSgHK7bgcZ0j2j5SO
27j4nltrbOR2PdHUjGLWoJd2Qu8tG0A03PyYCtVjiea/y1QPT/cqzn9sxxNtUJLSIZsSVcAbl7b9
suLRwEs4lzO2bgAyP5P6NNwIexEjl/uASogLzzWNz46B2ZrJMpf2xao5taTsYkWRgxtU6w==
`protect end_protected
