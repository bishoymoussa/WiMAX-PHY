��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$Rx�y�<��wA�*;�x���@�̦�W�X�fa�M-$u����n~�%���P�$��W��kYَ���P7�?UMfT��q�6�U��k�>����~�\N�(�����X�e���/6U|)�X2pF�]$h���d.���9E�	�IN�f"�\��e�z�y�b�����Oo2�?�qˁ'�͜k-�K�P|����y:����3�l�d���bl��ˢ_�d���kx�rq�mh�MذM�`aS�.�DW�mS�9���Y��+�>��!��!�T�uOB���,��\L�7m�O��W���6����'���j)n_�I����2:��$�K�2�Sʫ��l ��!���{�l����.�j4�	��很�̢=�����N��s���s5���_�R�>����ТP .W;������	�"�מԫ�����]�#7@O+?�⡾�Ԫ���e�O�\A�	�ͼ���ƹ�d�	@�nQ˰��E؁Bf���|D_�%au�-�'���w�*%��"AM$w�*�?ZxC!M*�l-ܵ\ka�2d�eA���q�y7�
8�8���0'lĵDJ�qC�i�5�A��nS7�$�3�kSQ՞F�U%O�_��o�h	��.����ډV�Ɖn�N��
�}���~y�����E�y����#/	ΖcՐ��nQ��-�Ki�1���t���A��0�U�z�]�J��	J��[���f�Es��R���_�֗k��Q���VM#y0 L��)�0���Ah�\��*XHGp�H6ɖ/Q��4�/9�	B���q}�-_h�,��hfPK�u�ӊrf�iܛ!�j��`՟�o-$%1�LGc��o������O���0ߤ�7��Q�7�<}�����(Rk�>���6���V��^@���l��꒞܆�dQ9*"O/�\�LI\��~"(��NA�eO�&���Rlz���'��}&x ��^�G�+��*�F��C������vj�E�>։J٢����&�����EZ�O����]�[5q���I>}YBYr+L��tC�/�+��]�k/=��c��$�����
�1s�o:��lOc�%�����b�}#������^1sJ-�[�c�ؓ�%�/{�uW'̜��ޭ����U����dI�����-R!�_�O�2�;N^u��%N��1wZ�&����?�?T�.����(�
(-Ԍ�^mR�yV��v�~�Rp�Z���\�StH�Rfʼ�1p|7�3~��-,G)Gu}���n���)�^��oJ��[7��^;ݟ�r�������5���7ei�üu��n�aM�^�YR�J��}�A�I�����������,'`��q���߰�R���v@���&J|$g���ͅ��+Q�
s�P�Uu:4����Bo�Tٯ���8~~U 
���׾�K��|���t�<�t��%Ľ��p\]���|+���ܝ�@Ĩ�D�������u=���d����S�V�8�+=�[��4/Oj��m��!,x{�p4��P�C�2=U#�T��^
t��y	��6Ph����7/��<����@�P��v�� )v�6���g�4�N�/�7M8��Ƿ�SR=uE��S� ĳ�w�����u��V����F=�:`�7E>��^�9��-$�m�qK�������`d�q?�A���U�T@�d�*���m��o�?�F�����39��9B[�[�rV�~�Kͱ��]��r";%4������i�&�/���Ô����"R�VX�{��w�{6C'��;�>�(ŬH�y����Nu��IЭ�n�D0�f���~�X-r�߻q�J�D�L���M�����(Ƒwy�}������
�9���71�E��2=����v��W\"EM�(Zd}�2n�1�ro��F:�@z��>��U��/��<�K���t���-���"ZpE�>��(ぐ�ׂ�A3y:R�uj��?�������ԘR���?�,�����}����rIȗμ����y? �0Hf �����4g.ڵ��>�x,�:��}�+0��b=�1H'�}h��;�H^n��Lz�z�f����B��^$�|�y�rV�5�0Vq����ɳ����B�
 ��B��%�ƷS*xz�S`x6}��U@6.�/���0���+(s��RF��Bv��V�I��
�*�:�s���]Uv��G��́Dq�`��oC�c� D%L�	�X�%�&B�B�����,臍���-��V�EfDPӗ��Fo,��"=[�]e1���\�7ɛ�[��"m��֝��	�g{��&�2�MN��h�����;±e
T_q�z�/{ډ�U!7�[W ��L���ÿL�"S"�@@o@oJ8�B��3����D��t��Y?9�p�m �u��e�Lp*a�&���z�3v l���|쐮�_�����D֗�@�Y�B� ܖ����s�F:�G�|be.H�]n=F�6
��K(�3n��e���m3���
�tA���W�ۡ�j�E���j��n�
�$�
���K�6.�nϾ���%��9�����N���s�4�>`A���'���!7H�g
�K�H]&�z�W"�u�p3��c<� �+��:��V������^A)�-'����_>�YZ��\ޥq�<w5����P��+����>�<q�6jb��,>2���h���j絹����'���%�	��Ѿ����`w�GbBC<���	�z�<_h�𥑈��g��������0��f�vu�5m��o	�to��i�m�dJ-sƸf�`eޓa� l�3�lZ�@dո��*�"�a���#����'~ל�y�ȸ�5?w��G�l��fs̔"ScJ�����炂�Y�"��&�ǰ��+�<��gžP����i��!��tG�6�Ӎs��9R[��e��8�$�+J���ȫ|'"��0GQ���4S^}����2nbm�]go�F�z+^l��(�wiX'/����f�<�B6�=��I��0b �U"�~_�C�cx�f���9��|E�}6�z[,Ɉ�#tY�|�I����uX�l��fM�f�
��A��0���m�O��<��~U�[�4��ZXsTN� �&�W"�۳ad�ɇ��!�xMa~�Ⅳ�>���[��:�R��c; G,H���v���dS�rǈq�r��U�p�ʪQ��F��H8W�������@W���픠�OGAI<��5��J�.��Tk�����y�I���-W�aoپ��gN$H�'�ӎџ�1?�-��h�l�h����踖U���H�a�K�hU��I�n�Eޮv����%���D{�s-�'��4�G5����#��B�:�����*��^���~�$� [��I�1��^�@�b8r��}N��J��`8�ȀT������ �e�c:�;��N N|b9��qakS�á�2D��>�M?J�Y,�<�Qt�.J��>f�+����U'�<�<�ׂ[q:%�}����t.ԇVν4��5zy@`��\mMs{��p`�N��!y��I5Ƙ�P�%����z�����wPЇ�є���'͎+��i׶��|��C1�P,���Q���-�~��
"��D���9/;1KHƆ�X�Ǎȋs��	�$�-�k
H���ہSl�=�j�����h<��r�篏Bщ�s�VQ���nŷ
it��6������?Y�z��i�HJ�
�2'���I'9wz"���^yN�4�)���?PַfLD`�-�?���H�6����@^�$�+wNr;�����u��\� �D!�i7�?~�s�I�SP���Bz���Hh��R���AI1Wp(�K��r�.L�Z7ͩr	�D���Vh�)1t�k1�g:���$�G�}�g���9_F����%�v���:�Z�?r��O�m4���~��4�ؓ\k╗쪂�8T��@��S<���3A��t,��(1�{�a� �^$Rkn���Q8��>_��u��iA}�²��Ue?x�=i��U�2x&���Ib\�BÞ�m�g�:�a�F����|������>'���P0��Y�D�iˑ]�'���ʹ��-C.������9�X�_��Հj�۰oIj�=���xEh}xط�@1τ�s$p#{��M}s'9ޏ��Lzu��d�ߗ���)`��������qRv	`�"FA�k�'W�S��R�����`�v�~ԐI� ��3t&�N��vprE�7��y�:�v~%�ש@S��;���ĸ��,uP�M�"�����`������LGa�a�>��;/.��t� xM  6���6g��Te�]��u��Y�`�Yv�i��>S!�C����j�b��Mi�1Z܌s�O3� ��檨��}Г{���d����Q*�Lb2e�{���+�臢�[�k�pE}Hli{�<�;�u���5��k%04VHd׀��i������َ�� 	��8u�D@J��c�)ߤyh[����0P>$k��+��JX*`��So��@@DK���S�Z�l?Z�4+��� ����v�
>G��\�����!T�#�^/~��c���B�P�Jk�.�����f�W�κc�>&RZ�A�]2�Y�ܦ�K��7N����#؇fA����F�� �V��̹��f�r pk���IB�va+_Xv���ba��e��&���@�$z�:�C��<�l��΃	ݤ�[��G|�J�hKF�CcA;�&�n<j=�p�T,��@��8[�@IT������В5`j��"j�� ladd��>�O7����0��B��8D��]G���2��e�C����]d�,��b���S����ť
^r�v6N��𕸺�S)�'����'���V�D��*�nb�^�R��U�i�l��L���<+-yt� �g��t�'�U�z��łl��"V�o�������)��������y���xͨ��Y�I(	7*�΍jO�!G6��W~�ܙ0L���t��	��R61=�����<V(*�3�O�kם�y�t>b�L���ǡw�HgI�J��W� ��9Z� ԣ�N������+aA}�&z��]��E��~�$�Imv�N����UI2O�Tc(�}@}죯w���@����e�xSI�2���1f;�['�~а� I�%:%��ޓH�8�%%�W=�S~`�e�����	�a�H��(���U|D�F�5�iě"f�* =�����md�4�C0�y�ť8fg4>�R�C}�?g^�Agm�5W�� Pm�8�@C1u�{���	���$�����d-ב�_ �Xa�'0�����	$��*y��m p����S�$u
T���;fe��d��E_2����L���*	#Xq���pE'8-đe"K��Q�!z����Dt�Z"i_��ek�Ў�%Or�&Ũ/�+V�%���R]R�`��"@q)�ئRu��?z��W�o��&�����=�.�b�Y�K��yr���T� G�&��e���G� �=�p3����*��`�����:xkB�����1w-���Z�7�9�7+�{�!�J�)��<�SL�~�a���C�P
��*I6���Tj ����E���݁�Ԉ�u��Ll��R��>\^ǈ�����v#���K����[)Џ��05u�g��^du��:ݞ�q`���{���kݼ�*��  ~.�v�n��q��֧Bvܱ�[��+���YLH>g{�?�����rs� �z���l`Dan�.��)T�����!�d;��r�'�GK���o��W9�WF���Z-Pò��1������cx�m��YPx9h�*�F��s�x�=�Ey,PU`OK�DU+�&\���sN0�͌G�M$Ɛ	��co�ȃQ�6�y�,��^j�"�y��,�
�q �q�x]��"2��Y�xW��i�x�l���� &���
;��f�u@�h�{z��r*Y8�<RPg����b�뇀c��8׃g��/��R��Ϸ��K�@��Ǡ{�
{��8ϙ;@�YAg���h{L-�5���Z������Ԩj5R~�q�c��
1�6)
���Y!Mju�ٮ=����d|z���Zg�m��i_�}>����ā��ٖZ��?�e$�.\�S��	)>��e^#��:��)���ە �$�X� r��ṽ���|���w�ۏz~�@�&2���.��K�$���-���$@�&f�6[yx0�;Q�b������҈K�2�f8���=m��"/]��� �!>��bgo�-�*�����;7��C}L�S>�܀��F$٩#�u�U�"�����ޤ�n�fk�,��!3�q���+�K��=T�T�Bnh7�ȣ��u��)4���F�B��'�����^wo��\9�]x@#diI����4��O;k�B�����T�y|g����U��2�wW���A �s����K?�FUY�����_�&�4�v?�˾��n��w����%��	�E�7$%�Rebڏ�뺰U\F��R!�WM��ũkw&��X����|GE`��5��+��V�O�>�c05搒�"���8��d�̤wu�Q�z�C����?�Y��g��!�
]���Hz���N���r#���F�Tʍ=��{䪩�8�~�Ss�CW�σu?_��W��z��~�7Lg�V�J�)Tm��ˑs�z���n���#�l�	b�J���w��|���,�\"Z����Oz��ޓ� ���IЌ��~8���R���f�p�I�PzX� ��`+\�1�����%Mcǉ��T�@ipD*\�%&��z�E�i�)��=��)��y*`[���IƗ�;9��Z�L$�; ,��&�D�3�t�{�������W�LF��J'l��?v�G]��HN4�Q��(��BEQ�w�
0�XK�~�����pVa�>�s�N������F�]������׺6\esy�<�Z��%��k�_X���p�ꮈs��@�cx��J��`�CNn��>���ͬ�J]k�`G.��\�*��-�ՀVD�t#�e�7�4-���~S�j@����_#-�K/�����uI-�v�9Q���|v��ϫ/!�Jx뷫2�VveY��#_R�����3�|��bZ�߯�s����L��:I&�u�r����ϕ����,��
�zڮ*.q�+uD��c 7����U�,#�T9EZ١��ͫ�鏕�X�>�D�޽�YsK��7�k�ǘ=a���y���ǧњ��/��5�}x K"_�ܸ+�4��Q�%-6P���p)f<	�}疡
��[7p������kX8c�؅1S� �kY��$���2aT@�Ξ�/2���3wT߳r��DY���w�g"	�G#���`S�l��{*�I,O��ot	х��?hX�N�����ܽ�6��>+���&���p�XD�:.�L����
�����ҟָ���81~}�����"�ۏ(E�Ւ�f���Ԁ�_���:�����Ar`�wi9��γC�"��� ��W���mK� }.٧�����L�,�V)�Z�g���d�$�{8�C�g�=��`G�����.N������Y���IC�1�?�.y���I?�8ѝW���Y���@B�
��N�C|!�~��7�:hv�Ke�1��^VzJ�čZ�-���ۋ��Hվ�3;c���~w������))貑�Lo���f��7�%��H0N
�1cv��i��i�ӝ{0��&4�@ee��@G�Ne�}�P�0g�3�b�>äi�ì����wӶ]����i��#������y����B�eQ��d��, �
�jG3�tЊH�K��� ��]�s#�Ö%��!�y���̔�?�(�@��z��ǻMv��ES�w@�\=�XИ/v�Z>��~ʦ��BC/WF������pE�8�`p��jb�u�ʚ[��89�� 0��3��'��v�4i��%,��ܾ�ˬ�3?�D-�6?��rA�2ŏn,2B光�����`XS]Ê�����t��S,��*�`��2�@T5E?{fX�����^�Ǜ��eY��Sk���s�`�슔P��MT�9��^�v63�%���
�����ϦgA�{��!�w��2!�e�f�dS�+H��)�2����J&�MX��0=�c����������|"�ޏm���pK �*|8K"lIK��^����������6�̽y��9��E�#���=6>����Z�S��вZ	R��?E�1 ͬm�VjJ��?v7���c���
�8��L�b���%$��Evr¢�釜�$ɪ�3��ԍ3J�l/Z�|m��M�W�џ�ذ�l��Ԭ��gӕ�0��G��e������j�{NR��`�2ϝ���5a;�Z^Kґ1�C���b6��B���>���)�2���J	��H=H�wB���i�x���V=��ވ{ ܺd��mܽ�Tu���cW��9�O��1@Oɓ/���%$W� �tR�a��&f$��X~�Ȧ���&G���0Ot!Ɯ͡���)�29�hi2�EP�Pd��m �.�{�����f��L���Ֆ�?����V|�����miأ���a�{��l�)!.0DC��g�s_%�39�� ՚x��ݡ�x���_�i�8�yJϗ�@����ɦ,@R�ؖ�Ҭٻ6�/�[�4RI��(I������[�v~l�NB��3�MØ��RԲ�h���`\ _�MM���`}(���o������C��a	X�"���F|�<��Of�r�V���9�FwȠ��I��l�]?@��pf�XUP7�b�,����nwQ��@���#X����ַ��'1,3�%�^z��o��E�~5�L��� {Y�(m{����F���	�%g��Oi���oR~�}h��q��I��Wk�6AYCX���A�K�E[w��&�,5���cI���!���x�$U��	���İ/��\l�y����q����/sxf�M8ůB��B.�X�*|��#N�'��r0�ȗ~��Mt�]d2��]^�Wj�2��E����ް�^-5��v�-�]h��/���|�$�*��~f����K���h�J��޽�~���c�{��Fku_I�g�����2�꜠-����M�[�]s�"9ݠ"0����۹�R��
:og$�!{B�͡��d6��]�p�!���O�޾�T*63����&k���`V���P�x��x��1�W7Y��l�
|����0}O prL�#:P0���Q������н�e�pH���D�XC�˴��=�|9bҏ@���͢�Ǆ��XF?���RR{�+ye;"�0��|��Q��zM��ݕ	\�#�������g�M@����H4��Y�9���t�����]r�ZǞ0��Ac	�B���n���3�ߜr8g����e�	_]�2町��;�H7�[�X 8�g��/F����P��w��:��_yi	`�E���?�R�S��/����o��k��,-����ěP++�X�j�MKC�6�ILe�An"B�XW�ұ������jQԬ���%����ю�0{�N�?���K]�Ն�7IqՀ����y�,-P�?|:��^mˍ��B+��sR��+�f��<Ȫ;
F���4��S�':i�)��3Ԫ�P��̯?W�M~oG񨘉(�$F�>i	[�1�y�|QZPZ�ALw�S���mb! P-�դ�d<�f�k�=����u/���=���X�՚>Uc��X����gjE6�c�]��t�B�Ũd9��* j+��D�E�3���}%�L��%,�Y�0���rgG;s����T~B�Gbtztr�7���Ru�- 
�d2(S���u�s�z����>���N���2@VQ"�L���^����4�Mg��FB�|e�D<�	�=�y��kJ6ci����J�ńi�;�k ΌdG7q;��\c�f���d��I�.�[E�$�f{ܴ�ZW�{�-g$�3�������p䛓�bb��Z��]��j'��ٹj!e�Dڞ�����UO����sɌ=�:41��"�Y8	^�Y�P(�?�IR�����b곪F~B��&K�j����%[�j���_���dL�:�ҝf�\`��08�7��/�v[Ԙui[KZO󛋧�w8P�����[�qӼM�[�X؟�Zpۯ��L�f�9��S�RB��>�q ��pj���W�{%w���"����n���0g�}�G�v����+L���� ��a�F���v�� �f���7
��j2f�l��S|�����p#ѻ�Z�!��]e�Іp�}�y��t�C1h<��gu�����f��f�ݥ�A�p\��?�W1��%ݩ�RF��;�9��7,�2��n���F���|���a�f:��-�K?Q��C�_��>2Z�=x��Zamc�Wt�s����YI��7pɺ��&�k�.PO�A��8�7U*��C�X8�����a�bR��� j$&.@ٛx��ȇ�g����[��y�)w0�=�W�,H;��%�2�8-��wr�jB�)�
�]���C{�D����]��T}B��5C��c�m-�;&hN�E<��ʖ̇uȽ�MP���o�}�9�A���p��'�G>������� 4��ЪV���`�m�2HX�*w(8�p1ƨ�P�[�c&�F��Эy�=
�1���;�s�:Zj��	�́���e��p`Ռ~�Ǹ1|嘵�`'��go��D9`}K9Z�@2�U��3[nh�/������p:=�3���.0�ȼ�L�`PeW��n��T��%+����b>� ��\�p�5&��U�5����A�J��Ŝ��",&|�|p���ET����(��HJ�hyK�x;��ƅ���8T:�$�Yf�U���o~�8�	.�<���Bv�	={��X�������5dp��=uҋ�}��E#حK;�`��05�,�m��!���L�X�����VձM
�X�����)�"�if��}K?�}�+�_@��c����WS�#|@�Pqt���{
\$Is.��1>	>�v!Q�?�/��8p��'$�
�ѤJ���B�`�K�d<#���(U\-kj��ý���8��=w"��*� �Hn�[��&�t%ݦ�-N�����M6Ċ����kY�.(}ܞ��`�� �s#���p]:��|����u`i�#D�]�%ӽ���vHtq�5 G�eV�� b�DNƓ�3ݚ}�5�kD�oS��8��8����� ;�7Y���ڰlҋ0��d�)=�����xq�����2�[��FDC1:���`�n����0f�~:g�E���h}�c(����e;G*��B/��{��g�e\��v��S&��F��˖	6�r�;���/�"k�QF��I��5����Q�s�:��
�б�!1�W�f�ݧ�n¿d]��r�q\mFB݉�|p&���#�Gk��3}�'0���k�ז���0.�t�kR�|�|�E�yC6l��v��~�y+r���l�Nm�X���Ҳ�xL<Ɇ;4��1�޺�o��Xj�Ч$��WR��R�^�$Ѝ��!yQ4R���Ft2"�����u D̀��%�cq�DL��,w�*Ā&}��3���;�-�6��l˭��
ǚk��F�ɬ�|F�E�{Ͻu��Ƃ�c��R��U)C���)R�'	�|�KߵӔf��z��M�, ���v+H����u����-K��IK�W5�r��S��OA<Z:ȣ8C�땬����d�/���&�k ����Z�QI�m
����F��?(�Km�O�u"L��ߘ|(��fԧ��$k&;/`ۭF� Y�e��њbH�� >#�Z����q�F:�F�q���h��o@��U�r���@i[h[���ɫ��o���R���)��-#�J�WudM,�\�\��ߨ[O�[����Bq�^�G=�Ø��"�8��ɿT(|ږ[n�h̺6�݄<�Aj�gr�R	�iE�q^)�'��ϋ��]FW �J�!��F�2��L�cǨ��}�0x��"��3ѯ|9���0aK�a�[/�(� f���	�v�@B�^�X�-	`?�OԐ&��ͩ��#�j���k������؟�zkv:���Mh(�p�gq,}��]<���cT��7�3+�˛�S!vM��:�G��\a����X�]�1Ɉ�vD�qa�IjT�9$&`#�1wy���l��o�@q�l�̐�G�F�d������y��^B�"��&/�$5�&�*�V�%j����
�c�n����Mn��Ê3]���J0bh\�K�U�jb���Q������梯 �\�� �o�sٸ��d��GT��v)ո5
�S�9A,��ڸY���[Q:�����dT��?q�!{���u��ndBh�7nz{��C�dSm��L�&�D,������C_�YA�P�I��Y�-ߩ<-q͠�[4Cl>%c��ĵ\ƅѠ�	np�1�`�4�(��J�GK���"�%����8]zI4��,
��W�R��G��#�¯�e�l�Gi�h�}.y7�p{�ˎ�Ƥ�l8� LF��\&#f��6o�p���T�����)������� �˼|�G�ڤ�&@�z�� T�m�m�?D���s���>�iB �H������]�W�<IT��}�G��;�R�T�tdJK ̘mEĊb�o���x�{�g���l�K6l�Uq �@�R�PH�+�>�X� d�<'�	v�e��a[��%�V�z[��8$5E�!ͽ�V9�2.��9��!6��6�'O�da�!3�F�
EmW���9*�.'
�)1�⇷�_ ���B^>�ࣝ"J�B���a
A�Ņ���e\�g���Eyhn�������
��埛ZK�B��A^��=�>7?+@�SL���i�E�4�����5@A5��2�kX�=�SɞJ�b�s�P�B v���haᒧX�a{��\����A���U�+m\ࠦ��e_���]��(?����BH�%�?�ek��3+`r�΄��I'`K �?�;�#��r �B'�½S>+3)����<��N���+�iL�
�*�� ��2s93LE����yyII�����o��oK����;l�W<���� �A��F.�O��r:�<RBq~K�*�y&��F�sK��:	�>]�?R��/Y�F�f��_1�V�L���@o�v<��H�Mͻl �2�v첞�^�xf���D���3n���'B�d��E�]�]N/ɂ����8�Z7��'�H�-LQ'�Jv�&t:b�&����Tz�+�s�N�FSoR��Ve�y��1�ga;�i���� (��q��������_#���x�Yii���iɂ�=(��p)��jd���(*HK��ej�ؓ5��(�^�*�Ġ��wڻ�[��o�bE��O�݉>&��OM��.���n�Z�`
�Ī�;��H2;ח�q YvT�:<�Y4P�Ѿdޢ�w��.LY�8�*�Jd\�G,����_P�/]�o���s�#z ���.���K̆E��v���t�?���l���c��ߦ>�	ز�2���X�Y�db�1۩��2��CT^,��i#�E�)��)2��DЎH���UJ�#�)����դ��jWC�e��(o��O^i7O�ԟ[�	x�m���T�KTB2�#;�kM�8p�a�@qL�/�Ap(�a�U2;P��ϥX�r�`��-F%m�����-�T�v�wϫ���/����ֲ�%���3�)�����Z���Z�p�:o}�6$��X*��GJ���ǧ�#�E�1�k��v�V��M�n���$�W^�(��0[�����ч��P+V�8ȾS��L��y��P�q�8�,�rU���^�:��	�d��=���U-/�W8�c�۰⣳ :�t��$%,	2��iS��3*�W5��٧#Y$(���x�����N��r���h�Z�Bh2L����|�c��|��$|��cxl<���j>�:��I1
�P9����!?�t�=�t�);�I���W�Ӗ�K���;
LeUy�o-?��>�~r����o�_����j�0_X��G#������]�KF�0�'t���rE�e����ǭ�?���$�I.]�O�ᒍ;�;�˲"��_|�zy�Aߏ�Cf弛d���9��i�s�����@�U;�	��բ�)[�7zl�Lr<a��9 �|��5�O���ί��0`H m
�p��]7�-��R\�z�?��f0U4�K�~��遶G�֝�L��w{8�Q�:��m������ΘS�.���r��a%�Nt�r%�d_�?����ub[P;�_tdO�ѮV����+z�P�*��(*\  ��j8v@����%�Ȏ�m�Ύ�x�4��%��6�y����\AڠG�f~�a\Eռ���*#� ZL����[�r���o��H1_�U����:��¯�^!��8��qYg�)XsCS�t�T���(�F�a	x������~Z�kAf��͋WO���q�Ԗ�Wjw!"�j-��@/�Q��w�/[8����~FX~":,��Y���)��f2Ŭ��Fߨ���1���jF�r��';�J��
�mm�U��
C��DqL����e6z�,��X�r�r��9��v;�+�w�+�JQ��ذ Zq��!ؔp�ݒ�����}[҆]^z�~l�~���2��# ���6�M�\s�V��t� Y���Qt�ⷶ�V�`J~�{&b����o���z�%��pI�;)S����ԃ����"�.���
ٸ�ٚ���5�"�ٚ��)����
 P,74�f��9t�R��=��X�`Ǘ��;�C$�"���ձk9׏Ǽm&
Р̱xwTD[IF��o�MT�����˻hk��"�Y��8�'y�$�~�z�Z����`�V����g��5=�^��&VƊ���^��߫���Q;~m�a�^p;b��[�2�Nhh��L;�#ы��L���ӄ��:b~�nc8�q��>�t��E�h���d{�g��Hw���f���L��Z�u(od���O"�]����I29fX>�N��v�M}��l��N>͂�3+�kwTl�*���t�W}���k+9����9O�� �'K���q�c�)D���,���`�oEq-�?���Q+e�] y:)��Tl�(��^�~��w�er7Ҕ�$B˱y�-�V�Ǧ�+)�� @����FY��K0򭾃��h��3Öz��W��H���t�DHh
��f�O/頛42w^@�:�q\�q�*�˝"HBN�(ҟA{��D��F��ږ��n��F�}�1�˚l|��E)v�5��{�'�'r�J��|N,�/.R�B�U��jR	]���lS��`7G�4Yr����)Qʓ�?�x��Àvle�Qgxf��? �S���~ԧ��i	�r>h8��8�i�_�Ȭד�M	J�Y��n_k�s3�7 )�!em�L1<2�%^N�(��),�]V����0Lۈ� �=`lI��D��Sߋ�__A@��~�?��ۮ��H�
ڣT���9g$�Ǿ~Yɼ����,��a&�IoA��iG�7T�;�,ѝ��٪��(_m���
�F#�������}*�2.�s�U��e�G��G��,�K0x�����G�A��0��H�������3�w3�g(�u��M;�	g�� �iA<#N]R���|3�B�)���0v���Ǣǭf���VM�d��T"QRA Ĝh�_��6����1��(�+)��)��Tq'a�i꼩�s A"��㋀.�71d�9��ԓǐ[�Ū�K��sd�/�P]�) �gu��vD�T�^�A�Q�����f���>��;t�I�K��qD�IhK����c]̹M��3O����� b��ˍOe&�L��D
�#څ)*�JRu�&)I�����m���u�0�~<tO�9��*�J�[��ee����a���p����or���ݿ׎	<]k�t��z���6B�r�I�m=��@��8T��H]��h�˥0pv��L�Yg�D���qL>F<�����F�2.��3O�v:�W[��^�	����g�cW�׻�u�DM?RHDG[������3AhrvI�� f�ݯ�}�g��k=d�i> �O�\���C��W$)�=Ҏ��#����GQ����P�ºc������˫�w�O��v`s�����E��$�� �R^����#��%�Su��Q�PC���5.�>+C��8�L�vQE���O������U=��&��!Q8���b�}�l���0��du�ä��Ԡ�ۡ�b���iP���*	c�)��*�>z-��`▜iȺ�C����0!S�=-k�_ξ��T'}N������kx7V�K�4�J�X;�qE|"��Ѻ����Ƅ�m���2iH��KLJ�]R
��Iv�0�uab%:Q��`���a�j������Gb�S_�_ʨ4�.z��)��`� <]A����ZϯZT5 ��d՞,tK ��)Ks�v�-HD>\F�a�b7A|Ex��i���ƷEv���88?�N�	q`�22�5K�ޮ�c��$r�Ia��~�?\�2P����]q�l)�4 EG�k�8�QZ�;ў¿��#�P@Y�b)��)�=X@+�lq(�wM���*�L�_��oL<d��4&���_%p;��f����ƯdY�E��i��Ցߠ�Z&U hk|����s��87�9�>i��_I��3��x<¯b�S?[�E�`U�4)�ׄ��-aYM>��ʖ���_�HOH4I�u�����EJ�U�o����#�[�UA���1ag�f����(q���U�[��B��ܨ�Y�9� �vӫ���m��a�$�p3ӌ�i�9��X����.���a����3B��E�┚� r�Ć]��Q-�'&�gI��3e�)����NH
v�#T��A7�T��'Yہ�G�\2VZVE,L�|Y��1��l8�8����o���0Qb��׈h(&+\�m��$�?.JQz���o��XH?*�"��������艳�:�ҍ}����
��O����˛u�a�/�Ȯ�e�ݖ{��-/��n�sv`��ojh��/:â�0���Py=���l���II�j�=��~U���sѸ���\�z�?���P�g��� G��iјFb�[:߿�S��@�Ֆ�=YiDG��d�bǹ��
�ʿ�0�}�]{KP�?BN	��l3T~z�?���w�Aj�Kn�]��K�^��@Þ�8���=�o�<�͔�$~�*߻$V����h3�8%�
&ꃏ�� &�v�7sv�m�艸�Ǹ��'87K���>0��8�~����U����Y��E��=Ь��W>���<j}z�0-Z��X����E�m��24�;�`$��\�-d�u���MϽ�6,��f���JJ��[ud�,�=��&q��#I��vRD�#��ձ�������@�[Ma�yØ����μ����@���l$�& ǣ�I�Mw^��L�B�S�'�CL�� <"� r;�O���f�K��W�pW1b9Ԕ��A�ΒD�a#�պ3P�����E�LR>ӽLo8v�aiL �B�6l:E	W��G����Xd�ُ�o��*C�!�Jaܭk����B�.j�n�,�����������x���
��j�U:{��_�w d��4�"&�г�ZJ?�a'���Hд �P`xl!�������m�� ˻O��@�I$���e\͒�h!�q����RL��=V�TY�'�v���̆ݺ������ǎ,�ğ�!�������\!G^����v
V��E\����D�����P��%��]5���=�8�%F���	�t�톁�U�����>?���9���%�<�s��ߔ��Fȥ0A��t�t8}�ܣ����3�)2,�F����}N!r�M�-�E�`��&f�%�����M6���#���l/�ZOm��i˧�$]�戦��@ߨ>�%�.{�h�c�D�2z�B$h�_�˃y���t9�#@P�_�fYN�վ��I��6�i:UD��>s���d�7	�jL��~�����=.��~a�p��wKR��ϵE
��7/��$lb�S�u�
����������ȬZx3'�[�Dv
L���O�O��k��\rj��ʮ�����j�B+�Νm-#�;�H���r�Ea�\���e�9�8���y̵qi���=�3l�,/��D����ʈ�����Ц��$^a�Z.sّ�>�0���*�
8�=��Qd���M��1�#@�E��|,�Q��ui�Q9"�Kǌu�#����W�M@��0\�`�T�"���֓�V�V���aX���ݻ�-.�d���'8��gb����g�e$g�>��QAG;�o�3�/�B�҈�����ߙ?	���:��p��Qw���Po�ϧK�^%���B�C�Y��LJ��x�_Tjo�Z��kc���7~ō
��q���|V9��CC�}�B�7D��|T��>f�
��׫�梶�+�����/�);����p6�����	�(j.�t;��{�?�)���h��Ų�[ ������m����������%��F�!2^�¤��0�#�>�
���'y���5�%!oљ�~��@Y�:;E�P�7$*�q1r�r�S熞�,�3��`�\w�@3��Kz�#p� Y�~Β��L4�'��C��A%{����MT|8�.�Zy��z+YN����@):Y1��*g*�*��7����^aSj��.��ܔIKJ��*I�y�̗D���J[�V��LV9R���D;���X|6k�?��x��j����$Q��k�U�З�� ���#R�6V�,7j{eǸʲ���R�d��ᙄ�U�Z�`�֐h�����F+v������<R�U<V���Ԣ�Y�v������ά��!�KE��,]�Y�iJ�ƈ�{����ug@A�|$Fpt�`@�Y�9��h��u����_���,��k����g���W���[�� 
��yP/��p'hbGƾ��l��h��żlzƞ�P�z����� �w��#�˩�J��(q�
�P&Yp+ۅ%YtC��.
s�o�:�'���W9ę