-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
hzBZ8Jv0VeYUnGi2qUg5Ao7Ge0yt1j3PvDn8rt44lJfVn1H3ESkN/lEH9AoPCdXqbrb4s4T0Nngb
CZbg81lQlLXTD8BB5UVHiRFlBIVqbx5CF+zjdmfZCJIr8gdRqEkNpx3loyxJ8xQS3gJs4c5uzqm0
ETW8ucr2sIMHQqlNldB+IicGQoR/axicuQ7vZBEps564DKAawwQE2m1NjvacU44SO/bCssXk6FMu
Ydw1LaYpxeK0otPVrS6nlIwfYAShSy2jkpyycoRnpULTWY2dyoDs9LKlQ30MaNYauhk/9/L++J7C
gU5O2Bhe6k1KGCLzSrD1S+iQOCRfgK4cwnAmqw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 10256)
`protect data_block
Ye7MDARxNERH6AdoZImN/i1g5wCSaybVxNM/UuaEXhk9SvdVHJZTF1BaEhzvApJP4AUjnP76BDcm
td7DkD79kCbcq31mhODM7XAYMdpnWXz1Yk4Kin7HrNkTpRfeWp0wYid39H8ZtYyvUYOgeK2JejH+
gqTeTiSb3905rAzWfGFlEo8HzEP6hk6hmtc0KDERlaVlyCnH1KxTc4SEVcJkuN2W3u/RdIKJocjg
Q7hNz8sP0Gr0WhIh37Hbnc+bKXg6RNI/+OXRnFR+tAqGW6sc+TFaVrHp9Fhv+tCK4aanFSSmIUti
oAiba8xNRFtuFBWO5TeJOgsa5MgEVRtJQnCnwxTU6nxXnLevhNL01lifbbzc9ecRoSPE0GcV23YY
Lnn5ElPawvkyOxsLvD5qhhM9kNphMEo2pMRj7eKD44tg4VWqdDvaD9X9BUQ8UJ+SrLgbb423+b1v
JoRVR1HBOTn85UrBGNlxWQ7ofjtW/u2T9ZE3quZK4I+ZhjKu99JpR310LMCwOjjnnZNBVUKPPI5l
YAxO4dVF7jalIhmtvjEGPPChjSl3Kbd/hI6OwdRxuRpE/hUjZ8DS7OHwfxoPY4+d20T8Eyj1zwmV
sLjiEnn3btrdw0Y/RpuP2F61wPaWu1DYgq8a8V4KKv6yg6lH/rdLEZQHUDTMYXEfd/uv8xmgEhiX
AcS3KA0Yw7oMjQwKh8sZ73vhuErlqh0lo2hYbR4EQdQa9mWKpazIPXgwS0FgcBWR8f6N9Ytfq5S/
UOrwv80kPVUbpgMMK9Ih4J4t6z3J2+WlV8FI7qj3/TW44fbuFATe8ydxKeVdoIjg99zn87ngaXTj
liKHvEI5P0jhr3goxOK6KBinzjxrZy0D1ArLCF4LJUMCwYX2KbeX+c6/14TsvDA4Yr2vCc48WVQ9
L6RM0bDuE/KGM0xtIwYN/W3DE3+SJm+mvj9VlSqAq585En2tFBWi8Y8IUpGO11GROhh9Fv7JjCF0
Z9uVaR/R6MhaaVIpF05EL8sJ3zK8IPi/xDZ31DrUASxOboii09JSopZPv22XnrNeCuEyf+sqSSvK
C/5pqPf+mr+FB0y1wtbvxwcJoQbImof6s0ceHZ/QTiGIK8GdtPfeaMTkm6TIIft56lSW4pB+CS48
i6i26ZOV6KJmTFjPfUZTD9JHl+LjCrQQBiwVbz/8bSHYheeP8TTTFhstK8+/nLI2oYMJmgN8IVAR
+uRGwe8ohXdnggdr5Xnx38EguVQ1/78BKC5eC+bCrML6kgoOQaR4G93fdWZVd3hnb20OkBMk18cO
TVmI7u/aUHAiZengaZ6QvXAETTuCUAyki3NQntRWtA02L20D7dxpUHCqx4FcY9Iej99AwfT6ZVJd
OlqOxfJYSxatfWgmqoYafGSUwwvJrKb41zEE4yv2/ZEmAfe5TEUGHZyfLnV03r68Tzis5NhRhd6M
+PJah//OrAFzdWuZ2an4I8c67XOZoI8m08333RHLON+liPEJi+tOaosNyrc761zCmVGsCk60aKDs
gC+JzckTf9r5Pv5s46jWGkEVjHz54VNkTtaT63zyQdVWYdsyHh5gHISXdQ8S3UVptiK5JXoJb/wL
/oj8PuQMekIUF4XUNx2dy+QM/p3CcpChzkr+XdHdTvcBCE+vQ+VlQBATQUME1PcehK1aF9CIfA9R
dxNvywoKu54NcyTRJjC9NkCzeIgob0T6H0QpM3yN9oIyxECkyMZ/KHRlhxdE0SgO7DX4NBNVtDVN
rbzeqzGoBVetPcksL7nKVbAnF3hMN99e8E4asSBN3YRzZG6JNZlKErgF4f8zEV8DBlpSg31Id5da
snhE3/1lGVtQ/7l5nIlS0mHQcH7u/V6b8s1NPVSc+1qPX6914HRrOiVCAU1VqpiDf0MoBVw+5yRX
GT2p+gGJYE/Ek3AJ7tdiauX+KD60tDh6axYcySetKFj7IE4WIgd8vaLxCUCadhUvcktRKhBJPAF4
sc4DWqJfZO65nvgXm56LONIbBQxOLGR2YG0PYebxjqHqNK/zr3wzPDO/2ivb14d1ZsoZu5NZo2hq
rtro3Ndc0zrhG33V8pyWeYowoYujBvbON5Q0hgC9qHrRyFaMJQs54g5aXvoQCF1BLI1HURFmSUHR
tMc1l8ViBKPSJss5qQpw9PVVeJGWJ3AXd11a/WrHP56wXRQmBP29dMs1PiPdE8HYGf9LU/T2ktMN
zw/7oy7rT9GJ+lGoA8G4FEUBeGtkVFP+0oDoyqllTRQe4GYbdkR0rkTSfCZQkAjQ5B0E9G2VTXFI
cDw7z7AKaV7OsYk1WvMxfca/BYcuz0tYxcvkek/NopuUri76Il0zO090e+Dra4DB5Px/VVm6C749
EK/ccvX4cY6khXcTUUtvmSPMaArKUYEAWAF+nKBx3N96iTiLNp449ABcEzafolkPJmUCf5myR7Ac
TABLeCnrbTj+1Hp7KAGLJK41BQUtXVm5E5M2XpqBjsBBaeu8tH13RlQmGNmyvMijMh7D0Dfcvja9
YNKfyU96Z9yogWZCfjvrm24thYQbCH/MDlSqB6EtD/XCHR6GNGkd+13L1GCwvIqGOP+pihyfOqly
wqJFn3tP3yIZ6ForZ6OEfgNNMb7vPw/9VRILcv5qA15NNgyK8o3ujr4NBymqN9kFNEU/JGORemN+
KTZ+SOsuMWTeTwuxRNQvdFlf01J2EB//pj4H3Vogxs5tiHAQwYlV0ZCyWYqh3axCV8kueUQOU7Md
8hGVB78SxjQOE1oUxvFZb55owBZCVbvg0WJ+BzedUjjnMaV8y7F3sR2w3sED1QI3OHkO0Mj4HjUP
e93GbQeM2c8ebznDyOBSnki41JHBP8aZ2LItMBeOGk7uI5vK9My6ISuQPIS997Gnbl757oTrvhzd
sTkzJrzwXjNRgo9PuGcLm+7Pp9lsrQsBcqjS/aInPKKf1PE0D4eNL/8UNBGnWD6IPa3j1bjeDIva
2zOMDmZEWlntChEpnikDXdUpmQGa3RMRSENmF7PF3xMenM+3jNuplK9+kF1kqyZqCduhwqeq981z
L7UNit7YFAfCIMFnpTrwq5NveQJd6pDk9LTyfcJTdpx0vTtDOaH45YVwpktOCnuqB7ZXFwHy+Ujn
YhpjW2X2MuAq9LsIrq2HaL5yMS0qRJ2gSShUCLHn135TYaCaRGVz8XmjTk6V3IQEhsj0bt02QFqB
RDEKg/KKJQ/5W3C+ePZZqmXnjthSg9xQsJla/og8TBKFv1ak4+5DNS/uXo1JhyZHkGul2juDMTj+
2p0o7TnlVUxSQ8oVGUFDaTNG0vnLDuZtIJGKnwUtZ3vYEe35M7ib1BEtSKC1NiPsWYucQKrpGayE
CR7j3m2lPjE6N5cEEc+IXYl+0ZUGq30HS1QF8UYp8hfVo6nKLnl3JR0BAJC6esSSWdiMhDATkWT+
AyiCvX3jwSk5tFTpL/wC3dRy8Y3a0QajsA7WJ43K0IpwKJiGGJOpIpm0WSogomtC3QEIZXxood6y
jwX739uECEEOFpRZN1w8lat22y14ni/SV10zAYzaMF7tYwOdnA5bVYY9wzA1HLf8msdOuDsuxal7
WVxyAAdKx7LBThFIc3dBXuOp2WDZ75lt4uYbPyM+5+0KO4sAHJ+kUtTOH3Es3wwNsJOoH5tXoHea
kfFNkTE7qI4olBMpxOSwdvfijqrbyGr924Q4weE1tTdOxKeoOMUvs61gRoJhfBFpZi1Y0UUNRUki
5/hXRYvt1JlCx0vxUdpB+3ci+cr+BQYWD7njzlKp7QdEjCaWAyWCq/ZFRUanJp+0iRNE49AZBii6
fAcPZtDvxC5cG978FDKX0maGkv2zl45iBNbkIF3O8ClRX5EA0LFiRdT1IWjP2Yd4qmd5MQwFTBQj
cjFjCx50H2nlIKY3p0sxwV5P0s0WKgquTd2iKslhURfNeXaNdV/Jr4+klu8Kt3YD0FTIPGRuaFJ1
uc1GAGFGjinf84oZ7iYy77xFICatGp6MF4PK58OmgA9kA0CtzjbdqxLHf7ZVy8/e/STu8YBG4gY/
8A5A60A7IGA/aYIlS/K9KGllJC5fLb6bH/UuM/+yqMOQo6U5SSGXGC5IgUYWT2IZnALDnaq2xBPz
ztzViatSIC0U6+4wn3ju55vZd6MNooWgBATSEiUGje4lfxF+5lIsKvYG+bCbVbV28ARHiqWdHHy+
3b4mV6Eq30WsnJizXIZJuxRjYVpu0ifqtYDXrBLa1IVZp46EkqD9WQ/D6TA3vhbeJfyydbNE2GdX
OTgvJbQOEBSb5Rw9ATjAHWwrPYJwSlSymsJ8v3hOdq4f3+c4d+4W8WxfX0VihUxmrtpRVQcQ+XXF
8Is/3Q59+HsfrWgBtQL6akCcamMTF1wXWsuCA0g9ULHju2CKMdDI3mJ8xma6Err83LTSSMvxMFII
hGyhJLlKQY+t6iHeIHLv3gStGUaJ0b2zJNsU2GTVKtOcf7b6JFDNc9Xke/pSzOgW+SZIJyiRLUCQ
mTdk+kML52HU1vCFLu3SDDfnOCS7XDFpUyidMO2Yxz8zcnX8JoQr99QphskqSnNeso17sGJMgzCW
QraC8W3t291UwfpwJ2HN+K2KgG+GgakS0KZKe1G4b83EmrnouqcCzR4MshSmDFM6Z9zyzyTJMoac
wBP4K+UOjTw3KZFuJ3IxmF1O1b3Ku0A3dgiVAdRgXQErCUf6PiLl1bg0/4k7lnY97l1wrD5MQ4Wa
M/N9Y/mZzBH64eY8Q2NfPKuxqccrmTRFAA/xpHfX60AVNHuc+ja9VIx8m4akWXu6W97gwtBGxNvz
LHPVDxUTkiJeHfKLEFjogATFe44Ng4AXypXPxrl6+XPtRSOG26RZbOyLlypw0zk/XOTn4rPMyGQC
EpApfZtxZ+YzB6meVg3iPvqiELkJORSosDaomz3H1q025C79Hgjuxce92jrJhwVUczLnhRqk2Bj4
8oRIHV5oWEeB7aThcASKXbai6tnXHzYQPzEr9JwCFUsZGqlxiwtqFO3IHoygqpvYfwFCNZfucw9a
612zOlhxjWpA5ztUyIQI3alhBhAVjsRY/DT9YxKZfVzJBvXFw3I/QRqvpTHC0Pnwt+4/INvrQbHa
VrvM1iquH89/2G91m2cdOg77CduaIAu4nhQh2lLFlPxy2INsJav/vRMdHiak8UyRGe+zYS0ldohq
tUBs+SftP6DANcI62DdoDFbPERc6uVfUdv1hpIWtrL+4r7/gmVcJKgHoug5XHahY+qGWLG6OqdBr
kZ7LjOpG1e3AwMrtNr0n7oClA4pwYD5U7zR7fdMttfF+b45qEGq5MTrnl1tYtvzQ53f/6kXGKE8+
72CSX/7Upjlnjo5Xdad2Gnd0+vRyt68Ice1bgHNOFkYoFtY5FAed0qUawqg0iFkjo3/Ysg8Lhcqz
jeQ/aIqskUxk8FvvSQzuj78fRWDLKKFqgTtKIcj/3WclY6wPnqam2ZZLEW+YPnOQL0Uiz5K5MS8p
vl7NMXYSVA59IwIdDJ0fNIuvSDLiA+3qH6GmkuDCy1nNHdqGx/rUCYoZiFNPCwgWOF1FrSgCULEY
CT5p/Xl3D+1SgLeHnMHxsYYN0Ayoyx0VZs5H1caJTx64ATPZaYLZRqAwWB1rz4Ttvc9ZrJwHBrfb
HaTlzvLvboSuW/qb//ZrsvIPVgsGpJ5yzBAx/oflU/WSb1s9kSdbUuyJXdji/jV29X8TT+RkVRJT
c2ECgXzXOHOmIR/L8AX5XVK2dChwHB/IYeaH1bOQrMgMkDMrk9VRhnRzC3nIOKHfcXj7dCkmS7Eq
VdyVoSvZz0rbNHY0miiuzYgyh1/YNFbYwbH1Xr7bSo2Lvsr3Se/LRyD67MEJu53XRxR2SUsuRa5y
FDpBnoe848yMhj+9efiPOKPTbcAWlGC7dizL1zB5yjftN5H48wL/SCuZcmBA82wfr5C5hZcx51+B
/JyWJfsPWfHHwYVQKZhPN93GMnwPGh/CrcUWLdCn1xu+eitXZt3wm4r7EOpgtl7LMdc+Ff7/etBy
jYIAeGibC+54sgEmRPZeoacReI8vnP3rR7Mr+jimN4zceyux8TiMsT6oTsELYqjBFZOK+fGg431H
GPCZgHvbNQrJ1KYFeLWffpjuNCWHwklhhvPXm34RbRv6DkROy+gtXPzIT8c7gjRh030M17wQcSiN
VMvlfne8b4ZLALTdz4BncDLncyPQkMzvz7pt4lifc1oBsiQxcUpN1o+OfkrPTtCKwSc/JnkELdvQ
q9JPByW2hwQhvBdk/FfPOlX982cEqV/lZG0L17hlSw214Zn0wPL1nOMfsZnFOViFyOhG5qdItAGn
I6XvAFby6VYEOUqGw4tvEqE6BppXTPsD14gCyB5FKDTE8MgPy5L4rYayMDVymi51xkaiqWPbGuOo
TKtyuI7Gw2GTC40R8/0S8KO8CIobtAIQLKB3HLpDfm0BczziguRvVK8Yvz+u93k3RdKkVnV9XRAt
YOUir41vbZlxvxJAVrvymmlHIIer6uoqXr3nAZeuuOnCwh0O1yeRQGZYnPwRlwDnmTcoEOyZDYI9
PYSsp2iSLShteA6p6+BQUum1vtyGCU/59uJ/2PW0eqkzci0gKF6QXI6S2KL/GnGMOfyYW0snrMKb
KEoJtTEjuPl81eTyBoWcp2IF+ueDPZEh1xnOq9QYZIDsciZ88MVNyWEcStyjr2q0wHKb/22n4812
DSVl5+eaoeDbTtbtyUD5HPyZIRZwRpTtxnzK2a90bJ88seykpL0gfd9Vt6GeZEDq53o2/98sEWu1
2WnRc7zujqh9NXsrp8CG5P3zQKCbiXJ3/NHEuRhyTReg2dq0cRuD2iNMHaKeW1tLpl2oHU7+rL/q
4jN9i9+WMsACCiKziB/65f2vA1X9My0g8Eo0n1kJHal2C4vmcH2QQUxABaWTKntBnJaqBR+OIRUL
Ipe9lMc7oqFpdqcDOxDGvi/gmNz7IMswD7NKKKtXrl/+GzRtxn7uNUWKKhbZdkIqfH3twq/Dyx3f
mH9p11EG9hmX7YTn3JtUYEnUtqUWWmzmrPfAA/sR+6wrPvbUuTBu7ObjQ+psti9HR8THJ/9SAoeG
4VOOLNlm5pQlISQBQvRIbIT3decUajWn2TLe/61/NIh7TGS3ZElrJFvg/xUjN014BHRyUHCp7uiJ
i6gbnSROsHAMyB1J0qEJ5y2P/jNR/kldt3X157N+t626XxNw2sJU3JcXfTEpWFqFO5J4w/RklAqT
+KrOKUwSMR7MyUrtMcnThh8NUcYAswODARuE1IZ72gE3RWlnvyb+p9bGSh5cbFkgzO8TAyiGbZA0
aQXRaalVcz/Bmsrpphwen4h+jf2fIjsEb4EvzKmvbcKhlAOjnsVlnaILhRIwH1FmGMENIQeKHjdc
NFCFtM16AvdUtlh6E48ancEmFTA/GfA7fuMEwHKAE+gwblYzzGVcE8CY8hgJLONOrc6jg+ZxrxXX
5zCFCAhzRSqN8QEZhPRxaQv/SagFcimpa8LlOVuQguPTfDUIKo5COSVJKw/XwjnF4iaKDIISyE/n
3OsRRVJfymqo0Jq/Rb2OifmL3iVsDAhVqGSXSxp/i19BlH7F4weShVfyEvVmJ11az3sPJovnwgdQ
3yG8no+TJh6vnpU5+pqM6Wg/4MSkivN3LvvrYIB/RAfcAVjKaL2ofUNAlqLS1r/AFG41RcOlsvvg
NaiBE5nPrzRGDzqsFFVDMyC1GCkHpI9GsBaw7NGmcNXTS+13oKcpHdtH61MpnOmZ7QItklnhLcSp
p6zJq/J8dZO6o5dQ0Ug27P4+9hNWR6h3WBeR4KGtAOrtr/TZXuYYcZwhNL0vEea1fLAHtCD49wRR
kyzpfdZ2spgfTP1OsGHxLPAyMY0o6LJD6SCe8zDqUC9LmjTlnT+uUKRCOW6s35ygcFvqCh2Qd8vM
oxiEcX6sRj8GlMl3E2R29zCg6wUMV213WCPcwHhmIs5QC113u/u/sjQ0Mo/aP2Hsx+PSIkFUWE3b
ShaX/ma65x9VbhRbpVIVslL3GFJgJjAwzR6rKFoztRMSSeWSnhZc3K3Vesg9o5eGF+01rhIvo2Bf
OslZWMUeEa3WK7Q0mItU1A11+71N3/9NOfBAcyHj5psS5/pv6mfgGImGFYjAJq1MqElRklD+ov7b
iwaSC8ndBL4foZtNnB4fhfY44pgmt4vTlXhY3/b66ZOwl65vK+81udDZgNb3T5bVSxwyFjHZvYbZ
fqYTMDsr5+78dWwjeD9oItG4OZDtFtKPjNNApLL36Kzm4QM7fifSPju/zEWoNQlAMUtWNV8pQKKf
mu+IumIKIoV87CkS9SjqyFP78cM+hzy4wtAUrylWiA9C4VHwRV5wc/dLcLu8s14uaIMRSxOtamk5
TFuHq9a8gkTAStY2fO3jyaBPoVHlcAPBzAuzbs/UtNTsHm8v8TlAMzdxL38H5viMgvEBxNfgo/o5
N3B9dqwoSjeJ7RkHGXTFpjCd4BsR/JAVfTHS9QveuPeHy4akR2dwBOXggTsAz5nWLNHTDCtOnZqU
BiEmIACDfMMOallAtTq+Gq63EA32JFJPZo0hXUARBRH1VPBSSy6pLhVmGv75g3wbnSmcZZFBfBZz
VdMuM6PKekvjfyOvrmmnYfsFcEvcrr5dza3IVkKsxIe3h3HA/01LBR6wQydb1T/3iJSG7OykcPUx
TJdoHaYMD1lneAq4cLptPVz26yMMw+Pwoyegu4OX/Bosnl/JwHmlDD21RrrhkKTQsHlY0OZL55wa
qc4R92rm2IEROSGKGic5UaGsIX52fn3HHYh/Hf/PAsh4cwZ9l9SEZm3EtNiEZUnyfn1UccD3QXM1
KxtxVtvKYYeuaqe30NA8K2BvQEI1uCFcAkNO90kSwlDzX401ioD8ZfhqKV6+OprsICWTcW3wUMQs
hiufS52dI9/4hOgNTHAgtne6ewoh3D3j1IlaZ4xukdbuK7MzLPCj7/mZS3c/dFSDMtJOzN3kj6Du
pbr2j/j660cPzoQmCkMZqWjRsTPVdsGdBp5D6uzMGdsxGL9zeMalbeO2jNHJ+EB+RIe/dPqs7LQp
5IDrfzQscppYd1MulniYoxWV+mWO4QfS42HfYN2j1qiLYwbHu0hg1x6bgUK/Ob03xE/nbAwUyr5w
IKG/K/QOqMNsClO9dxCO3WTFqNrgXW/SnpD3x55DaBkbMQRCKvAdgMayWlBzWCHtLSmHjYY03qcN
07wOqpgvUs9tLMXacBEe5X6NMlZoJGQOtqbQR1aMGoegr2y0pSgUzX3UXp3im9TJ0MUrR+0FqbVZ
79y0k1m0eaTXs6Lp5XQxnAX8d0iw0cbWPQYv+/XyUVUt+xv8PVPS+2kJibdmtmCWh7q8PNwrvSVg
I2eXy1eSU1jRGfKHrfTRABE/Re2nQAcNmV9OdmerGNqmAGTjtKY1pKKjiXE3DD4SCyig+EtXMcdF
aHjYIWijuT7BmIKyJqY57OQXQCAs/RaKJeCedsdHnJPf+N3QHlGuOEX9dPG8uQv0cDqFjJkM8rmq
b1998Z2NQTovhvoEPsUWuzCU81/C5cfHoJAl9KUM/8z17SL9IUvaPiRGmSjyceB0iNKtyPBjydXj
XG8TkM7M7buQe3azrOFkrkG0nDvLfmUIHT7Cx4tkkBvVVdasT3BAh1b5HEBNpS5Un2t4oqAdFQsA
FxfrvcTaoTv1NU/FlbmFSS6+Uqefz6LxkXGIsOhq4BRNCIHRdb19S1qV2xEmFRS3rB73aKAnRCrm
AqWEHYbA5waz/Ky4O4hl5oT9WW+s5o101bWyIRtPO2l/xxG4k6P88wUAGbfssX/rPBt9+07MqHxS
rUtlJFAnjMRkT9qDrpP+B1HvoAsvgXUMm0zDAroYoaoXR5MxXhGTJrRZKhVy5bs2GF9Y1VJ3OhHS
mYWb6NsTHPetVF9lGPZVh3XB51cm9Y5H69anYf4W9x0vH9ZmvO/I47j8BPOYGPc1fFd0ncqyqODU
3A9wTThDd0e1lhiLtOQySCxaKUh1wO61fB2+0o2mO3rgSnCCMMAKOdDDNeOFSmMcC/7LbgF4gH5f
qRDSR71Kc1s2u0KtW8ANRhbck3kM2s4b0Qjt1GHBtP+ZeyMQZKVkHErbZpLdmiVFkKbaNQFoZz3r
Bu7o6CENYq5z7MB33hHweIvQHwCacc+Y2ETL692+7Ds3iixWgS4WH4FtaDUEw+MKimo40bKoCqEj
bDeaCtLcP+2EY+OSrqTPZ4Fww0fOLrDeOv/ou4huqJ7bThMsruDol0VmErOZJhtXCxci3+2Qal/d
ZxQlMzbEFdSq/eeWIOUV0ys9VDqN4mvSQ3RD/LrDEMWmVmqqsrpx3c+uGPRNmvv8XXGJc0Oi8w10
rtT5oXK5P6KQvNxWuTowrpn5rOOjugta+hNj6vS0zC1y/yrncjRHMkqkFWYejnhweiWT8lmgkCFp
uKynEuCUZ4SbDwTP4ZiGRE/21Tj1pvhk6emuV083U9NZ4k6hQUsgxXuCdos5x5Le00p6FcVUdYQa
LRgclruFXS6ion7cA7BOSlRKI1eBmwl9N41Yzy+bPJVZF270/+BqF39yGsJTQ7aCyt85DxEB8Xed
OiPtWVtR5iRve2XliAaPglbfh7zZOASoHkUWHCkM3bkFbTvF0Yd8vibVPzV9Q0b/9qzXQ9y5DQMj
QLwMaHzpKk8RJHtPIykOxXi1IYWJ72j59SYxtLGK1IfgCa1K2CPu9xUxtBEDyWRxaqogJK7dC68h
zWNbKXfnASgvT9tF9RymhV16bAgcnny7DMk9xPln5xdf5I+Rkpf58uAJHVQwUxGDkWK2RupbSBTe
G4YF07X8G+8EW+0AACN4KKXDk7usaXhpO7FXHY973BBaJqUIW/v6KzaqH1o3MjBBplL+++/vHMeF
36Ea/XRtYMGTphzm5IEHkA/jnXl07kBixDSF4+47kXTtUCEJE0kUfTVy0qv7CikQVUcCKSJYO4Y2
c1iP4HK+vYRdSX3Dqe+/CczgnbEveuGIHZbj2K/y8TQUlPadVxQxZMg4+VtyRgK/SEAm/m3BurFd
rhwJigiWKQPmtR5FfTFkAXxkS03vlcIIMBxblHSOQaWkvcsEgDasnyv6gj39DUzY1gpb0KmDIGof
RZYfWLUklqcIs6ym22XirQVzuSja+UZZ3O5B+3XJtALEFtiaVjg3MqTF3U8Yvult0ZsjtvkK7YrC
i4Cft8py06BtymD6DwPIM2vkbsJhYEFy36kSqdPPTD8xCZgUYCmwU6NLIDEptAKfI3UZyPHk0vp8
dUMa3l9P8lxKAiiSTLw4tsJxXW1OeyVtWdOUTsacnwoCml3oiDBqGqSyatOlpXG7QDcBiBpa4PAO
xbDBEQdkcta3qVMYVYvZq06YNC+KJkSte06l6KTn2UdPxRU6L2PxHCtBGRFL+usX3ZSDVyOmyjq2
NAKgOF1TxrE/6k6koi+IHXaP0SnOCFvIWqGbWA4Uer5nxqC2PaAxtqc/JoU2PvbroDcgAaQ3qr4V
9hQOQlGElA7SC92IPbzutcqZGSt6O552oU/3dHtAbFZjbN7dCudmdeFlDlXnNkl89cT6daewLtJ4
oEMxdlP5uZGhaYsiDvw8fj6/aKq0jubTjHYicRKUv3ROJI3/+OWR0tf7d0tF/64/4yeo2irCQo32
v2dr59VXO6rKXjR0o3/5HmXSKORuoU7Hw8/6Vhl0CER1VYh24EJfydgxx5gj0mfQXMzpi0SK4+tE
z+u883epaiAk5vfDk+uDWPaejxS5/+Dq4VFy7FdSj7Gnos48v8ySPfWi9df7mYL8j0GZEIVMtRWc
tTTCWjIvpxvrOkj9TaHJ55ZSpeQu0/JFmBgQir5gmQFaQ3RFMQsCq/uCwTx3pQsfmjwZWsTEAINb
lHLZugSpDd6RvdzM0VP9oYNbeB3K/1xb2rI9QyV8n95e8S1gZqMr/i+YjBMOYSihzJUEa+WgEWxG
JEQBIvtvZgYoDFGvaUJJHpPp0ez1sW/4RMM9hxNJt5pMEL7NikagwsWDKn6Bv/uSfS8jeuWtZ0AE
iFOHNDcbUGWEfBhG+XjCTMni0pkBB6TztjcmmWQHrx19W2B1B3DGplxcrpl/S0Zq8F1WHk6b2BdR
wX+3mGnrtVb8rf3ddnqQPh2Ty12yF8hJ778zrG7JpsI5DKjio2ETCKQh7eQPgYphua+VsX5D95up
1pgl9NArIvmqSpj5bFu3j4IfyRi2UjB3qmFSlpUWCbBDVyrGnQtnpqEVebIb7o79qu1PyXsG5Pm2
4WRorT3QycgrtggHJp49deGlEDp7TiX1Me2IOd6U9GY0ku4SmVv7HYczUURWKLxcVYqKoAMy+ZPk
X86WTxx7Dm/7iUD/oF9DAhehX4pkrmespTCG+q3IqtEe4iBSlJSYCyt2ymTY8U8wTYaQRaIho9Q/
qSdcFHyN9AhOnE0zWwMnGTvmcFNxb9sTOs8gn/FxAXy3/feltrcWKN9Gzbck+J/OtQb7eK3JzUUo
H4ksJHwAFgdPVHwvDDszpiaLpaw2/TuoG7iXiHX7ad/s79/kzRIQTBbi1lC77T6RFkueASKMCFC5
4JZxE9OSnYXRgk4bavTtGX9px2cb0t6ZTADp7FopZRnAtB1sTvZe0w/80+31efXyRoh8GkRCTBsO
K8J65zXlH0egxbYzybrdxkjUfvN09f+6+yayj/GA0QFngYfwpPCGYIogZsR4fvS8lGyirFfFYWf/
nIT6rNX5skLMg3Y0vAM0iL/em8as+9azQW7fK2nOT9sZOR1K0MYwnwj2JXJs+Y1YZ1BLa16yEXO3
Hp2I/HF13/+alVLYOGtauLOCsJHlpGYd6nPY7TaluuSrvw6e3oFRVSYCWWfPGACyG8XWoSr+LRVI
k0hNp0n9/CvJWy4tfTiP0GoEUbKODOvcXUuvwHhbjhrhib/VqovJ6ARfVdUpB/21joMtn2IDJZqE
3MoqEW0TKTvoj9W27EFgAJp06Dc2iERoDPbYayUX2v0bPtUahBssb1VSU8JRsnmB3I1iY4b+rosA
cuM2DQeY0L69det7UMTLA6JKX1iAVh6oaJD2xWLhIY7BZCJmpXlxikmDMJUZgRoJ6ZHMisiDqX8G
a1axk6l42YuyhEmR3iz/A9EO+7ztHsSeaRjWCdsJuCxpUwtOBSNsgO5cKc7hENQD+T1PaozMvnoe
Effs1DknDxSmsY9gPdp1CGooRu+gAmCWgPYVyROaEfj0p1k4DexL3ufOy5RThQgG8sSqhI4iVmZi
TH3CaireBj9vWEXseKCBdalrAc8cjPN0Q+TyZWZ99pCo6AlPjTGQa2gq/LJOz0EqjBRxR3LYm3Ta
yAdAAwcDEVBwi+77rAB7cOGzLxaxpR3MHd6zHgR4Y7Q0NHq1B+XOsEEnFHvcdMIiy0Eb96FDs3IJ
IhNN4TMGb6e14p7sEQ14uo4vgxAMZBiuMhFzMgH02VkdauOaUF1PHanT/TruXDyFPpm3bda4qdLr
ba9t4sh/kVy+CkftCI2iTo2AONcPfhluqnFsad/wWdzHHSEPd2JCHS2qTQEktU+cRfCxm7A68z5i
NihjGG0Pvykj7Zyz4aPeOm2E190YbKp/U4hq1FwwLLluwSImI2aVzFKUjKmu4VAAcL4J9oN4vWgb
pcp8sMyFdXogtDnNsX5f2IfkxdImnYQIfFG9kE50OlieAyD7SQd/kYdcxKJGgzVYzQD861U=
`protect end_protected
