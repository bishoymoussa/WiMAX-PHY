-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
BoUsCE82Gb17lneq7HJb1omL/U9hlqlVgYjOX/MsM21ve5fBC4ilv+WA1lQADh5mdF5mnfCiHRzv
ftcEmdlBKAG8596d+wsmGxbH2A4P9mDPo3T4WU44NAQNqNouxaJHL7t7xOzawtBeBh10nQZZeSvl
4EKKD2nT++X/wW/kfrT2OVrFUTho06C2PSS1j5/m9mhIuy4GV/zgOiRqSQmiEe8uf1XQMwEiSxm4
evCMHgWNSYZ3cYOOe0pHo73O3bKRswB5mtV+ILUj0sW8VTHUAoNhJ8hb8ow2BgyF2mN1Hv597aqr
cMag7Y9QooQ7BopQz63PeH8Kr8QaXNg5VtYMJw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 82048)
`protect data_block
wT7lVa22rW9P/TD31YMvAXqqt0dick2bRIBk2z6Uu7cZFipG2SFQXZlMbIBinuq51MtFaCVSmDPx
oJVmDt6AxobWtF+o0UY4wkqtWB314OqkSkILv/ieIVflDBEgubRaqmsyDrhSjtrsGH3G5DSj6+bO
naYVMiXca5QY0+gy7nWrEJlUxk4H7RpzRBKo//AvEqUarrm/PoSb4zHgw4ZAnOtokfRGvSmqBrTl
RlMDA3FibXlmp4AAS2jkXOUDbLe7RpN2JXNacVsE7aE1hiBiDGxDSBqEXeVqjKoVKjzsLnO4YBAO
jiv4SyOOFBvpMhtNLoXT9ALv6WhHeSDnR8446agZSTED/ECPUrazMht4evF5Q6VfSKNZLaSeXHII
UrIY0Grp9uMRhIE3KNgMQLGksSFq9ys4cmTY+/qWz5jwY4DYtH424zDAiRLaEISAaEYwlcZp1sLl
4nJFpdr+X4NFSbx5CSaMu926yvlvUXeVU7k3g69U6tiPf6WNh+i/RY11z23f72IMqpHxKVfXbA1L
2NeiSbykqJM8IPv52Gt04hLJU0s30KNv41qEwS/1XGdLhdXkr19d0mAIFs4mnzjaxCNSpNy11Blv
yKVFKFzg+HKUC+EmISo7/m3yKlaGG7keqyG+RjMmW7wGuAUghODT4Q7mQGOQucb6cvP31recieow
hIB1Hy89JfTv+YWczTnKtIyUwwjuVsyq+gg1yS1A6YkBoKo6XbyhPR7vKqo2rBGb/yRLGP7dpyTo
I3IXbOXJxMNaBa2xxJXbmFUtHGVnWG0jC4Rxv/XNP4Kko6V/W78TX2Oi2+gjPLMGVD+2a/e6D1gs
YRrn5yH0md1uv9GoFM73tVXe9oapcPnj+tFyI4H4A5J9j+CIRo4syRTcvnVm/A2aY3s3D7vrdhxN
xx+grB34cVGCEU6LIJ5zkuzGt2dNBfbCjWEqf1aEpGsncr0pcLo2z7sTd4cn7GpJvUmHR93PHQfZ
azF4eh6974hJzp8td1VKyENtgIM3HUVA3rIZSZJ7N0Q7VmP04D52VYL1GAzE1+4eDu7xEtd+Xejw
g78v3inD2OqvTctP6TSMCsUGsr26gfICGmNeXhLmYCstjWAK76jBnW5d9rDZJTrjMiQWAZgXTpzS
k/mMfnXAAhxHG3mTfTPjfEr/UeZdhbzfV1cOTvi2DBpXp+8/GPyB8TUv69eYSmmipZnaDAJ29ZpY
Gtr9YW/ltu3Txm0QqTGdB/5ynqx1UMoRhjHz3g90SksY0eracGXvyLIVgk4Q2PBhPS8bAWG/vI5G
Fezw/WqpD/qHlIHlY8Q8Dn4blOOPyXAwUDJRBH1FQpntRcUFRsEh3oMfXp/mMRMw1st5bALVpM+k
sCXNADp9/RTpU0sNFjD4Q3CVnf8jp14VrF/WFpA251hqGoxg5010wu1O21qcFqnkiHCGTd0A+gWW
iTar6vGjUJz5wL5xOyj7Yc9hMfXAEhsRWakkv2lO6ORgHyNDZuGu6lgvgpAb4PxOFrUV//sbNNJd
OS34hvnTku0gWlQKmyujZB14BNkAcNqASwHgqfDJocSVezc0YtM+olfg/Kr0vpbQcp/NHYoZPCsh
mXzpuaOPYta3rwgO6uIalA200hl10a4/RqB4CHkUEz6aVNo20AtlAHYJwflCZZIT7tGO7Rio4i0q
PYJrGTxAtcu7JMjlCf4lyvl1k04y+EvCzYqy2mPsyHeWV+QgEyhnKEjBy0+ARBsuqzzM9dGxXGzm
prrgbPbVMxHyZx/i49xdcUcFK3JtGuy8RStXiM9G4SikNeH5cAOUpRkr8Zr3l6QSqGsd7iFBKI6/
gUok7blnKQksXWIw+AqBcje81uxsgpdIAZKJcSjk1WhRWHhifuxVBinJi9T4+zYIAoc3J83C94Cr
8hlrpqRyKYTbfWHwlPtn3TDzp9YFBHf38LWij+p/TP3nKrShIM0r5HyLI3O5tl2LVZIlIJKHJXtX
7GXhi53BTJMKvvyBghPzG3Gj/GGOoM0SWqLDLpucdR0OhfCqVrN/w1viHpGEPjsNCFYmgY678jVM
c7TwrRQ7VsRIrQ4e0AeXgYn1AIzguMbQ6qGi2hFbpKoNnwwf3XEHBNeCuobQTjYEsaSQ9PkYwAPX
e6U+yBUhIxTFisD28/gEcEpU2UW78sd+/rirSf5pUadV9xDMes8NIL9nPwFR0cqqMqPgnhHCG/vF
YUgtNLejb+eaw+daj9InZCHxiKzpUeCq0PJcV5dUVWpJHxe3deAJKP+DP9SnFA44A87CETeEOt/T
tbnmyIzNb+08cdBCN2QLKZh9Yag0zyUID6sjanzDCW0/gGSBoL8Sm+9vM6bdQ6+WGovhZO4crV+e
im7JYrYV0BJa9aX+Bt02fnbGzX2rroFgEJw387z1nZkm8S+VvK+Vf6U8EcCHlOiEM37JpbROGbFR
j7z147IxVsGAYuPa0m4vtBW+dDzfxGYEUJBF7qtluTBkPSEmp7VOuNK2BORpK2Wa5xtI3FFR1RmI
uprmJXb815GqYCqcyVQfDW4G737PNLOqUbDzdfRK0aWgiJDVVo1Lz3EYk04i4zzFVgFJKBVn2cRa
61aP7WaEiLbsRkaGaCHSpA9WlFsy/zzbWg2UzzUT4MGmmx67x6bPpbnYv5e5ebVug72upppumSes
CbA6QKconRe8gvNSX4YAPj/kOXQz/R9gaoD+ctly4NtT8H3zN8tgXCHSZrAwA8zUAYWmiO48+pgO
tl6T7keQcgW+zHGlgAP+Ux95XFO4rrP+hJ9e2VAkaHNjmSTCY5xabpcloyz5wGGymbtXzYz0dkWU
VhDEpdHJ+byyxmaFjNrtL6Iuc3vUhrFLjHCahRFfz169zoHSod7OeGawaqqD4om7ch4dZECzJE1+
HCtvFs15vQpsCwP6AluelnM9LgdzTe7jaLhlcN73s6PVHXLHjF6j9voVGOI0p/Z3F2WhbtpWLVCh
s6cqm5Pv9hYvR75d7ScKMjJmz1tQFZQI4F4mUHtoZyLA1ylCbE33Fd4ee6imG0mQTlExpzdv0sr+
sBUURv6VMzFM7C4eeGhdMYOOdioNquaX1uV6YvxzQaz3wSuQiO1FuadhMrGRgc3Fi9sntdZt5kDp
GN1Z4CJ6KVgKeCyW7FL9RG/194lne4bqo4HkI+P6VFWgRvmWUOBYy8LdBNBoLriNoGTP0yN5h1Ki
iF3zxVPjfPrVTs9uETPSp9Y+IpQMBC+9rKzrdFLkfXs2pbJwwnPIBlGfohfudGBH+4ayEAtdUtn4
nb9tGlT2SQildT7P+4qmy/5sqjsKAjCSW12DGgx6EoKi0aGMofcBOa97FHAg4b5hhzB//VwTtLpr
IZ1+LUh0etIXk3tOtvaVYkV64ub5DUVWXW4yRdjAJrShZTnyPF3+Gvr/OCd94TZUfWLR2KsKNF/j
+06/V9ui2YcC+T0E/3xeHnmA6jJqgEB6Ti03WPNF9aMSLziM/LqnnMDk0O69Cw3kXO5AFYi1AVxj
AD1NIAfbxVQsk6lwzxEIQDYSM+hPPZkmpHQWkA2HKeGI64+djcBB40V6ozDVexu1Xxizx4+8Jdtg
YVaE5VVH6moj/tB2kPqq8OY6CVxNLnuhDroOhSC9c+1Y6Q/bbk9mO5UzOcyndK7sLg3LfpcieUSx
1VACGJOP+4d5861sTve42JlCgr/leRFuRD+acZnyeZriVA7XgVjvhCkbD332eOi+mViTg2nQFMIw
ISdBZi1Ht3cYtTyMzAHJKpsk+8wf0LLbeFHAs5899vg1W4lHb1atcL7Y80CgGIYL0ZfQbOZlVnJ/
dCbJ/Dvu4FHWq6WKxHFt56EX1XBhEZlNIqFz0BNPDtiOqusKmQjGdzWdRt7pdYcQZWctkrWASt6H
bhXpJv/uAW4sovShn65LLqRjd01AoM9ZjPRABDWbj49CYE7JSFfTeZS4ym4GtHGh/4Eg25g1GAoJ
IvPO+araRwCTWVhjTwqb9DrFHt8fpzy1ZPob5XOkOTGvVw8sREkdtPHpsYHN2BBWin1OfAPhcZ64
zKsjyiVl0hek4oAl92SEOAUJEVJbS5IVbu626hf8+WMY/xLGBo4ZnRGW/MdqyNb11g3Z5QBKhEB/
yYZT1TEuihvk4esptxiJLTSrU7mEwMGiSdbjGt/rWXdftdo12W5kaslNmF+wn5RJYMg0rLAXEBCT
r61ROjXgTbrggEGEtJw8bTWVxt9r8fVHA9DFF2O1Mtwa8uFeu3Xi8NBJ5291I37w2X0p5ps/TcIf
O2nI3Aeq6OICvwUzIrGTYNxOe3FwEXLZMFUf8YrCOzMieRaBqIJJWYBj3RjiQAavtygbuG0+CVAT
beBxqNQ3PPhHbFoWAMbpykyiUQtiTCfy4Q6gO0O8DcYZ8VlZ8iijhqHpDgWJVny7JuGe8ZGwKzwq
SqvJMc+2E8yX6PZq5AbweoiuNjET9hAURGuoGq5gwU1XCZCdJgkqT9g2ItfVLzcF0rs57j55R12s
Qe2ahEGDoeYFnsczcrgn4cCOUBYumxbqVMg4C09g9QSu7u6+7AJFAYPFZoUfIOjpPwB8MtmsnH3U
p/OZyNqmT/a2jhzEPkZ2tyj/XIDOmk2UCVGhZGohdQzJp1wMfds9jtxOJkT75UniiYDlQFgYJfEg
1dyrHqte+6M74aK64XcVC9Lg5YrTaM5OlO8y0bZxAY1Jd4+ApwNO7p2i8HMJU0dL7HGhjFDBi9+k
BjFlfS1CTKEnJffySIIhGoTIe9KRv8GNo2LD9kK4PJVbygLZ6JF2U0W1k1cpRFyZKPB+WjhyqwKE
0mYDVvSyZBsQPJp1qHs47vAh5O7mQiIfaNWAPSI81WHr/RYG/Bccz18h5+eiJriez19tE5ei7XKJ
KW9Q4+Dq2WsvZ2teUv/66Np4t2art5Q5S20o36bK+o3o5/yF3UsUftTUBggdVLoW5SMlJVRmPTWG
nkwSuzq9T3edGhHBSo9ZyJMGwnkRRZMI6uSRpDHoHlTgaQlt/DuuwxuG2vU3Y/Oli6rZ6tK5UsVU
BepPjDJ7aRin9QMADQVmly/1+7Vmkngv5hv60su9O5z/uABDqWOiIEWDt+LDsTlIWkPB4T/og7BS
M0hmqAeXiekX/fZVQvZmdkTznqVIw1kCojZ7zZQ3NETzRR0uBxmLWluam05uZYu5dLMU0Q/pCl0p
7Zjz8J1m8RxCL6kHIKyOohBsNSy1GR+LMCP7DEb+2bA6xDEWNkElcxA7GvhZT/bjkLL8Z3CqMOKI
32e6Yrx1F5kX5JV1UwmcqKPvXQCtDRgQsnWhnHZ3OdGSLBXINnqljn4fvq5sV8TXuCdKIpfJpG9w
AJQkrqtcBh2BJaqW48WXZ2a8uWCvy3cF3RDE7Waxw5njSbojeldwAPzPXTkJb1PzXqhrf2yaWouk
idReOIg6G+ac7Yz4C6yT7XDNGIsm6zfaWqov11R+fA+QvaqZUuLk9jHPx6OT2gvD7K2LNixQjjTp
wPo0pOZUrfc5aTjLYF1vYmVnjJ9OJnd4krLpAQ80I339AusmRp+YerZ2rh7pWIO7M95sPlGoQTmV
04xCyCXdY17CmZ0ik6RyIFu5w4E45ZG2ya0z1rvT9xsWW4c0/yUdFSYDVYmwuMvODwwh6hDPmMi7
b/a7kKnmXjnYO4l8jEXR2Jumi8/Vrtla41AWeLOrXUtrapoxydeeaNxbCv4qBxrEmRGEtVwhCVNH
v3ZLuszEjEX8v+SKJLIkL3NdXQ1Eke+YiN5cBZWggUVKvzIVUsE7YwzrRTTdt9r6aLQbWDtuqXRi
ZKo391Ks3wmywla9e7KcJvstJyQwQV/QS872iBbSZ49h2cxnzwgd5umBW91PBxTw1TZTmDK39mOF
AUyTvLwCriGVQYvuLE4Ydqdl6OFAjw6gePyxJ4W4O5TKSBWt12yfGFvSBiwQ21uTJtsnLmJuQVk6
TuTSfoL/xRu589drkiuJoHssOESzGdwwPt36rgHse5/y18Tpp053XMTSwA78gRBdUvJVfEF8HcDx
lAjMZMnTrlHA7sBcDe8xZ1WUVp81dR4hgg3kybyC8ATm4zGzxvwGZ/lnYJeoEDK6OfUcH1ze+Dlt
gieRJWZk8jvZIFOsstnh8Bv52NjjFFaWI/kYgiIL8ncskeYLAwdyjhxUQWscLiE2SCxM2S0au9b9
8mRBZZyGOiSoacktPkuGMPEpXZDZwcXEy4q5q1sSAeI/FORl03ZK/E8s1r8VI/LBzy9FChQgrtl7
GNAnD6gdXNsLAonflYKxDaPSH7mcNdlhHiQXvAYf+RVU5gU5fVvdm0txslEOHxSWcBKk0hgpcKPh
i7Vv/n4l/TIdK9K1+FTInw/coHgBefCZJKZDr6esbA/vmoaKKdlCyOmkNqcA0P+Rm3rB3w8bQRM9
FHZbGFhUgAVUxTFzVkK1BVnAJ7uc61SX1cjmPZZq3+5TNavdguntEPL7srbQXXFjDhP/pSpco17Q
TmalX9rcpSQ5zDLH9/KmrSd5k8r/AZi5Qwci9we6vZC/xM4ZWBZXpPLp6JK/Jp6YR1BQxK5KZc0X
mRk5FfppJZR8mZ5jABanVuG6zAfnlNcazDGHHPJwAm9f8cF5m6kD//Zg92sLCKxrO+FsTFJ9TrJs
NY2oHaY7tsWvcYIn9SqnyaMqKvu/ZfFRrndo7suHhxzAmRf7KGhvDp7t33oVlG/uXiJUESe6+q3A
TFSD/Bo7Yix5Itw4JjCjYrWNHixHFX1Pdfqpo+cAFP19OlIwgDa0IrojPedj9Z7KBRO04FiwwSM2
6/7VZ1ku9mEeg8i+LBItUJjCKcVraiXeMGV/LGUibFiSyGIeOEhdN1RZCP53QCkMP9P4pWx6g8Ur
CPxKkxwi83Pg0+gctWKZRmgfq16SpxvyZstTnVN9HEvSXUoDKHRbu4rP5MvUBUqIXk2786kxVW6P
ThVPRbvM2VTY2vZNOpgdfbVfVn29dSU+AYENHSOzgH7gWf0zOIH0JwNLODiSyKI/siRbAiePrKLI
s5mTfDU9U2zmhtdmbtUrHg+ZmGYavs+r921M38lsE/M01mPCHwT6THRZffHnqwRMSVgf4jh3BpZF
mbHcbvcSrrjDPTP3603n6KcKcBVhqSru4csHbxUqW9d98BZZifM+y4+H1GU742DetWtYxuZqCkhJ
kGMDoiI+ipyjMZkGc/d6rPQrWEv/Hak2kFrQmXKfC1mOQNFJhiHZVgtVrVvMEs4IFlKqApbf3kd7
InFNeLBlBRnDSaSxA2XPCGX9EbylTvlKRKbfVAZQptFeb41ArO8DKriGyzM+14Mt2zAWNf6McwsY
XPKovF5HkTYigfS5vzaCNjHnPhIe+WtMPnCX0KHkVi1LgKk00H3PegkvqWrWuJE7Ng57DAmaAXAm
39tOdY1lBCOYV5zApw5VD0ETEr8UduLVWSj8bibWO7KfW/XaPKeXEYet1RURXuKpc2UVvOSC962y
ODF+rrQecPD45lTJ8amrIGhKAx8P4us/zrggPt35krGaCQIoQ8eYrwrbXPWkcmPD/W0YK7XWYzA6
6NcvUfGOF37uoN18/3YxshfAyPo5ygDaXhAvJz130GhzQ3kbD5447WV2K9txk0A/WGiu4g8xXPU0
vrQcn7DkN+VAUNSC9elQmnv2Di7O7UqrGcnn1z4D/bVLhfbaqm/icl52ComRr4v8z2pWgyN9gioN
kbOYy49wXGd78EuaAU0EgrfOL+H9X0smjwxFWqqvn2P3r04bc7tENS30gVKxMOH9HcYMbftsA+I6
eyINVLgEygd2jnNZbSe3ecSOwLF8gL2DbY1BTFUK86pVrmnPFA4jQXFzGI0uhbJdnzJsguWWG2KB
gdsdQfmeRINcykVkUAOxq3OWCHCIn3fnrwo3/3JPjn3jKPNv3NoxtcKRIpBxAxTKIs+wCSA7HGkF
iAdFJvmGTqKGJbacfewOOP6e1M+P403vJGIkpyV2Z47wg3frFhkG1Yv/hi6hcLoJ1KwiTEZUnHbX
poxwRUqTC1ivdO0eHVV1DI1ZZx4t++r/K6VJcSMoj8IwBIWTtbBroVvj/4Hk9bgm6moF1YcRHieg
Dd/UR173oBN8euOUPhn9VLiTTwbkk8gV7UfftpYzfMekb5WFJTq1W44T5qnCSOBVmJoFPjD21xCC
nSvYu8qoSJF3WfPfQRIe2LvqsPIOB9ZHNAiu3PV9tbCgaz7v/SWGCtdcCNq1VBv9kajyppIL1y8M
2d0xpGI0c9tKXH9yRjClFiynSeHmJ3lBPpUx/YtnSzh9+G8nRBntIRmssBx/hwPMmSxkNNUYS7hj
0l6p/Fm9NT0ai0sMYHJu+1yzpwl6oMocVusn4cyyTD0EZjGpE5+jpWPH5Ljbl7feDo3t+MWRGSHg
+3ZzmyXysBo+wpB68bkK7AfzaaDUhhQtDnuQ1BCZm+Vw0rhrG0bstQEy66TMwKOth+CMp3Ii5WQx
uWLQutpkhaMG93ET4loHB56EZBXOQ0V+HK6RMMSXna+egIXX/9zhfbYVaO6z2dAyyqUS2WDZiwUz
UICBMSGD22WwgISe98rwH7Gvs5505n/Jz/K5iRQg25rWH9qs+DZAhZj8PFca4xtKzjgNJqXsdPXQ
53ZRK0IynwDyXCH06J8M1et3sZ9danV6bAd3EWdQRw/59Hq3ZFV3t0ZpDnbH3WWEN1+UycaS8L/B
1m0WAACUN3sXTTJKYVVLMDMhsv8RF/gt1RzCViWx/5pNNeTkkakpUJr8w3YwnlCiJ9z4hf6rkGSP
zqGFsf/PSoaYLydwG76MiVaE7orpoNSmozPMdck3yP+R/8al8AgA70BAboES66IRksYOyP9kLSOT
aoXTHQUDAkQZi1g5KfIWQIDxm6kf/B570aAGiwUHV9gldJu7FUQ8nn+kzV14KTPFrgru60u/AKec
I4StvufvsCFkw7OT3JYZ9NADDVwGul2rF4cdm9OZ4eYr7TC4RUdQv8ZYEznZFP3SNYlPu8KKPiUd
1xFtmvMT1T12q2VNOP0+sQfPX+IZUipYVC0BhrQS8spsfmYevyorSlmg8mYGLVg4aMysF28bjJkH
hl6+RyG4guzTQtqJH5TmTIYv9NRsnoNXog4fsUf9IOZd17NyMik1Rh/CefeY+FEHkkSigGV+yCPo
brQh1A3et/S+270rOirbYHaNmDmbxZMlDl43xhWcrv1nDMkszLtTP3AslXMLFAf9M5oz35FdznlS
2I/uaYmWAA0fb2TUyI5r0+x0cgw57eo7hQBlEPNDBAhoqrGD8LdVug88p4bQRm8mYNeCpfG57Epd
tSm5Xs4PdzymUUg9WucV0qpby+NkenbHLLXeGTvJGI67pOvDEi+xfxJTPiNVbnaijHBZk7MVDwod
7nFQVJJUxXoIxMV5VDR7ilq5s/gOlOelIllWPC8vf+gNX7MHVIEGTQjPale88Sd+/k/c/c89O43t
/nSGY2gvNpfGiSpkHvHHDRKmEoPGH5aCUOudvGHxRH6uphsaJiVhxeVi1T58qtHs9O/pMqPv5qMx
GiZGuwqaw/TK6WPaMvmMQbETD11fNZoWZh5prVRktUT42VQ100MmS/Yq0MZ8LGihza5ZhSTFXTU7
FOgX37Mhcoromd2LhEA9OZjetg9f+qUe3bvYd9/Gu4dQEMBClwt9l/+GiWEh0msFHIq3ebTGKYg2
EGZeILrsWoepk4fZvRVDeOIGwKECHT5cj9TL4fF/jD48m3X9JspNPu7J5NS2MVQrXEInOqV3EYR5
DwgMhzbJEb2TfNpF372jBMAsnOfc3lvAKnTKyNuyctVeS61OmU9TtoPUDO4alZna3Fy+qEbGNnnI
eqjQkwdi7VJ+Gyw8c9T0U34x98OPd+YRn+pf96pLdMc6/lIGaKSI7AJE2gfZ1WV+M6+ODkWQZ+GD
Jf/B1OdZJsr0iD7+NpmHHZZp7KWlpFcloQlEr2AvT3PEiz8wSHVxMGH3q7eiOT5XDRrXEyb+cFjp
VT3K5CE4jrQYh352qGWOqCyK0evbWMyfCv0sfI1bohO1vCfQmLJ6eEnzLO+yvDNlNcev4n5bLnfg
povr3S3QV8By6FtCeP9kcOXwHkRigKcnw6zx+92wf8SBSC+4BuP6MezNPsYh/c2nKpE4eK+AtIsS
cfJ83YT6SUXEhVoWwAzlq8q3iD8coojjwjeZLE/6atDS9zRgmDCm42e5RTkstoX6wx1v+5P0BnMw
f5ASuOzmFeLKqRaOQoHJwNrso30hVxB2b9OU/DPZfq6TVkUEzd2/x9mLNLoKZ0I2xB0J+5AnZfxA
s2UjYOfq9K+mGFxYy92mKI8/JuqKaSXk2Xq/LL5R4QpP/w3Di9yEQOfozfmhN42jXr+/9lO2gUHb
qK6bAgObCBSDE9gp3vQQ/uVB7rQcUWKMsFMbXwYngY+ybKJjLdjg9NWDexSmZuWiBXFA9K/OZ9Q2
A7OALobQai1Eg7c3KVFGnyXVpXOqVX7b0NflaDGoQdbu9a7P/M+7igx1sYFxN6VNKjsI81hsKf6N
2ijNuZh687Ekh0m9Co1WbI8f0n3jjWvG1RcMXjfyo78Zlt6tJZNEvxkqZuf4tg4knPOOZuNkVZwi
EdqoxUUp6gO5buqRiSZQwv6T3Q3ua87mQ/iYx3cI35Cv25h/KUEVtz/g9FxBvYHWCRQMjoqHushe
/f+UgCp0oTNVpnAkiMhFXOVS4kkiWnH/ewXcpsFREVWPk1ZTG4/NEJ20uLd5wA+Z1b3nmb/FRQgx
YyD/AKzGjCPIlay/lltne8VSwP5pF/hWW4WJb/EGPZ4QYypoIE3K92ly+RPIXJhxFXSWierDxhQf
maBKM2KxAjW7Bi6Om6qIcxpLrHOpgTZGdvzNDxbgkHk2GAnVk7sJAGX69Nf95dyqP+Dd7NF8gJgo
ZFrm6OFJLXlLMsgdE5LQXG4gDGlfsHmMJ1RMRnUBpps+rikK6z6ucNx9U12HuGgBKhFoha0rZFw9
WI5P0R7cKi0nYOgHnYPBPoDULZDvqQP1fenotmQSiE0I5y2Qkk75YVxcE/2WCgSDN54RL9ZsbX7G
mNRM+kDmu0RBDeBHyFpB/gPUYbsxB+n6J6cUBEUiVDesycLNOypAtfJu+tkqbTyUQFBIK0GRJ7Ct
wEHrw+HUXvub8+ww8+iZtK18jGwgjXeEL2Kv+qIPY+Zg0XyojyffGjHyxmon/xrQ86YpebvwB8Er
LaPh+fwMyU48ng3Dd+a7arkLV+xB0nuZe8wosm6KcZZ09/hmfTbLHcN+CD4mASRABCMkA3Tw6eP+
TINyNhlQ/qlqV6VXDqZkZHjOYByAd8igkdvMWn7+2bvH7fKmIKj/+VfSECcSEEQuiYQy42p4c2uv
jpDMkvSBihnsaw2436Uqq6MfHkdVN0UX6oVtl5JGevYIqztYqi0S8zS/UhfEqF1f9na/v3/adD2p
gMCsshQ3/2s7ZC0X4Qh/tJXAuZkCS6vlT62M0+EAQ+bo50eeqEXPaFNJg6S+sqWYBsqzSIacRgXt
8yTHG1AJLDulCNGDgo/UZ2vkxg45lelLdCg+6OlpWVxEjWkYWiHKy/zqQ95GdEqRdzIFmvNTX0fc
Kij/DeIwYkIWgVFjkRSuN4tICud23dvvtJBYt5Kfhr4PMF9FbxvhGWvYfiAw1ra71ILobXlbPcBX
v7M/JrZ6z5QCYgwht4AiaGh9CzjcG9UUhpnLvJALcSrKMAk1/l+XqsC0ijSIEQV+KW1/RUq5uRuN
DdGs/tdA6arEKMRQf+Jd/5TKo8BH4mllFjSjs150KJABXxoMEYvevUa43nTKBet+SPCNlmx4JdKK
vvIYj+dP5rUPn2IsiYhfd9OMygXrZRvz1C8EtAFJtOoqtxsIi+XHU8SHwu08LdVnqW9qRyCiudXV
nsiUWV9rvbhOT1Fxq5oFGiBWvgOSxG8IHTxLdwu5tjpfY1eWnpfNqeteU0w9XUNr3CftmUKdbV7h
4oQSa3v31+ak919vcPa7NYEuiWkTYJILvkbZXF9KK6VTPaFKPHtxprRoGQmYuN3TE460FZFEPiYf
50KdTH1jH5a+zuBAU4a1s9MCkLFj4dbB+sr/e+HTo3fe9A6DgLs6SvPmY7WrRX84QQWQGAfDpLi9
9En1X3nEEnmqv18UBjyyVr9HM1r78Qm2Yu8EDtiMkHmUXel4IJsmRPARYRxfgDuZNRvOQmyAaVrg
H6GVb2NxzIO6MyglMT0eLUWTmOSsEOR2lEfnXuIBfD3Atq9/feN5oPu2ZtWS1BdsG0ACO7MYgYNF
lDKcKWYARq9Y2OYrKs6d2QWeWSPnVl91uhRLszovjilic+/p8v4pDLeZo4CeGfdmfd2zMtXFVp+N
aK2ocMk5FTtvmHTRTNOCtPsvtwCpzbhKtYYylbSAAbXcMMu4xmXzJBMEIfc6Q+xdf4Ao3wbJ/0wU
qDBMe9u/RDXMKqE1YZJ4lb16T/g5F2myiOkjjvvPyHV7VB/WbCgAgCfb7F8NRc+MxX4zGBq8qX8x
BTJP4gx/GGsp4Uxr3g1ylISA5XbrNAmntc9lVfusRaG8dDrkyxhfHSRrgakb6y7AVakGdcmisLES
lK2EZ2k8Ae39/Wacrk4FTtG6oR4+HvEV38fQlQRZ/SDvIlw62AnB8VlrTh0nt+b+K6L54xlF9dRL
NRNK6ATAeHqZjX9EZGlB7mcW/L852uwk4oNSU/uZ+STfvcS/3P4dETJ2AhSdli7CcavtVtu42vww
5pwd9uHNloVrFg90wMYP+AAJk3zv3p3H2UpvVnlu9/FdXZzi/Umlkih7U7ma991VtKJ+vmO7833y
qTTdQtCftxwZXVXcRCKQFZy6J1SEKdR8MKut89s4CA7gh6s/y6Yqed6FYAojIW7lzscbXlPmL4UD
uxyNbfvZ4Ybk/Ht9OJpHvBpzjGh2OjB1Ym2hpf0DMHiZZ9dzO8F7ioY1RtgZPB9YtfmkVPxIHVbh
jkCfEQFn0d1u2EADn/hdn7qg9Rege5d4qEfMD4iy8arxBeIrXbMr2OTpYvPty7hKUICnfVq/Krex
RHcITy3qjVI69GzuI8ZEP9Jioc4Y25/IQZ7TsmcxYjPDO4WQg3q1Q4LVMiwxV0IzX63bg82a4+nU
EW5q+vA3qucIQJvlojPfLLZx9f0EQdg3ly4s6bwUIZmGrPxMgFirUIb3m4kJ/YKVYgcXq5npFa7L
byBG1TPpfsoj2nm8VDV7tlCUAyIV9RErx8nNVcQmMBwvq4zjIFkfpACAX6BpfR1uUpsB+1DL0vCF
69+JMl2kfeQTEfhbm9KbHuZM771QncIJhTUZlvp9CO01HcNWeuSloTcSD/qJBt593aQezGpKnlZh
iD6+9mPkeAU3EqJ0VvZoxg6aAkUh+AwjnTvhInlScm88iFUxhgYVbdQrRKmmp1QZU2hDfvzLJMYL
6fpBwv0SgWt50uIKq4OrWEZYY1ZIeuWA0kv8hfr6g/wQxoSJ9AkFNUdMN6c3tisEN5zi5LH8UyMR
sJOfTg3aXbCjuC3sW8aeF7PqG11BgkFxpHYia2Inr14LSOuif/2kBlk8XZPs20oOKtzA0RJs20wj
fvAw7ZneTkajE714xDYUyBtKOWci8zjLCvIWkyeVI/iUX/2CSjZSdI/C5ZpvH9av36iImltn6+w6
Y8Yan0a0s19GGc8JD3+EHtEc/gn6Qhv7sHHIdloqH5kK99GEo1GynWLWGSqjVGGVS2kmPJ2TTe0g
AgoyqnS8hZjooJn5fdcBFqEX1+weqWlW6QGJY1j3bo2M2jbuQhfeB2XPPBHlQa+CX0vs3+VfIeS5
ttMdxXoMokQLTC59phuyZnT0/uvRln5Q5yvw6tpeG7s99Q4FRQaN7quzhP3JAKcWBP91m0nYs8Xb
6hBd8/gvU/QIcs5Uu1+25djaMzPDShEbL8LGgIZCK9O6MFvFsv1i5LGEszG5m0qkek3i6sh1UfYo
lZgth4LmmMqheJsxf5SWJL1eyd3VNlM37Gsx7rq0l1acNw+2caILTyD8OjeSdHU8HPCcgr5MqVXB
rJIC8+56+4WGqGT4CIWDSLX25CfLcDbllOTYNL05brqXhXRTb80UMX2WPwILHa+0tPIOLCxFeVEV
plkm9nP6GO4l7SbZjlp8MfLVecRnkqOkflKJ87jKWRvObPxWYX9Y45fll9PIKfmSATJvrLpRYCrn
QHIGYGZNdRcPOb8Gb5IEbVu2caYexYSl1XSzDCCNJqTJhbGWO2oTRaKYBk2RcBvtUGW3BdmiCYjC
Kr1pm2YyWBkkZvAvlprIrSZI8IY9M9Kn4B2uvRQgzdamwZ8Taefl71G80yet3wDUQdHg0VwIB0EP
a5sXueBirwN9ucsei+QP/CQuiFjUFr+C2Bhp0AyX1cXr2E8HmNoET/L5t/byHBa50hugxko4dqY5
xNbck+3UnixuY7hBkr6RtFyiqmVuO6yK16A+dgNnvwhfBdo9sxnVzM71FF1mzmlYlSsVkxyzkSji
SSDIcmUWEpnMLp82N3uV3aunSsL3o4KyeRgA4u9fgO380+cQ1RaN1r1/JDJGU8/CB8dJOlF0Coev
YXSbV7D3focSqY1zzDbKQ+qceG8a0jj2VZlbHXUUKlYQa7ALfW/tjeD9gLV0lb22vqPkw8xQvOA8
17s4oJIyg9+pS6Rlac8+vE4LfTFtnhC/4lA5K2igTwmubOETTfcYMEdlgpKiL9cthFt80k+Zba8i
aDcZD8cxshGsKV5kzg6Y9iUORvNSTkXBHSKTEqgbYi4fXIzEfD9oxW43cQ3lXF5JEi3NZUTLP6I/
U1IYZvOPigGJgYHhme/0yG83xlfJWRACv+eECAaao0we4eDiTRDIQYInHFx6c6B/JTIyxUUyEsUU
+giNZO9tt4stpM1Od9aZLFI+x2yaIFuRpssBmG5RASK3YC6rP2Yqv70S/LgccZG7J5Pf9ikmttIW
DJlSKMtjAL91AhhS58kKhuOkbIfn/YizCZZiPijRgmB6kkl2qeS+KwSFjtNcAo5wHSMJBJj38TDD
yQqDNOiz3SeA130nqDKDPQPwnkekGN1MxrNCBk3/cgw4x3+5W8QYyqfjX2XpjK2eS/pKBr5deD9l
ldbvAHRAELhY2drNc8/Vi3Yv//vyaUGe1K2kyu/pTfRxlrP8ApShCOPKhwGfXn9E11XYOZU2Zr71
2M3WYRFR0aopbOZTThV5RhHEa8Ut4BE0CuyLouUs6qr4J4SVuss5oGfJ+FnHg2e4ZRny+bFb75Aq
553bzifpr73EuYl/sBgliYD2IfjucFMlemAoCPte/2vmRQjMD3GR0dB9L4Rlj4tWFLmhyT0furVv
KwBrtJMhqdHGPECHbksUvm6VtTRJoCnFqe+4AsXmLnhnqsQFvhpeBgUJR9KCrPoVlElUarnEfPZf
nOK+m+EozVwAot93LDCuoUzHEVOy+/bRPgSAbL7U+J1t8J1n+vJTQWq2qQILFsJvaBooRnWc7pMT
C0fN4VG2ewh1Xyqi7njnkDTXiP1VWL5bkCwSphq24CBOQs/c6gQTogaY08U2DPqa9nszvpmwvroJ
8ojO4uvoATcLEIIL6rGdZKubaCiVL3gZnjGnraW+/pI75MPGxYQZo7o9nAgcTbNFZcluAU6lvVGn
meO4ze3W6YO594/L2zJquYsKvkLylj7NcIw/Km2tn0nHDfaon0CMCr6JuBeIgcAeWYjxo6XtsGyB
JhanVOBttLZOlnsxAdIS294fxSh/VaVa2P4lMSkXK8w2xlBYUdz40Q5S9iPsIZLfGZ90pSg6BwKk
O8XR5aRhhPK6lqvXOKs2dHRCLMBdZzHyujFeJgPAna53FPiNJDGHkMO3YB7SmS2uCYwH9CGQMNbB
WO1dq1Eoku3V4zA9qZEOlAFMlJMFEEdA24Z+Rw1clwuiUrDJQDhlByUZPz+JamjQ1FkeIauFWZBT
w03zEXvU7uJUHqaXTqLMuY7e9quHd8i1lVZGyZLMfw6stA7zVnkTGNtv9ZnlIa6b2AvLY8g1JZoC
16ZKaeVc+DmLE2c3an+t3KQfUS1xsud4ouOvJbTSv1+rM+LzWn0P8OMdoBlwgsor0TlkJ3jBYief
H+Xe53tSDpO/IEskZXaqG6i8lrki2AuOaXUmnL6CA9OitZaACN+cngxVFuv0pSz7Cu/3eW0+60oq
qsYm2qIVAoGnOqdzpCOGinfMjezWdgdSPaYijVfRe+L9lWrvrNqNCkAR+d2J7t0yutiD9aOUJQBs
y/L+zHcmWc3kFFjVBSDxq1i+dayHqrRHcaZ3BpHpI2vOuy9bptBFvt8VG5tH0EjesrNxD3LHaU/P
gajjIHMFsCkk4WfltZD1WgQ4744BRBk5u3/CtHrHDUKha7cUvHBRCnF/l+fEkqT62vfYk4Ehoi9f
QMQj0w+VLlCQvCLCyAcYhHA0MscJo2zpCOiQ8LSDUZ/Z2A9lQ5jDGvcyf8c4VPILWT/I0XmHh6N7
7xux+qXQeLYGS1i8biVLnGghxVfgpM7vYnVD+OE5VLI6OY3+NLjtaVbxh6mjTnq3oQb1oRh7ZrwZ
LQEknZy59siG1zLzdyTOBSk5ST5AqOnQspRZQo3x0/iJNYD2QdEOr47tc0IbSD/XegLhmfL+xC5z
4jnlHS+G0HDg08UQ4dgaFECqfX8WrDx1LpbZMnrs3gNZp/78z74joGOJrPSwVzjp/I4a0Rm6VsKi
58gLMBLA/sH4Atx2JY7MgVhIaxu4eq4xX1dg2LtXRRh/TqlSR4MsH2s8SXVor12raL8+Lyo9DccF
t7rXUm3jmErMVFocVhF4ADGfyjnuf7iqenNMEyx+bpkIm0TMiup8e3PZfcLULER8BAZJliz93NaW
5wOKYkuYdqPGEu360v3mRWiLAtCu2r+qihKeYYYOMSJe8MEtZ4xhyBQAwLO9U3WBzdISvJcuctRW
/aI+DLv/VgzSbp0aP8M3a5zujfMZUFdBXLG/mnSMDgKV+NRbYkkafBis7PybexTsddCi+jAhHt6B
spYUsfQbNHrBOyQv4zIRAMQ5gyAoJoy3KjAptUM2GbN2G9GTkOYRNyckFcp+E9Nw6n4xGYO+xLze
60iLZ7UEt5bcoitTDFTm6dCA6eqpU+1pd2JNaS2wrpgN//xwHJ/XzA8/2m5M/jE7wlHZ0uodJrN/
7pyu0xwQr1mzBkdlSddgHrcgaEuU2DqTEvUpX9qIsnuPBD2Q5dA+zKCRrvDvW/t2mOUQ2mXBu2IX
1M9z0eZpgQv2CY8HozYhwrvzcqgZ+uwbrjIyJaqARbFEucDQmE8sZNHagSwdpQjWZqHzvi3S3jne
ANxdzPR6wf8OilXTSY+gxzD20FX4KQudm98yR3xMBRqT+nEszNuadBDSTTDyTqua1sPPMqTgkX/q
LoGGqX6d/Ln2Gs+CTQisx8OzlEeYh+rqycw48ZQXfawiUERt2uGKlLZ49BFRoCP4lNMVDm8m3jnf
olTiFGPZ64vkHERPqiHGt19doLMIOEnH++vjEtqs37QL/uoihBK8kMFm1jYUrgmwJCS0u9voj/R8
XeIXsAy64RmhixfxrpDsSNHKgF30ppTDSztI7v2TtNQdvm5Jd1/KQ4ow6ZVFjRknAx4Tnae1Yr+6
MsxwdhpBV4zzYmEsEaaCWkGSfAlFdn3Vg/5Vmsk6RhyiFWHZQpxDtkAk3KJUQw5ExiEHjgY9eeKO
4KbN/yBpXSazAZ6BQeggZKr6IoFSWoJaYv4z8eylNQwI0VagmNDE+P6qSjAahjL43wqHP92/+1yW
eHrZh1266UqHdj+RuJ/rJbJGFRzN0DRkJs17C+rscEOvc+RjheRWDmwN0Y4b9ptifSO1AqOPSnXe
mjHKQQ9tnE3lA5AJJwRmhhv9LvobNphhqEC2eeox9rwzKxG26u5iEwtFFUfI2E9sAL7Fo71l0i6d
E+voDNF9P7hEA2UTtxb1cJ9Zc0bvMr1GWT7+M305++XuHAlmkBeFfs36K7OcyTdhagPgrl/Gcu0O
aImvbFbEoK46DbVSvVu4j8f+uDIAkgK++dRWHzAlFGTcOkyZYInDFPW2W75qmEDX1tmmbFwnNuHF
ZjU5cF7FsxQl+DZ5ssoY9ZRB1frsUZxld5NzR2slPune1a8POKPKwp86SIu1GaWlr5dmK6qM2dBL
mGPNZVtqsqedP5zMYGuAeMt7CE4rsO06Y8mqKFIdF85mQY/2EMJzHmrXkndZZCtgaazRVtXirbkD
WOyj3gF3mA0y1Zyjw0tzCTSm5T6IphXcUrLaEY3RpV5Z6FVG/0FLI4EHzI4s+AS1ZgwbValhMNdG
vDqExzgM8KOOlraO80KvO/mxyZ6KdsjpieoDHEUyar5mJH3/uBBn4ZCJMDearXMFFI1HeLpKjniJ
UhJoDrrs2Y7pgQh4LvvRPUFcJ4vf/4EhM81RRX1jSCbquuhkxNT7oHMjrGhOhoksybTpb1ZKZEL5
m08kgCg/TMqhx8INHjmdO4IMF0RJvDgQfUaaavCm6N3DXi04w1XHFcQubUUwzoBUZqL24XzJEaz+
CuRzxIUbIl+h4w/ikbCFyTDTq+nJa72+n8M3K6xUrzfklJges9ffstqwnzOdisF9ycgDuhD696bA
gyGlnUDtHLnL2bOsLnpxsRqX8HftXjD8kYJO3zM35TErPU1lavVVyQGBzboN4efos54gdwHfHte2
YiAGKzGt7LZ4jgLuOuy4LTWAJ1vVmePe3zUiFe2i3GkSDioiRh+xAv9hu+Z2hsvqynTuPtWXXn+T
Dof45aqO3R1FEhEXa5UyZP9P4AVSlQXGf93soKU6R2f2c4Wvre4gvMebWQ4nwnU87mnN2gnUyt7o
XV3QWUYcX+USw+4qoMAG3SZ3rd7ljRn0qCJ3I8p72gLZl4HYNqZByLmq5pGkA9PMMTJNAHYZdpHv
o6lVjAAhzQB928ueqdDHqBO5gKcqrxMs4HLEmMl7Me3JFqdohVjf6onD19eCb9xBxgWFl45wj8l0
pKdNC9ffbCBzmeCvUOpqaqG2QGpdTnEVKHq0WaoNJLLA2prqs17m53+X7Q5EtxFtuuwhhdLUBJJ5
MNfjqlnX6bS5MGDHKVerAhvwlHIm+ghKBXge0OxHesdHX23lWV972Ml4WPKMHicpeS6nolyqsGQh
otX69b38g38katnlts22YCvIgC9bSZJluT0mX2MZzssYoDl1NMEMxxumlBJdA8udcR6eQs5NJs+S
ejQKvXg48OI+A5N3WadnszNrrpdTCUa0U0snvEcietfF/jPHpHHw0HXECXxfgPeu7ZsreWPENN5B
XPRvfsF9EVI/uIFjwF10jDZXHyqKZ6nwX4Q4k/m944cOcCcpTEm+H4xD1b94eUWCkfwge3qgzBau
Fp6LFh720VHZDScoZpX2fz7VPhpzjgunJ/5Homf67yG8hFWf+eX28QUVYRDC1UK+OP4Bna88Hlv+
ADFAuCQgbx0oDdZRgzGgkXcR/DHOUqNv0uMXOZ28usoW2/eXGJkAGw7rPhe5xU4jvsNpTfCS6eKJ
4+mXV9WSSJRsNcu2LymXVqEaOpAxOd2JTp9eO79OPoD9Sq2vRFaeQfgfAiSPlZ3iuAf2fKZDBgTl
VAx5Dc1J3q27UxkN2+4k8FIsG4pNce2XaNIhQ7NS58W/gGN/uBjaSDTVJ+0MndUaFXIAwsEiUEZU
eynG4aGUK/sjJ9WhaI469eoUmjGYzM1cZa2d+i/DkZU9HsTJFBwb9XvkR4O00EppsmJF12xuP5+A
Huh+1yI5AnTfKGCf82lvS3d/f8Swk2EyICagKEweDvUK1Zc8Ie4j+917RfJC6vpFUv+DDiqagRZ3
NvF5gYNlM+pAU6MRxHY4dm0l5fWCwwct0SOs/trxjNiJDNXKmK7Ur32OuvzCIMWHVbzBrFLdcTcU
Gw/EK44eBhBtBtMCbatBKqZVSnPYv+UIGbrsVhBW4A0FltscdlBBCP5ULwZoZyHfSNxgzIzURNNB
Of2Zo1I/jNpSq4+4//O29ODzmK2vWFHmgDikArVVLt4K8nggFMQYJmhO8wPMhrsXJN6+1MEZ4AeT
8ihyH6a/I3DgIMjYPQdpnyIGQChfdaHtUb6Sumqn2hWYWMv7Oi5hey4Ny0qyl21qeuaZ4R5XKKBO
t/lC1bD5Ef1wHIUyTkQHolmi/kGtRe9tiSmBnOLMKJpWgOQ8jz+KhLmZkECiHHGuJQYB7CNkQgvx
AV1BQz7cYORAiIKjM8Ez2KuoxLjFLIB1mbIeSDWSJQUVXxo8bZq3GGm6co08XvRdUn10StYRtvlv
ZhubH7jDIHUQHCk2GASOfqhgRR5dy4EG62JdoHCM92BhBOr4Ug0ZjG1/2HFIeEZZsA0Xmoz0u1fh
1Gjn/+kEeL5Hi5XwOREQTXWULEb4ol7oHBa3i/73XSacLX7852Mrq3q2L1CNfGLFkWtr9G7JNKFT
Puc9j+qAOF4frnoakuqWpWLhWAkhM8jVomEmrGU1kwaUvrDmuBCPoWhrJnBoHjFiHnupLJgrHimI
7l42iZw8yHf00iBo522rCnqetqIQQMJC1JY3eEwvTosVYc1G5lE88Q1Ev39hWG6xmZfqL1nMOEWl
/93WEui4DosXQVma0p0LbJJavohdRlE3U9LzOQ6bLOR8updS/WtNlEMz1X7GLdxVGNh3C/jtZB1a
hGW0+CmgpZ/QjpFkNTr4n29lpwpEvouyflf8eTobgmxpwyeZe9AoP1ySYSyDXpGxCLNpkRA6Radz
UQOTkFMZM/MwAYTgUjwBu01ZX3LeCzELeszfV7CA7x5wCv5cp4Lkt89C8WurCbQnaxcN3MbgcDol
YkeivDvdaJBELctLIMiDkZeCui85/KYdQsLubDHCF5co52m/hY0ckibEyC8rNdnLoMo1OxH0Dp0L
yyJKCoAPLFDYi+FOZrt0GIL4ehmv/1zZ6ivz+DQ8P9r7rUYcZzzgS+1IBYpvnppD+kVQsQCkLnVR
vLFBBIy6ifYZ6Dj454O8xFvYIcIl5Bv2BRmWr4dazgQFN4uIJeZ7xmsxX9WtZZGfMxIKdUIlS6St
qRYT2+GBL7cpBupcsk95Vc4DsI/ROLKBs57A0AKKG642luRczRT4uTu5hJpKXnKzXnK5ibhIOTKT
UfM4opAwy6qpk0H/MKAr0nZKrf9MLak4RypKnk1699KWteL+4AOZmn5+FUtfJlO1XqO04A5Z6MMJ
plLggLbC4Qs/pjHeUJmScR3eF2Hh+EZQlAqnuKB/xOzfN3IMl0p7GionhGEItGVS3TABS9JVttSN
EaKQng46zgVn9zdVKbqKmcwkT+ZcEwhMZAA6zImLTiVPRheD3fcY1QQQURYMcid1K/RhQl58ZAW2
TMjR6B2fPRwVEt01XI/xNeYNkFcSjfc4naVt5LU91foyPLNuffI57lkQU1NT/HohRIn96tDvpAEf
6etRAvP1HiupLUeYn1tDxfh1xJUmSSiDbcfaMJjf37+ZfwfMvVXKOrGR+IO7HgxjTniad5+VtUnU
tB6MYcBB6LVdfs2F3I6iaDSmkdo53bnG9RVL8I0sVZ2sD5sSxYyaO/wD8LvTRKcQK+8Bm4FHxm0j
wn/letqwRjuko0T0PEfLX7zWswJwygkV0tBr7yMld8uZ+b1hoSeYTP+uzpBsFmg897mM6/WTqr50
eT91p5Sh1sOvZ/o61XoZonu5X5g9iIALmH075roQGQe9tQbEjEfQB4AcaJmPoyRABM7Oou6NaKMZ
qZq+xf5GCfd9oalcKM7pThanS3I9mEWBI0DBvTy9GXhbV8qVvL1/FePGxI5mads8ca09ekh07xMc
fMynbQ04+S1RUvJ8Qh8gQtLKUIMMm/vwHpIZdS4rjP63Aj82WCbxUPJzmD3dKPTTMpZ+YnUzh/3u
uSrMG4Js/ar9kvvyNk7sR1limJczHd1aV4mUz6bIbZPfukOMM0urXQbKZ/ZXpOHQg/1bN6A81SeH
VzBX8UeR3HbSvKBnQFB282iVBWPj6L7JcMbiGs4M4+4ooVCJwzlCjfZy4fd1M+iIi47wEDXqcBjU
m092Sq0NVhEwesfv4rL1cmGApl+0w4qybM1XvMRjttEQiBLskWDsp9zkUMdZ3Nk90dPkLb27tTwt
XZbznms+CVV7sMzKsKblGJDlan2xG1eLXRnSXnAnCAdeZ8NvwkSvimcyhX7yQp480aTfChlA9i4S
G7CldUsU5FmgYMegjLMEpE56ijMeI0ejzcH1p5lkchghFvucUUlmS7pTjcSnM2biWxJP55uC/wsp
+Hu5FDt0qggVt7xqnoj0LEZzOte8pOzzbkvRHc2WTfkByAQhh/c0+oqR8GBSRs4JxKs3pHTbWCXn
XkoihAtKhZbVusF4kiGvvXompneGEBWlHnxTuUYSTX72iy++luV0UqXs1SGkxHLdWCsZeU0LoeaV
JpZQHd7xmUkY38VwwCsXXJOylY5rf+MCzBbltXlUJM7WwJmIeWFnfhSqV3ua5pVbqtLYvOKeZms5
M0E/50q8W1kbF3p5MhiqpNqor8uaNMD63f7ehTfMH23J6E5JdQOB5YsGcZ1bXT7JPy+OYKHiwQ4s
q/IAKKzEulMADW1Gp8WqZgA3IsEL22IWPN2hDjRgfItZDm6WV5O70oGWweXEIuBwRgiZlMAq6l7i
XIl0EiZuEwSFPZGLIGBI2dX9QtvJlun5cUuLs0AVFBG7mhuZ41kni5+nPJXDr0NWjRPS24NP8DQW
lNuI2HigPlSgKOp04ljdB2ezwhdt6mTs7gtVYKyviDkZ07ynCxawutUz9AGNfaU9ICgcNM/ukTyf
o2Twjk7iK8DxLHQTFOEnc6zJZPpBINxdIFzmGsM90jkf2y8MubdNZCAUMjZEanHZH+SYTOOlzRpz
0hl/874vue+4zpJlo3WJ535Vu7tfeP6z6koSRRq5zlScS3lcQQJiiWBsD7ygmtUvVzcsmQg/mWCC
7d69/ZDhdmcaF+AsPWr1koGrAIIRSB8CWDy2XYvcpBMCl/fc9wkl/zQJR3MgqZtISXubPIw6U8P4
+7Wsj8nzuXya5a7gvED+zkV6vXlJc+A/V5VCr2lMIFuURiI07UDNhYeGNXIVRtFZCbcH8lIG7IZN
yHAdCZLlDoTqcWVXmjyzPhWd/MYm1bBuKxjasx/TFJO9O2/kv6ahV9mshGnRnkrbKSZjVDOjzFzU
LgA64fzRkacZYn04ybuH04JKQYl+iZns1tm1aTVQ0cPBRtpJ2Hv+gDDNmTp754+wErcejV1WSO4p
ZUArqIgrkbODqg9QN3pTuXtP3X9JJv8TlQEMDjxzCAoKVKAPNzaoMTTCex4Y1K3eR9acnngGi3DO
Zwr0WaUcK2W847ucrko+cqxmUF9gaBTp+cpRII7PCciqQu3zsrK63a0rGL7WewCQFpkDei9po/Al
f5t4Mhn3TzusHWoQtyvk+tce5+/V2HnI8Sd5FMTqtR2+9YxvTLLWdz7f3zMyDc2qNN33GqZqjeFC
2Dmy/ETYNSsrqvx2DDsJHCzB594oxkWZCRXccojtD+77bhNWibrPfx6M4hJVT8cTjKb/yaL6cz1I
C34gLPf6VIImbpvXRGmrNbxDrzNNHAY0DxX5gPpfuYVbzyVRycc6qoI+DCVZTC5PxvsKPKCsGteP
jgu5qgFB4UIkzDBtOcCQbwTWxcrcjf9HPCFM9cpc4d6nrvTGSnNvRPFLiB+3B+hCA+DbyBVMDgs6
zifv0T6IZHb2lhKcnvkWngVzF4z/KW5GYEyQt5Ld2SQGPmqCJSwOqNBb00p7FhEGZPEz8HZTC85U
MqeMBXiLnMkgQPvAaThB1M4G8FDlHWiQEY5SlKf6V0toKP2nisSRLi5wKBqd4bzrLeTH4EvcQSBG
nlDRPsWzzj0CLZSx6C67AQsiV8OkZnl4d6kL1x+v1OKcLRI8Dm3vPM9qrPljliHz91iPOMEx4ybN
Hf95bbZoLsONs7uuGqLEp679fvaxkafEXnFrMqxReCLZ2QD/87+Pi0gIX4DLYPiO7WGp4YECEG5p
cl9S2AuTsQauuh6zbxg40qESpYadAUMUdIYnwy0cc3kuXjOndAIh14bYYw1Uz6cflx++MVNn1NiW
v/FdeB9/xcH+bNEH9psU2UnfV6OIomJ5luFtvIev92U8fWl5J2CXRoq3a1U8OggmPCRROFSPyTTd
5Hbk7Dj8P2KxJ05/xsoTXeqjbqSbxWx1yF1UHV8CD2KaXGkZXC+xDi7/gyt5/zGu2PGKYGnQdi6r
oKK3CfbqTUiPqilq/qXScH7azZKecQn2MiwN6zZiYtjLee3O2s1yPeidux6uBOGNHabYukIHlfCC
I2L/H6pnqh3FiWZuwmUxOow7tljRMUTvENycG/b2BEtnBJHZPcVHWzyvFKEAeyCTUjkKydEwz+Fi
Nc9n5sD5q32WFrV5kyQWHck4ORNCalqbX3AOxHqY6k6+9MLFZGe1wo0CkSGY3yoHeA6CpX7lUTnS
GsN1R4E6F4A1YuPgFu8ESPfYu+0PoOCAJ8VZqm9LId71XEaZf43AXoiXGbvif01B+RAJVCOVn6OJ
DZQu2NyhtmeyGna88QneFjgArEmLiLT10D7m0/sioflJw15RHNTXExIn5OB0AAe85VGo4nLznGUf
t11pSujd3jB4bc/fvT9OA2MGy0CH8VuaDyFtun+GSbmy4tD3HDkTF5vVgLX7xNg1537HV8RVhqYO
DR7o7L6VGlHIhOp+S6F298X7yzqN6kvS+haTnqfz5bsuZZZc48JGYZD7X6RgZH4vraiTlRO2EPaY
H2bI7ch/fnBXXKMOrePCe2b+SUkVarJgZ3Q/JaxIPzdgl54NwsUCcNQb8mPemUkIvVvA8JnfWX4w
HymuiRaWzW0OcA16/BtJ7laNwqQVb2Xw2MbxHoz6GK69UyQ7/HmIYqPesf6to3GX9GPEeeB+fIxw
pBNv7/L6Vi+JPZU6Sx+Z82vTsr8YI6EBk51CVs+Wk/qNSgxpolgZMjUJGpbxqoEJsQSRK4UzHByr
GoUHFRBCRp/dZbpYCiCv2mNPyVl4WfY1KMzRHziqddihTWokAfY9khJhKbi3DKKI9QTCSC5NZ5av
LVHGfKtC3SVFxO1GmJH25ZRij+3HE9Q7mmxsP7ffw3lZ0BBwAaxfqUAsPOPBBjoyumVeoEI4lCFb
5ljx4JGNVdOau8mdmqzBoU+NivORSX1MxrHNnNFmlE74kp4kkCoKmeD/bL2rGTCgQY3kOt5/YSc/
V7ms4lT3qqcJu8nZjWdTN0h+ut9TStxzzDJzzJT4VjhuvBKM9DEZv78rcPkQYdaRcn4J2SDxkj0G
FrW5P5i2EkhD2fXh7DHIxz5iatO4qBxmRBd8BS2Ehz0Rwm7/GK1nSFbz1fsfrfNbJxUl7dUUgYQu
Yj+XbSd1WOmIvtKnSowHsMyBPndyNhcENmgt/oLpqebilXTcuQjvUPuhAuvjCy2cLxa1tfsASAUD
GxJTpC9cUODC/DufIvsEcUSyVrJsb4ayX2f5nmUdk1B1pBtyWja8n44rFvQ/3Ecf/ge9WSc6g5Km
FohDzvMjc+xFYb0mEdFo3RfKbGzsp3R8aE0SYCJMFe/GEJ8JuIKCT0jElztdD25dzv2GlWspG8HQ
dfMJ3U9daFhJl1LnnK7poQ98ljOaRwk5Z3TeSfAfEME8Jm7LiAab0hNDK3olzp/K9c17szLH95xz
pFZoOY53VlmQ6vzds67FMuoGWgLGu0zXRcA2jwd7B8MFhVzied27IBcgf9CNK9OGpXBZL90cubvW
B7Gp3m1Rha8DG2H9MZAjMKc1ADYjzfxuA/5X4AwT/ucIY/t5mHewtrYy7vKoxvtvHzzxDLLiRoES
egaMOso0wfUD6SXlWKPwS+D3TqkpiMZ00YnInqJ+xC4IwMz9T70lQ85OZ9d+4NjYWnNS2Ww4S0E9
XyE3TwHtNYlDKYBDBWPXOblVCdUKME5qjxfBD+ZucNapOSS/TZJm4VhFrPWYABBy41E0HAIoxLBo
yQM5yE51xWlzHM+9TI/YoGL5RjcmF8HDVdHOIFWDv5kSuSBUVbQEubytzH+zFNwGs1JeNv3vINlR
6sOvpmY+Z/WqsLnUyDEajqxYzKEp3WyaEYnoghvW/lHQGDZEx3XWDZ251BDAyuwelaKAqCFXImYQ
HJhX0CsQ+CptPq10YzF8P8h6+uvkErhpAw/ZNvPcfqgysRPztL1mWZ3zOzm7CCxYR39hy39H3hXJ
cCYb0ERDSd+CYKBxAFjKFlztiRM5fwjPkaneRpa0eFasf6SIXtfCtkWS4q/Qzxv9xjebv6ZVsJTv
eYdtSu37GuCNthLo1jABiyk68Jh1Fx3WCI2R/hLphMKVUMshLBANQ/0o9RRebuGZhf8wfYIvFyvP
C/ub1GwVoFuqMBZrbAc6NjBNR18ayJocRWvjlWrfZVWZMoOUFkiLe+lPyDs11LJ74OrBnzxNjAoV
x2z257qK3tuFLHs/9sIX3Of3JPy52MRGgNZwY8z/16PDTughFZ/qzRFfj6YW4nTnZKjA6RBl3pNk
qJ3ITtCMFedCrWAFP8/w6T0V/+gts5bdEp/CV3ldijh1ywMlhYQ2ZkIpAgK/8dC+DYhoQhkFRSol
IPLb2YzdS/F30NF2O6wWbGwAgw2b/MC/AwCBcgEcNnAX9DGjg7AhksHSNA0ZLW7UItAofypR3foj
Mopeie9mBI1LvkHGuxnS5O/rAyhdjExRnIhTy7sZJWRSGBCqj18oIE2AxEVHs299pPyOffx4U+p4
0p1owdAyM8AxBX1J27ex65F3KIKcesW+98ZOSBF8H7gXmR/gRDwZbLinPj60ynRsYiUCsQVt5QPw
z3VGyHV5zNwiG1nVwlBnxjJe8zISIHTnf9Jnx306SB+zTWbliPV4pII1p8DaCzYTptcyqGvReY9n
KB3+fyuyInSVdaWXYHpc5boY7QQcI2rtO5r7JygI6p74tdaMG78xxCXALMgHpIkn8bGWEZ9/mH41
fsiCggecyopuCa0c9mErzlLn2MYkTFJWvjvlHuHi4BZ9FTqS6lHl0vNN+6s9U6zD8NT9yMZB4Q2I
eX2XsRn20AmXWEGGuznlPJaANy6Ia57TDaf5BpErc7nF63Gk+wdRBj+lBx5T5jTGmPCd1fHOigk1
58vW4XEs8Z7u7e09Y2MdGtj1kyvDNPaV5GbvgjSvY+qd5GsZWFN8/awojiuP0a3hfoYxKukOaASh
0Xvd5DmsWnU77TT8buho444GqvE0fRlWRZ1n3olIT46hBoI1X42rOqhP+zWbDNeAjw7IUvAAOEYi
HWZepY+ciyjeJAzP4AYNSbaokHtoPxkqh+keYc9CMmpB/dXJJWbI9rZLHtjlY8nKA+bNx+DltcpF
HV4wCE6wpfJjPL/NAT0I6122sjY8PwzXJr1ecCi8fCl0bPPE0qypsO1E09RxZm+Xks+2OR25urSu
9b29XbhaNxMiUxDNxS2GjHlDN87lwAe8k4qazOd+E92B3PT5ApAlo6Fomw6oiYo0sx+NCGiJAt7W
MWf7MoFCFOun287Y/qs+Aa7Euew9JD0eYXZUpkmLdaI/Hnk0lsKYFoBaVqafZKN64TErN77faEw5
/c7LFBEg25FHQ6sOP1eMnE12VxBtAk/aTXl9tunWUqGMqUpJkOgdl+GDz9iE7CozdqnokhhfmYRe
mTq4NJLcCouESj6jIrpFLNmh8EncnCXeSzbKcM+7A3UJ5BLKq2EB2+WwdbvC51r5lPA01HqkmLov
aDI8BtrvZrDvOBskgD+jQhGqz3zVRnacywFP3lSACSISB60vUaOM/RBtqMJhECYX1xVY5sJ6a7R6
db17l+/gGTGYYu9Iwa4LU4MdW70Kt/ErGqFDO3VhhksCweAiI3Nw25cv/rMK4+uKzmmtbMRb4Bb6
Lj/M6llhq+/HN+k3y8uGBvk38sng4BtHiatINivJyCMwgvtqz1bBdwIAxD1xgqtslWcLiEQRlpTM
mRPeylx9S+KrL5nJJ95SsqLO3H6Fx0YvdKRFNkyWTLoYJBxzCNFMNuBw5X6VT6LR+DLJ1JGgas97
DhzYHA1eLv5XkfaLj7ojM0TLjXnS7fK6Sc3UKWsEJ5pj4SgAoFSCaHs9PLQxAdtWd70pS5uBBM8L
h1m24FjuDpxzkj7jv1H8QrIFTh0u7i+TfaRuPNzs/oc3QDMnTH4E32iAwgr/iLItX5PaeTKAEgqg
B7/annEXKW4vQ2bMgmUY2iSwyXbWEa9WIBlTgPnkI0B5sB/fpaRlk+B97YBo+edaXVRyBwc5d1y6
MVoqEqs1jnT2pYlE37XYVc8TuTXxvTIHfHE7Ifik9smXzs/db1K9iOx+dEoOLPj5eKTroHHaVvnZ
NTh41vEn4DSMhJxnvhFfUs+LKUi4KA1H1BPIM5KYexnC3U2u3qyfRqqS0QA2qtZDN1lpODJJ6xWU
bZWX4/0FZ4cGcYAV0vJK2kpOIecoZR1bbEgFu6Py2JP+nkybsvT9nkT29rdx/nOy5wHow8xvzOxv
Vd6CgaEb01ijtvsarEMMxPVji38EEmtu4R6+C3KJ4w5qR33nt9V68PvgvgV/SxY3ZF7rE/Voyc3O
K8Ehj9cwTncYkePurq9yFTxDVEeVtGN9uPL01J/QvKJdECcrSIgQp8ZdbIciPWpEuaVe1JGNgzNj
ZaFL0ET/hVjnwqkMwibPcaHCr1TpYiggk6jrCNSuYKw9BgPTYmDOdHRMH0ZE0yP2XPejsENaWJWl
mz7KfuxhfawJdpw8sofTu4gfHg4fDF2WN3YUmmhJXTqsdqZEllFVHZCB82CX5B/CpVfrEsF5KOF/
p5DHHvqSfwYLkmz9a2I5s/d8I68I2QwJxmAiCgDban4rywZUZRM2xn8e/dJHX1SwbYBrjon1vnQm
h0GO1zMOdpBywUwG0QcOkHq2Ae7M8SOsoqUfk+tE+MyslFgKf4+uZSgOpGc0fogETg+0KaqD2JZo
Juslin6ceNKhK3GySFKRaI/lyAHMil2+LYG0VlQu/JWRNk1+r3JqaKPobjKnNT+m8bsHq+lf1MmQ
yPPlRsMbAWiKOQH91quVzxCdu/Op3gYxFvPFHD3StzLS6f1/TTZPxfaWMJBdu5k2vVbgexqS0m7G
/qdrljydhZ/TcogCPOOf2NJRIhwBpmMflOtrIvPoKs3HbtICUN63OtmxiGPD2UcvRqVzzHrhkMWS
by5aoesZDDV/zppWA9xfl93LfM/S240MnVxllFyGHYXUPz2tOVuk2Iyg1D8TGj606e9pjAn37EtG
Oz1nL4t6D1WVQ8pOxM26NfNfsGF4ea8kPgrIokLLcjRah+oWhzsldL6N7w+KvmcMpJ46zefiSUDT
hfFelBd5GySA2CEBB6i1NO0fvsSVdVXQwDwBNpSSE7C46/sNXPDtEoa//MWrAusfnaZsHBzvpi6h
iIjkYlGW5thUCi7rPUxZm5LoeY+fMjOr8bKUpWVPn/4mHZYbHtvaEssmr3xnV2l7NDRZtw/lLdmc
9wpCCU2Dz+u6T9+REN6nBrvRhS3FVNY/f1fx6+RBFMU9y6QdwczWK6hwj0FOYLQ2cmz+6W0A7ICP
Gh5tJYmYY96oT3EANb48nM/ecuJ/w78SK8wpstPRCVn07ISUsxoBguQBij0mwDfDLVdV2RwyU0pY
P4PEDJnNz5bWLurs28fTjRwMs3rkIpFuAP14y8AMWGLhtpQ+Nhhn2hpUlLMMy2xlvFy6SNaySmQj
aEIdISoL3t6HUNmTTc1unuQMlAgsUP8mdvJPtzidvtah2d8jA9ois5isWLIj9WBHY+jAqWDYkqdR
6sQFHoLhN1hPIMKmRUXvDTrfqi44oKq57pwiGVUlDlR424GqBaADiRJ4uhu/MCK6JvYVLNBDuUS8
GbzcgahXjcUkBAYA1xR86ByJv1ASBxnk0JzgMoUsJsJZNwnkXhLB6qR+pHn4khvOTXDRUFP7gt2R
LRe57Bqf7rAcaMZh5bi0zemQQbuz/fsRwoWgCTVA4+6F/Mpt++p3uP5T9B5+x3jShNJumEzJqYzo
2WWGE70x3j+N6XtMGs0iHopTFjk2n48rJPqIPv5EpYCbac5uCfYVMMpht0/RGuEyGuYa8yPIztoZ
9adGnFbeTTkvsYO0+cMiz5Z9oXrYO0N2jsBRPVPVRBb+iKz9blLTOA+7N8HSZqWXO7HQrVSopu9c
IqSgmu1dfkWPHgfUd7tJb2g7yZlmThAFD7KCQ5Wa0sQU1407cmudD1hhe9R9A9IsXs7PmlsnC4PQ
H2ZI3LirvySA+3f873sn8xBMvk1fu5i5hpJLFO81u+aoRK9HQStIYstycGkiQmwQuyNNOrAPTvYD
Q3NObW+H/F0DyApMdfRdHZa0QciSXeXwcx5RGkVyjF7FhyUHRtLw1Xxe1TAfWb2/g71agqW9YfIH
A+1Yzr2ZfpvlWuhDcBdW1DzmRH3/T2rfaEbuKMugda83rubSHN4Aw3dHMdGlaZvx8YtkQ+fHAq2Z
fvjdKTKs3C/psEoJm5v2T0gV3a7oKdXFQ4SFSjTVfBxFAO3fS9YTOnVp0/UcbAtrB7VYuQSO9rMo
1k0eTbtbGCMowlB6+zz7kJV5YZEXfqVb0HadrlSCeJC4C1utGO1X5ufuLr15slTTdNjs80PuOPwf
VNPruEJFZ8Et5kEe5T9ehe/KV2IAqFt+stUHrxbnJoX78Llwrl5nxEED7LDKBsdP+bdcczMWFFeQ
Hor4Y8fat/+eA1mpqn+COVIwYLx/rCHDIUIw1qLRh2HgbFMHwIs75TgcSZOlzTSr9RUaeA/sEq+C
huM843cY6At3WiX6UhgyaC6Wx+KK+5v/3fHHv3KAbQ5kM02K6n/ijuUKRym7frtFTUN5Gedwpy/y
jD+D4hm2aYYMsDixk2u9I/zqiAo+4OaZAs+u1fG46P5Kp4XS1BdbFZPo6eUjYQLdaMIzUq865Pa8
Kn/lElwQxLFBg/vbpgkmEQRl8pq8z7N6Y5qEmBPTfkA+S9g5M0d6gEkUDwwuZTPNF8+IIX6If8YR
YVSq5SqyDDEJ17MHBOKgD6XvQ3VmirJxAZtZ/zv69xof7jMbS1qz/dLwrm9VnytRK+AiLc3MyKrp
XxBAlWSDnKNst2LpTNWKF67/vlKxli3gEl/N328uJPYVxTtqtk1NU7wr9erpOKoCIzvD+FJ+9mwc
zNKFxGJt5/TjusasJ1kr2NIIrFlnHR27/4e/bTCTiAmrzH/IPdqg3boeEF9gMiCgNNyMR3IUFqBk
Ti0dpmxDKqIBpI8rQrtPa4vZ3oS61dSXElcQ9LDm5MDA/rPIn1lkp/6L1ZmNyM+RRiUbNiae97Ke
7fKRETTskzkVDyTA2Rzk/tgS3YCSiSpQSl/7Gih4qbnOwf9MbFW9jMLOfQPV6VPXCs+CD6SA20SG
YnpCnhKnOGE3FgLQNDnKErQ6YjnSpmMRZryRYxb46vzgmnomKlJHVKDI4mvI6+SN9HMxogOY0YpB
GlmJNEHyWv2npITHS04otkSWg4V0Bm6OWyg74eMd20meK3UeTSY/Ix3VC+n+ybxsJ67DXZVQkUqV
uDcHhKQvtJamfXvZ7Fm+hMqN+0RPSHGqDDtGp1JNdQZpZkwU4b/vfwd1ReGF1Xy0VA5YQfzpi2Gn
HApx3dS679z98ek2P8HZV+HYveIMcY5lLPyPnBXPX0SLQ+tHzRDg8mh4337Y5RasdnXNa2w9KDKg
w0NXkrhIol1BayNzQK7TAif+QK9K1xk3FNLu4regswrLqEqWLQyxAUd3uMOXIB2h/cBH2IbRUotR
+xL7UtzgKs6kW9c1ibksV8hbupXeYnucsv65b3eLupgtcekY0AX/XbhrpZK1072LDsSOXpMF+4zK
fQ+a/UN87zGuxeR3+7+MQBqmgMYOh3/ergbebdnixJmXA10/pKOXZ57lZeosTlMB6GDTSpqCUerb
x15SObTrloE0R1+R1wjrIt2b2K9I0EfRz8i7Fbz+/TMbQH+CSsu4Xp/YMe6yvaxIVMqfWg9ScsJr
cSC4rDUX/mRh8thYZdwiWTb+iUkqq7ZOvawh03KYw2NrrXske1tHkyHwHS6s+mnGBl+ylobqyvL0
n/qhvpt6IGBuQ7cY1uyroNEoE2qmFy122YKaaQ/EbPx3s8KnF0asCyBIr7pM2yedTFxNLVtSwyM5
tkHJUvQD2eCePYgdD626Uz9DkcznVsM5LXKx8dYQ+x09FpL5ah6+5dgADMt2Qqp+FuWPoUP3eHRC
2E7ABSM8fhzxIn2WNO5YDiWPL2q34Q4Gyf7TjFOZSjr4jO6b5QWM6DTiXr+Su6g2Iyi1FJIw0/H3
xZd3JUva+4SHUoa9PknQCfS4PtwdK0zVqU9O5xrzWcdjJ6O2VHDsoJE7QmluHGMdSaZT+XSXFFfu
CH6TmvIbHdQG0I3//7RF1OMhwf21D/imLl0xH6vZ0KGX4qq9buG8bFzmmGDMRCcauyjJk3ZmYwWS
XGHwHixqDozcEiQhYVrEXgN6bBD8e8dEXKLwUCuixviwx2J1xrMRV4YYSC5sb6ywmy36UBVKu/pI
J/qV8yZ6PuA7/t6m7ODh4HWsWle9FxuPIhUZjYC2wW/bLohXNv2RYD90ODKDFnqkfNs1yEWt1RDK
bXnHpa06aVP0sBAXY44ViV1oW4DZaVhE1bgkTrifGgSRYn4jgWL7ccUigK9G5odVwpLeQoVB7j2h
ZvGiuIRZqApqdsksI4yRv/TFMij6mCuMVNa2lEf1b2q8vx9xR67To2q4zNaBd05Y9QKQpi1nXIFN
rP6peaJ8RycjoSrqxnSfX2HV3ZPxh3iWqjNItWpX60vDn3LzUKbJP89y6W+ynEtkCGmoWZAnDe51
owHey9LGw4WlDNaeWUXBISkW8wOUb9jVllQmu8YNOTbAda8WAcSos/QFLPmGQq0GGe8iK0WVgttB
lmGyex3TGJMFJ4hU7QRVSl0tcwKQP7qGRFh7eipcgK/YGkEiPvb/YuYz3u7VUjxrlPIRcvUwYgZO
9JoEmR6VEPKmq+h44wPMjs1A8GIUHixWYxXt0YKAzXeKyLCCN6vYpToxhc42YpnvWgIuO3jMMBKc
VRPb9QwgTiP83IwhLw5EbXJwHOtnuKUjst+6dfBya10NDtPjNDgmwSRMrUUhbdX0+ZIJC2QVhABd
BN6enEFQ250EVd2SiYac5YsdNY5O22vnBT+xHocJi2XUa6oXh3hiHY9UJZqJXPVkvyFuL9XIJrKb
3NfTYfryp2dhPYpP1hQEvdcl23D7s6vUROqyFzGmnrda5bbriRolgCcs4OmKihvauzoOJc8ol8T3
nH5cYPygWUU1nx0/figGny2e8qAQ6oYqIIYosrIkSw0VXmdqeNVDjOS4Nc43/EaSz9EB76F+FE0C
ZF9i5Lrp8iil6fdNOZrtkZpAbkFopp3c0bmRFbH8cw1PSINeyL+HpGPSc9YX2fVsEBMkjhsSFmF8
O0n78N8S6kpR1FYSdVV+Nq8MO+fYr3ScoX0I8jb5AkDonGxoRqqjuPyxzQNPmZIpEvCi/dVNPgwf
Nw1SVXhbF+BUZD7gvoEDvwM5KDbnZMw/vTaSwnONnOUP7b4olKyWKq40tTXJBl15KpIoijGpBVLM
5IMnH0/OE0g+3KVWF+R357zvzjRZeSAmcbzwfg947ObbHsxL4qpCLiIOZxe80rjtgbhj48PUlvUx
EKYSPgmQIm2OtVoyZPuAlcqjEXNIZpXGNqJH6xX3rkoLRrOvPKjOOOUHwALwYUQQdC5DwcSRcRcS
VQJ+ljqG72mzasCryYrd7i2pAHu3vr8n8XInzFIzA1Gj8OBKDVvbqlastzmcNvRwbDRh7rktmwgI
mEQd/l09Vc0iGDq3/RGYTbqzdA9KZFPnV3M3wTunYDuWnr+YLtTCuOUru3Jui6yD9lYhbKeSPvnf
NRP9KAMlmIpoqh+TC3HD19GnDtAvtlJkbLpB8XYRJbBIdIGVR1CMI9gxV1wcG5JHbGurP+YDU8We
vNcUNSfpevXE6HIYG1WzA02fmpx+P12V2sFGJ9uxtMoiuSNcvjiPHE/3Y69FcbOlxHvR8nHXkK39
2QWKiBDj5n9MQQ1WEKG/1i1ibRwt26VClw/TGeUSy1Diun49DlrRssxrIq0sfr1pUhFfpN1lIgaM
2RNbMKsThsO5QTReV26kBzkp2DlIMSrnbAtTQIBjE/Q2CAQMk+Sen4A4Yw5omLZ/Bx8r/plhPmh6
60vlHSeGlsyC/H9M0NPKPAPHjf6ZiiKQA6vqAaEgf+Q1rHt5TlEz5u3TVsBolAuvWiUHGQadt6kN
lu/s7zvibMzgDKX6ZLJVVRuOerP3CjtkEEKMVEAdLwSZD3sie9RILZ9gXEriDU7iaRQPiKh7GKBG
MGUMjbcGNXERijDJZ6qg0QYt8H+m6JkHhKMo/M+Bcjyo/TONnlSAz0ZuW0JZnJfdScXRapGcd7/b
HSwHoapYs+SO2WvSQRipvU390Ld2Mcg6Yi8v3l8ms9vgsObE4jerIAKlG5E5TRYCVIVA65PRbBH/
HO1pLsgVAjI1RI91jhUiDkDfjp+axrMs+kfiUaCc1/GWFFixW2HCvHIazXCd0puWdsR6kTg9d4/b
snP/AmEVBHrVxv054Ro1Pz+dXBT7GEJzZGM2K8FbYID4VSpz5CHYM8w2tGk9td/t4yooPk7LCxWL
1O9D7yGn/3nqvsLx2EJusurqH9EhCdfKT5/rTI3FnkoIfuFKeJhmeCzeYwNlsR70C7QCpOALUSXp
zXPiHhNs5ITKw/KlHthlpBsKH0dx2wOMb4sER2ReokbBJhsbHJFrfl6eqJRSd9APOR1qQD8qCN36
QWYjQqEJRrKfxrsO3vBbLRn6Qh4BC0CKGF2YVF/bYv1Y/5RaL6dIeQZrF+0lz+0yCWTRZ31QlbK/
1F/WxfZWauWgVINe7nBw9TlAFdwgqnrn/MzlCluobodkeY2ncho7gO8P7+qK6Pu7fnNUTyq7VhLg
4V/+BSuk6/mJx7xY+AWUZ8N+46HQR3TN958upPs+34gpPfzqtmJnJ0XLOMfrBHUF130QBHCjMCmL
Ik11fNCVGWx2fbDuv3JFiuVyZDaQFtTfurySpy8fhxHzs0NSvdkaiaapm+N49Ys0KknZHQolzd9f
LS323GQHwt8qx0HeQ1dvJRuYoX0GRFVB15XzlXO9QoltNqumcDNC8ibGHLEAzty5deCTK2iF16UD
gA2TbNpNb40+u+nS5GgNwcgL83n7kSJtnWbG5qX3b5ZXwYbszedYWbYLDnozFHjNEHxTWCmrh8To
iFBe5tGgEOPdsAVLTaHcqZX6QiEfBvPFeGggMYguq0QMzB1CMf62QqnVa8xJk9wMxu/YNzJ8byZB
SliJnGOuvBso3IKY9UtEEuxDOnFCnYlPLAMvA2z0Xn/vjqjNq2b4a0E7LS7zC1EegedFRz2ZXAuZ
EGIrC4jbzX4cgXV/ce7x1mwtqidaiEpzs2iMvQNjC7VyLxGpWWN6RlgpxlL5NY8HvDNUxku7MBup
MAFJHgJeOf92PhYCw8cWVgeQe8AryavNisJ0rpC+jTUvau8RYAz4ApjlOqbspAoZpELETpGpkCYU
ZCGWn3CdoGVWqmV738+hDe52VJ9CL1vXk2PWrN0rN+H+derNauIJbRg/B//9DvR2VDPXzcGlxQSe
PuENw4PlVv0ViFA8U66SiQ0RO6hYyN/DtJ/gOGgQCXqrJBtyK0dUYM8D1PEKFphQKBXgmtgREKT1
JyxCSy/KcIfW2WjYhVS3yVsO/f12PxV8rACFbNqz+tB77sM6LpSkC/ot8/zRpkszwKK5g6iJmoEI
LYxGFjS1nBRMtuIF+M+sjpeCvPrg8f08mCweyLJoOiqkN8CEANszi1FO++nNOK000V8PjECo7Xza
c5G95FX21C6EP+IWzU0778se+Xg22ChrUmaNu3cuceFE6PgzP61JbiUNyqZwaCu3L1VdsNty3sgF
yv0oKQQyZoS67RdL44LJ7tjaiet6X7kmDN6bizO5IS/l6JtCN9/TonO8f2vAQMdBlHDrFqy4vThi
jdgR97eaNlhFUmg9hIIrKAhVGrtCrFfrDk8G8r0CuqLUAo6X7fdbDWX+TpzHH5kS58lmnBKsLwuZ
fkiC3sS4+GAd9kPA2eUpQV08wtZaj1ByQ3RfQbgSd/3AA/jaBXQhs7beo9GTJ/CKjpfMZcw7zLvD
BErhDWOi/JVY6TRABV/glr5kKZUjgo7d5urz+us7jG/WUOgRQyq2FyCL725l9SUWT7jitCokwprA
6NufAn00u4P0cqv++jezX0KjLwwnx6U5qlI9/YeyYTYqCKMjV9hgCZys0pL78Duo3hxobroQhPZH
xM8KvQ47LcDRjq7kgC04r67MNspvpvxLZszk33y6UyJUcQyaTNlAgzwoOQTWf4EtiwaA/mAew95s
jkS8lF0qbm4qKUX3fuPPWV1xTYVzaFgCl2kkKg5qwVVNRkEwoIjL0q+m0Zpzq3M5kNKddx9mFwAa
2lFScexHqMXCMPgCX67Exe6NyewpajT35f5RMHSvedZ/eXbiRVZCCzIlEeXGQH2OEZpdOOr3a8qG
qgas1FfqPc/NfigVMg8ObUvsZxdc5x1Dmu6wNtvkafcls1/+AUFIc3iNRKXYcz3iIKAVJYGtBWuh
nAR60I0idrDsVJuuPmdwSEboKBu0aC9LAdKBC406hEZYF59GTAzaORSRBxkeCjPcEA/NdE2gEyYg
mzdIip9JVte42Ip7mYwF5QCBCSx01mwr2D+p7wjGv47e8gNajJAKbqBRBgohC+pEZFGTUKvnX9U+
ksT1r6YlGt7XOxMWG9msxBy+QVB8fn06rUW3GIN6bRQo90MF7prNIU3EhQ6Fe0kQrF8HdfXVGxl4
XbPA9raHf5FG7hFvaPS5MS23YG6LnT6NEoFCpE/zSZ08t+4AYudanvo2RJp7ZA9fFd5VVVewbTcw
LwzkNtUyxoZPmY+3tCTOz1PjkCnQTRHWH+Bl24UUFAaGRuWqjNfE61iX6oSZpE83iF2XcIGQtrs0
gw1hMfsbSmmIlNHg5179CNLjzuZLoMzZOao5LAvpTYKek7i6uH0g8quNcnngyX8lnAqJs2ohlJv3
nyq4ok63Q9WGOAZiy6li/KRp9A01qwA8KX4Zr3Lbgon+x/xizJC7Md1gw5/M2sCpcDCjavWtp2MY
3X6ypm6mDJvdy6SI6maHKn56hbIqSse+XtbfpOS5eNY1MkmgbDItd3J9TJzF76P5znbGX9jaPCxs
Cm3VhsK64Bcu6GgzFDw0LlCf7FKagdNZWSft+e06PS/+B4otGVK+17e9kpTVZ0K0a4Qu3BzlR+tZ
D8NHVXSw/xT2h4kM3mWfqBtlQv+gLk8lJ9wbj9OAJqUNKAh6isro5TQPMzg4lLo2dwf5sYfPq7CY
uVinTN0K01UcyPvxBkM6GMpB/ypHxE67zJkXD/8iB909PThO9WhGHsHeF0uKGAin/v3V6M2izvbP
kcscxYC1BzksSXwkdM0Or1XqcaYBb7GnB/yem4T/22i1dlWpSJSDFE6FMLufe4Wzp4DbbWeTaIFE
Kx+mcPjCALHNLWhrtbs4Zw2n2wrN1TqVdq79UMatTmMLrEMnC2akmKbunvFyswB82H+N8HrWJAq3
jjTQZh3b2Ej7z6CJKFkDbut7DHghwaVePBSUtB/pmL105rmNGglbtg/s8abntU17W7wjiL6JpW2h
5a6CeboA23fNRkg4IqPncclCSpisf+HxOWQXLkkyXxI6AEHuivtt/AFVCcf+aCO2m/3G+okrxqTB
A29Ni0VVxkv1IIWmp16E6orXAUsjae/4u09jd2vFzGqmZTe8VeTE61SHaYVV5iPwVzi3z6dEqf3K
68puXNhWqRSLpA6tKkvoHgh2ZikfB7sGqrEah4Ue/Av52rqq8uyWVEXPWahYIodsJjm+841TAOWZ
6zO7VQ3jR0nj5PhtwUTGtU2eTfDekfJYe2A/9u3eYN2GgYhFnF7liI84AxHDFVM8vt0R/2g/6DWa
WmEz6FB4nO7FGb32z/FH/H0kdic5HRuTD4Qh8fAcoxiiXQX1RLkZZI4lgdEbKabfZUrpcYh8bTLT
MHSfnq29k6fPPzclQo3CFTX8/qbAqI1AbDuOEDzq4UQWWAFOuNsHDpfa3HIcZb+1Im2IwtxbEyGc
kUuWQw+dzhoYZ8L3h8jdV3/5pkUfdSKilbhgoIQpY2am50+9PCYTsw1Bs/Xw9d3Ttcmz6jAK6+mq
Hu/v1Thvir3JtkiO43mzDCWfxojoo16rDwldB5LjxFqlr4XVP4QlB4aQiDicYAJJIEykPl9X6Ds5
VyUQoqRacVTNltKhCLhttg7d3yVE+3WswWlJ0Ot+0Ee0HyZ2pIsA1vPRfPQcP+lPfOoq3XXsqYS3
dt+YzQa7L0tSNCXlDWZ9tTxSAd/gDuM8DlCAWyaiEDEwMBe5pWzcfHpX3s89HKT1YQ86+rjTZp+J
Qp2UdZZbYJ0BySjAxYLBqn6kL+9mJRi3Xe1MW7COV6ZDaeQw/uu8FMMPR/kHZLqw40gAJm02hhTG
3fWxbQ2mECogTyrREZGguBu3QorR8GVacsxFRY6XGqQov/bP+iBwCQoxZAWQBKTI8SzQbUyyNWTc
mZpoGR6aiWzzk46IrNhCFugIPKVHCa6mMac72RWh1abCjlL57/PsHvyFv1fv/lBrOYLH1i31HvYI
nnWMJKvJXwRQG0Kgyjn4qCgP7ym6Lxt355BWgc2stf80W6Zj24MZ84GFQJ2Q8nj7+F1TCaAPXAB2
LgBoaNv0a7II/KlYqzq51W9uQmPV2ne6K97yhUoutoOCo9msF8+SqpR9MN0YsmP60XXiMyNLjMn4
H2bKmXqgL0g0wnJy3uipPihyvOv7ajnroDJuqIYyVr4qD08yhRefZnbYp3b84aBF688RaIzpye5G
Mh6SgWhHdCJXJ7SaTIYicUrxJZFbcPRqndaL4D8ycLQgFe6eROZd9u7O+O19WGyua+x+S6SB92LZ
/Ht3qPMU3l+hshmIApomq7/v0COTsKM8CDKvushU8/+Zn+MlwAZ20qB2vFjo5uuZDlLJKeZ42Qpd
EsbLxP4ZTk+KhA7qNa8l4h7V9R6ZOAwEJKM5YYLQX24+eYTW63aQfEvv9ilbfVQJAWdmL9ZvDAeX
39TuDqPKOxCpEe5faAhut697yg+7TCY8TdobgdAfNjSoX7xbHX0ErVNZkZ/bdDzO77enzRF0ZGS6
2695v6UDvs6y61gFX1woDlj//BbrIczaT4Mfe7q/AFc+GPhiwLH/q264gFCAP0RyOQq69uXnjQ//
vzcrKcQXpr/MM+M3fM6GjsasjgPa4bzQq8iTvxOX9uzfuliupC6tFlswPMgGQWrYQI/uGLFm32g/
fWVTk7n6UkmtCmbr8NGj88Kt5lA85o1TEqrYyFbknqn2RvgXItMK1vjU2nso3+G5JI2Sm6MfwUTr
DhgEEsUeeN7/HBj59eiaQ092MGrA9QR5yGdpoAU5WKHOv2O6+zwGTOv+AR+jo09tGWPVJkuSjWSP
ZMm65io6ezz4B5DcYyHNm4Vm/0KhC3j7+mnD7toWGPVrbL0ikEm4OGNpIdkccv3tu3BAa+Bk4Vfs
WEsZDsB9InzGkf0J/n9nr63ocnmH7Be986OmPeW3KITM4imrVqJ0yvcF2moJ6PvfE01mtQ6y8T8f
G5RmPel8Tkxcdg7tBeQOekpYR0ItduUExncOUiGaKghrCS9yx9mI2etbuBbgTeK3jw6IlbPfCsCt
Uz1xgdHgMBcPl0Xn6yQVS6LYEcMRfkkQ9ptlOApt0ktmhRlbj92Bh3v6DvzDlez4IrOpJhMwqswF
VPwsHr6gX0747oUBcZG0U4PA6NEqtTawr44CmHo7t9BGbI/DwjyzqtLjVMm+SoT6cA9IhjO/8Y3Z
Pwb07RladeAvwYpEwg7ty3OqW2PYmu/YfwZmeXucnDV64BBuV7vendrCBdPImH0CMAaGXCmjFfWz
Z8HTc6w+2jtjalaqI7sks1TNbFCfku9r7excTDzPPkuDlSjrimBkhVSJF5uwsfp5d4llUz9OLVrH
2NO6KwJxkxZ5ewwk7jt2gS3xj56MwOGWWAW+dG51passk4hi3wGrLUbbcOrFcgoC8DxFlviLK7HA
xIvzeGNwcXr9ozMG6ycMXHzUyI8/XLFn8SGJQAPyGWp9Gxl8E7OvfMK1cBpKFsiWwwqQIAUvWsZ/
yBELUyrkqS93PWOm2nSY1V76MH3GsCC2ekUOgctXgp7oWNbI1hYDkTIrJcr7wLB1QCW/I1axNn2l
dkRTZnWCeNBrNcSqty1bcIQ3zUmVWCfJhhevmLmEuAhFbg0UVgpaVGwT3hK7zuVrL+/FcsodXOqb
NijKcNSjGUJPDeFG3bbiPWuowNNECd8b6um5bPeG++wO0jHhn105oBdNR+C6RX/kBrEcaxMDOKhh
7rwPM8bcb6qNQ/uMqtekCfzwgqXzt19a/TzIOcDTjGx5tCkZr6w9IcD4JL3mp5dHCb1YPWHUOgr3
IP/3ekQXBHEMu2WlzmZDcO5o9Q1xJpZkH9GvBbPay8ycaqAy8x106rJE8gV1Hi6aPj97UQjerSLB
qDW6v4jjX8pVmoZp9DJZo0+S7I7yUVn0M1c7sDbIPx0dCkqECn3ZHMxjpR+20OipdrOuZXE9P94Z
68zpNwc1KcDzJ6q0//n4sw+jdWY3rTuSSO6kErA9h9PI0btLOpxAm5VfV8otVZuPvU4bKG9/mDj/
/eSP9HPDW6OGQXPMo0QZ1ZAczcKJtQ90wozzYvPl/q3NrRx02p+8KoOntW/g5jeZuPln2oRSvtKd
sT6FzTE3ZJ+JxQiuVmi8yyyf6iNZlUVEhV9psXyBsn3afq0b7BBQqcwx+Vkidn4IUipBNPRwSvcy
QJxFHK05U4rTAEtYJbg0ifwyuaWlwhRuUvgk49tXz1xhBkOGpflK0ujSymGvzS6hDuIwprHSIqSc
aR/n8kmBipgztcUqjo7r6aJLsMYMvck4blampKsBOjDH/ZjJmOoOyIqqBQRRBMzoJNhLblQ/EpNH
dlujBIf/Ov0GhM5f2s8zhyJqe3o6cDtBvvHN2MKsM3jYsO/nwJnzywppfYGrzwNDjDcH0CVW/394
WD9Ls3Fd8Xrs8I7pa4TiNLg1gGH42ufy2uF25wS+qKet2HcmEE3+vyvMHFoW8fOQNARcm5Gh28nf
RM1Etu85oPa5/kEX4nvkEAZ45KYuwrJAtpDHWJhBZCSNl2EDJFU1ZpdwV1+kmUE9r1kI7B/I6zz/
Rc2pX9mSUCLJAz0WtOzWAgOFu9208PV/CyrAnSARGqGpKrt6kwC1Uly9XgLCZnk9Lb7XICGYObAH
asjcFAgSH/dFvbbqMBKjbI0TXB7iwe9AgMWsKu+Ap3cq9kf18WCzKDX9ConGme9+cUKLnIPsuGgY
K4yZVBEr6cqnhq/QFNcEeJtV/LWJ0wctQ7+wQophto+znOnDiqY11lpGzuT1lgoyL46mCDqzAoeI
pbqpV2GW7Y3VrZt4WybVNSfy943nHqeIAsiGLZKZgNx6Eg5nKAXYGCnBPT+5uqjfDcYkxbGHcvxR
2EZbR+eO3wx4SqrNp9zfOp96bQNB6ClW0YsaS0A40sdk8ZqSSLHFIqHV2kldmGURy+owIHvUHCfy
SAfaS8gbkzwwbxWUs2WXCPFmzWY3mdcDrvT64JSR3qtBNSOhcTNYXEmnyajlJyJfjO/eNj9hzEoV
MnG67KBN6OaO2arBcHRo/+BoBuRJ5vwIhPhQoocVEscVWN26yYBz4DVekW5W7mP4jkzzbO26ebrU
CJkCEgNVnt7mZZf/mhUtZmnqEicF9we3TPVuw5NFviTtEs+TrNMEc7PkcQ5RH7J6Ir9HowTTEtE0
ChRGnw7YWKPuuWTiPpsZNVTuGyItNCoVKlRiChg5duSPGuXpnK6RuxBYjC4bxOOuUWN54Lles+la
i1ZNl5ZZT454YXazI4yhP83GgVMTE1kFV7snJpqkYsuzMDMPmPtdVYLZ/Mjxm80l4ptuvQi1PtDz
WFvb6Ff4JNGoGt5Exw0xUT9CtcdbZtJOQWQN9dOe+Jytfq3u3Ug8I8ZGh69/TtUUNeubSpu3ElJW
LiC90QfqMDTIyj7bGquY8lsVSAnNm1kCiynguKivRLsTgp6PwGtlTjqVsnqzL0xck5CfSwmRI2A8
DB51/yN2+jd0q869/B71ks6GwZet4+3baougxCVcOBiSnm+kgEsF2+E97vr8NX63+TEY4g0zlrsi
xsDaozZIn3bej8bDIv1Cz7NTqAlO+VjogXlgAzEGoEeOGHyCCt/mzvVZ4hI0rffI3NYQ2Nay4dzB
6w+17SnT2gJNmdS9LLcSVn25MwuoEq1J4T85FC79O5yBYeOsmKY3/7ANGnHdN+PZNTP0SYydlAjM
7723UFVDfe1sOxUmRgxdlNN61wsnUeWOuFEy00uHrhJQoAoJ5DMyzKXWeipactcWxtc2RlVBgfwY
wAO0o7WWYGQCL6scvHGZ7hPD80+1q04KE6+6XKCL38u2MOeHD4FrwN82PxDPfkDCw3fFzhiK8gUV
4yNJKEe1oTR+4El2qPt86d9KpL3A3/7ZBear/55VzFHp6KQl2cbDG+VNsu3R6igKwlkPFurHsSa6
UDGmUMcEaSoqIwe988EFJsxqtLgPWBVoDL24KilNGSuELB17GsNYmtmCk6WnqP3k/bwRDLXBmDYx
+Djbv2cti7cHdKcZBengErA/jt0eWmrEfx+6WjoVUmHtkD3rX7B9ihhT1/31OaOBb5stxL8gMj4y
2/K1XJE/mxvBEWqm0Ry938mk2lP/UTocnGPy5UDkjt+VxUkGfsiOmTlAZhwx1lNlpg481t82hxdH
EH4R4cb517s5RUlpnix7T4VKBZx0YT5FSFiAi+UryYiKxZNrVk1NtDpRmqQwuEdcaHcDY963oUbr
AjEoyN/xQ6yojDx+Fn4NFtpJPoS8HiL+g4VY/Zt1hmNyeCpDNSl8Q/DCUaop984GscxA7zaO+oC9
fgNoJ143zPGASYkBa3eobAm6oMHgc+ceZ0Mp5Qb+R77wciLjpPTamYWd2d6ZzrfnzoMmOk4v3Czu
EQz9fj3A6PEszqYhkCCYMAs1X44l5Z5LFqoVSXgXNec+JGXIbKP47PPgNWwPppJVN8Rb+/B0YH+L
wyfXIWAaqMaSQC/Zqt/JCBIXtd9TUdLyJ/iSSEUVK/LA/lvsZIjCslhv87jUCx+vULIC2AdVDoPr
IJXvQBtU08BQUMmK2p8NcQjq3bzlcD5OEt8xmPCprtGpMbrzWq9ChuPk7Z6r0nCmRNCyIg9O5iPv
Q6Yp4sM2ZXcrDI+KG5rns6Vofe83saT6DJKZl6OXhp2Bge3P8m2F0OmPlPypedYIG7Nqzn+fWgWF
pVTVPIP/Z8F8NjjM8syaFpMkWkksl94o+bLw45aWdOrnX/aBKdNfVtUl7vzIYi1VctRCUnHp+wMm
W40HCsfcao8Pv0Ud2w7v3vOalzReqHwhvEzqrtnDbIzrBRuxR0DrU3nYV4VQ31zFjw+tgXcRSptp
GIoyS9nEURUMkIz6oBa6r0rco5PTmjH5JcxvEfBAFwxhQuRCBT3vgGiY3P6IMtJOGgByk2RIRCQ+
H5AqS5acN/1zrGg4QRPJpV/yAQEjjlQyjkLacmGCeU51CLOgCuA2AfYm12PCzfGIWOTTUhh/7P9Q
mRvXvgL6Zx5HXc3NNIuzAV6P9TsdDTJlZTBg40RUpCvqvsZ6hnulchlcjLY3amKXWbQ89TLlikpb
Hy8hDNpv3gANiM29ZCY4skMhV9hPK5HN9UQgUZ24YDv+AL3oJYeWaAQ9oQ/mqNBcHDNkLbGRZOuq
V4n+MnQFBeCwcKzu5aSSWtGEu5pnYAMJACXymbflSsrPBIyu4IamV4u4JmPBtNTon0w07HJ2IX/Q
i45O7gZSSh/GlxZs3/znhdvi8lDmVxZaPbTineKcUxNebrgB6CG+eI16kMd8O5ihatGyWHGOQcNf
cyatg2paDTMGs66mpqYesArWPpOUUPSM4Y1jnYnh1PREB+cJfjMousVOW8rIsq0s6ibH9COEU4AL
RALafSg7SZ3otebgTiYf6G1PECn8eza59B+K4OIXy1yLf4AiwL0X7ohM91uiG0zooEylpcllSpxJ
YLRtqS2MhmVMC9GJuS2kxaNZMep17Vx6ym6k7qOjp1llwwq87qMMksHyn7RQR4w4/0tViumuXZ7C
GHvx+vo75qSNcqNU5IJNNWrUFKqhGCxxfaSC54MeoPkFyomwbEzEYwnw1j8oggm063r6QiS0Cro9
cbyjmFAB/VFG0w6vwpCmKAACcUu0Pku6Gy9Ep47Dh1/c1x25YX+2NPbMzMuEKPoNUatOQEr8LZHW
EW3C+Qd5AilTEwQavFVzKdzLx1GunO4bGiFrHfpbYSytGTSNZHDvSkrBC1Q0PC+GBvMgdQiiGXj/
ZCM1/QEkpoKmNDvYbV5MHNtzRN4BxbQmYw6HIB9nplUYZwY+D+P3Tt7Rh6+Cu84Vng7gG550gm6Z
vppFdaQgcKBTT60SBydKK5or4LW671PHhFjV2HiDLbGUXFoJydQkmzbvoyWbjqtu18PQNdGj4etE
sEaT5ul5lgWMvz66BCMN6ikU4Z30/KK2hmzcNG0Z68Z4F5tkMzH9aOVqi0xBM986ZG9mfz/f91ev
ReYXfFF3/KYwDPNgRcDnl0CO9zQ6LlCdvoUD/1OyGl8Xg0XXOvXDqJIUccG0NVaoEr7TfgZmhU50
iL8yPr2qEm6prW47YLXjMGKLfnBNKNjDOyb7FHaaSXqQ2lPjxUwYtw6UPYWvGVBugZrRYnhwoU9A
rvwciflvwIdZRYslRuY0Y1wiH2z69YWPJPnQKgswWC0jvGWRjMKvNzS3YFjoMTa22lUJje5Pcj0H
nPg6KdK0b1skpUaVVDq4nR8yQJC6XiSiGNxdpg76tUoP7NYCvBzaltCvNGQK6OBESVWU9dxzggr1
jKZzZTBZAzAO0U6ePKvMLi9aXZ3A6v8iZNBD0NbUPohmYTGAQP5+oOF7mOcbD0Q+0O9EHiNa5uI8
F3W1K+4uDTKoXDvhzFAZ68E6jPbFyenIGyAgHiOb3oF/8R5E5BPygdPcSA+82JczYutH8xdTE56S
dP+hw+J5gSd7VdcFVi+o9lkn3WW0VcPPXzc+e5Og0hlh0HZs/thuXcDmF4GQJakvEJdRcK0L38/A
aKHGbBnEVbd9HAsKdeEujpHtOQuJO9qTcxKKb8CF6lVZw74AKeQavZemCxETxSJtUREL3gBY7Ij8
4VqkiMOiRQG5pg+fVhd81bIClZLgm+sp/0ngzrW1rSi2KRd6R8kECTjOGZjioEDFWL5w6KgDwx0D
DX5rE0yjS4hfQ+D2AHHFkcE/4LQZb2LD6Ofo9gADyqmePvoDfrTVOLDwaVX1NovDG5Xd4ZG2jg2W
WMtHgTK8r1lBI/LeIlY0iHtTLUydAM9b7lwtueGZ+37th9NeuSbS9yn85UTPmnhrcS7kXW+hAZxh
HhIhqH6+v34DRdMFESq7rrznuLhYXwRq8GLjKYMy3vba+vrUpXnuJsiyMm2SuDIJmfg9ClCdHg3J
5BtDoB0tM7deDyquEbwuEsWNxoLyPx7wLEXtcGPSckrMVxbwIzquWWkJ7bruAISyFhQ6J3jH+9oU
hjSInUoj+znm79Sv8SO6XLo14UQPNnajIj6bUKQeACE1YVh5oy21cqz6X359xsSDHVOc7F6MuY93
nGLZXm30rZdY6hF0EYAR1dEXXKfnfoWFFGTl5heNKkWi2ErMLiVfhGXuRVIUa986HogTivsfm4hL
7h5G9GYrKsaDa7/0utllc8zDhBVdcSyDPhYgPJ8/PjlfI2XRTptE7o4bgUMnFpyMv/mPmIcpxgvo
XiUD+6lMOy6LzpagGFsYnFr97BwJnvFRypJPQGNN4GDMtQdw1ChK3/DyU21/3k8kJSpkF4EBFQkL
/DSYJKczaE278wsT2DvjoAFCXh8BBD+W5SH3D2QF2w3yudEv+MfaIuJEnc120sppb4g5k5sFf/wZ
dRJZYPEk5ndujP05cb8faNX5jCBkWez7xLqYiEuVHT26qn1xjtlMm40Ka6FcsqwHakbc5I/arnoL
ZFsojp4TPQ2sN2FFbCd5VJqdBCXy6OranJ7rtqB2MeeIguXw5qL5qJOni5qLhdW2xD3hLeNR8np4
sF3a/OZS1WWNtLQwJTolelS8jvyAuR/LLscuC32tCIQzTZoMRSITqfDfScV6OGvZHqq5uK/IjZ00
dvDTMhc065rvhlEwQ51NnAK/C84ly1mmFBXvMm5V98lZ0lhkfCcorG7F42ou15xFIw/HxxBdlFfX
00EpTVtiVJQ96NPDZJVV5V+agCtEr5BhPhlMKTGn5q9xV7iWf0GSey0cnFT/iN17goHtwwtBsImM
CAWN4EukS1g3TR8/wF+5ZdG1sqTA6otDA6hZpXto4M8s+smdtTWuKtSsVnhCkdnhNhTGFXMi6EpQ
cukEUrFKnz8VpYt5QMu5KgYYbLXOlnlfYsjLl+z6Q0ezDrACUqOrJfQoKKRDtbX0RmKon6jPgZPA
MytSoO/xIsn0ZqNvtUAh+IDyN8GQMSg628lSS7mYqqfT1RHD2GBOObgd/9gyIy9zpZHbg993X0Dq
5kukMJ0XeZ/g6V3VGA1AUC2hdQePkMxrJUwNA+z5WObYJFBR2yjzmWyKA7IuiLN96vNQ3GOU8Gcj
q5WIJnwwkKwjx9+pWg+kOJ0Rtr2x/avMIralCsMpzKjp8QQcMZFo1849UBBkCChCb8+w67w8jJC3
dkFjlBBhI+Hn5yj2vZTbLTgruJ6TQqk30B1v2u4WLcquGf0GsyumbSVjk+4jTGfYre+81x7pZLRR
XshGs1brp7dZwupeIfsEGCmJYx7bZK/ZzVqzgM7YpajMORdKCufkm0v9KMYxStxpDCFPFDnRE1AU
mqZ2u9lc87XAzK9wkQt/JfC8Y2SjTmZVQ3Z7lMMxUSZMt8V3scIBu5GjkeZ+eeVRlY6c3FuEnKJa
+ERz5uQyAmmAv4VAd0cywfqGRxr9CULPALwTaTeYItpjmOH14xiImBFvg5mVgQKB2k3acDCTrxln
JKK7BFVWWJeyBPhmEYHUQVkyj5t1fMKAIkHa8Z0cOIQOpwBWlWeCTdUXP4zo/X1Pk4ynAOhsPwBr
+JYeUdAvu6jkaQTTpKE/imjYC5a/pHZSNJlnAKG4h++dfpWDFAHcnmVqyBCKifpFFPU5097nIS4U
jRt1rQC/SonRJF47oCXooecLw7Ow4enbx+LqCg/JaiIh5fOm9wM+OB2fkaNDZC0ORADRcFfY9BRq
hjfvw/Pi+1TjBaUh79IGy88+2Twl+GRsCHZMTmCa3uRKKvDM2vX6JIF2hJP+jNOLwu8woUaHvr4m
3RN5pbHQfKntr3QywvWaJFIMErMQO/QaqJt1WFWaEby+VYyAbaH+TUB89N6WKVCIDz/PwO9bFYU2
47QvSRVxBDjVOfhvcgizBWhG/IkY1u1ZZVUj5MSaOhUfHyAG1G+FUO/xQBsZcQEJtWFHi9N6tVq2
/krAQuKpgbClzEz6fti2matAWvHPMnXWeNy61JUq4H9oBuJmRDi7JqGppCsH4ZiC8YO4iZq84wnP
U3Szn8zdrB6a4WRSi3sQvjqr86z8nBqNjCW/groXDhyywOrKx1d1rrRnr0VxjDGDf9113jSBYb30
zgCYJklkXY8Qc274mL/52FclrVMLlKINWwZeBvZQhI92UwOo7MVa+roemvHHpHLUxghy9BxWW6cu
Or7jkwLwV11pGIbT1H5A8mIAxtNlOtzpjDu3Gb5NNEGu4G/F0X1ddrRRWx90Gk+ZeITpwIVk+Qx4
zRT3BXD3roCpfK/kphjPgad7GX8RrLqoYcABBM7m8f7nQg++TkoRRhiicNdxVaxCy0g3VG0QrYLe
zCWfbxs9Wtq+pTZVXVijRiMT8ktKdLq0gMHTYOxR+i0uvOSJ60UdL37n3TMvx2DpXimX91FfTYmc
3bgLOGwqDkUmSjfDADerwlZj2xBf/8pquiIcFix2i1OBSsSshaNzJRFjsrUtcV3yEjaAfJKoFXtK
24IDKiXCkaOIAfA9pcQFscjLMjR7qURiYf5dEBiubvJc/Kgbd0rWPh6yK2s/NPLyftCZteqkDjwf
ROmZScL4/4gzuAc9SH/QjkNmxtv3vXF6bZ3+gq7iNIXI71yJAXdHjM0e+ySeRZeZgN116Qof1j4j
2rNuwuH5G045gGRLE+Q/MNk5iAWvZgcGyWQVOqOUQ+77VtJH5QiCUPLX5Q3Njsqvda4DzOeLpX8y
GGFnvYf2iukbbMUudEtuWFzhd1arHmCkktpougatG1FK8IMwyyvdiI6WtrpWfowQsXKt8dxbktAn
P+p3ij9dUxtwxF7+OIEqWF6G6Es+ja1Ce7db3CQ88OwxgQ1PAKt+3rFHfFrSRj+MLLY3R/anSD/C
AlVpMHgEIwYeuWXylOHBAxrQfI0PFg3ieCWnlJdnv6JBrrIUoDX4QmjEyfMz+Kci2eSc32FgHjHo
17SInI19DLJLjtRE6srXNjFx+aqFLxVjBa0sCakpCDxl1tGWL3ZJTiPieMQlCQMTijXy8TlV6YAX
ZlVaVZzsO/uptxDHBCsIJZ7GT6AbBU6nKlw2jO9ft2xPGV7TjFlWmM0IZek5UACGN0r54jDukSzo
10U0mQoZo+yntOIUBvd5Z+lDaf0FW6+/CztE+UkOqbQJm2QUlzLHCkx9TgHFpAOrwPYAkFuMUoQV
dBmMFEtzNH0DyYPUI9m1tiTtqDawPtqCqCuBirUyO6F4fk6ETtii8/sEQgdrIydVRwRuFkgfcPW/
XErrBMiTyCUBleYmxF+z796sFzbXV4WuhU5tUhGjMsXMln+Ickpc1ZIvb08xfN6OMvZ6t/G5tOo2
G/zqxfDTLDBVwvQi4j1mBVNofy1Q+lZ5I7oaTL7SXK3aC39Qftp+AqE/9CUOQnjUXpVDoMduSAN4
vjDkYgAqxksKAuoDLJsczYIiSoZhnvyEthNdRqbzN+lO/HZeGC71ohnauT4iOvO1tbzOsXO7QeYg
2ZyrEUj78Gs8Y9EaMmAJ+vNnAnaDiGh55+7WNKejRi3h1xpwUwaPd5/QJGsbMDg7iXQ5FgKbWXjB
Did0FvDC8Me3RW9zaVd/KgKPJaljXTaaooJNNug1iNH/rUsUSdFIe3VCRhfe1vONaKI/FdiCLQ77
4AL/RIqnAD/6mNS6ZUq2YlFNKMC9qGqZUPxbmQY5NlD0tFJTXce2IxTwZpCUqWQ+9N2mC3oCNK4Z
owIUyvhrUkEUv2DWhfH0cqt04F2mG4AsmXto57ZonwEq9PJisj+4ORr3W3L0WjZwgu8hR3KQGoqb
BIrDueyJUFY23te1oEl7mUYkoB00se+nnM5wuNm7fZu2eDUAxOB2SiUgGErTzHbhF2LFldzqhFPm
eStxiplr6l2cn09NlAmJeus9r06DuMc4GH9XKeQUZv+5IUGn+ROfzgr2qKwiwihJNwfkUYc86MkC
JylBZOgvS/5i7sMEYDlksS0rtmG2Qz3BCqumWUd70Ewu9AZ1xIWzjRUK//amlhpOwXXn6D9m73Zw
NiWzYauztRMH7+FHvjT+tJITW65KXnpzdEF4j7hpkYSt7PAxBh7LaeMY3+TNwXQ5PwbItFqjJC6f
ycBLLloKSzlRA5dV0LHp5f2vembXuO2cyNwc62A9eOvpj7srYLwJS0s7ahsCm9eNiAM4tSueP3jp
kUbi3hnZ1t6pxmfHqAKHLiZGsWlRgaAZPFOYebjo5NMB8R8O5lF3VqW9PI5e4V1XnZhzvDP2Hgmf
VfIW5+v2M8uXyfZ0XYAl7jPxWLLUA1JNMkD6wbYPDVH1U5nA6igdgm1KILfoVikfham/GKJhexgz
r3Z4htZ5iHYdoS0Ve6V8VEuAOQhLC167uSpoOO8pIe9pi5Yr/lkc68snQB3dtKQ5ZmCs0EhVKBVK
3kNaaHfr9sWpFMtSTDMWzHElSBtjGtpC4ru36iktFWsTzJfLRYLaC3zg9Q9BKRdVwrmdKaGoVcGb
NAGPLHPmW4dt8Xp3obJWl+a6hV09jXwtcBlmO90rrm1j00cJDdOQCE1Zj9qOuQQRLBjDcHdVwlk9
dlo2rNBciKR6afyvHdRIGfldN+qwFozJSzJnbcYSPK3haIcfTrGwehyCPjHDUNFbroZ0j2VV8vEV
rCpCpmq45eVgXbeVjoArh+MGGUqLnemmZ6ZO5EwDNBI5fjIWfEO7FHuj0n8Q/6EzL9u1Dy/lvlSD
Dl7Swgf87cvwYc4iX4Z24J0wGAkMLFQl+gGBVe4RjsDle0Q5e2whJAjCQ2474QCu4K17mRGFz+Jk
j+Y8jqisKVzm3bMO+nLACMVxMN5Pm1Yr6whIvI9ujlUKznArKUrnGytxb826Q/aHS/PYmg5y9UoQ
jDElOjNulRv17Ub7A/H5A0mueTKTp1RRaBa2MjqikQCp/I0av4uJr4Ujz0hBCPU0JOp6DzEut4n6
9jXUM04cVYtv7mqHEZ6ALXcd2IeQlWHNxlcHbacie6Vk+JyXFIFiVIXpw/ysXaqHZCf5n5uJzqeU
JbCJckrklTqDNSv15eLV2HBzV/j2MVjYp9Twr5lWen/ZgUVBwwP6NICYHpVyIY52z8FEjHsEVvJw
hbYTDCJqX8vJAlsRFW4NjOlpFXLNP3KeAUSzzCrqmUv0wHAvrUBXXrrgoxVlpXMnRxhohrha8soJ
j0e8tkbjTasq136tDdCbab4DStXy/hCTGibjNTkmDLdts3HL6Wapa9KkKuYrGMK3vAK/uwq0x5d/
sJWKNXY9LIvUgDvEYKdTOMgBed2YvTZOCiOnTQSvZx33l2nM6QuJOI80aQMcvkoAsucU1QycEw2P
TprZSxewD+aXkkIUH9zqfsd/Ku0mEZEDjUxwkldbXz2sJrq1Ev3pJpHJP47y014OhsvOtClO7Xnp
7QN6FO29mEUXi48atI2uxfaHzx59dNzWWm6YiCaVECbz4pzRuKAMnhgD9sU8NvJRMFUTfcRX4JbC
MzUCBVDPvkhLfL3IjO1RhRhJtgiSdYC9/yUuMqCdKIGncy/OA0wXL8F8XJyWrZ3xupJlSTR5F40i
wHtUEDBFAOAZby//64f9Zmim2N0eIX0OjYtz+jXUaolauvkSD4Ixb2XMI1k22mD6gW1WyX2b+fRc
CdjX401H49MfimLEWUndCPQLTx1aZQoRHFuYCu9pFSoLOgN+OrYzYo2ANN7JuEfCqnVUwix8/olS
/k4Ixi4rm1uFPX7HY7wGV0jGNyLbTA4cCP5dCozi1gzh88dVGKRumQE00v4TG4Q3rOBe4sxIHR5D
z+caddL6NmsNmphpMYyvd2a+9r/BLfm/Y/tPCJ/lkoXsL0xkith7gY/thpvpBm/uwiS5THT97KiJ
MtDrZ9ivEwWXVMwD1RbE2lgNGd8fNDkTQDOCWPiMd12zvQ2GoaAPgdh0tlq0sEhHIHv5jEf4NKCs
+DNzC0JgOUF0xHghvyDeYSctC6EcKwm51rjsbCCRWSrWgLZTtFoaIIVhiYXSpiOonOImaQVlS60R
sarJYTVjpAepIl0YQeJE+ix4ZUa2MgQRFn8aHyCyu3GQEYEBODsSUkhlzgWuir/DJ/pER4vDsrYs
5f6a7PPN52ugUNGagK5iMp06DoKX7EPMBMhNQrmngjXiOZJFO7Cq4gUoqmpjyMtzagwcgkJZXI6U
9opLZzYeJdFkEBN+tulnSLxjt8Nhw5oBWLFPDNYCnHwTVJC9WyaMJpvcx8zWUCvzKRN049PFOVEF
FuVZBMZ8uuKwKdMY47lp5rseNqr33XqOhlQJx52fbcVgu7S6Iu60UyfNrkHrohAgnxEpHQBkjCv2
uMIo5vjtjp2gIkF809D2MYfcN71TpyqS2mefaPo1/ZBb7W//13Zcc/Pveux5U9SpGCpnfo9J1FKB
0AG7UM/Zq8bI2ykf4oMathS1mV41TuYSvHABww6QD+4C7fAYpeBvmg0FWzZVoCr6MwxXRu/OCKQZ
lu1enFw4sqSgcaWGvJsuSoSOQfLH/dfQQp/zCw2UE4UNhQDdxPzExzzJHfyqgEehFUXDZkqq7nhi
z2NdGSoJh68NXPdw8sKJVwLeWoZDGLYKFz+sfv8uf6MgY75rVdRQHmhBFNnC7uIVeMLs8V1CND6W
iB6hrp9LlIHuohp7//Wz43oxBvvdO65Xo8izJmgs052eN78ize0TE05qpDsDjHQL7+UqfpyXnbdw
3v9N0qZhJE5LkfYLTvNdn5HUz3xD4j2PaCk3+CIt1nPWJRh8+7ixRx4+wJbtzHdidMx9kusxYHN9
CAbVlJ2/8YKOjSrpjkVbgrGQeLqzpmnWAlES8tEFLIwnVFed6ACfSD+Vmqb7bTJL1JAriKRXgMGd
PqnwIZrnub1a+zmpjHYKkdW8YJLVKFQ2u3elD6kFA0sz1uRyKpEPQhSYv1O6x3VEsSNapKpt9BF5
CDZBTyNJjZSpKv9kyUR5K6j2V0TJ1jhZzqwUZ6xRjjeE0zXKT+7mN4+iNZtUAGiijGCjdOZu4sA0
2spS5MBMt2hWcmyFT+QOC0WtFwx2qEgimVDqs9Us6+LX/vf56wYnlcJgfnBCUBpQX7/h8IystEYD
5vgGFqANI6wGpPH2Z7sORpzQss8gjiZVKKOuGlQUAzIQtv377xe5pjLBFz+go8WmY40GXxZU8kYE
K6aJyi4qDivVPzHvR/dC3dfaWn8sQgp57YJmKOgPGIrs61+TkGRg1yVCCi4/tT1ub0zb6sF/1Dry
tXKIMqx4wlHc1mOzvY2jpZmTaH98P8VFZQSiMg5Up5bVh9fvqlbWic2lTOxmF7F1Djlw3LwzLUZc
Yj3opTUXqb+dC5BJodb6AWZeAAfRf+UKfkLphYqqjkfnL9Kt0+5dCjfbxcIL/ET6SnvOJdrkA4zX
1tr5G4N4inC80YkvzspxEHsqRp2C/nTyWMvM1yqaXaUeOKhG4rTa7mwASe5i6zuaExXfBSxtvtnc
0v/9hz0f48GHOodN2u3/zeiCtDat21pteq73ihjnkC2hMgpebbETVtgFgQLjYIZYrpWwKh1koZUC
ZKiQYa+p8i4U2gVmELRfsjY7s+0mfcEBcMBAtvQi+Ii30nH6N29iYOXGVbgC/0SwT6gyr192KH8J
UaOdWTAq10vejUMBASwJh0Yb4qaDHUqqAW2HVciadan8zA0xHaXKrg7PXQccnwuF0awJQO5IHL8K
ylJ+vZUvd3uSp/YjBid3zxm34T1F7BsY8H7Ao3ZMVgqc9txl6hBpZi4upbnY0dm0Rktd98FFRGb1
zHLz+rBZgvTY5+pMKP+/GxrtOjQ75gvWbCXZBg5+9y2G9RUVb6N5CCBJd4WWZF0s0Uv9T06HJQVd
a8AYIyBP8ewe/pi0RJVG3GdMDGoD+8cKc6YJ22cqiKtVoV8U40pxSNcX6qSWk+v4ro4jY01b/hJf
6PCF+cVmBineP0GRrQ+3gcbSymN+iul2E6Yt5M05I4yNLB1V7MPsvPPdjny+OTswQc+WNTZfNKev
dPy+Fre0LxVpq/+jTpQiiTWI48UdIheOk3bTGWY981apEfDVr3lzfEEdV5I2ZVEaapYusQnwapnc
NasbUq1p5OyFaqx259GPaNhOMB0embqfT20bBFIP6u4nxAMWFgLf01dv1UMz7ckip0OVZFObKAkW
+b1f5qhXR5mzZqZzi7YmLYqiF3xkrmKtmd7PLWyLQZVSKcQ5UwQRl5fwKgsr1xHsPgdicNRFOn0M
QhcHVB+zP2JvrVte+3DH9zeGgIV3gguaCHXcD77WUwqeXOZ+CyBD66hi29fmpD1z7lYU2pE+lFWq
ZqpBefSuHYxLCuBiYwDOPmC/q05JbbwK2fuH7Tfv7svU2WROjg6+hf+Amtl9PBEB10Jd62Ywmc2K
/uE8HOzQSIMcVZnNIidOzrKr/7wx921kBckJaTv/kf5V5wmnM3BmdjDxg288AXcZVzBk/L+b0hLU
nZeQa1a5n7abRbnFAMR8BcQ/filffem4W/0SlLitPZvA2sg+WFp0Mvkgn12hPgQE4w/dqGLKYbOm
L2q/Gat092XDo1ZdAYw3MJJeSuUZJGeCFGHTNcWleLhyaBkp3FfgeU8FdVUV4gggC/yseCPNCzn+
Ut4Tv94M4x/OY+Es2oAIOMYJ+IjCJfb2qDfjTKlKukO1f1K6C/NbxwG0muoOKTJ3hqTM8+37eSPv
nR6NJ7J73DvFBTOxN6Jbj16AwdqhKJOY5aGYe2Jtadqss6SAuinsh5pFF6zT7A1MKojvsD8x140E
4wLoC5YzQSbk/ivqulURLpAOWbuliPWwbW3QwZMS3w1AKD0iGokZDlZYpJCIjeLbgk5oASnA7BWe
BVk84JFE6xj0QaD5W1EcI8cUaghWbPZxpc6ECzT8AsehUxumencl6emxFqUCE1XTqVuilHmCA/+n
sd2mGsQrgfdDEYJms7Ibfw3rYVKQNWdZ+i0Mi+4W05PSF1CuG+xaRhnbjimcqOk4SvEfKG3iYfvO
JblRD3Sk/S/MymJeCeGARGScMg4VVUn1L/uUpoeqsHlv3L0ddxCrHEiq+kXOhHM/GJST1YqnXtKv
kJl7QwugfMW/DbLzVXs8RsE3UYTr/k1GfzpnoMugYFK+d7b2QmNhQ5YomZ9xdm965mqHrb0beiKZ
fGzShKwvm4+iF6gzMY0wCr9RaD/kzjwhJsG4+jmUW49p+Pe9LD1YLAYiV9+NvsmPNFc1APlruGh1
KX5wdRxbT+wWKCUatO60HqEClVVS5orZnagEs/3wzK29KxuuZ2JiQpYYpLioOcA0GBbdH0gKtiag
iKXaQHkytsGRa/YugLJHUqtFUlUKUIeZWC7Mp4qNFuNav9AzGUcShEivG/VqXUtn14k6wNYJdx8v
+sWZA6M/0H/nIFq920GCHGsAXFYaO4W3azOGJc3uVBETJLtgeWqFvurCQogDwsMPQTEZBTPGSsu+
/k22WOH4eqF4KvTH8DYgA96qJNWO77zyx0O8kHLhvTMYnRKDeT3ZSnM4B71MBhdEBb7+vNof/Q79
Kh24YuFFC4oeKc4Kmy9JSFkOTnvBc/Cv6bLaceZP2Kl/k6HDQalR3E853zYZNPnc1Oq3QF/YEjw2
llk+Lcneke8O+cMT+25INioPeJ5ynkdHXWDLwuzCtjUTNoKkBeQyrjbo1nOVRKZS9dBYW+mRnPgX
hSVCFSjgE6cUyT8RS38d1JhzeMS0p/VoBtXRnjkKz3AUZoguhNWXIvUWN17NQvgz/eWEWvpBrP5/
mMG8Kaa/h8p2THpMVctd+HfM7c5Gva6uvbCPjudVySdwAqxeONrYx+Nz6FOCgVkew603i8mgcfmf
lKQl3yz9Cdn1ysMSvEYseJIv3g3ZqQKjRvZM7GTjDFmApuRU2OBDktWb8Na/vTTWJy632T2LH2fZ
skhQygJgPpZnO+ihe+RO78e+Z7eiCLP6ItM3bL2BOHIAMGMP24r3ccTiDSEA7ilWQv7/ktHji9nr
3QzjAIcXLuVOY9J0qspaQMVRDAKzqDPGkzoKV7jCR7zuus3CA8HzQkg/q+r6pBPCZ1J8L/SKNpGj
SeRd1whlVc0yguIkK7nIsrn0NuOVuEClcSm//dKn8XTNbrlFR6jD/RhA4cT89lf7lcibKijN2XdV
bfJg8dIglMlxhkWasBOgXawK2huA718eub3UEzkUvBB3jPGN2ptOh8PYm6gtI7Iopy8x9U3LrcyR
TKoDmWZkfxxe+Kmt1hDSdjLpZYx/pkrCU2p3q/w2YRWIeQjTRV9cu/TTWWa1AJy1TsDNd0YwvK6d
yNplUkz4ZXvNdg7j7dQoCLyNOgWLtTZ68p7n6b+902YjGwtYChtAVCT03PuYb/MeIpUaX8qjH467
zO3feue2sKhFF6qHRYgznet1PqVQIVSWb7FKigUHc9bDgaCr955b4wRR1cblvGDksNU489Dl9S28
CAN5SmMAhYDkRHAi7h4sJANUHKOvvW8Mkozt+4aZ3VvSDsvRjaP7/lA7uw06RJJSm4h30XxNH4z2
RcHYBwQ6LRAppbJNN+TMKuvFP2WbhR+ITobRazRHsuBBRl40gGdkq476YgpYeOLZek/nVoZiB7Pe
mcffXr9XAkuo27J1N82QNDHsenzw5AoFDyO4exD9IloIg+XBq0/cvrENhcD3ECmVUhMKdarVvcRe
jYAhm/SdneYgZDR+Sw6VaqzubjOTk3M+Eq+B/u4Z/AWuDPGz3uMTWIicPYfOfPyZL131TcyiEzgM
yA4hfc/tzlrGOKe37rQIziJtwWz5tmH9yyKq4DH9Mz6PbNG6FOAmvq8Ewgl7QxD/8rWKPrfHRkfP
uaJCW54spwHP81O3EbIzGDucInvhTpErRLf2qQiLJLAE+ZvAUSwcjhMDzBO4EdPfXj5rGZaKry7F
hYlcPHpdYisy1eX54U9zCNf9xk3/2WmW5+aGNugmjH+74S9TCfJ+11LeL6tKbPgexwmQKVLu9Ahf
oxUUn/2p+Uueo3YjVbJyVDP4GTyih13X8LaLOrFDAJ8E6tQq8xaHTM1OK+3+dtA/lUgp2X5TjxUx
FLrYjGaux5W7baiWltlKjEE8xbi/5soUY1f2Q3CFihFC/spJ8+c8dUH6qVoAbdTpTpkpcUc8lTCE
Tv1EAYbvpsmq0unzwGpCv7tqOK3TDx2BiVI177gBWzzcBdhdqBNVdKodaY8zkGiG5MvRTiXtqZFF
IkaNF1DY3DPmq6dgvLgLOffU/f9o1ThzJOQH5kv+ieBSxT+cGOu/D8Uk3t4WzcudgDUH6vu1sPK5
t0+5n3u3O5jozf9bsQO2FYj3Zb/3rm8C1zML4Y7Y51KxK5xxwawbWxfnPC7FAywZxp2hoIRyVcWV
XZIJ+IdoBjfrSOew5bmzU8lpo6X6FB5/kywsEu07Om3054KUTqiOUzyGXwBCRw7Om6RGpqgkdR7A
k92BXAlTrUB2rLpLwDVB576r90O6mndV7HF1t4TkDmrYE/jrrJperFBifTi7/0OzMDDDZ3t3F+f8
6eutrMLOBqL6wQOOTml87glxmkog6sMTVyzVDMXw5GIVEouhfKh8yVltEkt/ww5TA+KN7ibXLeSL
Hyk3f2ty7mxoLbwLprn+FuVNhessRr9VosLo2DlP4+STr8wUeDzSot+uASiB5GBaY0tcLMGb83oW
A1emPl23M/D8+1x8brLAWMIgBcBqze6aVT+CjFf/OGCYIBRWsXWWqSANwK/HTBgFgdOZSenobpeJ
z2Skwx+arLVo0BxCragxbP/RqemAD8NKWugkU1w4H+g/CKAgSM32zvcQOQmscbbnaC2xzzJLWJlx
WPLul0SnlKZwRfI1doYv5vQVjUv6BZ6OoPPde1XYOYPjH5/hqjdDuyoYGQXqOKqaWWW7Z53nAUtk
I2M0lZRgC8eE4VtwWHNtl1th9PdaoG6BPRNpu8Xeen4hZS7IzIaJXr3+PEFb92KrUr4aTjcVVNr2
NPp39cIlnzPblvSNglx6XWORvkRxfEPZ8kWRUHO3ASs4pqTh+Mn+tDcoI1i2tNPpafTSojy4FmAp
5lvYaa7JzFmzmeyaespREbDauflQ5+LvlVGkV0KYlUYpLdX+L3Ciz6qkxwx+nArjIFRLlOg/16x6
c+OWZnsPiIR1sfb6UD0+CARHRrF48Rh0hhVrxAeTejm+Q62cAe+7or2XKmLEVpKX/dRis8Ro+0Xa
o7Gq6BzFulk5JhN7xqays1TbVxIn3DLaRgNzL4/zf+ux57OYBvrQbUN8wu+7kMMS5qSFje/7FYCb
3Za91d9w9BKpCdj99cZCrcfAg6Pj/c7hmjfhNCBUtuOUTGPnO3sNTmf+89lU3t8T20Jg+vCxBzSL
ENShmUJ+qumdD+YQsV5iWsASL4CcMsvSoQB+IsluxlwsyXM4uvRXILkMVzaJ/E9MTxBFYa60TtH4
luo1lX1w/BzfTwq3wQg+7mzr0V1PHVXT6BZ3MWdUijAGg7j36gTCZhPUb9t6u1hOsXHm9oTvvpLy
mGL6mXiFFe+hSC9UY1QIahojG/YlA5S7Yan8kruLqjPQPMJ16PtDsTIOkPtddGJiL1TAtofqAGcy
OFo0qHhf80awli4kj1cOmWcfnvFUGCuMYTrCTlQAKxqUJpmj3Imk5Ms3mMhQQV+7GkUXdhAmUbvH
79eShuOYJsByMf6GgX8XRT7KkB/+pWYVYyBdnFtin9afXGVzVJAP28QoM23QYQLRltAoFKerclv8
3CGZikadIl8+vCDiA1n3VPrchzpSGNAACqHrAK+t84GvaL05u5XKb1V3afhnBpO0vmUNYTiDG7b5
1sJrHK7QMwku70VbAk/AeXCDQJcDEV4RZC1BUzLlWcCzzp4EA4twOBS3mt5W6PmzXfq2fkpX75Zc
WBZQSYqYKOukHgQBLy0P0E8sPFbvOPo3cUloP+wrbs6G07HUIT8aPZ+BpX3eYgSDngonZ132WTbU
mlHNusDOKGw//BcUW0vGDoVt9hfiu/988QLE6voo6D+PKU2Qbrk6zXKkofhOH9oEgNC8qjOax1XX
yrWrtLBjDNEDtKAcehGyWegyNuepEcnI/H34CWplpdQp5XBFoHHci/NQJYXwoSGsWyD3+air159w
oPnxzoJP1Fwhd3tYRtzSyfY+s1LQ2chWzKzjXNgT99vB7B3YiOIpSvAujlVCunYAbD77slmEgiMb
bBvGENMIS1YkJ6WRF7886iZyLcDSVT+hkbpxT1EKQgi4KfUr6irvE7yXw4CkzfzJ0inhASgsHLHi
XlrPemOK6YAJ+sLgI+D1F0y26x0MlikL9Wa9+KAOafGRmqQlBdY7iDJR+enFefUK2XDFmEeOPPkH
GdVSCjpB2F5rc9PuqV7Fi54M8EjN34/6dDy/iNOVqhGkksej/0FQt641nozKge2Kgh84pxBvXKRl
7OesoDpo/3V06a+rwVrsSZ1929VXqjP508k6QZoTykKIOdxGT9EKSush2RJv5pBGWInEXGt2eQkl
NywrpcoNAGLt7J4jIiMxXpeRy811DduPH29wK3R3D2hChKag3HwuJb6aTXPpqe33r8csYXhdfjJV
Ot0Deth41xbAUes7OjwhtTltlUK7zibOUzo1ZL0SXGcKycMUN3xq5X65xpqxbfJL/GnVvQA4VWYj
Wz6y6kVfimmniiVtjX9ZNU+lFPSOlJhfw5aBso6ComNCtzZBKfkvsvSWvZE1+3kIqT9h7l1HiFm3
SdWidm0fTUecc5gbMLwQuuhOMosxsgMBYV/JG8FtjrPlym1SLjuJTzm9BPz40Xcs5sTYGR4XIBeg
dxYtcZ3z3eQ77+UypH/WMbmD1W6VlJFIw5JvkQaOVIDGa0Mn+qEMNDLVnJ9g+UzY4mroPDSJzQ8c
3j/R5QhBL627vhtYk2IRD7HkAzoNHFomMf3TgS7ICbILBvnalBKT/De6QZdCOVLo0g/xtD2dMJUz
wRdWCtNaRyllWQFZKWu+4lRP72MsUO07whn2h9aq6bdUXgQb6mdRXbKFv0P34b1nP6KQFB1DKtHs
wLHnGzZb7brL5x9I9dSHrE9jABFaZE6hQnI7/ZG7df2LWcm86lUCP3D7Spok6kMsprYxVgWH/JnR
sjlPu12B97syqcYK3GP1TJjUAa3T+Di8qAgVTyhV498DPTrm9p8tJIMTL1kYBg+PHw3pF/YjxGEc
jzh5o9PRg1Nwj8x45GGA2CSoK2Je6+V3sZJjlAmMRAmE0CuuPlbM6Yjjzx+TNg5kgEJhYB7f4BXt
YSgmbLvmziXZ8lwr5GClBMqeS3l+0VLmWrD4GwOgX0PPlc/XKUP9XUaeHcw9bMMZMNSJrxEP16J8
ceuOvgHdXKCb/FLca8I/Bk3Qk2M9/T4kwKEmgW4A/QYTNuK1iFUSglSzky8FfYdKROuezhmT1Yzi
7tqLeCyuJg39PSkFXl3RfCZDCOCnVlplwxFlUv8K4EU/m83D+CqhlgX1HBQ5raDgbPaFIcm+0OOy
yMX2i5C9Ia2IErSVqgTe2mtPnPSP5HhNZAiEdHkbRyVts5ZcdHS1SIqtOb6kqIPVSd60tgAyjf1j
wojvgSy2t+rTDfCwnDpLnrRmQsW+KO83E8h2jOO4MM0xSe6rPsibJesI+eBYLv1Mjbnt0C5v52fN
nlohUVnydfglVRqIHyFn5aZ6n1yJn3S6imPpVx7Que+LBhiEbrg+ReGdKXIcuDg9AH5O4MAKrXmi
09JWwGjlwC8dq1v0y7QH1Q9NMFi/0zLYcJKpgKzGmVX88Zhr95DgCiTQMu+JLv05HpXD8w1xscg7
zZsuank+obA1FSh93lK6YBFDFdpeBEgiD4V39g8eK4ckt5rW3UNqjVz1nDwWArRCO8DF1W7Tmf3/
mR1tKGskYbzGqdEhPzr3JCvsXko7DijmHio3C7bSi628/Uhq09Mkj+cDI3F6K6kbDTUSLxOJBrBn
dU0xcoJVRdNUoaZsqcl8sbPyahqSdwdVHqO6TC2xxS3vhclgBVPhnvj+OdwB3snuvlfYRMKT6Ozr
VQpEIVJq9LfIICthFZHEU36m0b/rNUUZIee+x31q6L5EhcTGi4Mcb1IZ+2yNXy03sqjmWXeCZG5L
TBk7C6dXZFV2gw3oW6NKVIJufeh9x0iDxfz9JMdI2soCgG6bX1udkG48Ce2fNeH9jK5G/VhMgmS3
AEW41iBpYdP1j8xVhLs00R5y/TK8qaD7CjvR7j+k8AK40FxImltAngxS1y0liYId1BqC2YcVgX/A
uY6OgUNeG7jjiX6l/wYIo3XQ7rEs3LsVWpVTIKX3R0hvzLvgy++gtz5mMO3gZDMJcnbJMfduD8Kg
qaVOM0whZCpIFmvErHYcJQHv0SKKmmhoyAB2Lyo+donuV2hQgNGII/zPUkjOuc4i1aWgcpBgoGbt
eZsTHcxKBe2hifMvxbBxmOINiLH9LLrpQbdFdEFl6aWoOnVr+eQfA+/RHVFyNpcUEgR1eKTE35Nx
GYpfkWTJkjujgAPW6mi3v+yD44ZYOjaozP7zWiFpjJnYkZzl9ucwaXdgFJxnuoHdxv+ldaOcu42S
F0o2U/wxPUy/PqQ12u6bbQCHyVK9cIFQqJVptbjYQC3oQHTrSYrZaTpF+uJWwCd4+8Egz+bq0FTV
7IbBhleySqWN3bBLwrQkpHAlM3upLM2ste2MouyrC6z7YVBZC+GpwLAnAzk3I/fcIbaOJJOI/lQr
eNT02Mbnl9BSIszpEKbo7jXOYA5034r1UzRy6e5LlFq2yqu43VYoceo3jn/GHz9jMX9gZa5CdYrg
oFSM1obrr2hetL+Z3nz70DWLG2DuU4Cagr2saEs+pa/IJviKxV3/V3ysZ4ij+ZEoLQPFb2ISm4hH
yMWgBBlTr1Q2Pvk9Qo2AjooL8o2lBpGCnI8qM5/GjQhRwsZ/YgjDQMVxE+R5eSfaHdnSqRjit12g
+xuef/v8PPKVq4eaMPXrUvFDLOIp346lh/3fKzsREDMwsywz085bSBP2jvRuaAqSD2ujOEfceCCU
acfDioeouBFfgvJ7tEulOu0vt0HQEmrFymNDqRLyeR6vi7+OYFqeke35NVNPq3liI4IbcgyePpms
QSdpvOSGsdVXtE2mfinU9+yrOSV6IoShGx3k7Rd3CV+PK90sBb1ed0kYAXyBbM0Ktl4H5uGfGke9
aCjB8h/Qny2/G1ouPPXy0JnpvBzaqwcz8LzPSr6WO4cAKN3qYAIo/DdHZRvFwJ9eBbx44tjLWoxa
PIZM7XqYbEHv3sh1uyrJekLzevyFer41kuc8bTByMtzzwBTfe6zJPzSZ9zz2b6X+VNNWJ85aMP0G
lZ19pocp5HNINzdVf5TroFTID0ni3Tehk3q8pnCeSnptgAiQ1qPcs4TnyGQUQK/tLEUuvn3XFDMX
jJUWRaJib+96rVHkFbzzVMJMaSKewEut2EodEaZtOnJTxHqv5bAcZBuGHG9Sd4M9WrsGw6w7VaRv
QjLqZiv72tdBTUPfWOJVESSlD5UeqZwKWO9HWFGI746aUlWmJbwSdz74qfYYV/2qx1usL05SKzMH
sJ2YJKYehYVjon97m3bv46UiG/j5pCc69AraI0IdhC5zNJGzyLdkaJXfAOetzirkAx1q5YPK9UQ6
3kzm9rx3nNm9L2q2mLg7lTJEUNvFtZhW04XWtsukTWwpjj/jsbQ+LnQioEnwnkWxa2Yyib36bDtQ
52gRjbGxARNRGj3MtXGEVsbHl24SmPkZ9P4br5zX/jN7vxErguYNwlhPqvYNhQ9O7/QsCIle44J6
G2Hp+upciRLZKe6piwmonhFExF0DXB4QOcbndhQiKVbboQp1ik3GO3EQMhyTvXqQCBRiedVS79kj
hwtc6lgunUtioGzNGBs09pij8syOXJaUlGzC4eLuXFkP6qth2XQATyS7wq8j6yzB6/TnvYmvzKA+
O8WvRIkJqpOX/VAwFyrnvzG9xn85VC7JFKPzQRWq41KG+qQn62sOxUcMjlpaRpDFrw6lPQpkefxD
yNIfHRKGCgZLM7tSZGNY9t0BneFBD1+kek1YFkSUdoSAOxIeek1VJdvNGFRRHyTw2g07STy0vRTm
mvmzfkl4bRCuErtw0KGAwTqH6K4gJXvbRxD8Yg1Xr55K6vFYuKTmFTtg5FyWqr4eeUxF6dzVSAHC
7pZPll1zY0I7mL+kan82sDo8d+vYkSLSVHyYa0n8hTkpssvCsSFdd9ykamRMykUQ9YlHQSMHbAGN
ZobeKhObbULYuvJcPXPgNAtJQk+Z9VeUFcpQRaGezmEsd1x2/CumfsqlBZJwDTRJ5URqfa+wLYSw
+aFTjOJCqM1mx+DRJX0R//aqW+/rlQ5LBRXAcFQQkJkHihdFjOGk/lZ2Fbzp5RUSj7WuS53wvMOG
CqcC8OGtiyOkdMGYrjhtDOon+Cj/DHg/hWWtLIBiUgq6LMw/8+TWkw5BmdPlRGas7Sg/XmtNlgc5
VWyKKKchPJjk7BbDrcNg25Iesx/Go/fOxAJjrvbb6AndgWSARgSeKEtB1BQ0sZxMQz0ljhCu3/zi
NCPZUpVXtqaYvNNq6bU1Hzqho+3IGFUX/PQa2/y5u2fqaz7/O3MM7dquftdLkQHc2Wi9b9SjTVd4
/uaf7bWsMjiIMF7OXbQBgpjNckyBDq49+KeUb9msb9N2zvMF+s8txEElfY1MFG9E0UdjWgL1Z9us
TerGPs3QXrCbb7hXrHas/XT5aJg6emAvZsS7aYkLCnOneaFeOJ6fBi7UklQDGY6I+Qa6DqZA89aU
If2y6MS26VS7TItpNjIraDjmSj6/T+h1Op2xjsfVwTXzLreRllNViq8GUp5CA30zdiX/hL4CpkIv
0V8Frc5kIg3zg9cGGfUjwhr/SlZ0/WH0TE6zlA7xZVo2+lYtVGsGiYkXFMdI31ce46IWWKzjP1cQ
IP7X35y3vvT/Fxk24NZsLxdACfGwETxtib7tBP5g5gu6coVQ7/IBA8fw/EvvRP2jehUV4JtZ3l/u
U+60Ir+3YD3S9I/YtTVz93b4pAfZiyPkt2YeTduuxMRJqL9V+jFjPOa3POO5vJ7GK97fkl4GsNWh
RyfJJuUO8+9e5qnU6uN7T3fK8O3EkYWFwAK2WWBZVESvGdYGIqMFyRzOwnGvCgMSOHH9MDwTBDNm
NgxqrImnF1HKlnnTCr697oA8xLXpTa4JTxsVasCNFfYr+jGP0rD40K3YxZufq4u6ezR3kTwQgPIY
pFoptjvkW97un0GMichWXws7Z7UAICfxFFWP0WvhLuKt1kE5NXTgz7ESU29H8EyWwm0nA+iVf7+y
wdAWZhBioMLuzTiK3w9YEMWQF5v7HlodL8NvqJsMBqIvbPOY0zKxE3n2HcVZPDz4/q4uu2d0ILQF
ISpsHXqRTnUa6tjzmWMxR585nBx4HF14vKEFvzWHdGsM2uGHnloivrml6H94x5Ah2BpQgl41m45n
wiMjVjb0qDcghyjHwfBg9M9Pc/nlwM4qFVvyiQWr5hjFb+QTXwfrpepKcnU2nUP0givaXqjUeTlo
59zvjaXedJRbcPEIFySfhix/5uCRiTLUSQmhnsOsCiH00QuJ8Q6sYUuqPWZBpSOa6JlaOmTkmFum
gvgdlmGFvtYHPxy0S/0Wy1a9B3ClT7OL2TgeB6O3xa9xO2dit2Xf56xkYH12L0FXALtCnRSWcHx+
Lwi9bpBlLld94o9t9+eZtdcq/UA5EaPlNFxpdNspKITt0VwWdxn8bPBUhQUMEm1hjewtugpHo/wK
CQQ3vhKhvJWz8qgXpnW7Of1nErszrRf8N5YVgI7dm6jqjBvzaxMhavJngdrjDbDtxMzItHoKkhFL
o5k5GOeM0THJmT0Lv/N4BSTGsIAoeGPELPZidvABus+PVf3spkxHzshdAY+0wUwUe7nM4fIuPR2R
k0CEP4pYPkKHrFhMp5vyn+G2iiAHrp8xeHcPv/DXAYyCytbXWOLlVtA+eM2ttAAd5JUffKkErB1+
1KAhNqFMmQuxklQ3LaSqdZEyuuwwqc6GqwWKGMERzxSAlwZ8Ko0scxtTnUuQlRQO0bCjIusdiVL5
mgDJEkHqHVcqgsNf/9Wbq2kzheRxUrxB0I2+biPhM+leLU6RSL5q+f85H+vVurxIwfm2zjl/CnbW
foU3EgQAR5tJLZ39eSM5yqSAEk5g++8r5JnljnR1fcFP85+wMtoX29tv8VUUZcJYAVHUH66BpLCM
cnDbr3WIO4QMne3qCY4lcd2WFTp2aleHcAHFJ0cg4YUbzy2vPAYms+cx/zsfVAGB2nUv4QfXGK3T
fOkyxhkfAeJ5+yskPt6UhrbuKDSXo/aSwHcqCp/cM28bDx4RqW59tDepBtxpMiaZSG/uSQDzxIUX
lzHCppYJ5b1TU4Bn596fxbCq6z+8uoBRy91B72IuWwKX/T3K5jJ+rwRC5zKQesPvKcP5zqbemY8B
XYqwsdN4pWuQ912oBkEsQBZfns7ecuo95riNx4NYOeIw3S3brsVe9jTctZBLTuPQUIpt6ssXAcbk
wgG/9fZsZac6fo84+ng6uXASew01UsiaeL8wIVYl6WgCMUYABdoxY5DpzxODsWHF4OZJJxGPqh+f
ehibhJbW6LrW9qYMpIi2z3GZsRSzIIzzCFlx4F00asycXf1ftKA3iju6uZ+b321D/42MLqR5ZWgF
NEK3dbOvYqVozS708/2i5U0q+0jBjuFemHU0GkGLYeeZN0YUZiwDOotCqmeWSZb9POC/jOP7cAKO
pCc4boHbucvFNPPH9n+rywqaksGLpNFoxAKWfgrp4Ed3GT+1Tl2/3qgqYoHcnW+j4N5RTIMAwiET
lEaS4dvrz4+GG+wtD2Xef8qoEtWzaXV/9keGceZ/+T89liX0pO8esw5TyC+mwd4vAkoS2i7zfLak
GCt1O44dQrnJMI8RpqHOzDYFDTuGOhfVx5ji/3At5P72P36j+ebw6RKeDWiSJoJbFRoRRFY2C+2N
av3qhGxfBAGafftvW86EMEWAsXCeXxDSeOc9TSbJNJoUDtiG3ws1JZkxGjf2bMyzdj0+IYwOhu0W
GJ6d+tZ1wZu+58aJRY45CSlIMpM5sR7d3M5kMu0Sk8gUNwfAJua8TeXdUh9uc4O++Biu8vcpjWYF
37i7SYyIctx2bg7+RiXRWpZHGJU9OKwtW4ZR6kGVP+flSkCChmaBGc99l0GXOqH7Qaf9qD94521u
TcbAOP9FKZBBTdW9ZovaKkfmLQeufHQ0KrfxbcuWXNYAUyBRdJj3uBYjCt0rPzfUb9TkygV45xg1
Nowbo7Uv0d9kMmbgVdCcO/SZ++6CP9qrFiFimHUmER4BO1nHRz4iLtS0Lt+5JvzCfi/8CwSqiOpt
GX/YM3/0ouplC8ybkHUIqDnl/tBq87HQEgcj8VsSuEd5bfe9Q3nfDxNEJHp7BoAC2tMiOOO6BIRA
Ny7v4IMRNCITQRpZl6VTlIrN+dK1nSj82rF/6ZkpLNnoMQGQJNRYZqB4kUDROQogBfYjfjprxuYE
/Mofp1dWS1UEpjUTppm3DZNco/u6TniOV0HXQ+vdn7d7keO/i4jBQT2gZCiYGHFsL0kQhgzmY7Y7
Sq9dJm/7XdKtwna8aBpW80+s3zOzgXijVl3P3LadSuIt4yrQEuV9GKG9QXfr4uFvbur6NKZD6rMK
Qz6Yhi+l1Cr03oAQydlt515pLbCYyoraJLtjiecMm0SIk5BqYRqk1gtqTWwQxsBU+14hg/rdwdRc
cr+GH6o3LJQ6jdHrDCz6/m3ND2qbqo8ghevN/0uvufwBD7UxMXk1ZgXaaisQxV+/ey+7KT9Bd+Gf
WBa4dYQdQpvh5VA1mtQjHA7ytDV+AiHLbxU+63qQZq5KrrEk3XXEszPQ/pvcch+JjHTwx6zfsZUG
NVZTDu+IC7CQVKJxRC4Us4IRXpGT79kY2LLLhy8JYG7PTh9NlLOgKQQ1Hufrv+6YUmf11EmBaXL8
6/tLcLMC8zmC4FQGTlCYGThYzn0xl0jiyjs9S8ZwqWeQ9UCWAwgN8qJ7+tQ1HbCZKBXenqG0oS63
hpPV2ePl+TmRUuSrsahbw+21GYfiaYd39fmvMw4HYq8lOZfAuSwOPiTqetnqb62l1Z7W4qqU+Ehr
sxMIo2zoVVYqepv6877y8NFytgece3MdovyQziWArRxV0qXwEaNHHhzGAo01sC2zz8KcxVHzxicC
SphOOgHB89q2wboAwQklAgWL1oStHXqFmXNNIao4sr14jHYILDL66chA1JRMcxZTAJYxJ8NsUsbj
zBRcM1ANR/VGIhGMOOlJkhuUIjNyS9Mz+3Ca6dMLPHWwiHGRh28YCke1KoJ3nHmnku5YqPYfIV8L
u0haXeQhv87N3d6/Rh+gCpvl0f2kbDO0JG5/yd7r2Zq/T84RgJOmWOIkZNHwJTJEk2isebZJY7MO
c8c/YVepTGgwrAF4SOYIcBomrEhW4SGH/D+nhqPmEhRoBIY3skEBM0PTGe9eD6B8SX3VogmcgURb
919YL7i5LKxCRzbO8Vzuz3CHth1NPY2TLJbeqa52/t+Mt316CZSnqbvxWDOwTGj1bdnUS5rBg9vN
uEAkUNpYTT0lBs7BlBcoFMK2Li28I+kM3BFpaP5uV7Rv3q0RY4mkX3y59UsDzy2kyRWQu73zQaFP
y0kdO4JJz23k6KyqoCu3dJx3FoHdPqE9UiMgsVX2LHY/IBZ4fmwZUtIJa5MJdVaEpQKr3Jmicpkx
apzmOUiEpF+bZuiSD/piJNGDTWV3nC3zNw0fUsuZF4d0Gz2URYpwSigR9MtIWCVr5YDrCplUyeBr
+P5pHRordWb30O5w7S9N9nohXwE4ZKgq7ITwkERUekaOdhhnNJLrMZgu5sX+B2ElnoNgesPFtFCW
KtVv4rcSlDUZztaZG6OpTLlXUvfC69LbLNRmyEZqO/dFfKMm7/H9BA/jqPpNoR66YYUHGYn3ZphH
dUJN0T5lcM/EK971cWEzemIy0tkRvB8dIEDUQdAav3Gog8ToKFdlGiA3Y12qlnEsKH5DlJV6o5mR
52hOxRDLKs0Ym+475mWShLJjT70j4h54e/OZmxf1ywJZsSW9LLEcSUovaCCk64jjZyOEnwKyLlv3
I/t8x74fsExrggZEa8UsVjfV4lTpJqMXjr5H6HZMO3IU+VyT84/X96OR+DKyStnTuiRS4EnJot96
NY9sSa6Yj0hNhwgy/1zEcU8ch3/GGV5RCTm74RhntfRlR8uzpHfnF8dxt2OiiptEsR4ceyVb8Y55
l7yIRWNJ4hle4MeXQSn5Jc1ThN/ioUezEQXfk/Y1QaTyg4C+SdUhg2F+YHenT+R+PRfLoM9oR730
IsCn/RTmYN8qW+Tk8SRzGQaS8YxHAIxdM7O7fMhhqgpmnq6lib0nLAms0purGzQtOjmPlJ72zwom
TohUCzGssEdDqiEUYbaQvK5FsgKLhOXqmGoOu4sDhov/odnN4mSQO75dNk30O1OOjmq8fhdnCaXt
vpsPvarp9TMi5KirLhRLSNhn1L22vP5FYaIa6BrMkqLdlrYatUulhkMyTtnWKiBicEP4skmVNuS8
kUTrq2ERTW3qNctF03HzN8Z1CNkL9BLTAh6kD4twgQp5yM3aoT6+rTAMxxfNraEapsNTpmCAHKkb
EVwhpMWo6LPWDGyy5rbciiMHwF3j7Kj2oXG2uKeJCw5J4AjxGJpufm+cC+Ok0KGCXY8sQAATN6Zz
q4MKgUrK2wuw9LE6PYvAlJKlbVN+Y1Ae9h87Q6+i/JfF2ABzOUvumIj4llWm71MsxfDqId39Bj2S
jH5MOR3AzftBQeULo5VO84IbAws1NhiAwz2qnz5y5BICJJz3tuht3eVZ3V/rtmFmCE28XLSDPSNZ
eKn0yTrrC2adAthMvVypdwwpczlomk+cAVgaxTLMqd2cLTALPttq7vwDEd1gerXxSdMbKxVtbQye
8+pRJYehRVJBoCmz3K6aC/FwA6WHpC2VTFFNOWab6IiqP748O7uS0IePSBJooMx/x77ndipSKNV6
UniMNM8XV5gruhdrYJxIh9gr8KOvY7friUFVmOTBJJSR39x6JsdZ423lAwvEkdB1Ho3kYGIpRPEL
k4symEt0k/Y42CSYPtQvvun5OcP5XH1ja9quMra3dZV0+86SAnWA+Cb86hdgRF2qiTebO8U5XiYR
ukmbVMFDnpWMNdUOT8ndmlWZgipjsLWnFhb/EUg0+a8gbX81NTvHVueGpvXRY4wjsP1ebGM3/con
bUdbB5ZSptQDbRLe64RavFQd6U9TMitWV5KNshrkIwpxFhmgPktQ4WR98ZVYPxLDDGOrSKYhr6+a
o2cF1nkmfb4H6ujXKmPug65XG6IhiCEBF5XeOciJfKZyq03KxuTImUHmm8M8ONzNLQPMDsMroSBo
cVh31sxWAv1l1G0sF9HubFTjXQKesWov7NZPZOGSSNFfhjXEgqQwXD2Ng5W1bFU5/S/IGsIhPc1n
2FNmEV789NMcSyEpuvUyYaBJEuR05J9ubwJpPiW1TSDWIZ5QhU+mQcB3X2AhpiACvJNQgVuQncBV
412zrYbertpVHqmdunepiiolhLqtZ0xy7O2WB339XQ6AvYHXnV7a0bwrZ0Tezu3t89mvlKVXkvjX
1rA/HlRaEV3k+p0Kqxj9MZZis+SSxWSAUtbfp+bgKBTiGnx0rbWRzeqGNO3QGWGZ9wtv9Nw4FTeL
0p1RCsyPrAT23yY4yQm7janSswHuxXh9B2KbyrEMg5EGw289tan9huFnXqs+/P9wj0IJhUCVA0J/
vzPgc4nX2QGsbZ7HXjdl0JEOMdnRgh7ao6jiCtzC2HZWUGawr82BHK6ka1wAtcxtpqttCUKCv+IT
aNCPk+ALKY2FjFtaXSQ21aswY+Srnox6SkkwsKPmgQCG/iuvmo2MALDXWihpeLvxCAR3pHvpKApR
9ubtVmkBIP/SnSKvjFNVxvsaJkj+SRjG4DcvJrX1wyse4b6m9aRjgckGN8e6tAuBCULvkZ3Dkuey
43Beij1dvD/IHyS5j/gaBP3nZaqi1zPCxYrROXLAcx+mPJUQGaC95nEiL5Xud9bXsxEkH+TEwy+Z
2+rWKsS6nlzqcZca4Pdu+TDhBZHwC9sbk3S8v5Mz/DSEzQnrzldRNmnZi6+GfzY8kriPy9TQ/oaC
SXBJGTHYKfA1O/yLukob31RdfK3ZiAwZoBtnjnnxBCJFzRx+OJeRpsRGVdq411fs1t2JpZzVGj/D
/pEizDYnbqyVfDO35Gp6T45Nfmjbd/PoXhXKjanX6RjSr7+7H4vpoPqfQHxyaH84BGoQp4/8YqIX
/W6hrCOUttrPlgOpBE37PSs1Zn9TprKRo7KWzMAkvwv+QKOlVkW6Kws6k2s7cSe+qkw7XHkXOpSq
FuhNnh0wWggCyxHudMGFGqc4ShiZfPiAHnsWwelxmdMaVHfS3IglP4GXBXv0P5SiaEECSgzxEVRA
DH5E040HeSf8QakPJWCVMFTSKYSsOksbDLhLiG3zP+Q93fo4VLJxYYPhrxIlfgh7J3I6U2lQZpMN
Q1m24UlfyHPBrCimgHtXW9BjbTRrPzH/YOe7hA0Iknx0Oikius+UtgQeuJuxuqsGYn+HS1oBnOXh
GxFAoruDeuTUIQRYL+rep57OHg9pkKXDx3LzbIwXC5lmiCByjU7tA0jVTqR90ylvn4JGjlFlGdUQ
D48PQRCnAwMcwr/32oGSxrQzVgkcFnBlTcKYkIF119FN1juV7ui/bjfOagOPDMuchKmd7vGYTpa9
QKrWoJ4S4vyvtXYFVU40LdgEjTnzko2LZPtAU0ExSxrLLBw9Er9CIXH0E3iR7DPZp3H86VBvYUhR
VzLJ2oX7Ht6cSiiDC4TjMALZcpTvEcmX0JMvPin+RdFDisYYAAb+8w/UnBn9mrz2WNkNrOXMJprO
9CaIAlm9VrhwEb7EHML1TJScTQfdNYi+8y4ID43KaciynJ3dzUAp1SGyDv8RvYdS7s04xdJRSwoJ
NIggSy/ncnPnFwlWZ7xgMlv3dnWQX5eT48GwXjJW+fKuLuFKar+AKLy3yFQXWpSbdc/mOKNZ2J0+
XOHazD3ww6aF4RPLI5yrrkYYNuAo7z+yB3xKA5LLp2QwkzwYE0aFUy1YxW0i0kOsN+rXSY7MrRBz
j1ZFlQdEWfCPrAz7Kyiqz+cthykA09gVoVppPoQ9ZXmxrdVX2dN9pqOHTq8o34P++OJKEVRbyVoJ
M4welKnfEw2OGtJaPOfa2WuC4uWbbmQmtMKXgCWMYYCbShNF+iTCaBy1EwyodGMsBzFHqlwJdWE5
5SX8BQSu2nbdi8Drln9VzCqk4wD0CPwPgepKGgJPkYBoFqy5bnf1hVQrmS8tS6n4dZAHs++5RYP2
eEeDY5s/UIn+7IMcLe3BJSDof0PXuwackUYvTPOirtaPeuKxKA5QgcX5dc2e9tJTDt/JPxkgpKyA
XiHn9RzrKBNBQ/OYJ9e8QoO57c11yFXVzeS8NlCgWABhZRGcYp7Rvcqo6CcOE2t7jE8Y/rWKJagU
vGsLWD6+/Jf1Vg1QfNbGQ99c+mUL6+TP8RMZv8mPbZwBVYThhteM3+F4XMc80/3FiLKqeFy0e7BZ
tXfmwHQbhp5f55B3szQPi+K3QSfY8WtImhDtYzVaxw3qMb9h0PBSVt7N3fSmyRhtWItPWhXKxcZA
S//JVKu0HLiWxHAIAzTWKpTAu/vzeUvExjLKJnd40QIBTmkSKlgVS2Swn4sJbw5CmQFBtj6v2MDg
xnrIaNiI0BHYmitpSv7tvo/LxUBvWb0aiwfWgDEmrSgZMmV7WRvn0HVgT7AtsTm6BR8PlvoxGI4C
OT2iG5Z3QBbvj6VpdNzD69qJXqwmWFq5NFhU3p0v5NnfKDqZRHa7YITPmbOhw3tsvBum7J92TZk2
C5/gcMhD6uFtriYN6byoTdpr73LGspeeqS3YvQremaLLD4xhoYsG5t9kkusYH75ZHqv1pbjitweK
6G9KQ8rwnn+NuMg/aRg2b9lt4dYxgmKTHCjIiEoKVPmQyy4V0g6OHFh3fr6vAtP0bkx6/7snVdFy
yvYtJn+Zj4q7yzK+Qgrhu1owJajtYS+0dxeE0KMXqnTRFP4llmHDtYzpjLMFRy9Zi1fieBoQjHXY
Zp/UWJbEZNF9PQP1N7sF6mPdf4PLZPbOXa+3VUjcfoXc6yfxOZ4IMdZnkWwiRTeczDuZ8ig7briZ
jvrku9M/mcJLdNeSGj6IU/P97ggZTCaay2soGLKeTWkZQq/8xdKgs6BpkkQSSVUVDkubInUPOjc7
Bo4j3WOya2o8Fci5b+vy0yCz3rq/cukUkOjbJFZOb71Eqlh1cko6+62WlnnqwYBRx0WouUtvWP7H
IYjvNaZultn717M6OKbVNRAgiX/5aPDyk9Emfac3weMqMuxsnTjg7AV/Cb2l7WW0BBniCaYMoFtG
tpJKJUGdzQdTGc+75FbF8Q0Xt34D8qMxezbS6nTnAfWNqJ9ZDXmF3KUBxPhHpZqmVEaTrXVKFyR3
Csh998+eu6fyfHGum5bREaRyrE6EyNFZXlJKZBg2YfqRS5Te3i3yG3Dd1YOZbVtsvaQji6H4ynV1
c0ei/NNawOdkOQefjmCoBWJHjaZlFtd9TI5yBX++dON40MqQhx0eaD4Huu4nAgssnCLMmR+Zlhl2
QaQ1lQ1ZTdfzkc7BaUdFFjtdf/5+xNsU4HHJSeJci2TKACYHoKWJ0B5wyIgc8SGHeUZIGNKwJ/pj
cCHusSa3kVv8YaSX+4LDZoMecp4Tt7OlLAPEDTy3o670rvp4hhlxpExtjAG4OngGE8fYp0+ltiv5
hiXYoYeRqmwyIKx5wJQN9QfG5+e1PzfIRjG0JT1STlVaKiNNPCuBt/cb//IRo0byft4xxR27UMIb
F6Y44LE++EDcN6Wq9o2w1bdFcgl0XMly+E+Ijk07NYZgk3KLHVT7NTOCjMdEUx77hpExMdEJyDMU
eFaVTWW5X/Cdu01GVRbEDTRvdlqw9x4yZxyhZcw2g8zXjrQRVjmGbARMZSVwtplXcgTHzp9allMF
034Y59ENPANtgWlriPPYoagC/QtkutpiA6zgAJcCWzQ2rG3s0rbWRITbKPONWNT1NeNDhUq2CZ6h
MrCXww08oDRoLcTjLs1phXPrAWGdIflbkxFTbqXyVbi8X6oUW09JPPBg+9ErLRHzH3xBmweNXHji
qK2Og21sd0MpFx9D/JJ2VwKAdvPEM4KjPxZg2Vmz0aIEw8QLCRFCeIrQp861Hdr/JzWJxGTG0YiL
uWVHFoUOc5aKhKSESBkWK2mWrvovBVW6cNaZ4ZcIsWbcj4ewvYTl4lgI+GrtTCdOeQM6JKlhxCYh
YcYdjedX1vs2jXDUZYZyGboiNULpEogdkIZ9lbkIpX21v/O91alwtYyU0IWa+Ty4jWNL0a2ocLwx
+LpcnAaga6zDNz/3S4IPmBojd6mrpK7PIoTIfghkbCUZotxDc8+SMYGSyOV6bDqyTVAwBo+ODjBC
0Lw6WzTKQqdDugDGYRBv//hCKdvaFSXUIIQIyHWxgzg5aknIAIPUzaWBdRqcvhpBh9C2Ll+5jHXK
fYQzi5GleVLgzlB/sl4unM1livr+tKUUIqhwa3PkqkXuGmil6d2how1+8lKyBeG4f+0GXIUFxj5q
pGuCwTKIiJI5xsl5mJdUJweESAytKXwEodECxcCdTKgUzI4gxDL/2maNDG4BZbhx5I2w5ygQuIdY
Bt/yYzt2m1xGHD+xerZhIGk5byAPjwQlQ+MBpKNj18qf2NqrvWDGJ+ZxGlDk196GFEuHW6hf+6yC
FdOKR6xvHq/sNbIl1WoTSc558u6/ckfFzZuY3PCzUvfmCfG0Nt4d9UGYe22FbV+L5GsEV2LZakoQ
1gQL5Ur6+zb52vINNU08qwgN6ERoo8SfOmhnqcd17Fi57RSmQTGnPrpVsXekO3EpTZkb7rb1Rfd1
vPxW/RPJrmLni3TzjzVQhBRqqNhu6abBWfY80S6IvmlIKqisfv4SH80tlsudUNz8E55pE0iWHv7X
dhaHq/hXOiR6wurnDVHAR7Tv1Ed8qJ+77vLBl0hvPA1+tTf9loXBE+bC7tYgRKLdy2KcCq9/POQV
y5f5tpRzoZ6P6jOH0f+j/FuWQ3HRVGXLSRCtaHI2d8qNDqWdJZTuLDGe1zbKNQBbypH6Bc1JsL4+
65rLrJc548b0+ZPZHQ6BVGDXpXFowFaXnWuuYVMljXu8xTZhm4gjyEIi+AClL8iG5tJffkOXL4pI
ic/Qw3ZJz2crZdjJeV5pedWFjJ7JkBk+j6txROtoIIq0HNnHE8SBJ6UJ2CAVB/UwUrvaBybJzQsS
MXqQ4AaGjUTdXoXxBu9lzgmB1xTt/w9UfGoAIS9BW+wo6ZruX+1mujn+FSeWMySs09PHFIT8VLNM
Qp3/364e37gFlpglN/Kxh2kaPJJdkgvlSWkuFEmnBMcDZB2d70v8WIdIHxpJ/tZe0bmY5rarKP1I
JU+3j02zD0cbNitll1K1A7wqPjWF8TzQpI/WE0Vii4unieitSJokx09YVHcQXIzFQG53ZA7hk+E5
1TzDWffD3so4jS/p/CLe0wRrFOldeJT8AzQSgYi4lYtOETb7Lq3oMHVInK/l7e0Ki7IDfbqxiKao
zZKAh3/Ef2/LX7mrMtT4tBO5g3Aq5hPlsPWavJJOi36dmbnhilQx5U5n3HES3s3Vrc6MetqMn1HA
egawnFkqwrLNJvfFiFEoiNbDey+RVSpojjKWEBuQO8iqql1iHce7wX770sbCPq0Qzq47n5+e69aA
K01p5Z1GIg1PbUyqoS0ilsgE3fcg26vAPEs0FqvH8h6Vb38eYoEigBJCfKE+BiL9HLj/RYna0itG
2YvL70CtMcBkf/7Blf3SAoYYE38ewPYBCvhX727vyItdA6Catkj36jPyElhMS6LGtJqSzLB3iOPD
U8dKs+yB0Z0q1rpTcGrbbiwvgMCXxf0frszgN0ECxs8PSPLKdIWsQ7bW+U84m7ye4BbrCJW0OT4L
f5u9csp9RZ0k5PJMV58ufoApXFe6joZFeit6EABPBhfaYyeOM9kYzU2Pkg1HNsyz0DMm6q//6zo+
bKdYHCcf1sgpneRpHkRb4qynqlSYpVDUTElYmYKN9np2Jnflzw5+nFkvcBP6EaHiIybYusQj6DPi
pqCO5OGNgQ3VQ3EKCqezPIBk7vCNe5JUqwt5TkAjdzieesbOjfD3ZTLz2q6U1NqUaKaIc5RwW5a/
BoejdxHad9BZhf0l4CMk2NnD8VkcnZRIwh4hO8ofBqi8ejjFLoryGMaHi87HI75No6l2/9nzt1Tr
/yrh64QXMSW8vjoQNpsvh9ro+DrrXcCdSgDUv8QAVFJ3oerI0FSbKj07xidjHmAPmvOXxdeqzcEp
XApGqNMQ15UM7zBH3Bt3LEEOzfK4SZPvWeDFj9YgtF964r4oHIJ6fO/AKQF3d2z8cIVj3Kn2S2WW
/YA0w6lGbIdXoxRUXLLPfZPGFa+koq1BCl5Z1ck47lMI1l9FsMnpgCh7DmTDHwrFY79v0LLd4NVc
xQihilyHAFPlqp59JIQiZr+DLucFx4vUKmw7u90WInzzkw5YbjFKU4ViQ8B8+j5srmG4lfOzYT15
sHx4q5OFJlmjQblR17jYmoTCzNHZNEHeJdFn1osMWu4bWd3R0P/jZOeahoz1kzPFi/qtNGsAH5oc
mA827mbYmX/jKv7TfF+Tr4CJmSyRfKU0oDf8+hfoJ14YVe+E1TurRyIHiR7b+mTsTbwuV4X73ur2
I/lA8AtrZNEj1cBXcey7GiYhsauyLdLdWQb6f0QWmBZzdt0tlgkvm4NHbCdXvz9rSEPsVWUrx7h4
Z7uqk75d5dJmwot/dA9bHAe94EFDwRKP8aLQYjtMxhzLOBg5cW8Xf1NjbvMXOBUieYrpmNudfVDD
fINg/EC2uj7dAWwwY+gOWzPGhkqUNdy/p/A35tOzd/HrN9UWSX99zxvDwM4OANvJNNamB9nk8RZM
M5rdsNwmlnkKzIsGw2NGPEsVlmm7SBEtddxP7RGi+Iu74WIIWDtlhhsNdswqZLzXbpSp8DRc8SKv
KnUlA5B0n69/Y9l6D7Fe5n0jSYIXyzQFaO4R+O4I93UHC+d/86D5ixnjtWxDd/3pCNAVpQoh/rIn
7l7lVwUUUTA0VqUBhhNBd7/CJtZ3k8rdGXgTuK5mcyG+wNwbUMYqQKL4lSCxI/bVKUanYOrqam5e
m7YQbYbU+LC6xoQ6gt4FLqlUXW/XsuCRyj0e4/7QeYqUCWpnBKQRrqW+uj5/4Q/c8B1Xi9hI8Tn3
KsfgEOEv3hQk6IaFkkHVTcHqLBo93ZBdCwkE/gO0F+8fkMQqz/79ux3BidwgSbSdISS9EYMoZ7fX
1qYiaCIbJ4wRPLM43shY1we03/yWd3Nf29QRWCfzUzMQ4oSVFUlcIrUwu9Qi4OEk/muCQcfkUJtM
N1X7Tcl5soF39uqroUsjgoRApP9qoUfs4/lZiJvGTO4rQydYbD1FDTjHhxwggtkluGM5WgLuZdGE
gjUDn9IAwKcNfUWDTdJOzFcyD7MPtkhyzuy5WDv6GUsujz/xs+I/Ki4amm4vb2qVZy444FgAcbiv
O9vbeYuUWWlKeHjPimZPb/z/wwxdNMxhyaX5HMSoRwvdm0zlFZpEEGOZ/En7CrikV/InVj916rxZ
nu6c5dN+YZkPeVeprKHssUy7zDUvrWJ11pb6WJfYjEPcfeh9kmr4nNugZGdm0y/gP171hPBQg25i
GXWe41guzHBRaH9n1s9I9S5jPaleknxhZCddlvLJYFZKT6oTZN2MoJtCfeJtvc/HYxxpkUjn13Nk
A6oMRToDidx8iTDLDRNLDzGsuaQIYQ3LmYdILgiBsFt9UY5Y2+Ei8Oi/3tJLjMTPfi39rRrxyOmk
sKW527/4GFvxb04xhlaNAJi0OVUATYoJRecrmysdVPIa+2bMkIWrm+867WyJuRgaflgkt7EsV9E2
82iTrF5b7PL4UVaHlbD+jsGoFeZepV3IHDvZwML6yTDkEtqAchDm5jqA6BVIo6jtMezn6Q05Mvyo
1Bp6X6AYkb9WyZKpBUqVBwEatuNfmb4kTqwEMyL2S2rzZmACUQbFCPaAiDVaVal4RbfA3aFXLpY8
GQBnpTmgSHOrmWadKYgxO5E/XLDTh7VB5WFfoI+GmEVd43DU2/ArbuA5dFWwVHsH6sHcHjeoZUsI
Hrz15hVeD8Ps7/E62I9D1+U2nUvne3ouoDRFOWNmVZ/y4HwiYoETstndqkeUxBBPjJoBsx++7rYw
ayO+fa0+2P/M2egTdBPYgUkxa98mMiFekj8oHyljs1VigSb0ItgWrE/gISme4B9D9zQvJz82diAi
vfqpukVJYHbzDrT5N/KKXri64zI08LFFPpcO3quIBvtZP0e1hWz7sW8+2zZxcofi0qn7nUIBBhz5
/vB14ynq3lBc+NvoIjKSzPdOhgmHcvhPChFzzoP8OheHPnyBascxjj+ivmsmdOfefAaStyNNXhLD
tE5cXiGXZhDpdJvK0CUF+xi1tUrqahCjvJCeFOukAkPCE1YLvMOs/wM7VKL75WwB8pZspbm9mMHI
Wj8DB69uKhrxHOtrn76g5JPrumHwvrTuoTQJImsID9qTJ8HoazAX77NduI1nQ1wc9Z0Up22mwhiS
4W2X24hAQQ/Sah+/V/5cG99uUASDTVxW2ctR9XVwxDQQGl4tJE146mHuUrIMxkmTEYYt6WfiTKr4
oInw7ajHIoxJlWOTzAHdoznWlYso64y4ZTQZqMK8HHSoquLZgVvaSSOiKuO7xaOfQibCTC5NQQRP
sNhbl7RAeYM6MytFPenk0HBdjmd26QnFTgEyqaToCsa0uOF6IAOxaGl3l6jYGasIsnHt1Rf1HBaq
sYtIWgGravx3EpROnwKrP17BCooVlqsdAi6l/Nw8DPhR7Zu/FvKdy4tTIFzdBzNm7CVB6JvTQXGv
F6ctfUNjnWGD81zvsKQsSSB7OmPixAhsTPQy8jHJgITWBhXPm9Apwy+VYUy5VKexmT3ct9Jpc1Kg
khpSx+er5PaJOk+HC/6M8Lo8ki1yFtrusku1Zieu5Cym3mj3oTGl5GqGSBVayTjt8om6dMb0Z38P
0ZEH56JWKMe94jzvLW1jwbZQ9JemC22bfMQfnknB5qLR19y7ZhShDTPFu7h7PcpNWcgFiWgoBAqw
FRZRfQmlo0TVhZDsenPH9BaFes3PuPflj7xoFB8EdzBmPLDP/Q6N0BPj4mEaUrnRfVpzbB2skhHM
ru160vBltON0amwvHsXHqS7EmKYdNRZW8nuabSCN0wmUE97J8eZDdPTW8CfF7opTsEYuYlRffDVy
/QqA5YL+zMIjeDbwTeF89bPqC6LtQWw/O8WFFkp49dlU8fNo76Qn+rwbJa/phm6jsQ4tyhzlOOoX
mE9ejExpL3R8AHhaoKn+f2ww2UVmrpDxZiDiwp16Ny5YFiFGhmf0EJgy5tduhHU0ND79jrWI/MqE
kAPGwMYVdk+GiUV86VmE1NPhMxs3/3T3tvAF4jjUK4lZAhnfOFxXgtg80CvnPiSDAed0N3pPZUvZ
BWDp4GU5uHKL3ovpe1UYcgi3m0KtCmBDC5JMRU3fA1Sl60GinaMRofD81xUtm/CdpcTb+0l9HlGV
nZHJZ1kSbsGstusEZ1K31EbYHG4+pvDeUickLtR3qFicQCC+pLV7RcFMv9Ip8phesjGMkpL+eo7R
1V9CjweNBJ/2pVH2GVEfkgS1slRUwIsUXoJXKoqFk5gMsmEdBH8/9NIE22lOu+sihvrFfk0CXdKw
xfTxdGgxcWJQQ3xt5Hq1J1oN2mM7kYCODbeB4o4Ag+oUJc0FMOJi2YVcwp7Eks3ZTAgYpf8hUC7l
QkpZmKubX6wBSZGb3VPtCpYDT1+BR3n+fvCHJuCywQTalxJzUtfk0b+5lJyZg6CtWzEi2GojjAPz
oMaIQ3iO65e7prXU2UE4ArbueKzcok69IJzWrg1HCu3vdXKGeUxG+yuevaTx9Csp8/RGJiZU6gr7
8kONyItm47JcGujFIGeodp0q+AzSW+duv2h8SgmzRJuaMFYSVWuRL17fEuWwaKDT3xYmpSNv7ukC
EtC79QSRI1uJbNkvqHnzstinYtpU1zZEc9mwUmSm27V2wW692lkWNEvamCvmPgS7NmZV4NVUrIZg
reBczAW/fbUXixVQZBxOjCYbk9rT+YkrPSdxUwFupVd978Jf+sKjUIISJHpvTCT2gcHjyvZsdnpJ
8Go3Fbr1FTLHkgcK+OM+Dek4HcK0yGsrfUqLa/xL2JrMgRHuho4KjS7BVcwXNUUBfMfGXSnTarXp
SH89OJoB2OYkBsI0joloeqK6483RHazfDrY0L4gzMkn8uLFYx/W37Tux1eji+UR7At0U9jzKM0vL
QbtnVBxDOf8tKv+4u1wC+1Ogpkfs++wkd7SSHSHNszqwEtaG7HK2/ZWSF8c9VKXjUFz0vf0m1hqV
qWuk/S7nYTg0ZxS+x+caHebqcOkp3w50L/Y70fcP/As1Swya2MeHY76S/qq8LimC7tco2YzaFXgI
KdymeQ690uZ+YV8OxBeQbVDfanb+Q9vYkqrSChcp6NchYKk+haHJ8k9th7PjpEOhRY8JcZnaHvqk
qlgcVuQfzlafAJ346rdRpNqg7QVjeO4CFbylGdyEwUCr818CAqLd9rtFnrCuECSLZv1FZIPTGLon
91OSFF6aY0JGJkc3QW0uZOwF+9dUnnhV2mxbwaQ81v7jutI5hqQWC+cMbUerXDOzjQmWS4Z9QOMo
vYYIdQ4Pc/QI5CpY1EI7uqzCo2UVKnQT4ztnsbZvZc+qHhWHYBdvghgxIKg4D7NhDK6zDhp6PzQg
vNQJRuU8N1/Qrp/oDkqWEiKqV4WvNu64diJ4u+NtTpPUrTkKFQd0bnYxokb3ukS8eOkeMFlVhlXR
JIsxWnTbz2Mm91dQ45eolq7pw0ASFNIOq3To9C+WKueaHMO8XNZ59hNF0xBzDvCpuDj3hfFFPeSv
cG70pQ2+8aUZfcltEsGOT2ts2QbE6knxzIkB84JCAOivWfbwBbdIlc47cGYqWIoFCZSBb2ON5jfn
aeqbKWyn/o7GF1gP1dVqaGxeEC8LTzykEleQCjtIUOhIVSG/gM7QZcnLjqt6QSpD023UzeKt9bBH
/i0NnLFyzQ3DbU/oz1g8lLAHjBZBtu3V2HHO7Sv4kqfq1DTLLw8/5EjYFdNJPOkc30T0jN+cz8rW
1/dtx1sKGFtLQovRhTHQ3nK0y1F0hbRKyGsUCYF426DaOhg6UqwcPYQ5gMljC3SjfIwdQYXe/Vlf
vVgodiQteBnGakv+5AvY8u11MwRY+MOsOchLxZJ4c/zjhQ5psMzhpIMvzIt0JNksFGNc0FpRC93p
HrYjNyhzWVNPCSv7EhK9Dg+jUdnTBhQxJRqoqd6V1wgm1Q00+MCo+cQJBm4zoxF/PERfexeho4Mh
YZ0/uPJlAw3BfOmf7RkFlCIfB/Vd1kAeLVO6BAOkeWwsc1bq/bli+2b+lSTqf0+JLfc0OJ+nqid0
BBVqCpyMyWXMWtEg+jzRbEJSc1ROphcwqyNBvaZWDP11RcB8Vccovd6OoET35EEOPtPLVX8PiU24
hh2Uj5cre6Im/4s3GZKs098ddIKtLlMMbdrTgpOIhpBZ5o7YdJW9uHytYcy1p4ZNxkZ2vajGjMGz
v0zwlCs2remQlXIRuOTY9sfxp+hH5l/2s3zoTu6OxFaXrgDlHyyOAjZidPIpSIT8EhJYTCzsawjz
KUTJ4lyAFpekuKhV6coitMc//npyp49qpN8+aY/AEOEQeVgnrhXlq4oCSjfIXpuQnAqTEc2lK+zq
Gjep5wjvWzspLgwYRuBkhgIx6/gLjkDSyB0dyFu06X5KVwd+IDAunvDGHxVc7QdfhokBImcwajk3
IUh+z5Pac4kv6lU1wJgqD/Yy1nYHNTO7rtTUgIMs5sImwh5dVJyNbYbIYo1UpKxV01kqnWVkgnaA
PPc1e2pdXzxPX2xNckQqQjjLrnm4w0eHaXgsEhoFRpyclPOxZ1Ph87sWWDzMNc64psZHsRIeHke6
bfNeKNhoR8iJnyT8dVKw9wiNMuWzYK4Js+4GMcBwjZ9F85rbKnXAEZ8QEnXS52jWkOCpM2Ny4BM9
hU2G+KWgm1TP5/ZUUzlhuLctpUW80t1J+TqvoLgNp/9QE0NNeY+ahjLkNokPKiwbO9LNIp2NsU41
8l9zQprYyIJHYJlLfg8X021x93eE8J3BFhQamwEvmZrMffMJHLod+BKgSczMElFiPiXL45X+T/+u
KaQZHYSawHZwUhpUT7/aUnUdQvYp4lkde7uVG5jqUPp2Jh0R5sjKZRM7sVRA1ThUEZcY9jRyO7/h
73oiWH+G5YlBY+hLVtX6G+UwAx8So9hpNcFCCfJ1QwUbmvf5JncMbXyZj5yqNZ0vCSeETacHcpbV
AV0iByd9N1fPMaKVYnddMCVVHt/yxPxAEnqmgNKEWW6s739PSNoLdYJejf5QRE3yv8LomRnfQgUw
RZ1E3HLzOL2sCGLUB9uTK8fzf9CNsAJvcr4M4ggHraG2xHXRqIrhcaj2gHKChMNYnv2EuLyowDux
2BxYU1GRkM9h0iLQdrhyCyii3/Ha0u4Dd8B1VuPSPeS0eoVTIu03y5ia/tlhxiSaNKYrx/rNpzV0
42RYr+jWUaC1ioaaszxCd7wBj3Bqf8QdQZd4OXlruLtqkE469NTu0XwbcofmsrGH07oXonO70lBv
8kxHBeep6COoarUK5bAOpeiP89MB0yiBdOEM23l0pB+0nKXs0ujGaB5FsqvjEb4a/C0JAMJjTcGg
TEsTbdhxSrk7uyD8DlnSDwcF8ENzYZhZ8DwDIB9YAoCP0uhOQ5oEb0B0jWn/dWUrynLTvXmkxUZT
TaulHNycoGy4+YjJDZn3NFlxOrp6Al5kEtWhjHfZITd9sByT9n1aeRYGwD21uVSJtSrExJwvePRH
bfxlmFEsQ14cOqB7Ns8m2CD0w+tbA3FTxxU96SYRoLSRiMxEx9A7iuK6tbvjQKvGon/TVKv7vGIF
/A0PlWjDr5b7AS2rfQUOCbkPh/H/P4bE2e6kBmsO15Tnb7XBMk4bBzkg6F+HeROMzDCTQ43CljAW
tDAZLRhSCLOmtDHIz+snYDRzFy1F0R6psu72+du3niglv79h0s7OSBcIx/aHeYYOT1un0+UKzMVg
nOSKpdfIvg9QEbdpBst4KQDLL5TGpgZtVu18zwPWYBqQkbLM37qT0UYENZNp2AB71BEabSoO3QwA
iF4rAulOP0gXysn8o5ghmaKSsqQKGxpmcXUseIMgIRQVp/0+Q/OTVbJgLNqknnbF1RNAhEZtdNy8
Pq6klXJmOGQc4aIkc/0EwPCELZ32nhnMOPIcXJcKOwTibMrtME3l7BjmlqKXfq+/7nUJO+mhUzZU
DEJ97T7dM06OY+7Hnz5eBCfvugjUKvB0FJ14tkdwnwsGFXaXMOnojf2wrckmOh4sjEV6SogQPzbU
GB69kJGHgNuXF9NPs5nrxPtlRpfmPQMthHlayQZ0Omrq0p0fOl3xr3GoTD1ADztv8eL+s3FMkx+8
rQ11FwSTVlPGAXaiFHe8LKKUDoGwCgZgdKvrTZa5v31EiLIgB8xn3xG8ukqJ1xFoHJaXd05KhjbD
U26cQGKj1zqCkMG/1D9soDagl930+6PNakajQWz4ER0mfewZCz2/ebkTz/ZaxDoFg9NBNP7wTG2P
khEut59v9aBwKaalQurmWzTyjZkzf64sulQw/LaIUrpqu/ccD7hoGvi1edrX7mYgUEdRQG3oWNFp
Y0wPvYBhm8Ei2hlTYZauaSbDmXUJHCB/E3228Pa8RA58WVh22tiIeL2us7SpUx1u8H+aYrULjmNv
7+GiKLv+Op5UnlgDh/XrIzIDsLLXmUwv23iH1+siqyFzM5A0u5mpIsN0pCfB8jiFATZA+f/N2vmD
QtQA/FPU2aQXg+f68OthNV0SKPib/GeDWvN0xP88eJ73ITgo0ivo8e4oQledoRvNHW8CWP1iYyat
oU5GSbjiGopiueOu9QbQYmfacN72L9IA+LKwfS+WlPnf8sjW0tu6SIIb102mN+hv9tf1blgkRMWu
8RVEHUWOLnS10tVpPAZPoZegoHzoHMQfhiA30OZoSSkZ3+/nLkgKiYC/ke0zIofSsUMv4dBg3T2I
ZCeK216we8Vb0p5C2O/lo3DYtksKsBjccPOLQeTL1IQyX9D+7ZTYj29Ph5Ckl78iG15UwwUnOYJ0
jXbClgJR+pZlAloeuVbm+tN+ttoRPLMCsKSQ4RvYukk2yUM5n5TYKaZQnOtsa3LUV6euy/vgGyV1
+GqVaxPlvT8HnzfLHMm1IHLt7ZupyN0pvJ/LltmXrEEpO1jeJBvoIIW8mVcaf4viTIz2CdJP1tNA
0RWh8VP7qX2+m9VNUn2xdRSY+jhmGEeJPptSPZrwcw0atOV0D2eEcgdtKGsAHL2VtDAiTEI7gxB4
sD1HZ6AOJdVLd5Dhtqa94y7e0na3LyyhVHyZt2MxRK8U1VdaKnRaKTzx/iKuOmbc585QZxKyAyDv
ngG7ik2fEJtLsfkfTLsEuyUm6bClhcE+D5sV91qOUlP9NWofq+n+z5c8valrtw16HiWWJ68I77gk
CmHkJdY+e6A8NKb8+0YXxpeRwquV7S3g8zDhanTScVm2/4IOwQHKQ4fqnT6EWdxldZ6lTK34ngEo
NL5wDBQiGiAiLLazqDidSvD+i6MwrwkjcdaGbrPqDFxcdGF7ooxKSi1PTncfEbrCwUBTAwvjo0or
iRpo1NZ1uSrOOC1WPA1LJcL7V6uJeoBkqkTnTUCXdfJ/QTG6UPxwx14LPplGdCjjQVoveIgp5w0G
9EPInwoKgsJJUkUhmJxxzIqt5CiM9kRsLzk6zkfLprmt+xDqQ+kImNwGZcBhnGhr9CME6cOVze6S
1J5Rx+yzXE+hu0yDr/k4Hml1H2pgkjoGBP6TTsWZdzISjXYWhOHU/UfeA+S5CqVw9oe6elXCFHzk
fWonGkQZlcXRzfs3rRclod4b94lNLX3N75DdCycGeyybmWywMjvZ8ljlUmtQxrvhZvTSPk7zBMwJ
0dNA5Iozot6xYK1mk8deRo21/5lXvTsnViOdxoe+ek9Ds+K00pB8q9ljSlbmG2/cRiFCBTwpdm9I
kOCnH4AzVjCPV02QKj9QccxyYx1zb9BC+8piT4Y7FAhN/onjz7IlCp4cKKc6nu2vLKKivdp/kDpa
1qRLQnA4kMcifsOoFyw6UHe9LR8xOUarAh+UMPCscNjk/pnoG3LfLgIHJt47S/QpFTlNbGUT+BWa
sVsMfqvSgf2v5GNACdqO+cD6XjAXziPa3hCAml/VjbfDYaNVHNQQNwR9ed4GrMzz3k6Xbg9YeEeG
z8SvevKzdqpVQ0It6ogTm6rPhlnYNNDlgnyCCvLvdKIShE3KPWukN6ngfYvVcwPGhlGW4BFyDV80
4QhZ5unM7glnSPYcnpTQoNcWp6soN2V+asIT+Oev8TLXV/+x18EuF+odJXSXlrMWaz9IhGQmqKU5
FpsPlI9gGWzRzqy8gmrp9m7m4M2scXCQg6X6R0ygUuFM91i5Tsuviz7BYEASYAOEO/9QIHJKJZiE
QhR6oJs0xmP/MHMPgABaF6SeQVgnmI3XCVFbxB92iA2cSL55bFVVc7gURSigW6jIhh3/Liy8M1+z
GzHzA/qsRdLvHnLdmb5XMFRXau6Eh/hnr8OUT8TYTjKQCywIKg1w+TVqr+yIuA5K4nR3TZepDO5b
En3GAH6K8grPqGmbXD4I21mJcQ0RUl90Gfct0bCH9+7nNEpiEp1FxpKv1aby+gJMaLx1FxPDkLZz
yLqAXR+sS3V8pBD2cmCiPCdG+UsMgKfBVTEyVbNGnbp8xNNO5V/doYQwsZgXxwVUt3J5TGTdj+q5
AstQHK5GCis63vbh1MUMvbZ506TnTJosaZI1hqo38CJ4iuJ5x8QfkVZ8gZoxt2bOC5CP/I67jITH
1j4o/ec+obF+7nT10n3lza62BpjVX5Of4NzvqtSBaCEFBLi6WsCtpQQnddiY2pLBLf7yoD0eqgzI
zBgmXoos3MBJxF7o91aZPgVVIlLymOaKM+99Vh8ZIOUJatp+zWmjINHAVutMaf6SYmKIIRHz43wy
ncHpexRho5HOBJ+vTTD7UMxrWnOB4Of0PPsza2oJX5MMCRfhQWN+5HUBDMtOfSx7c35lkDQvNJkN
C/SgjGChwTzie8vqI1X72K5HYHkCEr2uPW2Z9Yv7o8TC14ZopZvF7FJlGlsgNzcr7+vBwG2J+icB
hGJT+IUxbbK85hOI/V6oLvuu4xZ+VFeo7XoCJR08LA6HSBDyuaC2KO2RRmOhjG53XCxJllVYuM46
p4KZwm+MUbvENABxl3A4eK91YI11UdyKkkzq+z30ZtRtmw942KzTMX7gVlAaaYkoBP9o+qPk2sHo
cg7Xq4wVrxs35/3PnPg6uJqwBFZBA4+sDfulurZWFhKLx6NW2ryjHLfknnNmbbaulBPv7oKUvIcL
alqDKWdXc2N1SPmQ5GnkP6gIPyccQNv0QqLOcHCyQ3dhbnKMo4Q+b2ZC9Bh8g2Wk2GJqBPzVLYXv
zCXlThHNZf2JTEbtsIFGz3NorsepOms905SAx92GPv/Qf1kLt/iyz0a1Elxly0TiKLBoyfo5b3oJ
EFLBy0kLmbO49Kl8emMWL+4kbiFbsJlSSrEqH/zrUNjg4y++/F+RQUH1aS0NufSEY4b/T3v6gO4W
1DICaemcsEmMle3D/K8KPLqjPz9XfshQleCvwCHLSK0lt6tBLUHj3uZ4tSh/IMgrctvDopzYeBp2
XhT5wmQ4ZuENDb/+wL5VoyBk9gvsxi4GXJNOaAUPFbPPfSB7/4B60N8j/cE+KuNiwtfExG7xC84E
zGhPIKM83AWp0jEGQe2hYAZB5H1mDWzzhfK8FqqmmvI2KmGQDWZIxlLq51WHr6mrJDvSdOa81oGM
jTyZwk7by9LTvGgXc+uXb1C9xiDqnBziK8/IuxfRFez4Zme5jFWp/Aa/5hD0QTW0DiliE+JHZ4ao
O+w8uxol5VyIArzhqVgtU6Onw1MiJZRcUZMlnHu0COoto5c4hV9bDq0Tpggfa8eoQqyx1cY7opDa
RwevLXWOgbKRDbreANxMlQHVxbPAOs/4rMattwrk9ROLE2PRM10fZFvKl7sv8aQ0tbFOucfnMa7g
m1hhYqSbNer1hpLYHCgEsdUq+Surl4nWO6UapDAp0qTFAYjMd79VIftMKhEo2XDmLBvpy1Kk2fBo
M3/dJaV5YtsgKlR+INuVGgFe+Sery3hNkdqxzg0BP6caJi185NFAtMvIOscjdo4pWE6kDGOzXv8W
dXlQLEahaIbOhEyIPOucN0TJrtgJdPuBXW4ufb4hfvd5KsIutNNQhnM3bz5hFlEUC0LgeNTWRNvG
Qr21v4agpR4aj5sTJ8jnZsIpzsqZURKhUCLBNMzXEfKSrkwoibYofz0fQyOSbw60rS6xgg3Ga9PQ
zVh9vBhGrp9sR0fJJJ0NQP6XRsXWQM30JaEeng09jXAAxIBE9tsTx61W0mc88ro+xlr2olYHepzz
xatR840b+dSK/u7lJpCCNQJv6T9CyIPdir/718rLi96sTmtgMg7bpPcKby98xvLTZoPnAIsD6G3i
bl7411YmX8seZnsajnCOuLI4EnewAA15jvCMHGhNCrTNQb3SBtkBJGViaEQkn5k7ixTFU/xvFheI
g89polvgYU66SkCiT7Yxm9M/cXklDccvuuC0dBRFeBx5eSUoH79lP0q6Edzjzps+l144uWOkOMtU
Q6gMg3JzCaKLKmOpjOkFEN73Aaa63pNlCt2jrPP3YDI/cHMm6WL4E0FfHOwieZW/RmsYyaWufnLg
1yxamj58jdb14g9NzfqR1h2CSMidRl5pFzZatR7zHLs6ZwkAOPmQnR7tBgvjBTVmeVLaQxpU7NsD
vqGH7T2P1ElhQA7KBKZkXb6DzLKTZt8oSf8SnKb0yLDhCAtvrdERRbuoX8VjY+WVnq1QHj3q8eqO
CuR3/N3YIhgwFjYd7BRttTjpd+C2UzgR1dnB10G3mXXPfyelxcf613lgTs9owyGr1pEnxtjSzc3g
1KYEfyXKgy2uK5lLSDvwCwUoHkX5I0r0Ak8At1tdP+7mL86qrq/VSodyVnWTIZcUyEAdMo/hnbZO
1A1Jdcvmchw1JhMdEjev3n74Xg0s+jXqTNTbgZ3vPLysb3RGFmnJaBsg6MuxSjQXByYqzDidmDDX
WWBx2vrDDNCkLQ8kvzN0DENb7UesgCa2NMlvIW1qwfcPobgxgusvng7tuGgSEwsM1vTtV5qw7qQP
kYF9Ac7YwD4MKYgeuzDE0T7VGnCOVPXenz3eEfBKMHJbrKyxE+2q3jqnncTNr3dAL+PwK6VqkrWI
kpeja0iT9wG4vuR7fZYbmzwxT2gRbzwJ4S+sZAkMybhMUhDe32asvvnkFDOucTMLR4+JVc0MjA+F
dW1tNNFUWWDza7DZ02eBzMuvrpuNsYcIB456ng2mYlNWt36Vzvc355CLz6fakwPLY0xDBB1BoU2V
AaqoJmPvIr3RPcZOyNi3TQtUVoE1G6ajmSlWqXMRC/tg8JKpDB0Qw0+Q3wWEWwG30bZeT4K9kBUF
HKxHcpacpU4Y6kJ9VN+9H8KvwNWQibP8GZpYlxjMq4EXmAa49CpAyr9MqSH2YaIP+XI7BEm/boFg
ZdsoknyLtgayZv/61vOpqznGGPdUbXoLgcVkd2Un8c6ejP7ul5yLckyxHsxvj0so5L0YQ5RbH5Sw
XaA+nfWxNSeVvTTqmjMV9tGerhaWzDU+FlqCtyxiiKoRlZ10SzqWLXBTw0412OsCAY7neE0Ay/YF
dLnB1j4uFu2IcSbZIig32QzciRl6bNz8cofxEbHI/bd5jZobQqyoEiDwnha+TmvkDe49lcsDzlKR
kz8tqtMYwkt3nVSJ3/gv5WzqRMIKiEP3UnvxhRL6JCN3irJ1diT+A+IXT+L6sk8cLvMsqbbqdnGL
sPYGT+EnTvej0QH9hTFAQrdqHoj6lVzycqMI0wYfJGDHo4LYx9C5+ypgLeoSDQ8+R0dp1yaIi/xL
hHWm2LB8Vs9snJh0GH3kC5T/Zsg8P3pST3zi/1a5s7W6l3d6UgNWANPNVG0dEEEQMDXrSTgCE2/b
Xv9z/8Qeo+acRaJ7ia+XRdGH2pBTX1qrh6uqMV1pN5TrZMeWTIfPVqZ3HCItvUrZDDXcRwaq5Bn8
tl8EcomIiVLlnpCG5xfobsM6coJlxy7fM9RF1tzZa8NQqrmz7DNgGMQ6D49nCzmZ/NiPdkOKAL+2
UuDzpGDOFfSAbXQCxkW635JXGN2TOUpodc2T3uFIZ/WXG7t+JPrJ2QFTddqYdbbMO/1YGT/jCNB2
/uEETM3uOPTmfmjQAv+ue/9o7J7wH0PGS1Qay9iA/3yJ2P2RjEYN4Wi9rFJDLFDw6ovegdNms6JH
cUlZP0+n/YuVJ1yW1YVIVnHQcvkptvq03MqPV38Xe1VM9x8/ACwzn3qnNrnbaDvNmhO+1hJtkPHR
//NqU58z8uznd70517OeQBtAj+t7xUf4UqRPU7dvUtpcZzcV8MIrljb35dfoeP3zdqujxayEOj1F
w9+ZCcddbm3rLGbjIAE4xXZH7v21UGxS4CjtxEW6+UKjJhQZJ1xOWmV/wnuNVFWD4Os7TPQZu37t
lXgSc6rhzfeZL7TQJPWdzqbZ4vRVSfwJSSQOM0wYrdl57n6RcNjq7aU2+JgnxUwcR6zp86tBSSyE
XTYmatsv0pXwGSsHKCUj3eMPKZdmDeOkz4QK1/9gvb74iewXy/P0ZBx4UIwjEHPK3B0ts/Yv84Kf
H2EBwDkvMocuBcCkUGBu+raQlzWCpI4YVrFmyznG52C2so0eEFgXbHyjklngOUxVrYa3AQ54UOye
6kE8cmESSb5eZfU+eJl8H9o8mMbojzD2L60KA4IIi5lNUUbGnpt5oa7iHZoeEGheoGzNeQ9UVl8l
Jq/Sj4LDgut+hu2h0oLaVECAKBrbVchXvj+qD3hNocnrJLy0ZRUDMsJkTh0vxg3g2WLyuIKnHP2f
Ez5xqoKKvxjSTUj6UK8/0N5ZCjyDBvPb2wuqFN70rMMg1mNWjReuslf9S2XzqF4bj1rVu2LNIYby
81foc0z2T4WC5YFZrLBnO2S1gVvUTqxvHWatYga9GQGPam+dwYu3nZFh7fW49XxHE2hjIVA2xxXo
piWgIMFZMYxKBUi6kqt+HAkT/Eakd/c4VRh02K9jm4oBiJ78UEsIH8y4Zk35moSkSO9ey+/UrU7B
ztrTUWl8Ioc2eGhg9Vu5qkQgPiYgw2HiYRrvRHfQ3OBYh2dJNhHQ0fTAEGewOuxWZ1Z6mmzAj1S0
ssehXya1IFfYpWj/e8ARPZR2fZ2sLAmLOGcZhZtlhdK1P4rRatcnGWKamo6nSf942ldS9/2LsER3
HsXbDW5moJ/VhBgNk9IgPyoJVXqUmL7uasoIStUaYJg5QeWm/si4gkO3ytf8rcdj8kSzxRzQ9mF0
IYy09KgxAObJ5ONoAe6frymS6Ctm4dv/lqXTyhRB1p3rz2JaOykVI4Sasg3pWL9bLpcBIEdoJqur
vVuwbsOIs95SKD4e9uVzUbHc0DI8C5KgbxEKlMTeY118QE5NaLXxSRErXcNbbiHhkKGgBHyQdCRV
xqILC4XLVNGlO1AMriffDk7zcZbuenoWZ3feO9LPS5J6WS6DmJBEdpCUDX93KLN2i3u4qPhnO1pt
G8ssIgVYj4F5nrAISUu9Q88CaXWXzGhNCGG3xof2GpOTXhYzk5tv8ejxKPkoGHDEqB//bfdg2fYs
ABd9bmf9bN/nFPqyJF/N1qfO6l/G2lxphSvWbXDcSw8O4Puy7zrhD4VAx3jLw36tbsowyVIIL7mz
kDwgQYqgQIHdiSqJZSzaHFUwlqjIqe1CMKNfc+kiOKiZqwvzR801zOEBGswFMuO3adNQsbro0Wod
IBUernNy2E5jVHSse3WKMIAH+qjZfXzDQPm5cGwsQxRWCZZWk1lm8KV7F7yElu6lf0rwoVwNpF8O
vFaphQ25EwoZfm5FPTY09m5G/OZ2pb7/h93F0mPM5uAMayAUgdhP/ut23v1GtYyVzP72cLR5sdS3
BuQalYgNFrg8kv5hUkT3Lw/yYNQ0avEl8kzr0texHFG7cn8qz/avPYfR0PsmSWUnRhQtzEWvDRi3
X2j6fYe5W5EU0TTMCa2hMj6okw09v0pXnN3hFgnfu2axVvc/AlbikYJF7RI7XMU88oAbDsRsjQbh
B3zdeBb0hm0hh+8HUnG/MEzyACRE98rLVdYwYLyPNUMIVU64jbbuFPv1v2qfHKstayIowVKAAySZ
5HEOR8V9AoiQe7pocqjvIO6pMAP6hCXcv/y8XhyaYNs4BLC7K/G+RDwM4sFe047fk3DDHyd+yqbi
H6XkLyjuF7qtW26XAuBIgkv7W9RLUlIHmQf7wp/T+gPDAi7uC2W203FkZtGPv2EQpdK5vPUq+Oi7
lE79DK0+818XntM8ekhetiHs+MzEe/+o+QiJuvE2untn+O+GOfCyDIbQQtNH+ngGRx8ZwV7bqVNE
A4obsmAXfBknNBBk8MuRXFzl91RXH+/QzGnh6HV9MXarDHj+GxgFF0nNv793DMJLJ10hsCv5LCuT
4UiUAEoxizMqVhIRJtoEmn6KMVht9pqncDs6bPbjWsXyuYqfN6a7bZpCkz2KjlauCP1R5gU4mPPU
tBC7mK1hwSOr2rX5nmNx9PeAIQMkGQk1Ah4N68hYCetBeVRZUG01CiZu5HcHl8NSBgzuoQ9VhcbB
12JDtEs3HV0SWvLoPZLpPlK0zw8E5G23ujBQPFIeCxrHu8ClbHM4Eni5XvSpBPdsMnlb51Wq7zKO
oz4thsdTXzJTAVVR9+jnM+OmtiW0OqVFn7hnhUsoLruoV4iM5fgOJjySO8CvZ87YSyzn9r86I47K
KZbZNoS7h7nv9BInLLPlypwZM4hBscL4nWUUltBxipEKd8dmvBD1KabvK1aR1L9WTv9K+pu3Wo3F
8VZFdlGy3ltMszCe4nZdQZvPgBM5B61uF2RU/5KiRbzKSGZrzNVv9PDKltf7HDD52U1VEL4o3Q33
58QrB48R9BBU6rbhOAZ1x21jk1ut0RUThdzhEYo8VVCaBael/Soxfk9dFF0n7zSuLKiaWTAC0x0k
6t2ovFt65q20yoZhVUMzFG8L6Qt3uSTFhVDxJkZXUshn9OrYc2k9gExoE8uo9jk5SZ/VW+t2x9O0
8UT7Sct9v156Mox1ybEe6CYksZOIjm9AOajx7t5wdaZJGGqmS/rdCkwjWv8dwKUC8ef/TNQC2CGA
89HZz0VUbVeu1AtpyWIfc0R7JmMRdMDSCpxVCsEjR5S3dtH98DjMJNj3gpKE3uufXaK3el/lpbEX
XcCm5UudmcHTNLRh3xGm4IJPT+ws3Om5vlAAq45Mh4Nd3gLSU+hO67f020I1FGQTGh2H/v7z/m17
fQThBT4j8X8hLfnpWIRke2K7m2LyKBfrlXjuYFz7Es8EgzLM3uPGaBPOhJQ2CrzLKccf1xgkeEXH
pYDpv5SEfvtOarJuOrkK6rQPe5y48uW4Kou9j6UVZfLLSXM9yS7ehAjthH2EZndhzS7LpnF7JCRn
fck05D2K46RC0FCXqfqH3Nd3Y+EDk+4JgyYQuWQcYA0j46uYqZEAtf/NQ/pNfEljhSZ9bQLTEjnK
BYPtT5oPCtMuTuHLjqQ68fRwe2G6K2iH+UtFAndA4rAexmbTmYTh/DBoCEn9jUXmW8Ang2ZFRqsv
f2OBsvcW9d6R6WzqM3zIuAa6EApdAukvQanHeDZQdAFEgGG+nv3e2IbVc+2kpsmIB9kr6ZTC7m+B
/57XcIfWV/m6kJMNmB979JPXXEtbsg0Ck6YTYuZlJIdaZzPf4QkW4Ni1BPOZeoDl6vOA5F1ojKdr
Aj5L7+DIjxoysUqwGIJ9a+94Rr9gSC1LRLkdliYMuAtpX62JQEkN7ukvuG35DaBaw/Fi3vl9nShx
cBIwvWWckidnPDDPLRxqmUvJm1t4bSyX+HCbkS6ZSboqCyLOw877QxjMjqUnRoEhWXtMVU1sMeSd
8dxh02iBUweJZvqnavVRgEtP37BRatMhBL54Synhfr7TIl+cVljQ9IXlHdjGgS9FQnev8hrdA8PA
90Zbnd6lyIttGZQeZhfim59vH5m1eXghbjjZEXVC32c+SDXeVLiC3Ti5tpYErhrnw0f2OoeNfKD1
10w6KM9LAz+fV5p7ef+6h79IR8KMTrrsa8wz8aBtmCGgR9feLhS7qMlTkuvnIjyQC4186cE07MTx
XL2UVtVoke96Ctoj9GGoCKCyCmW39Ff9syjGH9b2EOY7C6bUEZYKtzJZO/yuq1DM7wo20JDIe+Gn
PF/cBfbdDD8/zEl83chNImWiWpOLMR1xgY1umryEfmuKfQBHloVK4QUCWs/LAmLsVCFY/at8/1mf
qX/FpSFzUcGFj0ruqnNIbmLiqtzj+a3xc+uOn1PvSwzkMftUk+qex+i88f00Qo9Ja2rBn2g1YyZC
2/pdA0xSAEaPBatcK1232QxZtm7i6zefJ11Ge7QHdsQgVJ9+SwEU7vHV/EnA/pmKVov50EjVFd88
Q6TjeLHPA3QcC+fe7E5fAcZLEXWQWtUsbivtlG+fwZ+cQn397Lv+XwancU7o5Z7dj8/8owWv4+tu
8g2xuVzjfwVo5yeKmx/7OY3TRdPP73bDW6s8Nwy+ww4K6M38ayZ9UpIdZGyzCldslB0rt4SJenN7
QBKwX7KukVFypd+IEU/Ay3eVCo/Luz+mQ9XwBEbWC/+1wRfZl/LThoAYNt8QNhisXZR7TAvAsW+q
cU13wzVfIYdI70oAQ81b1GtDq0CsGQj0R0oLDQ5IMpYo6Xs0Oud3xI8K3OEXE9DE8jSp2zWBYRnZ
QCGkRpdvls/KIm8Y5nQoSbSdO1BbxQvCLM8etZEpDPuidE3lIrneKFSwn61tlyMl/zz8M1sBkpcU
qeZ0PZ7p4lkidesjka+au2hvml/oI47Lf3C3GcqoO0HBMx8Wc8U312TPiXdig7Rk8l7OysM75JQJ
UG8zvWyA91B3WftmdHSaQGCo3B9uW/Y3Cm/GptXlD1rJs7EAgSC2dm51R1WY0wp6tnIZHp4tU9lx
sZTu8q7V36Yds8ZM4S3slKb5iUkBfKSCUS5aiPvZc0XEjIKCnlKamSBDPcA7UVRAulTxPwS/jEZU
5hPmGIz642/BeyWn13DuXcIdU336u02U8GXG0ticuM0OykJLjNuEIA+rkHDwVC3p8u5EPFfk7FrR
C6zvIUzJ/Cdu4l+9he1ASUQQH4AfW4RnkGHfk1YPN3OfVWpGHtB9YLifN536WaFXrzs2dCHEuZuq
3qDDPdqQ4mPtyYQ8k7ZF2dj6ltwgHRRjpPrrdPZwwESMnylM88vsoRkvRmtHWLaNSj3PcsNDClbk
PW8gR5eUERASZKqBxQp54sBam4w6ge8WjJ193A+ybLWPTlkDLduOjEE4evMKmDDtLZzPj8LaDOqe
ClkMktWRazPf5M2zlFiJx+6+r7KnUfvW9beFhop67bqnbe+q/6D8x1a0lzuhxjTG0IbjVguqFZIQ
JNG7v43s4XCdiTmP4mbMozJ1bDaJt3exxzOs67pUqGw6RDKKRZaWnWIIO0ZsI3sKRwUdBUac/FPY
Ad+JtSw4Te8WoFxcA0PUKXu01sCsPI4l1eePdmGZzBae6l8mwm7/iVnSz23hMmtKvqrVciI2xf9R
y6LAirWDqOMfumi5UbfQwgCT/f2NgHx2HRKSwOrZuSERgOAKiq8vwru77DSGEX6fFuR1M22tL7VW
rpOodxq/1AR+T51a1BV+Mx14I51ckD3JKd/gg1Fe6N2O1xGfIWPOxdQPImWpmNq4HxkTXMdbE9cf
v4v20rMNsr32f1iXgPlVF4e+MmaQDP1bEHHmc4iIaSc4erDJxrEkiG2W4XULmgtaAeUc3aOO6XJl
6ee9lnMASMWzD0zG6nk6ZNqH8xRg9UUNVfbmzwhoD4kQYOuIJPq5Rk9lp3/CCBBu4dfkUuTwkaaS
y3wZ/TsvcmWzQeAOBToptOLLZhH75Dw655JuXljf+TZCjfVvw36pmkM/egTqd6oMkCued2/7z/r3
OowwwvQ0N1XP3ppGRqjqEmp5RnYXGTQKvjfkB8vfxYkMU6m/gOwhmjVgmG5VSZ+C7FcIkxU18Cf9
1ZIusaXgXtl5fqcOLJLR9hSb+JMWTzxTM3INU7RX9O8Tk5DcqkE3p7vyT7D23tOWpwZdNV6FFAx4
VIfarnUD1fq7XqEQjoJRpm+s8hlfQRwY5eS32QXtycsY1vty0yWuua7GvQ2VzJwf12ysG01dhncY
yn3zDKdyIoX+LMVduhITE2n6CdMoDeWztZwzl9KXq48xZgW/mB6afDd9c64ppCa5vJ9IGBkNzQDq
L11efxUuTD0VzWt8M/cjzaihpwPC7xKYhRx07B4w0YRbLc9a/swOJwUoNvZh7K567PqkyGHc3Mwt
5bFx6dXlNEFNI+N02FwMDAbHkoqr0xQv7zn2fdPfH5hlmRhcd0z3r5VuayUoBz3ciktoFvtJpdXO
d2WHdtZN/Rz8rOHKs5Ie+lJbjyvp+9QLYWBYNTbTWRBnb4Dvo0TUj8I9DDf3lBPwJK1SaH2uPPYQ
PEpdSufZ4NRmdZE+6HeX3S5QPUq+abd7EcOt05G3//Pg3GMq7fr4b7QslL+ImAZ9S9pOgTOaU4+E
gO82ELNmtWhhFaEPpL66FCKvLOBsBY9ZUriCC724RryBdac4qnvmNlS9XUMl+AglXDbdq6SibJCB
5hd2AY934ongUsBr77M2GmW0t301nzOExEDVMWVXxGIf0zd6f2kCsPfSl+7ISGyhsx6/kUvRDxmi
bqiHSbRhkftDfSFvQYyW+SckTd4PUzN7voKIIV9EPRAk6S1rwJHaUwJ+ryjcnKp06HqULn1f6rhT
Yu0+1W8dbnaXVssOyN7NrgQFGC9J0YDcfP0IfXyG8ER3hLMko37s5yYkofGv9mQpwQY2MGG8idkK
F5ZcV1qXDO5NHXcaNFbOpVCgH6h/+L3LfQ2NDllSll9Lovor1j9q/dk9ogUNF/bZQXiCLtgq9ft8
tXsgLoDmPCqExCPRh16v2YhMPqIsXiEm8iDIr87/U2f5pryjCADWtm+ffJjD90QxzAHCSNPX2ocE
w0B2KFghHmqPMlBU6GgRGTyc6IXNdltcTJe1U12lK+YVXP3mL4syTM/ISe5az+DqQMM42PZF/lJq
e6BMgr3t7JE3HGqxDgdn1CrstRKOIfKtxxP8V3YLFWBkk3clEUHwKixx1O9dgq62W8FIqMpUP31h
lBAJtNkUCQ6hRbzbCCbhV3358SRaDLRmryD8eyTidClSSLhM4+54SNwQWpfnc/2mC9B/AldAvSFt
5JIbQ6+bTJmL7XQ9QK9LCo1CWTLObS1rTQRpWLcH/98uQwalhkyC9InbyrKAZIWVt6UrW9M4E36p
hf6Mu9jASDGkoPwOB96NkJUqaRdOFQyhtjVjuy0kS/Tyzb9nSSVOieXCIn+bArqaVi8FN77fTOGv
EOIFfXtGnUISvmyl5lpZqBYVesj4Gg96eB58iAey7xJnA+qyw5+IynnCRfOlzKn6pX2tKJo+TbQF
NjD8/15rQkSyMToI3fDiWkyvdRBtVCQubsLhVp0JaqbRDIBfOp90BBX00rVIeLY5xfeepee5uOy3
CJ93bUoad6V/xWt8nSPfM8+0dxDdoUznIz4N1cJu3h3MTYUff9ggEazeISMWhPzMCTI/vkUWhJgc
TtI34XH+mxnn+v7orLTWbPRZ/T0JtzzbwUPda9+WOfqftIK6nJqbsrhUF6LKx7DOlONdR8/XUsdj
eYiVdLT+wl6zjkmBj6HaZhS3yWCmTrCzbR93GWP/Ghg6LtfCpVY+sOcMcq5xMeJX550r9vEhTtL9
AchoUjouvnCW+NT+fiKbzPSFZhFQMuCDUJxjjPJGwQuNjFD0+09fcF7iH0jAfRZ6zoQsvdUDRGiP
A7bUATk8y7/ly3MiHZgSRtcd2L5QlhYXwnpylXqApkxob+KfNLUVbJW5ZskU6+M2G3BjWY7+dv34
3FESaPX6njLeyFpUIkhixYKJWacfRm4z+fFxw3G5dX5mq06D7s6Bej3nPDSvs9W9N8vnpWrKI49L
w9R9eQ2bzWTjxlGF2qE/WjWh2QwvekvsGmGVzomUTXzMKpTyQMJrjsSzdPdPvrQGdeKfzy3ZFrpR
0C/KgzVeTGNsvx4FcxbXywxE2UacH6cK6qGDwtlCjh9zOD0g6fRlplwyf+G3IEYZDtKRmB790NM+
nemoRwaBGpCPELNj24gsjJWqH2o9xprrOb7IZblkvu3TLIEPswkHZgB3JC+XdG+aPLRzeMhfCk1m
3aKANSus+qMwNztWsoXuXzli8QzUBf4RaVSZVCN6la2yNnBFTPJYhFD7YxnIbRqK+EgaNE2xlrPx
pWkKkjFB8WJFFlWpMtUAGUzL2UzEZ3YIyA4C0GBdcPXG1qYpuMuqH1A51NMEaaky327OSoR0QdQn
PSQdp4ETws7gdEnIcPbSdnqp0lhULGCUKqgU4dA6S5XBzrGQK8EkvXSznaeRuOpGJI4YkacmZDCk
xNLRbLLQxIZqddT8LZuzQinDbqKEBvR1GGDic9XZdng50J8tXx0nYtlpdlAi2F0G7l4yByGoDeHN
WAh36+ReCS4acT4GNHuwo/dJszs8fsBcHwkBem7bVY1ZLdThbfXZ6rAXUZYjj71vasi56RL7pHgq
1Z6QYZfqjgyhXHFlbE/Qyx36KY6VMRRRH42Grjb8JUvbsWkiDSdbEqhDmjH7zRv4H+B7pyVnw7tX
1ZhMhMPAcBImdiDLh/MQDkIMNqr5D/jHNZYw/7Znb/xvNS3ude66UmvTU9NF4SSWMczNiOSmwS3h
lF70EByIwrn+/TXhGNDFlyPxCEYvGtAi6m7XSJqO71NCbU5XW0U8b6dOAPeAw1gcFEzB3iUEavvy
Jhfv3dHEbFTbczFFM/Rdm4fPTn5fumxoGLu79dr0n6HRIvh3ZteLGOEgN3eln5DGGoqmh70jhW/M
0FEbcSC9YSYXMctMu1DVC375/aWn1NhJF7FobUpvOAMDLr1eWWftY5GnyL3L4iKCKQgXU+ie41AU
1Pli6x7MPrP4OfVfpK8qebexb0luI8CbtrdADXDomuieYKyNe9raRSZ1TjxmNgnmiqlP//Tk2Hpz
AaJFty2/C6Z430Ik7xvOiAStW/a+Z0JQrSQLO0mEpfs62tSXeLnb6zOVq8vcs+jW3d17LgweEFJD
szyy6CWcNwkxe16hzc8s7jmmKvXd1ws9HJYlW7kZpOlUQqR8RrmfseFnX9cjANOlSv7hArHb8YGj
lLF6DaRzOH49fFM7zqFY+5THtNg1C4E4P02qk1ruIjKyxtQIxArmqhDOUU09eyvfUU5dmv5fM8tL
9CDdqLF5fEcHjfX1CzdvMTnCxSa+ehblTnEffER+hYUQlVcGqVNOEFoFDN32WEV6jgPxcCOMC3au
VKaoe7n470ODGb6UWuQ9JnkXkg2aI04l0vHdX1Ihsot2w4Xg4yQno5QVXhV+Mug/+7ouUw2sCBdZ
0kHq17VdjKLns2uOBPXiH9gdVMudcIiwwuQQ20G2wrnb89fjbNI8jivhIhDXEhQ/l+HLdQUmge/H
H7aVN6z5RNc8PhMJAXsQWZvhZDPrYTfjc/WBniHv//dBR6OQfDyk7vEFRws+R7AXCmdE53V7ebdL
HPTE7Zbnh8u46AnGKFrUB4suefSJ8GbD6uELNp/taBxmVytQBUwKdjGFOOw8Nv0nhfDlXbbINWHC
nOgsSYm1GEfO6t6kcIojMHv9NtF32uUWOSA50oqgAOnL+yRyya79sbUwMczIxC8vocS+Btn2YcvD
Ah2dJ/6MtUX40FquBo1bAPXm7F+66roDuknSPoRKio8dZIY9Qb8n5kFwfANQVFs8J0iQjfVCwmAe
yNqYbGjFWbKut0VvJ8tpMTmaTQYBe6tCdXOWEG+VFU0mcNPLDTfdMnltInhrHQLfNc45bVH0GVMS
ErTI7jmkyEjb2ANF+Sj471Me60ROxCWbvByB4l1FJsN/SxfDyS1CraXPd5FqI47wMPlUnmPK42n+
omH9R4U1Ft104rH5Zh0veJjFyrFG5YxUmbo0QjX2YfULySDi11lhNFmXzs+kYa2Jknj+L2MWCmgN
xZInjNzhF4N6IHSIaUox3Hl2j1BNu1dBpzxiaRru8rWa6QI2xtuAnCD7Dh1FE1duqU5EFyD7ShVk
+RdlokrHs+qWnByqyNYDm6arxWmYWhsn+xx15jvfCq0NP7HuPoNnFwzjj+N6DxP4htE7KOTSzHvC
DW6C25jzt7rksXEHFgPaO78N2m67EzIkk6Q9SouyXItT24QzDoQAAkLtj67s0n9kHrPCQ5bZ/cmY
s0wkO2b+YdmhCWuO397BwsFNn641zDoalkeNTZpcPCUDw7Q0MaO9wRZpy7BCdEVWkyX1MUVj1tXM
dv6kJJcifS+WBpejky69tmYKZ9eah6Ex8uqPIycVomw40xxRWQTxhb3Xdhsx79rP5f5bBO8m+oLZ
6U7loywd1rIOVaD9X315ePavHACXyvxfd3+jaJar7lYmwddK81amf8+mjZdoElRblQHoVmF+BlqP
uv21zzc130aMgC84fCIbUI8NYi1XvA8MPw9Cikw5cbHzUDxdT6Xnj+URP8NhBpvy4DacuIPXfCwD
WXswICuwKNBm5HrbJNEVCnwBcKe64triEYnJsSMkEHI9+kgTnCIXu9RCtsBJL1vfOH/NZhLzakBx
tpbrLSUizoGxsF6kkzOs4JuZYtSPPkVNLql3AU0EtIC3JGtun1aOuUuUOqvwyb4J9DTHPdM7PzvV
ypZIlvtphmyxb/JJG5xNokpRHCOlkt9Y/H2n9o6ejDHS3uEEqWFR8CYaNi97CVc6ojDmjOvZgL5H
Tyu5fY/D1QBB+H40FeqrIShRfMi05z7YkCL/Bd8HUzijNMz/8hYDm4SPvYhy45HMoPGcIuY98h1m
IVlooMQmk9H4nZdfuS2UjKOyOXqzWJoFQYQOo4gyGGZjAFuFUDksPmOyeSZRw8qjG9ep8poYMfQ9
uApb4li2PsS0OWoETEkkNi2JaPJO/mZeBjClsRTW/gAEqG0Sfs+NFM8ZJ9DVZ6ljt7glgWr2hTOv
C8Sgo9LOgxDnQDJ6onsAocuslbNABvGK0jqzjrv2rMAEmohenN9VZTP8u7gJdpZFntsByAD9uYgV
Xe0zspGlyLLDLSylROaMILZYri1W5j2TVvQJH26ubqIwS30d5JcdF0YqUR3M+dIu98ueRO+yDHC3
eTzaen+iieVj3pzgpznan3KO8z3tBgASJ3krJAhRrLAMEy2wd6g2Isy/c5HrXR3yXDMeC9cdWh7p
OO47LdJw+lYhpeAP/MksCokaGa70ohnZzzzMMzNQd1Mv/PeouDksgtCUTUFzpdWzQDHw2kWJM0PJ
seocF4GuH5eZyzPkQq6JTHEUA3GC9G1hNPrhuz80A+NdEDr4EQg/Ntnlfwgjd0uKqmAFMcWTXhHa
Nwh/8NO6Ina4P7cNWVNloFBRjkF4Yj3PQEIZB7znbSuPkJBkbLO+8vfi3ONoXiqeloH+v8Jm3lqK
Ftkh5nxFCrDn+YURpU4yjqP5yZqGoBFvpFY0UaVH9T3SCRUbWo3jx4EOpcPbSododK8Sfm1j+NUF
BxxdUnah/PvnkKKVShGKzOWZE6RLsr6mVT9FS+tQDZ9hA7IUQ/aKvhJ+lSXbDfaCF/C3IZQ18heS
LKsI0+Db98AiB+rz1mCKy0BdzF4vz/9v14jGUGRZmmlysVSZh8XdhnVE6xADGqO5hcIsYreglnqA
WvQuDi/aF3p1w6WVBGIWYVwkgTWmR7pfApUbKPVLqEe5tOYdcCOXB3D8xmaznw77ydUL+VQ6kNrH
K3G9W8BLoT+IeOfyGYxHU3H0y7Z4YCyPIad866bqfDrP2BDIoXJQzXjxACkmaEf9Vlx/23DXEI1A
aRuqXdFNUGXClUeb09t74s4USgsYHJht+Mpxl3nkdZfNfFV0ZHi90AFdZfy9/auQ6LyYRoBUoViT
gVzuGW6yDIzavjUu71qdCbKo5FD7Qtz/wYOfLGjpQSqpN2ogHFR6hEhEThgN1pC9JbloVUezXuq6
afd+azsNDa2XbwTVhTGk2O4zbtoTkVtklJDPBLq+GhDBHZS6+IRJEo+7xJ97bg6zF4FFHBmWn0OU
IjoTQ1+lqr0CwUsKn2Jg1E9IK2i6Mz4v27lpge8m8VPqi7uW/O7mUgznLW/LGESHDRAMukFliy9p
deadKoto5icWQz1Na2Q0bED3WUkNiPb/c3PjRyJyhmVimSKPCx1cflarpDZpXelWbrbtPPjjBCXY
k955stRjAgO5jbOex1p7fZXpoluGLIpZxGDNUZiI39qBO0FLEvKKhOjwFNauNTfchCmDQQStYOA6
vRzi/oxzyTStPbmFq9Nv3gqZVUma1g0xDUIt/bPzpNyWMhULSabGRNPo2cOPTR5IYD4IqIf7xi/y
VevkCbOKo8abYBUojoq79qLfTafWSLR+Vpb8KNex991uMjZtPO/52yztTKGlXcq8v7uSd2qfeIg2
pYcfEJr402bvomiwmaiZVeIH0ZezAtUPOqCliuKxL74KFx06L9ojgbVAi0BDsPWLsg/4j2zMAMC1
DIlYQtnTGhPmVAi7s1MCxULOVqwNb8eLikqPfsa608SX5dGgrARJj26hMLywLEmCRugLjR4XXkeT
DgfYV2UY0ZIYEam6cTkQ1BDKDP6c4g/dbH5KasRGO5NVpnyL3WJEsXufVNcaQVnjREjkR3shM2ko
V7LZqm1co+1Epx01QQ0gVFZQDusskc0NFT/Cv8tslbffOzSm5A++b6w8f+DWGnYxQpZDfK5EjAAV
A/p8DI/REZsxxxChBzphHghIooFvGxjhB2pWp0UioHRfXVjCkW0fyOMpzJg50FO/wDnBhYq+zM8F
nv5tVKBfmlg32M3+8jjXPVD7WrCLkGu6PAE34Ke+r6ZiXoQtF2XKlczoUKGJVGOhn2kTtLAASRob
OaMVeV+mglHsymGLwcKwksTWrhxRE+6lTSLZnN0kng5AVtodYcFu0xeOyn3pNR7OudofNKr6hL0G
uuZt0PjXv30XYhF02e6KQYbdk+xZ97ne1TwTlyzMBcGM96IYn0oZPt4CUPaY7mt20lgY9H/eWB0h
sbNIISdm2DaitV4OfGcSnxFFxjzUvwmEEO/vtEwZvRlebLxP2GBiKd22IBeN2gylodHoqi8vDMse
aVVTsWhQWGe2qUlerN53LaWul9yNmtUlg6Sr10IZ4ku7IjI++nOWnyGODorCbxMiiW/6oBpg+okE
98+OLl35tExPN+UKLwT5DkcYPK+LB2zkAyRo/4Y+XxJB+k5q1DRqUSSQWJQh2LfmXd9KOSyYm+qR
qphGLYTdWgmJKZKCClbXSCy5HI9hEXZcgcD4XY3GDMhnTJ4XYFJcGByv6r63RPHPWWH5lbSRlajH
TmTU9IH6yemO3Ot9coX+gmzOF9g3EWeeMF67XHPOq7cyMpNsrqXYG9K1d6IPJT/s7LZOSllPiTV1
vP2kiHbbrFpd7uPk2LCGH6yb/3J+unBNSuJCklY+XP59KG47kiZ845+1qgqVnjMLddb2AaE+yfNs
CypLcBTVa5xDsB1r+hsEsLvI8NwWLX08vOtVLFX7Vx55h7+TXTsrKh3mos1eN7eXHXEA9/TCOgev
D2bcJb5FbS/Tl4EfS2AS5vozRwiU9mY/rMPCoVr6WGD3LYvFg1jQ2qUQgl2b0LGDpWAme0PvtE2A
HPc7pQt2dS9t1v2CylwDXwFRMb+Mzf6zLwv+sJ2O3iReGlEMXyj5mstYzLRV5C57eU61aDB2Ic8i
gHx2DV5KQ9QMeiWXj5cj4jvhbCAsYhEeTXP7Q3z6QyMpx2rM83P3vaQweUOGupFKhftLSdKhh2pU
Utv23fsDE02JXvKmNth6CuweS4f08t0bfAu5A5dJ8eOL0SVJmqaGDSk5um52H8EbxhXQ7l8rGJt2
dubFyHDuRnTP/7K2wzjlfqDkdk1m198YdwjMyH28Zj3sjDjzsadf9br8HzpFwPcYDMU9UzFzIiU6
YswCR5FMT7EnLgB/XEk1GNURX7mmxShClH09pOTw9lgNTbD+5X44GfrhDxmDE7yy8sw1COySGNNA
WkEliRcvjAoKZRSQzrG3tM9PBirRmkslzjXpxlD2c+2gbiFeqbxqSjf3LU6xR8TdWyi78+VvI5gq
BQV5VRn8gaVKNL/pV8PQ0GUJOqm+0zVoWAnsqKqon6PJT518C8Di9KJh+vdRvi2HSdYc5+KEn7sP
jBFgnk7rwCaSMSwqBFKQW58mywrVQibd65bss9MFB0+utILI72az/gxSUcz0Z0bbIhrH43MbMGYc
Tm9hXGA+6F7uiEQjNYJBAoI25Hb2OPglbbOF3fGnWIPMC74ONWlC9eXOV22Sy4bzcyhhDYMyAS2I
X8i/DTXhR+j/Cpiz2IuDousyas2ZZEQteqfa4ugUFK9aao8dLIIM52uyZD9dAERVjvmZsX8KUUfR
7u2M4wGTEsxB3BXPfn84iHnCscvvPn9vfhVskp5jOtVhdjVwBg0Ld2xVs6pBavBrqa7O6nsPO2O2
Xgk0ToBmT1mBm7RB9JoeeJQ3XjfgSZVTtpPtL/53QFQRGGjQC1Yb8TVtCHxbPSsi0L6E6gKuHkpN
Tj6UTl3pFmnvRzEmbupynQ0aXryy3VJPUPjfelMqZ0uuL3uHiLiQbrGGUnPd23rOC/LLjHlOh+A1
iXyOptjIB9GN4jXALPJHwRHUZt4I5pKK1inJAZY6u1/HdLENW1yQZfbROZCUZ06d4XBSofUgvqsk
gd27O5+in+BQYzB740Sc6dZs7EuslyuYByb0NKg6+t+pGmwm0F1j+L5qS4MVjIFbAAWu27Jhjr2T
znvO58G3ylkDDlJqRT9Jr8PSYchZ3s9R9lHruloquujBCMU5leFx4C9mGgpYpqBOOETyltXBbcy4
AFmbB9UBMqgGlPO2UWmW5Ln8rdU836owxyku6uTPHzNrL4hnTzj8A8kDRbL59iaL7lDjGYNlqNiw
ZhOVuEaQCjS4u8X/OXgkahhfKOsbXacfp4pLJhklkiK2Z6NZjR+IWAjsmXV5dTyWQuCrpePHTL5Y
jrYcvKQ7JXrHTZiP2r9/1u41s8Plmv6c5G37rAFSUMh17/22be4Pr15VFRyo0dvled+NYXrALQZm
VDQRN2Pw0Ji9Nrqy6EHYYLez5/SddbpfBqwU48Y5Oyn4Q44SdYuN88s5W4V8x4aa27Elmqa6FDx2
xw227L6wLBldUkvAnvagQJwpIYl/6E2mqip0uTSDglHn57J4eblv8/SoNQg2OYfqgr+9riIN1NwZ
y4Dd67QHCGRbMMXdx0I2iazw9Vm/RQ2tarHOYDDfJva+TiXYpXyGLz1hh6bCyWCX9hYG+BlCVkXe
EHA3A8ADLfcIz6/KExAWKGRYRNw4p8O++5/uje6rj/K82aFr3JEKqh/HSwvrTrAB+IukYXpLXdMb
vOR2Kz3WTf6JNFi6kCblSDPiQhshVl61c2vXBG+6WjkzwGl1ZESY6viPh6nv3WjVGEIFTKSKfBXb
+eG93yVm2iD4W7wCF9m9Oy71qRzFQyVz9p0KMLBX3T9j4XNiduFtgPhv17CxPYond42C8j/Y265J
Ww/DbC0YTlWJvTPsRTDqAGSahnxetXhNYD4zvExSRX/3PL4ls67GnHhfU8/cDtDzS245HsLoPPOV
4bmO4ErZdgOZU8yMOlUFxz6xtdazocsRXYB26+6iUjgl+dL8wVQB6YOvDgiQQSPYjqD1vT0O4TL6
4n1VGgZDUxB4IWqWRdtc2e72PUSSxmt0W86KxuL+zKEq/tk5G8G/V0sJFCJt25Gq89YxaJdHTsIT
/aHZDdomb76xh/qnrzSyh2fFbTo9Lxi+qHL3HCnPgmeToMpZPjiP8kWl4ucHbbmE5lwf9Jo5tm8Y
4Tunhw1ZP0qHKmgU/hqb6D0ws8i5er/HmOqK3afwyM5CzLYrk94fHpVh6kjBaKq394TtFEIOOkOF
A849WYGOxSdnsL1Vlnl4hTBcFYdbcFVQWjCpJB3hunJoEL3k8pqvag0qpcrFEXQtXvL4si6ccOW2
wJIm5AMLhpbrlk+Ojx6mvKK5pHRR6zuvfwqATB6XR9VeMUdwujWV+oT77QG6htifpBK4omLni/GI
eq9+oO5si0DvtsqUMINx5r7GI6EC88WoKie1mwcBJ2xkk3imMxctZ3NQfvDgHaODmwSXFXPbiKC1
QIxrcdMoLCmG8HqQ0OJYzdM1eCK4T/N2FpZQaFvO1NrxCuWCBXpwVHo0ub7Foa2pb+QXFg29A18b
NheIBxQzYtYbaE9Fc3ajt5MYpNXu8Hk3ZgYZSAqBlcxLqO5V4AM6a1qC4jRFUTEoALysLpp4VBYr
J7D5dkLiUatdJfXSrWLMryH8kdiR9Oss1BhtPID/nzFLxuU6pJ5A3Hoq2Jwu3CavBUGVhR4wPGsj
gqa+qqFRmrigFs7ywoI6gcxjFK0cxKNBS+OF7UwMfGcbYI+7ckiFboRcLW0XBvv7cuGfu9+0zdo+
KrujuNPesyS2++IJu0rGaza3/PCDAjyWPPxv+NG4VYTcOsKgkCzrdOZywhQQyNDdtoUjKuluMITk
fiV/Xd3vrCFsLborL6EaqfX7L/TGeRbWrIsYWs7BjyO2iAmJlBL8zoNonYWB22SryS0EqOdqFkvc
D1p80Oi1ciRcSY4lTtRBx9Qz9N/WM8fV4LtLMCm2tryrm40/1CfXhzN1ZVIlM0CqGcOrNUeopnOQ
FozRjkjpUyAC3GC3u2QLgia5fv1QZEvgxSrV0VLZ1ee6tqUBAB+e9Ujq+sBll8UNB9BYZxuYj9bz
l4tMzoWB9CYRVzNlAACEbIK2iCNWBpCHdvyCShEvW/nnMqFAtN/d2JnzZerLMkY2GEF9HkO+6RF1
DKGiJ3SXVTa4IH9NSvPFuttKb4P0UpaVStnrIuIWCKszBx+23YfPvjverPIMgn5V/2nL7lHFqkil
OepVgOuylKw9bd/ZnCgab3354QEEqGnaQ8E57Q9Nm6kkB1C3BxykmQVxVsOz5knw34YRk91pO+7H
5b81Gy4j/ukSe6cFo558JSq0ypAVpcfXeyLRVmE4bde361M1Y6ShWFfJafySBOugZPjO6VjYAceL
slzz3oHeD6KhK6CbwwkoXrQULms9cEB1yH0vCfnb/l0JtM7DzvD8yY2JoxebsmCe+lJ4w+MKFqxX
syUYTmaQMzjP2pvLVhtL1e1j1kbWK8kMWkMMr6S6QAs+iNnDNNDU2k9MZ96cNs+eiJupdHAakN1c
sBQ5bVMQZJdfCd4PZxawKNf4geX17YjUlTeyNaqdQbMtuTpea1jr0Y2Y9x/We+MaOwv4RXjlJgwW
x2IQkYQyno55vdJRMWE+Yv3VIxCylKCbnlFbRAw0EF3vOOkMtuEoVTal7UBTHWQiK4nCrEv9yuIW
GyFYFSQ1K+n1EiKYtrZBRvmdKQgclxNH0E0HYxEMMpwUYq6tm5Np2vVbF2v/UGWRXuS2ucXLW6Uj
MmRsRHNPq5+oCBz55hdhAAY5V7HSyPq1QCi2ZGs8hPWw4VmKHKWrCwbwJE0hJgvJLw2xkY+5X1mt
y+iL8BVrq9pCOrjjl+TLciAzCmVRV6Npo3dldUl8Z6L5k8RXDqHG7FcrQsfFE7E7ADY0Nj1timVk
aLuDVgdqd6ZiKNaCqNPVclzqhCCTfYQuHJCGysw6kfZwfTDgs025rVrzz1zxBOJVc9PgfDRvYiH3
xc0+JtNthwOxhJpWqVn+3fr31+1teNPjzixPli3Ox0uBhj5cocgQAUBFGzn9RbTItP+/We/OrZz+
FTj16nqdSba+5Y8AURBr7t2sihtc92l9p47xkvSMAIe0Sfbr8C8IyTmuOCxmXFmuDQ7PQzdyqA1O
RsHURrMbWz9pD6n7be5goLhGlmh/SwHt//SspfE47zAwSO3GPZKf5kizvss38wT9jt2TzWU3N4+v
LEXlajsQLmPwFb3/kNJuuKBVJWPFxo6JiWJrDK024htgA1t4NzpM/AGpKOufYXH/6Mr4v9JOp5Cb
uUjlX3CKakOj9iJ6ixOzoAYwhjv502ksTm+DlNhKVRcPydU2PlGfKYBPux8CDYiGmc458Nb86H/d
U+aLBya+c6NoM04p/Tqm3U0a3ZZZctjR1d5EqYAVR8UM36fFUdJnAKIm47B7f4hxXVDhRUbLG852
v159ETyF6085YqdG1SYDXPO9Wl6afdPhfsj48j6aixMuDVl6Nq3l/FLkX7CtyDHD1LDxAMbSWLaa
5etALDZx0pHIHd7SILdzSMaJA76lC8VxxrIqY3o0N3BRHfa8Hw2q8UYWXyDLho4U4orC8plqGQw0
Tgvnw/rIxmpo7w3Nl3TylTFaRhJH9dk7h16cvGl/Yj9xSJ7BXsRbxgxNbekxkMZ/43cABUtaQWSU
LOeyj2c882TwvS2J/Mp99wwIaFreL3H/sIqJR5JShuvMn+ziVJSW+1B38eaoIZjc/Q5ZZQ5gyd+T
4KG/iBm38wduydWFcKjN5IFnj+vNwjsWW+unbbbA/hS6MaaAbJuluyQFC9qz+ZcdpV0U4sbtmKgY
b1M27JvI5WJKPGmxAwSo011PFchqgmWloxv8lMGtI1V2NALTckCPZrV5QywgL25QmESTzKTf6wJm
HN7L39+aHBs0hTI8R3+kYtjj/uON7id116Kx0SZhfufRpnqRcj7y0yMEf+fzY6L8k6cC3ZVmVJ4d
cTsH8L2sDVzDyzJFqi9QkF/In6TMINfn14yoL/8FvNbxC/UTiBE61Amm5z7zv799TIryic/NbmEW
CGHG4OLM1WY9fQ6UipIR0MeL/SbNGp1QZ/7MWD+gioD4GBmjo7vt3UqJB3uzH9/3O4ZRJ/LMIyqO
yYjPpNUd748CR2eCSZdE5KHdLbLrDoIwDQwZm1xsieCDQJzDrUQ5TXyg5rqf6JVsLPQ4sH/dUK9B
FTL1h7qKbn2MmbJYzPMGCBPUdgpj5Ew2++IYzh6CCXlAXEtKz9rscKcAOMvxB44rbxOdSHTUM3Gz
A9nkDI7KIcbYzoTqV78Iu2TZMETolEs55g6DP4QHzVk3XwJlnR6P/r/dQP2PJUpjg/Q8JB8/Lk7O
kNVbfcNK9Hpds/hwoRaAwlSSt+I4rICeMW0FJXPsYs6LXv5iYwwxbGn5Y5TU/PTNeGQrU+/m2zAZ
g8fO+nsz9yXQTQgHVSaZ6IKHQ6XuBpItAoqXJtRAPVCisxMQtouEztsZfxgvKPJPyxR9mL63kVU0
kxIj6XU+cXMPFlPdypaeasD+c9wghxwdkSLSRdnVMNHtD2b5/URzJE0UiUS//P98wyb2hiOioRs9
8HLHDDJzuja0JbMYFomLLXF+iH1zTsLGYl4Tre5C6z4XbmxMK+lkyEKCbCEJYW5KgXwuRs0HNdWj
W/vdC6GfwqIeW2Ufn98lGhIBzTlmZOf/Y0zGIVXhROQrThwuO0kmCFJDK1hcX+IRReX0Eao3Zcba
b7hBfNwMBKJhooaBLMRfHdOxQWXBjVMfDIQqO5/sac0mpZiZWMpIt2x0g4G1nhGCk6MLxX9b768t
rwmEL1ZOA32wJCPVI/E5yDmnMbLdkzN5H7CbQ2YSVoN0ssPOJN7z3NSWo6m9Vqc85AaD+iogbxB/
yUk/975MSbgXvecQ/fwLI1hUSOgLXhviPN01bljobWj7Vu32DBzrNDLIJD9UZvBsXoVw0JrCPA6g
2AMZhtIA7DuxuzFfbesh/zQTkIh12V8g/5lWoKff5xQ+icVsVfN5sbNz6Ml4o8U/wq0RIc7mNHiZ
B/CDKmVoBZlrawkjd/MQeDPGb0nFc5LkOj7omvyB3umMZuWd1QK4Z4i92lXZJn/Lvl5c8ZirP/K/
B0Q0uyBSvtYEL/aM48wKz35eJ7rtvpgCt91iq54WL845dhxvC16DQ+op4TYlGX4vMdNyB2L0+v3w
IbGYE9nRZJLaWjg1mxjoruCE+QWweinytqpP7NueS0mP0jdFOjaqEs8T8SLpmMLGaVQI9YjYUlhH
Ncy81IylKvHQ7jTP+XPQJRFbZqan6G1M+f4R3VpA6rUNZAuFv3vbBugfALWFQNc1W4hF65s3OfS9
RoTUR0HdHp8l/pkFtYXNIK4kV+QnU3wWlbsuOiPC38kjGYx9BP0YhMFgJRzeY19X6kESPko3zH9j
dzn1M+eVUJQFlO2YOoq1YMcc5PRcVfj0/zPVwacaQbpF90NHLRZn//kPVnNa9TNwzyUwkqyNBzL3
w1Hue4T++BVsbnvjNB1yjAt5WrJ1jEw8NrYCSPyTDORTpqZU0tMdlBhOc4CezxobX8CFzYdP5ffD
zULpIkx2UwyaRaT+h742DWRASB/9efhqP3ft9txNPqdHaXss0UN1Du5KZQ6+b8CWu8luVdZI4nDE
D8uOQCCnJrRTRM+LalEjfwtgoVpSCxLwutmpMMQTMcSELIHOTqGMD3qQ9RsHK8KzbDzn117uotu9
DZkbmLPzzxe7QFr3yL0BMDGct1OiSbfCxwoJv8hXlPaS+7w5EItTlfmhMzUvkXKEzf/9PRcIqw5c
c6QyB5jtxjsEB7M549nfaJZbD9HFiL5v3pvbs4OXnMbMMY0Nd/k0m4tD5KRbgrQB2yqIRx/rkVyU
XOBLpv90XYI+Xf/0Q08z4dQVOEU9PUT79t1uedl9wV0ybI3NQaARwMWFtpfiXMKhUTptqfrgD0IZ
YmAMgr/uPJeiDm0VZmTxTaxBVudU9wt5WbS+zJ5GCmOfxIZjCmu5OITthH7CKv7NmnrGYOZMJaMc
D5+aX+kJUOeMM5NqBxv39mfLd5EakIRmaGtie8Znk8V+4CFcExj8ojbk+wxyV680DgqHMf6LmNaF
1sC84Y0m5xN17D8QnxTHX3sAThCtvt66Cpsts68z0uWQv/gOqTP6UmrFBaj4Pl3eHBv/lXXFG7BO
muD4Ajzqh0ia8Nk4JIgKoffDA9ArW/uYproHScRUzGJ/zt9fGDnP/nm/ubyh9dKAIU8gvbn2AX1C
CqXTseHYxd0OVuoL2MDdpTtVKZ+IQ7vZ1MfkUG+286LWYZcVKQw2DY6YNbE87HKudV68wf7oojG6
auc2mJz8ys63rJqhffNqfSNupdez+Axv0O1zSX5UEIYnHbtHTX9yoELNLhr9hw+XbD5IUWHPVcaS
/6dzxIscM1G57RGHrGJdyWldSEJiFQsaBM/A22olsqqgXsUc54BQilnGItrs21eKxmJinFbWU0vf
M+7K3mqT2Ko78N7xiD9d9CH9eysMRZRvjLrY12OJoxMFFKQgsvGz10HpD0jSXGlr6xpYcRfF717a
Nt/ul89LkZ65XxWE5s9vcD4Op8gDn/vtLWrRWjtsI/fNFRjuHJgCxp7y/o97Ny822/vmo1+rdqa7
6+kz2xg5fHISpVEZoY8JkzKhXIOAlGBChgAd83otNpcvDemufx4hJCcMFz779kGRi/flymliHWVj
HTA5yMVO3mhB5ePFiiuDHjs8EXd0NTWSMzPW15NvVdDVkCebcimyQQem5xdBwd51hMPiBs4SZYrb
OfpFh4s5iukkamOyf41mn2/yjnXUyJi6aeyC0O9fYK4gG52gUx5d+FHFJuQxqRbU/AnhgZZZcv3A
Zyu2hS6V+AGWY+v9Z+Ggc1BVQKi2rgGcXg==
`protect end_protected
