��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$Rx�y�<��wA�*;�x���@�̦�W�X�fa�M-$u����n~�%���P�$��W��kYَ���P7�?UMfT��q�6�U��k�>����~�\N�(�����X�e���/6U|)�X2pF�]$h���d.���9E��WG��L�X"]�Ad����ľS���8od����e�GT?y	7�������ݵ�^��R�q^]�鍦�����s�ae���h��L��P_���ާ��YЭF���'\��68�b�[����w8�[X��V�F�0͘3����q諵�uW� �h�u\V�?@��_6G�_�*�G���B�絉�f������[�G��U&�����~�F��AׯK1�`c��[<��FY���4I� �#�G��x[X�=�Q1��`��R>(�w����R�O�?����7�,(�H\�#h(W�EH=�������yq��Ѿ��aF����:�U~m<|��.��0=�P/���4ǆ���T(����]�┎L1f���vp�W�i�A��\��2���{�˙���x����]��!6���$�&7��DaU��, ���Bַ�F(`�d3���*��t/����5_Z�"��wU4zE���J��q�����g3o����"��ܾ��I�n�SضM�@|��tE�KL�p�~�Ja��A��&\��Dݖ��#���{���� H/t��� �\��>���~�k�HI�����*��F��f���g]��c�.�!�^k	��C�I��TF��$�`���� �_�C���q�s��Gc�������X��*���g�>�хZw�8���oC��x��aI�hdv��Cy��~
�ࠡ~t���=��V�Z�'�ж�(��m�de �_xA�f>E�DDzzY#��R�;����^:�Pt-�1��'.�&����K�(h��P0�N��"D2Ip���҂4�ʈC���jQ�ȗ�@U����]/�P�@q݌�E^��%��ap���,.#� և��r�5�43��M���x�����v��R2���i�=ᤁ��'�==u�_���N�!jw{�n�!1*.ӗ鷡��p� �eT�CP$�*�!��]?SsU_��S�FzΟi7�k�o��
��$`ƛ��b��@�?��$�Ҹ�y���a|!�ـ��l�qWǭ{@cO��y����A��27X�ֶ��S�"8��.�>����X���&����@l��E�,E<�</_#�B�qEJ�����(%��&������`��#�Y_!�Q	�M% ��ɷ�m����+Q��<u>Eu	��|f�k2��Yĺ)�t[�<�xsHհ0|���,P.�U�[��.#�Y�5�k���+��B���6��β6Q��S`�����EU^;k�ϊw+WV�^�X㝼���Q�:��F0V��7ӹ�w8\(�3N�Z�h����9?��^�[��|�qz��z�|�@rf��8�;)洦#��Y����h��a�>4�S��p�o�gf������r��lc7Hc�wW��Y�a���g�Ux����	Z�ƴ+4�z2�II�a����a��-[N�Y"0�<�B(8������Kr�i� ֪M�`{ 8�����u= \Gِ��P��>�_� �O�*�?w��k�%P����y�E���X�o:��X�IBQ{��,�`�M��������#N_���j�x�)n��j�Zz�����;�� �Ԅ�� ����ô��� �����Z����L �A��S>E��r�!䑞`U2�XY MS�}�b��}��#��o(��Q@*�{�N���ɴ�W�6	j�uI�Z�ʰXL��C�
0'F�`ϗnAp@��O�M��Y,�f���ns@�l�0�s��&^1&�c�Xva�Й��r8[y���K9�G-�x\�=��O���������	��f~gQ�<��;�q�ߤ�^��n��N��oy4����46OF�e�Auܾ�%&;NG�����Q]�`��U;:m2��;�oW����'{S���U���"8�R�!6U#=��-�5u,�N���� bYT:�R�@wz�=~l�^.<�r�&|S�^��i�
8�t���;�n�v�bl-�A��V	�Nc���y]�k"�����6W&�����E$���3=�l�9VYDYy/��R�G�5��3j��`���0�;��D�?�u��V�[�aC��f�ܡi3�����ŧ��q,���?�G�FE|�)�~��˙��nA�́A��(Z�\𝟨�h�8��pS����ģu��m�&ЍɁH_�6�c�z_��o}5S�f-e�݂�4q����nبxh�#�AI*e��V��n���[�P��yO�����"z�[���Ց*�us3TYv=1����*aq_�����ig>j�=
W�J�P�1\�E���*���/+O_��ms ���o6�2;m�l,�ܲ;��^������:�W�a��x��$A��?ͥ� ������y���|���d3�(`;�&����-��Tn\�t��"D����W/��j��:�x��?W.t䪫LB�M�ϤE���Ci�	1Z�FY��S�y��{$gubM0�`�i��f͢4D���Dj��GN������,��_���aT��]��%������}�v8כ�J�4䰘3^pQ!c����d�����kݠ>���ky���i��J͠�p���c��H+��79z�Gه���v�>�,��Y�R}������l���徯�F�TP�r�^۳�!�Q�'�%f��(yB/�H�'j�Z��>�I�����tz�Q��k��l4�"�w�q�3�Q9�մt��h���P���U�K��R�3��6��ͽ�dz���#F�ҹ��Pϗ�fܱ?Ҭ7��s���3�8�������/�e������*?��Z�y��ѯ� D$�X���-���|����+r���wǷ�� '+_ǚ���Y6���J9���z�� ��O1Z��O�J���'��f�_7C�9,� �'']5-m,P�	�,����<��fmrm 0�qETx��������qμ��Y��]���{]���=`�n�һ1W�\����6,�_>�*Ӌ[����c��+?5�a�#q��� <�2��֎q� 8�p�B_w8�?���Gp�ۙ�']42���w��^j i�;18��å��Fq����?�v�&`��j�+,���K�5�qV�]?�IzuU�Q�H�4)���D	��C��@s��nR����n�ٝu�BϺ�L���2������9zkڌM�������EY]�����~e�2�]TD��,���C)"x��^3��3�����<r����a���D��Qmg�$�/�4M�ϩC�$rBG�b��f,�W:sI�%�kO̱U��H�C��ְ+6�Ǘ��Z$�*k"�l�:�E�7��Ci�dG�X��W�t�L�����{���7�I�hK>�꫌P�5R�/b����Y�^o/��u�vH(���ZG8���ΐ%�7�����kp�� �~���S���1XX�Րk_meWJ'��*�'�hǟ��-�Œ��δQ��y��6���/�t�Tl-�߿�NH�]8���%�>�G2�a6�͕����Bʲ(����q2���Z�	��eUc%�Fا�Ʀ�w3H�g˭J��p�ET��Z
�dOl�b�{XL}[�8h�u`��^�t�30p������~l�]=JD� ����vN��~��O���|0�BI�
��|;���-�Ԁ�,B@�B�K�!���I�h(0H�k����r^��7�Ǻ�ƻ�I��Q�=�=�{��;-��!Er��O�">K���Ά�o�A�c�x�����AFN2l��kF��&> ݺͬ��%xv����{�1��T�#2���� J-�B��P�1��_ʾ&�JOmٲS����|�&��a�ѡ�7m�(�F���X�#�(|M�B�%���;Y���j����e�f�$�h�ie0��&��!��N!a�W�}<�,!� �x?@��T\��h�*
�#��-gfʯSy˜{%^��!a����u,B[CV^fEđ��WLj��
*6|�k�f-�=�AU�l�t�#���l"�@� ѫe۪Ţ�X��BN�G����˚���˥Z9���:uxa���
�O6$L�j��u��&ڞ��xT5���0z���o�j"O{��6���|V�/w�x	��o��UرzTѼ8�1�!iu��O����li�Ɂ�������3�0_���ڞ' h�&�Y�|�
hmBKͨ�Y��?SQ�~����к������g�W1(���˘���S:�{g��2�ދ��B{����?��A62*�p�3[Ө�����d<��)�{��Mh�V�C{� T�NU�Ƶ����_��[�U��*E��|�-�C�:1Y~$9O�T��&��'	�A����؉�m�u��]�X�D�N����]9�a�@�.(���-�'0(����%�ZI�!WYe_��t'�����:���Ѐa�=�fԅ�h��""��
��.���;����Ga2ʢa������m�F�^�o�k^�S�W$�rIN�/@��y�i��� �.W�&�k'�.����"`�����@ 鷱}E����*��:[bm����a��t��vRm�*E�A���#��ac��]�c��=u�#�c���EB�:���P�J�҂����u��)���C*A:7g���� �9�w��F��$�y��i��{�J=����C�|�ScJ�S�)�(���=C�K7���G��p����ϴ��x���#��0u��pc�o�K�By(e�_��_�6�����sI��aK�o�/��^�Z��;��s9�H�VY9(LwDL�_=��'�R9]����X�v��䋪zھc^G�PE�#�T�_��":!g+bjw�>�W�L��b-3�X?�Y�p*���c-1&���AJ�͆��l�������G�-[]D�����|$$�%�SR1c�++������P��^s>ch𷰳a6d�L��*~�����@4��hK���$�I�L����{����n>�Q|m��'_օ���e�e��%��P��6M��$se�q�L55r&^�l���Y�װ����vR8�`������;�X5�A�&)e�}� �eJQ�x�˓*M�d�+��nr|�"Fj�[����K�����r9I����BxQw(ck��-�/vI����� /�Ǿ|��n�� �6&��'I���lI%vpS�g�<��S�r��|Т�����'ʭ������/�2�,�#���]'?!]�aw_��D�,���n��������TBe��.w R�_m�i.T����~���|�K번g����N��| ���F�s���r��� ����'?�Q��h+��\szV/|]��-���s��c��k��G���	���|Úw5s�h1ה���f���$ol�7�FP��7g�enoR��Ix�fw����� �t9̾��J�p���+lH۳��K�%�PA���g�����J�g��D�vO�s��1.�oW�5�u�L??��ѩ�q��-��IHs;7S��fm�
Q�u�{��EBsu��}�����Y�uM�	84Y�X��1i��u1�,.�~�ԡ�-0��֗��^5�z1Ϯt6@X���I�%��&����]���!�]th=�T����O?z��<L��}�k,�.7��9N���;�!C���'/��˹�2]~BL����{#�������#g!��6��O��� ��E/4�N��o��W�L@�p����$�ź���ӹgNyJ������~��� ��׎_��U�9B���������'��zd�lX�;%�䪙�)��V�=6�������8���{�a3��ۚg\�{��2g�-�]>�dn�
u�ȃ?@��#S
�@��4��>[�k4ȅ�u��j�T�����[(�S���I�9p��Kc([\�w��'�(�z�x"bl��LR�؋�q��u��C-�%�_k�B���n<���K�,c���e:1a�j��O	nrp�y�b���Ю'Lne���º�rR��I�v�
�"��xO(
��P#�N�Vxl�j�b��J*H�qy\�4YO �'QǮ��P�*���xD��5�Y0g��H��X�;�s�n�ֈ%�=�?�� [[U�b0�w�l>�;Kg�O�����-ڡ3�J4�~��V����k�>BW}r����q��S+�0;"rh����0o��3'��)�99]�y�&~CE�Gc�,���+,�6��n��W��М���#��,\�3���ė�Ǣ��˩�ғb��P
�Z�;og�8'V<����S� �Ny��[СH��J؍n��������x�]�O��9�V�Ul|��!�
H�Բ:M�b(o��C�Kil�2�dm��qE�$s�[Y��(}�73��r9< hLJM������md��p�5�(��2���5$_�N��0Z�I��p��Ⱥ���ӎP�<&}$/�2H��;�_.��FK�#W�O#���2!hkN.�P��lօ�NCvL�Y��l��O�e�"�&��J���s�$#�m�cg��~�Q�+a�j��R����垫�=�B�A("��B
����P���gS�>�M��kȁ>z��r�)�����\��S~U$LC�`�+^���M;����֤2t�S̀���^.ϱ��-l��:~��vu��?}�μ�dG�-D���C��T�m�?'�)#�L*�0�����=�a����wF.�@s/W��@�b����t�]{�v.t�"��i�6�Ճ�^�?�7(XU�s)�W��&������!�ӆ$��������\�ĳQ��r��|_l�^[�XˆN���t�����7@iw	v�Jc���X��WA�9��o��?�E'9����/���_z�m����D�3X�����76L�P�`dExR_�c��e�K�����f�Ƀ�znw.w�X�eI�s��|1���R�h(�Q��a8�Ƭt�����(E�c0�t�l�$?
}}8�1�	����''�~��6c�7ѫK@ĵQ��$��~ݟ����nI��9�����K��ͿG�b-e�v?mS���;`��6� 0�X��H����&`p�z@����x�l~9Qΐjϝ��u=u+�Q���A��U���6o��U2ǁ�hlE�`\�����|�ߎ�A������+��͐�֯(�b_��@Ǒvp.�g]"% �5I8g�FJ��ਤ/ǹ�)�����H�O�9^�f�#ޑ����G¨B��e}��P����T����h*}���ߏk�YB�߳b�b\��90���.&�gT6a���_�g,^$71�&�t�Z�	��pX\G��iy0�9��Q	�&X_6Շ?��!*���p�}j�j��X��3t�n�����7!���0���+ j
�M�,/�慦�Iɴ�$�7�I����t�!�g\a!��������3vݔr�����]=I*�Q��]Է�IQH0�M`פ��r`>�G�|���[J*��D�F?�m�|4u�/��-Ϡ��bt~��=���[���ϴ��+��V���%��\�Qkh�����������o#��i"����������	�����ܰ-�k��\?�>�����y�����K�=y"���E�s��'�<�j���y��t�j�yZ�c��=C?�D�2�nS����� �M|a�#�S��y59�N���&!�AP(�ZL�|-��!(h�(���-�_J� \� (��#�I��W��9a{�Q�E�`���2o3,�56.�p��d&k�d��ܰ ��
�p���Tǅ�(o���L�@_IT���n���Ѩ����V<uɠRp`�$g&�tC��X�hLj_�&n�.�a6�K1G4\R���0c�}���Ý�Q���KQ+�Ҧ�&c�U1�	� �Ʃ��k�ߙ���/�a��&z��v]W��%���,h��� ,=]fkX�ε�L��t����ż�Z3@��^��DK�~���G�@,�ǎ��9�����[��2Yyz�G(mt���Sɀ�4���]@����9yt9�P�&;�oV�W���-,�~�
E�����r�<��-�$���Cq2��6�ƽ��D� z�G�@�H�W�&�@Z��&���}���Np4�<���n�T��B�$�k����ĵ�kl�?+�mҗً��I��$�ő��k�|�˴�h��%�.� ���ͷ�Y���Z0�&���M�t��)
q����/�{���s��=;+�`DFԴL���Ad�EP�n�8.�r����+�,3<�:�C��o*��
�����
}�~3l�Mߦ8
(V3W9�ڸw�T��k-�9O�x(�DVCS*<nn�$Gl��L0A|U��}z�u�Gh/B�n�G��Z�(f�$��1���ï�|�&X3��*v�s�K�d���qh+�����PZ;�NMS�J�fχ�Ek�9fq�}��ى�m(߮O
/�]��-��E����$^�t������c%��/��������mHi��>2�y&��Иqo��,18,Z����<�߇�-���D��	�8���pa���J_�TEeI�M 3��,G����2!^9,OZ�Oi���s]��}�ȭ�%�Kh���.)����+8�C�;�5��)`v-YdҺ�Μ	rpA�a�Y�+�e� ��\���2��#71d�+9i��/`H��J	���RE��C��5�^�!�)@(�����TAVt��I��o@�sl�[�	,h���Z3�߁�
<`���ޒ�`��ǒk�E1`�/%e����d�1��s�X�u�_�W掔��I���.�ݲ�Tϖ�Qo����_uO�#�X�8UtT�4$��CIl�>-�2B�ȷ�������\��C�q~#%��lz���Ou�rо�n���;���;�T�
"e.�	�"N	��*��v��� �yDL;ѓ&{�9��O��������-E�wU���N��r�:ӎ�@#l�O����h��5�HV��c���qk~�*��x9U� �,�b�����mgN7|��bAuC	E�d�t����j��;���8���9�-ro�5.���F��3e��]�t`��KҺ�D�3T��������>�h��Ʊ��M*���wKX�jLE[�����G*1�L)*�%pi�|�w��<d"�����Y.�
@�9��V�� ��&�T.��Ar��q���