-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
iNwGQ8Q5QYC9R7jQla70YWBgop5D181TVBgORoUUkSNEdihvpANHuKUAMMbHwqBhoAUrCOV2Iana
QGSl46j6RsZW77opNfLHBx4bic/AC0PBXZX5rCKJbqY6TGHOiWmo2WWBLYlk7df4ekIWI6ZBDISt
NJe8wz5Jd8OPTyYYThkPS0WDbD4iru29Ap9T0AjW5qMwdjT5n7M1fyAb5r6x51rHsM4qolZuyCLm
iBNMgHeZoxtRXgiJZf7Ueu8nZFGlJVjlZSJsdV7rQTcL++ydrh8pYPRfgtDD3zjSj84mFeRhYV/G
SdQ/q+50vKQAiQTcRAP2U3O7cxw8+Yu9jHc2jg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 20544)
`protect data_block
k9s6Tf/XQA047DA36xx0h/mEoyuKkS+mP63lDpO1P3WBGrL+vSbbObPv/yUuS6SVmc8Bj60fshkX
CRhO5APc9iRCo3XywqB4AB7m+mYRjkcuU81Wrpr0f2ZMarWNT+LCPv0w3K7NyRo6eR1hEcjW0KmL
31GvhzXjm7uGxAbdixhT9hHa7hxREIW3rEy5jU5HXqSQ/dDKkAN8M9ITuR6Ij3elLu+0uFrY8SI9
TDrbstGe5bXBEMdySZmEUw0/IhD2jvJH+ThHvuwSZ+g1qqfdSGTIo1+7g3MFkY4AI70V1+4x5Uxe
ACpsnuwGD6SeT7GIuK42yiJLwR3QFGx/Cu8+8g8mEbXj5poLwvmHBxkzp6y65Rwr2QP62rh2sXmD
XelszH1D938rU4N6DxTsx2jN6sgVdDvHGII6HXIkZLmm8ZjajUHaV1VZTrPmN7GdhQLR+9rFfZ30
30PmtiTj3TcYpmjruKhKxaNeCxVBFoMJpTDpGSatSQJAzpT5sKX8hml0J1/LICt5p8Az1i8zxugG
7Le3W3sZ4V2ZYy8qG6sITTGPKgogEFpUSrZBErGSqNTBVonVs4J3shhPWDNyCpz0BuKZpoFipsJ6
04kkPZi/nuGJTT5/Oy1nR68G81nKSlT6HyYJBNz8d/tUY+avwVEJuuv2nEqsjcX2ii1/G/FqmJSt
BdoxfOVm6s4cAIxqfrLFC5bw0P7Y9mlLqXMACCD8LkaSyQCvHuSHYZO6S2zf7djddTLhYTtVjoLA
Sf7Gpzh/KrNNyOB+dWBf2ASPlQYAnRN5tzKKt7eNBGQo6Tl227tvxh8wK9PZFfqk7X6jaRHbHc0V
oQ4sIwg1Sqnmmvnkx94sLp262icR2NyccnaSxbiIF9S87JebDxDPOMoS/pbd72jKeF9q7Na71Vxh
PjRXNpABb0mYpLrkPxQxwY35V0RmkqRF1rqvbeg8Wm3EYnjeJ9om8S1Cjd7D9PviRMGKD28+Mjg1
nY73rsYqtHAE5wZXgD2xufy+ydiq27l7LeMSBXdr9w6aLpUbg3WADw5CBWiKGLw8bgLwl4Uoynse
ttAej89zBeT0e3InHtaWUPePAsSfmJ6aCVZ40/u1CA/MO9URbArJsTnDBr87SApxi+WWQMSRGKLC
gSF/0BvoIP/+IAvdV13zWijCZwZQVtXqNew0pNVTpdxwwzj93BQtjl2wvjRfTt+HHJapr3ypI9ZK
qEZeAYCyjluJCp6bcgeJToQSpDdsQmakQXRxq+2CsR2XZVkoN7urBmDmYICz/PmK1EHeTh8BNzfK
wlcYIPnduNtBW2rYpAQT32SvwwhP33NoVW/RlIaC70vVlhlnGgQqG2stOL8uUcuIAffZ6RKCHK24
53wDE8qTjsLZp0eXjpdyEvdXnXVdPs9gcp0VSdlcLL4ERiw+x5OfuTgvBSkq9fydfKYsJLfaY2dS
H+o0YmPJkTP7zpZO28vYSboSzClSQYxBqngV22Q/LmnsXTn3rIXloD46kjbHddCZPflpTdEC22Y6
ARzOioTiKU+6w+9rNC1ae2fwuOwWjYt6JVWNFZ9gLV8A0xnZpUgGigosDKLbRAPCdfu0nmlIuNaR
ROVTuLHEoC4btMbpCY0O2FAGpsE0IZLOKCg47xtWdE6aN6h5mR43A8etAn/kBn76AKFRshXlcVdt
U+oxdFaunxmp1U2lTk1TR+/EjUg+meYpX2pyG1EbqHTghoSliZHDNIol5mrQd3smksccrcJTXF76
Bfld6Egfuo7F3aZBJehB398FqOR40jq4oj5h/hBFA07PWYdDD40Cf2rRSqauiQnj3uNljrCnPO58
sWlnlhISmkl5Y6no1dPtuWpKvaqgunhRm7VbLABAHD5WGXOxdmKeOKp5dlsUFvCSWrpeg4Z0vny+
bHgNtWPX7OzI6dy8Y5a1a9KD3O2MZD5e1EiElcxw0oEGMuo+sz6zuDh+6UnXQhAS6VEgaeetVSIf
NEmRXaNx/IfriGiC5GcgIjPR+7xIb9NEEhNYAINEoin5tH1UvTxFIEHqDTqo72+XybAYoaj7rSFF
XRjpIwBA8PWcF6bh+uQhL/rigBKW9ob4ufqlcAJMFd7BJzXjpnXt17VV51QDMsn8kIkl0AEpv0A9
VtRSHn5Pp//oY9d7cY0Ml10IAqKFpR9Aq4uyLEDEg5Mb7qa0V1niWKFAR/dvpau7EZpKIPBSrvzy
X9SiwwSZ50R1Y1Sz+p4PHrG/hRWJWSBZbhQfjw6/jSwUSmFsd/i6QhwfCFBRBIYJSW8osTRCZ9VF
u+gA9ZpgnemSJgMPfmeQ9ge3d8/JzWDyMAzvs8l5AnyUKgw2A3gpV5RY4U25VIORzwyuqCnrLl0c
2A364Ccbp7HgmzlQsGrK7EeWYlLHilwyVBVXf7IdVz10pfsBZ4eTq1JY5ju+mfGcija4L28Yyq9p
2auUJM2mSnuQr1CgZSVNcK3oOAZDfRqZdb4Y6KunWKyJOf/a3SBcvpgImCEhcPKkWB0xMDqVONAK
zeJhNIG1eEnO/wMJuecKK7ym5Auz659qMyqWmc5cjHDL1KHbOMR5mvTys4/zJkm9SB39EEFpv5/z
R6UoBWWY/hzQzWIWsveDB5eyvgN5eCQgRAbyf9jlH3qHtFW47QPkGCnq3GoWwDbS+eqOrHujFdIA
n/rf6P8LN1cY6mFrqrllbR4FXW25/I2UhYA/2fOjgpY12Xf45YFZd5qxBYrgACXHyA9hay40kDiS
5b9FM6vJmU5lDjHA3tZdx8XWZrilJy7AgK/K3dvK7twcLj5ke9ccI4Np4819nXiLKjN6Tm96LDRP
/HwJFrqn0aFLTj+2ktQIDREc8O4ZbaabTYzcJDT5XgvbyAy9EEeSM5N92t+u6BUW8qn83/J26wS7
JkTZyuDx59KKL8XRuthDvXIOchYAq6KiiExU1eIQ69qdeYxbnpMHN++TAPL+8mGIOHstPzbTSupM
Q2Db/k9noqkcByvIi0R7kIxwRmCe94G4AjFG1YxxsWcPASYdWyWUU6rLJXw1Wz4DIKErbPQi2CcP
AMwK7VhEPrJicCX08+iAjSi80yIKdcTEMR3QeeWpYBLcACcxS83M46CQAIYsd1Wb49GbwxKoMehA
CPvCiVgy09ZEo6qRi1lztyy2xLqvPd7f7Mlr+/bx+Ex+R64zjy5Sx+fsBBpAr3V9XkaN4mOMAplY
N1tO/qv/P5bDVqLDGlhvyfsF5v4GxaJWvCnkQkIyRbiz7+3QhczGgyJnld6ze/yU+W4EMU5DWnrx
ckVZPAurQqXdpdYzulKkN+AhznwXYFF28XWjo4SIDZQl1hJokNSEVsEwE1yJm/yZfJRtSFNyUqNK
JHigDBLH5n6wKP1a5VzuRd5BVt7eUHd3cHngW9zZa+egtMg6HsmB4gJ3Doovww+O3Syni8CmWoiT
McqavDvgop6nhO4VmsulRpADXh8xW+DPV+TF37Q8ZrTxfvehK2RzOIGGxLWymXVQwCehjgISbH+X
JNh6HqJWzrhHbsY+kXyPpcv6w6bVkyHltFlnOr1GVUzrhyNsbgRvajCk4HYdzip0Uc0shPlqJUTI
+Gl3wI9v8nN0+dml3YJNG2KjvJlQ9Ml8rxp1ZutijWyLhRnup2cWf/7Xj9+CbL47xcKgFXKj/Yxo
dFX3NcoIR3QY0jKxhTz/N7LKa5mwH96xVDUMcRKgTWCxmdQn9PUWDuxJsLOw+HLBUX4/S/Y98k8e
DARPINnO97MUiheZ+z2QwTHudFeIjf3uqT90YbuwM2GJScOqcbJEJMT9w+4aQ0QrElrF1e36DUdg
NiS5rYtw/c0m9HSfVwdLV4Fcn4uMBzcz4lN5qyb75CK82Bch/zeDY6GdAKK/rF/uyNGslFmkDg8s
RQv5IbsiqXN8tA0qjsnIy//wLTT+/qb4qfZ3vASFvWoe5Tp3qwsWxmArB+zYUItxwPVWB1J+SjLA
ZJBOkfLHfdp5WZtnixVO4PLiWWL1G1z4wl81QZFMNrxXwBggNqHPeHlrlGG/xvAxD/uJFrns0C0/
H6kC/+fLR+QRZO1WTQKbWGrhlCA/uoGdAqIkf9nMiQCqjUJE2L+M/OcqcZUGxgzhEiLLlC8DYK2j
byJNeNckQgBE2Uzyz/RxHEHaWfXTmcmowYEKvfiJYRwgrzo5xLgJsf0bks7z7REP3QsEkTKJsAU9
y3a6BUyC5QmJz9hKMsrYgK9gd4q8H/Ft63hgn3GUAE/57lhtaHQkzRljW79TmsP7AzrPmDDSBX+8
qymZ7rae6F8in7GQbShs37JJLWWbkEFkeGr5DYKd0J+Rj+F3goAjiIDFYab1ezlMOsjuLM5M/yL2
8VyBrXN2jt7lurkREAKgMGh28zL/mpKQH1Ce9k8G/DEcSIqVnFOSYnoDvWkULKyTaxefdi0N7st0
TfFhdXMZeqamLPRxcDLo+kH44xLNcdTM+J08654QRSm8PTV7dk64nGGDpdwCfGLai8hnxNxHTNKR
pX09x1QVYZeBObUdZq6RLbnGZXe5ewwhroaDwn9pIdYqxNb8zpjJmRr/RFia3u8TsTln3CEBmZ0G
3YSeZ682Vy0KNsUzCaWDsOwdzbB2MouRfROb+jPGfHJIxYzaAKg0msZQZWaJP+47Kpsc9hdVV9dL
ZOfh+b4kmD0nluRD7k6BtSFopYXr9qpD77N6z4RgiWS4/upHlFNabA314sjob0jiAHnn4dgBGRLb
mB9arJvxhGnZNBe/fBITPejSSROscxIrNGMc8RpeOK2pd8mpQhBA6m5w9StHndG1QqTPvDTU9r2q
2eG+pWdA+//OviJm3Zoz7+a1R55jEzhmBHwqoSK2uk8SpSyWhqYmeKqTbPkKbSSNgmrEsGl5jDCe
PmI//MVeTkp3lb9bX4c+xTxXqg/EKnG96vPae/gfAfVkyOpT+wzL9K/sY7SdRROiFGDq8MypUSFa
wlK95BZVA4LkvRV3MOh5sY//1WbOJK1gglvPB35PFcbzNRRTEwwC4St/St8K9NSuMj1Z2AwzQJmg
VkR49BXZZZLUp8Xydm5wnXpYjmEEbIWF+hSeskN7jOEGx6jjSpsHVXaipnwKGhkMIOmRPEIMTyQA
RLKTzcIOWS75dRbvIWgKCJpKOXVdQqsOEApBKfevvTYmIEDiHFApfeM5tZ1SxhVkFUWn+CqQowxk
Z8Ru7rPUS4jueFZG30co5KgBBuuXXfUWnzymdDlI6qnoTPV5tRWyUF0ED5D3HnLF6/oe5RLL8YRe
dp8+af9Sx4OupC19J3ziMpnpWkFq3ucZCjnLLjasmuWTS/ceRqja3b4LEnwUPEiZ3BMk7X9WWsE0
DZPxkBM41vRAcf1S1kWj/dmTCv0J88ViLK8t9IIrh+imlArBRbA3e2y7Q8HNvKPBnuvz/6D8aNNF
SuDjQcFTA3/1wtn0a+eAomV47HMFATPsGo0tyhOovsFotLNOL/dhpwoy1oiDd2FNU6PIElmEt1e/
qLy3/X8MTyMwbcaS3SmEgM/WI/OOeVW54+YXqsS9O+A0t3TfXzgqLlVnKFU3UO2ktxqdTcLIqfL6
Dif0vzQuL1SgMkNaR1wUuOW++DUBAl9oLtp8QvgF3BIDmoRS4n5S9yHI0UIlTKichbJ1lBivQrtm
3JeEZ+v0i0xHV9iQ2yUU9bsvxPWhWQhnHaZN66JIGkKWn6mmw9xTdBSIDqD42Sx1vUhp/GzGQ6AR
JRM5hJq38wUr02LDdnVWuiO4HJIGsz98eobhaF+Hs4CAPpqVN8P3TiCsZcVei5Cm+1mOX4OHQGhC
fpQDPih9M2wT/Y9+dZhqPkzGWkareMfJnO8TQss0eykntnUyntv9f8RiKFHcspT5TDsAW2u7RJR/
llw3WRQ61PQ9PkKylI3mDJ1QtkdbFWbJMu0YDBl8MT5iRO9qkI2Ps+MQiRQEnw5BcTfguss8T6r1
LOe0/X+nvrh4WyVaVuUSL1tT8NL2B8/35ja+G+GafeUwMVdM4a0FFMTaqSOXLEow0BqF8fnYsrch
tlW7ysAltdQaj3d8kXa24bNf/8TOXs1hxtbNqqovOCHPJHlMqlVGY7Nqv68SqQ1p2BG1eLfgbdyg
z/rdsg2AX4/7ijjQbyps11yJj9ORaIZ+dsPjl3DMfcOQMMhmLGN4C/aa0zY91DYfypzv/mWIpsA7
ufg6OEMQwg0rqYU3q3phoYz/CtudlBtq8U8D5GKVqEg3O3RTLIrAN5Q5ZruMfuFqltrNCW4dpvMU
/xBaJxySt26R5fyiRQM6p1d3v/ZbeIUZwq6SWQnIgPYAWNiMBIGVPh381Wwqzm+/GLwz4L7em1cz
KcYSIYLVJFcMjrxXFQEQltCDCZu0VJTvrX8jTGebI7l7ud/p2iNAGfHeu2cG/rSI/4/rglo1q9Wg
mrt8U6TZ7/E5uDxPlTMB43A2+dj44JcQO4OzwXN1/R6lG6ca5cIpT3lvhpKODWGuK55kSKI4hCUg
KF93jC190nwXVrdAAAnQqssyFMH8G1HoLgdNPU9xO22HIwIhZR9Plozn0WS9jKaBU7F94G3XSTR3
vbwRTuQlD07gOEx27yMow7JFNvhgSzKRNX7DRE6sQFa12kCK7+JGqqTx2un8bakTTLoKSTJDyOwm
JnKZXl96om83HxhWGAoWN273C3RXlOk3bU9SFI+jWRjBhBvVbdBo1ftIbkapjyU8e+lki3DvdjmN
EF6Blvwp8q/XE1//sj8KH1p0pqehh6BRZEg03zLHzBVQz7OFqKZHGwL9eMgwzMCX4yyW1YtWsOIO
0ju519zWoX4tHXZNRqAWmutclYz53a4HsgJMQlqILc7LyZc5F5fuLj8D/5Qkl79K4F1t0YKkZSHe
+F69C+eYYRQ66t//rkxJ/fEvYN5o+3RXonq2CvWr3zfFRieZ8pa6NxSEouWC0S+cRjtNMe5OMcc8
Kpd0KhB/E///C/KVuzTEiH5mHJRFJpbEyKjI0qwGzxt9vKRFpLAKXhd3xay8ZpaWzWTZIQ/heoUK
wS0hkzXBPNtVQuQtfaWMxm9iNa9Kxj/SYF1VDnSEYBh3A4SFu0oySza0P8PMUFVTShETvuxbxccR
JoxGlO4xV6yuD9ljYwxfoeuO8H7Ek8/FLpwfb2NINyhtXSmcrbkRCB91Qm+y8Fv+/LcBZj0+F6f4
EbJezfYCBFoxQI9DkEjzc3tssx4VUCpwcL9Svnp0pc4YRp2LZ/QVZjoKRgYd+OuUE/Y7syBubr85
Mb5kTdyhOcTbqrEB5LuiFlsncj70RwYSLq+1MQW3G4R9/GavqdinrvUbZnozqH4vPUD1KbIBZNaq
wm27jfX5KEdJSsRj3i2iQZiIN+9K9IBH++sTUmRMN6plPJ+b0C6BlYoDn+n6JITfmlbq8WEKJLsY
G7Z3woSzJfyX+9sX015SMMQCjbF6Qrhvyu5jiMyfUlpMakRuaGf3ji+epNC937AyAdFajhoT8Xpr
GHTavjKV7Pl5CCVTLU6X+lyD5999Tw3GGdczZvpj2i8u6wJc7+cr9Y8VY7wNB14bQiHviWft8I0x
LAGPCmFAM+6hsw2LTUpXMYVkRrccoNPCcF3dQVyqamZszbB5Sf2emCaufyZ+qqZtgBEgEclLToTE
idAT96a2jmfgrSP8IpylGZSY2aL97CBiO2P+4rI2yzHihue31mrD9OBD7p/vsOnxM6z/LKZprw6A
q9T2muICaMGw15BNZu/JuBo0pTHlV1B1DjLyXKUYuin1eih1VwuGgyj/77Q9esouQv0fCkWGqJ78
YljSV9uhmRxev+1oztEac2D9dnzWzY+iE1E8pzv1+m+8kvMQzutYROMIdOQpnlCMQPGbiR5qHRNS
5Syqmi3bWjJluhvWnIWk0dnVQIaq/yDL/1nTj7vcaShVll8KB+jSoC2jYqySe+fNIvPRMrstaSt0
D3pxFB6RdEph+g6MbnKtMwDTuibhdUYlqAJm2apuGNPM2YLZporCpkJlMvs533X1UxcyWnuB6KEb
8oGZ4JLuH7sm+4PvUv2GBOvqiVKy0E6ucQ/Eu+mgPnn606kMDrDzgaFsz/e63kr8e8FXO7gtks3q
+qb8rSaB+XDlK7lJPTUkJCh/N8Y+YltdLVaqfsYj8oAZ+HLiGgv8yHW41/kas5NjoEW+KdITINBL
IqiSMQsnJzJR6JPoumZpwLoNnt9/gcXAuVO9X6t1RusWUDqPR0yK3ehdn1tslUdYybxlfsYRwpNe
TMIIwtvmvcIF+Z+UNzceONnxIJ9LD3u4anaSzCYrd/PdKJHqMqQszNmSSHRlRgezTv7XV92tvCO6
VdteMFrpQ9JpKv4QjuVBQDHoYWdy1SC0fStdMDPnqwwgnHzj4nZ6LDQCC0daIUDtK2bEKyxNE8Wk
DhOBp9S39LbsxdxkC3PP9/0hCB1QuME6XGpyUsDwqfGwyxkc2y90TgGgwicyeVZJbqHBYPHZcyYY
glPzX43WIRWhQ7b8f1qCE5dDx1bo6xtGP+2Jvdsd1VVwFf70/fm1IZQ9DxKIT3HUecQEi/JqnmpP
B+UJz08LHKEqBesmjB/wUZ5Ygq9Z62DtvAFckHzLS2KMIL3h50QXpYy+lunDRq9OjmSgdcRnDazW
gsDh3OZknm8oD4VHCUE6A+9GRvUd/zz8LOatbmAHUO11Frqjr9p8VfZCqVfkKdfrC8Gr67cqYpI9
xhvj+dJUAmo2pTjIR3kTsk2FGF50ieuYCgwSn+eO1HTeytSZ+TSHVPyUJkHg/b1SeaNK50ClR52P
IPMrLwp9CWUPTykySaw1G1SbdWNhankqco+WvjlXyrWQNsxMu+jqgnXR7FH5FDu7wwizw2Ocvkk1
76dyVZJv83jCBBLol+Nwd8+BYfzP+X9C69lk97GQKTJ90TGqKPZOCtjwu9vtOzBbjQgg9quYuB+R
qDIzdWyDUSFlJCJmJ6ACTQ38B+SJLhOENbc4lS138PcE0+isGww0b+2IP56cJ4qSG8zf+tLTdVvv
5d+2qEP1d+8NNw8P97+UA7E4Ch6vbQKhLMkupihOvwSvUQsBfuSbaVpSJSKqdY/FnjGJ7EZus5+K
vFMyNZqv+mfeU5pW+h+Q2jkxYe7zsOH+ElO7GQ1bYyAMXk1IFJ3LxqC+A5u1VZIVnjpbHil082MR
s3ApT8Ka/PKUVg4RMxKtx2ugCms4JcKvI9iAeVs6IKNNo7/fbuc/iHm3to/8pz+oXkL41IarfwUw
rffoSlXYuu00iTOIQRgcSbb+Gl9YoTcsfq5hlI6+RJ2BgDnsYnMcbt7VPaq+vnAoFWNO1U+bXQT6
S1P2+za2jv0dgDNQtMtcAsWdotADE+f+B5QN3yOH7txSznxI3R1amlss+hkMTaG1yxUDWLU+ynVs
JDEUYPTpXr4Tua0VqjxC/AeyK6MTA7Vw00HtuGbk30BqNoL7hjJTUoLQSKmhdsfP6TnKfc/VHbHf
GdziYhZk2hBgimzCX42QFHekywVf4mTAWwRh+ReExLhWWxGifriJi6J/gnzE8iMw6wBDHjvJyMEP
tHcs/DI0ZmgXvakjBTGX7VTn8MBH08Xy5+ii0RFSXFcx962vi6UL+qDLb1BRyQ+fPO/I7sTYQz8J
UQ5tIMLejSwKFUkNeufRQOwILrnDAWT2IrSpSktVNxA2Hm4pn0M0yCFvCZst52HjbYuVI5gFFwIG
R1Bp/StN8BjP1pXRDxS3jLYqwd4r1FeQmncpOSuUqpwRr+kHIupw5U03Uuc2z4dVJm0OcSaJukgl
yE8Kq1T6tbxYNVyG3R9yXrN9KuSk91A2Pawz+iOpBv9J9POd7dBBr7Th6IQdeIKe8KFcx1MfkrUB
/Ulea66j+3CRsRj2YQCea5WbOq7CYnkfQQ6eduiC0udqGQr8TXOenylkVhVlmwj1ITgt/snwUogC
Vr5LGiyN1ipAGdnwEWWVb3Mmp+OBLoki7ILE+lDWwmJ/RDtBPFhzoAK5B3ZZsv2d1Hl63EES9QyG
DhH98JJR/tGAIN2uFZM+dWTMyomZZOEXioG7MGmVbFkYr5F6BTfk09OsQCk8PMNgIew5YJTAvWt7
nftaCNDl8K3Uol6An0OpusKacseZzSYeDFjs98STSTRFPm+EIYl720GmrXU2BRgwceVqB9VcU5sX
ieo8Y634qruKLhpWbRJdYc+dPYphLxtdFebiZXg3fnDW5nF3fO3mS1EDuR6HiHxgniEoQaPrD3zg
iNeWs0RMIVXpZUoVprwUI6Og23wOiPzYRoFEDENnhm9+NYyXcwEtWeWpkplY0MKTMDe3wsPSl0Zv
pIqJeva1+EtGrH3sVrrp73m8SkeQhcyDuQvV3OM0rniA9vx/Sh7NYIz8LRUH19C0bA29n000Qs5y
hnnqdkj6N83QEPnYRZFT7kM9sGSuji27MOqW7e1ca0JvD0t2RwTOHJH8Nxc/uboWJrxtMrarOr4u
haFSXEJ6Q+tr9NqT00qyld0SviAPi6V9yK9vBxgQcT25b1oMCfPDb/j4DfPm02PxqRS2SkaHbdJA
qIpNRpLlFVkeUrLRYSH1mJdQziLTB7OmL01uZz58J/rw6umnrpe4Z0a4oYFYzxE3B67R//Qqzxwt
HnBKs4w1X0218qKYCKtVemmhdInL07X5fWksD4UXUyryzrPtjjABt2IW2riPP9j7VNG8DgXjRUoa
OFxUs4Io4uA4Bqeh9N3hItZWMnsByBRt7axZyUcHgx70py5zImjs2qeGBmU+Eq3yE8vvUCY+ayZc
14UdYgjxSh0NMxpi6c2nDUA1U88BBZzqb/UazZPPSK6f0ajC2RgT6B8aFP/X9pIHBWW6AGydj/Oe
M+vbVw4/P0Gr2AJ3CKHQ71FemtrcgA8jaOsTpt1nwof0G0HRMTxS0v/oOXLgP05EAJneNEW1kHdC
seHWWRTbEQaBzSYbWqQHICSPe7cNgDpEsM/Q+KlV9BP1rLPeDPJGnWwCfdjx/nw0viVpUsWQNguJ
3r90GQZZFoW/W0pA+91xql9bT8/a+GdqX/qeQPKfVMgEXky4xDFZeOJI6CWr+e6PdcJT3AHnKros
eKIcORfNv+ZsHDuM4Rj1qhT52++RfCVFl5/CQlKCOYSRM/S+7goVqnRiagZpcKHBQTAerrRgTzq/
ia8IoMQDNdtIy+s3D5IH5pkGYpruFVBbvhPEYMgB/F5ZXYsijkVgVe8dADMvdiRGEiN1AscWsm6U
3STxJeKwmqwjqhsOKluiKpz50bQMM118M/LaNYXk5uPiyFLJ85A66ORzldVoA4aXQyF20dgaXw8Z
cRpSgxdOR24zYK8qGkQKdhPHJyoKYEznEGJB5i0niQxyZWYpEtBoVK+qylSah+gbdtuZkzxUQqV+
tsRoZTePiMQUcYXEGf55WM2qzPfkOxeq23XCowC2dphOLuGxd7EWm+NY/rvLlGuevn8k8wNW2jcw
mXalXQYrtdSm/RRRABCXwzVORjhRXMd3Xk+OrJDUwyY00DqGUizdOb9mnJ4xe4zgptKt65+9xR5b
2mJ/sxKzRqaTpizppmSmP/RQMp5FoQMIXX9Q27MLhpWstkCeHXDTAWlz5d2w6XM4RovLeMyJvE1Z
QwB8JSkyuc8qxS3yGPRxnR5+n+WKQpQam+bTb81nRHAf88hNH0Z+M6qJZZ2fkmH9YMlFmVmeKtia
ROLz7nbRZAAEMtpauIeGpVF2kxr5Y3ECWoAx5+nmMFOAB2YWX1/+4AGdCxRDW9ZDrVwxhKjVHljw
8jQGJumg3e8MXUnZGaqQQQQuJ6tg5QpEwBiO5sW/RJ7ZbfWnNYKyzW6ZNYxCb1XSBzHD5jEUreLv
bnCzLIq5Q8Chw0QUq6l6i3o1ym8YyeAMQyifo3MOhoTTS/4Z+K6Ml4ta4cviIUsP9TutpjUmgGJX
fgBk+Jwhut2Spodp9P3binnvSCjxi5d4eUbze2mxBbRQuAQmjttgQSa9sCcPUybG7bQBYjDrhoQa
GB4vyRZLv5WVsnXr2asQmxkoSOODhLmzs3ebrA04sBx3YF3spWREMhxZudXD1vsu6MjPfMA2JE5i
JTM2dp9YknmXr0Vyqma5namk+Yy4eOCVB/Z/XSe4nI66xGVRXQGKMi80yTiQeTyMqb9PqYrP/y1z
BO63QI85qLuPADvVrjV4hibESvx2McFdSVem4g/1owWZct4NAocl11A8g/ETeS9UpOm8GMCygIzI
cgsJO8y/thePJun3AYdJ/1J+6c0qB4YrFsWDtkqgqnczSW3Tjli/mnue+EI/Z+WtotCrMCk/fGb8
ON1FgWNqNPQbWZQ3vRtUi+/U5MfnSLkpCBzFtm0kZDrxgyyjue0rg4C7lx122xIqpW/qlCCA/Ija
JYX/+Kk3/VIKA3zpSSTv9AcvAKWi9qcYJFfIrsTqTNAScgrXNFDvNwmbXyBJnBXCgWCwKk3FdAMh
/ztmpI4MSAWDq6UUf80UbIrs1Nr6mq4PWzC9rpTRCPR7rir8ZybBLgY/SW2px4PrlEOJ8gFgjGzm
/llrYzLzrj6rK8lZs8ceGu5uCfyQHPv0UbwmoculuurFOmW0EWBQNi6Cs+aTjzAm9wYRdN6ZWuV4
lUzaMbxiTRxxM22UniYClX6yRgrN3kox0eGAFOuhjnZmYKZ6wlmwJsrVH9Vke5UCdN3xtduvZnoM
LwFHYe12PTNKpgha+p0Za3KfbNmZxtgoLiP70jZefGQ9sVyoWFAYFDd0oxhNtJAflWLHZI+AXt8K
BsV3xJevFcklBW87m3a/XVmaCwR1vqFAm5LpuOIgj3UmTMpvbQgrukdM5vufIDkR832VKcv9x+nn
+nfsEwOMVxU71La24JqSKMb4WIQRxHh62rohbwnZxnvugXA1DNwEnWbnkMNFcPxSU62MAuRPJ2ZI
3dAleu7Fa1KwOekFq0PpXi/FVd9u10hPcveVxH2zJCrfbROKxNc3uxoRkPUXaNTDshakSf7LjiBo
yoNCfiPZOtw5C8JhMP8JQfcme8afM+ZLmNEUi0xXOrEKglX5wetxefKKjwkL9U7U1VP1aVSPPhzr
yBybIxG5Vf6PWGdZuA+vkc+FyOXvjaWo4o9mCdDIrndMHwS4fjOCTEvabN5PpMcvhERlc1migeyv
AyCgqH+c9LSWvMmcazC4Wg/1FNohGievlzykQ7vZj5fVzB3cU8TeTD1uokbf5BHk1x/Nk+msqAoV
LNOeexEMlV2DmBWnlFNgccCj/60GSGn1uIfbSB9rQyMB1n2dRMNO1Ve6xym3+uWrdc0coDuNLwAP
/j+5zXAoyDD3W/LRCYuuMjc8QvUKb6mmKFk9S1VSxRWKJctVhesbU7pQAl1RbkbXlleDamzDfRhY
F4XdCPqaObx2G09lykPWKHUk4ZCpunLea4w8XRFqcNuPEPKRhkS1D51xWYkiqokDnreiXI9VAiBQ
h3fkcWN6wc1F3HvnS9HAc3WmS3H+3djbgt6fnBVQTz8PkYFZjUkhwg9N2+RCemXDXdYoa0F6jzKn
+LxIQPyYmXAqOWST1MQ37xFY7YYwQuMR+7E/BIknumqYiWzSzCNpm5clfgHlVV7nrEyHbhSRgc3x
kdCQN5r0AWPUnbR5U2jrBKEmh1Y0mBbXWt3c7Cmes2wIJexTnJ7xylFEH6oycZzhYjmuPkOvp3u1
T0KDVNJEGVag8k603xip0UZFG4o+Jm9xWbuP8/XPJbIZQjYD1JFwIUDepuR/RUU99kLqxf7NkvLr
3iKq4hjJTUx21L6N4it1J5G94hatck2buOcldfle5auIbiIfTKExAmvGYuxRMHfzxHmK0Km8OlcG
b5Kxg9JpgGSZszz5f7DHt207vtKo/CJNXm1vZms9OsbzCe1nnlmLEW3WOPEhmh+YXyGvZFkiUxs9
+KcKrdhvvNYpUKOaQBmSL5VwVif4hidxlMcmY6Jt7Yj+Z6PBFkzUtptOa4Y1lXTfQ7UMFxRcWg7R
tWeB3zQjn2FIAuB/ffowhtSBanQ5Ch/QMoOnT8AAee3hlI2EKrGU6xZN5G/Mxb6Ou1rW11yikPaR
0x+4/dOxURO/MCZhiuBwjmj2tjZ0LUi+vJVOM2xvre+8mSRSpnWdHkPlgdHsiiM/pCWUMAAKdXnR
04KoJ6LlHMBMZhzYLGxinj+E/LRvtmAXO/HisnXRw60wLkLijgWBWI4ZvDlk7/W/hMqwx9EWt6Rv
cFiiG7zBnW9CiEtA0wSvoEzRhTx+XQ8tmBIqzNrpVQan2EKsW7w+PwVBSitRYbqqYLGSv3qvXMnH
e08eqBH8If4smMy2g22VdL/7wTP0gxNXeYgVw9ZFm1E7sedgNkntMSi586RwXRlFM5pf/yErSy4S
8iF7ucFhNvbafjmWLDgh9D5qBnFVjLviWg6DdS6LOesSf1x6uju3i+G1a7xxJvm6ehpt5ELW4cVg
q1caj8mQDpwxcg57CLNFTdm9NYI0LTJLQuXn5VkrdRhYjAg/vYcFXl4vBzs4JtMqunWE+CWsz/Wh
bgHgfyPtgC6caDFuWhpACw9Qz1HdZZYVHCT1++x1ZWGHwCJIlkcJMDy06QpjJoW8zj6CsWev8FmF
uBoFgRiEXyHwbWwDVFDtXtr58RJcc5Lqm5mP63zpcaHJqvNR7A97gcPWnC6mtECjTDl+ucONYfNI
G1h/ABEYe3WRQgWGotibxJH3ciGN/gpkaBNvCdEj4VmEUYwFxs/Oc06WYtPgEtrpxb9CjIZ34gJ5
gkZsuBpKfYWhDh+r/yiib0ChmEY/au2VNV3g2GFatU+8owh3zrhxdYOvQz5KtJqoN2N7Ml41kv7y
BRSJwXKtSasTgdGnU3MW9gUpnj9dra5TVmBKgeomFqmNYUFhOi1I7VYmvxmcwHzGizFwuRGmgsrk
QktawuviDFshhUq8HTc610S9PqvS9ruOOSTfDGk4I1KjiKAgpeG1SEWEzPLwdKHuLM1klqgay3YN
/HRkxJlih6ZLrKvC0hZbwIJgvwCspCEophPCbA8Ueqo9O1VwOvaeIuI6Ans1QiFll5MRF2rVrzoy
Umqs/aSgWfikdW5jEkqBJ/KAy5emX1ogwTbRiXRDc4mnpTuh1GCjbnco8NIwnoQ/xNH5BA710eG7
068ud4v+JZj/DihEpW6VHObWXgZuVqVBGloNEGUPi8DLv0evrIwiLRbxRaqWlB9MHrI1OeUbBPMX
tQB2qECmvnt92sFe8OoJajAB8kSiel2YDY7XpUyljgzIGjQ0/k22apQXGngKIPqaN+sn4jyrJvbc
xP+eRyl2Xrsy6qJsrehe//KIqH8QakayF2paSFRV39+Y5JIxdXdA5823W8ZqFyXGUGpwuyshp9c4
UNyIjrdK826WmyY4xGqoYhCd8zEpWQ1YtRNMq8VD22K6+QbHMWdp/np6aa4hkxh3JIEyYH7CLdEW
yViY3q2oOCvB/FWsdfvcN3Yd9zKWUhDosw7H8WFNQbziUgKOA5hNmuqo5uIS1eaeFQ8njH5o4jZr
pOg3kxHDQQe4qX9DUqj9B1afvDyRhm7Lz6MQjNep62XFtraL/NNtMywaC6AGVq1ogvA0m2qiwkyt
//q8BJxZZu4HsmD0b9BhraaNgqhN1LkLrUdIfh5ACJuwNZAfQnim6GE9hibncD1Gulm/F8SOtGjP
mmCtobw6qTBmm8rKUHck1Yl9KfGfek96xXGzmFuVdoCRTkOk+yVHbpLdjlQ53IHWpmcHlnb0zvaA
ssqtX6v3e5soA6K9SPAOrxo1NzpDr+9aZzpenDw8LEvy32n4KZLOIiVSlDz7qR145cLxP6Qji3Go
LdFU4bpz13PWp+39n96Ra/WM24Tn0G/bW4J1GSQfd0+WxtjnkRqe7eBVRWLB4ny1Bo8qNY6CI4NT
YIZ6KHlIwcyHft6I9gX8BFLOPsU5t8g2hjzsgxDNMNHWGHCWRi9Dieya97NH9sguoIhO/6KkzVG9
zIOSKG3GpDPVrxbYYF5oEtVHYco4HFR7dHxI78EM3wGXtebHnDmRd1CtW2dIf7GfUt/tNlZNMbqI
SslAo+ywWA/SCcmQuRW+bQoF7tR/ijI9lFjLaDoGl2RJx/kWlzkCuTGq43moz3DP5BVH8Ah46mCW
tI7Jy3dp1IBgnJb4Ig3irxcfQIiEFbmMb0BnK8vnmbgEU8J0+qcIcjdpz9fHIz7Xzeb7adlUPoD8
28P35XBsI5Y2losCVFfTJJ5gDkLNJEyYk77T8uqBdZEvz5kpbS3ePqS71aZnL4k1ptnI5sBLLq9T
Xk5fhyI2k9QmeiOkLuhuWkJDm837FOezFSNvst1bGXds+kWQ+uZbzd+NR+Dz//koXdYTY8Byke00
U793E38Apo4uSs92bANpUiUnXxQpQaxHvm3uRPr5iipxCFRWf/NJvJ/0sg7itZhBwNm8Z/223diF
elL7ArwMUrmVukXYJ6t+3JmlhCbLcVDyBrPfZeSQihrH8UKXm9dzD2yYa9TRIpyyMcsH01od4l/r
9rj3cawT0EnWF/CDxW8qGMSWkX46iErQ8qa0ZV4f6L/06yUFoAr1jG9grpZJAd/PdVm/YOy4Z7ik
JBxzjniPX0BrOwZFzkQT6VJtJ7jdX104xmKy4Xx+3V1HGnKHF7DK2OhIQB9mFdzdgYiDxYBZA6FN
oVtARpZns1yOpjxOB+aTll99zsxob+OqE6cq7BRNwQfn7ggSyxoS91ePRnGhVwyh8c1m2QJRFvNn
fNWCd4Ha4c6Owhc6vB6yTwdIJ5U2y/gZFyGPdkjlZQvBjaPdwdEz4hw4tbFhNr4MXCNiT5REhvxi
IwCkO6LnDIYtW4rkslhHJuvcxZmwdQt2DITgfG2tsFfPra2Ye/67hEacMYBZ9dfrCaDHkvDu6UpS
OH6Y6a9cYMFO0RqTNXfMNIJwElgA25eNNYiCUTMchENMKxaHY1E1XIzOw9kCMgsVdc3On8SvpSPI
y7+ywrRlqCKfu09M2GSpa4UTTJoxP9TzfLLIr8hIgztnKaJxpiD2BtgIuQkKXakCH60eE+XiwdOg
9MdPuYqLUS4BbwAktKFRx217a+Bg0kSagcvyu7PgtWD0KoBV7XOszgH9TTyN7dXxg8LWN6iMt/Bm
kWB7ehR2Zei147Z5u3vVxD5dEQtYo6Ouik1R0xvbfXXZYgCSBB0wWY/O6Q6V1WhFuypIafcPXRUg
G/G4Yk02x4mwn7fQJfNon0Cv8AKpNbzaTLr5nQFz4gg+5r6oMeczjTCtOsVOovbi5fHRq4OGkQmT
Yrj85yoigTlT9lSWzmZv27Iyu1U7pb8GOekpH3K9DK7uqaBZ80N9oYTJov6toRLhTrqivOcAfDE2
w7DJeAVCrPhLPwdHTIqz9V6bm5xZ0/aYIMIDBJcKL5jETbVI7kuCmXt0I4/byeDKggywjgZoUYG6
Djm47QY9h5eugsuSPEwtjkviyW8J0FqZYkgEZudJ5Pv0O2syb4fEvTecmLhVfxhtC3jrfk+ZEt1I
hbZEGjXhmowAjjZDKO+xxJKpmAPnI2EiB3sWsXwKMI5KgeZMCUDHgqvD+FuK1OpJjn7/FBSh6UTL
78pVhT44XgXZevS1QdvpTloRx20miv3XYKdyFgCah5+upI9vkfnsHoLxhxOmH4IyLXmtj7qGDbdr
Yf3mFj4SxitMsUkPs/KtVdutZEqA9BpjtWXR3zI3IYRQUTy/pavvJBvO7Bezy3JfqHEAcT4DPG7/
yQhz/yD8mvsSUDy+wqx0oP8I6K5oTdI3dtyirSOP0P9f3hJjh8s7nUFBdbdw2urA1H3oSt9e/Yxl
H3VqGNFQGaSgviScaFqgeyhIUWRTyr9/QJdcmql9oICM97ijtACXn53++WDt8Q7z6bVi/ij1oy6r
c3eVt9efh+T+2huGXEn/Sf0qrJzmVjY6jB4lPL9COtsCXXW7LBu8m5BcX+1mPkc6Ol8MGeKr1bk/
cHYqU0OEeA9VJ/+NQnx06i+80uU1p3a7te/BnM+hobvbDtTA7p0zS8oi/ns+wBqQZ7xTwmOqX1QK
3htOSFZSvh7wTPyfgPhoIAB24q2XCGt/uq9ZtEDRK6UxCJh/0IXX6TzBwBN0yd3oVmY5uUoMeP/M
5a/dcskRCLHr8RaqK+Jgu+3NgehYf/Sdq1/CraI0g85I7KUg524MCH17xqBQKjIeDItTbtQvEYLp
y/hADTCiwgYVBXp/7W6iKfIbhg61jWqQfre2QVDcsbf9fpRhDmGYwFP+VaI/LXrGF2zDu4TI3rYz
Vng2OF4DvScI3gaZ5bfpoULPBF4V3xNphmvkVyX3hGWh6nL7j750qMYFofaZ0owDa1rdU8aRX+hI
ksjhwo/0MgHV/E3Vv8qpqdS9Xrb2r+AmKLPjBVm6ER4IABHNdGXZEM4dzUtRlDxicaxLMaxFdz5c
OT1gtaZoXEDOPLpV+55a++BSQJ1/BxmN5w37ZdQoN6kRpfGkKKr1oan9H7PtHbqxPu2g3RPjmuat
B6Hy8UjiLsqU2e3ECFH1lyPORs64TFciA1/g55jec0Kk9RbMp7+JnDsJTdUVEsrippzuo6bUWrYR
UlZVIVRdcIc8gBms+mxz3RfVE/ZSPrWoEoszqKvw/5rM8AsOC4o9L9e8uktYaCAewZOtbe1sc0fK
ycPxLwT4nft9UiJ9IddyVTQKTTFGVB/XjjPp73kyEV5UvPU32KRL6vXN/xhp4CtMOqX016aTUFav
Bg/az1sDnkUxrQte+eQoWQR7+MTlgjF6D5TMKTmOkMZ/EEaB6RNUG4l+/03No5WE50oWAdDYHOQk
i02FSAe6dqq1k7Zh3D2fimP5eruyFFhKjZdhsm4XB0E3b42xPoF3o5ddBCmjNnMZ4CFli50JtsTS
5TXs89QRYZN+DM4aT1IVGR3cJRh1GYyXQ9QmpHgTp3UUM5+H513zBLi5fVh5njc4oM44ZYZms4up
G2CeOW9G/Its9LuYJyRYVPqdASjJOxf7R3jSrbJEBjyXS9jD6J1OSHfpayhcwWuIT9/qe0AQ7T4p
5pf9Hz4S0C87OTw+IhIFkdgFSrAxEMC4zz4rvS2u4azbrAF8CZPe4vxBCxWGFYRMzfgkaZ1+dhcQ
XFyNYb3mI6OedTwKyKVCUO37KRf/DmqSwhJfDtfV4zj0qeLdx0KCiQd/9SCjS1tvfg7gfa6UvG2/
y4sj/hwJabP6qN/3mp+F8wfE5N4xroc84dlT0+XcZiQH9JGdl4Mbft+I5pc2t+aO+3hCqIUdMQyJ
gv+Zyq0P9ttuQk9J7vaGRjBvXiX7IN7kst9lzpBoCXajOQhb7cp1TYKG2fg2eM8s+Ma0BqeHNQ97
hZaicW+tKRg3WQSOeAsMFq5TQtzDw8IK4yP2cMNXGYcsHsVlZodOfPy6GuU/M29vbEES2tVfyjM3
LH0jWJ86I0u+ltEbNdiKy0hriR1aGhog6hS5YhVPelDiRMRINVmWiRuv6B0YKnVnBS8jSgK6Yd7m
6/pVPQjJTLVaoTsWoPpMKnPa9/ZNSFa0bn0cDOd8dI9898rYfBMRYqF5FjDMd4jUqP9dmvUyWdnh
0F+LnT3E6nj5KelsZzOEPPdSrGIMOEaXsoqzjB0f8P9xrEIgU1RTcH1xTYYIxbSqZ25lt4qJEg/Z
YhhvBE0V3pFVqq7vqfeIRibhOn21nHwAJefYHaq2aIuHP3yq81GdigokvlE6Q5pjLJyWcQpsvJ+S
L+EdqX07xU5XKcysRhASCm4krmZP0vYD8VbnOvJ/D7rG0HVcw2t3u2JwST77/vFYQW9Xjw6pZ5mf
u39TiCIWBrKetPp6W6faJ/N8SQGtYTDOrohawn49XKOtFWBqyOsGd6Jvlfy9p+gi5D9KP5IJUp/e
EYmxLW+9Kuslb+DfyKYyX1/Hmuc2N61/b/MUFvQ6HiMgDWj9aiMvCdoy+30OcAT77SmdvtYpWYqx
WE098E0BOk3AXWXrn2vLtlp87gRDBqWtCYYysF9p3VYSQxGD1CWg+w8MUvey5sRtPSW3V8WfiR4T
OWZy74PksIBqgSCJl538ECKoZcqRBTILMQYQw+FvUTAPNNdUwfUO4Q5uC7AnbQdcN2JRXdMsGhI0
IpHbGF5BKmPX4/X2u0BCyQZWFggdM7nZ3tcgkdg7Qn1qpnby3XrJIBGqC6r/q10pIap83aLvwmEI
AVl4srQ4VhNu0ZA3L2cdImZIr5PaCCKrsPAe8mWUQxdFYdCMhpgREDox7Accw+nV69bALNLJuD+j
g7MvYf9DBmO0Bui+FkmGqSENDJzlHLZ4k4lb5wups9R9I0MwBouJHBFpX/gYpkiBAo2zSHIo1ouA
/ILsElunsg8vlUp6sgzpQwR5IKxxPJ7TEpgIxNnIgLCmL0YWnBrZuXnNtAPkMQwzroYYhrHf9v2k
t+5zm/OaAkSQ01eKmGijh5hz2eVxR52BS/RIkS3mM0/MuqoaoRoTEj46H5yFMmpNstiO6mHcht1B
UYk7HcJKr8wOZD9QTAx0AUuXwr+Lx0VE4IlxV8p/YYHP61i06RmwQH4tH9tmskL1WA2xM8Th6OtF
V0IL46lURg+cAehnAyk5+SFQ4w9YO4YBSm384Pei0rFx6yWsQLgZRpVEg7X9XeN1Pu8GrWrP21dB
Aep1/dN9TuwFSUn/vkzq6st8Y1SmC3upSPGdCSajuWQAwUIG2ou3w9XJ1dCJHHYpy9fKrlcUx/U5
NId0om3PrNhKG00bRjzAOMhP7Ph5++VSEA2kJ/iMG39eBb2YPLR1aIr3YjlP9nFMC8/kNObLqpib
wl/cq1EiVNid7LeTujX9Uxs8AtxRt5mVYe2sKsKpFWZ8i5hNSDWGR04KPJdCuSpqHPb/UUAnYyUY
Gjt8TyCfpC7bKEeH64bFdKIe+KkhxQkAfMKqQT8vebzpnJxMUbouveJx1y67o9U4zgdDTs4xk2/o
yyuDsBGSAGTZUidMHw/a1maiiC94FC+QGaWkp3XPXNTw44h1fX3DrfsntTz253efxUphcnD1n1TI
FZf7BUZ/4F7+EwifbKjp7dc2NgijfqNhO12sNNeYBqmVd5q+fd3HULPEAiQHyD63zmliERHFSv+z
Sk7GFbahGX6RjkyAJYxNe++uw1GmMiR66Nl2Mka6J4JBWFtKtvz80qa176GqQr+ifFU3BkVdOw26
RXDtBm0GpggBTk3TLy00Y/w15McYoTis4jXpS0uXwo/iOLV1vzleRHQ4siQMy6cq6JrrP3qoFEZB
Gn53fgigBFoj+9q/cdl2Xnh4PzCeex1yqvG8tiJMYxsatyldemG5tbbTu7C6C5b+iFAkQmqPHQxX
hxnwdGy/48KB7n9X88/dZaaycV/akfYugVxPPnlabybltsg87+54YIgutJCf/uqYxDjrA8W0U8ik
1Lo3pXNfbGJvEwDjUxKFdPgTUiexdgYYEJ/EUOE5OmyuCVWjuXsyrboBAV20bqxzfV19aZiyRWVB
/e7EGrUAATMgXBCAxbzWGGmDRBYgSJi3EztV79yOujKNFuUb052Wp0X2LWxJWZNB57qzKQUj7n94
kA2u/v7s8k1LeDrI0CpluVGbO9w9hQbKvN3icNByl3Hyv4D4sYIiph+zOpy/26bKX6soWfSdUCw2
hnuRrIkG8+KbknOc86f0TU1WxeCXAz9yYM7FRuks00xugWCXWT6cU63JofOEGs7lnxqyLpiWSp2m
I/SQ3kzAsEQGxkG8Svfl8d0wMyRL41Zvtmu6UIeiciW33Tz3PE7bHsJyT3DDVfnRHGPCGzSzBryL
I+zR66yRAbf70H/UrQwJ+3W10CsqRDRV/RAMSTR47qDZQJ3EtnizJR/rkW+v8iw3sJk6xaUlLI7r
XwVUOF2/MlaMmfrb5tMkyg9riGwUdtix087Is0b4eS36+rX+CQ4Lx/UlDs3GOJcvi7T6EuzH1NG5
M17ebYoQVQ4ODV9OrK6610k3iMw7GvYIbSkaQSbB4A5Hax1mZfEM1UqSHfWPICfldm0GnG0NBMS8
uNX3ahMsy7aX1rTEC5HUvNIdHPcR3QTpLzteYaRLc1+kdB1xSL6UWU8ZpYxnkpiD8h+1AjzXZMmt
TXu55s0m5u3qZaHW7GZaf6J0PtpX9WSTbyXX2OJniFfY/mjOnjV0uYTZerfM+KgmgSDXUWbGLngx
AZI5tnOoXkUdfCMov4b4x5NoGDW7o4p32mi2cHfvYLZA7pB09Any6U+Sf5Qq8xUDULP4dqF0VWyk
acsor3LOwiJ4z467qNdUHNbjwxjjaUGSnkHLrPX/1gWPwxGjLCif+LuDFbbd0MtPUYUD5wkr1peq
eqNuI7yhVPHTBbQPAAEutb2pF/fA7eMDgMOY3RebvGj/W2id40/GV7nULiKv5UBRonB31ERuZ6Fh
NZgW8WMSOig/Ui1Hko1LnRTLEflQ9LgdE6DUXTni02sUywHSCY9UJRwI4UeHhFHkJnup0MPXq2aW
o1OSp2FzZvU0GZ6+w7aUbrWzmmT+BqIGpEBkaGfX/k2XTwIz5ilaT83AZSbWbbIVQit3C4c91hWY
sbWhjyVkiIZYP6tFmL7l7WoUpJ88hlDmhJ2uj/sYbOFWWVjFl/DdS0XOkVr1VHor3XbHx/aLJDj0
Rl9SRbmifq9f1IZsJMIhCDd3xwO+HeAYfG72MW2TjRH/snKxRVONCtupWLPVNOjYtDJh2VGDhi6V
r6V6O9EFfVTRc5N5ogEq5cGX/ffnd3cqt5X5oxtjpzAI7epOnUuyiFTDg6fLUwPUf2Jd0gT7OcUr
Vy/vo5eGPhOYODrC0UTjUnjksXlYm8r2PTOqrS6Bozg+Iz0J9gT7JLHjoyyaDBBS07mmwDd4FJOS
fRQ/dwDsMV85fugY3zav+//yHgaTROq26SGnJg1ZqzdUuscuNMGacLzohDRFWse1bnhA/S/yeOob
hDoExN9AwKMcBbBcyvRTpJdjhuSpaFCwGcq9gXsZQv0GT7VFiDc9VJ6xN0wwz3SPvoIK9qCoeJa+
O1C+IK3Jc7B95e3bDhjOxQTF5YTnkyyYgYPctFYrIR2/TdxyOm0B3zh30l7wrFL6YoEag0/kUraD
Ap2b6y4O1d68wD3iBy8Y81V4zuH3v3FlpV76V3cezCpydkUQTrdMEe7ZL58rts/BMFgYEx4WZXAC
MasNKOREfq9PFLhncvHTW1CkAYtm4MP20MsZRQsC54TctRat+jOqPXhuZohwZygtIxBjZJDnJHLn
2LW2XFAvpxQoup9yQIxegawbbZx8ZkNAh/w8NcY+CHlKNOQwavVSQNhsXnEN8Ntk9sEFtyG2VFcn
JnXzit/tDR7y7SV3/4WkyMqC6bTrqoUrvD0zv3iSZ4gfHMMNcxp92kG3psf6UJQG2gOcmIYv/x/v
xqdmLT+ciPEVP5oTileP2SY/0zdNhGfbjQvck80I6wBCPPlOEhsYW2t5xREHxWzn5ULGQ68nhVMq
qUj85dThleiuVVVcyKdd8AaIW3bCvc3BuxoL9v2kFyRnYV0GxLhGmbxdrUh/kPVCF6oK9QiPRNTd
GC1wbB5H348braHvwTzjNotXCYxgP89xvLhgGLNuRt2eD/s24oz7KvNq0L3HMquUEqm7UIj2/AhX
zQlllFd1rdQxXOCjibN+W4x4tu2AqoulUXmJwR4hQsFGYT3aejSjkBMLbYQdmiU+HFapLGB6BrTR
dWX4Y2a9rUlFpnU+1JUQNKBNcK5oRaIErkd9fUBqwKZVgL8rs0Bj5d+LqeQM92m1hxZPkShhb0c3
pl5IavgEVYt9Nk1918HX75vnjx5V8duARRNUPgGmQ3HGTWNPceXi2G62JlULBIqTlp7peSKLr7hf
eaWzUHjjaCUskY/MJojQBVfIvOckK3ZyfkEECYS5Pq/sDyx4AjvX2H6bhYvAgF0jG+8TTbCsnKbi
Bka2b8G5VxvZi+ZSyLnQaanf7/43um+Cxzs14MnS8IWM9nihPcT2EZvl5eJTEOKbMqGeda2vR/Pn
PGTzc55zIuuUwY04LS/qZZqOTVVT/JLBolLF+Mo10Mojc2CXrxPE6yc3waUMp3m4LXM5UDJ/hKB9
VL9JcRDfw4BzRIrOgkmN0p5tW818J0JnzC+6dK8iEmLebLrwLTsoOiv00DCqzA6urtxapTWaaJIQ
YI90DCP4k4rXHctTQJ0QOXCx/9hPq3BmkFqLtz6kt2K44bhsdnvyfnHc1HZFHUitPNOkyltajsUv
ZnsorIUUnpthGSELnQZbsOTIftTS8Al+PgihseNAuzVf/jWoHd/ubdmgtc545CXjQV/qr+F7tz2e
YlBCd32Qd4zCFgXcmur8SxVYENI4DIMntUXDRDqI6K8fjjkEBEqo8NNFisszZsHZYbiWPU7LwzfO
BlYGPucBWUIYfTZ4BDbbxg8pL7ZNKofj3FK4ZDE+ZMJRXP5fAIewcL5t+tSpwpdcHAXIEE9zu/SN
T6xME9xRrZHMvtBoB18wT11VkN0pwMiqz4BkJmnc9hq+kWBt5t7SBXupPuP6VnOS0LpZYKyu/CwY
fiMXxtgNY72pFD/MoYoy5tvwtgM6zEY+U1uDj7DJtoN1erN9B5LoZ+PEBHUArQfuV+r9e0QggUXk
ofSLd1+JOINmsUakAQ/0KgflScjI6qhbOvwjtEwTqtsNbLhXCgYyczJg+GJaxHMCOKAkfX8IoGdY
4LCkTGpEbvg3TI3MTbtd0Xb3yEZDCWu+6uVfdbh4Bp1wqcAFsfvGz5ZmnSFOhxNoRAZe8he/WfRF
0iFSRMpeDlg7T9mKokY3MQiH0YbGLIakRIi/e/j0hztzrgFeBxkoedKXZQqbgiWwQoaPxyh0a1eM
Y0wO4qo3sU7hpdjgl2mxr7dnk2XGlDxCQJS7Gq+VUaEU89o/DtNtIWflH/eqPbuov1rQ5+BqDLbB
96/tIbpX9fkdQqSfPLKt1SVakjT56qvRNvpIh0PjaMU8Gseoyzh78j2Z4JBiNdxXgAWq8qC/kKWu
OVXRqgyDwCfjCcviij+WDdQal2a8bqzEqNBxmCiSw7iCuF8CR3NYqxeMFYcB2EvnqiiOwhafAbEo
+Jr86Z6exKyKjbN0ycxMuRuns2P+OoXSrtz8in/JnTL9TMw8IXRpsID+ZZAg83rbgOP6B9QYkXT2
6kJCX1qBcn4FJmW3oHI/uhPrRRr1z99k1pOtcgRew/MeJVImiWbfphsnj4P3J2cKjWcJQkM8S1zd
Upe3Jergy/5+JvdFTmsa45lCqbJECFELIAFt0sMpVdiIXCSs6DOBKR0Z29JOWUWufCueKYvWmFNN
ZESnVfEQHM1dXArfLQbTEocZXCt6aazB2VFTPLrztBHHYNOY9H3AO4g8r+vgZ9Jfdd4F+LZix/ZX
ugLyEFEYdW4vY0woCdqMcpsT+Fn/pHnoMJ2C24lZSkEoUZckepQmyJQB1lxnJdMPIih8YQbFCudp
Uv/8N4yWcntw+YA+OATZlfQ+gHUw1Jijew76BPbBSLovmKQ3gy9yo+limCOv9d/SriVr4tdf3Zde
mJcgAzT5aDkjD8nOyTvhwh/9WqJnREmUDZ9xRy/jaLe/LXhguW5V0Hl6m3h45Qm6EzdOOP99VxvK
e+zsOVNHpq+DFU50tJmAgLzodrG+nRI0llSiwYwJ+4PcmN38dEcNeFP4rMeeLbq5xjbFH1NH12lD
gGYnOzJC407ERNqgbr3bEaS17rdY9CHu40QR24Fg3bEqVX8geaRGa5NIaRmb+2e7ApovxW6tDKyx
aCdSRZmxmZLItBe43sSv9hMY2EZFOcAo7IK8B1vRbzEFIbT+JJ8hl4f4rOiUUdSEpOuMb8SHqMTZ
NVaBjggbp/aqJeD+JGZB4CYWNfFHSz5Iu+pZsczSC1l6MfBKDR/KmCj6jnjUwwYET/FE7MThQR09
DQZN0LQmc2a4bshUX1PhBnJKV4MHe6KDUrjCHliVkoepeT4AIhXZEgAkvH9YY+3Ahivplq2DmrNf
V4OYPcozeOIx6msqI+kav7OAonzKZsu17I0WFU5zFoALJkqRKfZaLgXUQLwobXXCac4gzN7RnpQG
VKwjH8BwNaMVXwuyHEWXziI0dsXmjOH9w69Czmc+qENjG0NRdV5bP96i3oGaIndA+U0ZDQ1erO2f
BJ9rmqPCrv7OFBBTVhFEa/tadS+dta/I/jC7CPmxqj/Dar09YtlTCPYdxDnYk9tiI1XukCn5Ff+o
uH4krJ7XfM9j4oPT5PilUqQaICv8kBDzI5SEqkq87ahAMTMob8nGo1pFbcHMVQeLyCduN/o6GUnb
/J7WrcXJiEwrWztATBuO9Nd0sELKbJQZslGrSEpTmDAJZ+PrYzR5s55o4E88mcgbk0oY1dsuPFy6
PYTFMWHMxAx+s9U6Z8qcf0FL1yvddVUHwjPq2YDUHtCAOyIGUi56Z0SYPwVgj3UmHniEpfEJ9TP8
NM5b1w79oo78h1opK/YiJA4/RjseCeJt90Ifa0svJmBHlOEEeqDeRlpwYteW1cTGpVRM1Orc5df1
VvJAgB1Rt/mNWmfYEbZ6AqiQCDZNM7ZQiZRKBgA+iN/zwWYjOC1OtlB6NCi1SqPAtm6VQUar1PjA
rw65QNp1dPgLPbiyE2REshg5s1cQDWXbexi1bWKG6TYCN6LBfsFzBK0uRPHXRJ9poyXAK20o2pku
kHrLCbDRT0TpREKCjOLY07c84t9cyT/+EsNZ7ed1kk4N5ShTddlYa9Iqrgl/cUW6lF5MKPslkgug
drMvwB9ZAWu3knfbcqBIZ/93190Sb7rnBJIokXznlIDpc9AHvySifx4vxURiAGAK5bF9GijKpuIe
cRNkvaioS2nkUmJdpXpldTJRRfE+qV9boVGjgvF43hPeoXqPh7ac4dobKip2+o7LcyyuA9lnERrt
NO95y8QXPX2DS0k+NJv36ociO+JtpkBJ7/Han3sxN77gqkJJVCQY3s822m4e7X3s/PsSOVfBr/+t
Qs+j/owqAnaiXLaGaIMap53bTJ13DGVAw4EWJTTc3rV8rlYkfNDNcCp3482AH/rotivEUs6Puq4X
5jyKFZl6PZhVkqmRH6Zs4i59YJTWXJA5y0kz82knhSMNVLWVzApeOlVnhBnZtUTztujDPi9x999w
gBVxQXUZqS6/MQv8dYT4T8NIRKOZoPeWpIl24cRHQQsNQ3Kz6MDBQQQF8WgrcM2dUaoC6zS/9/gi
PE0VVME5SPYYy0S7Ag3Muf5NH1COPaGaGNmwS3AtSKtuS+ZAac1yXwKn1vMIISOY1bcVH54FKaA+
UqN+d/NCuIYf6UQry7jndq57LEEpDwzVPh1/g2hqErK/xCsUK6ixyH/YKqabs7izsYF3i5FpLKtF
uWIAP0KjmzDTmf6nCAMNAn3nle1o1KslOtAZaLKckAGu1WHT2pnQDOTAvTzm0EfA1AWDihfrouXj
x5yL1GUfmvGnkYNAsOHGAKY79gjxltdeHynG7DAdlwJTpos/nnTZLVXC/zzQo5ZSNSeZLPM5rqZE
vGr8aDy+lzWblEpbztWUMOxrEg5xnzha
`protect end_protected
