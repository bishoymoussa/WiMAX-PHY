-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
EQHNPOFv2cCyclxWU41PZe8ndkxDunYw6FQH/qBUdQ2R7cTjjAj0KQg7Shg6Myvd9MWywFtGaq0L
ai8o2b/xbcUVDl9G598HUioVJmEbbNdCCiSubcB6LSm/YYxKO/ptBTjTwa9vHIBmlfkleokAPMBC
Es+7ZVa0oGWXNDgrDsg5yCviBbKSxHWCN0hH3oRrPZRAxZgLGf3V4FUUHLyJSaEp2L8mE5CNU5Yl
4UZvlOcsnnpcqvhvoM025eYF7aOSnw3V7miEScPKl/b7mn4ynxbJWd43bXRmwd9vv1wczY/Kr77f
I3lra9Qb3nzqghJ3lNc4eUt6XzkFcSwhlovPoQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 2736)
`protect data_block
8llBm5Uvjws7XEfATeiILPxWgPjl94RSS80Q7XLmvMmRwJyVsBObA/0HbyKKTT7jGjml7HUl1g+U
p5EBA6eWEQD1x9+uXPmNK93B1lIbMzvfS8gIyWQS/t+TxMEjbGVRMiCuJ3KPEaTwpaUkXUJSaTmf
ysPCd5Ls3MZChqLjrC49iUXOFWBk361z25N/HjX4RPrNkdHVmBS8w7VaeAjRGT3myg1rlS5qjYh6
TfvxOaFntbKdXD1wBG/mkcXUOx4ltZifIVqx6rVCrednppIKFvndJSRCKeLjc/cyylRU9XDuNmsv
VC1EJ57GGWlUVy52CJ6Az9RHwXtDR0PsgBN29S5iyqsBQwnVi0RRdZcEkaQN3blaWcomWkjVre62
wQe+8KZK/QoC7UiRwWzGO+yEXMmykASlKb+3Zdtx9YWBaLUV4SLhSEJTvE/tJB+Z80C1PfpCeAIK
TSsK+BR8KP9ZJpAc4OxgQ0o5iqFasPfgG3ZxVREXmwOXb3/b7yj/ev6pnuUlk7+OVDKsO566hRPD
T9lzzt2O2spiu97jKwZjMp5ypcsgYYrkFD9LZleNRGr+3391+sjj8Zs2gZoh4z7Lbi8miG9nh8+f
URhFCz5cG9fcn2hw9jCXgcTDNbThrphiSgzs58PYciEerpPiE7LCjwEi3u3Dit+mSsWunKpnoGKW
W1zKhQD3r1yvgxuQV95R+ECJFmLqgOJpl0YUm0FR09BdXpIHRUPTjnRmwGNcJUv1AqD18wAdEq4u
++O4Q3eNGHs4QvyS+RDe8IgBwzedvS9/me+Fvk3ekyPj7nr21H/UgYMCK+w+VvOzVuVpj/EqO17r
GLot54N74JdaBTj1uMnErmbqCa/jeEd3MSMsW9GRKFYG86oc8+yiDiUlAPGIlRtX/6s55sAcj+D7
H9RnhdFKU3SIlXxBPhJ7uBV2Y9TDDzMoLHQjtmuKtPWEXBfPNYlx4wJ/L05gs19VyIb48VGCrxci
q4/Zm6Buc0l91SY/lWW3PEDjQwBTtW7eMSBQQb2VXuJfpAsMpE5g/kvYp5WP1wrFYfQkYraxatz8
C/yiXXoISEpYpQArKQRziE7vs+4/wTVSQ48uNW5+8ZmGEAve8R5ILXsuZSxu1w+QDKaD778/h8hS
RssnqRTIoi1Eh1KxMK5HqMDFK4APSiyyCSM7VO/x1UunDjvakVJfumoTrO2J3+Ctq7VNbLW0vobT
C9h4Fi9uroIUMyM/VswupowJAlZOJfaiv122Q3mzhewMnZp7vBMSOL3h51kEchkfX64T0VF8lcf3
B0OXgXgN4c4ck7OetTygJgqWcyUxnfzDxgFcG6QVdPBUHScUhnm7Uo8FUKUgBjaLVScvQLpipNRw
nnAPIEB40RdD14fQ++qwf3w8ZbbcN9aXdAQ3SjF3AqjZVq9/9cihv05TitT9AmodBNDA9xeSHQZQ
rXfLFMfL1XgppbmabDf36/XbElBsHxphKB4mQ5ueFch04k3Meqj8Kh5mMKS9do2FQphCU6O0975S
2X2YTL/t3DVzynj9Cd50o9IFQUNFNIF9Dmril1ZVFaamhJjwWSQVHjtyqH4tIi0nsx2rryT3l127
K621wSPDPD7Ws9q5L5o9SWj2HqEzqjFfVBl1HwzKL+eyLVn5Cm64eFn2Hyav4V9jIuyp/xVLPYBa
2fcnrDe1Wji20YdQZsySIoFmp+igCbOmxm9e8APjWVLXFFLFaiYesYINXfJQxV08H0uc6RxHOahr
FharGxPn9dAzNIwtrIk9HaMhSX2LfrGHjozuyp9zznb66Wv2nJuHu3634IsI8aDOG0jaIDS3/aC1
lQy/h5h3/7C1fpRY5VH/7slFQa7Q6rTaJqjPmIMheYMBtzwmNELP2u0wBHPTAfpM7tyO3Tw5if6I
xx7HMcH++RjF8z+qzSKQECBZl8J8AwhVAl62COfjV9SsWZ7Sw5qKi48ui+14Mc77tFQM55SWLroh
uWLhRT2PgjbSaoHvDWF+VUWI0mAiO57pugthkdGyUtRGwbd/IZidy3AItPgJOYWfBy80x3OrTuDs
azU2SXX72xh78lLsPDOmNIVi4Eg2lXzTNSJuB0lWsJqpX/2A/magphYKb6dkfzmVCLatSPY1e3q+
ze/hhY17N0xKazWdL6XNEwAt/CiYZ3+ADz7KWmiveM8kRbtcrg2Pxnm8aqkWG4iJBx5E7vFfY2Pu
4RLPzzAtsGPMIvseJmyy+zdBZbV/a09AhEbmGlYeFNHWRcivJC/hyUEUxCP4vs8lXIyubcJymMzc
0Oh6cMVGFy9WqGKgVgKfr0K9tByH3DL0K8PK8mMS31psf0XKLOc2IM0sfraN7ic6XUVl2xhgn6C5
r1EHkM4bZ9AIWhAXmnyK66NG89Lr+yVKa2nLy6SEQ/DMiArB9FLWBCztSwpRav4Ofdx+RR1NiqHi
xTUB909L9Nig28M6TEUdNPWOAdhz/0pgylayDUTgiqw8oB2VoEBPHKjST42POlVzHEKORaunuBlc
vWtEQdcih5+5FwmgshERRYaccnt8v1l2pTQ/Bp8mzrOMRbfs51WZDs+8nhIhNb9efqahbZLFljNV
U5EGqE9yg03O87wLtd2OzBTjXmq49hgiavD3l3rma8g2OKEV9zD9cVy+SFlGhkMOeuhq9AstXazB
re9EWCdPJZyx+93aEiJ4eyWfK739NBp9tZGVSDRYaCOM9ac1c3YO2uXSxMlVTjBfviWl3Z0Z4ijj
iQzkY2QTM4td7pukCOy+aDWSXV6JqH0p+YCCDwL9thZdEuyqEgMMK2SoZ8w0QYiqt3eFXug9MHcF
/8/mqL9zUyKEcFYowSgdjvrQk1hN1X5wd0rR7wjcTyHeUuhL+WK8Nc/aHl00wBQT4mi5nsIQxXgJ
9t+qXidy0bvbqGDKUdv4lmEzHfoKE0l+ljmyg9fuqdNreNldNmTIidgxgTOz89XQbMvYiPsIAYWF
J0QvnoD3MejliuSmWWluqWwmHZ5XLpJ7SqCwUibQesRicNLRcvmd6Mr2fkbuYJ1wgr8CdaZmdWbX
LVvfD2+BtKkBjXpZMGvARChDbHG/UizINqSGjM+EEbm+tCG3IQaIu77pF7QJsPGL5G+B805NDXEh
+6UmRW+rkMx9JEEcx0VbhD0vRSGF7wlggVzYXfaFcBeXiN/VGsZceMUDNztWPMGviBjkW+qIj0/i
OzYXHkp6oN2LcYOh/WRTI47vRXcZyFmfHbZVlBPaBgTSpnQgLpqYgzHSqurB06bO6aNuTAUnyn8l
QsAPDQCH5d5cpqxOSZlbmnoDERqlAWOinPs68mmOtMEV1P+ebsEMrcOgTrum0FLatFDBNKKj724b
uhJ8Dm1R3+RczewCg6x5GuOnMW7+baHS0Oxgpv5Kxd7YUYi3l+ZtpfczILOQL5QKzaAwbR/2Ditc
gcGg1qWaOaOJA1J7Vyk5sv+no72mTmaWkBJ4wJg+d+eS+UO4ai/G0xUBP+hsBAkjwb+hTjYm2sV0
aPAQNdnErtSNh9Ff6ZLlwX+mEO1SKUg3ntgmqTi8TI5OBxOsx8DX8rxpAxsV64J23VBBi0ZUYs9j
SATdx0DO08ODDMOADYtTYZWU+G1rFtSE63lbzo+yvvMVEIVhe4IsMELXBwLENS1Ras/wzEHRW2sU
`protect end_protected
