��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$Rx�y�<��wA�*;�x���@�̦�W�X�fa�M-$u����n~�%���P�$��W��kYَ���P7�?UMfT��q�6�U��k�>����~�\N�(�����X�e���/6U|)�X2pF�]$h���d.���9E�	�IN�f"�\��e�z�y�b�����Oo2�?�qˁ'�͜k-�K�P|����y:����3�l�d���bl��ˢ_�d���kx�rq�mh�MذM�`aS�.�DW�mS�9���Y��+�>��!��!�T�uOB���,��\L�7m�O��W���6����'���j)n_�I����2:��$�K�2�Sʫ��l ��!���{�l����.�j4�	��很�̢=�����N��s���s5���_�R�>����ТP .W;������	�"�מԫ�����]�#7@O+?�⡾�Ԫ���e�O�\A�	�ͼ���ƹ�d�	@�nQ˰��E؁Bf���|D_�%au�-�'���w�*%��"AM$w�*�?ZxC!M�ߺV�;>%�A�0A��g�%��|���� $�B ��
��k�~%J�� �~֬���u3j:+�%�A��	]�,`a�d��e��nBL�_A5l��y�]�4v�{Q��f��[K��i+'�)1�O$+ ֬>�Ŷ���ܝlR�>73��h�������`���̌��w��ry�Te$1�n\E����UW�4+LF(v�q��9(��4���Eމ �1�Ѣ���)5���I�SI�pE���tM� �L݅�I+6O�A����|K�++����������aO Л��HR\�j���$���)��*�v�%!�T�tW��P�cDs
��Xn��sk�\re#,��ձt����i {8����>�J��z
6Ɍ�gt��{h���T�-��3O���|ػ޴pE�55��5V��3�J��7���q� =,e]o���S�+k�=Ikb�x���RkH3n,�c�)�{�Y���al��?VW�(.8qL<o����6�LV��RJ�
��P�(��!��{5��!�jbM�x.��`7�2��,P�_H�8w���Tb�Wͼ+%��$�TKw&�4�]�j�g���
y�¬hE�fw���S�p��ԟN�Ʈ� �\�z^-cV'�c!���FH�'uB��HP`+<��rJ�������
M�J��E\LL)c��i�����x�p4yxpغ	�����;�<��jX�܏�s�"�6|����1�h/.^����B�sY��$�"�-W��~��i�#@yۓ肖���a�k�&3ڱy�o1�I��e5T�t�t?�xe��ݑ;�jS!q���X���OL��hH8�7�����1v(>�E�evלX�.Eu"�J��\A�O0��>[0�>�f������(��+�#��^%�[��GF�?���W�M>Y��pv(������Hn�L��4 �cU�[��$��ݱl�q�� � G9S�x�v2�@��J���dn�
|{�^M�%�.T�o!0��������ܩ�t���>��3з5�u����r[aQ+|��6)�)���;vz6��P��<�5xS�qg< 8 0L@*���Z�,ҋN��:(��.���E4�e�v�]�}Ģ#�V��\yzGH�Y���kY��\-�}�ǜ�LE�!�\۴!�%��d���ul�O���;ـ��[3Hc*l<R4`�1U������c"`��X�fmy\|.i��+�f�5��v�@6 }Y��1���-6�J�%(1|4�� X{2��vR�%�J�xGzSV,P3�Ɛ'�B�I���f�����w}��k��,�@8k�/�؊@0plƅ��t ���OiZ����3@���q,FH8g��T��rJ��ڻ,���#�}4bz�qz@4���y[���K���;��bڤ��|FU�*SH��߿&�ڝ��+|B��V��%KCʱ��(�qV�n��uǃ���ac*��ݮI��� h�l������%T���Hv����?���Kl�Te�/����0W3��0�RQ7bV�A
�����'G"���m�Hat[ &������W��\^�)�_��?���C��s���k�Z��漏�iy�,o�Q�F�p���Z#�q(]	���P7d�ݡ�6�G?x���D{b$_�K���DL�/"�:��!G���Oi���
����#!�> ��kF��x�?�̅��W��@Ă@�҆����C�o��j��s�L�Oa!;r$��ϰ�O�U��n��<}B*оT<1�4MK�G�#4�q�R�d]�����8܎�Y^���F��0l�@嬎7�|2���!_ �A��s��-��+�,^de�.D�{�W����&�>yA�N��b����z�SvnÈ�(0�9�ف|�VB�ሞ|S�M��n�%�G�Π�������.��H��,WU��R�o�@C�I���s@	�-��`yB�1T3�yƺ 2<��:�Y#���["�'
�:���>VL�����0^O��P�d��Pl'�*Dp�W�s)����0�Q�a�HR?�]��g���n�L�>�����Sv�&�1yKޤzD�z��y	������t
so^jw���g{��Խ�m��njG�:+Ł��ʃ`0��6���IS ��o�t���zN���-aY䯠��	ԩ`\h�8�q#��DPuy�(.j���K��&�2L��Kk˾q0��%P��i�ڬ�:�T�I3�M�2>~�
�K��me���	��J/Fh�����$U������b-���5�-���G��Hl�V�9A�Gּ��cp<ڋPM�h|�� ���0ߨ\f�Nѓ9�J�����=�q}�-�<����{�P��(>���?�K�r*�m���ˌoR ԸW��{��������o�"�z[VD��_�uM���:|���3�*q�
�@~KVد-��a���!T���w�������Y�<&ә&�{�J��#:s0��8����;0��WF���2�2��L18�2�K��l6��5�2\0h�6���BZ��T,&	��l�Ns�Pwi����& ckK��K����3����2(�t�+��-8�m�=:>$���!"/�UC2�yV�A�j��������T�ȋ���x��g��3n4�G{թ�躴��fBŤ���\�*W�]�?v�N��R7�L��< �9�/�����b�I�e�W�G����EI��u8�ǂ�=G5�R�ʴh�R*�|_�:�4����J�AH!~���=M�̳"!� ���!sX���۠eS���t���eu�|�h8�6�[]�Q1�@3���� ~BiwZ���
��	�_w���%�q�ӣl�j�p�T���)�"*5�ka�Ԣ�78�v*�,����q��H6x��Eu�|0��V׸y�N�60�H��L=�ݫºd�91W针��["��y)	Ӿ@>	���x��1�:�۹콷���r�จ�Vk�&)�r_��#�|�yI�y�'z偻~S������⏊���MR��(Q}����ʍн�»���L��S�ڻ�c_�̯�nWJt�Q~�+�=,� �S����|������@*���#�i�GK���V�1�H���s�[���aO8c��D��o��T�pu���p�O~б�|{K>j2�
�WG�34�8����B�	H� ��);㩇�6<�T��"G�sX^Ң�J����6�W~7f��5�ݔ�����!u��^�[��>�'�[mpi�A�@���g�Qà"3_�Qq"=t^���x�� �y�X�t!g��x���y�e��?%n3X�q�6-S�X(OX��n��.�~H��A�!��2�J������VP%-�nt���K������3i[~��O�}r�!?6G؅2g�l��$.<LY�1n̼�+j���s	8��f8|��+�bO�-F%��[��.�)�l(�VX�! G��!��t��\�Ʀ*
�T�'�Kk�\����~�;ܹ�q{��~zg�f4t?��9����$�2v0̮Ε		S���!9���T ��Fʕ�̭s�M�8�$�V�90/$Zՠ yV�ghi�v�j���Τ+7�*o�nбaV ���#�CA�X	� �� >�X���mc� ��{��s�d����0h�|�.��g�r��4Φr$��*׀fd�8w��ַ���Ֆ�R�[�;����AE��#p��W�^�ti�ђk0 �T�q3�ؔ��vNG)'ή�{����e-~Du݈�GO��$]�O�6Z�]=R1SŠ	Q�o�;�PQ��SþF�1Y����Т|�?9�E���g����
Z��Gu眉vދ�8�8B�����O ߆�>y�����O�,r��v�.]������H�n��Wr>�mȗ�^9/!���|%���j�pv�ů�~ʃg]�-�W��oܠk���.�����@ ��[J�{6�p��-�6 �߿w/f�؁����Ԫ�2�MO�Ng�� ��OF����	˼z6h�s���@t�-D��͓c8��f� �t�R��Q2�k�8��"~��N�d�F��8U��#`q��y��0C���h��|x�F�����=`CƉ�˃BI��������]�#<8���{+=����Vm�+T����mԆI��o���M���.�<v LnF�;[�iTC�VQ�ť}����s��l3J��*����y��b�q�2^~�F�:�OB���|�%o!��l��y^���U�$��$��f��Q�Vب�5a�-�;���]+P���bӢ���o�08�S��YŉF��3���^�Vؓ�o\�?/�vv��*��D�R,P(��[9�?c�����̳4&�}Qr�ޕXm`U7hs��}�Am���k�M��:  }��g�� i�FŶط�)�HMK��&B�2[�\�D�7d�����������ᖝ=��wWL�X��`���?T�!/r�/h%��w�Rz�G�L¿.������Õ@����Э��P�Q��z�����O#�._�ޮ�F�`8~��a���p���\�о���4^����ГU>�ą�I�_�;��M��(��.��P��G��)���k�T�������/ZC��r�82^�%����	*h���7�8zw�/��΅�4�#�NA׻7�^W1��o`iRnp�C+��͈��K1�:��jѼ��՞+��ƞ��J ��W<�N�U��U	Ğ�F玔��PF�����ޛ&Z|��P���[��઀H �6���w�H��} t�bS"�9�Ƃt��w��+�/2�s&≋�ˮd3�,�aN^�Ԧ���0�s�0�0�5���
�Jp%/�*��v�1��3Mv{<U%Sw3=
���}��!_:~�J���ֽ�ƌ�kӷ�P�l݉,%CT��	c�[�mn!jDu#¡�TH�	Y��W�,�+�I�I�_v����c�]rnc����,�2^V�i�9��`�y��FG�!�/�Gsiy�4R&�ܑ����3�y�����P��c�+i[����1�v�f�!�^������Op;�N�.�sEN%�i��X�@������xCn�QU>��s��b��(H�@�>jZ�#�D��Xq$Ү�#��}�V�F����l��ĺ�]�pw�cufqc)@| ��/D�hDaؼEĤ�aqT~#6(��tL�w�1�t�O9[���n���Һ�����Y�ޮj+�����������M����P�AJ���ݖ��1c?��]����b�4�d��j��d�C:@H>o/�)�L�)�4|����3�k�XK���u�e:�����7��Sć�!й��)�vk*��3u�����ț/O�Z����#\�8Ql������yfCOkr�VUѭ���B���\F�rk��.��N�C��ւ��n r7.��D1��D��:ss��}x�3U����M�Ͷ4H)	��Q�����xQ��g��j�)���v���௓w�})t-��q�4a;:������&�P�q��X�E,�����S뿩�>��_���{�ɸ_u2x�1�jD���bʄs	�{m��̀�������TR�]C}��f�]l�61�����栐8�]dLb�}�p��o�R�mI	+V(#9FR?͎ŧ�rt�^���1J������.y��.Lz�k ���sO�lI7l��fSD���zN���s�q����c߽���.�<,�����~@ݱ�*�a��[�����^��a$ڙJ��gr$Q�g��kޯ)�|cX�M �d-��ْ�ٌ2�DGxJ���ʂ4�W��6���C���vV�O��!����2υ���o��ν���݀M�����L58 �\���־�C�{�a�K�ﲸ���:�}����^:��l"&c%�m���NS�ޗ�<:����!�8�$J�$��w�����2RF�+4ճ�{��M9�h��v��|��������]�S��̪4�,���Y��D.��#L�gsX�A�:+ k���B\G�p�[c�/z�XQ'lB\ S�z�l�t<ݛ���,��#]��0��T�nI��~�ehZ��4��R�@vkekK��e�&@�)�8��[6���
�H��s8�����-��Jغ�Ք�dG�~[��Q�8v����E|����G��}���=lJ��C�G���ė@5.>-.� ����ɿ7t�k,�}����.Ҟ�%��9x��u������>�0��(
���A3Tl~��ao*���� !*$��&|�,��k7�-԰P	!�8�I��#*���)b�R"��A�k�"QD�܉��:J��� ����r���*��7�y8ā��*K|�%*Hܩ�Z
'��"EuB@7�KqGN�>��p5��u�D���jF{�~Ԯ�.���^e��]4��:�S�,4E7�/�#zʵ#��\%�ųrKn�HU��(��˘l۸W=��T��[$.U\�T��'�Y����L����n�H:���IK��w����p?贕���/P@�]~�8T����$�dJ������Ha7x��SD����/����˛���W�W�����cQ��Ox�� 0�Ũ�зس��8=%P@�g�נ��U0V:�j����ni�1�|�*�C'�VPO�P3b�f5l�S��K��b�h'ޱVu�D/� �csGϋ�Ö�z���sQu��U+7����0����J��yW��O}�l!��2�E�l����e�,�{���m�%�|��Ji���.�����{v�7���j$�>Ru���!�lv��~��{!�'��Kkp�DC%��+�S��%}��
01[�R��x�/�Ef�.@X���$��|��AX��[O�E���L$�P�8��>Q�~����x�wt�9@�!3��4�}�k��>�7f@U�� �H&5t:�x�w=�A���耾��k�Ҧ&��+��t|ڧeͤ�UlS7����RT��аaE��cZ�9��1ҧ*I��ϰ��w/]�x�-;1����:d�CSjCB��s(���\�sy ������z�E����',����U��D�63�1�zsճL��Gq-,��9���n��p[�tD���H>�:��3E�J� ��iE4I~�%���T6�z�F�J�lf��6�j�yp�!�DgVu�"��B��t.�&<��_Q2��k���8�2���&� ����8�ێ�n���l�o��p���@1�рspЛ�L�cV��1@�1*}?�0Aj]�֮L�� /$>��k-M�=��u��%�V@�>�аa���'��P��n���\M�-:�֯@�}ssE��U�[Sj���C�+�)�ѳd��oғ�Tbf�܅�:���ټ	��O���p���1h��#��[��������(�
0A+O�A���{�"�Ԫ���)��U/!��^у�r�h��e��Kx���j��v�F�߂ �O�Q/�̟M�9a{���#q{����\ˆ�dt�u1.Wó�p������l9
(^�T;t�.������錵w.AB?ɇv8>R1ku��>��~��	К�@���BG����(!�2`�ڏn4�!�<�}�m�iP���O*4+s"���>+�0����	M�t���܈�7�]$���jt{�"TJ�STLv��|�@$ǿ.8e�!S�vt���g_3X|�Lx��,�Q�!��G�9b˘��O=�Jv�o:}�fы��wQ(�P���0!Q�1y�)�>K2�{�K& 8=?���൏)���^$��{���hH|�5=���U��^�� _�b�J6��eث_�ym�Uͺz�݅"�7�i����jc�!���1*�~v�!<H�pT>O?��ݭ�2�W@+g(�P��b򰲃ef,L���3�<Ow��#�u�x���q�L�!%b �`LC\��㺋�jdy�c�����-y%W��|����ç�n�F�U�ؔ)�grf���׭���L���`l刟-���*�澌3���3�U�BXF5��M� �BN�ziFub��/�i�`�
�v`*R��+z:���ʽ�\נׄ�Ws�\����&^�4�4&����>�gW~�ߟ׸�/>�
���q�d�1�`*��膯`rCD�+�Q�fT��bօ� ��׽r�Rz�L�N��r2�
P��jV�%�U�{F�;��}��%����D�e�(D��%�R8�Ǘ'.v�3�s�ұà5�X��wW�N6�wX�˲Ӱ��W��X)�f�������>.��������WkCQ��m�Pj�KlnQ�	�V��<�si����q
SQ�5�$�I���waa뚵P�y~\�5�DM����s���%0�����,%@P�O$�:H嗚�@i�P~Sg���*@�޻;sB�E���'��N�rV���E�gp�p���[�Y����{�"DN�l�}?�����LڹU�X����#���ctE���V�)\AN].�~��g�n�~OR
�9-��"��#x�a��ڴ�+������2U
���#��\�`�MP�٪?t�p->E.W�5��:Jb����発}�?]к�2��^��{x���3��g�-o]8��K�]�ΞV�gXbˮ����Ŝa�*�sfQ��k�8t9�C:�}V��xΓH�^�.��k�{��];������,(�����P?0q*���&v���	�~�V��Ol�>(C�u�^����N��5C�2�L��o��'��/6�Ў�9�j��4)���|c!�ki�N�L)4~SU|:x�=hV[�@�&��)�Y�;8���v��%��~���Ē����ì�*������C�)��Y��D���1<��=Iin�a�{�4�Q~%*�7+Q�]�$ ~]c��-���m�yxp���0y��\)b��YU@-�p+��z1�e��r�Rg��g�z?y[c�>��ч)x��SFa�����x��%w��d�T{�4��2��l��q��OxgQ�V1��������]�����j�I��48T9��{������D&yH��>MHNjU���U�h����=c��	���ӳڍ&Q�d�8�5h�/�F��h�r��O7���wx	m� A�>��<�3V�՚1���w�F���ք����`AM�Q@�r�Hf�KR��5`���ڎ��ǡ���ݢ*z���ҙ ��󐡟2�o.<�jL����1�w䝙�C�75Z.<����AZ�'��kN���0G�Z��u�n�&�	/���^��-�T�FJ�^�Q��y�E�>sTt}�����oMt��u�c��?,��[�Ra-ʥh@bd�7��%z84=�ϒ�X��w2��<ۣ�eXSF�	�n#~������·0mQ;���r�`��.�ѩ�)��aq�ihn�(�b��Z*�z����3�9 �O�^��2;\�p�q� ����ŏj(���ڋ���O�Q��l�isX��#��`;5M����ݾW�Y{h|D	�%�D�
R�!�%̵T���Y
�.'
�R#%��1�b�U:A��2�!�gI���$�0�UE-�2ޘ:��bdA����{5 �s��.P1߷8a0{��j��6�޼j9���vU�.� �5B�+90�I�gQ�#��v��/�Z#$�'�\�@��iROF�hh��{5��J���,�L�D
]��0i�]��F�r�z~�]��W1n���Xe�{��Ċ���xiz�r�V����PNR^a,W6l2�N�/y!Y	'4u�ȟ(�`ʆ���}k�[z1�N�W����-O BP�]����@&U����jڷ�2j� �t'���y9�GJ��B�J�	*+�{:��c�����=FX�VD��;J	�<���@���	��#/0�r���KA��,z�<3�Dj]w�}������;���&^������T�@!_;��&�J���5\B\�4�A´�ٯ��P����K�u�X)���;o���5�����S|~;����z��-�5��-C͞5z7�.BC\��	��~Tl���,C~2)���{�eYmR���O�8����b��Ϧ�;�
\�}_�HgɎ�,Tvہ��([�RX�7a����W-jVI��\�����!y%��76Ǵ�zW:g�P)rӜh� ;��v,�@&']*���Q	oK,�z/n�p�GS�H��:H�i���O�b&��6�Χ�{��4X�垼�3�9�)L����}���D(�[�aY�W�糍ƀ�2/������n :EgW�|g���H��'˪�k�L�ǟF�x=��ڶJN�`��]�Y=t�PpGuEY�P}�P�!��7w�yC6+���� Y<C���$��&�����G@<�7R�
�K�� X,�Z�ԝ�lÝ���A� �4km��њ��_��k���x�����o��Δ�+�Oo��@�B�����Y��_�`KlvIJ�����\
�AB�U:#�Ky������q78���6�v�j|V�-�C���z�<���,��w��E �DG9Gx���`y�(�A���K5g��e�K��l.��p���f�x�^t�;�۠?��uO�.��:��G��_%�.B���1^q�Hǜ�p�Ӝ�̀ͣ�&+C�80�W�x����ݭ���AZ����w�k�+�^)%X3a�T3q���?�4�b�A�p4CB1G���=��x��Q��q ���`�g�e�!�v!1k�U{1D?��Q|+�g���r�""T�m��L���%S[��E�7u�Î�aI�]@�P�I��/,O�KW��q)ݳ�:ʝKKO��כ��ik�;��j����fk9�w���'��^.X.�>.	XxاI�E],�ͷ4v�U%p/�A���ߋ�t����*J�>�GZ�jK~i3	��M*&�.�q�Hf ��O��
����{��m�o�"����R�1�	1�s\?�>�G�k?�C���R���۞��	#{��ĐI�����Ἲƶ���~K�%�1���j	�	u���MA�U����g�ǏQRȎ"U������OxP�MtM�SP��l�hY0�s�"vƮV��l'��>DJh��]�8%��xA~dሀg�w�B��kx�e�C3NÎ�?'�Y���CZ�#�½�c��`�q��#�KӉ;��T8����2!B�6��a�X��͙�E )����:hYX\�k*T��HŞ���VM���Bjy��eiȴ_E"��ǝ�R����~eN���5�T~�T�����;�^�,�~Q�NPd�t���_�^�Kc�\L'S��S�'������,"��kh'[�ϑ��E:��{�tP�ϔZ����V�SH�ЈXD��N����Z6�Z)��iul?l�f1A��3�2��U�I�1X�*�wi�h��-P��]��F��!�3��I�-_P�d�ԡUƟ;i���.� � ��~�7L�7��\��u����P��*+X��NWH��^�m��O�#� �|q�i�w5���0*x��9_�FT�Q��LR��t�ۅ"���`Y�y@��5��V�`���;P�hM��Ϟ�L�2:Z�b�b���*�&�:NH�Y�ɽ�Z�K�q�G�4)��z�"4p��|�s>m�+!�g}O��u=�v���2�� S� ��>%=(w��S�e��@��6@y
��x�ܛ ˚^ ��r�K�Xڙ�H?��hz�L7�f����"�NA�]f����\\�q�/�X�t�i��ry�:�uz�PՀSql�{�p�ui+,�S-$�o�; 8�j�;�V��}!��͡�#Ӑ��.^�&����]x�/�үp���&F���h�8f��J�,��S�zh4LM� ��L���f���p��@1�_k��K� �!c�,��"�o:u�k�`����hql��:*i(ۼ3�F,���m�R�霸��\A0XF���[\��!;�j���(�&�#K'?��(O�~���,�C���W��3r><�OZ�>\��F��}J\	�{�>��������x\�v�%C8DY���mh��0s:��k�*Q�6����5Æ�%m����'�&�i��c�"y��@S���Y��P���@������
�d���7y���3�X��)�iPD��o�I:�����U�t�����#��=��)�;�'�d��V l�?@�$�E>#�J�����C�qźv3�P�ȱv��z�8���	1,���mI E���xd%?����)#�WTA�91�M�/��~� ���9�p�Uڔ��3N�?C���%�ﺵnDR7P�"V[r��\L՞�����U�+���I԰�!��4��
�����F���+����1⦔	��>W�>�O�4 ��d%>��C��u���a�������R5�=��0tŲ�y��ı���KuIa��-�劊m�\[eE�\Wp�(PdV#e��B}I�iVN�"�x9גT�����%��l'��q���>5�h|!i��$����W����M�&�ő$~�D"���WX*�*^�	FAVk��l��mDs��\�����@�� �k@�u�V󚾜���pvX�릜���* #����n�s���c��t�v�9�����P?`����tC�t���6_4o]VD�*���;{Y�`z)��w0 YՁ.��B��v�-	N�j�f�?��n���o��0�����|�, 2}wW�<:'��+ȁj%�r$�.��a�����	�_g}��&���gjԩء<�7Ò4?�ki�R��2E�����|0fU�٭���~�3���+15S�����*�V�k�~ Јf_�b��	c�E��@�' ��A:�Mm��<X���ߣ�4*�L��|&�1^�7ɗ|���0��#�o'�I���_a��`�80B{^��������U�ɹ1 �������H�γ�^�_T�֫%����DuL'��h^���+��9�<d���?��*^Q�i��?���#Ѹf϶X;�C�����L�RtW-�-��uի�j���QR)�լga���<��p��|J��X�	���j�d����_G}b�g��۠'�Khx�L ~c� (u�w�6�O��:�����&NT�C������gX/�����c�.|��e�K��Vz��H*ؠ�6�G�y�BOX��d,����s�������W0ؗ9>Ә]YI��sb��O��Ќ^�����h�b�cU�E�E���8���鐈��Z���Ѡ;C
g�R�&S_?Hie#_j$䏀�)mx$��zTA<跕�m�AU��k�6�S��QH�q�̇/�=�]��=9�vp�q�A#��ޝi���d(mؔ��z#	�i�p!��m�!n���M���">I���Fl�/����\�]o��U!Us�ߨ�{i]Z �ٗ�MgJ&=���D�i��Y�"��{za!�͊0�5��c�i�Fo�����h8pz��.�]�[��=���>͖��J�����/sΨ��h{}X���3��� C�S-��EP�7E���zY��~�H?��Ė���
������r����.�Eu�@Z�A��^����BiYw�8��(nz����<+�q8Ք��ݥ�9��J����l�޷Yղp5��x�<�@�Z�b�p./�3����wE/Q�77���-����͚#�� ��/���}x#��ډ�K���$��`P,�`�Q����t���U�9�x�`�+�/�v��ښ�t?_����"��X�7iu1�䵅�-6Sy���=|�>��0ݴ;�X�^��p�jػʫ��Uҿ��3�VdF���+�w��;П�l����P�����eH�	O�e�za��@+��r�ȂSF�Yܓ��n(�j�) �*��//�M�p;�N��?�֧�]$�:Z�I	��	.S�R�f���c���(AezU�*�PHnJ��߈�u�ǿc �A��6�m�$1d*�-��O!dm�i��!�N�K< #���}���o&����a�����LM�(���Q	E��9i�5k@N�#r�u�6��q(Z��T��B
���<&�@;���ϦA��%�[Ye,@�����@�~GX���﮶~��#���� vU��0p���kyg@�twk`�Y��0�pr*gzq�3��`o�q| Z�A7m�6_��G�)2�ֱ��2D��i-rs#:0IX@���s����,!0q���-�aa-ι!�;/@��~�=z��-��E��< zmLx!�4H����.G��n��p9�O�����]�IF��$B�I�8s�f�u/�v�Qa�H��OС���h<����XT�������'M9,�X��	�G /�^&���{I�R��� �e��X�u��l�\Z��,��9{{�(����ݤ�f��_`��U%T
D����~��!�z�܄���f�����[M�7�.~�"����=��'� �h�R�AVnM����׾�$*`�����!2�@��8���U$����"�����ń��~I.���NMf���=�������)n�v@�jN|��������PiN�Hg��	���U���dX��-���oN�Y�*�6�fUw*��c�A�.��3SP�uߡ�%6��, ��V�Ҁ疍���
������h+�R��fgc�S�  s��L*	̂]%E�B�Y(�~H�?<M�_3�vE���2>t~;�Bz�aAY��Y~�F��]8U���E��(x*�Xaj:���A�C��q�]���T$-��v���Gk���_l���#\�2�]Ҕ�(�Y'D��p\s����D��"������aˢ"�}K�ɳ�fx�V��H��f���"n u���IL9߃~-+RNc����O�_��c���Kr!��<f. j��9�(���n��IZ�:����q#��C݃pK���"�S@e�w������S�&ۏ��Q��v�Y=�j,�D�7�Ln�s߷�<,<ߢ����@���qL(���]�-�w�a����?�/���@'��ؽR#'ª�-4���0,K$Y�;��܀��SbV�*V+T =1��X��_O��%�0�y�Y$z�w_~^]}�`��"���Wn��� =��\�f�|�a��&09���l,E���{���I��)�In�.i�y^A�0)9��������]>5��Y��{�����	���$n�|��LSƜ�J�\�9�"�T>"ͤ-��K�	B9�'*����h�ʣQ�w�v�(�����]>&g�KIO�%���鄆�������I$�ܺ$Y�6�̀@@���@C8��v���)��$SPW�2[��OHoɈ�3Xlڬ���҉�>�"���^i�Q9�c�o�b�f�傶5�&O��\�d�9x�>�X��,e��&:��.�h�����Dx�`X\�t �������M���̀�
�Ƈ�q�AF�ZSYApz|���	��g�1�c�m9Y�]�R��D�@{�[���������"��*��>�޸��@)��|�S���?��+k�G70�9�E�h����og��v�T�����6��sP����!�%G����֟�R���?�R�uW�'i��!��w�eM�!
������w�c��N0̈�5e�\� 8Ǉ��c����n'*K�/�l��}.ɥ���|[[��D1��ъ���7r�uN���2�����4�.׸�L-5��t!�&��B.��w�JI%���'����c��&��ã��>�L2�p�-b�L�lzu7��cO7��0_�M�%�T�Ko���������DR�:>ח:��a�ۈ(����u`�x�41/Y��^��'Pm�-�6,�U��NЁ�̾��R3�~�i�?��j���$g'��`K41�[���䖮r˪�xܟ��|};��oe�W�tHp�`�z�W���FXq�^�B 5�h����o�Za���kK5<�v7�RYy��R����c�'b}�y@4y�[V���\:Y&�8Y�3})��H���g@��J���Z;��;zW�U	�W���M���7�e���}t?��C��c�E�W�+��9��=��d��mc��T�}�p�ֿ��hɩ>pg�kN�7��I��Ǐ���XTDz�q���ٶko��a��M���P����ʯ��u}��q|S�un���go'�|�0�
76=Z�Sk8�����x��dՍpV�M��t$�fNRx����S`���Y�)�E [_�����ߖ>E�Si:tj��.�"�1��6���X�l�_{X�^x[�����Z2\L�X(����&�$z�F:ipVS������Rɔ���i�Ά�S�w L�h�~&�&D�_�4���-���9�8�j+��rbn�������@⤀c���S�s�V~�EծFT#߄18�K��������x1⠒v�.2 B�y����۫� >FL�."��73���t�}n�b��Ndk<K�J����n�\]n�=�cI*��x,ˆ���Y����j�����?� �t�f��~ء�* ��"d�+q�Z�0c�s�+��11���Ϝ\Zg��� ��¶α�*�&XJE���t��h{��GV?/��-��g�@�Sr<��M��nT-���<C彔6n鞰��0�"/�j������X�s�Lwg|=�����R� �b�MR:�q��19�QT߼�7fP¾�jC�l�V��p�z���u������\��?g�=����@���Fcj�Y2
�
GL�\�|��\ͺe��K��w��q�����`SDmV�sDH(S ��1���[[�Կ��薈�A��ԃ���s�E>ձw�p�,���ە��K&>�D��"`j���Ӓ3�8��/G��$/���C��7د���<@J�7oB�/�˹��hN���ޗ��>�Pl�G*y&?Kx�������	:��C 
��)�Y[&y�� ���t��S�j>�����כW ڝډ��W�{L� ��.�֫�P7/�qۦURj��$��Dq�H����.��������􀒚��}#6�8ˮ+2ڰã�Ic��ŭZ�"��}���������'s���>D-�G��3��״���Eņ��?�����Z�=C�6H��������8Rb(��K'�2	6�j n:�1Q�<Й�l�E����U��0��_�I�n|����;�0ZN���5<��X��u��Z���iKF� *T3V�ނ	>�p�αX���Rm�	y@Ke��%n����N�z�Qb*��!��wjDUG�y�_jo]�/�(4=I,N�?(�sū0�-ek,8���&�'`�L����^h(,�69	�Z���eΩ�xT+K�_ܬ@�~5y	b�n��������k�W��%�v����^�>o��Ѐ8w{�N�(��q��)1�׀ƕ��^$7��{����"�^���ӆd��L��WI��ුB��b>h��
Ή��H9�{���W��E�Yun�����F��<�]1mz%��$(��o�O�.vJ�j���h���ZS\����7���=Y��1�@����\�:�����,]�c,Y�����.�'��0��h��?}�@ڟ��ݍ���\o�tۧL%(��,s n�ƫey���O2�����th����rT���!4,-�glP�Yc"���"x.���}�	TeσG8�,0���[�ffYԾ�P�8+���p,�o��*�=ѧ��O�+��^��yx%�)?0�R�;?C���^���t��Nj]%a�����9I�?5�-%u=f��� o�$�f7����l}�q�`�.1s�K"��{;���=�Em�%Hv7}_:�O�k�3�Wzr�S���AE�W=P��ۅ�S ��\��K���R����h}kX���G�5��n�1�����O��7�˽ ��Y&bo���GG�Ʒ���R�o��o懨�i�	��x�M�p�����莎٘�w����%�-���4��D����bk�'lZ�)�IxF��!��~�;|���i�}A|7�I�1��5o�>M���|B�Yا�xȀD�K�������ڻ�d����Zv4n�>{r��<
,�;6���\��G��N�(d�����y,8�ܡ,x@Yݑ��~X�^iZMGtk˿�hZ����Td�MX�#C'����k�t�zoF
���;Ţ�{@+�(\����Ǜ��_^�y1�S&/�-�Q�s�PsU�c�m�����"܅ u�����ւ�7Yi	�'��bt@����.|2d�~�+����D�ܥ9�+��~�r�ꗊ�����큙)I�5�G�Eоh�a�!F5.�d�B/<�G-�U͖�UVy`�/�Z8�dF;%������e��.O�<�_c�v��A�W���ʔź����T��/:��4#cr:XH(�!=(�͙�P�iJ��`ը���m��<��݀���gj������ﬆs����0��j���[��[_���X-4Մ�ؑ{�8"��rYo.��wg�8��8���Љ�b��WU���?	U����"�y3��g��g`�1��/z�ȭ۸����M���v�X��2y�a�(pU����_�,���u>�Ϋ�3Z)Ic���������&�"�||�_Y���<�I�F+��-���%z���&o�Tߑ�ݩ�a}w�c�v̇~Bgl+~�=c�O���j�NL��~�V���+30F^;�Q2�.lZ�!���|��v[υ&�#z+
��z'~=;�}����ӄ~p��&Rךe`g�keoJ
�[�<�m�����NWJW�4Φ;�A�9ŵu+��E`X��TdKP8����$������:�|#�,
k�9�gp���,���p�q�M�}����6]{��b��|9A c��o��r���.��=Խg����4PS�륲�^�|IfMmhm����t��y�t�gg Lj֗​���k�^P����xO$&Nt��w6�>��G6rJ��� �PP�EAݼ3�� Ӄ'�d��I������Sb�u�0,��� �_
��Q��$[#݄�Ĵy~���&투�oS����.D2�e �y����l�)�{e�,@'�a5A�@�s:��Iy�h�!zDI���@d;w��$�
��֒��� ����F���䰍G�5��UE?�櫹'Dڐ������"�������[�>��X~K�ϵ�ڹ�iuq̡�[�as;��Z�<���;�o�������{m���Sߕ-���B��Wk�]�dQ����?��+�opB���,޲v�>�]����v5�-b����_8�QNN��1��kH�:���eɉϬ;B����8㰸������Ztu؅�M����t��Z��zQ�
��m��C�Uפ��F��K�g+�G'�&bW��4��`��w���n�W08�v��E���n��P�����i�����WglLR"���q�@��~%ݏ�|Я��%�,J!�������bӴ�[�Ѻu�YԸ�/���������ɬ��@ǖ��"���t1YʟL*��{�^~>�J�h��Q��D'ҝ��Z��,[�a�G�3�dkV�I�/��^���I������\�#E�SH��2����u����L��w6r�HL�^N�����"(�FaEOd��Ϫ��������\�@��`�����:��1�6,%�Xǋq��K�����Gn��,A1�iב'$dm~�I��K�SD�ڶ_��2�������_�a rw���~E� k��y��w��"SK8��p�����������ȜX���<�����-<}ah2io��L�i��x�'�x�&��y�.�_D+�M YK�;V�I������y��k�i(�,G�^=R���G0𭏊j�
�'!�[5���Z��'?���ۇO����hʀGХu��u_f@m��.���*�6�D
����I-�7˛��+Ȧ*�5K Dw����-P�:Tď�d \��$U��9��'H7W�/V=��
���R5|=D|�1���۴F�v~�$̖�
qoW�S|7P���d���6O�E�3��n[��gq��3��);*��{�c��w�i�]��?lb��+���<D��_�_��"��U2�>�Sc
\(j��&�_M��=�ӜN�<�{�-�Y�����b52���*�zZ�<���������@C�"�;X�</p�Ԥ�Z������o_#�"E/Z��G ��@�Ac�4P2	n�7��4��n��;��q��^���}��[�J�����7h�ᗙ����>����.�N�5�"UQ�k�R�U�q�i�\��y��Y�6�l��<�T䟓���?J�q�ΐ����1UoS>��	�@NN+(��p�,�������Y�2�W��	�.P�E���P}����SA�g ���W�L�.��2Y#{�#|N���w���
,���9�S���/�ޢf�ߍu���>�s�碉��"�\Lm��Э:�H�mC�w]WT8��-6]J6[�w�v ��ٶ1��'k�y쳻��U=��ňu�6M�hx��"Gy�N���Z�r*%�^NZ���Ϟ���׌�۪��;�Z7�a ���Ϟm7���o��N�9�n��֎�>E옹�����������Ig(�M�2j��)�*u�����a������K�q�ϻEL~"�/�]��ݦm����w#fu��n`�)ʬ����Ǆ�[/�e�^�����R�e ;��v
<�(���j\�^�G]L5|�4�qy��3�M�ڨ9IN�ddZ�;sgd�m�0���3�������f)��-%�uì�m1.0���J�}L?= kGN��F���̒¸E���:G���m�Ez�0��·�z�j��.����bLx��\;�ȺbT�Ɉ�t���(�C%9^8YR����b� �����k[��L�0�������tCcU���ݤ'.LTG6x�0�c:���w�@��!��ćBz�u�S˸o�&:�AO\s����1	c""�EH��厹�uI>�����o)�����_ti&�"^s*�;@%0�L3Q �M&�v�a~�*D��|������D�i�*���R�em)�B��w�z��:��DcVC�#�7"P���� H��׎��+��v܃*Z�ý��F5%D"��l��b}�;i�9
r`	`������~$hv*���;�醶fE�-��M��P�Y�@�J��7=קv ���v&p�̡7D3R��{<�����雪�����OOe&�bL[R�?����^6��]de�x������4���r��O��#B�s>�ɵo�G�z�xǵz�4�	\��J����)��Y*���3�w'�p�}I�����4���<� �c��
<����>Li����8����[�}6��5�cxa$�>�D��3Ƹ��oJ\a�ٿEi3#{���i�W�@Ð��?ڝ�!����w�S�<(�$��s&[W��U���p�o��1����N�]%�A�W�]�λ�S*���Z��4�0-��%�Î�@'��7�j$e�Aq(X���FN���@@��=���$��Z���l��Ǟ����r�oE\�I$��-D�8&�4%]�Ѥh��	����ae'1�N� �,qh��k��ES�0%IOtG�X]������Cl�5���$K�KZ�Ĉ�C���ط�+��U�궬����EW���8W6F$~ܔ�49y>rV�/��s0Z�<.xKe�%����Z'$(�T�Z�Y��D9\��z!�!D�:]���`��|��\�L�>�k���b�'��Z҉:3�V�փ}�E���7���g�P�.xĳ5��(A�B���''�㹱��l�r=!֣#lʡ��1^������|F��
Lu�c�E"���Z���|Q�Nw���
���h���v��gbD6������'�r�Y
Tyy\g=n�U/���]	2߶��ĝ�Ǟ���4�~�[�p!�7�1F�m\!yZx�9���n�u�>�f��;� ��UH�s];U�n�J�t4q=d��H��Vɫ�7.�I.���h�p�����Kteε5`{j�7���y���q���n����^�7�fU�GᜏE�Y�"V'p�;%�g��k`N 承ų8}�&A��\ ��&+���8ʒ��e�Ov�6�(�LNf���^w��c��h��b�2���-��j6A���:щ�����d�:y���3|�i�R�Ѣ]�o���k-B�G���-SS��Q�;��PI���&O�vʐ��5
�Z��8i�;�L�	��2���p�NVz�ȫ=�rCH�w�{x���Į5Wn��F�����@b���Y,�,�-"��D��G� �XR�IZk���K�]���Rg�Rz¬X�S�}���=���5��P�M��La�uck�(~)(�c;)k&ׯ�ds��(��q�'�g|����O,���L��������I4Qy���S�Y��3I?8w���Nq��߃��n HO�^́�^7;�q"���+�\�t�8���I�aw�綟�q�l��'��C��7���/ۭ]��Qc���y�；U��p�J��Цg�۱��-zT�/�"BQϾ��h��qE�t���;�I�cAI��b����[����BG��+�s���^�c>#���
�W����ږ��, P%��
��7")T��{&d73d�m�¼dm����;7�zzu�^�qh�}�hف�U"4�DLq�Q[���9���>������?Y�SPܟCN�+��c�eD`Gd�$�|hL�偞�ܤ%��\��1^$q��"T���ĝ�J�Z����y�JW�:l/��\-���*��r(��'��O� L.�i�_)�f *�6�+�K��4t*���Hi��fF�ȹ!c�������2g���`�|��Z]�>˧��eӒ�ϰ����;Z����O�Z�{]�iS�r��Jam�����V�w�@u�ƹF7�&�Ǚ�h��z�QC�| *�*�A2]<�'c;?���g��HS����4c450�|-��V�m(˶�o$���f�D`�^�����?܌?��lv#Α��^ g�Q���u�����e������8����T���������=�AG�*�n�p��04|s6��N��a�a2�:t���W��n�>t��j���B�o����?�J����W��n ���%f�W�� �x�*�c�����)�m<���\��z�Z�� ��SHL��6���S6u�IZF>��\��]������&�5�@�ђW��$��&��s1%���n)&�OK�G�$'W��%H�?�T,lYMg|Y}�qS�&�>�k��ycbȧ�K´����溙ҳ�~��՛��U�0a]�ܰ���	�|k�7s�*Ȇ�"q�"���A�̙��9���\ySn�O�.joj-F$؅˜����#D5#"��=5ߓ��[��
�<5F��H��b;v;	�w�q��D�tr���O�����[��\�*��L�����WDHp<�޾�[ 3�w��W�W�~�x��),��:�)�^�J�;���cȭ9A��r�#�tPy<�ya���������e(	ƨ�K���2�E�yr����m�9�O|�18���P�o�����?}L�ܡ�z��h���q�|N{�2&�()����]9W�k.��b)�-S��(��~v�zd�Q9b	���ǖ�b�-;Gг�s�8�"�,,*Z��o�	���y��P�`���Z���n��T��� z�����H_�͖{�N���؋;����[ ����vA.0�a���K�8�,�rï]����N���`1�v����Ц&_j`r�����ȅ�����)�i�����5�b
7�u(��^�j�Ւ#S��}�#�V4�N��N�0��j?��)ҋ�hb�*�~�M՜䦸'��y�����`[(����V�?��+���?1�݉b�xB�Q	�ʴ��$�OĶ�w2��!��h�>b���	���@����y���#��'��S�Hm��U�%F���u�E��;ٵG27:U�b�Zi�z,�����f�򩼀��l��	l*Χ���b�LI��ټk�!�xвh���!{�;�_����ߥX��J ��0E��y�(az�؇�K�f��X��Fܹ# W�SiXŐ��2�Z���ӣ���OI�;)�%5���9iR�)J�G}�]���%$���skH_[��5w؟��oN�X��-t7�j0��ak��"�ت��$@!Y����l��\����q��}m�O�'m�)G^��gb4�z,�dL��!�V���� 0�g�	�3�}qe'�ޥb��/����)�Ji�6�Թ
j�=xܣ7T�\����h�Rƍ1���L0ݏ�3�u٣˪ô8/�s��av��$�o�����w�g��h�q5*�-t���x��p�$�l��K��}�Û���d��]JO�*���F�3�C9%�n�q Q�諕)Q1GLo<،��Y�V
��.�D�g)ߊy�@R�_,�۫*e�"?li������59��sӹ�"��MuƖy�r����r�o#�j�D;,�?����*��l�9��lK�%6ɀu���';-@��C�_�cy�^R��������S?�\7��}t��Œ���5�r��Kg�-
1ܕ-G �}\�Qk��B�f�J�S��&�/Ep���T����
C�$ΊȪ�k���U�	��s�����u#����*݇��Ts��8����ܿ�R �S�\Y��СV�=��S~r8� ��*s��D��-�ˇ�2�̟���qF��o����I�C}�*��O�>��z��	�Y�bF��;�0<E��Կ�A��i��Z�ˉ��j��_�]XA?��4c/�yX�/��{'�S0W�65W{�F"{��zbu�b�G�F��XVQE܏8T�h��]�i����?�>p�l3�fq��E{8�6�������>nV�U���k�S����:�^}Χ��xS�b��Vԡz,y���ZԌ��&śD�;�I.׹�auv#7l�.�k�UЏ���إϗfQ�j�!�6Е����_�P:
Sx��]Ξ��Nzυ��(O�_tJ^ڏ5ڡ$:iGA��諜B%�[�r����mf�[�4��h�%2e�=��f<+����k���O����G��0�e��Jh�I�ӂwW����ѣ�Sz�5!���u<��T��v �jX8g��2[�����'ؕA�S�,�5���RfO�-��\>�7+����g{e��)_�#�5#w��<�����e'�B��ri�����h
d%�hqwF���`�ཛ�v��nT�!���	�����K�mQ�����d�G��!��][�s7��c��V)�ߥ(���S<��Җ��v�&�w������ǳt��������d�7hP�w�c5`4�� e$sPo "��{IE�A��W�d��l'��9ǵ�=-3�������6��jІ��T�Ω���8!j=�Y���N��͋	�IVW^C�H���m����������~�������/t�D���7�ru@�qA��d�V)Ŋ����h��T�����eC	v�Z�����F/�Ef��}��6����ߖBQ�w�L7C�xd=8�`��|%�Խ'�"�u�f�hm���$�Չvc�H����fz�!�ls�	��o���X����x:�)2FD����z��Tu�$�7׮�kؕFެ�9h^7�~�,%��q�`&N�ad�`H,m�����۶�m#}�,�l/y��`�O�i�yy3a��%��GN��lx�/+�=��DOIF;�͏{7�f�N�
hx4�bb�S%-�x��G�V�`S3]��a�;37���/M{!�D?`�BҙKQ5�����.ΰk9��t!BU-�]��*�(�,�VTs��.�A��Z��K�.�(�,�����O#jɨ�L�7c��BAV�τ,��N�{,�5�Ȯ��{rT�H1ܽ�}Q'����-��@�`�0b�B�����䐹�G�ի��#�-��4YvK��s�@����J&>��jʆ��Q���a�ٜv�sIoT��>�Ih�eI/KT�^Iq�H����K	��@���[�$3�9S��2	�9}�1Ҷ����)���]���/y��{�kX��ȟ�o��Z]��{�7�>���6�j	��.����ׇj71Fp�R��_I:���c�yC$�&�@�z6zwg��a�j�"����-Z�Et��:"ll>,ƣA	�?�!f��b=�x+�;*8Q�vw,�8U�J���	)���!+�6��ߒg�;��`i��ۖZ��\�7���v�C�H��ĕ[�g�����HJ�^�X���&�Y���D2S_KQ����l�n��U!�.D�`�$� :�QW��������K�3�d2z�S?T�*m�S��ٱv�p�XO���"*�=��V�A����^�9À���� H���d�2mi~E��6C��#��X��L������,D��\�K%��z�?������̞�$p�& ��þ��
�
�E�2T��&���9O7)�۬m�d���*_N���+�� .[$�1l�V��:�~�lȑ-tM��ڇ`�4��	����׻�����c]h�h�㏕�-��$$0S޻<����j�*��ېA�/�m׈8:f>���Ê���)�����;����W�\�-��(����(ú��gV��(��n������.�o�uq�x��/grpǯW��ͱ'�ʹHkŌ��5͎�b|���,`�|��:����Iv�N0���eRS��U�꥞/�?�p�F�U��߱S�����n�mMJa&��Ry?D���w��tLPae���P�����t![i=�PZq�: �g���Ԓ��ާ&�����u��w�Ħ�ݾS\�{rH>�Ș26o��h>�"��_Ł��y�9`a��j
���-K��RY��>�G���MD�1'��4�E��N�XЫ2.��r�6�.'`���X9�%�pY�lp�#3c�ۋ�C{��f�������ϵ>_��:�O�3ҭ����~�j)�W�Cľ$j�渥v9�����6c���z��<�E�� �@�)5��]�ae��5HX�ͮ3Y��4��4����K^�ߌ,�E�9X�/�UD揇��<jA����"֯��2o�%������]���g �q�/�{�8j�7	��V�9Y�4�u� Goi�( 
u��Z��
�O�G�ٟ._�E_&�{�?�)1�Vzix�h�]hIn�BY�DR�7��Y"�`a�}ά���!�IӀ� �8߾c�Δ�:@(�,��Zo�ZX��F������ƱG��3����L���	��_�k����i���O�p(F�Q�v�����DTU>�Fr�x��лuD�	^TQ#�h��>!�^�&ʁ5��}%u*���l�8��а�0���q�F&��lS�J�j�ևc���x� � �sZ���a�ϊT,���[�y[��no I/YɆiTX��>%8�k��Y��qæo�j��b'n�e�\�[3\�C�rY��|0N�B;��!:��R��%`q�믳�P�w�VA;����XjT�0v�$s *�ǋ�H��~ʪ���_1��L2a2�����}�b���tK���}�젽u*H��l�>q�]c~{m�A��7l�J�@R^��Es�&�)Z[��i���i�o��G+���G�&.om��/� ���m����g�>˔�(a��X]�2���C;]�EaTK�5����8������]�6�����
X%��|�u)-��F�-�����H��XQ�A1���{&�B|B�#��	�Q��o���8������X��渜�C�iڿU�Y������Z5�B�YC�����Ո��?��O
�.CD�UlR7�BGS���g�O�(&f݁�z���������N-T�L<*���8��2 ���KրO�.��vA`|D���߮*?h^7>U������e�i���|�+#���Y���a�J�1�?<��� ���]���C�L���v�|�0�+�!֏1M���	�����#XK�6�G=�����C	�RHc�eO����)5���]vN2G�T�A�����0a�g{���Vl�X����?�V[����#�T]��]��^u漽
���pcW`:�G0��䭵�:n*�X�\xF��f�^J�l�R�w�H&���s�N�>��aj�NF呋��`��0 ȅ�Rz�!�>��K�8�F��-�J���h������K ]�� "�c��w%�sgї%��GI��&1��K�v(����x��k[�,������ �rO�䱸7@�*�Sqqe����^����"_���mm���w�	:�X�H�����JK��෨|���Ȁ�T���[�ʠ����m���+ue-���#�x�bM���l���bno�]��A����d�!��{��?H�Z��9%�^��x�~���u�`Q���.;�^ש��?N���������a�\ޓeG7�U��/�����}#����@����T�ܛݵ��	pէ�j�������t���ߓHU3��Q�h�aqecߧ�UF�-���KAh6��Ü���VBO�渡��0J�}b��.]���kߺ���~9��Ly#�T��=�P$3=�b����|RE�wC�/84�?ç<���K`ܚ��d��Am�{�@β�t����q��fDlHU����|�њ0���V;�W��jiO�tzA��1�I�X.�@�%��N�!\b��a��x��fm��)i��L�d�e���ʞ�4جC�+�<��'#I�0ͤ�7�|A%�M�ǽot[���C�b�W9�^�[�k�v��P��N������~ɍ�c�Y�I���ˢ�����R3d	Xr��xb�nb�ԃ��J��d
�*��]|R;:{|�kTj� _�� P�7�B��!zg%�G�&δ�`�_����[�d_��fڌ��;��<�җ�zR�n�0v����; ��3�pU��AjD2J�>.����=C����ܟ�����Q�:Z��.]O�R�	�?)�fw��5���j��֙i��x�|<�B�������/P���f�nv���S�\���D<,�{K%yқ����F�v
}���^��-(�b�|��'��y
%��I�Q�oT��(w��Դ�v��G��a�j9��r�v����"�e���(��$H������%��OفYG���S���*��,x��ﱌ��F]���Y��t��+��{��+��rN���tX�xP	[�I
��Y�=3�,+{~�d3���m_���D��3@t�r<��g}�{ 6דU���b=Bʅe#K�?'�c;�T��k��KC���yX���{Zr	\}`���Υ�������� [l�h�܃@@sf��H��Y4�H�`nԏ�zq�<Fl]��;z�ML�C�h�gT:�P& G�W�����Z��Z�����؊�X Xzn^���N��	r�I>#殮s���O&ۄ�R H�Q�8���N���IX�3Ҽ�W)��N1t�"�If�&`4��|�B6v�|Ć��ˢX}�������hjw5����E�b�wx.�?`e"������d���vx%��r��u�Yӑ���f]퐹wraA�Ŧs�q̑[�m%�o��V�0��u�ь�h�@X�aj����P�1��Уqdq���U�t�&�>9��J,�d��x��/{A|0�R��A�6h��嚤a��hwt��m�K�������wdN�HN�ǆ���+.���|�mG@�m\�U�̤���q"?Q��B	d��4�I��N�\��e91*���1o/$���L:1�i� ��k��Yo��5�~�ed�׵s'���(�U��n�G�wΩ��T5�>w9�����!��/т�>�T �e��|��J��q���2����IDd���R�Ԏ��th�p�e)S���6�h:��
�S�������3D: �*5�[�*mh#�������c}�i����L~4�pmN��$V�̤��b�2b����HE?�.��/T��k�Q�#���"̘!�2����A��!l�Ð	�w�{�����*s��0zt����'&�$�;��-1|�ݙ��W�`Uqm����p��qI��&AÛf��i5�V��Sa���U�C�G8p{L���[ {��|@<.r�U���\0^Ӗ�w�q� ���:S梨�?d�Т�Z�x�>�3e��d��Q�y���|ǥ��ܣ~�"@e�	@]e��}�ru=��ep��b�*�6b"�+�E6I�j��m�Q��4�����Y��EC�Pϸ�!����bx=�/~o�rf��w8�a��rG/��a��+�X�ӳ!��=�[;ꏫ�v�Q�BHA���nY\r�lA��:M�29�}֊���a�J��2eռ�64�F}�y�������KVvQ7�;��,A#�AN,쪊�F����S��,�75��=�c�21?���ah��)�E�َqg?Ūp��ٹ��^�Z��t��.��e/Qm���\�+쮰z��:J����d�9���?e��q��j�KKl�Θ�A.�3%ͧ�H8.(�TZ.a�a�d���!v�9���?L*}��V�l�꿽:܏�uA|��Gi�A��g�2�����N��4p����,�"�ӓer�\�u^�� ����)����x�� bA��RZ2�XW�Ꮸ���P��6�-YH?�0^�c���,�PC�l��x2[�Ň� vԮ~�_�ޞ��Σh�S��<+xZ�q*[�u����8K�mihX[�H@v��	b��(������taC�ú�(�����^��ʣ�lŠ~�N̔4?<�[-S"Z|C��] �2���!1�n���*/JJ}�k2
T��Ǔ��Ë?F� El8m�v���-n<���[�eSg�l"�*�"@��L����b�Czr'������A!
,�[�&8���0�1g*)�(��X/:���"��T��;%kz� Q)��fk�."�i[�J�2���4�'b�B�*�vނ�̣�hg|���{�V�� *?�t!����R����t����0���&�S��6��?�Y�M�Ʌ��~HTR�7�0,�1�K�ō������g�Q�bb�lBu>�M�rA����#AOg��u�t.�8�T�6;�c!�tO+
��~$%����e!��3��������=W�:$p��R�Lc�˲`��l\�y�3�}$��I״C��8���!g~h�W���!���MV��N����M+m�AY�eКeS�^��W��X�k��� �Л������������
B�eSZ��Az����L���1��ߥ�ϗ���ͺ hY�czL��lH��K&i�躿'��֕>����Y��w�^O����|x�p� ��}##<qH�����+N]k�[3�(m�+�w�#*>��X\j�� ��j�fg"E�3�2��\�v]c�]|�����Y�L��xCZ<;>�:�>#�ԋ�U������k�c�߭sB��g&D�s{�N@P�`�W2�HD�ݪ���ץt��>���n���l�ژ��j#8��������`w�����]Q�<\+��Qű������ՄH*齉�-�:����l�4 ��/��i��-�ĴzuD=���3���@Ͷ���>�B6�mIl�#0�0��rMIK&��d�82���SE�cz���7���:�)T��K1��fݾ���≵��{lK��v� �լ��Ĺ�W�Hr&�Z�L_�<��dU���u��zfu zA%�\1�����Fg忇�J�]�ҫ[���W|�Ko����l���oE&�d��u��������d��o�ٛ�
�,,E'�q,���9o�=�b������s�N�t��&�3��e��'x���KG�x���.�ߣ���?��'��؄��?f�>z���"����q��h"�_Y�>ɗ��~�66k~��*ɉ�s���6Y�yt6
(������;�+��H�\�%'��^gA�r3u��	�ȟY��:��ʖ
��Ŝg y*X"c��Fk*��)��{�<~`����H�9k~��>8��[������ R�00
���9å�݌A��N�}+lKO�f��(>�6e��)qioz~k��xE�-'5m�U_Um���jHFh7jݦ*}��aMF�IA@�()1kN7ɢ��f��0:�6�P/���v�!E|�D\%9
�p��q��t���K���dw���_LafX���vDx����-x/�1�Ӗ�<'�2�)����5�}�=�Żm"!��cGk��";Dv2�r��)��y�X���"E���t�`���?.b2M�3�0��<�S�G:�l�®�w��wa���7�oO�٩9d�V�	���Y��b�j��@I��5��h��b��6���f��/c띂*4�&!║�g�'A ��S��%�26���qĚ��.��r����ߘ-�@A�s�U��ē���P��A7Ng��r:nG�%��?�iO�n
2���g�f�}�=P��U�w�����kt�l�2<�Nֈ?�����a�~V��� ��f�g����­{�y���I4#/��m�3��B���<���?��]�J���Fm�u�4	�V���  *��`N��w7�s{��6�|)��U�'^�٥��aZ��.���������ە`��g��zWZ\��Q���^e1i�����Pͱ716w|�_�%�s� �3lPD�5� g������p�)��)�����g$F8I��h���C����C;:����HG_&AJ�!��E�� Ձ�R�����3���R�.�y@�-��	����n���t�@<uź�w\��n8�7��s����R���"���"̽zDQ��C.>5�vb�}�~+}�l��_#��V��:�#@{s��QhN�D��yEn��z����AI@�:�1�Q2����$|M��yݏ���4�_������N�?���.�t>Lp�)��s�F��܄��;������ o#Ȝ�����Xgѐ���H~T��K���(�����O^ǺL|$�[��$����#�����U6Uqy�#������q)���f���EW���J4*��
V��^u	.�K_G���~<�"�����mPXQ��g�.*������p0��%��/b��B-#^y�Z^W����[ly�b,�9��F�@� sb�+�t�w`�.��G��<GG�ƍ��m�4�^Ŝs���9�D9L�Lh��DB1� �(�F"�"�ݩm�QpDa4��q_�5������P��!��y(��L�E�e�X��[:�dg�s|�������vLz���D��f�5W;�����8�IGF�����4a���E2�C�$'a�tuX�!^�����I�	�N�Мw)t�?����3������S^�����B	�7'I��{��_��p
-�K�k%�Vp����մ��(Mj�)K!�쭷��"G���Y���k��A�7�V
Y����nHچ���P5�%���!����l���~l���{IH�Ϸ��4M�O�n�Ӏ�W!�����P����߼��H/�T��\��z!q�
�Kq���.�T�PW��l�2�:�W���3Ձő'��<�Z7���P�)��,-B��4+��T�Q`��-���ai�uvl�S���:E^m�(���:$Al}�����_r# -�<�=lB}d��n�冦�d�#7v�x��`2�-b�O�|�_kbH	�����ײ�� D3�NT�	��K=z ���9Ĝ��^-W�R��]ŵ�pgpBBk�?�����<�Q���J�AB#L���^������)-WHn��<���oF��I!���&��{�t�ā>Y�PR�9����_q�&%�ۃ�0����!{�S	�-*�=�г���F.�1O���xGSH��6ejx�R<['�Aٌ�&Y��M�ma �����h(;����ˇ�Ɂ������h���#۹Yœ�4�Z$�2d)��'��K:?�G���=�J��U�~��Hե��W+��( Њ����7�1�t�
��)L���w.�}	"�g�;�4��d�`���TG�1�������@)�G9:����	m��f=�F�%�i�^"N>��mw���_���Z��ב�"EF℩�<'eA5��|C�]Gv��~
��Ժ�`4�G1˘ �F�Fk�i{JF���d�}�b1�	g=�?�*"����6�Ɋ����1^ؗ,1�	/'s����CSC֭K�6tR��'%e��T䬾���;*�$�h�gc���#E\��	�C�P�GəO�7����d�ĩ5G�s��`#�Q8�[7��]�h8��~���=�M�9���Wi�|�fᤘ�y�6�wuvH?t��my�3IUL��K��[h>�G�8eѥ�6\u$_�b�Z�#�A�H��L�F��5�y��cC�� uh����؜�i�7�<����ʙ�Y�R�H����jh;�����H�X�~8�=���nTմ��{D����y�#�r"��0ѫ�1�մ?��