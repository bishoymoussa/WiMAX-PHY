-- (C) 2001-2017 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 17.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
GxjeCqWEKAOs7Z/NMP9fyrfBFoto5jCKquVmU9evAZHxC9iz3ewc+4o7BihYRnHt6c5vbBUri/Pb
udSz9MD2dRnZ1g3jYkL3TILY/X5gmSTllmvz6jyxCw+0RnioMmNNOGVu4mDvcbTknfltwkzL4zJV
JNx1Tq3wnce/aytLmlRVEubBwkhrsqDtd3M7X5KhvMN4CQt4w+hH9NTbZL8n1Xr5/Ap27AhSqhCI
LRYYQF7lhbBamdcvjllqoo80ri9P6of0QLmFU8o1MMo9KXdRMyDIyg11mUsCruoltChgFPQsUmBS
8dyAAuewqiBlICLJFRecTJjin4oaWXuhOrcLKw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 26880)
`protect data_block
vpMPCpvbbtDiqPzq85VYXpYjRRByXxgDuSMN8SqCd0vh1WvCLLDPqL+IPPUqKFZAx6d2PSR6P7RR
Qo5LeZO6+9sCgbz6JutlqDDhfSb6mPvpEIAXoCwBl7wVu1fAvpoFNbti2tu3SKbhGzotpFeFOZiL
M0AwkWlNS11a5PVayMNtgXKEGT++53xwkISkJ0IJwbuz/40mSagNx3MrCnNU0gTLimKaeqBKdxvM
GZBdnF0KRth/dbNzrx5HK4DPs25pkF7A/PqMJG57Rd5TNFd20K6yhfR006qDoF4PCqEkLRQJramp
S8FnBAt1EyWLEbBkywP1xq5wnvRcgAx6yJHBiH1McqEaXatvpW/w+RaRR1F/MjYbsiLs0vzuRnaW
1NjS+quzh0nKxUzeW9qoUE0SaSTlOMgAVv45tqUOL4nGInTzy9yhNGZNAy9qczlJeIzhJr5wUy+A
9EHl0yY8njuGRXfYo8/LZ0ap/xKXu5ALQBQCO6caEWqfIFP4bydCxW06cp7DneHQT3eSHrH7j34T
dGT7ulKdo0LdC3csqtDXudBqHj2U+aWKySbXGheY0O6shYkQoX7YfUzRz8BMYsXBwF4V6IbF9uKq
q8TXDCY0ug5AIE6rbcaGENI/26AYzgvTYo79p39B3O4XXH+/zHUSShHLoOrNTbcjnPbbrW4MeLsF
nMK4fg2LGVyy/tn/N0KthXTikbd9r9pafzk5St2DjqAnwOu3guVWsb3KhYT6Xu1f6UVaZhk0oTgb
puZMAdV9VMGVoNKuEEr3U0sy86/DISjUkiUHyJ5RHPpWpDPbdTCquxXlF1dTdoRhz7rbmd72pPUp
VYtCw1pd/hmrCRpmm0Cnp/ea2Ih/ziRv4xMzMrLBZrywqb98RJciwoBh8dDI6yCbj1iIhAMfmXoU
GeiPp+Boru+M2yWfsuamWnU5/lSMDnQB1yoOr2Esul1nr1iNSB2ql2nEBs0QErURARKSMAa4GxzB
pfnADmAK8rAe+QlnJymw5OPQWQRrMz2yok28VD9uYuzZXHJ9SGRwacVGpW3qtSGBWwDFYjbGoqDr
4A0orZbwQlF3j6QauoeBy9WikbI+qcLmNL8OoUI/YPC9mgiFeEPzzTclMWVMJjnWiudGIYCTxp6d
Fs8vKXIxZPlAiQN8XVjPpUAU8TUhA4ySV9j1I7n++FVOD2uo3MjE6VmYRuir0rgWzHfe8ST75qPu
kKfcObKmN+/8D5shdm1qTEce8lt+xpFFbZocZqNF1tL/OzqFXX/uTyL8oLDH+X8Mt/0RxVo/hchQ
xsQeClKOeNpGG1QYA93QncmU1AaXlXxK4XJZ8aVoMXICgXXNM9U1IVLyEUwHA/z0OTNgH5jSgsDl
n9ACajtxh+xjBKzaqdNhTgrPqaLC4+yViG51jxGS7McS242y/OmBY2h1gUekWuHjv6oKv3Lk1w6E
eC85uQ3QkFb3kFTytwChwcbh8xloinYlFOlMADTPGXoR9dreu7j/u1Y7h+Y2ji2Rtxq5vgat9P46
CoXUsKwm7NCIcN7nHYWpNRSdvE13p5QngFrPEbpLg7ebkw4WAH/8tnIucKZzuVC7NYuegs/XjqAM
NgFCZZXIL6RyyL+PTnezavioG+ac7ywjnuCmT8/f/Q4yuv0Wq9UOztWGddeZqhZneb75zJaRvB99
ZKx4bLjrjSckOwBkHnqwexwD/yj5MGCdPzmXy/L8Ya0glCehQbYheOef0TowUVPTFnumF2tojnP7
Rn4vniwOnMOOXE+CbMQ53119PdiwoO7HrxVsqPAutYptCW+3O2gjHTTsmQfwWIHuj/i24wr+jo3k
xC+Ok791dzD/THqgaYGx8/VESbxQMysK+8UVp+swMvllP7tbJpfjhGEdbgau/qs89Zllbt1N+YT6
wFOmnZuA8fvsbmTV87ufxZX8cZOZXTLMwy1F3q6N+Qh0YsTvWItRF2YET/mDoViHOLwKhwjjTVf1
h1jawFvQFUocLtXMOxeikuArDex5siw1ByOtWqrFpd17XRBiUuke3nsF6Ar94tevGW1RuAg3wnKF
jPSL2ljRVhNNQlpbVnpQzw9+emXvQUmFljNQ2P87z/hI3Z0vya+tKOQMeKh6OSAWslvoqbgReTen
531eceH1OnF21mNtPdT6nqjhO3oVGXIaRZDMOzj1SNK4589V0u56uQaDhZ55RGKtsjs6J86SSINA
hXCTYy5g1BHc5fFKZLvwVyQek/3DMhII3t3GVmevj2XPqDRouWepWLTEYdYV3Lv5Vyjao52v03zv
LQKj5UVA0ORsJ5RZgU7ZwfCU6D7dIy9qUxaIFcWrd4szM31zj2Bc5RFNl3u/dxd2f2Q5flPAaXfm
AETD36fw+mTVzV/VDYTnIvJZ6NMJWSd1NPIN/NnG3oNMZ99hS8wAGkOF8rzPGSqvmI0YjZza8JSp
0kJ0mnnMamQEgNoBVwk+Pa4ysRjFIdmQxtJnF1/ww6kiaY8+OS0XNJp79Om3veJqoP4+wTAg9J8j
Xmv/jXI2I436uS/A1hoKnyBO3ZGz7GJ0D7DUv1SXBODa45UADcchS5PiE/LDANDvmzAI6HcNE1Tt
qlr6c6rhKYzf5VdtcqgdC0maq4dKy45hiBWFYWFnXYEqNnPS9LAlCWwwdQb5R+vbeq58onQvLg4h
aObAJ6pk7e91CYYo/L57tkV8F3O+HuISVrNS0FxsbBPI2MZJDYhOHisDmK9aDVQy4cnK2h7IoLP3
NYfqYPIoUW7McMHtbvrWdBfXrFmbtvFLokuLtDH6GxV+xa+yPJ1jEiMFBpdvazyJn80DZE3f1Ckq
Gm/zBq+LaKEOveO7FCg1hFDnMVaIvnw1gVHqLk4OHOXdmeZj+S2x6RsYHerCrsJcQYWhdfyWQjiR
4RVN8EJzz24GoLC9UlgpK/RDQgU2eixzUJlVUeUm3aue67IFhOWnNqF4001lTvOjPok2hIxgD7Bx
Y4SCJ2FUy/XFwmYbKq7JNUw4IYfzuCHEQhz14IzGQ6z3rqPKCqH1SvLkkoZ5f/WUovA6Bj0panLl
vzxqtOKENWORP6/djFvC2oVKT/xyBL5ekgetaPGC/+tlejUivTiCCT0oUc9/qrbbCRWsUunU42Nl
pBh+cbP4m7CloQ9eJUT+7iu2/Dfl/L4ycxYo51Xa3CHCq+6RVvI+ccZTJArvAfIeTDVn1+sj+LeH
mp1GRVOwTfTt+HJWl2qyp7f+fDTja+L1s9Vl4FsFXWJqT2IHzBDriV7hI7MFhmhIBhJEk8MhAz4h
EiCVqJpoHQp3+1Z15K8tvfqpXFn13P/eDCJoUegGPHAkiukUg6jL7UlNC/DHqUJv9GcvAPP6R2aV
TfzABG4wYcBHrKjYeHS/4YLhUJLO4fqDBmyj4kyhp/BRMcY0IFx5VA5TBSch4oHZfgTcn56odHwZ
VDQ4iM8eXWdnixNaMLYYTkT0UPwljGs2I1NBWLMUhqgjQjcwQLRnoYG6SVthrrLo3cnyhSBWq7KE
O68XGW7XYAW4Kxf0I80OpfFle2hUgGGR5tEcWEJRMP/81FhAtrmzuqeRMDhhX1qLVObSZ8pf7YVk
9q5vXygZ9Uzm72ADJ7aCtvqlCxkxVWcjyNC+ISdydLouF+FFjhBULeXJpMwAPoIn6IfasUNVmZ5k
sTO09RvrJ+vFWy1WYKBR5QX4PbyfwU6XIL2z7is8GRPMlF5IPp6h3nNhqTG7DMGkPgMkTRwzdG7U
5PGtxL8ro5Oy0yuLF+OHJm77ensi1SjJbpfF770vdSwY0qxeliNsFlMe4As2MuCmwrKYTDnvnf2p
XtNpVQ1wltMq3/x1o68qw4UrbOwcjm7pOzHBoJ2nOBHCxNDH4TyYbpuXV0+DjRxHhtJQzWgrnpsq
4g0drK7+seDntg2ZPOfRwvA9DiHM7Tb5rHf2T5n1CZ1ve1zgy17DZY5VIDPjNiaSG55DPUukCmio
vwuow+YoZdqVAal5ErYYJEEVA7ZlsWXYkpKncg8dyL5PhnU4F9ciyeAjf4YWcGDyteqQ1rCICsHX
3rX00+xHysN3h7seCJqZa6BxFNSav7KNs6BmnywUJqbdlmFwFk3JI70fHLLFZwI/ApOpS9MkhrIP
unCBZacrQIytaaYZlvByyksuQ+KNi6W3Tt/mrf56/2nibgQFpPOvZJMVfZ8A6U2lI1zXDSM5Y5NZ
k8aeqAwFggLTzDSPZcHbPyJMybR2TgkPAB9qDtehI+pH22YERc5Ho4L/Ujf1L2PLxkTwKkBDG8PX
8QxoHHZlsNAWXkkCZEvWGoUUt25Wc6urRjnGTQmysEZ/OdW9SYaHUB5sjag9QnQ3NU20FpVv8XhV
yJB9oaPVRPgPNvC5Et2y/CLpAqEu6/vEaLfehvycWo3SKkzd1DF7HKSJzdAQQl9nMHNjpriw1bYl
J4t8K0VTDroIRCx7n72ZXYN4xo3KSQj/CFJuUxeetsuuRlgrMMwhNKOqSehg82l78RQCm3PqqZsp
EFLi2LePt+W279BFN8kpIuIjHWhXsM2oIc79I4Jol8NHVxzPIRhfNRh0e/ylYv4qfq7Ipg3xcfzp
6cmwVbRPufzotkfyIn2SKaT7jajPq7fCqBjG3Mn7pHFUebPkeXkGT/GTB+xbH15jSpFxuzfrQB4U
gBE9ckjzBi2WEi1X4V12zqfWvGwdRpwks/E3y3YzLaEFEtUJLRR98tbhO+q8zCTnAxB63vBqCffd
v+dYAmyl79TdoW1Jf37Uq1CPTCXUL4SEvv4UTltUJzJ4fOFwebVVigALd2mIPwSzOc1Fnl42M9nW
kYxJvyFciCAQ/jkWiJsblYfbYmNci4WrnIURFsOB8LhFkTCrROOQZzY+QAV+Cqt5/6RYK2YP+fR8
jBHt+wifMX3w6kfozZyZJ4fp2yRJ2u8Gf/8TvqmDXA6Or1CWHraAkUGI2K40LElJ1bGST4fzv5nP
t3v0o/81oVPzarGam7gfNkYmm/W4kYmXy20BT+CshWbmyfnca7T6K4e2hCLMqv71PuRjBhUz3tbH
mDKHwg17GThP5MVd/vFiVW2FYBCDY0pS2W83E0jUVnfxUjKz79ST2NEoVc+aEQJCj52L6vaYfqOT
6HW7Rv69aQ6+3kkyUU6n9d7F9UeElbs+XCzX0v/0Wxjytwo0CjFaRSnh2hLODEo54UIkXa3KWAdF
SafPm7XA35Ytv8FBTCVbCi7OYkgZLqsXXV/IWTDKfLOntlSeWgs0+jGDKtbID3dA1NYRqZXBOk6C
1izs8f3wYh9OZ29USgn3IA4F3NoFnIdEAi89PbqINe486d5ZeVc3RazXhn0JVaHb9zF2vjZ4Bda3
MxN3Uc5l0KxRisqLRMgMYCr5I8fbF0CMGceCvRy7zES1sHZa3BxOR6yyy1j7z2WADblxG+sXCR0H
IJ6UkfmrPcuLl4He/h4vfC3M4IcNJpSrYiNSU+T7jBEecAOPynm8W88Md1Am6W4LtQMcKUkVY9rF
gK1kpufMk6jAqFhNvonZYgYO9YPRwitUe7jgfeqV719cvr0mcKf6QZ8BlwXB+w3gDr6vk9v/zjz4
UazDwYwV3CcOfHnyZzfYDeWKicGc5/+kV2ktznHJya4E4Eo7g1XKlulMVa894fyeMu6+8N1WF2kg
Cp9LHWGcv7VVRbqlIWXugqEt5dIz3i7dzuwao9gqcZEMQRvD3C9A4rcLqr14xuOY73egJL3e+MX4
uk4MMDVqaF8L6gvlW91iCNzrToUwGEQ65DKi4w7rj2co610PSNrY/yJHBD0hvm3JGF+pJ8oS9H0o
Mq1wlYLWtaKoxKqvNq0OnJDAybz7hyXTn+QXbpZo+FjyalWr3IkfVFE07YPZKEzmRYEyDnGbqzPH
zjB5mXcNexMWCri9nc/odgeWADh+B5vHeie8P5imYQsYPpI99AOLVo3Vlp3Wpqaf7rB6K/dXMbUL
U4dIWNFfOlwiMp/VSvtLHOqU+7EyoYlaHA+hpGyCc5nNGUZA0X7dPCZ0J57gJV7dRldDIvcQaBx/
ad0+TJSU0Xs157TlxbTYbfJ9DFPRlT6Z6yPAM/aED8Oity4C7yTJQRZtSTtxKrOrSwY0R5cMqAMq
JGCl6tZO9SNH5SRIrVo7cRv0TEnMrbELgtKjt7uqJRr5JITTHnPxVsRW0NGKZbd0dT9OfZJPDKMk
1ac2tT1CCEg4cfY7gWvGE8yl09Hx0+Qn2D0em0Mewn5L5GCvO3/hNsd3s4ObevyJdnozJ1I9GNFV
fiAREiT9NXkJkzGTo5rSkc2Q1tYoufdRsX5JV74FdZSvtKkH5MAds76tfHeri2K8L79UctbhsDQL
PI6yikuQqGYwHnGCagjxkhiz1pzZxugtnyDbY5lORGy6XEdgTbD8Nx1p2qqMIdYNB3qxSu3cel/m
Hu5F34gNVVtQH0Ihy8Yjt8bseni6Y4yD/YP5bDNm5wN4mFrY349ukgdqz++tOybEpjCgfwWlsVV/
cJ6V8sOykufUYi7eko0h5g+hlCsX5dPbWPbStk3vGs1/E7g6VnE9udbhnQJsks9Oirx9EcDpbfzh
LfZT+AZAFUreXZmlsK650CZ6kSnhBIdj+qk3xBU27O1QtF5KO83oWxGjRiPbw2XxEsd8SWQ24bXy
6WWAraNQkquOYbXxfiIoqSrfM+Tm7wEUIV283vkzc5ok+zBt86lRSuQXkXH5d2vv2RaJIQwaCt43
I0V4ACj9IECkKQ69E8VAh9HUxBr8LYLsdDsDpsqdCXWFvzJKxBuOawDt08zZd5iSXx6/GttNGPrU
Z8Nsd6TFiD4ltTMnmUziFosaiyZAgGY8IsYaTI5vsy88+lJTvhg3VUYun8TOSrStSmLjO3QPgcAy
YfllDHAxQhP5Z5kbmV/RddQwBhRKXRLKpoTPUyQXSK49yFSmJquNDkNOyNiN4I6CH8B+TPI5Lc/O
9V+HpToLBbKlGEr70Lyfnk6TQIZzAxuMjXKP6EqI8cL0USnZh2EC3RbS1jCsyFI++WVW3xjteUqN
tKvEVjFlDxej0QIjQq1Frwh6bR1fd+WjmB+ySkY3Y1fIoBzJWyI5TyEeNlbOnGjHjT5aP18ithn8
/fByOjnUc5KtksVNFG/RcTFxW4mujxHz5ULrKHdjy1VGj9IBwMtRl8Rt0K3qPneDtqK500WN5JBK
bNEVAN2cTgXaeg5C0s2aNSxTD4I9qAY7lVnP1sZ/XztfgpASjzdOsvupkSrALekUESE3F3QTAivB
X7I1d3gW1xDHOkkV0NIspBcuqyAeMAc4rBNziEJD+JtKwxPa/Co9I+GsFciZso5mouAO7PiNFj56
XLncZ1TxkrVKcCi5teRv/SaJ2U/Zgq48JLFayhJMxeZsU9Yb9cxDzWk0ulFKlM4fGmxC+B8c1pwk
3LvI2DLbgnVUn0myuoBuRmW/Vmm0238ZPq3AUlflTsPXywikOnlcsC04rOmYuasmpINOw6r3yVqF
7XnphwZkNRLHmB6//OlCgpYUkAvnnpm63cmWvoJJOQH55svtmsv1qOgoKX34YFQLgGf729anstrI
flZILkXOmLSFdT0lBK8PDhSgqv5t5pVYzU+VSJ+bz0pdr98qCz7b9QbfeWo6w0djAKR1H42IqWXV
MPXu5WKiYK3Br5TYhJHUwvqLmg52bYVIbXDzO+lBon5dWNd1qq/brJ7CrTfdHMRVQ0EHdtqwwcIM
YIVN9kRqgQIRnA11g1h+URAqYLPVEAo2ttvX9HPG4aLvHqreedgRapZ3PtGMPdt5ztXm3fExv34K
Zffqka9NYekr126qMtVXD6hDw80t5qW/kxUL3wS9bglOBCGodMPYoeLCHg5Wg5VSigX/0EGONeaO
b4CPyoD5k2wpDd85yARixncYFyaJalJlx8YJurJDryeW07xkeS4hmpknk1RKaL104XxfxJuumoTP
TJ9HD0oho/WdI1ffn7kdpphsH3kIMlt3XUPuPffpfpK5KlaVbF7F5GS9EDpDfOWqEQ18Eyu+aD0H
sO8hxu9V64KZkIZELSKv19pmyO0waugZpBnociztOELQUMdI1/qG0i0+AaAK37ZHH7ElRUEdqkcv
pMn64b0xk+p17No/J4eNetbfrK1GvZQ5UMelDTYWznXlIZTw5QyR4aj/2J/dBl5Z+9Ry/Cdtqjuf
LZXjoaHP8MLlaPiiVJBykswIoVQH01pr4yCUyvNDJXYhrZAYZsXzngd74W5H5ufo+eSFT9BjRC2n
Q87vrIQxjQe4D2I31z7Rdta7NY2w9MJJssgJ6FA9AyPUn7Bcwhwdbf0xUxymib2qmsjh9aXTGF4G
mwihX1PlZBincgwQ6DKhUn5nuoZtk+Gek6zDtWlhX55EwwWZahdCJaMuhVM2ol9T4vZ3NvwSJtFp
MEvokLGpi1rcPiC1UZ6yu6VrBqow84k4b3tR5H/enD0Y+9lLkT7fHex5LakHW65fSwOgQCVXt10H
Jx4TIMFlX2ugoUaOnKU+vm97BAJOkU++eoDKEiGtUbAtO6zaFkgcPcC1g6P411UXddRxVgXOzR9e
FEqU/lpJoUPzCal0ECoI0xQmj1tFtnk1ef7kzAHsjSYDIv2Y7pf2D6Gu5hSDlAk6oduBFf7xQ1zJ
aYPafyPlzc0pPoTVyT/gtHLtqHwya0H/KGX8nvHbqNR7iN9XI4W470gLLwE8drcJAJbvz+F9mji1
Ql+WdllzTdGUIpZHZnSrkhXrLPn3sewokJrUIBJI9/54qKzVsN9HcoIsiA7XsCkM4obiyVm0P1pu
apPH/+QLqbfKMMsD8CbsWpTLAY7OeAT6unbyRMIW5PrS4QmzbJtWaBK8BPBOhbKuGqhUt2WKYwgn
w3vUiqHH6zC+2wLH8pZd30jsoYs9Wrnfra7XLsoyGS/9Iw5huKnSB8tH/vvGshjlPw0VN827HU1g
VxnIvGwQst4yrezaQLrSKXm9PRAGkKuCCWcABRKhsTvGe8CoI2Hr01vz7YJp7IFY4JZC5M/39kBW
IN1C2z+brFT4sJerC7QVi60OFyggXG3JbR95AYfMboZC/WixBM5As6SNy5txp+/hVvRNdpdGKEW7
WhR6KPXNnhpJ5aeZgMZu+dLshhjSmmNh/l3c7kaTmC05RXrxnbLNp1QcO+MV+AKC4NMmyt1jPg5c
T2UL9FZZX2jpLzpr+C1kfqm5gHB+S6JAT+3rk7ub0UgvyzKHSJuwsCej9wocGjXCL3By0ehjpYyn
c8Djqqx4SydUNbJxfuie+TCQpR3KpMk+ug8qahlxr06K5ru6m80Fh5TDuqGxT0JMTNF98F6CrV5R
Nul5zZ614e1knQGHVIqeKhlbt0+X1uM6kvn7O2Nzn6ZiTAbtk8Qq3FZr6ldHKwxZgNR3/MM0DX3I
OtlWZrnNEzv6G6QJobB7u8ZrwiAXlKEBoj3wsEjQjkqpEsdlMEP72dWkAih2O08I+xppkF8jYxSU
YyatufqD1AK86r+2dj/0SE2PeBqfm8CADQBE1lW1Vu9Q4YKP7Egy8N6p+kh9fgRpAFneb+MdHs3y
10+nmCFlVISERZr7Qq274tBosA+d6HvhdK2AoVdexH8Sze/pf2cWLhVbnvPA9it0jOBqIB2NEnHS
1rGyU7eyxbR2O6gSXSqkMqJg1iDdKHsiy82UxmrtDpBYohlusB6EUxwww2bscv9js1ZXyMdS8SzC
2QDQGhBT+YfcDWQ1KxfiUj4p+pC6KP8cUSq1qSC23ks8AwoDD1RnBsRKDIb29mexmJmWn79Ix//Z
xfshKKa0ESY67qR37yhGsZ86OBToGQb9wU5ZJRKU5R71HOOZuc8HIauWaciIHfpXAzF306DI5RUO
Z10+ItXlTALcy/7QPrpaEamVeQE/zJoiST7x0buDdtrpO3lgVA40UbMZouJFsfXMpkdStyHVClnj
5FCxedXMmRbWoTMTHdirot7QppNVAyzJUdOuFvcCRWbUC60PPzDPhOSGlyetds9Z5GQmGONU7sU/
gRdlFzFGo8s3WyqtfmRNZlxlYPDIa4uHqkaJGL0y1pcIp8YOWX0o791n3B1VuATDq2zuvG0TdMk4
wYeD1iFqrcVhugw+G4bj7UDc/Xpn5/BfadhzqBmq9Y8GdD+1COgj8jLEikslj77OkPqHf6huReTq
xak860HNLubxgh/sohCc5xHipKepb3M3Vwb7sHwv/LcaTZllBpwe4xVK8z7cGD+Bg7RYaJAkjVmx
OLM5LzEBBNuEXZTW1ISqmarYOhClzRjPHg4Ndju67OSO8NfZkrRlneK+1myheGqVlQcqTFFXvDtE
Lvn3a9Jg9lvTHmU9NlsO3OE2N3CoTmuFP26eTvAwq0NP3QBzAt2qxetfC32WmmUH7tL/McW3AQZ2
3mp1D63SBnBNOtGU4/virlRlPfJAhF4Ta+zpWm7V6mEZH45tF7+KTL16zuQwfCq6gWoHJc3zety0
NsA/2xPcwyArOq9g1dWuu4wpLWpULFrb/FKjHwoTkN5JlytkGHbA/+h15J5+5STkrXheTS4LaBO4
IzrYhWEcrhwz1MlEOpsD/tqXEPND8y+8wPhe7kQZPvoVwKYilTcqLyJSnegWdNUrpHVuMEqpFj/d
kl4R78dSRppXHDzdEFqR7TtQyHIecCnYPBXHCLYMbh1ds3PaudtDaqzBfVH74dFYpwRvs46OFngJ
VVC0KAsWKGjOBoLoR48JMEs1vtkFCndt9I8Kc2TapE/I9DUUk8r/u4mQTHskRkyG0TESc7/icfTC
SYAFGcr5nhSS/JBkdyHWpURZG5VO7SgxvxuBQ26iE0FddQNU5WAuLIx32Nfa+Xr1TZWZ7mJf7U/l
AGNFPj6lh3gnG69HmiLTlLDSYogBgr0xt7AAKwqEYDlUe52NlY8P3GUQDpcHXA1jZf5FkUqCUmz8
7AZRqRrhA0OXhbRp1qLNIiqZAwp9sCCGzKB2iC5/jaqokay1yLx8l6mIMAhl9vWNb+QlOG4SNCRN
sWKQJQV6WyRRORGnKb5wiXgBRkGZA6aqy6w0rgbBGU9KXgG9Lrv1CRx0y/mfc0PttIdgh8IWJxXG
vbPNJYj07wb2jOljeuzT5VsI8rWDCc0YssLN+zid8Pr3j/WkEo/DhzqARYIK38AyLj8bqiaZmp6N
7osGAzCIIprNwIZq4+39I3L9eJGuS4Z5bc05wk07y4VQgUsx5GTVZZpRL6AvKt3tOxoCWyNmD1Z5
BvIMrf5t/g7LdBcRnzttXIfYvruiJyVwdhXKeawSrBAehX8Xo3zjvT0csCzEIlo/AZRjQmndUZI4
0tdt0cKuiDFn5IQjYsiUzNQ+ppA5jrxQSaCRj+AaU/N2BrHQC2NrppUOiL3CFGlvp2S5id9z52bf
M3LR6vlXdPpufRM5Xjar2L03XWovdv75Fa3BQ1ZWBU5uJFUQ4RpxaKB6KaHovMFCXupx5zFlO6+D
jBJVBC+o6fTYGZol5GS7wgiH6x1ttCcF5494uImQroeF6cAVFtjPboaSV9xou8EZEV7XqlCNrLTO
JF63Jw6ncks2dL9WNWm0M/XToBfZkiHdZcAfNMYNrNSoD4w7e5yxF61r7gZIYHq28qhwrz56VEsJ
x2C5H20qQX2z5i+axCHwETfOq/5cWqSVkXIxEXA6PF/aNjrT1szyt1u9DM4UYzWLRfdAtoBPybpc
NUCbo/Gch69w1xnAhA7oZB2ScVVeT3/c1RmiPfGoTMpgeanjke1JfOh/U8eZyzqxDvvBmw9Km8J1
1j0Rpr97tVVpTxBerR6amyycgnufq7EA+9PXhqw6exVTt1nECXrEONoeZ1b//NQCZ4I3TROF0lXs
c+81l9RS6m4l4Db9Y/e/lxSTFUPv4iISuJXBBktR0kIN0lMtLzHh3cXIoVZauC6i7S3r8HSSibvh
3+Az9Fei5RKS1aTjurF2hckGLngi4CYRDep8SPdl4FUJWdMz7Pt8c7se92VDFtmRU/Zo6oEu750E
n0R5zZlqblyKP8NSXsRQWxgsY80Q8mVl04gnj8ABChqrstSlnVvPFH+VhWzEwbFF9zsxECLPZgnf
DbRvMdAJ8lIMZjgxS0AyJeHvU630uc5+uWoK8BoE9NfDJN4jANh/TdCuXvilkfAY5k0puGMThE01
BhqA5XU43WH5DHd1gSsBUOD3idttc4V9pqtpefXYzTLMdPAwI5pCF1D0XfMe0Js0ysodGcl8uWFy
UIMbwQPDLjO46hF2EGPZvOIoIkRw4N0dUDIsVFbjf7Mtr3AzrrCpdrT8eOkK3WVN2uYGI4qSjMXF
zosFobEji/m9pIIHk1MSIaKbo6/aI9VoB64ZuIkNUx1Do8wrqWtVfheUafVtE45IT046CklAFOSc
H4ifIzV2oNp5oQlaqKJXLjdPyKLpfJMbot6NlWuNBrg0KCu8k/Nx/amMkMoRYgploQ+O0Vs4/km1
fWPUYBSSFGclwJ37pg4e2LkgiX2TEaKqzKxBmGijdAh3WRSlNfbpLKPJjYm82sPwoawuXfLQfY5p
Z7FIk2ZN/4vNzlAbWOQMnjrvEHjBDEKxDGgB1nN+TEEaBjVjNp1qtuDpm8u4J0n5uIuWpMIhAKol
P+eKWKoYZlUKx6PtcOYeHVuV1aYvN8nMBhmy/IT6sQ5deZRsY/Xv9YQeAfa0tCexI8utWbIjGknn
OL9Dgp/esMW0FIw8NF9HjQMouzZMxIZUgL3ZBJ+dW0ThwEqPmxLRHLyrXbcaYfmxzDcp+HRkplaV
Pt3PUf4ePlaqUoNDFT9F9CartJnIUktcHLHsnsKS1DzSZLtZR+4ByaJQHPlRbsl3IxNKOtgtqZGj
iXXhkHumcBUQhb+TPkv8gpYPjKtlzsyarpplmtoYpZAJhIRDkikHZNBsRAsWls7u985j9eUTgKoZ
JMv3B/UiBURPthGA2GU9SQnkvuzzWpuppLpPJLd5Sa+6Zqc+u+0EUUrssHg1OTlaHCHDYxqEklwn
pjVpODztAd90moUAEzowCEpPlhHFnM/WFKUdoAPwg3wgI4bCWgIaQkVl4ejFIgD7RIC/ZCgmLVR8
yLXffrctAWA7gWHeUKqN7YAWpx+tvjbtICuPx6p1uAd/540vYBC6qtx99C9V3vem5jjypQuW/dlv
43Aw3mIyhw8DH0mj1gNbkXOVBBTiRYEs7zf/iGN/XyzrwB4R9+orFNuz0c5+xFRjQV/AwNzq0axZ
TRrVw01R20c0cLMftEiJ6PII3qXmsQi9u9Qw2hXUV0Rc1P2AICZwax0MDIhM8R9LtmbAwXeG0QWj
6wYJ9Kti/xTTdW+AKl29q9D/PPMcZRQlLuz5ucmg1VCU0vbxLp9ML/eDuIDdTZoH40FVuX1IfNXZ
Dl/HfzOMCGaCNR+sVNt77TJxx8lCrQlZxeroz++Ea35AdRtVHCbeVY1E+Y+vq6m1wgBqDk2I5QV6
2wKaIIblrClIM6seLaSTTgdC83a33b/chin4xWyEtrrrBP1qgboHZwDhNrRIRC4SsNgsjYJ2AlSQ
ifEfpaxXUQ6YJa7WxYBl9QxYbfLqsvs94V6qOtjC7XcC3R9x9NbTzKB9fbfA+y4Sip8cceSJ1cWI
Z7ySgnH04C8MoV/4pYbubArMhYhP2iz1Vbnl4mEgBCGqjsoloSQuxcIf0dzMuMsAtYKjYawE6A/6
v5K7HE5VXj+XILBGTCx5pB8cvEzyyhhxEvSNpvmycebXRDQjwewvzP8nejMnCFZ+kp6GIM9S9PoS
1/imFTQ29wUXeADNp81Y6xCz8vw2+bak+IFYqUOMPW0sm8dB6jDJ4D3udn+duTh4ev/SPg5ixkX5
UVYlpwMt/DQAQpsnUoO98nxIr9ZbNN/mcuJFCozhvsLNnW2opnoMqewQBg8tZQhuR0y7YUMFX3iN
Af5UzJzdvl+ElZEuGDoJ8aoynjc8LhMj0gwBu5A9c3zNc/oZwcqSUJqXTdSt5dqzPWW1BkZqC8jF
yujevcHnFGbNKvSaaQY8o4J5TmdpyLFZPZ4hnxM+SOAZucXCIfNKScXa0ZEyw8dOGCgkbv+KQFnk
fQbHsV0kVY4GE3PbPiRthc1m2MtivNmskq8PU95A848wVmdNwrKMukBJyYK/RNumxmJEJ+2/wN+f
7wkfha6yamOCqka+mgfcWlVeEgBBST09WUg0jujT/RLFNlmxpTzn/SrUYdBMcNx3jbDe2kSpojIQ
zy/mAhYKDRD3l8dDV3Zm6bOxKStV9J/+7csQhrTvG+OU6O5MGARCEeUL9SDWbtuL4VU8nei1y98T
6L6nQ0oB4D69xZYtkZuXcyfyMiAI/0rLMq03qcvP3kPTe68dNiU0pXu1aXRnt4U4PFzBjNSMmkO/
bDEu7BaTa5SL+V/FTUMY3LxUAXT2q+7z8OzAHi2kGv2q/LtYAyLEWlQ62aPfw6mu7M0Aqo0VSgFZ
ETCIE80Z0ThB1ttF5aQDYbJDh20/4qDGCwM8eFOXMBqHA0EFLcaNSUbIlH6hFbOegAx4eWKzCnog
bQMBuoQgR6K0p5Jh6/pjz1VN2Lqi79lf9wvhsBtIGU9RcuT1GObYvpZn4jZ5uO3qCvrm84EFiSRK
DdReQu/VzkDKBBMiRRmTntlsDIq3N5OId/0O0gtltgeCL7hlORYdUiwx5Pfl+99CTlhDFK6+L0Id
h+gawSYL2g/8zMf0b+3TmnkS4sl5Gj9seoCo9CSkd6iX3G9AZaQ5cG+YProSKcx2105SUShNqdXT
+EEOTis52B24ODCl1QAA0QLlS+TkFhRlqay+0X/bSh/6fPMa4wcXLyd4mpsl54JFx48KPNWggkAX
VdMk6YK8bhk5h4MjgxA7qIvatAJa6uaw8glZP76yPcgcq8HOhCgY8+1GYQRp+yu48u9c2+GlFB+0
mrYWAbCpOjt+BrCArYnw5zIJfG53bi7LbtpUZVuYe5M8TZK2Njxzvbqvkp/RG9bzPM9dNALnISEs
Du6b9VjYO1KGG/DitoshzfFO93Dk/dN2BtYdGLy/q7BisCO4xEiEJ+Hw3A38fyCbdF7/vCJ5TlNA
DEmqziqH+EuJ/TVNLI9o2hCSatDr9ns0K3sEisiRdHbMqEFun3Xk42Gxzo01BYajZCxMurAVRMiq
XIA7ZX6jbJr4O2t1P14NZvGv5piS2J9FM3Ijwfu32hmJ7lv4VfYP1G3+qwtZu1N6m9/7WeOPV92F
3DqbGKH/cPzwzmphVQujLVHw7SnNyKN0O14Ld+iivb+4lCCCVokmiY6uZeySbLDHOvzwPY7QjJa5
ZFDORHJBd/xpv5jJPUWdrcrBNsKcVNzxy97+t/Mhn39u6ZwXAuBJmqDBKigylE9ydWUFcd0TQU/0
lXDkIN2P+1qxgV9L7ktVuOSH0Mpysw0kLkLjUWqSxxx9BRZZNbYq2WhVi8KRknKdOCT4vWEflf3H
bAa8jyJgbFR3D82nXxiH+tH0dYSo44h2qFSy/RbQjIGIGIRxetRG0k9jF2YvnPu04zSMcoU5wvJq
V8ApS1smarFTscTXQpBe20AQ1HwJgm5swMmmM+a8ZKCNugmG+K0UZgSXEYYi/I3/IF17Z2Gi0xBh
CWSPCwbPbGzt+lf4nRPsPNsSgmvbhwMgchRl3LBQ2sVQrjP3tQn5huqe29oXV7B8i2021QeqP8vJ
9dVssWa5ZVciJjpHurO6iR+Yi4jWMOZ6icWV2+I7iG39IcncsVWAb5bjzpTH6iOzWuuU/wmK/WkE
hhUYZciyjMGYhVxaSp6GmyEjb0anJKH3vDAkSJKZunBQZLRTWUTqsKDsRnIhJxDATAEfDjvSEc8Y
dES/KdFKXTC9E9WIfpaDfH682RwezHBRLRWahP2cL9Rxm43W24r5jHy0Iv4U6vULfyXc9ixtPjNt
two0+upntthojznzT4GjOIdVPNgiajfDF8UdlHxA+F4K3kE7T85twpC+Y7GxTB8uSWoPTcztRwFn
qBXeopGu93vl/4X70TXeFaUyD0Buk1XSdBZnEzfJeTp4A7M+fYsdVAObsm2kCGKztj99gJrZ9f+o
PP3hyTGvUPhoY/uC9grdhksI4hwdNRE8C+I8PE7FOnBWTySqFnWy0E+KNa+NloO6BsO3jm9WL2gd
LeJRgwbgl0vA4ASZb3/dbcjPb1OH8QpiZauG2su62u1vGAl1OXjGPhgjsNL+IYGbYl4j0txTg4fM
8OtmOQO3RHBvmS9Y+e2RRq6yimfkKDaBR0ZNevC5i2haT+opv/g5dBPJNl/Y4YFnOi+HETOnlrki
YvC2njOID4p4zKabyhXj66HwC8jOQBavg+RNcTEw/cAH5NkuIyVNTFunuulF8q77VEYNXNUglK/A
ChNWifZHOMMjLUJ5M4We2+AokHJLxwzAMJtUM3YWKlbTOZ3GXDW89+nGmwCsUt4h7HcaHPppCtbu
B3wSoElD3igelYOaylEr808bsUyOiH+PDmff+BcxvmHhr/AfU7jvyDqSbJg6icQaKUuBf7p4xsm9
mJwrkAOeeJm2mYTFymWrsWJFzeHc6snk3tzpDLibGZ9EPf3HqFEiS8660XY8KqvMT1rQJD000Faj
vE19nEUO7sFlbr6eVIowGE+Tr8I36lb9mn9Hb8Aji5W9JuQOPsN50ZxOUWilNLxZQviFGQZFIRQH
qAVYZGZ/Z+b9g8ED+ptuJTrgB8pjxirKwKcwZrAkSEedzfc1s1Xk2bv4qQk7J0qtfsryhpHZncW7
7a0KAyddtXN5YXtBe7/DCYRTvJ155n0duS+SD5OTuWlIF+BJlZB8HRhj2UG3Y+pLbt50tAivlIbL
EoMXbJwFADGHwZpvqnsOXq0rRSFrexqKoZ44mbAuyZPVrB6cVWKUw5HITPZa7XsEP/Apfa4Apvfn
lrCroVuWLYSRzR/SZIGUEGQtOfnKv3jygx9S+j/HjRF438zPxTzy7rioNpAt6r0kq7nZPEcZHVSE
S9kcNalhUjX5RqGJT2MRrh+1alPm4O7kzZ+CRbepHqn141Lawzfnk2o1tkur/Li6ZUvoOVvkUsU1
e5OGX0SB2xGiOruMHX8u7yxnKRFulriFUctSiw67uj2pKujLKBhVYRJoFHrdC6uhh6iyeY1W0Aeq
/EBoY6XnrzRhXodRzTxzAs9BroI7ZF4BuBIuAu7EhaqDL/US2LDjxDg67xEw2BAL8qABTwWp70Eb
a1aoFHvq5EY63WL9KCNHZLsEXsFQiGpQhBt9/Xr491PqZMPIFnIO0u7/nh9HlPWyn6iVSJCmLUwe
snQAXK1z/3tI52ENxQASWRCyapSZ1zFOcZoFLr7zcxWbxMWX9yLdunNjOePavWeWCsqNAo+PwzO+
JXkHvo+3jdDKOgbf2l396X2UP8cvVFS154WY34Y0yNXBipgpoEX1Q2mTpDtCUQ5r5Q+6kCAxcmRe
64v1BMiVGG5iV3O5uYe/t66GBbqwIUmRqFDcK+0B8FjkprnOyXTQO1IedQGqz8LkNW5drWGXHdIE
uhg5twxM4zNExK1LtwWiy4sTZHYlDzaVjMAy/D7WnRqUSvJrRmqMElOG59m0DpiHajN/VSBL9NNd
KBAyXpBp1Ys6peLp27FsRHILtlSopyAhSMNCV/na00qwDHRp56gzY0eLrjzKMnhh6YaLd9D/GdzL
we7qVxd/mWl2UKJOQRGdKm2hShfvQ35xbpZNi94JBdDgyArJvzbGKVh4G7KBlK/gvMuvWTkR7/NP
xLcn8QyTjoTVQnnl77E34VQ2mMrKtXsrI2+3ViiMRnKe3OBQg+cZZd4NaUeMD10779vjrNYbyzyg
oXe0lrvDSai7l8/mUQ1VOtxpsI8tesJBIt/dYeX5cansysYDav+fZ2XhCPinJQO3U9PLyOD8e84T
PVxa7O+ucaj5fw4CXRw93wWUoFCJlHpen2XMfDZwoMAicl3YGLg6+SODF6YrMabXdC7mGZ52/E07
Uu9K39cWiyA91RLaQdCif4bINjtjwlwyE2V+b3pfLWE1UJ0wvxvMfTxFQEs5333mWcuVH15myAfC
OBil2lWTxhXJVyItrka6N9MDthQ+qApCC/US6Z3EDDaIp0HcpExplwmmTcRJb79xgi7ojSRlw77P
UZvInYlBDwv9hLMnDvniw7gUsMFDB0wp6md7v7LPNhZGnAfuLZ3i45tyW8zKy+AaPBQsoydHY3Ao
dFnfskSNt2O5GwEZG6NzW0falI2pkJmeRwZ2LUCmrAlB4H0Mh/alHfvntQZPdzYD21QdkmOUJhAY
ApAjjh94pI7rn3XEJXOfEmlCTm8FajorkcdO5kF275jqGIKkaqc/9TVjkF396Ns38h2dJKZpb+ai
drAS3nepBkmqIQ3n0kocdl9ocLXRQ347SwuOxJLorwS1KpYlUcbKEgb45XIwU1jTt00f53XlXfch
74FZDHcM7sYfetBRgY3hCLKvlcMW0DbyXrpKA5RNEyd0bTaUBIRfffZ4odbZDEOi8fpTdUTIGU1b
QBVDtpT/ASaGoL/IImvIbWmmSwS4xgGZFh9yMciZh2+Vfj+yK24nQMOzMEwa4H6rIkBCAjA0riIA
kezilpYEEsYdXnBOFUpZ1gBvopr6woHaQYdW60nipkYwYSW2CS1V/5UnweCQUjrZdW05uAJ1SNps
sCr+OXOilKnIkevr920Q01U7NB2kiDHWq8n+PM9O3IAQi0siHd+yaGR5QoDNvFtpikgJ3XslIsLj
O1eRct3pN7f4U2H3rSnLFXnLocEfXzArwdofhrb9Zj+cXGaxm2CRk1iB/D48ij/HUyMHCoVoPtou
/oBrjS/dWTV7eab1DFlNeTtYJ1V+jOkymC2WUCnNUh23gjEnI3PLf6INqZTYAHwzb/ptYqh966Wc
90Fzl0ZY55JY2LBkG7533hgCCj24LMes1arGiW2pRaHn/qHVnotNvDDrbF8UFcjtAtvFWW8FbRY5
FYewXRPLY4dLhonb0rCPFc5wQnGbiehTkGq8xMyom5PoDS3elQywf6ZHOBqmwRKBzMEWTQf0/uh3
mTrFglB5767kWrC2Ryne/TbaxGM//pPoe510iLCVXw2UrfyER/9H8fwmvRDw/bgYdVvSrrjNLHeR
joeX6J8ZbVsBhBmqcghj2GkcNmtMnKvuUOf2J+rfs/oH80HoYs1cWYtE0HussaVgnt7hvbVlcq6m
q5Xi4WZ6yE6MFCNPa01QmsyEWuC0DrC3+8mT21hTxwQ5MLJz+QvQyeeaGsPODZq2FqH2LC11iBmJ
8/+E4JCc/0J2fMaAKCNQW95aW9QaRfZfAxZ+SYc+6imE/nrVO7qtvuIeZ8a4K6hwl39gY2JSOmg4
RRgdbHGWkXxvHfTlqzLTU6aNCJyieFLcx+ha/NaxWsWL+3CBFukQHLM10+cI3AAkv8fDvC4fXx1R
/yxHv/irdZ3D11PWCOoQ6r6yNE9dl/XE6k1505wia2XjWRSHjRIg+M0dduPL9weC6xqfHbQPAJ+g
d6gld6BVMy6Bm1i0pm49j+vgBBX8WzLxBHQJvRjLZ0EdR0wRJMbQUmV3E0/jjx8U0tiKlFGri6ad
w4+cZPS4xfks9DgIdKEw8XoXdHA9y1u56gprpwez8mx6cnyzw/MGMQwyDxdDMiF7Wq1ATXtdD8hO
dux2aaugePeYuzTcKYVrGK2Fun2Zd0UjqAL7tJq8tDvZv3aeweaVrAm3lwa529s+NaApDXA3du4d
qlCnVJ4vZyEa94MGrvT8Ro8BNYztpNckFIeQ9zpy6bggKZE/nIBDnYiFI+/jvbFVbZuYjgLs3nsH
yyD2+3+AtoID3kFecp7Wytmagl2mW5IyBPfKz/ujdCRVKbaHj5tSwiy34H5nHkc9PN6Sn+VegPRa
4bufxFQSsol+JkvHzmhFDqVjL4rq1KAeB0K2tO6+BHZ08YUIQqSgRK3W0ebTDb4UYLryoILI4hF8
H1Q7h8f5hCImf2rxG4hCBknecY0o9J4eEKZ+47hkuPlVeX1QFL9UWarWA3AMFVLTBLItdo6hW9y3
WVhTkRDo3N35e52ZzdmhZ6jcwfUf9grL7ifId+S8WR1bRkz9Cvb6nf6wTkxwbwtNMZph8wqINnXn
v8aqSkEYZAmynPSEgrFfod8QhheaZKUhpIJE0QQ9Fd9r1MI1idTnCMx8Q6DCzKW4gD4SVxDaXRPP
FrgW1qiNlWwkNQmL4NadNedl9QOoGhRIxDmUVZZVtOslcoDj8QB3WkJ+88bDtMXDHg/JlJ5EIbsW
bvPFbLnG7MhMUESa5Vuh4ZsZlTXbXtVeQvz46FxnqYnYZfoy1rRJvmigqM7pt2KWvytidudiBsmt
hWB9O1Ugvk1NXAYTzRU0bcEs6hZp6iNgz6Sdc+6MrJ7x+9IPxOVGKk8EAXEB4rwUrLYxXuxzz4Gm
YwLh2N4J15WZ7ebY+4X9xb3JXJdSPJTSviXI/cY1fL+k4N4eRzOQO9ncLRdpvVCDFGvyKCdtZCcs
6Cbs44Xhjo8t/0Y2JXXpJwbIQzM/pkMYV42miXA6Fo8Ev3ATF5z2JYNGJzJX6GNVS6QvmNd+Zc/0
yGUYIRzxmayOSY6oEn3RGRSRznUjzzFyKQRVvytfA+qZA1Y0Q+AE/5uZy3Z7qwTEn0gZkU5c1HSf
sG/tpZyIpPQc/HtbCBi3aX93aA5LDjkDOv+o0rIybUAsffVlRurlv5NlPlEurmO3mnhfxrok7Vp4
MMLVIV/q3qTV1ZqYdENcsVoiZ5rt4oG+yEUd17BzwY6VMyPVpIZf5BFVorI90exvEH5TwXyey0qW
vMEBRL+IqC8X34LQX8NMTFSTeAXpbCJ1RpC4GkgsDnK7pGJQ3POU1C+ZY9sEOfXYidIXsw+yPpVH
UWN65WZCQ/1cgYQ6SrINFXfr7690VmkoYyemBNSDdbDERwp6Puniuwzw4Dzt3ZXTRwqLFmutaACs
vidk3mcX4v5qg0D90vJKEPH57C2GD1h9GxjyGgQMKGF/c9sHUYB6s0cP6ZMCwYT6v6hfgtzvTHvz
gIg4dSEO2Vx/E6pOxZM5sD5KwJlQfIZ55r+UlizVDcWFXPC0N/6DcU8wd/e2+sN8gyah8ny+wSyD
35nee6Sb4GHOtpQPzAkU6ZfDmJk3LZAcB0oMAav1MnwgNSvl6eWN+F8QL7Drrrsjj0EPg+e9AaVa
FIeIzKa3oJjdgxKmn9+xNmBs0yrSCDizpv1SOQCAK8qxdWgASZ3g8n2H+Iie3p0W/iIXF4g0QiJt
KBAhbQ+O2l6IU4K1AEc82hj28+9dCx1hS4JScFvK4kX4U8/qHsjbOUNNieozt0k0t5lZo4xdg6cf
bjHfgm3CZbCEcc2W1ywDP+5YX6tVO4TPKldq1H67nmf+NU5XTS5N4zXzQbCSSfF1k7xgvmUG0ZBQ
ESONM80oAgw59v7X2judcN2TEptiEyBeXXgoV2DEiZFL7AQIxHLCVtGURv4oG1ItxwsESKX/8d8d
NfRN2tXr/qRuC0JPd+Vun08AKmpeeaFbsv0m8u/X0O61GpBG7cB+rKA6RcfA9hcPzb4wGBt2NQF6
45SQYFcssDpkS+DwrOmY9d5Sl+Y0uNeWZM6Pq9EmoFPeFGGldvbFdyEfEV9EVYGFN7QBc3/aaoku
uNYm2hnzpj+2IEYfBQWieAgR6VlaXMMyaF9sXBRR8f9gwNi2vKGnNL/86wSNkjgFSOrqhrQOV2JJ
mNeUJbUGss15yXqwtefq1QL1xoIejhunAUt0Qf/NkHvQf3dLwxPvrCPu0BPHfiJOctGdI6xcm3rj
D4ZKf6LE9vxfAN6hZj9T4zYuPdSTtXKynxEBaAnHOpdvLo1yBtu1631AStl8pGNWPbfRKY35pppA
LFv6ZcXjHJlxfrX2II2fbpWmdUVIVJdLoiNpxz2l/HSiz4CKxiD5MVDBcN9TVECgyiFzNqVzwmtn
IyyI4qER5nEMyYwBjpzzKDNMjrYAyVgwqHAVnkcjnxtzAUyaxjB4oLHDevYO2iGmq+HmPwP+AEuD
9rEDVOw75M++tNQNuAKzhqqlaZAfY3dG2vnRvcgvmB6966O5qUNIG4hAZaWpYTLhBJpKwIvp2Zhp
tthUE3ZxVtFnrb9MIvwCdUfnOSSPZ1RldcjRZRwaG6tzNckuNXQgIXj0zb/DqxbkSWpLAyLY4MFx
4xkhayfpF4pRDlqJcP4yzd+0ZJTyM1RRLfvqmozmYFbwjuMm4VQZX6hx52emeiiUhZGH4Ac0Pl+6
0EgAAaKw7gbmrP7DwET4m6JTKfuMa7xltbD3RAIrMIxqcDnW7dMqIdWTCH+uWX38XfCmWY8ogS0m
uaLTf0AuhiNEUNwB6nztKB2BWxUGPtmubfd3wqMqOJ1nsOYZdS6FvMLSlze6brvgrRbFlLDbwr1Q
zhnas3fqDBk+80cqOQ9pKPLssGWV7gPbIiBW8wMjawXiFtIe6bm76siXGJLYDcatNcXN7p6q+OxB
iY0nCr1u1MlGhJnCnYxE3Q+yLcY7Hj3YqeBHI+H2Bap5pzihW1piX84dPVlPkMtJZ7lgA5BYP8Dn
abUVnYM1khcHIY5QHGfuLmoCD9DuHqg8KoUm8Mlh8oSJ0JG6JpeOjTe8OZRfvcljrOvsSSagX4T7
CpTgCiWvcb8d8oFbs5NZdPsCRzeIAOH7qYSiDUE+xkeo3+posBuochgPTp014EsUr7wrNtt9TPas
XpvHqZRA621DYaGv7OFj4Gp7F9oyhN4oGCsn+0fMXxMgReUelolNFx/ik/+lqu3X/+zEYACgTwO8
iXKYyGy1wKPEOARY/gR4ONJiX8H5hQFVeRcGQPdWwnVAKVp1nbHTOP33lKv3t6r9tS9UmBlcsl52
Zz14pMuEa0QIOkUO7Jd1IEEwaR1wd53Ua1fUh/ouI13XqcfR1t4VfGdaFc2/jd3nPlOTnO5MKw6L
CSWFyLV8d8ZqUwV0eJ/RnePBkZFGMj9WdwBsxmioyRf6mi8t5sxf9Yfd11RsW4ZPJpa29hCv+azN
O5TA+2Tc8ZtTP2o/Peel1OvYrYNrK5F6IBVqyfQczJ2+kl9DtnFkGtcfiZbaJFLPt6WoGjKHkhpr
a/4oTobYjfGKeFDG/igmB9Thg67eBUIvIQRzJ2GHQx+YR7ewW49Xp2KykamRH1nIAq8oggm70Ast
sgGjiHG4Gq3tWjcqjyG5KEf10RAxMCoA2tqa7HuVlAee28Oiipo40llWypD3/qQA3HdsCA8Ft4cg
E+BS6azsmn2Y/Q8F5XTAc3kMDQ8SoWVw6hmvrord4B9EEBSe16IrMLUjSMWxH5sJB+glbwSunuJ2
mqApRJ0QSpUuKfuTn/CFgrOvmn1fkGou1wQtBkfUXJvfxABoNzdb5sao0fBMi6zaIMvPjbBs3Trv
LE1fcZDAftnOXm3dSBNu7J8oQh+Gi/Dh+1BkZiM9pOQsN4y3s+kOYEbzfDne5/k9vS5IeIeMDe3v
NmE8bGuGUvXQkNM7kciEx/Q9SCZ3piDQMajr5YD3TIS+P3PnG7odDIODKbCrdGmJai9u7bN9oPHT
TywkUa83FULb1qzZgwm8Sj1kyjDsUd519/s8imsZMp0RJXGomjokf9IJPLxNHX0+DgYR0Rtsa9UQ
atlU86O/jtWZRFme0qM4QRcmGy5LcyjH11KZL//0v91NELDDemYiV8JmH0yFCbheTOnG1Y67uYEr
5V096W9lNegwPPpysG7VzMjMtGF2bCFXqADd35MPNDbpvuC8/KZDlBhXCCM2PkElWBJRPFQbXQZl
bYUTvKyEeq2hwXSukqK+CCZRps1NrAGtDwRL4QjRi6NYPhAiJwmIf74NZORYN89wT3cvDuWXLpfv
6eN+k70wByiMmixV6wYCvLGoDL0WQvSM68T8IJQ5FJjIiB6kjoeLWC9N1BUi1WjsFVjiLYcxab+V
fXRmdspOVc5yljub+qyvkbl4fcU2iskHHYHziZJDqt+MR7tLtk/RMknWYg9tbEqjQ5ffEVXcSNML
Vefs4ULw5XIRzYHy/KYwMr6+2QYzZv3Im3JyBqW8sNE0ElRy1QXBcNsuOWQDrMObzLwLOOmygEbt
kRhJVNVP8QiC3OrpCEP8NLE4dfftQeuTit+XlkWtCmE1TXfm/p3H+KlKkfwx3NHxGu73AKn+iPRs
+84bbJdsoW8sVXxR30f9Dm46bpakKEenGDgsbY7VxUz7cEYgKjR5p24QYE/NtNV2k1fYMUTtAwt4
Dke/sdcMKZH1Pp+qHuttNHoHCjrcHYGL5TjrjU8msi0dYRfJV0GPOWknVH6IP73pUzSgpMI8OWgj
3wtJGTEGz+HbMHuu2hNXo499Z2N3WiE8XUAQgFR/ZmALIvicPJPTj6SBIZH3PBG/MtPtJ3Ng7ATJ
bfnK0TcrJ8+mPmHKCwwpnJfaPrKyTKKPUoN+LzNWocJvhhQxAAL1eAoIbJXPhYrk+96VAwqgA+qi
PCpxcS982pEZ9FONlmnXFk2jv4zI0Nv95/V6OEIRh/hZHTgVRkxtDfmrINr9rfpGAZDlMtLEljyk
6VKQo1le8TDBKh8bRvvDGDF19d9BAopzqpIjMw3lGNGMyC5kU/3nd4OBlFJHt5w09yBxFJWAS/oW
8A2YFUEan4L2z9/TpYnsME7ptFmHSA2LGqd8oSRt52vMw9dCspKv+RSVsAQYzqtU6vKGPjdsEnvh
ir2RQ7xxMk//fLENWMobHi1ega7M0tRhixOoW8mso9mqFWo9gxjcQbKLEg+CRhnaMxe1TFm+lzFP
LBiUr55u/8UCjYwYvUMP0/UFPfTLkslg/zLV3v9fxlle5Gul2b855B3BO/WoqzEg0lL8DRKp/ey/
omP1qi/dLs2qID9He7nX60sP5+AbamxReHBGK3UpRj9h9OMNHm1qK3ijMsVx2GALHipI5tsQ6R7y
pUvdZlhZorBUDE0yH4l+rLebIuz76we5cl2arx8zy7CnaqF/zKiCq89B6VriOc4Opd3K8yo58f54
lOd7TB7mOsMygzDUP81QAh8Q+6pOVYr//4VrNpn4fBGYYYg2VVpZbjuBikZ/sAKzEc4k9Y9+pe2p
91u9WPMNBirwIwJpSw5yBeprXpydHoetmJNdbRlL6HiXT2XhdqcHGoMFyEbydW+6MYjspK5DJFiV
YSj2ZDWfqXa0ayqsZepfKZWlvjbi83XknaB0Y60FSUDEhMLqhu+ZSHh9WSAtVpZlry6IJQdqslt3
COO7ujZMiCkueSXGnH0fWBj0XvfaEKFh0adCbgXM4x+iVUFaMFPlL3GpwP+Tlylv9GNRlXWbqr7V
OqDMdATCSVLQ9HMxDm3DfEt+VJB2IYbKVLCaP0KMMQKvUF46GTcu0zeLI7nItU+GqxtjPsaFBt9d
prTKmynjfSQJWcmsVle4WJOH6mOZkPSAoCuUwzi9/ayH+oFO5ktTykaasv566smDIgZDbcoTtYDC
O5vTV1dzokRZEDxKPTVhASM2T13uGzEa/sJ18rk5aoAW7caS2odKjFVK4f9OeM+XBnmhWfK2OjRt
UaHW6eTWkZaOWcCwm+DNama8UZb/ELpvRe7SUSNxfwtugqLHAmHz8mNwKVaP6F3B/Hvg/JTWiCKN
hGs/UMMNX1irHL5Mr4rj6+ZnsPr2l3eHrbJ0un9sQ43Pg3aN1pGdJ1nSFvJN6B0rhuBlHb/kJgVH
ALdx1Whizp/A0jNHGtf6e9STJDLaTdXg43+5GyYNbRSiIIcI4uIx+Lh0CptFFGrH3mcbCc0ynAiu
05pW7p4eKFrzki0LnuaRDfCzAG4myRfIcNKaiOq5j70tTeqF609S1LbdKzkGtH2oDaxSeme6VN1k
rSdCUwzMwkNW/dHRI8E6nfcahnEWQ4BVhtudB2IttluLmy0ONAphjtdiND+0cFBCkjmHwjPiWP4t
cl6/7hoHp1eRKrY8cmQQdfiGqX7SFaYaJWiN/iJBb/AZJiaZlzzfnHHqWQqOyjzSCLbhz5ShIuFF
w4mAXthxK/bbXRtm3DQZ5WwqzX8ksHE1zAGy5aNtL/NjcSmm2U4OofyKdUN5LIgQuVEKZ+8RI07p
MjKpfqBjekvo3E+BnXPG9gghG2sh2yD96chPprv4lcPPDI1Lz1nkxfJQKGS9TEYS6bAIGFIFzXwd
+ub8xB126dm/Pd30rIZCycALqeeYNwZrNXidh51BAHEcldb+jcvH5W9y6aZitUYdnrfKAW56BcAQ
iunRdMiihBkmryJY6wOal8W8Dq1m9KvFPUoutgX8CYLxW8U8vyPcXYd8uhY0/BQus0UVC4O92HeS
IU324hpH0LgCvZsW7FWCBLdcvfxaHPHsLnDZsuqfjVHk3ySZiIAOC2mmr4IzLW6IqLoYCJWqu8+n
sNuf4UXO1ogy8LIZzTtvlu7veT91UlDb/2AIytClkL8Ix/DZouUMLNZpOkBrG9ASb87IJa+8Gcz4
84iqR3Mabs1+dpQeuNpBwjLA1ykPm9jUrfxoB7K9MtzfvWOgNk/neryLkh6xSop4y5oAzOox7W9u
mWYoOqvIeQiRt1M8Y3AKCi8OVzIro/2qzBdoiICVr/oNBoNXGKIabX3VifQJgYRdY9FlPjFwHXfR
OORNDmAr+ItBHun/pJWjfjNmsnjr9AI5HEMTVLAPpbOFD2J5Z4fnNiCojlsH/Di5Hn9hm7FLCl3S
Nd5mhLD9Borc+bBpwo+//9yUZ6G8FVZgn/PEmTd3v0/+1rZdNvisKobWR8tgSAbhrFF82ZFALAVx
OGT7OY40mvogiKH/36v3Hwe6WajdOSA17yMSSvpHUuKwX7P5NrjSxkyk1B0e45jB0lGG09qX+0gY
JPGLp7yj8lq19rsYEcyhEGiHhWpeEvM0vwoMyh/JtV08mMLkyPsc9ONU7hDwGSW5wlWiD2ETALh9
n3CWGtevV21JaamG5KD375psePfWSUKA7FZYMrG0GqNlceQPRe1Zlp+NzxgQd7a/qyZUAF1vho8W
XSMMPEAOiOVytHxF8CaAXxcORV7R+aIOT4IainykDYOp+iM8o1Oc5Y6DbUBRnmsVcG2zYg6s96HT
c0p+x0ByDJAs2X3mvR+qA/qloc7tkur0q3pBI+CwU/a5tOOhdC2d9GB3rnVvKJxPpk0xRSoDVXqi
yeBYyFEUWs8GGLG5IeJBQ4JmiaAtTs0ZEBAn3LJu0ba4dVcZEmrr4igOd/9IZ9uSt5ImfGXYDKof
a91ZQ6NOVJZet/eiXMHEe4uQ/vzrZ8ZHfY6zicLo+MvqlG+BuH6/2f6T+qzqg/G4KUm2HOnGEzqw
kqCBbC/7Wxd3HIw2NhQnrcQAXa+3e+qAasn2GksDZvbCI+Xdf7aqQI1UB7OHO/UwhzuKb37SLbIA
cwmP6x4ETI3g9Ip8y96uyIXSn+Buw6bD5kIdmPIT+LLv2Sq5BcveD5t5JnxIAYfH+VWVxEfNYTWj
NKf6BrZm+Iob1Sp+iBM+4nue0Je6Nq0BS+KjoZ1xeULlYzuyjmqNjFxcoVpgynfELPpMrjum+INp
9qj1FSL3ig2jkU/ONPkAbjSgEdPi9eBz/81+keXDL+ZcffFwIyOC+B654nWZmeiwOQLBtx3cyy08
5XknRzlcpLh4/3x9ahUv+KouVWkc3gEKmt8rAnt8+BjFPbFDoazqgf4EixEW1KTEZy6pb3NGxJed
QB/O9wcK8NvtATdwxl4sNfU38Sjp2CkB35AK4B2xdT3bRmxa5EeAac+ytQl1DWXHBhQ3YWjCmjTD
pElHu84U64SVpSg4KpGQsp2+5I6Oa9EiC9puUhgZaYsgHQd6SjpZ8qePIxrQ79tUoDHBrWPwpKi/
u3Kv0EVrwtMAVYcYOjqqv5w/taSThkyT4nutXQTyRo0xYIVdQHYebhmLXF7tE7CfvVq2NiNuA5Jb
ciMd9K5HyIjh9SpdZqr7xtnhqUxqu8jWrB51/fyV+Ov3ur1CDOh44vvnsa2q+FcS3Gvy0KFfF78h
yWQgL6+endtx/LR35BVjtYTjFx3LVb/2xM9lLXy+fW1lUjk5VCY5rnlM0i9Sn9Y4vQ8RC0dfOkIv
ldicLGZuuQorA4NDTNiMBHr9uz06JCW1n/FoMzluoWLPMXqz2M0voC2dEsDziiHZUoI9U4Q8+x2Q
F51DdWWPmNb7DHxnkiX6hMkKn3c4hRXGfqohSScSCdKSxpol4uK0YORt34986S6yyayohBczuyrR
E5SPe/VMGsLRkY0xqMnXGeqcWKbubbvDxgTslfoZJ3c+roT+ebw1lXi5BUQLjZHPAAyc/H6PI9/y
Fz4ycnBqn77vXzstqC9tMxxpm1gfnX1yrVnx1ScsHhFWORXaYx65ip8cGMZMCGqQKAzcmxRTOTy6
nUZkl+7Em0N3NiN9qIKRh6ElKY2kyeH+R7EnJuQpRaJJPvCf+tKwcLaHqrnI9JXs2+fg7z7UD3+d
OHB/cgBoFZGZTN1FCe9nanFJ1vn4ee4Y251cKIwa4p3kMimSh1hE1yAROSJ/kYX3eVnKF+RJTpoP
RFAXH+wjn5xHYgSlLZt4k/YxO5WMZVdgnnJGIB+9N5lXnXoTOKlMJj/bufDIGFA5BC9qufENrCg2
BSNoWjonMF8z7P4YxUpnwYxpdmN/g6CQ9meOdfYeAjpZJU3hmR6/8WfnEKK5iL4/wh8JfVzbzLul
5sUktyAOfEoiXKciNoPMcRevsCjCCqUaO7dqKmik9qqIarsTpc9KL7CCaJ6+8LfGMkazcFrHI0AJ
qUb6jr6B/Prv62PJ06vPeEEIGtysAnESMTkceKJK9g2ctfpClz2TnmAlo554n740bTSYpaWnVCZZ
Q48f2zROWsgcoSG6QRD6lf48FB/dfaD92Bf928r0RkK7sK/n1Zr3DeiaxecKR/GUVpK4alrOLPhZ
iulmPG64jTE27UQzuya9qmKLHZpkHAxAW/pJ34uo4bNhTWBRZxDJb8JaRzLZSEKNPr65Yw0GidnB
UZWFSZBYJMcp99wc0mHJjqrRfZl89yYDwNfeuNWPsjIM9+UjRsGGnO6z3SE1Rmy37A9Y0+4sURZ4
3Vy41a3YnjTGUqpfc16hJtzRIbZBlSqXpeIa4MvCefQBAYrCCgErGynawrz4YwMw9cWbW8ZtPb6S
FWig+Fevu46xWTkPRtGek+UqvYxO8LX2Y1vmlCwlL+O6eSf8C8WLc0lbQRdPimqYlYzuGssq8qHz
O9Ou201YyZZ6gvSor7SdUAX46Kliw80rBwDpbYFYO/1ySxvPQl8t7TwBiIJbnjJq5XDQcs+CKQwc
90leWKAUDZq6eOXI6bFjDlUkcZ4Ioe5IgpgOGoEEzFNbSQ2fGKhn3mga9whR9whqXozUkUKmniYA
BUUG2tpHVJiF3+oAff78+V9LIWi291Rc4/KajDG88M5fydrhrlCW5SpKCyyG8hW2/vGc1LiG+yIo
/VYiXPZlBWhx2+L5gG3TjqRyKvm/WdqceZShDnkWvjNqzKlG6jVtOXW3BXNiSjSpx8KjG2LNPgJg
V611r13n+vHSJS2hPCbzHQ6sD+YpSffBIJ9mptKHySiArZEpdTav+r6b5DzYdZdeTVcs8P66fjGG
DRt0jGtlTMWJk1m9SotdBRQangyN1NG+7Zy/Op5Dh20/dFvt5+GU30LtjHEFzi7QBFSrQjGMdfyS
71UbsXEX21ochMjUgL0tzUoag9x8FkUOdkOB2ZgGXw2sWpFS+KE1StiE6oUXa4QnNWQRLKT0JQ7q
qYNzPvFT3Q8182VJ/WZeIOAuzIjzGnLALQozeUZYVtiOASTz87d6VDAaoyzqA6l+sE3bCzQe1xJA
TD65TKlyQnO1ym/S1Rx1KLVZZFFpovaacPbRYSWRSmtaTOh79JaFWg+9y/I6alDQBynBPJIpxsmi
ceGPYbyVWzxxS1fbqjQiqrrPCuhm5TXH1zJzWQJZe5JtddMIwzMyj5+LhhamP64U4+valWQIaqka
8x3m+jI+6mrU0QU6q6GgZz0NRsH75irHuCrNuOR457ijf2OAkD6e+eVQb+pzxNiQ9onmcLaO0sCb
UVkSM9hFoOTAhQKYM+DDsy4MZfouQXLCf3dbkb37mn8yhrE+7UzvEMcJrVQaVmvZe2iPFH5EzgKK
JgLKEPG0a6YqW4q1btd2ZaEInMyzQeTzocdOkKV6OzszaY4JgB7H7apx2U4sib1IEHmR74yql0KX
yYkfkUwQ4kMb9quGfnbQyxeZg0c1dj5Ec1CXsWVK6T9a8tnlmm2cl9An3gRyQ5ofGLIGh0iBWhzw
r9hA+td49/JrMJ2nFa3JyMo9h9XHQlDyNVOLnwkeseUvKFXbpr82pElr7nmfkhi0mPURyx+t91Mi
RgnX7RCbTs0eqwMlQAc9SVFu6KGIXC1pJY7j6pgAxcuu6DPwW3lEf1qViCtlaH67IKINhGtIh7Qe
GIu441/liupXgQwgW9hoVfv2MXphsiweNOjEGlnMatKnJBbkPVOwIiYFWeVk+WW4vmBKDD/yIcsi
Ng3f4Rf7SJEA64y1yWI+9Yc5fyvOPvXLZwcnQCGRXVcmTcVz6DNQvIJHRfP4MZ5fE28mT8Z7RaRE
C+nqaT6tTaWLN5iEV81aYutPu0Ebk2/HyO+CpOVadw84U83QsGlgFjNTZ44OTldPsRoJSDRpKJrV
HTT6U8t/BmxEsVtT0FEzdvXiqzqRUSw9IZc+7FcMoB7PS0dPiHQD5BjgcLMUFHB473I5qYQl8wNe
nem2s0PJl0NhMgDpfKnN3oFfvNgLPVk18hh1np7qwkcJqvmQmSARwvX0CavYkH9zNaydiIqpAd8s
pzsGjNKgIfuIvIqGMJ62Yfe6U+R3R4UezSMdPkwWSn8zah0nVDjsDu+HIos/X+29IdRPa8RGBYsi
+kcn6efLxD8GVZqZ6wtqIO+xzjsdApti7W1mePezC6EGV2xewVEfMY2UdUUHZKAaw63fTJyrhrJi
evfW2BTGidCpXF/1toAz8iSh3EuDcC23zsCcPXAA3EwtzvQYmEQ6ziKmiCI8qmjiXkrXVIkZRjob
lKCQBRQ8lunLaORgyu56DIvXeVVxyl8QXCVMYJlKzYhrsSdf+VH+Fa+hHLxknGmkjWfsEseLjeoh
b2kmbFk+2MAK+bOv/gDgoT9t2oceli14WsFe496YBEn6h7rdhxlOUZ/h1vLmh+XxBZaawJ87xKjf
Z0bOmocwrlueQEK/+wEbFR6boMMbfXwH8rXudhTczKf1LaYWKxOwyO8/Ws+qcRli58iZsuOpC4us
CQtLQUSaJD1+H1WionauVvHcUc7PQvvPd2VNdfst/i36/sZkp4CUJ8r9fRe6HdfhQrqKkXCCFbH5
sKxbKKaomudmakHx3a5WBbnf5AW6DOkTMY7TAOPHhwmzE2hI31gPySWSTJu/Lac3pcKt/8OqZ135
YR4uNxBCsuj+BO2oXOCZaPQ8SqJSt8ifkieWgys1SlRalgDOqBy5ygXLZNKgDkKVfck4nbKm4YuC
O03FBQUMvwS+KSCYzM9VJg3asNWecQitNCSAc5BzrfSY2DqHJevw1dKucwkeJzr9LWvyTp/plRFY
7PFsjYdwj3aO04dxtFYiSohpllalUx4Z08LpxqDcKrxBuGF1Qtq/1Sq2uP2Xe57t8mzTKEsmg1wt
UvxFA8BhfbV8N5GRNhH6wc+5XhutWww0zKvColKHmYzLKWY9ON9W7FN2bTzYKuPma5vaakI+fX7Z
5yM32+xQtJ5Htwh1eRqffHlCwAke+f9SxZaWtwz61fBQBLOe/KqMLVKDjHT2G3KpC+RvLIfruWjh
apgWnZo/YyfvmVflfcEjTz1o87Z9+EB0aDHusqJzB7O1xo6RyfInwTvx8eb+tXg8uUBNYOpwuHef
WDC6VXl5sjF32MqiXu9WsUXF26b5iYLehdaxiAI2nG3ezW8de7B5vfwqRyFhi8fx1ZMVgclXrhYf
f92/R3rBZNKKIMwGzVhK+akn4Xgko0cGshfyjpIZsHFD1TcTDXIPeG7g18WLwj5lOX5lxp/ZOosN
nRTSrzOgaY3oYu8gz8cbogl0SQQyUoKWHeBgGH62mrd2SxcguKcuU84IYJuijrZSA4cWKHogs1i3
1FGLwP66rYyjKyfTqRpKGEwnIDe6UHLprsOBjBmDuRcTKDmO/h6pk/Y/s83ghuDXdRzh5JYT4JBZ
gYeJf/Y5amWWtJg1FVjex006wVvl8ften/fCy1zlWF+YUKE34pquzwL3JuP8irN4QxsJs2XGVHKF
C2UxQZ7zLnhMQJW7X80hj5pUYPS/7vi8Pq8P6UNxFHDNOV/2IiVGjn5U9/UNuPwSFP85efHCQZ6V
E0E5UL0ty/XPP06mpNfJeWRe6jo4N9TJ/keu0+C8QTyHiQVEbzgqQq5EL/jqnNfj1s3b87tuC7Fc
ZZ3oM8RaS4eJsUiWJhh31mGpaQ/L8a2sgC7XYImoFDeKFer+JQYBJDFpJxLQNj/8UqMUcv/9qlE9
BZmUQ4GTW3DJMfSjfVR6OFX0cEWmXSeDW75VbEvYli4m3m+TTlTZtObnolZ49ok12EPWqzJD1alM
EfF8O6i9lPrYZ5vOwIIGi8P6HEQFgjVR9pUvj6wyHCc3rQPKuVDCV/Ig5+jm6NpMOO1h2RkNqxwH
trgYBDpRWAl+by0GqVJMj5sszAOVh1KM3gmWOKE1ZFTmxdEkx60MH5nPW1saFRFXjNTuJXXdM9HK
gZxp5Jv+MQIwtz6pwiK/7vEyg7RP38tng3JFQzwjlNWHeEU5n1nFAth4ViGQ4b6bFYXkAwb89Hdh
r7uvmRYjl0Ok+t8XCOyGixjJtx/y1uez5LPBl6rTAcTRiNFjVJutLKm+QzDN5qh10Jr56LjI7b+p
9h48ZqrqZlOz9zK5P1kHTYN9Js1uFkSDnBrUd7Hv1zfXEtIXl8WDV337ZKhamNT+7kQCWqtru+ld
Iwp0epUMh5x3MreDDq5W0BGFapre/BTmmdLJoClVYgMI8ikfyT+f70p88ExRsd1ChQeXk2KraGNn
WO9i4LLP2KLLeSfZF0+ZFiInNrAvehibzAJjob1VJf82y+nid0AI4jjLOKx9sdGg5uhheu3ku34i
ujgotV8jO7zKD4bhKAnGMRlgWOc9pEOD8J4T43fgo9/yWqvxT7CRkQsH8o7IMnw0kASV4J5jyTK5
Q8D5va+LFmCzwK4eTEibefnzc3RI6Z6/G3jUt8QMIjg0vdcy3GSAiktthns2hGzb14WZoox1VG1K
xYO0N77RfSOrRMG18rye8I31IqWvWejkwDK8Ig5wDkvpEDVDvo+UjBTXDyq1bDbKctM3ufSb+IQg
im71xSYZ4bgl4edMw2jo8jqM8B5ziTCgTnyC8e7zVy8VhGwj6rJo5V3PRZi8GHEECk3/5R6gAwcy
Lu3An/l0ammB8TcHx6s7qM2p71nEXKBzyZNKsHzRMVd8/h1S9ChfzoY4tX5BMEIYkr0lAte+kbxw
y+nNoyOZUQ+Ro1VLfCHdhq9+wFv/y7vdSrBKuI1FvQ7CEtAYf20F1TjqvBByLLbgqimfNXeTQRIC
FDOmEr7gEPSSoCLyM/yenFPXXFMpgjpesLzBbNambiJ35VRsAd1SafzZf87yJjVR3xwwmNuEbHlh
Dw5Jn9+7Iv2O9pX1REbLpu5i0dunacIEC4i0GDtQIMiIZzujixNK60CneYINp9TvAOanXf69A35+
vAlrPEhQmIjHjhDIaDM4KN4vsU6wqtDKhYU9uE6SbcQfN8sSrcPgwKHRg4dycbrilsuju2spVbsD
22DhFGGHFo7FV2PCvx8FJfd0NGns59ZM0640DAAAxvRsNLo4PGrdLGxKmu/bwegTsWrckjkBA63F
2K6TAyKp8u6Nu4Elr7cWbGF280Y1M5AfcsY0sujyOHIrQqZpNDD7R2iYcAFvahXohSagq+u0A2Lk
/eLQPf8i/AcVx/ADtaDnK2qzqth7Na+TV75oKsVTH9piAC3HBgoUdrUDv3QREcR/aGZ1TLcMKwt0
ForbNS0RKpWE6RlWThgLwrqSBLK+28GACB3Ppt0mJofy61Kkyey9osuAvdMG3sZ62tT7q2hpBqd5
vlp7oCKE7nShCZXtN4K3ImWUMlZV+6hHDukukMYUWS73auFVnE3k8HvAUqpAXXh8rFCCSHL38Oor
5uwWGHXFQtLbeA2QQtHDbSo0kDnrQO63PiD4Vm60owRIDkeP/Bq/EWVak36NLUpy98LHtoTEAWXN
q3iOGjWmpSai4rET+KZajRuti5Q8C3/BmMJuhFmfAeS373R/36eVAkO6bfz7cv3c8K/29m5rMJYw
VctRen6t5WAxqLNDN2NdJcdRYlC6ZrUxP/VHDp+FN3V4YhqcxDiM5RSIp0Cuy50AFdy8F6yZWWrn
CSvkKQVMEBClsefowY9+wbZsNa6Qo035iNhfG2qR/RUgFSJlwboIcfrMGrnBd2SGwX59nnymMore
magMGAvcVhyWOrq3pf6q1wZ93OJ/y+sO3pqVRUxNL6dwLUhRKh1g8p8KJuM2vcVOaKLJOrQB9iGi
+/vT+jIHWXBDHeKHZ8YW6tRJLrtHRKDS9DBD3B9oVFtf43lFoz5Guvyu6OMMiODe6sJRZ9/HKfds
XUbJTy1YXwlEGNDahY+nsq0h9sAYCZe9G7RLZr+E3GktNV0vgvkP7tkq4dF8QDDSf0r51TTTfO/X
D8QRfUCGoOsvQ4C35cDXjoh5BNDRZ66y1Z6W7v/beRODCMHb7NjYCl9etx2JGGd56hMlwIXok+gc
Fio7akxGcfEshlxkVgt+fgF8JUuZ5ZESUFJHs/XdljhSuV4c5UJ2CEw3xFsewbhRDTaOhePqKAAk
WZutwJ3WwbHFlAPzIgHK08QjhnWmZns326E3EKUxzUK+ed4YrUsinRG5cgNigphT2D1LVlfPTYuL
Y64TV83wd/PMcId74K/yBPijDzVjCKpJsxtjnLGaMA/pbD8rCEX8cdExwS1E/4KRt+6a/HNmHXSQ
UC+7yMi7rEw2O4H9Eud2l9I4GudSVWSzGOrUu1PI9zLTf+/NNsGiyX6A9RFFONWk6DZFNv/W3rZP
G5zozAD8cHuN99RB5VPBcMZNXIXc+czQxCRz0gwkdlvEPF0Ii8jZHUvmxrsUPnd/iq6gx4rbDTnR
oPUh2IvDyS5ar+gxsEGGbEpZ0lSu9rdxxmdNhBmvkDYoalGqhBPpylckhI+qOiPvrKi9uMMUC5fA
NRr2e11iW7kMlgTZMhgV2TGyJrJuWFkrahckwaOT17mx0cMUqtWSGwHXgZDUpf0a7rwySfGIMaaa
fjKDrHyrrle+tNF2Fnx7hLN4myPE3br6fJs5vnreLU44vmlyZ64LizO4PzQbGB4cOnPTM8gcTaiY
P7ZuS9H8Q63uCA8XQcwve97ec1fmfIg4KrYyH5kzs3Lk+4SZjxS4E5gC41mEiBdi9BW7d6mBzh7j
piMsjlYZpus8g0DaY668Zcx4fthdWE7uB/p7oiFSCZt0E5NCGUqAfc46EaaHj9w3x/50Bw1KtJs+
AtXlPoLBdRs+M0GJAqWVhGJj4zj80/uKiv86fUzepZlbY6rFps/qcu5fz8tfhAfQwSGMeyD3DW3p
lIZ5dB6KTgG/vR3mejBD9E1TD4z59rJD68Td4btuFRCHYpukkbRiTfzsxqIu0GmK4jHEnnVMy2dZ
9/XLbutifrGXvnnIywbzqRxt1MRvvgXjKfDPf6hJSam+0cL+lGuBcV5Upx3LjHuAXHI0zmvyCwoo
M1NSDLR4kc73Bu3HkCFdtakTAi426DSaHPed4E1YNcOlJ+0f3Pl48fQircpOxPxlhENvgmptsrfB
nEneQsxJ/wd355U+7xIz9st3Eftqjl73WYpOkIv88AytMtt45RGITEavd/V0H26L/vvsB7iq58y1
nD+4v9HqYkJeHn24G29Zg264iuEiew1HrM57IoJdqsZfkDmG5kWGPE+EEwQjJCAdMzhjMQPiJgtc
ISj4XX+NqeZUBAnAvg+qpmN8qZifzjmtf+l1O7vsIylL
`protect end_protected
