��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-�  �n2ҧJ����TZ���o{��-���	��wKm\������K]-��7�ŗ��q�	�q���r{����T�
Kf�ˠg,.���g/�z�Б�!f�Z!��ی�D��h._�t.��<m�ryN�� Mڔ����߁{-i0tV�~6�D��u�7 ����4qeJ��/�ʋ1�����W��y�k���l�/����
��.b��Ky�~�r�w޵�)Mf�
�ţ�^�p�܈�>��*����8 ��S���ۙ��f�{���?#�� ��0K#t,�-|���&<gL�#n�ua��פS�:P~��p�g� ��~���'�@���#�Y�/'i+�z�dk���W��AX��;j�b�^�%]E��\Gq5J�O�'r��H&��C���S�F��"�J2tcLq>l��P��`�I�=�4�c���&�És����7�?m��X��B���;+�v�y|.Sx�^�D0��7�3A{F��V5u�\T\:��e-d�Ӳ�<��	�T�En�TR��hs�fC����A�L����J�ภ�2��.���MW��L*mmݪP�%�{�>[@퓷��|��͓"k7!}BIl�C�{R>�}���I=om7.T���n��2A��=��99�5���L0Р{��;�Lh7�w.f��a�v��������������$��$��k8겆oU,�SI;�|���i���o�wkQ�|�])h��uvC�~�߇Ι'��F8g��SL�����):u�U�S��;$�
�Y}�t�#og���������On���u����ݺG�a2o�u8�6di����ސմ'ӄ$Rx�y�<��wA�*;�x���@�̦�W�X�fa�M-$u����n~�%���P�$��W��kYَ���P7�?UMfT��q�6�U��k�>����~�\N�(�����X�e���/6U|)�X2pF�]$h���d.���9E��WG��L�X"]�Ad����ľS���8od����e�GT?y	7�������ݵ�^��R�q^]�鍦�����s�ae���h��L��P_���ާ��YЭF���'\��68�b�[����w8�[X��V�F�0͘3����q諵�uW� �h�u\V�?@��_6G�_�*�G���B�絉�f������[�G��U&�����~�F��AׯK1�`c��[<��FY���4I� �#�G��x[X�=�Q1��`��R>(�w����R�O�?����7�,(�H\�#h(W�EH=�������yq��Ѿ��aF����:�U~m<|��.��0=�P/���4ǆ���T(��������0Z�"�2���j��˹{6� ��/�t5Q�؝է⌋�o�A	@����y��VE�7(�W��4�T�Y�{��Z��j�z��h�9%�d�@7!���"��|��~�@&��$D�☖w��3B@'�cu��;��M��%˄��?�5��:�|4V]ꊿFbQ&������V�I[�Z�O�@e	3�������YA�QPΠ��ͱ��~�h�/X����r���i]�E�/��¸lRU������ʗc�!��>(f/�n��F�s5; �!�+�T�#�7��h���"ݟ�!t��l�ſ�41�s�l��&~����a}�em;[���	��Lf$���\�,%��}c���.;2d��kH�%��ޛ�\�
8�T����>Gg�d�!<=͆���90��hZ�1���������4Aփ����p
�^�M&-�FP���
��Q����6W����Mh����I�v�w��d:�d=Ю)�4ٓ��0)��I�
#�ٗ�s@�W�-���#m8�5����=M����|fy��5r�t��0�N��d�B�IQo)�_oE�;�����}�Z�k6�O[�m�Ar�+�=���Lm_R��k˳\4R����:2&1��?�9Re(@У�z%쾿=�.�iZ5#p�q�P�k�?2���e`6y������&&����mM�ִ�,E�*�ښ;�Ȱ��i�#@x
^�����f@�K��ɁR@�fq��_P�<������[�+�6���>�^��CV����J���=xF��%�;ݛ<��Tx���T�C];''P���Y�8(wc�JD��Kw��G�Y��?G�M3�n-w��b�C���_bU
���K!8�K!��]T�)�G�6u��Ž��ծ꺕��̥�a�},�:���צ.�>��IT�s�i.D�@��n��i��K�mL����h�3�����|���o8�-���Z����[���@j_RA=	�����im����K�:�ǂ����>��{��݌�T�\��E̩�~^���T�?ۥ�|����Z�I|D��(s4T�����A�km��m��)��ȓ�՚��X{7��6�<��JB��dyT�z�ֆ����_c��wf�E���8b�2;���k�Oe��zހǏe�bf?PAf�H�)�o�7�+���p'�[\r���Fl��,�n�%�Đ�c��4�i)�M1�g��R�L_r�5V_-<�ў��lHI�>&#����|
�DG�˨�Tv��.<�{��aU�!5	�#���}��y��ǧ$���E��/�aXP�9�D�vr��ps����%^�ı%\pn��0,��5q�ʭ�r�}�b;682ן>6�2o[�����i��Ȩ�[�C̉W�5�-R�攦�g��)�t"��G�gY�#�X�|�r<QxK�/�� қl�䮬-�(�;��F^�|�h�JzA����CHB�����b�B��P7�2!rw[kױ,��R]u���/�����)TУ:��-�B�"i�7��Q�D�8�w���%֤��5d�hW;��_ub��|�Q���ͪm�� �=&y}��;��������Lu��F멮�U��c����!�sĿ��֣�w�:Ժ�|�7�tNA���:�-���c�����ǰ4M��@6*���;�rk����^q��2��a�9��<#ǯ���R�3U9 �h$���z�ߟ�sG,(���F�achF������[���!��cU�"�C�Q�x�{ͳ���	�1bd8ݰ8[�!u$g]c�C�ٝdU\]o-X��-'�kTףw6S��p_�Y�}����@��b�q�`6z�?����6KZ��E�d�� �4� sTK:��)���mL���2���_H=�39��򘽾ҨFD����*R��%6-��x�*���W.���@��Ƞ�]�mz[���s��Y��e���G[�6WLYn�i��1b�V�1�S�%�.=�BA���q��甃��v3�(�a�R�f'��m���w�����5����qSʠs�´3���]�ʫ	 ����.����P�D�Q^�Fp�+�d!Z"�}��&�k��5�@����6�.�8��T� �1���j4WMB�{>\���"���z���LJ�REgX�P���}�x�7p��n*R'=��/��;y���+��������#Z׃V
�8Ba�U:�����]�g�5o6�'��j'��f46��
ԛ_vK��d����"��v��Gz9��Pg>$��w�o8�:���+/&#��gX�����=ߗ�V����Z޼w䃛F�s�l��@��}�Cnۧ�s�#B�p�<xA�����z��!__��X{�m^�g�o�����CH������\���>?Xƛ�~-��8V��gZ˝���.�:e��L��<v����@�IRu��I�.é�ʊ!#�8w�&B�S*ԟ�ε2�XF1�є���rt���)�m�C�*�"9�Q�V�7���ۛ\6�<�s���p�{�{��s�H_B�����VY��ّ����+�4�[�0�g�f�٫6��n�g'�ux�x��S�9<y�I���JE�nt?�f�#�%i���S�T�|z�A���%��<W���&2ҫb�Y��j�d�M���_�?�����Qm�*`��)��[G� ��]��(�Oָ�@���U��C#�,M��B���uM�4�����Ԣ{u��^�?]A�{~[)7t��ވ6p��~}�}#)��'�T �*�j-45�����Q��K�3Y���w�@��5�܍��E���Ͻ����j�AB���C�B��V�} -��|�\"11 �rM�ZD6��%�L"r��t>�A��*o�oР��6��S��3�4���Xe8���N���{����m�)х�g�?�3��a�O�əm�� `gR�_����=��SԑQksn�kUJ���b����}ѽ�/�ۓw�p���(lk�*��E�U��,w�TZ���T4C���wTV��׀ӎ�.�db8�KS�v�ܢ	[�m����7`8�]�R�������
7N����:���:�7@0�#(�� ,����: :��.N��-X��P�c�ՆlS"����[����� �N���p	�R�ޙ����&|����T�-�կsB����|���O�B�k���q鏊svcP�ɘS�X�P:�g
Uz	���w�K� ����>%���0��������IN3S"!*�I�Kg�����&[�<�^C�#�Cc:.z4�`f���iB z�[$v��-R�����Y�p�b�GB��]�����溇�K@*�o"���d�Ǌ+�q�/�p9����U�t?�k$�hbk����9��Aw�9����r���~B��?1.� �V]U������7��@A�\�h&+g��R��߰RC���R[ܭh�ɣ���9�(ԼO�΄�	ȏ6�ȱ��'�̾q�d8��1��v~۹,�9{�h���b�8�Yna��=���'U�v�� ���~ɠz녹���
����Ul��ܡ���������)�{g��1�۞�W����C/�(����x���0�J�"Vq����D��j�r���-X���T�}���=3���A<�����\
?�h�QSZ�x�ppuY����F2�m� ����@��u�l�gt�I�{j'R�d��>������%@: IjK�С�>氳�s�g�7�����[�5쭼U���N6�',3ZMG,z	��s���'_��������L�`�5�ry�WRT�q	a[g܍س�/\%kn� è���u�ݠ*���%���_BΔ���������=�g��w�,y>�vū
�����n��sJA�5�<,s�yH�O��0�Jfs5�Ď����$1B���g��A=YoQEQ�V��R�F��t`ti]���6��m�_bF�
�@%���� �44��~N����iO��Aׁ�2�R��}�dy_y+���	\�R����K(y�ud3�K�9�3�?���n�<��ˇR1ђ��	O�E&��*�wJ��mF�Y6^����w�$�E�p��M���ٛq����!�!�R��¬�~�t-�"��+�
�n�ϣ��v���O�\�����+�A��,��mv��Z��eG_�UE>�w{*`�s�L<�h�Q���n�)e���i�9'�^uR�Aj%��������	&>E�g��&��Ň��*!ۡ)�XX 9�^���kK���T�嗥p-�L�H��D��=�P�~v��×ؘ��uK�\E��%�X�8?`�tf��1��,q��Ǜ�7^R���[JT��B�_��P�W&6!a�:�>������+�2;�vVM$���+�Jmw�04��,P�
�XY=���
�N��2u���k�i���3�E&c�]�WPPǿ|��C�t�L��FY&x�,�Z�Qp��J�8�_��;��!�'I#q�O����q���G[_��U���z�z�ΐ��h��#���RvS?��&�|�Ғ���?v�Bw<����ʾ�!+D�,	i���o8�z	��=�F�G�g���A�M
E��g���$],��Q���Q�xV�/��qW��f�r���a_<5� {�W��x���< ���䗥������/3�/%~�)o����Ud��;3��8p�2��4<U��9�}��P�Nǝ7�-x���^;_"3��7�Cτ�e���>���oM�̫Ȝ$��2�f�������WWf�C0����~�ի�YU<OF�%�ݿ�uszQ�m��ڊc��by*��#�A͆��1����{MbDM�L �!F�D�k���\9�UB�rZnm;JP�����ބ��-v�����0���Y���5�)�v�t �E�<�W�z8�� �Sqeou�Ac���`�B�=�_�C5G�B]�_q���y�@�d���Y����l�GD2{�}����aNȖ�y������F3$�Rė^�~
L�==�I���q���"/�JO�M��$è�rڊ�Ӟ�!��<�����Io{9��!� .�3J��b��M�j�5����vy��p+uk�Q� R�"�-���R>Z�i��֓�Z�R1�3L_�t�3���E5G��N'���`��8�~�Y�ϻ2��.��^�B�������=S�:#��[cd��|z:�![��_�O��4�|�!��H;��g��n^t/�]>�*�V�jCD��q��*M����_��^�9����4����nC4��&dVI6�*\�w��m���+���a�O+�{�whr���Ȁh����ă��9��V����I!���F.�_zdaP��5O�K��b�	Q [^�#���Dیq��r�(���)ӗB3.W9��Z�G�tl�D��lf�7�O�)�J�s��U+���hc���`1!�{rg�8���5��ug����R��������ݘ#��Y�)�����B}�
�D
 ��ȭyк �pkȈ��G3�P�vZ�mm���׆���mW����)-� l��p�(vk�W��ж�㰾�m����'K,Y=J�b�
.��V��9p׃%��)��ݐ��%���9������w�ޛ0Pa<F>��F/����������Q0��_��>�5��4vB�������l[ 3��Cx	36u�z� �[�Y������%�pM�T�]e�9>����avi���Cl4��3�AnD�fOX���r,�F�!�\���S�E���1�g�4�ؕU�y�O��1�����X�ߖ�핐����/��Nj˪D��:w���ZniOgv2iޡQ�֣v�S�0N���lO��f�s�HR�����h��FQ^��.+��O��,�B���D��ļ��30�q��ۜln���Yj���e¡*�Pd6j�����oƩ���Bq���L��UAK�-v09�Xp��v���C/N����Y�,?�xr��k�j��BM=%���c�~��к]~2ѫf��ސm�	����e�R �&
Q�}U{ �GZo�S��+]�./ZqU+�r���V�$���h�Z���4%1��M��j؛ڛ��>U9�ꖓ���2PU7�F��y�)��%� ��T�P6ӛ���-R0�*���h�����HC�g2��\ɋ
�w)�ZB
���ɟ�U�!�t7�I<�`�����>kJ ���ٔ�b��.N��C��o��qO�bd;Ⓚ)��qc�@w`ll��Z�f�I�;���S��ǌ��g�9�jﱇ�C��3�ԫ+e �yM2��'z�.�}�1t$�l&�d�)l�TB��i�z��5Z��K)ۻQBtq���P�8�Ofc�����R�G\M���^�P�S�&(ᴬ�S�t�ԍs�b��J�hl>ubadg<:*T�1��{g)Cs�ݶ盀+�@W.���x��i�fcC�.߫����z�ad�뜯q�1��f�aFR��W�DBhm$w�4� M(�Ofg%��m�Mm���D��Eh¾�4�yeI�k��B�0"���5Eq�R��O��#CX�D<`��CL�%�;�e~����v��G|�R�AzxqňZ�;���32_��-[|����;���(�aY�"f�y_��/X͚�v�ݒ;~3ǝ ��L]�F�Y��n��p��}�yH��_�A1�af,�W��3cxԿI����ӛ4�b���Ł���M_�~�h �2A��hZ4����G�b��q�|i�^"N����pu��ra��>���e3�	�f�L>��G�j�T�8�%I�S`���O?�h_���o5�o�%1z����
ݔT5���pN�ϓ���Q���ݼ��|	�=Z�Ϸ�Di�c�?���9>�g����xMs\Oee�8�յ.-���O�j�L@%~P,F��`���:$���ǻ��|gg����G�L��B�2��H�?�x�.)�.hb_i<�6K=2�����z0�����0	j��l~c�܋r/��W[� L�q�M�W�>H�`��n|W��r�Q0�p�?��ӊbTj����Bp'�oF�&u��j BMY9�z޷�3�}��g�n"��T6�]'��qwr��^�	ߏ�I;���e0'�X5�ɯjK�C��J|6�f4%۱A(�#k.K�)�z떕��N	��W�WW�>���
��4��=|㗯�;�M-<mM,f{ ll:*;�^X�;t�v���~�8�|kz(tm��n�S���D]���z����ɝJy���J-4�tLu�*-MY�KE��荧�^�Ft0�˂���%����-�����p�7��[��3ӟ�d������&Y8͇1D�"�vty�V�\|)�ˊ��W��x��ax�b�ظ�l~�@ƦU1:��N�������![^p�Ce^�}B��t����51=�J�~"Zu/��*���L!���me�e���ҽ�fv�V�!�*Fq`�aF�T�������q�8�m��0���"�mB�%�f��\G��2c��t|�e�v�,F���:0(��"]�x��k�l��T�O�a���H ѱ˸��uV_�f��B�TJU*�x�MPhwP&�x�k"�����׮9���˱h$mk���)�h������;0+7W:�#K�u���5h�ŏ�l����

���t3*����2�QvC1��eWZn���[&*���arr������f��u�HJImа�걪�_�)�<��#�k@1��ѩ D� �4�%�O򮏼�3�� a7!�v�e�QG�"*a�rB��:�'� �����0m$�d��u��'B��ʟV�k�Vi��j/#'�l��ܭCq���l���"��ښ����J #j5���Rױ�{��3��iuP��2�!c�*A�����H�V��3�#�����؁ Q�T6�OE���`\�B�� ��}�B�w��0��?\��9��Ԓ�i�T��K�G��u����M;}ߺ�E���dp�Q�c��{=z�q踟�`=r�V�!���z0���͘ߨ���ё^�J7(�"�gug)Nm��	��W��u"�.(�tG� �ʹ9��YN�1xi�45}gFX0���������f�>�����"���s�U��+It>o]OT>SO�4�`eݮ�ѿJ"(!E�������8��g9��^1l�6�k^c����9=e6��|�Lw �M�����'ǂ('������m�S��œo�Ļj����J�Zk�֜��"۪z�6�RJ���r;���ٝ��l��f]%�݇�R&T���n-FB$S�ڐv�GT�kY��ҭ51��
�>�+�p�a��Yd@BYFԳ�[�ᵗ�c��ߡ4�V1���kO43���6���%l�Cw1Id_P9<�����Z�q�ZE��Ȝ��NVFA������N���1f�n�6�/���D)6�~�	�q�ǀ��n�ӖtBU�����n��o��L�Ս�H�I<�<��PIGjT�*4攑�pW�dz�]dM�<�U�ü6�1���������Y�0�b5	MKdp�n`aL��F AӳB��G�D%�iy�u�U5�CI\�Q��a)(q��KR$~
T��"�ez�ia0��H%B<���}Pn�=n������D}g�s���TD#��W�9+x\�b���X�!����jS�N�K��m�l��g��=�W��nY�$�����'�aI�B*�&�E�ĝ<\S�E��"X��Z��bUQ�����_[G��m@�a'�O���+����1�O��-�J���Yhyi��o�u������>����0(��7�*�X�a��R��!p1戕�k	��.Ci� \�3���;7z]���c,a
>���þ�2<�Kv8�5�51��h���8�Y_|�B���L��<�FL�㔝������?2�&��$���+H)}"bͱ�vXa��S[R�~�G:�0x���X�m8�#V]�lݿK+��HXG�G����x�]����
)��<�}���,zp����V˾�~Y�5��j�=(v&����vGZ��ڵ�M���𰪒Ke���:�$�2����5�6V��G_�kluC9�4�@}��_���H��>������9�yM�jߞ�'3�E��0�w%Aa�fk��r�Bq�є��v0:�Ӛ}"��#`��Y17�H��T|�9�,rD�yA3��:�YG�"�hkH��S�� .^<d��[~<�z���-;N�$�2+�_�P���)��"�+��3�L���.0�غ��!Oy���^��,gzX$���P�)	�7{�|�Ql@%���O����X��T�@^��( �܈5ǭY��2��v�P�iCRc�$*U�;�X>+t?"{���."Kƶ�:z�sV����a�;�<P���5�lH#���u�����0�!�ǜ��ȧ�]�9��!E�l��,G�����*Rf�S�������q�㶫ղy
�,$	�R$&���S¤�V���H/���E��4�C�[�a�4�#�ݑ�2����Ӂ��R{�����b��c ���E�7��5�
�v@�}nW2%��%�A�l/?f�ǹ�v?����@�f�"�[�gHΗs(�H�����U�Ё�!�^��`����g�7��H��H�qeh8����Ì� (ʺ�U]�pe���O���)�`J�%�������w��G�Q��'|�
�}sз�)+��!�(+��9y���L�~��X������妣DyE�wb��zMbEF����'
>kF1�<ګR]��usQq[2QF*>��!rvw�����tɎfd챨{�}�ԑ/�޵� d���ȱo
~�Z������ �.*�t	�V���r<�C4��!{�b�|�1Q�~��|��͡F��8�i��M����l�A�q��iN��T�4K�Gö�\�H��<�Io�W]���`T}�d���!^ �$���Xsp@s�6q���L��Mt6�z�Ez(+����E��C��Bwq	�U��~c�f4o]�f����x>�Y���k��m$]��1�,<!m������W�������dQ)��C>F�[u�?��;�u3�>�0�8���L=ǁѸ���35?6�I����׻*[�^G�{��uĴt�����~^�S�߮vk�p(�Lo����W<��+A�����d��W"+��- w�QފH���� og<�A)_�L�]���\���'1����)�Ϸ��ؑ���}����g*N����j1fH��c��������"�+�I9�ԅj�I��b�C�Ǧ�B���݁�`��@Y��ǃ���<�Jg�+	�i�hܖ�4�Ar�V�ڠ+��O���Ť��.׀x�\#G̵Ơ�C�	'ҫb	��\c����z� �%��P��_��QaC�G��g�lV9�'����}���0Lſ�O���j�9�b�R�k+b��`J�x�R�#���hq�T7JS�e��.w/����Cƛ����R��1X��4�ZG�V%<CƊj��8{�Gˬ#���Θ�F���5��Í"�A��l�e��e$��E�T�Af$�{F�<�I�Cq�2��v� ,��,i-��Ao��nX&Vl7bz�ˈm��FSɯ�b�Kh
��=vA�Nܸ����Eu�^A����1�)�ֈ�`'�O�x��ܽ4y-n�xB>���C^X��Z��$=�x���Z�ϳi�������s�������E�z0�p,ڜ�*Pt��nWë\��O�)�S��ΜR�gk�@=D� �m�%�$��w=��H����S��K��)E0�!D͌��5�8�lkn~��g��Q$uLg�qM',�Q����L��(	��f��^��H�����A�>X�f]b�v��������7И���&2A�̈́1��Y��Oҕ���d�iv;��;,�ӶR��:�6�F0إ��b��y2�\��!I�j�/x,��Q�R�e�.�8��!f,R��--@D	)��;ͺtX�s�K��s��תpD��@飤gc�-�{��j x_ۑ�m�m��왩SI��m}I���}�0�ssW��?X�ojs��j��-W�R��;�'�zġ*���h_ �D�N�>�m��l:���;�.�' <]W\��rw;D�4���&����y#�������v�-[��SbO�h��7�k�W����&]7S��U6Q�$3?!H�]�C��G,�F����f1J��C�pvh���{hú_Xt��e�ܠWf��B�'�]UzL	�Ҋ��(݇�f����j+�dG*���/o����&m��@��c���T���)%qII���}�n:�p����eŖ%3ұ�8D��"J�8=�5ݸ\�^T
TW���]��4'?��Я��2}����x��r�ƤJ;_�?ǁ�$�Y�R������ǖ�z.7A��`��q��D���M�#�L�!"Ed)$rʟD���� �1M%$	�"�u���ަ���s��m�EUS�S�I�+�-��܀LS=�`�]��-ɭ�͉��'7J�nk����Jң����,D��Ao�oe��[R��	Y���ڥ�h��a}c_U"����1�}|	���K�<�B��^��3��V/�),/���_�̱EG7��o��p؉&e�O���1#?��"��jY����Ke�EtY��ҌM��cr��;*�T���@�`�ӡ��ۢY�I�d�R���7p�2ڀ1	X]��=q�&���*�;ޖ�mV]��o�IPĦ0$��If����t��L�΅9� �6s���o�hq+�!�i '٬����%�U���y�[kN�|�����C�!�*�!f��F.ZhMj���x�ak��G����ؼ$�-O��馀�כ*e3��Q&���RֻH��d�w;�%ˣ9)���$�h`G�D�d~�|HL٤��`"P��Ų\����e}x��0�nW�Tn�d�ց}�V
�g1�e�7�U׹l5H�/6�n���L��grņ=��Eo��s�S� �c�]�/-Ѡc顄����.}���J����(#)��A\�S2B�*U��\�Wnt�Gz� -.���ԃ��ޱ#R4��r�1��*Z� ��E�y��ΔW{RG�R��8�c���
>�?�z�b�m~_�j��#�"���C�4��C��7�wH,�5v/)�}�*]`��P3��qB�8��(b�5�^#�x��	o�Ы6ìP�J���0�XT��]����P�F7��NH�hǘ��Mo*q~����W�Ί	��ѩ0-"l�ټ1���)k��>���}����ش>����PE�
(o��U{X�P�m��3Վy��
���C42�����9f�e0s=�,��s��MN	[K̕��y꛸NH�[�=E�����w��X����uO�r7%��@U[>�Q���.��ߴW����<Uv�,:?8��ƆT�gCXˊz�e� �avV4vFB�|�����.?�D��Q�N��=O��f���H6ǿpt#(ɾ��H��3E�r~ �U�K�[ˀn+�	m�v�p~j�ꑤ���U��W&٘��S#��7-*�ⅼ��Don��~��]���
M���d+^�t��{G��H��V�,|�>`���̽��>�?����d��� � �% �1�:XC	�>��,_�k65�B��mT�03�.�4(�)'Q�EkR"0�J$����$MVx�4Y�.�t�@v�ڔ���r<�.���������Y�oB���ȉ�r��2���f���fP٪VΉ���Oh�y��r�ʢ��^��6	��MF[Ȯ|Ae�5�N�>Z�K`@qkA�<��3������M9��f�Sk������</eUd2��� �k-��#�=�' m*���)�o��nu�޹�=�g�����E�
����Yot�yX�n�^�0��H�����Y��Ҙ�8龜2��M,-/1y��-C5���W���n�~�Z�\Z��M��X]C#r �NG��8�xġ?��X�ǋwߢp�-�u gR���:O���J&�W�Q��f�ȤA�\�P>K&�=��p�+��8\�MwQ��Q@X>=ǁ���'MVAlu�;@#�#f�(��F:?�uV�g�ϕ/��0*B�n�a�����|"hˍ�uC�M�.<P���rQ׭�="����=����@���bz+�e$�t�˿J꣺QF�D���;��.���j������m^>@�;^I�vӐ{�ӗ;�~��*̘�y�m��L����lU�.ŋ��ѝy��Nځ�w�c�@s�y�z|R�r��%��o�)1� ���{�!9k��lj�$�:�sf���������s3C��-�,�w!�P��3�"��]��Y[�:KK/���R�Y[�ώ�����z�+BǾ��XqJΠb�g��͘b_�5���6��>���N�nF�GpY��2+���;N"�l����|�TeH���v�5�d9����_����o�V-����CI,}�M���kln�.3���Z�B�ޛ^��9�|�b�4��#)���.}�q׈���r�n��n�]9�15��ޫ��F�X؉@�H������B��G�.]�l�޾��3����֍i�a�����t,��m���SJ��(9��pzh���Ξg��i��yb!�a�t�f��`$5��vt�6<�*ԑ�W�^� `a��h�E�C7KX.�GG��� ��z�N�l]��D��wߜ��	��*��B��k�ݮMU	f�W�cA$i�.��D(r�8��_�"P��~��Jx���lnki˲U�.\x9��Y�Y^9�"<�N��.��TÌ�[#�(�$4����-ܴǜ�m�ت<L�3Z�8:1�6V�� ڝ1��7��O@����^W�k9I__��e�5w��;Bx�|8���{��mO���a�����%�`}��X_�w���c��\�w�cf�����V������t�뒰y�aIV�	��3��ܬqx��0Z'w1-�G�������	p@��;�y=ב��49�لX��aH�态&�ԏǈ�Ť�325\6���HU�y��b�+j'�"��~Z�0��	�f�+}�-��}#ŧ�gz��_d�**���V�e�1��\4G�@TERbLԂ��.~G�͢�5�=�wv$�$w:�v����vi�ļX��v��o����nWCBF�[�u;�_|I'_��s�L+o�tD�V�� i�H��Κּү��MP��d@x�Q�P6��˛B�X61,��)�j�t4�?���dc��}�O�ׇ>��}�*���t��u�b:�=����x3bo~q)O��������bA0!�0���7���P�D���ڞ*�@C.��-��C�������	�����V�V�)1H�`ﴸ��K�7V5}�ƴ3�m����O�Q��3e�s�;���y�-49�<V�ֿ�8l�X��A<GC-�ؾ��>�_)���������p~� ��1_� ��7ǋ��3dn�쾅�,�#�i�\w-�J�I�Ne�? �h�A(�`v@D�/tp�:��V:+�u�S� T+jk���p��@&r����m���@
��7B�ߜ�[[kOMՎ����3�G��W�I�N�ئ�Us� ��;/�D�M9rou��4���`xn�wv��ɽf����Ǐ�t���	)��v�]e=�E��!����6� 7�Ia[u�N_ !�i���t�,P��7�a���,k� �=Bf]�g�����[xR����8G�"y
�CE�[��-X3Δ�.	e�he��1��e`Qu<�R[�m�~|nu�Iz<����PS��I<glR�G��q�"6ko�|�g�A{F�Z��g�F��q�lhLˁ!\�l��Qr�l��R��`B��c�}TR~��X"o*n��L'�B��5�L�V�k����e�n��9^�x嵀(P��`[?�o�v���a��[�4��`������pg)��;
�$��cύ2����UMk"���1�ʦ�����_��ݿp1�N�	Q-
%U���PZ:����P;	ĺs�s5÷kɰ����bR��tq��Z��}�� ��H����h*	�J3+�5�w^��<-N�Q�!�ѝ`@��rPrߢ媺,�"��m�����m�g�׶`�k#�ɺp���V}��і[H���?�T�<�s�/�}�u9j�q3�Ġ��|�4ƿځ�y+[��<��_x`�+�ru��YPj�*�B9������#��q�f?��_�	�����m��ڭ̠�U�+��!�2��jɾ�f���S�(IZ�������3�#�i�{��g�s��Sc����#B��	RE��,F,H��cR�X�V�d���^��;�BgXP�ڼ���y�O�?Bz ��s<�F�5�/����L��)W��!ُb����a��-7U��S`%-���U�RR�ʞA��Y���su�@���}�T5+1����yv-��Ja�%*Z�T�7�
�U�R��h���lsV�k$u������<<�>(uUܐ������ԇ�P�\d?�H�z��� C5�jW�����'p�?ܲ����*C]k������!�������yK5.����7����h�o[��-8l7���OүW:�(fy\�l�Nm�7��;�h��M�;���@�~gi�� �Zpls_/8�`D@Ѐ;Jk������]��i�0C(k?M5�������2i�1�gw
���F_����F�3�ި(t��j���g���\�K�0�D��u�f������ �U�����]�L�?�Y�Q�<e�_b�����TsDx\0׭\����d�yg�h}���A��<��� �\�t��*� u�P��L�8b�/��[PL����vh.�xk~�!x�'a�FK:l�t���d�~'QI��s���	�uB�2�30�T�>�A������k3/���(�e7	`c\��3��(��H(�7[�Mϓ7<OK3�O2�7����[�u�ÌY;y��;��ܖ����%��ˎ���(�ս�N-y�4cݱ�d�`83~�ص�;�=�g�GlĵT�J�:g#e��':B�����&I̧Z�������)
������3����G�'�� 1$5C��qm�iwj������<�����7�
����X��
 *C<H�vgJ��g�ws��*Ȁx�MA����p��!���[�ddnS:
N��=Y<ˊ��OL�I}�7G�?��
�[.��xpz?c�S#���I�N�3�[�sB!��ѸbB��U� %��e�q�Oc]g���8�ǒ�e)>7g�Y��qI�O�	v����*��Z+9������ϊ;�	��#rO�5z �̚Cr�A����D��B�f,<o4�.�s�`��ۇE%ވ�5Z�bH�kӐt� L�k��%���
�b�{���'�mP��Н�-ߊ�~�fU(��!��LD�@_�k\`�fqd��E�2s(L-d�Q �x�̊��`����߿M�}���ܬVּ)�a�e�M�"9N��G=��bn����N�J8ӂ��׾2)CQW>;*�w,��[7�)�;F��oZ[P���~.-���f���#t�0WwMh� ����4V�,-<����-�-�_��_��w�(e.��r49�|y�Q)�d����n#�rs)��g�?�=�>��V��6��n���e*�m'#y��8��BF��Cn{�(���N����,s���8���1���hJ4��[24��aA���|��1�\�!!G����h�xPj�b7O��j��#. {�����x�E�;\mU�+Ԣ�����Q��������O���=�_c*2�4k�������e�:��{����H�h��~�U1|��n��+�Y���� r|����r�Q��&�A~���0�\Ќz�wd�@��{�i+�y�ɽG��j�7������ƈ�dt����aD٦��(
��(:}َ�o0N������ƪ2��5KM�ۂ<߶��ǩ���N�<�%�����Ab��4�[BժWG�>wҕLڮ!�����o�,ң��-��{
���]�z
o��0��q�OUp~�m_-��9��+�9>-������n=��s�n<3�c �;��E��u_&��5���apt��9ziK
�}�<��AV�L8랑��0&w�J���h��n�HH�J-�Go0s�#�~���9��7��sl{��eAO~w_�O����� 	��c�u�dC�|,���xB�����TJ�̀����N󫒢��-|� 6���>�p� �U��q~�5½&����|N���'bdMz�6r�w�=�� ����?fu�)�!veQ+��C%�������X,&����@9����j	$~����Ӊqֹ�fsM����d�*罜�*��np�j׮,3u��+�C]�^��(Wz���?e�l����Z��7e�}�� :��Bxӗ�Q��GHM���)��a7�ï����G�gוa��Py�bZ�v�8!�>D~}y��*�\4�FҤ��ղZP+���uw-���OeϩT)_>��xI�>��t~ފK�㔌�b�������i+�l���&�!��/q�� {G8��?J�ԔL�8�H���>=���:�1�&5D@��֡�*f��.,H�<	@D֮0MO�q������l�_�F�hǢI�%�Z��	0��\�k�>��E�]�@�ѣ����(KB�P��VԸ%�T�����1P�X�֟�'�GMԣ�v�\Tv?��G����m����^R� �LO�V���#{���Z�#H�cX��*Hi􎽲x'�T�H����W�q>:jK��̨�R9N��T��C���&��I��7L��Ё�����K��D�'�c��F0��W�w��e�\V�4>���;��Xd���b��1�ك�Qbd(o��U���1S���3�&}�#7u]�`+�b���i���TV��$����;�*�F�|�S��r��l�#���Ne��RR\h	!�� �Ȁ���p�x
/�H��p�~����s�)/[$q�i��Y�w3`T�����݋��,jm�o
4:@����^��w��i봿��t��%���>�Z�����a\�����2��
gdIL��Mf���83���ٺ&��u]|�S>��«N���;��OV��cMh=f�ܢՁ@`.�+�#������Q���Ǫ�	�����̼Þ�b��@~us�YÚ�^����/�p�����G�&����?�*$N�}����Y�{t��Z��!��a^�ࡓ0�>r�����5�i�u��^-ܕjE?B���mW��ܾ���f��"���(��B[0+������z���*�@��Nvx���ӿ�Vj�?NFz�=�D�W��!��rڜ���Ilp<�Ѡ�y�l	l�zĳ;C�!D>	�{�a���a�a��M��-s!�R�'��g+������y�ߛ��X4	3������Q�M@�
��?R09�N{m
�P�I��&c���)D���>->�s0��ē��§���(��I�J��^\}D�#a�w�!�'V�XtN�3�[(�FW�����"J\*���Q+��X=[H�đ*u,W	xM`���〔�(�bkQ�IK��5-%5T�_H��s��*���$� �0���ڃy��E�����ɕ���Ś?I�㶦�t����׏�X2��E��f��_UOX��GL����uR�'dD�C�< ����v���Xm�d�b�V�=N"hr����y �z�/0op�Lj�:�Lb�CY����P�h̉L��~�י�EnshpE��?Q��W�B���/xV��R���y��x�FC,�^@�B	���Ǚ�8lhL@�y
!���qE?��.�nZ!߄��*�p$�S͢���̈́|��-�C�k/n���6�A�t��j#"�j���5�M�w�u�y�����-�	��Q�䗁g����ϊ���:i��<�/ޗMc�a�D
䞛V�D�I6m�7�R+����k��P�C�����E�O/�I���]�zL�ٰ���%
%��SF&�Q�&Ѻ�|fՖ����d}Z%�A�� �Ҏ�bIx�p���������T�[�r��K[�lQ2�Iǁ���^����,�H[�	��*���?�o_�ܚ	9s�}I��%VՕ�ig�`��_�7�PB�i��2�7���<N5��������2�Ԡ�)�#贕�����\ƍ�P2՛�q�ԯ����U���2�ӝ+�������Y�/oz��WeyY��I �h�̫�Ar��+Jt�����j�'�'�5cݪ$�����@��k�UWE�,�DYf��w�'���p:ᩙt��1�j�NJ��Bx��5q��j�}����X�Ze5d��
\�5y^O��O�ؚ��m×e��I�*,u�>�U�����2ΛR�+r��$��%�����+���]�4a������v��0PD��$�aUDI�^Y�+�`�1�ZD�V.��LΐO�b_�)%���"M|P$O��5�ϰ�FtO�4�iSp���JՎ�
f�������)���IcXٱ���	_F��є�i�՜K"c
�'n���*���Q��=����z�_6��]lQozo"��w��ja�;8���8?�N��'��S�Q*����:�#gc�o�q����s��D2��_'��G���md)h�o�=����=��`�,|\(ؾ}˰:��T� ��E�����ng0�K�"�Kض�
�m"��i9��J{m�U�9Qj���q�HP�wQ�b,LI`��9l#���\ZI���$X��Zn|zͰ���d�R���V}<W�1=3lu:^ӣF���u���bIK�
�# Z]$�m��2�\O|+�	��E�����4����y��3�R�R�9���q~5>��v�ϡ3u�2���2N�=���-{��)bh"D���YHb�;K��Ä�;ݰ8���QiM� RI���csq��7�� oZ�_�`WH=�J��FD�ʓ�?:Z"H���	���w��?�Y2t�����i� �8��e�[� �t-��fB�#Cz�
���)�I�����i�=(�N6K�I�*�x4�����Ȣ?NT�ŇT������H�8�ݝ�Y�Lq���%s����7mZze���ؽ~��u��A���T�!��{*E�y�}��WD8y����i�}��&&������??Th�3{�Y�ǧ���H��y���"=��#��ƒS�oF���;��c�T7\�	��W!��q���T5�u(���2Uq�&�.ޙu���,1m�u`ys��M�U#k�c���"�u��*/�p������8����7U�4����^̦�/9�TYn=�.x�����n���QfT�ٓCG�>3�4%rʭ�U_���S^A���=�Byr5X)�/���-Z���~�����O��M������s�s���E֒z�>v�$l�sdqҿ���=���X�B�'���q������w�|~���Q�z �����'[��;*�GP)%� Y��N�7R�ez���O�ӶG�qA�Y�ݼ�gh���g$j}�����R(������h�:8j�����AY�´ ��L�ʺȮp��K$;�u��k���(s4�i4�`*�#	���4����|g����_OM�y�)i�M�y�B�	�aP*L�Gc��'A�}%�@�6`U���gnG�W��_�5U}�$L!�,�����!DE�5���|�XY���|@��f��{5D���`g�:yR^$����v�\if�u<W���q嗦��1� 	��vO���`�<$%_1{�:��>l��d�ȫ}�GS�� �x�����\�/����*\���Į$
4���suj��>+��[S�
)�1q�SbY'��o����k/%Q���)	Ŧ��M��PS��j6�u|Ȍ�lW�K����s��ݰ>#�Klh�	=�y#�|���HOZ�ÝJ|e_0E�
��s��z*;����$���Z?�1��G����id��D��Y��`������k�)�k�!��\p��6�����t�л��������;�w�fP�N9o
��D��*�ҧ�Ƅу)m��y�Vܮr�@E����p�D���J�$�p�/R��#�?���K^����P�mBZ{��׶X--6��XN7�f�Ų����o��o�����נ�"y��a���`/�P��!�W�
�;��Hv X�O�#��=Ok�7q������e{,�{Qf|��$�R�M�d��1]��8/��`�grȤ�!r[�ێ�"�B����3����<h����A^�_i �ԁV!҂����V�{ja(�l��V�^������F����4����?���������t/�[���,Xf����z��7�r�BN�k�m��e&ݜ>4=�ҽqԨ��i�"W���������*#�y �̃�t�g��j�mL�K�3/ۨd�m-���M[v~?b�z�Tp��X�ak�t�YS�S��1�qұ�'�Me���H@��?�]�9�T8�U���� T�S�0��-El��B4���M�<ؕ��u�
�k1������4�yz'*���%�pL(^[5��杙 BM;���H}4�lD;rJ2��#�T΅6����
�p�=�Op8�o���k"� ����as~��񕨚ב�6���S�&����M9�1zL��-�j,�}�:]� ��G�&8Ջ�S�`^���
$I���ʎ�@T�<3�$oDj�#�+$�ZR+����Y��mB�R�7�x3R�
+����*�'`� fT�nx�i])lk%H�������L�l�|���
�����T�D������h���A���#p��K�N���C��S~�0 x�.,>�%��f~���H�Jq2�s5U�_^���,������.���=7����͔��'����Pcn�B�X�#W@X�k��J*A�tb�x��v�g�BT|b��p�W�[���o;��
�l�O֒B&u��J�T�y�Y�.7�͗���_Z�,$Qb-������z2Uh���zj�}��Uk�w��4F��u�@/��<t2&=��}�iɓ{sIm)UX�#��R���Ҵ�����k�?R��G�8%DUͰi�R!�����k��X�_���)9�.��L��:�Tz�'�K.�2�"�zH�E(�A2K*��*z\��W?�����!��ʁ]�7#�>t�מ�Ш�'�8D�?�ίcM-Y���.9D<>��X61S��� �0��+����=�C^��\ɾ�h��R �U��!��,�("Is#�h�:d紻|9��m��To�2�]n��N��������Ⱦ,�G�<V ��/�/F}J+eP&Ƌ-F�)�΋
�=i�Âx�]9�G�~uA�@���e�(���D@��e�GQb������(q2G���B� ��:�O@A���/�zi�0c��.����$����������R���;V��Qs�/Oы��4hz.ES�w�EjE�C�#Z�..KN��WU�9���B߳��@٠��0�?��U0�8����Q�Ң:�F�}�;�0M%M%��P���x%����EF��A���X6p39�)��ݮ��s�RL6ů��ku�)#�Л��9>���0[�b	�2�lTH��N��0���Ò[{q�n���p��zA��9�J�Q���O�����������u�?���SL�NX�D���pv�a�e�~l���Z�L%A���4L�v;q/��w�T�ٍ��xT?�;���Z����e5�wኰK��b���Bn���s�sT�k�����G��bH�aK�{���f�F-�7a���hG5\��,%-SZ�'?H�6�vf;��1�:�����;��Ŭ����^+��џ����V�G�1��[�۵��&հ��|%�������Zŕ!1W��#�z�����{����Sp���:�Y����;D���y����F���wnI��$�"��JU���<xx�<��2u=u��r���}����:�4�ȲV�Z�Uw���r/�nq����YNJ��G:JZvm����wiYD��)S��5��¬����$�)WÉ��A��\oݠ[C��K�P��{@��^����Z%Ma'ɦgl;Y��i���
y1ǩXͮ���Q�M�]�i�O��`?>+�C��8)G���x���n82J��=��âo�VՔ@���^��]?$Ӈ��XGy�o�H�K��?�}�M���FB-*�����p��ͷEv)O/H�y(�2�$��Y�u^4a��Ct���9@��(��Gյ?�a��kO`�����3����:�u�����&%����iz� 0��	�O��+`�t��)l��E���kN꒞�g��8L��8uE���4N��q	Cv��0�C�X��M�s�fy��c�!|�;�9@��2����� e�>�ojIa+�\��4��'X����¹����rᇀ7��7��M@��moHÏJi���>+���[ԯ��
m���A�� ZG�N�Tb��c���|�
��s)h5�7ٲV:nQ�K��y>�qi�1�~e��2��m�)3{�� g����������w��z���?=ԏ��Jgӝ=�Br �	�AEAE5���9���y�P�ʢ1Y)��^iZ=���\v�|Z�/&�Z'o\s��TX|��>와�vb6ni����P~<�-���ᆅ|�S��m�����W@�,�}�&?gM+�~��]\�h6#�,�k`��{�����ݢ�:����mp�S���.~��:;Ӡ��_�y� ����y"����db���.á��@��^��|.-EnB�*=�3*��spJ������ŒS��ǩ;���������z�z���g��>-��zq��z��q����Z�F-��$�r�؏��?�B��=C��>���S̈:�@@p��@��?rٍ�lo�h˰�dN�8�����C|�mv�<�_�c!2{�?��?U�3�'��@gkږk��<?�!ӆǩ�^z	���g�.\�%ʹN�����_eb�H����2���n�(�,G`�QV[�Dޛ��Q��r9�&<�(yg����zCͶm��O_�4�N-�L��	�m�y�1w[A�Z�2�Cg�5�a�A	���l�={�=��8�Ǆ��b!C��;�oǫ8,�&j�͂<���5�忾������t��C��>-pe�V�jAT��B�����t�X�ͯ?�k�S�q�]u�^��:�p�.@@�eXb��l6>~Ѧ���j?K�Q��ǃ �:��|�Ò�6��P�������+�����8~����~en?uow�>y����t5��"�R�9[�Ӡ�|i��H�����6�$5�'��7tϘ��jOŗ�[$QI?�ϩ��34C�Bȟp��N���\CH:�`�M�pX�v������aJa��#�\���-_�|R1~?�Fнb뢺%*L����D$n�(��16�Ԩd�S�~�ܟ ש(>�L3n�"G�
죄[|:*(:s_�I�.�\;��I��"��8Npg3�g�(�b�I�Z����R:נ��3��L��1�3�\�l#�vg����#y�r�!��-AX�^��׵�C�5Ԩ�fbEџ�Jto����Z��^�DD���;�uo�珂��-"E����뤨���߮�\����0��pa��on�a����r��B.|��5��)w�{ZN����3�
>8�;�i��t����r��nE�@frK3��G�L-+��]�����r�!K����*����V�!�'���g��N	ruv3>8s���ZG�����c]�,��;������L��W��� �����)�6YA�f3�g�Ș����y��/
&�%Ɔ��/^�!;oõ���Hy ��3���p�2/�e�l�da�Wmj8=?Y�04w�!&��MW@c�lt�f�J���m�Y�:Eai
�Mm�`�a�f!g�]�{:��쵡�2&���I7�>B\ǘ`���x�/�e�ND޲`�� �o������)	d�������,�l ���2��(K0�2�zZ������%�'�n��.�
�c�� ��=����f,�?!�0���	h+�a�)��kJ˫��"�%��$�ё�����@n�3k��GEi['I*{O�W��i�oO����󐈁y���h�IQ�oD��y��ɚ�Θ'���~BD�H8�}k�!�U�	T��П�&!�����p�ڊt �&:D�Φ'(���v[���9�D���vQ�$����g�VfSY����[�%8��*g�2K]Ğ���I@כ��� ��N����O$����=��a�Z��o���Q�p�^��q~�����ڔrh�ȃ	/#6����].���V��0T9�2�{6|�k,�x��� �Ӷ�?^Q��=/	m��?�Mg<x�81��ͦTa�  �*x��a��{�����%2,�[\��X��4��iU�S��İ�	�Y$��tAɺ�݈̿x�����������&�z/KR·�~�M��>��{��[�ֵ�m�<��4Y�-����/�X  #�
7`6�d�?�e:0e��m9ܐ�,gζ��w�ÈE�p
�T~-�$�������"��|n�r���T�'��L�p�˺�ׇr���W�f��Sz~>E������*
k2�[���'O@��\)/�:������>���K�\�בj�&���=����̡6_�KE�o|�8_�4���gϱ��Q�Y�Xx0��bA����dn ��m�a��C����n@C�tV�s�߰����!��b��j1`��F-_�'g"��ENm鱉K}��lz���rW�& K�^���(>�0��s}�7G�5Ɩ�p�txf�Ŵb�Wsm�(�aaӬ��`u�[xz���0!�,�1�#��������x���N����},�L�j�� (���K����/@�;x����=05�W�~���Y�P�nlǂ�X���EX�~�U�]��e��{�~��&�/05"���|+y��<Dօ�� q%��G;h���lhϊ��%'ڝ[%ɾ'��:%�A'���L���~(p�a�2���L��ɤ�B�ش�� �Z�I�y\���+1(ʽ�i�N��*K�ԩ~��1��T�f*�K�j`آ�T�!궥m	 �� ��p�
׼�y;�� Bd���9jO^�����I@�����']*�@�X
Yw+�~�e��(�/�i���`�z���11��,�T9�#Y4Cr�˯^HO^�j�d�5h}�A�z/�v>���T3_�_�j@Ss���]G����۞?/7�'�1��@;Jg
s'�|&/B��H��QۯF�)`U�J��8��Aʙ����
14!��z�J���di�Q�Ш������L�0��Oϒ�7����� �
>%������zF5�rϧ9%K���O�˝��FJ�Vk-Y�M��J�6Q�,Ʈ''L(2ʬ��4;�XaB8���p��ހ���j�(�j{�+Q:�?Fj> fJ��=�~a)��_� ��'Β�5��D��b,c�y�wRs��4v/��W|A+��0E�T��Ϙ��V��$��{�&2�^4�1�D��1ډ�w}�f|hա�u'���{S��G9a���#��$\F��@��;�Y��I����+^!$WʼAsy���Ú��(����cW�7��`^�ZB��d,TOȰ���K��Aڏ���ԭ������� uR���sh��ަ��_o�j=5C��+ޒu4{�Į����T醥��.�K��j	"mػ��:�iz��n�< -����[�9"�(i���$m�6ч����.���[��,`��~X}:ќx�ȩ.��]$H�	G߫��2a7�fz�m�
�%˅�y�hR�ny�7����)�0�qLP�+ǐ�J&���&i��Y����� f�1:tP�lv���vvY�1�bٳzN�[[>��� =C8urs>��t˴�1ڿAKBO[^ƻ����R2A�&�oI��n/�KC����8�+�w<![��?P��9׬j�c�93�7#���X*�"���E[��� �����(��X,s/��)&�	��>� �䌬a����q����0�u� ��',��?��	X�=0*����Ǩq[�5�T��A貂�����ηS�����h��dy�	gy{%�'Lݯ�J\�ḝj z)I�'���B���,��"�v�0�?�/�<\�25Ԉa��p��P�����{��2�&.O�5-8zd�B��P���e�(���s�Ϯ�7��1ד�}���
��e��m@� #A;%����3�HE�^��C�;$���1-��8�}�T�'SQ/��& �Bwq��bJ��\�F-�.E&��XCs(ėk�A%4Ϡ�Ac�_���Od�:)�W�i��-�X��=�y��h�|>���iH���n�?L%���Z�Κaga�RW F%���yM�C��Ļ��5w���L�b�ں��Ӭ���ˬ�"�k��:r�����MW=���d�K���Dax��V�� ���n���nG(���,�&�C.��(XgG�[�B�c��D�Hy�ˑ��$��q�)�Y&"q.�RD�l��oiR�K���_��2����
ƚGJe�=k0��'����萡��+��_�fPX�T�1r